* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 CSoutput.t235 commonsourceibias.t80 gnd.t384 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 a_n1986_8322.t17 a_n1986_13878.t40 vdd.t166 vdd.t165 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X2 a_n1808_13878.t11 a_n1986_13878.t19 a_n1986_13878.t20 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X3 gnd.t383 commonsourceibias.t81 CSoutput.t234 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 vdd.t9 a_n7636_8799.t28 CSoutput.t4 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 CSoutput.t233 commonsourceibias.t82 gnd.t382 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 CSoutput.t232 commonsourceibias.t83 gnd.t381 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 gnd.t373 commonsourceibias.t84 CSoutput.t231 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 a_n1986_13878.t24 a_n1986_13878.t23 a_n1808_13878.t10 vdd.t144 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X9 vdd.t244 vdd.t242 vdd.t243 vdd.t220 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X10 CSoutput.t240 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X11 CSoutput.t5 a_n7636_8799.t29 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 a_n1808_13878.t9 a_n1986_13878.t21 a_n1986_13878.t22 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 a_n1808_13878.t19 a_n1986_13878.t41 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 vdd.t249 a_n7636_8799.t30 CSoutput.t76 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 CSoutput.t77 a_n7636_8799.t31 vdd.t250 vdd.t94 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 CSoutput.t230 commonsourceibias.t85 gnd.t380 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t44 a_n7636_8799.t32 vdd.t89 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 gnd.t379 commonsourceibias.t86 CSoutput.t229 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t228 commonsourceibias.t87 gnd.t378 gnd.t280 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 a_n7636_8799.t22 plus.t5 a_n2903_n3924.t28 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X21 gnd.t374 commonsourceibias.t88 CSoutput.t227 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X22 CSoutput.t226 commonsourceibias.t89 gnd.t377 gnd.t280 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t225 commonsourceibias.t90 gnd.t376 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 gnd.t375 commonsourceibias.t91 CSoutput.t224 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 gnd.t129 gnd.t126 gnd.t128 gnd.t127 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X26 gnd.t125 gnd.t123 gnd.t124 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X27 commonsourceibias.t79 commonsourceibias.t78 gnd.t372 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 vdd.t241 vdd.t239 vdd.t240 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X29 vdd.t21 CSoutput.t241 output.t15 gnd.t183 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X30 CSoutput.t223 commonsourceibias.t92 gnd.t371 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 a_n1986_8322.t1 a_n1986_13878.t42 a_n7636_8799.t18 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X32 gnd.t122 gnd.t120 gnd.t121 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X33 CSoutput.t45 a_n7636_8799.t33 vdd.t91 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 vdd.t33 a_n7636_8799.t34 CSoutput.t8 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 CSoutput.t222 commonsourceibias.t93 gnd.t370 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t369 commonsourceibias.t94 CSoutput.t221 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd.t119 gnd.t117 gnd.t118 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X38 a_n7636_8799.t5 plus.t6 a_n2903_n3924.t27 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X39 CSoutput.t220 commonsourceibias.t95 gnd.t368 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t219 commonsourceibias.t96 gnd.t367 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 vdd.t35 a_n7636_8799.t35 CSoutput.t9 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 CSoutput.t218 commonsourceibias.t97 gnd.t366 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 vdd.t290 a_n7636_8799.t36 CSoutput.t114 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 CSoutput.t115 a_n7636_8799.t37 vdd.t291 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 a_n7636_8799.t17 a_n1986_13878.t43 a_n1986_8322.t3 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X46 vdd.t55 a_n7636_8799.t38 CSoutput.t22 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 a_n2903_n3924.t8 diffpairibias.t16 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X48 gnd.t365 commonsourceibias.t98 CSoutput.t217 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X49 a_n2903_n3924.t33 minus.t5 a_n1986_13878.t37 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X50 CSoutput.t23 a_n7636_8799.t39 vdd.t56 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X51 gnd.t364 commonsourceibias.t99 CSoutput.t216 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 gnd.t116 gnd.t114 plus.t4 gnd.t115 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X53 a_n2903_n3924.t26 plus.t7 a_n7636_8799.t21 gnd.t144 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X54 CSoutput.t215 commonsourceibias.t100 gnd.t344 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t214 commonsourceibias.t101 gnd.t363 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X56 a_n1986_13878.t36 minus.t6 a_n2903_n3924.t32 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X57 gnd.t362 commonsourceibias.t2 commonsourceibias.t3 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 CSoutput.t213 commonsourceibias.t102 gnd.t361 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 a_n2903_n3924.t0 minus.t7 a_n1986_13878.t0 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X60 gnd.t360 commonsourceibias.t103 CSoutput.t212 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X61 vdd.t238 vdd.t236 vdd.t237 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X62 CSoutput.t84 a_n7636_8799.t40 vdd.t258 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 CSoutput.t85 a_n7636_8799.t41 vdd.t259 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 CSoutput.t211 commonsourceibias.t104 gnd.t359 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X65 CSoutput.t210 commonsourceibias.t105 gnd.t358 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 gnd.t357 commonsourceibias.t106 CSoutput.t209 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 CSoutput.t208 commonsourceibias.t107 gnd.t353 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 gnd.t356 commonsourceibias.t108 CSoutput.t207 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 vdd.t16 CSoutput.t242 output.t14 gnd.t184 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X70 CSoutput.t243 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X71 output.t13 CSoutput.t244 vdd.t26 gnd.t179 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X72 CSoutput.t82 a_n7636_8799.t42 vdd.t256 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X73 gnd.t355 commonsourceibias.t0 commonsourceibias.t1 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 a_n2903_n3924.t31 minus.t8 a_n1986_13878.t35 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X75 CSoutput.t206 commonsourceibias.t109 gnd.t354 gnd.t280 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 gnd.t113 gnd.t111 gnd.t112 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X77 CSoutput.t205 commonsourceibias.t110 gnd.t352 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X78 diffpairibias.t15 diffpairibias.t14 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 a_n1808_13878.t8 a_n1986_13878.t31 a_n1986_13878.t32 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X80 vdd.t235 vdd.t233 vdd.t234 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X81 gnd.t351 commonsourceibias.t111 CSoutput.t204 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 vdd.t257 a_n7636_8799.t43 CSoutput.t83 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t110 a_n7636_8799.t44 vdd.t286 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 a_n1986_13878.t26 a_n1986_13878.t25 a_n1808_13878.t7 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X85 CSoutput.t203 commonsourceibias.t112 gnd.t350 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X86 gnd.t110 gnd.t107 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X87 CSoutput.t202 commonsourceibias.t113 gnd.t349 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 gnd.t348 commonsourceibias.t114 CSoutput.t201 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t347 commonsourceibias.t115 CSoutput.t200 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t111 a_n7636_8799.t45 vdd.t287 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 vdd.t232 vdd.t230 vdd.t231 vdd.t205 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X92 gnd.t346 commonsourceibias.t116 CSoutput.t199 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 gnd.t106 gnd.t104 plus.t3 gnd.t105 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X94 vdd.t51 a_n7636_8799.t46 CSoutput.t20 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 minus.t4 gnd.t101 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X96 CSoutput.t198 commonsourceibias.t117 gnd.t345 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 diffpairibias.t13 diffpairibias.t12 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X98 gnd.t343 commonsourceibias.t8 commonsourceibias.t9 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t342 commonsourceibias.t118 CSoutput.t197 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 CSoutput.t196 commonsourceibias.t119 gnd.t341 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 gnd.t299 commonsourceibias.t120 CSoutput.t195 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X102 CSoutput.t194 commonsourceibias.t121 gnd.t340 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X103 CSoutput.t193 commonsourceibias.t122 gnd.t339 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 CSoutput.t21 a_n7636_8799.t47 vdd.t53 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 vdd.t292 a_n7636_8799.t48 CSoutput.t236 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X106 vdd.t293 a_n7636_8799.t49 CSoutput.t237 vdd.t265 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 CSoutput.t192 commonsourceibias.t123 gnd.t338 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t337 commonsourceibias.t124 CSoutput.t191 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 vdd.t294 a_n7636_8799.t50 CSoutput.t238 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 vdd.t295 a_n7636_8799.t51 CSoutput.t239 vdd.t271 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 CSoutput.t74 a_n7636_8799.t52 vdd.t247 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X112 CSoutput.t75 a_n7636_8799.t53 vdd.t248 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 gnd.t336 commonsourceibias.t6 commonsourceibias.t7 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 gnd.t335 commonsourceibias.t4 commonsourceibias.t5 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X115 CSoutput.t190 commonsourceibias.t125 gnd.t334 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 a_n7636_8799.t19 plus.t8 a_n2903_n3924.t25 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X117 CSoutput.t189 commonsourceibias.t126 gnd.t333 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 vdd.t116 a_n7636_8799.t54 CSoutput.t64 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X119 gnd.t332 commonsourceibias.t127 CSoutput.t188 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 CSoutput.t65 a_n7636_8799.t55 vdd.t117 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 output.t12 CSoutput.t245 vdd.t24 gnd.t180 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X122 a_n2903_n3924.t5 diffpairibias.t17 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X123 CSoutput.t62 a_n7636_8799.t56 vdd.t114 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 CSoutput.t63 a_n7636_8799.t57 vdd.t115 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X125 CSoutput.t246 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X126 vdd.t23 CSoutput.t247 output.t11 gnd.t175 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X127 CSoutput.t42 a_n7636_8799.t58 vdd.t86 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 gnd.t100 gnd.t98 gnd.t99 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X129 a_n2903_n3924.t4 minus.t9 a_n1986_13878.t4 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X130 gnd.t331 commonsourceibias.t128 CSoutput.t187 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 vdd.t87 a_n7636_8799.t59 CSoutput.t43 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X132 a_n1986_13878.t38 minus.t10 a_n2903_n3924.t34 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X133 gnd.t97 gnd.t95 gnd.t96 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X134 a_n2903_n3924.t24 plus.t9 a_n7636_8799.t6 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X135 gnd.t330 commonsourceibias.t129 CSoutput.t186 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 CSoutput.t185 commonsourceibias.t130 gnd.t329 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 vdd.t18 CSoutput.t248 output.t10 gnd.t176 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X138 vdd.t167 a_n7636_8799.t60 CSoutput.t70 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X139 commonsourceibias.t15 commonsourceibias.t14 gnd.t328 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 a_n1986_13878.t34 a_n1986_13878.t33 a_n1808_13878.t6 vdd.t161 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 vdd.t168 a_n7636_8799.t61 CSoutput.t71 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 vdd.t245 a_n7636_8799.t62 CSoutput.t72 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X143 a_n7636_8799.t16 a_n1986_13878.t44 a_n1986_8322.t2 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 a_n1986_13878.t28 a_n1986_13878.t27 a_n1808_13878.t5 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X145 gnd.t327 commonsourceibias.t131 CSoutput.t184 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 vdd.t246 a_n7636_8799.t63 CSoutput.t73 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X147 a_n2903_n3924.t29 minus.t11 a_n1986_13878.t9 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X148 gnd.t321 commonsourceibias.t132 CSoutput.t183 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 gnd.t326 commonsourceibias.t12 commonsourceibias.t13 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 gnd.t324 commonsourceibias.t133 CSoutput.t182 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 vdd.t280 a_n7636_8799.t64 CSoutput.t104 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 CSoutput.t105 a_n7636_8799.t65 vdd.t281 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X153 output.t9 CSoutput.t249 vdd.t27 gnd.t177 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X154 gnd.t94 gnd.t92 gnd.t93 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X155 CSoutput.t181 commonsourceibias.t134 gnd.t325 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X156 vdd.t229 vdd.t227 vdd.t228 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X157 vdd.t278 a_n7636_8799.t66 CSoutput.t102 vdd.t271 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X158 gnd.t323 commonsourceibias.t135 CSoutput.t180 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 a_n2903_n3924.t39 diffpairibias.t18 gnd.t398 gnd.t397 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X160 CSoutput.t103 a_n7636_8799.t67 vdd.t279 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 gnd.t322 commonsourceibias.t136 CSoutput.t179 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 a_n1986_13878.t1 minus.t12 a_n2903_n3924.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X163 vdd.t226 vdd.t223 vdd.t225 vdd.t224 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X164 gnd.t320 commonsourceibias.t10 commonsourceibias.t11 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 CSoutput.t178 commonsourceibias.t137 gnd.t319 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 gnd.t318 commonsourceibias.t138 CSoutput.t177 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 CSoutput.t176 commonsourceibias.t139 gnd.t317 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 CSoutput.t175 commonsourceibias.t140 gnd.t316 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X169 CSoutput.t174 commonsourceibias.t141 gnd.t315 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 vdd.t222 vdd.t219 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X171 output.t8 CSoutput.t250 vdd.t19 gnd.t178 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X172 a_n2903_n3924.t23 plus.t10 a_n7636_8799.t4 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X173 vdd.t218 vdd.t216 vdd.t217 vdd.t209 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X174 vdd.t160 a_n1986_13878.t45 a_n1986_8322.t16 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 a_n1986_8322.t15 a_n1986_13878.t46 vdd.t158 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 CSoutput.t60 a_n7636_8799.t68 vdd.t112 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X177 CSoutput.t61 a_n7636_8799.t69 vdd.t113 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 gnd.t91 gnd.t89 gnd.t90 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X179 vdd.t83 a_n7636_8799.t70 CSoutput.t40 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 vdd.t156 a_n1986_13878.t47 a_n1808_13878.t18 vdd.t155 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X181 a_n7636_8799.t23 plus.t11 a_n2903_n3924.t22 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X182 vdd.t215 vdd.t212 vdd.t214 vdd.t213 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X183 diffpairibias.t11 diffpairibias.t10 gnd.t388 gnd.t387 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X184 vdd.t211 vdd.t208 vdd.t210 vdd.t209 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X185 vdd.t84 a_n7636_8799.t71 CSoutput.t41 vdd.t34 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X186 CSoutput.t173 commonsourceibias.t142 gnd.t314 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 commonsourceibias.t21 commonsourceibias.t20 gnd.t313 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 gnd.t312 commonsourceibias.t143 CSoutput.t172 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 gnd.t311 commonsourceibias.t18 commonsourceibias.t19 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 vdd.t207 vdd.t204 vdd.t206 vdd.t205 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X191 a_n7636_8799.t15 a_n1986_13878.t48 a_n1986_8322.t5 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X192 a_n1986_8322.t14 a_n1986_13878.t49 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X193 CSoutput.t171 commonsourceibias.t144 gnd.t310 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 CSoutput.t38 a_n7636_8799.t72 vdd.t79 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X195 plus.t2 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X196 vdd.t81 a_n7636_8799.t73 CSoutput.t39 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 vdd.t5 a_n7636_8799.t74 CSoutput.t2 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X198 gnd.t85 gnd.t82 gnd.t84 gnd.t83 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X199 a_n1986_13878.t30 a_n1986_13878.t29 a_n1808_13878.t4 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X200 gnd.t81 gnd.t79 minus.t3 gnd.t80 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X201 a_n7636_8799.t14 a_n1986_13878.t50 a_n1986_8322.t4 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X202 CSoutput.t3 a_n7636_8799.t75 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 a_n1986_13878.t7 minus.t13 a_n2903_n3924.t9 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X204 CSoutput.t170 commonsourceibias.t145 gnd.t309 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 a_n1808_13878.t3 a_n1986_13878.t15 a_n1986_13878.t16 vdd.t151 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X206 gnd.t308 commonsourceibias.t146 CSoutput.t169 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 gnd.t307 commonsourceibias.t147 CSoutput.t168 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 gnd.t306 commonsourceibias.t148 CSoutput.t167 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 gnd.t305 commonsourceibias.t149 CSoutput.t166 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X210 vdd.t20 CSoutput.t251 output.t7 gnd.t162 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X211 commonsourceibias.t17 commonsourceibias.t16 gnd.t304 gnd.t303 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 gnd.t302 commonsourceibias.t150 CSoutput.t165 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 gnd.t78 gnd.t76 gnd.t77 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 gnd.t300 commonsourceibias.t151 CSoutput.t164 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X215 CSoutput.t66 a_n7636_8799.t76 vdd.t118 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 vdd.t150 a_n1986_13878.t51 a_n1986_8322.t13 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X217 vdd.t120 a_n7636_8799.t77 CSoutput.t67 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 CSoutput.t163 commonsourceibias.t152 gnd.t298 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 a_n2903_n3924.t12 diffpairibias.t19 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X220 gnd.t21 gnd.t18 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X221 a_n2903_n3924.t11 diffpairibias.t20 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X222 commonsourceibias.t35 commonsourceibias.t34 gnd.t297 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X223 a_n1986_13878.t5 minus.t14 a_n2903_n3924.t6 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X224 CSoutput.t68 a_n7636_8799.t78 vdd.t121 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 vdd.t122 a_n7636_8799.t79 CSoutput.t69 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X226 gnd.t75 gnd.t73 gnd.t74 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X227 vdd.t29 a_n7636_8799.t80 CSoutput.t6 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 CSoutput.t162 commonsourceibias.t153 gnd.t295 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X229 CSoutput.t161 commonsourceibias.t154 gnd.t294 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 commonsourceibias.t33 commonsourceibias.t32 gnd.t293 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 vdd.t31 a_n7636_8799.t81 CSoutput.t7 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 output.t16 outputibias.t8 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X233 vdd.t288 a_n7636_8799.t82 CSoutput.t112 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 CSoutput.t160 commonsourceibias.t155 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 commonsourceibias.t31 commonsourceibias.t30 gnd.t290 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 a_n1986_13878.t10 minus.t15 a_n2903_n3924.t30 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X237 CSoutput.t159 commonsourceibias.t156 gnd.t289 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X238 outputibias.t7 outputibias.t6 gnd.t394 gnd.t393 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X239 gnd.t288 commonsourceibias.t28 commonsourceibias.t29 gnd.t287 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 diffpairibias.t9 diffpairibias.t8 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X241 output.t17 outputibias.t9 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X242 CSoutput.t158 commonsourceibias.t157 gnd.t286 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 output.t6 CSoutput.t252 vdd.t13 gnd.t163 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X244 CSoutput.t157 commonsourceibias.t158 gnd.t285 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X245 CSoutput.t113 a_n7636_8799.t83 vdd.t289 vdd.t252 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 CSoutput.t156 commonsourceibias.t159 gnd.t284 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X247 a_n2903_n3924.t21 plus.t12 a_n7636_8799.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X248 gnd.t283 commonsourceibias.t26 commonsourceibias.t27 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t58 a_n7636_8799.t84 vdd.t109 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 CSoutput.t59 a_n7636_8799.t85 vdd.t110 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 outputibias.t5 outputibias.t4 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X252 commonsourceibias.t25 commonsourceibias.t24 gnd.t281 gnd.t280 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 gnd.t279 commonsourceibias.t160 CSoutput.t155 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t69 gnd.t67 gnd.t68 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X255 plus.t1 gnd.t70 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X256 a_n1808_13878.t17 a_n1986_13878.t52 vdd.t148 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X257 a_n2903_n3924.t20 plus.t13 a_n7636_8799.t3 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X258 vdd.t203 vdd.t201 vdd.t202 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X259 gnd.t278 commonsourceibias.t22 commonsourceibias.t23 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 gnd.t66 gnd.t64 gnd.t65 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X261 gnd.t63 gnd.t61 minus.t2 gnd.t62 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X262 vdd.t146 a_n1986_13878.t53 a_n1808_13878.t16 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X263 gnd.t259 commonsourceibias.t161 CSoutput.t154 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 vdd.t200 vdd.t198 vdd.t199 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X265 commonsourceibias.t49 commonsourceibias.t48 gnd.t277 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X266 CSoutput.t100 a_n7636_8799.t86 vdd.t276 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 vdd.t277 a_n7636_8799.t87 CSoutput.t101 vdd.t119 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 gnd.t276 commonsourceibias.t46 commonsourceibias.t47 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 vdd.t197 vdd.t195 vdd.t196 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X270 CSoutput.t153 commonsourceibias.t162 gnd.t275 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 diffpairibias.t7 diffpairibias.t6 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X272 commonsourceibias.t45 commonsourceibias.t44 gnd.t274 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 gnd.t60 gnd.t58 gnd.t59 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X274 CSoutput.t56 a_n7636_8799.t88 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 vdd.t108 a_n7636_8799.t89 CSoutput.t57 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X276 vdd.t75 a_n7636_8799.t90 CSoutput.t36 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 gnd.t273 commonsourceibias.t163 CSoutput.t152 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t14 CSoutput.t253 output.t5 gnd.t164 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X279 CSoutput.t37 a_n7636_8799.t91 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 a_n1986_8322.t9 a_n1986_13878.t54 a_n7636_8799.t13 vdd.t144 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X281 gnd.t272 commonsourceibias.t42 commonsourceibias.t43 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 CSoutput.t151 commonsourceibias.t164 gnd.t270 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 vdd.t274 a_n7636_8799.t92 CSoutput.t98 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X284 CSoutput.t99 a_n7636_8799.t93 vdd.t275 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 vdd.t272 a_n7636_8799.t94 CSoutput.t96 vdd.t271 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 vdd.t143 a_n1986_13878.t55 a_n1986_8322.t12 vdd.t142 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X287 vdd.t273 a_n7636_8799.t95 CSoutput.t97 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 vdd.t103 a_n7636_8799.t96 CSoutput.t54 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 gnd.t269 commonsourceibias.t165 CSoutput.t150 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 gnd.t57 gnd.t55 minus.t1 gnd.t56 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X291 gnd.t54 gnd.t51 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X292 output.t4 CSoutput.t254 vdd.t12 gnd.t165 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X293 a_n1808_13878.t15 a_n1986_13878.t56 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X294 a_n2903_n3924.t35 diffpairibias.t21 gnd.t390 gnd.t389 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X295 CSoutput.t255 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X296 gnd.t268 commonsourceibias.t40 commonsourceibias.t41 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 vdd.t104 a_n7636_8799.t97 CSoutput.t55 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 outputibias.t3 outputibias.t2 gnd.t167 gnd.t166 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X299 CSoutput.t34 a_n7636_8799.t98 vdd.t72 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 CSoutput.t35 a_n7636_8799.t99 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 vdd.t194 vdd.t191 vdd.t193 vdd.t192 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X302 output.t18 outputibias.t10 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X303 vdd.t190 vdd.t188 vdd.t189 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X304 a_n1986_8322.t8 a_n1986_13878.t57 a_n7636_8799.t12 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X305 vdd.t187 vdd.t184 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X306 vdd.t138 a_n1986_13878.t58 a_n1986_8322.t11 vdd.t137 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X307 CSoutput.t32 a_n7636_8799.t100 vdd.t70 vdd.t69 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 vdd.t71 a_n7636_8799.t101 CSoutput.t33 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 gnd.t267 commonsourceibias.t38 commonsourceibias.t39 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 a_n2903_n3924.t19 plus.t14 a_n7636_8799.t20 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X311 CSoutput.t0 a_n7636_8799.t102 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 CSoutput.t149 commonsourceibias.t166 gnd.t266 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 vdd.t3 a_n7636_8799.t103 CSoutput.t1 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X314 gnd.t50 gnd.t48 gnd.t49 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X315 a_n7636_8799.t27 plus.t15 a_n2903_n3924.t18 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X316 vdd.t100 a_n7636_8799.t104 CSoutput.t52 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 CSoutput.t148 commonsourceibias.t167 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X318 a_n2903_n3924.t2 minus.t16 a_n1986_13878.t2 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X319 diffpairibias.t5 diffpairibias.t4 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X320 CSoutput.t256 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X321 output.t3 CSoutput.t257 vdd.t22 gnd.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X322 a_n2903_n3924.t10 minus.t17 a_n1986_13878.t8 gnd.t144 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X323 a_n7636_8799.t2 plus.t16 a_n2903_n3924.t17 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X324 vdd.t183 vdd.t180 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X325 gnd.t47 gnd.t44 gnd.t46 gnd.t45 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X326 vdd.t101 a_n7636_8799.t105 CSoutput.t53 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X327 CSoutput.t94 a_n7636_8799.t106 vdd.t269 vdd.t111 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X328 CSoutput.t95 a_n7636_8799.t107 vdd.t270 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 gnd.t263 commonsourceibias.t36 commonsourceibias.t37 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 a_n1808_13878.t2 a_n1986_13878.t13 a_n1986_13878.t14 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 CSoutput.t147 commonsourceibias.t168 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 output.t2 CSoutput.t258 vdd.t17 gnd.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X333 a_n1986_8322.t20 a_n1986_13878.t59 a_n7636_8799.t11 vdd.t136 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X334 commonsourceibias.t63 commonsourceibias.t62 gnd.t258 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X335 a_n2903_n3924.t16 plus.t17 a_n7636_8799.t26 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X336 CSoutput.t50 a_n7636_8799.t108 vdd.t98 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t51 a_n7636_8799.t109 vdd.t99 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 gnd.t188 commonsourceibias.t169 CSoutput.t146 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 vdd.t66 a_n7636_8799.t110 CSoutput.t30 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 vdd.t68 a_n7636_8799.t111 CSoutput.t31 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X341 a_n1986_8322.t10 a_n1986_13878.t60 vdd.t135 vdd.t134 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X342 CSoutput.t92 a_n7636_8799.t112 vdd.t267 vdd.t73 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t257 commonsourceibias.t170 CSoutput.t145 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 a_n2903_n3924.t3 minus.t18 a_n1986_13878.t3 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X345 gnd.t256 commonsourceibias.t171 CSoutput.t144 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 vdd.t133 a_n1986_13878.t61 a_n1808_13878.t14 vdd.t132 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X347 commonsourceibias.t61 commonsourceibias.t60 gnd.t255 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 CSoutput.t93 a_n7636_8799.t113 vdd.t268 vdd.t90 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X349 CSoutput.t12 a_n7636_8799.t114 vdd.t39 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 vdd.t15 CSoutput.t259 output.t1 gnd.t181 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X351 gnd.t253 commonsourceibias.t172 CSoutput.t143 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 vdd.t40 a_n7636_8799.t115 CSoutput.t13 vdd.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 vdd.t63 a_n7636_8799.t116 CSoutput.t28 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 vdd.t179 vdd.t176 vdd.t178 vdd.t177 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X355 commonsourceibias.t59 commonsourceibias.t58 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 a_n1986_8322.t19 a_n1986_13878.t62 a_n7636_8799.t10 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X357 vdd.t175 vdd.t173 vdd.t174 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X358 gnd.t43 gnd.t40 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X359 CSoutput.t29 a_n7636_8799.t117 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X360 a_n7636_8799.t9 a_n1986_13878.t63 a_n1986_8322.t7 vdd.t131 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X361 gnd.t244 commonsourceibias.t173 CSoutput.t142 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 vdd.t264 a_n7636_8799.t118 CSoutput.t90 vdd.t102 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 commonsourceibias.t57 commonsourceibias.t56 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X364 a_n1808_13878.t13 a_n1986_13878.t64 vdd.t130 vdd.t129 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X365 gnd.t248 commonsourceibias.t174 CSoutput.t141 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 a_n1986_13878.t6 minus.t19 a_n2903_n3924.t7 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X367 CSoutput.t140 commonsourceibias.t175 gnd.t242 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 vdd.t266 a_n7636_8799.t119 CSoutput.t91 vdd.t265 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 gnd.t246 commonsourceibias.t54 commonsourceibias.t55 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 CSoutput.t88 a_n7636_8799.t120 vdd.t262 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 outputibias.t1 outputibias.t0 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X372 gnd.t245 commonsourceibias.t52 commonsourceibias.t53 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X373 commonsourceibias.t51 commonsourceibias.t50 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 gnd.t39 gnd.t36 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X375 gnd.t239 commonsourceibias.t176 CSoutput.t139 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 gnd.t238 commonsourceibias.t177 CSoutput.t138 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X377 vdd.t263 a_n7636_8799.t121 CSoutput.t89 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 CSoutput.t48 a_n7636_8799.t122 vdd.t96 vdd.t78 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 a_n7636_8799.t24 plus.t18 a_n2903_n3924.t15 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X380 CSoutput.t49 a_n7636_8799.t123 vdd.t97 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X381 CSoutput.t26 a_n7636_8799.t124 vdd.t61 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 CSoutput.t27 a_n7636_8799.t125 vdd.t62 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 a_n1808_13878.t1 a_n1986_13878.t17 a_n1986_13878.t18 vdd.t128 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X384 a_n2903_n3924.t36 diffpairibias.t22 gnd.t392 gnd.t391 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 gnd.t237 commonsourceibias.t178 CSoutput.t137 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X386 CSoutput.t136 commonsourceibias.t179 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 vdd.t93 a_n7636_8799.t126 CSoutput.t46 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 gnd.t227 commonsourceibias.t180 CSoutput.t135 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 CSoutput.t134 commonsourceibias.t181 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 gnd.t35 gnd.t32 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X391 a_n2903_n3924.t14 plus.t19 a_n7636_8799.t25 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X392 CSoutput.t47 a_n7636_8799.t127 vdd.t95 vdd.t94 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X393 CSoutput.t133 commonsourceibias.t182 gnd.t233 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 gnd.t232 commonsourceibias.t183 CSoutput.t132 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X395 commonsourceibias.t75 commonsourceibias.t74 gnd.t230 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X396 vdd.t57 a_n7636_8799.t128 CSoutput.t24 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 vdd.t59 a_n7636_8799.t129 CSoutput.t25 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X398 CSoutput.t131 commonsourceibias.t184 gnd.t226 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X399 gnd.t17 gnd.t14 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X400 diffpairibias.t3 diffpairibias.t2 gnd.t5 gnd.t4 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X401 CSoutput.t86 a_n7636_8799.t130 vdd.t260 vdd.t252 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X402 a_n1986_13878.t12 a_n1986_13878.t11 a_n1808_13878.t0 vdd.t127 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X403 CSoutput.t130 commonsourceibias.t185 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 gnd.t222 commonsourceibias.t186 CSoutput.t129 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 vdd.t261 a_n7636_8799.t131 CSoutput.t87 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X406 a_n7636_8799.t8 a_n1986_13878.t65 a_n1986_8322.t6 vdd.t126 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X407 CSoutput.t10 a_n7636_8799.t132 vdd.t37 vdd.t36 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X408 vdd.t38 a_n7636_8799.t133 CSoutput.t11 vdd.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X409 diffpairibias.t1 diffpairibias.t0 gnd.t156 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X410 gnd.t221 commonsourceibias.t187 CSoutput.t128 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 a_n7636_8799.t1 plus.t20 a_n2903_n3924.t13 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X412 CSoutput.t260 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X413 vdd.t49 a_n7636_8799.t134 CSoutput.t18 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 vdd.t172 vdd.t169 vdd.t171 vdd.t170 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X415 commonsourceibias.t73 commonsourceibias.t72 gnd.t219 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X416 gnd.t208 commonsourceibias.t188 CSoutput.t127 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X417 CSoutput.t19 a_n7636_8799.t135 vdd.t50 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X418 commonsourceibias.t71 commonsourceibias.t70 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X419 CSoutput.t126 commonsourceibias.t189 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X420 vdd.t284 a_n7636_8799.t136 CSoutput.t108 vdd.t265 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X421 gnd.t214 commonsourceibias.t68 commonsourceibias.t69 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X422 gnd.t212 commonsourceibias.t66 commonsourceibias.t67 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 gnd.t210 commonsourceibias.t190 CSoutput.t125 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 a_n1986_13878.t39 minus.t20 a_n2903_n3924.t37 gnd.t173 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X425 vdd.t125 a_n1986_13878.t66 a_n1808_13878.t12 vdd.t124 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X426 commonsourceibias.t65 commonsourceibias.t64 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 gnd.t205 commonsourceibias.t191 CSoutput.t124 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X428 gnd.t203 commonsourceibias.t192 CSoutput.t123 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X429 CSoutput.t109 a_n7636_8799.t137 vdd.t285 vdd.t60 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X430 gnd.t192 commonsourceibias.t193 CSoutput.t122 gnd.t191 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X431 CSoutput.t16 a_n7636_8799.t138 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X432 vdd.t25 CSoutput.t261 output.t0 gnd.t182 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X433 vdd.t48 a_n7636_8799.t139 CSoutput.t17 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X434 vdd.t254 a_n7636_8799.t140 CSoutput.t80 vdd.t92 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X435 output.t19 outputibias.t11 gnd.t386 gnd.t385 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X436 CSoutput.t81 a_n7636_8799.t141 vdd.t255 vdd.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X437 gnd.t31 gnd.t29 gnd.t30 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X438 gnd.t201 commonsourceibias.t194 CSoutput.t121 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X439 gnd.t28 gnd.t25 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X440 gnd.t24 gnd.t22 plus.t0 gnd.t23 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X441 gnd.t200 commonsourceibias.t195 CSoutput.t120 gnd.t199 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X442 CSoutput.t106 a_n7636_8799.t142 vdd.t282 vdd.t94 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X443 gnd.t190 commonsourceibias.t196 CSoutput.t119 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X444 CSoutput.t118 commonsourceibias.t197 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X445 commonsourceibias.t77 commonsourceibias.t76 gnd.t196 gnd.t195 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X446 CSoutput.t117 commonsourceibias.t198 gnd.t194 gnd.t193 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X447 a_n1986_8322.t18 a_n1986_13878.t67 a_n7636_8799.t7 vdd.t123 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X448 minus.t0 gnd.t11 gnd.t13 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X449 vdd.t283 a_n7636_8799.t143 CSoutput.t107 vdd.t58 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X450 vdd.t42 a_n7636_8799.t144 CSoutput.t14 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X451 a_n2903_n3924.t38 diffpairibias.t23 gnd.t396 gnd.t395 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X452 CSoutput.t15 a_n7636_8799.t145 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X453 vdd.t251 a_n7636_8799.t146 CSoutput.t78 vdd.t107 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X454 CSoutput.t79 a_n7636_8799.t147 vdd.t253 vdd.t252 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X455 gnd.t186 commonsourceibias.t199 CSoutput.t116 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
R0 commonsourceibias.n397 commonsourceibias.t184 222.032
R1 commonsourceibias.n281 commonsourceibias.t134 222.032
R2 commonsourceibias.n44 commonsourceibias.t62 222.032
R3 commonsourceibias.n166 commonsourceibias.t140 222.032
R4 commonsourceibias.n875 commonsourceibias.t191 222.032
R5 commonsourceibias.n759 commonsourceibias.t98 222.032
R6 commonsourceibias.n529 commonsourceibias.t4 222.032
R7 commonsourceibias.n645 commonsourceibias.t177 222.032
R8 commonsourceibias.n480 commonsourceibias.t183 207.983
R9 commonsourceibias.n364 commonsourceibias.t88 207.983
R10 commonsourceibias.n127 commonsourceibias.t52 207.983
R11 commonsourceibias.n249 commonsourceibias.t151 207.983
R12 commonsourceibias.n963 commonsourceibias.t101 207.983
R13 commonsourceibias.n847 commonsourceibias.t189 207.983
R14 commonsourceibias.n617 commonsourceibias.t48 207.983
R15 commonsourceibias.n732 commonsourceibias.t112 207.983
R16 commonsourceibias.n396 commonsourceibias.t150 168.701
R17 commonsourceibias.n402 commonsourceibias.t155 168.701
R18 commonsourceibias.n408 commonsourceibias.t199 168.701
R19 commonsourceibias.n392 commonsourceibias.t175 168.701
R20 commonsourceibias.n416 commonsourceibias.t165 168.701
R21 commonsourceibias.n422 commonsourceibias.t96 168.701
R22 commonsourceibias.n387 commonsourceibias.t187 168.701
R23 commonsourceibias.n430 commonsourceibias.t168 168.701
R24 commonsourceibias.n436 commonsourceibias.t172 168.701
R25 commonsourceibias.n382 commonsourceibias.t80 168.701
R26 commonsourceibias.n444 commonsourceibias.t173 168.701
R27 commonsourceibias.n450 commonsourceibias.t182 168.701
R28 commonsourceibias.n377 commonsourceibias.t149 168.701
R29 commonsourceibias.n458 commonsourceibias.t110 168.701
R30 commonsourceibias.n464 commonsourceibias.t194 168.701
R31 commonsourceibias.n372 commonsourceibias.t157 168.701
R32 commonsourceibias.n472 commonsourceibias.t163 168.701
R33 commonsourceibias.n478 commonsourceibias.t92 168.701
R34 commonsourceibias.n362 commonsourceibias.t198 168.701
R35 commonsourceibias.n356 commonsourceibias.t186 168.701
R36 commonsourceibias.n256 commonsourceibias.t95 168.701
R37 commonsourceibias.n348 commonsourceibias.t196 168.701
R38 commonsourceibias.n342 commonsourceibias.t105 168.701
R39 commonsourceibias.n261 commonsourceibias.t94 168.701
R40 commonsourceibias.n334 commonsourceibias.t197 168.701
R41 commonsourceibias.n328 commonsourceibias.t115 168.701
R42 commonsourceibias.n266 commonsourceibias.t141 168.701
R43 commonsourceibias.n320 commonsourceibias.t195 168.701
R44 commonsourceibias.n314 commonsourceibias.t113 168.701
R45 commonsourceibias.n271 commonsourceibias.t138 168.701
R46 commonsourceibias.n306 commonsourceibias.t130 168.701
R47 commonsourceibias.n300 commonsourceibias.t114 168.701
R48 commonsourceibias.n276 commonsourceibias.t139 168.701
R49 commonsourceibias.n292 commonsourceibias.t129 168.701
R50 commonsourceibias.n286 commonsourceibias.t125 168.701
R51 commonsourceibias.n280 commonsourceibias.t147 168.701
R52 commonsourceibias.n125 commonsourceibias.t20 168.701
R53 commonsourceibias.n119 commonsourceibias.t66 168.701
R54 commonsourceibias.n19 commonsourceibias.t50 168.701
R55 commonsourceibias.n111 commonsourceibias.t0 168.701
R56 commonsourceibias.n105 commonsourceibias.t56 168.701
R57 commonsourceibias.n24 commonsourceibias.t42 168.701
R58 commonsourceibias.n97 commonsourceibias.t72 168.701
R59 commonsourceibias.n91 commonsourceibias.t54 168.701
R60 commonsourceibias.n29 commonsourceibias.t34 168.701
R61 commonsourceibias.n83 commonsourceibias.t38 168.701
R62 commonsourceibias.n77 commonsourceibias.t44 168.701
R63 commonsourceibias.n34 commonsourceibias.t6 168.701
R64 commonsourceibias.n69 commonsourceibias.t58 168.701
R65 commonsourceibias.n63 commonsourceibias.t10 168.701
R66 commonsourceibias.n39 commonsourceibias.t76 168.701
R67 commonsourceibias.n55 commonsourceibias.t22 168.701
R68 commonsourceibias.n49 commonsourceibias.t32 168.701
R69 commonsourceibias.n43 commonsourceibias.t18 168.701
R70 commonsourceibias.n247 commonsourceibias.t83 168.701
R71 commonsourceibias.n241 commonsourceibias.t161 168.701
R72 commonsourceibias.n5 commonsourceibias.t152 168.701
R73 commonsourceibias.n233 commonsourceibias.t171 168.701
R74 commonsourceibias.n227 commonsourceibias.t145 168.701
R75 commonsourceibias.n10 commonsourceibias.t124 168.701
R76 commonsourceibias.n219 commonsourceibias.t158 168.701
R77 commonsourceibias.n213 commonsourceibias.t148 168.701
R78 commonsourceibias.n150 commonsourceibias.t93 168.701
R79 commonsourceibias.n151 commonsourceibias.t131 168.701
R80 commonsourceibias.n153 commonsourceibias.t117 168.701
R81 commonsourceibias.n155 commonsourceibias.t176 168.701
R82 commonsourceibias.n191 commonsourceibias.t144 168.701
R83 commonsourceibias.n185 commonsourceibias.t190 168.701
R84 commonsourceibias.n161 commonsourceibias.t164 168.701
R85 commonsourceibias.n177 commonsourceibias.t111 168.701
R86 commonsourceibias.n171 commonsourceibias.t100 168.701
R87 commonsourceibias.n165 commonsourceibias.t84 168.701
R88 commonsourceibias.n874 commonsourceibias.t156 168.701
R89 commonsourceibias.n880 commonsourceibias.t146 168.701
R90 commonsourceibias.n886 commonsourceibias.t126 168.701
R91 commonsourceibias.n888 commonsourceibias.t91 168.701
R92 commonsourceibias.n895 commonsourceibias.t181 168.701
R93 commonsourceibias.n901 commonsourceibias.t136 168.701
R94 commonsourceibias.n903 commonsourceibias.t107 168.701
R95 commonsourceibias.n910 commonsourceibias.t192 168.701
R96 commonsourceibias.n916 commonsourceibias.t167 168.701
R97 commonsourceibias.n918 commonsourceibias.t127 168.701
R98 commonsourceibias.n925 commonsourceibias.t87 168.701
R99 commonsourceibias.n931 commonsourceibias.t99 168.701
R100 commonsourceibias.n933 commonsourceibias.t137 168.701
R101 commonsourceibias.n940 commonsourceibias.t143 168.701
R102 commonsourceibias.n946 commonsourceibias.t122 168.701
R103 commonsourceibias.n948 commonsourceibias.t170 168.701
R104 commonsourceibias.n955 commonsourceibias.t153 168.701
R105 commonsourceibias.n961 commonsourceibias.t133 168.701
R106 commonsourceibias.n758 commonsourceibias.t123 168.701
R107 commonsourceibias.n764 commonsourceibias.t132 168.701
R108 commonsourceibias.n770 commonsourceibias.t104 168.701
R109 commonsourceibias.n772 commonsourceibias.t118 168.701
R110 commonsourceibias.n779 commonsourceibias.t85 168.701
R111 commonsourceibias.n785 commonsourceibias.t106 168.701
R112 commonsourceibias.n787 commonsourceibias.t119 168.701
R113 commonsourceibias.n794 commonsourceibias.t86 168.701
R114 commonsourceibias.n800 commonsourceibias.t97 168.701
R115 commonsourceibias.n802 commonsourceibias.t120 168.701
R116 commonsourceibias.n809 commonsourceibias.t89 168.701
R117 commonsourceibias.n815 commonsourceibias.t178 168.701
R118 commonsourceibias.n817 commonsourceibias.t121 168.701
R119 commonsourceibias.n824 commonsourceibias.t81 168.701
R120 commonsourceibias.n830 commonsourceibias.t179 168.701
R121 commonsourceibias.n832 commonsourceibias.t193 168.701
R122 commonsourceibias.n839 commonsourceibias.t82 168.701
R123 commonsourceibias.n845 commonsourceibias.t180 168.701
R124 commonsourceibias.n528 commonsourceibias.t70 168.701
R125 commonsourceibias.n534 commonsourceibias.t68 168.701
R126 commonsourceibias.n540 commonsourceibias.t14 168.701
R127 commonsourceibias.n542 commonsourceibias.t36 168.701
R128 commonsourceibias.n549 commonsourceibias.t78 168.701
R129 commonsourceibias.n555 commonsourceibias.t28 168.701
R130 commonsourceibias.n557 commonsourceibias.t64 168.701
R131 commonsourceibias.n564 commonsourceibias.t12 168.701
R132 commonsourceibias.n570 commonsourceibias.t30 168.701
R133 commonsourceibias.n572 commonsourceibias.t8 168.701
R134 commonsourceibias.n579 commonsourceibias.t24 168.701
R135 commonsourceibias.n585 commonsourceibias.t40 168.701
R136 commonsourceibias.n587 commonsourceibias.t16 168.701
R137 commonsourceibias.n594 commonsourceibias.t26 168.701
R138 commonsourceibias.n600 commonsourceibias.t74 168.701
R139 commonsourceibias.n602 commonsourceibias.t46 168.701
R140 commonsourceibias.n609 commonsourceibias.t60 168.701
R141 commonsourceibias.n615 commonsourceibias.t2 168.701
R142 commonsourceibias.n730 commonsourceibias.t169 168.701
R143 commonsourceibias.n724 commonsourceibias.t142 168.701
R144 commonsourceibias.n717 commonsourceibias.t116 168.701
R145 commonsourceibias.n715 commonsourceibias.t154 168.701
R146 commonsourceibias.n709 commonsourceibias.t108 168.701
R147 commonsourceibias.n702 commonsourceibias.t90 168.701
R148 commonsourceibias.n700 commonsourceibias.t128 168.701
R149 commonsourceibias.n694 commonsourceibias.t109 168.701
R150 commonsourceibias.n687 commonsourceibias.t174 168.701
R151 commonsourceibias.n644 commonsourceibias.t159 168.701
R152 commonsourceibias.n650 commonsourceibias.t160 168.701
R153 commonsourceibias.n656 commonsourceibias.t185 168.701
R154 commonsourceibias.n658 commonsourceibias.t135 168.701
R155 commonsourceibias.n665 commonsourceibias.t166 168.701
R156 commonsourceibias.n671 commonsourceibias.t103 168.701
R157 commonsourceibias.n635 commonsourceibias.t162 168.701
R158 commonsourceibias.n633 commonsourceibias.t188 168.701
R159 commonsourceibias.n631 commonsourceibias.t102 168.701
R160 commonsourceibias.n479 commonsourceibias.n367 161.3
R161 commonsourceibias.n477 commonsourceibias.n476 161.3
R162 commonsourceibias.n475 commonsourceibias.n368 161.3
R163 commonsourceibias.n474 commonsourceibias.n473 161.3
R164 commonsourceibias.n471 commonsourceibias.n369 161.3
R165 commonsourceibias.n470 commonsourceibias.n469 161.3
R166 commonsourceibias.n468 commonsourceibias.n370 161.3
R167 commonsourceibias.n467 commonsourceibias.n466 161.3
R168 commonsourceibias.n465 commonsourceibias.n371 161.3
R169 commonsourceibias.n463 commonsourceibias.n462 161.3
R170 commonsourceibias.n461 commonsourceibias.n373 161.3
R171 commonsourceibias.n460 commonsourceibias.n459 161.3
R172 commonsourceibias.n457 commonsourceibias.n374 161.3
R173 commonsourceibias.n456 commonsourceibias.n455 161.3
R174 commonsourceibias.n454 commonsourceibias.n375 161.3
R175 commonsourceibias.n453 commonsourceibias.n452 161.3
R176 commonsourceibias.n451 commonsourceibias.n376 161.3
R177 commonsourceibias.n449 commonsourceibias.n448 161.3
R178 commonsourceibias.n447 commonsourceibias.n378 161.3
R179 commonsourceibias.n446 commonsourceibias.n445 161.3
R180 commonsourceibias.n443 commonsourceibias.n379 161.3
R181 commonsourceibias.n442 commonsourceibias.n441 161.3
R182 commonsourceibias.n440 commonsourceibias.n380 161.3
R183 commonsourceibias.n439 commonsourceibias.n438 161.3
R184 commonsourceibias.n437 commonsourceibias.n381 161.3
R185 commonsourceibias.n435 commonsourceibias.n434 161.3
R186 commonsourceibias.n433 commonsourceibias.n383 161.3
R187 commonsourceibias.n432 commonsourceibias.n431 161.3
R188 commonsourceibias.n429 commonsourceibias.n384 161.3
R189 commonsourceibias.n428 commonsourceibias.n427 161.3
R190 commonsourceibias.n426 commonsourceibias.n385 161.3
R191 commonsourceibias.n425 commonsourceibias.n424 161.3
R192 commonsourceibias.n423 commonsourceibias.n386 161.3
R193 commonsourceibias.n421 commonsourceibias.n420 161.3
R194 commonsourceibias.n419 commonsourceibias.n388 161.3
R195 commonsourceibias.n418 commonsourceibias.n417 161.3
R196 commonsourceibias.n415 commonsourceibias.n389 161.3
R197 commonsourceibias.n414 commonsourceibias.n413 161.3
R198 commonsourceibias.n412 commonsourceibias.n390 161.3
R199 commonsourceibias.n411 commonsourceibias.n410 161.3
R200 commonsourceibias.n409 commonsourceibias.n391 161.3
R201 commonsourceibias.n407 commonsourceibias.n406 161.3
R202 commonsourceibias.n405 commonsourceibias.n393 161.3
R203 commonsourceibias.n404 commonsourceibias.n403 161.3
R204 commonsourceibias.n401 commonsourceibias.n394 161.3
R205 commonsourceibias.n400 commonsourceibias.n399 161.3
R206 commonsourceibias.n398 commonsourceibias.n395 161.3
R207 commonsourceibias.n282 commonsourceibias.n279 161.3
R208 commonsourceibias.n284 commonsourceibias.n283 161.3
R209 commonsourceibias.n285 commonsourceibias.n278 161.3
R210 commonsourceibias.n288 commonsourceibias.n287 161.3
R211 commonsourceibias.n289 commonsourceibias.n277 161.3
R212 commonsourceibias.n291 commonsourceibias.n290 161.3
R213 commonsourceibias.n293 commonsourceibias.n275 161.3
R214 commonsourceibias.n295 commonsourceibias.n294 161.3
R215 commonsourceibias.n296 commonsourceibias.n274 161.3
R216 commonsourceibias.n298 commonsourceibias.n297 161.3
R217 commonsourceibias.n299 commonsourceibias.n273 161.3
R218 commonsourceibias.n302 commonsourceibias.n301 161.3
R219 commonsourceibias.n303 commonsourceibias.n272 161.3
R220 commonsourceibias.n305 commonsourceibias.n304 161.3
R221 commonsourceibias.n307 commonsourceibias.n270 161.3
R222 commonsourceibias.n309 commonsourceibias.n308 161.3
R223 commonsourceibias.n310 commonsourceibias.n269 161.3
R224 commonsourceibias.n312 commonsourceibias.n311 161.3
R225 commonsourceibias.n313 commonsourceibias.n268 161.3
R226 commonsourceibias.n316 commonsourceibias.n315 161.3
R227 commonsourceibias.n317 commonsourceibias.n267 161.3
R228 commonsourceibias.n319 commonsourceibias.n318 161.3
R229 commonsourceibias.n321 commonsourceibias.n265 161.3
R230 commonsourceibias.n323 commonsourceibias.n322 161.3
R231 commonsourceibias.n324 commonsourceibias.n264 161.3
R232 commonsourceibias.n326 commonsourceibias.n325 161.3
R233 commonsourceibias.n327 commonsourceibias.n263 161.3
R234 commonsourceibias.n330 commonsourceibias.n329 161.3
R235 commonsourceibias.n331 commonsourceibias.n262 161.3
R236 commonsourceibias.n333 commonsourceibias.n332 161.3
R237 commonsourceibias.n335 commonsourceibias.n260 161.3
R238 commonsourceibias.n337 commonsourceibias.n336 161.3
R239 commonsourceibias.n338 commonsourceibias.n259 161.3
R240 commonsourceibias.n340 commonsourceibias.n339 161.3
R241 commonsourceibias.n341 commonsourceibias.n258 161.3
R242 commonsourceibias.n344 commonsourceibias.n343 161.3
R243 commonsourceibias.n345 commonsourceibias.n257 161.3
R244 commonsourceibias.n347 commonsourceibias.n346 161.3
R245 commonsourceibias.n349 commonsourceibias.n255 161.3
R246 commonsourceibias.n351 commonsourceibias.n350 161.3
R247 commonsourceibias.n352 commonsourceibias.n254 161.3
R248 commonsourceibias.n354 commonsourceibias.n353 161.3
R249 commonsourceibias.n355 commonsourceibias.n253 161.3
R250 commonsourceibias.n358 commonsourceibias.n357 161.3
R251 commonsourceibias.n359 commonsourceibias.n252 161.3
R252 commonsourceibias.n361 commonsourceibias.n360 161.3
R253 commonsourceibias.n363 commonsourceibias.n251 161.3
R254 commonsourceibias.n45 commonsourceibias.n42 161.3
R255 commonsourceibias.n47 commonsourceibias.n46 161.3
R256 commonsourceibias.n48 commonsourceibias.n41 161.3
R257 commonsourceibias.n51 commonsourceibias.n50 161.3
R258 commonsourceibias.n52 commonsourceibias.n40 161.3
R259 commonsourceibias.n54 commonsourceibias.n53 161.3
R260 commonsourceibias.n56 commonsourceibias.n38 161.3
R261 commonsourceibias.n58 commonsourceibias.n57 161.3
R262 commonsourceibias.n59 commonsourceibias.n37 161.3
R263 commonsourceibias.n61 commonsourceibias.n60 161.3
R264 commonsourceibias.n62 commonsourceibias.n36 161.3
R265 commonsourceibias.n65 commonsourceibias.n64 161.3
R266 commonsourceibias.n66 commonsourceibias.n35 161.3
R267 commonsourceibias.n68 commonsourceibias.n67 161.3
R268 commonsourceibias.n70 commonsourceibias.n33 161.3
R269 commonsourceibias.n72 commonsourceibias.n71 161.3
R270 commonsourceibias.n73 commonsourceibias.n32 161.3
R271 commonsourceibias.n75 commonsourceibias.n74 161.3
R272 commonsourceibias.n76 commonsourceibias.n31 161.3
R273 commonsourceibias.n79 commonsourceibias.n78 161.3
R274 commonsourceibias.n80 commonsourceibias.n30 161.3
R275 commonsourceibias.n82 commonsourceibias.n81 161.3
R276 commonsourceibias.n84 commonsourceibias.n28 161.3
R277 commonsourceibias.n86 commonsourceibias.n85 161.3
R278 commonsourceibias.n87 commonsourceibias.n27 161.3
R279 commonsourceibias.n89 commonsourceibias.n88 161.3
R280 commonsourceibias.n90 commonsourceibias.n26 161.3
R281 commonsourceibias.n93 commonsourceibias.n92 161.3
R282 commonsourceibias.n94 commonsourceibias.n25 161.3
R283 commonsourceibias.n96 commonsourceibias.n95 161.3
R284 commonsourceibias.n98 commonsourceibias.n23 161.3
R285 commonsourceibias.n100 commonsourceibias.n99 161.3
R286 commonsourceibias.n101 commonsourceibias.n22 161.3
R287 commonsourceibias.n103 commonsourceibias.n102 161.3
R288 commonsourceibias.n104 commonsourceibias.n21 161.3
R289 commonsourceibias.n107 commonsourceibias.n106 161.3
R290 commonsourceibias.n108 commonsourceibias.n20 161.3
R291 commonsourceibias.n110 commonsourceibias.n109 161.3
R292 commonsourceibias.n112 commonsourceibias.n18 161.3
R293 commonsourceibias.n114 commonsourceibias.n113 161.3
R294 commonsourceibias.n115 commonsourceibias.n17 161.3
R295 commonsourceibias.n117 commonsourceibias.n116 161.3
R296 commonsourceibias.n118 commonsourceibias.n16 161.3
R297 commonsourceibias.n121 commonsourceibias.n120 161.3
R298 commonsourceibias.n122 commonsourceibias.n15 161.3
R299 commonsourceibias.n124 commonsourceibias.n123 161.3
R300 commonsourceibias.n126 commonsourceibias.n14 161.3
R301 commonsourceibias.n167 commonsourceibias.n164 161.3
R302 commonsourceibias.n169 commonsourceibias.n168 161.3
R303 commonsourceibias.n170 commonsourceibias.n163 161.3
R304 commonsourceibias.n173 commonsourceibias.n172 161.3
R305 commonsourceibias.n174 commonsourceibias.n162 161.3
R306 commonsourceibias.n176 commonsourceibias.n175 161.3
R307 commonsourceibias.n178 commonsourceibias.n160 161.3
R308 commonsourceibias.n180 commonsourceibias.n179 161.3
R309 commonsourceibias.n181 commonsourceibias.n159 161.3
R310 commonsourceibias.n183 commonsourceibias.n182 161.3
R311 commonsourceibias.n184 commonsourceibias.n158 161.3
R312 commonsourceibias.n187 commonsourceibias.n186 161.3
R313 commonsourceibias.n188 commonsourceibias.n157 161.3
R314 commonsourceibias.n190 commonsourceibias.n189 161.3
R315 commonsourceibias.n192 commonsourceibias.n156 161.3
R316 commonsourceibias.n194 commonsourceibias.n193 161.3
R317 commonsourceibias.n196 commonsourceibias.n195 161.3
R318 commonsourceibias.n197 commonsourceibias.n154 161.3
R319 commonsourceibias.n199 commonsourceibias.n198 161.3
R320 commonsourceibias.n201 commonsourceibias.n200 161.3
R321 commonsourceibias.n202 commonsourceibias.n152 161.3
R322 commonsourceibias.n204 commonsourceibias.n203 161.3
R323 commonsourceibias.n206 commonsourceibias.n205 161.3
R324 commonsourceibias.n208 commonsourceibias.n207 161.3
R325 commonsourceibias.n209 commonsourceibias.n13 161.3
R326 commonsourceibias.n211 commonsourceibias.n210 161.3
R327 commonsourceibias.n212 commonsourceibias.n12 161.3
R328 commonsourceibias.n215 commonsourceibias.n214 161.3
R329 commonsourceibias.n216 commonsourceibias.n11 161.3
R330 commonsourceibias.n218 commonsourceibias.n217 161.3
R331 commonsourceibias.n220 commonsourceibias.n9 161.3
R332 commonsourceibias.n222 commonsourceibias.n221 161.3
R333 commonsourceibias.n223 commonsourceibias.n8 161.3
R334 commonsourceibias.n225 commonsourceibias.n224 161.3
R335 commonsourceibias.n226 commonsourceibias.n7 161.3
R336 commonsourceibias.n229 commonsourceibias.n228 161.3
R337 commonsourceibias.n230 commonsourceibias.n6 161.3
R338 commonsourceibias.n232 commonsourceibias.n231 161.3
R339 commonsourceibias.n234 commonsourceibias.n4 161.3
R340 commonsourceibias.n236 commonsourceibias.n235 161.3
R341 commonsourceibias.n237 commonsourceibias.n3 161.3
R342 commonsourceibias.n239 commonsourceibias.n238 161.3
R343 commonsourceibias.n240 commonsourceibias.n2 161.3
R344 commonsourceibias.n243 commonsourceibias.n242 161.3
R345 commonsourceibias.n244 commonsourceibias.n1 161.3
R346 commonsourceibias.n246 commonsourceibias.n245 161.3
R347 commonsourceibias.n248 commonsourceibias.n0 161.3
R348 commonsourceibias.n962 commonsourceibias.n850 161.3
R349 commonsourceibias.n960 commonsourceibias.n959 161.3
R350 commonsourceibias.n958 commonsourceibias.n851 161.3
R351 commonsourceibias.n957 commonsourceibias.n956 161.3
R352 commonsourceibias.n954 commonsourceibias.n852 161.3
R353 commonsourceibias.n953 commonsourceibias.n952 161.3
R354 commonsourceibias.n951 commonsourceibias.n853 161.3
R355 commonsourceibias.n950 commonsourceibias.n949 161.3
R356 commonsourceibias.n947 commonsourceibias.n854 161.3
R357 commonsourceibias.n945 commonsourceibias.n944 161.3
R358 commonsourceibias.n943 commonsourceibias.n855 161.3
R359 commonsourceibias.n942 commonsourceibias.n941 161.3
R360 commonsourceibias.n939 commonsourceibias.n856 161.3
R361 commonsourceibias.n938 commonsourceibias.n937 161.3
R362 commonsourceibias.n936 commonsourceibias.n857 161.3
R363 commonsourceibias.n935 commonsourceibias.n934 161.3
R364 commonsourceibias.n932 commonsourceibias.n858 161.3
R365 commonsourceibias.n930 commonsourceibias.n929 161.3
R366 commonsourceibias.n928 commonsourceibias.n859 161.3
R367 commonsourceibias.n927 commonsourceibias.n926 161.3
R368 commonsourceibias.n924 commonsourceibias.n860 161.3
R369 commonsourceibias.n923 commonsourceibias.n922 161.3
R370 commonsourceibias.n921 commonsourceibias.n861 161.3
R371 commonsourceibias.n920 commonsourceibias.n919 161.3
R372 commonsourceibias.n917 commonsourceibias.n862 161.3
R373 commonsourceibias.n915 commonsourceibias.n914 161.3
R374 commonsourceibias.n913 commonsourceibias.n863 161.3
R375 commonsourceibias.n912 commonsourceibias.n911 161.3
R376 commonsourceibias.n909 commonsourceibias.n864 161.3
R377 commonsourceibias.n908 commonsourceibias.n907 161.3
R378 commonsourceibias.n906 commonsourceibias.n865 161.3
R379 commonsourceibias.n905 commonsourceibias.n904 161.3
R380 commonsourceibias.n902 commonsourceibias.n866 161.3
R381 commonsourceibias.n900 commonsourceibias.n899 161.3
R382 commonsourceibias.n898 commonsourceibias.n867 161.3
R383 commonsourceibias.n897 commonsourceibias.n896 161.3
R384 commonsourceibias.n894 commonsourceibias.n868 161.3
R385 commonsourceibias.n893 commonsourceibias.n892 161.3
R386 commonsourceibias.n891 commonsourceibias.n869 161.3
R387 commonsourceibias.n890 commonsourceibias.n889 161.3
R388 commonsourceibias.n887 commonsourceibias.n870 161.3
R389 commonsourceibias.n885 commonsourceibias.n884 161.3
R390 commonsourceibias.n883 commonsourceibias.n871 161.3
R391 commonsourceibias.n882 commonsourceibias.n881 161.3
R392 commonsourceibias.n879 commonsourceibias.n872 161.3
R393 commonsourceibias.n878 commonsourceibias.n877 161.3
R394 commonsourceibias.n876 commonsourceibias.n873 161.3
R395 commonsourceibias.n846 commonsourceibias.n734 161.3
R396 commonsourceibias.n844 commonsourceibias.n843 161.3
R397 commonsourceibias.n842 commonsourceibias.n735 161.3
R398 commonsourceibias.n841 commonsourceibias.n840 161.3
R399 commonsourceibias.n838 commonsourceibias.n736 161.3
R400 commonsourceibias.n837 commonsourceibias.n836 161.3
R401 commonsourceibias.n835 commonsourceibias.n737 161.3
R402 commonsourceibias.n834 commonsourceibias.n833 161.3
R403 commonsourceibias.n831 commonsourceibias.n738 161.3
R404 commonsourceibias.n829 commonsourceibias.n828 161.3
R405 commonsourceibias.n827 commonsourceibias.n739 161.3
R406 commonsourceibias.n826 commonsourceibias.n825 161.3
R407 commonsourceibias.n823 commonsourceibias.n740 161.3
R408 commonsourceibias.n822 commonsourceibias.n821 161.3
R409 commonsourceibias.n820 commonsourceibias.n741 161.3
R410 commonsourceibias.n819 commonsourceibias.n818 161.3
R411 commonsourceibias.n816 commonsourceibias.n742 161.3
R412 commonsourceibias.n814 commonsourceibias.n813 161.3
R413 commonsourceibias.n812 commonsourceibias.n743 161.3
R414 commonsourceibias.n811 commonsourceibias.n810 161.3
R415 commonsourceibias.n808 commonsourceibias.n744 161.3
R416 commonsourceibias.n807 commonsourceibias.n806 161.3
R417 commonsourceibias.n805 commonsourceibias.n745 161.3
R418 commonsourceibias.n804 commonsourceibias.n803 161.3
R419 commonsourceibias.n801 commonsourceibias.n746 161.3
R420 commonsourceibias.n799 commonsourceibias.n798 161.3
R421 commonsourceibias.n797 commonsourceibias.n747 161.3
R422 commonsourceibias.n796 commonsourceibias.n795 161.3
R423 commonsourceibias.n793 commonsourceibias.n748 161.3
R424 commonsourceibias.n792 commonsourceibias.n791 161.3
R425 commonsourceibias.n790 commonsourceibias.n749 161.3
R426 commonsourceibias.n789 commonsourceibias.n788 161.3
R427 commonsourceibias.n786 commonsourceibias.n750 161.3
R428 commonsourceibias.n784 commonsourceibias.n783 161.3
R429 commonsourceibias.n782 commonsourceibias.n751 161.3
R430 commonsourceibias.n781 commonsourceibias.n780 161.3
R431 commonsourceibias.n778 commonsourceibias.n752 161.3
R432 commonsourceibias.n777 commonsourceibias.n776 161.3
R433 commonsourceibias.n775 commonsourceibias.n753 161.3
R434 commonsourceibias.n774 commonsourceibias.n773 161.3
R435 commonsourceibias.n771 commonsourceibias.n754 161.3
R436 commonsourceibias.n769 commonsourceibias.n768 161.3
R437 commonsourceibias.n767 commonsourceibias.n755 161.3
R438 commonsourceibias.n766 commonsourceibias.n765 161.3
R439 commonsourceibias.n763 commonsourceibias.n756 161.3
R440 commonsourceibias.n762 commonsourceibias.n761 161.3
R441 commonsourceibias.n760 commonsourceibias.n757 161.3
R442 commonsourceibias.n616 commonsourceibias.n504 161.3
R443 commonsourceibias.n614 commonsourceibias.n613 161.3
R444 commonsourceibias.n612 commonsourceibias.n505 161.3
R445 commonsourceibias.n611 commonsourceibias.n610 161.3
R446 commonsourceibias.n608 commonsourceibias.n506 161.3
R447 commonsourceibias.n607 commonsourceibias.n606 161.3
R448 commonsourceibias.n605 commonsourceibias.n507 161.3
R449 commonsourceibias.n604 commonsourceibias.n603 161.3
R450 commonsourceibias.n601 commonsourceibias.n508 161.3
R451 commonsourceibias.n599 commonsourceibias.n598 161.3
R452 commonsourceibias.n597 commonsourceibias.n509 161.3
R453 commonsourceibias.n596 commonsourceibias.n595 161.3
R454 commonsourceibias.n593 commonsourceibias.n510 161.3
R455 commonsourceibias.n592 commonsourceibias.n591 161.3
R456 commonsourceibias.n590 commonsourceibias.n511 161.3
R457 commonsourceibias.n589 commonsourceibias.n588 161.3
R458 commonsourceibias.n586 commonsourceibias.n512 161.3
R459 commonsourceibias.n584 commonsourceibias.n583 161.3
R460 commonsourceibias.n582 commonsourceibias.n513 161.3
R461 commonsourceibias.n581 commonsourceibias.n580 161.3
R462 commonsourceibias.n578 commonsourceibias.n514 161.3
R463 commonsourceibias.n577 commonsourceibias.n576 161.3
R464 commonsourceibias.n575 commonsourceibias.n515 161.3
R465 commonsourceibias.n574 commonsourceibias.n573 161.3
R466 commonsourceibias.n571 commonsourceibias.n516 161.3
R467 commonsourceibias.n569 commonsourceibias.n568 161.3
R468 commonsourceibias.n567 commonsourceibias.n517 161.3
R469 commonsourceibias.n566 commonsourceibias.n565 161.3
R470 commonsourceibias.n563 commonsourceibias.n518 161.3
R471 commonsourceibias.n562 commonsourceibias.n561 161.3
R472 commonsourceibias.n560 commonsourceibias.n519 161.3
R473 commonsourceibias.n559 commonsourceibias.n558 161.3
R474 commonsourceibias.n556 commonsourceibias.n520 161.3
R475 commonsourceibias.n554 commonsourceibias.n553 161.3
R476 commonsourceibias.n552 commonsourceibias.n521 161.3
R477 commonsourceibias.n551 commonsourceibias.n550 161.3
R478 commonsourceibias.n548 commonsourceibias.n522 161.3
R479 commonsourceibias.n547 commonsourceibias.n546 161.3
R480 commonsourceibias.n545 commonsourceibias.n523 161.3
R481 commonsourceibias.n544 commonsourceibias.n543 161.3
R482 commonsourceibias.n541 commonsourceibias.n524 161.3
R483 commonsourceibias.n539 commonsourceibias.n538 161.3
R484 commonsourceibias.n537 commonsourceibias.n525 161.3
R485 commonsourceibias.n536 commonsourceibias.n535 161.3
R486 commonsourceibias.n533 commonsourceibias.n526 161.3
R487 commonsourceibias.n532 commonsourceibias.n531 161.3
R488 commonsourceibias.n530 commonsourceibias.n527 161.3
R489 commonsourceibias.n686 commonsourceibias.n685 161.3
R490 commonsourceibias.n684 commonsourceibias.n683 161.3
R491 commonsourceibias.n682 commonsourceibias.n632 161.3
R492 commonsourceibias.n681 commonsourceibias.n680 161.3
R493 commonsourceibias.n679 commonsourceibias.n678 161.3
R494 commonsourceibias.n677 commonsourceibias.n634 161.3
R495 commonsourceibias.n676 commonsourceibias.n675 161.3
R496 commonsourceibias.n674 commonsourceibias.n673 161.3
R497 commonsourceibias.n672 commonsourceibias.n636 161.3
R498 commonsourceibias.n670 commonsourceibias.n669 161.3
R499 commonsourceibias.n668 commonsourceibias.n637 161.3
R500 commonsourceibias.n667 commonsourceibias.n666 161.3
R501 commonsourceibias.n664 commonsourceibias.n638 161.3
R502 commonsourceibias.n663 commonsourceibias.n662 161.3
R503 commonsourceibias.n661 commonsourceibias.n639 161.3
R504 commonsourceibias.n660 commonsourceibias.n659 161.3
R505 commonsourceibias.n657 commonsourceibias.n640 161.3
R506 commonsourceibias.n655 commonsourceibias.n654 161.3
R507 commonsourceibias.n653 commonsourceibias.n641 161.3
R508 commonsourceibias.n652 commonsourceibias.n651 161.3
R509 commonsourceibias.n649 commonsourceibias.n642 161.3
R510 commonsourceibias.n648 commonsourceibias.n647 161.3
R511 commonsourceibias.n646 commonsourceibias.n643 161.3
R512 commonsourceibias.n731 commonsourceibias.n483 161.3
R513 commonsourceibias.n729 commonsourceibias.n728 161.3
R514 commonsourceibias.n727 commonsourceibias.n484 161.3
R515 commonsourceibias.n726 commonsourceibias.n725 161.3
R516 commonsourceibias.n723 commonsourceibias.n485 161.3
R517 commonsourceibias.n722 commonsourceibias.n721 161.3
R518 commonsourceibias.n720 commonsourceibias.n486 161.3
R519 commonsourceibias.n719 commonsourceibias.n718 161.3
R520 commonsourceibias.n716 commonsourceibias.n487 161.3
R521 commonsourceibias.n714 commonsourceibias.n713 161.3
R522 commonsourceibias.n712 commonsourceibias.n488 161.3
R523 commonsourceibias.n711 commonsourceibias.n710 161.3
R524 commonsourceibias.n708 commonsourceibias.n489 161.3
R525 commonsourceibias.n707 commonsourceibias.n706 161.3
R526 commonsourceibias.n705 commonsourceibias.n490 161.3
R527 commonsourceibias.n704 commonsourceibias.n703 161.3
R528 commonsourceibias.n701 commonsourceibias.n491 161.3
R529 commonsourceibias.n699 commonsourceibias.n698 161.3
R530 commonsourceibias.n697 commonsourceibias.n492 161.3
R531 commonsourceibias.n696 commonsourceibias.n695 161.3
R532 commonsourceibias.n693 commonsourceibias.n493 161.3
R533 commonsourceibias.n692 commonsourceibias.n691 161.3
R534 commonsourceibias.n690 commonsourceibias.n494 161.3
R535 commonsourceibias.n689 commonsourceibias.n688 161.3
R536 commonsourceibias.n141 commonsourceibias.n139 81.5057
R537 commonsourceibias.n497 commonsourceibias.n495 81.5057
R538 commonsourceibias.n141 commonsourceibias.n140 80.9324
R539 commonsourceibias.n143 commonsourceibias.n142 80.9324
R540 commonsourceibias.n145 commonsourceibias.n144 80.9324
R541 commonsourceibias.n147 commonsourceibias.n146 80.9324
R542 commonsourceibias.n138 commonsourceibias.n137 80.9324
R543 commonsourceibias.n136 commonsourceibias.n135 80.9324
R544 commonsourceibias.n134 commonsourceibias.n133 80.9324
R545 commonsourceibias.n132 commonsourceibias.n131 80.9324
R546 commonsourceibias.n130 commonsourceibias.n129 80.9324
R547 commonsourceibias.n620 commonsourceibias.n619 80.9324
R548 commonsourceibias.n622 commonsourceibias.n621 80.9324
R549 commonsourceibias.n624 commonsourceibias.n623 80.9324
R550 commonsourceibias.n626 commonsourceibias.n625 80.9324
R551 commonsourceibias.n628 commonsourceibias.n627 80.9324
R552 commonsourceibias.n503 commonsourceibias.n502 80.9324
R553 commonsourceibias.n501 commonsourceibias.n500 80.9324
R554 commonsourceibias.n499 commonsourceibias.n498 80.9324
R555 commonsourceibias.n497 commonsourceibias.n496 80.9324
R556 commonsourceibias.n481 commonsourceibias.n480 80.6037
R557 commonsourceibias.n365 commonsourceibias.n364 80.6037
R558 commonsourceibias.n128 commonsourceibias.n127 80.6037
R559 commonsourceibias.n250 commonsourceibias.n249 80.6037
R560 commonsourceibias.n964 commonsourceibias.n963 80.6037
R561 commonsourceibias.n848 commonsourceibias.n847 80.6037
R562 commonsourceibias.n618 commonsourceibias.n617 80.6037
R563 commonsourceibias.n733 commonsourceibias.n732 80.6037
R564 commonsourceibias.n438 commonsourceibias.n437 56.5617
R565 commonsourceibias.n452 commonsourceibias.n451 56.5617
R566 commonsourceibias.n322 commonsourceibias.n321 56.5617
R567 commonsourceibias.n308 commonsourceibias.n307 56.5617
R568 commonsourceibias.n85 commonsourceibias.n84 56.5617
R569 commonsourceibias.n71 commonsourceibias.n70 56.5617
R570 commonsourceibias.n207 commonsourceibias.n206 56.5617
R571 commonsourceibias.n193 commonsourceibias.n192 56.5617
R572 commonsourceibias.n919 commonsourceibias.n917 56.5617
R573 commonsourceibias.n934 commonsourceibias.n932 56.5617
R574 commonsourceibias.n803 commonsourceibias.n801 56.5617
R575 commonsourceibias.n818 commonsourceibias.n816 56.5617
R576 commonsourceibias.n573 commonsourceibias.n571 56.5617
R577 commonsourceibias.n588 commonsourceibias.n586 56.5617
R578 commonsourceibias.n688 commonsourceibias.n686 56.5617
R579 commonsourceibias.n410 commonsourceibias.n409 56.5617
R580 commonsourceibias.n424 commonsourceibias.n423 56.5617
R581 commonsourceibias.n466 commonsourceibias.n465 56.5617
R582 commonsourceibias.n350 commonsourceibias.n349 56.5617
R583 commonsourceibias.n336 commonsourceibias.n335 56.5617
R584 commonsourceibias.n294 commonsourceibias.n293 56.5617
R585 commonsourceibias.n113 commonsourceibias.n112 56.5617
R586 commonsourceibias.n99 commonsourceibias.n98 56.5617
R587 commonsourceibias.n57 commonsourceibias.n56 56.5617
R588 commonsourceibias.n235 commonsourceibias.n234 56.5617
R589 commonsourceibias.n221 commonsourceibias.n220 56.5617
R590 commonsourceibias.n179 commonsourceibias.n178 56.5617
R591 commonsourceibias.n889 commonsourceibias.n887 56.5617
R592 commonsourceibias.n904 commonsourceibias.n902 56.5617
R593 commonsourceibias.n949 commonsourceibias.n947 56.5617
R594 commonsourceibias.n773 commonsourceibias.n771 56.5617
R595 commonsourceibias.n788 commonsourceibias.n786 56.5617
R596 commonsourceibias.n833 commonsourceibias.n831 56.5617
R597 commonsourceibias.n543 commonsourceibias.n541 56.5617
R598 commonsourceibias.n558 commonsourceibias.n556 56.5617
R599 commonsourceibias.n603 commonsourceibias.n601 56.5617
R600 commonsourceibias.n718 commonsourceibias.n716 56.5617
R601 commonsourceibias.n703 commonsourceibias.n701 56.5617
R602 commonsourceibias.n659 commonsourceibias.n657 56.5617
R603 commonsourceibias.n673 commonsourceibias.n672 56.5617
R604 commonsourceibias.n401 commonsourceibias.n400 51.2335
R605 commonsourceibias.n473 commonsourceibias.n368 51.2335
R606 commonsourceibias.n357 commonsourceibias.n252 51.2335
R607 commonsourceibias.n285 commonsourceibias.n284 51.2335
R608 commonsourceibias.n120 commonsourceibias.n15 51.2335
R609 commonsourceibias.n48 commonsourceibias.n47 51.2335
R610 commonsourceibias.n242 commonsourceibias.n1 51.2335
R611 commonsourceibias.n170 commonsourceibias.n169 51.2335
R612 commonsourceibias.n879 commonsourceibias.n878 51.2335
R613 commonsourceibias.n956 commonsourceibias.n851 51.2335
R614 commonsourceibias.n763 commonsourceibias.n762 51.2335
R615 commonsourceibias.n840 commonsourceibias.n735 51.2335
R616 commonsourceibias.n533 commonsourceibias.n532 51.2335
R617 commonsourceibias.n610 commonsourceibias.n505 51.2335
R618 commonsourceibias.n725 commonsourceibias.n484 51.2335
R619 commonsourceibias.n649 commonsourceibias.n648 51.2335
R620 commonsourceibias.n480 commonsourceibias.n479 50.9056
R621 commonsourceibias.n364 commonsourceibias.n363 50.9056
R622 commonsourceibias.n127 commonsourceibias.n126 50.9056
R623 commonsourceibias.n249 commonsourceibias.n248 50.9056
R624 commonsourceibias.n963 commonsourceibias.n962 50.9056
R625 commonsourceibias.n847 commonsourceibias.n846 50.9056
R626 commonsourceibias.n617 commonsourceibias.n616 50.9056
R627 commonsourceibias.n732 commonsourceibias.n731 50.9056
R628 commonsourceibias.n415 commonsourceibias.n414 50.2647
R629 commonsourceibias.n459 commonsourceibias.n373 50.2647
R630 commonsourceibias.n343 commonsourceibias.n257 50.2647
R631 commonsourceibias.n299 commonsourceibias.n298 50.2647
R632 commonsourceibias.n106 commonsourceibias.n20 50.2647
R633 commonsourceibias.n62 commonsourceibias.n61 50.2647
R634 commonsourceibias.n228 commonsourceibias.n6 50.2647
R635 commonsourceibias.n184 commonsourceibias.n183 50.2647
R636 commonsourceibias.n894 commonsourceibias.n893 50.2647
R637 commonsourceibias.n941 commonsourceibias.n855 50.2647
R638 commonsourceibias.n778 commonsourceibias.n777 50.2647
R639 commonsourceibias.n825 commonsourceibias.n739 50.2647
R640 commonsourceibias.n548 commonsourceibias.n547 50.2647
R641 commonsourceibias.n595 commonsourceibias.n509 50.2647
R642 commonsourceibias.n710 commonsourceibias.n488 50.2647
R643 commonsourceibias.n664 commonsourceibias.n663 50.2647
R644 commonsourceibias.n397 commonsourceibias.n396 49.9027
R645 commonsourceibias.n281 commonsourceibias.n280 49.9027
R646 commonsourceibias.n44 commonsourceibias.n43 49.9027
R647 commonsourceibias.n166 commonsourceibias.n165 49.9027
R648 commonsourceibias.n875 commonsourceibias.n874 49.9027
R649 commonsourceibias.n759 commonsourceibias.n758 49.9027
R650 commonsourceibias.n529 commonsourceibias.n528 49.9027
R651 commonsourceibias.n645 commonsourceibias.n644 49.9027
R652 commonsourceibias.n429 commonsourceibias.n428 49.296
R653 commonsourceibias.n445 commonsourceibias.n378 49.296
R654 commonsourceibias.n329 commonsourceibias.n262 49.296
R655 commonsourceibias.n313 commonsourceibias.n312 49.296
R656 commonsourceibias.n92 commonsourceibias.n25 49.296
R657 commonsourceibias.n76 commonsourceibias.n75 49.296
R658 commonsourceibias.n214 commonsourceibias.n11 49.296
R659 commonsourceibias.n198 commonsourceibias.n197 49.296
R660 commonsourceibias.n909 commonsourceibias.n908 49.296
R661 commonsourceibias.n926 commonsourceibias.n859 49.296
R662 commonsourceibias.n793 commonsourceibias.n792 49.296
R663 commonsourceibias.n810 commonsourceibias.n743 49.296
R664 commonsourceibias.n563 commonsourceibias.n562 49.296
R665 commonsourceibias.n580 commonsourceibias.n513 49.296
R666 commonsourceibias.n695 commonsourceibias.n492 49.296
R667 commonsourceibias.n678 commonsourceibias.n677 49.296
R668 commonsourceibias.n431 commonsourceibias.n383 48.3272
R669 commonsourceibias.n443 commonsourceibias.n442 48.3272
R670 commonsourceibias.n327 commonsourceibias.n326 48.3272
R671 commonsourceibias.n315 commonsourceibias.n267 48.3272
R672 commonsourceibias.n90 commonsourceibias.n89 48.3272
R673 commonsourceibias.n78 commonsourceibias.n30 48.3272
R674 commonsourceibias.n212 commonsourceibias.n211 48.3272
R675 commonsourceibias.n202 commonsourceibias.n201 48.3272
R676 commonsourceibias.n911 commonsourceibias.n863 48.3272
R677 commonsourceibias.n924 commonsourceibias.n923 48.3272
R678 commonsourceibias.n795 commonsourceibias.n747 48.3272
R679 commonsourceibias.n808 commonsourceibias.n807 48.3272
R680 commonsourceibias.n565 commonsourceibias.n517 48.3272
R681 commonsourceibias.n578 commonsourceibias.n577 48.3272
R682 commonsourceibias.n693 commonsourceibias.n692 48.3272
R683 commonsourceibias.n682 commonsourceibias.n681 48.3272
R684 commonsourceibias.n417 commonsourceibias.n388 47.3584
R685 commonsourceibias.n457 commonsourceibias.n456 47.3584
R686 commonsourceibias.n341 commonsourceibias.n340 47.3584
R687 commonsourceibias.n301 commonsourceibias.n272 47.3584
R688 commonsourceibias.n104 commonsourceibias.n103 47.3584
R689 commonsourceibias.n64 commonsourceibias.n35 47.3584
R690 commonsourceibias.n226 commonsourceibias.n225 47.3584
R691 commonsourceibias.n186 commonsourceibias.n157 47.3584
R692 commonsourceibias.n896 commonsourceibias.n867 47.3584
R693 commonsourceibias.n939 commonsourceibias.n938 47.3584
R694 commonsourceibias.n780 commonsourceibias.n751 47.3584
R695 commonsourceibias.n823 commonsourceibias.n822 47.3584
R696 commonsourceibias.n550 commonsourceibias.n521 47.3584
R697 commonsourceibias.n593 commonsourceibias.n592 47.3584
R698 commonsourceibias.n708 commonsourceibias.n707 47.3584
R699 commonsourceibias.n666 commonsourceibias.n637 47.3584
R700 commonsourceibias.n403 commonsourceibias.n393 46.3896
R701 commonsourceibias.n471 commonsourceibias.n470 46.3896
R702 commonsourceibias.n355 commonsourceibias.n354 46.3896
R703 commonsourceibias.n287 commonsourceibias.n277 46.3896
R704 commonsourceibias.n118 commonsourceibias.n117 46.3896
R705 commonsourceibias.n50 commonsourceibias.n40 46.3896
R706 commonsourceibias.n240 commonsourceibias.n239 46.3896
R707 commonsourceibias.n172 commonsourceibias.n162 46.3896
R708 commonsourceibias.n881 commonsourceibias.n871 46.3896
R709 commonsourceibias.n954 commonsourceibias.n953 46.3896
R710 commonsourceibias.n765 commonsourceibias.n755 46.3896
R711 commonsourceibias.n838 commonsourceibias.n837 46.3896
R712 commonsourceibias.n535 commonsourceibias.n525 46.3896
R713 commonsourceibias.n608 commonsourceibias.n607 46.3896
R714 commonsourceibias.n723 commonsourceibias.n722 46.3896
R715 commonsourceibias.n651 commonsourceibias.n641 46.3896
R716 commonsourceibias.n398 commonsourceibias.n397 44.7059
R717 commonsourceibias.n876 commonsourceibias.n875 44.7059
R718 commonsourceibias.n760 commonsourceibias.n759 44.7059
R719 commonsourceibias.n530 commonsourceibias.n529 44.7059
R720 commonsourceibias.n646 commonsourceibias.n645 44.7059
R721 commonsourceibias.n282 commonsourceibias.n281 44.7059
R722 commonsourceibias.n45 commonsourceibias.n44 44.7059
R723 commonsourceibias.n167 commonsourceibias.n166 44.7059
R724 commonsourceibias.n407 commonsourceibias.n393 34.7644
R725 commonsourceibias.n470 commonsourceibias.n370 34.7644
R726 commonsourceibias.n354 commonsourceibias.n254 34.7644
R727 commonsourceibias.n291 commonsourceibias.n277 34.7644
R728 commonsourceibias.n117 commonsourceibias.n17 34.7644
R729 commonsourceibias.n54 commonsourceibias.n40 34.7644
R730 commonsourceibias.n239 commonsourceibias.n3 34.7644
R731 commonsourceibias.n176 commonsourceibias.n162 34.7644
R732 commonsourceibias.n885 commonsourceibias.n871 34.7644
R733 commonsourceibias.n953 commonsourceibias.n853 34.7644
R734 commonsourceibias.n769 commonsourceibias.n755 34.7644
R735 commonsourceibias.n837 commonsourceibias.n737 34.7644
R736 commonsourceibias.n539 commonsourceibias.n525 34.7644
R737 commonsourceibias.n607 commonsourceibias.n507 34.7644
R738 commonsourceibias.n722 commonsourceibias.n486 34.7644
R739 commonsourceibias.n655 commonsourceibias.n641 34.7644
R740 commonsourceibias.n421 commonsourceibias.n388 33.7956
R741 commonsourceibias.n456 commonsourceibias.n375 33.7956
R742 commonsourceibias.n340 commonsourceibias.n259 33.7956
R743 commonsourceibias.n305 commonsourceibias.n272 33.7956
R744 commonsourceibias.n103 commonsourceibias.n22 33.7956
R745 commonsourceibias.n68 commonsourceibias.n35 33.7956
R746 commonsourceibias.n225 commonsourceibias.n8 33.7956
R747 commonsourceibias.n190 commonsourceibias.n157 33.7956
R748 commonsourceibias.n900 commonsourceibias.n867 33.7956
R749 commonsourceibias.n938 commonsourceibias.n857 33.7956
R750 commonsourceibias.n784 commonsourceibias.n751 33.7956
R751 commonsourceibias.n822 commonsourceibias.n741 33.7956
R752 commonsourceibias.n554 commonsourceibias.n521 33.7956
R753 commonsourceibias.n592 commonsourceibias.n511 33.7956
R754 commonsourceibias.n707 commonsourceibias.n490 33.7956
R755 commonsourceibias.n670 commonsourceibias.n637 33.7956
R756 commonsourceibias.n435 commonsourceibias.n383 32.8269
R757 commonsourceibias.n442 commonsourceibias.n380 32.8269
R758 commonsourceibias.n326 commonsourceibias.n264 32.8269
R759 commonsourceibias.n319 commonsourceibias.n267 32.8269
R760 commonsourceibias.n89 commonsourceibias.n27 32.8269
R761 commonsourceibias.n82 commonsourceibias.n30 32.8269
R762 commonsourceibias.n211 commonsourceibias.n13 32.8269
R763 commonsourceibias.n203 commonsourceibias.n202 32.8269
R764 commonsourceibias.n915 commonsourceibias.n863 32.8269
R765 commonsourceibias.n923 commonsourceibias.n861 32.8269
R766 commonsourceibias.n799 commonsourceibias.n747 32.8269
R767 commonsourceibias.n807 commonsourceibias.n745 32.8269
R768 commonsourceibias.n569 commonsourceibias.n517 32.8269
R769 commonsourceibias.n577 commonsourceibias.n515 32.8269
R770 commonsourceibias.n692 commonsourceibias.n494 32.8269
R771 commonsourceibias.n683 commonsourceibias.n682 32.8269
R772 commonsourceibias.n428 commonsourceibias.n385 31.8581
R773 commonsourceibias.n449 commonsourceibias.n378 31.8581
R774 commonsourceibias.n333 commonsourceibias.n262 31.8581
R775 commonsourceibias.n312 commonsourceibias.n269 31.8581
R776 commonsourceibias.n96 commonsourceibias.n25 31.8581
R777 commonsourceibias.n75 commonsourceibias.n32 31.8581
R778 commonsourceibias.n218 commonsourceibias.n11 31.8581
R779 commonsourceibias.n197 commonsourceibias.n196 31.8581
R780 commonsourceibias.n908 commonsourceibias.n865 31.8581
R781 commonsourceibias.n930 commonsourceibias.n859 31.8581
R782 commonsourceibias.n792 commonsourceibias.n749 31.8581
R783 commonsourceibias.n814 commonsourceibias.n743 31.8581
R784 commonsourceibias.n562 commonsourceibias.n519 31.8581
R785 commonsourceibias.n584 commonsourceibias.n513 31.8581
R786 commonsourceibias.n699 commonsourceibias.n492 31.8581
R787 commonsourceibias.n677 commonsourceibias.n676 31.8581
R788 commonsourceibias.n414 commonsourceibias.n390 30.8893
R789 commonsourceibias.n463 commonsourceibias.n373 30.8893
R790 commonsourceibias.n347 commonsourceibias.n257 30.8893
R791 commonsourceibias.n298 commonsourceibias.n274 30.8893
R792 commonsourceibias.n110 commonsourceibias.n20 30.8893
R793 commonsourceibias.n61 commonsourceibias.n37 30.8893
R794 commonsourceibias.n232 commonsourceibias.n6 30.8893
R795 commonsourceibias.n183 commonsourceibias.n159 30.8893
R796 commonsourceibias.n893 commonsourceibias.n869 30.8893
R797 commonsourceibias.n945 commonsourceibias.n855 30.8893
R798 commonsourceibias.n777 commonsourceibias.n753 30.8893
R799 commonsourceibias.n829 commonsourceibias.n739 30.8893
R800 commonsourceibias.n547 commonsourceibias.n523 30.8893
R801 commonsourceibias.n599 commonsourceibias.n509 30.8893
R802 commonsourceibias.n714 commonsourceibias.n488 30.8893
R803 commonsourceibias.n663 commonsourceibias.n639 30.8893
R804 commonsourceibias.n400 commonsourceibias.n395 29.9206
R805 commonsourceibias.n477 commonsourceibias.n368 29.9206
R806 commonsourceibias.n361 commonsourceibias.n252 29.9206
R807 commonsourceibias.n284 commonsourceibias.n279 29.9206
R808 commonsourceibias.n124 commonsourceibias.n15 29.9206
R809 commonsourceibias.n47 commonsourceibias.n42 29.9206
R810 commonsourceibias.n246 commonsourceibias.n1 29.9206
R811 commonsourceibias.n169 commonsourceibias.n164 29.9206
R812 commonsourceibias.n878 commonsourceibias.n873 29.9206
R813 commonsourceibias.n960 commonsourceibias.n851 29.9206
R814 commonsourceibias.n762 commonsourceibias.n757 29.9206
R815 commonsourceibias.n844 commonsourceibias.n735 29.9206
R816 commonsourceibias.n532 commonsourceibias.n527 29.9206
R817 commonsourceibias.n614 commonsourceibias.n505 29.9206
R818 commonsourceibias.n729 commonsourceibias.n484 29.9206
R819 commonsourceibias.n648 commonsourceibias.n643 29.9206
R820 commonsourceibias.n479 commonsourceibias.n478 21.8872
R821 commonsourceibias.n363 commonsourceibias.n362 21.8872
R822 commonsourceibias.n126 commonsourceibias.n125 21.8872
R823 commonsourceibias.n248 commonsourceibias.n247 21.8872
R824 commonsourceibias.n962 commonsourceibias.n961 21.8872
R825 commonsourceibias.n846 commonsourceibias.n845 21.8872
R826 commonsourceibias.n616 commonsourceibias.n615 21.8872
R827 commonsourceibias.n731 commonsourceibias.n730 21.8872
R828 commonsourceibias.n410 commonsourceibias.n392 21.3954
R829 commonsourceibias.n465 commonsourceibias.n464 21.3954
R830 commonsourceibias.n349 commonsourceibias.n348 21.3954
R831 commonsourceibias.n294 commonsourceibias.n276 21.3954
R832 commonsourceibias.n112 commonsourceibias.n111 21.3954
R833 commonsourceibias.n57 commonsourceibias.n39 21.3954
R834 commonsourceibias.n234 commonsourceibias.n233 21.3954
R835 commonsourceibias.n179 commonsourceibias.n161 21.3954
R836 commonsourceibias.n889 commonsourceibias.n888 21.3954
R837 commonsourceibias.n947 commonsourceibias.n946 21.3954
R838 commonsourceibias.n773 commonsourceibias.n772 21.3954
R839 commonsourceibias.n831 commonsourceibias.n830 21.3954
R840 commonsourceibias.n543 commonsourceibias.n542 21.3954
R841 commonsourceibias.n601 commonsourceibias.n600 21.3954
R842 commonsourceibias.n716 commonsourceibias.n715 21.3954
R843 commonsourceibias.n659 commonsourceibias.n658 21.3954
R844 commonsourceibias.n424 commonsourceibias.n387 20.9036
R845 commonsourceibias.n451 commonsourceibias.n450 20.9036
R846 commonsourceibias.n335 commonsourceibias.n334 20.9036
R847 commonsourceibias.n308 commonsourceibias.n271 20.9036
R848 commonsourceibias.n98 commonsourceibias.n97 20.9036
R849 commonsourceibias.n71 commonsourceibias.n34 20.9036
R850 commonsourceibias.n220 commonsourceibias.n219 20.9036
R851 commonsourceibias.n193 commonsourceibias.n155 20.9036
R852 commonsourceibias.n904 commonsourceibias.n903 20.9036
R853 commonsourceibias.n932 commonsourceibias.n931 20.9036
R854 commonsourceibias.n788 commonsourceibias.n787 20.9036
R855 commonsourceibias.n816 commonsourceibias.n815 20.9036
R856 commonsourceibias.n558 commonsourceibias.n557 20.9036
R857 commonsourceibias.n586 commonsourceibias.n585 20.9036
R858 commonsourceibias.n701 commonsourceibias.n700 20.9036
R859 commonsourceibias.n673 commonsourceibias.n635 20.9036
R860 commonsourceibias.n437 commonsourceibias.n436 20.4117
R861 commonsourceibias.n438 commonsourceibias.n382 20.4117
R862 commonsourceibias.n322 commonsourceibias.n266 20.4117
R863 commonsourceibias.n321 commonsourceibias.n320 20.4117
R864 commonsourceibias.n85 commonsourceibias.n29 20.4117
R865 commonsourceibias.n84 commonsourceibias.n83 20.4117
R866 commonsourceibias.n207 commonsourceibias.n150 20.4117
R867 commonsourceibias.n206 commonsourceibias.n151 20.4117
R868 commonsourceibias.n917 commonsourceibias.n916 20.4117
R869 commonsourceibias.n919 commonsourceibias.n918 20.4117
R870 commonsourceibias.n801 commonsourceibias.n800 20.4117
R871 commonsourceibias.n803 commonsourceibias.n802 20.4117
R872 commonsourceibias.n571 commonsourceibias.n570 20.4117
R873 commonsourceibias.n573 commonsourceibias.n572 20.4117
R874 commonsourceibias.n688 commonsourceibias.n687 20.4117
R875 commonsourceibias.n686 commonsourceibias.n631 20.4117
R876 commonsourceibias.n423 commonsourceibias.n422 19.9199
R877 commonsourceibias.n452 commonsourceibias.n377 19.9199
R878 commonsourceibias.n336 commonsourceibias.n261 19.9199
R879 commonsourceibias.n307 commonsourceibias.n306 19.9199
R880 commonsourceibias.n99 commonsourceibias.n24 19.9199
R881 commonsourceibias.n70 commonsourceibias.n69 19.9199
R882 commonsourceibias.n221 commonsourceibias.n10 19.9199
R883 commonsourceibias.n192 commonsourceibias.n191 19.9199
R884 commonsourceibias.n902 commonsourceibias.n901 19.9199
R885 commonsourceibias.n934 commonsourceibias.n933 19.9199
R886 commonsourceibias.n786 commonsourceibias.n785 19.9199
R887 commonsourceibias.n818 commonsourceibias.n817 19.9199
R888 commonsourceibias.n556 commonsourceibias.n555 19.9199
R889 commonsourceibias.n588 commonsourceibias.n587 19.9199
R890 commonsourceibias.n703 commonsourceibias.n702 19.9199
R891 commonsourceibias.n672 commonsourceibias.n671 19.9199
R892 commonsourceibias.n409 commonsourceibias.n408 19.4281
R893 commonsourceibias.n466 commonsourceibias.n372 19.4281
R894 commonsourceibias.n350 commonsourceibias.n256 19.4281
R895 commonsourceibias.n293 commonsourceibias.n292 19.4281
R896 commonsourceibias.n113 commonsourceibias.n19 19.4281
R897 commonsourceibias.n56 commonsourceibias.n55 19.4281
R898 commonsourceibias.n235 commonsourceibias.n5 19.4281
R899 commonsourceibias.n178 commonsourceibias.n177 19.4281
R900 commonsourceibias.n887 commonsourceibias.n886 19.4281
R901 commonsourceibias.n949 commonsourceibias.n948 19.4281
R902 commonsourceibias.n771 commonsourceibias.n770 19.4281
R903 commonsourceibias.n833 commonsourceibias.n832 19.4281
R904 commonsourceibias.n541 commonsourceibias.n540 19.4281
R905 commonsourceibias.n603 commonsourceibias.n602 19.4281
R906 commonsourceibias.n718 commonsourceibias.n717 19.4281
R907 commonsourceibias.n657 commonsourceibias.n656 19.4281
R908 commonsourceibias.n402 commonsourceibias.n401 13.526
R909 commonsourceibias.n473 commonsourceibias.n472 13.526
R910 commonsourceibias.n357 commonsourceibias.n356 13.526
R911 commonsourceibias.n286 commonsourceibias.n285 13.526
R912 commonsourceibias.n120 commonsourceibias.n119 13.526
R913 commonsourceibias.n49 commonsourceibias.n48 13.526
R914 commonsourceibias.n242 commonsourceibias.n241 13.526
R915 commonsourceibias.n171 commonsourceibias.n170 13.526
R916 commonsourceibias.n880 commonsourceibias.n879 13.526
R917 commonsourceibias.n956 commonsourceibias.n955 13.526
R918 commonsourceibias.n764 commonsourceibias.n763 13.526
R919 commonsourceibias.n840 commonsourceibias.n839 13.526
R920 commonsourceibias.n534 commonsourceibias.n533 13.526
R921 commonsourceibias.n610 commonsourceibias.n609 13.526
R922 commonsourceibias.n725 commonsourceibias.n724 13.526
R923 commonsourceibias.n650 commonsourceibias.n649 13.526
R924 commonsourceibias.n130 commonsourceibias.n128 13.2322
R925 commonsourceibias.n620 commonsourceibias.n618 13.2322
R926 commonsourceibias.n416 commonsourceibias.n415 13.0342
R927 commonsourceibias.n459 commonsourceibias.n458 13.0342
R928 commonsourceibias.n343 commonsourceibias.n342 13.0342
R929 commonsourceibias.n300 commonsourceibias.n299 13.0342
R930 commonsourceibias.n106 commonsourceibias.n105 13.0342
R931 commonsourceibias.n63 commonsourceibias.n62 13.0342
R932 commonsourceibias.n228 commonsourceibias.n227 13.0342
R933 commonsourceibias.n185 commonsourceibias.n184 13.0342
R934 commonsourceibias.n895 commonsourceibias.n894 13.0342
R935 commonsourceibias.n941 commonsourceibias.n940 13.0342
R936 commonsourceibias.n779 commonsourceibias.n778 13.0342
R937 commonsourceibias.n825 commonsourceibias.n824 13.0342
R938 commonsourceibias.n549 commonsourceibias.n548 13.0342
R939 commonsourceibias.n595 commonsourceibias.n594 13.0342
R940 commonsourceibias.n710 commonsourceibias.n709 13.0342
R941 commonsourceibias.n665 commonsourceibias.n664 13.0342
R942 commonsourceibias.n430 commonsourceibias.n429 12.5423
R943 commonsourceibias.n445 commonsourceibias.n444 12.5423
R944 commonsourceibias.n329 commonsourceibias.n328 12.5423
R945 commonsourceibias.n314 commonsourceibias.n313 12.5423
R946 commonsourceibias.n92 commonsourceibias.n91 12.5423
R947 commonsourceibias.n77 commonsourceibias.n76 12.5423
R948 commonsourceibias.n214 commonsourceibias.n213 12.5423
R949 commonsourceibias.n198 commonsourceibias.n153 12.5423
R950 commonsourceibias.n910 commonsourceibias.n909 12.5423
R951 commonsourceibias.n926 commonsourceibias.n925 12.5423
R952 commonsourceibias.n794 commonsourceibias.n793 12.5423
R953 commonsourceibias.n810 commonsourceibias.n809 12.5423
R954 commonsourceibias.n564 commonsourceibias.n563 12.5423
R955 commonsourceibias.n580 commonsourceibias.n579 12.5423
R956 commonsourceibias.n695 commonsourceibias.n694 12.5423
R957 commonsourceibias.n678 commonsourceibias.n633 12.5423
R958 commonsourceibias.n431 commonsourceibias.n430 12.0505
R959 commonsourceibias.n444 commonsourceibias.n443 12.0505
R960 commonsourceibias.n328 commonsourceibias.n327 12.0505
R961 commonsourceibias.n315 commonsourceibias.n314 12.0505
R962 commonsourceibias.n91 commonsourceibias.n90 12.0505
R963 commonsourceibias.n78 commonsourceibias.n77 12.0505
R964 commonsourceibias.n213 commonsourceibias.n212 12.0505
R965 commonsourceibias.n201 commonsourceibias.n153 12.0505
R966 commonsourceibias.n911 commonsourceibias.n910 12.0505
R967 commonsourceibias.n925 commonsourceibias.n924 12.0505
R968 commonsourceibias.n795 commonsourceibias.n794 12.0505
R969 commonsourceibias.n809 commonsourceibias.n808 12.0505
R970 commonsourceibias.n565 commonsourceibias.n564 12.0505
R971 commonsourceibias.n579 commonsourceibias.n578 12.0505
R972 commonsourceibias.n694 commonsourceibias.n693 12.0505
R973 commonsourceibias.n681 commonsourceibias.n633 12.0505
R974 commonsourceibias.n417 commonsourceibias.n416 11.5587
R975 commonsourceibias.n458 commonsourceibias.n457 11.5587
R976 commonsourceibias.n342 commonsourceibias.n341 11.5587
R977 commonsourceibias.n301 commonsourceibias.n300 11.5587
R978 commonsourceibias.n105 commonsourceibias.n104 11.5587
R979 commonsourceibias.n64 commonsourceibias.n63 11.5587
R980 commonsourceibias.n227 commonsourceibias.n226 11.5587
R981 commonsourceibias.n186 commonsourceibias.n185 11.5587
R982 commonsourceibias.n896 commonsourceibias.n895 11.5587
R983 commonsourceibias.n940 commonsourceibias.n939 11.5587
R984 commonsourceibias.n780 commonsourceibias.n779 11.5587
R985 commonsourceibias.n824 commonsourceibias.n823 11.5587
R986 commonsourceibias.n550 commonsourceibias.n549 11.5587
R987 commonsourceibias.n594 commonsourceibias.n593 11.5587
R988 commonsourceibias.n709 commonsourceibias.n708 11.5587
R989 commonsourceibias.n666 commonsourceibias.n665 11.5587
R990 commonsourceibias.n403 commonsourceibias.n402 11.0668
R991 commonsourceibias.n472 commonsourceibias.n471 11.0668
R992 commonsourceibias.n356 commonsourceibias.n355 11.0668
R993 commonsourceibias.n287 commonsourceibias.n286 11.0668
R994 commonsourceibias.n119 commonsourceibias.n118 11.0668
R995 commonsourceibias.n50 commonsourceibias.n49 11.0668
R996 commonsourceibias.n241 commonsourceibias.n240 11.0668
R997 commonsourceibias.n172 commonsourceibias.n171 11.0668
R998 commonsourceibias.n881 commonsourceibias.n880 11.0668
R999 commonsourceibias.n955 commonsourceibias.n954 11.0668
R1000 commonsourceibias.n765 commonsourceibias.n764 11.0668
R1001 commonsourceibias.n839 commonsourceibias.n838 11.0668
R1002 commonsourceibias.n535 commonsourceibias.n534 11.0668
R1003 commonsourceibias.n609 commonsourceibias.n608 11.0668
R1004 commonsourceibias.n724 commonsourceibias.n723 11.0668
R1005 commonsourceibias.n651 commonsourceibias.n650 11.0668
R1006 commonsourceibias.n966 commonsourceibias.n482 10.122
R1007 commonsourceibias.n149 commonsourceibias.n148 9.50363
R1008 commonsourceibias.n630 commonsourceibias.n629 9.50363
R1009 commonsourceibias.n366 commonsourceibias.n250 8.76042
R1010 commonsourceibias.n849 commonsourceibias.n733 8.76042
R1011 commonsourceibias.n966 commonsourceibias.n965 8.46921
R1012 commonsourceibias.n408 commonsourceibias.n407 5.16479
R1013 commonsourceibias.n372 commonsourceibias.n370 5.16479
R1014 commonsourceibias.n256 commonsourceibias.n254 5.16479
R1015 commonsourceibias.n292 commonsourceibias.n291 5.16479
R1016 commonsourceibias.n19 commonsourceibias.n17 5.16479
R1017 commonsourceibias.n55 commonsourceibias.n54 5.16479
R1018 commonsourceibias.n5 commonsourceibias.n3 5.16479
R1019 commonsourceibias.n177 commonsourceibias.n176 5.16479
R1020 commonsourceibias.n886 commonsourceibias.n885 5.16479
R1021 commonsourceibias.n948 commonsourceibias.n853 5.16479
R1022 commonsourceibias.n770 commonsourceibias.n769 5.16479
R1023 commonsourceibias.n832 commonsourceibias.n737 5.16479
R1024 commonsourceibias.n540 commonsourceibias.n539 5.16479
R1025 commonsourceibias.n602 commonsourceibias.n507 5.16479
R1026 commonsourceibias.n717 commonsourceibias.n486 5.16479
R1027 commonsourceibias.n656 commonsourceibias.n655 5.16479
R1028 commonsourceibias.n482 commonsourceibias.n481 5.03125
R1029 commonsourceibias.n366 commonsourceibias.n365 5.03125
R1030 commonsourceibias.n965 commonsourceibias.n964 5.03125
R1031 commonsourceibias.n849 commonsourceibias.n848 5.03125
R1032 commonsourceibias.n422 commonsourceibias.n421 4.67295
R1033 commonsourceibias.n377 commonsourceibias.n375 4.67295
R1034 commonsourceibias.n261 commonsourceibias.n259 4.67295
R1035 commonsourceibias.n306 commonsourceibias.n305 4.67295
R1036 commonsourceibias.n24 commonsourceibias.n22 4.67295
R1037 commonsourceibias.n69 commonsourceibias.n68 4.67295
R1038 commonsourceibias.n10 commonsourceibias.n8 4.67295
R1039 commonsourceibias.n191 commonsourceibias.n190 4.67295
R1040 commonsourceibias.n901 commonsourceibias.n900 4.67295
R1041 commonsourceibias.n933 commonsourceibias.n857 4.67295
R1042 commonsourceibias.n785 commonsourceibias.n784 4.67295
R1043 commonsourceibias.n817 commonsourceibias.n741 4.67295
R1044 commonsourceibias.n555 commonsourceibias.n554 4.67295
R1045 commonsourceibias.n587 commonsourceibias.n511 4.67295
R1046 commonsourceibias.n702 commonsourceibias.n490 4.67295
R1047 commonsourceibias.n671 commonsourceibias.n670 4.67295
R1048 commonsourceibias commonsourceibias.n966 4.20978
R1049 commonsourceibias.n436 commonsourceibias.n435 4.18111
R1050 commonsourceibias.n382 commonsourceibias.n380 4.18111
R1051 commonsourceibias.n266 commonsourceibias.n264 4.18111
R1052 commonsourceibias.n320 commonsourceibias.n319 4.18111
R1053 commonsourceibias.n29 commonsourceibias.n27 4.18111
R1054 commonsourceibias.n83 commonsourceibias.n82 4.18111
R1055 commonsourceibias.n150 commonsourceibias.n13 4.18111
R1056 commonsourceibias.n203 commonsourceibias.n151 4.18111
R1057 commonsourceibias.n916 commonsourceibias.n915 4.18111
R1058 commonsourceibias.n918 commonsourceibias.n861 4.18111
R1059 commonsourceibias.n800 commonsourceibias.n799 4.18111
R1060 commonsourceibias.n802 commonsourceibias.n745 4.18111
R1061 commonsourceibias.n570 commonsourceibias.n569 4.18111
R1062 commonsourceibias.n572 commonsourceibias.n515 4.18111
R1063 commonsourceibias.n687 commonsourceibias.n494 4.18111
R1064 commonsourceibias.n683 commonsourceibias.n631 4.18111
R1065 commonsourceibias.n482 commonsourceibias.n366 3.72967
R1066 commonsourceibias.n965 commonsourceibias.n849 3.72967
R1067 commonsourceibias.n387 commonsourceibias.n385 3.68928
R1068 commonsourceibias.n450 commonsourceibias.n449 3.68928
R1069 commonsourceibias.n334 commonsourceibias.n333 3.68928
R1070 commonsourceibias.n271 commonsourceibias.n269 3.68928
R1071 commonsourceibias.n97 commonsourceibias.n96 3.68928
R1072 commonsourceibias.n34 commonsourceibias.n32 3.68928
R1073 commonsourceibias.n219 commonsourceibias.n218 3.68928
R1074 commonsourceibias.n196 commonsourceibias.n155 3.68928
R1075 commonsourceibias.n903 commonsourceibias.n865 3.68928
R1076 commonsourceibias.n931 commonsourceibias.n930 3.68928
R1077 commonsourceibias.n787 commonsourceibias.n749 3.68928
R1078 commonsourceibias.n815 commonsourceibias.n814 3.68928
R1079 commonsourceibias.n557 commonsourceibias.n519 3.68928
R1080 commonsourceibias.n585 commonsourceibias.n584 3.68928
R1081 commonsourceibias.n700 commonsourceibias.n699 3.68928
R1082 commonsourceibias.n676 commonsourceibias.n635 3.68928
R1083 commonsourceibias.n392 commonsourceibias.n390 3.19744
R1084 commonsourceibias.n464 commonsourceibias.n463 3.19744
R1085 commonsourceibias.n348 commonsourceibias.n347 3.19744
R1086 commonsourceibias.n276 commonsourceibias.n274 3.19744
R1087 commonsourceibias.n111 commonsourceibias.n110 3.19744
R1088 commonsourceibias.n39 commonsourceibias.n37 3.19744
R1089 commonsourceibias.n233 commonsourceibias.n232 3.19744
R1090 commonsourceibias.n161 commonsourceibias.n159 3.19744
R1091 commonsourceibias.n888 commonsourceibias.n869 3.19744
R1092 commonsourceibias.n946 commonsourceibias.n945 3.19744
R1093 commonsourceibias.n772 commonsourceibias.n753 3.19744
R1094 commonsourceibias.n830 commonsourceibias.n829 3.19744
R1095 commonsourceibias.n542 commonsourceibias.n523 3.19744
R1096 commonsourceibias.n600 commonsourceibias.n599 3.19744
R1097 commonsourceibias.n715 commonsourceibias.n714 3.19744
R1098 commonsourceibias.n658 commonsourceibias.n639 3.19744
R1099 commonsourceibias.n139 commonsourceibias.t19 2.82907
R1100 commonsourceibias.n139 commonsourceibias.t63 2.82907
R1101 commonsourceibias.n140 commonsourceibias.t23 2.82907
R1102 commonsourceibias.n140 commonsourceibias.t33 2.82907
R1103 commonsourceibias.n142 commonsourceibias.t11 2.82907
R1104 commonsourceibias.n142 commonsourceibias.t77 2.82907
R1105 commonsourceibias.n144 commonsourceibias.t7 2.82907
R1106 commonsourceibias.n144 commonsourceibias.t59 2.82907
R1107 commonsourceibias.n146 commonsourceibias.t39 2.82907
R1108 commonsourceibias.n146 commonsourceibias.t45 2.82907
R1109 commonsourceibias.n137 commonsourceibias.t55 2.82907
R1110 commonsourceibias.n137 commonsourceibias.t35 2.82907
R1111 commonsourceibias.n135 commonsourceibias.t43 2.82907
R1112 commonsourceibias.n135 commonsourceibias.t73 2.82907
R1113 commonsourceibias.n133 commonsourceibias.t1 2.82907
R1114 commonsourceibias.n133 commonsourceibias.t57 2.82907
R1115 commonsourceibias.n131 commonsourceibias.t67 2.82907
R1116 commonsourceibias.n131 commonsourceibias.t51 2.82907
R1117 commonsourceibias.n129 commonsourceibias.t53 2.82907
R1118 commonsourceibias.n129 commonsourceibias.t21 2.82907
R1119 commonsourceibias.n619 commonsourceibias.t3 2.82907
R1120 commonsourceibias.n619 commonsourceibias.t49 2.82907
R1121 commonsourceibias.n621 commonsourceibias.t47 2.82907
R1122 commonsourceibias.n621 commonsourceibias.t61 2.82907
R1123 commonsourceibias.n623 commonsourceibias.t27 2.82907
R1124 commonsourceibias.n623 commonsourceibias.t75 2.82907
R1125 commonsourceibias.n625 commonsourceibias.t41 2.82907
R1126 commonsourceibias.n625 commonsourceibias.t17 2.82907
R1127 commonsourceibias.n627 commonsourceibias.t9 2.82907
R1128 commonsourceibias.n627 commonsourceibias.t25 2.82907
R1129 commonsourceibias.n502 commonsourceibias.t13 2.82907
R1130 commonsourceibias.n502 commonsourceibias.t31 2.82907
R1131 commonsourceibias.n500 commonsourceibias.t29 2.82907
R1132 commonsourceibias.n500 commonsourceibias.t65 2.82907
R1133 commonsourceibias.n498 commonsourceibias.t37 2.82907
R1134 commonsourceibias.n498 commonsourceibias.t79 2.82907
R1135 commonsourceibias.n496 commonsourceibias.t69 2.82907
R1136 commonsourceibias.n496 commonsourceibias.t15 2.82907
R1137 commonsourceibias.n495 commonsourceibias.t5 2.82907
R1138 commonsourceibias.n495 commonsourceibias.t71 2.82907
R1139 commonsourceibias.n396 commonsourceibias.n395 2.7056
R1140 commonsourceibias.n478 commonsourceibias.n477 2.7056
R1141 commonsourceibias.n362 commonsourceibias.n361 2.7056
R1142 commonsourceibias.n280 commonsourceibias.n279 2.7056
R1143 commonsourceibias.n125 commonsourceibias.n124 2.7056
R1144 commonsourceibias.n43 commonsourceibias.n42 2.7056
R1145 commonsourceibias.n247 commonsourceibias.n246 2.7056
R1146 commonsourceibias.n165 commonsourceibias.n164 2.7056
R1147 commonsourceibias.n874 commonsourceibias.n873 2.7056
R1148 commonsourceibias.n961 commonsourceibias.n960 2.7056
R1149 commonsourceibias.n758 commonsourceibias.n757 2.7056
R1150 commonsourceibias.n845 commonsourceibias.n844 2.7056
R1151 commonsourceibias.n528 commonsourceibias.n527 2.7056
R1152 commonsourceibias.n615 commonsourceibias.n614 2.7056
R1153 commonsourceibias.n730 commonsourceibias.n729 2.7056
R1154 commonsourceibias.n644 commonsourceibias.n643 2.7056
R1155 commonsourceibias.n132 commonsourceibias.n130 0.573776
R1156 commonsourceibias.n134 commonsourceibias.n132 0.573776
R1157 commonsourceibias.n136 commonsourceibias.n134 0.573776
R1158 commonsourceibias.n138 commonsourceibias.n136 0.573776
R1159 commonsourceibias.n147 commonsourceibias.n145 0.573776
R1160 commonsourceibias.n145 commonsourceibias.n143 0.573776
R1161 commonsourceibias.n143 commonsourceibias.n141 0.573776
R1162 commonsourceibias.n499 commonsourceibias.n497 0.573776
R1163 commonsourceibias.n501 commonsourceibias.n499 0.573776
R1164 commonsourceibias.n503 commonsourceibias.n501 0.573776
R1165 commonsourceibias.n628 commonsourceibias.n626 0.573776
R1166 commonsourceibias.n626 commonsourceibias.n624 0.573776
R1167 commonsourceibias.n624 commonsourceibias.n622 0.573776
R1168 commonsourceibias.n622 commonsourceibias.n620 0.573776
R1169 commonsourceibias.n148 commonsourceibias.n138 0.287138
R1170 commonsourceibias.n148 commonsourceibias.n147 0.287138
R1171 commonsourceibias.n629 commonsourceibias.n503 0.287138
R1172 commonsourceibias.n629 commonsourceibias.n628 0.287138
R1173 commonsourceibias.n481 commonsourceibias.n367 0.285035
R1174 commonsourceibias.n365 commonsourceibias.n251 0.285035
R1175 commonsourceibias.n128 commonsourceibias.n14 0.285035
R1176 commonsourceibias.n250 commonsourceibias.n0 0.285035
R1177 commonsourceibias.n964 commonsourceibias.n850 0.285035
R1178 commonsourceibias.n848 commonsourceibias.n734 0.285035
R1179 commonsourceibias.n618 commonsourceibias.n504 0.285035
R1180 commonsourceibias.n733 commonsourceibias.n483 0.285035
R1181 commonsourceibias.n476 commonsourceibias.n367 0.189894
R1182 commonsourceibias.n476 commonsourceibias.n475 0.189894
R1183 commonsourceibias.n475 commonsourceibias.n474 0.189894
R1184 commonsourceibias.n474 commonsourceibias.n369 0.189894
R1185 commonsourceibias.n469 commonsourceibias.n369 0.189894
R1186 commonsourceibias.n469 commonsourceibias.n468 0.189894
R1187 commonsourceibias.n468 commonsourceibias.n467 0.189894
R1188 commonsourceibias.n467 commonsourceibias.n371 0.189894
R1189 commonsourceibias.n462 commonsourceibias.n371 0.189894
R1190 commonsourceibias.n462 commonsourceibias.n461 0.189894
R1191 commonsourceibias.n461 commonsourceibias.n460 0.189894
R1192 commonsourceibias.n460 commonsourceibias.n374 0.189894
R1193 commonsourceibias.n455 commonsourceibias.n374 0.189894
R1194 commonsourceibias.n455 commonsourceibias.n454 0.189894
R1195 commonsourceibias.n454 commonsourceibias.n453 0.189894
R1196 commonsourceibias.n453 commonsourceibias.n376 0.189894
R1197 commonsourceibias.n448 commonsourceibias.n376 0.189894
R1198 commonsourceibias.n448 commonsourceibias.n447 0.189894
R1199 commonsourceibias.n447 commonsourceibias.n446 0.189894
R1200 commonsourceibias.n446 commonsourceibias.n379 0.189894
R1201 commonsourceibias.n441 commonsourceibias.n379 0.189894
R1202 commonsourceibias.n441 commonsourceibias.n440 0.189894
R1203 commonsourceibias.n440 commonsourceibias.n439 0.189894
R1204 commonsourceibias.n439 commonsourceibias.n381 0.189894
R1205 commonsourceibias.n434 commonsourceibias.n381 0.189894
R1206 commonsourceibias.n434 commonsourceibias.n433 0.189894
R1207 commonsourceibias.n433 commonsourceibias.n432 0.189894
R1208 commonsourceibias.n432 commonsourceibias.n384 0.189894
R1209 commonsourceibias.n427 commonsourceibias.n384 0.189894
R1210 commonsourceibias.n427 commonsourceibias.n426 0.189894
R1211 commonsourceibias.n426 commonsourceibias.n425 0.189894
R1212 commonsourceibias.n425 commonsourceibias.n386 0.189894
R1213 commonsourceibias.n420 commonsourceibias.n386 0.189894
R1214 commonsourceibias.n420 commonsourceibias.n419 0.189894
R1215 commonsourceibias.n419 commonsourceibias.n418 0.189894
R1216 commonsourceibias.n418 commonsourceibias.n389 0.189894
R1217 commonsourceibias.n413 commonsourceibias.n389 0.189894
R1218 commonsourceibias.n413 commonsourceibias.n412 0.189894
R1219 commonsourceibias.n412 commonsourceibias.n411 0.189894
R1220 commonsourceibias.n411 commonsourceibias.n391 0.189894
R1221 commonsourceibias.n406 commonsourceibias.n391 0.189894
R1222 commonsourceibias.n406 commonsourceibias.n405 0.189894
R1223 commonsourceibias.n405 commonsourceibias.n404 0.189894
R1224 commonsourceibias.n404 commonsourceibias.n394 0.189894
R1225 commonsourceibias.n399 commonsourceibias.n394 0.189894
R1226 commonsourceibias.n399 commonsourceibias.n398 0.189894
R1227 commonsourceibias.n360 commonsourceibias.n251 0.189894
R1228 commonsourceibias.n360 commonsourceibias.n359 0.189894
R1229 commonsourceibias.n359 commonsourceibias.n358 0.189894
R1230 commonsourceibias.n358 commonsourceibias.n253 0.189894
R1231 commonsourceibias.n353 commonsourceibias.n253 0.189894
R1232 commonsourceibias.n353 commonsourceibias.n352 0.189894
R1233 commonsourceibias.n352 commonsourceibias.n351 0.189894
R1234 commonsourceibias.n351 commonsourceibias.n255 0.189894
R1235 commonsourceibias.n346 commonsourceibias.n255 0.189894
R1236 commonsourceibias.n346 commonsourceibias.n345 0.189894
R1237 commonsourceibias.n345 commonsourceibias.n344 0.189894
R1238 commonsourceibias.n344 commonsourceibias.n258 0.189894
R1239 commonsourceibias.n339 commonsourceibias.n258 0.189894
R1240 commonsourceibias.n339 commonsourceibias.n338 0.189894
R1241 commonsourceibias.n338 commonsourceibias.n337 0.189894
R1242 commonsourceibias.n337 commonsourceibias.n260 0.189894
R1243 commonsourceibias.n332 commonsourceibias.n260 0.189894
R1244 commonsourceibias.n332 commonsourceibias.n331 0.189894
R1245 commonsourceibias.n331 commonsourceibias.n330 0.189894
R1246 commonsourceibias.n330 commonsourceibias.n263 0.189894
R1247 commonsourceibias.n325 commonsourceibias.n263 0.189894
R1248 commonsourceibias.n325 commonsourceibias.n324 0.189894
R1249 commonsourceibias.n324 commonsourceibias.n323 0.189894
R1250 commonsourceibias.n323 commonsourceibias.n265 0.189894
R1251 commonsourceibias.n318 commonsourceibias.n265 0.189894
R1252 commonsourceibias.n318 commonsourceibias.n317 0.189894
R1253 commonsourceibias.n317 commonsourceibias.n316 0.189894
R1254 commonsourceibias.n316 commonsourceibias.n268 0.189894
R1255 commonsourceibias.n311 commonsourceibias.n268 0.189894
R1256 commonsourceibias.n311 commonsourceibias.n310 0.189894
R1257 commonsourceibias.n310 commonsourceibias.n309 0.189894
R1258 commonsourceibias.n309 commonsourceibias.n270 0.189894
R1259 commonsourceibias.n304 commonsourceibias.n270 0.189894
R1260 commonsourceibias.n304 commonsourceibias.n303 0.189894
R1261 commonsourceibias.n303 commonsourceibias.n302 0.189894
R1262 commonsourceibias.n302 commonsourceibias.n273 0.189894
R1263 commonsourceibias.n297 commonsourceibias.n273 0.189894
R1264 commonsourceibias.n297 commonsourceibias.n296 0.189894
R1265 commonsourceibias.n296 commonsourceibias.n295 0.189894
R1266 commonsourceibias.n295 commonsourceibias.n275 0.189894
R1267 commonsourceibias.n290 commonsourceibias.n275 0.189894
R1268 commonsourceibias.n290 commonsourceibias.n289 0.189894
R1269 commonsourceibias.n289 commonsourceibias.n288 0.189894
R1270 commonsourceibias.n288 commonsourceibias.n278 0.189894
R1271 commonsourceibias.n283 commonsourceibias.n278 0.189894
R1272 commonsourceibias.n283 commonsourceibias.n282 0.189894
R1273 commonsourceibias.n123 commonsourceibias.n14 0.189894
R1274 commonsourceibias.n123 commonsourceibias.n122 0.189894
R1275 commonsourceibias.n122 commonsourceibias.n121 0.189894
R1276 commonsourceibias.n121 commonsourceibias.n16 0.189894
R1277 commonsourceibias.n116 commonsourceibias.n16 0.189894
R1278 commonsourceibias.n116 commonsourceibias.n115 0.189894
R1279 commonsourceibias.n115 commonsourceibias.n114 0.189894
R1280 commonsourceibias.n114 commonsourceibias.n18 0.189894
R1281 commonsourceibias.n109 commonsourceibias.n18 0.189894
R1282 commonsourceibias.n109 commonsourceibias.n108 0.189894
R1283 commonsourceibias.n108 commonsourceibias.n107 0.189894
R1284 commonsourceibias.n107 commonsourceibias.n21 0.189894
R1285 commonsourceibias.n102 commonsourceibias.n21 0.189894
R1286 commonsourceibias.n102 commonsourceibias.n101 0.189894
R1287 commonsourceibias.n101 commonsourceibias.n100 0.189894
R1288 commonsourceibias.n100 commonsourceibias.n23 0.189894
R1289 commonsourceibias.n95 commonsourceibias.n23 0.189894
R1290 commonsourceibias.n95 commonsourceibias.n94 0.189894
R1291 commonsourceibias.n94 commonsourceibias.n93 0.189894
R1292 commonsourceibias.n93 commonsourceibias.n26 0.189894
R1293 commonsourceibias.n88 commonsourceibias.n26 0.189894
R1294 commonsourceibias.n88 commonsourceibias.n87 0.189894
R1295 commonsourceibias.n87 commonsourceibias.n86 0.189894
R1296 commonsourceibias.n86 commonsourceibias.n28 0.189894
R1297 commonsourceibias.n81 commonsourceibias.n28 0.189894
R1298 commonsourceibias.n81 commonsourceibias.n80 0.189894
R1299 commonsourceibias.n80 commonsourceibias.n79 0.189894
R1300 commonsourceibias.n79 commonsourceibias.n31 0.189894
R1301 commonsourceibias.n74 commonsourceibias.n31 0.189894
R1302 commonsourceibias.n74 commonsourceibias.n73 0.189894
R1303 commonsourceibias.n73 commonsourceibias.n72 0.189894
R1304 commonsourceibias.n72 commonsourceibias.n33 0.189894
R1305 commonsourceibias.n67 commonsourceibias.n33 0.189894
R1306 commonsourceibias.n67 commonsourceibias.n66 0.189894
R1307 commonsourceibias.n66 commonsourceibias.n65 0.189894
R1308 commonsourceibias.n65 commonsourceibias.n36 0.189894
R1309 commonsourceibias.n60 commonsourceibias.n36 0.189894
R1310 commonsourceibias.n60 commonsourceibias.n59 0.189894
R1311 commonsourceibias.n59 commonsourceibias.n58 0.189894
R1312 commonsourceibias.n58 commonsourceibias.n38 0.189894
R1313 commonsourceibias.n53 commonsourceibias.n38 0.189894
R1314 commonsourceibias.n53 commonsourceibias.n52 0.189894
R1315 commonsourceibias.n52 commonsourceibias.n51 0.189894
R1316 commonsourceibias.n51 commonsourceibias.n41 0.189894
R1317 commonsourceibias.n46 commonsourceibias.n41 0.189894
R1318 commonsourceibias.n46 commonsourceibias.n45 0.189894
R1319 commonsourceibias.n205 commonsourceibias.n204 0.189894
R1320 commonsourceibias.n204 commonsourceibias.n152 0.189894
R1321 commonsourceibias.n200 commonsourceibias.n152 0.189894
R1322 commonsourceibias.n200 commonsourceibias.n199 0.189894
R1323 commonsourceibias.n199 commonsourceibias.n154 0.189894
R1324 commonsourceibias.n195 commonsourceibias.n154 0.189894
R1325 commonsourceibias.n195 commonsourceibias.n194 0.189894
R1326 commonsourceibias.n194 commonsourceibias.n156 0.189894
R1327 commonsourceibias.n189 commonsourceibias.n156 0.189894
R1328 commonsourceibias.n189 commonsourceibias.n188 0.189894
R1329 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1330 commonsourceibias.n187 commonsourceibias.n158 0.189894
R1331 commonsourceibias.n182 commonsourceibias.n158 0.189894
R1332 commonsourceibias.n182 commonsourceibias.n181 0.189894
R1333 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1334 commonsourceibias.n180 commonsourceibias.n160 0.189894
R1335 commonsourceibias.n175 commonsourceibias.n160 0.189894
R1336 commonsourceibias.n175 commonsourceibias.n174 0.189894
R1337 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1338 commonsourceibias.n173 commonsourceibias.n163 0.189894
R1339 commonsourceibias.n168 commonsourceibias.n163 0.189894
R1340 commonsourceibias.n168 commonsourceibias.n167 0.189894
R1341 commonsourceibias.n245 commonsourceibias.n0 0.189894
R1342 commonsourceibias.n245 commonsourceibias.n244 0.189894
R1343 commonsourceibias.n244 commonsourceibias.n243 0.189894
R1344 commonsourceibias.n243 commonsourceibias.n2 0.189894
R1345 commonsourceibias.n238 commonsourceibias.n2 0.189894
R1346 commonsourceibias.n238 commonsourceibias.n237 0.189894
R1347 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1348 commonsourceibias.n236 commonsourceibias.n4 0.189894
R1349 commonsourceibias.n231 commonsourceibias.n4 0.189894
R1350 commonsourceibias.n231 commonsourceibias.n230 0.189894
R1351 commonsourceibias.n230 commonsourceibias.n229 0.189894
R1352 commonsourceibias.n229 commonsourceibias.n7 0.189894
R1353 commonsourceibias.n224 commonsourceibias.n7 0.189894
R1354 commonsourceibias.n224 commonsourceibias.n223 0.189894
R1355 commonsourceibias.n223 commonsourceibias.n222 0.189894
R1356 commonsourceibias.n222 commonsourceibias.n9 0.189894
R1357 commonsourceibias.n217 commonsourceibias.n9 0.189894
R1358 commonsourceibias.n217 commonsourceibias.n216 0.189894
R1359 commonsourceibias.n216 commonsourceibias.n215 0.189894
R1360 commonsourceibias.n215 commonsourceibias.n12 0.189894
R1361 commonsourceibias.n210 commonsourceibias.n12 0.189894
R1362 commonsourceibias.n210 commonsourceibias.n209 0.189894
R1363 commonsourceibias.n209 commonsourceibias.n208 0.189894
R1364 commonsourceibias.n877 commonsourceibias.n876 0.189894
R1365 commonsourceibias.n877 commonsourceibias.n872 0.189894
R1366 commonsourceibias.n882 commonsourceibias.n872 0.189894
R1367 commonsourceibias.n883 commonsourceibias.n882 0.189894
R1368 commonsourceibias.n884 commonsourceibias.n883 0.189894
R1369 commonsourceibias.n884 commonsourceibias.n870 0.189894
R1370 commonsourceibias.n890 commonsourceibias.n870 0.189894
R1371 commonsourceibias.n891 commonsourceibias.n890 0.189894
R1372 commonsourceibias.n892 commonsourceibias.n891 0.189894
R1373 commonsourceibias.n892 commonsourceibias.n868 0.189894
R1374 commonsourceibias.n897 commonsourceibias.n868 0.189894
R1375 commonsourceibias.n898 commonsourceibias.n897 0.189894
R1376 commonsourceibias.n899 commonsourceibias.n898 0.189894
R1377 commonsourceibias.n899 commonsourceibias.n866 0.189894
R1378 commonsourceibias.n905 commonsourceibias.n866 0.189894
R1379 commonsourceibias.n906 commonsourceibias.n905 0.189894
R1380 commonsourceibias.n907 commonsourceibias.n906 0.189894
R1381 commonsourceibias.n907 commonsourceibias.n864 0.189894
R1382 commonsourceibias.n912 commonsourceibias.n864 0.189894
R1383 commonsourceibias.n913 commonsourceibias.n912 0.189894
R1384 commonsourceibias.n914 commonsourceibias.n913 0.189894
R1385 commonsourceibias.n914 commonsourceibias.n862 0.189894
R1386 commonsourceibias.n920 commonsourceibias.n862 0.189894
R1387 commonsourceibias.n921 commonsourceibias.n920 0.189894
R1388 commonsourceibias.n922 commonsourceibias.n921 0.189894
R1389 commonsourceibias.n922 commonsourceibias.n860 0.189894
R1390 commonsourceibias.n927 commonsourceibias.n860 0.189894
R1391 commonsourceibias.n928 commonsourceibias.n927 0.189894
R1392 commonsourceibias.n929 commonsourceibias.n928 0.189894
R1393 commonsourceibias.n929 commonsourceibias.n858 0.189894
R1394 commonsourceibias.n935 commonsourceibias.n858 0.189894
R1395 commonsourceibias.n936 commonsourceibias.n935 0.189894
R1396 commonsourceibias.n937 commonsourceibias.n936 0.189894
R1397 commonsourceibias.n937 commonsourceibias.n856 0.189894
R1398 commonsourceibias.n942 commonsourceibias.n856 0.189894
R1399 commonsourceibias.n943 commonsourceibias.n942 0.189894
R1400 commonsourceibias.n944 commonsourceibias.n943 0.189894
R1401 commonsourceibias.n944 commonsourceibias.n854 0.189894
R1402 commonsourceibias.n950 commonsourceibias.n854 0.189894
R1403 commonsourceibias.n951 commonsourceibias.n950 0.189894
R1404 commonsourceibias.n952 commonsourceibias.n951 0.189894
R1405 commonsourceibias.n952 commonsourceibias.n852 0.189894
R1406 commonsourceibias.n957 commonsourceibias.n852 0.189894
R1407 commonsourceibias.n958 commonsourceibias.n957 0.189894
R1408 commonsourceibias.n959 commonsourceibias.n958 0.189894
R1409 commonsourceibias.n959 commonsourceibias.n850 0.189894
R1410 commonsourceibias.n761 commonsourceibias.n760 0.189894
R1411 commonsourceibias.n761 commonsourceibias.n756 0.189894
R1412 commonsourceibias.n766 commonsourceibias.n756 0.189894
R1413 commonsourceibias.n767 commonsourceibias.n766 0.189894
R1414 commonsourceibias.n768 commonsourceibias.n767 0.189894
R1415 commonsourceibias.n768 commonsourceibias.n754 0.189894
R1416 commonsourceibias.n774 commonsourceibias.n754 0.189894
R1417 commonsourceibias.n775 commonsourceibias.n774 0.189894
R1418 commonsourceibias.n776 commonsourceibias.n775 0.189894
R1419 commonsourceibias.n776 commonsourceibias.n752 0.189894
R1420 commonsourceibias.n781 commonsourceibias.n752 0.189894
R1421 commonsourceibias.n782 commonsourceibias.n781 0.189894
R1422 commonsourceibias.n783 commonsourceibias.n782 0.189894
R1423 commonsourceibias.n783 commonsourceibias.n750 0.189894
R1424 commonsourceibias.n789 commonsourceibias.n750 0.189894
R1425 commonsourceibias.n790 commonsourceibias.n789 0.189894
R1426 commonsourceibias.n791 commonsourceibias.n790 0.189894
R1427 commonsourceibias.n791 commonsourceibias.n748 0.189894
R1428 commonsourceibias.n796 commonsourceibias.n748 0.189894
R1429 commonsourceibias.n797 commonsourceibias.n796 0.189894
R1430 commonsourceibias.n798 commonsourceibias.n797 0.189894
R1431 commonsourceibias.n798 commonsourceibias.n746 0.189894
R1432 commonsourceibias.n804 commonsourceibias.n746 0.189894
R1433 commonsourceibias.n805 commonsourceibias.n804 0.189894
R1434 commonsourceibias.n806 commonsourceibias.n805 0.189894
R1435 commonsourceibias.n806 commonsourceibias.n744 0.189894
R1436 commonsourceibias.n811 commonsourceibias.n744 0.189894
R1437 commonsourceibias.n812 commonsourceibias.n811 0.189894
R1438 commonsourceibias.n813 commonsourceibias.n812 0.189894
R1439 commonsourceibias.n813 commonsourceibias.n742 0.189894
R1440 commonsourceibias.n819 commonsourceibias.n742 0.189894
R1441 commonsourceibias.n820 commonsourceibias.n819 0.189894
R1442 commonsourceibias.n821 commonsourceibias.n820 0.189894
R1443 commonsourceibias.n821 commonsourceibias.n740 0.189894
R1444 commonsourceibias.n826 commonsourceibias.n740 0.189894
R1445 commonsourceibias.n827 commonsourceibias.n826 0.189894
R1446 commonsourceibias.n828 commonsourceibias.n827 0.189894
R1447 commonsourceibias.n828 commonsourceibias.n738 0.189894
R1448 commonsourceibias.n834 commonsourceibias.n738 0.189894
R1449 commonsourceibias.n835 commonsourceibias.n834 0.189894
R1450 commonsourceibias.n836 commonsourceibias.n835 0.189894
R1451 commonsourceibias.n836 commonsourceibias.n736 0.189894
R1452 commonsourceibias.n841 commonsourceibias.n736 0.189894
R1453 commonsourceibias.n842 commonsourceibias.n841 0.189894
R1454 commonsourceibias.n843 commonsourceibias.n842 0.189894
R1455 commonsourceibias.n843 commonsourceibias.n734 0.189894
R1456 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1457 commonsourceibias.n531 commonsourceibias.n526 0.189894
R1458 commonsourceibias.n536 commonsourceibias.n526 0.189894
R1459 commonsourceibias.n537 commonsourceibias.n536 0.189894
R1460 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1461 commonsourceibias.n538 commonsourceibias.n524 0.189894
R1462 commonsourceibias.n544 commonsourceibias.n524 0.189894
R1463 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1464 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1465 commonsourceibias.n546 commonsourceibias.n522 0.189894
R1466 commonsourceibias.n551 commonsourceibias.n522 0.189894
R1467 commonsourceibias.n552 commonsourceibias.n551 0.189894
R1468 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1469 commonsourceibias.n553 commonsourceibias.n520 0.189894
R1470 commonsourceibias.n559 commonsourceibias.n520 0.189894
R1471 commonsourceibias.n560 commonsourceibias.n559 0.189894
R1472 commonsourceibias.n561 commonsourceibias.n560 0.189894
R1473 commonsourceibias.n561 commonsourceibias.n518 0.189894
R1474 commonsourceibias.n566 commonsourceibias.n518 0.189894
R1475 commonsourceibias.n567 commonsourceibias.n566 0.189894
R1476 commonsourceibias.n568 commonsourceibias.n567 0.189894
R1477 commonsourceibias.n568 commonsourceibias.n516 0.189894
R1478 commonsourceibias.n574 commonsourceibias.n516 0.189894
R1479 commonsourceibias.n575 commonsourceibias.n574 0.189894
R1480 commonsourceibias.n576 commonsourceibias.n575 0.189894
R1481 commonsourceibias.n576 commonsourceibias.n514 0.189894
R1482 commonsourceibias.n581 commonsourceibias.n514 0.189894
R1483 commonsourceibias.n582 commonsourceibias.n581 0.189894
R1484 commonsourceibias.n583 commonsourceibias.n582 0.189894
R1485 commonsourceibias.n583 commonsourceibias.n512 0.189894
R1486 commonsourceibias.n589 commonsourceibias.n512 0.189894
R1487 commonsourceibias.n590 commonsourceibias.n589 0.189894
R1488 commonsourceibias.n591 commonsourceibias.n590 0.189894
R1489 commonsourceibias.n591 commonsourceibias.n510 0.189894
R1490 commonsourceibias.n596 commonsourceibias.n510 0.189894
R1491 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1492 commonsourceibias.n598 commonsourceibias.n597 0.189894
R1493 commonsourceibias.n598 commonsourceibias.n508 0.189894
R1494 commonsourceibias.n604 commonsourceibias.n508 0.189894
R1495 commonsourceibias.n605 commonsourceibias.n604 0.189894
R1496 commonsourceibias.n606 commonsourceibias.n605 0.189894
R1497 commonsourceibias.n606 commonsourceibias.n506 0.189894
R1498 commonsourceibias.n611 commonsourceibias.n506 0.189894
R1499 commonsourceibias.n612 commonsourceibias.n611 0.189894
R1500 commonsourceibias.n613 commonsourceibias.n612 0.189894
R1501 commonsourceibias.n613 commonsourceibias.n504 0.189894
R1502 commonsourceibias.n647 commonsourceibias.n646 0.189894
R1503 commonsourceibias.n647 commonsourceibias.n642 0.189894
R1504 commonsourceibias.n652 commonsourceibias.n642 0.189894
R1505 commonsourceibias.n653 commonsourceibias.n652 0.189894
R1506 commonsourceibias.n654 commonsourceibias.n653 0.189894
R1507 commonsourceibias.n654 commonsourceibias.n640 0.189894
R1508 commonsourceibias.n660 commonsourceibias.n640 0.189894
R1509 commonsourceibias.n661 commonsourceibias.n660 0.189894
R1510 commonsourceibias.n662 commonsourceibias.n661 0.189894
R1511 commonsourceibias.n662 commonsourceibias.n638 0.189894
R1512 commonsourceibias.n667 commonsourceibias.n638 0.189894
R1513 commonsourceibias.n668 commonsourceibias.n667 0.189894
R1514 commonsourceibias.n669 commonsourceibias.n668 0.189894
R1515 commonsourceibias.n669 commonsourceibias.n636 0.189894
R1516 commonsourceibias.n674 commonsourceibias.n636 0.189894
R1517 commonsourceibias.n675 commonsourceibias.n674 0.189894
R1518 commonsourceibias.n675 commonsourceibias.n634 0.189894
R1519 commonsourceibias.n679 commonsourceibias.n634 0.189894
R1520 commonsourceibias.n680 commonsourceibias.n679 0.189894
R1521 commonsourceibias.n680 commonsourceibias.n632 0.189894
R1522 commonsourceibias.n684 commonsourceibias.n632 0.189894
R1523 commonsourceibias.n685 commonsourceibias.n684 0.189894
R1524 commonsourceibias.n690 commonsourceibias.n689 0.189894
R1525 commonsourceibias.n691 commonsourceibias.n690 0.189894
R1526 commonsourceibias.n691 commonsourceibias.n493 0.189894
R1527 commonsourceibias.n696 commonsourceibias.n493 0.189894
R1528 commonsourceibias.n697 commonsourceibias.n696 0.189894
R1529 commonsourceibias.n698 commonsourceibias.n697 0.189894
R1530 commonsourceibias.n698 commonsourceibias.n491 0.189894
R1531 commonsourceibias.n704 commonsourceibias.n491 0.189894
R1532 commonsourceibias.n705 commonsourceibias.n704 0.189894
R1533 commonsourceibias.n706 commonsourceibias.n705 0.189894
R1534 commonsourceibias.n706 commonsourceibias.n489 0.189894
R1535 commonsourceibias.n711 commonsourceibias.n489 0.189894
R1536 commonsourceibias.n712 commonsourceibias.n711 0.189894
R1537 commonsourceibias.n713 commonsourceibias.n712 0.189894
R1538 commonsourceibias.n713 commonsourceibias.n487 0.189894
R1539 commonsourceibias.n719 commonsourceibias.n487 0.189894
R1540 commonsourceibias.n720 commonsourceibias.n719 0.189894
R1541 commonsourceibias.n721 commonsourceibias.n720 0.189894
R1542 commonsourceibias.n721 commonsourceibias.n485 0.189894
R1543 commonsourceibias.n726 commonsourceibias.n485 0.189894
R1544 commonsourceibias.n727 commonsourceibias.n726 0.189894
R1545 commonsourceibias.n728 commonsourceibias.n727 0.189894
R1546 commonsourceibias.n728 commonsourceibias.n483 0.189894
R1547 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R1548 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R1549 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R1550 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R1551 gnd.n2773 gnd.n2772 1148.88
R1552 gnd.n4727 gnd.n4726 939.716
R1553 gnd.n5836 gnd.n1477 771.183
R1554 gnd.n6860 gnd.n766 771.183
R1555 gnd.n5840 gnd.n1459 771.183
R1556 gnd.n6862 gnd.n762 771.183
R1557 gnd.n4634 gnd.n1820 766.379
R1558 gnd.n4637 gnd.n4636 766.379
R1559 gnd.n3875 gnd.n3778 766.379
R1560 gnd.n3871 gnd.n3776 766.379
R1561 gnd.n4725 gnd.n1842 756.769
R1562 gnd.n4628 gnd.n4627 756.769
R1563 gnd.n3968 gnd.n3685 756.769
R1564 gnd.n3966 gnd.n3688 756.769
R1565 gnd.n3109 gnd.n2098 756.769
R1566 gnd.n2771 gnd.n2431 756.769
R1567 gnd.n2601 gnd.n357 756.769
R1568 gnd.n1974 gnd.n1973 756.769
R1569 gnd.n251 gnd.n241 751.963
R1570 gnd.n7449 gnd.n7448 751.963
R1571 gnd.n627 gnd.n571 751.963
R1572 gnd.n7067 gnd.n573 751.963
R1573 gnd.n5700 gnd.n5699 751.963
R1574 gnd.n5766 gnd.n1454 751.963
R1575 gnd.n4783 gnd.n4729 751.963
R1576 gnd.n5042 gnd.n4731 751.963
R1577 gnd.n7661 gnd.n245 696.707
R1578 gnd.n7537 gnd.n7536 696.707
R1579 gnd.n691 gnd.n570 696.707
R1580 gnd.n7069 gnd.n568 696.707
R1581 gnd.n5959 gnd.n1431 696.707
R1582 gnd.n5974 gnd.n1419 696.707
R1583 gnd.n5030 gnd.n4728 696.707
R1584 gnd.n5044 gnd.n1818 696.707
R1585 gnd.n7349 gnd.n357 589.749
R1586 gnd.n1973 gnd.n1972 589.749
R1587 gnd.n2098 gnd.n2097 585
R1588 gnd.n3111 gnd.n2098 585
R1589 gnd.n3114 gnd.n3113 585
R1590 gnd.n3113 gnd.n3112 585
R1591 gnd.n2095 gnd.n2094 585
R1592 gnd.n2094 gnd.n2093 585
R1593 gnd.n3119 gnd.n3118 585
R1594 gnd.n3120 gnd.n3119 585
R1595 gnd.n2092 gnd.n2091 585
R1596 gnd.n3121 gnd.n2092 585
R1597 gnd.n3124 gnd.n3123 585
R1598 gnd.n3123 gnd.n3122 585
R1599 gnd.n2089 gnd.n2088 585
R1600 gnd.n2088 gnd.n2087 585
R1601 gnd.n3129 gnd.n3128 585
R1602 gnd.n3130 gnd.n3129 585
R1603 gnd.n2086 gnd.n2085 585
R1604 gnd.n3131 gnd.n2086 585
R1605 gnd.n3134 gnd.n3133 585
R1606 gnd.n3133 gnd.n3132 585
R1607 gnd.n2083 gnd.n2082 585
R1608 gnd.n2082 gnd.n2081 585
R1609 gnd.n3139 gnd.n3138 585
R1610 gnd.n3140 gnd.n3139 585
R1611 gnd.n2080 gnd.n2079 585
R1612 gnd.n3141 gnd.n2080 585
R1613 gnd.n3144 gnd.n3143 585
R1614 gnd.n3143 gnd.n3142 585
R1615 gnd.n2077 gnd.n2076 585
R1616 gnd.n2076 gnd.n2075 585
R1617 gnd.n3149 gnd.n3148 585
R1618 gnd.n3150 gnd.n3149 585
R1619 gnd.n2074 gnd.n2073 585
R1620 gnd.n3151 gnd.n2074 585
R1621 gnd.n3154 gnd.n3153 585
R1622 gnd.n3153 gnd.n3152 585
R1623 gnd.n2071 gnd.n2070 585
R1624 gnd.n2070 gnd.n2069 585
R1625 gnd.n3159 gnd.n3158 585
R1626 gnd.n3160 gnd.n3159 585
R1627 gnd.n2068 gnd.n2067 585
R1628 gnd.n3161 gnd.n2068 585
R1629 gnd.n3164 gnd.n3163 585
R1630 gnd.n3163 gnd.n3162 585
R1631 gnd.n2065 gnd.n2064 585
R1632 gnd.n2064 gnd.n2063 585
R1633 gnd.n3169 gnd.n3168 585
R1634 gnd.n3170 gnd.n3169 585
R1635 gnd.n2062 gnd.n2061 585
R1636 gnd.n3171 gnd.n2062 585
R1637 gnd.n3174 gnd.n3173 585
R1638 gnd.n3173 gnd.n3172 585
R1639 gnd.n2059 gnd.n2058 585
R1640 gnd.n2058 gnd.n2057 585
R1641 gnd.n3179 gnd.n3178 585
R1642 gnd.n3180 gnd.n3179 585
R1643 gnd.n2056 gnd.n2055 585
R1644 gnd.n3181 gnd.n2056 585
R1645 gnd.n3184 gnd.n3183 585
R1646 gnd.n3183 gnd.n3182 585
R1647 gnd.n2053 gnd.n2052 585
R1648 gnd.n2052 gnd.n2051 585
R1649 gnd.n3189 gnd.n3188 585
R1650 gnd.n3190 gnd.n3189 585
R1651 gnd.n2050 gnd.n2049 585
R1652 gnd.n3191 gnd.n2050 585
R1653 gnd.n3194 gnd.n3193 585
R1654 gnd.n3193 gnd.n3192 585
R1655 gnd.n2047 gnd.n2046 585
R1656 gnd.n2046 gnd.n2045 585
R1657 gnd.n3199 gnd.n3198 585
R1658 gnd.n3200 gnd.n3199 585
R1659 gnd.n2044 gnd.n2043 585
R1660 gnd.n3201 gnd.n2044 585
R1661 gnd.n3204 gnd.n3203 585
R1662 gnd.n3203 gnd.n3202 585
R1663 gnd.n2041 gnd.n2040 585
R1664 gnd.n2040 gnd.n2039 585
R1665 gnd.n3209 gnd.n3208 585
R1666 gnd.n3210 gnd.n3209 585
R1667 gnd.n2038 gnd.n2037 585
R1668 gnd.n3211 gnd.n2038 585
R1669 gnd.n3214 gnd.n3213 585
R1670 gnd.n3213 gnd.n3212 585
R1671 gnd.n2035 gnd.n2034 585
R1672 gnd.n2034 gnd.n2033 585
R1673 gnd.n3219 gnd.n3218 585
R1674 gnd.n3220 gnd.n3219 585
R1675 gnd.n2032 gnd.n2031 585
R1676 gnd.n3221 gnd.n2032 585
R1677 gnd.n3224 gnd.n3223 585
R1678 gnd.n3223 gnd.n3222 585
R1679 gnd.n2029 gnd.n2028 585
R1680 gnd.n2028 gnd.n2027 585
R1681 gnd.n3229 gnd.n3228 585
R1682 gnd.n3230 gnd.n3229 585
R1683 gnd.n2026 gnd.n2025 585
R1684 gnd.n3231 gnd.n2026 585
R1685 gnd.n3234 gnd.n3233 585
R1686 gnd.n3233 gnd.n3232 585
R1687 gnd.n2023 gnd.n2022 585
R1688 gnd.n2022 gnd.n2021 585
R1689 gnd.n3239 gnd.n3238 585
R1690 gnd.n3240 gnd.n3239 585
R1691 gnd.n2020 gnd.n2019 585
R1692 gnd.n3241 gnd.n2020 585
R1693 gnd.n3244 gnd.n3243 585
R1694 gnd.n3243 gnd.n3242 585
R1695 gnd.n2017 gnd.n2016 585
R1696 gnd.n2016 gnd.n2015 585
R1697 gnd.n3249 gnd.n3248 585
R1698 gnd.n3250 gnd.n3249 585
R1699 gnd.n2014 gnd.n2013 585
R1700 gnd.n3251 gnd.n2014 585
R1701 gnd.n3254 gnd.n3253 585
R1702 gnd.n3253 gnd.n3252 585
R1703 gnd.n2011 gnd.n2010 585
R1704 gnd.n2010 gnd.n2009 585
R1705 gnd.n3259 gnd.n3258 585
R1706 gnd.n3260 gnd.n3259 585
R1707 gnd.n2008 gnd.n2007 585
R1708 gnd.n3261 gnd.n2008 585
R1709 gnd.n3264 gnd.n3263 585
R1710 gnd.n3263 gnd.n3262 585
R1711 gnd.n2005 gnd.n2004 585
R1712 gnd.n2004 gnd.n2003 585
R1713 gnd.n3269 gnd.n3268 585
R1714 gnd.n3270 gnd.n3269 585
R1715 gnd.n2002 gnd.n2001 585
R1716 gnd.n3271 gnd.n2002 585
R1717 gnd.n3274 gnd.n3273 585
R1718 gnd.n3273 gnd.n3272 585
R1719 gnd.n1999 gnd.n1998 585
R1720 gnd.n1998 gnd.n1997 585
R1721 gnd.n3279 gnd.n3278 585
R1722 gnd.n3280 gnd.n3279 585
R1723 gnd.n1996 gnd.n1995 585
R1724 gnd.n3281 gnd.n1996 585
R1725 gnd.n3284 gnd.n3283 585
R1726 gnd.n3283 gnd.n3282 585
R1727 gnd.n1993 gnd.n1992 585
R1728 gnd.n1992 gnd.n1991 585
R1729 gnd.n3289 gnd.n3288 585
R1730 gnd.n3290 gnd.n3289 585
R1731 gnd.n1990 gnd.n1989 585
R1732 gnd.n3291 gnd.n1990 585
R1733 gnd.n3294 gnd.n3293 585
R1734 gnd.n3293 gnd.n3292 585
R1735 gnd.n1987 gnd.n1986 585
R1736 gnd.n1986 gnd.n1985 585
R1737 gnd.n3299 gnd.n3298 585
R1738 gnd.n3300 gnd.n3299 585
R1739 gnd.n1984 gnd.n1983 585
R1740 gnd.n3301 gnd.n1984 585
R1741 gnd.n3304 gnd.n3303 585
R1742 gnd.n3303 gnd.n3302 585
R1743 gnd.n1981 gnd.n1980 585
R1744 gnd.n1980 gnd.n1979 585
R1745 gnd.n3309 gnd.n3308 585
R1746 gnd.n3310 gnd.n3309 585
R1747 gnd.n1978 gnd.n1977 585
R1748 gnd.n3311 gnd.n1978 585
R1749 gnd.n3314 gnd.n3313 585
R1750 gnd.n3313 gnd.n3312 585
R1751 gnd.n1975 gnd.n1911 585
R1752 gnd.n1911 gnd.n1910 585
R1753 gnd.n3321 gnd.n3320 585
R1754 gnd.n3322 gnd.n3321 585
R1755 gnd.n3109 gnd.n3108 585
R1756 gnd.n3110 gnd.n3109 585
R1757 gnd.n2101 gnd.n2100 585
R1758 gnd.n2100 gnd.n2099 585
R1759 gnd.n3104 gnd.n3103 585
R1760 gnd.n3103 gnd.n3102 585
R1761 gnd.n2104 gnd.n2103 585
R1762 gnd.n3101 gnd.n2104 585
R1763 gnd.n3099 gnd.n3098 585
R1764 gnd.n3100 gnd.n3099 585
R1765 gnd.n3097 gnd.n2106 585
R1766 gnd.n2106 gnd.n2105 585
R1767 gnd.n3096 gnd.n3095 585
R1768 gnd.n3095 gnd.n3094 585
R1769 gnd.n2111 gnd.n2110 585
R1770 gnd.n3093 gnd.n2111 585
R1771 gnd.n3091 gnd.n3090 585
R1772 gnd.n3092 gnd.n3091 585
R1773 gnd.n3089 gnd.n2113 585
R1774 gnd.n2113 gnd.n2112 585
R1775 gnd.n3088 gnd.n3087 585
R1776 gnd.n3087 gnd.n3086 585
R1777 gnd.n2119 gnd.n2118 585
R1778 gnd.n3085 gnd.n2119 585
R1779 gnd.n3083 gnd.n3082 585
R1780 gnd.n3084 gnd.n3083 585
R1781 gnd.n3081 gnd.n2121 585
R1782 gnd.n2121 gnd.n2120 585
R1783 gnd.n3080 gnd.n3079 585
R1784 gnd.n3079 gnd.n3078 585
R1785 gnd.n2127 gnd.n2126 585
R1786 gnd.n3077 gnd.n2127 585
R1787 gnd.n3075 gnd.n3074 585
R1788 gnd.n3076 gnd.n3075 585
R1789 gnd.n3073 gnd.n2129 585
R1790 gnd.n2129 gnd.n2128 585
R1791 gnd.n3072 gnd.n3071 585
R1792 gnd.n3071 gnd.n3070 585
R1793 gnd.n2135 gnd.n2134 585
R1794 gnd.n3069 gnd.n2135 585
R1795 gnd.n3067 gnd.n3066 585
R1796 gnd.n3068 gnd.n3067 585
R1797 gnd.n3065 gnd.n2137 585
R1798 gnd.n2137 gnd.n2136 585
R1799 gnd.n3064 gnd.n3063 585
R1800 gnd.n3063 gnd.n3062 585
R1801 gnd.n2143 gnd.n2142 585
R1802 gnd.n3061 gnd.n2143 585
R1803 gnd.n3059 gnd.n3058 585
R1804 gnd.n3060 gnd.n3059 585
R1805 gnd.n3057 gnd.n2145 585
R1806 gnd.n2145 gnd.n2144 585
R1807 gnd.n3056 gnd.n3055 585
R1808 gnd.n3055 gnd.n3054 585
R1809 gnd.n2151 gnd.n2150 585
R1810 gnd.n3053 gnd.n2151 585
R1811 gnd.n3051 gnd.n3050 585
R1812 gnd.n3052 gnd.n3051 585
R1813 gnd.n3049 gnd.n2153 585
R1814 gnd.n2153 gnd.n2152 585
R1815 gnd.n3048 gnd.n3047 585
R1816 gnd.n3047 gnd.n3046 585
R1817 gnd.n2159 gnd.n2158 585
R1818 gnd.n3045 gnd.n2159 585
R1819 gnd.n3043 gnd.n3042 585
R1820 gnd.n3044 gnd.n3043 585
R1821 gnd.n3041 gnd.n2161 585
R1822 gnd.n2161 gnd.n2160 585
R1823 gnd.n3040 gnd.n3039 585
R1824 gnd.n3039 gnd.n3038 585
R1825 gnd.n2167 gnd.n2166 585
R1826 gnd.n3037 gnd.n2167 585
R1827 gnd.n3035 gnd.n3034 585
R1828 gnd.n3036 gnd.n3035 585
R1829 gnd.n3033 gnd.n2169 585
R1830 gnd.n2169 gnd.n2168 585
R1831 gnd.n3032 gnd.n3031 585
R1832 gnd.n3031 gnd.n3030 585
R1833 gnd.n2175 gnd.n2174 585
R1834 gnd.n3029 gnd.n2175 585
R1835 gnd.n3027 gnd.n3026 585
R1836 gnd.n3028 gnd.n3027 585
R1837 gnd.n3025 gnd.n2177 585
R1838 gnd.n2177 gnd.n2176 585
R1839 gnd.n3024 gnd.n3023 585
R1840 gnd.n3023 gnd.n3022 585
R1841 gnd.n2183 gnd.n2182 585
R1842 gnd.n3021 gnd.n2183 585
R1843 gnd.n3019 gnd.n3018 585
R1844 gnd.n3020 gnd.n3019 585
R1845 gnd.n3017 gnd.n2185 585
R1846 gnd.n2185 gnd.n2184 585
R1847 gnd.n3016 gnd.n3015 585
R1848 gnd.n3015 gnd.n3014 585
R1849 gnd.n2191 gnd.n2190 585
R1850 gnd.n3013 gnd.n2191 585
R1851 gnd.n3011 gnd.n3010 585
R1852 gnd.n3012 gnd.n3011 585
R1853 gnd.n3009 gnd.n2193 585
R1854 gnd.n2193 gnd.n2192 585
R1855 gnd.n3008 gnd.n3007 585
R1856 gnd.n3007 gnd.n3006 585
R1857 gnd.n2199 gnd.n2198 585
R1858 gnd.n3005 gnd.n2199 585
R1859 gnd.n3003 gnd.n3002 585
R1860 gnd.n3004 gnd.n3003 585
R1861 gnd.n3001 gnd.n2201 585
R1862 gnd.n2201 gnd.n2200 585
R1863 gnd.n3000 gnd.n2999 585
R1864 gnd.n2999 gnd.n2998 585
R1865 gnd.n2207 gnd.n2206 585
R1866 gnd.n2997 gnd.n2207 585
R1867 gnd.n2995 gnd.n2994 585
R1868 gnd.n2996 gnd.n2995 585
R1869 gnd.n2993 gnd.n2209 585
R1870 gnd.n2209 gnd.n2208 585
R1871 gnd.n2992 gnd.n2991 585
R1872 gnd.n2991 gnd.n2990 585
R1873 gnd.n2215 gnd.n2214 585
R1874 gnd.n2989 gnd.n2215 585
R1875 gnd.n2987 gnd.n2986 585
R1876 gnd.n2988 gnd.n2987 585
R1877 gnd.n2985 gnd.n2217 585
R1878 gnd.n2217 gnd.n2216 585
R1879 gnd.n2984 gnd.n2983 585
R1880 gnd.n2983 gnd.n2982 585
R1881 gnd.n2223 gnd.n2222 585
R1882 gnd.n2981 gnd.n2223 585
R1883 gnd.n2979 gnd.n2978 585
R1884 gnd.n2980 gnd.n2979 585
R1885 gnd.n2977 gnd.n2225 585
R1886 gnd.n2225 gnd.n2224 585
R1887 gnd.n2976 gnd.n2975 585
R1888 gnd.n2975 gnd.n2974 585
R1889 gnd.n2231 gnd.n2230 585
R1890 gnd.n2973 gnd.n2231 585
R1891 gnd.n2971 gnd.n2970 585
R1892 gnd.n2972 gnd.n2971 585
R1893 gnd.n2969 gnd.n2233 585
R1894 gnd.n2233 gnd.n2232 585
R1895 gnd.n2968 gnd.n2967 585
R1896 gnd.n2967 gnd.n2966 585
R1897 gnd.n2239 gnd.n2238 585
R1898 gnd.n2965 gnd.n2239 585
R1899 gnd.n2963 gnd.n2962 585
R1900 gnd.n2964 gnd.n2963 585
R1901 gnd.n2961 gnd.n2241 585
R1902 gnd.n2241 gnd.n2240 585
R1903 gnd.n2960 gnd.n2959 585
R1904 gnd.n2959 gnd.n2958 585
R1905 gnd.n2247 gnd.n2246 585
R1906 gnd.n2957 gnd.n2247 585
R1907 gnd.n2955 gnd.n2954 585
R1908 gnd.n2956 gnd.n2955 585
R1909 gnd.n2953 gnd.n2249 585
R1910 gnd.n2249 gnd.n2248 585
R1911 gnd.n2952 gnd.n2951 585
R1912 gnd.n2951 gnd.n2950 585
R1913 gnd.n2255 gnd.n2254 585
R1914 gnd.n2949 gnd.n2255 585
R1915 gnd.n2947 gnd.n2946 585
R1916 gnd.n2948 gnd.n2947 585
R1917 gnd.n2945 gnd.n2257 585
R1918 gnd.n2257 gnd.n2256 585
R1919 gnd.n2944 gnd.n2943 585
R1920 gnd.n2943 gnd.n2942 585
R1921 gnd.n2263 gnd.n2262 585
R1922 gnd.n2941 gnd.n2263 585
R1923 gnd.n2939 gnd.n2938 585
R1924 gnd.n2940 gnd.n2939 585
R1925 gnd.n2937 gnd.n2265 585
R1926 gnd.n2265 gnd.n2264 585
R1927 gnd.n2936 gnd.n2935 585
R1928 gnd.n2935 gnd.n2934 585
R1929 gnd.n2271 gnd.n2270 585
R1930 gnd.n2933 gnd.n2271 585
R1931 gnd.n2931 gnd.n2930 585
R1932 gnd.n2932 gnd.n2931 585
R1933 gnd.n2929 gnd.n2273 585
R1934 gnd.n2273 gnd.n2272 585
R1935 gnd.n2928 gnd.n2927 585
R1936 gnd.n2927 gnd.n2926 585
R1937 gnd.n2279 gnd.n2278 585
R1938 gnd.n2925 gnd.n2279 585
R1939 gnd.n2923 gnd.n2922 585
R1940 gnd.n2924 gnd.n2923 585
R1941 gnd.n2921 gnd.n2281 585
R1942 gnd.n2281 gnd.n2280 585
R1943 gnd.n2920 gnd.n2919 585
R1944 gnd.n2919 gnd.n2918 585
R1945 gnd.n2287 gnd.n2286 585
R1946 gnd.n2917 gnd.n2287 585
R1947 gnd.n2915 gnd.n2914 585
R1948 gnd.n2916 gnd.n2915 585
R1949 gnd.n2913 gnd.n2289 585
R1950 gnd.n2289 gnd.n2288 585
R1951 gnd.n2912 gnd.n2911 585
R1952 gnd.n2911 gnd.n2910 585
R1953 gnd.n2295 gnd.n2294 585
R1954 gnd.n2909 gnd.n2295 585
R1955 gnd.n2907 gnd.n2906 585
R1956 gnd.n2908 gnd.n2907 585
R1957 gnd.n2905 gnd.n2297 585
R1958 gnd.n2297 gnd.n2296 585
R1959 gnd.n2904 gnd.n2903 585
R1960 gnd.n2903 gnd.n2902 585
R1961 gnd.n2303 gnd.n2302 585
R1962 gnd.n2901 gnd.n2303 585
R1963 gnd.n2899 gnd.n2898 585
R1964 gnd.n2900 gnd.n2899 585
R1965 gnd.n2897 gnd.n2305 585
R1966 gnd.n2305 gnd.n2304 585
R1967 gnd.n2896 gnd.n2895 585
R1968 gnd.n2895 gnd.n2894 585
R1969 gnd.n2311 gnd.n2310 585
R1970 gnd.n2893 gnd.n2311 585
R1971 gnd.n2891 gnd.n2890 585
R1972 gnd.n2892 gnd.n2891 585
R1973 gnd.n2889 gnd.n2313 585
R1974 gnd.n2313 gnd.n2312 585
R1975 gnd.n2888 gnd.n2887 585
R1976 gnd.n2887 gnd.n2886 585
R1977 gnd.n2319 gnd.n2318 585
R1978 gnd.n2885 gnd.n2319 585
R1979 gnd.n2883 gnd.n2882 585
R1980 gnd.n2884 gnd.n2883 585
R1981 gnd.n2881 gnd.n2321 585
R1982 gnd.n2321 gnd.n2320 585
R1983 gnd.n2880 gnd.n2879 585
R1984 gnd.n2879 gnd.n2878 585
R1985 gnd.n2327 gnd.n2326 585
R1986 gnd.n2877 gnd.n2327 585
R1987 gnd.n2875 gnd.n2874 585
R1988 gnd.n2876 gnd.n2875 585
R1989 gnd.n2873 gnd.n2329 585
R1990 gnd.n2329 gnd.n2328 585
R1991 gnd.n2872 gnd.n2871 585
R1992 gnd.n2871 gnd.n2870 585
R1993 gnd.n2335 gnd.n2334 585
R1994 gnd.n2869 gnd.n2335 585
R1995 gnd.n2867 gnd.n2866 585
R1996 gnd.n2868 gnd.n2867 585
R1997 gnd.n2865 gnd.n2337 585
R1998 gnd.n2337 gnd.n2336 585
R1999 gnd.n2864 gnd.n2863 585
R2000 gnd.n2863 gnd.n2862 585
R2001 gnd.n2343 gnd.n2342 585
R2002 gnd.n2861 gnd.n2343 585
R2003 gnd.n2859 gnd.n2858 585
R2004 gnd.n2860 gnd.n2859 585
R2005 gnd.n2857 gnd.n2345 585
R2006 gnd.n2345 gnd.n2344 585
R2007 gnd.n2856 gnd.n2855 585
R2008 gnd.n2855 gnd.n2854 585
R2009 gnd.n2351 gnd.n2350 585
R2010 gnd.n2853 gnd.n2351 585
R2011 gnd.n2851 gnd.n2850 585
R2012 gnd.n2852 gnd.n2851 585
R2013 gnd.n2849 gnd.n2353 585
R2014 gnd.n2353 gnd.n2352 585
R2015 gnd.n2848 gnd.n2847 585
R2016 gnd.n2847 gnd.n2846 585
R2017 gnd.n2359 gnd.n2358 585
R2018 gnd.n2845 gnd.n2359 585
R2019 gnd.n2843 gnd.n2842 585
R2020 gnd.n2844 gnd.n2843 585
R2021 gnd.n2841 gnd.n2361 585
R2022 gnd.n2361 gnd.n2360 585
R2023 gnd.n2840 gnd.n2839 585
R2024 gnd.n2839 gnd.n2838 585
R2025 gnd.n2367 gnd.n2366 585
R2026 gnd.n2837 gnd.n2367 585
R2027 gnd.n2835 gnd.n2834 585
R2028 gnd.n2836 gnd.n2835 585
R2029 gnd.n2833 gnd.n2369 585
R2030 gnd.n2369 gnd.n2368 585
R2031 gnd.n2832 gnd.n2831 585
R2032 gnd.n2831 gnd.n2830 585
R2033 gnd.n2375 gnd.n2374 585
R2034 gnd.n2829 gnd.n2375 585
R2035 gnd.n2827 gnd.n2826 585
R2036 gnd.n2828 gnd.n2827 585
R2037 gnd.n2825 gnd.n2377 585
R2038 gnd.n2377 gnd.n2376 585
R2039 gnd.n2824 gnd.n2823 585
R2040 gnd.n2823 gnd.n2822 585
R2041 gnd.n2383 gnd.n2382 585
R2042 gnd.n2821 gnd.n2383 585
R2043 gnd.n2819 gnd.n2818 585
R2044 gnd.n2820 gnd.n2819 585
R2045 gnd.n2817 gnd.n2385 585
R2046 gnd.n2385 gnd.n2384 585
R2047 gnd.n2816 gnd.n2815 585
R2048 gnd.n2815 gnd.n2814 585
R2049 gnd.n2391 gnd.n2390 585
R2050 gnd.n2813 gnd.n2391 585
R2051 gnd.n2811 gnd.n2810 585
R2052 gnd.n2812 gnd.n2811 585
R2053 gnd.n2809 gnd.n2393 585
R2054 gnd.n2393 gnd.n2392 585
R2055 gnd.n2808 gnd.n2807 585
R2056 gnd.n2807 gnd.n2806 585
R2057 gnd.n2399 gnd.n2398 585
R2058 gnd.n2805 gnd.n2399 585
R2059 gnd.n2803 gnd.n2802 585
R2060 gnd.n2804 gnd.n2803 585
R2061 gnd.n2801 gnd.n2401 585
R2062 gnd.n2401 gnd.n2400 585
R2063 gnd.n2800 gnd.n2799 585
R2064 gnd.n2799 gnd.n2798 585
R2065 gnd.n2407 gnd.n2406 585
R2066 gnd.n2797 gnd.n2407 585
R2067 gnd.n2795 gnd.n2794 585
R2068 gnd.n2796 gnd.n2795 585
R2069 gnd.n2793 gnd.n2409 585
R2070 gnd.n2409 gnd.n2408 585
R2071 gnd.n2792 gnd.n2791 585
R2072 gnd.n2791 gnd.n2790 585
R2073 gnd.n2415 gnd.n2414 585
R2074 gnd.n2789 gnd.n2415 585
R2075 gnd.n2787 gnd.n2786 585
R2076 gnd.n2788 gnd.n2787 585
R2077 gnd.n2785 gnd.n2417 585
R2078 gnd.n2417 gnd.n2416 585
R2079 gnd.n2784 gnd.n2783 585
R2080 gnd.n2783 gnd.n2782 585
R2081 gnd.n2423 gnd.n2422 585
R2082 gnd.n2781 gnd.n2423 585
R2083 gnd.n2779 gnd.n2778 585
R2084 gnd.n2780 gnd.n2779 585
R2085 gnd.n2777 gnd.n2425 585
R2086 gnd.n2425 gnd.n2424 585
R2087 gnd.n2776 gnd.n2775 585
R2088 gnd.n2775 gnd.n2774 585
R2089 gnd.n2431 gnd.n2430 585
R2090 gnd.n2773 gnd.n2431 585
R2091 gnd.n2605 gnd.n2604 585
R2092 gnd.n2604 gnd.n2603 585
R2093 gnd.n2606 gnd.n2594 585
R2094 gnd.n2594 gnd.n2593 585
R2095 gnd.n2608 gnd.n2607 585
R2096 gnd.n2609 gnd.n2608 585
R2097 gnd.n2592 gnd.n2591 585
R2098 gnd.n2610 gnd.n2592 585
R2099 gnd.n2613 gnd.n2612 585
R2100 gnd.n2612 gnd.n2611 585
R2101 gnd.n2614 gnd.n2586 585
R2102 gnd.n2586 gnd.n2585 585
R2103 gnd.n2616 gnd.n2615 585
R2104 gnd.n2617 gnd.n2616 585
R2105 gnd.n2584 gnd.n2583 585
R2106 gnd.n2618 gnd.n2584 585
R2107 gnd.n2621 gnd.n2620 585
R2108 gnd.n2620 gnd.n2619 585
R2109 gnd.n2622 gnd.n2578 585
R2110 gnd.n2578 gnd.n2577 585
R2111 gnd.n2624 gnd.n2623 585
R2112 gnd.n2625 gnd.n2624 585
R2113 gnd.n2576 gnd.n2575 585
R2114 gnd.n2626 gnd.n2576 585
R2115 gnd.n2629 gnd.n2628 585
R2116 gnd.n2628 gnd.n2627 585
R2117 gnd.n2630 gnd.n2570 585
R2118 gnd.n2570 gnd.n2569 585
R2119 gnd.n2632 gnd.n2631 585
R2120 gnd.n2633 gnd.n2632 585
R2121 gnd.n2568 gnd.n2567 585
R2122 gnd.n2634 gnd.n2568 585
R2123 gnd.n2637 gnd.n2636 585
R2124 gnd.n2636 gnd.n2635 585
R2125 gnd.n2638 gnd.n2562 585
R2126 gnd.n2562 gnd.n2561 585
R2127 gnd.n2640 gnd.n2639 585
R2128 gnd.n2641 gnd.n2640 585
R2129 gnd.n2560 gnd.n2559 585
R2130 gnd.n2642 gnd.n2560 585
R2131 gnd.n2645 gnd.n2644 585
R2132 gnd.n2644 gnd.n2643 585
R2133 gnd.n2646 gnd.n2554 585
R2134 gnd.n2554 gnd.n2553 585
R2135 gnd.n2648 gnd.n2647 585
R2136 gnd.n2649 gnd.n2648 585
R2137 gnd.n2552 gnd.n2551 585
R2138 gnd.n2650 gnd.n2552 585
R2139 gnd.n2653 gnd.n2652 585
R2140 gnd.n2652 gnd.n2651 585
R2141 gnd.n2654 gnd.n2546 585
R2142 gnd.n2546 gnd.n2545 585
R2143 gnd.n2656 gnd.n2655 585
R2144 gnd.n2657 gnd.n2656 585
R2145 gnd.n2544 gnd.n2543 585
R2146 gnd.n2658 gnd.n2544 585
R2147 gnd.n2661 gnd.n2660 585
R2148 gnd.n2660 gnd.n2659 585
R2149 gnd.n2662 gnd.n2538 585
R2150 gnd.n2538 gnd.n2537 585
R2151 gnd.n2664 gnd.n2663 585
R2152 gnd.n2665 gnd.n2664 585
R2153 gnd.n2536 gnd.n2535 585
R2154 gnd.n2666 gnd.n2536 585
R2155 gnd.n2669 gnd.n2668 585
R2156 gnd.n2668 gnd.n2667 585
R2157 gnd.n2670 gnd.n2530 585
R2158 gnd.n2530 gnd.n2529 585
R2159 gnd.n2672 gnd.n2671 585
R2160 gnd.n2673 gnd.n2672 585
R2161 gnd.n2528 gnd.n2527 585
R2162 gnd.n2674 gnd.n2528 585
R2163 gnd.n2677 gnd.n2676 585
R2164 gnd.n2676 gnd.n2675 585
R2165 gnd.n2678 gnd.n2522 585
R2166 gnd.n2522 gnd.n2521 585
R2167 gnd.n2680 gnd.n2679 585
R2168 gnd.n2681 gnd.n2680 585
R2169 gnd.n2520 gnd.n2519 585
R2170 gnd.n2682 gnd.n2520 585
R2171 gnd.n2685 gnd.n2684 585
R2172 gnd.n2684 gnd.n2683 585
R2173 gnd.n2686 gnd.n2514 585
R2174 gnd.n2514 gnd.n2513 585
R2175 gnd.n2688 gnd.n2687 585
R2176 gnd.n2689 gnd.n2688 585
R2177 gnd.n2512 gnd.n2511 585
R2178 gnd.n2690 gnd.n2512 585
R2179 gnd.n2693 gnd.n2692 585
R2180 gnd.n2692 gnd.n2691 585
R2181 gnd.n2694 gnd.n2506 585
R2182 gnd.n2506 gnd.n2505 585
R2183 gnd.n2696 gnd.n2695 585
R2184 gnd.n2697 gnd.n2696 585
R2185 gnd.n2504 gnd.n2503 585
R2186 gnd.n2698 gnd.n2504 585
R2187 gnd.n2701 gnd.n2700 585
R2188 gnd.n2700 gnd.n2699 585
R2189 gnd.n2702 gnd.n2498 585
R2190 gnd.n2498 gnd.n2497 585
R2191 gnd.n2704 gnd.n2703 585
R2192 gnd.n2705 gnd.n2704 585
R2193 gnd.n2496 gnd.n2495 585
R2194 gnd.n2706 gnd.n2496 585
R2195 gnd.n2709 gnd.n2708 585
R2196 gnd.n2708 gnd.n2707 585
R2197 gnd.n2710 gnd.n2490 585
R2198 gnd.n2490 gnd.n2489 585
R2199 gnd.n2712 gnd.n2711 585
R2200 gnd.n2713 gnd.n2712 585
R2201 gnd.n2488 gnd.n2487 585
R2202 gnd.n2714 gnd.n2488 585
R2203 gnd.n2717 gnd.n2716 585
R2204 gnd.n2716 gnd.n2715 585
R2205 gnd.n2718 gnd.n2482 585
R2206 gnd.n2482 gnd.n2481 585
R2207 gnd.n2720 gnd.n2719 585
R2208 gnd.n2721 gnd.n2720 585
R2209 gnd.n2480 gnd.n2479 585
R2210 gnd.n2722 gnd.n2480 585
R2211 gnd.n2725 gnd.n2724 585
R2212 gnd.n2724 gnd.n2723 585
R2213 gnd.n2726 gnd.n2474 585
R2214 gnd.n2474 gnd.n2473 585
R2215 gnd.n2728 gnd.n2727 585
R2216 gnd.n2729 gnd.n2728 585
R2217 gnd.n2472 gnd.n2471 585
R2218 gnd.n2730 gnd.n2472 585
R2219 gnd.n2733 gnd.n2732 585
R2220 gnd.n2732 gnd.n2731 585
R2221 gnd.n2734 gnd.n2466 585
R2222 gnd.n2466 gnd.n2465 585
R2223 gnd.n2736 gnd.n2735 585
R2224 gnd.n2737 gnd.n2736 585
R2225 gnd.n2464 gnd.n2463 585
R2226 gnd.n2738 gnd.n2464 585
R2227 gnd.n2741 gnd.n2740 585
R2228 gnd.n2740 gnd.n2739 585
R2229 gnd.n2742 gnd.n2458 585
R2230 gnd.n2458 gnd.n2457 585
R2231 gnd.n2744 gnd.n2743 585
R2232 gnd.n2745 gnd.n2744 585
R2233 gnd.n2456 gnd.n2455 585
R2234 gnd.n2746 gnd.n2456 585
R2235 gnd.n2749 gnd.n2748 585
R2236 gnd.n2748 gnd.n2747 585
R2237 gnd.n2750 gnd.n2450 585
R2238 gnd.n2450 gnd.n2449 585
R2239 gnd.n2752 gnd.n2751 585
R2240 gnd.n2753 gnd.n2752 585
R2241 gnd.n2448 gnd.n2447 585
R2242 gnd.n2754 gnd.n2448 585
R2243 gnd.n2757 gnd.n2756 585
R2244 gnd.n2756 gnd.n2755 585
R2245 gnd.n2758 gnd.n2443 585
R2246 gnd.n2443 gnd.n2442 585
R2247 gnd.n2760 gnd.n2759 585
R2248 gnd.n2761 gnd.n2760 585
R2249 gnd.n2440 gnd.n2438 585
R2250 gnd.n2762 gnd.n2440 585
R2251 gnd.n2765 gnd.n2764 585
R2252 gnd.n2764 gnd.n2763 585
R2253 gnd.n2439 gnd.n2436 585
R2254 gnd.n2441 gnd.n2439 585
R2255 gnd.n2769 gnd.n2433 585
R2256 gnd.n2433 gnd.n2432 585
R2257 gnd.n2771 gnd.n2770 585
R2258 gnd.n2772 gnd.n2771 585
R2259 gnd.n5699 gnd.n1423 585
R2260 gnd.n5699 gnd.n5698 585
R2261 gnd.n5860 gnd.n1429 585
R2262 gnd.n5966 gnd.n1429 585
R2263 gnd.n5861 gnd.n1441 585
R2264 gnd.n1452 gnd.n1441 585
R2265 gnd.n5863 gnd.n5862 585
R2266 gnd.n5864 gnd.n5863 585
R2267 gnd.n1442 gnd.n1440 585
R2268 gnd.n5854 gnd.n1440 585
R2269 gnd.n5440 gnd.n1499 585
R2270 gnd.n5452 gnd.n1499 585
R2271 gnd.n5441 gnd.n1510 585
R2272 gnd.n1510 gnd.n1498 585
R2273 gnd.n5443 gnd.n5442 585
R2274 gnd.n5444 gnd.n5443 585
R2275 gnd.n1511 gnd.n1509 585
R2276 gnd.n5432 gnd.n1509 585
R2277 gnd.n5405 gnd.n5404 585
R2278 gnd.n5404 gnd.n5403 585
R2279 gnd.n5406 gnd.n1525 585
R2280 gnd.n5420 gnd.n1525 585
R2281 gnd.n5407 gnd.n1537 585
R2282 gnd.n5353 gnd.n1537 585
R2283 gnd.n5409 gnd.n5408 585
R2284 gnd.n5410 gnd.n5409 585
R2285 gnd.n1538 gnd.n1536 585
R2286 gnd.n5386 gnd.n1536 585
R2287 gnd.n5362 gnd.n5361 585
R2288 gnd.n5361 gnd.n1550 585
R2289 gnd.n5363 gnd.n1561 585
R2290 gnd.n5377 gnd.n1561 585
R2291 gnd.n5364 gnd.n1573 585
R2292 gnd.n5348 gnd.n1573 585
R2293 gnd.n5366 gnd.n5365 585
R2294 gnd.n5367 gnd.n5366 585
R2295 gnd.n1574 gnd.n1572 585
R2296 gnd.n5344 gnd.n1572 585
R2297 gnd.n5320 gnd.n5319 585
R2298 gnd.n5319 gnd.n5318 585
R2299 gnd.n5321 gnd.n1592 585
R2300 gnd.n5335 gnd.n1592 585
R2301 gnd.n5322 gnd.n1604 585
R2302 gnd.n5312 gnd.n1604 585
R2303 gnd.n5324 gnd.n5323 585
R2304 gnd.n5325 gnd.n5324 585
R2305 gnd.n1605 gnd.n1603 585
R2306 gnd.n5308 gnd.n1603 585
R2307 gnd.n5284 gnd.n5283 585
R2308 gnd.n5283 gnd.n5282 585
R2309 gnd.n5285 gnd.n1621 585
R2310 gnd.n5299 gnd.n1621 585
R2311 gnd.n5286 gnd.n1639 585
R2312 gnd.n5276 gnd.n1639 585
R2313 gnd.n5288 gnd.n5287 585
R2314 gnd.n5289 gnd.n5288 585
R2315 gnd.n1640 gnd.n1638 585
R2316 gnd.n5272 gnd.n1638 585
R2317 gnd.n5257 gnd.n5256 585
R2318 gnd.n5258 gnd.n5257 585
R2319 gnd.n1658 gnd.n1655 585
R2320 gnd.n5263 gnd.n1655 585
R2321 gnd.n5249 gnd.n5248 585
R2322 gnd.n5250 gnd.n5249 585
R2323 gnd.n5247 gnd.n1663 585
R2324 gnd.n5237 gnd.n1663 585
R2325 gnd.n1671 gnd.n1664 585
R2326 gnd.n5242 gnd.n1671 585
R2327 gnd.n5228 gnd.n5227 585
R2328 gnd.n5229 gnd.n5228 585
R2329 gnd.n5226 gnd.n1680 585
R2330 gnd.n5222 gnd.n1680 585
R2331 gnd.n5216 gnd.n1681 585
R2332 gnd.n5217 gnd.n5216 585
R2333 gnd.n5215 gnd.n1690 585
R2334 gnd.n5215 gnd.n5214 585
R2335 gnd.n5189 gnd.n1689 585
R2336 gnd.n5185 gnd.n1689 585
R2337 gnd.n5190 gnd.n1700 585
R2338 gnd.n5204 gnd.n1700 585
R2339 gnd.n5191 gnd.n1710 585
R2340 gnd.n1710 gnd.n1698 585
R2341 gnd.n5193 gnd.n5192 585
R2342 gnd.n5194 gnd.n5193 585
R2343 gnd.n1711 gnd.n1709 585
R2344 gnd.n5177 gnd.n1709 585
R2345 gnd.n5152 gnd.n5151 585
R2346 gnd.n5151 gnd.n1719 585
R2347 gnd.n5153 gnd.n1727 585
R2348 gnd.n5167 gnd.n1727 585
R2349 gnd.n5154 gnd.n1737 585
R2350 gnd.n1737 gnd.n1725 585
R2351 gnd.n5156 gnd.n5155 585
R2352 gnd.n5157 gnd.n5156 585
R2353 gnd.n1738 gnd.n1736 585
R2354 gnd.n5142 gnd.n1736 585
R2355 gnd.n5117 gnd.n5116 585
R2356 gnd.n5116 gnd.n1744 585
R2357 gnd.n5118 gnd.n1751 585
R2358 gnd.n5132 gnd.n1751 585
R2359 gnd.n5119 gnd.n1762 585
R2360 gnd.n1762 gnd.n1760 585
R2361 gnd.n5121 gnd.n5120 585
R2362 gnd.n5122 gnd.n5121 585
R2363 gnd.n1763 gnd.n1761 585
R2364 gnd.n5107 gnd.n1761 585
R2365 gnd.n5082 gnd.n5081 585
R2366 gnd.n5081 gnd.n1769 585
R2367 gnd.n5083 gnd.n1776 585
R2368 gnd.n5097 gnd.n1776 585
R2369 gnd.n5084 gnd.n1788 585
R2370 gnd.n1788 gnd.n1786 585
R2371 gnd.n5086 gnd.n5085 585
R2372 gnd.n5087 gnd.n5086 585
R2373 gnd.n1789 gnd.n1787 585
R2374 gnd.n1787 gnd.n1783 585
R2375 gnd.n5059 gnd.n1797 585
R2376 gnd.n5071 gnd.n1797 585
R2377 gnd.n5060 gnd.n1807 585
R2378 gnd.n1807 gnd.n1795 585
R2379 gnd.n5062 gnd.n5061 585
R2380 gnd.n5063 gnd.n5062 585
R2381 gnd.n1808 gnd.n1806 585
R2382 gnd.n1806 gnd.n1803 585
R2383 gnd.n5035 gnd.n1814 585
R2384 gnd.n5051 gnd.n1814 585
R2385 gnd.n5040 gnd.n4732 585
R2386 gnd.n4732 gnd.n4730 585
R2387 gnd.n5042 gnd.n5041 585
R2388 gnd.n5043 gnd.n5042 585
R2389 gnd.n4820 gnd.n4731 585
R2390 gnd.n4819 gnd.n4818 585
R2391 gnd.n4816 gnd.n4734 585
R2392 gnd.n4814 gnd.n4813 585
R2393 gnd.n4812 gnd.n4735 585
R2394 gnd.n4811 gnd.n4810 585
R2395 gnd.n4808 gnd.n4740 585
R2396 gnd.n4806 gnd.n4805 585
R2397 gnd.n4804 gnd.n4741 585
R2398 gnd.n4803 gnd.n4802 585
R2399 gnd.n4800 gnd.n4746 585
R2400 gnd.n4798 gnd.n4797 585
R2401 gnd.n4796 gnd.n4747 585
R2402 gnd.n4795 gnd.n4794 585
R2403 gnd.n4792 gnd.n4752 585
R2404 gnd.n4790 gnd.n4789 585
R2405 gnd.n4788 gnd.n4753 585
R2406 gnd.n4782 gnd.n4758 585
R2407 gnd.n4784 gnd.n4783 585
R2408 gnd.n4783 gnd.n4727 585
R2409 gnd.n5767 gnd.n5766 585
R2410 gnd.n5768 gnd.n5764 585
R2411 gnd.n5779 gnd.n5761 585
R2412 gnd.n5780 gnd.n5759 585
R2413 gnd.n5758 gnd.n5751 585
R2414 gnd.n5787 gnd.n5750 585
R2415 gnd.n5788 gnd.n5749 585
R2416 gnd.n5747 gnd.n5739 585
R2417 gnd.n5795 gnd.n5738 585
R2418 gnd.n5796 gnd.n5736 585
R2419 gnd.n5735 gnd.n5728 585
R2420 gnd.n5803 gnd.n5727 585
R2421 gnd.n5804 gnd.n5726 585
R2422 gnd.n5724 gnd.n5716 585
R2423 gnd.n5811 gnd.n5715 585
R2424 gnd.n5812 gnd.n5713 585
R2425 gnd.n5712 gnd.n5702 585
R2426 gnd.n5819 gnd.n5701 585
R2427 gnd.n5820 gnd.n5700 585
R2428 gnd.n5700 gnd.n1369 585
R2429 gnd.n5846 gnd.n1454 585
R2430 gnd.n5698 gnd.n1454 585
R2431 gnd.n5847 gnd.n1427 585
R2432 gnd.n5966 gnd.n1427 585
R2433 gnd.n5848 gnd.n1453 585
R2434 gnd.n1453 gnd.n1452 585
R2435 gnd.n1449 gnd.n1438 585
R2436 gnd.n5864 gnd.n1438 585
R2437 gnd.n5853 gnd.n5852 585
R2438 gnd.n5854 gnd.n5853 585
R2439 gnd.n1448 gnd.n1447 585
R2440 gnd.n5452 gnd.n1447 585
R2441 gnd.n5426 gnd.n5425 585
R2442 gnd.n5425 gnd.n1498 585
R2443 gnd.n1519 gnd.n1507 585
R2444 gnd.n5444 gnd.n1507 585
R2445 gnd.n5431 gnd.n5430 585
R2446 gnd.n5432 gnd.n5431 585
R2447 gnd.n1518 gnd.n1517 585
R2448 gnd.n5403 gnd.n1517 585
R2449 gnd.n5422 gnd.n5421 585
R2450 gnd.n5421 gnd.n5420 585
R2451 gnd.n1522 gnd.n1521 585
R2452 gnd.n5353 gnd.n1522 585
R2453 gnd.n1554 gnd.n1534 585
R2454 gnd.n5410 gnd.n1534 585
R2455 gnd.n5385 gnd.n5384 585
R2456 gnd.n5386 gnd.n5385 585
R2457 gnd.n1553 gnd.n1552 585
R2458 gnd.n1552 gnd.n1550 585
R2459 gnd.n5379 gnd.n5378 585
R2460 gnd.n5378 gnd.n5377 585
R2461 gnd.n1557 gnd.n1556 585
R2462 gnd.n5348 gnd.n1557 585
R2463 gnd.n1585 gnd.n1570 585
R2464 gnd.n5367 gnd.n1570 585
R2465 gnd.n5343 gnd.n5342 585
R2466 gnd.n5344 gnd.n5343 585
R2467 gnd.n1584 gnd.n1583 585
R2468 gnd.n5318 gnd.n1583 585
R2469 gnd.n5337 gnd.n5336 585
R2470 gnd.n5336 gnd.n5335 585
R2471 gnd.n1588 gnd.n1587 585
R2472 gnd.n5312 gnd.n1588 585
R2473 gnd.n1614 gnd.n1601 585
R2474 gnd.n5325 gnd.n1601 585
R2475 gnd.n5307 gnd.n5306 585
R2476 gnd.n5308 gnd.n5307 585
R2477 gnd.n1613 gnd.n1612 585
R2478 gnd.n5282 gnd.n1612 585
R2479 gnd.n5301 gnd.n5300 585
R2480 gnd.n5300 gnd.n5299 585
R2481 gnd.n1617 gnd.n1616 585
R2482 gnd.n5276 gnd.n1617 585
R2483 gnd.n1648 gnd.n1636 585
R2484 gnd.n5289 gnd.n1636 585
R2485 gnd.n5271 gnd.n5270 585
R2486 gnd.n5272 gnd.n5271 585
R2487 gnd.n1647 gnd.n1646 585
R2488 gnd.n5258 gnd.n1646 585
R2489 gnd.n5265 gnd.n5264 585
R2490 gnd.n5264 gnd.n5263 585
R2491 gnd.n1651 gnd.n1650 585
R2492 gnd.n5250 gnd.n1651 585
R2493 gnd.n5236 gnd.n5235 585
R2494 gnd.n5237 gnd.n5236 585
R2495 gnd.n1675 gnd.n1669 585
R2496 gnd.n5242 gnd.n1669 585
R2497 gnd.n5231 gnd.n5230 585
R2498 gnd.n5230 gnd.n5229 585
R2499 gnd.n1678 gnd.n1677 585
R2500 gnd.n5222 gnd.n1678 585
R2501 gnd.n5211 gnd.n1688 585
R2502 gnd.n5217 gnd.n1688 585
R2503 gnd.n5213 gnd.n5212 585
R2504 gnd.n5214 gnd.n5213 585
R2505 gnd.n1694 gnd.n1693 585
R2506 gnd.n5185 gnd.n1693 585
R2507 gnd.n5206 gnd.n5205 585
R2508 gnd.n5205 gnd.n5204 585
R2509 gnd.n1697 gnd.n1696 585
R2510 gnd.n1698 gnd.n1697 585
R2511 gnd.n5174 gnd.n1708 585
R2512 gnd.n5194 gnd.n1708 585
R2513 gnd.n5176 gnd.n5175 585
R2514 gnd.n5177 gnd.n5176 585
R2515 gnd.n1721 gnd.n1720 585
R2516 gnd.n1720 gnd.n1719 585
R2517 gnd.n5169 gnd.n5168 585
R2518 gnd.n5168 gnd.n5167 585
R2519 gnd.n1724 gnd.n1723 585
R2520 gnd.n1725 gnd.n1724 585
R2521 gnd.n5139 gnd.n1735 585
R2522 gnd.n5157 gnd.n1735 585
R2523 gnd.n5141 gnd.n5140 585
R2524 gnd.n5142 gnd.n5141 585
R2525 gnd.n1746 gnd.n1745 585
R2526 gnd.n1745 gnd.n1744 585
R2527 gnd.n5134 gnd.n5133 585
R2528 gnd.n5133 gnd.n5132 585
R2529 gnd.n1749 gnd.n1748 585
R2530 gnd.n1760 gnd.n1749 585
R2531 gnd.n5104 gnd.n1759 585
R2532 gnd.n5122 gnd.n1759 585
R2533 gnd.n5106 gnd.n5105 585
R2534 gnd.n5107 gnd.n5106 585
R2535 gnd.n1771 gnd.n1770 585
R2536 gnd.n1770 gnd.n1769 585
R2537 gnd.n5099 gnd.n5098 585
R2538 gnd.n5098 gnd.n5097 585
R2539 gnd.n1774 gnd.n1773 585
R2540 gnd.n1786 gnd.n1774 585
R2541 gnd.n4767 gnd.n1785 585
R2542 gnd.n5087 gnd.n1785 585
R2543 gnd.n4769 gnd.n4768 585
R2544 gnd.n4768 gnd.n1783 585
R2545 gnd.n4770 gnd.n1796 585
R2546 gnd.n5071 gnd.n1796 585
R2547 gnd.n4772 gnd.n4771 585
R2548 gnd.n4771 gnd.n1795 585
R2549 gnd.n4773 gnd.n1805 585
R2550 gnd.n5063 gnd.n1805 585
R2551 gnd.n4775 gnd.n4774 585
R2552 gnd.n4774 gnd.n1803 585
R2553 gnd.n4776 gnd.n1813 585
R2554 gnd.n5051 gnd.n1813 585
R2555 gnd.n4778 gnd.n4777 585
R2556 gnd.n4777 gnd.n4730 585
R2557 gnd.n4779 gnd.n4729 585
R2558 gnd.n5043 gnd.n4729 585
R2559 gnd.n4634 gnd.n4633 585
R2560 gnd.n4635 gnd.n4634 585
R2561 gnd.n1895 gnd.n1894 585
R2562 gnd.n1901 gnd.n1894 585
R2563 gnd.n4608 gnd.n3326 585
R2564 gnd.n3326 gnd.n1900 585
R2565 gnd.n4610 gnd.n4609 585
R2566 gnd.n4611 gnd.n4610 585
R2567 gnd.n3327 gnd.n3325 585
R2568 gnd.n3325 gnd.n1908 585
R2569 gnd.n4342 gnd.n4341 585
R2570 gnd.n4341 gnd.n4340 585
R2571 gnd.n3332 gnd.n3331 585
R2572 gnd.n4311 gnd.n3332 585
R2573 gnd.n4331 gnd.n4330 585
R2574 gnd.n4330 gnd.n4329 585
R2575 gnd.n3339 gnd.n3338 585
R2576 gnd.n4317 gnd.n3339 585
R2577 gnd.n4287 gnd.n3359 585
R2578 gnd.n3359 gnd.n3358 585
R2579 gnd.n4289 gnd.n4288 585
R2580 gnd.n4290 gnd.n4289 585
R2581 gnd.n3360 gnd.n3357 585
R2582 gnd.n3368 gnd.n3357 585
R2583 gnd.n4265 gnd.n3380 585
R2584 gnd.n3380 gnd.n3367 585
R2585 gnd.n4267 gnd.n4266 585
R2586 gnd.n4268 gnd.n4267 585
R2587 gnd.n3381 gnd.n3379 585
R2588 gnd.n3379 gnd.n3375 585
R2589 gnd.n4253 gnd.n4252 585
R2590 gnd.n4252 gnd.n4251 585
R2591 gnd.n3386 gnd.n3385 585
R2592 gnd.n3396 gnd.n3386 585
R2593 gnd.n4242 gnd.n4241 585
R2594 gnd.n4241 gnd.n4240 585
R2595 gnd.n3393 gnd.n3392 585
R2596 gnd.n4228 gnd.n3393 585
R2597 gnd.n4202 gnd.n3414 585
R2598 gnd.n3414 gnd.n3403 585
R2599 gnd.n4204 gnd.n4203 585
R2600 gnd.n4205 gnd.n4204 585
R2601 gnd.n3415 gnd.n3413 585
R2602 gnd.n3423 gnd.n3413 585
R2603 gnd.n4180 gnd.n3435 585
R2604 gnd.n3435 gnd.n3422 585
R2605 gnd.n4182 gnd.n4181 585
R2606 gnd.n4183 gnd.n4182 585
R2607 gnd.n3436 gnd.n3434 585
R2608 gnd.n3434 gnd.n3430 585
R2609 gnd.n4168 gnd.n4167 585
R2610 gnd.n4167 gnd.n4166 585
R2611 gnd.n3441 gnd.n3440 585
R2612 gnd.n3450 gnd.n3441 585
R2613 gnd.n4157 gnd.n4156 585
R2614 gnd.n4156 gnd.n4155 585
R2615 gnd.n3448 gnd.n3447 585
R2616 gnd.n4143 gnd.n3448 585
R2617 gnd.n3581 gnd.n3580 585
R2618 gnd.n3581 gnd.n3457 585
R2619 gnd.n4100 gnd.n4099 585
R2620 gnd.n4099 gnd.n4098 585
R2621 gnd.n4101 gnd.n3575 585
R2622 gnd.n3586 gnd.n3575 585
R2623 gnd.n4103 gnd.n4102 585
R2624 gnd.n4104 gnd.n4103 585
R2625 gnd.n3576 gnd.n3574 585
R2626 gnd.n3599 gnd.n3574 585
R2627 gnd.n3559 gnd.n3558 585
R2628 gnd.n3562 gnd.n3559 585
R2629 gnd.n4114 gnd.n4113 585
R2630 gnd.n4113 gnd.n4112 585
R2631 gnd.n4115 gnd.n3553 585
R2632 gnd.n4074 gnd.n3553 585
R2633 gnd.n4117 gnd.n4116 585
R2634 gnd.n4118 gnd.n4117 585
R2635 gnd.n3554 gnd.n3552 585
R2636 gnd.n3613 gnd.n3552 585
R2637 gnd.n4066 gnd.n4065 585
R2638 gnd.n4065 gnd.n4064 585
R2639 gnd.n3610 gnd.n3609 585
R2640 gnd.n4048 gnd.n3610 585
R2641 gnd.n4035 gnd.n3629 585
R2642 gnd.n3629 gnd.n3628 585
R2643 gnd.n4037 gnd.n4036 585
R2644 gnd.n4038 gnd.n4037 585
R2645 gnd.n3630 gnd.n3627 585
R2646 gnd.n3636 gnd.n3627 585
R2647 gnd.n4016 gnd.n4015 585
R2648 gnd.n4017 gnd.n4016 585
R2649 gnd.n3647 gnd.n3646 585
R2650 gnd.n3646 gnd.n3642 585
R2651 gnd.n4006 gnd.n4005 585
R2652 gnd.n4007 gnd.n4006 585
R2653 gnd.n3657 gnd.n3656 585
R2654 gnd.n3662 gnd.n3656 585
R2655 gnd.n3984 gnd.n3675 585
R2656 gnd.n3675 gnd.n3661 585
R2657 gnd.n3986 gnd.n3985 585
R2658 gnd.n3987 gnd.n3986 585
R2659 gnd.n3676 gnd.n3674 585
R2660 gnd.n3674 gnd.n3670 585
R2661 gnd.n3975 gnd.n3974 585
R2662 gnd.n3976 gnd.n3975 585
R2663 gnd.n3683 gnd.n3682 585
R2664 gnd.n3687 gnd.n3682 585
R2665 gnd.n3952 gnd.n3704 585
R2666 gnd.n3704 gnd.n3686 585
R2667 gnd.n3954 gnd.n3953 585
R2668 gnd.n3955 gnd.n3954 585
R2669 gnd.n3705 gnd.n3703 585
R2670 gnd.n3703 gnd.n3694 585
R2671 gnd.n3947 gnd.n3946 585
R2672 gnd.n3946 gnd.n3945 585
R2673 gnd.n3752 gnd.n3751 585
R2674 gnd.n3753 gnd.n3752 585
R2675 gnd.n3906 gnd.n3905 585
R2676 gnd.n3907 gnd.n3906 585
R2677 gnd.n3762 gnd.n3761 585
R2678 gnd.n3761 gnd.n3760 585
R2679 gnd.n3901 gnd.n3900 585
R2680 gnd.n3900 gnd.n3899 585
R2681 gnd.n3765 gnd.n3764 585
R2682 gnd.n3766 gnd.n3765 585
R2683 gnd.n3890 gnd.n3889 585
R2684 gnd.n3891 gnd.n3890 585
R2685 gnd.n3773 gnd.n3772 585
R2686 gnd.n3882 gnd.n3772 585
R2687 gnd.n3885 gnd.n3884 585
R2688 gnd.n3884 gnd.n3883 585
R2689 gnd.n3776 gnd.n3775 585
R2690 gnd.n3777 gnd.n3776 585
R2691 gnd.n3871 gnd.n3870 585
R2692 gnd.n3869 gnd.n3795 585
R2693 gnd.n3868 gnd.n3794 585
R2694 gnd.n3873 gnd.n3794 585
R2695 gnd.n3867 gnd.n3866 585
R2696 gnd.n3865 gnd.n3864 585
R2697 gnd.n3863 gnd.n3862 585
R2698 gnd.n3861 gnd.n3860 585
R2699 gnd.n3859 gnd.n3858 585
R2700 gnd.n3857 gnd.n3856 585
R2701 gnd.n3855 gnd.n3854 585
R2702 gnd.n3853 gnd.n3852 585
R2703 gnd.n3851 gnd.n3850 585
R2704 gnd.n3849 gnd.n3848 585
R2705 gnd.n3847 gnd.n3846 585
R2706 gnd.n3845 gnd.n3844 585
R2707 gnd.n3843 gnd.n3842 585
R2708 gnd.n3841 gnd.n3840 585
R2709 gnd.n3839 gnd.n3838 585
R2710 gnd.n3837 gnd.n3836 585
R2711 gnd.n3835 gnd.n3834 585
R2712 gnd.n3833 gnd.n3832 585
R2713 gnd.n3831 gnd.n3830 585
R2714 gnd.n3829 gnd.n3828 585
R2715 gnd.n3827 gnd.n3826 585
R2716 gnd.n3825 gnd.n3824 585
R2717 gnd.n3782 gnd.n3781 585
R2718 gnd.n3876 gnd.n3875 585
R2719 gnd.n4638 gnd.n4637 585
R2720 gnd.n4640 gnd.n4639 585
R2721 gnd.n4642 gnd.n4641 585
R2722 gnd.n4644 gnd.n4643 585
R2723 gnd.n4646 gnd.n4645 585
R2724 gnd.n4648 gnd.n4647 585
R2725 gnd.n4650 gnd.n4649 585
R2726 gnd.n4652 gnd.n4651 585
R2727 gnd.n4654 gnd.n4653 585
R2728 gnd.n4656 gnd.n4655 585
R2729 gnd.n4658 gnd.n4657 585
R2730 gnd.n4660 gnd.n4659 585
R2731 gnd.n4662 gnd.n4661 585
R2732 gnd.n4664 gnd.n4663 585
R2733 gnd.n4666 gnd.n4665 585
R2734 gnd.n4668 gnd.n4667 585
R2735 gnd.n4670 gnd.n4669 585
R2736 gnd.n4672 gnd.n4671 585
R2737 gnd.n4674 gnd.n4673 585
R2738 gnd.n4676 gnd.n4675 585
R2739 gnd.n4678 gnd.n4677 585
R2740 gnd.n4680 gnd.n4679 585
R2741 gnd.n4682 gnd.n4681 585
R2742 gnd.n4684 gnd.n4683 585
R2743 gnd.n4686 gnd.n4685 585
R2744 gnd.n4687 gnd.n1862 585
R2745 gnd.n4688 gnd.n1820 585
R2746 gnd.n4726 gnd.n1820 585
R2747 gnd.n4636 gnd.n1892 585
R2748 gnd.n4636 gnd.n4635 585
R2749 gnd.n4304 gnd.n1891 585
R2750 gnd.n1901 gnd.n1891 585
R2751 gnd.n4306 gnd.n4305 585
R2752 gnd.n4305 gnd.n1900 585
R2753 gnd.n4307 gnd.n3323 585
R2754 gnd.n4611 gnd.n3323 585
R2755 gnd.n4309 gnd.n4308 585
R2756 gnd.n4308 gnd.n1908 585
R2757 gnd.n4310 gnd.n3334 585
R2758 gnd.n4340 gnd.n3334 585
R2759 gnd.n4313 gnd.n4312 585
R2760 gnd.n4312 gnd.n4311 585
R2761 gnd.n4314 gnd.n3341 585
R2762 gnd.n4329 gnd.n3341 585
R2763 gnd.n4316 gnd.n4315 585
R2764 gnd.n4317 gnd.n4316 585
R2765 gnd.n3351 gnd.n3350 585
R2766 gnd.n3358 gnd.n3350 585
R2767 gnd.n4292 gnd.n4291 585
R2768 gnd.n4291 gnd.n4290 585
R2769 gnd.n3354 gnd.n3353 585
R2770 gnd.n3368 gnd.n3354 585
R2771 gnd.n4218 gnd.n4217 585
R2772 gnd.n4217 gnd.n3367 585
R2773 gnd.n4219 gnd.n3377 585
R2774 gnd.n4268 gnd.n3377 585
R2775 gnd.n4221 gnd.n4220 585
R2776 gnd.n4220 gnd.n3375 585
R2777 gnd.n4222 gnd.n3388 585
R2778 gnd.n4251 gnd.n3388 585
R2779 gnd.n4224 gnd.n4223 585
R2780 gnd.n4223 gnd.n3396 585
R2781 gnd.n4225 gnd.n3395 585
R2782 gnd.n4240 gnd.n3395 585
R2783 gnd.n4227 gnd.n4226 585
R2784 gnd.n4228 gnd.n4227 585
R2785 gnd.n3407 gnd.n3406 585
R2786 gnd.n3406 gnd.n3403 585
R2787 gnd.n4207 gnd.n4206 585
R2788 gnd.n4206 gnd.n4205 585
R2789 gnd.n3410 gnd.n3409 585
R2790 gnd.n3423 gnd.n3410 585
R2791 gnd.n4131 gnd.n4130 585
R2792 gnd.n4130 gnd.n3422 585
R2793 gnd.n4132 gnd.n3432 585
R2794 gnd.n4183 gnd.n3432 585
R2795 gnd.n4134 gnd.n4133 585
R2796 gnd.n4133 gnd.n3430 585
R2797 gnd.n4135 gnd.n3443 585
R2798 gnd.n4166 gnd.n3443 585
R2799 gnd.n4137 gnd.n4136 585
R2800 gnd.n4136 gnd.n3450 585
R2801 gnd.n4138 gnd.n3449 585
R2802 gnd.n4155 gnd.n3449 585
R2803 gnd.n4140 gnd.n4139 585
R2804 gnd.n4143 gnd.n4140 585
R2805 gnd.n3460 gnd.n3459 585
R2806 gnd.n3459 gnd.n3457 585
R2807 gnd.n3583 gnd.n3582 585
R2808 gnd.n4098 gnd.n3582 585
R2809 gnd.n3585 gnd.n3584 585
R2810 gnd.n3586 gnd.n3585 585
R2811 gnd.n3596 gnd.n3572 585
R2812 gnd.n4104 gnd.n3572 585
R2813 gnd.n3598 gnd.n3597 585
R2814 gnd.n3599 gnd.n3598 585
R2815 gnd.n3595 gnd.n3594 585
R2816 gnd.n3595 gnd.n3562 585
R2817 gnd.n3593 gnd.n3560 585
R2818 gnd.n4112 gnd.n3560 585
R2819 gnd.n3549 gnd.n3547 585
R2820 gnd.n4074 gnd.n3549 585
R2821 gnd.n4120 gnd.n4119 585
R2822 gnd.n4119 gnd.n4118 585
R2823 gnd.n3548 gnd.n3546 585
R2824 gnd.n3613 gnd.n3548 585
R2825 gnd.n4045 gnd.n3612 585
R2826 gnd.n4064 gnd.n3612 585
R2827 gnd.n4047 gnd.n4046 585
R2828 gnd.n4048 gnd.n4047 585
R2829 gnd.n3622 gnd.n3621 585
R2830 gnd.n3628 gnd.n3621 585
R2831 gnd.n4040 gnd.n4039 585
R2832 gnd.n4039 gnd.n4038 585
R2833 gnd.n3625 gnd.n3624 585
R2834 gnd.n3636 gnd.n3625 585
R2835 gnd.n3925 gnd.n3644 585
R2836 gnd.n4017 gnd.n3644 585
R2837 gnd.n3927 gnd.n3926 585
R2838 gnd.n3926 gnd.n3642 585
R2839 gnd.n3928 gnd.n3655 585
R2840 gnd.n4007 gnd.n3655 585
R2841 gnd.n3930 gnd.n3929 585
R2842 gnd.n3930 gnd.n3662 585
R2843 gnd.n3932 gnd.n3931 585
R2844 gnd.n3931 gnd.n3661 585
R2845 gnd.n3933 gnd.n3672 585
R2846 gnd.n3987 gnd.n3672 585
R2847 gnd.n3935 gnd.n3934 585
R2848 gnd.n3934 gnd.n3670 585
R2849 gnd.n3936 gnd.n3681 585
R2850 gnd.n3976 gnd.n3681 585
R2851 gnd.n3938 gnd.n3937 585
R2852 gnd.n3938 gnd.n3687 585
R2853 gnd.n3940 gnd.n3939 585
R2854 gnd.n3939 gnd.n3686 585
R2855 gnd.n3941 gnd.n3702 585
R2856 gnd.n3955 gnd.n3702 585
R2857 gnd.n3942 gnd.n3755 585
R2858 gnd.n3755 gnd.n3694 585
R2859 gnd.n3944 gnd.n3943 585
R2860 gnd.n3945 gnd.n3944 585
R2861 gnd.n3756 gnd.n3754 585
R2862 gnd.n3754 gnd.n3753 585
R2863 gnd.n3909 gnd.n3908 585
R2864 gnd.n3908 gnd.n3907 585
R2865 gnd.n3759 gnd.n3758 585
R2866 gnd.n3760 gnd.n3759 585
R2867 gnd.n3898 gnd.n3897 585
R2868 gnd.n3899 gnd.n3898 585
R2869 gnd.n3768 gnd.n3767 585
R2870 gnd.n3767 gnd.n3766 585
R2871 gnd.n3893 gnd.n3892 585
R2872 gnd.n3892 gnd.n3891 585
R2873 gnd.n3771 gnd.n3770 585
R2874 gnd.n3882 gnd.n3771 585
R2875 gnd.n3881 gnd.n3880 585
R2876 gnd.n3883 gnd.n3881 585
R2877 gnd.n3779 gnd.n3778 585
R2878 gnd.n3778 gnd.n3777 585
R2879 gnd.n241 gnd.n240 585
R2880 gnd.n244 gnd.n241 585
R2881 gnd.n7670 gnd.n7669 585
R2882 gnd.n7669 gnd.n7668 585
R2883 gnd.n7671 gnd.n236 585
R2884 gnd.n236 gnd.n235 585
R2885 gnd.n7673 gnd.n7672 585
R2886 gnd.n7674 gnd.n7673 585
R2887 gnd.n221 gnd.n220 585
R2888 gnd.n225 gnd.n221 585
R2889 gnd.n7682 gnd.n7681 585
R2890 gnd.n7681 gnd.n7680 585
R2891 gnd.n7683 gnd.n216 585
R2892 gnd.n222 gnd.n216 585
R2893 gnd.n7685 gnd.n7684 585
R2894 gnd.n7686 gnd.n7685 585
R2895 gnd.n203 gnd.n202 585
R2896 gnd.n206 gnd.n203 585
R2897 gnd.n7694 gnd.n7693 585
R2898 gnd.n7693 gnd.n7692 585
R2899 gnd.n7695 gnd.n198 585
R2900 gnd.n198 gnd.n197 585
R2901 gnd.n7697 gnd.n7696 585
R2902 gnd.n7698 gnd.n7697 585
R2903 gnd.n183 gnd.n182 585
R2904 gnd.n194 gnd.n183 585
R2905 gnd.n7706 gnd.n7705 585
R2906 gnd.n7705 gnd.n7704 585
R2907 gnd.n7707 gnd.n178 585
R2908 gnd.n184 gnd.n178 585
R2909 gnd.n7709 gnd.n7708 585
R2910 gnd.n7710 gnd.n7709 585
R2911 gnd.n165 gnd.n164 585
R2912 gnd.n168 gnd.n165 585
R2913 gnd.n7718 gnd.n7717 585
R2914 gnd.n7717 gnd.n7716 585
R2915 gnd.n7719 gnd.n160 585
R2916 gnd.n160 gnd.n159 585
R2917 gnd.n7721 gnd.n7720 585
R2918 gnd.n7722 gnd.n7721 585
R2919 gnd.n145 gnd.n144 585
R2920 gnd.n156 gnd.n145 585
R2921 gnd.n7730 gnd.n7729 585
R2922 gnd.n7729 gnd.n7728 585
R2923 gnd.n7731 gnd.n140 585
R2924 gnd.n146 gnd.n140 585
R2925 gnd.n7733 gnd.n7732 585
R2926 gnd.n7734 gnd.n7733 585
R2927 gnd.n128 gnd.n127 585
R2928 gnd.n131 gnd.n128 585
R2929 gnd.n7742 gnd.n7741 585
R2930 gnd.n7741 gnd.n7740 585
R2931 gnd.n7743 gnd.n122 585
R2932 gnd.n7490 gnd.n122 585
R2933 gnd.n7745 gnd.n7744 585
R2934 gnd.n7746 gnd.n7745 585
R2935 gnd.n123 gnd.n121 585
R2936 gnd.n7360 gnd.n121 585
R2937 gnd.n7355 gnd.n7354 585
R2938 gnd.n7354 gnd.n7353 585
R2939 gnd.n355 gnd.n103 585
R2940 gnd.n7754 gnd.n103 585
R2941 gnd.n7342 gnd.n7341 585
R2942 gnd.n7343 gnd.n7342 585
R2943 gnd.n363 gnd.n362 585
R2944 gnd.n7335 gnd.n362 585
R2945 gnd.n7329 gnd.n7328 585
R2946 gnd.n7330 gnd.n7329 585
R2947 gnd.n374 gnd.n373 585
R2948 gnd.n7323 gnd.n373 585
R2949 gnd.n7304 gnd.n385 585
R2950 gnd.n7312 gnd.n385 585
R2951 gnd.n7306 gnd.n7305 585
R2952 gnd.n7307 gnd.n7306 585
R2953 gnd.n391 gnd.n390 585
R2954 gnd.n7299 gnd.n390 585
R2955 gnd.n7270 gnd.n7269 585
R2956 gnd.n7269 gnd.n7268 585
R2957 gnd.n7271 gnd.n405 585
R2958 gnd.n7285 gnd.n405 585
R2959 gnd.n7272 gnd.n416 585
R2960 gnd.n7262 gnd.n416 585
R2961 gnd.n7274 gnd.n7273 585
R2962 gnd.n7275 gnd.n7274 585
R2963 gnd.n417 gnd.n415 585
R2964 gnd.n7258 gnd.n415 585
R2965 gnd.n7224 gnd.n433 585
R2966 gnd.n7236 gnd.n433 585
R2967 gnd.n7225 gnd.n444 585
R2968 gnd.n444 gnd.n431 585
R2969 gnd.n7227 gnd.n7226 585
R2970 gnd.n7228 gnd.n7227 585
R2971 gnd.n445 gnd.n443 585
R2972 gnd.n7216 gnd.n443 585
R2973 gnd.n7183 gnd.n7182 585
R2974 gnd.n7182 gnd.n7181 585
R2975 gnd.n7184 gnd.n459 585
R2976 gnd.n7198 gnd.n459 585
R2977 gnd.n7185 gnd.n471 585
R2978 gnd.n509 gnd.n471 585
R2979 gnd.n7187 gnd.n7186 585
R2980 gnd.n7188 gnd.n7187 585
R2981 gnd.n472 gnd.n470 585
R2982 gnd.n7144 gnd.n470 585
R2983 gnd.n7149 gnd.n491 585
R2984 gnd.n7161 gnd.n491 585
R2985 gnd.n7150 gnd.n501 585
R2986 gnd.n501 gnd.n487 585
R2987 gnd.n7152 gnd.n7151 585
R2988 gnd.n7153 gnd.n7152 585
R2989 gnd.n502 gnd.n500 585
R2990 gnd.n543 gnd.n500 585
R2991 gnd.n7113 gnd.n7112 585
R2992 gnd.n7112 gnd.n7111 585
R2993 gnd.n7114 gnd.n524 585
R2994 gnd.n7128 gnd.n524 585
R2995 gnd.n7115 gnd.n536 585
R2996 gnd.n7099 gnd.n536 585
R2997 gnd.n7117 gnd.n7116 585
R2998 gnd.n7118 gnd.n7117 585
R2999 gnd.n537 gnd.n535 585
R3000 gnd.n7087 gnd.n535 585
R3001 gnd.n579 gnd.n578 585
R3002 gnd.n578 gnd.n577 585
R3003 gnd.n576 gnd.n563 585
R3004 gnd.n7078 gnd.n563 585
R3005 gnd.n7065 gnd.n574 585
R3006 gnd.n7060 gnd.n574 585
R3007 gnd.n7067 gnd.n7066 585
R3008 gnd.n7068 gnd.n7067 585
R3009 gnd.n704 gnd.n573 585
R3010 gnd.n6918 gnd.n705 585
R3011 gnd.n6917 gnd.n706 585
R3012 gnd.n713 gnd.n707 585
R3013 gnd.n6910 gnd.n714 585
R3014 gnd.n6909 gnd.n715 585
R3015 gnd.n717 gnd.n716 585
R3016 gnd.n6902 gnd.n723 585
R3017 gnd.n6901 gnd.n724 585
R3018 gnd.n731 gnd.n725 585
R3019 gnd.n6894 gnd.n732 585
R3020 gnd.n6893 gnd.n733 585
R3021 gnd.n735 gnd.n734 585
R3022 gnd.n6886 gnd.n741 585
R3023 gnd.n6885 gnd.n742 585
R3024 gnd.n751 gnd.n743 585
R3025 gnd.n6878 gnd.n752 585
R3026 gnd.n6877 gnd.n6874 585
R3027 gnd.n753 gnd.n627 585
R3028 gnd.n7041 gnd.n627 585
R3029 gnd.n7448 gnd.n7447 585
R3030 gnd.n7441 gnd.n7394 585
R3031 gnd.n7443 gnd.n7442 585
R3032 gnd.n7440 gnd.n7439 585
R3033 gnd.n7438 gnd.n7437 585
R3034 gnd.n7431 gnd.n7396 585
R3035 gnd.n7433 gnd.n7432 585
R3036 gnd.n7430 gnd.n7429 585
R3037 gnd.n7428 gnd.n7427 585
R3038 gnd.n7421 gnd.n7398 585
R3039 gnd.n7423 gnd.n7422 585
R3040 gnd.n7420 gnd.n7419 585
R3041 gnd.n7418 gnd.n7417 585
R3042 gnd.n7411 gnd.n7400 585
R3043 gnd.n7413 gnd.n7412 585
R3044 gnd.n7410 gnd.n7409 585
R3045 gnd.n7408 gnd.n7407 585
R3046 gnd.n7404 gnd.n7403 585
R3047 gnd.n7402 gnd.n251 585
R3048 gnd.n7660 gnd.n251 585
R3049 gnd.n7450 gnd.n7449 585
R3050 gnd.n7449 gnd.n244 585
R3051 gnd.n7451 gnd.n243 585
R3052 gnd.n7668 gnd.n243 585
R3053 gnd.n7453 gnd.n7452 585
R3054 gnd.n7452 gnd.n235 585
R3055 gnd.n7454 gnd.n234 585
R3056 gnd.n7674 gnd.n234 585
R3057 gnd.n7456 gnd.n7455 585
R3058 gnd.n7455 gnd.n225 585
R3059 gnd.n7457 gnd.n224 585
R3060 gnd.n7680 gnd.n224 585
R3061 gnd.n7459 gnd.n7458 585
R3062 gnd.n7458 gnd.n222 585
R3063 gnd.n7460 gnd.n215 585
R3064 gnd.n7686 gnd.n215 585
R3065 gnd.n7462 gnd.n7461 585
R3066 gnd.n7461 gnd.n206 585
R3067 gnd.n7463 gnd.n205 585
R3068 gnd.n7692 gnd.n205 585
R3069 gnd.n7465 gnd.n7464 585
R3070 gnd.n7464 gnd.n197 585
R3071 gnd.n7466 gnd.n196 585
R3072 gnd.n7698 gnd.n196 585
R3073 gnd.n7468 gnd.n7467 585
R3074 gnd.n7467 gnd.n194 585
R3075 gnd.n7469 gnd.n186 585
R3076 gnd.n7704 gnd.n186 585
R3077 gnd.n7471 gnd.n7470 585
R3078 gnd.n7470 gnd.n184 585
R3079 gnd.n7472 gnd.n177 585
R3080 gnd.n7710 gnd.n177 585
R3081 gnd.n7474 gnd.n7473 585
R3082 gnd.n7473 gnd.n168 585
R3083 gnd.n7475 gnd.n167 585
R3084 gnd.n7716 gnd.n167 585
R3085 gnd.n7477 gnd.n7476 585
R3086 gnd.n7476 gnd.n159 585
R3087 gnd.n7478 gnd.n158 585
R3088 gnd.n7722 gnd.n158 585
R3089 gnd.n7480 gnd.n7479 585
R3090 gnd.n7479 gnd.n156 585
R3091 gnd.n7481 gnd.n148 585
R3092 gnd.n7728 gnd.n148 585
R3093 gnd.n7483 gnd.n7482 585
R3094 gnd.n7482 gnd.n146 585
R3095 gnd.n7484 gnd.n139 585
R3096 gnd.n7734 gnd.n139 585
R3097 gnd.n7486 gnd.n7485 585
R3098 gnd.n7485 gnd.n131 585
R3099 gnd.n7487 gnd.n130 585
R3100 gnd.n7740 gnd.n130 585
R3101 gnd.n7489 gnd.n7488 585
R3102 gnd.n7490 gnd.n7489 585
R3103 gnd.n350 gnd.n119 585
R3104 gnd.n7746 gnd.n119 585
R3105 gnd.n7362 gnd.n7361 585
R3106 gnd.n7361 gnd.n7360 585
R3107 gnd.n100 gnd.n99 585
R3108 gnd.n7353 gnd.n100 585
R3109 gnd.n7756 gnd.n7755 585
R3110 gnd.n7755 gnd.n7754 585
R3111 gnd.n7757 gnd.n98 585
R3112 gnd.n7343 gnd.n98 585
R3113 gnd.n368 gnd.n96 585
R3114 gnd.n7335 gnd.n368 585
R3115 gnd.n7291 gnd.n372 585
R3116 gnd.n7330 gnd.n372 585
R3117 gnd.n7292 gnd.n379 585
R3118 gnd.n7323 gnd.n379 585
R3119 gnd.n7293 gnd.n384 585
R3120 gnd.n7312 gnd.n384 585
R3121 gnd.n398 gnd.n389 585
R3122 gnd.n7307 gnd.n389 585
R3123 gnd.n7298 gnd.n7297 585
R3124 gnd.n7299 gnd.n7298 585
R3125 gnd.n397 gnd.n396 585
R3126 gnd.n7268 gnd.n396 585
R3127 gnd.n7287 gnd.n7286 585
R3128 gnd.n7286 gnd.n7285 585
R3129 gnd.n401 gnd.n400 585
R3130 gnd.n7262 gnd.n401 585
R3131 gnd.n7205 gnd.n413 585
R3132 gnd.n7275 gnd.n413 585
R3133 gnd.n7208 gnd.n424 585
R3134 gnd.n7258 gnd.n424 585
R3135 gnd.n7209 gnd.n432 585
R3136 gnd.n7236 gnd.n432 585
R3137 gnd.n7210 gnd.n7204 585
R3138 gnd.n7204 gnd.n431 585
R3139 gnd.n452 gnd.n441 585
R3140 gnd.n7228 gnd.n441 585
R3141 gnd.n7215 gnd.n7214 585
R3142 gnd.n7216 gnd.n7215 585
R3143 gnd.n451 gnd.n450 585
R3144 gnd.n7181 gnd.n450 585
R3145 gnd.n7200 gnd.n7199 585
R3146 gnd.n7199 gnd.n7198 585
R3147 gnd.n455 gnd.n454 585
R3148 gnd.n509 gnd.n455 585
R3149 gnd.n514 gnd.n468 585
R3150 gnd.n7188 gnd.n468 585
R3151 gnd.n7143 gnd.n7142 585
R3152 gnd.n7144 gnd.n7143 585
R3153 gnd.n513 gnd.n489 585
R3154 gnd.n7161 gnd.n489 585
R3155 gnd.n7137 gnd.n7136 585
R3156 gnd.n7136 gnd.n487 585
R3157 gnd.n7135 gnd.n498 585
R3158 gnd.n7153 gnd.n498 585
R3159 gnd.n7134 gnd.n517 585
R3160 gnd.n543 gnd.n517 585
R3161 gnd.n521 gnd.n516 585
R3162 gnd.n7111 gnd.n521 585
R3163 gnd.n7130 gnd.n7129 585
R3164 gnd.n7129 gnd.n7128 585
R3165 gnd.n520 gnd.n519 585
R3166 gnd.n7099 gnd.n520 585
R3167 gnd.n557 gnd.n533 585
R3168 gnd.n7118 gnd.n533 585
R3169 gnd.n7086 gnd.n7085 585
R3170 gnd.n7087 gnd.n7086 585
R3171 gnd.n556 gnd.n555 585
R3172 gnd.n577 gnd.n555 585
R3173 gnd.n7080 gnd.n7079 585
R3174 gnd.n7079 gnd.n7078 585
R3175 gnd.n560 gnd.n559 585
R3176 gnd.n7060 gnd.n560 585
R3177 gnd.n6866 gnd.n571 585
R3178 gnd.n7068 gnd.n571 585
R3179 gnd.n4621 gnd.n1842 585
R3180 gnd.n1842 gnd.n1819 585
R3181 gnd.n4622 gnd.n1903 585
R3182 gnd.n1903 gnd.n1893 585
R3183 gnd.n4624 gnd.n4623 585
R3184 gnd.n4625 gnd.n4624 585
R3185 gnd.n1904 gnd.n1902 585
R3186 gnd.n3324 gnd.n1902 585
R3187 gnd.n4615 gnd.n4614 585
R3188 gnd.n4614 gnd.n4613 585
R3189 gnd.n1907 gnd.n1906 585
R3190 gnd.n4339 gnd.n1907 585
R3191 gnd.n4325 gnd.n3343 585
R3192 gnd.n3343 gnd.n3333 585
R3193 gnd.n4327 gnd.n4326 585
R3194 gnd.n4328 gnd.n4327 585
R3195 gnd.n3344 gnd.n3342 585
R3196 gnd.n3342 gnd.n3340 585
R3197 gnd.n4320 gnd.n4319 585
R3198 gnd.n4319 gnd.n4318 585
R3199 gnd.n3347 gnd.n3346 585
R3200 gnd.n3356 gnd.n3347 585
R3201 gnd.n4276 gnd.n3370 585
R3202 gnd.n3370 gnd.n3355 585
R3203 gnd.n4278 gnd.n4277 585
R3204 gnd.n4279 gnd.n4278 585
R3205 gnd.n3371 gnd.n3369 585
R3206 gnd.n3378 gnd.n3369 585
R3207 gnd.n4271 gnd.n4270 585
R3208 gnd.n4270 gnd.n4269 585
R3209 gnd.n3374 gnd.n3373 585
R3210 gnd.n4250 gnd.n3374 585
R3211 gnd.n4236 gnd.n3398 585
R3212 gnd.n3398 gnd.n3387 585
R3213 gnd.n4238 gnd.n4237 585
R3214 gnd.n4239 gnd.n4238 585
R3215 gnd.n3399 gnd.n3397 585
R3216 gnd.n3397 gnd.n3394 585
R3217 gnd.n4231 gnd.n4230 585
R3218 gnd.n4230 gnd.n4229 585
R3219 gnd.n3402 gnd.n3401 585
R3220 gnd.n3412 gnd.n3402 585
R3221 gnd.n4191 gnd.n3425 585
R3222 gnd.n3425 gnd.n3411 585
R3223 gnd.n4193 gnd.n4192 585
R3224 gnd.n4194 gnd.n4193 585
R3225 gnd.n3426 gnd.n3424 585
R3226 gnd.n3433 gnd.n3424 585
R3227 gnd.n4186 gnd.n4185 585
R3228 gnd.n4185 gnd.n4184 585
R3229 gnd.n3429 gnd.n3428 585
R3230 gnd.n4165 gnd.n3429 585
R3231 gnd.n4151 gnd.n3452 585
R3232 gnd.n3452 gnd.n3442 585
R3233 gnd.n4153 gnd.n4152 585
R3234 gnd.n4154 gnd.n4153 585
R3235 gnd.n3453 gnd.n3451 585
R3236 gnd.n4142 gnd.n3451 585
R3237 gnd.n4146 gnd.n4145 585
R3238 gnd.n4145 gnd.n4144 585
R3239 gnd.n3456 gnd.n3455 585
R3240 gnd.n4097 gnd.n3456 585
R3241 gnd.n3590 gnd.n3589 585
R3242 gnd.n3591 gnd.n3590 585
R3243 gnd.n3570 gnd.n3569 585
R3244 gnd.n3573 gnd.n3570 585
R3245 gnd.n4107 gnd.n4106 585
R3246 gnd.n4106 gnd.n4105 585
R3247 gnd.n4108 gnd.n3564 585
R3248 gnd.n3600 gnd.n3564 585
R3249 gnd.n4110 gnd.n4109 585
R3250 gnd.n4111 gnd.n4110 585
R3251 gnd.n3565 gnd.n3563 585
R3252 gnd.n4075 gnd.n3563 585
R3253 gnd.n4059 gnd.n4058 585
R3254 gnd.n4058 gnd.n3551 585
R3255 gnd.n4060 gnd.n3615 585
R3256 gnd.n3615 gnd.n3550 585
R3257 gnd.n4062 gnd.n4061 585
R3258 gnd.n4063 gnd.n4062 585
R3259 gnd.n3616 gnd.n3614 585
R3260 gnd.n3614 gnd.n3611 585
R3261 gnd.n4051 gnd.n4050 585
R3262 gnd.n4050 gnd.n4049 585
R3263 gnd.n3619 gnd.n3618 585
R3264 gnd.n3626 gnd.n3619 585
R3265 gnd.n4025 gnd.n4024 585
R3266 gnd.n4026 gnd.n4025 585
R3267 gnd.n3638 gnd.n3637 585
R3268 gnd.n3645 gnd.n3637 585
R3269 gnd.n4020 gnd.n4019 585
R3270 gnd.n4019 gnd.n4018 585
R3271 gnd.n3641 gnd.n3640 585
R3272 gnd.n4008 gnd.n3641 585
R3273 gnd.n3995 gnd.n3665 585
R3274 gnd.n3665 gnd.n3664 585
R3275 gnd.n3997 gnd.n3996 585
R3276 gnd.n3998 gnd.n3997 585
R3277 gnd.n3666 gnd.n3663 585
R3278 gnd.n3673 gnd.n3663 585
R3279 gnd.n3990 gnd.n3989 585
R3280 gnd.n3989 gnd.n3988 585
R3281 gnd.n3669 gnd.n3668 585
R3282 gnd.n3977 gnd.n3669 585
R3283 gnd.n3964 gnd.n3690 585
R3284 gnd.n3690 gnd.n3689 585
R3285 gnd.n3966 gnd.n3965 585
R3286 gnd.n3967 gnd.n3966 585
R3287 gnd.n3960 gnd.n3688 585
R3288 gnd.n3959 gnd.n3958 585
R3289 gnd.n3693 gnd.n3692 585
R3290 gnd.n3956 gnd.n3693 585
R3291 gnd.n3715 gnd.n3714 585
R3292 gnd.n3718 gnd.n3717 585
R3293 gnd.n3716 gnd.n3711 585
R3294 gnd.n3723 gnd.n3722 585
R3295 gnd.n3725 gnd.n3724 585
R3296 gnd.n3728 gnd.n3727 585
R3297 gnd.n3726 gnd.n3709 585
R3298 gnd.n3733 gnd.n3732 585
R3299 gnd.n3735 gnd.n3734 585
R3300 gnd.n3738 gnd.n3737 585
R3301 gnd.n3736 gnd.n3707 585
R3302 gnd.n3743 gnd.n3742 585
R3303 gnd.n3747 gnd.n3744 585
R3304 gnd.n3748 gnd.n3685 585
R3305 gnd.n4627 gnd.n1857 585
R3306 gnd.n4694 gnd.n4693 585
R3307 gnd.n4696 gnd.n4695 585
R3308 gnd.n4698 gnd.n4697 585
R3309 gnd.n4700 gnd.n4699 585
R3310 gnd.n4702 gnd.n4701 585
R3311 gnd.n4704 gnd.n4703 585
R3312 gnd.n4706 gnd.n4705 585
R3313 gnd.n4708 gnd.n4707 585
R3314 gnd.n4710 gnd.n4709 585
R3315 gnd.n4712 gnd.n4711 585
R3316 gnd.n4714 gnd.n4713 585
R3317 gnd.n4716 gnd.n4715 585
R3318 gnd.n4719 gnd.n4718 585
R3319 gnd.n4717 gnd.n1845 585
R3320 gnd.n4723 gnd.n1843 585
R3321 gnd.n4725 gnd.n4724 585
R3322 gnd.n4726 gnd.n4725 585
R3323 gnd.n4628 gnd.n1898 585
R3324 gnd.n4628 gnd.n1819 585
R3325 gnd.n4630 gnd.n4629 585
R3326 gnd.n4629 gnd.n1893 585
R3327 gnd.n4626 gnd.n1897 585
R3328 gnd.n4626 gnd.n4625 585
R3329 gnd.n4604 gnd.n1899 585
R3330 gnd.n3324 gnd.n1899 585
R3331 gnd.n4603 gnd.n1909 585
R3332 gnd.n4613 gnd.n1909 585
R3333 gnd.n4338 gnd.n3329 585
R3334 gnd.n4339 gnd.n4338 585
R3335 gnd.n4337 gnd.n4336 585
R3336 gnd.n4337 gnd.n3333 585
R3337 gnd.n4335 gnd.n3335 585
R3338 gnd.n4328 gnd.n3335 585
R3339 gnd.n3348 gnd.n3336 585
R3340 gnd.n3348 gnd.n3340 585
R3341 gnd.n4284 gnd.n3349 585
R3342 gnd.n4318 gnd.n3349 585
R3343 gnd.n4283 gnd.n4282 585
R3344 gnd.n4282 gnd.n3356 585
R3345 gnd.n4281 gnd.n3364 585
R3346 gnd.n4281 gnd.n3355 585
R3347 gnd.n4280 gnd.n3366 585
R3348 gnd.n4280 gnd.n4279 585
R3349 gnd.n4259 gnd.n3365 585
R3350 gnd.n3378 gnd.n3365 585
R3351 gnd.n4258 gnd.n3376 585
R3352 gnd.n4269 gnd.n3376 585
R3353 gnd.n4249 gnd.n3383 585
R3354 gnd.n4250 gnd.n4249 585
R3355 gnd.n4248 gnd.n4247 585
R3356 gnd.n4248 gnd.n3387 585
R3357 gnd.n4246 gnd.n3389 585
R3358 gnd.n4239 gnd.n3389 585
R3359 gnd.n3404 gnd.n3390 585
R3360 gnd.n3404 gnd.n3394 585
R3361 gnd.n4199 gnd.n3405 585
R3362 gnd.n4229 gnd.n3405 585
R3363 gnd.n4198 gnd.n4197 585
R3364 gnd.n4197 gnd.n3412 585
R3365 gnd.n4196 gnd.n3419 585
R3366 gnd.n4196 gnd.n3411 585
R3367 gnd.n4195 gnd.n3421 585
R3368 gnd.n4195 gnd.n4194 585
R3369 gnd.n4174 gnd.n3420 585
R3370 gnd.n3433 gnd.n3420 585
R3371 gnd.n4173 gnd.n3431 585
R3372 gnd.n4184 gnd.n3431 585
R3373 gnd.n4164 gnd.n3438 585
R3374 gnd.n4165 gnd.n4164 585
R3375 gnd.n4163 gnd.n4162 585
R3376 gnd.n4163 gnd.n3442 585
R3377 gnd.n4161 gnd.n3444 585
R3378 gnd.n4154 gnd.n3444 585
R3379 gnd.n4141 gnd.n3445 585
R3380 gnd.n4142 gnd.n4141 585
R3381 gnd.n4094 gnd.n3458 585
R3382 gnd.n4144 gnd.n3458 585
R3383 gnd.n4096 gnd.n4095 585
R3384 gnd.n4097 gnd.n4096 585
R3385 gnd.n4089 gnd.n3592 585
R3386 gnd.n3592 gnd.n3591 585
R3387 gnd.n4087 gnd.n4086 585
R3388 gnd.n4086 gnd.n3573 585
R3389 gnd.n4084 gnd.n3571 585
R3390 gnd.n4105 gnd.n3571 585
R3391 gnd.n3602 gnd.n3601 585
R3392 gnd.n3601 gnd.n3600 585
R3393 gnd.n4078 gnd.n3561 585
R3394 gnd.n4111 gnd.n3561 585
R3395 gnd.n4077 gnd.n4076 585
R3396 gnd.n4076 gnd.n4075 585
R3397 gnd.n4073 gnd.n3604 585
R3398 gnd.n4073 gnd.n3551 585
R3399 gnd.n4072 gnd.n4071 585
R3400 gnd.n4072 gnd.n3550 585
R3401 gnd.n3607 gnd.n3606 585
R3402 gnd.n4063 gnd.n3606 585
R3403 gnd.n4031 gnd.n4030 585
R3404 gnd.n4030 gnd.n3611 585
R3405 gnd.n4032 gnd.n3620 585
R3406 gnd.n4049 gnd.n3620 585
R3407 gnd.n4029 gnd.n4028 585
R3408 gnd.n4028 gnd.n3626 585
R3409 gnd.n4027 gnd.n3634 585
R3410 gnd.n4027 gnd.n4026 585
R3411 gnd.n4012 gnd.n3635 585
R3412 gnd.n3645 gnd.n3635 585
R3413 gnd.n4011 gnd.n3643 585
R3414 gnd.n4018 gnd.n3643 585
R3415 gnd.n4010 gnd.n4009 585
R3416 gnd.n4009 gnd.n4008 585
R3417 gnd.n3654 gnd.n3651 585
R3418 gnd.n3664 gnd.n3654 585
R3419 gnd.n4000 gnd.n3999 585
R3420 gnd.n3999 gnd.n3998 585
R3421 gnd.n3660 gnd.n3659 585
R3422 gnd.n3673 gnd.n3660 585
R3423 gnd.n3980 gnd.n3671 585
R3424 gnd.n3988 gnd.n3671 585
R3425 gnd.n3979 gnd.n3978 585
R3426 gnd.n3978 gnd.n3977 585
R3427 gnd.n3680 gnd.n3678 585
R3428 gnd.n3689 gnd.n3680 585
R3429 gnd.n3969 gnd.n3968 585
R3430 gnd.n3968 gnd.n3967 585
R3431 gnd.n6640 gnd.n935 585
R3432 gnd.n935 gnd.n891 585
R3433 gnd.n6642 gnd.n6641 585
R3434 gnd.n6643 gnd.n6642 585
R3435 gnd.n6551 gnd.n934 585
R3436 gnd.n6518 gnd.n934 585
R3437 gnd.n6550 gnd.n6549 585
R3438 gnd.n6549 gnd.n6548 585
R3439 gnd.n937 gnd.n936 585
R3440 gnd.n6471 gnd.n937 585
R3441 gnd.n6537 gnd.n6536 585
R3442 gnd.n6538 gnd.n6537 585
R3443 gnd.n6535 gnd.n949 585
R3444 gnd.n949 gnd.n945 585
R3445 gnd.n6534 gnd.n6533 585
R3446 gnd.n6533 gnd.n6532 585
R3447 gnd.n951 gnd.n950 585
R3448 gnd.n6481 gnd.n951 585
R3449 gnd.n6461 gnd.n997 585
R3450 gnd.n997 gnd.n991 585
R3451 gnd.n6463 gnd.n6462 585
R3452 gnd.n6464 gnd.n6463 585
R3453 gnd.n6460 gnd.n996 585
R3454 gnd.n996 gnd.n972 585
R3455 gnd.n6459 gnd.n6458 585
R3456 gnd.n6458 gnd.n6457 585
R3457 gnd.n999 gnd.n998 585
R3458 gnd.n1001 gnd.n999 585
R3459 gnd.n6446 gnd.n1008 585
R3460 gnd.n1008 gnd.n981 585
R3461 gnd.n6448 gnd.n6447 585
R3462 gnd.n6449 gnd.n6448 585
R3463 gnd.n6445 gnd.n1007 585
R3464 gnd.n1013 gnd.n1007 585
R3465 gnd.n6444 gnd.n6443 585
R3466 gnd.n6443 gnd.n6442 585
R3467 gnd.n1010 gnd.n1009 585
R3468 gnd.n6418 gnd.n1010 585
R3469 gnd.n6431 gnd.n6430 585
R3470 gnd.n6432 gnd.n6431 585
R3471 gnd.n6429 gnd.n1023 585
R3472 gnd.n1028 gnd.n1023 585
R3473 gnd.n6428 gnd.n6427 585
R3474 gnd.n6427 gnd.n6426 585
R3475 gnd.n1025 gnd.n1024 585
R3476 gnd.n6407 gnd.n1025 585
R3477 gnd.n6392 gnd.n6391 585
R3478 gnd.n6391 gnd.n1042 585
R3479 gnd.n6393 gnd.n1054 585
R3480 gnd.n6379 gnd.n1054 585
R3481 gnd.n6395 gnd.n6394 585
R3482 gnd.n6396 gnd.n6395 585
R3483 gnd.n6390 gnd.n1053 585
R3484 gnd.n1053 gnd.n1049 585
R3485 gnd.n6389 gnd.n6388 585
R3486 gnd.n6388 gnd.n6387 585
R3487 gnd.n1056 gnd.n1055 585
R3488 gnd.n6370 gnd.n1056 585
R3489 gnd.n6355 gnd.n6354 585
R3490 gnd.n6354 gnd.n1069 585
R3491 gnd.n6356 gnd.n1081 585
R3492 gnd.n6341 gnd.n1081 585
R3493 gnd.n6358 gnd.n6357 585
R3494 gnd.n6359 gnd.n6358 585
R3495 gnd.n6353 gnd.n1080 585
R3496 gnd.n1080 gnd.n1076 585
R3497 gnd.n6352 gnd.n6351 585
R3498 gnd.n6351 gnd.n6350 585
R3499 gnd.n1083 gnd.n1082 585
R3500 gnd.n1101 gnd.n1083 585
R3501 gnd.n6293 gnd.n6292 585
R3502 gnd.n6292 gnd.n1099 585
R3503 gnd.n6294 gnd.n1111 585
R3504 gnd.n6278 gnd.n1111 585
R3505 gnd.n6296 gnd.n6295 585
R3506 gnd.n6297 gnd.n6296 585
R3507 gnd.n6291 gnd.n1110 585
R3508 gnd.n1117 gnd.n1110 585
R3509 gnd.n6290 gnd.n6289 585
R3510 gnd.n6289 gnd.n6288 585
R3511 gnd.n1113 gnd.n1112 585
R3512 gnd.n6261 gnd.n1113 585
R3513 gnd.n6247 gnd.n6246 585
R3514 gnd.n6246 gnd.n1128 585
R3515 gnd.n6248 gnd.n1139 585
R3516 gnd.n6234 gnd.n1139 585
R3517 gnd.n6250 gnd.n6249 585
R3518 gnd.n6251 gnd.n6250 585
R3519 gnd.n6245 gnd.n1138 585
R3520 gnd.n6240 gnd.n1138 585
R3521 gnd.n6244 gnd.n6243 585
R3522 gnd.n6243 gnd.n6242 585
R3523 gnd.n1141 gnd.n1140 585
R3524 gnd.n6221 gnd.n1141 585
R3525 gnd.n6212 gnd.n1161 585
R3526 gnd.n1161 gnd.n1160 585
R3527 gnd.n6214 gnd.n6213 585
R3528 gnd.n6215 gnd.n6214 585
R3529 gnd.n6211 gnd.n1158 585
R3530 gnd.n1166 gnd.n1158 585
R3531 gnd.n6210 gnd.n6209 585
R3532 gnd.n6209 gnd.n6208 585
R3533 gnd.n1163 gnd.n1162 585
R3534 gnd.n1206 gnd.n1163 585
R3535 gnd.n6170 gnd.n6169 585
R3536 gnd.n6170 gnd.n1176 585
R3537 gnd.n6172 gnd.n6171 585
R3538 gnd.n6171 gnd.n1174 585
R3539 gnd.n6173 gnd.n1188 585
R3540 gnd.n6146 gnd.n1188 585
R3541 gnd.n6175 gnd.n6174 585
R3542 gnd.n6176 gnd.n6175 585
R3543 gnd.n6168 gnd.n1187 585
R3544 gnd.n6163 gnd.n1187 585
R3545 gnd.n6167 gnd.n6166 585
R3546 gnd.n6166 gnd.n6165 585
R3547 gnd.n1190 gnd.n1189 585
R3548 gnd.t87 gnd.n1190 585
R3549 gnd.n1287 gnd.n1286 585
R3550 gnd.n1286 gnd.n1200 585
R3551 gnd.n1288 gnd.n1265 585
R3552 gnd.n1265 gnd.n1218 585
R3553 gnd.n6097 gnd.n6096 585
R3554 gnd.n6095 gnd.n1264 585
R3555 gnd.n6094 gnd.n1263 585
R3556 gnd.n6099 gnd.n1263 585
R3557 gnd.n6093 gnd.n6092 585
R3558 gnd.n6091 gnd.n6090 585
R3559 gnd.n6089 gnd.n6088 585
R3560 gnd.n6087 gnd.n6086 585
R3561 gnd.n6085 gnd.n6084 585
R3562 gnd.n6083 gnd.n6082 585
R3563 gnd.n6081 gnd.n6080 585
R3564 gnd.n6079 gnd.n6078 585
R3565 gnd.n6077 gnd.n6076 585
R3566 gnd.n6075 gnd.n6074 585
R3567 gnd.n6073 gnd.n6072 585
R3568 gnd.n6071 gnd.n6070 585
R3569 gnd.n6069 gnd.n6068 585
R3570 gnd.n6067 gnd.n6066 585
R3571 gnd.n6065 gnd.n6064 585
R3572 gnd.n6063 gnd.n6062 585
R3573 gnd.n6061 gnd.n6060 585
R3574 gnd.n6059 gnd.n6058 585
R3575 gnd.n6057 gnd.n6056 585
R3576 gnd.n6055 gnd.n6054 585
R3577 gnd.n6053 gnd.n6052 585
R3578 gnd.n6051 gnd.n6050 585
R3579 gnd.n6049 gnd.n6048 585
R3580 gnd.n6047 gnd.n6046 585
R3581 gnd.n6045 gnd.n6044 585
R3582 gnd.n6043 gnd.n6042 585
R3583 gnd.n6041 gnd.n6040 585
R3584 gnd.n6039 gnd.n6038 585
R3585 gnd.n6037 gnd.n6036 585
R3586 gnd.n6035 gnd.n6034 585
R3587 gnd.n6033 gnd.n1360 585
R3588 gnd.n1359 gnd.n1358 585
R3589 gnd.n1357 gnd.n1356 585
R3590 gnd.n1354 gnd.n1353 585
R3591 gnd.n1352 gnd.n1351 585
R3592 gnd.n1350 gnd.n1349 585
R3593 gnd.n1348 gnd.n1347 585
R3594 gnd.n1346 gnd.n1345 585
R3595 gnd.n1344 gnd.n1343 585
R3596 gnd.n1342 gnd.n1341 585
R3597 gnd.n1340 gnd.n1339 585
R3598 gnd.n1338 gnd.n1337 585
R3599 gnd.n1336 gnd.n1335 585
R3600 gnd.n1334 gnd.n1333 585
R3601 gnd.n1332 gnd.n1331 585
R3602 gnd.n1330 gnd.n1329 585
R3603 gnd.n1328 gnd.n1327 585
R3604 gnd.n1326 gnd.n1325 585
R3605 gnd.n1324 gnd.n1323 585
R3606 gnd.n1322 gnd.n1321 585
R3607 gnd.n1320 gnd.n1319 585
R3608 gnd.n1318 gnd.n1317 585
R3609 gnd.n1316 gnd.n1315 585
R3610 gnd.n1314 gnd.n1313 585
R3611 gnd.n1312 gnd.n1311 585
R3612 gnd.n1310 gnd.n1309 585
R3613 gnd.n1308 gnd.n1307 585
R3614 gnd.n1306 gnd.n1305 585
R3615 gnd.n1304 gnd.n1303 585
R3616 gnd.n1302 gnd.n1301 585
R3617 gnd.n1300 gnd.n1299 585
R3618 gnd.n1298 gnd.n1297 585
R3619 gnd.n6647 gnd.n6646 585
R3620 gnd.n6649 gnd.n6648 585
R3621 gnd.n6651 gnd.n6650 585
R3622 gnd.n6653 gnd.n6652 585
R3623 gnd.n6655 gnd.n6654 585
R3624 gnd.n6657 gnd.n6656 585
R3625 gnd.n6659 gnd.n6658 585
R3626 gnd.n6661 gnd.n6660 585
R3627 gnd.n6663 gnd.n6662 585
R3628 gnd.n6665 gnd.n6664 585
R3629 gnd.n6667 gnd.n6666 585
R3630 gnd.n6669 gnd.n6668 585
R3631 gnd.n6671 gnd.n6670 585
R3632 gnd.n6673 gnd.n6672 585
R3633 gnd.n6675 gnd.n6674 585
R3634 gnd.n6677 gnd.n6676 585
R3635 gnd.n6679 gnd.n6678 585
R3636 gnd.n6681 gnd.n6680 585
R3637 gnd.n6683 gnd.n6682 585
R3638 gnd.n6685 gnd.n6684 585
R3639 gnd.n6687 gnd.n6686 585
R3640 gnd.n6689 gnd.n6688 585
R3641 gnd.n6691 gnd.n6690 585
R3642 gnd.n6693 gnd.n6692 585
R3643 gnd.n6695 gnd.n6694 585
R3644 gnd.n6697 gnd.n6696 585
R3645 gnd.n6699 gnd.n6698 585
R3646 gnd.n6701 gnd.n6700 585
R3647 gnd.n6703 gnd.n6702 585
R3648 gnd.n6706 gnd.n6705 585
R3649 gnd.n6708 gnd.n6707 585
R3650 gnd.n6710 gnd.n6709 585
R3651 gnd.n6712 gnd.n6711 585
R3652 gnd.n6573 gnd.n657 585
R3653 gnd.n6575 gnd.n6574 585
R3654 gnd.n6577 gnd.n6576 585
R3655 gnd.n6579 gnd.n6578 585
R3656 gnd.n6582 gnd.n6581 585
R3657 gnd.n6584 gnd.n6583 585
R3658 gnd.n6586 gnd.n6585 585
R3659 gnd.n6588 gnd.n6587 585
R3660 gnd.n6590 gnd.n6589 585
R3661 gnd.n6592 gnd.n6591 585
R3662 gnd.n6594 gnd.n6593 585
R3663 gnd.n6596 gnd.n6595 585
R3664 gnd.n6598 gnd.n6597 585
R3665 gnd.n6600 gnd.n6599 585
R3666 gnd.n6602 gnd.n6601 585
R3667 gnd.n6604 gnd.n6603 585
R3668 gnd.n6606 gnd.n6605 585
R3669 gnd.n6608 gnd.n6607 585
R3670 gnd.n6610 gnd.n6609 585
R3671 gnd.n6612 gnd.n6611 585
R3672 gnd.n6614 gnd.n6613 585
R3673 gnd.n6616 gnd.n6615 585
R3674 gnd.n6618 gnd.n6617 585
R3675 gnd.n6620 gnd.n6619 585
R3676 gnd.n6622 gnd.n6621 585
R3677 gnd.n6624 gnd.n6623 585
R3678 gnd.n6626 gnd.n6625 585
R3679 gnd.n6628 gnd.n6627 585
R3680 gnd.n6630 gnd.n6629 585
R3681 gnd.n6632 gnd.n6631 585
R3682 gnd.n6634 gnd.n6633 585
R3683 gnd.n6636 gnd.n6635 585
R3684 gnd.n6638 gnd.n6637 585
R3685 gnd.n6645 gnd.n929 585
R3686 gnd.n6645 gnd.n891 585
R3687 gnd.n6644 gnd.n931 585
R3688 gnd.n6644 gnd.n6643 585
R3689 gnd.n6468 gnd.n930 585
R3690 gnd.n6518 gnd.n930 585
R3691 gnd.n6469 gnd.n939 585
R3692 gnd.n6548 gnd.n939 585
R3693 gnd.n6473 gnd.n6472 585
R3694 gnd.n6472 gnd.n6471 585
R3695 gnd.n6474 gnd.n946 585
R3696 gnd.n6538 gnd.n946 585
R3697 gnd.n6476 gnd.n6475 585
R3698 gnd.n6475 gnd.n945 585
R3699 gnd.n6477 gnd.n953 585
R3700 gnd.n6532 gnd.n953 585
R3701 gnd.n6479 gnd.n6478 585
R3702 gnd.n6481 gnd.n6479 585
R3703 gnd.n6467 gnd.n992 585
R3704 gnd.n992 gnd.n991 585
R3705 gnd.n6466 gnd.n6465 585
R3706 gnd.n6465 gnd.n6464 585
R3707 gnd.n994 gnd.n993 585
R3708 gnd.n994 gnd.n972 585
R3709 gnd.n6455 gnd.n6454 585
R3710 gnd.n6457 gnd.n6455 585
R3711 gnd.n6453 gnd.n1002 585
R3712 gnd.n1002 gnd.n1001 585
R3713 gnd.n6452 gnd.n6451 585
R3714 gnd.n6451 gnd.n981 585
R3715 gnd.n6450 gnd.n1003 585
R3716 gnd.n6450 gnd.n6449 585
R3717 gnd.n6414 gnd.n1004 585
R3718 gnd.n1013 gnd.n1004 585
R3719 gnd.n6415 gnd.n1011 585
R3720 gnd.n6442 gnd.n1011 585
R3721 gnd.n6417 gnd.n6416 585
R3722 gnd.n6418 gnd.n6417 585
R3723 gnd.n6413 gnd.n1021 585
R3724 gnd.n6432 gnd.n1021 585
R3725 gnd.n6412 gnd.n6411 585
R3726 gnd.n6411 gnd.n1028 585
R3727 gnd.n6410 gnd.n1027 585
R3728 gnd.n6426 gnd.n1027 585
R3729 gnd.n6409 gnd.n6408 585
R3730 gnd.n6408 gnd.n6407 585
R3731 gnd.n1041 gnd.n1040 585
R3732 gnd.n1042 gnd.n1041 585
R3733 gnd.n6378 gnd.n6377 585
R3734 gnd.n6379 gnd.n6378 585
R3735 gnd.n6376 gnd.n1051 585
R3736 gnd.n6396 gnd.n1051 585
R3737 gnd.n6375 gnd.n6374 585
R3738 gnd.n6374 gnd.n1049 585
R3739 gnd.n6373 gnd.n1058 585
R3740 gnd.n6387 gnd.n1058 585
R3741 gnd.n6372 gnd.n6371 585
R3742 gnd.n6371 gnd.n6370 585
R3743 gnd.n1068 gnd.n1067 585
R3744 gnd.n1069 gnd.n1068 585
R3745 gnd.n6268 gnd.n1093 585
R3746 gnd.n6341 gnd.n1093 585
R3747 gnd.n6269 gnd.n1078 585
R3748 gnd.n6359 gnd.n1078 585
R3749 gnd.n6271 gnd.n6270 585
R3750 gnd.n6270 gnd.n1076 585
R3751 gnd.n6272 gnd.n1084 585
R3752 gnd.n6350 gnd.n1084 585
R3753 gnd.n6274 gnd.n6273 585
R3754 gnd.n6273 gnd.n1101 585
R3755 gnd.n6275 gnd.n1125 585
R3756 gnd.n1125 gnd.n1099 585
R3757 gnd.n6277 gnd.n6276 585
R3758 gnd.n6278 gnd.n6277 585
R3759 gnd.n6267 gnd.n1108 585
R3760 gnd.n6297 gnd.n1108 585
R3761 gnd.n6266 gnd.n6265 585
R3762 gnd.n6265 gnd.n1117 585
R3763 gnd.n6264 gnd.n1115 585
R3764 gnd.n6288 gnd.n1115 585
R3765 gnd.n6263 gnd.n6262 585
R3766 gnd.n6262 gnd.n6261 585
R3767 gnd.n1127 gnd.n1126 585
R3768 gnd.n1128 gnd.n1127 585
R3769 gnd.n6236 gnd.n6235 585
R3770 gnd.n6235 gnd.n6234 585
R3771 gnd.n6237 gnd.n1137 585
R3772 gnd.n6251 gnd.n1137 585
R3773 gnd.n6239 gnd.n6238 585
R3774 gnd.n6240 gnd.n6239 585
R3775 gnd.n1144 gnd.n1142 585
R3776 gnd.n6242 gnd.n1142 585
R3777 gnd.n6220 gnd.n6219 585
R3778 gnd.n6221 gnd.n6220 585
R3779 gnd.n6218 gnd.n1153 585
R3780 gnd.n1160 gnd.n1153 585
R3781 gnd.n6217 gnd.n6216 585
R3782 gnd.n6216 gnd.n6215 585
R3783 gnd.n1155 gnd.n1154 585
R3784 gnd.n1166 gnd.n1155 585
R3785 gnd.n1208 gnd.n1165 585
R3786 gnd.n6208 gnd.n1165 585
R3787 gnd.n1209 gnd.n1207 585
R3788 gnd.n1207 gnd.n1206 585
R3789 gnd.n1211 gnd.n1210 585
R3790 gnd.n1211 gnd.n1176 585
R3791 gnd.n1212 gnd.n1204 585
R3792 gnd.n1212 gnd.n1174 585
R3793 gnd.n6148 gnd.n6147 585
R3794 gnd.n6147 gnd.n6146 585
R3795 gnd.n6149 gnd.n1184 585
R3796 gnd.n6176 gnd.n1184 585
R3797 gnd.n6150 gnd.n1194 585
R3798 gnd.n6163 gnd.n1194 585
R3799 gnd.n6151 gnd.n1192 585
R3800 gnd.n6165 gnd.n1192 585
R3801 gnd.n6153 gnd.n6152 585
R3802 gnd.t87 gnd.n6153 585
R3803 gnd.n1203 gnd.n1202 585
R3804 gnd.n1202 gnd.n1200 585
R3805 gnd.n1296 gnd.n1295 585
R3806 gnd.n1296 gnd.n1218 585
R3807 gnd.n5963 gnd.n1431 585
R3808 gnd.n5698 gnd.n1431 585
R3809 gnd.n5965 gnd.n5964 585
R3810 gnd.n5966 gnd.n5965 585
R3811 gnd.n1432 gnd.n1430 585
R3812 gnd.n1452 gnd.n1430 585
R3813 gnd.n5866 gnd.n5865 585
R3814 gnd.n5865 gnd.n5864 585
R3815 gnd.n1435 gnd.n1434 585
R3816 gnd.n5854 gnd.n1435 585
R3817 gnd.n5451 gnd.n5450 585
R3818 gnd.n5452 gnd.n5451 585
R3819 gnd.n1501 gnd.n1500 585
R3820 gnd.n1500 gnd.n1498 585
R3821 gnd.n5446 gnd.n5445 585
R3822 gnd.n5445 gnd.n5444 585
R3823 gnd.n1504 gnd.n1503 585
R3824 gnd.n5432 gnd.n1504 585
R3825 gnd.n5417 gnd.n1527 585
R3826 gnd.n5403 gnd.n1527 585
R3827 gnd.n5419 gnd.n5418 585
R3828 gnd.n5420 gnd.n5419 585
R3829 gnd.n1528 gnd.n1526 585
R3830 gnd.n5353 gnd.n1526 585
R3831 gnd.n5412 gnd.n5411 585
R3832 gnd.n5411 gnd.n5410 585
R3833 gnd.n1531 gnd.n1530 585
R3834 gnd.n5386 gnd.n1531 585
R3835 gnd.n5374 gnd.n1563 585
R3836 gnd.n1563 gnd.n1550 585
R3837 gnd.n5376 gnd.n5375 585
R3838 gnd.n5377 gnd.n5376 585
R3839 gnd.n1564 gnd.n1562 585
R3840 gnd.n5348 gnd.n1562 585
R3841 gnd.n5369 gnd.n5368 585
R3842 gnd.n5368 gnd.n5367 585
R3843 gnd.n1567 gnd.n1566 585
R3844 gnd.n5344 gnd.n1567 585
R3845 gnd.n5332 gnd.n1594 585
R3846 gnd.n5318 gnd.n1594 585
R3847 gnd.n5334 gnd.n5333 585
R3848 gnd.n5335 gnd.n5334 585
R3849 gnd.n1595 gnd.n1593 585
R3850 gnd.n5312 gnd.n1593 585
R3851 gnd.n5327 gnd.n5326 585
R3852 gnd.n5326 gnd.n5325 585
R3853 gnd.n1598 gnd.n1597 585
R3854 gnd.n5308 gnd.n1598 585
R3855 gnd.n5296 gnd.n1623 585
R3856 gnd.n5282 gnd.n1623 585
R3857 gnd.n5298 gnd.n5297 585
R3858 gnd.n5299 gnd.n5298 585
R3859 gnd.n1624 gnd.n1622 585
R3860 gnd.n5276 gnd.n1622 585
R3861 gnd.n5291 gnd.n5290 585
R3862 gnd.n5290 gnd.n5289 585
R3863 gnd.n1633 gnd.n1632 585
R3864 gnd.n5272 gnd.n1633 585
R3865 gnd.n5260 gnd.n5259 585
R3866 gnd.n5259 gnd.n5258 585
R3867 gnd.n5262 gnd.n5261 585
R3868 gnd.n5263 gnd.n5262 585
R3869 gnd.n1673 gnd.n1656 585
R3870 gnd.n5250 gnd.n1656 585
R3871 gnd.n5238 gnd.n1674 585
R3872 gnd.n5238 gnd.n5237 585
R3873 gnd.n5241 gnd.n5240 585
R3874 gnd.n5242 gnd.n5241 585
R3875 gnd.n5239 gnd.n1672 585
R3876 gnd.n5229 gnd.n1672 585
R3877 gnd.n5221 gnd.n5220 585
R3878 gnd.n5222 gnd.n5221 585
R3879 gnd.n5219 gnd.n5218 585
R3880 gnd.n5218 gnd.n5217 585
R3881 gnd.n5200 gnd.n1686 585
R3882 gnd.n5214 gnd.n1686 585
R3883 gnd.n5201 gnd.n1702 585
R3884 gnd.n5185 gnd.n1702 585
R3885 gnd.n5203 gnd.n5202 585
R3886 gnd.n5204 gnd.n5203 585
R3887 gnd.n1703 gnd.n1701 585
R3888 gnd.n1701 gnd.n1698 585
R3889 gnd.n5196 gnd.n5195 585
R3890 gnd.n5195 gnd.n5194 585
R3891 gnd.n1706 gnd.n1705 585
R3892 gnd.n5177 gnd.n1706 585
R3893 gnd.n5164 gnd.n1729 585
R3894 gnd.n1729 gnd.n1719 585
R3895 gnd.n5166 gnd.n5165 585
R3896 gnd.n5167 gnd.n5166 585
R3897 gnd.n1730 gnd.n1728 585
R3898 gnd.n1728 gnd.n1725 585
R3899 gnd.n5159 gnd.n5158 585
R3900 gnd.n5158 gnd.n5157 585
R3901 gnd.n1733 gnd.n1732 585
R3902 gnd.n5142 gnd.n1733 585
R3903 gnd.n5129 gnd.n1753 585
R3904 gnd.n1753 gnd.n1744 585
R3905 gnd.n5131 gnd.n5130 585
R3906 gnd.n5132 gnd.n5131 585
R3907 gnd.n1754 gnd.n1752 585
R3908 gnd.n1760 gnd.n1752 585
R3909 gnd.n5124 gnd.n5123 585
R3910 gnd.n5123 gnd.n5122 585
R3911 gnd.n1757 gnd.n1756 585
R3912 gnd.n5107 gnd.n1757 585
R3913 gnd.n5094 gnd.n1778 585
R3914 gnd.n1778 gnd.n1769 585
R3915 gnd.n5096 gnd.n5095 585
R3916 gnd.n5097 gnd.n5096 585
R3917 gnd.n1779 gnd.n1777 585
R3918 gnd.n1786 gnd.n1777 585
R3919 gnd.n5089 gnd.n5088 585
R3920 gnd.n5088 gnd.n5087 585
R3921 gnd.n1782 gnd.n1781 585
R3922 gnd.n1783 gnd.n1782 585
R3923 gnd.n5070 gnd.n5069 585
R3924 gnd.n5071 gnd.n5070 585
R3925 gnd.n1799 gnd.n1798 585
R3926 gnd.n1798 gnd.n1795 585
R3927 gnd.n5065 gnd.n5064 585
R3928 gnd.n5064 gnd.n5063 585
R3929 gnd.n1802 gnd.n1801 585
R3930 gnd.n1803 gnd.n1802 585
R3931 gnd.n5050 gnd.n5049 585
R3932 gnd.n5051 gnd.n5050 585
R3933 gnd.n1816 gnd.n1815 585
R3934 gnd.n4730 gnd.n1815 585
R3935 gnd.n5045 gnd.n5044 585
R3936 gnd.n5044 gnd.n5043 585
R3937 gnd.n4884 gnd.n1818 585
R3938 gnd.n4887 gnd.n4886 585
R3939 gnd.n4883 gnd.n4882 585
R3940 gnd.n4882 gnd.n4727 585
R3941 gnd.n4892 gnd.n4891 585
R3942 gnd.n4894 gnd.n4881 585
R3943 gnd.n4897 gnd.n4896 585
R3944 gnd.n4879 gnd.n4878 585
R3945 gnd.n4902 gnd.n4901 585
R3946 gnd.n4904 gnd.n4877 585
R3947 gnd.n4907 gnd.n4906 585
R3948 gnd.n4875 gnd.n4874 585
R3949 gnd.n4912 gnd.n4911 585
R3950 gnd.n4914 gnd.n4873 585
R3951 gnd.n4917 gnd.n4916 585
R3952 gnd.n4871 gnd.n4870 585
R3953 gnd.n4922 gnd.n4921 585
R3954 gnd.n4924 gnd.n4866 585
R3955 gnd.n4927 gnd.n4926 585
R3956 gnd.n4864 gnd.n4863 585
R3957 gnd.n4932 gnd.n4931 585
R3958 gnd.n4934 gnd.n4862 585
R3959 gnd.n4937 gnd.n4936 585
R3960 gnd.n4860 gnd.n4859 585
R3961 gnd.n4942 gnd.n4941 585
R3962 gnd.n4944 gnd.n4858 585
R3963 gnd.n4947 gnd.n4946 585
R3964 gnd.n4856 gnd.n4855 585
R3965 gnd.n4952 gnd.n4951 585
R3966 gnd.n4954 gnd.n4854 585
R3967 gnd.n4957 gnd.n4956 585
R3968 gnd.n4852 gnd.n4851 585
R3969 gnd.n4962 gnd.n4961 585
R3970 gnd.n4964 gnd.n4850 585
R3971 gnd.n4967 gnd.n4966 585
R3972 gnd.n4848 gnd.n4847 585
R3973 gnd.n4972 gnd.n4971 585
R3974 gnd.n4974 gnd.n4846 585
R3975 gnd.n4979 gnd.n4976 585
R3976 gnd.n4844 gnd.n4843 585
R3977 gnd.n4984 gnd.n4983 585
R3978 gnd.n4986 gnd.n4842 585
R3979 gnd.n4989 gnd.n4988 585
R3980 gnd.n4840 gnd.n4839 585
R3981 gnd.n4994 gnd.n4993 585
R3982 gnd.n4996 gnd.n4838 585
R3983 gnd.n4999 gnd.n4998 585
R3984 gnd.n4836 gnd.n4835 585
R3985 gnd.n5004 gnd.n5003 585
R3986 gnd.n5006 gnd.n4834 585
R3987 gnd.n5009 gnd.n5008 585
R3988 gnd.n4832 gnd.n4831 585
R3989 gnd.n5014 gnd.n5013 585
R3990 gnd.n5016 gnd.n4830 585
R3991 gnd.n5019 gnd.n5018 585
R3992 gnd.n4828 gnd.n4827 585
R3993 gnd.n5025 gnd.n5024 585
R3994 gnd.n5027 gnd.n4826 585
R3995 gnd.n5028 gnd.n4825 585
R3996 gnd.n5031 gnd.n5030 585
R3997 gnd.n5974 gnd.n5973 585
R3998 gnd.n5976 gnd.n1417 585
R3999 gnd.n5978 gnd.n5977 585
R4000 gnd.n5979 gnd.n1410 585
R4001 gnd.n5981 gnd.n5980 585
R4002 gnd.n5983 gnd.n1408 585
R4003 gnd.n5985 gnd.n5984 585
R4004 gnd.n5986 gnd.n1403 585
R4005 gnd.n5988 gnd.n5987 585
R4006 gnd.n5990 gnd.n1401 585
R4007 gnd.n5992 gnd.n5991 585
R4008 gnd.n5993 gnd.n1396 585
R4009 gnd.n5995 gnd.n5994 585
R4010 gnd.n5997 gnd.n1394 585
R4011 gnd.n5999 gnd.n5998 585
R4012 gnd.n6000 gnd.n1389 585
R4013 gnd.n6002 gnd.n6001 585
R4014 gnd.n6004 gnd.n1388 585
R4015 gnd.n6005 gnd.n1385 585
R4016 gnd.n6008 gnd.n6007 585
R4017 gnd.n1387 gnd.n1381 585
R4018 gnd.n6012 gnd.n1378 585
R4019 gnd.n6014 gnd.n6013 585
R4020 gnd.n6016 gnd.n1376 585
R4021 gnd.n6018 gnd.n6017 585
R4022 gnd.n6019 gnd.n1371 585
R4023 gnd.n6021 gnd.n6020 585
R4024 gnd.n6023 gnd.n1370 585
R4025 gnd.n6024 gnd.n1366 585
R4026 gnd.n6027 gnd.n6026 585
R4027 gnd.n1367 gnd.n1361 585
R4028 gnd.n5916 gnd.n1362 585
R4029 gnd.n5918 gnd.n5917 585
R4030 gnd.n5919 gnd.n5909 585
R4031 gnd.n5921 gnd.n5920 585
R4032 gnd.n5923 gnd.n5907 585
R4033 gnd.n5925 gnd.n5924 585
R4034 gnd.n5926 gnd.n5899 585
R4035 gnd.n5928 gnd.n5927 585
R4036 gnd.n5930 gnd.n5897 585
R4037 gnd.n5932 gnd.n5931 585
R4038 gnd.n5933 gnd.n5892 585
R4039 gnd.n5935 gnd.n5934 585
R4040 gnd.n5937 gnd.n5890 585
R4041 gnd.n5939 gnd.n5938 585
R4042 gnd.n5940 gnd.n5885 585
R4043 gnd.n5942 gnd.n5941 585
R4044 gnd.n5944 gnd.n5883 585
R4045 gnd.n5946 gnd.n5945 585
R4046 gnd.n5947 gnd.n5878 585
R4047 gnd.n5949 gnd.n5948 585
R4048 gnd.n5951 gnd.n5876 585
R4049 gnd.n5953 gnd.n5952 585
R4050 gnd.n5954 gnd.n5872 585
R4051 gnd.n5956 gnd.n5955 585
R4052 gnd.n5958 gnd.n5871 585
R4053 gnd.n5960 gnd.n5959 585
R4054 gnd.n5959 gnd.n1369 585
R4055 gnd.n5969 gnd.n1419 585
R4056 gnd.n5698 gnd.n1419 585
R4057 gnd.n5968 gnd.n5967 585
R4058 gnd.n5967 gnd.n5966 585
R4059 gnd.n1425 gnd.n1424 585
R4060 gnd.n1452 gnd.n1425 585
R4061 gnd.n5857 gnd.n1437 585
R4062 gnd.n5864 gnd.n1437 585
R4063 gnd.n5856 gnd.n5855 585
R4064 gnd.n5855 gnd.n5854 585
R4065 gnd.n1445 gnd.n1444 585
R4066 gnd.n5452 gnd.n1445 585
R4067 gnd.n5437 gnd.n5436 585
R4068 gnd.n5436 gnd.n1498 585
R4069 gnd.n5435 gnd.n1506 585
R4070 gnd.n5444 gnd.n1506 585
R4071 gnd.n5434 gnd.n5433 585
R4072 gnd.n5433 gnd.n5432 585
R4073 gnd.n1515 gnd.n1513 585
R4074 gnd.n5403 gnd.n1515 585
R4075 gnd.n5352 gnd.n1524 585
R4076 gnd.n5420 gnd.n1524 585
R4077 gnd.n5355 gnd.n5354 585
R4078 gnd.n5354 gnd.n5353 585
R4079 gnd.n5356 gnd.n1533 585
R4080 gnd.n5410 gnd.n1533 585
R4081 gnd.n5357 gnd.n1551 585
R4082 gnd.n5386 gnd.n1551 585
R4083 gnd.n5359 gnd.n5358 585
R4084 gnd.n5358 gnd.n1550 585
R4085 gnd.n5351 gnd.n1559 585
R4086 gnd.n5377 gnd.n1559 585
R4087 gnd.n5350 gnd.n5349 585
R4088 gnd.n5349 gnd.n5348 585
R4089 gnd.n5347 gnd.n1569 585
R4090 gnd.n5367 gnd.n1569 585
R4091 gnd.n5346 gnd.n5345 585
R4092 gnd.n5345 gnd.n5344 585
R4093 gnd.n1581 gnd.n1579 585
R4094 gnd.n5318 gnd.n1581 585
R4095 gnd.n5315 gnd.n1590 585
R4096 gnd.n5335 gnd.n1590 585
R4097 gnd.n5314 gnd.n5313 585
R4098 gnd.n5313 gnd.n5312 585
R4099 gnd.n5311 gnd.n1600 585
R4100 gnd.n5325 gnd.n1600 585
R4101 gnd.n5310 gnd.n5309 585
R4102 gnd.n5309 gnd.n5308 585
R4103 gnd.n1610 gnd.n1608 585
R4104 gnd.n5282 gnd.n1610 585
R4105 gnd.n5279 gnd.n1619 585
R4106 gnd.n5299 gnd.n1619 585
R4107 gnd.n5278 gnd.n5277 585
R4108 gnd.n5277 gnd.n5276 585
R4109 gnd.n5275 gnd.n1635 585
R4110 gnd.n5289 gnd.n1635 585
R4111 gnd.n5274 gnd.n5273 585
R4112 gnd.n5273 gnd.n5272 585
R4113 gnd.n1645 gnd.n1643 585
R4114 gnd.n5258 gnd.n1645 585
R4115 gnd.n5253 gnd.n1653 585
R4116 gnd.n5263 gnd.n1653 585
R4117 gnd.n5252 gnd.n5251 585
R4118 gnd.n5251 gnd.n5250 585
R4119 gnd.n1661 gnd.n1660 585
R4120 gnd.n5237 gnd.n1661 585
R4121 gnd.n5244 gnd.n5243 585
R4122 gnd.n5243 gnd.n5242 585
R4123 gnd.n1667 gnd.n1666 585
R4124 gnd.n5229 gnd.n1667 585
R4125 gnd.n5224 gnd.n5223 585
R4126 gnd.n5223 gnd.n5222 585
R4127 gnd.n1684 gnd.n1683 585
R4128 gnd.n5217 gnd.n1684 585
R4129 gnd.n5184 gnd.n1692 585
R4130 gnd.n5214 gnd.n1692 585
R4131 gnd.n5187 gnd.n5186 585
R4132 gnd.n5186 gnd.n5185 585
R4133 gnd.n5183 gnd.n1699 585
R4134 gnd.n5204 gnd.n1699 585
R4135 gnd.n5182 gnd.n5181 585
R4136 gnd.n5181 gnd.n1698 585
R4137 gnd.n5180 gnd.n1707 585
R4138 gnd.n5194 gnd.n1707 585
R4139 gnd.n5179 gnd.n5178 585
R4140 gnd.n5178 gnd.n5177 585
R4141 gnd.n1718 gnd.n1716 585
R4142 gnd.n1719 gnd.n1718 585
R4143 gnd.n5148 gnd.n1726 585
R4144 gnd.n5167 gnd.n1726 585
R4145 gnd.n5147 gnd.n5146 585
R4146 gnd.n5146 gnd.n1725 585
R4147 gnd.n5145 gnd.n1734 585
R4148 gnd.n5157 gnd.n1734 585
R4149 gnd.n5144 gnd.n5143 585
R4150 gnd.n5143 gnd.n5142 585
R4151 gnd.n1743 gnd.n1741 585
R4152 gnd.n1744 gnd.n1743 585
R4153 gnd.n5113 gnd.n1750 585
R4154 gnd.n5132 gnd.n1750 585
R4155 gnd.n5112 gnd.n5111 585
R4156 gnd.n5111 gnd.n1760 585
R4157 gnd.n5110 gnd.n1758 585
R4158 gnd.n5122 gnd.n1758 585
R4159 gnd.n5109 gnd.n5108 585
R4160 gnd.n5108 gnd.n5107 585
R4161 gnd.n1768 gnd.n1766 585
R4162 gnd.n1769 gnd.n1768 585
R4163 gnd.n5078 gnd.n1775 585
R4164 gnd.n5097 gnd.n1775 585
R4165 gnd.n5077 gnd.n5076 585
R4166 gnd.n5076 gnd.n1786 585
R4167 gnd.n5075 gnd.n1784 585
R4168 gnd.n5087 gnd.n1784 585
R4169 gnd.n5074 gnd.n5073 585
R4170 gnd.n5073 gnd.n1783 585
R4171 gnd.n5072 gnd.n1792 585
R4172 gnd.n5072 gnd.n5071 585
R4173 gnd.n5056 gnd.n1794 585
R4174 gnd.n1795 gnd.n1794 585
R4175 gnd.n5055 gnd.n1804 585
R4176 gnd.n5063 gnd.n1804 585
R4177 gnd.n5054 gnd.n5053 585
R4178 gnd.n5053 gnd.n1803 585
R4179 gnd.n5052 gnd.n1810 585
R4180 gnd.n5052 gnd.n5051 585
R4181 gnd.n5038 gnd.n1812 585
R4182 gnd.n4730 gnd.n1812 585
R4183 gnd.n5037 gnd.n4728 585
R4184 gnd.n5043 gnd.n4728 585
R4185 gnd.n7665 gnd.n245 585
R4186 gnd.n245 gnd.n244 585
R4187 gnd.n7667 gnd.n7666 585
R4188 gnd.n7668 gnd.n7667 585
R4189 gnd.n232 gnd.n231 585
R4190 gnd.n235 gnd.n232 585
R4191 gnd.n7676 gnd.n7675 585
R4192 gnd.n7675 gnd.n7674 585
R4193 gnd.n7677 gnd.n226 585
R4194 gnd.n226 gnd.n225 585
R4195 gnd.n7679 gnd.n7678 585
R4196 gnd.n7680 gnd.n7679 585
R4197 gnd.n213 gnd.n212 585
R4198 gnd.n222 gnd.n213 585
R4199 gnd.n7688 gnd.n7687 585
R4200 gnd.n7687 gnd.n7686 585
R4201 gnd.n7689 gnd.n207 585
R4202 gnd.n207 gnd.n206 585
R4203 gnd.n7691 gnd.n7690 585
R4204 gnd.n7692 gnd.n7691 585
R4205 gnd.n193 gnd.n192 585
R4206 gnd.n197 gnd.n193 585
R4207 gnd.n7700 gnd.n7699 585
R4208 gnd.n7699 gnd.n7698 585
R4209 gnd.n7701 gnd.n187 585
R4210 gnd.n194 gnd.n187 585
R4211 gnd.n7703 gnd.n7702 585
R4212 gnd.n7704 gnd.n7703 585
R4213 gnd.n175 gnd.n174 585
R4214 gnd.n184 gnd.n175 585
R4215 gnd.n7712 gnd.n7711 585
R4216 gnd.n7711 gnd.n7710 585
R4217 gnd.n7713 gnd.n169 585
R4218 gnd.n169 gnd.n168 585
R4219 gnd.n7715 gnd.n7714 585
R4220 gnd.n7716 gnd.n7715 585
R4221 gnd.n155 gnd.n154 585
R4222 gnd.n159 gnd.n155 585
R4223 gnd.n7724 gnd.n7723 585
R4224 gnd.n7723 gnd.n7722 585
R4225 gnd.n7725 gnd.n149 585
R4226 gnd.n156 gnd.n149 585
R4227 gnd.n7727 gnd.n7726 585
R4228 gnd.n7728 gnd.n7727 585
R4229 gnd.n137 gnd.n136 585
R4230 gnd.n146 gnd.n137 585
R4231 gnd.n7736 gnd.n7735 585
R4232 gnd.n7735 gnd.n7734 585
R4233 gnd.n7737 gnd.n132 585
R4234 gnd.n132 gnd.n131 585
R4235 gnd.n7739 gnd.n7738 585
R4236 gnd.n7740 gnd.n7739 585
R4237 gnd.n116 gnd.n114 585
R4238 gnd.n7490 gnd.n116 585
R4239 gnd.n7748 gnd.n7747 585
R4240 gnd.n7747 gnd.n7746 585
R4241 gnd.n115 gnd.n107 585
R4242 gnd.n7360 gnd.n115 585
R4243 gnd.n7751 gnd.n105 585
R4244 gnd.n7353 gnd.n105 585
R4245 gnd.n7753 gnd.n7752 585
R4246 gnd.n7754 gnd.n7753 585
R4247 gnd.n7332 gnd.n104 585
R4248 gnd.n7343 gnd.n104 585
R4249 gnd.n7334 gnd.n7333 585
R4250 gnd.n7335 gnd.n7334 585
R4251 gnd.n7331 gnd.n371 585
R4252 gnd.n7331 gnd.n7330 585
R4253 gnd.n370 gnd.n369 585
R4254 gnd.n7323 gnd.n369 585
R4255 gnd.n7311 gnd.n7310 585
R4256 gnd.n7312 gnd.n7311 585
R4257 gnd.n7309 gnd.n7308 585
R4258 gnd.n7308 gnd.n7307 585
R4259 gnd.n7281 gnd.n386 585
R4260 gnd.n7299 gnd.n386 585
R4261 gnd.n7282 gnd.n407 585
R4262 gnd.n7268 gnd.n407 585
R4263 gnd.n7284 gnd.n7283 585
R4264 gnd.n7285 gnd.n7284 585
R4265 gnd.n408 gnd.n406 585
R4266 gnd.n7262 gnd.n406 585
R4267 gnd.n7277 gnd.n7276 585
R4268 gnd.n7276 gnd.n7275 585
R4269 gnd.n411 gnd.n410 585
R4270 gnd.n7258 gnd.n411 585
R4271 gnd.n7235 gnd.n7234 585
R4272 gnd.n7236 gnd.n7235 585
R4273 gnd.n435 gnd.n434 585
R4274 gnd.n434 gnd.n431 585
R4275 gnd.n7230 gnd.n7229 585
R4276 gnd.n7229 gnd.n7228 585
R4277 gnd.n438 gnd.n437 585
R4278 gnd.n7216 gnd.n438 585
R4279 gnd.n7195 gnd.n461 585
R4280 gnd.n7181 gnd.n461 585
R4281 gnd.n7197 gnd.n7196 585
R4282 gnd.n7198 gnd.n7197 585
R4283 gnd.n462 gnd.n460 585
R4284 gnd.n509 gnd.n460 585
R4285 gnd.n7190 gnd.n7189 585
R4286 gnd.n7189 gnd.n7188 585
R4287 gnd.n465 gnd.n464 585
R4288 gnd.n7144 gnd.n465 585
R4289 gnd.n7160 gnd.n7159 585
R4290 gnd.n7161 gnd.n7160 585
R4291 gnd.n493 gnd.n492 585
R4292 gnd.n492 gnd.n487 585
R4293 gnd.n7155 gnd.n7154 585
R4294 gnd.n7154 gnd.n7153 585
R4295 gnd.n496 gnd.n495 585
R4296 gnd.n543 gnd.n496 585
R4297 gnd.n7125 gnd.n526 585
R4298 gnd.n7111 gnd.n526 585
R4299 gnd.n7127 gnd.n7126 585
R4300 gnd.n7128 gnd.n7127 585
R4301 gnd.n527 gnd.n525 585
R4302 gnd.n7099 gnd.n525 585
R4303 gnd.n7120 gnd.n7119 585
R4304 gnd.n7119 gnd.n7118 585
R4305 gnd.n530 gnd.n529 585
R4306 gnd.n7087 gnd.n530 585
R4307 gnd.n7075 gnd.n565 585
R4308 gnd.n577 gnd.n565 585
R4309 gnd.n7077 gnd.n7076 585
R4310 gnd.n7078 gnd.n7077 585
R4311 gnd.n566 gnd.n564 585
R4312 gnd.n7060 gnd.n564 585
R4313 gnd.n7070 gnd.n7069 585
R4314 gnd.n7069 gnd.n7068 585
R4315 gnd.n629 gnd.n568 585
R4316 gnd.n7039 gnd.n7038 585
R4317 gnd.n7037 gnd.n628 585
R4318 gnd.n7041 gnd.n628 585
R4319 gnd.n7036 gnd.n7035 585
R4320 gnd.n7034 gnd.n7033 585
R4321 gnd.n7032 gnd.n7031 585
R4322 gnd.n7030 gnd.n7029 585
R4323 gnd.n7028 gnd.n7027 585
R4324 gnd.n7026 gnd.n7025 585
R4325 gnd.n7024 gnd.n7023 585
R4326 gnd.n7022 gnd.n7021 585
R4327 gnd.n7020 gnd.n7019 585
R4328 gnd.n7018 gnd.n7017 585
R4329 gnd.n7016 gnd.n7015 585
R4330 gnd.n7014 gnd.n7013 585
R4331 gnd.n7012 gnd.n7011 585
R4332 gnd.n7010 gnd.n7009 585
R4333 gnd.n7008 gnd.n7007 585
R4334 gnd.n7005 gnd.n7004 585
R4335 gnd.n7003 gnd.n7002 585
R4336 gnd.n7001 gnd.n7000 585
R4337 gnd.n6999 gnd.n6998 585
R4338 gnd.n6997 gnd.n6996 585
R4339 gnd.n6995 gnd.n6994 585
R4340 gnd.n6993 gnd.n6992 585
R4341 gnd.n6991 gnd.n6990 585
R4342 gnd.n6988 gnd.n6987 585
R4343 gnd.n6986 gnd.n6985 585
R4344 gnd.n6984 gnd.n6983 585
R4345 gnd.n6982 gnd.n6981 585
R4346 gnd.n6980 gnd.n6979 585
R4347 gnd.n6978 gnd.n6977 585
R4348 gnd.n6976 gnd.n6975 585
R4349 gnd.n6974 gnd.n6973 585
R4350 gnd.n6972 gnd.n6971 585
R4351 gnd.n6970 gnd.n6969 585
R4352 gnd.n6968 gnd.n6967 585
R4353 gnd.n6966 gnd.n6965 585
R4354 gnd.n6964 gnd.n6963 585
R4355 gnd.n6962 gnd.n6961 585
R4356 gnd.n6960 gnd.n6959 585
R4357 gnd.n6958 gnd.n6957 585
R4358 gnd.n6956 gnd.n6955 585
R4359 gnd.n6954 gnd.n6953 585
R4360 gnd.n6952 gnd.n6951 585
R4361 gnd.n6950 gnd.n6949 585
R4362 gnd.n6948 gnd.n6947 585
R4363 gnd.n6946 gnd.n6945 585
R4364 gnd.n6944 gnd.n6943 585
R4365 gnd.n6942 gnd.n6941 585
R4366 gnd.n6940 gnd.n6939 585
R4367 gnd.n6938 gnd.n6937 585
R4368 gnd.n6936 gnd.n6935 585
R4369 gnd.n6934 gnd.n6933 585
R4370 gnd.n6932 gnd.n6931 585
R4371 gnd.n6930 gnd.n6929 585
R4372 gnd.n692 gnd.n691 585
R4373 gnd.n7536 gnd.n345 585
R4374 gnd.n7544 gnd.n7543 585
R4375 gnd.n7546 gnd.n7545 585
R4376 gnd.n7548 gnd.n7547 585
R4377 gnd.n7550 gnd.n7549 585
R4378 gnd.n7552 gnd.n7551 585
R4379 gnd.n7554 gnd.n7553 585
R4380 gnd.n7556 gnd.n7555 585
R4381 gnd.n7558 gnd.n7557 585
R4382 gnd.n7560 gnd.n7559 585
R4383 gnd.n7562 gnd.n7561 585
R4384 gnd.n7564 gnd.n7563 585
R4385 gnd.n7566 gnd.n7565 585
R4386 gnd.n7568 gnd.n7567 585
R4387 gnd.n7570 gnd.n7569 585
R4388 gnd.n7572 gnd.n7571 585
R4389 gnd.n7574 gnd.n7573 585
R4390 gnd.n7576 gnd.n7575 585
R4391 gnd.n7578 gnd.n7577 585
R4392 gnd.n7581 gnd.n7580 585
R4393 gnd.n7579 gnd.n325 585
R4394 gnd.n7586 gnd.n7585 585
R4395 gnd.n7588 gnd.n7587 585
R4396 gnd.n7590 gnd.n7589 585
R4397 gnd.n7592 gnd.n7591 585
R4398 gnd.n7594 gnd.n7593 585
R4399 gnd.n7596 gnd.n7595 585
R4400 gnd.n7598 gnd.n7597 585
R4401 gnd.n7600 gnd.n7599 585
R4402 gnd.n7602 gnd.n7601 585
R4403 gnd.n7604 gnd.n7603 585
R4404 gnd.n7606 gnd.n7605 585
R4405 gnd.n7608 gnd.n7607 585
R4406 gnd.n7610 gnd.n7609 585
R4407 gnd.n7612 gnd.n7611 585
R4408 gnd.n7614 gnd.n7613 585
R4409 gnd.n7616 gnd.n7615 585
R4410 gnd.n7618 gnd.n7617 585
R4411 gnd.n7620 gnd.n7619 585
R4412 gnd.n7622 gnd.n7621 585
R4413 gnd.n7624 gnd.n7623 585
R4414 gnd.n7629 gnd.n7628 585
R4415 gnd.n7631 gnd.n7630 585
R4416 gnd.n7633 gnd.n7632 585
R4417 gnd.n7635 gnd.n7634 585
R4418 gnd.n7637 gnd.n7636 585
R4419 gnd.n7639 gnd.n7638 585
R4420 gnd.n7641 gnd.n7640 585
R4421 gnd.n7643 gnd.n7642 585
R4422 gnd.n7645 gnd.n7644 585
R4423 gnd.n7647 gnd.n7646 585
R4424 gnd.n7649 gnd.n7648 585
R4425 gnd.n7651 gnd.n7650 585
R4426 gnd.n7653 gnd.n7652 585
R4427 gnd.n7655 gnd.n7654 585
R4428 gnd.n7656 gnd.n289 585
R4429 gnd.n7658 gnd.n7657 585
R4430 gnd.n250 gnd.n249 585
R4431 gnd.n7662 gnd.n7661 585
R4432 gnd.n7661 gnd.n7660 585
R4433 gnd.n7538 gnd.n7537 585
R4434 gnd.n7537 gnd.n244 585
R4435 gnd.n7535 gnd.n242 585
R4436 gnd.n7668 gnd.n242 585
R4437 gnd.n7534 gnd.n7533 585
R4438 gnd.n7533 gnd.n235 585
R4439 gnd.n7532 gnd.n233 585
R4440 gnd.n7674 gnd.n233 585
R4441 gnd.n7531 gnd.n7530 585
R4442 gnd.n7530 gnd.n225 585
R4443 gnd.n7528 gnd.n223 585
R4444 gnd.n7680 gnd.n223 585
R4445 gnd.n7527 gnd.n7526 585
R4446 gnd.n7526 gnd.n222 585
R4447 gnd.n7525 gnd.n214 585
R4448 gnd.n7686 gnd.n214 585
R4449 gnd.n7524 gnd.n7523 585
R4450 gnd.n7523 gnd.n206 585
R4451 gnd.n7521 gnd.n204 585
R4452 gnd.n7692 gnd.n204 585
R4453 gnd.n7520 gnd.n7519 585
R4454 gnd.n7519 gnd.n197 585
R4455 gnd.n7518 gnd.n195 585
R4456 gnd.n7698 gnd.n195 585
R4457 gnd.n7517 gnd.n7516 585
R4458 gnd.n7516 gnd.n194 585
R4459 gnd.n7514 gnd.n185 585
R4460 gnd.n7704 gnd.n185 585
R4461 gnd.n7513 gnd.n7512 585
R4462 gnd.n7512 gnd.n184 585
R4463 gnd.n7511 gnd.n176 585
R4464 gnd.n7710 gnd.n176 585
R4465 gnd.n7510 gnd.n7509 585
R4466 gnd.n7509 gnd.n168 585
R4467 gnd.n7507 gnd.n166 585
R4468 gnd.n7716 gnd.n166 585
R4469 gnd.n7506 gnd.n7505 585
R4470 gnd.n7505 gnd.n159 585
R4471 gnd.n7504 gnd.n157 585
R4472 gnd.n7722 gnd.n157 585
R4473 gnd.n7503 gnd.n7502 585
R4474 gnd.n7502 gnd.n156 585
R4475 gnd.n7500 gnd.n147 585
R4476 gnd.n7728 gnd.n147 585
R4477 gnd.n7499 gnd.n7498 585
R4478 gnd.n7498 gnd.n146 585
R4479 gnd.n7497 gnd.n138 585
R4480 gnd.n7734 gnd.n138 585
R4481 gnd.n7496 gnd.n7495 585
R4482 gnd.n7495 gnd.n131 585
R4483 gnd.n7493 gnd.n129 585
R4484 gnd.n7740 gnd.n129 585
R4485 gnd.n7492 gnd.n7491 585
R4486 gnd.n7491 gnd.n7490 585
R4487 gnd.n349 gnd.n118 585
R4488 gnd.n7746 gnd.n118 585
R4489 gnd.n7359 gnd.n7358 585
R4490 gnd.n7360 gnd.n7359 585
R4491 gnd.n353 gnd.n352 585
R4492 gnd.n7353 gnd.n352 585
R4493 gnd.n7338 gnd.n101 585
R4494 gnd.n7754 gnd.n101 585
R4495 gnd.n7339 gnd.n361 585
R4496 gnd.n7343 gnd.n361 585
R4497 gnd.n7337 gnd.n7336 585
R4498 gnd.n7336 gnd.n7335 585
R4499 gnd.n366 gnd.n365 585
R4500 gnd.n7330 gnd.n366 585
R4501 gnd.n7325 gnd.n7324 585
R4502 gnd.n7324 gnd.n7323 585
R4503 gnd.n377 gnd.n376 585
R4504 gnd.n7312 gnd.n377 585
R4505 gnd.n7302 gnd.n388 585
R4506 gnd.n7307 gnd.n388 585
R4507 gnd.n7301 gnd.n7300 585
R4508 gnd.n7300 gnd.n7299 585
R4509 gnd.n394 gnd.n393 585
R4510 gnd.n7268 gnd.n394 585
R4511 gnd.n7265 gnd.n403 585
R4512 gnd.n7285 gnd.n403 585
R4513 gnd.n7264 gnd.n7263 585
R4514 gnd.n7263 gnd.n7262 585
R4515 gnd.n7261 gnd.n412 585
R4516 gnd.n7275 gnd.n412 585
R4517 gnd.n7260 gnd.n7259 585
R4518 gnd.n7259 gnd.n7258 585
R4519 gnd.n422 gnd.n420 585
R4520 gnd.n7236 gnd.n422 585
R4521 gnd.n7221 gnd.n7220 585
R4522 gnd.n7220 gnd.n431 585
R4523 gnd.n7219 gnd.n440 585
R4524 gnd.n7228 gnd.n440 585
R4525 gnd.n7218 gnd.n7217 585
R4526 gnd.n7217 gnd.n7216 585
R4527 gnd.n449 gnd.n447 585
R4528 gnd.n7181 gnd.n449 585
R4529 gnd.n508 gnd.n457 585
R4530 gnd.n7198 gnd.n457 585
R4531 gnd.n511 gnd.n510 585
R4532 gnd.n510 gnd.n509 585
R4533 gnd.n512 gnd.n467 585
R4534 gnd.n7188 gnd.n467 585
R4535 gnd.n7146 gnd.n7145 585
R4536 gnd.n7145 gnd.n7144 585
R4537 gnd.n7147 gnd.n488 585
R4538 gnd.n7161 gnd.n488 585
R4539 gnd.n507 gnd.n506 585
R4540 gnd.n506 gnd.n487 585
R4541 gnd.n7092 gnd.n497 585
R4542 gnd.n7153 gnd.n497 585
R4543 gnd.n7094 gnd.n7093 585
R4544 gnd.n7093 gnd.n543 585
R4545 gnd.n7095 gnd.n542 585
R4546 gnd.n7111 gnd.n542 585
R4547 gnd.n7096 gnd.n522 585
R4548 gnd.n7128 gnd.n522 585
R4549 gnd.n7098 gnd.n7097 585
R4550 gnd.n7099 gnd.n7098 585
R4551 gnd.n7090 gnd.n532 585
R4552 gnd.n7118 gnd.n532 585
R4553 gnd.n7089 gnd.n7088 585
R4554 gnd.n7088 gnd.n7087 585
R4555 gnd.n553 gnd.n551 585
R4556 gnd.n577 gnd.n553 585
R4557 gnd.n7062 gnd.n561 585
R4558 gnd.n7078 gnd.n561 585
R4559 gnd.n7063 gnd.n7061 585
R4560 gnd.n7061 gnd.n7060 585
R4561 gnd.n582 gnd.n570 585
R4562 gnd.n7068 gnd.n570 585
R4563 gnd.n3319 gnd.n1974 585
R4564 gnd.n1974 gnd.n1691 585
R4565 gnd.n2601 gnd.n2600 585
R4566 gnd.n2601 gnd.n120 585
R4567 gnd.n357 gnd.n117 585
R4568 gnd.n7351 gnd.n7350 585
R4569 gnd.n7352 gnd.n7351 585
R4570 gnd.n7348 gnd.n356 585
R4571 gnd.n356 gnd.n102 585
R4572 gnd.n7346 gnd.n7345 585
R4573 gnd.n7345 gnd.n7344 585
R4574 gnd.n359 gnd.n358 585
R4575 gnd.n360 gnd.n359 585
R4576 gnd.n7319 gnd.n381 585
R4577 gnd.n381 gnd.n367 585
R4578 gnd.n7321 gnd.n7320 585
R4579 gnd.n7322 gnd.n7321 585
R4580 gnd.n7316 gnd.n380 585
R4581 gnd.n380 gnd.n378 585
R4582 gnd.n7315 gnd.n7314 585
R4583 gnd.n7314 gnd.n7313 585
R4584 gnd.n7248 gnd.n383 585
R4585 gnd.n387 gnd.n383 585
R4586 gnd.n7250 gnd.n7249 585
R4587 gnd.n7250 gnd.n395 585
R4588 gnd.n7251 gnd.n7245 585
R4589 gnd.n7251 gnd.n404 585
R4590 gnd.n7253 gnd.n7252 585
R4591 gnd.n7252 gnd.n402 585
R4592 gnd.n7254 gnd.n426 585
R4593 gnd.n426 gnd.n414 585
R4594 gnd.n7256 gnd.n7255 585
R4595 gnd.n7257 gnd.n7256 585
R4596 gnd.n427 gnd.n425 585
R4597 gnd.n425 gnd.n423 585
R4598 gnd.n7239 gnd.n7238 585
R4599 gnd.n7238 gnd.n7237 585
R4600 gnd.n430 gnd.n429 585
R4601 gnd.n442 gnd.n430 585
R4602 gnd.n7177 gnd.n478 585
R4603 gnd.n478 gnd.n439 585
R4604 gnd.n7179 gnd.n7178 585
R4605 gnd.n7180 gnd.n7179 585
R4606 gnd.n479 gnd.n477 585
R4607 gnd.n477 gnd.n458 585
R4608 gnd.n7172 gnd.n7171 585
R4609 gnd.n7171 gnd.n456 585
R4610 gnd.n7170 gnd.n481 585
R4611 gnd.n7170 gnd.n469 585
R4612 gnd.n7169 gnd.n7168 585
R4613 gnd.n7169 gnd.n466 585
R4614 gnd.n483 gnd.n482 585
R4615 gnd.n490 gnd.n482 585
R4616 gnd.n7164 gnd.n7163 585
R4617 gnd.n7163 gnd.n7162 585
R4618 gnd.n486 gnd.n485 585
R4619 gnd.n499 gnd.n486 585
R4620 gnd.n7107 gnd.n546 585
R4621 gnd.n546 gnd.n545 585
R4622 gnd.n7109 gnd.n7108 585
R4623 gnd.n7110 gnd.n7109 585
R4624 gnd.n547 gnd.n544 585
R4625 gnd.n544 gnd.n523 585
R4626 gnd.n7102 gnd.n7101 585
R4627 gnd.n7101 gnd.n7100 585
R4628 gnd.n550 gnd.n549 585
R4629 gnd.n550 gnd.n534 585
R4630 gnd.n7053 gnd.n7052 585
R4631 gnd.n7053 gnd.n531 585
R4632 gnd.n7055 gnd.n7054 585
R4633 gnd.n7054 gnd.n554 585
R4634 gnd.n7056 gnd.n584 585
R4635 gnd.n584 gnd.n562 585
R4636 gnd.n7058 gnd.n7057 585
R4637 gnd.n7059 gnd.n7058 585
R4638 gnd.n585 gnd.n583 585
R4639 gnd.n583 gnd.n572 585
R4640 gnd.n7045 gnd.n7044 585
R4641 gnd.n7044 gnd.n569 585
R4642 gnd.n7043 gnd.n587 585
R4643 gnd.n7043 gnd.n7042 585
R4644 gnd.n6841 gnd.n588 585
R4645 gnd.n589 gnd.n588 585
R4646 gnd.n6843 gnd.n6842 585
R4647 gnd.n6844 gnd.n6843 585
R4648 gnd.n797 gnd.n796 585
R4649 gnd.n796 gnd.n776 585
R4650 gnd.n6836 gnd.n6835 585
R4651 gnd.n6835 gnd.n764 585
R4652 gnd.n6834 gnd.n799 585
R4653 gnd.n6834 gnd.n763 585
R4654 gnd.n6833 gnd.n801 585
R4655 gnd.n6833 gnd.n6832 585
R4656 gnd.n6818 gnd.n800 585
R4657 gnd.n802 gnd.n800 585
R4658 gnd.n6820 gnd.n6819 585
R4659 gnd.n6821 gnd.n6820 585
R4660 gnd.n813 gnd.n812 585
R4661 gnd.n812 gnd.n809 585
R4662 gnd.n6812 gnd.n6811 585
R4663 gnd.n6811 gnd.n6810 585
R4664 gnd.n816 gnd.n815 585
R4665 gnd.n825 gnd.n816 585
R4666 gnd.n6782 gnd.n837 585
R4667 gnd.n837 gnd.n824 585
R4668 gnd.n6784 gnd.n6783 585
R4669 gnd.n6785 gnd.n6784 585
R4670 gnd.n838 gnd.n836 585
R4671 gnd.n836 gnd.n833 585
R4672 gnd.n6777 gnd.n6776 585
R4673 gnd.n6776 gnd.n6775 585
R4674 gnd.n841 gnd.n840 585
R4675 gnd.n849 gnd.n841 585
R4676 gnd.n6752 gnd.n862 585
R4677 gnd.n862 gnd.n848 585
R4678 gnd.n6754 gnd.n6753 585
R4679 gnd.n6755 gnd.n6754 585
R4680 gnd.n863 gnd.n861 585
R4681 gnd.n861 gnd.n858 585
R4682 gnd.n6747 gnd.n6746 585
R4683 gnd.n6746 gnd.n6745 585
R4684 gnd.n866 gnd.n865 585
R4685 gnd.n874 gnd.n866 585
R4686 gnd.n6722 gnd.n886 585
R4687 gnd.n886 gnd.n873 585
R4688 gnd.n6724 gnd.n6723 585
R4689 gnd.n6725 gnd.n6724 585
R4690 gnd.n887 gnd.n885 585
R4691 gnd.n6713 gnd.n885 585
R4692 gnd.n6717 gnd.n6716 585
R4693 gnd.n6716 gnd.n6715 585
R4694 gnd.n890 gnd.n889 585
R4695 gnd.n932 gnd.n890 585
R4696 gnd.n6546 gnd.n6545 585
R4697 gnd.n6547 gnd.n6546 585
R4698 gnd.n941 gnd.n940 585
R4699 gnd.n6470 gnd.n940 585
R4700 gnd.n6541 gnd.n6540 585
R4701 gnd.n6540 gnd.n6539 585
R4702 gnd.n944 gnd.n943 585
R4703 gnd.n952 gnd.n944 585
R4704 gnd.n6483 gnd.n990 585
R4705 gnd.n6483 gnd.n6482 585
R4706 gnd.n6485 gnd.n6484 585
R4707 gnd.n6484 gnd.n973 585
R4708 gnd.n6486 gnd.n984 585
R4709 gnd.n6456 gnd.n984 585
R4710 gnd.n6488 gnd.n6487 585
R4711 gnd.n6489 gnd.n6488 585
R4712 gnd.n985 gnd.n983 585
R4713 gnd.n1006 gnd.n983 585
R4714 gnd.n1038 gnd.n1037 585
R4715 gnd.n1038 gnd.n1014 585
R4716 gnd.n6421 gnd.n6420 585
R4717 gnd.n6420 gnd.n6419 585
R4718 gnd.n6422 gnd.n1030 585
R4719 gnd.n1030 gnd.n1022 585
R4720 gnd.n6424 gnd.n6423 585
R4721 gnd.n6425 gnd.n6424 585
R4722 gnd.n1031 gnd.n1029 585
R4723 gnd.n6406 gnd.n1029 585
R4724 gnd.n6382 gnd.n6381 585
R4725 gnd.n6381 gnd.n6380 585
R4726 gnd.n6383 gnd.n1060 585
R4727 gnd.n1060 gnd.n1052 585
R4728 gnd.n6385 gnd.n6384 585
R4729 gnd.n6386 gnd.n6385 585
R4730 gnd.n1061 gnd.n1059 585
R4731 gnd.n6369 gnd.n1059 585
R4732 gnd.n6344 gnd.n6343 585
R4733 gnd.n6343 gnd.n6342 585
R4734 gnd.n6345 gnd.n1087 585
R4735 gnd.n1087 gnd.n1079 585
R4736 gnd.n6347 gnd.n6346 585
R4737 gnd.n6348 gnd.n6347 585
R4738 gnd.n1088 gnd.n1086 585
R4739 gnd.n1100 gnd.n1086 585
R4740 gnd.n6282 gnd.n6281 585
R4741 gnd.n6281 gnd.n6280 585
R4742 gnd.n6283 gnd.n1119 585
R4743 gnd.n1119 gnd.n1109 585
R4744 gnd.n6285 gnd.n6284 585
R4745 gnd.n6286 gnd.n6285 585
R4746 gnd.n1120 gnd.n1118 585
R4747 gnd.n1118 gnd.n1114 585
R4748 gnd.n6231 gnd.n6230 585
R4749 gnd.n6232 gnd.n6231 585
R4750 gnd.n1148 gnd.n1147 585
R4751 gnd.n1147 gnd.n1145 585
R4752 gnd.n6225 gnd.n6224 585
R4753 gnd.n6224 gnd.n1135 585
R4754 gnd.n6223 gnd.n1150 585
R4755 gnd.n6223 gnd.n6222 585
R4756 gnd.n6203 gnd.n1151 585
R4757 gnd.n1159 gnd.n1151 585
R4758 gnd.n6204 gnd.n1169 585
R4759 gnd.n1169 gnd.n1156 585
R4760 gnd.n6206 gnd.n6205 585
R4761 gnd.n6207 gnd.n6206 585
R4762 gnd.n1170 gnd.n1168 585
R4763 gnd.n1205 gnd.n1168 585
R4764 gnd.n6197 gnd.n6196 585
R4765 gnd.n6196 gnd.n6195 585
R4766 gnd.n1173 gnd.n1172 585
R4767 gnd.n1186 gnd.n1173 585
R4768 gnd.n6161 gnd.n6160 585
R4769 gnd.n6162 gnd.n6161 585
R4770 gnd.n1196 gnd.n1195 585
R4771 gnd.n1195 gnd.n1191 585
R4772 gnd.n6156 gnd.n6155 585
R4773 gnd.n6155 gnd.n6154 585
R4774 gnd.n1199 gnd.n1198 585
R4775 gnd.n1260 gnd.n1199 585
R4776 gnd.n5648 gnd.n5647 585
R4777 gnd.n5647 gnd.n1262 585
R4778 gnd.n5649 gnd.n5507 585
R4779 gnd.n5507 gnd.n1226 585
R4780 gnd.n5651 gnd.n5650 585
R4781 gnd.n5652 gnd.n5651 585
R4782 gnd.n5508 gnd.n5506 585
R4783 gnd.n5506 gnd.n5503 585
R4784 gnd.n5641 gnd.n5640 585
R4785 gnd.n5640 gnd.n5639 585
R4786 gnd.n5511 gnd.n5510 585
R4787 gnd.n5619 gnd.n5511 585
R4788 gnd.n5617 gnd.n5616 585
R4789 gnd.n5618 gnd.n5617 585
R4790 gnd.n5521 gnd.n5520 585
R4791 gnd.n5608 gnd.n5520 585
R4792 gnd.n5612 gnd.n5611 585
R4793 gnd.n5611 gnd.n5610 585
R4794 gnd.n5524 gnd.n5523 585
R4795 gnd.n5598 gnd.n5524 585
R4796 gnd.n5596 gnd.n5595 585
R4797 gnd.n5597 gnd.n5596 585
R4798 gnd.n5533 gnd.n5532 585
R4799 gnd.n5587 gnd.n5532 585
R4800 gnd.n5591 gnd.n5590 585
R4801 gnd.n5590 gnd.n5589 585
R4802 gnd.n5536 gnd.n5535 585
R4803 gnd.n5577 gnd.n5536 585
R4804 gnd.n5575 gnd.n5574 585
R4805 gnd.n5576 gnd.n5575 585
R4806 gnd.n5545 gnd.n5544 585
R4807 gnd.n5566 gnd.n5544 585
R4808 gnd.n5570 gnd.n5569 585
R4809 gnd.n5569 gnd.n5568 585
R4810 gnd.n5549 gnd.n5548 585
R4811 gnd.n5557 gnd.n5549 585
R4812 gnd.n5476 gnd.n5475 585
R4813 gnd.n5480 gnd.n5476 585
R4814 gnd.n5685 gnd.n5684 585
R4815 gnd.n5684 gnd.n5683 585
R4816 gnd.n5686 gnd.n5470 585
R4817 gnd.n5477 gnd.n5470 585
R4818 gnd.n5688 gnd.n5687 585
R4819 gnd.n5688 gnd.n1474 585
R4820 gnd.n5689 gnd.n5469 585
R4821 gnd.n5689 gnd.n1460 585
R4822 gnd.n5693 gnd.n5692 585
R4823 gnd.n5692 gnd.n5691 585
R4824 gnd.n5694 gnd.n1489 585
R4825 gnd.n5690 gnd.n1489 585
R4826 gnd.n5696 gnd.n5695 585
R4827 gnd.n5697 gnd.n5696 585
R4828 gnd.n1490 gnd.n1488 585
R4829 gnd.n1488 gnd.n1428 585
R4830 gnd.n5463 gnd.n5462 585
R4831 gnd.n5462 gnd.n1426 585
R4832 gnd.n5461 gnd.n1492 585
R4833 gnd.n5461 gnd.n1439 585
R4834 gnd.n5460 gnd.n5459 585
R4835 gnd.n5460 gnd.n1436 585
R4836 gnd.n1494 gnd.n1493 585
R4837 gnd.n1493 gnd.n1446 585
R4838 gnd.n5455 gnd.n5454 585
R4839 gnd.n5454 gnd.n5453 585
R4840 gnd.n1497 gnd.n1496 585
R4841 gnd.n1508 gnd.n1497 585
R4842 gnd.n5398 gnd.n5397 585
R4843 gnd.n5397 gnd.n1505 585
R4844 gnd.n5399 gnd.n1544 585
R4845 gnd.n1544 gnd.n1516 585
R4846 gnd.n5401 gnd.n5400 585
R4847 gnd.n5402 gnd.n5401 585
R4848 gnd.n1545 gnd.n1543 585
R4849 gnd.n1543 gnd.n1523 585
R4850 gnd.n5391 gnd.n5390 585
R4851 gnd.n5390 gnd.n1535 585
R4852 gnd.n5389 gnd.n1547 585
R4853 gnd.n5389 gnd.n1532 585
R4854 gnd.n5388 gnd.n1549 585
R4855 gnd.n5388 gnd.n5387 585
R4856 gnd.n1939 gnd.n1548 585
R4857 gnd.n1560 gnd.n1548 585
R4858 gnd.n1940 gnd.n1933 585
R4859 gnd.n1933 gnd.n1558 585
R4860 gnd.n1942 gnd.n1941 585
R4861 gnd.n1942 gnd.n1571 585
R4862 gnd.n1943 gnd.n1932 585
R4863 gnd.n1943 gnd.n1568 585
R4864 gnd.n1945 gnd.n1944 585
R4865 gnd.n1944 gnd.n1582 585
R4866 gnd.n1946 gnd.n1927 585
R4867 gnd.n1927 gnd.n1591 585
R4868 gnd.n1948 gnd.n1947 585
R4869 gnd.n1948 gnd.n1589 585
R4870 gnd.n1949 gnd.n1926 585
R4871 gnd.n1949 gnd.n1602 585
R4872 gnd.n1951 gnd.n1950 585
R4873 gnd.n1950 gnd.n1599 585
R4874 gnd.n1952 gnd.n1921 585
R4875 gnd.n1921 gnd.n1611 585
R4876 gnd.n1954 gnd.n1953 585
R4877 gnd.n1954 gnd.n1620 585
R4878 gnd.n1955 gnd.n1920 585
R4879 gnd.n1955 gnd.n1618 585
R4880 gnd.n1957 gnd.n1956 585
R4881 gnd.n1956 gnd.n1637 585
R4882 gnd.n1958 gnd.n1917 585
R4883 gnd.n1917 gnd.n1634 585
R4884 gnd.n1960 gnd.n1959 585
R4885 gnd.n1960 gnd.n1657 585
R4886 gnd.n1961 gnd.n1916 585
R4887 gnd.n1961 gnd.n1654 585
R4888 gnd.n1963 gnd.n1962 585
R4889 gnd.n1962 gnd.n1652 585
R4890 gnd.n1965 gnd.n1914 585
R4891 gnd.n1914 gnd.n1662 585
R4892 gnd.n1967 gnd.n1966 585
R4893 gnd.n1967 gnd.n1670 585
R4894 gnd.n1968 gnd.n1913 585
R4895 gnd.n1968 gnd.n1668 585
R4896 gnd.n1970 gnd.n1969 585
R4897 gnd.n1969 gnd.n1679 585
R4898 gnd.n1971 gnd.n1912 585
R4899 gnd.n1912 gnd.n1685 585
R4900 gnd.n1973 gnd.n1687 585
R4901 gnd.n6860 gnd.n6859 585
R4902 gnd.n6861 gnd.n6860 585
R4903 gnd.n767 gnd.n765 585
R4904 gnd.n6831 gnd.n765 585
R4905 gnd.n6829 gnd.n6828 585
R4906 gnd.n6830 gnd.n6829 585
R4907 gnd.n805 gnd.n804 585
R4908 gnd.n811 gnd.n804 585
R4909 gnd.n6824 gnd.n6823 585
R4910 gnd.n6823 gnd.n6822 585
R4911 gnd.n808 gnd.n807 585
R4912 gnd.n6809 gnd.n808 585
R4913 gnd.n829 gnd.n827 585
R4914 gnd.n827 gnd.n817 585
R4915 gnd.n6794 gnd.n6793 585
R4916 gnd.n6795 gnd.n6794 585
R4917 gnd.n828 gnd.n826 585
R4918 gnd.n835 gnd.n826 585
R4919 gnd.n6788 gnd.n6787 585
R4920 gnd.n6787 gnd.n6786 585
R4921 gnd.n832 gnd.n831 585
R4922 gnd.n6774 gnd.n832 585
R4923 gnd.n854 gnd.n852 585
R4924 gnd.n852 gnd.n851 585
R4925 gnd.n6764 gnd.n6763 585
R4926 gnd.n6765 gnd.n6764 585
R4927 gnd.n853 gnd.n850 585
R4928 gnd.n860 gnd.n850 585
R4929 gnd.n6758 gnd.n6757 585
R4930 gnd.n6757 gnd.n6756 585
R4931 gnd.n857 gnd.n856 585
R4932 gnd.n6744 gnd.n857 585
R4933 gnd.n879 gnd.n877 585
R4934 gnd.n877 gnd.n876 585
R4935 gnd.n6734 gnd.n6733 585
R4936 gnd.n6735 gnd.n6734 585
R4937 gnd.n878 gnd.n875 585
R4938 gnd.n884 gnd.n875 585
R4939 gnd.n6728 gnd.n6727 585
R4940 gnd.n6727 gnd.n6726 585
R4941 gnd.n882 gnd.n881 585
R4942 gnd.n6714 gnd.n882 585
R4943 gnd.n6523 gnd.n6521 585
R4944 gnd.n6521 gnd.n933 585
R4945 gnd.n6524 gnd.n6520 585
R4946 gnd.n6520 gnd.n6519 585
R4947 gnd.n6525 gnd.n960 585
R4948 gnd.n960 gnd.n938 585
R4949 gnd.n957 gnd.n948 585
R4950 gnd.n6538 gnd.n948 585
R4951 gnd.n6530 gnd.n6529 585
R4952 gnd.n6531 gnd.n6530 585
R4953 gnd.n956 gnd.n955 585
R4954 gnd.n6480 gnd.n955 585
R4955 gnd.n977 gnd.n975 585
R4956 gnd.n995 gnd.n975 585
R4957 gnd.n6498 gnd.n6497 585
R4958 gnd.n6499 gnd.n6498 585
R4959 gnd.n976 gnd.n974 585
R4960 gnd.n1000 gnd.n974 585
R4961 gnd.n6492 gnd.n6491 585
R4962 gnd.n6491 gnd.n6490 585
R4963 gnd.n980 gnd.n979 585
R4964 gnd.n1005 gnd.n980 585
R4965 gnd.n6440 gnd.n6439 585
R4966 gnd.n6441 gnd.n6440 585
R4967 gnd.n1016 gnd.n1015 585
R4968 gnd.n1039 gnd.n1015 585
R4969 gnd.n6435 gnd.n6434 585
R4970 gnd.n6434 gnd.n6433 585
R4971 gnd.n1019 gnd.n1018 585
R4972 gnd.n1026 gnd.n1019 585
R4973 gnd.n6404 gnd.n6403 585
R4974 gnd.n6405 gnd.n6404 585
R4975 gnd.n1045 gnd.n1044 585
R4976 gnd.n1066 gnd.n1044 585
R4977 gnd.n6399 gnd.n6398 585
R4978 gnd.n6398 gnd.n6397 585
R4979 gnd.n1048 gnd.n1047 585
R4980 gnd.n1057 gnd.n1048 585
R4981 gnd.n6367 gnd.n6366 585
R4982 gnd.n6368 gnd.n6367 585
R4983 gnd.n1072 gnd.n1071 585
R4984 gnd.n6341 gnd.n1071 585
R4985 gnd.n6362 gnd.n6361 585
R4986 gnd.n6361 gnd.n6360 585
R4987 gnd.n1075 gnd.n1074 585
R4988 gnd.n6349 gnd.n1075 585
R4989 gnd.n6305 gnd.n6304 585
R4990 gnd.n6306 gnd.n6305 585
R4991 gnd.n1103 gnd.n1102 585
R4992 gnd.n6279 gnd.n1102 585
R4993 gnd.n6300 gnd.n6299 585
R4994 gnd.n6299 gnd.n6298 585
R4995 gnd.n1106 gnd.n1105 585
R4996 gnd.n6287 gnd.n1106 585
R4997 gnd.n6259 gnd.n6258 585
R4998 gnd.n6260 gnd.n6259 585
R4999 gnd.n1131 gnd.n1130 585
R5000 gnd.n6233 gnd.n1130 585
R5001 gnd.n6254 gnd.n6253 585
R5002 gnd.n6253 gnd.n6252 585
R5003 gnd.n1134 gnd.n1133 585
R5004 gnd.n6241 gnd.n1134 585
R5005 gnd.n6186 gnd.n6184 585
R5006 gnd.n6184 gnd.n1152 585
R5007 gnd.n6187 gnd.n6183 585
R5008 gnd.n6183 gnd.n1157 585
R5009 gnd.n6188 gnd.n6182 585
R5010 gnd.n6182 gnd.n1167 585
R5011 gnd.n1180 gnd.n1178 585
R5012 gnd.n1178 gnd.n1164 585
R5013 gnd.n6193 gnd.n6192 585
R5014 gnd.n6194 gnd.n6193 585
R5015 gnd.n1179 gnd.n1177 585
R5016 gnd.n6145 gnd.n1177 585
R5017 gnd.n6178 gnd.n6177 585
R5018 gnd.n6177 gnd.n6176 585
R5019 gnd.n1183 gnd.n1182 585
R5020 gnd.n6164 gnd.n1183 585
R5021 gnd.n1222 gnd.n1220 585
R5022 gnd.n1220 gnd.n1201 585
R5023 gnd.n6108 gnd.n6107 585
R5024 gnd.n6109 gnd.n6108 585
R5025 gnd.n1221 gnd.n1219 585
R5026 gnd.n1261 gnd.n1219 585
R5027 gnd.n6102 gnd.n6101 585
R5028 gnd.n6101 gnd.n6100 585
R5029 gnd.n1225 gnd.n1224 585
R5030 gnd.n5505 gnd.n1225 585
R5031 gnd.n5656 gnd.n5654 585
R5032 gnd.n5654 gnd.n5653 585
R5033 gnd.n5657 gnd.n5502 585
R5034 gnd.n5638 gnd.n5502 585
R5035 gnd.n5658 gnd.n5501 585
R5036 gnd.n5512 gnd.n5501 585
R5037 gnd.n5620 gnd.n5499 585
R5038 gnd.n5621 gnd.n5620 585
R5039 gnd.n5662 gnd.n5498 585
R5040 gnd.n5519 gnd.n5498 585
R5041 gnd.n5663 gnd.n5497 585
R5042 gnd.n5609 gnd.n5497 585
R5043 gnd.n5664 gnd.n5496 585
R5044 gnd.n5525 gnd.n5496 585
R5045 gnd.n5599 gnd.n5494 585
R5046 gnd.n5600 gnd.n5599 585
R5047 gnd.n5668 gnd.n5493 585
R5048 gnd.n5531 gnd.n5493 585
R5049 gnd.n5669 gnd.n5492 585
R5050 gnd.n5588 gnd.n5492 585
R5051 gnd.n5670 gnd.n5491 585
R5052 gnd.n5537 gnd.n5491 585
R5053 gnd.n5578 gnd.n5489 585
R5054 gnd.n5579 gnd.n5578 585
R5055 gnd.n5674 gnd.n5488 585
R5056 gnd.n5543 gnd.n5488 585
R5057 gnd.n5675 gnd.n5487 585
R5058 gnd.n5567 gnd.n5487 585
R5059 gnd.n5676 gnd.n5486 585
R5060 gnd.n5550 gnd.n5486 585
R5061 gnd.n5483 gnd.n5481 585
R5062 gnd.n5558 gnd.n5481 585
R5063 gnd.n5681 gnd.n5680 585
R5064 gnd.n5682 gnd.n5681 585
R5065 gnd.n5482 gnd.n1477 585
R5066 gnd.n5478 gnd.n1477 585
R5067 gnd.n5836 gnd.n5835 585
R5068 gnd.n5834 gnd.n1476 585
R5069 gnd.n1479 gnd.n1475 585
R5070 gnd.n5838 gnd.n1475 585
R5071 gnd.n5830 gnd.n1481 585
R5072 gnd.n5829 gnd.n1482 585
R5073 gnd.n5828 gnd.n1483 585
R5074 gnd.n5825 gnd.n1484 585
R5075 gnd.n5824 gnd.n1485 585
R5076 gnd.n5704 gnd.n1486 585
R5077 gnd.n5706 gnd.n5705 585
R5078 gnd.n5816 gnd.n5707 585
R5079 gnd.n5815 gnd.n5708 585
R5080 gnd.n5718 gnd.n5709 585
R5081 gnd.n5808 gnd.n5719 585
R5082 gnd.n5807 gnd.n5720 585
R5083 gnd.n5722 gnd.n5721 585
R5084 gnd.n5800 gnd.n5730 585
R5085 gnd.n5799 gnd.n5731 585
R5086 gnd.n5741 gnd.n5732 585
R5087 gnd.n5792 gnd.n5742 585
R5088 gnd.n5791 gnd.n5743 585
R5089 gnd.n5745 gnd.n5744 585
R5090 gnd.n5784 gnd.n5753 585
R5091 gnd.n5783 gnd.n5754 585
R5092 gnd.n5774 gnd.n5755 585
R5093 gnd.n5776 gnd.n5775 585
R5094 gnd.n1472 gnd.n1457 585
R5095 gnd.n5842 gnd.n1458 585
R5096 gnd.n5841 gnd.n5840 585
R5097 gnd.n6863 gnd.n6862 585
R5098 gnd.n6862 gnd.n6861 585
R5099 gnd.n761 gnd.n760 585
R5100 gnd.n6831 gnd.n761 585
R5101 gnd.n6802 gnd.n803 585
R5102 gnd.n6830 gnd.n803 585
R5103 gnd.n6803 gnd.n6801 585
R5104 gnd.n6801 gnd.n811 585
R5105 gnd.n820 gnd.n810 585
R5106 gnd.n6822 gnd.n810 585
R5107 gnd.n6808 gnd.n6807 585
R5108 gnd.n6809 gnd.n6808 585
R5109 gnd.n819 gnd.n818 585
R5110 gnd.n818 gnd.n817 585
R5111 gnd.n6797 gnd.n6796 585
R5112 gnd.n6796 gnd.n6795 585
R5113 gnd.n823 gnd.n822 585
R5114 gnd.n835 gnd.n823 585
R5115 gnd.n844 gnd.n834 585
R5116 gnd.n6786 gnd.n834 585
R5117 gnd.n6773 gnd.n6772 585
R5118 gnd.n6774 gnd.n6773 585
R5119 gnd.n843 gnd.n842 585
R5120 gnd.n851 gnd.n842 585
R5121 gnd.n6767 gnd.n6766 585
R5122 gnd.n6766 gnd.n6765 585
R5123 gnd.n847 gnd.n846 585
R5124 gnd.n860 gnd.n847 585
R5125 gnd.n869 gnd.n859 585
R5126 gnd.n6756 gnd.n859 585
R5127 gnd.n6743 gnd.n6742 585
R5128 gnd.n6744 gnd.n6743 585
R5129 gnd.n868 gnd.n867 585
R5130 gnd.n876 gnd.n867 585
R5131 gnd.n6737 gnd.n6736 585
R5132 gnd.n6736 gnd.n6735 585
R5133 gnd.n872 gnd.n871 585
R5134 gnd.n884 gnd.n872 585
R5135 gnd.n6511 gnd.n883 585
R5136 gnd.n6726 gnd.n883 585
R5137 gnd.n6512 gnd.n892 585
R5138 gnd.n6714 gnd.n892 585
R5139 gnd.n964 gnd.n962 585
R5140 gnd.n962 gnd.n933 585
R5141 gnd.n6517 gnd.n6516 585
R5142 gnd.n6519 gnd.n6517 585
R5143 gnd.n963 gnd.n961 585
R5144 gnd.n961 gnd.n938 585
R5145 gnd.n6507 gnd.n947 585
R5146 gnd.n6538 gnd.n947 585
R5147 gnd.n6506 gnd.n954 585
R5148 gnd.n6531 gnd.n954 585
R5149 gnd.n6505 gnd.n967 585
R5150 gnd.n6480 gnd.n967 585
R5151 gnd.n971 gnd.n966 585
R5152 gnd.n995 gnd.n971 585
R5153 gnd.n6501 gnd.n6500 585
R5154 gnd.n6500 gnd.n6499 585
R5155 gnd.n970 gnd.n969 585
R5156 gnd.n1000 gnd.n970 585
R5157 gnd.n6322 gnd.n982 585
R5158 gnd.n6490 gnd.n982 585
R5159 gnd.n6323 gnd.n6321 585
R5160 gnd.n6321 gnd.n1005 585
R5161 gnd.n6319 gnd.n1012 585
R5162 gnd.n6441 gnd.n1012 585
R5163 gnd.n6327 gnd.n6318 585
R5164 gnd.n6318 gnd.n1039 585
R5165 gnd.n6328 gnd.n1020 585
R5166 gnd.n6433 gnd.n1020 585
R5167 gnd.n6329 gnd.n6317 585
R5168 gnd.n6317 gnd.n1026 585
R5169 gnd.n6315 gnd.n1043 585
R5170 gnd.n6405 gnd.n1043 585
R5171 gnd.n6333 gnd.n6314 585
R5172 gnd.n6314 gnd.n1066 585
R5173 gnd.n6334 gnd.n1050 585
R5174 gnd.n6397 gnd.n1050 585
R5175 gnd.n6335 gnd.n6313 585
R5176 gnd.n6313 gnd.n1057 585
R5177 gnd.n1095 gnd.n1070 585
R5178 gnd.n6368 gnd.n1070 585
R5179 gnd.n6340 gnd.n6339 585
R5180 gnd.n6341 gnd.n6340 585
R5181 gnd.n1094 gnd.n1077 585
R5182 gnd.n6360 gnd.n1077 585
R5183 gnd.n6309 gnd.n1085 585
R5184 gnd.n6349 gnd.n1085 585
R5185 gnd.n6308 gnd.n6307 585
R5186 gnd.n6307 gnd.n6306 585
R5187 gnd.n1098 gnd.n1097 585
R5188 gnd.n6279 gnd.n1098 585
R5189 gnd.n6126 gnd.n1107 585
R5190 gnd.n6298 gnd.n1107 585
R5191 gnd.n6127 gnd.n1116 585
R5192 gnd.n6287 gnd.n1116 585
R5193 gnd.n6123 gnd.n1129 585
R5194 gnd.n6260 gnd.n1129 585
R5195 gnd.n6131 gnd.n1146 585
R5196 gnd.n6233 gnd.n1146 585
R5197 gnd.n6132 gnd.n1136 585
R5198 gnd.n6252 gnd.n1136 585
R5199 gnd.n6133 gnd.n1143 585
R5200 gnd.n6241 gnd.n1143 585
R5201 gnd.n6121 gnd.n6120 585
R5202 gnd.n6120 gnd.n1152 585
R5203 gnd.n6137 gnd.n6119 585
R5204 gnd.n6119 gnd.n1157 585
R5205 gnd.n6138 gnd.n6118 585
R5206 gnd.n6118 gnd.n1167 585
R5207 gnd.n6139 gnd.n6117 585
R5208 gnd.n6117 gnd.n1164 585
R5209 gnd.n1214 gnd.n1175 585
R5210 gnd.n6194 gnd.n1175 585
R5211 gnd.n6144 gnd.n6143 585
R5212 gnd.n6145 gnd.n6144 585
R5213 gnd.n1213 gnd.n1185 585
R5214 gnd.n6176 gnd.n1185 585
R5215 gnd.n6113 gnd.n1193 585
R5216 gnd.n6164 gnd.n1193 585
R5217 gnd.n6112 gnd.n6111 585
R5218 gnd.n6111 gnd.n1201 585
R5219 gnd.n6110 gnd.n1216 585
R5220 gnd.n6110 gnd.n6109 585
R5221 gnd.n5630 gnd.n1217 585
R5222 gnd.n1261 gnd.n1217 585
R5223 gnd.n5631 gnd.n1227 585
R5224 gnd.n6100 gnd.n1227 585
R5225 gnd.n5632 gnd.n5627 585
R5226 gnd.n5627 gnd.n5505 585
R5227 gnd.n5515 gnd.n5504 585
R5228 gnd.n5653 gnd.n5504 585
R5229 gnd.n5637 gnd.n5636 585
R5230 gnd.n5638 gnd.n5637 585
R5231 gnd.n5514 gnd.n5513 585
R5232 gnd.n5513 gnd.n5512 585
R5233 gnd.n5623 gnd.n5622 585
R5234 gnd.n5622 gnd.n5621 585
R5235 gnd.n5518 gnd.n5517 585
R5236 gnd.n5519 gnd.n5518 585
R5237 gnd.n5607 gnd.n5606 585
R5238 gnd.n5609 gnd.n5607 585
R5239 gnd.n5527 gnd.n5526 585
R5240 gnd.n5526 gnd.n5525 585
R5241 gnd.n5602 gnd.n5601 585
R5242 gnd.n5601 gnd.n5600 585
R5243 gnd.n5530 gnd.n5529 585
R5244 gnd.n5531 gnd.n5530 585
R5245 gnd.n5586 gnd.n5585 585
R5246 gnd.n5588 gnd.n5586 585
R5247 gnd.n5539 gnd.n5538 585
R5248 gnd.n5538 gnd.n5537 585
R5249 gnd.n5581 gnd.n5580 585
R5250 gnd.n5580 gnd.n5579 585
R5251 gnd.n5542 gnd.n5541 585
R5252 gnd.n5543 gnd.n5542 585
R5253 gnd.n5565 gnd.n5564 585
R5254 gnd.n5567 gnd.n5565 585
R5255 gnd.n5552 gnd.n5551 585
R5256 gnd.n5551 gnd.n5550 585
R5257 gnd.n5560 gnd.n5559 585
R5258 gnd.n5559 gnd.n5558 585
R5259 gnd.n5556 gnd.n5479 585
R5260 gnd.n5682 gnd.n5479 585
R5261 gnd.n5555 gnd.n1459 585
R5262 gnd.n5478 gnd.n1459 585
R5263 gnd.n6881 gnd.n746 585
R5264 gnd.n6845 gnd.n746 585
R5265 gnd.n6882 gnd.n745 585
R5266 gnd.n791 gnd.n739 585
R5267 gnd.n6889 gnd.n738 585
R5268 gnd.n6890 gnd.n737 585
R5269 gnd.n788 gnd.n729 585
R5270 gnd.n6897 gnd.n728 585
R5271 gnd.n6898 gnd.n727 585
R5272 gnd.n786 gnd.n721 585
R5273 gnd.n6905 gnd.n720 585
R5274 gnd.n6906 gnd.n719 585
R5275 gnd.n783 gnd.n711 585
R5276 gnd.n6913 gnd.n710 585
R5277 gnd.n6914 gnd.n709 585
R5278 gnd.n781 gnd.n701 585
R5279 gnd.n6921 gnd.n700 585
R5280 gnd.n6922 gnd.n699 585
R5281 gnd.n6923 gnd.n698 585
R5282 gnd.n6847 gnd.n697 585
R5283 gnd.n6849 gnd.n6848 585
R5284 gnd.n6850 gnd.n774 585
R5285 gnd.n778 gnd.n772 585
R5286 gnd.n6854 gnd.n771 585
R5287 gnd.n6855 gnd.n770 585
R5288 gnd.n6856 gnd.n766 585
R5289 gnd.n762 gnd.n758 585
R5290 gnd.n6870 gnd.n757 585
R5291 gnd.n6871 gnd.n756 585
R5292 gnd.n793 gnd.n755 585
R5293 gnd.n1293 gnd.t29 543.808
R5294 gnd.n927 gnd.t25 543.808
R5295 gnd.n1290 gnd.t67 543.808
R5296 gnd.n6571 gnd.t64 543.808
R5297 gnd.n6637 gnd.n935 497.305
R5298 gnd.n6646 gnd.n6645 497.305
R5299 gnd.n1297 gnd.n1296 497.305
R5300 gnd.n6097 gnd.n1265 497.305
R5301 gnd.n3111 gnd.n3110 462.966
R5302 gnd.n5771 gnd.t18 371.625
R5303 gnd.n6875 gnd.t98 371.625
R5304 gnd.n5762 gnd.t117 371.625
R5305 gnd.n647 gnd.t95 371.625
R5306 gnd.n670 gnd.t89 371.625
R5307 gnd.n693 gnd.t32 371.625
R5308 gnd.n346 gnd.t123 371.625
R5309 gnd.n326 gnd.t40 371.625
R5310 gnd.n7625 gnd.t58 371.625
R5311 gnd.n7392 gnd.t76 371.625
R5312 gnd.n4867 gnd.t92 371.625
R5313 gnd.n4977 gnd.t36 371.625
R5314 gnd.n4823 gnd.t48 371.625
R5315 gnd.n4756 gnd.t120 371.625
R5316 gnd.n5900 gnd.t111 371.625
R5317 gnd.n1415 gnd.t44 371.625
R5318 gnd.n1382 gnd.t73 371.625
R5319 gnd.n747 gnd.t51 371.625
R5320 gnd.n3745 gnd.t82 323.425
R5321 gnd.n1858 gnd.t107 323.425
R5322 gnd.n4593 gnd.n4567 289.615
R5323 gnd.n4561 gnd.n4535 289.615
R5324 gnd.n4529 gnd.n4503 289.615
R5325 gnd.n4498 gnd.n4472 289.615
R5326 gnd.n4466 gnd.n4440 289.615
R5327 gnd.n4434 gnd.n4408 289.615
R5328 gnd.n4402 gnd.n4376 289.615
R5329 gnd.n4371 gnd.n4345 289.615
R5330 gnd.n3819 gnd.t14 279.217
R5331 gnd.n1884 gnd.t126 279.217
R5332 gnd.n1272 gnd.t106 260.649
R5333 gnd.n6563 gnd.t63 260.649
R5334 gnd.n6099 gnd.n6098 256.663
R5335 gnd.n6099 gnd.n1228 256.663
R5336 gnd.n6099 gnd.n1229 256.663
R5337 gnd.n6099 gnd.n1230 256.663
R5338 gnd.n6099 gnd.n1231 256.663
R5339 gnd.n6099 gnd.n1232 256.663
R5340 gnd.n6099 gnd.n1233 256.663
R5341 gnd.n6099 gnd.n1234 256.663
R5342 gnd.n6099 gnd.n1235 256.663
R5343 gnd.n6099 gnd.n1236 256.663
R5344 gnd.n6099 gnd.n1237 256.663
R5345 gnd.n6099 gnd.n1238 256.663
R5346 gnd.n6099 gnd.n1239 256.663
R5347 gnd.n6099 gnd.n1240 256.663
R5348 gnd.n6099 gnd.n1241 256.663
R5349 gnd.n6099 gnd.n1242 256.663
R5350 gnd.n6035 gnd.n6032 256.663
R5351 gnd.n6099 gnd.n1243 256.663
R5352 gnd.n6099 gnd.n1244 256.663
R5353 gnd.n6099 gnd.n1245 256.663
R5354 gnd.n6099 gnd.n1246 256.663
R5355 gnd.n6099 gnd.n1247 256.663
R5356 gnd.n6099 gnd.n1248 256.663
R5357 gnd.n6099 gnd.n1249 256.663
R5358 gnd.n6099 gnd.n1250 256.663
R5359 gnd.n6099 gnd.n1251 256.663
R5360 gnd.n6099 gnd.n1252 256.663
R5361 gnd.n6099 gnd.n1253 256.663
R5362 gnd.n6099 gnd.n1254 256.663
R5363 gnd.n6099 gnd.n1255 256.663
R5364 gnd.n6099 gnd.n1256 256.663
R5365 gnd.n6099 gnd.n1257 256.663
R5366 gnd.n6099 gnd.n1258 256.663
R5367 gnd.n6099 gnd.n1259 256.663
R5368 gnd.n6712 gnd.n910 256.663
R5369 gnd.n6712 gnd.n911 256.663
R5370 gnd.n6712 gnd.n912 256.663
R5371 gnd.n6712 gnd.n913 256.663
R5372 gnd.n6712 gnd.n914 256.663
R5373 gnd.n6712 gnd.n915 256.663
R5374 gnd.n6712 gnd.n916 256.663
R5375 gnd.n6712 gnd.n917 256.663
R5376 gnd.n6712 gnd.n918 256.663
R5377 gnd.n6712 gnd.n919 256.663
R5378 gnd.n6712 gnd.n920 256.663
R5379 gnd.n6712 gnd.n921 256.663
R5380 gnd.n6712 gnd.n922 256.663
R5381 gnd.n6712 gnd.n923 256.663
R5382 gnd.n6712 gnd.n924 256.663
R5383 gnd.n6712 gnd.n925 256.663
R5384 gnd.n926 gnd.n657 256.663
R5385 gnd.n6712 gnd.n909 256.663
R5386 gnd.n6712 gnd.n908 256.663
R5387 gnd.n6712 gnd.n907 256.663
R5388 gnd.n6712 gnd.n906 256.663
R5389 gnd.n6712 gnd.n905 256.663
R5390 gnd.n6712 gnd.n904 256.663
R5391 gnd.n6712 gnd.n903 256.663
R5392 gnd.n6712 gnd.n902 256.663
R5393 gnd.n6712 gnd.n901 256.663
R5394 gnd.n6712 gnd.n900 256.663
R5395 gnd.n6712 gnd.n899 256.663
R5396 gnd.n6712 gnd.n898 256.663
R5397 gnd.n6712 gnd.n897 256.663
R5398 gnd.n6712 gnd.n896 256.663
R5399 gnd.n6712 gnd.n895 256.663
R5400 gnd.n6712 gnd.n894 256.663
R5401 gnd.n6712 gnd.n893 256.663
R5402 gnd.n4817 gnd.n4727 242.672
R5403 gnd.n4815 gnd.n4727 242.672
R5404 gnd.n4809 gnd.n4727 242.672
R5405 gnd.n4807 gnd.n4727 242.672
R5406 gnd.n4801 gnd.n4727 242.672
R5407 gnd.n4799 gnd.n4727 242.672
R5408 gnd.n4793 gnd.n4727 242.672
R5409 gnd.n4791 gnd.n4727 242.672
R5410 gnd.n4781 gnd.n4727 242.672
R5411 gnd.n5765 gnd.n1369 242.672
R5412 gnd.n5760 gnd.n1369 242.672
R5413 gnd.n5757 gnd.n1369 242.672
R5414 gnd.n5748 gnd.n1369 242.672
R5415 gnd.n5737 gnd.n1369 242.672
R5416 gnd.n5734 gnd.n1369 242.672
R5417 gnd.n5725 gnd.n1369 242.672
R5418 gnd.n5714 gnd.n1369 242.672
R5419 gnd.n5711 gnd.n1369 242.672
R5420 gnd.n3873 gnd.n3872 242.672
R5421 gnd.n3873 gnd.n3783 242.672
R5422 gnd.n3873 gnd.n3784 242.672
R5423 gnd.n3873 gnd.n3785 242.672
R5424 gnd.n3873 gnd.n3786 242.672
R5425 gnd.n3873 gnd.n3787 242.672
R5426 gnd.n3873 gnd.n3788 242.672
R5427 gnd.n3873 gnd.n3789 242.672
R5428 gnd.n3873 gnd.n3790 242.672
R5429 gnd.n3873 gnd.n3791 242.672
R5430 gnd.n3873 gnd.n3792 242.672
R5431 gnd.n3873 gnd.n3793 242.672
R5432 gnd.n3874 gnd.n3873 242.672
R5433 gnd.n4726 gnd.n1833 242.672
R5434 gnd.n4726 gnd.n1832 242.672
R5435 gnd.n4726 gnd.n1831 242.672
R5436 gnd.n4726 gnd.n1830 242.672
R5437 gnd.n4726 gnd.n1829 242.672
R5438 gnd.n4726 gnd.n1828 242.672
R5439 gnd.n4726 gnd.n1827 242.672
R5440 gnd.n4726 gnd.n1826 242.672
R5441 gnd.n4726 gnd.n1825 242.672
R5442 gnd.n4726 gnd.n1824 242.672
R5443 gnd.n4726 gnd.n1823 242.672
R5444 gnd.n4726 gnd.n1822 242.672
R5445 gnd.n4726 gnd.n1821 242.672
R5446 gnd.n7041 gnd.n618 242.672
R5447 gnd.n7041 gnd.n619 242.672
R5448 gnd.n7041 gnd.n620 242.672
R5449 gnd.n7041 gnd.n621 242.672
R5450 gnd.n7041 gnd.n622 242.672
R5451 gnd.n7041 gnd.n623 242.672
R5452 gnd.n7041 gnd.n624 242.672
R5453 gnd.n7041 gnd.n625 242.672
R5454 gnd.n7041 gnd.n626 242.672
R5455 gnd.n7660 gnd.n260 242.672
R5456 gnd.n7660 gnd.n259 242.672
R5457 gnd.n7660 gnd.n258 242.672
R5458 gnd.n7660 gnd.n257 242.672
R5459 gnd.n7660 gnd.n256 242.672
R5460 gnd.n7660 gnd.n255 242.672
R5461 gnd.n7660 gnd.n254 242.672
R5462 gnd.n7660 gnd.n253 242.672
R5463 gnd.n7660 gnd.n252 242.672
R5464 gnd.n3957 gnd.n3956 242.672
R5465 gnd.n3956 gnd.n3695 242.672
R5466 gnd.n3956 gnd.n3696 242.672
R5467 gnd.n3956 gnd.n3697 242.672
R5468 gnd.n3956 gnd.n3698 242.672
R5469 gnd.n3956 gnd.n3699 242.672
R5470 gnd.n3956 gnd.n3700 242.672
R5471 gnd.n3956 gnd.n3701 242.672
R5472 gnd.n4726 gnd.n1834 242.672
R5473 gnd.n4726 gnd.n1835 242.672
R5474 gnd.n4726 gnd.n1836 242.672
R5475 gnd.n4726 gnd.n1837 242.672
R5476 gnd.n4726 gnd.n1838 242.672
R5477 gnd.n4726 gnd.n1839 242.672
R5478 gnd.n4726 gnd.n1840 242.672
R5479 gnd.n4726 gnd.n1841 242.672
R5480 gnd.n4885 gnd.n4727 242.672
R5481 gnd.n4893 gnd.n4727 242.672
R5482 gnd.n4895 gnd.n4727 242.672
R5483 gnd.n4903 gnd.n4727 242.672
R5484 gnd.n4905 gnd.n4727 242.672
R5485 gnd.n4913 gnd.n4727 242.672
R5486 gnd.n4915 gnd.n4727 242.672
R5487 gnd.n4923 gnd.n4727 242.672
R5488 gnd.n4925 gnd.n4727 242.672
R5489 gnd.n4933 gnd.n4727 242.672
R5490 gnd.n4935 gnd.n4727 242.672
R5491 gnd.n4943 gnd.n4727 242.672
R5492 gnd.n4945 gnd.n4727 242.672
R5493 gnd.n4953 gnd.n4727 242.672
R5494 gnd.n4955 gnd.n4727 242.672
R5495 gnd.n4963 gnd.n4727 242.672
R5496 gnd.n4965 gnd.n4727 242.672
R5497 gnd.n4973 gnd.n4727 242.672
R5498 gnd.n4975 gnd.n4727 242.672
R5499 gnd.n4985 gnd.n4727 242.672
R5500 gnd.n4987 gnd.n4727 242.672
R5501 gnd.n4995 gnd.n4727 242.672
R5502 gnd.n4997 gnd.n4727 242.672
R5503 gnd.n5005 gnd.n4727 242.672
R5504 gnd.n5007 gnd.n4727 242.672
R5505 gnd.n5015 gnd.n4727 242.672
R5506 gnd.n5017 gnd.n4727 242.672
R5507 gnd.n5026 gnd.n4727 242.672
R5508 gnd.n5029 gnd.n4727 242.672
R5509 gnd.n5975 gnd.n1369 242.672
R5510 gnd.n1418 gnd.n1369 242.672
R5511 gnd.n5982 gnd.n1369 242.672
R5512 gnd.n1409 gnd.n1369 242.672
R5513 gnd.n5989 gnd.n1369 242.672
R5514 gnd.n1402 gnd.n1369 242.672
R5515 gnd.n5996 gnd.n1369 242.672
R5516 gnd.n1395 gnd.n1369 242.672
R5517 gnd.n6003 gnd.n1369 242.672
R5518 gnd.n6006 gnd.n1369 242.672
R5519 gnd.n1386 gnd.n1369 242.672
R5520 gnd.n6015 gnd.n1369 242.672
R5521 gnd.n1377 gnd.n1369 242.672
R5522 gnd.n6022 gnd.n1369 242.672
R5523 gnd.n6025 gnd.n1369 242.672
R5524 gnd.n1369 gnd.n1368 242.672
R5525 gnd.n6031 gnd.n1363 242.672
R5526 gnd.n5915 gnd.n1369 242.672
R5527 gnd.n5914 gnd.n1369 242.672
R5528 gnd.n5922 gnd.n1369 242.672
R5529 gnd.n5908 gnd.n1369 242.672
R5530 gnd.n5929 gnd.n1369 242.672
R5531 gnd.n5898 gnd.n1369 242.672
R5532 gnd.n5936 gnd.n1369 242.672
R5533 gnd.n5891 gnd.n1369 242.672
R5534 gnd.n5943 gnd.n1369 242.672
R5535 gnd.n5884 gnd.n1369 242.672
R5536 gnd.n5950 gnd.n1369 242.672
R5537 gnd.n5877 gnd.n1369 242.672
R5538 gnd.n5957 gnd.n1369 242.672
R5539 gnd.n7041 gnd.n7040 242.672
R5540 gnd.n7041 gnd.n590 242.672
R5541 gnd.n7041 gnd.n591 242.672
R5542 gnd.n7041 gnd.n592 242.672
R5543 gnd.n7041 gnd.n593 242.672
R5544 gnd.n7041 gnd.n594 242.672
R5545 gnd.n7041 gnd.n595 242.672
R5546 gnd.n7041 gnd.n596 242.672
R5547 gnd.n7041 gnd.n597 242.672
R5548 gnd.n7041 gnd.n598 242.672
R5549 gnd.n7041 gnd.n599 242.672
R5550 gnd.n7041 gnd.n600 242.672
R5551 gnd.n7041 gnd.n601 242.672
R5552 gnd.n6989 gnd.n658 242.672
R5553 gnd.n7041 gnd.n602 242.672
R5554 gnd.n7041 gnd.n603 242.672
R5555 gnd.n7041 gnd.n604 242.672
R5556 gnd.n7041 gnd.n605 242.672
R5557 gnd.n7041 gnd.n606 242.672
R5558 gnd.n7041 gnd.n607 242.672
R5559 gnd.n7041 gnd.n608 242.672
R5560 gnd.n7041 gnd.n609 242.672
R5561 gnd.n7041 gnd.n610 242.672
R5562 gnd.n7041 gnd.n611 242.672
R5563 gnd.n7041 gnd.n612 242.672
R5564 gnd.n7041 gnd.n613 242.672
R5565 gnd.n7041 gnd.n614 242.672
R5566 gnd.n7041 gnd.n615 242.672
R5567 gnd.n7041 gnd.n616 242.672
R5568 gnd.n7041 gnd.n617 242.672
R5569 gnd.n7660 gnd.n261 242.672
R5570 gnd.n7660 gnd.n262 242.672
R5571 gnd.n7660 gnd.n263 242.672
R5572 gnd.n7660 gnd.n264 242.672
R5573 gnd.n7660 gnd.n265 242.672
R5574 gnd.n7660 gnd.n266 242.672
R5575 gnd.n7660 gnd.n267 242.672
R5576 gnd.n7660 gnd.n268 242.672
R5577 gnd.n7660 gnd.n269 242.672
R5578 gnd.n7660 gnd.n270 242.672
R5579 gnd.n7660 gnd.n271 242.672
R5580 gnd.n7660 gnd.n272 242.672
R5581 gnd.n7660 gnd.n273 242.672
R5582 gnd.n7660 gnd.n274 242.672
R5583 gnd.n7660 gnd.n275 242.672
R5584 gnd.n7660 gnd.n276 242.672
R5585 gnd.n7660 gnd.n277 242.672
R5586 gnd.n7660 gnd.n278 242.672
R5587 gnd.n7660 gnd.n279 242.672
R5588 gnd.n7660 gnd.n280 242.672
R5589 gnd.n7660 gnd.n281 242.672
R5590 gnd.n7660 gnd.n282 242.672
R5591 gnd.n7660 gnd.n283 242.672
R5592 gnd.n7660 gnd.n284 242.672
R5593 gnd.n7660 gnd.n285 242.672
R5594 gnd.n7660 gnd.n286 242.672
R5595 gnd.n7660 gnd.n287 242.672
R5596 gnd.n7660 gnd.n288 242.672
R5597 gnd.n7660 gnd.n7659 242.672
R5598 gnd.n5838 gnd.n5837 242.672
R5599 gnd.n5838 gnd.n1461 242.672
R5600 gnd.n5838 gnd.n1462 242.672
R5601 gnd.n5838 gnd.n1463 242.672
R5602 gnd.n5838 gnd.n1464 242.672
R5603 gnd.n5838 gnd.n1465 242.672
R5604 gnd.n5838 gnd.n1466 242.672
R5605 gnd.n5838 gnd.n1467 242.672
R5606 gnd.n5838 gnd.n1468 242.672
R5607 gnd.n5838 gnd.n1469 242.672
R5608 gnd.n5838 gnd.n1470 242.672
R5609 gnd.n5838 gnd.n1471 242.672
R5610 gnd.n5838 gnd.n1473 242.672
R5611 gnd.n5839 gnd.n5838 242.672
R5612 gnd.n6845 gnd.n792 242.672
R5613 gnd.n6845 gnd.n790 242.672
R5614 gnd.n6845 gnd.n789 242.672
R5615 gnd.n6845 gnd.n787 242.672
R5616 gnd.n6845 gnd.n785 242.672
R5617 gnd.n6845 gnd.n784 242.672
R5618 gnd.n6845 gnd.n782 242.672
R5619 gnd.n6845 gnd.n780 242.672
R5620 gnd.n6846 gnd.n6845 242.672
R5621 gnd.n6845 gnd.n775 242.672
R5622 gnd.n6845 gnd.n779 242.672
R5623 gnd.n6845 gnd.n777 242.672
R5624 gnd.n6845 gnd.n795 242.672
R5625 gnd.n6845 gnd.n794 242.672
R5626 gnd.n7661 gnd.n250 240.244
R5627 gnd.n7658 gnd.n289 240.244
R5628 gnd.n7654 gnd.n7653 240.244
R5629 gnd.n7650 gnd.n7649 240.244
R5630 gnd.n7646 gnd.n7645 240.244
R5631 gnd.n7642 gnd.n7641 240.244
R5632 gnd.n7638 gnd.n7637 240.244
R5633 gnd.n7634 gnd.n7633 240.244
R5634 gnd.n7630 gnd.n7629 240.244
R5635 gnd.n7623 gnd.n7622 240.244
R5636 gnd.n7619 gnd.n7618 240.244
R5637 gnd.n7615 gnd.n7614 240.244
R5638 gnd.n7611 gnd.n7610 240.244
R5639 gnd.n7607 gnd.n7606 240.244
R5640 gnd.n7603 gnd.n7602 240.244
R5641 gnd.n7599 gnd.n7598 240.244
R5642 gnd.n7595 gnd.n7594 240.244
R5643 gnd.n7591 gnd.n7590 240.244
R5644 gnd.n7587 gnd.n7586 240.244
R5645 gnd.n7580 gnd.n7579 240.244
R5646 gnd.n7577 gnd.n7576 240.244
R5647 gnd.n7573 gnd.n7572 240.244
R5648 gnd.n7569 gnd.n7568 240.244
R5649 gnd.n7565 gnd.n7564 240.244
R5650 gnd.n7561 gnd.n7560 240.244
R5651 gnd.n7557 gnd.n7556 240.244
R5652 gnd.n7553 gnd.n7552 240.244
R5653 gnd.n7549 gnd.n7548 240.244
R5654 gnd.n7545 gnd.n7544 240.244
R5655 gnd.n7061 gnd.n570 240.244
R5656 gnd.n7061 gnd.n561 240.244
R5657 gnd.n561 gnd.n553 240.244
R5658 gnd.n7088 gnd.n553 240.244
R5659 gnd.n7088 gnd.n532 240.244
R5660 gnd.n7098 gnd.n532 240.244
R5661 gnd.n7098 gnd.n522 240.244
R5662 gnd.n542 gnd.n522 240.244
R5663 gnd.n7093 gnd.n542 240.244
R5664 gnd.n7093 gnd.n497 240.244
R5665 gnd.n506 gnd.n497 240.244
R5666 gnd.n506 gnd.n488 240.244
R5667 gnd.n7145 gnd.n488 240.244
R5668 gnd.n7145 gnd.n467 240.244
R5669 gnd.n510 gnd.n467 240.244
R5670 gnd.n510 gnd.n457 240.244
R5671 gnd.n457 gnd.n449 240.244
R5672 gnd.n7217 gnd.n449 240.244
R5673 gnd.n7217 gnd.n440 240.244
R5674 gnd.n7220 gnd.n440 240.244
R5675 gnd.n7220 gnd.n422 240.244
R5676 gnd.n7259 gnd.n422 240.244
R5677 gnd.n7259 gnd.n412 240.244
R5678 gnd.n7263 gnd.n412 240.244
R5679 gnd.n7263 gnd.n403 240.244
R5680 gnd.n403 gnd.n394 240.244
R5681 gnd.n7300 gnd.n394 240.244
R5682 gnd.n7300 gnd.n388 240.244
R5683 gnd.n388 gnd.n377 240.244
R5684 gnd.n7324 gnd.n377 240.244
R5685 gnd.n7324 gnd.n366 240.244
R5686 gnd.n7336 gnd.n366 240.244
R5687 gnd.n7336 gnd.n361 240.244
R5688 gnd.n361 gnd.n101 240.244
R5689 gnd.n352 gnd.n101 240.244
R5690 gnd.n7359 gnd.n352 240.244
R5691 gnd.n7359 gnd.n118 240.244
R5692 gnd.n7491 gnd.n118 240.244
R5693 gnd.n7491 gnd.n129 240.244
R5694 gnd.n7495 gnd.n129 240.244
R5695 gnd.n7495 gnd.n138 240.244
R5696 gnd.n7498 gnd.n138 240.244
R5697 gnd.n7498 gnd.n147 240.244
R5698 gnd.n7502 gnd.n147 240.244
R5699 gnd.n7502 gnd.n157 240.244
R5700 gnd.n7505 gnd.n157 240.244
R5701 gnd.n7505 gnd.n166 240.244
R5702 gnd.n7509 gnd.n166 240.244
R5703 gnd.n7509 gnd.n176 240.244
R5704 gnd.n7512 gnd.n176 240.244
R5705 gnd.n7512 gnd.n185 240.244
R5706 gnd.n7516 gnd.n185 240.244
R5707 gnd.n7516 gnd.n195 240.244
R5708 gnd.n7519 gnd.n195 240.244
R5709 gnd.n7519 gnd.n204 240.244
R5710 gnd.n7523 gnd.n204 240.244
R5711 gnd.n7523 gnd.n214 240.244
R5712 gnd.n7526 gnd.n214 240.244
R5713 gnd.n7526 gnd.n223 240.244
R5714 gnd.n7530 gnd.n223 240.244
R5715 gnd.n7530 gnd.n233 240.244
R5716 gnd.n7533 gnd.n233 240.244
R5717 gnd.n7533 gnd.n242 240.244
R5718 gnd.n7537 gnd.n242 240.244
R5719 gnd.n7039 gnd.n628 240.244
R5720 gnd.n7035 gnd.n628 240.244
R5721 gnd.n7033 gnd.n7032 240.244
R5722 gnd.n7029 gnd.n7028 240.244
R5723 gnd.n7025 gnd.n7024 240.244
R5724 gnd.n7021 gnd.n7020 240.244
R5725 gnd.n7017 gnd.n7016 240.244
R5726 gnd.n7013 gnd.n7012 240.244
R5727 gnd.n7009 gnd.n7008 240.244
R5728 gnd.n7004 gnd.n7003 240.244
R5729 gnd.n7000 gnd.n6999 240.244
R5730 gnd.n6996 gnd.n6995 240.244
R5731 gnd.n6992 gnd.n6991 240.244
R5732 gnd.n6987 gnd.n6986 240.244
R5733 gnd.n6983 gnd.n6982 240.244
R5734 gnd.n6979 gnd.n6978 240.244
R5735 gnd.n6975 gnd.n6974 240.244
R5736 gnd.n6971 gnd.n6970 240.244
R5737 gnd.n6967 gnd.n6966 240.244
R5738 gnd.n6963 gnd.n6962 240.244
R5739 gnd.n6959 gnd.n6958 240.244
R5740 gnd.n6955 gnd.n6954 240.244
R5741 gnd.n6951 gnd.n6950 240.244
R5742 gnd.n6947 gnd.n6946 240.244
R5743 gnd.n6943 gnd.n6942 240.244
R5744 gnd.n6939 gnd.n6938 240.244
R5745 gnd.n6935 gnd.n6934 240.244
R5746 gnd.n6931 gnd.n6930 240.244
R5747 gnd.n7069 gnd.n564 240.244
R5748 gnd.n7077 gnd.n564 240.244
R5749 gnd.n7077 gnd.n565 240.244
R5750 gnd.n565 gnd.n530 240.244
R5751 gnd.n7119 gnd.n530 240.244
R5752 gnd.n7119 gnd.n525 240.244
R5753 gnd.n7127 gnd.n525 240.244
R5754 gnd.n7127 gnd.n526 240.244
R5755 gnd.n526 gnd.n496 240.244
R5756 gnd.n7154 gnd.n496 240.244
R5757 gnd.n7154 gnd.n492 240.244
R5758 gnd.n7160 gnd.n492 240.244
R5759 gnd.n7160 gnd.n465 240.244
R5760 gnd.n7189 gnd.n465 240.244
R5761 gnd.n7189 gnd.n460 240.244
R5762 gnd.n7197 gnd.n460 240.244
R5763 gnd.n7197 gnd.n461 240.244
R5764 gnd.n461 gnd.n438 240.244
R5765 gnd.n7229 gnd.n438 240.244
R5766 gnd.n7229 gnd.n434 240.244
R5767 gnd.n7235 gnd.n434 240.244
R5768 gnd.n7235 gnd.n411 240.244
R5769 gnd.n7276 gnd.n411 240.244
R5770 gnd.n7276 gnd.n406 240.244
R5771 gnd.n7284 gnd.n406 240.244
R5772 gnd.n7284 gnd.n407 240.244
R5773 gnd.n407 gnd.n386 240.244
R5774 gnd.n7308 gnd.n386 240.244
R5775 gnd.n7311 gnd.n7308 240.244
R5776 gnd.n7311 gnd.n369 240.244
R5777 gnd.n7331 gnd.n369 240.244
R5778 gnd.n7334 gnd.n7331 240.244
R5779 gnd.n7334 gnd.n104 240.244
R5780 gnd.n7753 gnd.n104 240.244
R5781 gnd.n7753 gnd.n105 240.244
R5782 gnd.n115 gnd.n105 240.244
R5783 gnd.n7747 gnd.n115 240.244
R5784 gnd.n7747 gnd.n116 240.244
R5785 gnd.n7739 gnd.n116 240.244
R5786 gnd.n7739 gnd.n132 240.244
R5787 gnd.n7735 gnd.n132 240.244
R5788 gnd.n7735 gnd.n137 240.244
R5789 gnd.n7727 gnd.n137 240.244
R5790 gnd.n7727 gnd.n149 240.244
R5791 gnd.n7723 gnd.n149 240.244
R5792 gnd.n7723 gnd.n155 240.244
R5793 gnd.n7715 gnd.n155 240.244
R5794 gnd.n7715 gnd.n169 240.244
R5795 gnd.n7711 gnd.n169 240.244
R5796 gnd.n7711 gnd.n175 240.244
R5797 gnd.n7703 gnd.n175 240.244
R5798 gnd.n7703 gnd.n187 240.244
R5799 gnd.n7699 gnd.n187 240.244
R5800 gnd.n7699 gnd.n193 240.244
R5801 gnd.n7691 gnd.n193 240.244
R5802 gnd.n7691 gnd.n207 240.244
R5803 gnd.n7687 gnd.n207 240.244
R5804 gnd.n7687 gnd.n213 240.244
R5805 gnd.n7679 gnd.n213 240.244
R5806 gnd.n7679 gnd.n226 240.244
R5807 gnd.n7675 gnd.n226 240.244
R5808 gnd.n7675 gnd.n232 240.244
R5809 gnd.n7667 gnd.n232 240.244
R5810 gnd.n7667 gnd.n245 240.244
R5811 gnd.n5959 gnd.n5958 240.244
R5812 gnd.n5956 gnd.n5872 240.244
R5813 gnd.n5952 gnd.n5951 240.244
R5814 gnd.n5949 gnd.n5878 240.244
R5815 gnd.n5945 gnd.n5944 240.244
R5816 gnd.n5942 gnd.n5885 240.244
R5817 gnd.n5938 gnd.n5937 240.244
R5818 gnd.n5935 gnd.n5892 240.244
R5819 gnd.n5931 gnd.n5930 240.244
R5820 gnd.n5928 gnd.n5899 240.244
R5821 gnd.n5924 gnd.n5923 240.244
R5822 gnd.n5921 gnd.n5909 240.244
R5823 gnd.n5917 gnd.n5916 240.244
R5824 gnd.n6026 gnd.n1367 240.244
R5825 gnd.n6024 gnd.n6023 240.244
R5826 gnd.n6021 gnd.n1371 240.244
R5827 gnd.n6017 gnd.n6016 240.244
R5828 gnd.n6014 gnd.n1378 240.244
R5829 gnd.n6007 gnd.n1387 240.244
R5830 gnd.n6005 gnd.n6004 240.244
R5831 gnd.n6002 gnd.n1389 240.244
R5832 gnd.n5998 gnd.n5997 240.244
R5833 gnd.n5995 gnd.n1396 240.244
R5834 gnd.n5991 gnd.n5990 240.244
R5835 gnd.n5988 gnd.n1403 240.244
R5836 gnd.n5984 gnd.n5983 240.244
R5837 gnd.n5981 gnd.n1410 240.244
R5838 gnd.n5977 gnd.n5976 240.244
R5839 gnd.n4728 gnd.n1812 240.244
R5840 gnd.n5052 gnd.n1812 240.244
R5841 gnd.n5053 gnd.n5052 240.244
R5842 gnd.n5053 gnd.n1804 240.244
R5843 gnd.n1804 gnd.n1794 240.244
R5844 gnd.n5072 gnd.n1794 240.244
R5845 gnd.n5073 gnd.n5072 240.244
R5846 gnd.n5073 gnd.n1784 240.244
R5847 gnd.n5076 gnd.n1784 240.244
R5848 gnd.n5076 gnd.n1775 240.244
R5849 gnd.n1775 gnd.n1768 240.244
R5850 gnd.n5108 gnd.n1768 240.244
R5851 gnd.n5108 gnd.n1758 240.244
R5852 gnd.n5111 gnd.n1758 240.244
R5853 gnd.n5111 gnd.n1750 240.244
R5854 gnd.n1750 gnd.n1743 240.244
R5855 gnd.n5143 gnd.n1743 240.244
R5856 gnd.n5143 gnd.n1734 240.244
R5857 gnd.n5146 gnd.n1734 240.244
R5858 gnd.n5146 gnd.n1726 240.244
R5859 gnd.n1726 gnd.n1718 240.244
R5860 gnd.n5178 gnd.n1718 240.244
R5861 gnd.n5178 gnd.n1707 240.244
R5862 gnd.n5181 gnd.n1707 240.244
R5863 gnd.n5181 gnd.n1699 240.244
R5864 gnd.n5186 gnd.n1699 240.244
R5865 gnd.n5186 gnd.n1692 240.244
R5866 gnd.n1692 gnd.n1684 240.244
R5867 gnd.n5223 gnd.n1684 240.244
R5868 gnd.n5223 gnd.n1667 240.244
R5869 gnd.n5243 gnd.n1667 240.244
R5870 gnd.n5243 gnd.n1661 240.244
R5871 gnd.n5251 gnd.n1661 240.244
R5872 gnd.n5251 gnd.n1653 240.244
R5873 gnd.n1653 gnd.n1645 240.244
R5874 gnd.n5273 gnd.n1645 240.244
R5875 gnd.n5273 gnd.n1635 240.244
R5876 gnd.n5277 gnd.n1635 240.244
R5877 gnd.n5277 gnd.n1619 240.244
R5878 gnd.n1619 gnd.n1610 240.244
R5879 gnd.n5309 gnd.n1610 240.244
R5880 gnd.n5309 gnd.n1600 240.244
R5881 gnd.n5313 gnd.n1600 240.244
R5882 gnd.n5313 gnd.n1590 240.244
R5883 gnd.n1590 gnd.n1581 240.244
R5884 gnd.n5345 gnd.n1581 240.244
R5885 gnd.n5345 gnd.n1569 240.244
R5886 gnd.n5349 gnd.n1569 240.244
R5887 gnd.n5349 gnd.n1559 240.244
R5888 gnd.n5358 gnd.n1559 240.244
R5889 gnd.n5358 gnd.n1551 240.244
R5890 gnd.n1551 gnd.n1533 240.244
R5891 gnd.n5354 gnd.n1533 240.244
R5892 gnd.n5354 gnd.n1524 240.244
R5893 gnd.n1524 gnd.n1515 240.244
R5894 gnd.n5433 gnd.n1515 240.244
R5895 gnd.n5433 gnd.n1506 240.244
R5896 gnd.n5436 gnd.n1506 240.244
R5897 gnd.n5436 gnd.n1445 240.244
R5898 gnd.n5855 gnd.n1445 240.244
R5899 gnd.n5855 gnd.n1437 240.244
R5900 gnd.n1437 gnd.n1425 240.244
R5901 gnd.n5967 gnd.n1425 240.244
R5902 gnd.n5967 gnd.n1419 240.244
R5903 gnd.n4886 gnd.n4882 240.244
R5904 gnd.n4892 gnd.n4882 240.244
R5905 gnd.n4896 gnd.n4894 240.244
R5906 gnd.n4902 gnd.n4878 240.244
R5907 gnd.n4906 gnd.n4904 240.244
R5908 gnd.n4912 gnd.n4874 240.244
R5909 gnd.n4916 gnd.n4914 240.244
R5910 gnd.n4922 gnd.n4870 240.244
R5911 gnd.n4926 gnd.n4924 240.244
R5912 gnd.n4932 gnd.n4863 240.244
R5913 gnd.n4936 gnd.n4934 240.244
R5914 gnd.n4942 gnd.n4859 240.244
R5915 gnd.n4946 gnd.n4944 240.244
R5916 gnd.n4952 gnd.n4855 240.244
R5917 gnd.n4956 gnd.n4954 240.244
R5918 gnd.n4962 gnd.n4851 240.244
R5919 gnd.n4966 gnd.n4964 240.244
R5920 gnd.n4972 gnd.n4847 240.244
R5921 gnd.n4976 gnd.n4974 240.244
R5922 gnd.n4984 gnd.n4843 240.244
R5923 gnd.n4988 gnd.n4986 240.244
R5924 gnd.n4994 gnd.n4839 240.244
R5925 gnd.n4998 gnd.n4996 240.244
R5926 gnd.n5004 gnd.n4835 240.244
R5927 gnd.n5008 gnd.n5006 240.244
R5928 gnd.n5014 gnd.n4831 240.244
R5929 gnd.n5018 gnd.n5016 240.244
R5930 gnd.n5025 gnd.n4827 240.244
R5931 gnd.n5028 gnd.n5027 240.244
R5932 gnd.n5044 gnd.n1815 240.244
R5933 gnd.n5050 gnd.n1815 240.244
R5934 gnd.n5050 gnd.n1802 240.244
R5935 gnd.n5064 gnd.n1802 240.244
R5936 gnd.n5064 gnd.n1798 240.244
R5937 gnd.n5070 gnd.n1798 240.244
R5938 gnd.n5070 gnd.n1782 240.244
R5939 gnd.n5088 gnd.n1782 240.244
R5940 gnd.n5088 gnd.n1777 240.244
R5941 gnd.n5096 gnd.n1777 240.244
R5942 gnd.n5096 gnd.n1778 240.244
R5943 gnd.n1778 gnd.n1757 240.244
R5944 gnd.n5123 gnd.n1757 240.244
R5945 gnd.n5123 gnd.n1752 240.244
R5946 gnd.n5131 gnd.n1752 240.244
R5947 gnd.n5131 gnd.n1753 240.244
R5948 gnd.n1753 gnd.n1733 240.244
R5949 gnd.n5158 gnd.n1733 240.244
R5950 gnd.n5158 gnd.n1728 240.244
R5951 gnd.n5166 gnd.n1728 240.244
R5952 gnd.n5166 gnd.n1729 240.244
R5953 gnd.n1729 gnd.n1706 240.244
R5954 gnd.n5195 gnd.n1706 240.244
R5955 gnd.n5195 gnd.n1701 240.244
R5956 gnd.n5203 gnd.n1701 240.244
R5957 gnd.n5203 gnd.n1702 240.244
R5958 gnd.n1702 gnd.n1686 240.244
R5959 gnd.n5218 gnd.n1686 240.244
R5960 gnd.n5221 gnd.n5218 240.244
R5961 gnd.n5221 gnd.n1672 240.244
R5962 gnd.n5241 gnd.n1672 240.244
R5963 gnd.n5241 gnd.n5238 240.244
R5964 gnd.n5238 gnd.n1656 240.244
R5965 gnd.n5262 gnd.n1656 240.244
R5966 gnd.n5262 gnd.n5259 240.244
R5967 gnd.n5259 gnd.n1633 240.244
R5968 gnd.n5290 gnd.n1633 240.244
R5969 gnd.n5290 gnd.n1622 240.244
R5970 gnd.n5298 gnd.n1622 240.244
R5971 gnd.n5298 gnd.n1623 240.244
R5972 gnd.n1623 gnd.n1598 240.244
R5973 gnd.n5326 gnd.n1598 240.244
R5974 gnd.n5326 gnd.n1593 240.244
R5975 gnd.n5334 gnd.n1593 240.244
R5976 gnd.n5334 gnd.n1594 240.244
R5977 gnd.n1594 gnd.n1567 240.244
R5978 gnd.n5368 gnd.n1567 240.244
R5979 gnd.n5368 gnd.n1562 240.244
R5980 gnd.n5376 gnd.n1562 240.244
R5981 gnd.n5376 gnd.n1563 240.244
R5982 gnd.n1563 gnd.n1531 240.244
R5983 gnd.n5411 gnd.n1531 240.244
R5984 gnd.n5411 gnd.n1526 240.244
R5985 gnd.n5419 gnd.n1526 240.244
R5986 gnd.n5419 gnd.n1527 240.244
R5987 gnd.n1527 gnd.n1504 240.244
R5988 gnd.n5445 gnd.n1504 240.244
R5989 gnd.n5445 gnd.n1500 240.244
R5990 gnd.n5451 gnd.n1500 240.244
R5991 gnd.n5451 gnd.n1435 240.244
R5992 gnd.n5865 gnd.n1435 240.244
R5993 gnd.n5865 gnd.n1430 240.244
R5994 gnd.n5965 gnd.n1430 240.244
R5995 gnd.n5965 gnd.n1431 240.244
R5996 gnd.n4725 gnd.n1843 240.244
R5997 gnd.n4718 gnd.n4717 240.244
R5998 gnd.n4715 gnd.n4714 240.244
R5999 gnd.n4711 gnd.n4710 240.244
R6000 gnd.n4707 gnd.n4706 240.244
R6001 gnd.n4703 gnd.n4702 240.244
R6002 gnd.n4699 gnd.n4698 240.244
R6003 gnd.n4695 gnd.n4694 240.244
R6004 gnd.n3968 gnd.n3680 240.244
R6005 gnd.n3978 gnd.n3680 240.244
R6006 gnd.n3978 gnd.n3671 240.244
R6007 gnd.n3671 gnd.n3660 240.244
R6008 gnd.n3999 gnd.n3660 240.244
R6009 gnd.n3999 gnd.n3654 240.244
R6010 gnd.n4009 gnd.n3654 240.244
R6011 gnd.n4009 gnd.n3643 240.244
R6012 gnd.n3643 gnd.n3635 240.244
R6013 gnd.n4027 gnd.n3635 240.244
R6014 gnd.n4028 gnd.n4027 240.244
R6015 gnd.n4028 gnd.n3620 240.244
R6016 gnd.n4030 gnd.n3620 240.244
R6017 gnd.n4030 gnd.n3606 240.244
R6018 gnd.n4072 gnd.n3606 240.244
R6019 gnd.n4073 gnd.n4072 240.244
R6020 gnd.n4076 gnd.n4073 240.244
R6021 gnd.n4076 gnd.n3561 240.244
R6022 gnd.n3601 gnd.n3561 240.244
R6023 gnd.n3601 gnd.n3571 240.244
R6024 gnd.n4086 gnd.n3571 240.244
R6025 gnd.n4086 gnd.n3592 240.244
R6026 gnd.n4096 gnd.n3592 240.244
R6027 gnd.n4096 gnd.n3458 240.244
R6028 gnd.n4141 gnd.n3458 240.244
R6029 gnd.n4141 gnd.n3444 240.244
R6030 gnd.n4163 gnd.n3444 240.244
R6031 gnd.n4164 gnd.n4163 240.244
R6032 gnd.n4164 gnd.n3431 240.244
R6033 gnd.n3431 gnd.n3420 240.244
R6034 gnd.n4195 gnd.n3420 240.244
R6035 gnd.n4196 gnd.n4195 240.244
R6036 gnd.n4197 gnd.n4196 240.244
R6037 gnd.n4197 gnd.n3405 240.244
R6038 gnd.n3405 gnd.n3404 240.244
R6039 gnd.n3404 gnd.n3389 240.244
R6040 gnd.n4248 gnd.n3389 240.244
R6041 gnd.n4249 gnd.n4248 240.244
R6042 gnd.n4249 gnd.n3376 240.244
R6043 gnd.n3376 gnd.n3365 240.244
R6044 gnd.n4280 gnd.n3365 240.244
R6045 gnd.n4281 gnd.n4280 240.244
R6046 gnd.n4282 gnd.n4281 240.244
R6047 gnd.n4282 gnd.n3349 240.244
R6048 gnd.n3349 gnd.n3348 240.244
R6049 gnd.n3348 gnd.n3335 240.244
R6050 gnd.n4337 gnd.n3335 240.244
R6051 gnd.n4338 gnd.n4337 240.244
R6052 gnd.n4338 gnd.n1909 240.244
R6053 gnd.n1909 gnd.n1899 240.244
R6054 gnd.n4626 gnd.n1899 240.244
R6055 gnd.n4629 gnd.n4626 240.244
R6056 gnd.n4629 gnd.n4628 240.244
R6057 gnd.n3958 gnd.n3693 240.244
R6058 gnd.n3714 gnd.n3693 240.244
R6059 gnd.n3717 gnd.n3716 240.244
R6060 gnd.n3724 gnd.n3723 240.244
R6061 gnd.n3727 gnd.n3726 240.244
R6062 gnd.n3734 gnd.n3733 240.244
R6063 gnd.n3737 gnd.n3736 240.244
R6064 gnd.n3744 gnd.n3743 240.244
R6065 gnd.n3966 gnd.n3690 240.244
R6066 gnd.n3690 gnd.n3669 240.244
R6067 gnd.n3989 gnd.n3669 240.244
R6068 gnd.n3989 gnd.n3663 240.244
R6069 gnd.n3997 gnd.n3663 240.244
R6070 gnd.n3997 gnd.n3665 240.244
R6071 gnd.n3665 gnd.n3641 240.244
R6072 gnd.n4019 gnd.n3641 240.244
R6073 gnd.n4019 gnd.n3637 240.244
R6074 gnd.n4025 gnd.n3637 240.244
R6075 gnd.n4025 gnd.n3619 240.244
R6076 gnd.n4050 gnd.n3619 240.244
R6077 gnd.n4050 gnd.n3614 240.244
R6078 gnd.n4062 gnd.n3614 240.244
R6079 gnd.n4062 gnd.n3615 240.244
R6080 gnd.n4058 gnd.n3615 240.244
R6081 gnd.n4058 gnd.n3563 240.244
R6082 gnd.n4110 gnd.n3563 240.244
R6083 gnd.n4110 gnd.n3564 240.244
R6084 gnd.n4106 gnd.n3564 240.244
R6085 gnd.n4106 gnd.n3570 240.244
R6086 gnd.n3590 gnd.n3570 240.244
R6087 gnd.n3590 gnd.n3456 240.244
R6088 gnd.n4145 gnd.n3456 240.244
R6089 gnd.n4145 gnd.n3451 240.244
R6090 gnd.n4153 gnd.n3451 240.244
R6091 gnd.n4153 gnd.n3452 240.244
R6092 gnd.n3452 gnd.n3429 240.244
R6093 gnd.n4185 gnd.n3429 240.244
R6094 gnd.n4185 gnd.n3424 240.244
R6095 gnd.n4193 gnd.n3424 240.244
R6096 gnd.n4193 gnd.n3425 240.244
R6097 gnd.n3425 gnd.n3402 240.244
R6098 gnd.n4230 gnd.n3402 240.244
R6099 gnd.n4230 gnd.n3397 240.244
R6100 gnd.n4238 gnd.n3397 240.244
R6101 gnd.n4238 gnd.n3398 240.244
R6102 gnd.n3398 gnd.n3374 240.244
R6103 gnd.n4270 gnd.n3374 240.244
R6104 gnd.n4270 gnd.n3369 240.244
R6105 gnd.n4278 gnd.n3369 240.244
R6106 gnd.n4278 gnd.n3370 240.244
R6107 gnd.n3370 gnd.n3347 240.244
R6108 gnd.n4319 gnd.n3347 240.244
R6109 gnd.n4319 gnd.n3342 240.244
R6110 gnd.n4327 gnd.n3342 240.244
R6111 gnd.n4327 gnd.n3343 240.244
R6112 gnd.n3343 gnd.n1907 240.244
R6113 gnd.n4614 gnd.n1907 240.244
R6114 gnd.n4614 gnd.n1902 240.244
R6115 gnd.n4624 gnd.n1902 240.244
R6116 gnd.n4624 gnd.n1903 240.244
R6117 gnd.n1903 gnd.n1842 240.244
R6118 gnd.n7403 gnd.n251 240.244
R6119 gnd.n7409 gnd.n7408 240.244
R6120 gnd.n7412 gnd.n7411 240.244
R6121 gnd.n7419 gnd.n7418 240.244
R6122 gnd.n7422 gnd.n7421 240.244
R6123 gnd.n7429 gnd.n7428 240.244
R6124 gnd.n7432 gnd.n7431 240.244
R6125 gnd.n7439 gnd.n7438 240.244
R6126 gnd.n7442 gnd.n7441 240.244
R6127 gnd.n571 gnd.n560 240.244
R6128 gnd.n7079 gnd.n560 240.244
R6129 gnd.n7079 gnd.n555 240.244
R6130 gnd.n7086 gnd.n555 240.244
R6131 gnd.n7086 gnd.n533 240.244
R6132 gnd.n533 gnd.n520 240.244
R6133 gnd.n7129 gnd.n520 240.244
R6134 gnd.n7129 gnd.n521 240.244
R6135 gnd.n521 gnd.n517 240.244
R6136 gnd.n517 gnd.n498 240.244
R6137 gnd.n7136 gnd.n498 240.244
R6138 gnd.n7136 gnd.n489 240.244
R6139 gnd.n7143 gnd.n489 240.244
R6140 gnd.n7143 gnd.n468 240.244
R6141 gnd.n468 gnd.n455 240.244
R6142 gnd.n7199 gnd.n455 240.244
R6143 gnd.n7199 gnd.n450 240.244
R6144 gnd.n7215 gnd.n450 240.244
R6145 gnd.n7215 gnd.n441 240.244
R6146 gnd.n7204 gnd.n441 240.244
R6147 gnd.n7204 gnd.n432 240.244
R6148 gnd.n432 gnd.n424 240.244
R6149 gnd.n424 gnd.n413 240.244
R6150 gnd.n413 gnd.n401 240.244
R6151 gnd.n7286 gnd.n401 240.244
R6152 gnd.n7286 gnd.n396 240.244
R6153 gnd.n7298 gnd.n396 240.244
R6154 gnd.n7298 gnd.n389 240.244
R6155 gnd.n389 gnd.n384 240.244
R6156 gnd.n384 gnd.n379 240.244
R6157 gnd.n379 gnd.n372 240.244
R6158 gnd.n372 gnd.n368 240.244
R6159 gnd.n368 gnd.n98 240.244
R6160 gnd.n7755 gnd.n98 240.244
R6161 gnd.n7755 gnd.n100 240.244
R6162 gnd.n7361 gnd.n100 240.244
R6163 gnd.n7361 gnd.n119 240.244
R6164 gnd.n7489 gnd.n119 240.244
R6165 gnd.n7489 gnd.n130 240.244
R6166 gnd.n7485 gnd.n130 240.244
R6167 gnd.n7485 gnd.n139 240.244
R6168 gnd.n7482 gnd.n139 240.244
R6169 gnd.n7482 gnd.n148 240.244
R6170 gnd.n7479 gnd.n148 240.244
R6171 gnd.n7479 gnd.n158 240.244
R6172 gnd.n7476 gnd.n158 240.244
R6173 gnd.n7476 gnd.n167 240.244
R6174 gnd.n7473 gnd.n167 240.244
R6175 gnd.n7473 gnd.n177 240.244
R6176 gnd.n7470 gnd.n177 240.244
R6177 gnd.n7470 gnd.n186 240.244
R6178 gnd.n7467 gnd.n186 240.244
R6179 gnd.n7467 gnd.n196 240.244
R6180 gnd.n7464 gnd.n196 240.244
R6181 gnd.n7464 gnd.n205 240.244
R6182 gnd.n7461 gnd.n205 240.244
R6183 gnd.n7461 gnd.n215 240.244
R6184 gnd.n7458 gnd.n215 240.244
R6185 gnd.n7458 gnd.n224 240.244
R6186 gnd.n7455 gnd.n224 240.244
R6187 gnd.n7455 gnd.n234 240.244
R6188 gnd.n7452 gnd.n234 240.244
R6189 gnd.n7452 gnd.n243 240.244
R6190 gnd.n7449 gnd.n243 240.244
R6191 gnd.n706 gnd.n705 240.244
R6192 gnd.n714 gnd.n713 240.244
R6193 gnd.n716 gnd.n715 240.244
R6194 gnd.n724 gnd.n723 240.244
R6195 gnd.n732 gnd.n731 240.244
R6196 gnd.n734 gnd.n733 240.244
R6197 gnd.n742 gnd.n741 240.244
R6198 gnd.n752 gnd.n751 240.244
R6199 gnd.n6874 gnd.n627 240.244
R6200 gnd.n7067 gnd.n574 240.244
R6201 gnd.n574 gnd.n563 240.244
R6202 gnd.n578 gnd.n563 240.244
R6203 gnd.n578 gnd.n535 240.244
R6204 gnd.n7117 gnd.n535 240.244
R6205 gnd.n7117 gnd.n536 240.244
R6206 gnd.n536 gnd.n524 240.244
R6207 gnd.n7112 gnd.n524 240.244
R6208 gnd.n7112 gnd.n500 240.244
R6209 gnd.n7152 gnd.n500 240.244
R6210 gnd.n7152 gnd.n501 240.244
R6211 gnd.n501 gnd.n491 240.244
R6212 gnd.n491 gnd.n470 240.244
R6213 gnd.n7187 gnd.n470 240.244
R6214 gnd.n7187 gnd.n471 240.244
R6215 gnd.n471 gnd.n459 240.244
R6216 gnd.n7182 gnd.n459 240.244
R6217 gnd.n7182 gnd.n443 240.244
R6218 gnd.n7227 gnd.n443 240.244
R6219 gnd.n7227 gnd.n444 240.244
R6220 gnd.n444 gnd.n433 240.244
R6221 gnd.n433 gnd.n415 240.244
R6222 gnd.n7274 gnd.n415 240.244
R6223 gnd.n7274 gnd.n416 240.244
R6224 gnd.n416 gnd.n405 240.244
R6225 gnd.n7269 gnd.n405 240.244
R6226 gnd.n7269 gnd.n390 240.244
R6227 gnd.n7306 gnd.n390 240.244
R6228 gnd.n7306 gnd.n385 240.244
R6229 gnd.n385 gnd.n373 240.244
R6230 gnd.n7329 gnd.n373 240.244
R6231 gnd.n7329 gnd.n362 240.244
R6232 gnd.n7342 gnd.n362 240.244
R6233 gnd.n7342 gnd.n103 240.244
R6234 gnd.n7354 gnd.n103 240.244
R6235 gnd.n7354 gnd.n121 240.244
R6236 gnd.n7745 gnd.n121 240.244
R6237 gnd.n7745 gnd.n122 240.244
R6238 gnd.n7741 gnd.n122 240.244
R6239 gnd.n7741 gnd.n128 240.244
R6240 gnd.n7733 gnd.n128 240.244
R6241 gnd.n7733 gnd.n140 240.244
R6242 gnd.n7729 gnd.n140 240.244
R6243 gnd.n7729 gnd.n145 240.244
R6244 gnd.n7721 gnd.n145 240.244
R6245 gnd.n7721 gnd.n160 240.244
R6246 gnd.n7717 gnd.n160 240.244
R6247 gnd.n7717 gnd.n165 240.244
R6248 gnd.n7709 gnd.n165 240.244
R6249 gnd.n7709 gnd.n178 240.244
R6250 gnd.n7705 gnd.n178 240.244
R6251 gnd.n7705 gnd.n183 240.244
R6252 gnd.n7697 gnd.n183 240.244
R6253 gnd.n7697 gnd.n198 240.244
R6254 gnd.n7693 gnd.n198 240.244
R6255 gnd.n7693 gnd.n203 240.244
R6256 gnd.n7685 gnd.n203 240.244
R6257 gnd.n7685 gnd.n216 240.244
R6258 gnd.n7681 gnd.n216 240.244
R6259 gnd.n7681 gnd.n221 240.244
R6260 gnd.n7673 gnd.n221 240.244
R6261 gnd.n7673 gnd.n236 240.244
R6262 gnd.n7669 gnd.n236 240.244
R6263 gnd.n7669 gnd.n241 240.244
R6264 gnd.n1862 gnd.n1820 240.244
R6265 gnd.n4685 gnd.n4684 240.244
R6266 gnd.n4681 gnd.n4680 240.244
R6267 gnd.n4677 gnd.n4676 240.244
R6268 gnd.n4673 gnd.n4672 240.244
R6269 gnd.n4669 gnd.n4668 240.244
R6270 gnd.n4665 gnd.n4664 240.244
R6271 gnd.n4661 gnd.n4660 240.244
R6272 gnd.n4657 gnd.n4656 240.244
R6273 gnd.n4653 gnd.n4652 240.244
R6274 gnd.n4649 gnd.n4648 240.244
R6275 gnd.n4645 gnd.n4644 240.244
R6276 gnd.n4641 gnd.n4640 240.244
R6277 gnd.n3881 gnd.n3778 240.244
R6278 gnd.n3881 gnd.n3771 240.244
R6279 gnd.n3892 gnd.n3771 240.244
R6280 gnd.n3892 gnd.n3767 240.244
R6281 gnd.n3898 gnd.n3767 240.244
R6282 gnd.n3898 gnd.n3759 240.244
R6283 gnd.n3908 gnd.n3759 240.244
R6284 gnd.n3908 gnd.n3754 240.244
R6285 gnd.n3944 gnd.n3754 240.244
R6286 gnd.n3944 gnd.n3755 240.244
R6287 gnd.n3755 gnd.n3702 240.244
R6288 gnd.n3939 gnd.n3702 240.244
R6289 gnd.n3939 gnd.n3938 240.244
R6290 gnd.n3938 gnd.n3681 240.244
R6291 gnd.n3934 gnd.n3681 240.244
R6292 gnd.n3934 gnd.n3672 240.244
R6293 gnd.n3931 gnd.n3672 240.244
R6294 gnd.n3931 gnd.n3930 240.244
R6295 gnd.n3930 gnd.n3655 240.244
R6296 gnd.n3926 gnd.n3655 240.244
R6297 gnd.n3926 gnd.n3644 240.244
R6298 gnd.n3644 gnd.n3625 240.244
R6299 gnd.n4039 gnd.n3625 240.244
R6300 gnd.n4039 gnd.n3621 240.244
R6301 gnd.n4047 gnd.n3621 240.244
R6302 gnd.n4047 gnd.n3612 240.244
R6303 gnd.n3612 gnd.n3548 240.244
R6304 gnd.n4119 gnd.n3548 240.244
R6305 gnd.n4119 gnd.n3549 240.244
R6306 gnd.n3560 gnd.n3549 240.244
R6307 gnd.n3595 gnd.n3560 240.244
R6308 gnd.n3598 gnd.n3595 240.244
R6309 gnd.n3598 gnd.n3572 240.244
R6310 gnd.n3585 gnd.n3572 240.244
R6311 gnd.n3585 gnd.n3582 240.244
R6312 gnd.n3582 gnd.n3459 240.244
R6313 gnd.n4140 gnd.n3459 240.244
R6314 gnd.n4140 gnd.n3449 240.244
R6315 gnd.n4136 gnd.n3449 240.244
R6316 gnd.n4136 gnd.n3443 240.244
R6317 gnd.n4133 gnd.n3443 240.244
R6318 gnd.n4133 gnd.n3432 240.244
R6319 gnd.n4130 gnd.n3432 240.244
R6320 gnd.n4130 gnd.n3410 240.244
R6321 gnd.n4206 gnd.n3410 240.244
R6322 gnd.n4206 gnd.n3406 240.244
R6323 gnd.n4227 gnd.n3406 240.244
R6324 gnd.n4227 gnd.n3395 240.244
R6325 gnd.n4223 gnd.n3395 240.244
R6326 gnd.n4223 gnd.n3388 240.244
R6327 gnd.n4220 gnd.n3388 240.244
R6328 gnd.n4220 gnd.n3377 240.244
R6329 gnd.n4217 gnd.n3377 240.244
R6330 gnd.n4217 gnd.n3354 240.244
R6331 gnd.n4291 gnd.n3354 240.244
R6332 gnd.n4291 gnd.n3350 240.244
R6333 gnd.n4316 gnd.n3350 240.244
R6334 gnd.n4316 gnd.n3341 240.244
R6335 gnd.n4312 gnd.n3341 240.244
R6336 gnd.n4312 gnd.n3334 240.244
R6337 gnd.n4308 gnd.n3334 240.244
R6338 gnd.n4308 gnd.n3323 240.244
R6339 gnd.n4305 gnd.n3323 240.244
R6340 gnd.n4305 gnd.n1891 240.244
R6341 gnd.n4636 gnd.n1891 240.244
R6342 gnd.n3795 gnd.n3794 240.244
R6343 gnd.n3866 gnd.n3794 240.244
R6344 gnd.n3864 gnd.n3863 240.244
R6345 gnd.n3860 gnd.n3859 240.244
R6346 gnd.n3856 gnd.n3855 240.244
R6347 gnd.n3852 gnd.n3851 240.244
R6348 gnd.n3848 gnd.n3847 240.244
R6349 gnd.n3844 gnd.n3843 240.244
R6350 gnd.n3840 gnd.n3839 240.244
R6351 gnd.n3836 gnd.n3835 240.244
R6352 gnd.n3832 gnd.n3831 240.244
R6353 gnd.n3828 gnd.n3827 240.244
R6354 gnd.n3824 gnd.n3782 240.244
R6355 gnd.n3884 gnd.n3776 240.244
R6356 gnd.n3884 gnd.n3772 240.244
R6357 gnd.n3890 gnd.n3772 240.244
R6358 gnd.n3890 gnd.n3765 240.244
R6359 gnd.n3900 gnd.n3765 240.244
R6360 gnd.n3900 gnd.n3761 240.244
R6361 gnd.n3906 gnd.n3761 240.244
R6362 gnd.n3906 gnd.n3752 240.244
R6363 gnd.n3946 gnd.n3752 240.244
R6364 gnd.n3946 gnd.n3703 240.244
R6365 gnd.n3954 gnd.n3703 240.244
R6366 gnd.n3954 gnd.n3704 240.244
R6367 gnd.n3704 gnd.n3682 240.244
R6368 gnd.n3975 gnd.n3682 240.244
R6369 gnd.n3975 gnd.n3674 240.244
R6370 gnd.n3986 gnd.n3674 240.244
R6371 gnd.n3986 gnd.n3675 240.244
R6372 gnd.n3675 gnd.n3656 240.244
R6373 gnd.n4006 gnd.n3656 240.244
R6374 gnd.n4006 gnd.n3646 240.244
R6375 gnd.n4016 gnd.n3646 240.244
R6376 gnd.n4016 gnd.n3627 240.244
R6377 gnd.n4037 gnd.n3627 240.244
R6378 gnd.n4037 gnd.n3629 240.244
R6379 gnd.n3629 gnd.n3610 240.244
R6380 gnd.n4065 gnd.n3610 240.244
R6381 gnd.n4065 gnd.n3552 240.244
R6382 gnd.n4117 gnd.n3552 240.244
R6383 gnd.n4117 gnd.n3553 240.244
R6384 gnd.n4113 gnd.n3553 240.244
R6385 gnd.n4113 gnd.n3559 240.244
R6386 gnd.n3574 gnd.n3559 240.244
R6387 gnd.n4103 gnd.n3574 240.244
R6388 gnd.n4103 gnd.n3575 240.244
R6389 gnd.n4099 gnd.n3575 240.244
R6390 gnd.n4099 gnd.n3581 240.244
R6391 gnd.n3581 gnd.n3448 240.244
R6392 gnd.n4156 gnd.n3448 240.244
R6393 gnd.n4156 gnd.n3441 240.244
R6394 gnd.n4167 gnd.n3441 240.244
R6395 gnd.n4167 gnd.n3434 240.244
R6396 gnd.n4182 gnd.n3434 240.244
R6397 gnd.n4182 gnd.n3435 240.244
R6398 gnd.n3435 gnd.n3413 240.244
R6399 gnd.n4204 gnd.n3413 240.244
R6400 gnd.n4204 gnd.n3414 240.244
R6401 gnd.n3414 gnd.n3393 240.244
R6402 gnd.n4241 gnd.n3393 240.244
R6403 gnd.n4241 gnd.n3386 240.244
R6404 gnd.n4252 gnd.n3386 240.244
R6405 gnd.n4252 gnd.n3379 240.244
R6406 gnd.n4267 gnd.n3379 240.244
R6407 gnd.n4267 gnd.n3380 240.244
R6408 gnd.n3380 gnd.n3357 240.244
R6409 gnd.n4289 gnd.n3357 240.244
R6410 gnd.n4289 gnd.n3359 240.244
R6411 gnd.n3359 gnd.n3339 240.244
R6412 gnd.n4330 gnd.n3339 240.244
R6413 gnd.n4330 gnd.n3332 240.244
R6414 gnd.n4341 gnd.n3332 240.244
R6415 gnd.n4341 gnd.n3325 240.244
R6416 gnd.n4610 gnd.n3325 240.244
R6417 gnd.n4610 gnd.n3326 240.244
R6418 gnd.n3326 gnd.n1894 240.244
R6419 gnd.n4634 gnd.n1894 240.244
R6420 gnd.n5701 gnd.n5700 240.244
R6421 gnd.n5713 gnd.n5712 240.244
R6422 gnd.n5724 gnd.n5715 240.244
R6423 gnd.n5727 gnd.n5726 240.244
R6424 gnd.n5736 gnd.n5735 240.244
R6425 gnd.n5747 gnd.n5738 240.244
R6426 gnd.n5750 gnd.n5749 240.244
R6427 gnd.n5759 gnd.n5758 240.244
R6428 gnd.n5764 gnd.n5761 240.244
R6429 gnd.n4777 gnd.n4729 240.244
R6430 gnd.n4777 gnd.n1813 240.244
R6431 gnd.n4774 gnd.n1813 240.244
R6432 gnd.n4774 gnd.n1805 240.244
R6433 gnd.n4771 gnd.n1805 240.244
R6434 gnd.n4771 gnd.n1796 240.244
R6435 gnd.n4768 gnd.n1796 240.244
R6436 gnd.n4768 gnd.n1785 240.244
R6437 gnd.n1785 gnd.n1774 240.244
R6438 gnd.n5098 gnd.n1774 240.244
R6439 gnd.n5098 gnd.n1770 240.244
R6440 gnd.n5106 gnd.n1770 240.244
R6441 gnd.n5106 gnd.n1759 240.244
R6442 gnd.n1759 gnd.n1749 240.244
R6443 gnd.n5133 gnd.n1749 240.244
R6444 gnd.n5133 gnd.n1745 240.244
R6445 gnd.n5141 gnd.n1745 240.244
R6446 gnd.n5141 gnd.n1735 240.244
R6447 gnd.n1735 gnd.n1724 240.244
R6448 gnd.n5168 gnd.n1724 240.244
R6449 gnd.n5168 gnd.n1720 240.244
R6450 gnd.n5176 gnd.n1720 240.244
R6451 gnd.n5176 gnd.n1708 240.244
R6452 gnd.n1708 gnd.n1697 240.244
R6453 gnd.n5205 gnd.n1697 240.244
R6454 gnd.n5205 gnd.n1693 240.244
R6455 gnd.n5213 gnd.n1693 240.244
R6456 gnd.n5213 gnd.n1688 240.244
R6457 gnd.n1688 gnd.n1678 240.244
R6458 gnd.n5230 gnd.n1678 240.244
R6459 gnd.n5230 gnd.n1669 240.244
R6460 gnd.n5236 gnd.n1669 240.244
R6461 gnd.n5236 gnd.n1651 240.244
R6462 gnd.n5264 gnd.n1651 240.244
R6463 gnd.n5264 gnd.n1646 240.244
R6464 gnd.n5271 gnd.n1646 240.244
R6465 gnd.n5271 gnd.n1636 240.244
R6466 gnd.n1636 gnd.n1617 240.244
R6467 gnd.n5300 gnd.n1617 240.244
R6468 gnd.n5300 gnd.n1612 240.244
R6469 gnd.n5307 gnd.n1612 240.244
R6470 gnd.n5307 gnd.n1601 240.244
R6471 gnd.n1601 gnd.n1588 240.244
R6472 gnd.n5336 gnd.n1588 240.244
R6473 gnd.n5336 gnd.n1583 240.244
R6474 gnd.n5343 gnd.n1583 240.244
R6475 gnd.n5343 gnd.n1570 240.244
R6476 gnd.n1570 gnd.n1557 240.244
R6477 gnd.n5378 gnd.n1557 240.244
R6478 gnd.n5378 gnd.n1552 240.244
R6479 gnd.n5385 gnd.n1552 240.244
R6480 gnd.n5385 gnd.n1534 240.244
R6481 gnd.n1534 gnd.n1522 240.244
R6482 gnd.n5421 gnd.n1522 240.244
R6483 gnd.n5421 gnd.n1517 240.244
R6484 gnd.n5431 gnd.n1517 240.244
R6485 gnd.n5431 gnd.n1507 240.244
R6486 gnd.n5425 gnd.n1507 240.244
R6487 gnd.n5425 gnd.n1447 240.244
R6488 gnd.n5853 gnd.n1447 240.244
R6489 gnd.n5853 gnd.n1438 240.244
R6490 gnd.n1453 gnd.n1438 240.244
R6491 gnd.n1453 gnd.n1427 240.244
R6492 gnd.n1454 gnd.n1427 240.244
R6493 gnd.n4818 gnd.n4816 240.244
R6494 gnd.n4814 gnd.n4735 240.244
R6495 gnd.n4810 gnd.n4808 240.244
R6496 gnd.n4806 gnd.n4741 240.244
R6497 gnd.n4802 gnd.n4800 240.244
R6498 gnd.n4798 gnd.n4747 240.244
R6499 gnd.n4794 gnd.n4792 240.244
R6500 gnd.n4790 gnd.n4753 240.244
R6501 gnd.n4783 gnd.n4782 240.244
R6502 gnd.n5042 gnd.n4732 240.244
R6503 gnd.n4732 gnd.n1814 240.244
R6504 gnd.n1814 gnd.n1806 240.244
R6505 gnd.n5062 gnd.n1806 240.244
R6506 gnd.n5062 gnd.n1807 240.244
R6507 gnd.n1807 gnd.n1797 240.244
R6508 gnd.n1797 gnd.n1787 240.244
R6509 gnd.n5086 gnd.n1787 240.244
R6510 gnd.n5086 gnd.n1788 240.244
R6511 gnd.n1788 gnd.n1776 240.244
R6512 gnd.n5081 gnd.n1776 240.244
R6513 gnd.n5081 gnd.n1761 240.244
R6514 gnd.n5121 gnd.n1761 240.244
R6515 gnd.n5121 gnd.n1762 240.244
R6516 gnd.n1762 gnd.n1751 240.244
R6517 gnd.n5116 gnd.n1751 240.244
R6518 gnd.n5116 gnd.n1736 240.244
R6519 gnd.n5156 gnd.n1736 240.244
R6520 gnd.n5156 gnd.n1737 240.244
R6521 gnd.n1737 gnd.n1727 240.244
R6522 gnd.n5151 gnd.n1727 240.244
R6523 gnd.n5151 gnd.n1709 240.244
R6524 gnd.n5193 gnd.n1709 240.244
R6525 gnd.n5193 gnd.n1710 240.244
R6526 gnd.n1710 gnd.n1700 240.244
R6527 gnd.n1700 gnd.n1689 240.244
R6528 gnd.n5215 gnd.n1689 240.244
R6529 gnd.n5216 gnd.n5215 240.244
R6530 gnd.n5216 gnd.n1680 240.244
R6531 gnd.n5228 gnd.n1680 240.244
R6532 gnd.n5228 gnd.n1671 240.244
R6533 gnd.n1671 gnd.n1663 240.244
R6534 gnd.n5249 gnd.n1663 240.244
R6535 gnd.n5249 gnd.n1655 240.244
R6536 gnd.n5257 gnd.n1655 240.244
R6537 gnd.n5257 gnd.n1638 240.244
R6538 gnd.n5288 gnd.n1638 240.244
R6539 gnd.n5288 gnd.n1639 240.244
R6540 gnd.n1639 gnd.n1621 240.244
R6541 gnd.n5283 gnd.n1621 240.244
R6542 gnd.n5283 gnd.n1603 240.244
R6543 gnd.n5324 gnd.n1603 240.244
R6544 gnd.n5324 gnd.n1604 240.244
R6545 gnd.n1604 gnd.n1592 240.244
R6546 gnd.n5319 gnd.n1592 240.244
R6547 gnd.n5319 gnd.n1572 240.244
R6548 gnd.n5366 gnd.n1572 240.244
R6549 gnd.n5366 gnd.n1573 240.244
R6550 gnd.n1573 gnd.n1561 240.244
R6551 gnd.n5361 gnd.n1561 240.244
R6552 gnd.n5361 gnd.n1536 240.244
R6553 gnd.n5409 gnd.n1536 240.244
R6554 gnd.n5409 gnd.n1537 240.244
R6555 gnd.n1537 gnd.n1525 240.244
R6556 gnd.n5404 gnd.n1525 240.244
R6557 gnd.n5404 gnd.n1509 240.244
R6558 gnd.n5443 gnd.n1509 240.244
R6559 gnd.n5443 gnd.n1510 240.244
R6560 gnd.n1510 gnd.n1499 240.244
R6561 gnd.n1499 gnd.n1440 240.244
R6562 gnd.n5863 gnd.n1440 240.244
R6563 gnd.n5863 gnd.n1441 240.244
R6564 gnd.n1441 gnd.n1429 240.244
R6565 gnd.n5699 gnd.n1429 240.244
R6566 gnd.n3109 gnd.n2100 240.244
R6567 gnd.n3103 gnd.n2100 240.244
R6568 gnd.n3103 gnd.n2104 240.244
R6569 gnd.n3099 gnd.n2104 240.244
R6570 gnd.n3099 gnd.n2106 240.244
R6571 gnd.n3095 gnd.n2106 240.244
R6572 gnd.n3095 gnd.n2111 240.244
R6573 gnd.n3091 gnd.n2111 240.244
R6574 gnd.n3091 gnd.n2113 240.244
R6575 gnd.n3087 gnd.n2113 240.244
R6576 gnd.n3087 gnd.n2119 240.244
R6577 gnd.n3083 gnd.n2119 240.244
R6578 gnd.n3083 gnd.n2121 240.244
R6579 gnd.n3079 gnd.n2121 240.244
R6580 gnd.n3079 gnd.n2127 240.244
R6581 gnd.n3075 gnd.n2127 240.244
R6582 gnd.n3075 gnd.n2129 240.244
R6583 gnd.n3071 gnd.n2129 240.244
R6584 gnd.n3071 gnd.n2135 240.244
R6585 gnd.n3067 gnd.n2135 240.244
R6586 gnd.n3067 gnd.n2137 240.244
R6587 gnd.n3063 gnd.n2137 240.244
R6588 gnd.n3063 gnd.n2143 240.244
R6589 gnd.n3059 gnd.n2143 240.244
R6590 gnd.n3059 gnd.n2145 240.244
R6591 gnd.n3055 gnd.n2145 240.244
R6592 gnd.n3055 gnd.n2151 240.244
R6593 gnd.n3051 gnd.n2151 240.244
R6594 gnd.n3051 gnd.n2153 240.244
R6595 gnd.n3047 gnd.n2153 240.244
R6596 gnd.n3047 gnd.n2159 240.244
R6597 gnd.n3043 gnd.n2159 240.244
R6598 gnd.n3043 gnd.n2161 240.244
R6599 gnd.n3039 gnd.n2161 240.244
R6600 gnd.n3039 gnd.n2167 240.244
R6601 gnd.n3035 gnd.n2167 240.244
R6602 gnd.n3035 gnd.n2169 240.244
R6603 gnd.n3031 gnd.n2169 240.244
R6604 gnd.n3031 gnd.n2175 240.244
R6605 gnd.n3027 gnd.n2175 240.244
R6606 gnd.n3027 gnd.n2177 240.244
R6607 gnd.n3023 gnd.n2177 240.244
R6608 gnd.n3023 gnd.n2183 240.244
R6609 gnd.n3019 gnd.n2183 240.244
R6610 gnd.n3019 gnd.n2185 240.244
R6611 gnd.n3015 gnd.n2185 240.244
R6612 gnd.n3015 gnd.n2191 240.244
R6613 gnd.n3011 gnd.n2191 240.244
R6614 gnd.n3011 gnd.n2193 240.244
R6615 gnd.n3007 gnd.n2193 240.244
R6616 gnd.n3007 gnd.n2199 240.244
R6617 gnd.n3003 gnd.n2199 240.244
R6618 gnd.n3003 gnd.n2201 240.244
R6619 gnd.n2999 gnd.n2201 240.244
R6620 gnd.n2999 gnd.n2207 240.244
R6621 gnd.n2995 gnd.n2207 240.244
R6622 gnd.n2995 gnd.n2209 240.244
R6623 gnd.n2991 gnd.n2209 240.244
R6624 gnd.n2991 gnd.n2215 240.244
R6625 gnd.n2987 gnd.n2215 240.244
R6626 gnd.n2987 gnd.n2217 240.244
R6627 gnd.n2983 gnd.n2217 240.244
R6628 gnd.n2983 gnd.n2223 240.244
R6629 gnd.n2979 gnd.n2223 240.244
R6630 gnd.n2979 gnd.n2225 240.244
R6631 gnd.n2975 gnd.n2225 240.244
R6632 gnd.n2975 gnd.n2231 240.244
R6633 gnd.n2971 gnd.n2231 240.244
R6634 gnd.n2971 gnd.n2233 240.244
R6635 gnd.n2967 gnd.n2233 240.244
R6636 gnd.n2967 gnd.n2239 240.244
R6637 gnd.n2963 gnd.n2239 240.244
R6638 gnd.n2963 gnd.n2241 240.244
R6639 gnd.n2959 gnd.n2241 240.244
R6640 gnd.n2959 gnd.n2247 240.244
R6641 gnd.n2955 gnd.n2247 240.244
R6642 gnd.n2955 gnd.n2249 240.244
R6643 gnd.n2951 gnd.n2249 240.244
R6644 gnd.n2951 gnd.n2255 240.244
R6645 gnd.n2947 gnd.n2255 240.244
R6646 gnd.n2947 gnd.n2257 240.244
R6647 gnd.n2943 gnd.n2257 240.244
R6648 gnd.n2943 gnd.n2263 240.244
R6649 gnd.n2939 gnd.n2263 240.244
R6650 gnd.n2939 gnd.n2265 240.244
R6651 gnd.n2935 gnd.n2265 240.244
R6652 gnd.n2935 gnd.n2271 240.244
R6653 gnd.n2931 gnd.n2271 240.244
R6654 gnd.n2931 gnd.n2273 240.244
R6655 gnd.n2927 gnd.n2273 240.244
R6656 gnd.n2927 gnd.n2279 240.244
R6657 gnd.n2923 gnd.n2279 240.244
R6658 gnd.n2923 gnd.n2281 240.244
R6659 gnd.n2919 gnd.n2281 240.244
R6660 gnd.n2919 gnd.n2287 240.244
R6661 gnd.n2915 gnd.n2287 240.244
R6662 gnd.n2915 gnd.n2289 240.244
R6663 gnd.n2911 gnd.n2289 240.244
R6664 gnd.n2911 gnd.n2295 240.244
R6665 gnd.n2907 gnd.n2295 240.244
R6666 gnd.n2907 gnd.n2297 240.244
R6667 gnd.n2903 gnd.n2297 240.244
R6668 gnd.n2903 gnd.n2303 240.244
R6669 gnd.n2899 gnd.n2303 240.244
R6670 gnd.n2899 gnd.n2305 240.244
R6671 gnd.n2895 gnd.n2305 240.244
R6672 gnd.n2895 gnd.n2311 240.244
R6673 gnd.n2891 gnd.n2311 240.244
R6674 gnd.n2891 gnd.n2313 240.244
R6675 gnd.n2887 gnd.n2313 240.244
R6676 gnd.n2887 gnd.n2319 240.244
R6677 gnd.n2883 gnd.n2319 240.244
R6678 gnd.n2883 gnd.n2321 240.244
R6679 gnd.n2879 gnd.n2321 240.244
R6680 gnd.n2879 gnd.n2327 240.244
R6681 gnd.n2875 gnd.n2327 240.244
R6682 gnd.n2875 gnd.n2329 240.244
R6683 gnd.n2871 gnd.n2329 240.244
R6684 gnd.n2871 gnd.n2335 240.244
R6685 gnd.n2867 gnd.n2335 240.244
R6686 gnd.n2867 gnd.n2337 240.244
R6687 gnd.n2863 gnd.n2337 240.244
R6688 gnd.n2863 gnd.n2343 240.244
R6689 gnd.n2859 gnd.n2343 240.244
R6690 gnd.n2859 gnd.n2345 240.244
R6691 gnd.n2855 gnd.n2345 240.244
R6692 gnd.n2855 gnd.n2351 240.244
R6693 gnd.n2851 gnd.n2351 240.244
R6694 gnd.n2851 gnd.n2353 240.244
R6695 gnd.n2847 gnd.n2353 240.244
R6696 gnd.n2847 gnd.n2359 240.244
R6697 gnd.n2843 gnd.n2359 240.244
R6698 gnd.n2843 gnd.n2361 240.244
R6699 gnd.n2839 gnd.n2361 240.244
R6700 gnd.n2839 gnd.n2367 240.244
R6701 gnd.n2835 gnd.n2367 240.244
R6702 gnd.n2835 gnd.n2369 240.244
R6703 gnd.n2831 gnd.n2369 240.244
R6704 gnd.n2831 gnd.n2375 240.244
R6705 gnd.n2827 gnd.n2375 240.244
R6706 gnd.n2827 gnd.n2377 240.244
R6707 gnd.n2823 gnd.n2377 240.244
R6708 gnd.n2823 gnd.n2383 240.244
R6709 gnd.n2819 gnd.n2383 240.244
R6710 gnd.n2819 gnd.n2385 240.244
R6711 gnd.n2815 gnd.n2385 240.244
R6712 gnd.n2815 gnd.n2391 240.244
R6713 gnd.n2811 gnd.n2391 240.244
R6714 gnd.n2811 gnd.n2393 240.244
R6715 gnd.n2807 gnd.n2393 240.244
R6716 gnd.n2807 gnd.n2399 240.244
R6717 gnd.n2803 gnd.n2399 240.244
R6718 gnd.n2803 gnd.n2401 240.244
R6719 gnd.n2799 gnd.n2401 240.244
R6720 gnd.n2799 gnd.n2407 240.244
R6721 gnd.n2795 gnd.n2407 240.244
R6722 gnd.n2795 gnd.n2409 240.244
R6723 gnd.n2791 gnd.n2409 240.244
R6724 gnd.n2791 gnd.n2415 240.244
R6725 gnd.n2787 gnd.n2415 240.244
R6726 gnd.n2787 gnd.n2417 240.244
R6727 gnd.n2783 gnd.n2417 240.244
R6728 gnd.n2783 gnd.n2423 240.244
R6729 gnd.n2779 gnd.n2423 240.244
R6730 gnd.n2779 gnd.n2425 240.244
R6731 gnd.n2775 gnd.n2425 240.244
R6732 gnd.n2775 gnd.n2431 240.244
R6733 gnd.n2771 gnd.n2433 240.244
R6734 gnd.n2439 gnd.n2433 240.244
R6735 gnd.n2764 gnd.n2439 240.244
R6736 gnd.n2764 gnd.n2440 240.244
R6737 gnd.n2760 gnd.n2440 240.244
R6738 gnd.n2760 gnd.n2443 240.244
R6739 gnd.n2756 gnd.n2443 240.244
R6740 gnd.n2756 gnd.n2448 240.244
R6741 gnd.n2752 gnd.n2448 240.244
R6742 gnd.n2752 gnd.n2450 240.244
R6743 gnd.n2748 gnd.n2450 240.244
R6744 gnd.n2748 gnd.n2456 240.244
R6745 gnd.n2744 gnd.n2456 240.244
R6746 gnd.n2744 gnd.n2458 240.244
R6747 gnd.n2740 gnd.n2458 240.244
R6748 gnd.n2740 gnd.n2464 240.244
R6749 gnd.n2736 gnd.n2464 240.244
R6750 gnd.n2736 gnd.n2466 240.244
R6751 gnd.n2732 gnd.n2466 240.244
R6752 gnd.n2732 gnd.n2472 240.244
R6753 gnd.n2728 gnd.n2472 240.244
R6754 gnd.n2728 gnd.n2474 240.244
R6755 gnd.n2724 gnd.n2474 240.244
R6756 gnd.n2724 gnd.n2480 240.244
R6757 gnd.n2720 gnd.n2480 240.244
R6758 gnd.n2720 gnd.n2482 240.244
R6759 gnd.n2716 gnd.n2482 240.244
R6760 gnd.n2716 gnd.n2488 240.244
R6761 gnd.n2712 gnd.n2488 240.244
R6762 gnd.n2712 gnd.n2490 240.244
R6763 gnd.n2708 gnd.n2490 240.244
R6764 gnd.n2708 gnd.n2496 240.244
R6765 gnd.n2704 gnd.n2496 240.244
R6766 gnd.n2704 gnd.n2498 240.244
R6767 gnd.n2700 gnd.n2498 240.244
R6768 gnd.n2700 gnd.n2504 240.244
R6769 gnd.n2696 gnd.n2504 240.244
R6770 gnd.n2696 gnd.n2506 240.244
R6771 gnd.n2692 gnd.n2506 240.244
R6772 gnd.n2692 gnd.n2512 240.244
R6773 gnd.n2688 gnd.n2512 240.244
R6774 gnd.n2688 gnd.n2514 240.244
R6775 gnd.n2684 gnd.n2514 240.244
R6776 gnd.n2684 gnd.n2520 240.244
R6777 gnd.n2680 gnd.n2520 240.244
R6778 gnd.n2680 gnd.n2522 240.244
R6779 gnd.n2676 gnd.n2522 240.244
R6780 gnd.n2676 gnd.n2528 240.244
R6781 gnd.n2672 gnd.n2528 240.244
R6782 gnd.n2672 gnd.n2530 240.244
R6783 gnd.n2668 gnd.n2530 240.244
R6784 gnd.n2668 gnd.n2536 240.244
R6785 gnd.n2664 gnd.n2536 240.244
R6786 gnd.n2664 gnd.n2538 240.244
R6787 gnd.n2660 gnd.n2538 240.244
R6788 gnd.n2660 gnd.n2544 240.244
R6789 gnd.n2656 gnd.n2544 240.244
R6790 gnd.n2656 gnd.n2546 240.244
R6791 gnd.n2652 gnd.n2546 240.244
R6792 gnd.n2652 gnd.n2552 240.244
R6793 gnd.n2648 gnd.n2552 240.244
R6794 gnd.n2648 gnd.n2554 240.244
R6795 gnd.n2644 gnd.n2554 240.244
R6796 gnd.n2644 gnd.n2560 240.244
R6797 gnd.n2640 gnd.n2560 240.244
R6798 gnd.n2640 gnd.n2562 240.244
R6799 gnd.n2636 gnd.n2562 240.244
R6800 gnd.n2636 gnd.n2568 240.244
R6801 gnd.n2632 gnd.n2568 240.244
R6802 gnd.n2632 gnd.n2570 240.244
R6803 gnd.n2628 gnd.n2570 240.244
R6804 gnd.n2628 gnd.n2576 240.244
R6805 gnd.n2624 gnd.n2576 240.244
R6806 gnd.n2624 gnd.n2578 240.244
R6807 gnd.n2620 gnd.n2578 240.244
R6808 gnd.n2620 gnd.n2584 240.244
R6809 gnd.n2616 gnd.n2584 240.244
R6810 gnd.n2616 gnd.n2586 240.244
R6811 gnd.n2612 gnd.n2586 240.244
R6812 gnd.n2612 gnd.n2592 240.244
R6813 gnd.n2608 gnd.n2592 240.244
R6814 gnd.n2608 gnd.n2594 240.244
R6815 gnd.n2604 gnd.n2594 240.244
R6816 gnd.n2604 gnd.n2601 240.244
R6817 gnd.n1973 gnd.n1912 240.244
R6818 gnd.n1969 gnd.n1912 240.244
R6819 gnd.n1969 gnd.n1968 240.244
R6820 gnd.n1968 gnd.n1967 240.244
R6821 gnd.n1967 gnd.n1914 240.244
R6822 gnd.n1962 gnd.n1914 240.244
R6823 gnd.n1962 gnd.n1961 240.244
R6824 gnd.n1961 gnd.n1960 240.244
R6825 gnd.n1960 gnd.n1917 240.244
R6826 gnd.n1956 gnd.n1917 240.244
R6827 gnd.n1956 gnd.n1955 240.244
R6828 gnd.n1955 gnd.n1954 240.244
R6829 gnd.n1954 gnd.n1921 240.244
R6830 gnd.n1950 gnd.n1921 240.244
R6831 gnd.n1950 gnd.n1949 240.244
R6832 gnd.n1949 gnd.n1948 240.244
R6833 gnd.n1948 gnd.n1927 240.244
R6834 gnd.n1944 gnd.n1927 240.244
R6835 gnd.n1944 gnd.n1943 240.244
R6836 gnd.n1943 gnd.n1942 240.244
R6837 gnd.n1942 gnd.n1933 240.244
R6838 gnd.n1933 gnd.n1548 240.244
R6839 gnd.n5388 gnd.n1548 240.244
R6840 gnd.n5389 gnd.n5388 240.244
R6841 gnd.n5390 gnd.n5389 240.244
R6842 gnd.n5390 gnd.n1543 240.244
R6843 gnd.n5401 gnd.n1543 240.244
R6844 gnd.n5401 gnd.n1544 240.244
R6845 gnd.n5397 gnd.n1544 240.244
R6846 gnd.n5397 gnd.n1497 240.244
R6847 gnd.n5454 gnd.n1497 240.244
R6848 gnd.n5454 gnd.n1493 240.244
R6849 gnd.n5460 gnd.n1493 240.244
R6850 gnd.n5461 gnd.n5460 240.244
R6851 gnd.n5462 gnd.n5461 240.244
R6852 gnd.n5462 gnd.n1488 240.244
R6853 gnd.n5696 gnd.n1488 240.244
R6854 gnd.n5696 gnd.n1489 240.244
R6855 gnd.n5692 gnd.n1489 240.244
R6856 gnd.n5692 gnd.n5689 240.244
R6857 gnd.n5689 gnd.n5688 240.244
R6858 gnd.n5688 gnd.n5470 240.244
R6859 gnd.n5684 gnd.n5470 240.244
R6860 gnd.n5684 gnd.n5476 240.244
R6861 gnd.n5549 gnd.n5476 240.244
R6862 gnd.n5569 gnd.n5549 240.244
R6863 gnd.n5569 gnd.n5544 240.244
R6864 gnd.n5575 gnd.n5544 240.244
R6865 gnd.n5575 gnd.n5536 240.244
R6866 gnd.n5590 gnd.n5536 240.244
R6867 gnd.n5590 gnd.n5532 240.244
R6868 gnd.n5596 gnd.n5532 240.244
R6869 gnd.n5596 gnd.n5524 240.244
R6870 gnd.n5611 gnd.n5524 240.244
R6871 gnd.n5611 gnd.n5520 240.244
R6872 gnd.n5617 gnd.n5520 240.244
R6873 gnd.n5617 gnd.n5511 240.244
R6874 gnd.n5640 gnd.n5511 240.244
R6875 gnd.n5640 gnd.n5506 240.244
R6876 gnd.n5651 gnd.n5506 240.244
R6877 gnd.n5651 gnd.n5507 240.244
R6878 gnd.n5647 gnd.n5507 240.244
R6879 gnd.n5647 gnd.n1199 240.244
R6880 gnd.n6155 gnd.n1199 240.244
R6881 gnd.n6155 gnd.n1195 240.244
R6882 gnd.n6161 gnd.n1195 240.244
R6883 gnd.n6161 gnd.n1173 240.244
R6884 gnd.n6196 gnd.n1173 240.244
R6885 gnd.n6196 gnd.n1168 240.244
R6886 gnd.n6206 gnd.n1168 240.244
R6887 gnd.n6206 gnd.n1169 240.244
R6888 gnd.n1169 gnd.n1151 240.244
R6889 gnd.n6223 gnd.n1151 240.244
R6890 gnd.n6224 gnd.n6223 240.244
R6891 gnd.n6224 gnd.n1147 240.244
R6892 gnd.n6231 gnd.n1147 240.244
R6893 gnd.n6231 gnd.n1118 240.244
R6894 gnd.n6285 gnd.n1118 240.244
R6895 gnd.n6285 gnd.n1119 240.244
R6896 gnd.n6281 gnd.n1119 240.244
R6897 gnd.n6281 gnd.n1086 240.244
R6898 gnd.n6347 gnd.n1086 240.244
R6899 gnd.n6347 gnd.n1087 240.244
R6900 gnd.n6343 gnd.n1087 240.244
R6901 gnd.n6343 gnd.n1059 240.244
R6902 gnd.n6385 gnd.n1059 240.244
R6903 gnd.n6385 gnd.n1060 240.244
R6904 gnd.n6381 gnd.n1060 240.244
R6905 gnd.n6381 gnd.n1029 240.244
R6906 gnd.n6424 gnd.n1029 240.244
R6907 gnd.n6424 gnd.n1030 240.244
R6908 gnd.n6420 gnd.n1030 240.244
R6909 gnd.n6420 gnd.n1038 240.244
R6910 gnd.n1038 gnd.n983 240.244
R6911 gnd.n6488 gnd.n983 240.244
R6912 gnd.n6488 gnd.n984 240.244
R6913 gnd.n6484 gnd.n984 240.244
R6914 gnd.n6484 gnd.n6483 240.244
R6915 gnd.n6483 gnd.n944 240.244
R6916 gnd.n6540 gnd.n944 240.244
R6917 gnd.n6540 gnd.n940 240.244
R6918 gnd.n6546 gnd.n940 240.244
R6919 gnd.n6546 gnd.n890 240.244
R6920 gnd.n6716 gnd.n890 240.244
R6921 gnd.n6716 gnd.n885 240.244
R6922 gnd.n6724 gnd.n885 240.244
R6923 gnd.n6724 gnd.n886 240.244
R6924 gnd.n886 gnd.n866 240.244
R6925 gnd.n6746 gnd.n866 240.244
R6926 gnd.n6746 gnd.n861 240.244
R6927 gnd.n6754 gnd.n861 240.244
R6928 gnd.n6754 gnd.n862 240.244
R6929 gnd.n862 gnd.n841 240.244
R6930 gnd.n6776 gnd.n841 240.244
R6931 gnd.n6776 gnd.n836 240.244
R6932 gnd.n6784 gnd.n836 240.244
R6933 gnd.n6784 gnd.n837 240.244
R6934 gnd.n837 gnd.n816 240.244
R6935 gnd.n6811 gnd.n816 240.244
R6936 gnd.n6811 gnd.n812 240.244
R6937 gnd.n6820 gnd.n812 240.244
R6938 gnd.n6820 gnd.n800 240.244
R6939 gnd.n6833 gnd.n800 240.244
R6940 gnd.n6834 gnd.n6833 240.244
R6941 gnd.n6835 gnd.n6834 240.244
R6942 gnd.n6835 gnd.n796 240.244
R6943 gnd.n6843 gnd.n796 240.244
R6944 gnd.n6843 gnd.n588 240.244
R6945 gnd.n7043 gnd.n588 240.244
R6946 gnd.n7044 gnd.n7043 240.244
R6947 gnd.n7044 gnd.n583 240.244
R6948 gnd.n7058 gnd.n583 240.244
R6949 gnd.n7058 gnd.n584 240.244
R6950 gnd.n7054 gnd.n584 240.244
R6951 gnd.n7054 gnd.n7053 240.244
R6952 gnd.n7053 gnd.n550 240.244
R6953 gnd.n7101 gnd.n550 240.244
R6954 gnd.n7101 gnd.n544 240.244
R6955 gnd.n7109 gnd.n544 240.244
R6956 gnd.n7109 gnd.n546 240.244
R6957 gnd.n546 gnd.n486 240.244
R6958 gnd.n7163 gnd.n486 240.244
R6959 gnd.n7163 gnd.n482 240.244
R6960 gnd.n7169 gnd.n482 240.244
R6961 gnd.n7170 gnd.n7169 240.244
R6962 gnd.n7171 gnd.n7170 240.244
R6963 gnd.n7171 gnd.n477 240.244
R6964 gnd.n7179 gnd.n477 240.244
R6965 gnd.n7179 gnd.n478 240.244
R6966 gnd.n478 gnd.n430 240.244
R6967 gnd.n7238 gnd.n430 240.244
R6968 gnd.n7238 gnd.n425 240.244
R6969 gnd.n7256 gnd.n425 240.244
R6970 gnd.n7256 gnd.n426 240.244
R6971 gnd.n7252 gnd.n426 240.244
R6972 gnd.n7252 gnd.n7251 240.244
R6973 gnd.n7251 gnd.n7250 240.244
R6974 gnd.n7250 gnd.n383 240.244
R6975 gnd.n7314 gnd.n383 240.244
R6976 gnd.n7314 gnd.n380 240.244
R6977 gnd.n7321 gnd.n380 240.244
R6978 gnd.n7321 gnd.n381 240.244
R6979 gnd.n381 gnd.n359 240.244
R6980 gnd.n7345 gnd.n359 240.244
R6981 gnd.n7345 gnd.n356 240.244
R6982 gnd.n7351 gnd.n356 240.244
R6983 gnd.n7351 gnd.n357 240.244
R6984 gnd.n3113 gnd.n2098 240.244
R6985 gnd.n3113 gnd.n2094 240.244
R6986 gnd.n3119 gnd.n2094 240.244
R6987 gnd.n3119 gnd.n2092 240.244
R6988 gnd.n3123 gnd.n2092 240.244
R6989 gnd.n3123 gnd.n2088 240.244
R6990 gnd.n3129 gnd.n2088 240.244
R6991 gnd.n3129 gnd.n2086 240.244
R6992 gnd.n3133 gnd.n2086 240.244
R6993 gnd.n3133 gnd.n2082 240.244
R6994 gnd.n3139 gnd.n2082 240.244
R6995 gnd.n3139 gnd.n2080 240.244
R6996 gnd.n3143 gnd.n2080 240.244
R6997 gnd.n3143 gnd.n2076 240.244
R6998 gnd.n3149 gnd.n2076 240.244
R6999 gnd.n3149 gnd.n2074 240.244
R7000 gnd.n3153 gnd.n2074 240.244
R7001 gnd.n3153 gnd.n2070 240.244
R7002 gnd.n3159 gnd.n2070 240.244
R7003 gnd.n3159 gnd.n2068 240.244
R7004 gnd.n3163 gnd.n2068 240.244
R7005 gnd.n3163 gnd.n2064 240.244
R7006 gnd.n3169 gnd.n2064 240.244
R7007 gnd.n3169 gnd.n2062 240.244
R7008 gnd.n3173 gnd.n2062 240.244
R7009 gnd.n3173 gnd.n2058 240.244
R7010 gnd.n3179 gnd.n2058 240.244
R7011 gnd.n3179 gnd.n2056 240.244
R7012 gnd.n3183 gnd.n2056 240.244
R7013 gnd.n3183 gnd.n2052 240.244
R7014 gnd.n3189 gnd.n2052 240.244
R7015 gnd.n3189 gnd.n2050 240.244
R7016 gnd.n3193 gnd.n2050 240.244
R7017 gnd.n3193 gnd.n2046 240.244
R7018 gnd.n3199 gnd.n2046 240.244
R7019 gnd.n3199 gnd.n2044 240.244
R7020 gnd.n3203 gnd.n2044 240.244
R7021 gnd.n3203 gnd.n2040 240.244
R7022 gnd.n3209 gnd.n2040 240.244
R7023 gnd.n3209 gnd.n2038 240.244
R7024 gnd.n3213 gnd.n2038 240.244
R7025 gnd.n3213 gnd.n2034 240.244
R7026 gnd.n3219 gnd.n2034 240.244
R7027 gnd.n3219 gnd.n2032 240.244
R7028 gnd.n3223 gnd.n2032 240.244
R7029 gnd.n3223 gnd.n2028 240.244
R7030 gnd.n3229 gnd.n2028 240.244
R7031 gnd.n3229 gnd.n2026 240.244
R7032 gnd.n3233 gnd.n2026 240.244
R7033 gnd.n3233 gnd.n2022 240.244
R7034 gnd.n3239 gnd.n2022 240.244
R7035 gnd.n3239 gnd.n2020 240.244
R7036 gnd.n3243 gnd.n2020 240.244
R7037 gnd.n3243 gnd.n2016 240.244
R7038 gnd.n3249 gnd.n2016 240.244
R7039 gnd.n3249 gnd.n2014 240.244
R7040 gnd.n3253 gnd.n2014 240.244
R7041 gnd.n3253 gnd.n2010 240.244
R7042 gnd.n3259 gnd.n2010 240.244
R7043 gnd.n3259 gnd.n2008 240.244
R7044 gnd.n3263 gnd.n2008 240.244
R7045 gnd.n3263 gnd.n2004 240.244
R7046 gnd.n3269 gnd.n2004 240.244
R7047 gnd.n3269 gnd.n2002 240.244
R7048 gnd.n3273 gnd.n2002 240.244
R7049 gnd.n3273 gnd.n1998 240.244
R7050 gnd.n3279 gnd.n1998 240.244
R7051 gnd.n3279 gnd.n1996 240.244
R7052 gnd.n3283 gnd.n1996 240.244
R7053 gnd.n3283 gnd.n1992 240.244
R7054 gnd.n3289 gnd.n1992 240.244
R7055 gnd.n3289 gnd.n1990 240.244
R7056 gnd.n3293 gnd.n1990 240.244
R7057 gnd.n3293 gnd.n1986 240.244
R7058 gnd.n3299 gnd.n1986 240.244
R7059 gnd.n3299 gnd.n1984 240.244
R7060 gnd.n3303 gnd.n1984 240.244
R7061 gnd.n3303 gnd.n1980 240.244
R7062 gnd.n3309 gnd.n1980 240.244
R7063 gnd.n3309 gnd.n1978 240.244
R7064 gnd.n3313 gnd.n1978 240.244
R7065 gnd.n3313 gnd.n1911 240.244
R7066 gnd.n3321 gnd.n1911 240.244
R7067 gnd.n3321 gnd.n1974 240.244
R7068 gnd.n5681 gnd.n1477 240.244
R7069 gnd.n5681 gnd.n5481 240.244
R7070 gnd.n5486 gnd.n5481 240.244
R7071 gnd.n5487 gnd.n5486 240.244
R7072 gnd.n5488 gnd.n5487 240.244
R7073 gnd.n5578 gnd.n5488 240.244
R7074 gnd.n5578 gnd.n5491 240.244
R7075 gnd.n5492 gnd.n5491 240.244
R7076 gnd.n5493 gnd.n5492 240.244
R7077 gnd.n5599 gnd.n5493 240.244
R7078 gnd.n5599 gnd.n5496 240.244
R7079 gnd.n5497 gnd.n5496 240.244
R7080 gnd.n5498 gnd.n5497 240.244
R7081 gnd.n5620 gnd.n5498 240.244
R7082 gnd.n5620 gnd.n5501 240.244
R7083 gnd.n5502 gnd.n5501 240.244
R7084 gnd.n5654 gnd.n5502 240.244
R7085 gnd.n5654 gnd.n1225 240.244
R7086 gnd.n6101 gnd.n1225 240.244
R7087 gnd.n6101 gnd.n1219 240.244
R7088 gnd.n6108 gnd.n1219 240.244
R7089 gnd.n6108 gnd.n1220 240.244
R7090 gnd.n1220 gnd.n1183 240.244
R7091 gnd.n6177 gnd.n1183 240.244
R7092 gnd.n6177 gnd.n1177 240.244
R7093 gnd.n6193 gnd.n1177 240.244
R7094 gnd.n6193 gnd.n1178 240.244
R7095 gnd.n6182 gnd.n1178 240.244
R7096 gnd.n6183 gnd.n6182 240.244
R7097 gnd.n6184 gnd.n6183 240.244
R7098 gnd.n6184 gnd.n1134 240.244
R7099 gnd.n6253 gnd.n1134 240.244
R7100 gnd.n6253 gnd.n1130 240.244
R7101 gnd.n6259 gnd.n1130 240.244
R7102 gnd.n6259 gnd.n1106 240.244
R7103 gnd.n6299 gnd.n1106 240.244
R7104 gnd.n6299 gnd.n1102 240.244
R7105 gnd.n6305 gnd.n1102 240.244
R7106 gnd.n6305 gnd.n1075 240.244
R7107 gnd.n6361 gnd.n1075 240.244
R7108 gnd.n6361 gnd.n1071 240.244
R7109 gnd.n6367 gnd.n1071 240.244
R7110 gnd.n6367 gnd.n1048 240.244
R7111 gnd.n6398 gnd.n1048 240.244
R7112 gnd.n6398 gnd.n1044 240.244
R7113 gnd.n6404 gnd.n1044 240.244
R7114 gnd.n6404 gnd.n1019 240.244
R7115 gnd.n6434 gnd.n1019 240.244
R7116 gnd.n6434 gnd.n1015 240.244
R7117 gnd.n6440 gnd.n1015 240.244
R7118 gnd.n6440 gnd.n980 240.244
R7119 gnd.n6491 gnd.n980 240.244
R7120 gnd.n6491 gnd.n974 240.244
R7121 gnd.n6498 gnd.n974 240.244
R7122 gnd.n6498 gnd.n975 240.244
R7123 gnd.n975 gnd.n955 240.244
R7124 gnd.n6530 gnd.n955 240.244
R7125 gnd.n6530 gnd.n948 240.244
R7126 gnd.n960 gnd.n948 240.244
R7127 gnd.n6520 gnd.n960 240.244
R7128 gnd.n6521 gnd.n6520 240.244
R7129 gnd.n6521 gnd.n882 240.244
R7130 gnd.n6727 gnd.n882 240.244
R7131 gnd.n6727 gnd.n875 240.244
R7132 gnd.n6734 gnd.n875 240.244
R7133 gnd.n6734 gnd.n877 240.244
R7134 gnd.n877 gnd.n857 240.244
R7135 gnd.n6757 gnd.n857 240.244
R7136 gnd.n6757 gnd.n850 240.244
R7137 gnd.n6764 gnd.n850 240.244
R7138 gnd.n6764 gnd.n852 240.244
R7139 gnd.n852 gnd.n832 240.244
R7140 gnd.n6787 gnd.n832 240.244
R7141 gnd.n6787 gnd.n826 240.244
R7142 gnd.n6794 gnd.n826 240.244
R7143 gnd.n6794 gnd.n827 240.244
R7144 gnd.n827 gnd.n808 240.244
R7145 gnd.n6823 gnd.n808 240.244
R7146 gnd.n6823 gnd.n804 240.244
R7147 gnd.n6829 gnd.n804 240.244
R7148 gnd.n6829 gnd.n765 240.244
R7149 gnd.n6860 gnd.n765 240.244
R7150 gnd.n1476 gnd.n1475 240.244
R7151 gnd.n1481 gnd.n1475 240.244
R7152 gnd.n1483 gnd.n1482 240.244
R7153 gnd.n1485 gnd.n1484 240.244
R7154 gnd.n5705 gnd.n5704 240.244
R7155 gnd.n5708 gnd.n5707 240.244
R7156 gnd.n5719 gnd.n5718 240.244
R7157 gnd.n5721 gnd.n5720 240.244
R7158 gnd.n5731 gnd.n5730 240.244
R7159 gnd.n5742 gnd.n5741 240.244
R7160 gnd.n5744 gnd.n5743 240.244
R7161 gnd.n5754 gnd.n5753 240.244
R7162 gnd.n5775 gnd.n5774 240.244
R7163 gnd.n1472 gnd.n1458 240.244
R7164 gnd.n5479 gnd.n1459 240.244
R7165 gnd.n5559 gnd.n5479 240.244
R7166 gnd.n5559 gnd.n5551 240.244
R7167 gnd.n5565 gnd.n5551 240.244
R7168 gnd.n5565 gnd.n5542 240.244
R7169 gnd.n5580 gnd.n5542 240.244
R7170 gnd.n5580 gnd.n5538 240.244
R7171 gnd.n5586 gnd.n5538 240.244
R7172 gnd.n5586 gnd.n5530 240.244
R7173 gnd.n5601 gnd.n5530 240.244
R7174 gnd.n5601 gnd.n5526 240.244
R7175 gnd.n5607 gnd.n5526 240.244
R7176 gnd.n5607 gnd.n5518 240.244
R7177 gnd.n5622 gnd.n5518 240.244
R7178 gnd.n5622 gnd.n5513 240.244
R7179 gnd.n5637 gnd.n5513 240.244
R7180 gnd.n5637 gnd.n5504 240.244
R7181 gnd.n5627 gnd.n5504 240.244
R7182 gnd.n5627 gnd.n1227 240.244
R7183 gnd.n1227 gnd.n1217 240.244
R7184 gnd.n6110 gnd.n1217 240.244
R7185 gnd.n6111 gnd.n6110 240.244
R7186 gnd.n6111 gnd.n1193 240.244
R7187 gnd.n1193 gnd.n1185 240.244
R7188 gnd.n6144 gnd.n1185 240.244
R7189 gnd.n6144 gnd.n1175 240.244
R7190 gnd.n6117 gnd.n1175 240.244
R7191 gnd.n6118 gnd.n6117 240.244
R7192 gnd.n6119 gnd.n6118 240.244
R7193 gnd.n6120 gnd.n6119 240.244
R7194 gnd.n6120 gnd.n1143 240.244
R7195 gnd.n1143 gnd.n1136 240.244
R7196 gnd.n1146 gnd.n1136 240.244
R7197 gnd.n1146 gnd.n1129 240.244
R7198 gnd.n1129 gnd.n1116 240.244
R7199 gnd.n1116 gnd.n1107 240.244
R7200 gnd.n1107 gnd.n1098 240.244
R7201 gnd.n6307 gnd.n1098 240.244
R7202 gnd.n6307 gnd.n1085 240.244
R7203 gnd.n1085 gnd.n1077 240.244
R7204 gnd.n6340 gnd.n1077 240.244
R7205 gnd.n6340 gnd.n1070 240.244
R7206 gnd.n6313 gnd.n1070 240.244
R7207 gnd.n6313 gnd.n1050 240.244
R7208 gnd.n6314 gnd.n1050 240.244
R7209 gnd.n6314 gnd.n1043 240.244
R7210 gnd.n6317 gnd.n1043 240.244
R7211 gnd.n6317 gnd.n1020 240.244
R7212 gnd.n6318 gnd.n1020 240.244
R7213 gnd.n6318 gnd.n1012 240.244
R7214 gnd.n6321 gnd.n1012 240.244
R7215 gnd.n6321 gnd.n982 240.244
R7216 gnd.n982 gnd.n970 240.244
R7217 gnd.n6500 gnd.n970 240.244
R7218 gnd.n6500 gnd.n971 240.244
R7219 gnd.n971 gnd.n967 240.244
R7220 gnd.n967 gnd.n954 240.244
R7221 gnd.n954 gnd.n947 240.244
R7222 gnd.n961 gnd.n947 240.244
R7223 gnd.n6517 gnd.n961 240.244
R7224 gnd.n6517 gnd.n962 240.244
R7225 gnd.n962 gnd.n892 240.244
R7226 gnd.n892 gnd.n883 240.244
R7227 gnd.n883 gnd.n872 240.244
R7228 gnd.n6736 gnd.n872 240.244
R7229 gnd.n6736 gnd.n867 240.244
R7230 gnd.n6743 gnd.n867 240.244
R7231 gnd.n6743 gnd.n859 240.244
R7232 gnd.n859 gnd.n847 240.244
R7233 gnd.n6766 gnd.n847 240.244
R7234 gnd.n6766 gnd.n842 240.244
R7235 gnd.n6773 gnd.n842 240.244
R7236 gnd.n6773 gnd.n834 240.244
R7237 gnd.n834 gnd.n823 240.244
R7238 gnd.n6796 gnd.n823 240.244
R7239 gnd.n6796 gnd.n818 240.244
R7240 gnd.n6808 gnd.n818 240.244
R7241 gnd.n6808 gnd.n810 240.244
R7242 gnd.n6801 gnd.n810 240.244
R7243 gnd.n6801 gnd.n803 240.244
R7244 gnd.n803 gnd.n761 240.244
R7245 gnd.n6862 gnd.n761 240.244
R7246 gnd.n771 gnd.n770 240.244
R7247 gnd.n778 gnd.n774 240.244
R7248 gnd.n6848 gnd.n6847 240.244
R7249 gnd.n699 gnd.n698 240.244
R7250 gnd.n781 gnd.n700 240.244
R7251 gnd.n710 gnd.n709 240.244
R7252 gnd.n783 gnd.n719 240.244
R7253 gnd.n786 gnd.n720 240.244
R7254 gnd.n728 gnd.n727 240.244
R7255 gnd.n788 gnd.n737 240.244
R7256 gnd.n791 gnd.n738 240.244
R7257 gnd.n746 gnd.n745 240.244
R7258 gnd.n793 gnd.n746 240.244
R7259 gnd.n757 gnd.n756 240.244
R7260 gnd.n1272 gnd.n1271 240.132
R7261 gnd.n6563 gnd.n6562 240.132
R7262 gnd.n3110 gnd.n2099 225.874
R7263 gnd.n3102 gnd.n2099 225.874
R7264 gnd.n3102 gnd.n3101 225.874
R7265 gnd.n3101 gnd.n3100 225.874
R7266 gnd.n3100 gnd.n2105 225.874
R7267 gnd.n3094 gnd.n2105 225.874
R7268 gnd.n3094 gnd.n3093 225.874
R7269 gnd.n3093 gnd.n3092 225.874
R7270 gnd.n3092 gnd.n2112 225.874
R7271 gnd.n3086 gnd.n2112 225.874
R7272 gnd.n3086 gnd.n3085 225.874
R7273 gnd.n3085 gnd.n3084 225.874
R7274 gnd.n3084 gnd.n2120 225.874
R7275 gnd.n3078 gnd.n2120 225.874
R7276 gnd.n3078 gnd.n3077 225.874
R7277 gnd.n3077 gnd.n3076 225.874
R7278 gnd.n3076 gnd.n2128 225.874
R7279 gnd.n3070 gnd.n2128 225.874
R7280 gnd.n3070 gnd.n3069 225.874
R7281 gnd.n3069 gnd.n3068 225.874
R7282 gnd.n3068 gnd.n2136 225.874
R7283 gnd.n3062 gnd.n2136 225.874
R7284 gnd.n3062 gnd.n3061 225.874
R7285 gnd.n3061 gnd.n3060 225.874
R7286 gnd.n3060 gnd.n2144 225.874
R7287 gnd.n3054 gnd.n2144 225.874
R7288 gnd.n3054 gnd.n3053 225.874
R7289 gnd.n3053 gnd.n3052 225.874
R7290 gnd.n3052 gnd.n2152 225.874
R7291 gnd.n3046 gnd.n2152 225.874
R7292 gnd.n3046 gnd.n3045 225.874
R7293 gnd.n3045 gnd.n3044 225.874
R7294 gnd.n3044 gnd.n2160 225.874
R7295 gnd.n3038 gnd.n2160 225.874
R7296 gnd.n3038 gnd.n3037 225.874
R7297 gnd.n3037 gnd.n3036 225.874
R7298 gnd.n3036 gnd.n2168 225.874
R7299 gnd.n3030 gnd.n2168 225.874
R7300 gnd.n3030 gnd.n3029 225.874
R7301 gnd.n3029 gnd.n3028 225.874
R7302 gnd.n3028 gnd.n2176 225.874
R7303 gnd.n3022 gnd.n2176 225.874
R7304 gnd.n3022 gnd.n3021 225.874
R7305 gnd.n3021 gnd.n3020 225.874
R7306 gnd.n3020 gnd.n2184 225.874
R7307 gnd.n3014 gnd.n2184 225.874
R7308 gnd.n3014 gnd.n3013 225.874
R7309 gnd.n3013 gnd.n3012 225.874
R7310 gnd.n3012 gnd.n2192 225.874
R7311 gnd.n3006 gnd.n2192 225.874
R7312 gnd.n3006 gnd.n3005 225.874
R7313 gnd.n3005 gnd.n3004 225.874
R7314 gnd.n3004 gnd.n2200 225.874
R7315 gnd.n2998 gnd.n2200 225.874
R7316 gnd.n2998 gnd.n2997 225.874
R7317 gnd.n2997 gnd.n2996 225.874
R7318 gnd.n2996 gnd.n2208 225.874
R7319 gnd.n2990 gnd.n2208 225.874
R7320 gnd.n2990 gnd.n2989 225.874
R7321 gnd.n2989 gnd.n2988 225.874
R7322 gnd.n2988 gnd.n2216 225.874
R7323 gnd.n2982 gnd.n2216 225.874
R7324 gnd.n2982 gnd.n2981 225.874
R7325 gnd.n2981 gnd.n2980 225.874
R7326 gnd.n2980 gnd.n2224 225.874
R7327 gnd.n2974 gnd.n2224 225.874
R7328 gnd.n2974 gnd.n2973 225.874
R7329 gnd.n2973 gnd.n2972 225.874
R7330 gnd.n2972 gnd.n2232 225.874
R7331 gnd.n2966 gnd.n2232 225.874
R7332 gnd.n2966 gnd.n2965 225.874
R7333 gnd.n2965 gnd.n2964 225.874
R7334 gnd.n2964 gnd.n2240 225.874
R7335 gnd.n2958 gnd.n2240 225.874
R7336 gnd.n2958 gnd.n2957 225.874
R7337 gnd.n2957 gnd.n2956 225.874
R7338 gnd.n2956 gnd.n2248 225.874
R7339 gnd.n2950 gnd.n2248 225.874
R7340 gnd.n2950 gnd.n2949 225.874
R7341 gnd.n2949 gnd.n2948 225.874
R7342 gnd.n2948 gnd.n2256 225.874
R7343 gnd.n2942 gnd.n2256 225.874
R7344 gnd.n2942 gnd.n2941 225.874
R7345 gnd.n2941 gnd.n2940 225.874
R7346 gnd.n2940 gnd.n2264 225.874
R7347 gnd.n2934 gnd.n2264 225.874
R7348 gnd.n2934 gnd.n2933 225.874
R7349 gnd.n2933 gnd.n2932 225.874
R7350 gnd.n2932 gnd.n2272 225.874
R7351 gnd.n2926 gnd.n2272 225.874
R7352 gnd.n2926 gnd.n2925 225.874
R7353 gnd.n2925 gnd.n2924 225.874
R7354 gnd.n2924 gnd.n2280 225.874
R7355 gnd.n2918 gnd.n2280 225.874
R7356 gnd.n2918 gnd.n2917 225.874
R7357 gnd.n2917 gnd.n2916 225.874
R7358 gnd.n2916 gnd.n2288 225.874
R7359 gnd.n2910 gnd.n2288 225.874
R7360 gnd.n2910 gnd.n2909 225.874
R7361 gnd.n2909 gnd.n2908 225.874
R7362 gnd.n2908 gnd.n2296 225.874
R7363 gnd.n2902 gnd.n2296 225.874
R7364 gnd.n2902 gnd.n2901 225.874
R7365 gnd.n2901 gnd.n2900 225.874
R7366 gnd.n2900 gnd.n2304 225.874
R7367 gnd.n2894 gnd.n2304 225.874
R7368 gnd.n2894 gnd.n2893 225.874
R7369 gnd.n2893 gnd.n2892 225.874
R7370 gnd.n2892 gnd.n2312 225.874
R7371 gnd.n2886 gnd.n2312 225.874
R7372 gnd.n2886 gnd.n2885 225.874
R7373 gnd.n2885 gnd.n2884 225.874
R7374 gnd.n2884 gnd.n2320 225.874
R7375 gnd.n2878 gnd.n2320 225.874
R7376 gnd.n2878 gnd.n2877 225.874
R7377 gnd.n2877 gnd.n2876 225.874
R7378 gnd.n2876 gnd.n2328 225.874
R7379 gnd.n2870 gnd.n2328 225.874
R7380 gnd.n2870 gnd.n2869 225.874
R7381 gnd.n2869 gnd.n2868 225.874
R7382 gnd.n2868 gnd.n2336 225.874
R7383 gnd.n2862 gnd.n2336 225.874
R7384 gnd.n2862 gnd.n2861 225.874
R7385 gnd.n2861 gnd.n2860 225.874
R7386 gnd.n2860 gnd.n2344 225.874
R7387 gnd.n2854 gnd.n2344 225.874
R7388 gnd.n2854 gnd.n2853 225.874
R7389 gnd.n2853 gnd.n2852 225.874
R7390 gnd.n2852 gnd.n2352 225.874
R7391 gnd.n2846 gnd.n2352 225.874
R7392 gnd.n2846 gnd.n2845 225.874
R7393 gnd.n2845 gnd.n2844 225.874
R7394 gnd.n2844 gnd.n2360 225.874
R7395 gnd.n2838 gnd.n2360 225.874
R7396 gnd.n2838 gnd.n2837 225.874
R7397 gnd.n2837 gnd.n2836 225.874
R7398 gnd.n2836 gnd.n2368 225.874
R7399 gnd.n2830 gnd.n2368 225.874
R7400 gnd.n2830 gnd.n2829 225.874
R7401 gnd.n2829 gnd.n2828 225.874
R7402 gnd.n2828 gnd.n2376 225.874
R7403 gnd.n2822 gnd.n2376 225.874
R7404 gnd.n2822 gnd.n2821 225.874
R7405 gnd.n2821 gnd.n2820 225.874
R7406 gnd.n2820 gnd.n2384 225.874
R7407 gnd.n2814 gnd.n2384 225.874
R7408 gnd.n2814 gnd.n2813 225.874
R7409 gnd.n2813 gnd.n2812 225.874
R7410 gnd.n2812 gnd.n2392 225.874
R7411 gnd.n2806 gnd.n2392 225.874
R7412 gnd.n2806 gnd.n2805 225.874
R7413 gnd.n2805 gnd.n2804 225.874
R7414 gnd.n2804 gnd.n2400 225.874
R7415 gnd.n2798 gnd.n2400 225.874
R7416 gnd.n2798 gnd.n2797 225.874
R7417 gnd.n2797 gnd.n2796 225.874
R7418 gnd.n2796 gnd.n2408 225.874
R7419 gnd.n2790 gnd.n2408 225.874
R7420 gnd.n2790 gnd.n2789 225.874
R7421 gnd.n2789 gnd.n2788 225.874
R7422 gnd.n2788 gnd.n2416 225.874
R7423 gnd.n2782 gnd.n2416 225.874
R7424 gnd.n2782 gnd.n2781 225.874
R7425 gnd.n2781 gnd.n2780 225.874
R7426 gnd.n2780 gnd.n2424 225.874
R7427 gnd.n2774 gnd.n2424 225.874
R7428 gnd.n2774 gnd.n2773 225.874
R7429 gnd.n3819 gnd.t17 224.174
R7430 gnd.n1884 gnd.t128 224.174
R7431 gnd.n658 gnd.n601 199.319
R7432 gnd.n658 gnd.n602 199.319
R7433 gnd.n5915 gnd.n1363 199.319
R7434 gnd.n1368 gnd.n1363 199.319
R7435 gnd.n1273 gnd.n1270 186.49
R7436 gnd.n6564 gnd.n6561 186.49
R7437 gnd.n4594 gnd.n4593 185
R7438 gnd.n4592 gnd.n4591 185
R7439 gnd.n4571 gnd.n4570 185
R7440 gnd.n4586 gnd.n4585 185
R7441 gnd.n4584 gnd.n4583 185
R7442 gnd.n4575 gnd.n4574 185
R7443 gnd.n4578 gnd.n4577 185
R7444 gnd.n4562 gnd.n4561 185
R7445 gnd.n4560 gnd.n4559 185
R7446 gnd.n4539 gnd.n4538 185
R7447 gnd.n4554 gnd.n4553 185
R7448 gnd.n4552 gnd.n4551 185
R7449 gnd.n4543 gnd.n4542 185
R7450 gnd.n4546 gnd.n4545 185
R7451 gnd.n4530 gnd.n4529 185
R7452 gnd.n4528 gnd.n4527 185
R7453 gnd.n4507 gnd.n4506 185
R7454 gnd.n4522 gnd.n4521 185
R7455 gnd.n4520 gnd.n4519 185
R7456 gnd.n4511 gnd.n4510 185
R7457 gnd.n4514 gnd.n4513 185
R7458 gnd.n4499 gnd.n4498 185
R7459 gnd.n4497 gnd.n4496 185
R7460 gnd.n4476 gnd.n4475 185
R7461 gnd.n4491 gnd.n4490 185
R7462 gnd.n4489 gnd.n4488 185
R7463 gnd.n4480 gnd.n4479 185
R7464 gnd.n4483 gnd.n4482 185
R7465 gnd.n4467 gnd.n4466 185
R7466 gnd.n4465 gnd.n4464 185
R7467 gnd.n4444 gnd.n4443 185
R7468 gnd.n4459 gnd.n4458 185
R7469 gnd.n4457 gnd.n4456 185
R7470 gnd.n4448 gnd.n4447 185
R7471 gnd.n4451 gnd.n4450 185
R7472 gnd.n4435 gnd.n4434 185
R7473 gnd.n4433 gnd.n4432 185
R7474 gnd.n4412 gnd.n4411 185
R7475 gnd.n4427 gnd.n4426 185
R7476 gnd.n4425 gnd.n4424 185
R7477 gnd.n4416 gnd.n4415 185
R7478 gnd.n4419 gnd.n4418 185
R7479 gnd.n4403 gnd.n4402 185
R7480 gnd.n4401 gnd.n4400 185
R7481 gnd.n4380 gnd.n4379 185
R7482 gnd.n4395 gnd.n4394 185
R7483 gnd.n4393 gnd.n4392 185
R7484 gnd.n4384 gnd.n4383 185
R7485 gnd.n4387 gnd.n4386 185
R7486 gnd.n4372 gnd.n4371 185
R7487 gnd.n4370 gnd.n4369 185
R7488 gnd.n4349 gnd.n4348 185
R7489 gnd.n4364 gnd.n4363 185
R7490 gnd.n4362 gnd.n4361 185
R7491 gnd.n4353 gnd.n4352 185
R7492 gnd.n4356 gnd.n4355 185
R7493 gnd.n3820 gnd.t16 178.987
R7494 gnd.n1885 gnd.t129 178.987
R7495 gnd.n1 gnd.t390 170.774
R7496 gnd.n7 gnd.t398 170.103
R7497 gnd.n6 gnd.t392 170.103
R7498 gnd.n5 gnd.t148 170.103
R7499 gnd.n4 gnd.t396 170.103
R7500 gnd.n3 gnd.t150 170.103
R7501 gnd.n2 gnd.t138 170.103
R7502 gnd.n1 gnd.t132 170.103
R7503 gnd.n6635 gnd.n6634 163.367
R7504 gnd.n6631 gnd.n6630 163.367
R7505 gnd.n6627 gnd.n6626 163.367
R7506 gnd.n6623 gnd.n6622 163.367
R7507 gnd.n6619 gnd.n6618 163.367
R7508 gnd.n6615 gnd.n6614 163.367
R7509 gnd.n6611 gnd.n6610 163.367
R7510 gnd.n6607 gnd.n6606 163.367
R7511 gnd.n6603 gnd.n6602 163.367
R7512 gnd.n6599 gnd.n6598 163.367
R7513 gnd.n6595 gnd.n6594 163.367
R7514 gnd.n6591 gnd.n6590 163.367
R7515 gnd.n6587 gnd.n6586 163.367
R7516 gnd.n6583 gnd.n6582 163.367
R7517 gnd.n6578 gnd.n6577 163.367
R7518 gnd.n6574 gnd.n6573 163.367
R7519 gnd.n6711 gnd.n6710 163.367
R7520 gnd.n6707 gnd.n6706 163.367
R7521 gnd.n6702 gnd.n6701 163.367
R7522 gnd.n6698 gnd.n6697 163.367
R7523 gnd.n6694 gnd.n6693 163.367
R7524 gnd.n6690 gnd.n6689 163.367
R7525 gnd.n6686 gnd.n6685 163.367
R7526 gnd.n6682 gnd.n6681 163.367
R7527 gnd.n6678 gnd.n6677 163.367
R7528 gnd.n6674 gnd.n6673 163.367
R7529 gnd.n6670 gnd.n6669 163.367
R7530 gnd.n6666 gnd.n6665 163.367
R7531 gnd.n6662 gnd.n6661 163.367
R7532 gnd.n6658 gnd.n6657 163.367
R7533 gnd.n6654 gnd.n6653 163.367
R7534 gnd.n6650 gnd.n6649 163.367
R7535 gnd.n1296 gnd.n1202 163.367
R7536 gnd.n6153 gnd.n1202 163.367
R7537 gnd.n6153 gnd.n1192 163.367
R7538 gnd.n1194 gnd.n1192 163.367
R7539 gnd.n1194 gnd.n1184 163.367
R7540 gnd.n6147 gnd.n1184 163.367
R7541 gnd.n6147 gnd.n1212 163.367
R7542 gnd.n1212 gnd.n1211 163.367
R7543 gnd.n1211 gnd.n1207 163.367
R7544 gnd.n1207 gnd.n1165 163.367
R7545 gnd.n1165 gnd.n1155 163.367
R7546 gnd.n6216 gnd.n1155 163.367
R7547 gnd.n6216 gnd.n1153 163.367
R7548 gnd.n6220 gnd.n1153 163.367
R7549 gnd.n6220 gnd.n1142 163.367
R7550 gnd.n6239 gnd.n1142 163.367
R7551 gnd.n6239 gnd.n1137 163.367
R7552 gnd.n6235 gnd.n1137 163.367
R7553 gnd.n6235 gnd.n1127 163.367
R7554 gnd.n6262 gnd.n1127 163.367
R7555 gnd.n6262 gnd.n1115 163.367
R7556 gnd.n6265 gnd.n1115 163.367
R7557 gnd.n6265 gnd.n1108 163.367
R7558 gnd.n6277 gnd.n1108 163.367
R7559 gnd.n6277 gnd.n1125 163.367
R7560 gnd.n6273 gnd.n1125 163.367
R7561 gnd.n6273 gnd.n1084 163.367
R7562 gnd.n6270 gnd.n1084 163.367
R7563 gnd.n6270 gnd.n1078 163.367
R7564 gnd.n1093 gnd.n1078 163.367
R7565 gnd.n1093 gnd.n1068 163.367
R7566 gnd.n6371 gnd.n1068 163.367
R7567 gnd.n6371 gnd.n1058 163.367
R7568 gnd.n6374 gnd.n1058 163.367
R7569 gnd.n6374 gnd.n1051 163.367
R7570 gnd.n6378 gnd.n1051 163.367
R7571 gnd.n6378 gnd.n1041 163.367
R7572 gnd.n6408 gnd.n1041 163.367
R7573 gnd.n6408 gnd.n1027 163.367
R7574 gnd.n6411 gnd.n1027 163.367
R7575 gnd.n6411 gnd.n1021 163.367
R7576 gnd.n6417 gnd.n1021 163.367
R7577 gnd.n6417 gnd.n1011 163.367
R7578 gnd.n1011 gnd.n1004 163.367
R7579 gnd.n6450 gnd.n1004 163.367
R7580 gnd.n6451 gnd.n6450 163.367
R7581 gnd.n6451 gnd.n1002 163.367
R7582 gnd.n6455 gnd.n1002 163.367
R7583 gnd.n6455 gnd.n994 163.367
R7584 gnd.n6465 gnd.n994 163.367
R7585 gnd.n6465 gnd.n992 163.367
R7586 gnd.n6479 gnd.n992 163.367
R7587 gnd.n6479 gnd.n953 163.367
R7588 gnd.n6475 gnd.n953 163.367
R7589 gnd.n6475 gnd.n946 163.367
R7590 gnd.n6472 gnd.n946 163.367
R7591 gnd.n6472 gnd.n939 163.367
R7592 gnd.n939 gnd.n930 163.367
R7593 gnd.n6644 gnd.n930 163.367
R7594 gnd.n6645 gnd.n6644 163.367
R7595 gnd.n1264 gnd.n1263 163.367
R7596 gnd.n6092 gnd.n1263 163.367
R7597 gnd.n6090 gnd.n6089 163.367
R7598 gnd.n6086 gnd.n6085 163.367
R7599 gnd.n6082 gnd.n6081 163.367
R7600 gnd.n6078 gnd.n6077 163.367
R7601 gnd.n6074 gnd.n6073 163.367
R7602 gnd.n6070 gnd.n6069 163.367
R7603 gnd.n6066 gnd.n6065 163.367
R7604 gnd.n6062 gnd.n6061 163.367
R7605 gnd.n6058 gnd.n6057 163.367
R7606 gnd.n6054 gnd.n6053 163.367
R7607 gnd.n6050 gnd.n6049 163.367
R7608 gnd.n6046 gnd.n6045 163.367
R7609 gnd.n6042 gnd.n6041 163.367
R7610 gnd.n6038 gnd.n6037 163.367
R7611 gnd.n6034 gnd.n6033 163.367
R7612 gnd.n1358 gnd.n1357 163.367
R7613 gnd.n1353 gnd.n1352 163.367
R7614 gnd.n1349 gnd.n1348 163.367
R7615 gnd.n1345 gnd.n1344 163.367
R7616 gnd.n1341 gnd.n1340 163.367
R7617 gnd.n1337 gnd.n1336 163.367
R7618 gnd.n1333 gnd.n1332 163.367
R7619 gnd.n1329 gnd.n1328 163.367
R7620 gnd.n1325 gnd.n1324 163.367
R7621 gnd.n1321 gnd.n1320 163.367
R7622 gnd.n1317 gnd.n1316 163.367
R7623 gnd.n1313 gnd.n1312 163.367
R7624 gnd.n1309 gnd.n1308 163.367
R7625 gnd.n1305 gnd.n1304 163.367
R7626 gnd.n1301 gnd.n1300 163.367
R7627 gnd.n1286 gnd.n1265 163.367
R7628 gnd.n1286 gnd.n1190 163.367
R7629 gnd.n6166 gnd.n1190 163.367
R7630 gnd.n6166 gnd.n1187 163.367
R7631 gnd.n6175 gnd.n1187 163.367
R7632 gnd.n6175 gnd.n1188 163.367
R7633 gnd.n6171 gnd.n1188 163.367
R7634 gnd.n6171 gnd.n6170 163.367
R7635 gnd.n6170 gnd.n1163 163.367
R7636 gnd.n6209 gnd.n1163 163.367
R7637 gnd.n6209 gnd.n1158 163.367
R7638 gnd.n6214 gnd.n1158 163.367
R7639 gnd.n6214 gnd.n1161 163.367
R7640 gnd.n1161 gnd.n1141 163.367
R7641 gnd.n6243 gnd.n1141 163.367
R7642 gnd.n6243 gnd.n1138 163.367
R7643 gnd.n6250 gnd.n1138 163.367
R7644 gnd.n6250 gnd.n1139 163.367
R7645 gnd.n6246 gnd.n1139 163.367
R7646 gnd.n6246 gnd.n1113 163.367
R7647 gnd.n6289 gnd.n1113 163.367
R7648 gnd.n6289 gnd.n1110 163.367
R7649 gnd.n6296 gnd.n1110 163.367
R7650 gnd.n6296 gnd.n1111 163.367
R7651 gnd.n6292 gnd.n1111 163.367
R7652 gnd.n6292 gnd.n1083 163.367
R7653 gnd.n6351 gnd.n1083 163.367
R7654 gnd.n6351 gnd.n1080 163.367
R7655 gnd.n6358 gnd.n1080 163.367
R7656 gnd.n6358 gnd.n1081 163.367
R7657 gnd.n6354 gnd.n1081 163.367
R7658 gnd.n6354 gnd.n1056 163.367
R7659 gnd.n6388 gnd.n1056 163.367
R7660 gnd.n6388 gnd.n1053 163.367
R7661 gnd.n6395 gnd.n1053 163.367
R7662 gnd.n6395 gnd.n1054 163.367
R7663 gnd.n6391 gnd.n1054 163.367
R7664 gnd.n6391 gnd.n1025 163.367
R7665 gnd.n6427 gnd.n1025 163.367
R7666 gnd.n6427 gnd.n1023 163.367
R7667 gnd.n6431 gnd.n1023 163.367
R7668 gnd.n6431 gnd.n1010 163.367
R7669 gnd.n6443 gnd.n1010 163.367
R7670 gnd.n6443 gnd.n1007 163.367
R7671 gnd.n6448 gnd.n1007 163.367
R7672 gnd.n6448 gnd.n1008 163.367
R7673 gnd.n1008 gnd.n999 163.367
R7674 gnd.n6458 gnd.n999 163.367
R7675 gnd.n6458 gnd.n996 163.367
R7676 gnd.n6463 gnd.n996 163.367
R7677 gnd.n6463 gnd.n997 163.367
R7678 gnd.n997 gnd.n951 163.367
R7679 gnd.n6533 gnd.n951 163.367
R7680 gnd.n6533 gnd.n949 163.367
R7681 gnd.n6537 gnd.n949 163.367
R7682 gnd.n6537 gnd.n937 163.367
R7683 gnd.n6549 gnd.n937 163.367
R7684 gnd.n6549 gnd.n934 163.367
R7685 gnd.n6642 gnd.n934 163.367
R7686 gnd.n6642 gnd.n935 163.367
R7687 gnd.n6570 gnd.n6569 156.462
R7688 gnd.n6989 gnd.n657 154.689
R7689 gnd.n6035 gnd.n6031 154.689
R7690 gnd.n4534 gnd.n4502 153.042
R7691 gnd.n4598 gnd.n4597 152.079
R7692 gnd.n4566 gnd.n4565 152.079
R7693 gnd.n4534 gnd.n4533 152.079
R7694 gnd.n1278 gnd.n1277 152
R7695 gnd.n1279 gnd.n1268 152
R7696 gnd.n1281 gnd.n1280 152
R7697 gnd.n1283 gnd.n1266 152
R7698 gnd.n1285 gnd.n1284 152
R7699 gnd.n6568 gnd.n6552 152
R7700 gnd.n6560 gnd.n6553 152
R7701 gnd.n6559 gnd.n6558 152
R7702 gnd.n6557 gnd.n6554 152
R7703 gnd.n6555 gnd.t61 150.546
R7704 gnd.t152 gnd.n4576 147.661
R7705 gnd.t158 gnd.n4544 147.661
R7706 gnd.t386 gnd.n4512 147.661
R7707 gnd.t154 gnd.n4481 147.661
R7708 gnd.t394 gnd.n4449 147.661
R7709 gnd.t134 gnd.n4417 147.661
R7710 gnd.t167 gnd.n4385 147.661
R7711 gnd.t161 gnd.n4354 147.661
R7712 gnd.n926 gnd.n909 143.351
R7713 gnd.n6032 gnd.n1242 143.351
R7714 gnd.n6032 gnd.n1243 143.351
R7715 gnd.n1275 gnd.t114 130.484
R7716 gnd.n1284 gnd.t104 126.766
R7717 gnd.n1282 gnd.t86 126.766
R7718 gnd.n1268 gnd.t22 126.766
R7719 gnd.n1276 gnd.t70 126.766
R7720 gnd.n6556 gnd.t11 126.766
R7721 gnd.n6558 gnd.t79 126.766
R7722 gnd.n6567 gnd.t101 126.766
R7723 gnd.n6569 gnd.t55 126.766
R7724 gnd.n4593 gnd.n4592 104.615
R7725 gnd.n4592 gnd.n4570 104.615
R7726 gnd.n4585 gnd.n4570 104.615
R7727 gnd.n4585 gnd.n4584 104.615
R7728 gnd.n4584 gnd.n4574 104.615
R7729 gnd.n4577 gnd.n4574 104.615
R7730 gnd.n4561 gnd.n4560 104.615
R7731 gnd.n4560 gnd.n4538 104.615
R7732 gnd.n4553 gnd.n4538 104.615
R7733 gnd.n4553 gnd.n4552 104.615
R7734 gnd.n4552 gnd.n4542 104.615
R7735 gnd.n4545 gnd.n4542 104.615
R7736 gnd.n4529 gnd.n4528 104.615
R7737 gnd.n4528 gnd.n4506 104.615
R7738 gnd.n4521 gnd.n4506 104.615
R7739 gnd.n4521 gnd.n4520 104.615
R7740 gnd.n4520 gnd.n4510 104.615
R7741 gnd.n4513 gnd.n4510 104.615
R7742 gnd.n4498 gnd.n4497 104.615
R7743 gnd.n4497 gnd.n4475 104.615
R7744 gnd.n4490 gnd.n4475 104.615
R7745 gnd.n4490 gnd.n4489 104.615
R7746 gnd.n4489 gnd.n4479 104.615
R7747 gnd.n4482 gnd.n4479 104.615
R7748 gnd.n4466 gnd.n4465 104.615
R7749 gnd.n4465 gnd.n4443 104.615
R7750 gnd.n4458 gnd.n4443 104.615
R7751 gnd.n4458 gnd.n4457 104.615
R7752 gnd.n4457 gnd.n4447 104.615
R7753 gnd.n4450 gnd.n4447 104.615
R7754 gnd.n4434 gnd.n4433 104.615
R7755 gnd.n4433 gnd.n4411 104.615
R7756 gnd.n4426 gnd.n4411 104.615
R7757 gnd.n4426 gnd.n4425 104.615
R7758 gnd.n4425 gnd.n4415 104.615
R7759 gnd.n4418 gnd.n4415 104.615
R7760 gnd.n4402 gnd.n4401 104.615
R7761 gnd.n4401 gnd.n4379 104.615
R7762 gnd.n4394 gnd.n4379 104.615
R7763 gnd.n4394 gnd.n4393 104.615
R7764 gnd.n4393 gnd.n4383 104.615
R7765 gnd.n4386 gnd.n4383 104.615
R7766 gnd.n4371 gnd.n4370 104.615
R7767 gnd.n4370 gnd.n4348 104.615
R7768 gnd.n4363 gnd.n4348 104.615
R7769 gnd.n4363 gnd.n4362 104.615
R7770 gnd.n4362 gnd.n4352 104.615
R7771 gnd.n4355 gnd.n4352 104.615
R7772 gnd.n2772 gnd.n2432 103.311
R7773 gnd.n2441 gnd.n2432 103.311
R7774 gnd.n2763 gnd.n2441 103.311
R7775 gnd.n2763 gnd.n2762 103.311
R7776 gnd.n2762 gnd.n2761 103.311
R7777 gnd.n2761 gnd.n2442 103.311
R7778 gnd.n2755 gnd.n2442 103.311
R7779 gnd.n2755 gnd.n2754 103.311
R7780 gnd.n2754 gnd.n2753 103.311
R7781 gnd.n2753 gnd.n2449 103.311
R7782 gnd.n2747 gnd.n2449 103.311
R7783 gnd.n2747 gnd.n2746 103.311
R7784 gnd.n2746 gnd.n2745 103.311
R7785 gnd.n2745 gnd.n2457 103.311
R7786 gnd.n2739 gnd.n2457 103.311
R7787 gnd.n2739 gnd.n2738 103.311
R7788 gnd.n2738 gnd.n2737 103.311
R7789 gnd.n2737 gnd.n2465 103.311
R7790 gnd.n2731 gnd.n2465 103.311
R7791 gnd.n2731 gnd.n2730 103.311
R7792 gnd.n2730 gnd.n2729 103.311
R7793 gnd.n2729 gnd.n2473 103.311
R7794 gnd.n2723 gnd.n2473 103.311
R7795 gnd.n2723 gnd.n2722 103.311
R7796 gnd.n2722 gnd.n2721 103.311
R7797 gnd.n2721 gnd.n2481 103.311
R7798 gnd.n2715 gnd.n2481 103.311
R7799 gnd.n2715 gnd.n2714 103.311
R7800 gnd.n2714 gnd.n2713 103.311
R7801 gnd.n2713 gnd.n2489 103.311
R7802 gnd.n2707 gnd.n2489 103.311
R7803 gnd.n2707 gnd.n2706 103.311
R7804 gnd.n2706 gnd.n2705 103.311
R7805 gnd.n2705 gnd.n2497 103.311
R7806 gnd.n2699 gnd.n2497 103.311
R7807 gnd.n2699 gnd.n2698 103.311
R7808 gnd.n2698 gnd.n2697 103.311
R7809 gnd.n2697 gnd.n2505 103.311
R7810 gnd.n2691 gnd.n2505 103.311
R7811 gnd.n2691 gnd.n2690 103.311
R7812 gnd.n2690 gnd.n2689 103.311
R7813 gnd.n2689 gnd.n2513 103.311
R7814 gnd.n2683 gnd.n2513 103.311
R7815 gnd.n2683 gnd.n2682 103.311
R7816 gnd.n2682 gnd.n2681 103.311
R7817 gnd.n2681 gnd.n2521 103.311
R7818 gnd.n2675 gnd.n2521 103.311
R7819 gnd.n2675 gnd.n2674 103.311
R7820 gnd.n2674 gnd.n2673 103.311
R7821 gnd.n2673 gnd.n2529 103.311
R7822 gnd.n2667 gnd.n2529 103.311
R7823 gnd.n2667 gnd.n2666 103.311
R7824 gnd.n2666 gnd.n2665 103.311
R7825 gnd.n2665 gnd.n2537 103.311
R7826 gnd.n2659 gnd.n2537 103.311
R7827 gnd.n2659 gnd.n2658 103.311
R7828 gnd.n2658 gnd.n2657 103.311
R7829 gnd.n2657 gnd.n2545 103.311
R7830 gnd.n2651 gnd.n2545 103.311
R7831 gnd.n2651 gnd.n2650 103.311
R7832 gnd.n2650 gnd.n2649 103.311
R7833 gnd.n2649 gnd.n2553 103.311
R7834 gnd.n2643 gnd.n2553 103.311
R7835 gnd.n2643 gnd.n2642 103.311
R7836 gnd.n2642 gnd.n2641 103.311
R7837 gnd.n2641 gnd.n2561 103.311
R7838 gnd.n2635 gnd.n2561 103.311
R7839 gnd.n2635 gnd.n2634 103.311
R7840 gnd.n2634 gnd.n2633 103.311
R7841 gnd.n2633 gnd.n2569 103.311
R7842 gnd.n2627 gnd.n2569 103.311
R7843 gnd.n2627 gnd.n2626 103.311
R7844 gnd.n2626 gnd.n2625 103.311
R7845 gnd.n2625 gnd.n2577 103.311
R7846 gnd.n2619 gnd.n2577 103.311
R7847 gnd.n2619 gnd.n2618 103.311
R7848 gnd.n2618 gnd.n2617 103.311
R7849 gnd.n2617 gnd.n2585 103.311
R7850 gnd.n2611 gnd.n2585 103.311
R7851 gnd.n2611 gnd.n2610 103.311
R7852 gnd.n2610 gnd.n2609 103.311
R7853 gnd.n2609 gnd.n2593 103.311
R7854 gnd.n2603 gnd.n2593 103.311
R7855 gnd.n3745 gnd.t85 100.632
R7856 gnd.n1858 gnd.t109 100.632
R7857 gnd.n7659 gnd.n7658 99.6594
R7858 gnd.n7654 gnd.n288 99.6594
R7859 gnd.n7650 gnd.n287 99.6594
R7860 gnd.n7646 gnd.n286 99.6594
R7861 gnd.n7642 gnd.n285 99.6594
R7862 gnd.n7638 gnd.n284 99.6594
R7863 gnd.n7634 gnd.n283 99.6594
R7864 gnd.n7630 gnd.n282 99.6594
R7865 gnd.n7623 gnd.n281 99.6594
R7866 gnd.n7619 gnd.n280 99.6594
R7867 gnd.n7615 gnd.n279 99.6594
R7868 gnd.n7611 gnd.n278 99.6594
R7869 gnd.n7607 gnd.n277 99.6594
R7870 gnd.n7603 gnd.n276 99.6594
R7871 gnd.n7599 gnd.n275 99.6594
R7872 gnd.n7595 gnd.n274 99.6594
R7873 gnd.n7591 gnd.n273 99.6594
R7874 gnd.n7587 gnd.n272 99.6594
R7875 gnd.n7579 gnd.n271 99.6594
R7876 gnd.n7577 gnd.n270 99.6594
R7877 gnd.n7573 gnd.n269 99.6594
R7878 gnd.n7569 gnd.n268 99.6594
R7879 gnd.n7565 gnd.n267 99.6594
R7880 gnd.n7561 gnd.n266 99.6594
R7881 gnd.n7557 gnd.n265 99.6594
R7882 gnd.n7553 gnd.n264 99.6594
R7883 gnd.n7549 gnd.n263 99.6594
R7884 gnd.n7545 gnd.n262 99.6594
R7885 gnd.n7536 gnd.n261 99.6594
R7886 gnd.n7040 gnd.n568 99.6594
R7887 gnd.n7035 gnd.n590 99.6594
R7888 gnd.n7032 gnd.n591 99.6594
R7889 gnd.n7028 gnd.n592 99.6594
R7890 gnd.n7024 gnd.n593 99.6594
R7891 gnd.n7020 gnd.n594 99.6594
R7892 gnd.n7016 gnd.n595 99.6594
R7893 gnd.n7012 gnd.n596 99.6594
R7894 gnd.n7008 gnd.n597 99.6594
R7895 gnd.n7003 gnd.n598 99.6594
R7896 gnd.n6999 gnd.n599 99.6594
R7897 gnd.n6995 gnd.n600 99.6594
R7898 gnd.n6991 gnd.n601 99.6594
R7899 gnd.n6986 gnd.n603 99.6594
R7900 gnd.n6982 gnd.n604 99.6594
R7901 gnd.n6978 gnd.n605 99.6594
R7902 gnd.n6974 gnd.n606 99.6594
R7903 gnd.n6970 gnd.n607 99.6594
R7904 gnd.n6966 gnd.n608 99.6594
R7905 gnd.n6962 gnd.n609 99.6594
R7906 gnd.n6958 gnd.n610 99.6594
R7907 gnd.n6954 gnd.n611 99.6594
R7908 gnd.n6950 gnd.n612 99.6594
R7909 gnd.n6946 gnd.n613 99.6594
R7910 gnd.n6942 gnd.n614 99.6594
R7911 gnd.n6938 gnd.n615 99.6594
R7912 gnd.n6934 gnd.n616 99.6594
R7913 gnd.n6930 gnd.n617 99.6594
R7914 gnd.n5957 gnd.n5956 99.6594
R7915 gnd.n5952 gnd.n5877 99.6594
R7916 gnd.n5950 gnd.n5949 99.6594
R7917 gnd.n5945 gnd.n5884 99.6594
R7918 gnd.n5943 gnd.n5942 99.6594
R7919 gnd.n5938 gnd.n5891 99.6594
R7920 gnd.n5936 gnd.n5935 99.6594
R7921 gnd.n5931 gnd.n5898 99.6594
R7922 gnd.n5929 gnd.n5928 99.6594
R7923 gnd.n5924 gnd.n5908 99.6594
R7924 gnd.n5922 gnd.n5921 99.6594
R7925 gnd.n5917 gnd.n5914 99.6594
R7926 gnd.n1368 gnd.n1367 99.6594
R7927 gnd.n6025 gnd.n6024 99.6594
R7928 gnd.n6022 gnd.n6021 99.6594
R7929 gnd.n6017 gnd.n1377 99.6594
R7930 gnd.n6015 gnd.n6014 99.6594
R7931 gnd.n1387 gnd.n1386 99.6594
R7932 gnd.n6006 gnd.n6005 99.6594
R7933 gnd.n6003 gnd.n6002 99.6594
R7934 gnd.n5998 gnd.n1395 99.6594
R7935 gnd.n5996 gnd.n5995 99.6594
R7936 gnd.n5991 gnd.n1402 99.6594
R7937 gnd.n5989 gnd.n5988 99.6594
R7938 gnd.n5984 gnd.n1409 99.6594
R7939 gnd.n5982 gnd.n5981 99.6594
R7940 gnd.n5977 gnd.n1418 99.6594
R7941 gnd.n5975 gnd.n5974 99.6594
R7942 gnd.n4885 gnd.n1818 99.6594
R7943 gnd.n4893 gnd.n4892 99.6594
R7944 gnd.n4896 gnd.n4895 99.6594
R7945 gnd.n4903 gnd.n4902 99.6594
R7946 gnd.n4906 gnd.n4905 99.6594
R7947 gnd.n4913 gnd.n4912 99.6594
R7948 gnd.n4916 gnd.n4915 99.6594
R7949 gnd.n4923 gnd.n4922 99.6594
R7950 gnd.n4926 gnd.n4925 99.6594
R7951 gnd.n4933 gnd.n4932 99.6594
R7952 gnd.n4936 gnd.n4935 99.6594
R7953 gnd.n4943 gnd.n4942 99.6594
R7954 gnd.n4946 gnd.n4945 99.6594
R7955 gnd.n4953 gnd.n4952 99.6594
R7956 gnd.n4956 gnd.n4955 99.6594
R7957 gnd.n4963 gnd.n4962 99.6594
R7958 gnd.n4966 gnd.n4965 99.6594
R7959 gnd.n4973 gnd.n4972 99.6594
R7960 gnd.n4976 gnd.n4975 99.6594
R7961 gnd.n4985 gnd.n4984 99.6594
R7962 gnd.n4988 gnd.n4987 99.6594
R7963 gnd.n4995 gnd.n4994 99.6594
R7964 gnd.n4998 gnd.n4997 99.6594
R7965 gnd.n5005 gnd.n5004 99.6594
R7966 gnd.n5008 gnd.n5007 99.6594
R7967 gnd.n5015 gnd.n5014 99.6594
R7968 gnd.n5018 gnd.n5017 99.6594
R7969 gnd.n5026 gnd.n5025 99.6594
R7970 gnd.n5029 gnd.n5028 99.6594
R7971 gnd.n4717 gnd.n1841 99.6594
R7972 gnd.n4715 gnd.n1840 99.6594
R7973 gnd.n4711 gnd.n1839 99.6594
R7974 gnd.n4707 gnd.n1838 99.6594
R7975 gnd.n4703 gnd.n1837 99.6594
R7976 gnd.n4699 gnd.n1836 99.6594
R7977 gnd.n4695 gnd.n1835 99.6594
R7978 gnd.n4627 gnd.n1834 99.6594
R7979 gnd.n3957 gnd.n3688 99.6594
R7980 gnd.n3714 gnd.n3695 99.6594
R7981 gnd.n3716 gnd.n3696 99.6594
R7982 gnd.n3724 gnd.n3697 99.6594
R7983 gnd.n3726 gnd.n3698 99.6594
R7984 gnd.n3734 gnd.n3699 99.6594
R7985 gnd.n3736 gnd.n3700 99.6594
R7986 gnd.n3744 gnd.n3701 99.6594
R7987 gnd.n7408 gnd.n252 99.6594
R7988 gnd.n7412 gnd.n253 99.6594
R7989 gnd.n7418 gnd.n254 99.6594
R7990 gnd.n7422 gnd.n255 99.6594
R7991 gnd.n7428 gnd.n256 99.6594
R7992 gnd.n7432 gnd.n257 99.6594
R7993 gnd.n7438 gnd.n258 99.6594
R7994 gnd.n7442 gnd.n259 99.6594
R7995 gnd.n7448 gnd.n260 99.6594
R7996 gnd.n618 gnd.n573 99.6594
R7997 gnd.n706 gnd.n619 99.6594
R7998 gnd.n714 gnd.n620 99.6594
R7999 gnd.n716 gnd.n621 99.6594
R8000 gnd.n724 gnd.n622 99.6594
R8001 gnd.n732 gnd.n623 99.6594
R8002 gnd.n734 gnd.n624 99.6594
R8003 gnd.n742 gnd.n625 99.6594
R8004 gnd.n752 gnd.n626 99.6594
R8005 gnd.n4685 gnd.n1821 99.6594
R8006 gnd.n4681 gnd.n1822 99.6594
R8007 gnd.n4677 gnd.n1823 99.6594
R8008 gnd.n4673 gnd.n1824 99.6594
R8009 gnd.n4669 gnd.n1825 99.6594
R8010 gnd.n4665 gnd.n1826 99.6594
R8011 gnd.n4661 gnd.n1827 99.6594
R8012 gnd.n4657 gnd.n1828 99.6594
R8013 gnd.n4653 gnd.n1829 99.6594
R8014 gnd.n4649 gnd.n1830 99.6594
R8015 gnd.n4645 gnd.n1831 99.6594
R8016 gnd.n4641 gnd.n1832 99.6594
R8017 gnd.n4637 gnd.n1833 99.6594
R8018 gnd.n3872 gnd.n3871 99.6594
R8019 gnd.n3866 gnd.n3783 99.6594
R8020 gnd.n3863 gnd.n3784 99.6594
R8021 gnd.n3859 gnd.n3785 99.6594
R8022 gnd.n3855 gnd.n3786 99.6594
R8023 gnd.n3851 gnd.n3787 99.6594
R8024 gnd.n3847 gnd.n3788 99.6594
R8025 gnd.n3843 gnd.n3789 99.6594
R8026 gnd.n3839 gnd.n3790 99.6594
R8027 gnd.n3835 gnd.n3791 99.6594
R8028 gnd.n3831 gnd.n3792 99.6594
R8029 gnd.n3827 gnd.n3793 99.6594
R8030 gnd.n3874 gnd.n3782 99.6594
R8031 gnd.n5712 gnd.n5711 99.6594
R8032 gnd.n5715 gnd.n5714 99.6594
R8033 gnd.n5726 gnd.n5725 99.6594
R8034 gnd.n5735 gnd.n5734 99.6594
R8035 gnd.n5738 gnd.n5737 99.6594
R8036 gnd.n5749 gnd.n5748 99.6594
R8037 gnd.n5758 gnd.n5757 99.6594
R8038 gnd.n5761 gnd.n5760 99.6594
R8039 gnd.n5766 gnd.n5765 99.6594
R8040 gnd.n4817 gnd.n4731 99.6594
R8041 gnd.n4816 gnd.n4815 99.6594
R8042 gnd.n4809 gnd.n4735 99.6594
R8043 gnd.n4808 gnd.n4807 99.6594
R8044 gnd.n4801 gnd.n4741 99.6594
R8045 gnd.n4800 gnd.n4799 99.6594
R8046 gnd.n4793 gnd.n4747 99.6594
R8047 gnd.n4792 gnd.n4791 99.6594
R8048 gnd.n4781 gnd.n4753 99.6594
R8049 gnd.n4818 gnd.n4817 99.6594
R8050 gnd.n4815 gnd.n4814 99.6594
R8051 gnd.n4810 gnd.n4809 99.6594
R8052 gnd.n4807 gnd.n4806 99.6594
R8053 gnd.n4802 gnd.n4801 99.6594
R8054 gnd.n4799 gnd.n4798 99.6594
R8055 gnd.n4794 gnd.n4793 99.6594
R8056 gnd.n4791 gnd.n4790 99.6594
R8057 gnd.n4782 gnd.n4781 99.6594
R8058 gnd.n5765 gnd.n5764 99.6594
R8059 gnd.n5760 gnd.n5759 99.6594
R8060 gnd.n5757 gnd.n5750 99.6594
R8061 gnd.n5748 gnd.n5747 99.6594
R8062 gnd.n5737 gnd.n5736 99.6594
R8063 gnd.n5734 gnd.n5727 99.6594
R8064 gnd.n5725 gnd.n5724 99.6594
R8065 gnd.n5714 gnd.n5713 99.6594
R8066 gnd.n5711 gnd.n5701 99.6594
R8067 gnd.n3872 gnd.n3795 99.6594
R8068 gnd.n3864 gnd.n3783 99.6594
R8069 gnd.n3860 gnd.n3784 99.6594
R8070 gnd.n3856 gnd.n3785 99.6594
R8071 gnd.n3852 gnd.n3786 99.6594
R8072 gnd.n3848 gnd.n3787 99.6594
R8073 gnd.n3844 gnd.n3788 99.6594
R8074 gnd.n3840 gnd.n3789 99.6594
R8075 gnd.n3836 gnd.n3790 99.6594
R8076 gnd.n3832 gnd.n3791 99.6594
R8077 gnd.n3828 gnd.n3792 99.6594
R8078 gnd.n3824 gnd.n3793 99.6594
R8079 gnd.n3875 gnd.n3874 99.6594
R8080 gnd.n4640 gnd.n1833 99.6594
R8081 gnd.n4644 gnd.n1832 99.6594
R8082 gnd.n4648 gnd.n1831 99.6594
R8083 gnd.n4652 gnd.n1830 99.6594
R8084 gnd.n4656 gnd.n1829 99.6594
R8085 gnd.n4660 gnd.n1828 99.6594
R8086 gnd.n4664 gnd.n1827 99.6594
R8087 gnd.n4668 gnd.n1826 99.6594
R8088 gnd.n4672 gnd.n1825 99.6594
R8089 gnd.n4676 gnd.n1824 99.6594
R8090 gnd.n4680 gnd.n1823 99.6594
R8091 gnd.n4684 gnd.n1822 99.6594
R8092 gnd.n1862 gnd.n1821 99.6594
R8093 gnd.n705 gnd.n618 99.6594
R8094 gnd.n713 gnd.n619 99.6594
R8095 gnd.n715 gnd.n620 99.6594
R8096 gnd.n723 gnd.n621 99.6594
R8097 gnd.n731 gnd.n622 99.6594
R8098 gnd.n733 gnd.n623 99.6594
R8099 gnd.n741 gnd.n624 99.6594
R8100 gnd.n751 gnd.n625 99.6594
R8101 gnd.n6874 gnd.n626 99.6594
R8102 gnd.n7441 gnd.n260 99.6594
R8103 gnd.n7439 gnd.n259 99.6594
R8104 gnd.n7431 gnd.n258 99.6594
R8105 gnd.n7429 gnd.n257 99.6594
R8106 gnd.n7421 gnd.n256 99.6594
R8107 gnd.n7419 gnd.n255 99.6594
R8108 gnd.n7411 gnd.n254 99.6594
R8109 gnd.n7409 gnd.n253 99.6594
R8110 gnd.n7403 gnd.n252 99.6594
R8111 gnd.n3958 gnd.n3957 99.6594
R8112 gnd.n3717 gnd.n3695 99.6594
R8113 gnd.n3723 gnd.n3696 99.6594
R8114 gnd.n3727 gnd.n3697 99.6594
R8115 gnd.n3733 gnd.n3698 99.6594
R8116 gnd.n3737 gnd.n3699 99.6594
R8117 gnd.n3743 gnd.n3700 99.6594
R8118 gnd.n3701 gnd.n3685 99.6594
R8119 gnd.n4694 gnd.n1834 99.6594
R8120 gnd.n4698 gnd.n1835 99.6594
R8121 gnd.n4702 gnd.n1836 99.6594
R8122 gnd.n4706 gnd.n1837 99.6594
R8123 gnd.n4710 gnd.n1838 99.6594
R8124 gnd.n4714 gnd.n1839 99.6594
R8125 gnd.n4718 gnd.n1840 99.6594
R8126 gnd.n1843 gnd.n1841 99.6594
R8127 gnd.n4886 gnd.n4885 99.6594
R8128 gnd.n4894 gnd.n4893 99.6594
R8129 gnd.n4895 gnd.n4878 99.6594
R8130 gnd.n4904 gnd.n4903 99.6594
R8131 gnd.n4905 gnd.n4874 99.6594
R8132 gnd.n4914 gnd.n4913 99.6594
R8133 gnd.n4915 gnd.n4870 99.6594
R8134 gnd.n4924 gnd.n4923 99.6594
R8135 gnd.n4925 gnd.n4863 99.6594
R8136 gnd.n4934 gnd.n4933 99.6594
R8137 gnd.n4935 gnd.n4859 99.6594
R8138 gnd.n4944 gnd.n4943 99.6594
R8139 gnd.n4945 gnd.n4855 99.6594
R8140 gnd.n4954 gnd.n4953 99.6594
R8141 gnd.n4955 gnd.n4851 99.6594
R8142 gnd.n4964 gnd.n4963 99.6594
R8143 gnd.n4965 gnd.n4847 99.6594
R8144 gnd.n4974 gnd.n4973 99.6594
R8145 gnd.n4975 gnd.n4843 99.6594
R8146 gnd.n4986 gnd.n4985 99.6594
R8147 gnd.n4987 gnd.n4839 99.6594
R8148 gnd.n4996 gnd.n4995 99.6594
R8149 gnd.n4997 gnd.n4835 99.6594
R8150 gnd.n5006 gnd.n5005 99.6594
R8151 gnd.n5007 gnd.n4831 99.6594
R8152 gnd.n5016 gnd.n5015 99.6594
R8153 gnd.n5017 gnd.n4827 99.6594
R8154 gnd.n5027 gnd.n5026 99.6594
R8155 gnd.n5030 gnd.n5029 99.6594
R8156 gnd.n5976 gnd.n5975 99.6594
R8157 gnd.n1418 gnd.n1410 99.6594
R8158 gnd.n5983 gnd.n5982 99.6594
R8159 gnd.n1409 gnd.n1403 99.6594
R8160 gnd.n5990 gnd.n5989 99.6594
R8161 gnd.n1402 gnd.n1396 99.6594
R8162 gnd.n5997 gnd.n5996 99.6594
R8163 gnd.n1395 gnd.n1389 99.6594
R8164 gnd.n6004 gnd.n6003 99.6594
R8165 gnd.n6007 gnd.n6006 99.6594
R8166 gnd.n1386 gnd.n1378 99.6594
R8167 gnd.n6016 gnd.n6015 99.6594
R8168 gnd.n1377 gnd.n1371 99.6594
R8169 gnd.n6023 gnd.n6022 99.6594
R8170 gnd.n6026 gnd.n6025 99.6594
R8171 gnd.n5916 gnd.n5915 99.6594
R8172 gnd.n5914 gnd.n5909 99.6594
R8173 gnd.n5923 gnd.n5922 99.6594
R8174 gnd.n5908 gnd.n5899 99.6594
R8175 gnd.n5930 gnd.n5929 99.6594
R8176 gnd.n5898 gnd.n5892 99.6594
R8177 gnd.n5937 gnd.n5936 99.6594
R8178 gnd.n5891 gnd.n5885 99.6594
R8179 gnd.n5944 gnd.n5943 99.6594
R8180 gnd.n5884 gnd.n5878 99.6594
R8181 gnd.n5951 gnd.n5950 99.6594
R8182 gnd.n5877 gnd.n5872 99.6594
R8183 gnd.n5958 gnd.n5957 99.6594
R8184 gnd.n7040 gnd.n7039 99.6594
R8185 gnd.n7033 gnd.n590 99.6594
R8186 gnd.n7029 gnd.n591 99.6594
R8187 gnd.n7025 gnd.n592 99.6594
R8188 gnd.n7021 gnd.n593 99.6594
R8189 gnd.n7017 gnd.n594 99.6594
R8190 gnd.n7013 gnd.n595 99.6594
R8191 gnd.n7009 gnd.n596 99.6594
R8192 gnd.n7004 gnd.n597 99.6594
R8193 gnd.n7000 gnd.n598 99.6594
R8194 gnd.n6996 gnd.n599 99.6594
R8195 gnd.n6992 gnd.n600 99.6594
R8196 gnd.n6987 gnd.n602 99.6594
R8197 gnd.n6983 gnd.n603 99.6594
R8198 gnd.n6979 gnd.n604 99.6594
R8199 gnd.n6975 gnd.n605 99.6594
R8200 gnd.n6971 gnd.n606 99.6594
R8201 gnd.n6967 gnd.n607 99.6594
R8202 gnd.n6963 gnd.n608 99.6594
R8203 gnd.n6959 gnd.n609 99.6594
R8204 gnd.n6955 gnd.n610 99.6594
R8205 gnd.n6951 gnd.n611 99.6594
R8206 gnd.n6947 gnd.n612 99.6594
R8207 gnd.n6943 gnd.n613 99.6594
R8208 gnd.n6939 gnd.n614 99.6594
R8209 gnd.n6935 gnd.n615 99.6594
R8210 gnd.n6931 gnd.n616 99.6594
R8211 gnd.n691 gnd.n617 99.6594
R8212 gnd.n7544 gnd.n261 99.6594
R8213 gnd.n7548 gnd.n262 99.6594
R8214 gnd.n7552 gnd.n263 99.6594
R8215 gnd.n7556 gnd.n264 99.6594
R8216 gnd.n7560 gnd.n265 99.6594
R8217 gnd.n7564 gnd.n266 99.6594
R8218 gnd.n7568 gnd.n267 99.6594
R8219 gnd.n7572 gnd.n268 99.6594
R8220 gnd.n7576 gnd.n269 99.6594
R8221 gnd.n7580 gnd.n270 99.6594
R8222 gnd.n7586 gnd.n271 99.6594
R8223 gnd.n7590 gnd.n272 99.6594
R8224 gnd.n7594 gnd.n273 99.6594
R8225 gnd.n7598 gnd.n274 99.6594
R8226 gnd.n7602 gnd.n275 99.6594
R8227 gnd.n7606 gnd.n276 99.6594
R8228 gnd.n7610 gnd.n277 99.6594
R8229 gnd.n7614 gnd.n278 99.6594
R8230 gnd.n7618 gnd.n279 99.6594
R8231 gnd.n7622 gnd.n280 99.6594
R8232 gnd.n7629 gnd.n281 99.6594
R8233 gnd.n7633 gnd.n282 99.6594
R8234 gnd.n7637 gnd.n283 99.6594
R8235 gnd.n7641 gnd.n284 99.6594
R8236 gnd.n7645 gnd.n285 99.6594
R8237 gnd.n7649 gnd.n286 99.6594
R8238 gnd.n7653 gnd.n287 99.6594
R8239 gnd.n289 gnd.n288 99.6594
R8240 gnd.n7659 gnd.n250 99.6594
R8241 gnd.n5837 gnd.n5836 99.6594
R8242 gnd.n1481 gnd.n1461 99.6594
R8243 gnd.n1483 gnd.n1462 99.6594
R8244 gnd.n1485 gnd.n1463 99.6594
R8245 gnd.n5705 gnd.n1464 99.6594
R8246 gnd.n5708 gnd.n1465 99.6594
R8247 gnd.n5719 gnd.n1466 99.6594
R8248 gnd.n5721 gnd.n1467 99.6594
R8249 gnd.n5731 gnd.n1468 99.6594
R8250 gnd.n5742 gnd.n1469 99.6594
R8251 gnd.n5744 gnd.n1470 99.6594
R8252 gnd.n5754 gnd.n1471 99.6594
R8253 gnd.n5775 gnd.n1473 99.6594
R8254 gnd.n5839 gnd.n1458 99.6594
R8255 gnd.n5837 gnd.n1476 99.6594
R8256 gnd.n1482 gnd.n1461 99.6594
R8257 gnd.n1484 gnd.n1462 99.6594
R8258 gnd.n5704 gnd.n1463 99.6594
R8259 gnd.n5707 gnd.n1464 99.6594
R8260 gnd.n5718 gnd.n1465 99.6594
R8261 gnd.n5720 gnd.n1466 99.6594
R8262 gnd.n5730 gnd.n1467 99.6594
R8263 gnd.n5741 gnd.n1468 99.6594
R8264 gnd.n5743 gnd.n1469 99.6594
R8265 gnd.n5753 gnd.n1470 99.6594
R8266 gnd.n5774 gnd.n1471 99.6594
R8267 gnd.n1473 gnd.n1472 99.6594
R8268 gnd.n5840 gnd.n5839 99.6594
R8269 gnd.n777 gnd.n770 99.6594
R8270 gnd.n779 gnd.n778 99.6594
R8271 gnd.n6848 gnd.n775 99.6594
R8272 gnd.n6846 gnd.n698 99.6594
R8273 gnd.n780 gnd.n700 99.6594
R8274 gnd.n782 gnd.n709 99.6594
R8275 gnd.n784 gnd.n783 99.6594
R8276 gnd.n785 gnd.n720 99.6594
R8277 gnd.n787 gnd.n727 99.6594
R8278 gnd.n789 gnd.n788 99.6594
R8279 gnd.n790 gnd.n738 99.6594
R8280 gnd.n792 gnd.n745 99.6594
R8281 gnd.n794 gnd.n793 99.6594
R8282 gnd.n795 gnd.n757 99.6594
R8283 gnd.n792 gnd.n791 99.6594
R8284 gnd.n790 gnd.n737 99.6594
R8285 gnd.n789 gnd.n728 99.6594
R8286 gnd.n787 gnd.n786 99.6594
R8287 gnd.n785 gnd.n719 99.6594
R8288 gnd.n784 gnd.n710 99.6594
R8289 gnd.n782 gnd.n781 99.6594
R8290 gnd.n780 gnd.n699 99.6594
R8291 gnd.n6847 gnd.n6846 99.6594
R8292 gnd.n775 gnd.n774 99.6594
R8293 gnd.n779 gnd.n771 99.6594
R8294 gnd.n777 gnd.n766 99.6594
R8295 gnd.n795 gnd.n762 99.6594
R8296 gnd.n794 gnd.n756 99.6594
R8297 gnd.n5771 gnd.t21 98.63
R8298 gnd.n6875 gnd.t100 98.63
R8299 gnd.n5762 gnd.t118 98.63
R8300 gnd.n647 gnd.t97 98.63
R8301 gnd.n670 gnd.t91 98.63
R8302 gnd.n693 gnd.t35 98.63
R8303 gnd.n346 gnd.t124 98.63
R8304 gnd.n326 gnd.t42 98.63
R8305 gnd.n7625 gnd.t59 98.63
R8306 gnd.n7392 gnd.t77 98.63
R8307 gnd.n4867 gnd.t94 98.63
R8308 gnd.n4977 gnd.t39 98.63
R8309 gnd.n4823 gnd.t50 98.63
R8310 gnd.n4756 gnd.t122 98.63
R8311 gnd.n5900 gnd.t112 98.63
R8312 gnd.n1415 gnd.t46 98.63
R8313 gnd.n1382 gnd.t74 98.63
R8314 gnd.n747 gnd.t53 98.63
R8315 gnd.n1293 gnd.t31 88.9408
R8316 gnd.n927 gnd.t27 88.9408
R8317 gnd.n1290 gnd.t69 88.933
R8318 gnd.n6571 gnd.t65 88.933
R8319 gnd.n1275 gnd.n1274 81.8399
R8320 gnd.n3746 gnd.t84 74.8376
R8321 gnd.n1859 gnd.t110 74.8376
R8322 gnd.n1294 gnd.t30 72.8438
R8323 gnd.n928 gnd.t28 72.8438
R8324 gnd.n1276 gnd.n1269 72.8411
R8325 gnd.n1282 gnd.n1267 72.8411
R8326 gnd.n6567 gnd.n6566 72.8411
R8327 gnd.n5772 gnd.t20 72.836
R8328 gnd.n1291 gnd.t68 72.836
R8329 gnd.n6572 gnd.t66 72.836
R8330 gnd.n6876 gnd.t99 72.836
R8331 gnd.n5763 gnd.t119 72.836
R8332 gnd.n648 gnd.t96 72.836
R8333 gnd.n671 gnd.t90 72.836
R8334 gnd.n694 gnd.t34 72.836
R8335 gnd.n347 gnd.t125 72.836
R8336 gnd.n327 gnd.t43 72.836
R8337 gnd.n7626 gnd.t60 72.836
R8338 gnd.n7393 gnd.t78 72.836
R8339 gnd.n4868 gnd.t93 72.836
R8340 gnd.n4978 gnd.t38 72.836
R8341 gnd.n4824 gnd.t49 72.836
R8342 gnd.n4757 gnd.t121 72.836
R8343 gnd.n5901 gnd.t113 72.836
R8344 gnd.n1416 gnd.t47 72.836
R8345 gnd.n1383 gnd.t75 72.836
R8346 gnd.n748 gnd.t54 72.836
R8347 gnd.n6635 gnd.n893 71.676
R8348 gnd.n6631 gnd.n894 71.676
R8349 gnd.n6627 gnd.n895 71.676
R8350 gnd.n6623 gnd.n896 71.676
R8351 gnd.n6619 gnd.n897 71.676
R8352 gnd.n6615 gnd.n898 71.676
R8353 gnd.n6611 gnd.n899 71.676
R8354 gnd.n6607 gnd.n900 71.676
R8355 gnd.n6603 gnd.n901 71.676
R8356 gnd.n6599 gnd.n902 71.676
R8357 gnd.n6595 gnd.n903 71.676
R8358 gnd.n6591 gnd.n904 71.676
R8359 gnd.n6587 gnd.n905 71.676
R8360 gnd.n6583 gnd.n906 71.676
R8361 gnd.n6578 gnd.n907 71.676
R8362 gnd.n6574 gnd.n908 71.676
R8363 gnd.n6711 gnd.n926 71.676
R8364 gnd.n6707 gnd.n925 71.676
R8365 gnd.n6702 gnd.n924 71.676
R8366 gnd.n6698 gnd.n923 71.676
R8367 gnd.n6694 gnd.n922 71.676
R8368 gnd.n6690 gnd.n921 71.676
R8369 gnd.n6686 gnd.n920 71.676
R8370 gnd.n6682 gnd.n919 71.676
R8371 gnd.n6678 gnd.n918 71.676
R8372 gnd.n6674 gnd.n917 71.676
R8373 gnd.n6670 gnd.n916 71.676
R8374 gnd.n6666 gnd.n915 71.676
R8375 gnd.n6662 gnd.n914 71.676
R8376 gnd.n6658 gnd.n913 71.676
R8377 gnd.n6654 gnd.n912 71.676
R8378 gnd.n6650 gnd.n911 71.676
R8379 gnd.n6646 gnd.n910 71.676
R8380 gnd.n6098 gnd.n6097 71.676
R8381 gnd.n6092 gnd.n1228 71.676
R8382 gnd.n6089 gnd.n1229 71.676
R8383 gnd.n6085 gnd.n1230 71.676
R8384 gnd.n6081 gnd.n1231 71.676
R8385 gnd.n6077 gnd.n1232 71.676
R8386 gnd.n6073 gnd.n1233 71.676
R8387 gnd.n6069 gnd.n1234 71.676
R8388 gnd.n6065 gnd.n1235 71.676
R8389 gnd.n6061 gnd.n1236 71.676
R8390 gnd.n6057 gnd.n1237 71.676
R8391 gnd.n6053 gnd.n1238 71.676
R8392 gnd.n6049 gnd.n1239 71.676
R8393 gnd.n6045 gnd.n1240 71.676
R8394 gnd.n6041 gnd.n1241 71.676
R8395 gnd.n6037 gnd.n1242 71.676
R8396 gnd.n6033 gnd.n1244 71.676
R8397 gnd.n1357 gnd.n1245 71.676
R8398 gnd.n1352 gnd.n1246 71.676
R8399 gnd.n1348 gnd.n1247 71.676
R8400 gnd.n1344 gnd.n1248 71.676
R8401 gnd.n1340 gnd.n1249 71.676
R8402 gnd.n1336 gnd.n1250 71.676
R8403 gnd.n1332 gnd.n1251 71.676
R8404 gnd.n1328 gnd.n1252 71.676
R8405 gnd.n1324 gnd.n1253 71.676
R8406 gnd.n1320 gnd.n1254 71.676
R8407 gnd.n1316 gnd.n1255 71.676
R8408 gnd.n1312 gnd.n1256 71.676
R8409 gnd.n1308 gnd.n1257 71.676
R8410 gnd.n1304 gnd.n1258 71.676
R8411 gnd.n1300 gnd.n1259 71.676
R8412 gnd.n6098 gnd.n1264 71.676
R8413 gnd.n6090 gnd.n1228 71.676
R8414 gnd.n6086 gnd.n1229 71.676
R8415 gnd.n6082 gnd.n1230 71.676
R8416 gnd.n6078 gnd.n1231 71.676
R8417 gnd.n6074 gnd.n1232 71.676
R8418 gnd.n6070 gnd.n1233 71.676
R8419 gnd.n6066 gnd.n1234 71.676
R8420 gnd.n6062 gnd.n1235 71.676
R8421 gnd.n6058 gnd.n1236 71.676
R8422 gnd.n6054 gnd.n1237 71.676
R8423 gnd.n6050 gnd.n1238 71.676
R8424 gnd.n6046 gnd.n1239 71.676
R8425 gnd.n6042 gnd.n1240 71.676
R8426 gnd.n6038 gnd.n1241 71.676
R8427 gnd.n6034 gnd.n1243 71.676
R8428 gnd.n1358 gnd.n1244 71.676
R8429 gnd.n1353 gnd.n1245 71.676
R8430 gnd.n1349 gnd.n1246 71.676
R8431 gnd.n1345 gnd.n1247 71.676
R8432 gnd.n1341 gnd.n1248 71.676
R8433 gnd.n1337 gnd.n1249 71.676
R8434 gnd.n1333 gnd.n1250 71.676
R8435 gnd.n1329 gnd.n1251 71.676
R8436 gnd.n1325 gnd.n1252 71.676
R8437 gnd.n1321 gnd.n1253 71.676
R8438 gnd.n1317 gnd.n1254 71.676
R8439 gnd.n1313 gnd.n1255 71.676
R8440 gnd.n1309 gnd.n1256 71.676
R8441 gnd.n1305 gnd.n1257 71.676
R8442 gnd.n1301 gnd.n1258 71.676
R8443 gnd.n1297 gnd.n1259 71.676
R8444 gnd.n6649 gnd.n910 71.676
R8445 gnd.n6653 gnd.n911 71.676
R8446 gnd.n6657 gnd.n912 71.676
R8447 gnd.n6661 gnd.n913 71.676
R8448 gnd.n6665 gnd.n914 71.676
R8449 gnd.n6669 gnd.n915 71.676
R8450 gnd.n6673 gnd.n916 71.676
R8451 gnd.n6677 gnd.n917 71.676
R8452 gnd.n6681 gnd.n918 71.676
R8453 gnd.n6685 gnd.n919 71.676
R8454 gnd.n6689 gnd.n920 71.676
R8455 gnd.n6693 gnd.n921 71.676
R8456 gnd.n6697 gnd.n922 71.676
R8457 gnd.n6701 gnd.n923 71.676
R8458 gnd.n6706 gnd.n924 71.676
R8459 gnd.n6710 gnd.n925 71.676
R8460 gnd.n6573 gnd.n909 71.676
R8461 gnd.n6577 gnd.n908 71.676
R8462 gnd.n6582 gnd.n907 71.676
R8463 gnd.n6586 gnd.n906 71.676
R8464 gnd.n6590 gnd.n905 71.676
R8465 gnd.n6594 gnd.n904 71.676
R8466 gnd.n6598 gnd.n903 71.676
R8467 gnd.n6602 gnd.n902 71.676
R8468 gnd.n6606 gnd.n901 71.676
R8469 gnd.n6610 gnd.n900 71.676
R8470 gnd.n6614 gnd.n899 71.676
R8471 gnd.n6618 gnd.n898 71.676
R8472 gnd.n6622 gnd.n897 71.676
R8473 gnd.n6626 gnd.n896 71.676
R8474 gnd.n6630 gnd.n895 71.676
R8475 gnd.n6634 gnd.n894 71.676
R8476 gnd.n6637 gnd.n893 71.676
R8477 gnd.n8 gnd.t169 69.1507
R8478 gnd.n14 gnd.t156 68.4792
R8479 gnd.n13 gnd.t146 68.4792
R8480 gnd.n12 gnd.t388 68.4792
R8481 gnd.n11 gnd.t171 68.4792
R8482 gnd.n10 gnd.t5 68.4792
R8483 gnd.n9 gnd.t140 68.4792
R8484 gnd.n8 gnd.t142 68.4792
R8485 gnd.n3873 gnd.n3777 64.369
R8486 gnd.n2603 gnd.n2602 61.9869
R8487 gnd.n1355 gnd.n1294 59.5399
R8488 gnd.n6704 gnd.n928 59.5399
R8489 gnd.n1292 gnd.n1291 59.5399
R8490 gnd.n6580 gnd.n6572 59.5399
R8491 gnd.n1289 gnd.n1285 59.1804
R8492 gnd.n4726 gnd.n1819 57.3586
R8493 gnd.n3524 gnd.t277 56.407
R8494 gnd.n3465 gnd.t363 56.407
R8495 gnd.n3484 gnd.t216 56.407
R8496 gnd.n3504 gnd.t350 56.407
R8497 gnd.n76 gnd.t245 56.407
R8498 gnd.n17 gnd.t232 56.407
R8499 gnd.n36 gnd.t374 56.407
R8500 gnd.n56 gnd.t300 56.407
R8501 gnd.n3541 gnd.t335 55.8337
R8502 gnd.n3482 gnd.t205 55.8337
R8503 gnd.n3501 gnd.t365 55.8337
R8504 gnd.n3521 gnd.t238 55.8337
R8505 gnd.n93 gnd.t258 55.8337
R8506 gnd.n34 gnd.t226 55.8337
R8507 gnd.n53 gnd.t325 55.8337
R8508 gnd.n73 gnd.t316 55.8337
R8509 gnd.n1273 gnd.n1272 54.358
R8510 gnd.n6564 gnd.n6563 54.358
R8511 gnd.n3524 gnd.n3523 53.0052
R8512 gnd.n3526 gnd.n3525 53.0052
R8513 gnd.n3528 gnd.n3527 53.0052
R8514 gnd.n3530 gnd.n3529 53.0052
R8515 gnd.n3532 gnd.n3531 53.0052
R8516 gnd.n3534 gnd.n3533 53.0052
R8517 gnd.n3536 gnd.n3535 53.0052
R8518 gnd.n3538 gnd.n3537 53.0052
R8519 gnd.n3540 gnd.n3539 53.0052
R8520 gnd.n3465 gnd.n3464 53.0052
R8521 gnd.n3467 gnd.n3466 53.0052
R8522 gnd.n3469 gnd.n3468 53.0052
R8523 gnd.n3471 gnd.n3470 53.0052
R8524 gnd.n3473 gnd.n3472 53.0052
R8525 gnd.n3475 gnd.n3474 53.0052
R8526 gnd.n3477 gnd.n3476 53.0052
R8527 gnd.n3479 gnd.n3478 53.0052
R8528 gnd.n3481 gnd.n3480 53.0052
R8529 gnd.n3484 gnd.n3483 53.0052
R8530 gnd.n3486 gnd.n3485 53.0052
R8531 gnd.n3488 gnd.n3487 53.0052
R8532 gnd.n3490 gnd.n3489 53.0052
R8533 gnd.n3492 gnd.n3491 53.0052
R8534 gnd.n3494 gnd.n3493 53.0052
R8535 gnd.n3496 gnd.n3495 53.0052
R8536 gnd.n3498 gnd.n3497 53.0052
R8537 gnd.n3500 gnd.n3499 53.0052
R8538 gnd.n3504 gnd.n3503 53.0052
R8539 gnd.n3506 gnd.n3505 53.0052
R8540 gnd.n3508 gnd.n3507 53.0052
R8541 gnd.n3510 gnd.n3509 53.0052
R8542 gnd.n3512 gnd.n3511 53.0052
R8543 gnd.n3514 gnd.n3513 53.0052
R8544 gnd.n3516 gnd.n3515 53.0052
R8545 gnd.n3518 gnd.n3517 53.0052
R8546 gnd.n3520 gnd.n3519 53.0052
R8547 gnd.n92 gnd.n91 53.0052
R8548 gnd.n90 gnd.n89 53.0052
R8549 gnd.n88 gnd.n87 53.0052
R8550 gnd.n86 gnd.n85 53.0052
R8551 gnd.n84 gnd.n83 53.0052
R8552 gnd.n82 gnd.n81 53.0052
R8553 gnd.n80 gnd.n79 53.0052
R8554 gnd.n78 gnd.n77 53.0052
R8555 gnd.n76 gnd.n75 53.0052
R8556 gnd.n33 gnd.n32 53.0052
R8557 gnd.n31 gnd.n30 53.0052
R8558 gnd.n29 gnd.n28 53.0052
R8559 gnd.n27 gnd.n26 53.0052
R8560 gnd.n25 gnd.n24 53.0052
R8561 gnd.n23 gnd.n22 53.0052
R8562 gnd.n21 gnd.n20 53.0052
R8563 gnd.n19 gnd.n18 53.0052
R8564 gnd.n17 gnd.n16 53.0052
R8565 gnd.n52 gnd.n51 53.0052
R8566 gnd.n50 gnd.n49 53.0052
R8567 gnd.n48 gnd.n47 53.0052
R8568 gnd.n46 gnd.n45 53.0052
R8569 gnd.n44 gnd.n43 53.0052
R8570 gnd.n42 gnd.n41 53.0052
R8571 gnd.n40 gnd.n39 53.0052
R8572 gnd.n38 gnd.n37 53.0052
R8573 gnd.n36 gnd.n35 53.0052
R8574 gnd.n72 gnd.n71 53.0052
R8575 gnd.n70 gnd.n69 53.0052
R8576 gnd.n68 gnd.n67 53.0052
R8577 gnd.n66 gnd.n65 53.0052
R8578 gnd.n64 gnd.n63 53.0052
R8579 gnd.n62 gnd.n61 53.0052
R8580 gnd.n60 gnd.n59 53.0052
R8581 gnd.n58 gnd.n57 53.0052
R8582 gnd.n56 gnd.n55 53.0052
R8583 gnd.n6555 gnd.n6554 52.4801
R8584 gnd.n4577 gnd.t152 52.3082
R8585 gnd.n4545 gnd.t158 52.3082
R8586 gnd.n4513 gnd.t386 52.3082
R8587 gnd.n4482 gnd.t154 52.3082
R8588 gnd.n4450 gnd.t394 52.3082
R8589 gnd.n4418 gnd.t134 52.3082
R8590 gnd.n4386 gnd.t167 52.3082
R8591 gnd.n4355 gnd.t161 52.3082
R8592 gnd.n5043 gnd.n4727 51.6227
R8593 gnd.n7660 gnd.n244 51.6227
R8594 gnd.n4407 gnd.n4375 51.4173
R8595 gnd.n4471 gnd.n4470 50.455
R8596 gnd.n4439 gnd.n4438 50.455
R8597 gnd.n4407 gnd.n4406 50.455
R8598 gnd.n3820 gnd.n3819 45.1884
R8599 gnd.n1885 gnd.n1884 45.1884
R8600 gnd.n6639 gnd.n6570 44.3322
R8601 gnd.n1276 gnd.n1275 44.3189
R8602 gnd.n5773 gnd.n5772 42.2793
R8603 gnd.n6877 gnd.n6876 42.2793
R8604 gnd.n3821 gnd.n3820 42.2793
R8605 gnd.n1886 gnd.n1885 42.2793
R8606 gnd.n3747 gnd.n3746 42.2793
R8607 gnd.n4693 gnd.n1859 42.2793
R8608 gnd.n5768 gnd.n5763 42.2793
R8609 gnd.n7006 gnd.n648 42.2793
R8610 gnd.n6969 gnd.n671 42.2793
R8611 gnd.n6929 gnd.n694 42.2793
R8612 gnd.n7543 gnd.n347 42.2793
R8613 gnd.n7585 gnd.n327 42.2793
R8614 gnd.n7627 gnd.n7626 42.2793
R8615 gnd.n7394 gnd.n7393 42.2793
R8616 gnd.n4869 gnd.n4868 42.2793
R8617 gnd.n4979 gnd.n4978 42.2793
R8618 gnd.n4825 gnd.n4824 42.2793
R8619 gnd.n4758 gnd.n4757 42.2793
R8620 gnd.n5902 gnd.n5901 42.2793
R8621 gnd.n1417 gnd.n1416 42.2793
R8622 gnd.n6012 gnd.n1383 42.2793
R8623 gnd.n749 gnd.n748 42.2793
R8624 gnd.n1274 gnd.n1273 41.6274
R8625 gnd.n6565 gnd.n6564 41.6274
R8626 gnd.n1283 gnd.n1282 40.8975
R8627 gnd.n6568 gnd.n6567 40.8975
R8628 gnd.n1282 gnd.n1281 35.055
R8629 gnd.n1277 gnd.n1276 35.055
R8630 gnd.n6557 gnd.n6556 35.055
R8631 gnd.n6567 gnd.n6553 35.055
R8632 gnd.n3112 gnd.n3111 34.3058
R8633 gnd.n3112 gnd.n2093 34.3058
R8634 gnd.n3120 gnd.n2093 34.3058
R8635 gnd.n3121 gnd.n3120 34.3058
R8636 gnd.n3122 gnd.n3121 34.3058
R8637 gnd.n3122 gnd.n2087 34.3058
R8638 gnd.n3130 gnd.n2087 34.3058
R8639 gnd.n3131 gnd.n3130 34.3058
R8640 gnd.n3132 gnd.n3131 34.3058
R8641 gnd.n3132 gnd.n2081 34.3058
R8642 gnd.n3140 gnd.n2081 34.3058
R8643 gnd.n3141 gnd.n3140 34.3058
R8644 gnd.n3142 gnd.n3141 34.3058
R8645 gnd.n3142 gnd.n2075 34.3058
R8646 gnd.n3150 gnd.n2075 34.3058
R8647 gnd.n3151 gnd.n3150 34.3058
R8648 gnd.n3152 gnd.n3151 34.3058
R8649 gnd.n3152 gnd.n2069 34.3058
R8650 gnd.n3160 gnd.n2069 34.3058
R8651 gnd.n3161 gnd.n3160 34.3058
R8652 gnd.n3162 gnd.n3161 34.3058
R8653 gnd.n3162 gnd.n2063 34.3058
R8654 gnd.n3170 gnd.n2063 34.3058
R8655 gnd.n3171 gnd.n3170 34.3058
R8656 gnd.n3172 gnd.n3171 34.3058
R8657 gnd.n3172 gnd.n2057 34.3058
R8658 gnd.n3180 gnd.n2057 34.3058
R8659 gnd.n3181 gnd.n3180 34.3058
R8660 gnd.n3182 gnd.n3181 34.3058
R8661 gnd.n3182 gnd.n2051 34.3058
R8662 gnd.n3190 gnd.n2051 34.3058
R8663 gnd.n3191 gnd.n3190 34.3058
R8664 gnd.n3192 gnd.n3191 34.3058
R8665 gnd.n3192 gnd.n2045 34.3058
R8666 gnd.n3200 gnd.n2045 34.3058
R8667 gnd.n3201 gnd.n3200 34.3058
R8668 gnd.n3202 gnd.n3201 34.3058
R8669 gnd.n3202 gnd.n2039 34.3058
R8670 gnd.n3210 gnd.n2039 34.3058
R8671 gnd.n3211 gnd.n3210 34.3058
R8672 gnd.n3212 gnd.n3211 34.3058
R8673 gnd.n3212 gnd.n2033 34.3058
R8674 gnd.n3220 gnd.n2033 34.3058
R8675 gnd.n3221 gnd.n3220 34.3058
R8676 gnd.n3222 gnd.n3221 34.3058
R8677 gnd.n3222 gnd.n2027 34.3058
R8678 gnd.n3230 gnd.n2027 34.3058
R8679 gnd.n3231 gnd.n3230 34.3058
R8680 gnd.n3232 gnd.n3231 34.3058
R8681 gnd.n3232 gnd.n2021 34.3058
R8682 gnd.n3240 gnd.n2021 34.3058
R8683 gnd.n3241 gnd.n3240 34.3058
R8684 gnd.n3242 gnd.n3241 34.3058
R8685 gnd.n3242 gnd.n2015 34.3058
R8686 gnd.n3250 gnd.n2015 34.3058
R8687 gnd.n3251 gnd.n3250 34.3058
R8688 gnd.n3252 gnd.n3251 34.3058
R8689 gnd.n3252 gnd.n2009 34.3058
R8690 gnd.n3260 gnd.n2009 34.3058
R8691 gnd.n3261 gnd.n3260 34.3058
R8692 gnd.n3262 gnd.n3261 34.3058
R8693 gnd.n3262 gnd.n2003 34.3058
R8694 gnd.n3270 gnd.n2003 34.3058
R8695 gnd.n3271 gnd.n3270 34.3058
R8696 gnd.n3272 gnd.n3271 34.3058
R8697 gnd.n3272 gnd.n1997 34.3058
R8698 gnd.n3280 gnd.n1997 34.3058
R8699 gnd.n3281 gnd.n3280 34.3058
R8700 gnd.n3282 gnd.n3281 34.3058
R8701 gnd.n3282 gnd.n1991 34.3058
R8702 gnd.n3290 gnd.n1991 34.3058
R8703 gnd.n3291 gnd.n3290 34.3058
R8704 gnd.n3292 gnd.n3291 34.3058
R8705 gnd.n3292 gnd.n1985 34.3058
R8706 gnd.n3300 gnd.n1985 34.3058
R8707 gnd.n3301 gnd.n3300 34.3058
R8708 gnd.n3302 gnd.n3301 34.3058
R8709 gnd.n3302 gnd.n1979 34.3058
R8710 gnd.n3310 gnd.n1979 34.3058
R8711 gnd.n3311 gnd.n3310 34.3058
R8712 gnd.n3312 gnd.n3311 34.3058
R8713 gnd.n3312 gnd.n1910 34.3058
R8714 gnd.n3322 gnd.n1910 34.3058
R8715 gnd.n6647 gnd.n929 32.3127
R8716 gnd.n1298 gnd.n1295 32.3127
R8717 gnd.n3883 gnd.n3777 31.8661
R8718 gnd.n3883 gnd.n3882 31.8661
R8719 gnd.n3891 gnd.n3766 31.8661
R8720 gnd.n3899 gnd.n3766 31.8661
R8721 gnd.n3899 gnd.n3760 31.8661
R8722 gnd.n3907 gnd.n3760 31.8661
R8723 gnd.n3907 gnd.n3753 31.8661
R8724 gnd.n3945 gnd.n3753 31.8661
R8725 gnd.n3955 gnd.n3686 31.8661
R8726 gnd.n5043 gnd.n4730 31.8661
R8727 gnd.n5051 gnd.n1803 31.8661
R8728 gnd.n5063 gnd.n1803 31.8661
R8729 gnd.n5063 gnd.n1795 31.8661
R8730 gnd.n5071 gnd.n1795 31.8661
R8731 gnd.n5087 gnd.n1783 31.8661
R8732 gnd.n5087 gnd.n1786 31.8661
R8733 gnd.n5097 gnd.n1769 31.8661
R8734 gnd.n5107 gnd.n1769 31.8661
R8735 gnd.n5122 gnd.n1760 31.8661
R8736 gnd.n5132 gnd.n1744 31.8661
R8737 gnd.n5142 gnd.n1744 31.8661
R8738 gnd.n5157 gnd.n1725 31.8661
R8739 gnd.n5167 gnd.n1725 31.8661
R8740 gnd.n5177 gnd.n1719 31.8661
R8741 gnd.n5194 gnd.n1698 31.8661
R8742 gnd.n5204 gnd.n1698 31.8661
R8743 gnd.n5691 gnd.n5690 31.8661
R8744 gnd.n5691 gnd.n1460 31.8661
R8745 gnd.n5477 gnd.n1474 31.8661
R8746 gnd.n776 gnd.n764 31.8661
R8747 gnd.n6844 gnd.n589 31.8661
R8748 gnd.n7042 gnd.n589 31.8661
R8749 gnd.n7740 gnd.n131 31.8661
R8750 gnd.n7734 gnd.n131 31.8661
R8751 gnd.n7728 gnd.n146 31.8661
R8752 gnd.n7722 gnd.n156 31.8661
R8753 gnd.n7722 gnd.n159 31.8661
R8754 gnd.n7716 gnd.n168 31.8661
R8755 gnd.n7710 gnd.n168 31.8661
R8756 gnd.n7704 gnd.n184 31.8661
R8757 gnd.n7698 gnd.n194 31.8661
R8758 gnd.n7698 gnd.n197 31.8661
R8759 gnd.n7692 gnd.n206 31.8661
R8760 gnd.n7686 gnd.n206 31.8661
R8761 gnd.n7680 gnd.n222 31.8661
R8762 gnd.n7680 gnd.n225 31.8661
R8763 gnd.n7674 gnd.n225 31.8661
R8764 gnd.n7674 gnd.n235 31.8661
R8765 gnd.n7668 gnd.n244 31.8661
R8766 gnd.n5214 gnd.n1687 31.2288
R8767 gnd.n5222 gnd.n1679 31.2288
R8768 gnd.n5242 gnd.n1670 31.2288
R8769 gnd.n5237 gnd.n1662 31.2288
R8770 gnd.n5263 gnd.n1654 31.2288
R8771 gnd.n5258 gnd.n1657 31.2288
R8772 gnd.n5272 gnd.n1634 31.2288
R8773 gnd.n5289 gnd.n1637 31.2288
R8774 gnd.n5299 gnd.n1620 31.2288
R8775 gnd.n5282 gnd.n1611 31.2288
R8776 gnd.n5325 gnd.n1602 31.2288
R8777 gnd.n5335 gnd.n1591 31.2288
R8778 gnd.n5318 gnd.n1582 31.2288
R8779 gnd.n5367 gnd.n1571 31.2288
R8780 gnd.n5348 gnd.n1558 31.2288
R8781 gnd.n5387 gnd.n1550 31.2288
R8782 gnd.n5410 gnd.n1535 31.2288
R8783 gnd.n5353 gnd.n1523 31.2288
R8784 gnd.n5403 gnd.n1516 31.2288
R8785 gnd.n5432 gnd.n1505 31.2288
R8786 gnd.n5453 gnd.n1498 31.2288
R8787 gnd.n5452 gnd.n1446 31.2288
R8788 gnd.n5854 gnd.n1436 31.2288
R8789 gnd.n5864 gnd.n1439 31.2288
R8790 gnd.n5966 gnd.n1428 31.2288
R8791 gnd.n5698 gnd.n5697 31.2288
R8792 gnd.n7068 gnd.n569 31.2288
R8793 gnd.n7060 gnd.n572 31.2288
R8794 gnd.n577 gnd.n562 31.2288
R8795 gnd.n7087 gnd.n554 31.2288
R8796 gnd.n7118 gnd.n531 31.2288
R8797 gnd.n7099 gnd.n534 31.2288
R8798 gnd.n7111 gnd.n523 31.2288
R8799 gnd.n7110 gnd.n543 31.2288
R8800 gnd.n499 gnd.n487 31.2288
R8801 gnd.n7162 gnd.n7161 31.2288
R8802 gnd.n7188 gnd.n466 31.2288
R8803 gnd.n7198 gnd.n456 31.2288
R8804 gnd.n7181 gnd.n458 31.2288
R8805 gnd.n7228 gnd.n439 31.2288
R8806 gnd.n442 gnd.n431 31.2288
R8807 gnd.n7258 gnd.n423 31.2288
R8808 gnd.n7262 gnd.n414 31.2288
R8809 gnd.n7285 gnd.n402 31.2288
R8810 gnd.n7299 gnd.n395 31.2288
R8811 gnd.n7307 gnd.n387 31.2288
R8812 gnd.n7313 gnd.n7312 31.2288
R8813 gnd.n7323 gnd.n378 31.2288
R8814 gnd.n7335 gnd.n367 31.2288
R8815 gnd.n7343 gnd.n360 31.2288
R8816 gnd.n7353 gnd.n102 31.2288
R8817 gnd.n7746 gnd.n117 31.2288
R8818 gnd.t234 gnd.n1719 30.9101
R8819 gnd.n5214 gnd.n1691 30.9101
R8820 gnd.t202 gnd.n1685 30.9101
R8821 gnd.n5312 gnd.t282 30.9101
R8822 gnd.t249 gnd.n7236 30.9101
R8823 gnd.n7352 gnd.t260 30.9101
R8824 gnd.n7746 gnd.n120 30.9101
R8825 gnd.n7728 gnd.t209 30.9101
R8826 gnd.n5122 gnd.t213 30.2728
R8827 gnd.n5386 gnd.t254 30.2728
R8828 gnd.n7144 gnd.t211 30.2728
R8829 gnd.n7704 gnd.t291 30.2728
R8830 gnd.n4730 gnd.t37 28.3609
R8831 gnd.n7668 gnd.t41 28.3609
R8832 gnd.t45 gnd.n1426 27.7236
R8833 gnd.n7059 gnd.t33 27.7236
R8834 gnd.n5772 gnd.n5771 25.7944
R8835 gnd.n6876 gnd.n6875 25.7944
R8836 gnd.n3746 gnd.n3745 25.7944
R8837 gnd.n1859 gnd.n1858 25.7944
R8838 gnd.n5763 gnd.n5762 25.7944
R8839 gnd.n648 gnd.n647 25.7944
R8840 gnd.n671 gnd.n670 25.7944
R8841 gnd.n694 gnd.n693 25.7944
R8842 gnd.n347 gnd.n346 25.7944
R8843 gnd.n327 gnd.n326 25.7944
R8844 gnd.n7626 gnd.n7625 25.7944
R8845 gnd.n7393 gnd.n7392 25.7944
R8846 gnd.n4868 gnd.n4867 25.7944
R8847 gnd.n4978 gnd.n4977 25.7944
R8848 gnd.n4824 gnd.n4823 25.7944
R8849 gnd.n4757 gnd.n4756 25.7944
R8850 gnd.n5901 gnd.n5900 25.7944
R8851 gnd.n1416 gnd.n1415 25.7944
R8852 gnd.n1383 gnd.n1382 25.7944
R8853 gnd.n748 gnd.n747 25.7944
R8854 gnd.n3967 gnd.n3687 24.8557
R8855 gnd.n3977 gnd.n3670 24.8557
R8856 gnd.n3673 gnd.n3661 24.8557
R8857 gnd.n3998 gnd.n3662 24.8557
R8858 gnd.n4008 gnd.n3642 24.8557
R8859 gnd.n4018 gnd.n4017 24.8557
R8860 gnd.n3628 gnd.n3626 24.8557
R8861 gnd.n4049 gnd.n4048 24.8557
R8862 gnd.n4064 gnd.n3611 24.8557
R8863 gnd.n4118 gnd.n3550 24.8557
R8864 gnd.n4074 gnd.n3551 24.8557
R8865 gnd.n4111 gnd.n3562 24.8557
R8866 gnd.n3600 gnd.n3599 24.8557
R8867 gnd.n4105 gnd.n4104 24.8557
R8868 gnd.n3586 gnd.n3573 24.8557
R8869 gnd.n4144 gnd.n4143 24.8557
R8870 gnd.n4154 gnd.n3450 24.8557
R8871 gnd.n4166 gnd.n3442 24.8557
R8872 gnd.n4165 gnd.n3430 24.8557
R8873 gnd.n4184 gnd.n4183 24.8557
R8874 gnd.n4194 gnd.n3423 24.8557
R8875 gnd.n4205 gnd.n3411 24.8557
R8876 gnd.n4229 gnd.n4228 24.8557
R8877 gnd.n4240 gnd.n3394 24.8557
R8878 gnd.n4239 gnd.n3396 24.8557
R8879 gnd.n4251 gnd.n3387 24.8557
R8880 gnd.n4269 gnd.n4268 24.8557
R8881 gnd.n3378 gnd.n3367 24.8557
R8882 gnd.n4290 gnd.n3355 24.8557
R8883 gnd.n4318 gnd.n4317 24.8557
R8884 gnd.n4329 gnd.n3340 24.8557
R8885 gnd.n4340 gnd.n3333 24.8557
R8886 gnd.n4339 gnd.n1908 24.8557
R8887 gnd.n4635 gnd.n1893 24.8557
R8888 gnd.n3988 gnd.t160 23.2624
R8889 gnd.n5071 gnd.t204 23.2624
R8890 gnd.n3689 gnd.t83 22.6251
R8891 gnd.n1760 gnd.t223 22.6251
R8892 gnd.t215 gnd.n1508 22.6251
R8893 gnd.n7100 gnd.t231 22.6251
R8894 gnd.n184 gnd.t185 22.6251
R8895 gnd.n5177 gnd.t287 21.9878
R8896 gnd.t191 gnd.n1560 21.9878
R8897 gnd.t240 gnd.n469 21.9878
R8898 gnd.n146 gnd.t251 21.9878
R8899 gnd.t153 gnd.n3694 21.3504
R8900 gnd.n5229 gnd.t264 21.3504
R8901 gnd.t303 gnd.n1599 21.3504
R8902 gnd.n7257 gnd.t271 21.3504
R8903 gnd.n7754 gnd.t199 21.3504
R8904 gnd.t175 gnd.n3368 20.7131
R8905 gnd.n5185 gnd.t206 20.7131
R8906 gnd.t247 gnd.n1652 20.7131
R8907 gnd.n5276 gnd.t236 20.7131
R8908 gnd.n7268 gnd.t197 20.7131
R8909 gnd.n7322 gnd.t296 20.7131
R8910 gnd.n7490 gnd.t220 20.7131
R8911 gnd.n4612 gnd.n3322 20.5837
R8912 gnd.n5697 gnd.n1369 20.3945
R8913 gnd.n7041 gnd.n569 20.3945
R8914 gnd.n1289 gnd.n1288 20.1371
R8915 gnd.n6640 gnd.n6639 20.1371
R8916 gnd.t179 gnd.n3403 20.0758
R8917 gnd.n5157 gnd.t262 20.0758
R8918 gnd.n5344 gnd.t228 20.0758
R8919 gnd.n7216 gnd.t189 20.0758
R8920 gnd.t195 gnd.n159 20.0758
R8921 gnd.n1271 gnd.t88 19.8005
R8922 gnd.n1271 gnd.t24 19.8005
R8923 gnd.n1270 gnd.t72 19.8005
R8924 gnd.n1270 gnd.t116 19.8005
R8925 gnd.n6562 gnd.t13 19.8005
R8926 gnd.n6562 gnd.t81 19.8005
R8927 gnd.n6561 gnd.t103 19.8005
R8928 gnd.n6561 gnd.t57 19.8005
R8929 gnd.n1267 gnd.n1266 19.5087
R8930 gnd.n1280 gnd.n1267 19.5087
R8931 gnd.n1278 gnd.n1269 19.5087
R8932 gnd.n6566 gnd.n6560 19.5087
R8933 gnd.n4155 gnd.t183 19.4385
R8934 gnd.n5097 gnd.t217 19.4385
R8935 gnd.n5420 gnd.t187 19.4385
R8936 gnd.n7153 gnd.t193 19.4385
R8937 gnd.t301 gnd.n197 19.4385
R8938 gnd.n5556 gnd.n5555 19.3944
R8939 gnd.n5560 gnd.n5556 19.3944
R8940 gnd.n5560 gnd.n5552 19.3944
R8941 gnd.n5564 gnd.n5552 19.3944
R8942 gnd.n5564 gnd.n5541 19.3944
R8943 gnd.n5581 gnd.n5541 19.3944
R8944 gnd.n5581 gnd.n5539 19.3944
R8945 gnd.n5585 gnd.n5539 19.3944
R8946 gnd.n5585 gnd.n5529 19.3944
R8947 gnd.n5602 gnd.n5529 19.3944
R8948 gnd.n5602 gnd.n5527 19.3944
R8949 gnd.n5606 gnd.n5527 19.3944
R8950 gnd.n5606 gnd.n5517 19.3944
R8951 gnd.n5623 gnd.n5517 19.3944
R8952 gnd.n5623 gnd.n5514 19.3944
R8953 gnd.n5636 gnd.n5514 19.3944
R8954 gnd.n5636 gnd.n5515 19.3944
R8955 gnd.n5632 gnd.n5515 19.3944
R8956 gnd.n5632 gnd.n5631 19.3944
R8957 gnd.n5631 gnd.n5630 19.3944
R8958 gnd.n5630 gnd.n1216 19.3944
R8959 gnd.n6112 gnd.n1216 19.3944
R8960 gnd.n6113 gnd.n6112 19.3944
R8961 gnd.n6113 gnd.n1213 19.3944
R8962 gnd.n6143 gnd.n1213 19.3944
R8963 gnd.n6143 gnd.n1214 19.3944
R8964 gnd.n6139 gnd.n1214 19.3944
R8965 gnd.n6139 gnd.n6138 19.3944
R8966 gnd.n6138 gnd.n6137 19.3944
R8967 gnd.n6137 gnd.n6121 19.3944
R8968 gnd.n6133 gnd.n6121 19.3944
R8969 gnd.n6133 gnd.n6132 19.3944
R8970 gnd.n6132 gnd.n6131 19.3944
R8971 gnd.n6131 gnd.n6123 19.3944
R8972 gnd.n6127 gnd.n6123 19.3944
R8973 gnd.n6127 gnd.n6126 19.3944
R8974 gnd.n6126 gnd.n1097 19.3944
R8975 gnd.n6308 gnd.n1097 19.3944
R8976 gnd.n6309 gnd.n6308 19.3944
R8977 gnd.n6309 gnd.n1094 19.3944
R8978 gnd.n6339 gnd.n1094 19.3944
R8979 gnd.n6339 gnd.n1095 19.3944
R8980 gnd.n6335 gnd.n1095 19.3944
R8981 gnd.n6335 gnd.n6334 19.3944
R8982 gnd.n6334 gnd.n6333 19.3944
R8983 gnd.n6333 gnd.n6315 19.3944
R8984 gnd.n6329 gnd.n6315 19.3944
R8985 gnd.n6329 gnd.n6328 19.3944
R8986 gnd.n6328 gnd.n6327 19.3944
R8987 gnd.n6327 gnd.n6319 19.3944
R8988 gnd.n6323 gnd.n6319 19.3944
R8989 gnd.n6323 gnd.n6322 19.3944
R8990 gnd.n6322 gnd.n969 19.3944
R8991 gnd.n6501 gnd.n969 19.3944
R8992 gnd.n6501 gnd.n966 19.3944
R8993 gnd.n6505 gnd.n966 19.3944
R8994 gnd.n6506 gnd.n6505 19.3944
R8995 gnd.n6507 gnd.n6506 19.3944
R8996 gnd.n6507 gnd.n963 19.3944
R8997 gnd.n6516 gnd.n963 19.3944
R8998 gnd.n6516 gnd.n964 19.3944
R8999 gnd.n6512 gnd.n964 19.3944
R9000 gnd.n6512 gnd.n6511 19.3944
R9001 gnd.n6511 gnd.n871 19.3944
R9002 gnd.n6737 gnd.n871 19.3944
R9003 gnd.n6737 gnd.n868 19.3944
R9004 gnd.n6742 gnd.n868 19.3944
R9005 gnd.n6742 gnd.n869 19.3944
R9006 gnd.n869 gnd.n846 19.3944
R9007 gnd.n6767 gnd.n846 19.3944
R9008 gnd.n6767 gnd.n843 19.3944
R9009 gnd.n6772 gnd.n843 19.3944
R9010 gnd.n6772 gnd.n844 19.3944
R9011 gnd.n844 gnd.n822 19.3944
R9012 gnd.n6797 gnd.n822 19.3944
R9013 gnd.n6797 gnd.n819 19.3944
R9014 gnd.n6807 gnd.n819 19.3944
R9015 gnd.n6807 gnd.n820 19.3944
R9016 gnd.n6803 gnd.n820 19.3944
R9017 gnd.n6803 gnd.n6802 19.3944
R9018 gnd.n6802 gnd.n760 19.3944
R9019 gnd.n6863 gnd.n760 19.3944
R9020 gnd.n5776 gnd.n1457 19.3944
R9021 gnd.n5842 gnd.n1457 19.3944
R9022 gnd.n5842 gnd.n5841 19.3944
R9023 gnd.n5835 gnd.n5834 19.3944
R9024 gnd.n5834 gnd.n1479 19.3944
R9025 gnd.n5830 gnd.n1479 19.3944
R9026 gnd.n5830 gnd.n5829 19.3944
R9027 gnd.n5829 gnd.n5828 19.3944
R9028 gnd.n5828 gnd.n5825 19.3944
R9029 gnd.n5825 gnd.n5824 19.3944
R9030 gnd.n5824 gnd.n1486 19.3944
R9031 gnd.n5706 gnd.n1486 19.3944
R9032 gnd.n5816 gnd.n5706 19.3944
R9033 gnd.n5816 gnd.n5815 19.3944
R9034 gnd.n5815 gnd.n5709 19.3944
R9035 gnd.n5808 gnd.n5709 19.3944
R9036 gnd.n5808 gnd.n5807 19.3944
R9037 gnd.n5807 gnd.n5722 19.3944
R9038 gnd.n5800 gnd.n5722 19.3944
R9039 gnd.n5800 gnd.n5799 19.3944
R9040 gnd.n5799 gnd.n5732 19.3944
R9041 gnd.n5792 gnd.n5732 19.3944
R9042 gnd.n5792 gnd.n5791 19.3944
R9043 gnd.n5791 gnd.n5745 19.3944
R9044 gnd.n5784 gnd.n5745 19.3944
R9045 gnd.n5784 gnd.n5783 19.3944
R9046 gnd.n5783 gnd.n5755 19.3944
R9047 gnd.n6918 gnd.n704 19.3944
R9048 gnd.n6918 gnd.n6917 19.3944
R9049 gnd.n6917 gnd.n707 19.3944
R9050 gnd.n6910 gnd.n707 19.3944
R9051 gnd.n6910 gnd.n6909 19.3944
R9052 gnd.n6909 gnd.n717 19.3944
R9053 gnd.n6902 gnd.n717 19.3944
R9054 gnd.n6902 gnd.n6901 19.3944
R9055 gnd.n6901 gnd.n725 19.3944
R9056 gnd.n6894 gnd.n725 19.3944
R9057 gnd.n6894 gnd.n6893 19.3944
R9058 gnd.n6893 gnd.n735 19.3944
R9059 gnd.n6886 gnd.n735 19.3944
R9060 gnd.n6886 gnd.n6885 19.3944
R9061 gnd.n6885 gnd.n743 19.3944
R9062 gnd.n6878 gnd.n743 19.3944
R9063 gnd.n3870 gnd.n3869 19.3944
R9064 gnd.n3869 gnd.n3868 19.3944
R9065 gnd.n3868 gnd.n3867 19.3944
R9066 gnd.n3867 gnd.n3865 19.3944
R9067 gnd.n3865 gnd.n3862 19.3944
R9068 gnd.n3862 gnd.n3861 19.3944
R9069 gnd.n3861 gnd.n3858 19.3944
R9070 gnd.n3858 gnd.n3857 19.3944
R9071 gnd.n3857 gnd.n3854 19.3944
R9072 gnd.n3854 gnd.n3853 19.3944
R9073 gnd.n3853 gnd.n3850 19.3944
R9074 gnd.n3850 gnd.n3849 19.3944
R9075 gnd.n3849 gnd.n3846 19.3944
R9076 gnd.n3846 gnd.n3845 19.3944
R9077 gnd.n3845 gnd.n3842 19.3944
R9078 gnd.n3842 gnd.n3841 19.3944
R9079 gnd.n3841 gnd.n3838 19.3944
R9080 gnd.n3838 gnd.n3837 19.3944
R9081 gnd.n3837 gnd.n3834 19.3944
R9082 gnd.n3834 gnd.n3833 19.3944
R9083 gnd.n3833 gnd.n3830 19.3944
R9084 gnd.n3830 gnd.n3829 19.3944
R9085 gnd.n3826 gnd.n3825 19.3944
R9086 gnd.n3825 gnd.n3781 19.3944
R9087 gnd.n3876 gnd.n3781 19.3944
R9088 gnd.n4643 gnd.n4642 19.3944
R9089 gnd.n4642 gnd.n4639 19.3944
R9090 gnd.n4639 gnd.n4638 19.3944
R9091 gnd.n4688 gnd.n4687 19.3944
R9092 gnd.n4687 gnd.n4686 19.3944
R9093 gnd.n4686 gnd.n4683 19.3944
R9094 gnd.n4683 gnd.n4682 19.3944
R9095 gnd.n4682 gnd.n4679 19.3944
R9096 gnd.n4679 gnd.n4678 19.3944
R9097 gnd.n4678 gnd.n4675 19.3944
R9098 gnd.n4675 gnd.n4674 19.3944
R9099 gnd.n4674 gnd.n4671 19.3944
R9100 gnd.n4671 gnd.n4670 19.3944
R9101 gnd.n4670 gnd.n4667 19.3944
R9102 gnd.n4667 gnd.n4666 19.3944
R9103 gnd.n4666 gnd.n4663 19.3944
R9104 gnd.n4663 gnd.n4662 19.3944
R9105 gnd.n4662 gnd.n4659 19.3944
R9106 gnd.n4659 gnd.n4658 19.3944
R9107 gnd.n4658 gnd.n4655 19.3944
R9108 gnd.n4655 gnd.n4654 19.3944
R9109 gnd.n4654 gnd.n4651 19.3944
R9110 gnd.n4651 gnd.n4650 19.3944
R9111 gnd.n4650 gnd.n4647 19.3944
R9112 gnd.n4647 gnd.n4646 19.3944
R9113 gnd.n3969 gnd.n3678 19.3944
R9114 gnd.n3979 gnd.n3678 19.3944
R9115 gnd.n3980 gnd.n3979 19.3944
R9116 gnd.n3980 gnd.n3659 19.3944
R9117 gnd.n4000 gnd.n3659 19.3944
R9118 gnd.n4000 gnd.n3651 19.3944
R9119 gnd.n4010 gnd.n3651 19.3944
R9120 gnd.n4011 gnd.n4010 19.3944
R9121 gnd.n4012 gnd.n4011 19.3944
R9122 gnd.n4012 gnd.n3634 19.3944
R9123 gnd.n4029 gnd.n3634 19.3944
R9124 gnd.n4032 gnd.n4029 19.3944
R9125 gnd.n4032 gnd.n4031 19.3944
R9126 gnd.n4031 gnd.n3607 19.3944
R9127 gnd.n4071 gnd.n3607 19.3944
R9128 gnd.n4071 gnd.n3604 19.3944
R9129 gnd.n4077 gnd.n3604 19.3944
R9130 gnd.n4078 gnd.n4077 19.3944
R9131 gnd.n4078 gnd.n3602 19.3944
R9132 gnd.n4084 gnd.n3602 19.3944
R9133 gnd.n4087 gnd.n4084 19.3944
R9134 gnd.n4089 gnd.n4087 19.3944
R9135 gnd.n4095 gnd.n4089 19.3944
R9136 gnd.n4095 gnd.n4094 19.3944
R9137 gnd.n4094 gnd.n3445 19.3944
R9138 gnd.n4161 gnd.n3445 19.3944
R9139 gnd.n4162 gnd.n4161 19.3944
R9140 gnd.n4162 gnd.n3438 19.3944
R9141 gnd.n4173 gnd.n3438 19.3944
R9142 gnd.n4174 gnd.n4173 19.3944
R9143 gnd.n4174 gnd.n3421 19.3944
R9144 gnd.n3421 gnd.n3419 19.3944
R9145 gnd.n4198 gnd.n3419 19.3944
R9146 gnd.n4199 gnd.n4198 19.3944
R9147 gnd.n4199 gnd.n3390 19.3944
R9148 gnd.n4246 gnd.n3390 19.3944
R9149 gnd.n4247 gnd.n4246 19.3944
R9150 gnd.n4247 gnd.n3383 19.3944
R9151 gnd.n4258 gnd.n3383 19.3944
R9152 gnd.n4259 gnd.n4258 19.3944
R9153 gnd.n4259 gnd.n3366 19.3944
R9154 gnd.n3366 gnd.n3364 19.3944
R9155 gnd.n4283 gnd.n3364 19.3944
R9156 gnd.n4284 gnd.n4283 19.3944
R9157 gnd.n4284 gnd.n3336 19.3944
R9158 gnd.n4335 gnd.n3336 19.3944
R9159 gnd.n4336 gnd.n4335 19.3944
R9160 gnd.n4336 gnd.n3329 19.3944
R9161 gnd.n4603 gnd.n3329 19.3944
R9162 gnd.n4604 gnd.n4603 19.3944
R9163 gnd.n4604 gnd.n1897 19.3944
R9164 gnd.n4630 gnd.n1897 19.3944
R9165 gnd.n4630 gnd.n1898 19.3944
R9166 gnd.n3960 gnd.n3959 19.3944
R9167 gnd.n3959 gnd.n3692 19.3944
R9168 gnd.n3715 gnd.n3692 19.3944
R9169 gnd.n3718 gnd.n3715 19.3944
R9170 gnd.n3718 gnd.n3711 19.3944
R9171 gnd.n3722 gnd.n3711 19.3944
R9172 gnd.n3725 gnd.n3722 19.3944
R9173 gnd.n3728 gnd.n3725 19.3944
R9174 gnd.n3728 gnd.n3709 19.3944
R9175 gnd.n3732 gnd.n3709 19.3944
R9176 gnd.n3735 gnd.n3732 19.3944
R9177 gnd.n3738 gnd.n3735 19.3944
R9178 gnd.n3738 gnd.n3707 19.3944
R9179 gnd.n3742 gnd.n3707 19.3944
R9180 gnd.n3965 gnd.n3964 19.3944
R9181 gnd.n3964 gnd.n3668 19.3944
R9182 gnd.n3990 gnd.n3668 19.3944
R9183 gnd.n3990 gnd.n3666 19.3944
R9184 gnd.n3996 gnd.n3666 19.3944
R9185 gnd.n3996 gnd.n3995 19.3944
R9186 gnd.n3995 gnd.n3640 19.3944
R9187 gnd.n4020 gnd.n3640 19.3944
R9188 gnd.n4020 gnd.n3638 19.3944
R9189 gnd.n4024 gnd.n3638 19.3944
R9190 gnd.n4024 gnd.n3618 19.3944
R9191 gnd.n4051 gnd.n3618 19.3944
R9192 gnd.n4051 gnd.n3616 19.3944
R9193 gnd.n4061 gnd.n3616 19.3944
R9194 gnd.n4061 gnd.n4060 19.3944
R9195 gnd.n4060 gnd.n4059 19.3944
R9196 gnd.n4059 gnd.n3565 19.3944
R9197 gnd.n4109 gnd.n3565 19.3944
R9198 gnd.n4109 gnd.n4108 19.3944
R9199 gnd.n4108 gnd.n4107 19.3944
R9200 gnd.n4107 gnd.n3569 19.3944
R9201 gnd.n3589 gnd.n3569 19.3944
R9202 gnd.n3589 gnd.n3455 19.3944
R9203 gnd.n4146 gnd.n3455 19.3944
R9204 gnd.n4146 gnd.n3453 19.3944
R9205 gnd.n4152 gnd.n3453 19.3944
R9206 gnd.n4152 gnd.n4151 19.3944
R9207 gnd.n4151 gnd.n3428 19.3944
R9208 gnd.n4186 gnd.n3428 19.3944
R9209 gnd.n4186 gnd.n3426 19.3944
R9210 gnd.n4192 gnd.n3426 19.3944
R9211 gnd.n4192 gnd.n4191 19.3944
R9212 gnd.n4191 gnd.n3401 19.3944
R9213 gnd.n4231 gnd.n3401 19.3944
R9214 gnd.n4231 gnd.n3399 19.3944
R9215 gnd.n4237 gnd.n3399 19.3944
R9216 gnd.n4237 gnd.n4236 19.3944
R9217 gnd.n4236 gnd.n3373 19.3944
R9218 gnd.n4271 gnd.n3373 19.3944
R9219 gnd.n4271 gnd.n3371 19.3944
R9220 gnd.n4277 gnd.n3371 19.3944
R9221 gnd.n4277 gnd.n4276 19.3944
R9222 gnd.n4276 gnd.n3346 19.3944
R9223 gnd.n4320 gnd.n3346 19.3944
R9224 gnd.n4320 gnd.n3344 19.3944
R9225 gnd.n4326 gnd.n3344 19.3944
R9226 gnd.n4326 gnd.n4325 19.3944
R9227 gnd.n4325 gnd.n1906 19.3944
R9228 gnd.n4615 gnd.n1906 19.3944
R9229 gnd.n4615 gnd.n1904 19.3944
R9230 gnd.n4623 gnd.n1904 19.3944
R9231 gnd.n4623 gnd.n4622 19.3944
R9232 gnd.n4622 gnd.n4621 19.3944
R9233 gnd.n4724 gnd.n4723 19.3944
R9234 gnd.n4723 gnd.n1845 19.3944
R9235 gnd.n4719 gnd.n1845 19.3944
R9236 gnd.n4719 gnd.n4716 19.3944
R9237 gnd.n4716 gnd.n4713 19.3944
R9238 gnd.n4713 gnd.n4712 19.3944
R9239 gnd.n4712 gnd.n4709 19.3944
R9240 gnd.n4709 gnd.n4708 19.3944
R9241 gnd.n4708 gnd.n4705 19.3944
R9242 gnd.n4705 gnd.n4704 19.3944
R9243 gnd.n4704 gnd.n4701 19.3944
R9244 gnd.n4701 gnd.n4700 19.3944
R9245 gnd.n4700 gnd.n4697 19.3944
R9246 gnd.n4697 gnd.n4696 19.3944
R9247 gnd.n3880 gnd.n3779 19.3944
R9248 gnd.n3880 gnd.n3770 19.3944
R9249 gnd.n3893 gnd.n3770 19.3944
R9250 gnd.n3893 gnd.n3768 19.3944
R9251 gnd.n3897 gnd.n3768 19.3944
R9252 gnd.n3897 gnd.n3758 19.3944
R9253 gnd.n3909 gnd.n3758 19.3944
R9254 gnd.n3909 gnd.n3756 19.3944
R9255 gnd.n3943 gnd.n3756 19.3944
R9256 gnd.n3943 gnd.n3942 19.3944
R9257 gnd.n3942 gnd.n3941 19.3944
R9258 gnd.n3941 gnd.n3940 19.3944
R9259 gnd.n3940 gnd.n3937 19.3944
R9260 gnd.n3937 gnd.n3936 19.3944
R9261 gnd.n3936 gnd.n3935 19.3944
R9262 gnd.n3935 gnd.n3933 19.3944
R9263 gnd.n3933 gnd.n3932 19.3944
R9264 gnd.n3932 gnd.n3929 19.3944
R9265 gnd.n3929 gnd.n3928 19.3944
R9266 gnd.n3928 gnd.n3927 19.3944
R9267 gnd.n3927 gnd.n3925 19.3944
R9268 gnd.n3925 gnd.n3624 19.3944
R9269 gnd.n4040 gnd.n3624 19.3944
R9270 gnd.n4040 gnd.n3622 19.3944
R9271 gnd.n4046 gnd.n3622 19.3944
R9272 gnd.n4046 gnd.n4045 19.3944
R9273 gnd.n4045 gnd.n3546 19.3944
R9274 gnd.n4120 gnd.n3546 19.3944
R9275 gnd.n4120 gnd.n3547 19.3944
R9276 gnd.n3594 gnd.n3593 19.3944
R9277 gnd.n3597 gnd.n3596 19.3944
R9278 gnd.n3584 gnd.n3583 19.3944
R9279 gnd.n4139 gnd.n3460 19.3944
R9280 gnd.n4139 gnd.n4138 19.3944
R9281 gnd.n4138 gnd.n4137 19.3944
R9282 gnd.n4137 gnd.n4135 19.3944
R9283 gnd.n4135 gnd.n4134 19.3944
R9284 gnd.n4134 gnd.n4132 19.3944
R9285 gnd.n4132 gnd.n4131 19.3944
R9286 gnd.n4131 gnd.n3409 19.3944
R9287 gnd.n4207 gnd.n3409 19.3944
R9288 gnd.n4207 gnd.n3407 19.3944
R9289 gnd.n4226 gnd.n3407 19.3944
R9290 gnd.n4226 gnd.n4225 19.3944
R9291 gnd.n4225 gnd.n4224 19.3944
R9292 gnd.n4224 gnd.n4222 19.3944
R9293 gnd.n4222 gnd.n4221 19.3944
R9294 gnd.n4221 gnd.n4219 19.3944
R9295 gnd.n4219 gnd.n4218 19.3944
R9296 gnd.n4218 gnd.n3353 19.3944
R9297 gnd.n4292 gnd.n3353 19.3944
R9298 gnd.n4292 gnd.n3351 19.3944
R9299 gnd.n4315 gnd.n3351 19.3944
R9300 gnd.n4315 gnd.n4314 19.3944
R9301 gnd.n4314 gnd.n4313 19.3944
R9302 gnd.n4313 gnd.n4310 19.3944
R9303 gnd.n4310 gnd.n4309 19.3944
R9304 gnd.n4309 gnd.n4307 19.3944
R9305 gnd.n4307 gnd.n4306 19.3944
R9306 gnd.n4306 gnd.n4304 19.3944
R9307 gnd.n4304 gnd.n1892 19.3944
R9308 gnd.n3885 gnd.n3775 19.3944
R9309 gnd.n3885 gnd.n3773 19.3944
R9310 gnd.n3889 gnd.n3773 19.3944
R9311 gnd.n3889 gnd.n3764 19.3944
R9312 gnd.n3901 gnd.n3764 19.3944
R9313 gnd.n3901 gnd.n3762 19.3944
R9314 gnd.n3905 gnd.n3762 19.3944
R9315 gnd.n3905 gnd.n3751 19.3944
R9316 gnd.n3947 gnd.n3751 19.3944
R9317 gnd.n3947 gnd.n3705 19.3944
R9318 gnd.n3953 gnd.n3705 19.3944
R9319 gnd.n3953 gnd.n3952 19.3944
R9320 gnd.n3952 gnd.n3683 19.3944
R9321 gnd.n3974 gnd.n3683 19.3944
R9322 gnd.n3974 gnd.n3676 19.3944
R9323 gnd.n3985 gnd.n3676 19.3944
R9324 gnd.n3985 gnd.n3984 19.3944
R9325 gnd.n3984 gnd.n3657 19.3944
R9326 gnd.n4005 gnd.n3657 19.3944
R9327 gnd.n4005 gnd.n3647 19.3944
R9328 gnd.n4015 gnd.n3647 19.3944
R9329 gnd.n4015 gnd.n3630 19.3944
R9330 gnd.n4036 gnd.n3630 19.3944
R9331 gnd.n4036 gnd.n4035 19.3944
R9332 gnd.n4035 gnd.n3609 19.3944
R9333 gnd.n4066 gnd.n3609 19.3944
R9334 gnd.n4066 gnd.n3554 19.3944
R9335 gnd.n4116 gnd.n3554 19.3944
R9336 gnd.n4116 gnd.n4115 19.3944
R9337 gnd.n4115 gnd.n4114 19.3944
R9338 gnd.n4114 gnd.n3558 19.3944
R9339 gnd.n3576 gnd.n3558 19.3944
R9340 gnd.n4102 gnd.n3576 19.3944
R9341 gnd.n4102 gnd.n4101 19.3944
R9342 gnd.n4101 gnd.n4100 19.3944
R9343 gnd.n4100 gnd.n3580 19.3944
R9344 gnd.n3580 gnd.n3447 19.3944
R9345 gnd.n4157 gnd.n3447 19.3944
R9346 gnd.n4157 gnd.n3440 19.3944
R9347 gnd.n4168 gnd.n3440 19.3944
R9348 gnd.n4168 gnd.n3436 19.3944
R9349 gnd.n4181 gnd.n3436 19.3944
R9350 gnd.n4181 gnd.n4180 19.3944
R9351 gnd.n4180 gnd.n3415 19.3944
R9352 gnd.n4203 gnd.n3415 19.3944
R9353 gnd.n4203 gnd.n4202 19.3944
R9354 gnd.n4202 gnd.n3392 19.3944
R9355 gnd.n4242 gnd.n3392 19.3944
R9356 gnd.n4242 gnd.n3385 19.3944
R9357 gnd.n4253 gnd.n3385 19.3944
R9358 gnd.n4253 gnd.n3381 19.3944
R9359 gnd.n4266 gnd.n3381 19.3944
R9360 gnd.n4266 gnd.n4265 19.3944
R9361 gnd.n4265 gnd.n3360 19.3944
R9362 gnd.n4288 gnd.n3360 19.3944
R9363 gnd.n4288 gnd.n4287 19.3944
R9364 gnd.n4287 gnd.n3338 19.3944
R9365 gnd.n4331 gnd.n3338 19.3944
R9366 gnd.n4331 gnd.n3331 19.3944
R9367 gnd.n4342 gnd.n3331 19.3944
R9368 gnd.n4342 gnd.n3327 19.3944
R9369 gnd.n4609 gnd.n3327 19.3944
R9370 gnd.n4609 gnd.n4608 19.3944
R9371 gnd.n4608 gnd.n1895 19.3944
R9372 gnd.n4633 gnd.n1895 19.3944
R9373 gnd.n5820 gnd.n5819 19.3944
R9374 gnd.n5819 gnd.n5702 19.3944
R9375 gnd.n5812 gnd.n5702 19.3944
R9376 gnd.n5812 gnd.n5811 19.3944
R9377 gnd.n5811 gnd.n5716 19.3944
R9378 gnd.n5804 gnd.n5716 19.3944
R9379 gnd.n5804 gnd.n5803 19.3944
R9380 gnd.n5803 gnd.n5728 19.3944
R9381 gnd.n5796 gnd.n5728 19.3944
R9382 gnd.n5796 gnd.n5795 19.3944
R9383 gnd.n5795 gnd.n5739 19.3944
R9384 gnd.n5788 gnd.n5739 19.3944
R9385 gnd.n5788 gnd.n5787 19.3944
R9386 gnd.n5787 gnd.n5751 19.3944
R9387 gnd.n5780 gnd.n5751 19.3944
R9388 gnd.n5780 gnd.n5779 19.3944
R9389 gnd.n2770 gnd.n2769 19.3944
R9390 gnd.n2769 gnd.n2436 19.3944
R9391 gnd.n2765 gnd.n2436 19.3944
R9392 gnd.n2765 gnd.n2438 19.3944
R9393 gnd.n2759 gnd.n2438 19.3944
R9394 gnd.n2759 gnd.n2758 19.3944
R9395 gnd.n2758 gnd.n2757 19.3944
R9396 gnd.n2757 gnd.n2447 19.3944
R9397 gnd.n2751 gnd.n2447 19.3944
R9398 gnd.n2751 gnd.n2750 19.3944
R9399 gnd.n2750 gnd.n2749 19.3944
R9400 gnd.n2749 gnd.n2455 19.3944
R9401 gnd.n2743 gnd.n2455 19.3944
R9402 gnd.n2743 gnd.n2742 19.3944
R9403 gnd.n2742 gnd.n2741 19.3944
R9404 gnd.n2741 gnd.n2463 19.3944
R9405 gnd.n2735 gnd.n2463 19.3944
R9406 gnd.n2735 gnd.n2734 19.3944
R9407 gnd.n2734 gnd.n2733 19.3944
R9408 gnd.n2733 gnd.n2471 19.3944
R9409 gnd.n2727 gnd.n2471 19.3944
R9410 gnd.n2727 gnd.n2726 19.3944
R9411 gnd.n2726 gnd.n2725 19.3944
R9412 gnd.n2725 gnd.n2479 19.3944
R9413 gnd.n2719 gnd.n2479 19.3944
R9414 gnd.n2719 gnd.n2718 19.3944
R9415 gnd.n2718 gnd.n2717 19.3944
R9416 gnd.n2717 gnd.n2487 19.3944
R9417 gnd.n2711 gnd.n2487 19.3944
R9418 gnd.n2711 gnd.n2710 19.3944
R9419 gnd.n2710 gnd.n2709 19.3944
R9420 gnd.n2709 gnd.n2495 19.3944
R9421 gnd.n2703 gnd.n2495 19.3944
R9422 gnd.n2703 gnd.n2702 19.3944
R9423 gnd.n2702 gnd.n2701 19.3944
R9424 gnd.n2701 gnd.n2503 19.3944
R9425 gnd.n2695 gnd.n2503 19.3944
R9426 gnd.n2695 gnd.n2694 19.3944
R9427 gnd.n2694 gnd.n2693 19.3944
R9428 gnd.n2693 gnd.n2511 19.3944
R9429 gnd.n2687 gnd.n2511 19.3944
R9430 gnd.n2687 gnd.n2686 19.3944
R9431 gnd.n2686 gnd.n2685 19.3944
R9432 gnd.n2685 gnd.n2519 19.3944
R9433 gnd.n2679 gnd.n2519 19.3944
R9434 gnd.n2679 gnd.n2678 19.3944
R9435 gnd.n2678 gnd.n2677 19.3944
R9436 gnd.n2677 gnd.n2527 19.3944
R9437 gnd.n2671 gnd.n2527 19.3944
R9438 gnd.n2671 gnd.n2670 19.3944
R9439 gnd.n2670 gnd.n2669 19.3944
R9440 gnd.n2669 gnd.n2535 19.3944
R9441 gnd.n2663 gnd.n2535 19.3944
R9442 gnd.n2663 gnd.n2662 19.3944
R9443 gnd.n2662 gnd.n2661 19.3944
R9444 gnd.n2661 gnd.n2543 19.3944
R9445 gnd.n2655 gnd.n2543 19.3944
R9446 gnd.n2655 gnd.n2654 19.3944
R9447 gnd.n2654 gnd.n2653 19.3944
R9448 gnd.n2653 gnd.n2551 19.3944
R9449 gnd.n2647 gnd.n2551 19.3944
R9450 gnd.n2647 gnd.n2646 19.3944
R9451 gnd.n2646 gnd.n2645 19.3944
R9452 gnd.n2645 gnd.n2559 19.3944
R9453 gnd.n2639 gnd.n2559 19.3944
R9454 gnd.n2639 gnd.n2638 19.3944
R9455 gnd.n2638 gnd.n2637 19.3944
R9456 gnd.n2637 gnd.n2567 19.3944
R9457 gnd.n2631 gnd.n2567 19.3944
R9458 gnd.n2631 gnd.n2630 19.3944
R9459 gnd.n2630 gnd.n2629 19.3944
R9460 gnd.n2629 gnd.n2575 19.3944
R9461 gnd.n2623 gnd.n2575 19.3944
R9462 gnd.n2623 gnd.n2622 19.3944
R9463 gnd.n2622 gnd.n2621 19.3944
R9464 gnd.n2621 gnd.n2583 19.3944
R9465 gnd.n2615 gnd.n2583 19.3944
R9466 gnd.n2615 gnd.n2614 19.3944
R9467 gnd.n2614 gnd.n2613 19.3944
R9468 gnd.n2613 gnd.n2591 19.3944
R9469 gnd.n2607 gnd.n2591 19.3944
R9470 gnd.n2607 gnd.n2606 19.3944
R9471 gnd.n2606 gnd.n2605 19.3944
R9472 gnd.n2605 gnd.n2600 19.3944
R9473 gnd.n3108 gnd.n2101 19.3944
R9474 gnd.n3104 gnd.n2101 19.3944
R9475 gnd.n3104 gnd.n2103 19.3944
R9476 gnd.n3098 gnd.n2103 19.3944
R9477 gnd.n3098 gnd.n3097 19.3944
R9478 gnd.n3097 gnd.n3096 19.3944
R9479 gnd.n3096 gnd.n2110 19.3944
R9480 gnd.n3090 gnd.n2110 19.3944
R9481 gnd.n3090 gnd.n3089 19.3944
R9482 gnd.n3089 gnd.n3088 19.3944
R9483 gnd.n3088 gnd.n2118 19.3944
R9484 gnd.n3082 gnd.n2118 19.3944
R9485 gnd.n3082 gnd.n3081 19.3944
R9486 gnd.n3081 gnd.n3080 19.3944
R9487 gnd.n3080 gnd.n2126 19.3944
R9488 gnd.n3074 gnd.n2126 19.3944
R9489 gnd.n3074 gnd.n3073 19.3944
R9490 gnd.n3073 gnd.n3072 19.3944
R9491 gnd.n3072 gnd.n2134 19.3944
R9492 gnd.n3066 gnd.n2134 19.3944
R9493 gnd.n3066 gnd.n3065 19.3944
R9494 gnd.n3065 gnd.n3064 19.3944
R9495 gnd.n3064 gnd.n2142 19.3944
R9496 gnd.n3058 gnd.n2142 19.3944
R9497 gnd.n3058 gnd.n3057 19.3944
R9498 gnd.n3057 gnd.n3056 19.3944
R9499 gnd.n3056 gnd.n2150 19.3944
R9500 gnd.n3050 gnd.n2150 19.3944
R9501 gnd.n3050 gnd.n3049 19.3944
R9502 gnd.n3049 gnd.n3048 19.3944
R9503 gnd.n3048 gnd.n2158 19.3944
R9504 gnd.n3042 gnd.n2158 19.3944
R9505 gnd.n3042 gnd.n3041 19.3944
R9506 gnd.n3041 gnd.n3040 19.3944
R9507 gnd.n3040 gnd.n2166 19.3944
R9508 gnd.n3034 gnd.n2166 19.3944
R9509 gnd.n3034 gnd.n3033 19.3944
R9510 gnd.n3033 gnd.n3032 19.3944
R9511 gnd.n3032 gnd.n2174 19.3944
R9512 gnd.n3026 gnd.n2174 19.3944
R9513 gnd.n3026 gnd.n3025 19.3944
R9514 gnd.n3025 gnd.n3024 19.3944
R9515 gnd.n3024 gnd.n2182 19.3944
R9516 gnd.n3018 gnd.n2182 19.3944
R9517 gnd.n3018 gnd.n3017 19.3944
R9518 gnd.n3017 gnd.n3016 19.3944
R9519 gnd.n3016 gnd.n2190 19.3944
R9520 gnd.n3010 gnd.n2190 19.3944
R9521 gnd.n3010 gnd.n3009 19.3944
R9522 gnd.n3009 gnd.n3008 19.3944
R9523 gnd.n3008 gnd.n2198 19.3944
R9524 gnd.n3002 gnd.n2198 19.3944
R9525 gnd.n3002 gnd.n3001 19.3944
R9526 gnd.n3001 gnd.n3000 19.3944
R9527 gnd.n3000 gnd.n2206 19.3944
R9528 gnd.n2994 gnd.n2206 19.3944
R9529 gnd.n2994 gnd.n2993 19.3944
R9530 gnd.n2993 gnd.n2992 19.3944
R9531 gnd.n2992 gnd.n2214 19.3944
R9532 gnd.n2986 gnd.n2214 19.3944
R9533 gnd.n2986 gnd.n2985 19.3944
R9534 gnd.n2985 gnd.n2984 19.3944
R9535 gnd.n2984 gnd.n2222 19.3944
R9536 gnd.n2978 gnd.n2222 19.3944
R9537 gnd.n2978 gnd.n2977 19.3944
R9538 gnd.n2977 gnd.n2976 19.3944
R9539 gnd.n2976 gnd.n2230 19.3944
R9540 gnd.n2970 gnd.n2230 19.3944
R9541 gnd.n2970 gnd.n2969 19.3944
R9542 gnd.n2969 gnd.n2968 19.3944
R9543 gnd.n2968 gnd.n2238 19.3944
R9544 gnd.n2962 gnd.n2238 19.3944
R9545 gnd.n2962 gnd.n2961 19.3944
R9546 gnd.n2961 gnd.n2960 19.3944
R9547 gnd.n2960 gnd.n2246 19.3944
R9548 gnd.n2954 gnd.n2246 19.3944
R9549 gnd.n2954 gnd.n2953 19.3944
R9550 gnd.n2953 gnd.n2952 19.3944
R9551 gnd.n2952 gnd.n2254 19.3944
R9552 gnd.n2946 gnd.n2254 19.3944
R9553 gnd.n2946 gnd.n2945 19.3944
R9554 gnd.n2945 gnd.n2944 19.3944
R9555 gnd.n2944 gnd.n2262 19.3944
R9556 gnd.n2938 gnd.n2262 19.3944
R9557 gnd.n2938 gnd.n2937 19.3944
R9558 gnd.n2937 gnd.n2936 19.3944
R9559 gnd.n2936 gnd.n2270 19.3944
R9560 gnd.n2930 gnd.n2270 19.3944
R9561 gnd.n2930 gnd.n2929 19.3944
R9562 gnd.n2929 gnd.n2928 19.3944
R9563 gnd.n2928 gnd.n2278 19.3944
R9564 gnd.n2922 gnd.n2278 19.3944
R9565 gnd.n2922 gnd.n2921 19.3944
R9566 gnd.n2921 gnd.n2920 19.3944
R9567 gnd.n2920 gnd.n2286 19.3944
R9568 gnd.n2914 gnd.n2286 19.3944
R9569 gnd.n2914 gnd.n2913 19.3944
R9570 gnd.n2913 gnd.n2912 19.3944
R9571 gnd.n2912 gnd.n2294 19.3944
R9572 gnd.n2906 gnd.n2294 19.3944
R9573 gnd.n2906 gnd.n2905 19.3944
R9574 gnd.n2905 gnd.n2904 19.3944
R9575 gnd.n2904 gnd.n2302 19.3944
R9576 gnd.n2898 gnd.n2302 19.3944
R9577 gnd.n2898 gnd.n2897 19.3944
R9578 gnd.n2897 gnd.n2896 19.3944
R9579 gnd.n2896 gnd.n2310 19.3944
R9580 gnd.n2890 gnd.n2310 19.3944
R9581 gnd.n2890 gnd.n2889 19.3944
R9582 gnd.n2889 gnd.n2888 19.3944
R9583 gnd.n2888 gnd.n2318 19.3944
R9584 gnd.n2882 gnd.n2318 19.3944
R9585 gnd.n2882 gnd.n2881 19.3944
R9586 gnd.n2881 gnd.n2880 19.3944
R9587 gnd.n2880 gnd.n2326 19.3944
R9588 gnd.n2874 gnd.n2326 19.3944
R9589 gnd.n2874 gnd.n2873 19.3944
R9590 gnd.n2873 gnd.n2872 19.3944
R9591 gnd.n2872 gnd.n2334 19.3944
R9592 gnd.n2866 gnd.n2334 19.3944
R9593 gnd.n2866 gnd.n2865 19.3944
R9594 gnd.n2865 gnd.n2864 19.3944
R9595 gnd.n2864 gnd.n2342 19.3944
R9596 gnd.n2858 gnd.n2342 19.3944
R9597 gnd.n2858 gnd.n2857 19.3944
R9598 gnd.n2857 gnd.n2856 19.3944
R9599 gnd.n2856 gnd.n2350 19.3944
R9600 gnd.n2850 gnd.n2350 19.3944
R9601 gnd.n2850 gnd.n2849 19.3944
R9602 gnd.n2849 gnd.n2848 19.3944
R9603 gnd.n2848 gnd.n2358 19.3944
R9604 gnd.n2842 gnd.n2358 19.3944
R9605 gnd.n2842 gnd.n2841 19.3944
R9606 gnd.n2841 gnd.n2840 19.3944
R9607 gnd.n2840 gnd.n2366 19.3944
R9608 gnd.n2834 gnd.n2366 19.3944
R9609 gnd.n2834 gnd.n2833 19.3944
R9610 gnd.n2833 gnd.n2832 19.3944
R9611 gnd.n2832 gnd.n2374 19.3944
R9612 gnd.n2826 gnd.n2374 19.3944
R9613 gnd.n2826 gnd.n2825 19.3944
R9614 gnd.n2825 gnd.n2824 19.3944
R9615 gnd.n2824 gnd.n2382 19.3944
R9616 gnd.n2818 gnd.n2382 19.3944
R9617 gnd.n2818 gnd.n2817 19.3944
R9618 gnd.n2817 gnd.n2816 19.3944
R9619 gnd.n2816 gnd.n2390 19.3944
R9620 gnd.n2810 gnd.n2390 19.3944
R9621 gnd.n2810 gnd.n2809 19.3944
R9622 gnd.n2809 gnd.n2808 19.3944
R9623 gnd.n2808 gnd.n2398 19.3944
R9624 gnd.n2802 gnd.n2398 19.3944
R9625 gnd.n2802 gnd.n2801 19.3944
R9626 gnd.n2801 gnd.n2800 19.3944
R9627 gnd.n2800 gnd.n2406 19.3944
R9628 gnd.n2794 gnd.n2406 19.3944
R9629 gnd.n2794 gnd.n2793 19.3944
R9630 gnd.n2793 gnd.n2792 19.3944
R9631 gnd.n2792 gnd.n2414 19.3944
R9632 gnd.n2786 gnd.n2414 19.3944
R9633 gnd.n2786 gnd.n2785 19.3944
R9634 gnd.n2785 gnd.n2784 19.3944
R9635 gnd.n2784 gnd.n2422 19.3944
R9636 gnd.n2778 gnd.n2422 19.3944
R9637 gnd.n2778 gnd.n2777 19.3944
R9638 gnd.n2777 gnd.n2776 19.3944
R9639 gnd.n2776 gnd.n2430 19.3944
R9640 gnd.n7038 gnd.n629 19.3944
R9641 gnd.n7038 gnd.n7037 19.3944
R9642 gnd.n7037 gnd.n7036 19.3944
R9643 gnd.n7036 gnd.n7034 19.3944
R9644 gnd.n7034 gnd.n7031 19.3944
R9645 gnd.n7031 gnd.n7030 19.3944
R9646 gnd.n7030 gnd.n7027 19.3944
R9647 gnd.n7027 gnd.n7026 19.3944
R9648 gnd.n7026 gnd.n7023 19.3944
R9649 gnd.n7023 gnd.n7022 19.3944
R9650 gnd.n7022 gnd.n7019 19.3944
R9651 gnd.n7019 gnd.n7018 19.3944
R9652 gnd.n7018 gnd.n7015 19.3944
R9653 gnd.n7015 gnd.n7014 19.3944
R9654 gnd.n7014 gnd.n7011 19.3944
R9655 gnd.n7011 gnd.n7010 19.3944
R9656 gnd.n7010 gnd.n7007 19.3944
R9657 gnd.n7005 gnd.n7002 19.3944
R9658 gnd.n7002 gnd.n7001 19.3944
R9659 gnd.n7001 gnd.n6998 19.3944
R9660 gnd.n6998 gnd.n6997 19.3944
R9661 gnd.n6997 gnd.n6994 19.3944
R9662 gnd.n6994 gnd.n6993 19.3944
R9663 gnd.n6993 gnd.n6990 19.3944
R9664 gnd.n6988 gnd.n6985 19.3944
R9665 gnd.n6985 gnd.n6984 19.3944
R9666 gnd.n6984 gnd.n6981 19.3944
R9667 gnd.n6981 gnd.n6980 19.3944
R9668 gnd.n6980 gnd.n6977 19.3944
R9669 gnd.n6977 gnd.n6976 19.3944
R9670 gnd.n6976 gnd.n6973 19.3944
R9671 gnd.n6973 gnd.n6972 19.3944
R9672 gnd.n6968 gnd.n6965 19.3944
R9673 gnd.n6965 gnd.n6964 19.3944
R9674 gnd.n6964 gnd.n6961 19.3944
R9675 gnd.n6961 gnd.n6960 19.3944
R9676 gnd.n6960 gnd.n6957 19.3944
R9677 gnd.n6957 gnd.n6956 19.3944
R9678 gnd.n6956 gnd.n6953 19.3944
R9679 gnd.n6953 gnd.n6952 19.3944
R9680 gnd.n6952 gnd.n6949 19.3944
R9681 gnd.n6949 gnd.n6948 19.3944
R9682 gnd.n6948 gnd.n6945 19.3944
R9683 gnd.n6945 gnd.n6944 19.3944
R9684 gnd.n6944 gnd.n6941 19.3944
R9685 gnd.n6941 gnd.n6940 19.3944
R9686 gnd.n6940 gnd.n6937 19.3944
R9687 gnd.n6937 gnd.n6936 19.3944
R9688 gnd.n6936 gnd.n6933 19.3944
R9689 gnd.n6933 gnd.n6932 19.3944
R9690 gnd.n7063 gnd.n582 19.3944
R9691 gnd.n7063 gnd.n7062 19.3944
R9692 gnd.n7062 gnd.n551 19.3944
R9693 gnd.n7089 gnd.n551 19.3944
R9694 gnd.n7090 gnd.n7089 19.3944
R9695 gnd.n7097 gnd.n7090 19.3944
R9696 gnd.n7097 gnd.n7096 19.3944
R9697 gnd.n7096 gnd.n7095 19.3944
R9698 gnd.n7095 gnd.n7094 19.3944
R9699 gnd.n7094 gnd.n7092 19.3944
R9700 gnd.n7092 gnd.n507 19.3944
R9701 gnd.n7147 gnd.n507 19.3944
R9702 gnd.n7147 gnd.n7146 19.3944
R9703 gnd.n7146 gnd.n512 19.3944
R9704 gnd.n512 gnd.n511 19.3944
R9705 gnd.n511 gnd.n508 19.3944
R9706 gnd.n508 gnd.n447 19.3944
R9707 gnd.n7218 gnd.n447 19.3944
R9708 gnd.n7219 gnd.n7218 19.3944
R9709 gnd.n7221 gnd.n7219 19.3944
R9710 gnd.n7221 gnd.n420 19.3944
R9711 gnd.n7260 gnd.n420 19.3944
R9712 gnd.n7261 gnd.n7260 19.3944
R9713 gnd.n7264 gnd.n7261 19.3944
R9714 gnd.n7265 gnd.n7264 19.3944
R9715 gnd.n7265 gnd.n393 19.3944
R9716 gnd.n7301 gnd.n393 19.3944
R9717 gnd.n7302 gnd.n7301 19.3944
R9718 gnd.n7302 gnd.n376 19.3944
R9719 gnd.n7325 gnd.n376 19.3944
R9720 gnd.n7325 gnd.n365 19.3944
R9721 gnd.n7337 gnd.n365 19.3944
R9722 gnd.n7339 gnd.n7337 19.3944
R9723 gnd.n7339 gnd.n7338 19.3944
R9724 gnd.n7338 gnd.n353 19.3944
R9725 gnd.n7358 gnd.n353 19.3944
R9726 gnd.n7358 gnd.n349 19.3944
R9727 gnd.n7492 gnd.n349 19.3944
R9728 gnd.n7493 gnd.n7492 19.3944
R9729 gnd.n7496 gnd.n7493 19.3944
R9730 gnd.n7497 gnd.n7496 19.3944
R9731 gnd.n7499 gnd.n7497 19.3944
R9732 gnd.n7500 gnd.n7499 19.3944
R9733 gnd.n7503 gnd.n7500 19.3944
R9734 gnd.n7504 gnd.n7503 19.3944
R9735 gnd.n7506 gnd.n7504 19.3944
R9736 gnd.n7507 gnd.n7506 19.3944
R9737 gnd.n7510 gnd.n7507 19.3944
R9738 gnd.n7511 gnd.n7510 19.3944
R9739 gnd.n7513 gnd.n7511 19.3944
R9740 gnd.n7514 gnd.n7513 19.3944
R9741 gnd.n7517 gnd.n7514 19.3944
R9742 gnd.n7518 gnd.n7517 19.3944
R9743 gnd.n7520 gnd.n7518 19.3944
R9744 gnd.n7521 gnd.n7520 19.3944
R9745 gnd.n7524 gnd.n7521 19.3944
R9746 gnd.n7525 gnd.n7524 19.3944
R9747 gnd.n7527 gnd.n7525 19.3944
R9748 gnd.n7528 gnd.n7527 19.3944
R9749 gnd.n7531 gnd.n7528 19.3944
R9750 gnd.n7532 gnd.n7531 19.3944
R9751 gnd.n7534 gnd.n7532 19.3944
R9752 gnd.n7535 gnd.n7534 19.3944
R9753 gnd.n7538 gnd.n7535 19.3944
R9754 gnd.n7066 gnd.n7065 19.3944
R9755 gnd.n7065 gnd.n576 19.3944
R9756 gnd.n579 gnd.n576 19.3944
R9757 gnd.n579 gnd.n537 19.3944
R9758 gnd.n7116 gnd.n537 19.3944
R9759 gnd.n7116 gnd.n7115 19.3944
R9760 gnd.n7115 gnd.n7114 19.3944
R9761 gnd.n7114 gnd.n7113 19.3944
R9762 gnd.n7113 gnd.n502 19.3944
R9763 gnd.n7151 gnd.n502 19.3944
R9764 gnd.n7151 gnd.n7150 19.3944
R9765 gnd.n7150 gnd.n7149 19.3944
R9766 gnd.n7149 gnd.n472 19.3944
R9767 gnd.n7186 gnd.n472 19.3944
R9768 gnd.n7186 gnd.n7185 19.3944
R9769 gnd.n7185 gnd.n7184 19.3944
R9770 gnd.n7184 gnd.n7183 19.3944
R9771 gnd.n7183 gnd.n445 19.3944
R9772 gnd.n7226 gnd.n445 19.3944
R9773 gnd.n7226 gnd.n7225 19.3944
R9774 gnd.n7225 gnd.n7224 19.3944
R9775 gnd.n7224 gnd.n417 19.3944
R9776 gnd.n7273 gnd.n417 19.3944
R9777 gnd.n7273 gnd.n7272 19.3944
R9778 gnd.n7272 gnd.n7271 19.3944
R9779 gnd.n7271 gnd.n7270 19.3944
R9780 gnd.n7270 gnd.n391 19.3944
R9781 gnd.n7305 gnd.n391 19.3944
R9782 gnd.n7305 gnd.n7304 19.3944
R9783 gnd.n7304 gnd.n374 19.3944
R9784 gnd.n7328 gnd.n374 19.3944
R9785 gnd.n7328 gnd.n363 19.3944
R9786 gnd.n7341 gnd.n363 19.3944
R9787 gnd.n7341 gnd.n355 19.3944
R9788 gnd.n7355 gnd.n355 19.3944
R9789 gnd.n7355 gnd.n123 19.3944
R9790 gnd.n7744 gnd.n123 19.3944
R9791 gnd.n7744 gnd.n7743 19.3944
R9792 gnd.n7743 gnd.n7742 19.3944
R9793 gnd.n7742 gnd.n127 19.3944
R9794 gnd.n7732 gnd.n127 19.3944
R9795 gnd.n7732 gnd.n7731 19.3944
R9796 gnd.n7731 gnd.n7730 19.3944
R9797 gnd.n7730 gnd.n144 19.3944
R9798 gnd.n7720 gnd.n144 19.3944
R9799 gnd.n7720 gnd.n7719 19.3944
R9800 gnd.n7719 gnd.n7718 19.3944
R9801 gnd.n7718 gnd.n164 19.3944
R9802 gnd.n7708 gnd.n164 19.3944
R9803 gnd.n7708 gnd.n7707 19.3944
R9804 gnd.n7707 gnd.n7706 19.3944
R9805 gnd.n7706 gnd.n182 19.3944
R9806 gnd.n7696 gnd.n182 19.3944
R9807 gnd.n7696 gnd.n7695 19.3944
R9808 gnd.n7695 gnd.n7694 19.3944
R9809 gnd.n7694 gnd.n202 19.3944
R9810 gnd.n7684 gnd.n202 19.3944
R9811 gnd.n7684 gnd.n7683 19.3944
R9812 gnd.n7683 gnd.n7682 19.3944
R9813 gnd.n7682 gnd.n220 19.3944
R9814 gnd.n7672 gnd.n220 19.3944
R9815 gnd.n7672 gnd.n7671 19.3944
R9816 gnd.n7671 gnd.n7670 19.3944
R9817 gnd.n7670 gnd.n240 19.3944
R9818 gnd.n7581 gnd.n325 19.3944
R9819 gnd.n7581 gnd.n7578 19.3944
R9820 gnd.n7578 gnd.n7575 19.3944
R9821 gnd.n7575 gnd.n7574 19.3944
R9822 gnd.n7574 gnd.n7571 19.3944
R9823 gnd.n7571 gnd.n7570 19.3944
R9824 gnd.n7570 gnd.n7567 19.3944
R9825 gnd.n7567 gnd.n7566 19.3944
R9826 gnd.n7566 gnd.n7563 19.3944
R9827 gnd.n7563 gnd.n7562 19.3944
R9828 gnd.n7562 gnd.n7559 19.3944
R9829 gnd.n7559 gnd.n7558 19.3944
R9830 gnd.n7558 gnd.n7555 19.3944
R9831 gnd.n7555 gnd.n7554 19.3944
R9832 gnd.n7554 gnd.n7551 19.3944
R9833 gnd.n7551 gnd.n7550 19.3944
R9834 gnd.n7550 gnd.n7547 19.3944
R9835 gnd.n7547 gnd.n7546 19.3944
R9836 gnd.n7624 gnd.n7621 19.3944
R9837 gnd.n7621 gnd.n7620 19.3944
R9838 gnd.n7620 gnd.n7617 19.3944
R9839 gnd.n7617 gnd.n7616 19.3944
R9840 gnd.n7616 gnd.n7613 19.3944
R9841 gnd.n7613 gnd.n7612 19.3944
R9842 gnd.n7612 gnd.n7609 19.3944
R9843 gnd.n7609 gnd.n7608 19.3944
R9844 gnd.n7608 gnd.n7605 19.3944
R9845 gnd.n7605 gnd.n7604 19.3944
R9846 gnd.n7604 gnd.n7601 19.3944
R9847 gnd.n7601 gnd.n7600 19.3944
R9848 gnd.n7600 gnd.n7597 19.3944
R9849 gnd.n7597 gnd.n7596 19.3944
R9850 gnd.n7596 gnd.n7593 19.3944
R9851 gnd.n7593 gnd.n7592 19.3944
R9852 gnd.n7592 gnd.n7589 19.3944
R9853 gnd.n7589 gnd.n7588 19.3944
R9854 gnd.n7662 gnd.n249 19.3944
R9855 gnd.n7657 gnd.n249 19.3944
R9856 gnd.n7657 gnd.n7656 19.3944
R9857 gnd.n7656 gnd.n7655 19.3944
R9858 gnd.n7655 gnd.n7652 19.3944
R9859 gnd.n7652 gnd.n7651 19.3944
R9860 gnd.n7651 gnd.n7648 19.3944
R9861 gnd.n7648 gnd.n7647 19.3944
R9862 gnd.n7647 gnd.n7644 19.3944
R9863 gnd.n7644 gnd.n7643 19.3944
R9864 gnd.n7643 gnd.n7640 19.3944
R9865 gnd.n7640 gnd.n7639 19.3944
R9866 gnd.n7639 gnd.n7636 19.3944
R9867 gnd.n7636 gnd.n7635 19.3944
R9868 gnd.n7635 gnd.n7632 19.3944
R9869 gnd.n7632 gnd.n7631 19.3944
R9870 gnd.n7631 gnd.n7628 19.3944
R9871 gnd.n7404 gnd.n7402 19.3944
R9872 gnd.n7407 gnd.n7404 19.3944
R9873 gnd.n7410 gnd.n7407 19.3944
R9874 gnd.n7413 gnd.n7410 19.3944
R9875 gnd.n7413 gnd.n7400 19.3944
R9876 gnd.n7417 gnd.n7400 19.3944
R9877 gnd.n7420 gnd.n7417 19.3944
R9878 gnd.n7423 gnd.n7420 19.3944
R9879 gnd.n7423 gnd.n7398 19.3944
R9880 gnd.n7427 gnd.n7398 19.3944
R9881 gnd.n7430 gnd.n7427 19.3944
R9882 gnd.n7433 gnd.n7430 19.3944
R9883 gnd.n7433 gnd.n7396 19.3944
R9884 gnd.n7437 gnd.n7396 19.3944
R9885 gnd.n7440 gnd.n7437 19.3944
R9886 gnd.n7443 gnd.n7440 19.3944
R9887 gnd.n6866 gnd.n559 19.3944
R9888 gnd.n7080 gnd.n559 19.3944
R9889 gnd.n7080 gnd.n556 19.3944
R9890 gnd.n7085 gnd.n556 19.3944
R9891 gnd.n7085 gnd.n557 19.3944
R9892 gnd.n557 gnd.n519 19.3944
R9893 gnd.n7130 gnd.n519 19.3944
R9894 gnd.n7130 gnd.n516 19.3944
R9895 gnd.n7134 gnd.n516 19.3944
R9896 gnd.n7135 gnd.n7134 19.3944
R9897 gnd.n7137 gnd.n7135 19.3944
R9898 gnd.n7137 gnd.n513 19.3944
R9899 gnd.n7142 gnd.n513 19.3944
R9900 gnd.n7142 gnd.n514 19.3944
R9901 gnd.n514 gnd.n454 19.3944
R9902 gnd.n7200 gnd.n454 19.3944
R9903 gnd.n7200 gnd.n451 19.3944
R9904 gnd.n7214 gnd.n451 19.3944
R9905 gnd.n7214 gnd.n452 19.3944
R9906 gnd.n7210 gnd.n452 19.3944
R9907 gnd.n7210 gnd.n7209 19.3944
R9908 gnd.n7209 gnd.n7208 19.3944
R9909 gnd.n7208 gnd.n7205 19.3944
R9910 gnd.n7205 gnd.n400 19.3944
R9911 gnd.n7287 gnd.n400 19.3944
R9912 gnd.n7287 gnd.n397 19.3944
R9913 gnd.n7297 gnd.n397 19.3944
R9914 gnd.n7297 gnd.n398 19.3944
R9915 gnd.n7293 gnd.n398 19.3944
R9916 gnd.n7293 gnd.n7292 19.3944
R9917 gnd.n7292 gnd.n7291 19.3944
R9918 gnd.n7291 gnd.n96 19.3944
R9919 gnd.n7757 gnd.n96 19.3944
R9920 gnd.n7757 gnd.n7756 19.3944
R9921 gnd.n7756 gnd.n99 19.3944
R9922 gnd.n7362 gnd.n99 19.3944
R9923 gnd.n7362 gnd.n350 19.3944
R9924 gnd.n7488 gnd.n350 19.3944
R9925 gnd.n7488 gnd.n7487 19.3944
R9926 gnd.n7487 gnd.n7486 19.3944
R9927 gnd.n7486 gnd.n7484 19.3944
R9928 gnd.n7484 gnd.n7483 19.3944
R9929 gnd.n7483 gnd.n7481 19.3944
R9930 gnd.n7481 gnd.n7480 19.3944
R9931 gnd.n7480 gnd.n7478 19.3944
R9932 gnd.n7478 gnd.n7477 19.3944
R9933 gnd.n7477 gnd.n7475 19.3944
R9934 gnd.n7475 gnd.n7474 19.3944
R9935 gnd.n7474 gnd.n7472 19.3944
R9936 gnd.n7472 gnd.n7471 19.3944
R9937 gnd.n7471 gnd.n7469 19.3944
R9938 gnd.n7469 gnd.n7468 19.3944
R9939 gnd.n7468 gnd.n7466 19.3944
R9940 gnd.n7466 gnd.n7465 19.3944
R9941 gnd.n7465 gnd.n7463 19.3944
R9942 gnd.n7463 gnd.n7462 19.3944
R9943 gnd.n7462 gnd.n7460 19.3944
R9944 gnd.n7460 gnd.n7459 19.3944
R9945 gnd.n7459 gnd.n7457 19.3944
R9946 gnd.n7457 gnd.n7456 19.3944
R9947 gnd.n7456 gnd.n7454 19.3944
R9948 gnd.n7454 gnd.n7453 19.3944
R9949 gnd.n7453 gnd.n7451 19.3944
R9950 gnd.n7451 gnd.n7450 19.3944
R9951 gnd.n7070 gnd.n566 19.3944
R9952 gnd.n7076 gnd.n566 19.3944
R9953 gnd.n7076 gnd.n7075 19.3944
R9954 gnd.n7075 gnd.n529 19.3944
R9955 gnd.n7120 gnd.n529 19.3944
R9956 gnd.n7120 gnd.n527 19.3944
R9957 gnd.n7126 gnd.n527 19.3944
R9958 gnd.n7126 gnd.n7125 19.3944
R9959 gnd.n7125 gnd.n495 19.3944
R9960 gnd.n7155 gnd.n495 19.3944
R9961 gnd.n7155 gnd.n493 19.3944
R9962 gnd.n7159 gnd.n493 19.3944
R9963 gnd.n7159 gnd.n464 19.3944
R9964 gnd.n7190 gnd.n464 19.3944
R9965 gnd.n7190 gnd.n462 19.3944
R9966 gnd.n7196 gnd.n462 19.3944
R9967 gnd.n7196 gnd.n7195 19.3944
R9968 gnd.n7195 gnd.n437 19.3944
R9969 gnd.n7230 gnd.n437 19.3944
R9970 gnd.n7230 gnd.n435 19.3944
R9971 gnd.n7234 gnd.n435 19.3944
R9972 gnd.n7234 gnd.n410 19.3944
R9973 gnd.n7277 gnd.n410 19.3944
R9974 gnd.n7277 gnd.n408 19.3944
R9975 gnd.n7283 gnd.n408 19.3944
R9976 gnd.n7283 gnd.n7282 19.3944
R9977 gnd.n7282 gnd.n7281 19.3944
R9978 gnd.n7310 gnd.n7309 19.3944
R9979 gnd.n371 gnd.n370 19.3944
R9980 gnd.n7333 gnd.n7332 19.3944
R9981 gnd.n7752 gnd.n7751 19.3944
R9982 gnd.n7748 gnd.n107 19.3944
R9983 gnd.n7748 gnd.n114 19.3944
R9984 gnd.n7738 gnd.n114 19.3944
R9985 gnd.n7738 gnd.n7737 19.3944
R9986 gnd.n7737 gnd.n7736 19.3944
R9987 gnd.n7736 gnd.n136 19.3944
R9988 gnd.n7726 gnd.n136 19.3944
R9989 gnd.n7726 gnd.n7725 19.3944
R9990 gnd.n7725 gnd.n7724 19.3944
R9991 gnd.n7724 gnd.n154 19.3944
R9992 gnd.n7714 gnd.n154 19.3944
R9993 gnd.n7714 gnd.n7713 19.3944
R9994 gnd.n7713 gnd.n7712 19.3944
R9995 gnd.n7712 gnd.n174 19.3944
R9996 gnd.n7702 gnd.n174 19.3944
R9997 gnd.n7702 gnd.n7701 19.3944
R9998 gnd.n7701 gnd.n7700 19.3944
R9999 gnd.n7700 gnd.n192 19.3944
R10000 gnd.n7690 gnd.n192 19.3944
R10001 gnd.n7690 gnd.n7689 19.3944
R10002 gnd.n7689 gnd.n7688 19.3944
R10003 gnd.n7688 gnd.n212 19.3944
R10004 gnd.n7678 gnd.n212 19.3944
R10005 gnd.n7678 gnd.n7677 19.3944
R10006 gnd.n7677 gnd.n7676 19.3944
R10007 gnd.n7676 gnd.n231 19.3944
R10008 gnd.n7666 gnd.n231 19.3944
R10009 gnd.n7666 gnd.n7665 19.3944
R10010 gnd.n1971 gnd.n1970 19.3944
R10011 gnd.n1970 gnd.n1913 19.3944
R10012 gnd.n1966 gnd.n1965 19.3944
R10013 gnd.n1963 gnd.n1916 19.3944
R10014 gnd.n1959 gnd.n1958 19.3944
R10015 gnd.n1958 gnd.n1957 19.3944
R10016 gnd.n1957 gnd.n1920 19.3944
R10017 gnd.n1953 gnd.n1920 19.3944
R10018 gnd.n1953 gnd.n1952 19.3944
R10019 gnd.n1952 gnd.n1951 19.3944
R10020 gnd.n1951 gnd.n1926 19.3944
R10021 gnd.n1947 gnd.n1926 19.3944
R10022 gnd.n1947 gnd.n1946 19.3944
R10023 gnd.n1946 gnd.n1945 19.3944
R10024 gnd.n1945 gnd.n1932 19.3944
R10025 gnd.n1941 gnd.n1932 19.3944
R10026 gnd.n1941 gnd.n1940 19.3944
R10027 gnd.n1940 gnd.n1939 19.3944
R10028 gnd.n1939 gnd.n1549 19.3944
R10029 gnd.n1549 gnd.n1547 19.3944
R10030 gnd.n5391 gnd.n1547 19.3944
R10031 gnd.n5391 gnd.n1545 19.3944
R10032 gnd.n5400 gnd.n1545 19.3944
R10033 gnd.n5400 gnd.n5399 19.3944
R10034 gnd.n5399 gnd.n5398 19.3944
R10035 gnd.n5398 gnd.n1496 19.3944
R10036 gnd.n5455 gnd.n1496 19.3944
R10037 gnd.n5455 gnd.n1494 19.3944
R10038 gnd.n5459 gnd.n1494 19.3944
R10039 gnd.n5459 gnd.n1492 19.3944
R10040 gnd.n5463 gnd.n1492 19.3944
R10041 gnd.n5463 gnd.n1490 19.3944
R10042 gnd.n5695 gnd.n1490 19.3944
R10043 gnd.n5695 gnd.n5694 19.3944
R10044 gnd.n5694 gnd.n5693 19.3944
R10045 gnd.n5693 gnd.n5469 19.3944
R10046 gnd.n5687 gnd.n5469 19.3944
R10047 gnd.n5687 gnd.n5686 19.3944
R10048 gnd.n5686 gnd.n5685 19.3944
R10049 gnd.n5685 gnd.n5475 19.3944
R10050 gnd.n5548 gnd.n5475 19.3944
R10051 gnd.n5570 gnd.n5548 19.3944
R10052 gnd.n5570 gnd.n5545 19.3944
R10053 gnd.n5574 gnd.n5545 19.3944
R10054 gnd.n5574 gnd.n5535 19.3944
R10055 gnd.n5591 gnd.n5535 19.3944
R10056 gnd.n5591 gnd.n5533 19.3944
R10057 gnd.n5595 gnd.n5533 19.3944
R10058 gnd.n5595 gnd.n5523 19.3944
R10059 gnd.n5612 gnd.n5523 19.3944
R10060 gnd.n5612 gnd.n5521 19.3944
R10061 gnd.n5616 gnd.n5521 19.3944
R10062 gnd.n5616 gnd.n5510 19.3944
R10063 gnd.n5641 gnd.n5510 19.3944
R10064 gnd.n5641 gnd.n5508 19.3944
R10065 gnd.n5650 gnd.n5508 19.3944
R10066 gnd.n5650 gnd.n5649 19.3944
R10067 gnd.n5649 gnd.n5648 19.3944
R10068 gnd.n5648 gnd.n1198 19.3944
R10069 gnd.n6156 gnd.n1198 19.3944
R10070 gnd.n6156 gnd.n1196 19.3944
R10071 gnd.n6160 gnd.n1196 19.3944
R10072 gnd.n6160 gnd.n1172 19.3944
R10073 gnd.n6197 gnd.n1172 19.3944
R10074 gnd.n6197 gnd.n1170 19.3944
R10075 gnd.n6205 gnd.n1170 19.3944
R10076 gnd.n6205 gnd.n6204 19.3944
R10077 gnd.n6204 gnd.n6203 19.3944
R10078 gnd.n6203 gnd.n1150 19.3944
R10079 gnd.n6225 gnd.n1150 19.3944
R10080 gnd.n6225 gnd.n1148 19.3944
R10081 gnd.n6230 gnd.n1148 19.3944
R10082 gnd.n6230 gnd.n1120 19.3944
R10083 gnd.n6284 gnd.n1120 19.3944
R10084 gnd.n6284 gnd.n6283 19.3944
R10085 gnd.n6283 gnd.n6282 19.3944
R10086 gnd.n6282 gnd.n1088 19.3944
R10087 gnd.n6346 gnd.n1088 19.3944
R10088 gnd.n6346 gnd.n6345 19.3944
R10089 gnd.n6345 gnd.n6344 19.3944
R10090 gnd.n6344 gnd.n1061 19.3944
R10091 gnd.n6384 gnd.n1061 19.3944
R10092 gnd.n6384 gnd.n6383 19.3944
R10093 gnd.n6383 gnd.n6382 19.3944
R10094 gnd.n6382 gnd.n1031 19.3944
R10095 gnd.n6423 gnd.n1031 19.3944
R10096 gnd.n6423 gnd.n6422 19.3944
R10097 gnd.n6422 gnd.n6421 19.3944
R10098 gnd.n6421 gnd.n1037 19.3944
R10099 gnd.n1037 gnd.n985 19.3944
R10100 gnd.n6487 gnd.n985 19.3944
R10101 gnd.n6487 gnd.n6486 19.3944
R10102 gnd.n6486 gnd.n6485 19.3944
R10103 gnd.n6485 gnd.n990 19.3944
R10104 gnd.n990 gnd.n943 19.3944
R10105 gnd.n6541 gnd.n943 19.3944
R10106 gnd.n6541 gnd.n941 19.3944
R10107 gnd.n6545 gnd.n941 19.3944
R10108 gnd.n6545 gnd.n889 19.3944
R10109 gnd.n6717 gnd.n889 19.3944
R10110 gnd.n6717 gnd.n887 19.3944
R10111 gnd.n6723 gnd.n887 19.3944
R10112 gnd.n6723 gnd.n6722 19.3944
R10113 gnd.n6722 gnd.n865 19.3944
R10114 gnd.n6747 gnd.n865 19.3944
R10115 gnd.n6747 gnd.n863 19.3944
R10116 gnd.n6753 gnd.n863 19.3944
R10117 gnd.n6753 gnd.n6752 19.3944
R10118 gnd.n6752 gnd.n840 19.3944
R10119 gnd.n6777 gnd.n840 19.3944
R10120 gnd.n6777 gnd.n838 19.3944
R10121 gnd.n6783 gnd.n838 19.3944
R10122 gnd.n6783 gnd.n6782 19.3944
R10123 gnd.n6782 gnd.n815 19.3944
R10124 gnd.n6812 gnd.n815 19.3944
R10125 gnd.n6812 gnd.n813 19.3944
R10126 gnd.n6819 gnd.n813 19.3944
R10127 gnd.n6819 gnd.n6818 19.3944
R10128 gnd.n6818 gnd.n801 19.3944
R10129 gnd.n801 gnd.n799 19.3944
R10130 gnd.n6836 gnd.n799 19.3944
R10131 gnd.n6836 gnd.n797 19.3944
R10132 gnd.n6842 gnd.n797 19.3944
R10133 gnd.n6842 gnd.n6841 19.3944
R10134 gnd.n6841 gnd.n587 19.3944
R10135 gnd.n7045 gnd.n587 19.3944
R10136 gnd.n7045 gnd.n585 19.3944
R10137 gnd.n7057 gnd.n585 19.3944
R10138 gnd.n7057 gnd.n7056 19.3944
R10139 gnd.n7056 gnd.n7055 19.3944
R10140 gnd.n7055 gnd.n7052 19.3944
R10141 gnd.n7052 gnd.n549 19.3944
R10142 gnd.n7102 gnd.n549 19.3944
R10143 gnd.n7102 gnd.n547 19.3944
R10144 gnd.n7108 gnd.n547 19.3944
R10145 gnd.n7108 gnd.n7107 19.3944
R10146 gnd.n7107 gnd.n485 19.3944
R10147 gnd.n7164 gnd.n485 19.3944
R10148 gnd.n7164 gnd.n483 19.3944
R10149 gnd.n7168 gnd.n483 19.3944
R10150 gnd.n7168 gnd.n481 19.3944
R10151 gnd.n7172 gnd.n481 19.3944
R10152 gnd.n7172 gnd.n479 19.3944
R10153 gnd.n7178 gnd.n479 19.3944
R10154 gnd.n7178 gnd.n7177 19.3944
R10155 gnd.n7177 gnd.n429 19.3944
R10156 gnd.n7239 gnd.n429 19.3944
R10157 gnd.n7239 gnd.n427 19.3944
R10158 gnd.n7255 gnd.n427 19.3944
R10159 gnd.n7255 gnd.n7254 19.3944
R10160 gnd.n7254 gnd.n7253 19.3944
R10161 gnd.n7253 gnd.n7245 19.3944
R10162 gnd.n7249 gnd.n7245 19.3944
R10163 gnd.n7249 gnd.n7248 19.3944
R10164 gnd.n7316 gnd.n7315 19.3944
R10165 gnd.n7320 gnd.n7319 19.3944
R10166 gnd.n7346 gnd.n358 19.3944
R10167 gnd.n7350 gnd.n7348 19.3944
R10168 gnd.n4887 gnd.n4884 19.3944
R10169 gnd.n4887 gnd.n4883 19.3944
R10170 gnd.n4891 gnd.n4883 19.3944
R10171 gnd.n4891 gnd.n4881 19.3944
R10172 gnd.n4897 gnd.n4881 19.3944
R10173 gnd.n4897 gnd.n4879 19.3944
R10174 gnd.n4901 gnd.n4879 19.3944
R10175 gnd.n4901 gnd.n4877 19.3944
R10176 gnd.n4907 gnd.n4877 19.3944
R10177 gnd.n4907 gnd.n4875 19.3944
R10178 gnd.n4911 gnd.n4875 19.3944
R10179 gnd.n4911 gnd.n4873 19.3944
R10180 gnd.n4917 gnd.n4873 19.3944
R10181 gnd.n4917 gnd.n4871 19.3944
R10182 gnd.n4921 gnd.n4871 19.3944
R10183 gnd.n4921 gnd.n4866 19.3944
R10184 gnd.n4927 gnd.n4866 19.3944
R10185 gnd.n4931 gnd.n4864 19.3944
R10186 gnd.n4931 gnd.n4862 19.3944
R10187 gnd.n4937 gnd.n4862 19.3944
R10188 gnd.n4937 gnd.n4860 19.3944
R10189 gnd.n4941 gnd.n4860 19.3944
R10190 gnd.n4941 gnd.n4858 19.3944
R10191 gnd.n4947 gnd.n4858 19.3944
R10192 gnd.n4947 gnd.n4856 19.3944
R10193 gnd.n4951 gnd.n4856 19.3944
R10194 gnd.n4951 gnd.n4854 19.3944
R10195 gnd.n4957 gnd.n4854 19.3944
R10196 gnd.n4957 gnd.n4852 19.3944
R10197 gnd.n4961 gnd.n4852 19.3944
R10198 gnd.n4961 gnd.n4850 19.3944
R10199 gnd.n4967 gnd.n4850 19.3944
R10200 gnd.n4967 gnd.n4848 19.3944
R10201 gnd.n4971 gnd.n4848 19.3944
R10202 gnd.n4971 gnd.n4846 19.3944
R10203 gnd.n4983 gnd.n4844 19.3944
R10204 gnd.n4983 gnd.n4842 19.3944
R10205 gnd.n4989 gnd.n4842 19.3944
R10206 gnd.n4989 gnd.n4840 19.3944
R10207 gnd.n4993 gnd.n4840 19.3944
R10208 gnd.n4993 gnd.n4838 19.3944
R10209 gnd.n4999 gnd.n4838 19.3944
R10210 gnd.n4999 gnd.n4836 19.3944
R10211 gnd.n5003 gnd.n4836 19.3944
R10212 gnd.n5003 gnd.n4834 19.3944
R10213 gnd.n5009 gnd.n4834 19.3944
R10214 gnd.n5009 gnd.n4832 19.3944
R10215 gnd.n5013 gnd.n4832 19.3944
R10216 gnd.n5013 gnd.n4830 19.3944
R10217 gnd.n5019 gnd.n4830 19.3944
R10218 gnd.n5019 gnd.n4828 19.3944
R10219 gnd.n5024 gnd.n4828 19.3944
R10220 gnd.n5024 gnd.n4826 19.3944
R10221 gnd.n4820 gnd.n4819 19.3944
R10222 gnd.n4819 gnd.n4734 19.3944
R10223 gnd.n4813 gnd.n4734 19.3944
R10224 gnd.n4813 gnd.n4812 19.3944
R10225 gnd.n4812 gnd.n4811 19.3944
R10226 gnd.n4811 gnd.n4740 19.3944
R10227 gnd.n4805 gnd.n4740 19.3944
R10228 gnd.n4805 gnd.n4804 19.3944
R10229 gnd.n4804 gnd.n4803 19.3944
R10230 gnd.n4803 gnd.n4746 19.3944
R10231 gnd.n4797 gnd.n4746 19.3944
R10232 gnd.n4797 gnd.n4796 19.3944
R10233 gnd.n4796 gnd.n4795 19.3944
R10234 gnd.n4795 gnd.n4752 19.3944
R10235 gnd.n4789 gnd.n4752 19.3944
R10236 gnd.n4789 gnd.n4788 19.3944
R10237 gnd.n4779 gnd.n4778 19.3944
R10238 gnd.n4778 gnd.n4776 19.3944
R10239 gnd.n4776 gnd.n4775 19.3944
R10240 gnd.n4775 gnd.n4773 19.3944
R10241 gnd.n4773 gnd.n4772 19.3944
R10242 gnd.n4772 gnd.n4770 19.3944
R10243 gnd.n4770 gnd.n4769 19.3944
R10244 gnd.n4769 gnd.n4767 19.3944
R10245 gnd.n4767 gnd.n1773 19.3944
R10246 gnd.n5099 gnd.n1773 19.3944
R10247 gnd.n5099 gnd.n1771 19.3944
R10248 gnd.n5105 gnd.n1771 19.3944
R10249 gnd.n5105 gnd.n5104 19.3944
R10250 gnd.n5104 gnd.n1748 19.3944
R10251 gnd.n5134 gnd.n1748 19.3944
R10252 gnd.n5134 gnd.n1746 19.3944
R10253 gnd.n5140 gnd.n1746 19.3944
R10254 gnd.n5140 gnd.n5139 19.3944
R10255 gnd.n5139 gnd.n1723 19.3944
R10256 gnd.n5169 gnd.n1723 19.3944
R10257 gnd.n5169 gnd.n1721 19.3944
R10258 gnd.n5175 gnd.n1721 19.3944
R10259 gnd.n5175 gnd.n5174 19.3944
R10260 gnd.n5174 gnd.n1696 19.3944
R10261 gnd.n5206 gnd.n1696 19.3944
R10262 gnd.n5206 gnd.n1694 19.3944
R10263 gnd.n5212 gnd.n1694 19.3944
R10264 gnd.n5212 gnd.n5211 19.3944
R10265 gnd.n5211 gnd.n1677 19.3944
R10266 gnd.n5231 gnd.n1677 19.3944
R10267 gnd.n5231 gnd.n1675 19.3944
R10268 gnd.n5235 gnd.n1675 19.3944
R10269 gnd.n5235 gnd.n1650 19.3944
R10270 gnd.n5265 gnd.n1650 19.3944
R10271 gnd.n5265 gnd.n1647 19.3944
R10272 gnd.n5270 gnd.n1647 19.3944
R10273 gnd.n5270 gnd.n1648 19.3944
R10274 gnd.n1648 gnd.n1616 19.3944
R10275 gnd.n5301 gnd.n1616 19.3944
R10276 gnd.n5301 gnd.n1613 19.3944
R10277 gnd.n5306 gnd.n1613 19.3944
R10278 gnd.n5306 gnd.n1614 19.3944
R10279 gnd.n1614 gnd.n1587 19.3944
R10280 gnd.n5337 gnd.n1587 19.3944
R10281 gnd.n5337 gnd.n1584 19.3944
R10282 gnd.n5342 gnd.n1584 19.3944
R10283 gnd.n5342 gnd.n1585 19.3944
R10284 gnd.n1585 gnd.n1556 19.3944
R10285 gnd.n5379 gnd.n1556 19.3944
R10286 gnd.n5379 gnd.n1553 19.3944
R10287 gnd.n5384 gnd.n1553 19.3944
R10288 gnd.n5384 gnd.n1554 19.3944
R10289 gnd.n1554 gnd.n1521 19.3944
R10290 gnd.n5422 gnd.n1521 19.3944
R10291 gnd.n5422 gnd.n1518 19.3944
R10292 gnd.n5430 gnd.n1518 19.3944
R10293 gnd.n5430 gnd.n1519 19.3944
R10294 gnd.n5426 gnd.n1519 19.3944
R10295 gnd.n5426 gnd.n1448 19.3944
R10296 gnd.n5852 gnd.n1448 19.3944
R10297 gnd.n5852 gnd.n1449 19.3944
R10298 gnd.n5848 gnd.n1449 19.3944
R10299 gnd.n5848 gnd.n5847 19.3944
R10300 gnd.n5847 gnd.n5846 19.3944
R10301 gnd.n5038 gnd.n5037 19.3944
R10302 gnd.n5038 gnd.n1810 19.3944
R10303 gnd.n5054 gnd.n1810 19.3944
R10304 gnd.n5055 gnd.n5054 19.3944
R10305 gnd.n5056 gnd.n5055 19.3944
R10306 gnd.n5056 gnd.n1792 19.3944
R10307 gnd.n5074 gnd.n1792 19.3944
R10308 gnd.n5075 gnd.n5074 19.3944
R10309 gnd.n5077 gnd.n5075 19.3944
R10310 gnd.n5078 gnd.n5077 19.3944
R10311 gnd.n5078 gnd.n1766 19.3944
R10312 gnd.n5109 gnd.n1766 19.3944
R10313 gnd.n5110 gnd.n5109 19.3944
R10314 gnd.n5112 gnd.n5110 19.3944
R10315 gnd.n5113 gnd.n5112 19.3944
R10316 gnd.n5113 gnd.n1741 19.3944
R10317 gnd.n5144 gnd.n1741 19.3944
R10318 gnd.n5145 gnd.n5144 19.3944
R10319 gnd.n5147 gnd.n5145 19.3944
R10320 gnd.n5148 gnd.n5147 19.3944
R10321 gnd.n5148 gnd.n1716 19.3944
R10322 gnd.n5179 gnd.n1716 19.3944
R10323 gnd.n5180 gnd.n5179 19.3944
R10324 gnd.n5182 gnd.n5180 19.3944
R10325 gnd.n5183 gnd.n5182 19.3944
R10326 gnd.n5187 gnd.n5183 19.3944
R10327 gnd.n5187 gnd.n5184 19.3944
R10328 gnd.n5184 gnd.n1683 19.3944
R10329 gnd.n5224 gnd.n1683 19.3944
R10330 gnd.n5224 gnd.n1666 19.3944
R10331 gnd.n5244 gnd.n1666 19.3944
R10332 gnd.n5244 gnd.n1660 19.3944
R10333 gnd.n5252 gnd.n1660 19.3944
R10334 gnd.n5253 gnd.n5252 19.3944
R10335 gnd.n5253 gnd.n1643 19.3944
R10336 gnd.n5274 gnd.n1643 19.3944
R10337 gnd.n5275 gnd.n5274 19.3944
R10338 gnd.n5278 gnd.n5275 19.3944
R10339 gnd.n5279 gnd.n5278 19.3944
R10340 gnd.n5279 gnd.n1608 19.3944
R10341 gnd.n5310 gnd.n1608 19.3944
R10342 gnd.n5311 gnd.n5310 19.3944
R10343 gnd.n5314 gnd.n5311 19.3944
R10344 gnd.n5315 gnd.n5314 19.3944
R10345 gnd.n5315 gnd.n1579 19.3944
R10346 gnd.n5346 gnd.n1579 19.3944
R10347 gnd.n5347 gnd.n5346 19.3944
R10348 gnd.n5350 gnd.n5347 19.3944
R10349 gnd.n5351 gnd.n5350 19.3944
R10350 gnd.n5359 gnd.n5351 19.3944
R10351 gnd.n5359 gnd.n5357 19.3944
R10352 gnd.n5357 gnd.n5356 19.3944
R10353 gnd.n5356 gnd.n5355 19.3944
R10354 gnd.n5355 gnd.n5352 19.3944
R10355 gnd.n5352 gnd.n1513 19.3944
R10356 gnd.n5434 gnd.n1513 19.3944
R10357 gnd.n5435 gnd.n5434 19.3944
R10358 gnd.n5437 gnd.n5435 19.3944
R10359 gnd.n5437 gnd.n1444 19.3944
R10360 gnd.n5856 gnd.n1444 19.3944
R10361 gnd.n5857 gnd.n5856 19.3944
R10362 gnd.n5857 gnd.n1424 19.3944
R10363 gnd.n5968 gnd.n1424 19.3944
R10364 gnd.n5969 gnd.n5968 19.3944
R10365 gnd.n5041 gnd.n5040 19.3944
R10366 gnd.n5040 gnd.n5035 19.3944
R10367 gnd.n5035 gnd.n1808 19.3944
R10368 gnd.n5061 gnd.n1808 19.3944
R10369 gnd.n5061 gnd.n5060 19.3944
R10370 gnd.n5060 gnd.n5059 19.3944
R10371 gnd.n5059 gnd.n1789 19.3944
R10372 gnd.n5085 gnd.n1789 19.3944
R10373 gnd.n5085 gnd.n5084 19.3944
R10374 gnd.n5084 gnd.n5083 19.3944
R10375 gnd.n5083 gnd.n5082 19.3944
R10376 gnd.n5082 gnd.n1763 19.3944
R10377 gnd.n5120 gnd.n1763 19.3944
R10378 gnd.n5120 gnd.n5119 19.3944
R10379 gnd.n5119 gnd.n5118 19.3944
R10380 gnd.n5118 gnd.n5117 19.3944
R10381 gnd.n5117 gnd.n1738 19.3944
R10382 gnd.n5155 gnd.n1738 19.3944
R10383 gnd.n5155 gnd.n5154 19.3944
R10384 gnd.n5154 gnd.n5153 19.3944
R10385 gnd.n5153 gnd.n5152 19.3944
R10386 gnd.n5152 gnd.n1711 19.3944
R10387 gnd.n5192 gnd.n1711 19.3944
R10388 gnd.n5192 gnd.n5191 19.3944
R10389 gnd.n5191 gnd.n5190 19.3944
R10390 gnd.n5190 gnd.n5189 19.3944
R10391 gnd.n5189 gnd.n1690 19.3944
R10392 gnd.n1690 gnd.n1681 19.3944
R10393 gnd.n5226 gnd.n1681 19.3944
R10394 gnd.n5227 gnd.n5226 19.3944
R10395 gnd.n5227 gnd.n1664 19.3944
R10396 gnd.n5247 gnd.n1664 19.3944
R10397 gnd.n5248 gnd.n5247 19.3944
R10398 gnd.n5248 gnd.n1658 19.3944
R10399 gnd.n5256 gnd.n1658 19.3944
R10400 gnd.n5256 gnd.n1640 19.3944
R10401 gnd.n5287 gnd.n1640 19.3944
R10402 gnd.n5287 gnd.n5286 19.3944
R10403 gnd.n5286 gnd.n5285 19.3944
R10404 gnd.n5285 gnd.n5284 19.3944
R10405 gnd.n5284 gnd.n1605 19.3944
R10406 gnd.n5323 gnd.n1605 19.3944
R10407 gnd.n5323 gnd.n5322 19.3944
R10408 gnd.n5322 gnd.n5321 19.3944
R10409 gnd.n5321 gnd.n5320 19.3944
R10410 gnd.n5320 gnd.n1574 19.3944
R10411 gnd.n5365 gnd.n1574 19.3944
R10412 gnd.n5365 gnd.n5364 19.3944
R10413 gnd.n5364 gnd.n5363 19.3944
R10414 gnd.n5363 gnd.n5362 19.3944
R10415 gnd.n5362 gnd.n1538 19.3944
R10416 gnd.n5408 gnd.n1538 19.3944
R10417 gnd.n5408 gnd.n5407 19.3944
R10418 gnd.n5407 gnd.n5406 19.3944
R10419 gnd.n5406 gnd.n5405 19.3944
R10420 gnd.n5405 gnd.n1511 19.3944
R10421 gnd.n5442 gnd.n1511 19.3944
R10422 gnd.n5442 gnd.n5441 19.3944
R10423 gnd.n5441 gnd.n5440 19.3944
R10424 gnd.n5440 gnd.n1442 19.3944
R10425 gnd.n5862 gnd.n1442 19.3944
R10426 gnd.n5862 gnd.n5861 19.3944
R10427 gnd.n5861 gnd.n5860 19.3944
R10428 gnd.n5860 gnd.n1423 19.3944
R10429 gnd.n5960 gnd.n5871 19.3944
R10430 gnd.n5955 gnd.n5871 19.3944
R10431 gnd.n5955 gnd.n5954 19.3944
R10432 gnd.n5954 gnd.n5953 19.3944
R10433 gnd.n5953 gnd.n5876 19.3944
R10434 gnd.n5948 gnd.n5876 19.3944
R10435 gnd.n5948 gnd.n5947 19.3944
R10436 gnd.n5947 gnd.n5946 19.3944
R10437 gnd.n5946 gnd.n5883 19.3944
R10438 gnd.n5941 gnd.n5883 19.3944
R10439 gnd.n5941 gnd.n5940 19.3944
R10440 gnd.n5940 gnd.n5939 19.3944
R10441 gnd.n5939 gnd.n5890 19.3944
R10442 gnd.n5934 gnd.n5890 19.3944
R10443 gnd.n5934 gnd.n5933 19.3944
R10444 gnd.n5933 gnd.n5932 19.3944
R10445 gnd.n5932 gnd.n5897 19.3944
R10446 gnd.n6008 gnd.n1381 19.3944
R10447 gnd.n6008 gnd.n1385 19.3944
R10448 gnd.n1388 gnd.n1385 19.3944
R10449 gnd.n6001 gnd.n1388 19.3944
R10450 gnd.n6001 gnd.n6000 19.3944
R10451 gnd.n6000 gnd.n5999 19.3944
R10452 gnd.n5999 gnd.n1394 19.3944
R10453 gnd.n5994 gnd.n1394 19.3944
R10454 gnd.n5994 gnd.n5993 19.3944
R10455 gnd.n5993 gnd.n5992 19.3944
R10456 gnd.n5992 gnd.n1401 19.3944
R10457 gnd.n5987 gnd.n1401 19.3944
R10458 gnd.n5987 gnd.n5986 19.3944
R10459 gnd.n5986 gnd.n5985 19.3944
R10460 gnd.n5985 gnd.n1408 19.3944
R10461 gnd.n5980 gnd.n1408 19.3944
R10462 gnd.n5980 gnd.n5979 19.3944
R10463 gnd.n5979 gnd.n5978 19.3944
R10464 gnd.n6027 gnd.n1361 19.3944
R10465 gnd.n6027 gnd.n1366 19.3944
R10466 gnd.n1370 gnd.n1366 19.3944
R10467 gnd.n6020 gnd.n1370 19.3944
R10468 gnd.n6020 gnd.n6019 19.3944
R10469 gnd.n6019 gnd.n6018 19.3944
R10470 gnd.n6018 gnd.n1376 19.3944
R10471 gnd.n6013 gnd.n1376 19.3944
R10472 gnd.n5927 gnd.n5926 19.3944
R10473 gnd.n5926 gnd.n5925 19.3944
R10474 gnd.n5925 gnd.n5907 19.3944
R10475 gnd.n5920 gnd.n5907 19.3944
R10476 gnd.n5920 gnd.n5919 19.3944
R10477 gnd.n5919 gnd.n5918 19.3944
R10478 gnd.n5918 gnd.n1362 19.3944
R10479 gnd.n5045 gnd.n1816 19.3944
R10480 gnd.n5049 gnd.n1816 19.3944
R10481 gnd.n5049 gnd.n1801 19.3944
R10482 gnd.n5065 gnd.n1801 19.3944
R10483 gnd.n5065 gnd.n1799 19.3944
R10484 gnd.n5069 gnd.n1799 19.3944
R10485 gnd.n5069 gnd.n1781 19.3944
R10486 gnd.n5089 gnd.n1781 19.3944
R10487 gnd.n5089 gnd.n1779 19.3944
R10488 gnd.n5095 gnd.n1779 19.3944
R10489 gnd.n5095 gnd.n5094 19.3944
R10490 gnd.n5094 gnd.n1756 19.3944
R10491 gnd.n5124 gnd.n1756 19.3944
R10492 gnd.n5124 gnd.n1754 19.3944
R10493 gnd.n5130 gnd.n1754 19.3944
R10494 gnd.n5130 gnd.n5129 19.3944
R10495 gnd.n5129 gnd.n1732 19.3944
R10496 gnd.n5159 gnd.n1732 19.3944
R10497 gnd.n5159 gnd.n1730 19.3944
R10498 gnd.n5165 gnd.n1730 19.3944
R10499 gnd.n5165 gnd.n5164 19.3944
R10500 gnd.n5164 gnd.n1705 19.3944
R10501 gnd.n5196 gnd.n1705 19.3944
R10502 gnd.n5196 gnd.n1703 19.3944
R10503 gnd.n5202 gnd.n1703 19.3944
R10504 gnd.n5202 gnd.n5201 19.3944
R10505 gnd.n5201 gnd.n5200 19.3944
R10506 gnd.n5220 gnd.n5219 19.3944
R10507 gnd.n5240 gnd.n5239 19.3944
R10508 gnd.n1674 gnd.n1673 19.3944
R10509 gnd.n5261 gnd.n5260 19.3944
R10510 gnd.n5291 gnd.n1632 19.3944
R10511 gnd.n5291 gnd.n1624 19.3944
R10512 gnd.n5297 gnd.n1624 19.3944
R10513 gnd.n5297 gnd.n5296 19.3944
R10514 gnd.n5296 gnd.n1597 19.3944
R10515 gnd.n5327 gnd.n1597 19.3944
R10516 gnd.n5327 gnd.n1595 19.3944
R10517 gnd.n5333 gnd.n1595 19.3944
R10518 gnd.n5333 gnd.n5332 19.3944
R10519 gnd.n5332 gnd.n1566 19.3944
R10520 gnd.n5369 gnd.n1566 19.3944
R10521 gnd.n5369 gnd.n1564 19.3944
R10522 gnd.n5375 gnd.n1564 19.3944
R10523 gnd.n5375 gnd.n5374 19.3944
R10524 gnd.n5374 gnd.n1530 19.3944
R10525 gnd.n5412 gnd.n1530 19.3944
R10526 gnd.n5412 gnd.n1528 19.3944
R10527 gnd.n5418 gnd.n1528 19.3944
R10528 gnd.n5418 gnd.n5417 19.3944
R10529 gnd.n5417 gnd.n1503 19.3944
R10530 gnd.n5446 gnd.n1503 19.3944
R10531 gnd.n5446 gnd.n1501 19.3944
R10532 gnd.n5450 gnd.n1501 19.3944
R10533 gnd.n5450 gnd.n1434 19.3944
R10534 gnd.n5866 gnd.n1434 19.3944
R10535 gnd.n5866 gnd.n1432 19.3944
R10536 gnd.n5964 gnd.n1432 19.3944
R10537 gnd.n5964 gnd.n5963 19.3944
R10538 gnd.n3114 gnd.n2097 19.3944
R10539 gnd.n3114 gnd.n2095 19.3944
R10540 gnd.n3118 gnd.n2095 19.3944
R10541 gnd.n3118 gnd.n2091 19.3944
R10542 gnd.n3124 gnd.n2091 19.3944
R10543 gnd.n3124 gnd.n2089 19.3944
R10544 gnd.n3128 gnd.n2089 19.3944
R10545 gnd.n3128 gnd.n2085 19.3944
R10546 gnd.n3134 gnd.n2085 19.3944
R10547 gnd.n3134 gnd.n2083 19.3944
R10548 gnd.n3138 gnd.n2083 19.3944
R10549 gnd.n3138 gnd.n2079 19.3944
R10550 gnd.n3144 gnd.n2079 19.3944
R10551 gnd.n3144 gnd.n2077 19.3944
R10552 gnd.n3148 gnd.n2077 19.3944
R10553 gnd.n3148 gnd.n2073 19.3944
R10554 gnd.n3154 gnd.n2073 19.3944
R10555 gnd.n3154 gnd.n2071 19.3944
R10556 gnd.n3158 gnd.n2071 19.3944
R10557 gnd.n3158 gnd.n2067 19.3944
R10558 gnd.n3164 gnd.n2067 19.3944
R10559 gnd.n3164 gnd.n2065 19.3944
R10560 gnd.n3168 gnd.n2065 19.3944
R10561 gnd.n3168 gnd.n2061 19.3944
R10562 gnd.n3174 gnd.n2061 19.3944
R10563 gnd.n3174 gnd.n2059 19.3944
R10564 gnd.n3178 gnd.n2059 19.3944
R10565 gnd.n3178 gnd.n2055 19.3944
R10566 gnd.n3184 gnd.n2055 19.3944
R10567 gnd.n3184 gnd.n2053 19.3944
R10568 gnd.n3188 gnd.n2053 19.3944
R10569 gnd.n3188 gnd.n2049 19.3944
R10570 gnd.n3194 gnd.n2049 19.3944
R10571 gnd.n3194 gnd.n2047 19.3944
R10572 gnd.n3198 gnd.n2047 19.3944
R10573 gnd.n3198 gnd.n2043 19.3944
R10574 gnd.n3204 gnd.n2043 19.3944
R10575 gnd.n3204 gnd.n2041 19.3944
R10576 gnd.n3208 gnd.n2041 19.3944
R10577 gnd.n3208 gnd.n2037 19.3944
R10578 gnd.n3214 gnd.n2037 19.3944
R10579 gnd.n3214 gnd.n2035 19.3944
R10580 gnd.n3218 gnd.n2035 19.3944
R10581 gnd.n3218 gnd.n2031 19.3944
R10582 gnd.n3224 gnd.n2031 19.3944
R10583 gnd.n3224 gnd.n2029 19.3944
R10584 gnd.n3228 gnd.n2029 19.3944
R10585 gnd.n3228 gnd.n2025 19.3944
R10586 gnd.n3234 gnd.n2025 19.3944
R10587 gnd.n3234 gnd.n2023 19.3944
R10588 gnd.n3238 gnd.n2023 19.3944
R10589 gnd.n3238 gnd.n2019 19.3944
R10590 gnd.n3244 gnd.n2019 19.3944
R10591 gnd.n3244 gnd.n2017 19.3944
R10592 gnd.n3248 gnd.n2017 19.3944
R10593 gnd.n3248 gnd.n2013 19.3944
R10594 gnd.n3254 gnd.n2013 19.3944
R10595 gnd.n3254 gnd.n2011 19.3944
R10596 gnd.n3258 gnd.n2011 19.3944
R10597 gnd.n3258 gnd.n2007 19.3944
R10598 gnd.n3264 gnd.n2007 19.3944
R10599 gnd.n3264 gnd.n2005 19.3944
R10600 gnd.n3268 gnd.n2005 19.3944
R10601 gnd.n3268 gnd.n2001 19.3944
R10602 gnd.n3274 gnd.n2001 19.3944
R10603 gnd.n3274 gnd.n1999 19.3944
R10604 gnd.n3278 gnd.n1999 19.3944
R10605 gnd.n3278 gnd.n1995 19.3944
R10606 gnd.n3284 gnd.n1995 19.3944
R10607 gnd.n3284 gnd.n1993 19.3944
R10608 gnd.n3288 gnd.n1993 19.3944
R10609 gnd.n3288 gnd.n1989 19.3944
R10610 gnd.n3294 gnd.n1989 19.3944
R10611 gnd.n3294 gnd.n1987 19.3944
R10612 gnd.n3298 gnd.n1987 19.3944
R10613 gnd.n3298 gnd.n1983 19.3944
R10614 gnd.n3304 gnd.n1983 19.3944
R10615 gnd.n3304 gnd.n1981 19.3944
R10616 gnd.n3308 gnd.n1981 19.3944
R10617 gnd.n3308 gnd.n1977 19.3944
R10618 gnd.n3314 gnd.n1977 19.3944
R10619 gnd.n3314 gnd.n1975 19.3944
R10620 gnd.n3320 gnd.n1975 19.3944
R10621 gnd.n3320 gnd.n3319 19.3944
R10622 gnd.n5680 gnd.n5482 19.3944
R10623 gnd.n5680 gnd.n5483 19.3944
R10624 gnd.n5676 gnd.n5483 19.3944
R10625 gnd.n5676 gnd.n5675 19.3944
R10626 gnd.n5675 gnd.n5674 19.3944
R10627 gnd.n5674 gnd.n5489 19.3944
R10628 gnd.n5670 gnd.n5489 19.3944
R10629 gnd.n5670 gnd.n5669 19.3944
R10630 gnd.n5669 gnd.n5668 19.3944
R10631 gnd.n5668 gnd.n5494 19.3944
R10632 gnd.n5664 gnd.n5494 19.3944
R10633 gnd.n5664 gnd.n5663 19.3944
R10634 gnd.n5663 gnd.n5662 19.3944
R10635 gnd.n5662 gnd.n5499 19.3944
R10636 gnd.n5658 gnd.n5499 19.3944
R10637 gnd.n5658 gnd.n5657 19.3944
R10638 gnd.n5657 gnd.n5656 19.3944
R10639 gnd.n5656 gnd.n1224 19.3944
R10640 gnd.n6102 gnd.n1224 19.3944
R10641 gnd.n6102 gnd.n1221 19.3944
R10642 gnd.n6107 gnd.n1221 19.3944
R10643 gnd.n6107 gnd.n1222 19.3944
R10644 gnd.n1222 gnd.n1182 19.3944
R10645 gnd.n6178 gnd.n1182 19.3944
R10646 gnd.n6178 gnd.n1179 19.3944
R10647 gnd.n6192 gnd.n1179 19.3944
R10648 gnd.n6192 gnd.n1180 19.3944
R10649 gnd.n6188 gnd.n1180 19.3944
R10650 gnd.n6188 gnd.n6187 19.3944
R10651 gnd.n6187 gnd.n6186 19.3944
R10652 gnd.n6186 gnd.n1133 19.3944
R10653 gnd.n6254 gnd.n1133 19.3944
R10654 gnd.n6254 gnd.n1131 19.3944
R10655 gnd.n6258 gnd.n1131 19.3944
R10656 gnd.n6258 gnd.n1105 19.3944
R10657 gnd.n6300 gnd.n1105 19.3944
R10658 gnd.n6300 gnd.n1103 19.3944
R10659 gnd.n6304 gnd.n1103 19.3944
R10660 gnd.n6304 gnd.n1074 19.3944
R10661 gnd.n6362 gnd.n1074 19.3944
R10662 gnd.n6362 gnd.n1072 19.3944
R10663 gnd.n6366 gnd.n1072 19.3944
R10664 gnd.n6366 gnd.n1047 19.3944
R10665 gnd.n6399 gnd.n1047 19.3944
R10666 gnd.n6399 gnd.n1045 19.3944
R10667 gnd.n6403 gnd.n1045 19.3944
R10668 gnd.n6403 gnd.n1018 19.3944
R10669 gnd.n6435 gnd.n1018 19.3944
R10670 gnd.n6435 gnd.n1016 19.3944
R10671 gnd.n6439 gnd.n1016 19.3944
R10672 gnd.n6439 gnd.n979 19.3944
R10673 gnd.n6492 gnd.n979 19.3944
R10674 gnd.n6492 gnd.n976 19.3944
R10675 gnd.n6497 gnd.n976 19.3944
R10676 gnd.n6497 gnd.n977 19.3944
R10677 gnd.n977 gnd.n956 19.3944
R10678 gnd.n6529 gnd.n956 19.3944
R10679 gnd.n6529 gnd.n957 19.3944
R10680 gnd.n6525 gnd.n957 19.3944
R10681 gnd.n6525 gnd.n6524 19.3944
R10682 gnd.n6524 gnd.n6523 19.3944
R10683 gnd.n6523 gnd.n881 19.3944
R10684 gnd.n6728 gnd.n881 19.3944
R10685 gnd.n6728 gnd.n878 19.3944
R10686 gnd.n6733 gnd.n878 19.3944
R10687 gnd.n6733 gnd.n879 19.3944
R10688 gnd.n879 gnd.n856 19.3944
R10689 gnd.n6758 gnd.n856 19.3944
R10690 gnd.n6758 gnd.n853 19.3944
R10691 gnd.n6763 gnd.n853 19.3944
R10692 gnd.n6763 gnd.n854 19.3944
R10693 gnd.n854 gnd.n831 19.3944
R10694 gnd.n6788 gnd.n831 19.3944
R10695 gnd.n6788 gnd.n828 19.3944
R10696 gnd.n6793 gnd.n828 19.3944
R10697 gnd.n6793 gnd.n829 19.3944
R10698 gnd.n829 gnd.n807 19.3944
R10699 gnd.n6824 gnd.n807 19.3944
R10700 gnd.n6824 gnd.n805 19.3944
R10701 gnd.n6828 gnd.n805 19.3944
R10702 gnd.n6828 gnd.n767 19.3944
R10703 gnd.n6859 gnd.n767 19.3944
R10704 gnd.n6856 gnd.n6855 19.3944
R10705 gnd.n6855 gnd.n6854 19.3944
R10706 gnd.n6854 gnd.n772 19.3944
R10707 gnd.n6850 gnd.n772 19.3944
R10708 gnd.n6850 gnd.n6849 19.3944
R10709 gnd.n6849 gnd.n697 19.3944
R10710 gnd.n6923 gnd.n697 19.3944
R10711 gnd.n6923 gnd.n6922 19.3944
R10712 gnd.n6922 gnd.n6921 19.3944
R10713 gnd.n6921 gnd.n701 19.3944
R10714 gnd.n6914 gnd.n701 19.3944
R10715 gnd.n6914 gnd.n6913 19.3944
R10716 gnd.n6913 gnd.n711 19.3944
R10717 gnd.n6906 gnd.n711 19.3944
R10718 gnd.n6906 gnd.n6905 19.3944
R10719 gnd.n6905 gnd.n721 19.3944
R10720 gnd.n6898 gnd.n721 19.3944
R10721 gnd.n6898 gnd.n6897 19.3944
R10722 gnd.n6897 gnd.n729 19.3944
R10723 gnd.n6890 gnd.n729 19.3944
R10724 gnd.n6890 gnd.n6889 19.3944
R10725 gnd.n6889 gnd.n739 19.3944
R10726 gnd.n6882 gnd.n739 19.3944
R10727 gnd.n6882 gnd.n6881 19.3944
R10728 gnd.n6871 gnd.n755 19.3944
R10729 gnd.n6871 gnd.n6870 19.3944
R10730 gnd.n6870 gnd.n758 19.3944
R10731 gnd.n4112 gnd.t165 18.8012
R10732 gnd.n4097 gnd.t157 18.8012
R10733 gnd.n2602 gnd.t225 18.8012
R10734 gnd.n3956 gnd.n3955 18.4825
R10735 gnd.n6990 gnd.n6989 18.4247
R10736 gnd.n6031 gnd.n1362 18.4247
R10737 gnd.n6878 gnd.n6877 18.2308
R10738 gnd.n5779 gnd.n5768 18.2308
R10739 gnd.n7443 gnd.n7394 18.2308
R10740 gnd.n4788 gnd.n4758 18.2308
R10741 gnd.t176 gnd.n3636 18.1639
R10742 gnd.n4612 gnd.n4611 17.8452
R10743 gnd.n3664 gnd.t9 17.5266
R10744 gnd.n4063 gnd.t184 16.8893
R10745 gnd.n6972 gnd.n6969 16.6793
R10746 gnd.n7588 gnd.n7585 16.6793
R10747 gnd.n4979 gnd.n4846 16.6793
R10748 gnd.n6013 gnd.n6012 16.6793
R10749 gnd.n3891 gnd.t15 16.2519
R10750 gnd.n3591 gnd.t180 16.2519
R10751 gnd.n1294 gnd.n1293 16.0975
R10752 gnd.n928 gnd.n927 16.0975
R10753 gnd.n1291 gnd.n1290 16.0975
R10754 gnd.n6572 gnd.n6571 16.0975
R10755 gnd.n5838 gnd.n1460 15.9333
R10756 gnd.n5838 gnd.n1474 15.9333
R10757 gnd.n5478 gnd.n5477 15.9333
R10758 gnd.n5683 gnd.n5478 15.9333
R10759 gnd.n5683 gnd.n5682 15.9333
R10760 gnd.n5682 gnd.n5480 15.9333
R10761 gnd.n5558 gnd.n5557 15.9333
R10762 gnd.n5557 gnd.n5550 15.9333
R10763 gnd.n5568 gnd.n5550 15.9333
R10764 gnd.n5568 gnd.n5567 15.9333
R10765 gnd.n5567 gnd.n5566 15.9333
R10766 gnd.n5566 gnd.n5543 15.9333
R10767 gnd.n5576 gnd.n5543 15.9333
R10768 gnd.n5579 gnd.n5576 15.9333
R10769 gnd.n5577 gnd.n5537 15.9333
R10770 gnd.n5589 gnd.n5537 15.9333
R10771 gnd.n5589 gnd.n5588 15.9333
R10772 gnd.n5588 gnd.n5587 15.9333
R10773 gnd.n5587 gnd.n5531 15.9333
R10774 gnd.n5597 gnd.n5531 15.9333
R10775 gnd.n5600 gnd.n5597 15.9333
R10776 gnd.n5600 gnd.n5598 15.9333
R10777 gnd.n5610 gnd.n5525 15.9333
R10778 gnd.n5610 gnd.n5609 15.9333
R10779 gnd.n5609 gnd.n5608 15.9333
R10780 gnd.n5608 gnd.n5519 15.9333
R10781 gnd.n5618 gnd.n5519 15.9333
R10782 gnd.n5621 gnd.n5618 15.9333
R10783 gnd.n5621 gnd.n5619 15.9333
R10784 gnd.n5619 gnd.n5512 15.9333
R10785 gnd.n5639 gnd.n5512 15.9333
R10786 gnd.n5638 gnd.n5503 15.9333
R10787 gnd.n5653 gnd.n5503 15.9333
R10788 gnd.n5653 gnd.n5652 15.9333
R10789 gnd.n5652 gnd.n5505 15.9333
R10790 gnd.n5505 gnd.n1226 15.9333
R10791 gnd.n6100 gnd.n1226 15.9333
R10792 gnd.n1262 gnd.n1261 15.9333
R10793 gnd.n1201 gnd.n1191 15.9333
R10794 gnd.n6176 gnd.n1186 15.9333
R10795 gnd.n6195 gnd.n6194 15.9333
R10796 gnd.n6207 gnd.n1167 15.9333
R10797 gnd.n1159 gnd.n1152 15.9333
R10798 gnd.n6252 gnd.n1135 15.9333
R10799 gnd.n6233 gnd.n6232 15.9333
R10800 gnd.n6287 gnd.n6286 15.9333
R10801 gnd.n6341 gnd.n1079 15.9333
R10802 gnd.n6342 gnd.n6341 15.9333
R10803 gnd.n6406 gnd.n1026 15.9333
R10804 gnd.n1039 gnd.n1022 15.9333
R10805 gnd.n6441 gnd.n1014 15.9333
R10806 gnd.n6490 gnd.n6489 15.9333
R10807 gnd.n6499 gnd.n973 15.9333
R10808 gnd.n6714 gnd.n6713 15.9333
R10809 gnd.n6726 gnd.n6725 15.9333
R10810 gnd.n6725 gnd.n884 15.9333
R10811 gnd.n884 gnd.n873 15.9333
R10812 gnd.n6735 gnd.n873 15.9333
R10813 gnd.n6735 gnd.n874 15.9333
R10814 gnd.n876 gnd.n874 15.9333
R10815 gnd.n6745 gnd.n6744 15.9333
R10816 gnd.n6744 gnd.n858 15.9333
R10817 gnd.n6756 gnd.n858 15.9333
R10818 gnd.n6756 gnd.n6755 15.9333
R10819 gnd.n6755 gnd.n860 15.9333
R10820 gnd.n860 gnd.n848 15.9333
R10821 gnd.n6765 gnd.n848 15.9333
R10822 gnd.n6765 gnd.n849 15.9333
R10823 gnd.n851 gnd.n849 15.9333
R10824 gnd.n6775 gnd.n6774 15.9333
R10825 gnd.n6774 gnd.n833 15.9333
R10826 gnd.n6786 gnd.n833 15.9333
R10827 gnd.n6786 gnd.n6785 15.9333
R10828 gnd.n6785 gnd.n835 15.9333
R10829 gnd.n835 gnd.n824 15.9333
R10830 gnd.n6795 gnd.n824 15.9333
R10831 gnd.n6795 gnd.n825 15.9333
R10832 gnd.n6810 gnd.n817 15.9333
R10833 gnd.n6810 gnd.n6809 15.9333
R10834 gnd.n6809 gnd.n809 15.9333
R10835 gnd.n6822 gnd.n809 15.9333
R10836 gnd.n6822 gnd.n6821 15.9333
R10837 gnd.n6821 gnd.n811 15.9333
R10838 gnd.n811 gnd.n802 15.9333
R10839 gnd.n6830 gnd.n802 15.9333
R10840 gnd.n6832 gnd.n6831 15.9333
R10841 gnd.n6831 gnd.n763 15.9333
R10842 gnd.n6861 gnd.n763 15.9333
R10843 gnd.n6861 gnd.n764 15.9333
R10844 gnd.n6845 gnd.n776 15.9333
R10845 gnd.n6845 gnd.n6844 15.9333
R10846 gnd.n4578 gnd.n4576 15.6674
R10847 gnd.n4546 gnd.n4544 15.6674
R10848 gnd.n4514 gnd.n4512 15.6674
R10849 gnd.n4483 gnd.n4481 15.6674
R10850 gnd.n4451 gnd.n4449 15.6674
R10851 gnd.n4419 gnd.n4417 15.6674
R10852 gnd.n4387 gnd.n4385 15.6674
R10853 gnd.n4356 gnd.n4354 15.6674
R10854 gnd.n3882 gnd.t15 15.6146
R10855 gnd.t127 gnd.n1900 15.6146
R10856 gnd.t108 gnd.n1901 15.6146
R10857 gnd.n5558 gnd.t19 15.6146
R10858 gnd.t52 gnd.n6830 15.6146
R10859 gnd.n6929 gnd.n692 15.3217
R10860 gnd.n7543 gnd.n345 15.3217
R10861 gnd.n5031 gnd.n4825 15.3217
R10862 gnd.n5973 gnd.n1417 15.3217
R10863 gnd.n6241 gnd.n6240 15.296
R10864 gnd.n6260 gnd.n1128 15.296
R10865 gnd.n6433 gnd.n6432 15.296
R10866 gnd.n1013 gnd.n1005 15.296
R10867 gnd.n6519 gnd.t80 15.296
R10868 gnd.n6556 gnd.n6555 15.0827
R10869 gnd.n1274 gnd.n1269 15.0481
R10870 gnd.n6566 gnd.n6565 15.0481
R10871 gnd.n4250 gnd.t8 14.9773
R10872 gnd.n5598 gnd.t168 14.9773
R10873 gnd.n6775 gnd.t397 14.9773
R10874 gnd.n6154 gnd.t87 14.6587
R10875 gnd.n1205 gnd.n1176 14.6587
R10876 gnd.n6482 gnd.n6481 14.6587
R10877 gnd.n6518 gnd.n932 14.6587
R10878 gnd.t393 gnd.n3356 14.34
R10879 gnd.n4328 gnd.t181 14.34
R10880 gnd.n4038 gnd.t385 13.7027
R10881 gnd.n3748 gnd.n3747 13.5763
R10882 gnd.n4693 gnd.n1857 13.5763
R10883 gnd.n3956 gnd.n3694 13.384
R10884 gnd.n1166 gnd.n1156 13.384
R10885 gnd.n6278 gnd.n1109 13.384
R10886 gnd.t1 gnd.n6279 13.384
R10887 gnd.t173 gnd.n6348 13.384
R10888 gnd.n6369 gnd.t159 13.384
R10889 gnd.n1066 gnd.t135 13.384
R10890 gnd.n6380 gnd.n6379 13.384
R10891 gnd.n6456 gnd.n972 13.384
R10892 gnd.n1285 gnd.n1266 13.1884
R10893 gnd.n1280 gnd.n1279 13.1884
R10894 gnd.n1279 gnd.n1278 13.1884
R10895 gnd.n6559 gnd.n6554 13.1884
R10896 gnd.n6560 gnd.n6559 13.1884
R10897 gnd.n1281 gnd.n1268 13.146
R10898 gnd.n1277 gnd.n1268 13.146
R10899 gnd.n6558 gnd.n6557 13.146
R10900 gnd.n6558 gnd.n6553 13.146
R10901 gnd.t131 gnd.n5638 13.0654
R10902 gnd.n876 gnd.t145 13.0654
R10903 gnd.n4579 gnd.n4575 12.8005
R10904 gnd.n4547 gnd.n4543 12.8005
R10905 gnd.n4515 gnd.n4511 12.8005
R10906 gnd.n4484 gnd.n4480 12.8005
R10907 gnd.n4452 gnd.n4448 12.8005
R10908 gnd.n4420 gnd.n4416 12.8005
R10909 gnd.n4388 gnd.n4384 12.8005
R10910 gnd.n4357 gnd.n4353 12.8005
R10911 gnd.n6109 gnd.n1218 12.7467
R10912 gnd.n6208 gnd.n1164 12.7467
R10913 gnd.n6306 gnd.n1099 12.7467
R10914 gnd.n6397 gnd.n6396 12.7467
R10915 gnd.n6464 gnd.n995 12.7467
R10916 gnd.n1786 gnd.t217 12.4281
R10917 gnd.n7692 gnd.t301 12.4281
R10918 gnd.n3747 gnd.n3742 12.4126
R10919 gnd.n4696 gnd.n4693 12.4126
R10920 gnd.n6096 gnd.n1289 12.1761
R10921 gnd.n6639 gnd.n6638 12.1761
R10922 gnd.n6176 gnd.t23 12.1094
R10923 gnd.n6222 gnd.n6221 12.1094
R10924 gnd.n6288 gnd.n1114 12.1094
R10925 gnd.n6426 gnd.n6425 12.1094
R10926 gnd.n1006 gnd.n981 12.1094
R10927 gnd.n6538 gnd.t26 12.1094
R10928 gnd.n4583 gnd.n4582 12.0247
R10929 gnd.n4551 gnd.n4550 12.0247
R10930 gnd.n4519 gnd.n4518 12.0247
R10931 gnd.n4488 gnd.n4487 12.0247
R10932 gnd.n4456 gnd.n4455 12.0247
R10933 gnd.n4424 gnd.n4423 12.0247
R10934 gnd.n4392 gnd.n4391 12.0247
R10935 gnd.n4361 gnd.n4360 12.0247
R10936 gnd.n5142 gnd.t262 11.7908
R10937 gnd.n5402 gnd.t187 11.7908
R10938 gnd.n545 gnd.t193 11.7908
R10939 gnd.n7716 gnd.t195 11.7908
R10940 gnd.n5690 gnd.n1369 11.4721
R10941 gnd.n6165 gnd.n6164 11.4721
R10942 gnd.n6360 gnd.n1076 11.4721
R10943 gnd.n6370 gnd.n6368 11.4721
R10944 gnd.n6532 gnd.n6531 11.4721
R10945 gnd.n6539 gnd.t12 11.4721
R10946 gnd.n6548 gnd.n938 11.4721
R10947 gnd.n7042 gnd.n7041 11.4721
R10948 gnd.n4586 gnd.n4573 11.249
R10949 gnd.n4554 gnd.n4541 11.249
R10950 gnd.n4522 gnd.n4509 11.249
R10951 gnd.n4491 gnd.n4478 11.249
R10952 gnd.n4459 gnd.n4446 11.249
R10953 gnd.n4427 gnd.n4414 11.249
R10954 gnd.n4395 gnd.n4382 11.249
R10955 gnd.n4364 gnd.n4351 11.249
R10956 gnd.n4026 gnd.t385 11.1535
R10957 gnd.n5204 gnd.t206 11.1535
R10958 gnd.t228 gnd.n1568 11.1535
R10959 gnd.n5579 gnd.t389 11.1535
R10960 gnd.t155 gnd.n817 11.1535
R10961 gnd.n7180 gnd.t189 11.1535
R10962 gnd.n7740 gnd.t220 11.1535
R10963 gnd.n6234 gnd.n1145 10.8348
R10964 gnd.n6419 gnd.n6418 10.8348
R10965 gnd.n6932 gnd.n6929 10.6672
R10966 gnd.n7546 gnd.n7543 10.6672
R10967 gnd.n4826 gnd.n4825 10.6672
R10968 gnd.n5978 gnd.n1417 10.6672
R10969 gnd.n6709 gnd.n6708 10.6151
R10970 gnd.n6708 gnd.n6705 10.6151
R10971 gnd.n6703 gnd.n6700 10.6151
R10972 gnd.n6700 gnd.n6699 10.6151
R10973 gnd.n6699 gnd.n6696 10.6151
R10974 gnd.n6696 gnd.n6695 10.6151
R10975 gnd.n6695 gnd.n6692 10.6151
R10976 gnd.n6692 gnd.n6691 10.6151
R10977 gnd.n6691 gnd.n6688 10.6151
R10978 gnd.n6688 gnd.n6687 10.6151
R10979 gnd.n6687 gnd.n6684 10.6151
R10980 gnd.n6684 gnd.n6683 10.6151
R10981 gnd.n6683 gnd.n6680 10.6151
R10982 gnd.n6680 gnd.n6679 10.6151
R10983 gnd.n6679 gnd.n6676 10.6151
R10984 gnd.n6676 gnd.n6675 10.6151
R10985 gnd.n6675 gnd.n6672 10.6151
R10986 gnd.n6672 gnd.n6671 10.6151
R10987 gnd.n6671 gnd.n6668 10.6151
R10988 gnd.n6668 gnd.n6667 10.6151
R10989 gnd.n6667 gnd.n6664 10.6151
R10990 gnd.n6664 gnd.n6663 10.6151
R10991 gnd.n6663 gnd.n6660 10.6151
R10992 gnd.n6660 gnd.n6659 10.6151
R10993 gnd.n6659 gnd.n6656 10.6151
R10994 gnd.n6656 gnd.n6655 10.6151
R10995 gnd.n6655 gnd.n6652 10.6151
R10996 gnd.n6652 gnd.n6651 10.6151
R10997 gnd.n6651 gnd.n6648 10.6151
R10998 gnd.n6648 gnd.n6647 10.6151
R10999 gnd.n1295 gnd.n1203 10.6151
R11000 gnd.n6152 gnd.n1203 10.6151
R11001 gnd.n6152 gnd.n6151 10.6151
R11002 gnd.n6151 gnd.n6150 10.6151
R11003 gnd.n6150 gnd.n6149 10.6151
R11004 gnd.n6149 gnd.n6148 10.6151
R11005 gnd.n6148 gnd.n1204 10.6151
R11006 gnd.n1210 gnd.n1204 10.6151
R11007 gnd.n1210 gnd.n1209 10.6151
R11008 gnd.n1209 gnd.n1208 10.6151
R11009 gnd.n1208 gnd.n1154 10.6151
R11010 gnd.n6217 gnd.n1154 10.6151
R11011 gnd.n6218 gnd.n6217 10.6151
R11012 gnd.n6219 gnd.n6218 10.6151
R11013 gnd.n6219 gnd.n1144 10.6151
R11014 gnd.n6238 gnd.n1144 10.6151
R11015 gnd.n6238 gnd.n6237 10.6151
R11016 gnd.n6237 gnd.n6236 10.6151
R11017 gnd.n6236 gnd.n1126 10.6151
R11018 gnd.n6263 gnd.n1126 10.6151
R11019 gnd.n6264 gnd.n6263 10.6151
R11020 gnd.n6266 gnd.n6264 10.6151
R11021 gnd.n6267 gnd.n6266 10.6151
R11022 gnd.n6276 gnd.n6267 10.6151
R11023 gnd.n6276 gnd.n6275 10.6151
R11024 gnd.n6275 gnd.n6274 10.6151
R11025 gnd.n6274 gnd.n6272 10.6151
R11026 gnd.n6272 gnd.n6271 10.6151
R11027 gnd.n6271 gnd.n6269 10.6151
R11028 gnd.n6269 gnd.n6268 10.6151
R11029 gnd.n6268 gnd.n1067 10.6151
R11030 gnd.n6372 gnd.n1067 10.6151
R11031 gnd.n6373 gnd.n6372 10.6151
R11032 gnd.n6375 gnd.n6373 10.6151
R11033 gnd.n6376 gnd.n6375 10.6151
R11034 gnd.n6377 gnd.n6376 10.6151
R11035 gnd.n6377 gnd.n1040 10.6151
R11036 gnd.n6409 gnd.n1040 10.6151
R11037 gnd.n6410 gnd.n6409 10.6151
R11038 gnd.n6412 gnd.n6410 10.6151
R11039 gnd.n6413 gnd.n6412 10.6151
R11040 gnd.n6416 gnd.n6413 10.6151
R11041 gnd.n6416 gnd.n6415 10.6151
R11042 gnd.n6415 gnd.n6414 10.6151
R11043 gnd.n6414 gnd.n1003 10.6151
R11044 gnd.n6452 gnd.n1003 10.6151
R11045 gnd.n6453 gnd.n6452 10.6151
R11046 gnd.n6454 gnd.n6453 10.6151
R11047 gnd.n6454 gnd.n993 10.6151
R11048 gnd.n6466 gnd.n993 10.6151
R11049 gnd.n6467 gnd.n6466 10.6151
R11050 gnd.n6478 gnd.n6467 10.6151
R11051 gnd.n6478 gnd.n6477 10.6151
R11052 gnd.n6477 gnd.n6476 10.6151
R11053 gnd.n6476 gnd.n6474 10.6151
R11054 gnd.n6474 gnd.n6473 10.6151
R11055 gnd.n6473 gnd.n6469 10.6151
R11056 gnd.n6469 gnd.n6468 10.6151
R11057 gnd.n6468 gnd.n931 10.6151
R11058 gnd.n931 gnd.n929 10.6151
R11059 gnd.n1360 gnd.n1359 10.6151
R11060 gnd.n1359 gnd.n1356 10.6151
R11061 gnd.n1354 gnd.n1351 10.6151
R11062 gnd.n1351 gnd.n1350 10.6151
R11063 gnd.n1350 gnd.n1347 10.6151
R11064 gnd.n1347 gnd.n1346 10.6151
R11065 gnd.n1346 gnd.n1343 10.6151
R11066 gnd.n1343 gnd.n1342 10.6151
R11067 gnd.n1342 gnd.n1339 10.6151
R11068 gnd.n1339 gnd.n1338 10.6151
R11069 gnd.n1338 gnd.n1335 10.6151
R11070 gnd.n1335 gnd.n1334 10.6151
R11071 gnd.n1334 gnd.n1331 10.6151
R11072 gnd.n1331 gnd.n1330 10.6151
R11073 gnd.n1330 gnd.n1327 10.6151
R11074 gnd.n1327 gnd.n1326 10.6151
R11075 gnd.n1326 gnd.n1323 10.6151
R11076 gnd.n1323 gnd.n1322 10.6151
R11077 gnd.n1322 gnd.n1319 10.6151
R11078 gnd.n1319 gnd.n1318 10.6151
R11079 gnd.n1318 gnd.n1315 10.6151
R11080 gnd.n1315 gnd.n1314 10.6151
R11081 gnd.n1314 gnd.n1311 10.6151
R11082 gnd.n1311 gnd.n1310 10.6151
R11083 gnd.n1310 gnd.n1307 10.6151
R11084 gnd.n1307 gnd.n1306 10.6151
R11085 gnd.n1306 gnd.n1303 10.6151
R11086 gnd.n1303 gnd.n1302 10.6151
R11087 gnd.n1302 gnd.n1299 10.6151
R11088 gnd.n1299 gnd.n1298 10.6151
R11089 gnd.n6096 gnd.n6095 10.6151
R11090 gnd.n6095 gnd.n6094 10.6151
R11091 gnd.n6094 gnd.n6093 10.6151
R11092 gnd.n6093 gnd.n6091 10.6151
R11093 gnd.n6091 gnd.n6088 10.6151
R11094 gnd.n6088 gnd.n6087 10.6151
R11095 gnd.n6087 gnd.n6084 10.6151
R11096 gnd.n6084 gnd.n6083 10.6151
R11097 gnd.n6083 gnd.n6080 10.6151
R11098 gnd.n6080 gnd.n6079 10.6151
R11099 gnd.n6079 gnd.n6076 10.6151
R11100 gnd.n6076 gnd.n6075 10.6151
R11101 gnd.n6075 gnd.n6072 10.6151
R11102 gnd.n6072 gnd.n6071 10.6151
R11103 gnd.n6071 gnd.n6068 10.6151
R11104 gnd.n6068 gnd.n6067 10.6151
R11105 gnd.n6067 gnd.n6064 10.6151
R11106 gnd.n6064 gnd.n6063 10.6151
R11107 gnd.n6063 gnd.n6060 10.6151
R11108 gnd.n6060 gnd.n6059 10.6151
R11109 gnd.n6059 gnd.n6056 10.6151
R11110 gnd.n6056 gnd.n6055 10.6151
R11111 gnd.n6055 gnd.n6052 10.6151
R11112 gnd.n6052 gnd.n6051 10.6151
R11113 gnd.n6051 gnd.n6048 10.6151
R11114 gnd.n6048 gnd.n6047 10.6151
R11115 gnd.n6047 gnd.n6044 10.6151
R11116 gnd.n6044 gnd.n6043 10.6151
R11117 gnd.n6040 gnd.n6039 10.6151
R11118 gnd.n6039 gnd.n6036 10.6151
R11119 gnd.n6638 gnd.n6636 10.6151
R11120 gnd.n6636 gnd.n6633 10.6151
R11121 gnd.n6633 gnd.n6632 10.6151
R11122 gnd.n6632 gnd.n6629 10.6151
R11123 gnd.n6629 gnd.n6628 10.6151
R11124 gnd.n6628 gnd.n6625 10.6151
R11125 gnd.n6625 gnd.n6624 10.6151
R11126 gnd.n6624 gnd.n6621 10.6151
R11127 gnd.n6621 gnd.n6620 10.6151
R11128 gnd.n6620 gnd.n6617 10.6151
R11129 gnd.n6617 gnd.n6616 10.6151
R11130 gnd.n6616 gnd.n6613 10.6151
R11131 gnd.n6613 gnd.n6612 10.6151
R11132 gnd.n6612 gnd.n6609 10.6151
R11133 gnd.n6609 gnd.n6608 10.6151
R11134 gnd.n6608 gnd.n6605 10.6151
R11135 gnd.n6605 gnd.n6604 10.6151
R11136 gnd.n6604 gnd.n6601 10.6151
R11137 gnd.n6601 gnd.n6600 10.6151
R11138 gnd.n6600 gnd.n6597 10.6151
R11139 gnd.n6597 gnd.n6596 10.6151
R11140 gnd.n6596 gnd.n6593 10.6151
R11141 gnd.n6593 gnd.n6592 10.6151
R11142 gnd.n6592 gnd.n6589 10.6151
R11143 gnd.n6589 gnd.n6588 10.6151
R11144 gnd.n6588 gnd.n6585 10.6151
R11145 gnd.n6585 gnd.n6584 10.6151
R11146 gnd.n6584 gnd.n6581 10.6151
R11147 gnd.n6579 gnd.n6576 10.6151
R11148 gnd.n6576 gnd.n6575 10.6151
R11149 gnd.n1288 gnd.n1287 10.6151
R11150 gnd.n1287 gnd.n1189 10.6151
R11151 gnd.n6167 gnd.n1189 10.6151
R11152 gnd.n6168 gnd.n6167 10.6151
R11153 gnd.n6174 gnd.n6168 10.6151
R11154 gnd.n6174 gnd.n6173 10.6151
R11155 gnd.n6173 gnd.n6172 10.6151
R11156 gnd.n6172 gnd.n6169 10.6151
R11157 gnd.n6169 gnd.n1162 10.6151
R11158 gnd.n6210 gnd.n1162 10.6151
R11159 gnd.n6211 gnd.n6210 10.6151
R11160 gnd.n6213 gnd.n6211 10.6151
R11161 gnd.n6213 gnd.n6212 10.6151
R11162 gnd.n6212 gnd.n1140 10.6151
R11163 gnd.n6244 gnd.n1140 10.6151
R11164 gnd.n6245 gnd.n6244 10.6151
R11165 gnd.n6249 gnd.n6245 10.6151
R11166 gnd.n6249 gnd.n6248 10.6151
R11167 gnd.n6248 gnd.n6247 10.6151
R11168 gnd.n6247 gnd.n1112 10.6151
R11169 gnd.n6290 gnd.n1112 10.6151
R11170 gnd.n6291 gnd.n6290 10.6151
R11171 gnd.n6295 gnd.n6291 10.6151
R11172 gnd.n6295 gnd.n6294 10.6151
R11173 gnd.n6294 gnd.n6293 10.6151
R11174 gnd.n6293 gnd.n1082 10.6151
R11175 gnd.n6352 gnd.n1082 10.6151
R11176 gnd.n6353 gnd.n6352 10.6151
R11177 gnd.n6357 gnd.n6353 10.6151
R11178 gnd.n6357 gnd.n6356 10.6151
R11179 gnd.n6356 gnd.n6355 10.6151
R11180 gnd.n6355 gnd.n1055 10.6151
R11181 gnd.n6389 gnd.n1055 10.6151
R11182 gnd.n6390 gnd.n6389 10.6151
R11183 gnd.n6394 gnd.n6390 10.6151
R11184 gnd.n6394 gnd.n6393 10.6151
R11185 gnd.n6393 gnd.n6392 10.6151
R11186 gnd.n6392 gnd.n1024 10.6151
R11187 gnd.n6428 gnd.n1024 10.6151
R11188 gnd.n6429 gnd.n6428 10.6151
R11189 gnd.n6430 gnd.n6429 10.6151
R11190 gnd.n6430 gnd.n1009 10.6151
R11191 gnd.n6444 gnd.n1009 10.6151
R11192 gnd.n6445 gnd.n6444 10.6151
R11193 gnd.n6447 gnd.n6445 10.6151
R11194 gnd.n6447 gnd.n6446 10.6151
R11195 gnd.n6446 gnd.n998 10.6151
R11196 gnd.n6459 gnd.n998 10.6151
R11197 gnd.n6460 gnd.n6459 10.6151
R11198 gnd.n6462 gnd.n6460 10.6151
R11199 gnd.n6462 gnd.n6461 10.6151
R11200 gnd.n6461 gnd.n950 10.6151
R11201 gnd.n6534 gnd.n950 10.6151
R11202 gnd.n6535 gnd.n6534 10.6151
R11203 gnd.n6536 gnd.n6535 10.6151
R11204 gnd.n6536 gnd.n936 10.6151
R11205 gnd.n6550 gnd.n936 10.6151
R11206 gnd.n6551 gnd.n6550 10.6151
R11207 gnd.n6641 gnd.n6551 10.6151
R11208 gnd.n6641 gnd.n6640 10.6151
R11209 gnd.n3945 gnd.t153 10.5161
R11210 gnd.n3358 gnd.t393 10.5161
R11211 gnd.n4311 gnd.t181 10.5161
R11212 gnd.n5250 gnd.t247 10.5161
R11213 gnd.t236 gnd.n1618 10.5161
R11214 gnd.t197 gnd.n404 10.5161
R11215 gnd.n7330 gnd.t296 10.5161
R11216 gnd.n4587 gnd.n4571 10.4732
R11217 gnd.n4555 gnd.n4539 10.4732
R11218 gnd.n4523 gnd.n4507 10.4732
R11219 gnd.n4492 gnd.n4476 10.4732
R11220 gnd.n4460 gnd.n4444 10.4732
R11221 gnd.n4428 gnd.n4412 10.4732
R11222 gnd.n4396 gnd.n4380 10.4732
R11223 gnd.n4365 gnd.n4349 10.4732
R11224 gnd.n6164 gnd.n6163 10.1975
R11225 gnd.n1160 gnd.t174 10.1975
R11226 gnd.n6360 gnd.n6359 10.1975
R11227 gnd.n6368 gnd.n1069 10.1975
R11228 gnd.n1001 gnd.t6 10.1975
R11229 gnd.n6471 gnd.n938 10.1975
R11230 gnd.t8 gnd.n3375 9.87883
R11231 gnd.n5194 gnd.t287 9.87883
R11232 gnd.t264 gnd.n1668 9.87883
R11233 gnd.n5308 gnd.t303 9.87883
R11234 gnd.n6100 gnd.n6099 9.87883
R11235 gnd.n7275 gnd.t271 9.87883
R11236 gnd.n7344 gnd.t199 9.87883
R11237 gnd.n7734 gnd.t251 9.87883
R11238 gnd.n4591 gnd.n4590 9.69747
R11239 gnd.n4559 gnd.n4558 9.69747
R11240 gnd.n4527 gnd.n4526 9.69747
R11241 gnd.n4496 gnd.n4495 9.69747
R11242 gnd.n4464 gnd.n4463 9.69747
R11243 gnd.n4432 gnd.n4431 9.69747
R11244 gnd.n4400 gnd.n4399 9.69747
R11245 gnd.n4369 gnd.n4368 9.69747
R11246 gnd.n6261 gnd.n1114 9.56018
R11247 gnd.n6425 gnd.n1028 9.56018
R11248 gnd.t62 gnd.n952 9.56018
R11249 gnd.n4597 gnd.n4596 9.45567
R11250 gnd.n4565 gnd.n4564 9.45567
R11251 gnd.n4533 gnd.n4532 9.45567
R11252 gnd.n4502 gnd.n4501 9.45567
R11253 gnd.n4470 gnd.n4469 9.45567
R11254 gnd.n4438 gnd.n4437 9.45567
R11255 gnd.n4406 gnd.n4405 9.45567
R11256 gnd.n4375 gnd.n4374 9.45567
R11257 gnd.n6969 gnd.n6968 9.30959
R11258 gnd.n7585 gnd.n325 9.30959
R11259 gnd.n4979 gnd.n4844 9.30959
R11260 gnd.n6012 gnd.n1381 9.30959
R11261 gnd.n4596 gnd.n4595 9.3005
R11262 gnd.n4569 gnd.n4568 9.3005
R11263 gnd.n4590 gnd.n4589 9.3005
R11264 gnd.n4588 gnd.n4587 9.3005
R11265 gnd.n4573 gnd.n4572 9.3005
R11266 gnd.n4582 gnd.n4581 9.3005
R11267 gnd.n4580 gnd.n4579 9.3005
R11268 gnd.n4564 gnd.n4563 9.3005
R11269 gnd.n4537 gnd.n4536 9.3005
R11270 gnd.n4558 gnd.n4557 9.3005
R11271 gnd.n4556 gnd.n4555 9.3005
R11272 gnd.n4541 gnd.n4540 9.3005
R11273 gnd.n4550 gnd.n4549 9.3005
R11274 gnd.n4548 gnd.n4547 9.3005
R11275 gnd.n4532 gnd.n4531 9.3005
R11276 gnd.n4505 gnd.n4504 9.3005
R11277 gnd.n4526 gnd.n4525 9.3005
R11278 gnd.n4524 gnd.n4523 9.3005
R11279 gnd.n4509 gnd.n4508 9.3005
R11280 gnd.n4518 gnd.n4517 9.3005
R11281 gnd.n4516 gnd.n4515 9.3005
R11282 gnd.n4501 gnd.n4500 9.3005
R11283 gnd.n4474 gnd.n4473 9.3005
R11284 gnd.n4495 gnd.n4494 9.3005
R11285 gnd.n4493 gnd.n4492 9.3005
R11286 gnd.n4478 gnd.n4477 9.3005
R11287 gnd.n4487 gnd.n4486 9.3005
R11288 gnd.n4485 gnd.n4484 9.3005
R11289 gnd.n4469 gnd.n4468 9.3005
R11290 gnd.n4442 gnd.n4441 9.3005
R11291 gnd.n4463 gnd.n4462 9.3005
R11292 gnd.n4461 gnd.n4460 9.3005
R11293 gnd.n4446 gnd.n4445 9.3005
R11294 gnd.n4455 gnd.n4454 9.3005
R11295 gnd.n4453 gnd.n4452 9.3005
R11296 gnd.n4437 gnd.n4436 9.3005
R11297 gnd.n4410 gnd.n4409 9.3005
R11298 gnd.n4431 gnd.n4430 9.3005
R11299 gnd.n4429 gnd.n4428 9.3005
R11300 gnd.n4414 gnd.n4413 9.3005
R11301 gnd.n4423 gnd.n4422 9.3005
R11302 gnd.n4421 gnd.n4420 9.3005
R11303 gnd.n4405 gnd.n4404 9.3005
R11304 gnd.n4378 gnd.n4377 9.3005
R11305 gnd.n4399 gnd.n4398 9.3005
R11306 gnd.n4397 gnd.n4396 9.3005
R11307 gnd.n4382 gnd.n4381 9.3005
R11308 gnd.n4391 gnd.n4390 9.3005
R11309 gnd.n4389 gnd.n4388 9.3005
R11310 gnd.n4374 gnd.n4373 9.3005
R11311 gnd.n4347 gnd.n4346 9.3005
R11312 gnd.n4368 gnd.n4367 9.3005
R11313 gnd.n4366 gnd.n4365 9.3005
R11314 gnd.n4351 gnd.n4350 9.3005
R11315 gnd.n4360 gnd.n4359 9.3005
R11316 gnd.n4358 gnd.n4357 9.3005
R11317 gnd.n4723 gnd.n4722 9.3005
R11318 gnd.n4721 gnd.n1845 9.3005
R11319 gnd.n4720 gnd.n4719 9.3005
R11320 gnd.n4716 gnd.n1846 9.3005
R11321 gnd.n4713 gnd.n1847 9.3005
R11322 gnd.n4712 gnd.n1848 9.3005
R11323 gnd.n4709 gnd.n1849 9.3005
R11324 gnd.n4708 gnd.n1850 9.3005
R11325 gnd.n4705 gnd.n1851 9.3005
R11326 gnd.n4704 gnd.n1852 9.3005
R11327 gnd.n4701 gnd.n1853 9.3005
R11328 gnd.n4700 gnd.n1854 9.3005
R11329 gnd.n4697 gnd.n1855 9.3005
R11330 gnd.n4696 gnd.n1856 9.3005
R11331 gnd.n4693 gnd.n4692 9.3005
R11332 gnd.n4691 gnd.n1857 9.3005
R11333 gnd.n4724 gnd.n1844 9.3005
R11334 gnd.n3964 gnd.n3963 9.3005
R11335 gnd.n3668 gnd.n3667 9.3005
R11336 gnd.n3991 gnd.n3990 9.3005
R11337 gnd.n3992 gnd.n3666 9.3005
R11338 gnd.n3996 gnd.n3993 9.3005
R11339 gnd.n3995 gnd.n3994 9.3005
R11340 gnd.n3640 gnd.n3639 9.3005
R11341 gnd.n4021 gnd.n4020 9.3005
R11342 gnd.n4022 gnd.n3638 9.3005
R11343 gnd.n4024 gnd.n4023 9.3005
R11344 gnd.n3618 gnd.n3617 9.3005
R11345 gnd.n4052 gnd.n4051 9.3005
R11346 gnd.n4053 gnd.n3616 9.3005
R11347 gnd.n4061 gnd.n4054 9.3005
R11348 gnd.n4060 gnd.n4055 9.3005
R11349 gnd.n4059 gnd.n4057 9.3005
R11350 gnd.n4056 gnd.n3565 9.3005
R11351 gnd.n4109 gnd.n3566 9.3005
R11352 gnd.n4108 gnd.n3567 9.3005
R11353 gnd.n4107 gnd.n3568 9.3005
R11354 gnd.n3587 gnd.n3569 9.3005
R11355 gnd.n3589 gnd.n3588 9.3005
R11356 gnd.n3455 gnd.n3454 9.3005
R11357 gnd.n4147 gnd.n4146 9.3005
R11358 gnd.n4148 gnd.n3453 9.3005
R11359 gnd.n4152 gnd.n4149 9.3005
R11360 gnd.n4151 gnd.n4150 9.3005
R11361 gnd.n3428 gnd.n3427 9.3005
R11362 gnd.n4187 gnd.n4186 9.3005
R11363 gnd.n4188 gnd.n3426 9.3005
R11364 gnd.n4192 gnd.n4189 9.3005
R11365 gnd.n4191 gnd.n4190 9.3005
R11366 gnd.n3401 gnd.n3400 9.3005
R11367 gnd.n4232 gnd.n4231 9.3005
R11368 gnd.n4233 gnd.n3399 9.3005
R11369 gnd.n4237 gnd.n4234 9.3005
R11370 gnd.n4236 gnd.n4235 9.3005
R11371 gnd.n3373 gnd.n3372 9.3005
R11372 gnd.n4272 gnd.n4271 9.3005
R11373 gnd.n4273 gnd.n3371 9.3005
R11374 gnd.n4277 gnd.n4274 9.3005
R11375 gnd.n4276 gnd.n4275 9.3005
R11376 gnd.n3346 gnd.n3345 9.3005
R11377 gnd.n4321 gnd.n4320 9.3005
R11378 gnd.n4322 gnd.n3344 9.3005
R11379 gnd.n4326 gnd.n4323 9.3005
R11380 gnd.n4325 gnd.n4324 9.3005
R11381 gnd.n1906 gnd.n1905 9.3005
R11382 gnd.n4616 gnd.n4615 9.3005
R11383 gnd.n4617 gnd.n1904 9.3005
R11384 gnd.n4623 gnd.n4618 9.3005
R11385 gnd.n4622 gnd.n4619 9.3005
R11386 gnd.n4621 gnd.n4620 9.3005
R11387 gnd.n3965 gnd.n3962 9.3005
R11388 gnd.n3747 gnd.n3706 9.3005
R11389 gnd.n3742 gnd.n3741 9.3005
R11390 gnd.n3740 gnd.n3707 9.3005
R11391 gnd.n3739 gnd.n3738 9.3005
R11392 gnd.n3735 gnd.n3708 9.3005
R11393 gnd.n3732 gnd.n3731 9.3005
R11394 gnd.n3730 gnd.n3709 9.3005
R11395 gnd.n3729 gnd.n3728 9.3005
R11396 gnd.n3725 gnd.n3710 9.3005
R11397 gnd.n3722 gnd.n3721 9.3005
R11398 gnd.n3720 gnd.n3711 9.3005
R11399 gnd.n3719 gnd.n3718 9.3005
R11400 gnd.n3715 gnd.n3713 9.3005
R11401 gnd.n3712 gnd.n3692 9.3005
R11402 gnd.n3959 gnd.n3691 9.3005
R11403 gnd.n3961 gnd.n3960 9.3005
R11404 gnd.n3749 gnd.n3748 9.3005
R11405 gnd.n3972 gnd.n3678 9.3005
R11406 gnd.n3979 gnd.n3679 9.3005
R11407 gnd.n3981 gnd.n3980 9.3005
R11408 gnd.n3982 gnd.n3659 9.3005
R11409 gnd.n4001 gnd.n4000 9.3005
R11410 gnd.n4003 gnd.n3651 9.3005
R11411 gnd.n4010 gnd.n3653 9.3005
R11412 gnd.n4011 gnd.n3648 9.3005
R11413 gnd.n4013 gnd.n4012 9.3005
R11414 gnd.n3649 gnd.n3634 9.3005
R11415 gnd.n4029 gnd.n3632 9.3005
R11416 gnd.n4033 gnd.n4032 9.3005
R11417 gnd.n4031 gnd.n3608 9.3005
R11418 gnd.n4068 gnd.n3607 9.3005
R11419 gnd.n4071 gnd.n4070 9.3005
R11420 gnd.n3604 gnd.n3603 9.3005
R11421 gnd.n4077 gnd.n3605 9.3005
R11422 gnd.n4079 gnd.n4078 9.3005
R11423 gnd.n4081 gnd.n3602 9.3005
R11424 gnd.n4084 gnd.n4083 9.3005
R11425 gnd.n4087 gnd.n4085 9.3005
R11426 gnd.n4089 gnd.n4088 9.3005
R11427 gnd.n4095 gnd.n4090 9.3005
R11428 gnd.n4094 gnd.n4093 9.3005
R11429 gnd.n3446 gnd.n3445 9.3005
R11430 gnd.n4161 gnd.n4160 9.3005
R11431 gnd.n4162 gnd.n3439 9.3005
R11432 gnd.n4170 gnd.n3438 9.3005
R11433 gnd.n4173 gnd.n4172 9.3005
R11434 gnd.n4175 gnd.n4174 9.3005
R11435 gnd.n4178 gnd.n3421 9.3005
R11436 gnd.n4176 gnd.n3419 9.3005
R11437 gnd.n4198 gnd.n3417 9.3005
R11438 gnd.n4200 gnd.n4199 9.3005
R11439 gnd.n3391 gnd.n3390 9.3005
R11440 gnd.n4246 gnd.n4245 9.3005
R11441 gnd.n4247 gnd.n3384 9.3005
R11442 gnd.n4255 gnd.n3383 9.3005
R11443 gnd.n4258 gnd.n4257 9.3005
R11444 gnd.n4260 gnd.n4259 9.3005
R11445 gnd.n4263 gnd.n3366 9.3005
R11446 gnd.n4261 gnd.n3364 9.3005
R11447 gnd.n4283 gnd.n3362 9.3005
R11448 gnd.n4285 gnd.n4284 9.3005
R11449 gnd.n3337 gnd.n3336 9.3005
R11450 gnd.n4335 gnd.n4334 9.3005
R11451 gnd.n4336 gnd.n3330 9.3005
R11452 gnd.n4344 gnd.n3329 9.3005
R11453 gnd.n4603 gnd.n4602 9.3005
R11454 gnd.n4605 gnd.n4604 9.3005
R11455 gnd.n4606 gnd.n1897 9.3005
R11456 gnd.n4631 gnd.n4630 9.3005
R11457 gnd.n1898 gnd.n1860 9.3005
R11458 gnd.n3970 gnd.n3969 9.3005
R11459 gnd.n4687 gnd.n1861 9.3005
R11460 gnd.n4686 gnd.n1863 9.3005
R11461 gnd.n4683 gnd.n1864 9.3005
R11462 gnd.n4682 gnd.n1865 9.3005
R11463 gnd.n4679 gnd.n1866 9.3005
R11464 gnd.n4678 gnd.n1867 9.3005
R11465 gnd.n4675 gnd.n1868 9.3005
R11466 gnd.n4674 gnd.n1869 9.3005
R11467 gnd.n4671 gnd.n1870 9.3005
R11468 gnd.n4670 gnd.n1871 9.3005
R11469 gnd.n4667 gnd.n1872 9.3005
R11470 gnd.n4666 gnd.n1873 9.3005
R11471 gnd.n4663 gnd.n1874 9.3005
R11472 gnd.n4662 gnd.n1875 9.3005
R11473 gnd.n4659 gnd.n1876 9.3005
R11474 gnd.n4658 gnd.n1877 9.3005
R11475 gnd.n4655 gnd.n1878 9.3005
R11476 gnd.n4654 gnd.n1879 9.3005
R11477 gnd.n4651 gnd.n1880 9.3005
R11478 gnd.n4650 gnd.n1881 9.3005
R11479 gnd.n4647 gnd.n1882 9.3005
R11480 gnd.n4646 gnd.n1883 9.3005
R11481 gnd.n4643 gnd.n1887 9.3005
R11482 gnd.n4642 gnd.n1888 9.3005
R11483 gnd.n4639 gnd.n1889 9.3005
R11484 gnd.n4638 gnd.n1890 9.3005
R11485 gnd.n4689 gnd.n4688 9.3005
R11486 gnd.n4139 gnd.n4123 9.3005
R11487 gnd.n4138 gnd.n4124 9.3005
R11488 gnd.n4137 gnd.n4125 9.3005
R11489 gnd.n4135 gnd.n4126 9.3005
R11490 gnd.n4134 gnd.n4127 9.3005
R11491 gnd.n4132 gnd.n4128 9.3005
R11492 gnd.n4131 gnd.n4129 9.3005
R11493 gnd.n3409 gnd.n3408 9.3005
R11494 gnd.n4208 gnd.n4207 9.3005
R11495 gnd.n4209 gnd.n3407 9.3005
R11496 gnd.n4226 gnd.n4210 9.3005
R11497 gnd.n4225 gnd.n4211 9.3005
R11498 gnd.n4224 gnd.n4212 9.3005
R11499 gnd.n4222 gnd.n4213 9.3005
R11500 gnd.n4221 gnd.n4214 9.3005
R11501 gnd.n4219 gnd.n4215 9.3005
R11502 gnd.n4218 gnd.n4216 9.3005
R11503 gnd.n3353 gnd.n3352 9.3005
R11504 gnd.n4293 gnd.n4292 9.3005
R11505 gnd.n4294 gnd.n3351 9.3005
R11506 gnd.n4315 gnd.n4295 9.3005
R11507 gnd.n4314 gnd.n4296 9.3005
R11508 gnd.n4313 gnd.n4297 9.3005
R11509 gnd.n4310 gnd.n4298 9.3005
R11510 gnd.n4309 gnd.n4299 9.3005
R11511 gnd.n4307 gnd.n4300 9.3005
R11512 gnd.n4306 gnd.n4301 9.3005
R11513 gnd.n4304 gnd.n4303 9.3005
R11514 gnd.n4302 gnd.n1892 9.3005
R11515 gnd.n3880 gnd.n3879 9.3005
R11516 gnd.n3770 gnd.n3769 9.3005
R11517 gnd.n3894 gnd.n3893 9.3005
R11518 gnd.n3895 gnd.n3768 9.3005
R11519 gnd.n3897 gnd.n3896 9.3005
R11520 gnd.n3758 gnd.n3757 9.3005
R11521 gnd.n3910 gnd.n3909 9.3005
R11522 gnd.n3911 gnd.n3756 9.3005
R11523 gnd.n3943 gnd.n3912 9.3005
R11524 gnd.n3942 gnd.n3913 9.3005
R11525 gnd.n3941 gnd.n3914 9.3005
R11526 gnd.n3940 gnd.n3915 9.3005
R11527 gnd.n3937 gnd.n3916 9.3005
R11528 gnd.n3936 gnd.n3917 9.3005
R11529 gnd.n3935 gnd.n3918 9.3005
R11530 gnd.n3933 gnd.n3919 9.3005
R11531 gnd.n3932 gnd.n3920 9.3005
R11532 gnd.n3929 gnd.n3921 9.3005
R11533 gnd.n3928 gnd.n3922 9.3005
R11534 gnd.n3927 gnd.n3923 9.3005
R11535 gnd.n3925 gnd.n3924 9.3005
R11536 gnd.n3624 gnd.n3623 9.3005
R11537 gnd.n4041 gnd.n4040 9.3005
R11538 gnd.n4042 gnd.n3622 9.3005
R11539 gnd.n4046 gnd.n4043 9.3005
R11540 gnd.n4045 gnd.n4044 9.3005
R11541 gnd.n3546 gnd.n3545 9.3005
R11542 gnd.n4121 gnd.n4120 9.3005
R11543 gnd.n3878 gnd.n3779 9.3005
R11544 gnd.n3781 gnd.n3780 9.3005
R11545 gnd.n3825 gnd.n3823 9.3005
R11546 gnd.n3826 gnd.n3822 9.3005
R11547 gnd.n3829 gnd.n3818 9.3005
R11548 gnd.n3830 gnd.n3817 9.3005
R11549 gnd.n3833 gnd.n3816 9.3005
R11550 gnd.n3834 gnd.n3815 9.3005
R11551 gnd.n3837 gnd.n3814 9.3005
R11552 gnd.n3838 gnd.n3813 9.3005
R11553 gnd.n3841 gnd.n3812 9.3005
R11554 gnd.n3842 gnd.n3811 9.3005
R11555 gnd.n3845 gnd.n3810 9.3005
R11556 gnd.n3846 gnd.n3809 9.3005
R11557 gnd.n3849 gnd.n3808 9.3005
R11558 gnd.n3850 gnd.n3807 9.3005
R11559 gnd.n3853 gnd.n3806 9.3005
R11560 gnd.n3854 gnd.n3805 9.3005
R11561 gnd.n3857 gnd.n3804 9.3005
R11562 gnd.n3858 gnd.n3803 9.3005
R11563 gnd.n3861 gnd.n3802 9.3005
R11564 gnd.n3862 gnd.n3801 9.3005
R11565 gnd.n3865 gnd.n3800 9.3005
R11566 gnd.n3867 gnd.n3799 9.3005
R11567 gnd.n3868 gnd.n3798 9.3005
R11568 gnd.n3869 gnd.n3797 9.3005
R11569 gnd.n3870 gnd.n3796 9.3005
R11570 gnd.n3877 gnd.n3876 9.3005
R11571 gnd.n3886 gnd.n3885 9.3005
R11572 gnd.n3887 gnd.n3773 9.3005
R11573 gnd.n3889 gnd.n3888 9.3005
R11574 gnd.n3764 gnd.n3763 9.3005
R11575 gnd.n3902 gnd.n3901 9.3005
R11576 gnd.n3903 gnd.n3762 9.3005
R11577 gnd.n3905 gnd.n3904 9.3005
R11578 gnd.n3751 gnd.n3750 9.3005
R11579 gnd.n3948 gnd.n3947 9.3005
R11580 gnd.n3949 gnd.n3705 9.3005
R11581 gnd.n3953 gnd.n3951 9.3005
R11582 gnd.n3952 gnd.n3684 9.3005
R11583 gnd.n3971 gnd.n3683 9.3005
R11584 gnd.n3974 gnd.n3973 9.3005
R11585 gnd.n3677 gnd.n3676 9.3005
R11586 gnd.n3985 gnd.n3983 9.3005
R11587 gnd.n3984 gnd.n3658 9.3005
R11588 gnd.n4002 gnd.n3657 9.3005
R11589 gnd.n4005 gnd.n4004 9.3005
R11590 gnd.n3652 gnd.n3647 9.3005
R11591 gnd.n4015 gnd.n4014 9.3005
R11592 gnd.n3650 gnd.n3630 9.3005
R11593 gnd.n4036 gnd.n3631 9.3005
R11594 gnd.n4035 gnd.n4034 9.3005
R11595 gnd.n3633 gnd.n3609 9.3005
R11596 gnd.n4067 gnd.n4066 9.3005
R11597 gnd.n4069 gnd.n3554 9.3005
R11598 gnd.n4116 gnd.n3555 9.3005
R11599 gnd.n4115 gnd.n3556 9.3005
R11600 gnd.n4114 gnd.n3557 9.3005
R11601 gnd.n4080 gnd.n3558 9.3005
R11602 gnd.n4082 gnd.n3576 9.3005
R11603 gnd.n4102 gnd.n3577 9.3005
R11604 gnd.n4101 gnd.n3578 9.3005
R11605 gnd.n4100 gnd.n3579 9.3005
R11606 gnd.n4091 gnd.n3580 9.3005
R11607 gnd.n4092 gnd.n3447 9.3005
R11608 gnd.n4158 gnd.n4157 9.3005
R11609 gnd.n4159 gnd.n3440 9.3005
R11610 gnd.n4169 gnd.n4168 9.3005
R11611 gnd.n4171 gnd.n3436 9.3005
R11612 gnd.n4181 gnd.n3437 9.3005
R11613 gnd.n4180 gnd.n4179 9.3005
R11614 gnd.n4177 gnd.n3415 9.3005
R11615 gnd.n4203 gnd.n3416 9.3005
R11616 gnd.n4202 gnd.n4201 9.3005
R11617 gnd.n3418 gnd.n3392 9.3005
R11618 gnd.n4243 gnd.n4242 9.3005
R11619 gnd.n4244 gnd.n3385 9.3005
R11620 gnd.n4254 gnd.n4253 9.3005
R11621 gnd.n4256 gnd.n3381 9.3005
R11622 gnd.n4266 gnd.n3382 9.3005
R11623 gnd.n4265 gnd.n4264 9.3005
R11624 gnd.n4262 gnd.n3360 9.3005
R11625 gnd.n4288 gnd.n3361 9.3005
R11626 gnd.n4287 gnd.n4286 9.3005
R11627 gnd.n3363 gnd.n3338 9.3005
R11628 gnd.n4332 gnd.n4331 9.3005
R11629 gnd.n4333 gnd.n3331 9.3005
R11630 gnd.n4343 gnd.n4342 9.3005
R11631 gnd.n4601 gnd.n3327 9.3005
R11632 gnd.n4609 gnd.n3328 9.3005
R11633 gnd.n4608 gnd.n4607 9.3005
R11634 gnd.n1896 gnd.n1895 9.3005
R11635 gnd.n4633 gnd.n4632 9.3005
R11636 gnd.n3775 gnd.n3774 9.3005
R11637 gnd.n3108 gnd.n3107 9.3005
R11638 gnd.n3106 gnd.n2101 9.3005
R11639 gnd.n3105 gnd.n3104 9.3005
R11640 gnd.n2103 gnd.n2102 9.3005
R11641 gnd.n3098 gnd.n2107 9.3005
R11642 gnd.n3097 gnd.n2108 9.3005
R11643 gnd.n3096 gnd.n2109 9.3005
R11644 gnd.n2114 gnd.n2110 9.3005
R11645 gnd.n3090 gnd.n2115 9.3005
R11646 gnd.n3089 gnd.n2116 9.3005
R11647 gnd.n3088 gnd.n2117 9.3005
R11648 gnd.n2122 gnd.n2118 9.3005
R11649 gnd.n3082 gnd.n2123 9.3005
R11650 gnd.n3081 gnd.n2124 9.3005
R11651 gnd.n3080 gnd.n2125 9.3005
R11652 gnd.n2130 gnd.n2126 9.3005
R11653 gnd.n3074 gnd.n2131 9.3005
R11654 gnd.n3073 gnd.n2132 9.3005
R11655 gnd.n3072 gnd.n2133 9.3005
R11656 gnd.n2138 gnd.n2134 9.3005
R11657 gnd.n3066 gnd.n2139 9.3005
R11658 gnd.n3065 gnd.n2140 9.3005
R11659 gnd.n3064 gnd.n2141 9.3005
R11660 gnd.n2146 gnd.n2142 9.3005
R11661 gnd.n3058 gnd.n2147 9.3005
R11662 gnd.n3057 gnd.n2148 9.3005
R11663 gnd.n3056 gnd.n2149 9.3005
R11664 gnd.n2154 gnd.n2150 9.3005
R11665 gnd.n3050 gnd.n2155 9.3005
R11666 gnd.n3049 gnd.n2156 9.3005
R11667 gnd.n3048 gnd.n2157 9.3005
R11668 gnd.n2162 gnd.n2158 9.3005
R11669 gnd.n3042 gnd.n2163 9.3005
R11670 gnd.n3041 gnd.n2164 9.3005
R11671 gnd.n3040 gnd.n2165 9.3005
R11672 gnd.n2170 gnd.n2166 9.3005
R11673 gnd.n3034 gnd.n2171 9.3005
R11674 gnd.n3033 gnd.n2172 9.3005
R11675 gnd.n3032 gnd.n2173 9.3005
R11676 gnd.n2178 gnd.n2174 9.3005
R11677 gnd.n3026 gnd.n2179 9.3005
R11678 gnd.n3025 gnd.n2180 9.3005
R11679 gnd.n3024 gnd.n2181 9.3005
R11680 gnd.n2186 gnd.n2182 9.3005
R11681 gnd.n3018 gnd.n2187 9.3005
R11682 gnd.n3017 gnd.n2188 9.3005
R11683 gnd.n3016 gnd.n2189 9.3005
R11684 gnd.n2194 gnd.n2190 9.3005
R11685 gnd.n3010 gnd.n2195 9.3005
R11686 gnd.n3009 gnd.n2196 9.3005
R11687 gnd.n3008 gnd.n2197 9.3005
R11688 gnd.n2202 gnd.n2198 9.3005
R11689 gnd.n3002 gnd.n2203 9.3005
R11690 gnd.n3001 gnd.n2204 9.3005
R11691 gnd.n3000 gnd.n2205 9.3005
R11692 gnd.n2210 gnd.n2206 9.3005
R11693 gnd.n2994 gnd.n2211 9.3005
R11694 gnd.n2993 gnd.n2212 9.3005
R11695 gnd.n2992 gnd.n2213 9.3005
R11696 gnd.n2218 gnd.n2214 9.3005
R11697 gnd.n2986 gnd.n2219 9.3005
R11698 gnd.n2985 gnd.n2220 9.3005
R11699 gnd.n2984 gnd.n2221 9.3005
R11700 gnd.n2226 gnd.n2222 9.3005
R11701 gnd.n2978 gnd.n2227 9.3005
R11702 gnd.n2977 gnd.n2228 9.3005
R11703 gnd.n2976 gnd.n2229 9.3005
R11704 gnd.n2234 gnd.n2230 9.3005
R11705 gnd.n2970 gnd.n2235 9.3005
R11706 gnd.n2969 gnd.n2236 9.3005
R11707 gnd.n2968 gnd.n2237 9.3005
R11708 gnd.n2242 gnd.n2238 9.3005
R11709 gnd.n2962 gnd.n2243 9.3005
R11710 gnd.n2961 gnd.n2244 9.3005
R11711 gnd.n2960 gnd.n2245 9.3005
R11712 gnd.n2250 gnd.n2246 9.3005
R11713 gnd.n2954 gnd.n2251 9.3005
R11714 gnd.n2953 gnd.n2252 9.3005
R11715 gnd.n2952 gnd.n2253 9.3005
R11716 gnd.n2258 gnd.n2254 9.3005
R11717 gnd.n2946 gnd.n2259 9.3005
R11718 gnd.n2945 gnd.n2260 9.3005
R11719 gnd.n2944 gnd.n2261 9.3005
R11720 gnd.n2266 gnd.n2262 9.3005
R11721 gnd.n2938 gnd.n2267 9.3005
R11722 gnd.n2937 gnd.n2268 9.3005
R11723 gnd.n2936 gnd.n2269 9.3005
R11724 gnd.n2274 gnd.n2270 9.3005
R11725 gnd.n2930 gnd.n2275 9.3005
R11726 gnd.n2929 gnd.n2276 9.3005
R11727 gnd.n2928 gnd.n2277 9.3005
R11728 gnd.n2282 gnd.n2278 9.3005
R11729 gnd.n2922 gnd.n2283 9.3005
R11730 gnd.n2921 gnd.n2284 9.3005
R11731 gnd.n2920 gnd.n2285 9.3005
R11732 gnd.n2290 gnd.n2286 9.3005
R11733 gnd.n2914 gnd.n2291 9.3005
R11734 gnd.n2913 gnd.n2292 9.3005
R11735 gnd.n2912 gnd.n2293 9.3005
R11736 gnd.n2298 gnd.n2294 9.3005
R11737 gnd.n2906 gnd.n2299 9.3005
R11738 gnd.n2905 gnd.n2300 9.3005
R11739 gnd.n2904 gnd.n2301 9.3005
R11740 gnd.n2306 gnd.n2302 9.3005
R11741 gnd.n2898 gnd.n2307 9.3005
R11742 gnd.n2897 gnd.n2308 9.3005
R11743 gnd.n2896 gnd.n2309 9.3005
R11744 gnd.n2314 gnd.n2310 9.3005
R11745 gnd.n2890 gnd.n2315 9.3005
R11746 gnd.n2889 gnd.n2316 9.3005
R11747 gnd.n2888 gnd.n2317 9.3005
R11748 gnd.n2322 gnd.n2318 9.3005
R11749 gnd.n2882 gnd.n2323 9.3005
R11750 gnd.n2881 gnd.n2324 9.3005
R11751 gnd.n2880 gnd.n2325 9.3005
R11752 gnd.n2330 gnd.n2326 9.3005
R11753 gnd.n2874 gnd.n2331 9.3005
R11754 gnd.n2873 gnd.n2332 9.3005
R11755 gnd.n2872 gnd.n2333 9.3005
R11756 gnd.n2338 gnd.n2334 9.3005
R11757 gnd.n2866 gnd.n2339 9.3005
R11758 gnd.n2865 gnd.n2340 9.3005
R11759 gnd.n2864 gnd.n2341 9.3005
R11760 gnd.n2346 gnd.n2342 9.3005
R11761 gnd.n2858 gnd.n2347 9.3005
R11762 gnd.n2857 gnd.n2348 9.3005
R11763 gnd.n2856 gnd.n2349 9.3005
R11764 gnd.n2354 gnd.n2350 9.3005
R11765 gnd.n2850 gnd.n2355 9.3005
R11766 gnd.n2849 gnd.n2356 9.3005
R11767 gnd.n2848 gnd.n2357 9.3005
R11768 gnd.n2362 gnd.n2358 9.3005
R11769 gnd.n2842 gnd.n2363 9.3005
R11770 gnd.n2841 gnd.n2364 9.3005
R11771 gnd.n2840 gnd.n2365 9.3005
R11772 gnd.n2370 gnd.n2366 9.3005
R11773 gnd.n2834 gnd.n2371 9.3005
R11774 gnd.n2833 gnd.n2372 9.3005
R11775 gnd.n2832 gnd.n2373 9.3005
R11776 gnd.n2378 gnd.n2374 9.3005
R11777 gnd.n2826 gnd.n2379 9.3005
R11778 gnd.n2825 gnd.n2380 9.3005
R11779 gnd.n2824 gnd.n2381 9.3005
R11780 gnd.n2386 gnd.n2382 9.3005
R11781 gnd.n2818 gnd.n2387 9.3005
R11782 gnd.n2817 gnd.n2388 9.3005
R11783 gnd.n2816 gnd.n2389 9.3005
R11784 gnd.n2394 gnd.n2390 9.3005
R11785 gnd.n2810 gnd.n2395 9.3005
R11786 gnd.n2809 gnd.n2396 9.3005
R11787 gnd.n2808 gnd.n2397 9.3005
R11788 gnd.n2402 gnd.n2398 9.3005
R11789 gnd.n2802 gnd.n2403 9.3005
R11790 gnd.n2801 gnd.n2404 9.3005
R11791 gnd.n2800 gnd.n2405 9.3005
R11792 gnd.n2410 gnd.n2406 9.3005
R11793 gnd.n2794 gnd.n2411 9.3005
R11794 gnd.n2793 gnd.n2412 9.3005
R11795 gnd.n2792 gnd.n2413 9.3005
R11796 gnd.n2418 gnd.n2414 9.3005
R11797 gnd.n2786 gnd.n2419 9.3005
R11798 gnd.n2785 gnd.n2420 9.3005
R11799 gnd.n2784 gnd.n2421 9.3005
R11800 gnd.n2426 gnd.n2422 9.3005
R11801 gnd.n2778 gnd.n2427 9.3005
R11802 gnd.n2777 gnd.n2428 9.3005
R11803 gnd.n2776 gnd.n2429 9.3005
R11804 gnd.n2434 gnd.n2430 9.3005
R11805 gnd.n2769 gnd.n2768 9.3005
R11806 gnd.n2767 gnd.n2436 9.3005
R11807 gnd.n2766 gnd.n2765 9.3005
R11808 gnd.n2438 gnd.n2437 9.3005
R11809 gnd.n2759 gnd.n2444 9.3005
R11810 gnd.n2758 gnd.n2445 9.3005
R11811 gnd.n2757 gnd.n2446 9.3005
R11812 gnd.n2451 gnd.n2447 9.3005
R11813 gnd.n2751 gnd.n2452 9.3005
R11814 gnd.n2750 gnd.n2453 9.3005
R11815 gnd.n2749 gnd.n2454 9.3005
R11816 gnd.n2459 gnd.n2455 9.3005
R11817 gnd.n2743 gnd.n2460 9.3005
R11818 gnd.n2742 gnd.n2461 9.3005
R11819 gnd.n2741 gnd.n2462 9.3005
R11820 gnd.n2467 gnd.n2463 9.3005
R11821 gnd.n2735 gnd.n2468 9.3005
R11822 gnd.n2734 gnd.n2469 9.3005
R11823 gnd.n2733 gnd.n2470 9.3005
R11824 gnd.n2475 gnd.n2471 9.3005
R11825 gnd.n2727 gnd.n2476 9.3005
R11826 gnd.n2726 gnd.n2477 9.3005
R11827 gnd.n2725 gnd.n2478 9.3005
R11828 gnd.n2483 gnd.n2479 9.3005
R11829 gnd.n2719 gnd.n2484 9.3005
R11830 gnd.n2718 gnd.n2485 9.3005
R11831 gnd.n2717 gnd.n2486 9.3005
R11832 gnd.n2491 gnd.n2487 9.3005
R11833 gnd.n2711 gnd.n2492 9.3005
R11834 gnd.n2710 gnd.n2493 9.3005
R11835 gnd.n2709 gnd.n2494 9.3005
R11836 gnd.n2499 gnd.n2495 9.3005
R11837 gnd.n2703 gnd.n2500 9.3005
R11838 gnd.n2702 gnd.n2501 9.3005
R11839 gnd.n2701 gnd.n2502 9.3005
R11840 gnd.n2507 gnd.n2503 9.3005
R11841 gnd.n2695 gnd.n2508 9.3005
R11842 gnd.n2694 gnd.n2509 9.3005
R11843 gnd.n2693 gnd.n2510 9.3005
R11844 gnd.n2515 gnd.n2511 9.3005
R11845 gnd.n2687 gnd.n2516 9.3005
R11846 gnd.n2686 gnd.n2517 9.3005
R11847 gnd.n2685 gnd.n2518 9.3005
R11848 gnd.n2523 gnd.n2519 9.3005
R11849 gnd.n2679 gnd.n2524 9.3005
R11850 gnd.n2678 gnd.n2525 9.3005
R11851 gnd.n2677 gnd.n2526 9.3005
R11852 gnd.n2531 gnd.n2527 9.3005
R11853 gnd.n2671 gnd.n2532 9.3005
R11854 gnd.n2670 gnd.n2533 9.3005
R11855 gnd.n2669 gnd.n2534 9.3005
R11856 gnd.n2539 gnd.n2535 9.3005
R11857 gnd.n2663 gnd.n2540 9.3005
R11858 gnd.n2662 gnd.n2541 9.3005
R11859 gnd.n2661 gnd.n2542 9.3005
R11860 gnd.n2547 gnd.n2543 9.3005
R11861 gnd.n2655 gnd.n2548 9.3005
R11862 gnd.n2654 gnd.n2549 9.3005
R11863 gnd.n2653 gnd.n2550 9.3005
R11864 gnd.n2555 gnd.n2551 9.3005
R11865 gnd.n2647 gnd.n2556 9.3005
R11866 gnd.n2646 gnd.n2557 9.3005
R11867 gnd.n2645 gnd.n2558 9.3005
R11868 gnd.n2563 gnd.n2559 9.3005
R11869 gnd.n2639 gnd.n2564 9.3005
R11870 gnd.n2638 gnd.n2565 9.3005
R11871 gnd.n2637 gnd.n2566 9.3005
R11872 gnd.n2571 gnd.n2567 9.3005
R11873 gnd.n2631 gnd.n2572 9.3005
R11874 gnd.n2630 gnd.n2573 9.3005
R11875 gnd.n2629 gnd.n2574 9.3005
R11876 gnd.n2579 gnd.n2575 9.3005
R11877 gnd.n2623 gnd.n2580 9.3005
R11878 gnd.n2622 gnd.n2581 9.3005
R11879 gnd.n2621 gnd.n2582 9.3005
R11880 gnd.n2587 gnd.n2583 9.3005
R11881 gnd.n2615 gnd.n2588 9.3005
R11882 gnd.n2614 gnd.n2589 9.3005
R11883 gnd.n2613 gnd.n2590 9.3005
R11884 gnd.n2595 gnd.n2591 9.3005
R11885 gnd.n2607 gnd.n2596 9.3005
R11886 gnd.n2606 gnd.n2597 9.3005
R11887 gnd.n2605 gnd.n2598 9.3005
R11888 gnd.n2600 gnd.n2599 9.3005
R11889 gnd.n2770 gnd.n2435 9.3005
R11890 gnd.n7758 gnd.n7757 9.3005
R11891 gnd.n7756 gnd.n97 9.3005
R11892 gnd.n351 gnd.n99 9.3005
R11893 gnd.n7363 gnd.n7362 9.3005
R11894 gnd.n7364 gnd.n350 9.3005
R11895 gnd.n7488 gnd.n7365 9.3005
R11896 gnd.n7487 gnd.n7366 9.3005
R11897 gnd.n7486 gnd.n7367 9.3005
R11898 gnd.n7484 gnd.n7368 9.3005
R11899 gnd.n7483 gnd.n7369 9.3005
R11900 gnd.n7481 gnd.n7370 9.3005
R11901 gnd.n7480 gnd.n7371 9.3005
R11902 gnd.n7478 gnd.n7372 9.3005
R11903 gnd.n7477 gnd.n7373 9.3005
R11904 gnd.n7475 gnd.n7374 9.3005
R11905 gnd.n7474 gnd.n7375 9.3005
R11906 gnd.n7472 gnd.n7376 9.3005
R11907 gnd.n7471 gnd.n7377 9.3005
R11908 gnd.n7469 gnd.n7378 9.3005
R11909 gnd.n7468 gnd.n7379 9.3005
R11910 gnd.n7466 gnd.n7380 9.3005
R11911 gnd.n7465 gnd.n7381 9.3005
R11912 gnd.n7463 gnd.n7382 9.3005
R11913 gnd.n7462 gnd.n7383 9.3005
R11914 gnd.n7460 gnd.n7384 9.3005
R11915 gnd.n7459 gnd.n7385 9.3005
R11916 gnd.n7457 gnd.n7386 9.3005
R11917 gnd.n7456 gnd.n7387 9.3005
R11918 gnd.n7454 gnd.n7388 9.3005
R11919 gnd.n7453 gnd.n7389 9.3005
R11920 gnd.n7451 gnd.n7390 9.3005
R11921 gnd.n7450 gnd.n7391 9.3005
R11922 gnd.n7405 gnd.n7404 9.3005
R11923 gnd.n7407 gnd.n7406 9.3005
R11924 gnd.n7410 gnd.n7401 9.3005
R11925 gnd.n7414 gnd.n7413 9.3005
R11926 gnd.n7415 gnd.n7400 9.3005
R11927 gnd.n7417 gnd.n7416 9.3005
R11928 gnd.n7420 gnd.n7399 9.3005
R11929 gnd.n7424 gnd.n7423 9.3005
R11930 gnd.n7425 gnd.n7398 9.3005
R11931 gnd.n7427 gnd.n7426 9.3005
R11932 gnd.n7430 gnd.n7397 9.3005
R11933 gnd.n7434 gnd.n7433 9.3005
R11934 gnd.n7435 gnd.n7396 9.3005
R11935 gnd.n7437 gnd.n7436 9.3005
R11936 gnd.n7440 gnd.n7395 9.3005
R11937 gnd.n7444 gnd.n7443 9.3005
R11938 gnd.n7445 gnd.n7394 9.3005
R11939 gnd.n7447 gnd.n7446 9.3005
R11940 gnd.n7402 gnd.n348 9.3005
R11941 gnd.n249 gnd.n248 9.3005
R11942 gnd.n7657 gnd.n290 9.3005
R11943 gnd.n7656 gnd.n291 9.3005
R11944 gnd.n7655 gnd.n292 9.3005
R11945 gnd.n7652 gnd.n293 9.3005
R11946 gnd.n7651 gnd.n294 9.3005
R11947 gnd.n7648 gnd.n295 9.3005
R11948 gnd.n7647 gnd.n296 9.3005
R11949 gnd.n7644 gnd.n297 9.3005
R11950 gnd.n7643 gnd.n298 9.3005
R11951 gnd.n7640 gnd.n299 9.3005
R11952 gnd.n7639 gnd.n300 9.3005
R11953 gnd.n7636 gnd.n301 9.3005
R11954 gnd.n7635 gnd.n302 9.3005
R11955 gnd.n7632 gnd.n303 9.3005
R11956 gnd.n7631 gnd.n304 9.3005
R11957 gnd.n7628 gnd.n305 9.3005
R11958 gnd.n7624 gnd.n306 9.3005
R11959 gnd.n7621 gnd.n307 9.3005
R11960 gnd.n7620 gnd.n308 9.3005
R11961 gnd.n7617 gnd.n309 9.3005
R11962 gnd.n7616 gnd.n310 9.3005
R11963 gnd.n7613 gnd.n311 9.3005
R11964 gnd.n7612 gnd.n312 9.3005
R11965 gnd.n7609 gnd.n313 9.3005
R11966 gnd.n7608 gnd.n314 9.3005
R11967 gnd.n7605 gnd.n315 9.3005
R11968 gnd.n7604 gnd.n316 9.3005
R11969 gnd.n7601 gnd.n317 9.3005
R11970 gnd.n7600 gnd.n318 9.3005
R11971 gnd.n7597 gnd.n319 9.3005
R11972 gnd.n7596 gnd.n320 9.3005
R11973 gnd.n7593 gnd.n321 9.3005
R11974 gnd.n7592 gnd.n322 9.3005
R11975 gnd.n7589 gnd.n323 9.3005
R11976 gnd.n7588 gnd.n324 9.3005
R11977 gnd.n7585 gnd.n7584 9.3005
R11978 gnd.n7583 gnd.n325 9.3005
R11979 gnd.n7582 gnd.n7581 9.3005
R11980 gnd.n7578 gnd.n328 9.3005
R11981 gnd.n7575 gnd.n329 9.3005
R11982 gnd.n7574 gnd.n330 9.3005
R11983 gnd.n7571 gnd.n331 9.3005
R11984 gnd.n7570 gnd.n332 9.3005
R11985 gnd.n7567 gnd.n333 9.3005
R11986 gnd.n7566 gnd.n334 9.3005
R11987 gnd.n7563 gnd.n335 9.3005
R11988 gnd.n7562 gnd.n336 9.3005
R11989 gnd.n7559 gnd.n337 9.3005
R11990 gnd.n7558 gnd.n338 9.3005
R11991 gnd.n7555 gnd.n339 9.3005
R11992 gnd.n7554 gnd.n340 9.3005
R11993 gnd.n7551 gnd.n341 9.3005
R11994 gnd.n7550 gnd.n342 9.3005
R11995 gnd.n7547 gnd.n343 9.3005
R11996 gnd.n7546 gnd.n344 9.3005
R11997 gnd.n7543 gnd.n7542 9.3005
R11998 gnd.n7541 gnd.n345 9.3005
R11999 gnd.n7663 gnd.n7662 9.3005
R12000 gnd.n7065 gnd.n7064 9.3005
R12001 gnd.n581 gnd.n576 9.3005
R12002 gnd.n580 gnd.n579 9.3005
R12003 gnd.n552 gnd.n537 9.3005
R12004 gnd.n7116 gnd.n538 9.3005
R12005 gnd.n7115 gnd.n539 9.3005
R12006 gnd.n7114 gnd.n540 9.3005
R12007 gnd.n7113 gnd.n541 9.3005
R12008 gnd.n7091 gnd.n502 9.3005
R12009 gnd.n7151 gnd.n503 9.3005
R12010 gnd.n7150 gnd.n504 9.3005
R12011 gnd.n7149 gnd.n7148 9.3005
R12012 gnd.n505 gnd.n472 9.3005
R12013 gnd.n7186 gnd.n473 9.3005
R12014 gnd.n7185 gnd.n474 9.3005
R12015 gnd.n7184 gnd.n475 9.3005
R12016 gnd.n7183 gnd.n476 9.3005
R12017 gnd.n448 gnd.n445 9.3005
R12018 gnd.n7226 gnd.n446 9.3005
R12019 gnd.n7225 gnd.n7222 9.3005
R12020 gnd.n7224 gnd.n7223 9.3005
R12021 gnd.n421 gnd.n417 9.3005
R12022 gnd.n7273 gnd.n418 9.3005
R12023 gnd.n7272 gnd.n419 9.3005
R12024 gnd.n7271 gnd.n7266 9.3005
R12025 gnd.n7270 gnd.n7267 9.3005
R12026 gnd.n392 gnd.n391 9.3005
R12027 gnd.n7305 gnd.n7303 9.3005
R12028 gnd.n7304 gnd.n375 9.3005
R12029 gnd.n7326 gnd.n374 9.3005
R12030 gnd.n7328 gnd.n7327 9.3005
R12031 gnd.n364 gnd.n363 9.3005
R12032 gnd.n7341 gnd.n7340 9.3005
R12033 gnd.n355 gnd.n354 9.3005
R12034 gnd.n7356 gnd.n7355 9.3005
R12035 gnd.n7357 gnd.n123 9.3005
R12036 gnd.n7744 gnd.n124 9.3005
R12037 gnd.n7743 gnd.n125 9.3005
R12038 gnd.n7742 gnd.n126 9.3005
R12039 gnd.n7494 gnd.n127 9.3005
R12040 gnd.n7732 gnd.n141 9.3005
R12041 gnd.n7731 gnd.n142 9.3005
R12042 gnd.n7730 gnd.n143 9.3005
R12043 gnd.n7501 gnd.n144 9.3005
R12044 gnd.n7720 gnd.n161 9.3005
R12045 gnd.n7719 gnd.n162 9.3005
R12046 gnd.n7718 gnd.n163 9.3005
R12047 gnd.n7508 gnd.n164 9.3005
R12048 gnd.n7708 gnd.n179 9.3005
R12049 gnd.n7707 gnd.n180 9.3005
R12050 gnd.n7706 gnd.n181 9.3005
R12051 gnd.n7515 gnd.n182 9.3005
R12052 gnd.n7696 gnd.n199 9.3005
R12053 gnd.n7695 gnd.n200 9.3005
R12054 gnd.n7694 gnd.n201 9.3005
R12055 gnd.n7522 gnd.n202 9.3005
R12056 gnd.n7684 gnd.n217 9.3005
R12057 gnd.n7683 gnd.n218 9.3005
R12058 gnd.n7682 gnd.n219 9.3005
R12059 gnd.n7529 gnd.n220 9.3005
R12060 gnd.n7672 gnd.n237 9.3005
R12061 gnd.n7671 gnd.n238 9.3005
R12062 gnd.n7670 gnd.n239 9.3005
R12063 gnd.n7539 gnd.n240 9.3005
R12064 gnd.n7066 gnd.n575 9.3005
R12065 gnd.n7064 gnd.n7063 9.3005
R12066 gnd.n7062 gnd.n581 9.3005
R12067 gnd.n580 gnd.n551 9.3005
R12068 gnd.n7089 gnd.n552 9.3005
R12069 gnd.n7090 gnd.n538 9.3005
R12070 gnd.n7097 gnd.n539 9.3005
R12071 gnd.n7096 gnd.n540 9.3005
R12072 gnd.n7095 gnd.n541 9.3005
R12073 gnd.n7094 gnd.n7091 9.3005
R12074 gnd.n7092 gnd.n503 9.3005
R12075 gnd.n507 gnd.n504 9.3005
R12076 gnd.n7148 gnd.n7147 9.3005
R12077 gnd.n7146 gnd.n505 9.3005
R12078 gnd.n512 gnd.n473 9.3005
R12079 gnd.n511 gnd.n474 9.3005
R12080 gnd.n508 gnd.n475 9.3005
R12081 gnd.n476 gnd.n447 9.3005
R12082 gnd.n7218 gnd.n448 9.3005
R12083 gnd.n7219 gnd.n446 9.3005
R12084 gnd.n7222 gnd.n7221 9.3005
R12085 gnd.n7223 gnd.n420 9.3005
R12086 gnd.n7260 gnd.n421 9.3005
R12087 gnd.n7261 gnd.n418 9.3005
R12088 gnd.n7264 gnd.n419 9.3005
R12089 gnd.n7266 gnd.n7265 9.3005
R12090 gnd.n7267 gnd.n393 9.3005
R12091 gnd.n7301 gnd.n392 9.3005
R12092 gnd.n7303 gnd.n7302 9.3005
R12093 gnd.n376 gnd.n375 9.3005
R12094 gnd.n7326 gnd.n7325 9.3005
R12095 gnd.n7327 gnd.n365 9.3005
R12096 gnd.n7337 gnd.n364 9.3005
R12097 gnd.n7340 gnd.n7339 9.3005
R12098 gnd.n7338 gnd.n354 9.3005
R12099 gnd.n7356 gnd.n353 9.3005
R12100 gnd.n7358 gnd.n7357 9.3005
R12101 gnd.n349 gnd.n124 9.3005
R12102 gnd.n7492 gnd.n125 9.3005
R12103 gnd.n7493 gnd.n126 9.3005
R12104 gnd.n7496 gnd.n7494 9.3005
R12105 gnd.n7497 gnd.n141 9.3005
R12106 gnd.n7499 gnd.n142 9.3005
R12107 gnd.n7500 gnd.n143 9.3005
R12108 gnd.n7503 gnd.n7501 9.3005
R12109 gnd.n7504 gnd.n161 9.3005
R12110 gnd.n7506 gnd.n162 9.3005
R12111 gnd.n7507 gnd.n163 9.3005
R12112 gnd.n7510 gnd.n7508 9.3005
R12113 gnd.n7511 gnd.n179 9.3005
R12114 gnd.n7513 gnd.n180 9.3005
R12115 gnd.n7514 gnd.n181 9.3005
R12116 gnd.n7517 gnd.n7515 9.3005
R12117 gnd.n7518 gnd.n199 9.3005
R12118 gnd.n7520 gnd.n200 9.3005
R12119 gnd.n7521 gnd.n201 9.3005
R12120 gnd.n7524 gnd.n7522 9.3005
R12121 gnd.n7525 gnd.n217 9.3005
R12122 gnd.n7527 gnd.n218 9.3005
R12123 gnd.n7528 gnd.n219 9.3005
R12124 gnd.n7531 gnd.n7529 9.3005
R12125 gnd.n7532 gnd.n237 9.3005
R12126 gnd.n7534 gnd.n238 9.3005
R12127 gnd.n7535 gnd.n239 9.3005
R12128 gnd.n7539 gnd.n7538 9.3005
R12129 gnd.n582 gnd.n575 9.3005
R12130 gnd.n6929 gnd.n6928 9.3005
R12131 gnd.n6932 gnd.n690 9.3005
R12132 gnd.n6933 gnd.n689 9.3005
R12133 gnd.n6936 gnd.n688 9.3005
R12134 gnd.n6937 gnd.n687 9.3005
R12135 gnd.n6940 gnd.n686 9.3005
R12136 gnd.n6941 gnd.n685 9.3005
R12137 gnd.n6944 gnd.n684 9.3005
R12138 gnd.n6945 gnd.n683 9.3005
R12139 gnd.n6948 gnd.n682 9.3005
R12140 gnd.n6949 gnd.n681 9.3005
R12141 gnd.n6952 gnd.n680 9.3005
R12142 gnd.n6953 gnd.n679 9.3005
R12143 gnd.n6956 gnd.n678 9.3005
R12144 gnd.n6957 gnd.n677 9.3005
R12145 gnd.n6960 gnd.n676 9.3005
R12146 gnd.n6961 gnd.n675 9.3005
R12147 gnd.n6964 gnd.n674 9.3005
R12148 gnd.n6965 gnd.n673 9.3005
R12149 gnd.n6968 gnd.n672 9.3005
R12150 gnd.n6972 gnd.n668 9.3005
R12151 gnd.n6973 gnd.n667 9.3005
R12152 gnd.n6976 gnd.n666 9.3005
R12153 gnd.n6977 gnd.n665 9.3005
R12154 gnd.n6980 gnd.n664 9.3005
R12155 gnd.n6981 gnd.n663 9.3005
R12156 gnd.n6984 gnd.n662 9.3005
R12157 gnd.n6985 gnd.n661 9.3005
R12158 gnd.n6988 gnd.n660 9.3005
R12159 gnd.n6990 gnd.n656 9.3005
R12160 gnd.n6993 gnd.n655 9.3005
R12161 gnd.n6994 gnd.n654 9.3005
R12162 gnd.n6997 gnd.n653 9.3005
R12163 gnd.n6998 gnd.n652 9.3005
R12164 gnd.n7001 gnd.n651 9.3005
R12165 gnd.n7002 gnd.n650 9.3005
R12166 gnd.n7005 gnd.n649 9.3005
R12167 gnd.n7007 gnd.n646 9.3005
R12168 gnd.n7010 gnd.n645 9.3005
R12169 gnd.n7011 gnd.n644 9.3005
R12170 gnd.n7014 gnd.n643 9.3005
R12171 gnd.n7015 gnd.n642 9.3005
R12172 gnd.n7018 gnd.n641 9.3005
R12173 gnd.n7019 gnd.n640 9.3005
R12174 gnd.n7022 gnd.n639 9.3005
R12175 gnd.n7023 gnd.n638 9.3005
R12176 gnd.n7026 gnd.n637 9.3005
R12177 gnd.n7027 gnd.n636 9.3005
R12178 gnd.n7030 gnd.n635 9.3005
R12179 gnd.n7031 gnd.n634 9.3005
R12180 gnd.n7034 gnd.n633 9.3005
R12181 gnd.n7036 gnd.n632 9.3005
R12182 gnd.n7037 gnd.n631 9.3005
R12183 gnd.n7038 gnd.n630 9.3005
R12184 gnd.n629 gnd.n567 9.3005
R12185 gnd.n6969 gnd.n669 9.3005
R12186 gnd.n6927 gnd.n692 9.3005
R12187 gnd.n7072 gnd.n566 9.3005
R12188 gnd.n7076 gnd.n7073 9.3005
R12189 gnd.n7075 gnd.n7074 9.3005
R12190 gnd.n529 gnd.n528 9.3005
R12191 gnd.n7121 gnd.n7120 9.3005
R12192 gnd.n7122 gnd.n527 9.3005
R12193 gnd.n7126 gnd.n7123 9.3005
R12194 gnd.n7125 gnd.n7124 9.3005
R12195 gnd.n495 gnd.n494 9.3005
R12196 gnd.n7156 gnd.n7155 9.3005
R12197 gnd.n7157 gnd.n493 9.3005
R12198 gnd.n7159 gnd.n7158 9.3005
R12199 gnd.n464 gnd.n463 9.3005
R12200 gnd.n7191 gnd.n7190 9.3005
R12201 gnd.n7192 gnd.n462 9.3005
R12202 gnd.n7196 gnd.n7193 9.3005
R12203 gnd.n7195 gnd.n7194 9.3005
R12204 gnd.n437 gnd.n436 9.3005
R12205 gnd.n7231 gnd.n7230 9.3005
R12206 gnd.n7232 gnd.n435 9.3005
R12207 gnd.n7234 gnd.n7233 9.3005
R12208 gnd.n410 gnd.n409 9.3005
R12209 gnd.n7278 gnd.n7277 9.3005
R12210 gnd.n7279 gnd.n408 9.3005
R12211 gnd.n7283 gnd.n7280 9.3005
R12212 gnd.n7282 gnd.n109 9.3005
R12213 gnd.n114 gnd.n108 9.3005
R12214 gnd.n7738 gnd.n133 9.3005
R12215 gnd.n7737 gnd.n134 9.3005
R12216 gnd.n7736 gnd.n135 9.3005
R12217 gnd.n150 gnd.n136 9.3005
R12218 gnd.n7726 gnd.n151 9.3005
R12219 gnd.n7725 gnd.n152 9.3005
R12220 gnd.n7724 gnd.n153 9.3005
R12221 gnd.n170 gnd.n154 9.3005
R12222 gnd.n7714 gnd.n171 9.3005
R12223 gnd.n7713 gnd.n172 9.3005
R12224 gnd.n7712 gnd.n173 9.3005
R12225 gnd.n188 gnd.n174 9.3005
R12226 gnd.n7702 gnd.n189 9.3005
R12227 gnd.n7701 gnd.n190 9.3005
R12228 gnd.n7700 gnd.n191 9.3005
R12229 gnd.n208 gnd.n192 9.3005
R12230 gnd.n7690 gnd.n209 9.3005
R12231 gnd.n7689 gnd.n210 9.3005
R12232 gnd.n7688 gnd.n211 9.3005
R12233 gnd.n227 gnd.n212 9.3005
R12234 gnd.n7678 gnd.n228 9.3005
R12235 gnd.n7677 gnd.n229 9.3005
R12236 gnd.n7676 gnd.n230 9.3005
R12237 gnd.n246 gnd.n231 9.3005
R12238 gnd.n7666 gnd.n247 9.3005
R12239 gnd.n7665 gnd.n7664 9.3005
R12240 gnd.n7071 gnd.n7070 9.3005
R12241 gnd.n7749 gnd.n7748 9.3005
R12242 gnd.n1957 gnd.n1919 9.3005
R12243 gnd.n1922 gnd.n1920 9.3005
R12244 gnd.n1953 gnd.n1923 9.3005
R12245 gnd.n1952 gnd.n1924 9.3005
R12246 gnd.n1951 gnd.n1925 9.3005
R12247 gnd.n1928 gnd.n1926 9.3005
R12248 gnd.n1947 gnd.n1929 9.3005
R12249 gnd.n1946 gnd.n1930 9.3005
R12250 gnd.n1945 gnd.n1931 9.3005
R12251 gnd.n1934 gnd.n1932 9.3005
R12252 gnd.n1941 gnd.n1935 9.3005
R12253 gnd.n1940 gnd.n1936 9.3005
R12254 gnd.n1939 gnd.n1938 9.3005
R12255 gnd.n1937 gnd.n1549 9.3005
R12256 gnd.n1547 gnd.n1546 9.3005
R12257 gnd.n5392 gnd.n5391 9.3005
R12258 gnd.n5393 gnd.n1545 9.3005
R12259 gnd.n5400 gnd.n5394 9.3005
R12260 gnd.n5399 gnd.n5395 9.3005
R12261 gnd.n5398 gnd.n5396 9.3005
R12262 gnd.n1496 gnd.n1495 9.3005
R12263 gnd.n5456 gnd.n5455 9.3005
R12264 gnd.n5457 gnd.n1494 9.3005
R12265 gnd.n5459 gnd.n5458 9.3005
R12266 gnd.n1492 gnd.n1491 9.3005
R12267 gnd.n5464 gnd.n5463 9.3005
R12268 gnd.n5465 gnd.n1490 9.3005
R12269 gnd.n5695 gnd.n5466 9.3005
R12270 gnd.n5694 gnd.n5467 9.3005
R12271 gnd.n5693 gnd.n5468 9.3005
R12272 gnd.n5471 gnd.n5469 9.3005
R12273 gnd.n5687 gnd.n5472 9.3005
R12274 gnd.n5686 gnd.n5473 9.3005
R12275 gnd.n5685 gnd.n5474 9.3005
R12276 gnd.n5546 gnd.n5475 9.3005
R12277 gnd.n5548 gnd.n5547 9.3005
R12278 gnd.n5571 gnd.n5570 9.3005
R12279 gnd.n5572 gnd.n5545 9.3005
R12280 gnd.n5574 gnd.n5573 9.3005
R12281 gnd.n5535 gnd.n5534 9.3005
R12282 gnd.n5592 gnd.n5591 9.3005
R12283 gnd.n5593 gnd.n5533 9.3005
R12284 gnd.n5595 gnd.n5594 9.3005
R12285 gnd.n5523 gnd.n5522 9.3005
R12286 gnd.n5613 gnd.n5612 9.3005
R12287 gnd.n5614 gnd.n5521 9.3005
R12288 gnd.n5616 gnd.n5615 9.3005
R12289 gnd.n5510 gnd.n5509 9.3005
R12290 gnd.n5642 gnd.n5641 9.3005
R12291 gnd.n5643 gnd.n5508 9.3005
R12292 gnd.n5650 gnd.n5644 9.3005
R12293 gnd.n5649 gnd.n5645 9.3005
R12294 gnd.n5648 gnd.n5646 9.3005
R12295 gnd.n1198 gnd.n1197 9.3005
R12296 gnd.n6157 gnd.n6156 9.3005
R12297 gnd.n6158 gnd.n1196 9.3005
R12298 gnd.n6160 gnd.n6159 9.3005
R12299 gnd.n1172 gnd.n1171 9.3005
R12300 gnd.n6198 gnd.n6197 9.3005
R12301 gnd.n6199 gnd.n1170 9.3005
R12302 gnd.n6205 gnd.n6200 9.3005
R12303 gnd.n6204 gnd.n6201 9.3005
R12304 gnd.n6203 gnd.n6202 9.3005
R12305 gnd.n1150 gnd.n1149 9.3005
R12306 gnd.n6226 gnd.n6225 9.3005
R12307 gnd.n6227 gnd.n1148 9.3005
R12308 gnd.n6230 gnd.n6229 9.3005
R12309 gnd.n6228 gnd.n1120 9.3005
R12310 gnd.n6284 gnd.n1121 9.3005
R12311 gnd.n6283 gnd.n1122 9.3005
R12312 gnd.n6282 gnd.n1124 9.3005
R12313 gnd.n1123 gnd.n1088 9.3005
R12314 gnd.n6346 gnd.n1089 9.3005
R12315 gnd.n6345 gnd.n1090 9.3005
R12316 gnd.n6344 gnd.n1092 9.3005
R12317 gnd.n1091 gnd.n1061 9.3005
R12318 gnd.n6384 gnd.n1062 9.3005
R12319 gnd.n6383 gnd.n1063 9.3005
R12320 gnd.n6382 gnd.n1065 9.3005
R12321 gnd.n1064 gnd.n1031 9.3005
R12322 gnd.n6423 gnd.n1032 9.3005
R12323 gnd.n6422 gnd.n1033 9.3005
R12324 gnd.n6421 gnd.n1034 9.3005
R12325 gnd.n1037 gnd.n1036 9.3005
R12326 gnd.n1035 gnd.n985 9.3005
R12327 gnd.n6487 gnd.n986 9.3005
R12328 gnd.n6486 gnd.n987 9.3005
R12329 gnd.n6485 gnd.n988 9.3005
R12330 gnd.n990 gnd.n989 9.3005
R12331 gnd.n943 gnd.n942 9.3005
R12332 gnd.n6542 gnd.n6541 9.3005
R12333 gnd.n6543 gnd.n941 9.3005
R12334 gnd.n6545 gnd.n6544 9.3005
R12335 gnd.n889 gnd.n888 9.3005
R12336 gnd.n6718 gnd.n6717 9.3005
R12337 gnd.n6719 gnd.n887 9.3005
R12338 gnd.n6723 gnd.n6720 9.3005
R12339 gnd.n6722 gnd.n6721 9.3005
R12340 gnd.n865 gnd.n864 9.3005
R12341 gnd.n6748 gnd.n6747 9.3005
R12342 gnd.n6749 gnd.n863 9.3005
R12343 gnd.n6753 gnd.n6750 9.3005
R12344 gnd.n6752 gnd.n6751 9.3005
R12345 gnd.n840 gnd.n839 9.3005
R12346 gnd.n6778 gnd.n6777 9.3005
R12347 gnd.n6779 gnd.n838 9.3005
R12348 gnd.n6783 gnd.n6780 9.3005
R12349 gnd.n6782 gnd.n6781 9.3005
R12350 gnd.n815 gnd.n814 9.3005
R12351 gnd.n6813 gnd.n6812 9.3005
R12352 gnd.n6814 gnd.n813 9.3005
R12353 gnd.n6819 gnd.n6815 9.3005
R12354 gnd.n6818 gnd.n6817 9.3005
R12355 gnd.n6816 gnd.n801 9.3005
R12356 gnd.n799 gnd.n798 9.3005
R12357 gnd.n6837 gnd.n6836 9.3005
R12358 gnd.n6838 gnd.n797 9.3005
R12359 gnd.n6842 gnd.n6839 9.3005
R12360 gnd.n6841 gnd.n6840 9.3005
R12361 gnd.n587 gnd.n586 9.3005
R12362 gnd.n7046 gnd.n7045 9.3005
R12363 gnd.n7047 gnd.n585 9.3005
R12364 gnd.n7057 gnd.n7048 9.3005
R12365 gnd.n7056 gnd.n7049 9.3005
R12366 gnd.n7055 gnd.n7050 9.3005
R12367 gnd.n7052 gnd.n7051 9.3005
R12368 gnd.n549 gnd.n548 9.3005
R12369 gnd.n7103 gnd.n7102 9.3005
R12370 gnd.n7104 gnd.n547 9.3005
R12371 gnd.n7108 gnd.n7105 9.3005
R12372 gnd.n7107 gnd.n7106 9.3005
R12373 gnd.n485 gnd.n484 9.3005
R12374 gnd.n7165 gnd.n7164 9.3005
R12375 gnd.n7166 gnd.n483 9.3005
R12376 gnd.n7168 gnd.n7167 9.3005
R12377 gnd.n481 gnd.n480 9.3005
R12378 gnd.n7173 gnd.n7172 9.3005
R12379 gnd.n7174 gnd.n479 9.3005
R12380 gnd.n7178 gnd.n7175 9.3005
R12381 gnd.n7177 gnd.n7176 9.3005
R12382 gnd.n429 gnd.n428 9.3005
R12383 gnd.n7240 gnd.n7239 9.3005
R12384 gnd.n7241 gnd.n427 9.3005
R12385 gnd.n7255 gnd.n7242 9.3005
R12386 gnd.n7254 gnd.n7243 9.3005
R12387 gnd.n7253 gnd.n7244 9.3005
R12388 gnd.n7246 gnd.n7245 9.3005
R12389 gnd.n7249 gnd.n7247 9.3005
R12390 gnd.n5235 gnd.n5234 9.3005
R12391 gnd.n4778 gnd.n4759 9.3005
R12392 gnd.n4776 gnd.n4760 9.3005
R12393 gnd.n4775 gnd.n4761 9.3005
R12394 gnd.n4773 gnd.n4762 9.3005
R12395 gnd.n4772 gnd.n4763 9.3005
R12396 gnd.n4770 gnd.n4764 9.3005
R12397 gnd.n4769 gnd.n4765 9.3005
R12398 gnd.n4767 gnd.n4766 9.3005
R12399 gnd.n1773 gnd.n1772 9.3005
R12400 gnd.n5100 gnd.n5099 9.3005
R12401 gnd.n5101 gnd.n1771 9.3005
R12402 gnd.n5105 gnd.n5102 9.3005
R12403 gnd.n5104 gnd.n5103 9.3005
R12404 gnd.n1748 gnd.n1747 9.3005
R12405 gnd.n5135 gnd.n5134 9.3005
R12406 gnd.n5136 gnd.n1746 9.3005
R12407 gnd.n5140 gnd.n5137 9.3005
R12408 gnd.n5139 gnd.n5138 9.3005
R12409 gnd.n1723 gnd.n1722 9.3005
R12410 gnd.n5170 gnd.n5169 9.3005
R12411 gnd.n5171 gnd.n1721 9.3005
R12412 gnd.n5175 gnd.n5172 9.3005
R12413 gnd.n5174 gnd.n5173 9.3005
R12414 gnd.n1696 gnd.n1695 9.3005
R12415 gnd.n5207 gnd.n5206 9.3005
R12416 gnd.n5208 gnd.n1694 9.3005
R12417 gnd.n5212 gnd.n5209 9.3005
R12418 gnd.n5211 gnd.n5210 9.3005
R12419 gnd.n1677 gnd.n1676 9.3005
R12420 gnd.n5232 gnd.n5231 9.3005
R12421 gnd.n5233 gnd.n1675 9.3005
R12422 gnd.n4780 gnd.n4779 9.3005
R12423 gnd.n4788 gnd.n4787 9.3005
R12424 gnd.n4789 gnd.n4755 9.3005
R12425 gnd.n4754 gnd.n4752 9.3005
R12426 gnd.n4795 gnd.n4751 9.3005
R12427 gnd.n4796 gnd.n4750 9.3005
R12428 gnd.n4797 gnd.n4749 9.3005
R12429 gnd.n4748 gnd.n4746 9.3005
R12430 gnd.n4803 gnd.n4745 9.3005
R12431 gnd.n4804 gnd.n4744 9.3005
R12432 gnd.n4805 gnd.n4743 9.3005
R12433 gnd.n4742 gnd.n4740 9.3005
R12434 gnd.n4811 gnd.n4739 9.3005
R12435 gnd.n4812 gnd.n4738 9.3005
R12436 gnd.n4813 gnd.n4737 9.3005
R12437 gnd.n4736 gnd.n4734 9.3005
R12438 gnd.n4819 gnd.n4733 9.3005
R12439 gnd.n4821 gnd.n4820 9.3005
R12440 gnd.n4786 gnd.n4758 9.3005
R12441 gnd.n4785 gnd.n4784 9.3005
R12442 gnd.n1364 gnd.n1362 9.3005
R12443 gnd.n5918 gnd.n5913 9.3005
R12444 gnd.n5919 gnd.n5912 9.3005
R12445 gnd.n5920 gnd.n5911 9.3005
R12446 gnd.n5910 gnd.n5907 9.3005
R12447 gnd.n5925 gnd.n5906 9.3005
R12448 gnd.n5926 gnd.n5905 9.3005
R12449 gnd.n5927 gnd.n5904 9.3005
R12450 gnd.n5903 gnd.n5897 9.3005
R12451 gnd.n5932 gnd.n5896 9.3005
R12452 gnd.n5933 gnd.n5895 9.3005
R12453 gnd.n5934 gnd.n5894 9.3005
R12454 gnd.n5893 gnd.n5890 9.3005
R12455 gnd.n5939 gnd.n5889 9.3005
R12456 gnd.n5940 gnd.n5888 9.3005
R12457 gnd.n5941 gnd.n5887 9.3005
R12458 gnd.n5886 gnd.n5883 9.3005
R12459 gnd.n5946 gnd.n5882 9.3005
R12460 gnd.n5947 gnd.n5881 9.3005
R12461 gnd.n5948 gnd.n5880 9.3005
R12462 gnd.n5879 gnd.n5876 9.3005
R12463 gnd.n5953 gnd.n5875 9.3005
R12464 gnd.n5954 gnd.n5874 9.3005
R12465 gnd.n5955 gnd.n5873 9.3005
R12466 gnd.n5871 gnd.n5870 9.3005
R12467 gnd.n5961 gnd.n5960 9.3005
R12468 gnd.n6028 gnd.n6027 9.3005
R12469 gnd.n1366 gnd.n1365 9.3005
R12470 gnd.n1372 gnd.n1370 9.3005
R12471 gnd.n6020 gnd.n1373 9.3005
R12472 gnd.n6019 gnd.n1374 9.3005
R12473 gnd.n6018 gnd.n1375 9.3005
R12474 gnd.n1379 gnd.n1376 9.3005
R12475 gnd.n6013 gnd.n1380 9.3005
R12476 gnd.n6012 gnd.n6011 9.3005
R12477 gnd.n6010 gnd.n1381 9.3005
R12478 gnd.n6009 gnd.n6008 9.3005
R12479 gnd.n1385 gnd.n1384 9.3005
R12480 gnd.n1390 gnd.n1388 9.3005
R12481 gnd.n6001 gnd.n1391 9.3005
R12482 gnd.n6000 gnd.n1392 9.3005
R12483 gnd.n5999 gnd.n1393 9.3005
R12484 gnd.n1397 gnd.n1394 9.3005
R12485 gnd.n5994 gnd.n1398 9.3005
R12486 gnd.n5993 gnd.n1399 9.3005
R12487 gnd.n5992 gnd.n1400 9.3005
R12488 gnd.n1404 gnd.n1401 9.3005
R12489 gnd.n5987 gnd.n1405 9.3005
R12490 gnd.n5986 gnd.n1406 9.3005
R12491 gnd.n5985 gnd.n1407 9.3005
R12492 gnd.n1411 gnd.n1408 9.3005
R12493 gnd.n5980 gnd.n1412 9.3005
R12494 gnd.n5979 gnd.n1413 9.3005
R12495 gnd.n5978 gnd.n1414 9.3005
R12496 gnd.n1420 gnd.n1417 9.3005
R12497 gnd.n5973 gnd.n5972 9.3005
R12498 gnd.n6029 gnd.n1361 9.3005
R12499 gnd.n5040 gnd.n5039 9.3005
R12500 gnd.n5036 gnd.n5035 9.3005
R12501 gnd.n1811 gnd.n1808 9.3005
R12502 gnd.n5061 gnd.n1809 9.3005
R12503 gnd.n5060 gnd.n5057 9.3005
R12504 gnd.n5059 gnd.n5058 9.3005
R12505 gnd.n1793 gnd.n1789 9.3005
R12506 gnd.n5085 gnd.n1790 9.3005
R12507 gnd.n5084 gnd.n1791 9.3005
R12508 gnd.n5083 gnd.n5079 9.3005
R12509 gnd.n5082 gnd.n5080 9.3005
R12510 gnd.n1767 gnd.n1763 9.3005
R12511 gnd.n5120 gnd.n1764 9.3005
R12512 gnd.n5119 gnd.n1765 9.3005
R12513 gnd.n5118 gnd.n5114 9.3005
R12514 gnd.n5117 gnd.n5115 9.3005
R12515 gnd.n1742 gnd.n1738 9.3005
R12516 gnd.n5155 gnd.n1739 9.3005
R12517 gnd.n5154 gnd.n1740 9.3005
R12518 gnd.n5153 gnd.n5149 9.3005
R12519 gnd.n5152 gnd.n5150 9.3005
R12520 gnd.n1717 gnd.n1711 9.3005
R12521 gnd.n5192 gnd.n1712 9.3005
R12522 gnd.n5191 gnd.n1713 9.3005
R12523 gnd.n5190 gnd.n1714 9.3005
R12524 gnd.n5189 gnd.n5188 9.3005
R12525 gnd.n1715 gnd.n1690 9.3005
R12526 gnd.n1682 gnd.n1681 9.3005
R12527 gnd.n5226 gnd.n5225 9.3005
R12528 gnd.n5227 gnd.n1665 9.3005
R12529 gnd.n5245 gnd.n1664 9.3005
R12530 gnd.n5247 gnd.n5246 9.3005
R12531 gnd.n5248 gnd.n1659 9.3005
R12532 gnd.n5254 gnd.n1658 9.3005
R12533 gnd.n5256 gnd.n5255 9.3005
R12534 gnd.n1644 gnd.n1640 9.3005
R12535 gnd.n5287 gnd.n1641 9.3005
R12536 gnd.n5286 gnd.n1642 9.3005
R12537 gnd.n5285 gnd.n5280 9.3005
R12538 gnd.n5284 gnd.n5281 9.3005
R12539 gnd.n1609 gnd.n1605 9.3005
R12540 gnd.n5323 gnd.n1606 9.3005
R12541 gnd.n5322 gnd.n1607 9.3005
R12542 gnd.n5321 gnd.n5316 9.3005
R12543 gnd.n5320 gnd.n5317 9.3005
R12544 gnd.n1580 gnd.n1574 9.3005
R12545 gnd.n5365 gnd.n1575 9.3005
R12546 gnd.n5364 gnd.n1576 9.3005
R12547 gnd.n5363 gnd.n1577 9.3005
R12548 gnd.n5362 gnd.n5360 9.3005
R12549 gnd.n1578 gnd.n1538 9.3005
R12550 gnd.n5408 gnd.n1539 9.3005
R12551 gnd.n5407 gnd.n1540 9.3005
R12552 gnd.n5406 gnd.n1541 9.3005
R12553 gnd.n5405 gnd.n1542 9.3005
R12554 gnd.n1514 gnd.n1511 9.3005
R12555 gnd.n5442 gnd.n1512 9.3005
R12556 gnd.n5441 gnd.n5438 9.3005
R12557 gnd.n5440 gnd.n5439 9.3005
R12558 gnd.n1443 gnd.n1442 9.3005
R12559 gnd.n5862 gnd.n5858 9.3005
R12560 gnd.n5861 gnd.n5859 9.3005
R12561 gnd.n5860 gnd.n1422 9.3005
R12562 gnd.n5970 gnd.n1423 9.3005
R12563 gnd.n5041 gnd.n5034 9.3005
R12564 gnd.n5039 gnd.n5038 9.3005
R12565 gnd.n5036 gnd.n1810 9.3005
R12566 gnd.n5054 gnd.n1811 9.3005
R12567 gnd.n5055 gnd.n1809 9.3005
R12568 gnd.n5057 gnd.n5056 9.3005
R12569 gnd.n5058 gnd.n1792 9.3005
R12570 gnd.n5074 gnd.n1793 9.3005
R12571 gnd.n5075 gnd.n1790 9.3005
R12572 gnd.n5077 gnd.n1791 9.3005
R12573 gnd.n5079 gnd.n5078 9.3005
R12574 gnd.n5080 gnd.n1766 9.3005
R12575 gnd.n5109 gnd.n1767 9.3005
R12576 gnd.n5110 gnd.n1764 9.3005
R12577 gnd.n5112 gnd.n1765 9.3005
R12578 gnd.n5114 gnd.n5113 9.3005
R12579 gnd.n5115 gnd.n1741 9.3005
R12580 gnd.n5144 gnd.n1742 9.3005
R12581 gnd.n5145 gnd.n1739 9.3005
R12582 gnd.n5147 gnd.n1740 9.3005
R12583 gnd.n5149 gnd.n5148 9.3005
R12584 gnd.n5150 gnd.n1716 9.3005
R12585 gnd.n5179 gnd.n1717 9.3005
R12586 gnd.n5180 gnd.n1712 9.3005
R12587 gnd.n5182 gnd.n1713 9.3005
R12588 gnd.n5183 gnd.n1714 9.3005
R12589 gnd.n5188 gnd.n5187 9.3005
R12590 gnd.n5184 gnd.n1715 9.3005
R12591 gnd.n1683 gnd.n1682 9.3005
R12592 gnd.n5225 gnd.n5224 9.3005
R12593 gnd.n1666 gnd.n1665 9.3005
R12594 gnd.n5245 gnd.n5244 9.3005
R12595 gnd.n5246 gnd.n1660 9.3005
R12596 gnd.n5252 gnd.n1659 9.3005
R12597 gnd.n5254 gnd.n5253 9.3005
R12598 gnd.n5255 gnd.n1643 9.3005
R12599 gnd.n5274 gnd.n1644 9.3005
R12600 gnd.n5275 gnd.n1641 9.3005
R12601 gnd.n5278 gnd.n1642 9.3005
R12602 gnd.n5280 gnd.n5279 9.3005
R12603 gnd.n5281 gnd.n1608 9.3005
R12604 gnd.n5310 gnd.n1609 9.3005
R12605 gnd.n5311 gnd.n1606 9.3005
R12606 gnd.n5314 gnd.n1607 9.3005
R12607 gnd.n5316 gnd.n5315 9.3005
R12608 gnd.n5317 gnd.n1579 9.3005
R12609 gnd.n5346 gnd.n1580 9.3005
R12610 gnd.n5347 gnd.n1575 9.3005
R12611 gnd.n5350 gnd.n1576 9.3005
R12612 gnd.n5351 gnd.n1577 9.3005
R12613 gnd.n5360 gnd.n5359 9.3005
R12614 gnd.n5357 gnd.n1578 9.3005
R12615 gnd.n5356 gnd.n1539 9.3005
R12616 gnd.n5355 gnd.n1540 9.3005
R12617 gnd.n5352 gnd.n1541 9.3005
R12618 gnd.n1542 gnd.n1513 9.3005
R12619 gnd.n5434 gnd.n1514 9.3005
R12620 gnd.n5435 gnd.n1512 9.3005
R12621 gnd.n5438 gnd.n5437 9.3005
R12622 gnd.n5439 gnd.n1444 9.3005
R12623 gnd.n5856 gnd.n1443 9.3005
R12624 gnd.n5858 gnd.n5857 9.3005
R12625 gnd.n5859 gnd.n1424 9.3005
R12626 gnd.n5968 gnd.n1422 9.3005
R12627 gnd.n5970 gnd.n5969 9.3005
R12628 gnd.n5037 gnd.n5034 9.3005
R12629 gnd.n4825 gnd.n4822 9.3005
R12630 gnd.n5022 gnd.n4826 9.3005
R12631 gnd.n5024 gnd.n5023 9.3005
R12632 gnd.n5021 gnd.n4828 9.3005
R12633 gnd.n5020 gnd.n5019 9.3005
R12634 gnd.n4830 gnd.n4829 9.3005
R12635 gnd.n5013 gnd.n5012 9.3005
R12636 gnd.n5011 gnd.n4832 9.3005
R12637 gnd.n5010 gnd.n5009 9.3005
R12638 gnd.n4834 gnd.n4833 9.3005
R12639 gnd.n5003 gnd.n5002 9.3005
R12640 gnd.n5001 gnd.n4836 9.3005
R12641 gnd.n5000 gnd.n4999 9.3005
R12642 gnd.n4838 gnd.n4837 9.3005
R12643 gnd.n4993 gnd.n4992 9.3005
R12644 gnd.n4991 gnd.n4840 9.3005
R12645 gnd.n4990 gnd.n4989 9.3005
R12646 gnd.n4842 gnd.n4841 9.3005
R12647 gnd.n4983 gnd.n4982 9.3005
R12648 gnd.n4981 gnd.n4844 9.3005
R12649 gnd.n4846 gnd.n4845 9.3005
R12650 gnd.n4971 gnd.n4970 9.3005
R12651 gnd.n4969 gnd.n4848 9.3005
R12652 gnd.n4968 gnd.n4967 9.3005
R12653 gnd.n4850 gnd.n4849 9.3005
R12654 gnd.n4961 gnd.n4960 9.3005
R12655 gnd.n4959 gnd.n4852 9.3005
R12656 gnd.n4958 gnd.n4957 9.3005
R12657 gnd.n4854 gnd.n4853 9.3005
R12658 gnd.n4951 gnd.n4950 9.3005
R12659 gnd.n4949 gnd.n4856 9.3005
R12660 gnd.n4948 gnd.n4947 9.3005
R12661 gnd.n4858 gnd.n4857 9.3005
R12662 gnd.n4941 gnd.n4940 9.3005
R12663 gnd.n4939 gnd.n4860 9.3005
R12664 gnd.n4938 gnd.n4937 9.3005
R12665 gnd.n4862 gnd.n4861 9.3005
R12666 gnd.n4931 gnd.n4930 9.3005
R12667 gnd.n4929 gnd.n4864 9.3005
R12668 gnd.n4928 gnd.n4927 9.3005
R12669 gnd.n4866 gnd.n4865 9.3005
R12670 gnd.n4921 gnd.n4920 9.3005
R12671 gnd.n4919 gnd.n4871 9.3005
R12672 gnd.n4918 gnd.n4917 9.3005
R12673 gnd.n4873 gnd.n4872 9.3005
R12674 gnd.n4911 gnd.n4910 9.3005
R12675 gnd.n4909 gnd.n4875 9.3005
R12676 gnd.n4908 gnd.n4907 9.3005
R12677 gnd.n4877 gnd.n4876 9.3005
R12678 gnd.n4901 gnd.n4900 9.3005
R12679 gnd.n4899 gnd.n4879 9.3005
R12680 gnd.n4898 gnd.n4897 9.3005
R12681 gnd.n4881 gnd.n4880 9.3005
R12682 gnd.n4891 gnd.n4890 9.3005
R12683 gnd.n4889 gnd.n4883 9.3005
R12684 gnd.n4888 gnd.n4887 9.3005
R12685 gnd.n4884 gnd.n1817 9.3005
R12686 gnd.n4980 gnd.n4979 9.3005
R12687 gnd.n5032 gnd.n5031 9.3005
R12688 gnd.n5047 gnd.n1816 9.3005
R12689 gnd.n5049 gnd.n5048 9.3005
R12690 gnd.n1801 gnd.n1800 9.3005
R12691 gnd.n5066 gnd.n5065 9.3005
R12692 gnd.n5067 gnd.n1799 9.3005
R12693 gnd.n5069 gnd.n5068 9.3005
R12694 gnd.n1781 gnd.n1780 9.3005
R12695 gnd.n5090 gnd.n5089 9.3005
R12696 gnd.n5091 gnd.n1779 9.3005
R12697 gnd.n5095 gnd.n5092 9.3005
R12698 gnd.n5094 gnd.n5093 9.3005
R12699 gnd.n1756 gnd.n1755 9.3005
R12700 gnd.n5125 gnd.n5124 9.3005
R12701 gnd.n5126 gnd.n1754 9.3005
R12702 gnd.n5130 gnd.n5127 9.3005
R12703 gnd.n5129 gnd.n5128 9.3005
R12704 gnd.n1732 gnd.n1731 9.3005
R12705 gnd.n5160 gnd.n5159 9.3005
R12706 gnd.n5161 gnd.n1730 9.3005
R12707 gnd.n5165 gnd.n5162 9.3005
R12708 gnd.n5164 gnd.n5163 9.3005
R12709 gnd.n1705 gnd.n1704 9.3005
R12710 gnd.n5197 gnd.n5196 9.3005
R12711 gnd.n5198 gnd.n1703 9.3005
R12712 gnd.n5202 gnd.n5199 9.3005
R12713 gnd.n5201 gnd.n1625 9.3005
R12714 gnd.n5293 gnd.n1624 9.3005
R12715 gnd.n5297 gnd.n5294 9.3005
R12716 gnd.n5296 gnd.n5295 9.3005
R12717 gnd.n1597 gnd.n1596 9.3005
R12718 gnd.n5328 gnd.n5327 9.3005
R12719 gnd.n5329 gnd.n1595 9.3005
R12720 gnd.n5333 gnd.n5330 9.3005
R12721 gnd.n5332 gnd.n5331 9.3005
R12722 gnd.n1566 gnd.n1565 9.3005
R12723 gnd.n5370 gnd.n5369 9.3005
R12724 gnd.n5371 gnd.n1564 9.3005
R12725 gnd.n5375 gnd.n5372 9.3005
R12726 gnd.n5374 gnd.n5373 9.3005
R12727 gnd.n1530 gnd.n1529 9.3005
R12728 gnd.n5413 gnd.n5412 9.3005
R12729 gnd.n5414 gnd.n1528 9.3005
R12730 gnd.n5418 gnd.n5415 9.3005
R12731 gnd.n5417 gnd.n5416 9.3005
R12732 gnd.n1503 gnd.n1502 9.3005
R12733 gnd.n5447 gnd.n5446 9.3005
R12734 gnd.n5448 gnd.n1501 9.3005
R12735 gnd.n5450 gnd.n5449 9.3005
R12736 gnd.n1434 gnd.n1433 9.3005
R12737 gnd.n5867 gnd.n5866 9.3005
R12738 gnd.n5868 gnd.n1432 9.3005
R12739 gnd.n5964 gnd.n5869 9.3005
R12740 gnd.n5963 gnd.n5962 9.3005
R12741 gnd.n5046 gnd.n5045 9.3005
R12742 gnd.n5292 gnd.n5291 9.3005
R12743 gnd.n1970 gnd.n1626 9.3005
R12744 gnd.n1958 gnd.n1626 9.3005
R12745 gnd.n3320 gnd.n3317 9.3005
R12746 gnd.n3316 gnd.n1975 9.3005
R12747 gnd.n3315 gnd.n3314 9.3005
R12748 gnd.n1977 gnd.n1976 9.3005
R12749 gnd.n3308 gnd.n3307 9.3005
R12750 gnd.n3306 gnd.n1981 9.3005
R12751 gnd.n3305 gnd.n3304 9.3005
R12752 gnd.n1983 gnd.n1982 9.3005
R12753 gnd.n3298 gnd.n3297 9.3005
R12754 gnd.n3296 gnd.n1987 9.3005
R12755 gnd.n3295 gnd.n3294 9.3005
R12756 gnd.n1989 gnd.n1988 9.3005
R12757 gnd.n3288 gnd.n3287 9.3005
R12758 gnd.n3286 gnd.n1993 9.3005
R12759 gnd.n3285 gnd.n3284 9.3005
R12760 gnd.n1995 gnd.n1994 9.3005
R12761 gnd.n3278 gnd.n3277 9.3005
R12762 gnd.n3276 gnd.n1999 9.3005
R12763 gnd.n3275 gnd.n3274 9.3005
R12764 gnd.n2001 gnd.n2000 9.3005
R12765 gnd.n3268 gnd.n3267 9.3005
R12766 gnd.n3266 gnd.n2005 9.3005
R12767 gnd.n3265 gnd.n3264 9.3005
R12768 gnd.n2007 gnd.n2006 9.3005
R12769 gnd.n3258 gnd.n3257 9.3005
R12770 gnd.n3256 gnd.n2011 9.3005
R12771 gnd.n3255 gnd.n3254 9.3005
R12772 gnd.n2013 gnd.n2012 9.3005
R12773 gnd.n3248 gnd.n3247 9.3005
R12774 gnd.n3246 gnd.n2017 9.3005
R12775 gnd.n3245 gnd.n3244 9.3005
R12776 gnd.n2019 gnd.n2018 9.3005
R12777 gnd.n3238 gnd.n3237 9.3005
R12778 gnd.n3236 gnd.n2023 9.3005
R12779 gnd.n3235 gnd.n3234 9.3005
R12780 gnd.n2025 gnd.n2024 9.3005
R12781 gnd.n3228 gnd.n3227 9.3005
R12782 gnd.n3226 gnd.n2029 9.3005
R12783 gnd.n3225 gnd.n3224 9.3005
R12784 gnd.n2031 gnd.n2030 9.3005
R12785 gnd.n3218 gnd.n3217 9.3005
R12786 gnd.n3216 gnd.n2035 9.3005
R12787 gnd.n3215 gnd.n3214 9.3005
R12788 gnd.n2037 gnd.n2036 9.3005
R12789 gnd.n3208 gnd.n3207 9.3005
R12790 gnd.n3206 gnd.n2041 9.3005
R12791 gnd.n3205 gnd.n3204 9.3005
R12792 gnd.n2043 gnd.n2042 9.3005
R12793 gnd.n3198 gnd.n3197 9.3005
R12794 gnd.n3196 gnd.n2047 9.3005
R12795 gnd.n3195 gnd.n3194 9.3005
R12796 gnd.n2049 gnd.n2048 9.3005
R12797 gnd.n3188 gnd.n3187 9.3005
R12798 gnd.n3186 gnd.n2053 9.3005
R12799 gnd.n3185 gnd.n3184 9.3005
R12800 gnd.n2055 gnd.n2054 9.3005
R12801 gnd.n3178 gnd.n3177 9.3005
R12802 gnd.n3176 gnd.n2059 9.3005
R12803 gnd.n3175 gnd.n3174 9.3005
R12804 gnd.n2061 gnd.n2060 9.3005
R12805 gnd.n3168 gnd.n3167 9.3005
R12806 gnd.n3166 gnd.n2065 9.3005
R12807 gnd.n3165 gnd.n3164 9.3005
R12808 gnd.n2067 gnd.n2066 9.3005
R12809 gnd.n3158 gnd.n3157 9.3005
R12810 gnd.n3156 gnd.n2071 9.3005
R12811 gnd.n3155 gnd.n3154 9.3005
R12812 gnd.n2073 gnd.n2072 9.3005
R12813 gnd.n3148 gnd.n3147 9.3005
R12814 gnd.n3146 gnd.n2077 9.3005
R12815 gnd.n3145 gnd.n3144 9.3005
R12816 gnd.n2079 gnd.n2078 9.3005
R12817 gnd.n3138 gnd.n3137 9.3005
R12818 gnd.n3136 gnd.n2083 9.3005
R12819 gnd.n3135 gnd.n3134 9.3005
R12820 gnd.n2085 gnd.n2084 9.3005
R12821 gnd.n3128 gnd.n3127 9.3005
R12822 gnd.n3126 gnd.n2089 9.3005
R12823 gnd.n3125 gnd.n3124 9.3005
R12824 gnd.n2091 gnd.n2090 9.3005
R12825 gnd.n3118 gnd.n3117 9.3005
R12826 gnd.n3116 gnd.n2095 9.3005
R12827 gnd.n3115 gnd.n3114 9.3005
R12828 gnd.n2097 gnd.n2096 9.3005
R12829 gnd.n3319 gnd.n3318 9.3005
R12830 gnd.n6865 gnd.n758 9.3005
R12831 gnd.n5556 gnd.n5553 9.3005
R12832 gnd.n5561 gnd.n5560 9.3005
R12833 gnd.n5562 gnd.n5552 9.3005
R12834 gnd.n5564 gnd.n5563 9.3005
R12835 gnd.n5541 gnd.n5540 9.3005
R12836 gnd.n5582 gnd.n5581 9.3005
R12837 gnd.n5583 gnd.n5539 9.3005
R12838 gnd.n5585 gnd.n5584 9.3005
R12839 gnd.n5529 gnd.n5528 9.3005
R12840 gnd.n5603 gnd.n5602 9.3005
R12841 gnd.n5604 gnd.n5527 9.3005
R12842 gnd.n5606 gnd.n5605 9.3005
R12843 gnd.n5517 gnd.n5516 9.3005
R12844 gnd.n5624 gnd.n5623 9.3005
R12845 gnd.n5625 gnd.n5514 9.3005
R12846 gnd.n5636 gnd.n5635 9.3005
R12847 gnd.n5634 gnd.n5515 9.3005
R12848 gnd.n5633 gnd.n5632 9.3005
R12849 gnd.n5631 gnd.n5626 9.3005
R12850 gnd.n5630 gnd.n5629 9.3005
R12851 gnd.n5628 gnd.n1216 9.3005
R12852 gnd.n6112 gnd.n1215 9.3005
R12853 gnd.n6114 gnd.n6113 9.3005
R12854 gnd.n6115 gnd.n1213 9.3005
R12855 gnd.n6143 gnd.n6142 9.3005
R12856 gnd.n6141 gnd.n1214 9.3005
R12857 gnd.n6140 gnd.n6139 9.3005
R12858 gnd.n6138 gnd.n6116 9.3005
R12859 gnd.n6137 gnd.n6136 9.3005
R12860 gnd.n6135 gnd.n6121 9.3005
R12861 gnd.n6134 gnd.n6133 9.3005
R12862 gnd.n6132 gnd.n6122 9.3005
R12863 gnd.n6131 gnd.n6130 9.3005
R12864 gnd.n6129 gnd.n6123 9.3005
R12865 gnd.n6128 gnd.n6127 9.3005
R12866 gnd.n6126 gnd.n6125 9.3005
R12867 gnd.n6124 gnd.n1097 9.3005
R12868 gnd.n6308 gnd.n1096 9.3005
R12869 gnd.n6310 gnd.n6309 9.3005
R12870 gnd.n6311 gnd.n1094 9.3005
R12871 gnd.n6339 gnd.n6338 9.3005
R12872 gnd.n6337 gnd.n1095 9.3005
R12873 gnd.n6336 gnd.n6335 9.3005
R12874 gnd.n6334 gnd.n6312 9.3005
R12875 gnd.n6333 gnd.n6332 9.3005
R12876 gnd.n6331 gnd.n6315 9.3005
R12877 gnd.n6330 gnd.n6329 9.3005
R12878 gnd.n6328 gnd.n6316 9.3005
R12879 gnd.n6327 gnd.n6326 9.3005
R12880 gnd.n6325 gnd.n6319 9.3005
R12881 gnd.n6324 gnd.n6323 9.3005
R12882 gnd.n6322 gnd.n6320 9.3005
R12883 gnd.n969 gnd.n968 9.3005
R12884 gnd.n6502 gnd.n6501 9.3005
R12885 gnd.n6503 gnd.n966 9.3005
R12886 gnd.n6505 gnd.n6504 9.3005
R12887 gnd.n6506 gnd.n965 9.3005
R12888 gnd.n6508 gnd.n6507 9.3005
R12889 gnd.n6509 gnd.n963 9.3005
R12890 gnd.n6516 gnd.n6515 9.3005
R12891 gnd.n6514 gnd.n964 9.3005
R12892 gnd.n6513 gnd.n6512 9.3005
R12893 gnd.n6511 gnd.n6510 9.3005
R12894 gnd.n871 gnd.n870 9.3005
R12895 gnd.n6738 gnd.n6737 9.3005
R12896 gnd.n6739 gnd.n868 9.3005
R12897 gnd.n6742 gnd.n6741 9.3005
R12898 gnd.n6740 gnd.n869 9.3005
R12899 gnd.n846 gnd.n845 9.3005
R12900 gnd.n6768 gnd.n6767 9.3005
R12901 gnd.n6769 gnd.n843 9.3005
R12902 gnd.n6772 gnd.n6771 9.3005
R12903 gnd.n6770 gnd.n844 9.3005
R12904 gnd.n822 gnd.n821 9.3005
R12905 gnd.n6798 gnd.n6797 9.3005
R12906 gnd.n6799 gnd.n819 9.3005
R12907 gnd.n6807 gnd.n6806 9.3005
R12908 gnd.n6805 gnd.n820 9.3005
R12909 gnd.n6804 gnd.n6803 9.3005
R12910 gnd.n6802 gnd.n6800 9.3005
R12911 gnd.n760 gnd.n759 9.3005
R12912 gnd.n6864 gnd.n6863 9.3005
R12913 gnd.n5555 gnd.n5554 9.3005
R12914 gnd.n5841 gnd.n1455 9.3005
R12915 gnd.n1650 gnd.n1649 9.3005
R12916 gnd.n5266 gnd.n5265 9.3005
R12917 gnd.n5267 gnd.n1647 9.3005
R12918 gnd.n5270 gnd.n5269 9.3005
R12919 gnd.n5268 gnd.n1648 9.3005
R12920 gnd.n1616 gnd.n1615 9.3005
R12921 gnd.n5302 gnd.n5301 9.3005
R12922 gnd.n5303 gnd.n1613 9.3005
R12923 gnd.n5306 gnd.n5305 9.3005
R12924 gnd.n5304 gnd.n1614 9.3005
R12925 gnd.n1587 gnd.n1586 9.3005
R12926 gnd.n5338 gnd.n5337 9.3005
R12927 gnd.n5339 gnd.n1584 9.3005
R12928 gnd.n5342 gnd.n5341 9.3005
R12929 gnd.n5340 gnd.n1585 9.3005
R12930 gnd.n1556 gnd.n1555 9.3005
R12931 gnd.n5380 gnd.n5379 9.3005
R12932 gnd.n5381 gnd.n1553 9.3005
R12933 gnd.n5384 gnd.n5383 9.3005
R12934 gnd.n5382 gnd.n1554 9.3005
R12935 gnd.n1521 gnd.n1520 9.3005
R12936 gnd.n5423 gnd.n5422 9.3005
R12937 gnd.n5424 gnd.n1518 9.3005
R12938 gnd.n5430 gnd.n5429 9.3005
R12939 gnd.n5428 gnd.n1519 9.3005
R12940 gnd.n5427 gnd.n5426 9.3005
R12941 gnd.n1450 gnd.n1448 9.3005
R12942 gnd.n5852 gnd.n5851 9.3005
R12943 gnd.n5850 gnd.n1449 9.3005
R12944 gnd.n5849 gnd.n5848 9.3005
R12945 gnd.n5847 gnd.n1451 9.3005
R12946 gnd.n5846 gnd.n5845 9.3005
R12947 gnd.n5819 gnd.n5818 9.3005
R12948 gnd.n5703 gnd.n5702 9.3005
R12949 gnd.n5813 gnd.n5812 9.3005
R12950 gnd.n5811 gnd.n5810 9.3005
R12951 gnd.n5717 gnd.n5716 9.3005
R12952 gnd.n5805 gnd.n5804 9.3005
R12953 gnd.n5803 gnd.n5802 9.3005
R12954 gnd.n5729 gnd.n5728 9.3005
R12955 gnd.n5797 gnd.n5796 9.3005
R12956 gnd.n5795 gnd.n5794 9.3005
R12957 gnd.n5740 gnd.n5739 9.3005
R12958 gnd.n5789 gnd.n5788 9.3005
R12959 gnd.n5787 gnd.n5786 9.3005
R12960 gnd.n5752 gnd.n5751 9.3005
R12961 gnd.n5781 gnd.n5780 9.3005
R12962 gnd.n5779 gnd.n5778 9.3005
R12963 gnd.n5770 gnd.n5768 9.3005
R12964 gnd.n5767 gnd.n1456 9.3005
R12965 gnd.n5821 gnd.n5820 9.3005
R12966 gnd.n5843 gnd.n5842 9.3005
R12967 gnd.n5769 gnd.n1457 9.3005
R12968 gnd.n5777 gnd.n5776 9.3005
R12969 gnd.n5756 gnd.n5755 9.3005
R12970 gnd.n5783 gnd.n5782 9.3005
R12971 gnd.n5785 gnd.n5784 9.3005
R12972 gnd.n5746 gnd.n5745 9.3005
R12973 gnd.n5791 gnd.n5790 9.3005
R12974 gnd.n5793 gnd.n5792 9.3005
R12975 gnd.n5733 gnd.n5732 9.3005
R12976 gnd.n5799 gnd.n5798 9.3005
R12977 gnd.n5801 gnd.n5800 9.3005
R12978 gnd.n5723 gnd.n5722 9.3005
R12979 gnd.n5807 gnd.n5806 9.3005
R12980 gnd.n5809 gnd.n5808 9.3005
R12981 gnd.n5710 gnd.n5709 9.3005
R12982 gnd.n5815 gnd.n5814 9.3005
R12983 gnd.n5817 gnd.n5816 9.3005
R12984 gnd.n5706 gnd.n1487 9.3005
R12985 gnd.n5822 gnd.n1486 9.3005
R12986 gnd.n5824 gnd.n5823 9.3005
R12987 gnd.n5826 gnd.n5825 9.3005
R12988 gnd.n5828 gnd.n5827 9.3005
R12989 gnd.n5829 gnd.n1480 9.3005
R12990 gnd.n5831 gnd.n5830 9.3005
R12991 gnd.n5832 gnd.n1479 9.3005
R12992 gnd.n5834 gnd.n5833 9.3005
R12993 gnd.n5835 gnd.n1478 9.3005
R12994 gnd.n5680 gnd.n5679 9.3005
R12995 gnd.n5678 gnd.n5483 9.3005
R12996 gnd.n5677 gnd.n5676 9.3005
R12997 gnd.n5675 gnd.n5485 9.3005
R12998 gnd.n5674 gnd.n5673 9.3005
R12999 gnd.n5672 gnd.n5489 9.3005
R13000 gnd.n5671 gnd.n5670 9.3005
R13001 gnd.n5669 gnd.n5490 9.3005
R13002 gnd.n5668 gnd.n5667 9.3005
R13003 gnd.n5666 gnd.n5494 9.3005
R13004 gnd.n5665 gnd.n5664 9.3005
R13005 gnd.n5663 gnd.n5495 9.3005
R13006 gnd.n5662 gnd.n5661 9.3005
R13007 gnd.n5660 gnd.n5499 9.3005
R13008 gnd.n5659 gnd.n5658 9.3005
R13009 gnd.n5657 gnd.n5500 9.3005
R13010 gnd.n5656 gnd.n5655 9.3005
R13011 gnd.n1224 gnd.n1223 9.3005
R13012 gnd.n6103 gnd.n6102 9.3005
R13013 gnd.n6104 gnd.n1221 9.3005
R13014 gnd.n6107 gnd.n6106 9.3005
R13015 gnd.n6105 gnd.n1222 9.3005
R13016 gnd.n1182 gnd.n1181 9.3005
R13017 gnd.n6179 gnd.n6178 9.3005
R13018 gnd.n6180 gnd.n1179 9.3005
R13019 gnd.n6192 gnd.n6191 9.3005
R13020 gnd.n6190 gnd.n1180 9.3005
R13021 gnd.n6189 gnd.n6188 9.3005
R13022 gnd.n6187 gnd.n6181 9.3005
R13023 gnd.n6186 gnd.n6185 9.3005
R13024 gnd.n1133 gnd.n1132 9.3005
R13025 gnd.n6255 gnd.n6254 9.3005
R13026 gnd.n6256 gnd.n1131 9.3005
R13027 gnd.n6258 gnd.n6257 9.3005
R13028 gnd.n1105 gnd.n1104 9.3005
R13029 gnd.n6301 gnd.n6300 9.3005
R13030 gnd.n6302 gnd.n1103 9.3005
R13031 gnd.n6304 gnd.n6303 9.3005
R13032 gnd.n1074 gnd.n1073 9.3005
R13033 gnd.n6363 gnd.n6362 9.3005
R13034 gnd.n6364 gnd.n1072 9.3005
R13035 gnd.n6366 gnd.n6365 9.3005
R13036 gnd.n1047 gnd.n1046 9.3005
R13037 gnd.n6400 gnd.n6399 9.3005
R13038 gnd.n6401 gnd.n1045 9.3005
R13039 gnd.n6403 gnd.n6402 9.3005
R13040 gnd.n1018 gnd.n1017 9.3005
R13041 gnd.n6436 gnd.n6435 9.3005
R13042 gnd.n6437 gnd.n1016 9.3005
R13043 gnd.n6439 gnd.n6438 9.3005
R13044 gnd.n979 gnd.n978 9.3005
R13045 gnd.n6493 gnd.n6492 9.3005
R13046 gnd.n6494 gnd.n976 9.3005
R13047 gnd.n6497 gnd.n6496 9.3005
R13048 gnd.n6495 gnd.n977 9.3005
R13049 gnd.n958 gnd.n956 9.3005
R13050 gnd.n6529 gnd.n6528 9.3005
R13051 gnd.n6527 gnd.n957 9.3005
R13052 gnd.n6526 gnd.n6525 9.3005
R13053 gnd.n6524 gnd.n959 9.3005
R13054 gnd.n6523 gnd.n6522 9.3005
R13055 gnd.n881 gnd.n880 9.3005
R13056 gnd.n6729 gnd.n6728 9.3005
R13057 gnd.n6730 gnd.n878 9.3005
R13058 gnd.n6733 gnd.n6732 9.3005
R13059 gnd.n6731 gnd.n879 9.3005
R13060 gnd.n856 gnd.n855 9.3005
R13061 gnd.n6759 gnd.n6758 9.3005
R13062 gnd.n6760 gnd.n853 9.3005
R13063 gnd.n6763 gnd.n6762 9.3005
R13064 gnd.n6761 gnd.n854 9.3005
R13065 gnd.n831 gnd.n830 9.3005
R13066 gnd.n6789 gnd.n6788 9.3005
R13067 gnd.n6790 gnd.n828 9.3005
R13068 gnd.n6793 gnd.n6792 9.3005
R13069 gnd.n6791 gnd.n829 9.3005
R13070 gnd.n807 gnd.n806 9.3005
R13071 gnd.n6825 gnd.n6824 9.3005
R13072 gnd.n6826 gnd.n805 9.3005
R13073 gnd.n6828 gnd.n6827 9.3005
R13074 gnd.n768 gnd.n767 9.3005
R13075 gnd.n6859 gnd.n6858 9.3005
R13076 gnd.n5484 gnd.n5482 9.3005
R13077 gnd.n6855 gnd.n769 9.3005
R13078 gnd.n6854 gnd.n6853 9.3005
R13079 gnd.n6852 gnd.n772 9.3005
R13080 gnd.n6851 gnd.n6850 9.3005
R13081 gnd.n6849 gnd.n773 9.3005
R13082 gnd.n697 gnd.n695 9.3005
R13083 gnd.n6857 gnd.n6856 9.3005
R13084 gnd.n6879 gnd.n6878 9.3005
R13085 gnd.n744 gnd.n743 9.3005
R13086 gnd.n6885 gnd.n6884 9.3005
R13087 gnd.n6887 gnd.n6886 9.3005
R13088 gnd.n736 gnd.n735 9.3005
R13089 gnd.n6893 gnd.n6892 9.3005
R13090 gnd.n6895 gnd.n6894 9.3005
R13091 gnd.n726 gnd.n725 9.3005
R13092 gnd.n6901 gnd.n6900 9.3005
R13093 gnd.n6903 gnd.n6902 9.3005
R13094 gnd.n718 gnd.n717 9.3005
R13095 gnd.n6909 gnd.n6908 9.3005
R13096 gnd.n6911 gnd.n6910 9.3005
R13097 gnd.n708 gnd.n707 9.3005
R13098 gnd.n6917 gnd.n6916 9.3005
R13099 gnd.n6919 gnd.n6918 9.3005
R13100 gnd.n704 gnd.n702 9.3005
R13101 gnd.n6877 gnd.n6873 9.3005
R13102 gnd.n754 gnd.n753 9.3005
R13103 gnd.n6924 gnd.n6923 9.3005
R13104 gnd.n6922 gnd.n696 9.3005
R13105 gnd.n6921 gnd.n6920 9.3005
R13106 gnd.n703 gnd.n701 9.3005
R13107 gnd.n6915 gnd.n6914 9.3005
R13108 gnd.n6913 gnd.n6912 9.3005
R13109 gnd.n712 gnd.n711 9.3005
R13110 gnd.n6907 gnd.n6906 9.3005
R13111 gnd.n6905 gnd.n6904 9.3005
R13112 gnd.n722 gnd.n721 9.3005
R13113 gnd.n6899 gnd.n6898 9.3005
R13114 gnd.n6897 gnd.n6896 9.3005
R13115 gnd.n730 gnd.n729 9.3005
R13116 gnd.n6891 gnd.n6890 9.3005
R13117 gnd.n6889 gnd.n6888 9.3005
R13118 gnd.n740 gnd.n739 9.3005
R13119 gnd.n6883 gnd.n6882 9.3005
R13120 gnd.n6881 gnd.n6880 9.3005
R13121 gnd.n755 gnd.n750 9.3005
R13122 gnd.n6872 gnd.n6871 9.3005
R13123 gnd.n6870 gnd.n6869 9.3005
R13124 gnd.n559 gnd.n558 9.3005
R13125 gnd.n7081 gnd.n7080 9.3005
R13126 gnd.n7082 gnd.n556 9.3005
R13127 gnd.n7085 gnd.n7084 9.3005
R13128 gnd.n7083 gnd.n557 9.3005
R13129 gnd.n519 gnd.n518 9.3005
R13130 gnd.n7131 gnd.n7130 9.3005
R13131 gnd.n7132 gnd.n516 9.3005
R13132 gnd.n7134 gnd.n7133 9.3005
R13133 gnd.n7135 gnd.n515 9.3005
R13134 gnd.n7138 gnd.n7137 9.3005
R13135 gnd.n7139 gnd.n513 9.3005
R13136 gnd.n7142 gnd.n7141 9.3005
R13137 gnd.n7140 gnd.n514 9.3005
R13138 gnd.n454 gnd.n453 9.3005
R13139 gnd.n7201 gnd.n7200 9.3005
R13140 gnd.n7202 gnd.n451 9.3005
R13141 gnd.n7214 gnd.n7213 9.3005
R13142 gnd.n7212 gnd.n452 9.3005
R13143 gnd.n7211 gnd.n7210 9.3005
R13144 gnd.n7209 gnd.n7203 9.3005
R13145 gnd.n7208 gnd.n7207 9.3005
R13146 gnd.n7206 gnd.n7205 9.3005
R13147 gnd.n400 gnd.n399 9.3005
R13148 gnd.n7288 gnd.n7287 9.3005
R13149 gnd.n7289 gnd.n397 9.3005
R13150 gnd.n7297 gnd.n7296 9.3005
R13151 gnd.n7295 gnd.n398 9.3005
R13152 gnd.n7294 gnd.n7293 9.3005
R13153 gnd.n7292 gnd.n7290 9.3005
R13154 gnd.n7291 gnd.n95 9.3005
R13155 gnd.n6867 gnd.n6866 9.3005
R13156 gnd.n7759 gnd.n96 9.3005
R13157 gnd.t164 gnd.n3422 9.24152
R13158 gnd.n3324 gnd.t127 9.24152
R13159 gnd.n4625 gnd.t108 9.24152
R13160 gnd.n5132 gnd.t223 9.24152
R13161 gnd.n5377 gnd.t191 9.24152
R13162 gnd.n6715 gnd.t391 9.24152
R13163 gnd.n509 gnd.t240 9.24152
R13164 gnd.n7710 gnd.t185 9.24152
R13165 gnd.t133 gnd.t164 8.92286
R13166 gnd.n6109 gnd.n1200 8.92286
R13167 gnd.n6145 gnd.t71 8.92286
R13168 gnd.n6222 gnd.t0 8.92286
R13169 gnd.n6251 gnd.t143 8.92286
R13170 gnd.n6306 gnd.n1101 8.92286
R13171 gnd.n6397 gnd.n1049 8.92286
R13172 gnd.n6442 gnd.t7 8.92286
R13173 gnd.t130 gnd.n1006 8.92286
R13174 gnd.n995 gnd.n991 8.92286
R13175 gnd.n6643 gnd.n933 8.92286
R13176 gnd.n4594 gnd.n4569 8.92171
R13177 gnd.n4562 gnd.n4537 8.92171
R13178 gnd.n4530 gnd.n4505 8.92171
R13179 gnd.n4499 gnd.n4474 8.92171
R13180 gnd.n4467 gnd.n4442 8.92171
R13181 gnd.n4435 gnd.n4410 8.92171
R13182 gnd.n4403 gnd.n4378 8.92171
R13183 gnd.n4372 gnd.n4347 8.92171
R13184 gnd.n6570 gnd.n6552 8.72777
R13185 gnd.n4098 gnd.t180 8.60421
R13186 gnd.t204 gnd.n1783 8.60421
R13187 gnd.n5444 gnd.t215 8.60421
R13188 gnd.n6350 gnd.t4 8.60421
R13189 gnd.n6387 gnd.t395 8.60421
R13190 gnd.n7128 gnd.t231 8.60421
R13191 gnd.n7686 gnd.t225 8.60421
R13192 gnd.n3502 gnd.n3482 8.43656
R13193 gnd.n54 gnd.n34 8.43656
R13194 gnd.n6215 gnd.n1156 8.28555
R13195 gnd.n6297 gnd.n1109 8.28555
R13196 gnd.n6380 gnd.n1042 8.28555
R13197 gnd.n6457 gnd.n6456 8.28555
R13198 gnd.n4595 gnd.n4567 8.14595
R13199 gnd.n4563 gnd.n4535 8.14595
R13200 gnd.n4531 gnd.n4503 8.14595
R13201 gnd.n4500 gnd.n4472 8.14595
R13202 gnd.n4468 gnd.n4440 8.14595
R13203 gnd.n4436 gnd.n4408 8.14595
R13204 gnd.n4404 gnd.n4376 8.14595
R13205 gnd.n4373 gnd.n4345 8.14595
R13206 gnd.n5234 gnd.n0 8.10675
R13207 gnd.n7760 gnd.n7759 8.10675
R13208 gnd.n4600 gnd.n4599 7.97301
R13209 gnd.t184 gnd.n3613 7.9669
R13210 gnd.n7760 gnd.n94 7.95236
R13211 gnd.n6877 gnd.n753 7.75808
R13212 gnd.n5768 gnd.n5767 7.75808
R13213 gnd.n7447 gnd.n7394 7.75808
R13214 gnd.n4784 gnd.n4758 7.75808
R13215 gnd.n6215 gnd.n1157 7.64824
R13216 gnd.n6298 gnd.t136 7.64824
R13217 gnd.n6298 gnd.n6297 7.64824
R13218 gnd.n6405 gnd.n1042 7.64824
R13219 gnd.t172 gnd.n6405 7.64824
R13220 gnd.n6457 gnd.n1000 7.64824
R13221 gnd.n3543 gnd.n3542 7.53171
R13222 gnd.n4007 gnd.t9 7.32958
R13223 gnd.n1284 gnd.n1283 7.30353
R13224 gnd.n6569 gnd.n6568 7.30353
R13225 gnd.n3967 gnd.n3686 7.01093
R13226 gnd.n3689 gnd.n3687 7.01093
R13227 gnd.n3977 gnd.n3976 7.01093
R13228 gnd.n3988 gnd.n3670 7.01093
R13229 gnd.n3987 gnd.n3673 7.01093
R13230 gnd.n3998 gnd.n3661 7.01093
R13231 gnd.n3664 gnd.n3662 7.01093
R13232 gnd.n4008 gnd.n4007 7.01093
R13233 gnd.n4018 gnd.n3642 7.01093
R13234 gnd.n4017 gnd.n3645 7.01093
R13235 gnd.n4026 gnd.n3636 7.01093
R13236 gnd.n4038 gnd.n3626 7.01093
R13237 gnd.n4048 gnd.n3611 7.01093
R13238 gnd.n4064 gnd.n4063 7.01093
R13239 gnd.n3613 gnd.n3550 7.01093
R13240 gnd.n4118 gnd.n3551 7.01093
R13241 gnd.n4112 gnd.n4111 7.01093
R13242 gnd.n3600 gnd.n3562 7.01093
R13243 gnd.n4104 gnd.n3573 7.01093
R13244 gnd.n3591 gnd.n3586 7.01093
R13245 gnd.n4098 gnd.n4097 7.01093
R13246 gnd.n4144 gnd.n3457 7.01093
R13247 gnd.n4143 gnd.n4142 7.01093
R13248 gnd.n4155 gnd.n4154 7.01093
R13249 gnd.n3450 gnd.n3442 7.01093
R13250 gnd.n4184 gnd.n3430 7.01093
R13251 gnd.n4183 gnd.n3433 7.01093
R13252 gnd.n4194 gnd.n3422 7.01093
R13253 gnd.n3423 gnd.n3411 7.01093
R13254 gnd.n4205 gnd.n3412 7.01093
R13255 gnd.n4229 gnd.n3403 7.01093
R13256 gnd.n4228 gnd.n3394 7.01093
R13257 gnd.n4251 gnd.n4250 7.01093
R13258 gnd.n4269 gnd.n3375 7.01093
R13259 gnd.n4268 gnd.n3378 7.01093
R13260 gnd.n4279 gnd.n3367 7.01093
R13261 gnd.n3368 gnd.n3355 7.01093
R13262 gnd.n4290 gnd.n3356 7.01093
R13263 gnd.n4317 gnd.n3340 7.01093
R13264 gnd.n4329 gnd.n4328 7.01093
R13265 gnd.n4311 gnd.n3333 7.01093
R13266 gnd.n4340 gnd.n4339 7.01093
R13267 gnd.n4613 gnd.n1908 7.01093
R13268 gnd.n4613 gnd.n4612 7.01093
R13269 gnd.n4611 gnd.n3324 7.01093
R13270 gnd.n4625 gnd.n1900 7.01093
R13271 gnd.n1901 gnd.n1893 7.01093
R13272 gnd.n4635 gnd.n1819 7.01093
R13273 gnd.n6154 gnd.n1200 7.01093
R13274 gnd.n1206 gnd.n1205 7.01093
R13275 gnd.n1206 gnd.t115 7.01093
R13276 gnd.n1101 gnd.n1100 7.01093
R13277 gnd.n6386 gnd.n1049 7.01093
R13278 gnd.n6482 gnd.n991 7.01093
R13279 gnd.n6643 gnd.n932 7.01093
R13280 gnd.t102 gnd.n891 7.01093
R13281 gnd.n3645 gnd.t176 6.69227
R13282 gnd.n3433 gnd.t133 6.69227
R13283 gnd.n4318 gnd.t177 6.69227
R13284 gnd.n1261 gnd.t141 6.69227
R13285 gnd.t391 gnd.n6714 6.69227
R13286 gnd.n6705 gnd.n6704 6.5566
R13287 gnd.n1356 gnd.n1355 6.5566
R13288 gnd.n6040 gnd.n1292 6.5566
R13289 gnd.n6580 gnd.n6579 6.5566
R13290 gnd.t105 gnd.n1260 6.37362
R13291 gnd.n6242 gnd.n6241 6.37362
R13292 gnd.n1117 gnd.t136 6.37362
R13293 gnd.n6407 gnd.t172 6.37362
R13294 gnd.n6449 gnd.n1005 6.37362
R13295 gnd.n6480 gnd.t62 6.37362
R13296 gnd.n5776 gnd.n5773 6.20656
R13297 gnd.n755 gnd.n749 6.20656
R13298 gnd.t166 gnd.n4074 6.05496
R13299 gnd.n4075 gnd.t165 6.05496
R13300 gnd.t157 gnd.n3457 6.05496
R13301 gnd.t182 gnd.n4239 6.05496
R13302 gnd.n6099 gnd.n1262 6.05496
R13303 gnd.n1100 gnd.t4 6.05496
R13304 gnd.t395 gnd.n6386 6.05496
R13305 gnd.n6713 gnd.n6712 6.05496
R13306 gnd.n4597 gnd.n4567 5.81868
R13307 gnd.n4565 gnd.n4535 5.81868
R13308 gnd.n4533 gnd.n4503 5.81868
R13309 gnd.n4502 gnd.n4472 5.81868
R13310 gnd.n4470 gnd.n4440 5.81868
R13311 gnd.n4438 gnd.n4408 5.81868
R13312 gnd.n4406 gnd.n4376 5.81868
R13313 gnd.n4375 gnd.n4345 5.81868
R13314 gnd.n6163 gnd.n6162 5.73631
R13315 gnd.n6146 gnd.n1186 5.73631
R13316 gnd.n6359 gnd.n1079 5.73631
R13317 gnd.n6342 gnd.n1069 5.73631
R13318 gnd.n6539 gnd.n945 5.73631
R13319 gnd.n6471 gnd.n6470 5.73631
R13320 gnd.n933 gnd.t102 5.73631
R13321 gnd.n6709 gnd.n657 5.62001
R13322 gnd.n6035 gnd.n1360 5.62001
R13323 gnd.n6036 gnd.n6035 5.62001
R13324 gnd.n6575 gnd.n657 5.62001
R13325 gnd.n3826 gnd.n3821 5.4308
R13326 gnd.n4643 gnd.n1886 5.4308
R13327 gnd.n4142 gnd.t183 5.41765
R13328 gnd.t163 gnd.n4165 5.41765
R13329 gnd.t151 gnd.n3387 5.41765
R13330 gnd.t137 gnd.n6145 5.41765
R13331 gnd.n6531 gnd.t387 5.41765
R13332 gnd.n6252 gnd.n6251 5.09899
R13333 gnd.n6234 gnd.n6233 5.09899
R13334 gnd.n6418 gnd.n1039 5.09899
R13335 gnd.n6442 gnd.n6441 5.09899
R13336 gnd.n6726 gnd.t56 5.09899
R13337 gnd.n4595 gnd.n4594 5.04292
R13338 gnd.n4563 gnd.n4562 5.04292
R13339 gnd.n4531 gnd.n4530 5.04292
R13340 gnd.n4500 gnd.n4499 5.04292
R13341 gnd.n4468 gnd.n4467 5.04292
R13342 gnd.n4436 gnd.n4435 5.04292
R13343 gnd.n4404 gnd.n4403 5.04292
R13344 gnd.n4373 gnd.n4372 5.04292
R13345 gnd.n4105 gnd.t162 4.78034
R13346 gnd.n3412 gnd.t179 4.78034
R13347 gnd.t389 gnd.n5577 4.78034
R13348 gnd.n6146 gnd.t137 4.78034
R13349 gnd.t387 gnd.n945 4.78034
R13350 gnd.n6712 gnd.t56 4.78034
R13351 gnd.n825 gnd.t155 4.78034
R13352 gnd.n3547 gnd.n3544 4.74817
R13353 gnd.n3597 gnd.n3463 4.74817
R13354 gnd.n3584 gnd.n3462 4.74817
R13355 gnd.n3461 gnd.n3460 4.74817
R13356 gnd.n3593 gnd.n3544 4.74817
R13357 gnd.n3594 gnd.n3463 4.74817
R13358 gnd.n3596 gnd.n3462 4.74817
R13359 gnd.n3583 gnd.n3461 4.74817
R13360 gnd.n7309 gnd.n113 4.74817
R13361 gnd.n370 gnd.n112 4.74817
R13362 gnd.n7333 gnd.n111 4.74817
R13363 gnd.n7752 gnd.n106 4.74817
R13364 gnd.n7750 gnd.n107 4.74817
R13365 gnd.n7281 gnd.n113 4.74817
R13366 gnd.n7310 gnd.n112 4.74817
R13367 gnd.n371 gnd.n111 4.74817
R13368 gnd.n7332 gnd.n106 4.74817
R13369 gnd.n7751 gnd.n7750 4.74817
R13370 gnd.n1972 gnd.n1971 4.74817
R13371 gnd.n1966 gnd.n1915 4.74817
R13372 gnd.n1964 gnd.n1963 4.74817
R13373 gnd.n1959 gnd.n1918 4.74817
R13374 gnd.n7315 gnd.n382 4.74817
R13375 gnd.n7320 gnd.n7317 4.74817
R13376 gnd.n7318 gnd.n358 4.74817
R13377 gnd.n7348 gnd.n7347 4.74817
R13378 gnd.n7248 gnd.n382 4.74817
R13379 gnd.n7317 gnd.n7316 4.74817
R13380 gnd.n7319 gnd.n7318 4.74817
R13381 gnd.n7347 gnd.n7346 4.74817
R13382 gnd.n7350 gnd.n7349 4.74817
R13383 gnd.n5219 gnd.n1631 4.74817
R13384 gnd.n5239 gnd.n1630 4.74817
R13385 gnd.n1674 gnd.n1629 4.74817
R13386 gnd.n5261 gnd.n1628 4.74817
R13387 gnd.n1632 gnd.n1627 4.74817
R13388 gnd.n5200 gnd.n1631 4.74817
R13389 gnd.n5220 gnd.n1630 4.74817
R13390 gnd.n5240 gnd.n1629 4.74817
R13391 gnd.n1673 gnd.n1628 4.74817
R13392 gnd.n5260 gnd.n1627 4.74817
R13393 gnd.n1915 gnd.n1913 4.74817
R13394 gnd.n1965 gnd.n1964 4.74817
R13395 gnd.n1918 gnd.n1916 4.74817
R13396 gnd.n3542 gnd.n3541 4.74296
R13397 gnd.n94 gnd.n93 4.74296
R13398 gnd.n3502 gnd.n3501 4.7074
R13399 gnd.n3522 gnd.n3521 4.7074
R13400 gnd.n54 gnd.n53 4.7074
R13401 gnd.n74 gnd.n73 4.7074
R13402 gnd.n3542 gnd.n3522 4.65959
R13403 gnd.n94 gnd.n74 4.65959
R13404 gnd.n6989 gnd.n659 4.6132
R13405 gnd.n6031 gnd.n6030 4.6132
R13406 gnd.n6165 gnd.n1191 4.46168
R13407 gnd.n6195 gnd.n1174 4.46168
R13408 gnd.n6348 gnd.n1076 4.46168
R13409 gnd.n6370 gnd.n6369 4.46168
R13410 gnd.n6532 gnd.n952 4.46168
R13411 gnd.t12 gnd.n6538 4.46168
R13412 gnd.n6548 gnd.n6547 4.46168
R13413 gnd.n2602 gnd.n222 4.46168
R13414 gnd.n6565 gnd.n6552 4.46111
R13415 gnd.n4580 gnd.n4576 4.38594
R13416 gnd.n4548 gnd.n4544 4.38594
R13417 gnd.n4516 gnd.n4512 4.38594
R13418 gnd.n4485 gnd.n4481 4.38594
R13419 gnd.n4453 gnd.n4449 4.38594
R13420 gnd.n4421 gnd.n4417 4.38594
R13421 gnd.n4389 gnd.n4385 4.38594
R13422 gnd.n4358 gnd.n4354 4.38594
R13423 gnd.n4591 gnd.n4569 4.26717
R13424 gnd.n4559 gnd.n4537 4.26717
R13425 gnd.n4527 gnd.n4505 4.26717
R13426 gnd.n4496 gnd.n4474 4.26717
R13427 gnd.n4464 gnd.n4442 4.26717
R13428 gnd.n4432 gnd.n4410 4.26717
R13429 gnd.n4400 gnd.n4378 4.26717
R13430 gnd.n4369 gnd.n4347 4.26717
R13431 gnd.n4049 gnd.t178 4.14303
R13432 gnd.n4279 gnd.t175 4.14303
R13433 gnd.n4599 gnd.n4598 4.08274
R13434 gnd.n6704 gnd.n6703 4.05904
R13435 gnd.n1355 gnd.n1354 4.05904
R13436 gnd.n6043 gnd.n1292 4.05904
R13437 gnd.n6581 gnd.n6580 4.05904
R13438 gnd.n15 gnd.n7 3.99943
R13439 gnd.n6162 gnd.t23 3.82437
R13440 gnd.t174 gnd.n1157 3.82437
R13441 gnd.n6221 gnd.n1152 3.82437
R13442 gnd.n6288 gnd.n6287 3.82437
R13443 gnd.n6426 gnd.n1026 3.82437
R13444 gnd.n6490 gnd.n981 3.82437
R13445 gnd.t6 gnd.n1000 3.82437
R13446 gnd.n6470 gnd.t26 3.82437
R13447 gnd.n4122 gnd.n3543 3.81325
R13448 gnd.n3522 gnd.n3502 3.72967
R13449 gnd.n74 gnd.n54 3.72967
R13450 gnd.n4599 gnd.n4471 3.70378
R13451 gnd.n15 gnd.n14 3.60163
R13452 gnd.n5051 gnd.t37 3.50571
R13453 gnd.n1452 gnd.t45 3.50571
R13454 gnd.n7078 gnd.t33 3.50571
R13455 gnd.t41 gnd.n235 3.50571
R13456 gnd.n4590 gnd.n4571 3.49141
R13457 gnd.n4558 gnd.n4539 3.49141
R13458 gnd.n4526 gnd.n4507 3.49141
R13459 gnd.n4495 gnd.n4476 3.49141
R13460 gnd.n4463 gnd.n4444 3.49141
R13461 gnd.n4431 gnd.n4412 3.49141
R13462 gnd.n4399 gnd.n4380 3.49141
R13463 gnd.n4368 gnd.n4349 3.49141
R13464 gnd.n7007 gnd.n7006 3.29747
R13465 gnd.n7006 gnd.n7005 3.29747
R13466 gnd.n7627 gnd.n7624 3.29747
R13467 gnd.n7628 gnd.n7627 3.29747
R13468 gnd.n4927 gnd.n4869 3.29747
R13469 gnd.n4869 gnd.n4864 3.29747
R13470 gnd.n5902 gnd.n5897 3.29747
R13471 gnd.n5927 gnd.n5902 3.29747
R13472 gnd.n1260 gnd.n1218 3.18706
R13473 gnd.n6261 gnd.t10 3.18706
R13474 gnd.n6280 gnd.n1099 3.18706
R13475 gnd.n6396 gnd.n1052 3.18706
R13476 gnd.n1028 gnd.t2 3.18706
R13477 gnd.n6715 gnd.n891 3.18706
R13478 gnd.n3628 gnd.t178 2.8684
R13479 gnd.n5639 gnd.t131 2.8684
R13480 gnd.t141 gnd.t105 2.8684
R13481 gnd.n6745 gnd.t145 2.8684
R13482 gnd.n3523 gnd.t255 2.82907
R13483 gnd.n3523 gnd.t362 2.82907
R13484 gnd.n3525 gnd.t230 2.82907
R13485 gnd.n3525 gnd.t276 2.82907
R13486 gnd.n3527 gnd.t304 2.82907
R13487 gnd.n3527 gnd.t283 2.82907
R13488 gnd.n3529 gnd.t281 2.82907
R13489 gnd.n3529 gnd.t268 2.82907
R13490 gnd.n3531 gnd.t290 2.82907
R13491 gnd.n3531 gnd.t343 2.82907
R13492 gnd.n3533 gnd.t207 2.82907
R13493 gnd.n3533 gnd.t326 2.82907
R13494 gnd.n3535 gnd.t372 2.82907
R13495 gnd.n3535 gnd.t288 2.82907
R13496 gnd.n3537 gnd.t328 2.82907
R13497 gnd.n3537 gnd.t263 2.82907
R13498 gnd.n3539 gnd.t218 2.82907
R13499 gnd.n3539 gnd.t214 2.82907
R13500 gnd.n3464 gnd.t295 2.82907
R13501 gnd.n3464 gnd.t324 2.82907
R13502 gnd.n3466 gnd.t339 2.82907
R13503 gnd.n3466 gnd.t257 2.82907
R13504 gnd.n3468 gnd.t319 2.82907
R13505 gnd.n3468 gnd.t312 2.82907
R13506 gnd.n3470 gnd.t378 2.82907
R13507 gnd.n3470 gnd.t364 2.82907
R13508 gnd.n3472 gnd.t265 2.82907
R13509 gnd.n3472 gnd.t332 2.82907
R13510 gnd.n3474 gnd.t353 2.82907
R13511 gnd.n3474 gnd.t203 2.82907
R13512 gnd.n3476 gnd.t235 2.82907
R13513 gnd.n3476 gnd.t322 2.82907
R13514 gnd.n3478 gnd.t333 2.82907
R13515 gnd.n3478 gnd.t375 2.82907
R13516 gnd.n3480 gnd.t289 2.82907
R13517 gnd.n3480 gnd.t308 2.82907
R13518 gnd.n3483 gnd.t382 2.82907
R13519 gnd.n3483 gnd.t227 2.82907
R13520 gnd.n3485 gnd.t229 2.82907
R13521 gnd.n3485 gnd.t192 2.82907
R13522 gnd.n3487 gnd.t340 2.82907
R13523 gnd.n3487 gnd.t383 2.82907
R13524 gnd.n3489 gnd.t377 2.82907
R13525 gnd.n3489 gnd.t237 2.82907
R13526 gnd.n3491 gnd.t366 2.82907
R13527 gnd.n3491 gnd.t299 2.82907
R13528 gnd.n3493 gnd.t341 2.82907
R13529 gnd.n3493 gnd.t379 2.82907
R13530 gnd.n3495 gnd.t380 2.82907
R13531 gnd.n3495 gnd.t357 2.82907
R13532 gnd.n3497 gnd.t359 2.82907
R13533 gnd.n3497 gnd.t342 2.82907
R13534 gnd.n3499 gnd.t338 2.82907
R13535 gnd.n3499 gnd.t321 2.82907
R13536 gnd.n3503 gnd.t314 2.82907
R13537 gnd.n3503 gnd.t188 2.82907
R13538 gnd.n3505 gnd.t294 2.82907
R13539 gnd.n3505 gnd.t346 2.82907
R13540 gnd.n3507 gnd.t376 2.82907
R13541 gnd.n3507 gnd.t356 2.82907
R13542 gnd.n3509 gnd.t354 2.82907
R13543 gnd.n3509 gnd.t331 2.82907
R13544 gnd.n3511 gnd.t361 2.82907
R13545 gnd.n3511 gnd.t248 2.82907
R13546 gnd.n3513 gnd.t275 2.82907
R13547 gnd.n3513 gnd.t208 2.82907
R13548 gnd.n3515 gnd.t266 2.82907
R13549 gnd.n3515 gnd.t360 2.82907
R13550 gnd.n3517 gnd.t224 2.82907
R13551 gnd.n3517 gnd.t323 2.82907
R13552 gnd.n3519 gnd.t284 2.82907
R13553 gnd.n3519 gnd.t279 2.82907
R13554 gnd.n91 gnd.t293 2.82907
R13555 gnd.n91 gnd.t311 2.82907
R13556 gnd.n89 gnd.t196 2.82907
R13557 gnd.n89 gnd.t278 2.82907
R13558 gnd.n87 gnd.t252 2.82907
R13559 gnd.n87 gnd.t320 2.82907
R13560 gnd.n85 gnd.t274 2.82907
R13561 gnd.n85 gnd.t336 2.82907
R13562 gnd.n83 gnd.t297 2.82907
R13563 gnd.n83 gnd.t267 2.82907
R13564 gnd.n81 gnd.t219 2.82907
R13565 gnd.n81 gnd.t246 2.82907
R13566 gnd.n79 gnd.t250 2.82907
R13567 gnd.n79 gnd.t272 2.82907
R13568 gnd.n77 gnd.t241 2.82907
R13569 gnd.n77 gnd.t355 2.82907
R13570 gnd.n75 gnd.t313 2.82907
R13571 gnd.n75 gnd.t212 2.82907
R13572 gnd.n32 gnd.t292 2.82907
R13573 gnd.n32 gnd.t302 2.82907
R13574 gnd.n30 gnd.t242 2.82907
R13575 gnd.n30 gnd.t186 2.82907
R13576 gnd.n28 gnd.t367 2.82907
R13577 gnd.n28 gnd.t269 2.82907
R13578 gnd.n26 gnd.t261 2.82907
R13579 gnd.n26 gnd.t221 2.82907
R13580 gnd.n24 gnd.t384 2.82907
R13581 gnd.n24 gnd.t253 2.82907
R13582 gnd.n22 gnd.t233 2.82907
R13583 gnd.n22 gnd.t244 2.82907
R13584 gnd.n20 gnd.t352 2.82907
R13585 gnd.n20 gnd.t305 2.82907
R13586 gnd.n18 gnd.t286 2.82907
R13587 gnd.n18 gnd.t201 2.82907
R13588 gnd.n16 gnd.t371 2.82907
R13589 gnd.n16 gnd.t273 2.82907
R13590 gnd.n51 gnd.t334 2.82907
R13591 gnd.n51 gnd.t307 2.82907
R13592 gnd.n49 gnd.t317 2.82907
R13593 gnd.n49 gnd.t330 2.82907
R13594 gnd.n47 gnd.t329 2.82907
R13595 gnd.n47 gnd.t348 2.82907
R13596 gnd.n45 gnd.t349 2.82907
R13597 gnd.n45 gnd.t318 2.82907
R13598 gnd.n43 gnd.t315 2.82907
R13599 gnd.n43 gnd.t200 2.82907
R13600 gnd.n41 gnd.t198 2.82907
R13601 gnd.n41 gnd.t347 2.82907
R13602 gnd.n39 gnd.t358 2.82907
R13603 gnd.n39 gnd.t369 2.82907
R13604 gnd.n37 gnd.t368 2.82907
R13605 gnd.n37 gnd.t190 2.82907
R13606 gnd.n35 gnd.t194 2.82907
R13607 gnd.n35 gnd.t222 2.82907
R13608 gnd.n71 gnd.t344 2.82907
R13609 gnd.n71 gnd.t373 2.82907
R13610 gnd.n69 gnd.t270 2.82907
R13611 gnd.n69 gnd.t351 2.82907
R13612 gnd.n67 gnd.t310 2.82907
R13613 gnd.n67 gnd.t210 2.82907
R13614 gnd.n65 gnd.t345 2.82907
R13615 gnd.n65 gnd.t239 2.82907
R13616 gnd.n63 gnd.t370 2.82907
R13617 gnd.n63 gnd.t327 2.82907
R13618 gnd.n61 gnd.t285 2.82907
R13619 gnd.n61 gnd.t306 2.82907
R13620 gnd.n59 gnd.t309 2.82907
R13621 gnd.n59 gnd.t337 2.82907
R13622 gnd.n57 gnd.t298 2.82907
R13623 gnd.n57 gnd.t256 2.82907
R13624 gnd.n55 gnd.t381 2.82907
R13625 gnd.n55 gnd.t259 2.82907
R13626 gnd.n4587 gnd.n4586 2.71565
R13627 gnd.n4555 gnd.n4554 2.71565
R13628 gnd.n4523 gnd.n4522 2.71565
R13629 gnd.n4492 gnd.n4491 2.71565
R13630 gnd.n4460 gnd.n4459 2.71565
R13631 gnd.n4428 gnd.n4427 2.71565
R13632 gnd.n4396 gnd.n4395 2.71565
R13633 gnd.n4365 gnd.n4364 2.71565
R13634 gnd.t71 gnd.n1174 2.54975
R13635 gnd.n1167 gnd.n1166 2.54975
R13636 gnd.n6279 gnd.n6278 2.54975
R13637 gnd.n6280 gnd.t1 2.54975
R13638 gnd.n6349 gnd.t173 2.54975
R13639 gnd.t159 gnd.n1057 2.54975
R13640 gnd.t135 gnd.n1052 2.54975
R13641 gnd.n6379 gnd.n1066 2.54975
R13642 gnd.n6499 gnd.n972 2.54975
R13643 gnd.n4122 gnd.n3544 2.27742
R13644 gnd.n4122 gnd.n3463 2.27742
R13645 gnd.n4122 gnd.n3462 2.27742
R13646 gnd.n4122 gnd.n3461 2.27742
R13647 gnd.n7749 gnd.n113 2.27742
R13648 gnd.n7749 gnd.n112 2.27742
R13649 gnd.n7749 gnd.n111 2.27742
R13650 gnd.n7749 gnd.n106 2.27742
R13651 gnd.n7750 gnd.n7749 2.27742
R13652 gnd.n382 gnd.n110 2.27742
R13653 gnd.n7317 gnd.n110 2.27742
R13654 gnd.n7318 gnd.n110 2.27742
R13655 gnd.n7347 gnd.n110 2.27742
R13656 gnd.n7349 gnd.n110 2.27742
R13657 gnd.n5292 gnd.n1631 2.27742
R13658 gnd.n5292 gnd.n1630 2.27742
R13659 gnd.n5292 gnd.n1629 2.27742
R13660 gnd.n5292 gnd.n1628 2.27742
R13661 gnd.n5292 gnd.n1627 2.27742
R13662 gnd.n1972 gnd.n1626 2.27742
R13663 gnd.n1915 gnd.n1626 2.27742
R13664 gnd.n1964 gnd.n1626 2.27742
R13665 gnd.n1918 gnd.n1626 2.27742
R13666 gnd.n3976 gnd.t83 2.23109
R13667 gnd.n3599 gnd.t162 2.23109
R13668 gnd.t149 gnd.n6260 2.23109
R13669 gnd.n6433 gnd.t170 2.23109
R13670 gnd.n4583 gnd.n4573 1.93989
R13671 gnd.n4551 gnd.n4541 1.93989
R13672 gnd.n4519 gnd.n4509 1.93989
R13673 gnd.n4488 gnd.n4478 1.93989
R13674 gnd.n4456 gnd.n4446 1.93989
R13675 gnd.n4424 gnd.n4414 1.93989
R13676 gnd.n4392 gnd.n4382 1.93989
R13677 gnd.n4361 gnd.n4351 1.93989
R13678 gnd.t115 gnd.n1164 1.91244
R13679 gnd.n6208 gnd.t144 1.91244
R13680 gnd.n1145 gnd.t143 1.91244
R13681 gnd.n6286 gnd.n1117 1.91244
R13682 gnd.n6407 gnd.n6406 1.91244
R13683 gnd.n6419 gnd.t7 1.91244
R13684 gnd.n6464 gnd.t3 1.91244
R13685 gnd.t160 gnd.n3987 1.59378
R13686 gnd.n4166 gnd.t163 1.59378
R13687 gnd.n3396 gnd.t151 1.59378
R13688 gnd.n5107 gnd.t213 1.59378
R13689 gnd.t139 gnd.n1159 1.59378
R13690 gnd.n6489 gnd.t147 1.59378
R13691 gnd.n194 gnd.t291 1.59378
R13692 gnd.t87 gnd.n1201 1.27512
R13693 gnd.n6194 gnd.n1176 1.27512
R13694 gnd.t144 gnd.n6207 1.27512
R13695 gnd.n6350 gnd.n6349 1.27512
R13696 gnd.n6387 gnd.n1057 1.27512
R13697 gnd.t3 gnd.n973 1.27512
R13698 gnd.n6481 gnd.n6480 1.27512
R13699 gnd.n6519 gnd.n6518 1.27512
R13700 gnd.n3829 gnd.n3821 1.16414
R13701 gnd.n4646 gnd.n1886 1.16414
R13702 gnd.n4582 gnd.n4575 1.16414
R13703 gnd.n4550 gnd.n4543 1.16414
R13704 gnd.n4518 gnd.n4511 1.16414
R13705 gnd.n4487 gnd.n4480 1.16414
R13706 gnd.n4455 gnd.n4448 1.16414
R13707 gnd.n4423 gnd.n4416 1.16414
R13708 gnd.n4391 gnd.n4384 1.16414
R13709 gnd.n4360 gnd.n4353 1.16414
R13710 gnd.n6989 gnd.n6988 0.970197
R13711 gnd.n6031 gnd.n1361 0.970197
R13712 gnd.n4566 gnd.n4534 0.962709
R13713 gnd.n4598 gnd.n4566 0.962709
R13714 gnd.n4439 gnd.n4407 0.962709
R13715 gnd.n4471 gnd.n4439 0.962709
R13716 gnd.n4075 gnd.t166 0.956468
R13717 gnd.n4240 gnd.t182 0.956468
R13718 gnd.n5167 gnd.t234 0.956468
R13719 gnd.n5185 gnd.n1691 0.956468
R13720 gnd.t254 gnd.n1532 0.956468
R13721 gnd.t168 gnd.n5525 0.956468
R13722 gnd.t10 gnd.t149 0.956468
R13723 gnd.t2 gnd.t170 0.956468
R13724 gnd.n851 gnd.t397 0.956468
R13725 gnd.t211 gnd.n490 0.956468
R13726 gnd.n7490 gnd.n120 0.956468
R13727 gnd.n156 gnd.t209 0.956468
R13728 gnd.n2 gnd.n1 0.672012
R13729 gnd.n3 gnd.n2 0.672012
R13730 gnd.n4 gnd.n3 0.672012
R13731 gnd.n5 gnd.n4 0.672012
R13732 gnd.n6 gnd.n5 0.672012
R13733 gnd.n7 gnd.n6 0.672012
R13734 gnd.n9 gnd.n8 0.672012
R13735 gnd.n10 gnd.n9 0.672012
R13736 gnd.n11 gnd.n10 0.672012
R13737 gnd.n12 gnd.n11 0.672012
R13738 gnd.n13 gnd.n12 0.672012
R13739 gnd.n14 gnd.n13 0.672012
R13740 gnd.n5217 gnd.n1687 0.637812
R13741 gnd.n5222 gnd.n1685 0.637812
R13742 gnd.n5229 gnd.n1679 0.637812
R13743 gnd.n5242 gnd.n1668 0.637812
R13744 gnd.n5237 gnd.n1670 0.637812
R13745 gnd.n5250 gnd.n1662 0.637812
R13746 gnd.n5263 gnd.n1652 0.637812
R13747 gnd.n5258 gnd.n1654 0.637812
R13748 gnd.n5289 gnd.n1634 0.637812
R13749 gnd.n5276 gnd.n1637 0.637812
R13750 gnd.n5299 gnd.n1618 0.637812
R13751 gnd.n5282 gnd.n1620 0.637812
R13752 gnd.n5308 gnd.n1611 0.637812
R13753 gnd.n5325 gnd.n1599 0.637812
R13754 gnd.n5312 gnd.n1602 0.637812
R13755 gnd.n5335 gnd.n1589 0.637812
R13756 gnd.n5318 gnd.n1591 0.637812
R13757 gnd.n5344 gnd.n1582 0.637812
R13758 gnd.n5367 gnd.n1568 0.637812
R13759 gnd.n5348 gnd.n1571 0.637812
R13760 gnd.n5377 gnd.n1558 0.637812
R13761 gnd.n1560 gnd.n1550 0.637812
R13762 gnd.n5387 gnd.n5386 0.637812
R13763 gnd.n5410 gnd.n1532 0.637812
R13764 gnd.n5353 gnd.n1535 0.637812
R13765 gnd.n5420 gnd.n1523 0.637812
R13766 gnd.n5403 gnd.n5402 0.637812
R13767 gnd.n5432 gnd.n1516 0.637812
R13768 gnd.n5444 gnd.n1505 0.637812
R13769 gnd.n1508 gnd.n1498 0.637812
R13770 gnd.n5453 gnd.n5452 0.637812
R13771 gnd.n5854 gnd.n1446 0.637812
R13772 gnd.n5864 gnd.n1436 0.637812
R13773 gnd.n1452 gnd.n1439 0.637812
R13774 gnd.n5966 gnd.n1426 0.637812
R13775 gnd.n5698 gnd.n1428 0.637812
R13776 gnd.n6242 gnd.t0 0.637812
R13777 gnd.n6240 gnd.n1135 0.637812
R13778 gnd.n6232 gnd.n1128 0.637812
R13779 gnd.n6432 gnd.n1022 0.637812
R13780 gnd.n1014 gnd.n1013 0.637812
R13781 gnd.n6449 gnd.t130 0.637812
R13782 gnd.n6547 gnd.t80 0.637812
R13783 gnd.n7068 gnd.n572 0.637812
R13784 gnd.n7060 gnd.n7059 0.637812
R13785 gnd.n7078 gnd.n562 0.637812
R13786 gnd.n577 gnd.n554 0.637812
R13787 gnd.n7087 gnd.n531 0.637812
R13788 gnd.n7118 gnd.n534 0.637812
R13789 gnd.n7100 gnd.n7099 0.637812
R13790 gnd.n7128 gnd.n523 0.637812
R13791 gnd.n7111 gnd.n7110 0.637812
R13792 gnd.n545 gnd.n543 0.637812
R13793 gnd.n7153 gnd.n499 0.637812
R13794 gnd.n7162 gnd.n487 0.637812
R13795 gnd.n7161 gnd.n490 0.637812
R13796 gnd.n7144 gnd.n466 0.637812
R13797 gnd.n7188 gnd.n469 0.637812
R13798 gnd.n509 gnd.n456 0.637812
R13799 gnd.n7198 gnd.n458 0.637812
R13800 gnd.n7181 gnd.n7180 0.637812
R13801 gnd.n7216 gnd.n439 0.637812
R13802 gnd.n7228 gnd.n442 0.637812
R13803 gnd.n7237 gnd.n431 0.637812
R13804 gnd.n7236 gnd.n423 0.637812
R13805 gnd.n7258 gnd.n7257 0.637812
R13806 gnd.n7275 gnd.n414 0.637812
R13807 gnd.n7262 gnd.n402 0.637812
R13808 gnd.n7285 gnd.n404 0.637812
R13809 gnd.n7268 gnd.n395 0.637812
R13810 gnd.n7299 gnd.n387 0.637812
R13811 gnd.n7312 gnd.n378 0.637812
R13812 gnd.n7323 gnd.n7322 0.637812
R13813 gnd.n7330 gnd.n367 0.637812
R13814 gnd.n7335 gnd.n360 0.637812
R13815 gnd.n7344 gnd.n7343 0.637812
R13816 gnd.n7754 gnd.n102 0.637812
R13817 gnd.n7353 gnd.n7352 0.637812
R13818 gnd.n7360 gnd.n117 0.637812
R13819 gnd.n7761 gnd.n7760 0.63688
R13820 gnd gnd.n0 0.634843
R13821 gnd.n3541 gnd.n3540 0.573776
R13822 gnd.n3540 gnd.n3538 0.573776
R13823 gnd.n3538 gnd.n3536 0.573776
R13824 gnd.n3536 gnd.n3534 0.573776
R13825 gnd.n3534 gnd.n3532 0.573776
R13826 gnd.n3532 gnd.n3530 0.573776
R13827 gnd.n3530 gnd.n3528 0.573776
R13828 gnd.n3528 gnd.n3526 0.573776
R13829 gnd.n3526 gnd.n3524 0.573776
R13830 gnd.n3482 gnd.n3481 0.573776
R13831 gnd.n3481 gnd.n3479 0.573776
R13832 gnd.n3479 gnd.n3477 0.573776
R13833 gnd.n3477 gnd.n3475 0.573776
R13834 gnd.n3475 gnd.n3473 0.573776
R13835 gnd.n3473 gnd.n3471 0.573776
R13836 gnd.n3471 gnd.n3469 0.573776
R13837 gnd.n3469 gnd.n3467 0.573776
R13838 gnd.n3467 gnd.n3465 0.573776
R13839 gnd.n3501 gnd.n3500 0.573776
R13840 gnd.n3500 gnd.n3498 0.573776
R13841 gnd.n3498 gnd.n3496 0.573776
R13842 gnd.n3496 gnd.n3494 0.573776
R13843 gnd.n3494 gnd.n3492 0.573776
R13844 gnd.n3492 gnd.n3490 0.573776
R13845 gnd.n3490 gnd.n3488 0.573776
R13846 gnd.n3488 gnd.n3486 0.573776
R13847 gnd.n3486 gnd.n3484 0.573776
R13848 gnd.n3521 gnd.n3520 0.573776
R13849 gnd.n3520 gnd.n3518 0.573776
R13850 gnd.n3518 gnd.n3516 0.573776
R13851 gnd.n3516 gnd.n3514 0.573776
R13852 gnd.n3514 gnd.n3512 0.573776
R13853 gnd.n3512 gnd.n3510 0.573776
R13854 gnd.n3510 gnd.n3508 0.573776
R13855 gnd.n3508 gnd.n3506 0.573776
R13856 gnd.n3506 gnd.n3504 0.573776
R13857 gnd.n78 gnd.n76 0.573776
R13858 gnd.n80 gnd.n78 0.573776
R13859 gnd.n82 gnd.n80 0.573776
R13860 gnd.n84 gnd.n82 0.573776
R13861 gnd.n86 gnd.n84 0.573776
R13862 gnd.n88 gnd.n86 0.573776
R13863 gnd.n90 gnd.n88 0.573776
R13864 gnd.n92 gnd.n90 0.573776
R13865 gnd.n93 gnd.n92 0.573776
R13866 gnd.n19 gnd.n17 0.573776
R13867 gnd.n21 gnd.n19 0.573776
R13868 gnd.n23 gnd.n21 0.573776
R13869 gnd.n25 gnd.n23 0.573776
R13870 gnd.n27 gnd.n25 0.573776
R13871 gnd.n29 gnd.n27 0.573776
R13872 gnd.n31 gnd.n29 0.573776
R13873 gnd.n33 gnd.n31 0.573776
R13874 gnd.n34 gnd.n33 0.573776
R13875 gnd.n38 gnd.n36 0.573776
R13876 gnd.n40 gnd.n38 0.573776
R13877 gnd.n42 gnd.n40 0.573776
R13878 gnd.n44 gnd.n42 0.573776
R13879 gnd.n46 gnd.n44 0.573776
R13880 gnd.n48 gnd.n46 0.573776
R13881 gnd.n50 gnd.n48 0.573776
R13882 gnd.n52 gnd.n50 0.573776
R13883 gnd.n53 gnd.n52 0.573776
R13884 gnd.n58 gnd.n56 0.573776
R13885 gnd.n60 gnd.n58 0.573776
R13886 gnd.n62 gnd.n60 0.573776
R13887 gnd.n64 gnd.n62 0.573776
R13888 gnd.n66 gnd.n64 0.573776
R13889 gnd.n68 gnd.n66 0.573776
R13890 gnd.n70 gnd.n68 0.573776
R13891 gnd.n72 gnd.n70 0.573776
R13892 gnd.n73 gnd.n72 0.573776
R13893 gnd.n6865 gnd.n6864 0.489829
R13894 gnd.n5554 gnd.n1455 0.489829
R13895 gnd.n5484 gnd.n1478 0.489829
R13896 gnd.n6858 gnd.n6857 0.489829
R13897 gnd.n4302 gnd.n1890 0.486781
R13898 gnd.n3878 gnd.n3877 0.48678
R13899 gnd.n4620 gnd.n1844 0.480683
R13900 gnd.n3962 gnd.n3961 0.480683
R13901 gnd.n3107 gnd.n2096 0.480683
R13902 gnd.n2435 gnd.n2434 0.480683
R13903 gnd.n7446 gnd.n7391 0.477634
R13904 gnd.n4785 gnd.n4780 0.477634
R13905 gnd.n7664 gnd.n7663 0.442573
R13906 gnd.n7071 gnd.n567 0.442573
R13907 gnd.n5962 gnd.n5961 0.442573
R13908 gnd.n5046 gnd.n1817 0.442573
R13909 gnd.n7749 gnd.n110 0.4255
R13910 gnd.n5292 gnd.n1626 0.4255
R13911 gnd.n5773 gnd.n5755 0.388379
R13912 gnd.n4579 gnd.n4578 0.388379
R13913 gnd.n4547 gnd.n4546 0.388379
R13914 gnd.n4515 gnd.n4514 0.388379
R13915 gnd.n4484 gnd.n4483 0.388379
R13916 gnd.n4452 gnd.n4451 0.388379
R13917 gnd.n4420 gnd.n4419 0.388379
R13918 gnd.n4388 gnd.n4387 0.388379
R13919 gnd.n4357 gnd.n4356 0.388379
R13920 gnd.n6881 gnd.n749 0.388379
R13921 gnd.n7761 gnd.n15 0.374463
R13922 gnd.n2599 gnd.n110 0.331293
R13923 gnd.n3318 gnd.n1626 0.331293
R13924 gnd.n3358 gnd.t177 0.319156
R13925 gnd.n5217 gnd.t202 0.319156
R13926 gnd.n1657 gnd.t280 0.319156
R13927 gnd.n5272 gnd.t280 0.319156
R13928 gnd.t282 gnd.n1589 0.319156
R13929 gnd.t19 gnd.n5480 0.319156
R13930 gnd.n1160 gnd.t139 0.319156
R13931 gnd.n1001 gnd.t147 0.319156
R13932 gnd.n6832 gnd.t52 0.319156
R13933 gnd.n7237 gnd.t249 0.319156
R13934 gnd.n7307 gnd.t243 0.319156
R13935 gnd.n7313 gnd.t243 0.319156
R13936 gnd.n7360 gnd.t260 0.319156
R13937 gnd.n3796 gnd.n3774 0.311721
R13938 gnd gnd.n7761 0.295112
R13939 gnd.n7540 gnd.n348 0.293183
R13940 gnd.n5033 gnd.n4821 0.293183
R13941 gnd.n4691 gnd.n4690 0.268793
R13942 gnd.n7541 gnd.n7540 0.258122
R13943 gnd.n6927 gnd.n6926 0.258122
R13944 gnd.n5972 gnd.n5971 0.258122
R13945 gnd.n5033 gnd.n5032 0.258122
R13946 gnd.n5845 gnd.n5844 0.247451
R13947 gnd.n6868 gnd.n6867 0.247451
R13948 gnd.n4690 gnd.n4689 0.241354
R13949 gnd.n659 gnd.n656 0.229039
R13950 gnd.n660 gnd.n659 0.229039
R13951 gnd.n6030 gnd.n1364 0.229039
R13952 gnd.n6030 gnd.n6029 0.229039
R13953 gnd.n3543 gnd.n0 0.210825
R13954 gnd.n3950 gnd.n3749 0.206293
R13955 gnd.n4596 gnd.n4568 0.155672
R13956 gnd.n4589 gnd.n4568 0.155672
R13957 gnd.n4589 gnd.n4588 0.155672
R13958 gnd.n4588 gnd.n4572 0.155672
R13959 gnd.n4581 gnd.n4572 0.155672
R13960 gnd.n4581 gnd.n4580 0.155672
R13961 gnd.n4564 gnd.n4536 0.155672
R13962 gnd.n4557 gnd.n4536 0.155672
R13963 gnd.n4557 gnd.n4556 0.155672
R13964 gnd.n4556 gnd.n4540 0.155672
R13965 gnd.n4549 gnd.n4540 0.155672
R13966 gnd.n4549 gnd.n4548 0.155672
R13967 gnd.n4532 gnd.n4504 0.155672
R13968 gnd.n4525 gnd.n4504 0.155672
R13969 gnd.n4525 gnd.n4524 0.155672
R13970 gnd.n4524 gnd.n4508 0.155672
R13971 gnd.n4517 gnd.n4508 0.155672
R13972 gnd.n4517 gnd.n4516 0.155672
R13973 gnd.n4501 gnd.n4473 0.155672
R13974 gnd.n4494 gnd.n4473 0.155672
R13975 gnd.n4494 gnd.n4493 0.155672
R13976 gnd.n4493 gnd.n4477 0.155672
R13977 gnd.n4486 gnd.n4477 0.155672
R13978 gnd.n4486 gnd.n4485 0.155672
R13979 gnd.n4469 gnd.n4441 0.155672
R13980 gnd.n4462 gnd.n4441 0.155672
R13981 gnd.n4462 gnd.n4461 0.155672
R13982 gnd.n4461 gnd.n4445 0.155672
R13983 gnd.n4454 gnd.n4445 0.155672
R13984 gnd.n4454 gnd.n4453 0.155672
R13985 gnd.n4437 gnd.n4409 0.155672
R13986 gnd.n4430 gnd.n4409 0.155672
R13987 gnd.n4430 gnd.n4429 0.155672
R13988 gnd.n4429 gnd.n4413 0.155672
R13989 gnd.n4422 gnd.n4413 0.155672
R13990 gnd.n4422 gnd.n4421 0.155672
R13991 gnd.n4405 gnd.n4377 0.155672
R13992 gnd.n4398 gnd.n4377 0.155672
R13993 gnd.n4398 gnd.n4397 0.155672
R13994 gnd.n4397 gnd.n4381 0.155672
R13995 gnd.n4390 gnd.n4381 0.155672
R13996 gnd.n4390 gnd.n4389 0.155672
R13997 gnd.n4374 gnd.n4346 0.155672
R13998 gnd.n4367 gnd.n4346 0.155672
R13999 gnd.n4367 gnd.n4366 0.155672
R14000 gnd.n4366 gnd.n4350 0.155672
R14001 gnd.n4359 gnd.n4350 0.155672
R14002 gnd.n4359 gnd.n4358 0.155672
R14003 gnd.n4722 gnd.n1844 0.152939
R14004 gnd.n4722 gnd.n4721 0.152939
R14005 gnd.n4721 gnd.n4720 0.152939
R14006 gnd.n4720 gnd.n1846 0.152939
R14007 gnd.n1847 gnd.n1846 0.152939
R14008 gnd.n1848 gnd.n1847 0.152939
R14009 gnd.n1849 gnd.n1848 0.152939
R14010 gnd.n1850 gnd.n1849 0.152939
R14011 gnd.n1851 gnd.n1850 0.152939
R14012 gnd.n1852 gnd.n1851 0.152939
R14013 gnd.n1853 gnd.n1852 0.152939
R14014 gnd.n1854 gnd.n1853 0.152939
R14015 gnd.n1855 gnd.n1854 0.152939
R14016 gnd.n1856 gnd.n1855 0.152939
R14017 gnd.n4692 gnd.n1856 0.152939
R14018 gnd.n4692 gnd.n4691 0.152939
R14019 gnd.n3963 gnd.n3962 0.152939
R14020 gnd.n3963 gnd.n3667 0.152939
R14021 gnd.n3991 gnd.n3667 0.152939
R14022 gnd.n3992 gnd.n3991 0.152939
R14023 gnd.n3993 gnd.n3992 0.152939
R14024 gnd.n3994 gnd.n3993 0.152939
R14025 gnd.n3994 gnd.n3639 0.152939
R14026 gnd.n4021 gnd.n3639 0.152939
R14027 gnd.n4022 gnd.n4021 0.152939
R14028 gnd.n4023 gnd.n4022 0.152939
R14029 gnd.n4023 gnd.n3617 0.152939
R14030 gnd.n4052 gnd.n3617 0.152939
R14031 gnd.n4053 gnd.n4052 0.152939
R14032 gnd.n4054 gnd.n4053 0.152939
R14033 gnd.n4055 gnd.n4054 0.152939
R14034 gnd.n4057 gnd.n4055 0.152939
R14035 gnd.n4057 gnd.n4056 0.152939
R14036 gnd.n4056 gnd.n3566 0.152939
R14037 gnd.n3567 gnd.n3566 0.152939
R14038 gnd.n3568 gnd.n3567 0.152939
R14039 gnd.n3587 gnd.n3568 0.152939
R14040 gnd.n3588 gnd.n3587 0.152939
R14041 gnd.n3588 gnd.n3454 0.152939
R14042 gnd.n4147 gnd.n3454 0.152939
R14043 gnd.n4148 gnd.n4147 0.152939
R14044 gnd.n4149 gnd.n4148 0.152939
R14045 gnd.n4150 gnd.n4149 0.152939
R14046 gnd.n4150 gnd.n3427 0.152939
R14047 gnd.n4187 gnd.n3427 0.152939
R14048 gnd.n4188 gnd.n4187 0.152939
R14049 gnd.n4189 gnd.n4188 0.152939
R14050 gnd.n4190 gnd.n4189 0.152939
R14051 gnd.n4190 gnd.n3400 0.152939
R14052 gnd.n4232 gnd.n3400 0.152939
R14053 gnd.n4233 gnd.n4232 0.152939
R14054 gnd.n4234 gnd.n4233 0.152939
R14055 gnd.n4235 gnd.n4234 0.152939
R14056 gnd.n4235 gnd.n3372 0.152939
R14057 gnd.n4272 gnd.n3372 0.152939
R14058 gnd.n4273 gnd.n4272 0.152939
R14059 gnd.n4274 gnd.n4273 0.152939
R14060 gnd.n4275 gnd.n4274 0.152939
R14061 gnd.n4275 gnd.n3345 0.152939
R14062 gnd.n4321 gnd.n3345 0.152939
R14063 gnd.n4322 gnd.n4321 0.152939
R14064 gnd.n4323 gnd.n4322 0.152939
R14065 gnd.n4324 gnd.n4323 0.152939
R14066 gnd.n4324 gnd.n1905 0.152939
R14067 gnd.n4616 gnd.n1905 0.152939
R14068 gnd.n4617 gnd.n4616 0.152939
R14069 gnd.n4618 gnd.n4617 0.152939
R14070 gnd.n4619 gnd.n4618 0.152939
R14071 gnd.n4620 gnd.n4619 0.152939
R14072 gnd.n3961 gnd.n3691 0.152939
R14073 gnd.n3712 gnd.n3691 0.152939
R14074 gnd.n3713 gnd.n3712 0.152939
R14075 gnd.n3719 gnd.n3713 0.152939
R14076 gnd.n3720 gnd.n3719 0.152939
R14077 gnd.n3721 gnd.n3720 0.152939
R14078 gnd.n3721 gnd.n3710 0.152939
R14079 gnd.n3729 gnd.n3710 0.152939
R14080 gnd.n3730 gnd.n3729 0.152939
R14081 gnd.n3731 gnd.n3730 0.152939
R14082 gnd.n3731 gnd.n3708 0.152939
R14083 gnd.n3739 gnd.n3708 0.152939
R14084 gnd.n3740 gnd.n3739 0.152939
R14085 gnd.n3741 gnd.n3740 0.152939
R14086 gnd.n3741 gnd.n3706 0.152939
R14087 gnd.n3749 gnd.n3706 0.152939
R14088 gnd.n4689 gnd.n1861 0.152939
R14089 gnd.n1863 gnd.n1861 0.152939
R14090 gnd.n1864 gnd.n1863 0.152939
R14091 gnd.n1865 gnd.n1864 0.152939
R14092 gnd.n1866 gnd.n1865 0.152939
R14093 gnd.n1867 gnd.n1866 0.152939
R14094 gnd.n1868 gnd.n1867 0.152939
R14095 gnd.n1869 gnd.n1868 0.152939
R14096 gnd.n1870 gnd.n1869 0.152939
R14097 gnd.n1871 gnd.n1870 0.152939
R14098 gnd.n1872 gnd.n1871 0.152939
R14099 gnd.n1873 gnd.n1872 0.152939
R14100 gnd.n1874 gnd.n1873 0.152939
R14101 gnd.n1875 gnd.n1874 0.152939
R14102 gnd.n1876 gnd.n1875 0.152939
R14103 gnd.n1877 gnd.n1876 0.152939
R14104 gnd.n1878 gnd.n1877 0.152939
R14105 gnd.n1879 gnd.n1878 0.152939
R14106 gnd.n1880 gnd.n1879 0.152939
R14107 gnd.n1881 gnd.n1880 0.152939
R14108 gnd.n1882 gnd.n1881 0.152939
R14109 gnd.n1883 gnd.n1882 0.152939
R14110 gnd.n1887 gnd.n1883 0.152939
R14111 gnd.n1888 gnd.n1887 0.152939
R14112 gnd.n1889 gnd.n1888 0.152939
R14113 gnd.n1890 gnd.n1889 0.152939
R14114 gnd.n4124 gnd.n4123 0.152939
R14115 gnd.n4125 gnd.n4124 0.152939
R14116 gnd.n4126 gnd.n4125 0.152939
R14117 gnd.n4127 gnd.n4126 0.152939
R14118 gnd.n4128 gnd.n4127 0.152939
R14119 gnd.n4129 gnd.n4128 0.152939
R14120 gnd.n4129 gnd.n3408 0.152939
R14121 gnd.n4208 gnd.n3408 0.152939
R14122 gnd.n4209 gnd.n4208 0.152939
R14123 gnd.n4210 gnd.n4209 0.152939
R14124 gnd.n4211 gnd.n4210 0.152939
R14125 gnd.n4212 gnd.n4211 0.152939
R14126 gnd.n4213 gnd.n4212 0.152939
R14127 gnd.n4214 gnd.n4213 0.152939
R14128 gnd.n4215 gnd.n4214 0.152939
R14129 gnd.n4216 gnd.n4215 0.152939
R14130 gnd.n4216 gnd.n3352 0.152939
R14131 gnd.n4293 gnd.n3352 0.152939
R14132 gnd.n4294 gnd.n4293 0.152939
R14133 gnd.n4295 gnd.n4294 0.152939
R14134 gnd.n4296 gnd.n4295 0.152939
R14135 gnd.n4297 gnd.n4296 0.152939
R14136 gnd.n4298 gnd.n4297 0.152939
R14137 gnd.n4299 gnd.n4298 0.152939
R14138 gnd.n4300 gnd.n4299 0.152939
R14139 gnd.n4301 gnd.n4300 0.152939
R14140 gnd.n4303 gnd.n4301 0.152939
R14141 gnd.n4303 gnd.n4302 0.152939
R14142 gnd.n3879 gnd.n3878 0.152939
R14143 gnd.n3879 gnd.n3769 0.152939
R14144 gnd.n3894 gnd.n3769 0.152939
R14145 gnd.n3895 gnd.n3894 0.152939
R14146 gnd.n3896 gnd.n3895 0.152939
R14147 gnd.n3896 gnd.n3757 0.152939
R14148 gnd.n3910 gnd.n3757 0.152939
R14149 gnd.n3911 gnd.n3910 0.152939
R14150 gnd.n3912 gnd.n3911 0.152939
R14151 gnd.n3913 gnd.n3912 0.152939
R14152 gnd.n3914 gnd.n3913 0.152939
R14153 gnd.n3915 gnd.n3914 0.152939
R14154 gnd.n3916 gnd.n3915 0.152939
R14155 gnd.n3917 gnd.n3916 0.152939
R14156 gnd.n3918 gnd.n3917 0.152939
R14157 gnd.n3919 gnd.n3918 0.152939
R14158 gnd.n3920 gnd.n3919 0.152939
R14159 gnd.n3921 gnd.n3920 0.152939
R14160 gnd.n3922 gnd.n3921 0.152939
R14161 gnd.n3923 gnd.n3922 0.152939
R14162 gnd.n3924 gnd.n3923 0.152939
R14163 gnd.n3924 gnd.n3623 0.152939
R14164 gnd.n4041 gnd.n3623 0.152939
R14165 gnd.n4042 gnd.n4041 0.152939
R14166 gnd.n4043 gnd.n4042 0.152939
R14167 gnd.n4044 gnd.n4043 0.152939
R14168 gnd.n4044 gnd.n3545 0.152939
R14169 gnd.n4121 gnd.n3545 0.152939
R14170 gnd.n3797 gnd.n3796 0.152939
R14171 gnd.n3798 gnd.n3797 0.152939
R14172 gnd.n3799 gnd.n3798 0.152939
R14173 gnd.n3800 gnd.n3799 0.152939
R14174 gnd.n3801 gnd.n3800 0.152939
R14175 gnd.n3802 gnd.n3801 0.152939
R14176 gnd.n3803 gnd.n3802 0.152939
R14177 gnd.n3804 gnd.n3803 0.152939
R14178 gnd.n3805 gnd.n3804 0.152939
R14179 gnd.n3806 gnd.n3805 0.152939
R14180 gnd.n3807 gnd.n3806 0.152939
R14181 gnd.n3808 gnd.n3807 0.152939
R14182 gnd.n3809 gnd.n3808 0.152939
R14183 gnd.n3810 gnd.n3809 0.152939
R14184 gnd.n3811 gnd.n3810 0.152939
R14185 gnd.n3812 gnd.n3811 0.152939
R14186 gnd.n3813 gnd.n3812 0.152939
R14187 gnd.n3814 gnd.n3813 0.152939
R14188 gnd.n3815 gnd.n3814 0.152939
R14189 gnd.n3816 gnd.n3815 0.152939
R14190 gnd.n3817 gnd.n3816 0.152939
R14191 gnd.n3818 gnd.n3817 0.152939
R14192 gnd.n3822 gnd.n3818 0.152939
R14193 gnd.n3823 gnd.n3822 0.152939
R14194 gnd.n3823 gnd.n3780 0.152939
R14195 gnd.n3877 gnd.n3780 0.152939
R14196 gnd.n3107 gnd.n3106 0.152939
R14197 gnd.n3106 gnd.n3105 0.152939
R14198 gnd.n3105 gnd.n2102 0.152939
R14199 gnd.n2107 gnd.n2102 0.152939
R14200 gnd.n2108 gnd.n2107 0.152939
R14201 gnd.n2109 gnd.n2108 0.152939
R14202 gnd.n2114 gnd.n2109 0.152939
R14203 gnd.n2115 gnd.n2114 0.152939
R14204 gnd.n2116 gnd.n2115 0.152939
R14205 gnd.n2117 gnd.n2116 0.152939
R14206 gnd.n2122 gnd.n2117 0.152939
R14207 gnd.n2123 gnd.n2122 0.152939
R14208 gnd.n2124 gnd.n2123 0.152939
R14209 gnd.n2125 gnd.n2124 0.152939
R14210 gnd.n2130 gnd.n2125 0.152939
R14211 gnd.n2131 gnd.n2130 0.152939
R14212 gnd.n2132 gnd.n2131 0.152939
R14213 gnd.n2133 gnd.n2132 0.152939
R14214 gnd.n2138 gnd.n2133 0.152939
R14215 gnd.n2139 gnd.n2138 0.152939
R14216 gnd.n2140 gnd.n2139 0.152939
R14217 gnd.n2141 gnd.n2140 0.152939
R14218 gnd.n2146 gnd.n2141 0.152939
R14219 gnd.n2147 gnd.n2146 0.152939
R14220 gnd.n2148 gnd.n2147 0.152939
R14221 gnd.n2149 gnd.n2148 0.152939
R14222 gnd.n2154 gnd.n2149 0.152939
R14223 gnd.n2155 gnd.n2154 0.152939
R14224 gnd.n2156 gnd.n2155 0.152939
R14225 gnd.n2157 gnd.n2156 0.152939
R14226 gnd.n2162 gnd.n2157 0.152939
R14227 gnd.n2163 gnd.n2162 0.152939
R14228 gnd.n2164 gnd.n2163 0.152939
R14229 gnd.n2165 gnd.n2164 0.152939
R14230 gnd.n2170 gnd.n2165 0.152939
R14231 gnd.n2171 gnd.n2170 0.152939
R14232 gnd.n2172 gnd.n2171 0.152939
R14233 gnd.n2173 gnd.n2172 0.152939
R14234 gnd.n2178 gnd.n2173 0.152939
R14235 gnd.n2179 gnd.n2178 0.152939
R14236 gnd.n2180 gnd.n2179 0.152939
R14237 gnd.n2181 gnd.n2180 0.152939
R14238 gnd.n2186 gnd.n2181 0.152939
R14239 gnd.n2187 gnd.n2186 0.152939
R14240 gnd.n2188 gnd.n2187 0.152939
R14241 gnd.n2189 gnd.n2188 0.152939
R14242 gnd.n2194 gnd.n2189 0.152939
R14243 gnd.n2195 gnd.n2194 0.152939
R14244 gnd.n2196 gnd.n2195 0.152939
R14245 gnd.n2197 gnd.n2196 0.152939
R14246 gnd.n2202 gnd.n2197 0.152939
R14247 gnd.n2203 gnd.n2202 0.152939
R14248 gnd.n2204 gnd.n2203 0.152939
R14249 gnd.n2205 gnd.n2204 0.152939
R14250 gnd.n2210 gnd.n2205 0.152939
R14251 gnd.n2211 gnd.n2210 0.152939
R14252 gnd.n2212 gnd.n2211 0.152939
R14253 gnd.n2213 gnd.n2212 0.152939
R14254 gnd.n2218 gnd.n2213 0.152939
R14255 gnd.n2219 gnd.n2218 0.152939
R14256 gnd.n2220 gnd.n2219 0.152939
R14257 gnd.n2221 gnd.n2220 0.152939
R14258 gnd.n2226 gnd.n2221 0.152939
R14259 gnd.n2227 gnd.n2226 0.152939
R14260 gnd.n2228 gnd.n2227 0.152939
R14261 gnd.n2229 gnd.n2228 0.152939
R14262 gnd.n2234 gnd.n2229 0.152939
R14263 gnd.n2235 gnd.n2234 0.152939
R14264 gnd.n2236 gnd.n2235 0.152939
R14265 gnd.n2237 gnd.n2236 0.152939
R14266 gnd.n2242 gnd.n2237 0.152939
R14267 gnd.n2243 gnd.n2242 0.152939
R14268 gnd.n2244 gnd.n2243 0.152939
R14269 gnd.n2245 gnd.n2244 0.152939
R14270 gnd.n2250 gnd.n2245 0.152939
R14271 gnd.n2251 gnd.n2250 0.152939
R14272 gnd.n2252 gnd.n2251 0.152939
R14273 gnd.n2253 gnd.n2252 0.152939
R14274 gnd.n2258 gnd.n2253 0.152939
R14275 gnd.n2259 gnd.n2258 0.152939
R14276 gnd.n2260 gnd.n2259 0.152939
R14277 gnd.n2261 gnd.n2260 0.152939
R14278 gnd.n2266 gnd.n2261 0.152939
R14279 gnd.n2267 gnd.n2266 0.152939
R14280 gnd.n2268 gnd.n2267 0.152939
R14281 gnd.n2269 gnd.n2268 0.152939
R14282 gnd.n2274 gnd.n2269 0.152939
R14283 gnd.n2275 gnd.n2274 0.152939
R14284 gnd.n2276 gnd.n2275 0.152939
R14285 gnd.n2277 gnd.n2276 0.152939
R14286 gnd.n2282 gnd.n2277 0.152939
R14287 gnd.n2283 gnd.n2282 0.152939
R14288 gnd.n2284 gnd.n2283 0.152939
R14289 gnd.n2285 gnd.n2284 0.152939
R14290 gnd.n2290 gnd.n2285 0.152939
R14291 gnd.n2291 gnd.n2290 0.152939
R14292 gnd.n2292 gnd.n2291 0.152939
R14293 gnd.n2293 gnd.n2292 0.152939
R14294 gnd.n2298 gnd.n2293 0.152939
R14295 gnd.n2299 gnd.n2298 0.152939
R14296 gnd.n2300 gnd.n2299 0.152939
R14297 gnd.n2301 gnd.n2300 0.152939
R14298 gnd.n2306 gnd.n2301 0.152939
R14299 gnd.n2307 gnd.n2306 0.152939
R14300 gnd.n2308 gnd.n2307 0.152939
R14301 gnd.n2309 gnd.n2308 0.152939
R14302 gnd.n2314 gnd.n2309 0.152939
R14303 gnd.n2315 gnd.n2314 0.152939
R14304 gnd.n2316 gnd.n2315 0.152939
R14305 gnd.n2317 gnd.n2316 0.152939
R14306 gnd.n2322 gnd.n2317 0.152939
R14307 gnd.n2323 gnd.n2322 0.152939
R14308 gnd.n2324 gnd.n2323 0.152939
R14309 gnd.n2325 gnd.n2324 0.152939
R14310 gnd.n2330 gnd.n2325 0.152939
R14311 gnd.n2331 gnd.n2330 0.152939
R14312 gnd.n2332 gnd.n2331 0.152939
R14313 gnd.n2333 gnd.n2332 0.152939
R14314 gnd.n2338 gnd.n2333 0.152939
R14315 gnd.n2339 gnd.n2338 0.152939
R14316 gnd.n2340 gnd.n2339 0.152939
R14317 gnd.n2341 gnd.n2340 0.152939
R14318 gnd.n2346 gnd.n2341 0.152939
R14319 gnd.n2347 gnd.n2346 0.152939
R14320 gnd.n2348 gnd.n2347 0.152939
R14321 gnd.n2349 gnd.n2348 0.152939
R14322 gnd.n2354 gnd.n2349 0.152939
R14323 gnd.n2355 gnd.n2354 0.152939
R14324 gnd.n2356 gnd.n2355 0.152939
R14325 gnd.n2357 gnd.n2356 0.152939
R14326 gnd.n2362 gnd.n2357 0.152939
R14327 gnd.n2363 gnd.n2362 0.152939
R14328 gnd.n2364 gnd.n2363 0.152939
R14329 gnd.n2365 gnd.n2364 0.152939
R14330 gnd.n2370 gnd.n2365 0.152939
R14331 gnd.n2371 gnd.n2370 0.152939
R14332 gnd.n2372 gnd.n2371 0.152939
R14333 gnd.n2373 gnd.n2372 0.152939
R14334 gnd.n2378 gnd.n2373 0.152939
R14335 gnd.n2379 gnd.n2378 0.152939
R14336 gnd.n2380 gnd.n2379 0.152939
R14337 gnd.n2381 gnd.n2380 0.152939
R14338 gnd.n2386 gnd.n2381 0.152939
R14339 gnd.n2387 gnd.n2386 0.152939
R14340 gnd.n2388 gnd.n2387 0.152939
R14341 gnd.n2389 gnd.n2388 0.152939
R14342 gnd.n2394 gnd.n2389 0.152939
R14343 gnd.n2395 gnd.n2394 0.152939
R14344 gnd.n2396 gnd.n2395 0.152939
R14345 gnd.n2397 gnd.n2396 0.152939
R14346 gnd.n2402 gnd.n2397 0.152939
R14347 gnd.n2403 gnd.n2402 0.152939
R14348 gnd.n2404 gnd.n2403 0.152939
R14349 gnd.n2405 gnd.n2404 0.152939
R14350 gnd.n2410 gnd.n2405 0.152939
R14351 gnd.n2411 gnd.n2410 0.152939
R14352 gnd.n2412 gnd.n2411 0.152939
R14353 gnd.n2413 gnd.n2412 0.152939
R14354 gnd.n2418 gnd.n2413 0.152939
R14355 gnd.n2419 gnd.n2418 0.152939
R14356 gnd.n2420 gnd.n2419 0.152939
R14357 gnd.n2421 gnd.n2420 0.152939
R14358 gnd.n2426 gnd.n2421 0.152939
R14359 gnd.n2427 gnd.n2426 0.152939
R14360 gnd.n2428 gnd.n2427 0.152939
R14361 gnd.n2429 gnd.n2428 0.152939
R14362 gnd.n2434 gnd.n2429 0.152939
R14363 gnd.n2768 gnd.n2435 0.152939
R14364 gnd.n2768 gnd.n2767 0.152939
R14365 gnd.n2767 gnd.n2766 0.152939
R14366 gnd.n2766 gnd.n2437 0.152939
R14367 gnd.n2444 gnd.n2437 0.152939
R14368 gnd.n2445 gnd.n2444 0.152939
R14369 gnd.n2446 gnd.n2445 0.152939
R14370 gnd.n2451 gnd.n2446 0.152939
R14371 gnd.n2452 gnd.n2451 0.152939
R14372 gnd.n2453 gnd.n2452 0.152939
R14373 gnd.n2454 gnd.n2453 0.152939
R14374 gnd.n2459 gnd.n2454 0.152939
R14375 gnd.n2460 gnd.n2459 0.152939
R14376 gnd.n2461 gnd.n2460 0.152939
R14377 gnd.n2462 gnd.n2461 0.152939
R14378 gnd.n2467 gnd.n2462 0.152939
R14379 gnd.n2468 gnd.n2467 0.152939
R14380 gnd.n2469 gnd.n2468 0.152939
R14381 gnd.n2470 gnd.n2469 0.152939
R14382 gnd.n2475 gnd.n2470 0.152939
R14383 gnd.n2476 gnd.n2475 0.152939
R14384 gnd.n2477 gnd.n2476 0.152939
R14385 gnd.n2478 gnd.n2477 0.152939
R14386 gnd.n2483 gnd.n2478 0.152939
R14387 gnd.n2484 gnd.n2483 0.152939
R14388 gnd.n2485 gnd.n2484 0.152939
R14389 gnd.n2486 gnd.n2485 0.152939
R14390 gnd.n2491 gnd.n2486 0.152939
R14391 gnd.n2492 gnd.n2491 0.152939
R14392 gnd.n2493 gnd.n2492 0.152939
R14393 gnd.n2494 gnd.n2493 0.152939
R14394 gnd.n2499 gnd.n2494 0.152939
R14395 gnd.n2500 gnd.n2499 0.152939
R14396 gnd.n2501 gnd.n2500 0.152939
R14397 gnd.n2502 gnd.n2501 0.152939
R14398 gnd.n2507 gnd.n2502 0.152939
R14399 gnd.n2508 gnd.n2507 0.152939
R14400 gnd.n2509 gnd.n2508 0.152939
R14401 gnd.n2510 gnd.n2509 0.152939
R14402 gnd.n2515 gnd.n2510 0.152939
R14403 gnd.n2516 gnd.n2515 0.152939
R14404 gnd.n2517 gnd.n2516 0.152939
R14405 gnd.n2518 gnd.n2517 0.152939
R14406 gnd.n2523 gnd.n2518 0.152939
R14407 gnd.n2524 gnd.n2523 0.152939
R14408 gnd.n2525 gnd.n2524 0.152939
R14409 gnd.n2526 gnd.n2525 0.152939
R14410 gnd.n2531 gnd.n2526 0.152939
R14411 gnd.n2532 gnd.n2531 0.152939
R14412 gnd.n2533 gnd.n2532 0.152939
R14413 gnd.n2534 gnd.n2533 0.152939
R14414 gnd.n2539 gnd.n2534 0.152939
R14415 gnd.n2540 gnd.n2539 0.152939
R14416 gnd.n2541 gnd.n2540 0.152939
R14417 gnd.n2542 gnd.n2541 0.152939
R14418 gnd.n2547 gnd.n2542 0.152939
R14419 gnd.n2548 gnd.n2547 0.152939
R14420 gnd.n2549 gnd.n2548 0.152939
R14421 gnd.n2550 gnd.n2549 0.152939
R14422 gnd.n2555 gnd.n2550 0.152939
R14423 gnd.n2556 gnd.n2555 0.152939
R14424 gnd.n2557 gnd.n2556 0.152939
R14425 gnd.n2558 gnd.n2557 0.152939
R14426 gnd.n2563 gnd.n2558 0.152939
R14427 gnd.n2564 gnd.n2563 0.152939
R14428 gnd.n2565 gnd.n2564 0.152939
R14429 gnd.n2566 gnd.n2565 0.152939
R14430 gnd.n2571 gnd.n2566 0.152939
R14431 gnd.n2572 gnd.n2571 0.152939
R14432 gnd.n2573 gnd.n2572 0.152939
R14433 gnd.n2574 gnd.n2573 0.152939
R14434 gnd.n2579 gnd.n2574 0.152939
R14435 gnd.n2580 gnd.n2579 0.152939
R14436 gnd.n2581 gnd.n2580 0.152939
R14437 gnd.n2582 gnd.n2581 0.152939
R14438 gnd.n2587 gnd.n2582 0.152939
R14439 gnd.n2588 gnd.n2587 0.152939
R14440 gnd.n2589 gnd.n2588 0.152939
R14441 gnd.n2590 gnd.n2589 0.152939
R14442 gnd.n2595 gnd.n2590 0.152939
R14443 gnd.n2596 gnd.n2595 0.152939
R14444 gnd.n2597 gnd.n2596 0.152939
R14445 gnd.n2598 gnd.n2597 0.152939
R14446 gnd.n2599 gnd.n2598 0.152939
R14447 gnd.n7749 gnd.n108 0.152939
R14448 gnd.n133 gnd.n108 0.152939
R14449 gnd.n134 gnd.n133 0.152939
R14450 gnd.n135 gnd.n134 0.152939
R14451 gnd.n150 gnd.n135 0.152939
R14452 gnd.n151 gnd.n150 0.152939
R14453 gnd.n152 gnd.n151 0.152939
R14454 gnd.n153 gnd.n152 0.152939
R14455 gnd.n170 gnd.n153 0.152939
R14456 gnd.n171 gnd.n170 0.152939
R14457 gnd.n172 gnd.n171 0.152939
R14458 gnd.n173 gnd.n172 0.152939
R14459 gnd.n188 gnd.n173 0.152939
R14460 gnd.n189 gnd.n188 0.152939
R14461 gnd.n190 gnd.n189 0.152939
R14462 gnd.n191 gnd.n190 0.152939
R14463 gnd.n208 gnd.n191 0.152939
R14464 gnd.n209 gnd.n208 0.152939
R14465 gnd.n210 gnd.n209 0.152939
R14466 gnd.n211 gnd.n210 0.152939
R14467 gnd.n227 gnd.n211 0.152939
R14468 gnd.n228 gnd.n227 0.152939
R14469 gnd.n229 gnd.n228 0.152939
R14470 gnd.n230 gnd.n229 0.152939
R14471 gnd.n246 gnd.n230 0.152939
R14472 gnd.n247 gnd.n246 0.152939
R14473 gnd.n7664 gnd.n247 0.152939
R14474 gnd.n7758 gnd.n97 0.152939
R14475 gnd.n351 gnd.n97 0.152939
R14476 gnd.n7363 gnd.n351 0.152939
R14477 gnd.n7364 gnd.n7363 0.152939
R14478 gnd.n7365 gnd.n7364 0.152939
R14479 gnd.n7366 gnd.n7365 0.152939
R14480 gnd.n7367 gnd.n7366 0.152939
R14481 gnd.n7368 gnd.n7367 0.152939
R14482 gnd.n7369 gnd.n7368 0.152939
R14483 gnd.n7370 gnd.n7369 0.152939
R14484 gnd.n7371 gnd.n7370 0.152939
R14485 gnd.n7372 gnd.n7371 0.152939
R14486 gnd.n7373 gnd.n7372 0.152939
R14487 gnd.n7374 gnd.n7373 0.152939
R14488 gnd.n7375 gnd.n7374 0.152939
R14489 gnd.n7376 gnd.n7375 0.152939
R14490 gnd.n7377 gnd.n7376 0.152939
R14491 gnd.n7378 gnd.n7377 0.152939
R14492 gnd.n7379 gnd.n7378 0.152939
R14493 gnd.n7380 gnd.n7379 0.152939
R14494 gnd.n7381 gnd.n7380 0.152939
R14495 gnd.n7382 gnd.n7381 0.152939
R14496 gnd.n7383 gnd.n7382 0.152939
R14497 gnd.n7384 gnd.n7383 0.152939
R14498 gnd.n7385 gnd.n7384 0.152939
R14499 gnd.n7386 gnd.n7385 0.152939
R14500 gnd.n7387 gnd.n7386 0.152939
R14501 gnd.n7388 gnd.n7387 0.152939
R14502 gnd.n7389 gnd.n7388 0.152939
R14503 gnd.n7390 gnd.n7389 0.152939
R14504 gnd.n7391 gnd.n7390 0.152939
R14505 gnd.n7405 gnd.n348 0.152939
R14506 gnd.n7406 gnd.n7405 0.152939
R14507 gnd.n7406 gnd.n7401 0.152939
R14508 gnd.n7414 gnd.n7401 0.152939
R14509 gnd.n7415 gnd.n7414 0.152939
R14510 gnd.n7416 gnd.n7415 0.152939
R14511 gnd.n7416 gnd.n7399 0.152939
R14512 gnd.n7424 gnd.n7399 0.152939
R14513 gnd.n7425 gnd.n7424 0.152939
R14514 gnd.n7426 gnd.n7425 0.152939
R14515 gnd.n7426 gnd.n7397 0.152939
R14516 gnd.n7434 gnd.n7397 0.152939
R14517 gnd.n7435 gnd.n7434 0.152939
R14518 gnd.n7436 gnd.n7435 0.152939
R14519 gnd.n7436 gnd.n7395 0.152939
R14520 gnd.n7444 gnd.n7395 0.152939
R14521 gnd.n7445 gnd.n7444 0.152939
R14522 gnd.n7446 gnd.n7445 0.152939
R14523 gnd.n7663 gnd.n248 0.152939
R14524 gnd.n290 gnd.n248 0.152939
R14525 gnd.n291 gnd.n290 0.152939
R14526 gnd.n292 gnd.n291 0.152939
R14527 gnd.n293 gnd.n292 0.152939
R14528 gnd.n294 gnd.n293 0.152939
R14529 gnd.n295 gnd.n294 0.152939
R14530 gnd.n296 gnd.n295 0.152939
R14531 gnd.n297 gnd.n296 0.152939
R14532 gnd.n298 gnd.n297 0.152939
R14533 gnd.n299 gnd.n298 0.152939
R14534 gnd.n300 gnd.n299 0.152939
R14535 gnd.n301 gnd.n300 0.152939
R14536 gnd.n302 gnd.n301 0.152939
R14537 gnd.n303 gnd.n302 0.152939
R14538 gnd.n304 gnd.n303 0.152939
R14539 gnd.n305 gnd.n304 0.152939
R14540 gnd.n306 gnd.n305 0.152939
R14541 gnd.n307 gnd.n306 0.152939
R14542 gnd.n308 gnd.n307 0.152939
R14543 gnd.n309 gnd.n308 0.152939
R14544 gnd.n310 gnd.n309 0.152939
R14545 gnd.n311 gnd.n310 0.152939
R14546 gnd.n312 gnd.n311 0.152939
R14547 gnd.n313 gnd.n312 0.152939
R14548 gnd.n314 gnd.n313 0.152939
R14549 gnd.n315 gnd.n314 0.152939
R14550 gnd.n316 gnd.n315 0.152939
R14551 gnd.n317 gnd.n316 0.152939
R14552 gnd.n318 gnd.n317 0.152939
R14553 gnd.n319 gnd.n318 0.152939
R14554 gnd.n320 gnd.n319 0.152939
R14555 gnd.n321 gnd.n320 0.152939
R14556 gnd.n322 gnd.n321 0.152939
R14557 gnd.n323 gnd.n322 0.152939
R14558 gnd.n324 gnd.n323 0.152939
R14559 gnd.n7584 gnd.n324 0.152939
R14560 gnd.n7584 gnd.n7583 0.152939
R14561 gnd.n7583 gnd.n7582 0.152939
R14562 gnd.n7582 gnd.n328 0.152939
R14563 gnd.n329 gnd.n328 0.152939
R14564 gnd.n330 gnd.n329 0.152939
R14565 gnd.n331 gnd.n330 0.152939
R14566 gnd.n332 gnd.n331 0.152939
R14567 gnd.n333 gnd.n332 0.152939
R14568 gnd.n334 gnd.n333 0.152939
R14569 gnd.n335 gnd.n334 0.152939
R14570 gnd.n336 gnd.n335 0.152939
R14571 gnd.n337 gnd.n336 0.152939
R14572 gnd.n338 gnd.n337 0.152939
R14573 gnd.n339 gnd.n338 0.152939
R14574 gnd.n340 gnd.n339 0.152939
R14575 gnd.n341 gnd.n340 0.152939
R14576 gnd.n342 gnd.n341 0.152939
R14577 gnd.n343 gnd.n342 0.152939
R14578 gnd.n344 gnd.n343 0.152939
R14579 gnd.n7542 gnd.n344 0.152939
R14580 gnd.n7542 gnd.n7541 0.152939
R14581 gnd.n630 gnd.n567 0.152939
R14582 gnd.n631 gnd.n630 0.152939
R14583 gnd.n632 gnd.n631 0.152939
R14584 gnd.n633 gnd.n632 0.152939
R14585 gnd.n634 gnd.n633 0.152939
R14586 gnd.n635 gnd.n634 0.152939
R14587 gnd.n636 gnd.n635 0.152939
R14588 gnd.n637 gnd.n636 0.152939
R14589 gnd.n638 gnd.n637 0.152939
R14590 gnd.n639 gnd.n638 0.152939
R14591 gnd.n640 gnd.n639 0.152939
R14592 gnd.n641 gnd.n640 0.152939
R14593 gnd.n642 gnd.n641 0.152939
R14594 gnd.n643 gnd.n642 0.152939
R14595 gnd.n644 gnd.n643 0.152939
R14596 gnd.n645 gnd.n644 0.152939
R14597 gnd.n646 gnd.n645 0.152939
R14598 gnd.n649 gnd.n646 0.152939
R14599 gnd.n650 gnd.n649 0.152939
R14600 gnd.n651 gnd.n650 0.152939
R14601 gnd.n652 gnd.n651 0.152939
R14602 gnd.n653 gnd.n652 0.152939
R14603 gnd.n654 gnd.n653 0.152939
R14604 gnd.n655 gnd.n654 0.152939
R14605 gnd.n656 gnd.n655 0.152939
R14606 gnd.n661 gnd.n660 0.152939
R14607 gnd.n662 gnd.n661 0.152939
R14608 gnd.n663 gnd.n662 0.152939
R14609 gnd.n664 gnd.n663 0.152939
R14610 gnd.n665 gnd.n664 0.152939
R14611 gnd.n666 gnd.n665 0.152939
R14612 gnd.n667 gnd.n666 0.152939
R14613 gnd.n668 gnd.n667 0.152939
R14614 gnd.n669 gnd.n668 0.152939
R14615 gnd.n672 gnd.n669 0.152939
R14616 gnd.n673 gnd.n672 0.152939
R14617 gnd.n674 gnd.n673 0.152939
R14618 gnd.n675 gnd.n674 0.152939
R14619 gnd.n676 gnd.n675 0.152939
R14620 gnd.n677 gnd.n676 0.152939
R14621 gnd.n678 gnd.n677 0.152939
R14622 gnd.n679 gnd.n678 0.152939
R14623 gnd.n680 gnd.n679 0.152939
R14624 gnd.n681 gnd.n680 0.152939
R14625 gnd.n682 gnd.n681 0.152939
R14626 gnd.n683 gnd.n682 0.152939
R14627 gnd.n684 gnd.n683 0.152939
R14628 gnd.n685 gnd.n684 0.152939
R14629 gnd.n686 gnd.n685 0.152939
R14630 gnd.n687 gnd.n686 0.152939
R14631 gnd.n688 gnd.n687 0.152939
R14632 gnd.n689 gnd.n688 0.152939
R14633 gnd.n690 gnd.n689 0.152939
R14634 gnd.n6928 gnd.n690 0.152939
R14635 gnd.n6928 gnd.n6927 0.152939
R14636 gnd.n7072 gnd.n7071 0.152939
R14637 gnd.n7073 gnd.n7072 0.152939
R14638 gnd.n7074 gnd.n7073 0.152939
R14639 gnd.n7074 gnd.n528 0.152939
R14640 gnd.n7121 gnd.n528 0.152939
R14641 gnd.n7122 gnd.n7121 0.152939
R14642 gnd.n7123 gnd.n7122 0.152939
R14643 gnd.n7124 gnd.n7123 0.152939
R14644 gnd.n7124 gnd.n494 0.152939
R14645 gnd.n7156 gnd.n494 0.152939
R14646 gnd.n7157 gnd.n7156 0.152939
R14647 gnd.n7158 gnd.n7157 0.152939
R14648 gnd.n7158 gnd.n463 0.152939
R14649 gnd.n7191 gnd.n463 0.152939
R14650 gnd.n7192 gnd.n7191 0.152939
R14651 gnd.n7193 gnd.n7192 0.152939
R14652 gnd.n7194 gnd.n7193 0.152939
R14653 gnd.n7194 gnd.n436 0.152939
R14654 gnd.n7231 gnd.n436 0.152939
R14655 gnd.n7232 gnd.n7231 0.152939
R14656 gnd.n7233 gnd.n7232 0.152939
R14657 gnd.n7233 gnd.n409 0.152939
R14658 gnd.n7278 gnd.n409 0.152939
R14659 gnd.n7279 gnd.n7278 0.152939
R14660 gnd.n7280 gnd.n7279 0.152939
R14661 gnd.n7280 gnd.n109 0.152939
R14662 gnd.n7749 gnd.n109 0.152939
R14663 gnd.n1922 gnd.n1919 0.152939
R14664 gnd.n1923 gnd.n1922 0.152939
R14665 gnd.n1924 gnd.n1923 0.152939
R14666 gnd.n1925 gnd.n1924 0.152939
R14667 gnd.n1928 gnd.n1925 0.152939
R14668 gnd.n1929 gnd.n1928 0.152939
R14669 gnd.n1930 gnd.n1929 0.152939
R14670 gnd.n1931 gnd.n1930 0.152939
R14671 gnd.n1934 gnd.n1931 0.152939
R14672 gnd.n1935 gnd.n1934 0.152939
R14673 gnd.n1936 gnd.n1935 0.152939
R14674 gnd.n1938 gnd.n1936 0.152939
R14675 gnd.n1938 gnd.n1937 0.152939
R14676 gnd.n1937 gnd.n1546 0.152939
R14677 gnd.n5392 gnd.n1546 0.152939
R14678 gnd.n5393 gnd.n5392 0.152939
R14679 gnd.n5394 gnd.n5393 0.152939
R14680 gnd.n5395 gnd.n5394 0.152939
R14681 gnd.n5396 gnd.n5395 0.152939
R14682 gnd.n5396 gnd.n1495 0.152939
R14683 gnd.n5456 gnd.n1495 0.152939
R14684 gnd.n5457 gnd.n5456 0.152939
R14685 gnd.n5458 gnd.n5457 0.152939
R14686 gnd.n5458 gnd.n1491 0.152939
R14687 gnd.n5464 gnd.n1491 0.152939
R14688 gnd.n5465 gnd.n5464 0.152939
R14689 gnd.n5466 gnd.n5465 0.152939
R14690 gnd.n5467 gnd.n5466 0.152939
R14691 gnd.n5468 gnd.n5467 0.152939
R14692 gnd.n5471 gnd.n5468 0.152939
R14693 gnd.n5472 gnd.n5471 0.152939
R14694 gnd.n5473 gnd.n5472 0.152939
R14695 gnd.n5474 gnd.n5473 0.152939
R14696 gnd.n5546 gnd.n5474 0.152939
R14697 gnd.n5547 gnd.n5546 0.152939
R14698 gnd.n5571 gnd.n5547 0.152939
R14699 gnd.n5572 gnd.n5571 0.152939
R14700 gnd.n5573 gnd.n5572 0.152939
R14701 gnd.n5573 gnd.n5534 0.152939
R14702 gnd.n5592 gnd.n5534 0.152939
R14703 gnd.n5593 gnd.n5592 0.152939
R14704 gnd.n5594 gnd.n5593 0.152939
R14705 gnd.n5594 gnd.n5522 0.152939
R14706 gnd.n5613 gnd.n5522 0.152939
R14707 gnd.n5614 gnd.n5613 0.152939
R14708 gnd.n5615 gnd.n5614 0.152939
R14709 gnd.n5615 gnd.n5509 0.152939
R14710 gnd.n5642 gnd.n5509 0.152939
R14711 gnd.n5643 gnd.n5642 0.152939
R14712 gnd.n5644 gnd.n5643 0.152939
R14713 gnd.n5645 gnd.n5644 0.152939
R14714 gnd.n5646 gnd.n5645 0.152939
R14715 gnd.n5646 gnd.n1197 0.152939
R14716 gnd.n6157 gnd.n1197 0.152939
R14717 gnd.n6158 gnd.n6157 0.152939
R14718 gnd.n6159 gnd.n6158 0.152939
R14719 gnd.n6159 gnd.n1171 0.152939
R14720 gnd.n6198 gnd.n1171 0.152939
R14721 gnd.n6199 gnd.n6198 0.152939
R14722 gnd.n6200 gnd.n6199 0.152939
R14723 gnd.n6201 gnd.n6200 0.152939
R14724 gnd.n6202 gnd.n6201 0.152939
R14725 gnd.n6202 gnd.n1149 0.152939
R14726 gnd.n6226 gnd.n1149 0.152939
R14727 gnd.n6227 gnd.n6226 0.152939
R14728 gnd.n6229 gnd.n6227 0.152939
R14729 gnd.n6229 gnd.n6228 0.152939
R14730 gnd.n6228 gnd.n1121 0.152939
R14731 gnd.n1122 gnd.n1121 0.152939
R14732 gnd.n1124 gnd.n1122 0.152939
R14733 gnd.n1124 gnd.n1123 0.152939
R14734 gnd.n1123 gnd.n1089 0.152939
R14735 gnd.n1090 gnd.n1089 0.152939
R14736 gnd.n1092 gnd.n1090 0.152939
R14737 gnd.n1092 gnd.n1091 0.152939
R14738 gnd.n1091 gnd.n1062 0.152939
R14739 gnd.n1063 gnd.n1062 0.152939
R14740 gnd.n1065 gnd.n1063 0.152939
R14741 gnd.n1065 gnd.n1064 0.152939
R14742 gnd.n1064 gnd.n1032 0.152939
R14743 gnd.n1033 gnd.n1032 0.152939
R14744 gnd.n1034 gnd.n1033 0.152939
R14745 gnd.n1036 gnd.n1034 0.152939
R14746 gnd.n1036 gnd.n1035 0.152939
R14747 gnd.n1035 gnd.n986 0.152939
R14748 gnd.n987 gnd.n986 0.152939
R14749 gnd.n988 gnd.n987 0.152939
R14750 gnd.n989 gnd.n988 0.152939
R14751 gnd.n989 gnd.n942 0.152939
R14752 gnd.n6542 gnd.n942 0.152939
R14753 gnd.n6543 gnd.n6542 0.152939
R14754 gnd.n6544 gnd.n6543 0.152939
R14755 gnd.n6544 gnd.n888 0.152939
R14756 gnd.n6718 gnd.n888 0.152939
R14757 gnd.n6719 gnd.n6718 0.152939
R14758 gnd.n6720 gnd.n6719 0.152939
R14759 gnd.n6721 gnd.n6720 0.152939
R14760 gnd.n6721 gnd.n864 0.152939
R14761 gnd.n6748 gnd.n864 0.152939
R14762 gnd.n6749 gnd.n6748 0.152939
R14763 gnd.n6750 gnd.n6749 0.152939
R14764 gnd.n6751 gnd.n6750 0.152939
R14765 gnd.n6751 gnd.n839 0.152939
R14766 gnd.n6778 gnd.n839 0.152939
R14767 gnd.n6779 gnd.n6778 0.152939
R14768 gnd.n6780 gnd.n6779 0.152939
R14769 gnd.n6781 gnd.n6780 0.152939
R14770 gnd.n6781 gnd.n814 0.152939
R14771 gnd.n6813 gnd.n814 0.152939
R14772 gnd.n6814 gnd.n6813 0.152939
R14773 gnd.n6815 gnd.n6814 0.152939
R14774 gnd.n6817 gnd.n6815 0.152939
R14775 gnd.n6817 gnd.n6816 0.152939
R14776 gnd.n6816 gnd.n798 0.152939
R14777 gnd.n6837 gnd.n798 0.152939
R14778 gnd.n6838 gnd.n6837 0.152939
R14779 gnd.n6839 gnd.n6838 0.152939
R14780 gnd.n6840 gnd.n6839 0.152939
R14781 gnd.n6840 gnd.n586 0.152939
R14782 gnd.n7046 gnd.n586 0.152939
R14783 gnd.n7047 gnd.n7046 0.152939
R14784 gnd.n7048 gnd.n7047 0.152939
R14785 gnd.n7049 gnd.n7048 0.152939
R14786 gnd.n7050 gnd.n7049 0.152939
R14787 gnd.n7051 gnd.n7050 0.152939
R14788 gnd.n7051 gnd.n548 0.152939
R14789 gnd.n7103 gnd.n548 0.152939
R14790 gnd.n7104 gnd.n7103 0.152939
R14791 gnd.n7105 gnd.n7104 0.152939
R14792 gnd.n7106 gnd.n7105 0.152939
R14793 gnd.n7106 gnd.n484 0.152939
R14794 gnd.n7165 gnd.n484 0.152939
R14795 gnd.n7166 gnd.n7165 0.152939
R14796 gnd.n7167 gnd.n7166 0.152939
R14797 gnd.n7167 gnd.n480 0.152939
R14798 gnd.n7173 gnd.n480 0.152939
R14799 gnd.n7174 gnd.n7173 0.152939
R14800 gnd.n7175 gnd.n7174 0.152939
R14801 gnd.n7176 gnd.n7175 0.152939
R14802 gnd.n7176 gnd.n428 0.152939
R14803 gnd.n7240 gnd.n428 0.152939
R14804 gnd.n7241 gnd.n7240 0.152939
R14805 gnd.n7242 gnd.n7241 0.152939
R14806 gnd.n7243 gnd.n7242 0.152939
R14807 gnd.n7244 gnd.n7243 0.152939
R14808 gnd.n7246 gnd.n7244 0.152939
R14809 gnd.n7247 gnd.n7246 0.152939
R14810 gnd.n4780 gnd.n4759 0.152939
R14811 gnd.n4760 gnd.n4759 0.152939
R14812 gnd.n4761 gnd.n4760 0.152939
R14813 gnd.n4762 gnd.n4761 0.152939
R14814 gnd.n4763 gnd.n4762 0.152939
R14815 gnd.n4764 gnd.n4763 0.152939
R14816 gnd.n4765 gnd.n4764 0.152939
R14817 gnd.n4766 gnd.n4765 0.152939
R14818 gnd.n4766 gnd.n1772 0.152939
R14819 gnd.n5100 gnd.n1772 0.152939
R14820 gnd.n5101 gnd.n5100 0.152939
R14821 gnd.n5102 gnd.n5101 0.152939
R14822 gnd.n5103 gnd.n5102 0.152939
R14823 gnd.n5103 gnd.n1747 0.152939
R14824 gnd.n5135 gnd.n1747 0.152939
R14825 gnd.n5136 gnd.n5135 0.152939
R14826 gnd.n5137 gnd.n5136 0.152939
R14827 gnd.n5138 gnd.n5137 0.152939
R14828 gnd.n5138 gnd.n1722 0.152939
R14829 gnd.n5170 gnd.n1722 0.152939
R14830 gnd.n5171 gnd.n5170 0.152939
R14831 gnd.n5172 gnd.n5171 0.152939
R14832 gnd.n5173 gnd.n5172 0.152939
R14833 gnd.n5173 gnd.n1695 0.152939
R14834 gnd.n5207 gnd.n1695 0.152939
R14835 gnd.n5208 gnd.n5207 0.152939
R14836 gnd.n5209 gnd.n5208 0.152939
R14837 gnd.n5210 gnd.n5209 0.152939
R14838 gnd.n5210 gnd.n1676 0.152939
R14839 gnd.n5232 gnd.n1676 0.152939
R14840 gnd.n5233 gnd.n5232 0.152939
R14841 gnd.n4821 gnd.n4733 0.152939
R14842 gnd.n4736 gnd.n4733 0.152939
R14843 gnd.n4737 gnd.n4736 0.152939
R14844 gnd.n4738 gnd.n4737 0.152939
R14845 gnd.n4739 gnd.n4738 0.152939
R14846 gnd.n4742 gnd.n4739 0.152939
R14847 gnd.n4743 gnd.n4742 0.152939
R14848 gnd.n4744 gnd.n4743 0.152939
R14849 gnd.n4745 gnd.n4744 0.152939
R14850 gnd.n4748 gnd.n4745 0.152939
R14851 gnd.n4749 gnd.n4748 0.152939
R14852 gnd.n4750 gnd.n4749 0.152939
R14853 gnd.n4751 gnd.n4750 0.152939
R14854 gnd.n4754 gnd.n4751 0.152939
R14855 gnd.n4755 gnd.n4754 0.152939
R14856 gnd.n4787 gnd.n4755 0.152939
R14857 gnd.n4787 gnd.n4786 0.152939
R14858 gnd.n4786 gnd.n4785 0.152939
R14859 gnd.n5293 gnd.n5292 0.152939
R14860 gnd.n5294 gnd.n5293 0.152939
R14861 gnd.n5295 gnd.n5294 0.152939
R14862 gnd.n5295 gnd.n1596 0.152939
R14863 gnd.n5328 gnd.n1596 0.152939
R14864 gnd.n5329 gnd.n5328 0.152939
R14865 gnd.n5330 gnd.n5329 0.152939
R14866 gnd.n5331 gnd.n5330 0.152939
R14867 gnd.n5331 gnd.n1565 0.152939
R14868 gnd.n5370 gnd.n1565 0.152939
R14869 gnd.n5371 gnd.n5370 0.152939
R14870 gnd.n5372 gnd.n5371 0.152939
R14871 gnd.n5373 gnd.n5372 0.152939
R14872 gnd.n5373 gnd.n1529 0.152939
R14873 gnd.n5413 gnd.n1529 0.152939
R14874 gnd.n5414 gnd.n5413 0.152939
R14875 gnd.n5415 gnd.n5414 0.152939
R14876 gnd.n5416 gnd.n5415 0.152939
R14877 gnd.n5416 gnd.n1502 0.152939
R14878 gnd.n5447 gnd.n1502 0.152939
R14879 gnd.n5448 gnd.n5447 0.152939
R14880 gnd.n5449 gnd.n5448 0.152939
R14881 gnd.n5449 gnd.n1433 0.152939
R14882 gnd.n5867 gnd.n1433 0.152939
R14883 gnd.n5868 gnd.n5867 0.152939
R14884 gnd.n5869 gnd.n5868 0.152939
R14885 gnd.n5962 gnd.n5869 0.152939
R14886 gnd.n5961 gnd.n5870 0.152939
R14887 gnd.n5873 gnd.n5870 0.152939
R14888 gnd.n5874 gnd.n5873 0.152939
R14889 gnd.n5875 gnd.n5874 0.152939
R14890 gnd.n5879 gnd.n5875 0.152939
R14891 gnd.n5880 gnd.n5879 0.152939
R14892 gnd.n5881 gnd.n5880 0.152939
R14893 gnd.n5882 gnd.n5881 0.152939
R14894 gnd.n5886 gnd.n5882 0.152939
R14895 gnd.n5887 gnd.n5886 0.152939
R14896 gnd.n5888 gnd.n5887 0.152939
R14897 gnd.n5889 gnd.n5888 0.152939
R14898 gnd.n5893 gnd.n5889 0.152939
R14899 gnd.n5894 gnd.n5893 0.152939
R14900 gnd.n5895 gnd.n5894 0.152939
R14901 gnd.n5896 gnd.n5895 0.152939
R14902 gnd.n5903 gnd.n5896 0.152939
R14903 gnd.n5904 gnd.n5903 0.152939
R14904 gnd.n5905 gnd.n5904 0.152939
R14905 gnd.n5906 gnd.n5905 0.152939
R14906 gnd.n5910 gnd.n5906 0.152939
R14907 gnd.n5911 gnd.n5910 0.152939
R14908 gnd.n5912 gnd.n5911 0.152939
R14909 gnd.n5913 gnd.n5912 0.152939
R14910 gnd.n5913 gnd.n1364 0.152939
R14911 gnd.n6029 gnd.n6028 0.152939
R14912 gnd.n6028 gnd.n1365 0.152939
R14913 gnd.n1372 gnd.n1365 0.152939
R14914 gnd.n1373 gnd.n1372 0.152939
R14915 gnd.n1374 gnd.n1373 0.152939
R14916 gnd.n1375 gnd.n1374 0.152939
R14917 gnd.n1379 gnd.n1375 0.152939
R14918 gnd.n1380 gnd.n1379 0.152939
R14919 gnd.n6011 gnd.n1380 0.152939
R14920 gnd.n6011 gnd.n6010 0.152939
R14921 gnd.n6010 gnd.n6009 0.152939
R14922 gnd.n6009 gnd.n1384 0.152939
R14923 gnd.n1390 gnd.n1384 0.152939
R14924 gnd.n1391 gnd.n1390 0.152939
R14925 gnd.n1392 gnd.n1391 0.152939
R14926 gnd.n1393 gnd.n1392 0.152939
R14927 gnd.n1397 gnd.n1393 0.152939
R14928 gnd.n1398 gnd.n1397 0.152939
R14929 gnd.n1399 gnd.n1398 0.152939
R14930 gnd.n1400 gnd.n1399 0.152939
R14931 gnd.n1404 gnd.n1400 0.152939
R14932 gnd.n1405 gnd.n1404 0.152939
R14933 gnd.n1406 gnd.n1405 0.152939
R14934 gnd.n1407 gnd.n1406 0.152939
R14935 gnd.n1411 gnd.n1407 0.152939
R14936 gnd.n1412 gnd.n1411 0.152939
R14937 gnd.n1413 gnd.n1412 0.152939
R14938 gnd.n1414 gnd.n1413 0.152939
R14939 gnd.n1420 gnd.n1414 0.152939
R14940 gnd.n5972 gnd.n1420 0.152939
R14941 gnd.n4888 gnd.n1817 0.152939
R14942 gnd.n4889 gnd.n4888 0.152939
R14943 gnd.n4890 gnd.n4889 0.152939
R14944 gnd.n4890 gnd.n4880 0.152939
R14945 gnd.n4898 gnd.n4880 0.152939
R14946 gnd.n4899 gnd.n4898 0.152939
R14947 gnd.n4900 gnd.n4899 0.152939
R14948 gnd.n4900 gnd.n4876 0.152939
R14949 gnd.n4908 gnd.n4876 0.152939
R14950 gnd.n4909 gnd.n4908 0.152939
R14951 gnd.n4910 gnd.n4909 0.152939
R14952 gnd.n4910 gnd.n4872 0.152939
R14953 gnd.n4918 gnd.n4872 0.152939
R14954 gnd.n4919 gnd.n4918 0.152939
R14955 gnd.n4920 gnd.n4919 0.152939
R14956 gnd.n4920 gnd.n4865 0.152939
R14957 gnd.n4928 gnd.n4865 0.152939
R14958 gnd.n4929 gnd.n4928 0.152939
R14959 gnd.n4930 gnd.n4929 0.152939
R14960 gnd.n4930 gnd.n4861 0.152939
R14961 gnd.n4938 gnd.n4861 0.152939
R14962 gnd.n4939 gnd.n4938 0.152939
R14963 gnd.n4940 gnd.n4939 0.152939
R14964 gnd.n4940 gnd.n4857 0.152939
R14965 gnd.n4948 gnd.n4857 0.152939
R14966 gnd.n4949 gnd.n4948 0.152939
R14967 gnd.n4950 gnd.n4949 0.152939
R14968 gnd.n4950 gnd.n4853 0.152939
R14969 gnd.n4958 gnd.n4853 0.152939
R14970 gnd.n4959 gnd.n4958 0.152939
R14971 gnd.n4960 gnd.n4959 0.152939
R14972 gnd.n4960 gnd.n4849 0.152939
R14973 gnd.n4968 gnd.n4849 0.152939
R14974 gnd.n4969 gnd.n4968 0.152939
R14975 gnd.n4970 gnd.n4969 0.152939
R14976 gnd.n4970 gnd.n4845 0.152939
R14977 gnd.n4980 gnd.n4845 0.152939
R14978 gnd.n4981 gnd.n4980 0.152939
R14979 gnd.n4982 gnd.n4981 0.152939
R14980 gnd.n4982 gnd.n4841 0.152939
R14981 gnd.n4990 gnd.n4841 0.152939
R14982 gnd.n4991 gnd.n4990 0.152939
R14983 gnd.n4992 gnd.n4991 0.152939
R14984 gnd.n4992 gnd.n4837 0.152939
R14985 gnd.n5000 gnd.n4837 0.152939
R14986 gnd.n5001 gnd.n5000 0.152939
R14987 gnd.n5002 gnd.n5001 0.152939
R14988 gnd.n5002 gnd.n4833 0.152939
R14989 gnd.n5010 gnd.n4833 0.152939
R14990 gnd.n5011 gnd.n5010 0.152939
R14991 gnd.n5012 gnd.n5011 0.152939
R14992 gnd.n5012 gnd.n4829 0.152939
R14993 gnd.n5020 gnd.n4829 0.152939
R14994 gnd.n5021 gnd.n5020 0.152939
R14995 gnd.n5023 gnd.n5021 0.152939
R14996 gnd.n5023 gnd.n5022 0.152939
R14997 gnd.n5022 gnd.n4822 0.152939
R14998 gnd.n5032 gnd.n4822 0.152939
R14999 gnd.n5047 gnd.n5046 0.152939
R15000 gnd.n5048 gnd.n5047 0.152939
R15001 gnd.n5048 gnd.n1800 0.152939
R15002 gnd.n5066 gnd.n1800 0.152939
R15003 gnd.n5067 gnd.n5066 0.152939
R15004 gnd.n5068 gnd.n5067 0.152939
R15005 gnd.n5068 gnd.n1780 0.152939
R15006 gnd.n5090 gnd.n1780 0.152939
R15007 gnd.n5091 gnd.n5090 0.152939
R15008 gnd.n5092 gnd.n5091 0.152939
R15009 gnd.n5093 gnd.n5092 0.152939
R15010 gnd.n5093 gnd.n1755 0.152939
R15011 gnd.n5125 gnd.n1755 0.152939
R15012 gnd.n5126 gnd.n5125 0.152939
R15013 gnd.n5127 gnd.n5126 0.152939
R15014 gnd.n5128 gnd.n5127 0.152939
R15015 gnd.n5128 gnd.n1731 0.152939
R15016 gnd.n5160 gnd.n1731 0.152939
R15017 gnd.n5161 gnd.n5160 0.152939
R15018 gnd.n5162 gnd.n5161 0.152939
R15019 gnd.n5163 gnd.n5162 0.152939
R15020 gnd.n5163 gnd.n1704 0.152939
R15021 gnd.n5197 gnd.n1704 0.152939
R15022 gnd.n5198 gnd.n5197 0.152939
R15023 gnd.n5199 gnd.n5198 0.152939
R15024 gnd.n5199 gnd.n1625 0.152939
R15025 gnd.n5292 gnd.n1625 0.152939
R15026 gnd.n3115 gnd.n2096 0.152939
R15027 gnd.n3116 gnd.n3115 0.152939
R15028 gnd.n3117 gnd.n3116 0.152939
R15029 gnd.n3117 gnd.n2090 0.152939
R15030 gnd.n3125 gnd.n2090 0.152939
R15031 gnd.n3126 gnd.n3125 0.152939
R15032 gnd.n3127 gnd.n3126 0.152939
R15033 gnd.n3127 gnd.n2084 0.152939
R15034 gnd.n3135 gnd.n2084 0.152939
R15035 gnd.n3136 gnd.n3135 0.152939
R15036 gnd.n3137 gnd.n3136 0.152939
R15037 gnd.n3137 gnd.n2078 0.152939
R15038 gnd.n3145 gnd.n2078 0.152939
R15039 gnd.n3146 gnd.n3145 0.152939
R15040 gnd.n3147 gnd.n3146 0.152939
R15041 gnd.n3147 gnd.n2072 0.152939
R15042 gnd.n3155 gnd.n2072 0.152939
R15043 gnd.n3156 gnd.n3155 0.152939
R15044 gnd.n3157 gnd.n3156 0.152939
R15045 gnd.n3157 gnd.n2066 0.152939
R15046 gnd.n3165 gnd.n2066 0.152939
R15047 gnd.n3166 gnd.n3165 0.152939
R15048 gnd.n3167 gnd.n3166 0.152939
R15049 gnd.n3167 gnd.n2060 0.152939
R15050 gnd.n3175 gnd.n2060 0.152939
R15051 gnd.n3176 gnd.n3175 0.152939
R15052 gnd.n3177 gnd.n3176 0.152939
R15053 gnd.n3177 gnd.n2054 0.152939
R15054 gnd.n3185 gnd.n2054 0.152939
R15055 gnd.n3186 gnd.n3185 0.152939
R15056 gnd.n3187 gnd.n3186 0.152939
R15057 gnd.n3187 gnd.n2048 0.152939
R15058 gnd.n3195 gnd.n2048 0.152939
R15059 gnd.n3196 gnd.n3195 0.152939
R15060 gnd.n3197 gnd.n3196 0.152939
R15061 gnd.n3197 gnd.n2042 0.152939
R15062 gnd.n3205 gnd.n2042 0.152939
R15063 gnd.n3206 gnd.n3205 0.152939
R15064 gnd.n3207 gnd.n3206 0.152939
R15065 gnd.n3207 gnd.n2036 0.152939
R15066 gnd.n3215 gnd.n2036 0.152939
R15067 gnd.n3216 gnd.n3215 0.152939
R15068 gnd.n3217 gnd.n3216 0.152939
R15069 gnd.n3217 gnd.n2030 0.152939
R15070 gnd.n3225 gnd.n2030 0.152939
R15071 gnd.n3226 gnd.n3225 0.152939
R15072 gnd.n3227 gnd.n3226 0.152939
R15073 gnd.n3227 gnd.n2024 0.152939
R15074 gnd.n3235 gnd.n2024 0.152939
R15075 gnd.n3236 gnd.n3235 0.152939
R15076 gnd.n3237 gnd.n3236 0.152939
R15077 gnd.n3237 gnd.n2018 0.152939
R15078 gnd.n3245 gnd.n2018 0.152939
R15079 gnd.n3246 gnd.n3245 0.152939
R15080 gnd.n3247 gnd.n3246 0.152939
R15081 gnd.n3247 gnd.n2012 0.152939
R15082 gnd.n3255 gnd.n2012 0.152939
R15083 gnd.n3256 gnd.n3255 0.152939
R15084 gnd.n3257 gnd.n3256 0.152939
R15085 gnd.n3257 gnd.n2006 0.152939
R15086 gnd.n3265 gnd.n2006 0.152939
R15087 gnd.n3266 gnd.n3265 0.152939
R15088 gnd.n3267 gnd.n3266 0.152939
R15089 gnd.n3267 gnd.n2000 0.152939
R15090 gnd.n3275 gnd.n2000 0.152939
R15091 gnd.n3276 gnd.n3275 0.152939
R15092 gnd.n3277 gnd.n3276 0.152939
R15093 gnd.n3277 gnd.n1994 0.152939
R15094 gnd.n3285 gnd.n1994 0.152939
R15095 gnd.n3286 gnd.n3285 0.152939
R15096 gnd.n3287 gnd.n3286 0.152939
R15097 gnd.n3287 gnd.n1988 0.152939
R15098 gnd.n3295 gnd.n1988 0.152939
R15099 gnd.n3296 gnd.n3295 0.152939
R15100 gnd.n3297 gnd.n3296 0.152939
R15101 gnd.n3297 gnd.n1982 0.152939
R15102 gnd.n3305 gnd.n1982 0.152939
R15103 gnd.n3306 gnd.n3305 0.152939
R15104 gnd.n3307 gnd.n3306 0.152939
R15105 gnd.n3307 gnd.n1976 0.152939
R15106 gnd.n3315 gnd.n1976 0.152939
R15107 gnd.n3316 gnd.n3315 0.152939
R15108 gnd.n3317 gnd.n3316 0.152939
R15109 gnd.n3318 gnd.n3317 0.152939
R15110 gnd.n5554 gnd.n5553 0.152939
R15111 gnd.n5561 gnd.n5553 0.152939
R15112 gnd.n5562 gnd.n5561 0.152939
R15113 gnd.n5563 gnd.n5562 0.152939
R15114 gnd.n5563 gnd.n5540 0.152939
R15115 gnd.n5582 gnd.n5540 0.152939
R15116 gnd.n5583 gnd.n5582 0.152939
R15117 gnd.n5584 gnd.n5583 0.152939
R15118 gnd.n5584 gnd.n5528 0.152939
R15119 gnd.n5603 gnd.n5528 0.152939
R15120 gnd.n5604 gnd.n5603 0.152939
R15121 gnd.n5605 gnd.n5604 0.152939
R15122 gnd.n5605 gnd.n5516 0.152939
R15123 gnd.n5624 gnd.n5516 0.152939
R15124 gnd.n5625 gnd.n5624 0.152939
R15125 gnd.n5635 gnd.n5625 0.152939
R15126 gnd.n5635 gnd.n5634 0.152939
R15127 gnd.n5634 gnd.n5633 0.152939
R15128 gnd.n5633 gnd.n5626 0.152939
R15129 gnd.n5629 gnd.n5626 0.152939
R15130 gnd.n5629 gnd.n5628 0.152939
R15131 gnd.n5628 gnd.n1215 0.152939
R15132 gnd.n6114 gnd.n1215 0.152939
R15133 gnd.n6115 gnd.n6114 0.152939
R15134 gnd.n6142 gnd.n6115 0.152939
R15135 gnd.n6142 gnd.n6141 0.152939
R15136 gnd.n6141 gnd.n6140 0.152939
R15137 gnd.n6140 gnd.n6116 0.152939
R15138 gnd.n6136 gnd.n6116 0.152939
R15139 gnd.n6136 gnd.n6135 0.152939
R15140 gnd.n6135 gnd.n6134 0.152939
R15141 gnd.n6134 gnd.n6122 0.152939
R15142 gnd.n6130 gnd.n6122 0.152939
R15143 gnd.n6130 gnd.n6129 0.152939
R15144 gnd.n6129 gnd.n6128 0.152939
R15145 gnd.n6128 gnd.n6125 0.152939
R15146 gnd.n6125 gnd.n6124 0.152939
R15147 gnd.n6124 gnd.n1096 0.152939
R15148 gnd.n6310 gnd.n1096 0.152939
R15149 gnd.n6311 gnd.n6310 0.152939
R15150 gnd.n6338 gnd.n6311 0.152939
R15151 gnd.n6338 gnd.n6337 0.152939
R15152 gnd.n6337 gnd.n6336 0.152939
R15153 gnd.n6336 gnd.n6312 0.152939
R15154 gnd.n6332 gnd.n6312 0.152939
R15155 gnd.n6332 gnd.n6331 0.152939
R15156 gnd.n6331 gnd.n6330 0.152939
R15157 gnd.n6330 gnd.n6316 0.152939
R15158 gnd.n6326 gnd.n6316 0.152939
R15159 gnd.n6326 gnd.n6325 0.152939
R15160 gnd.n6325 gnd.n6324 0.152939
R15161 gnd.n6324 gnd.n6320 0.152939
R15162 gnd.n6320 gnd.n968 0.152939
R15163 gnd.n6502 gnd.n968 0.152939
R15164 gnd.n6503 gnd.n6502 0.152939
R15165 gnd.n6504 gnd.n6503 0.152939
R15166 gnd.n6504 gnd.n965 0.152939
R15167 gnd.n6508 gnd.n965 0.152939
R15168 gnd.n6509 gnd.n6508 0.152939
R15169 gnd.n6515 gnd.n6509 0.152939
R15170 gnd.n6515 gnd.n6514 0.152939
R15171 gnd.n6514 gnd.n6513 0.152939
R15172 gnd.n6513 gnd.n6510 0.152939
R15173 gnd.n6510 gnd.n870 0.152939
R15174 gnd.n6738 gnd.n870 0.152939
R15175 gnd.n6739 gnd.n6738 0.152939
R15176 gnd.n6741 gnd.n6739 0.152939
R15177 gnd.n6741 gnd.n6740 0.152939
R15178 gnd.n6740 gnd.n845 0.152939
R15179 gnd.n6768 gnd.n845 0.152939
R15180 gnd.n6769 gnd.n6768 0.152939
R15181 gnd.n6771 gnd.n6769 0.152939
R15182 gnd.n6771 gnd.n6770 0.152939
R15183 gnd.n6770 gnd.n821 0.152939
R15184 gnd.n6798 gnd.n821 0.152939
R15185 gnd.n6799 gnd.n6798 0.152939
R15186 gnd.n6806 gnd.n6799 0.152939
R15187 gnd.n6806 gnd.n6805 0.152939
R15188 gnd.n6805 gnd.n6804 0.152939
R15189 gnd.n6804 gnd.n6800 0.152939
R15190 gnd.n6800 gnd.n759 0.152939
R15191 gnd.n6864 gnd.n759 0.152939
R15192 gnd.n5266 gnd.n1649 0.152939
R15193 gnd.n5267 gnd.n5266 0.152939
R15194 gnd.n5269 gnd.n5267 0.152939
R15195 gnd.n5269 gnd.n5268 0.152939
R15196 gnd.n5268 gnd.n1615 0.152939
R15197 gnd.n5302 gnd.n1615 0.152939
R15198 gnd.n5303 gnd.n5302 0.152939
R15199 gnd.n5305 gnd.n5303 0.152939
R15200 gnd.n5305 gnd.n5304 0.152939
R15201 gnd.n5304 gnd.n1586 0.152939
R15202 gnd.n5338 gnd.n1586 0.152939
R15203 gnd.n5339 gnd.n5338 0.152939
R15204 gnd.n5341 gnd.n5339 0.152939
R15205 gnd.n5341 gnd.n5340 0.152939
R15206 gnd.n5340 gnd.n1555 0.152939
R15207 gnd.n5380 gnd.n1555 0.152939
R15208 gnd.n5381 gnd.n5380 0.152939
R15209 gnd.n5383 gnd.n5381 0.152939
R15210 gnd.n5383 gnd.n5382 0.152939
R15211 gnd.n5382 gnd.n1520 0.152939
R15212 gnd.n5423 gnd.n1520 0.152939
R15213 gnd.n5424 gnd.n5423 0.152939
R15214 gnd.n5429 gnd.n5424 0.152939
R15215 gnd.n5429 gnd.n5428 0.152939
R15216 gnd.n5428 gnd.n5427 0.152939
R15217 gnd.n5427 gnd.n1450 0.152939
R15218 gnd.n5851 gnd.n1450 0.152939
R15219 gnd.n5851 gnd.n5850 0.152939
R15220 gnd.n5850 gnd.n5849 0.152939
R15221 gnd.n5849 gnd.n1451 0.152939
R15222 gnd.n5845 gnd.n1451 0.152939
R15223 gnd.n5833 gnd.n1478 0.152939
R15224 gnd.n5833 gnd.n5832 0.152939
R15225 gnd.n5832 gnd.n5831 0.152939
R15226 gnd.n5831 gnd.n1480 0.152939
R15227 gnd.n5827 gnd.n1480 0.152939
R15228 gnd.n5827 gnd.n5826 0.152939
R15229 gnd.n5679 gnd.n5484 0.152939
R15230 gnd.n5679 gnd.n5678 0.152939
R15231 gnd.n5678 gnd.n5677 0.152939
R15232 gnd.n5677 gnd.n5485 0.152939
R15233 gnd.n5673 gnd.n5485 0.152939
R15234 gnd.n5673 gnd.n5672 0.152939
R15235 gnd.n5672 gnd.n5671 0.152939
R15236 gnd.n5671 gnd.n5490 0.152939
R15237 gnd.n5667 gnd.n5490 0.152939
R15238 gnd.n5667 gnd.n5666 0.152939
R15239 gnd.n5666 gnd.n5665 0.152939
R15240 gnd.n5665 gnd.n5495 0.152939
R15241 gnd.n5661 gnd.n5495 0.152939
R15242 gnd.n5661 gnd.n5660 0.152939
R15243 gnd.n5660 gnd.n5659 0.152939
R15244 gnd.n5659 gnd.n5500 0.152939
R15245 gnd.n5655 gnd.n5500 0.152939
R15246 gnd.n5655 gnd.n1223 0.152939
R15247 gnd.n6103 gnd.n1223 0.152939
R15248 gnd.n6104 gnd.n6103 0.152939
R15249 gnd.n6106 gnd.n6104 0.152939
R15250 gnd.n6106 gnd.n6105 0.152939
R15251 gnd.n6105 gnd.n1181 0.152939
R15252 gnd.n6179 gnd.n1181 0.152939
R15253 gnd.n6180 gnd.n6179 0.152939
R15254 gnd.n6191 gnd.n6180 0.152939
R15255 gnd.n6191 gnd.n6190 0.152939
R15256 gnd.n6190 gnd.n6189 0.152939
R15257 gnd.n6189 gnd.n6181 0.152939
R15258 gnd.n6185 gnd.n6181 0.152939
R15259 gnd.n6185 gnd.n1132 0.152939
R15260 gnd.n6255 gnd.n1132 0.152939
R15261 gnd.n6256 gnd.n6255 0.152939
R15262 gnd.n6257 gnd.n6256 0.152939
R15263 gnd.n6257 gnd.n1104 0.152939
R15264 gnd.n6301 gnd.n1104 0.152939
R15265 gnd.n6302 gnd.n6301 0.152939
R15266 gnd.n6303 gnd.n6302 0.152939
R15267 gnd.n6303 gnd.n1073 0.152939
R15268 gnd.n6363 gnd.n1073 0.152939
R15269 gnd.n6364 gnd.n6363 0.152939
R15270 gnd.n6365 gnd.n6364 0.152939
R15271 gnd.n6365 gnd.n1046 0.152939
R15272 gnd.n6400 gnd.n1046 0.152939
R15273 gnd.n6401 gnd.n6400 0.152939
R15274 gnd.n6402 gnd.n6401 0.152939
R15275 gnd.n6402 gnd.n1017 0.152939
R15276 gnd.n6436 gnd.n1017 0.152939
R15277 gnd.n6437 gnd.n6436 0.152939
R15278 gnd.n6438 gnd.n6437 0.152939
R15279 gnd.n6438 gnd.n978 0.152939
R15280 gnd.n6493 gnd.n978 0.152939
R15281 gnd.n6494 gnd.n6493 0.152939
R15282 gnd.n6496 gnd.n6494 0.152939
R15283 gnd.n6496 gnd.n6495 0.152939
R15284 gnd.n6495 gnd.n958 0.152939
R15285 gnd.n6528 gnd.n958 0.152939
R15286 gnd.n6528 gnd.n6527 0.152939
R15287 gnd.n6527 gnd.n6526 0.152939
R15288 gnd.n6526 gnd.n959 0.152939
R15289 gnd.n6522 gnd.n959 0.152939
R15290 gnd.n6522 gnd.n880 0.152939
R15291 gnd.n6729 gnd.n880 0.152939
R15292 gnd.n6730 gnd.n6729 0.152939
R15293 gnd.n6732 gnd.n6730 0.152939
R15294 gnd.n6732 gnd.n6731 0.152939
R15295 gnd.n6731 gnd.n855 0.152939
R15296 gnd.n6759 gnd.n855 0.152939
R15297 gnd.n6760 gnd.n6759 0.152939
R15298 gnd.n6762 gnd.n6760 0.152939
R15299 gnd.n6762 gnd.n6761 0.152939
R15300 gnd.n6761 gnd.n830 0.152939
R15301 gnd.n6789 gnd.n830 0.152939
R15302 gnd.n6790 gnd.n6789 0.152939
R15303 gnd.n6792 gnd.n6790 0.152939
R15304 gnd.n6792 gnd.n6791 0.152939
R15305 gnd.n6791 gnd.n806 0.152939
R15306 gnd.n6825 gnd.n806 0.152939
R15307 gnd.n6826 gnd.n6825 0.152939
R15308 gnd.n6827 gnd.n6826 0.152939
R15309 gnd.n6827 gnd.n768 0.152939
R15310 gnd.n6858 gnd.n768 0.152939
R15311 gnd.n6857 gnd.n769 0.152939
R15312 gnd.n6853 gnd.n769 0.152939
R15313 gnd.n6853 gnd.n6852 0.152939
R15314 gnd.n6852 gnd.n6851 0.152939
R15315 gnd.n6851 gnd.n773 0.152939
R15316 gnd.n773 gnd.n695 0.152939
R15317 gnd.n6867 gnd.n558 0.152939
R15318 gnd.n7081 gnd.n558 0.152939
R15319 gnd.n7082 gnd.n7081 0.152939
R15320 gnd.n7084 gnd.n7082 0.152939
R15321 gnd.n7084 gnd.n7083 0.152939
R15322 gnd.n7083 gnd.n518 0.152939
R15323 gnd.n7131 gnd.n518 0.152939
R15324 gnd.n7132 gnd.n7131 0.152939
R15325 gnd.n7133 gnd.n7132 0.152939
R15326 gnd.n7133 gnd.n515 0.152939
R15327 gnd.n7138 gnd.n515 0.152939
R15328 gnd.n7139 gnd.n7138 0.152939
R15329 gnd.n7141 gnd.n7139 0.152939
R15330 gnd.n7141 gnd.n7140 0.152939
R15331 gnd.n7140 gnd.n453 0.152939
R15332 gnd.n7201 gnd.n453 0.152939
R15333 gnd.n7202 gnd.n7201 0.152939
R15334 gnd.n7213 gnd.n7202 0.152939
R15335 gnd.n7213 gnd.n7212 0.152939
R15336 gnd.n7212 gnd.n7211 0.152939
R15337 gnd.n7211 gnd.n7203 0.152939
R15338 gnd.n7207 gnd.n7203 0.152939
R15339 gnd.n7207 gnd.n7206 0.152939
R15340 gnd.n7206 gnd.n399 0.152939
R15341 gnd.n7288 gnd.n399 0.152939
R15342 gnd.n7289 gnd.n7288 0.152939
R15343 gnd.n7296 gnd.n7289 0.152939
R15344 gnd.n7296 gnd.n7295 0.152939
R15345 gnd.n7295 gnd.n7294 0.152939
R15346 gnd.n7294 gnd.n7290 0.152939
R15347 gnd.n7290 gnd.n95 0.152939
R15348 gnd.n1919 gnd.n1626 0.14989
R15349 gnd.n7247 gnd.n110 0.14989
R15350 gnd.n7759 gnd.n7758 0.145814
R15351 gnd.n5234 gnd.n5233 0.145814
R15352 gnd.n5234 gnd.n1649 0.145814
R15353 gnd.n7759 gnd.n95 0.145814
R15354 gnd.n5826 gnd.n1421 0.128549
R15355 gnd.n6925 gnd.n695 0.128549
R15356 gnd.n4123 gnd.n4122 0.0767195
R15357 gnd.n4122 gnd.n4121 0.0767195
R15358 gnd.n5971 gnd.n1421 0.063
R15359 gnd.n6926 gnd.n6925 0.063
R15360 gnd.n4690 gnd.n1860 0.0477147
R15361 gnd.n3886 gnd.n3774 0.0442063
R15362 gnd.n3887 gnd.n3886 0.0442063
R15363 gnd.n3888 gnd.n3887 0.0442063
R15364 gnd.n3888 gnd.n3763 0.0442063
R15365 gnd.n3902 gnd.n3763 0.0442063
R15366 gnd.n3903 gnd.n3902 0.0442063
R15367 gnd.n3904 gnd.n3903 0.0442063
R15368 gnd.n3904 gnd.n3750 0.0442063
R15369 gnd.n3948 gnd.n3750 0.0442063
R15370 gnd.n3949 gnd.n3948 0.0442063
R15371 gnd.n6926 gnd.n575 0.0416005
R15372 gnd.n7540 gnd.n7539 0.0416005
R15373 gnd.n5034 gnd.n5033 0.0416005
R15374 gnd.n5971 gnd.n5970 0.0416005
R15375 gnd.n3951 gnd.n3684 0.0344674
R15376 gnd.n7064 gnd.n575 0.0344674
R15377 gnd.n7064 gnd.n581 0.0344674
R15378 gnd.n581 gnd.n580 0.0344674
R15379 gnd.n580 gnd.n552 0.0344674
R15380 gnd.n552 gnd.n538 0.0344674
R15381 gnd.n539 gnd.n538 0.0344674
R15382 gnd.n540 gnd.n539 0.0344674
R15383 gnd.n541 gnd.n540 0.0344674
R15384 gnd.n7091 gnd.n541 0.0344674
R15385 gnd.n7091 gnd.n503 0.0344674
R15386 gnd.n504 gnd.n503 0.0344674
R15387 gnd.n7148 gnd.n504 0.0344674
R15388 gnd.n7148 gnd.n505 0.0344674
R15389 gnd.n505 gnd.n473 0.0344674
R15390 gnd.n474 gnd.n473 0.0344674
R15391 gnd.n475 gnd.n474 0.0344674
R15392 gnd.n476 gnd.n475 0.0344674
R15393 gnd.n476 gnd.n448 0.0344674
R15394 gnd.n448 gnd.n446 0.0344674
R15395 gnd.n7222 gnd.n446 0.0344674
R15396 gnd.n7223 gnd.n7222 0.0344674
R15397 gnd.n7223 gnd.n421 0.0344674
R15398 gnd.n421 gnd.n418 0.0344674
R15399 gnd.n419 gnd.n418 0.0344674
R15400 gnd.n7266 gnd.n419 0.0344674
R15401 gnd.n7267 gnd.n7266 0.0344674
R15402 gnd.n7267 gnd.n392 0.0344674
R15403 gnd.n7303 gnd.n392 0.0344674
R15404 gnd.n7303 gnd.n375 0.0344674
R15405 gnd.n7326 gnd.n375 0.0344674
R15406 gnd.n7327 gnd.n7326 0.0344674
R15407 gnd.n7327 gnd.n364 0.0344674
R15408 gnd.n7340 gnd.n364 0.0344674
R15409 gnd.n7340 gnd.n354 0.0344674
R15410 gnd.n7356 gnd.n354 0.0344674
R15411 gnd.n7357 gnd.n7356 0.0344674
R15412 gnd.n7357 gnd.n124 0.0344674
R15413 gnd.n125 gnd.n124 0.0344674
R15414 gnd.n126 gnd.n125 0.0344674
R15415 gnd.n7494 gnd.n126 0.0344674
R15416 gnd.n7494 gnd.n141 0.0344674
R15417 gnd.n142 gnd.n141 0.0344674
R15418 gnd.n143 gnd.n142 0.0344674
R15419 gnd.n7501 gnd.n143 0.0344674
R15420 gnd.n7501 gnd.n161 0.0344674
R15421 gnd.n162 gnd.n161 0.0344674
R15422 gnd.n163 gnd.n162 0.0344674
R15423 gnd.n7508 gnd.n163 0.0344674
R15424 gnd.n7508 gnd.n179 0.0344674
R15425 gnd.n180 gnd.n179 0.0344674
R15426 gnd.n181 gnd.n180 0.0344674
R15427 gnd.n7515 gnd.n181 0.0344674
R15428 gnd.n7515 gnd.n199 0.0344674
R15429 gnd.n200 gnd.n199 0.0344674
R15430 gnd.n201 gnd.n200 0.0344674
R15431 gnd.n7522 gnd.n201 0.0344674
R15432 gnd.n7522 gnd.n217 0.0344674
R15433 gnd.n218 gnd.n217 0.0344674
R15434 gnd.n219 gnd.n218 0.0344674
R15435 gnd.n7529 gnd.n219 0.0344674
R15436 gnd.n7529 gnd.n237 0.0344674
R15437 gnd.n238 gnd.n237 0.0344674
R15438 gnd.n239 gnd.n238 0.0344674
R15439 gnd.n7539 gnd.n239 0.0344674
R15440 gnd.n5039 gnd.n5034 0.0344674
R15441 gnd.n5039 gnd.n5036 0.0344674
R15442 gnd.n5036 gnd.n1811 0.0344674
R15443 gnd.n1811 gnd.n1809 0.0344674
R15444 gnd.n5057 gnd.n1809 0.0344674
R15445 gnd.n5058 gnd.n5057 0.0344674
R15446 gnd.n5058 gnd.n1793 0.0344674
R15447 gnd.n1793 gnd.n1790 0.0344674
R15448 gnd.n1791 gnd.n1790 0.0344674
R15449 gnd.n5079 gnd.n1791 0.0344674
R15450 gnd.n5080 gnd.n5079 0.0344674
R15451 gnd.n5080 gnd.n1767 0.0344674
R15452 gnd.n1767 gnd.n1764 0.0344674
R15453 gnd.n1765 gnd.n1764 0.0344674
R15454 gnd.n5114 gnd.n1765 0.0344674
R15455 gnd.n5115 gnd.n5114 0.0344674
R15456 gnd.n5115 gnd.n1742 0.0344674
R15457 gnd.n1742 gnd.n1739 0.0344674
R15458 gnd.n1740 gnd.n1739 0.0344674
R15459 gnd.n5149 gnd.n1740 0.0344674
R15460 gnd.n5150 gnd.n5149 0.0344674
R15461 gnd.n5150 gnd.n1717 0.0344674
R15462 gnd.n1717 gnd.n1712 0.0344674
R15463 gnd.n1713 gnd.n1712 0.0344674
R15464 gnd.n1714 gnd.n1713 0.0344674
R15465 gnd.n5188 gnd.n1714 0.0344674
R15466 gnd.n5188 gnd.n1715 0.0344674
R15467 gnd.n1715 gnd.n1682 0.0344674
R15468 gnd.n5225 gnd.n1682 0.0344674
R15469 gnd.n5225 gnd.n1665 0.0344674
R15470 gnd.n5245 gnd.n1665 0.0344674
R15471 gnd.n5246 gnd.n5245 0.0344674
R15472 gnd.n5246 gnd.n1659 0.0344674
R15473 gnd.n5254 gnd.n1659 0.0344674
R15474 gnd.n5255 gnd.n5254 0.0344674
R15475 gnd.n5255 gnd.n1644 0.0344674
R15476 gnd.n1644 gnd.n1641 0.0344674
R15477 gnd.n1642 gnd.n1641 0.0344674
R15478 gnd.n5280 gnd.n1642 0.0344674
R15479 gnd.n5281 gnd.n5280 0.0344674
R15480 gnd.n5281 gnd.n1609 0.0344674
R15481 gnd.n1609 gnd.n1606 0.0344674
R15482 gnd.n1607 gnd.n1606 0.0344674
R15483 gnd.n5316 gnd.n1607 0.0344674
R15484 gnd.n5317 gnd.n5316 0.0344674
R15485 gnd.n5317 gnd.n1580 0.0344674
R15486 gnd.n1580 gnd.n1575 0.0344674
R15487 gnd.n1576 gnd.n1575 0.0344674
R15488 gnd.n1577 gnd.n1576 0.0344674
R15489 gnd.n5360 gnd.n1577 0.0344674
R15490 gnd.n5360 gnd.n1578 0.0344674
R15491 gnd.n1578 gnd.n1539 0.0344674
R15492 gnd.n1540 gnd.n1539 0.0344674
R15493 gnd.n1541 gnd.n1540 0.0344674
R15494 gnd.n1542 gnd.n1541 0.0344674
R15495 gnd.n1542 gnd.n1514 0.0344674
R15496 gnd.n1514 gnd.n1512 0.0344674
R15497 gnd.n5438 gnd.n1512 0.0344674
R15498 gnd.n5439 gnd.n5438 0.0344674
R15499 gnd.n5439 gnd.n1443 0.0344674
R15500 gnd.n5858 gnd.n1443 0.0344674
R15501 gnd.n5859 gnd.n5858 0.0344674
R15502 gnd.n5859 gnd.n1422 0.0344674
R15503 gnd.n5970 gnd.n1422 0.0344674
R15504 gnd.n5823 gnd.n5822 0.0344674
R15505 gnd.n6924 gnd.n696 0.0344674
R15506 gnd.n5844 gnd.n5843 0.029712
R15507 gnd.n6869 gnd.n6868 0.029712
R15508 gnd.n3971 gnd.n3970 0.0269946
R15509 gnd.n3973 gnd.n3972 0.0269946
R15510 gnd.n3679 gnd.n3677 0.0269946
R15511 gnd.n3983 gnd.n3981 0.0269946
R15512 gnd.n3982 gnd.n3658 0.0269946
R15513 gnd.n4002 gnd.n4001 0.0269946
R15514 gnd.n4004 gnd.n4003 0.0269946
R15515 gnd.n3653 gnd.n3652 0.0269946
R15516 gnd.n4014 gnd.n3648 0.0269946
R15517 gnd.n4013 gnd.n3650 0.0269946
R15518 gnd.n3649 gnd.n3631 0.0269946
R15519 gnd.n4034 gnd.n3632 0.0269946
R15520 gnd.n4033 gnd.n3633 0.0269946
R15521 gnd.n4067 gnd.n3608 0.0269946
R15522 gnd.n4069 gnd.n4068 0.0269946
R15523 gnd.n4070 gnd.n3555 0.0269946
R15524 gnd.n3603 gnd.n3556 0.0269946
R15525 gnd.n3605 gnd.n3557 0.0269946
R15526 gnd.n4080 gnd.n4079 0.0269946
R15527 gnd.n4082 gnd.n4081 0.0269946
R15528 gnd.n4083 gnd.n3577 0.0269946
R15529 gnd.n4085 gnd.n3578 0.0269946
R15530 gnd.n4088 gnd.n3579 0.0269946
R15531 gnd.n4091 gnd.n4090 0.0269946
R15532 gnd.n4093 gnd.n4092 0.0269946
R15533 gnd.n4158 gnd.n3446 0.0269946
R15534 gnd.n4160 gnd.n4159 0.0269946
R15535 gnd.n4169 gnd.n3439 0.0269946
R15536 gnd.n4171 gnd.n4170 0.0269946
R15537 gnd.n4172 gnd.n3437 0.0269946
R15538 gnd.n4179 gnd.n4175 0.0269946
R15539 gnd.n4178 gnd.n4177 0.0269946
R15540 gnd.n4176 gnd.n3416 0.0269946
R15541 gnd.n4201 gnd.n3417 0.0269946
R15542 gnd.n4200 gnd.n3418 0.0269946
R15543 gnd.n4243 gnd.n3391 0.0269946
R15544 gnd.n4245 gnd.n4244 0.0269946
R15545 gnd.n4254 gnd.n3384 0.0269946
R15546 gnd.n4256 gnd.n4255 0.0269946
R15547 gnd.n4257 gnd.n3382 0.0269946
R15548 gnd.n4264 gnd.n4260 0.0269946
R15549 gnd.n4263 gnd.n4262 0.0269946
R15550 gnd.n4261 gnd.n3361 0.0269946
R15551 gnd.n4286 gnd.n3362 0.0269946
R15552 gnd.n4285 gnd.n3363 0.0269946
R15553 gnd.n4332 gnd.n3337 0.0269946
R15554 gnd.n4334 gnd.n4333 0.0269946
R15555 gnd.n4343 gnd.n3330 0.0269946
R15556 gnd.n4602 gnd.n3328 0.0269946
R15557 gnd.n4607 gnd.n4605 0.0269946
R15558 gnd.n4606 gnd.n1896 0.0269946
R15559 gnd.n4632 gnd.n4631 0.0269946
R15560 gnd.n5821 gnd.n1487 0.0225788
R15561 gnd.n5818 gnd.n5817 0.0225788
R15562 gnd.n5814 gnd.n5703 0.0225788
R15563 gnd.n5813 gnd.n5710 0.0225788
R15564 gnd.n5810 gnd.n5809 0.0225788
R15565 gnd.n5806 gnd.n5717 0.0225788
R15566 gnd.n5805 gnd.n5723 0.0225788
R15567 gnd.n5802 gnd.n5801 0.0225788
R15568 gnd.n5798 gnd.n5729 0.0225788
R15569 gnd.n5797 gnd.n5733 0.0225788
R15570 gnd.n5794 gnd.n5793 0.0225788
R15571 gnd.n5790 gnd.n5740 0.0225788
R15572 gnd.n5789 gnd.n5746 0.0225788
R15573 gnd.n5786 gnd.n5785 0.0225788
R15574 gnd.n5782 gnd.n5752 0.0225788
R15575 gnd.n5781 gnd.n5756 0.0225788
R15576 gnd.n5778 gnd.n5777 0.0225788
R15577 gnd.n5770 gnd.n5769 0.0225788
R15578 gnd.n5843 gnd.n1456 0.0225788
R15579 gnd.n6920 gnd.n702 0.0225788
R15580 gnd.n6919 gnd.n703 0.0225788
R15581 gnd.n6916 gnd.n6915 0.0225788
R15582 gnd.n6912 gnd.n708 0.0225788
R15583 gnd.n6911 gnd.n712 0.0225788
R15584 gnd.n6908 gnd.n6907 0.0225788
R15585 gnd.n6904 gnd.n718 0.0225788
R15586 gnd.n6903 gnd.n722 0.0225788
R15587 gnd.n6900 gnd.n6899 0.0225788
R15588 gnd.n6896 gnd.n726 0.0225788
R15589 gnd.n6895 gnd.n730 0.0225788
R15590 gnd.n6892 gnd.n6891 0.0225788
R15591 gnd.n6888 gnd.n736 0.0225788
R15592 gnd.n6887 gnd.n740 0.0225788
R15593 gnd.n6884 gnd.n6883 0.0225788
R15594 gnd.n6880 gnd.n744 0.0225788
R15595 gnd.n6879 gnd.n750 0.0225788
R15596 gnd.n6873 gnd.n6872 0.0225788
R15597 gnd.n6869 gnd.n754 0.0225788
R15598 gnd.n6868 gnd.n6865 0.0218415
R15599 gnd.n5844 gnd.n1455 0.0218415
R15600 gnd.n3951 gnd.n3950 0.0202011
R15601 gnd.n3950 gnd.n3949 0.0148637
R15602 gnd.n4600 gnd.n4344 0.0144266
R15603 gnd.n4601 gnd.n4600 0.0130679
R15604 gnd.n5822 gnd.n5821 0.0123886
R15605 gnd.n5818 gnd.n1487 0.0123886
R15606 gnd.n5817 gnd.n5703 0.0123886
R15607 gnd.n5814 gnd.n5813 0.0123886
R15608 gnd.n5810 gnd.n5710 0.0123886
R15609 gnd.n5809 gnd.n5717 0.0123886
R15610 gnd.n5806 gnd.n5805 0.0123886
R15611 gnd.n5802 gnd.n5723 0.0123886
R15612 gnd.n5801 gnd.n5729 0.0123886
R15613 gnd.n5798 gnd.n5797 0.0123886
R15614 gnd.n5794 gnd.n5733 0.0123886
R15615 gnd.n5793 gnd.n5740 0.0123886
R15616 gnd.n5790 gnd.n5789 0.0123886
R15617 gnd.n5786 gnd.n5746 0.0123886
R15618 gnd.n5785 gnd.n5752 0.0123886
R15619 gnd.n5782 gnd.n5781 0.0123886
R15620 gnd.n5778 gnd.n5756 0.0123886
R15621 gnd.n5777 gnd.n5770 0.0123886
R15622 gnd.n5769 gnd.n1456 0.0123886
R15623 gnd.n702 gnd.n696 0.0123886
R15624 gnd.n6920 gnd.n6919 0.0123886
R15625 gnd.n6916 gnd.n703 0.0123886
R15626 gnd.n6915 gnd.n708 0.0123886
R15627 gnd.n6912 gnd.n6911 0.0123886
R15628 gnd.n6908 gnd.n712 0.0123886
R15629 gnd.n6907 gnd.n718 0.0123886
R15630 gnd.n6904 gnd.n6903 0.0123886
R15631 gnd.n6900 gnd.n722 0.0123886
R15632 gnd.n6899 gnd.n726 0.0123886
R15633 gnd.n6896 gnd.n6895 0.0123886
R15634 gnd.n6892 gnd.n730 0.0123886
R15635 gnd.n6891 gnd.n736 0.0123886
R15636 gnd.n6888 gnd.n6887 0.0123886
R15637 gnd.n6884 gnd.n740 0.0123886
R15638 gnd.n6883 gnd.n744 0.0123886
R15639 gnd.n6880 gnd.n6879 0.0123886
R15640 gnd.n6873 gnd.n750 0.0123886
R15641 gnd.n6872 gnd.n754 0.0123886
R15642 gnd.n3970 gnd.n3684 0.00797283
R15643 gnd.n3972 gnd.n3971 0.00797283
R15644 gnd.n3973 gnd.n3679 0.00797283
R15645 gnd.n3981 gnd.n3677 0.00797283
R15646 gnd.n3983 gnd.n3982 0.00797283
R15647 gnd.n4001 gnd.n3658 0.00797283
R15648 gnd.n4003 gnd.n4002 0.00797283
R15649 gnd.n4004 gnd.n3653 0.00797283
R15650 gnd.n3652 gnd.n3648 0.00797283
R15651 gnd.n4014 gnd.n4013 0.00797283
R15652 gnd.n3650 gnd.n3649 0.00797283
R15653 gnd.n3632 gnd.n3631 0.00797283
R15654 gnd.n4034 gnd.n4033 0.00797283
R15655 gnd.n3633 gnd.n3608 0.00797283
R15656 gnd.n4068 gnd.n4067 0.00797283
R15657 gnd.n4070 gnd.n4069 0.00797283
R15658 gnd.n3603 gnd.n3555 0.00797283
R15659 gnd.n3605 gnd.n3556 0.00797283
R15660 gnd.n4079 gnd.n3557 0.00797283
R15661 gnd.n4081 gnd.n4080 0.00797283
R15662 gnd.n4083 gnd.n4082 0.00797283
R15663 gnd.n4085 gnd.n3577 0.00797283
R15664 gnd.n4088 gnd.n3578 0.00797283
R15665 gnd.n4090 gnd.n3579 0.00797283
R15666 gnd.n4093 gnd.n4091 0.00797283
R15667 gnd.n4092 gnd.n3446 0.00797283
R15668 gnd.n4160 gnd.n4158 0.00797283
R15669 gnd.n4159 gnd.n3439 0.00797283
R15670 gnd.n4170 gnd.n4169 0.00797283
R15671 gnd.n4172 gnd.n4171 0.00797283
R15672 gnd.n4175 gnd.n3437 0.00797283
R15673 gnd.n4179 gnd.n4178 0.00797283
R15674 gnd.n4177 gnd.n4176 0.00797283
R15675 gnd.n3417 gnd.n3416 0.00797283
R15676 gnd.n4201 gnd.n4200 0.00797283
R15677 gnd.n3418 gnd.n3391 0.00797283
R15678 gnd.n4245 gnd.n4243 0.00797283
R15679 gnd.n4244 gnd.n3384 0.00797283
R15680 gnd.n4255 gnd.n4254 0.00797283
R15681 gnd.n4257 gnd.n4256 0.00797283
R15682 gnd.n4260 gnd.n3382 0.00797283
R15683 gnd.n4264 gnd.n4263 0.00797283
R15684 gnd.n4262 gnd.n4261 0.00797283
R15685 gnd.n3362 gnd.n3361 0.00797283
R15686 gnd.n4286 gnd.n4285 0.00797283
R15687 gnd.n3363 gnd.n3337 0.00797283
R15688 gnd.n4334 gnd.n4332 0.00797283
R15689 gnd.n4333 gnd.n3330 0.00797283
R15690 gnd.n4344 gnd.n4343 0.00797283
R15691 gnd.n4602 gnd.n4601 0.00797283
R15692 gnd.n4605 gnd.n3328 0.00797283
R15693 gnd.n4607 gnd.n4606 0.00797283
R15694 gnd.n4631 gnd.n1896 0.00797283
R15695 gnd.n4632 gnd.n1860 0.00797283
R15696 gnd.n5823 gnd.n1421 0.00593478
R15697 gnd.n6925 gnd.n6924 0.00593478
R15698 CSoutput.n19 CSoutput.t258 184.661
R15699 CSoutput.n78 CSoutput.n77 165.8
R15700 CSoutput.n76 CSoutput.n0 165.8
R15701 CSoutput.n75 CSoutput.n74 165.8
R15702 CSoutput.n73 CSoutput.n72 165.8
R15703 CSoutput.n71 CSoutput.n2 165.8
R15704 CSoutput.n69 CSoutput.n68 165.8
R15705 CSoutput.n67 CSoutput.n3 165.8
R15706 CSoutput.n66 CSoutput.n65 165.8
R15707 CSoutput.n63 CSoutput.n4 165.8
R15708 CSoutput.n61 CSoutput.n60 165.8
R15709 CSoutput.n59 CSoutput.n5 165.8
R15710 CSoutput.n58 CSoutput.n57 165.8
R15711 CSoutput.n55 CSoutput.n6 165.8
R15712 CSoutput.n54 CSoutput.n53 165.8
R15713 CSoutput.n52 CSoutput.n51 165.8
R15714 CSoutput.n50 CSoutput.n8 165.8
R15715 CSoutput.n48 CSoutput.n47 165.8
R15716 CSoutput.n46 CSoutput.n9 165.8
R15717 CSoutput.n45 CSoutput.n44 165.8
R15718 CSoutput.n42 CSoutput.n10 165.8
R15719 CSoutput.n41 CSoutput.n40 165.8
R15720 CSoutput.n39 CSoutput.n38 165.8
R15721 CSoutput.n37 CSoutput.n12 165.8
R15722 CSoutput.n35 CSoutput.n34 165.8
R15723 CSoutput.n33 CSoutput.n13 165.8
R15724 CSoutput.n32 CSoutput.n31 165.8
R15725 CSoutput.n29 CSoutput.n14 165.8
R15726 CSoutput.n28 CSoutput.n27 165.8
R15727 CSoutput.n26 CSoutput.n25 165.8
R15728 CSoutput.n24 CSoutput.n16 165.8
R15729 CSoutput.n22 CSoutput.n21 165.8
R15730 CSoutput.n20 CSoutput.n17 165.8
R15731 CSoutput.n77 CSoutput.t259 162.194
R15732 CSoutput.n18 CSoutput.t248 120.501
R15733 CSoutput.n23 CSoutput.t250 120.501
R15734 CSoutput.n15 CSoutput.t242 120.501
R15735 CSoutput.n30 CSoutput.t254 120.501
R15736 CSoutput.n36 CSoutput.t251 120.501
R15737 CSoutput.n11 CSoutput.t245 120.501
R15738 CSoutput.n43 CSoutput.t241 120.501
R15739 CSoutput.n49 CSoutput.t252 120.501
R15740 CSoutput.n7 CSoutput.t253 120.501
R15741 CSoutput.n56 CSoutput.t244 120.501
R15742 CSoutput.n62 CSoutput.t261 120.501
R15743 CSoutput.n64 CSoutput.t257 120.501
R15744 CSoutput.n70 CSoutput.t247 120.501
R15745 CSoutput.n1 CSoutput.t249 120.501
R15746 CSoutput.n330 CSoutput.n328 103.469
R15747 CSoutput.n310 CSoutput.n308 103.469
R15748 CSoutput.n291 CSoutput.n289 103.469
R15749 CSoutput.n120 CSoutput.n118 103.469
R15750 CSoutput.n100 CSoutput.n98 103.469
R15751 CSoutput.n81 CSoutput.n79 103.469
R15752 CSoutput.n344 CSoutput.n343 103.111
R15753 CSoutput.n342 CSoutput.n341 103.111
R15754 CSoutput.n340 CSoutput.n339 103.111
R15755 CSoutput.n338 CSoutput.n337 103.111
R15756 CSoutput.n336 CSoutput.n335 103.111
R15757 CSoutput.n334 CSoutput.n333 103.111
R15758 CSoutput.n332 CSoutput.n331 103.111
R15759 CSoutput.n330 CSoutput.n329 103.111
R15760 CSoutput.n326 CSoutput.n325 103.111
R15761 CSoutput.n324 CSoutput.n323 103.111
R15762 CSoutput.n322 CSoutput.n321 103.111
R15763 CSoutput.n320 CSoutput.n319 103.111
R15764 CSoutput.n318 CSoutput.n317 103.111
R15765 CSoutput.n316 CSoutput.n315 103.111
R15766 CSoutput.n314 CSoutput.n313 103.111
R15767 CSoutput.n312 CSoutput.n311 103.111
R15768 CSoutput.n310 CSoutput.n309 103.111
R15769 CSoutput.n307 CSoutput.n306 103.111
R15770 CSoutput.n305 CSoutput.n304 103.111
R15771 CSoutput.n303 CSoutput.n302 103.111
R15772 CSoutput.n301 CSoutput.n300 103.111
R15773 CSoutput.n299 CSoutput.n298 103.111
R15774 CSoutput.n297 CSoutput.n296 103.111
R15775 CSoutput.n295 CSoutput.n294 103.111
R15776 CSoutput.n293 CSoutput.n292 103.111
R15777 CSoutput.n291 CSoutput.n290 103.111
R15778 CSoutput.n120 CSoutput.n119 103.111
R15779 CSoutput.n122 CSoutput.n121 103.111
R15780 CSoutput.n124 CSoutput.n123 103.111
R15781 CSoutput.n126 CSoutput.n125 103.111
R15782 CSoutput.n128 CSoutput.n127 103.111
R15783 CSoutput.n130 CSoutput.n129 103.111
R15784 CSoutput.n132 CSoutput.n131 103.111
R15785 CSoutput.n134 CSoutput.n133 103.111
R15786 CSoutput.n136 CSoutput.n135 103.111
R15787 CSoutput.n100 CSoutput.n99 103.111
R15788 CSoutput.n102 CSoutput.n101 103.111
R15789 CSoutput.n104 CSoutput.n103 103.111
R15790 CSoutput.n106 CSoutput.n105 103.111
R15791 CSoutput.n108 CSoutput.n107 103.111
R15792 CSoutput.n110 CSoutput.n109 103.111
R15793 CSoutput.n112 CSoutput.n111 103.111
R15794 CSoutput.n114 CSoutput.n113 103.111
R15795 CSoutput.n116 CSoutput.n115 103.111
R15796 CSoutput.n81 CSoutput.n80 103.111
R15797 CSoutput.n83 CSoutput.n82 103.111
R15798 CSoutput.n85 CSoutput.n84 103.111
R15799 CSoutput.n87 CSoutput.n86 103.111
R15800 CSoutput.n89 CSoutput.n88 103.111
R15801 CSoutput.n91 CSoutput.n90 103.111
R15802 CSoutput.n93 CSoutput.n92 103.111
R15803 CSoutput.n95 CSoutput.n94 103.111
R15804 CSoutput.n97 CSoutput.n96 103.111
R15805 CSoutput.n346 CSoutput.n345 103.111
R15806 CSoutput.n390 CSoutput.n388 81.5057
R15807 CSoutput.n370 CSoutput.n368 81.5057
R15808 CSoutput.n351 CSoutput.n349 81.5057
R15809 CSoutput.n450 CSoutput.n448 81.5057
R15810 CSoutput.n430 CSoutput.n428 81.5057
R15811 CSoutput.n411 CSoutput.n409 81.5057
R15812 CSoutput.n406 CSoutput.n405 80.9324
R15813 CSoutput.n404 CSoutput.n403 80.9324
R15814 CSoutput.n402 CSoutput.n401 80.9324
R15815 CSoutput.n400 CSoutput.n399 80.9324
R15816 CSoutput.n398 CSoutput.n397 80.9324
R15817 CSoutput.n396 CSoutput.n395 80.9324
R15818 CSoutput.n394 CSoutput.n393 80.9324
R15819 CSoutput.n392 CSoutput.n391 80.9324
R15820 CSoutput.n390 CSoutput.n389 80.9324
R15821 CSoutput.n386 CSoutput.n385 80.9324
R15822 CSoutput.n384 CSoutput.n383 80.9324
R15823 CSoutput.n382 CSoutput.n381 80.9324
R15824 CSoutput.n380 CSoutput.n379 80.9324
R15825 CSoutput.n378 CSoutput.n377 80.9324
R15826 CSoutput.n376 CSoutput.n375 80.9324
R15827 CSoutput.n374 CSoutput.n373 80.9324
R15828 CSoutput.n372 CSoutput.n371 80.9324
R15829 CSoutput.n370 CSoutput.n369 80.9324
R15830 CSoutput.n367 CSoutput.n366 80.9324
R15831 CSoutput.n365 CSoutput.n364 80.9324
R15832 CSoutput.n363 CSoutput.n362 80.9324
R15833 CSoutput.n361 CSoutput.n360 80.9324
R15834 CSoutput.n359 CSoutput.n358 80.9324
R15835 CSoutput.n357 CSoutput.n356 80.9324
R15836 CSoutput.n355 CSoutput.n354 80.9324
R15837 CSoutput.n353 CSoutput.n352 80.9324
R15838 CSoutput.n351 CSoutput.n350 80.9324
R15839 CSoutput.n450 CSoutput.n449 80.9324
R15840 CSoutput.n452 CSoutput.n451 80.9324
R15841 CSoutput.n454 CSoutput.n453 80.9324
R15842 CSoutput.n456 CSoutput.n455 80.9324
R15843 CSoutput.n458 CSoutput.n457 80.9324
R15844 CSoutput.n460 CSoutput.n459 80.9324
R15845 CSoutput.n462 CSoutput.n461 80.9324
R15846 CSoutput.n464 CSoutput.n463 80.9324
R15847 CSoutput.n466 CSoutput.n465 80.9324
R15848 CSoutput.n430 CSoutput.n429 80.9324
R15849 CSoutput.n432 CSoutput.n431 80.9324
R15850 CSoutput.n434 CSoutput.n433 80.9324
R15851 CSoutput.n436 CSoutput.n435 80.9324
R15852 CSoutput.n438 CSoutput.n437 80.9324
R15853 CSoutput.n440 CSoutput.n439 80.9324
R15854 CSoutput.n442 CSoutput.n441 80.9324
R15855 CSoutput.n444 CSoutput.n443 80.9324
R15856 CSoutput.n446 CSoutput.n445 80.9324
R15857 CSoutput.n411 CSoutput.n410 80.9324
R15858 CSoutput.n413 CSoutput.n412 80.9324
R15859 CSoutput.n415 CSoutput.n414 80.9324
R15860 CSoutput.n417 CSoutput.n416 80.9324
R15861 CSoutput.n419 CSoutput.n418 80.9324
R15862 CSoutput.n421 CSoutput.n420 80.9324
R15863 CSoutput.n423 CSoutput.n422 80.9324
R15864 CSoutput.n425 CSoutput.n424 80.9324
R15865 CSoutput.n427 CSoutput.n426 80.9324
R15866 CSoutput.n25 CSoutput.n24 48.1486
R15867 CSoutput.n69 CSoutput.n3 48.1486
R15868 CSoutput.n38 CSoutput.n37 48.1486
R15869 CSoutput.n42 CSoutput.n41 48.1486
R15870 CSoutput.n51 CSoutput.n50 48.1486
R15871 CSoutput.n55 CSoutput.n54 48.1486
R15872 CSoutput.n22 CSoutput.n17 46.462
R15873 CSoutput.n72 CSoutput.n71 46.462
R15874 CSoutput.n20 CSoutput.n19 44.9055
R15875 CSoutput.n29 CSoutput.n28 43.7635
R15876 CSoutput.n65 CSoutput.n63 43.7635
R15877 CSoutput.n35 CSoutput.n13 41.7396
R15878 CSoutput.n57 CSoutput.n5 41.7396
R15879 CSoutput.n44 CSoutput.n9 37.0171
R15880 CSoutput.n48 CSoutput.n9 37.0171
R15881 CSoutput.n76 CSoutput.n75 34.9932
R15882 CSoutput.n31 CSoutput.n13 32.2947
R15883 CSoutput.n61 CSoutput.n5 32.2947
R15884 CSoutput.n30 CSoutput.n29 29.6014
R15885 CSoutput.n63 CSoutput.n62 29.6014
R15886 CSoutput.n19 CSoutput.n18 28.4085
R15887 CSoutput.n18 CSoutput.n17 25.1176
R15888 CSoutput.n72 CSoutput.n1 25.1176
R15889 CSoutput.n43 CSoutput.n42 22.0922
R15890 CSoutput.n50 CSoutput.n49 22.0922
R15891 CSoutput.n77 CSoutput.n76 21.8586
R15892 CSoutput.n37 CSoutput.n36 18.9681
R15893 CSoutput.n56 CSoutput.n55 18.9681
R15894 CSoutput.n25 CSoutput.n15 17.6292
R15895 CSoutput.n64 CSoutput.n3 17.6292
R15896 CSoutput.n24 CSoutput.n23 15.844
R15897 CSoutput.n70 CSoutput.n69 15.844
R15898 CSoutput.n38 CSoutput.n11 14.5051
R15899 CSoutput.n54 CSoutput.n7 14.5051
R15900 CSoutput.n469 CSoutput.n78 11.4982
R15901 CSoutput.n41 CSoutput.n11 11.3811
R15902 CSoutput.n51 CSoutput.n7 11.3811
R15903 CSoutput.n23 CSoutput.n22 10.0422
R15904 CSoutput.n71 CSoutput.n70 10.0422
R15905 CSoutput.n327 CSoutput.n307 9.25285
R15906 CSoutput.n117 CSoutput.n97 9.25285
R15907 CSoutput.n387 CSoutput.n367 8.98182
R15908 CSoutput.n447 CSoutput.n427 8.98182
R15909 CSoutput.n408 CSoutput.n348 8.9496
R15910 CSoutput.n28 CSoutput.n15 8.25698
R15911 CSoutput.n65 CSoutput.n64 8.25698
R15912 CSoutput.n348 CSoutput.n347 7.12641
R15913 CSoutput.n138 CSoutput.n137 7.12641
R15914 CSoutput.n36 CSoutput.n35 6.91809
R15915 CSoutput.n57 CSoutput.n56 6.91809
R15916 CSoutput.n408 CSoutput.n407 6.02792
R15917 CSoutput.n468 CSoutput.n467 6.02792
R15918 CSoutput.n469 CSoutput.n138 5.35716
R15919 CSoutput.n407 CSoutput.n406 5.25266
R15920 CSoutput.n387 CSoutput.n386 5.25266
R15921 CSoutput.n467 CSoutput.n466 5.25266
R15922 CSoutput.n447 CSoutput.n446 5.25266
R15923 CSoutput.n347 CSoutput.n346 5.1449
R15924 CSoutput.n327 CSoutput.n326 5.1449
R15925 CSoutput.n137 CSoutput.n136 5.1449
R15926 CSoutput.n117 CSoutput.n116 5.1449
R15927 CSoutput.n229 CSoutput.n182 4.5005
R15928 CSoutput.n198 CSoutput.n182 4.5005
R15929 CSoutput.n193 CSoutput.n177 4.5005
R15930 CSoutput.n193 CSoutput.n179 4.5005
R15931 CSoutput.n193 CSoutput.n176 4.5005
R15932 CSoutput.n193 CSoutput.n180 4.5005
R15933 CSoutput.n193 CSoutput.n175 4.5005
R15934 CSoutput.n193 CSoutput.t260 4.5005
R15935 CSoutput.n193 CSoutput.n174 4.5005
R15936 CSoutput.n193 CSoutput.n181 4.5005
R15937 CSoutput.n193 CSoutput.n182 4.5005
R15938 CSoutput.n191 CSoutput.n177 4.5005
R15939 CSoutput.n191 CSoutput.n179 4.5005
R15940 CSoutput.n191 CSoutput.n176 4.5005
R15941 CSoutput.n191 CSoutput.n180 4.5005
R15942 CSoutput.n191 CSoutput.n175 4.5005
R15943 CSoutput.n191 CSoutput.t260 4.5005
R15944 CSoutput.n191 CSoutput.n174 4.5005
R15945 CSoutput.n191 CSoutput.n181 4.5005
R15946 CSoutput.n191 CSoutput.n182 4.5005
R15947 CSoutput.n190 CSoutput.n177 4.5005
R15948 CSoutput.n190 CSoutput.n179 4.5005
R15949 CSoutput.n190 CSoutput.n176 4.5005
R15950 CSoutput.n190 CSoutput.n180 4.5005
R15951 CSoutput.n190 CSoutput.n175 4.5005
R15952 CSoutput.n190 CSoutput.t260 4.5005
R15953 CSoutput.n190 CSoutput.n174 4.5005
R15954 CSoutput.n190 CSoutput.n181 4.5005
R15955 CSoutput.n190 CSoutput.n182 4.5005
R15956 CSoutput.n275 CSoutput.n177 4.5005
R15957 CSoutput.n275 CSoutput.n179 4.5005
R15958 CSoutput.n275 CSoutput.n176 4.5005
R15959 CSoutput.n275 CSoutput.n180 4.5005
R15960 CSoutput.n275 CSoutput.n175 4.5005
R15961 CSoutput.n275 CSoutput.t260 4.5005
R15962 CSoutput.n275 CSoutput.n174 4.5005
R15963 CSoutput.n275 CSoutput.n181 4.5005
R15964 CSoutput.n275 CSoutput.n182 4.5005
R15965 CSoutput.n273 CSoutput.n177 4.5005
R15966 CSoutput.n273 CSoutput.n179 4.5005
R15967 CSoutput.n273 CSoutput.n176 4.5005
R15968 CSoutput.n273 CSoutput.n180 4.5005
R15969 CSoutput.n273 CSoutput.n175 4.5005
R15970 CSoutput.n273 CSoutput.t260 4.5005
R15971 CSoutput.n273 CSoutput.n174 4.5005
R15972 CSoutput.n273 CSoutput.n181 4.5005
R15973 CSoutput.n271 CSoutput.n177 4.5005
R15974 CSoutput.n271 CSoutput.n179 4.5005
R15975 CSoutput.n271 CSoutput.n176 4.5005
R15976 CSoutput.n271 CSoutput.n180 4.5005
R15977 CSoutput.n271 CSoutput.n175 4.5005
R15978 CSoutput.n271 CSoutput.t260 4.5005
R15979 CSoutput.n271 CSoutput.n174 4.5005
R15980 CSoutput.n271 CSoutput.n181 4.5005
R15981 CSoutput.n201 CSoutput.n177 4.5005
R15982 CSoutput.n201 CSoutput.n179 4.5005
R15983 CSoutput.n201 CSoutput.n176 4.5005
R15984 CSoutput.n201 CSoutput.n180 4.5005
R15985 CSoutput.n201 CSoutput.n175 4.5005
R15986 CSoutput.n201 CSoutput.t260 4.5005
R15987 CSoutput.n201 CSoutput.n174 4.5005
R15988 CSoutput.n201 CSoutput.n181 4.5005
R15989 CSoutput.n201 CSoutput.n182 4.5005
R15990 CSoutput.n200 CSoutput.n177 4.5005
R15991 CSoutput.n200 CSoutput.n179 4.5005
R15992 CSoutput.n200 CSoutput.n176 4.5005
R15993 CSoutput.n200 CSoutput.n180 4.5005
R15994 CSoutput.n200 CSoutput.n175 4.5005
R15995 CSoutput.n200 CSoutput.t260 4.5005
R15996 CSoutput.n200 CSoutput.n174 4.5005
R15997 CSoutput.n200 CSoutput.n181 4.5005
R15998 CSoutput.n200 CSoutput.n182 4.5005
R15999 CSoutput.n204 CSoutput.n177 4.5005
R16000 CSoutput.n204 CSoutput.n179 4.5005
R16001 CSoutput.n204 CSoutput.n176 4.5005
R16002 CSoutput.n204 CSoutput.n180 4.5005
R16003 CSoutput.n204 CSoutput.n175 4.5005
R16004 CSoutput.n204 CSoutput.t260 4.5005
R16005 CSoutput.n204 CSoutput.n174 4.5005
R16006 CSoutput.n204 CSoutput.n181 4.5005
R16007 CSoutput.n204 CSoutput.n182 4.5005
R16008 CSoutput.n203 CSoutput.n177 4.5005
R16009 CSoutput.n203 CSoutput.n179 4.5005
R16010 CSoutput.n203 CSoutput.n176 4.5005
R16011 CSoutput.n203 CSoutput.n180 4.5005
R16012 CSoutput.n203 CSoutput.n175 4.5005
R16013 CSoutput.n203 CSoutput.t260 4.5005
R16014 CSoutput.n203 CSoutput.n174 4.5005
R16015 CSoutput.n203 CSoutput.n181 4.5005
R16016 CSoutput.n203 CSoutput.n182 4.5005
R16017 CSoutput.n186 CSoutput.n177 4.5005
R16018 CSoutput.n186 CSoutput.n179 4.5005
R16019 CSoutput.n186 CSoutput.n176 4.5005
R16020 CSoutput.n186 CSoutput.n180 4.5005
R16021 CSoutput.n186 CSoutput.n175 4.5005
R16022 CSoutput.n186 CSoutput.t260 4.5005
R16023 CSoutput.n186 CSoutput.n174 4.5005
R16024 CSoutput.n186 CSoutput.n181 4.5005
R16025 CSoutput.n186 CSoutput.n182 4.5005
R16026 CSoutput.n278 CSoutput.n177 4.5005
R16027 CSoutput.n278 CSoutput.n179 4.5005
R16028 CSoutput.n278 CSoutput.n176 4.5005
R16029 CSoutput.n278 CSoutput.n180 4.5005
R16030 CSoutput.n278 CSoutput.n175 4.5005
R16031 CSoutput.n278 CSoutput.t260 4.5005
R16032 CSoutput.n278 CSoutput.n174 4.5005
R16033 CSoutput.n278 CSoutput.n181 4.5005
R16034 CSoutput.n278 CSoutput.n182 4.5005
R16035 CSoutput.n265 CSoutput.n236 4.5005
R16036 CSoutput.n265 CSoutput.n242 4.5005
R16037 CSoutput.n223 CSoutput.n212 4.5005
R16038 CSoutput.n223 CSoutput.n214 4.5005
R16039 CSoutput.n223 CSoutput.n211 4.5005
R16040 CSoutput.n223 CSoutput.n215 4.5005
R16041 CSoutput.n223 CSoutput.n210 4.5005
R16042 CSoutput.n223 CSoutput.t256 4.5005
R16043 CSoutput.n223 CSoutput.n209 4.5005
R16044 CSoutput.n223 CSoutput.n216 4.5005
R16045 CSoutput.n265 CSoutput.n223 4.5005
R16046 CSoutput.n244 CSoutput.n212 4.5005
R16047 CSoutput.n244 CSoutput.n214 4.5005
R16048 CSoutput.n244 CSoutput.n211 4.5005
R16049 CSoutput.n244 CSoutput.n215 4.5005
R16050 CSoutput.n244 CSoutput.n210 4.5005
R16051 CSoutput.n244 CSoutput.t256 4.5005
R16052 CSoutput.n244 CSoutput.n209 4.5005
R16053 CSoutput.n244 CSoutput.n216 4.5005
R16054 CSoutput.n265 CSoutput.n244 4.5005
R16055 CSoutput.n222 CSoutput.n212 4.5005
R16056 CSoutput.n222 CSoutput.n214 4.5005
R16057 CSoutput.n222 CSoutput.n211 4.5005
R16058 CSoutput.n222 CSoutput.n215 4.5005
R16059 CSoutput.n222 CSoutput.n210 4.5005
R16060 CSoutput.n222 CSoutput.t256 4.5005
R16061 CSoutput.n222 CSoutput.n209 4.5005
R16062 CSoutput.n222 CSoutput.n216 4.5005
R16063 CSoutput.n265 CSoutput.n222 4.5005
R16064 CSoutput.n246 CSoutput.n212 4.5005
R16065 CSoutput.n246 CSoutput.n214 4.5005
R16066 CSoutput.n246 CSoutput.n211 4.5005
R16067 CSoutput.n246 CSoutput.n215 4.5005
R16068 CSoutput.n246 CSoutput.n210 4.5005
R16069 CSoutput.n246 CSoutput.t256 4.5005
R16070 CSoutput.n246 CSoutput.n209 4.5005
R16071 CSoutput.n246 CSoutput.n216 4.5005
R16072 CSoutput.n265 CSoutput.n246 4.5005
R16073 CSoutput.n212 CSoutput.n207 4.5005
R16074 CSoutput.n214 CSoutput.n207 4.5005
R16075 CSoutput.n211 CSoutput.n207 4.5005
R16076 CSoutput.n215 CSoutput.n207 4.5005
R16077 CSoutput.n210 CSoutput.n207 4.5005
R16078 CSoutput.t256 CSoutput.n207 4.5005
R16079 CSoutput.n209 CSoutput.n207 4.5005
R16080 CSoutput.n216 CSoutput.n207 4.5005
R16081 CSoutput.n268 CSoutput.n212 4.5005
R16082 CSoutput.n268 CSoutput.n214 4.5005
R16083 CSoutput.n268 CSoutput.n211 4.5005
R16084 CSoutput.n268 CSoutput.n215 4.5005
R16085 CSoutput.n268 CSoutput.n210 4.5005
R16086 CSoutput.n268 CSoutput.t256 4.5005
R16087 CSoutput.n268 CSoutput.n209 4.5005
R16088 CSoutput.n268 CSoutput.n216 4.5005
R16089 CSoutput.n266 CSoutput.n212 4.5005
R16090 CSoutput.n266 CSoutput.n214 4.5005
R16091 CSoutput.n266 CSoutput.n211 4.5005
R16092 CSoutput.n266 CSoutput.n215 4.5005
R16093 CSoutput.n266 CSoutput.n210 4.5005
R16094 CSoutput.n266 CSoutput.t256 4.5005
R16095 CSoutput.n266 CSoutput.n209 4.5005
R16096 CSoutput.n266 CSoutput.n216 4.5005
R16097 CSoutput.n266 CSoutput.n265 4.5005
R16098 CSoutput.n248 CSoutput.n212 4.5005
R16099 CSoutput.n248 CSoutput.n214 4.5005
R16100 CSoutput.n248 CSoutput.n211 4.5005
R16101 CSoutput.n248 CSoutput.n215 4.5005
R16102 CSoutput.n248 CSoutput.n210 4.5005
R16103 CSoutput.n248 CSoutput.t256 4.5005
R16104 CSoutput.n248 CSoutput.n209 4.5005
R16105 CSoutput.n248 CSoutput.n216 4.5005
R16106 CSoutput.n265 CSoutput.n248 4.5005
R16107 CSoutput.n220 CSoutput.n212 4.5005
R16108 CSoutput.n220 CSoutput.n214 4.5005
R16109 CSoutput.n220 CSoutput.n211 4.5005
R16110 CSoutput.n220 CSoutput.n215 4.5005
R16111 CSoutput.n220 CSoutput.n210 4.5005
R16112 CSoutput.n220 CSoutput.t256 4.5005
R16113 CSoutput.n220 CSoutput.n209 4.5005
R16114 CSoutput.n220 CSoutput.n216 4.5005
R16115 CSoutput.n265 CSoutput.n220 4.5005
R16116 CSoutput.n250 CSoutput.n212 4.5005
R16117 CSoutput.n250 CSoutput.n214 4.5005
R16118 CSoutput.n250 CSoutput.n211 4.5005
R16119 CSoutput.n250 CSoutput.n215 4.5005
R16120 CSoutput.n250 CSoutput.n210 4.5005
R16121 CSoutput.n250 CSoutput.t256 4.5005
R16122 CSoutput.n250 CSoutput.n209 4.5005
R16123 CSoutput.n250 CSoutput.n216 4.5005
R16124 CSoutput.n265 CSoutput.n250 4.5005
R16125 CSoutput.n219 CSoutput.n212 4.5005
R16126 CSoutput.n219 CSoutput.n214 4.5005
R16127 CSoutput.n219 CSoutput.n211 4.5005
R16128 CSoutput.n219 CSoutput.n215 4.5005
R16129 CSoutput.n219 CSoutput.n210 4.5005
R16130 CSoutput.n219 CSoutput.t256 4.5005
R16131 CSoutput.n219 CSoutput.n209 4.5005
R16132 CSoutput.n219 CSoutput.n216 4.5005
R16133 CSoutput.n265 CSoutput.n219 4.5005
R16134 CSoutput.n264 CSoutput.n212 4.5005
R16135 CSoutput.n264 CSoutput.n214 4.5005
R16136 CSoutput.n264 CSoutput.n211 4.5005
R16137 CSoutput.n264 CSoutput.n215 4.5005
R16138 CSoutput.n264 CSoutput.n210 4.5005
R16139 CSoutput.n264 CSoutput.t256 4.5005
R16140 CSoutput.n264 CSoutput.n209 4.5005
R16141 CSoutput.n264 CSoutput.n216 4.5005
R16142 CSoutput.n265 CSoutput.n264 4.5005
R16143 CSoutput.n263 CSoutput.n148 4.5005
R16144 CSoutput.n164 CSoutput.n148 4.5005
R16145 CSoutput.n159 CSoutput.n143 4.5005
R16146 CSoutput.n159 CSoutput.n145 4.5005
R16147 CSoutput.n159 CSoutput.n142 4.5005
R16148 CSoutput.n159 CSoutput.n146 4.5005
R16149 CSoutput.n159 CSoutput.n141 4.5005
R16150 CSoutput.n159 CSoutput.t255 4.5005
R16151 CSoutput.n159 CSoutput.n140 4.5005
R16152 CSoutput.n159 CSoutput.n147 4.5005
R16153 CSoutput.n159 CSoutput.n148 4.5005
R16154 CSoutput.n157 CSoutput.n143 4.5005
R16155 CSoutput.n157 CSoutput.n145 4.5005
R16156 CSoutput.n157 CSoutput.n142 4.5005
R16157 CSoutput.n157 CSoutput.n146 4.5005
R16158 CSoutput.n157 CSoutput.n141 4.5005
R16159 CSoutput.n157 CSoutput.t255 4.5005
R16160 CSoutput.n157 CSoutput.n140 4.5005
R16161 CSoutput.n157 CSoutput.n147 4.5005
R16162 CSoutput.n157 CSoutput.n148 4.5005
R16163 CSoutput.n156 CSoutput.n143 4.5005
R16164 CSoutput.n156 CSoutput.n145 4.5005
R16165 CSoutput.n156 CSoutput.n142 4.5005
R16166 CSoutput.n156 CSoutput.n146 4.5005
R16167 CSoutput.n156 CSoutput.n141 4.5005
R16168 CSoutput.n156 CSoutput.t255 4.5005
R16169 CSoutput.n156 CSoutput.n140 4.5005
R16170 CSoutput.n156 CSoutput.n147 4.5005
R16171 CSoutput.n156 CSoutput.n148 4.5005
R16172 CSoutput.n285 CSoutput.n143 4.5005
R16173 CSoutput.n285 CSoutput.n145 4.5005
R16174 CSoutput.n285 CSoutput.n142 4.5005
R16175 CSoutput.n285 CSoutput.n146 4.5005
R16176 CSoutput.n285 CSoutput.n141 4.5005
R16177 CSoutput.n285 CSoutput.t255 4.5005
R16178 CSoutput.n285 CSoutput.n140 4.5005
R16179 CSoutput.n285 CSoutput.n147 4.5005
R16180 CSoutput.n285 CSoutput.n148 4.5005
R16181 CSoutput.n283 CSoutput.n143 4.5005
R16182 CSoutput.n283 CSoutput.n145 4.5005
R16183 CSoutput.n283 CSoutput.n142 4.5005
R16184 CSoutput.n283 CSoutput.n146 4.5005
R16185 CSoutput.n283 CSoutput.n141 4.5005
R16186 CSoutput.n283 CSoutput.t255 4.5005
R16187 CSoutput.n283 CSoutput.n140 4.5005
R16188 CSoutput.n283 CSoutput.n147 4.5005
R16189 CSoutput.n281 CSoutput.n143 4.5005
R16190 CSoutput.n281 CSoutput.n145 4.5005
R16191 CSoutput.n281 CSoutput.n142 4.5005
R16192 CSoutput.n281 CSoutput.n146 4.5005
R16193 CSoutput.n281 CSoutput.n141 4.5005
R16194 CSoutput.n281 CSoutput.t255 4.5005
R16195 CSoutput.n281 CSoutput.n140 4.5005
R16196 CSoutput.n281 CSoutput.n147 4.5005
R16197 CSoutput.n167 CSoutput.n143 4.5005
R16198 CSoutput.n167 CSoutput.n145 4.5005
R16199 CSoutput.n167 CSoutput.n142 4.5005
R16200 CSoutput.n167 CSoutput.n146 4.5005
R16201 CSoutput.n167 CSoutput.n141 4.5005
R16202 CSoutput.n167 CSoutput.t255 4.5005
R16203 CSoutput.n167 CSoutput.n140 4.5005
R16204 CSoutput.n167 CSoutput.n147 4.5005
R16205 CSoutput.n167 CSoutput.n148 4.5005
R16206 CSoutput.n166 CSoutput.n143 4.5005
R16207 CSoutput.n166 CSoutput.n145 4.5005
R16208 CSoutput.n166 CSoutput.n142 4.5005
R16209 CSoutput.n166 CSoutput.n146 4.5005
R16210 CSoutput.n166 CSoutput.n141 4.5005
R16211 CSoutput.n166 CSoutput.t255 4.5005
R16212 CSoutput.n166 CSoutput.n140 4.5005
R16213 CSoutput.n166 CSoutput.n147 4.5005
R16214 CSoutput.n166 CSoutput.n148 4.5005
R16215 CSoutput.n170 CSoutput.n143 4.5005
R16216 CSoutput.n170 CSoutput.n145 4.5005
R16217 CSoutput.n170 CSoutput.n142 4.5005
R16218 CSoutput.n170 CSoutput.n146 4.5005
R16219 CSoutput.n170 CSoutput.n141 4.5005
R16220 CSoutput.n170 CSoutput.t255 4.5005
R16221 CSoutput.n170 CSoutput.n140 4.5005
R16222 CSoutput.n170 CSoutput.n147 4.5005
R16223 CSoutput.n170 CSoutput.n148 4.5005
R16224 CSoutput.n169 CSoutput.n143 4.5005
R16225 CSoutput.n169 CSoutput.n145 4.5005
R16226 CSoutput.n169 CSoutput.n142 4.5005
R16227 CSoutput.n169 CSoutput.n146 4.5005
R16228 CSoutput.n169 CSoutput.n141 4.5005
R16229 CSoutput.n169 CSoutput.t255 4.5005
R16230 CSoutput.n169 CSoutput.n140 4.5005
R16231 CSoutput.n169 CSoutput.n147 4.5005
R16232 CSoutput.n169 CSoutput.n148 4.5005
R16233 CSoutput.n152 CSoutput.n143 4.5005
R16234 CSoutput.n152 CSoutput.n145 4.5005
R16235 CSoutput.n152 CSoutput.n142 4.5005
R16236 CSoutput.n152 CSoutput.n146 4.5005
R16237 CSoutput.n152 CSoutput.n141 4.5005
R16238 CSoutput.n152 CSoutput.t255 4.5005
R16239 CSoutput.n152 CSoutput.n140 4.5005
R16240 CSoutput.n152 CSoutput.n147 4.5005
R16241 CSoutput.n152 CSoutput.n148 4.5005
R16242 CSoutput.n288 CSoutput.n143 4.5005
R16243 CSoutput.n288 CSoutput.n145 4.5005
R16244 CSoutput.n288 CSoutput.n142 4.5005
R16245 CSoutput.n288 CSoutput.n146 4.5005
R16246 CSoutput.n288 CSoutput.n141 4.5005
R16247 CSoutput.n288 CSoutput.t255 4.5005
R16248 CSoutput.n288 CSoutput.n140 4.5005
R16249 CSoutput.n288 CSoutput.n147 4.5005
R16250 CSoutput.n288 CSoutput.n148 4.5005
R16251 CSoutput.n347 CSoutput.n327 4.10845
R16252 CSoutput.n137 CSoutput.n117 4.10845
R16253 CSoutput.n345 CSoutput.t7 4.06363
R16254 CSoutput.n345 CSoutput.t63 4.06363
R16255 CSoutput.n343 CSoutput.t114 4.06363
R16256 CSoutput.n343 CSoutput.t49 4.06363
R16257 CSoutput.n341 CSoutput.t91 4.06363
R16258 CSoutput.n341 CSoutput.t75 4.06363
R16259 CSoutput.n339 CSoutput.t8 4.06363
R16260 CSoutput.n339 CSoutput.t45 4.06363
R16261 CSoutput.n337 CSoutput.t1 4.06363
R16262 CSoutput.n337 CSoutput.t0 4.06363
R16263 CSoutput.n335 CSoutput.t55 4.06363
R16264 CSoutput.n335 CSoutput.t44 4.06363
R16265 CSoutput.n333 CSoutput.t11 4.06363
R16266 CSoutput.n333 CSoutput.t35 4.06363
R16267 CSoutput.n331 CSoutput.t112 4.06363
R16268 CSoutput.n331 CSoutput.t42 4.06363
R16269 CSoutput.n329 CSoutput.t239 4.06363
R16270 CSoutput.n329 CSoutput.t47 4.06363
R16271 CSoutput.n328 CSoutput.t69 4.06363
R16272 CSoutput.n328 CSoutput.t68 4.06363
R16273 CSoutput.n325 CSoutput.t97 4.06363
R16274 CSoutput.n325 CSoutput.t60 4.06363
R16275 CSoutput.n323 CSoutput.t236 4.06363
R16276 CSoutput.n323 CSoutput.t109 4.06363
R16277 CSoutput.n321 CSoutput.t108 4.06363
R16278 CSoutput.n321 CSoutput.t103 4.06363
R16279 CSoutput.n319 CSoutput.t20 4.06363
R16280 CSoutput.n319 CSoutput.t111 4.06363
R16281 CSoutput.n317 CSoutput.t13 4.06363
R16282 CSoutput.n317 CSoutput.t12 4.06363
R16283 CSoutput.n315 CSoutput.t31 4.06363
R16284 CSoutput.n315 CSoutput.t82 4.06363
R16285 CSoutput.n313 CSoutput.t4 4.06363
R16286 CSoutput.n313 CSoutput.t92 4.06363
R16287 CSoutput.n311 CSoutput.t54 4.06363
R16288 CSoutput.n311 CSoutput.t61 4.06363
R16289 CSoutput.n309 CSoutput.t102 4.06363
R16290 CSoutput.n309 CSoutput.t106 4.06363
R16291 CSoutput.n308 CSoutput.t57 4.06363
R16292 CSoutput.n308 CSoutput.t56 4.06363
R16293 CSoutput.n306 CSoutput.t70 4.06363
R16294 CSoutput.n306 CSoutput.t94 4.06363
R16295 CSoutput.n304 CSoutput.t39 4.06363
R16296 CSoutput.n304 CSoutput.t26 4.06363
R16297 CSoutput.n302 CSoutput.t237 4.06363
R16298 CSoutput.n302 CSoutput.t10 4.06363
R16299 CSoutput.n300 CSoutput.t98 4.06363
R16300 CSoutput.n300 CSoutput.t93 4.06363
R16301 CSoutput.n298 CSoutput.t30 4.06363
R16302 CSoutput.n298 CSoutput.t19 4.06363
R16303 CSoutput.n296 CSoutput.t71 4.06363
R16304 CSoutput.n296 CSoutput.t81 4.06363
R16305 CSoutput.n294 CSoutput.t33 4.06363
R16306 CSoutput.n294 CSoutput.t115 4.06363
R16307 CSoutput.n292 CSoutput.t90 4.06363
R16308 CSoutput.n292 CSoutput.t65 4.06363
R16309 CSoutput.n290 CSoutput.t96 4.06363
R16310 CSoutput.n290 CSoutput.t77 4.06363
R16311 CSoutput.n289 CSoutput.t78 4.06363
R16312 CSoutput.n289 CSoutput.t110 4.06363
R16313 CSoutput.n118 CSoutput.t22 4.06363
R16314 CSoutput.n118 CSoutput.t23 4.06363
R16315 CSoutput.n119 CSoutput.t43 4.06363
R16316 CSoutput.n119 CSoutput.t27 4.06363
R16317 CSoutput.n121 CSoutput.t24 4.06363
R16318 CSoutput.n121 CSoutput.t85 4.06363
R16319 CSoutput.n123 CSoutput.t72 4.06363
R16320 CSoutput.n123 CSoutput.t59 4.06363
R16321 CSoutput.n125 CSoutput.t52 4.06363
R16322 CSoutput.n125 CSoutput.t5 4.06363
R16323 CSoutput.n127 CSoutput.t104 4.06363
R16324 CSoutput.n127 CSoutput.t105 4.06363
R16325 CSoutput.n129 CSoutput.t67 4.06363
R16326 CSoutput.n129 CSoutput.t95 4.06363
R16327 CSoutput.n131 CSoutput.t46 4.06363
R16328 CSoutput.n131 CSoutput.t66 4.06363
R16329 CSoutput.n133 CSoutput.t6 4.06363
R16330 CSoutput.n133 CSoutput.t51 4.06363
R16331 CSoutput.n135 CSoutput.t25 4.06363
R16332 CSoutput.n135 CSoutput.t86 4.06363
R16333 CSoutput.n98 CSoutput.t238 4.06363
R16334 CSoutput.n98 CSoutput.t74 4.06363
R16335 CSoutput.n99 CSoutput.t40 4.06363
R16336 CSoutput.n99 CSoutput.t16 4.06363
R16337 CSoutput.n101 CSoutput.t14 4.06363
R16338 CSoutput.n101 CSoutput.t62 4.06363
R16339 CSoutput.n103 CSoutput.t41 4.06363
R16340 CSoutput.n103 CSoutput.t34 4.06363
R16341 CSoutput.n105 CSoutput.t28 4.06363
R16342 CSoutput.n105 CSoutput.t84 4.06363
R16343 CSoutput.n107 CSoutput.t2 4.06363
R16344 CSoutput.n107 CSoutput.t3 4.06363
R16345 CSoutput.n109 CSoutput.t101 4.06363
R16346 CSoutput.n109 CSoutput.t88 4.06363
R16347 CSoutput.n111 CSoutput.t80 4.06363
R16348 CSoutput.n111 CSoutput.t100 4.06363
R16349 CSoutput.n113 CSoutput.t36 4.06363
R16350 CSoutput.n113 CSoutput.t48 4.06363
R16351 CSoutput.n115 CSoutput.t107 4.06363
R16352 CSoutput.n115 CSoutput.t79 4.06363
R16353 CSoutput.n79 CSoutput.t83 4.06363
R16354 CSoutput.n79 CSoutput.t15 4.06363
R16355 CSoutput.n80 CSoutput.t73 4.06363
R16356 CSoutput.n80 CSoutput.t99 4.06363
R16357 CSoutput.n82 CSoutput.t64 4.06363
R16358 CSoutput.n82 CSoutput.t29 4.06363
R16359 CSoutput.n84 CSoutput.t9 4.06363
R16360 CSoutput.n84 CSoutput.t32 4.06363
R16361 CSoutput.n86 CSoutput.t17 4.06363
R16362 CSoutput.n86 CSoutput.t58 4.06363
R16363 CSoutput.n88 CSoutput.t18 4.06363
R16364 CSoutput.n88 CSoutput.t50 4.06363
R16365 CSoutput.n90 CSoutput.t76 4.06363
R16366 CSoutput.n90 CSoutput.t37 4.06363
R16367 CSoutput.n92 CSoutput.t87 4.06363
R16368 CSoutput.n92 CSoutput.t21 4.06363
R16369 CSoutput.n94 CSoutput.t89 4.06363
R16370 CSoutput.n94 CSoutput.t38 4.06363
R16371 CSoutput.n96 CSoutput.t53 4.06363
R16372 CSoutput.n96 CSoutput.t113 4.06363
R16373 CSoutput.n44 CSoutput.n43 3.79402
R16374 CSoutput.n49 CSoutput.n48 3.79402
R16375 CSoutput.n407 CSoutput.n387 3.72967
R16376 CSoutput.n467 CSoutput.n447 3.72967
R16377 CSoutput.n469 CSoutput.n468 3.57343
R16378 CSoutput.n468 CSoutput.n408 3.42304
R16379 CSoutput.n405 CSoutput.t165 2.82907
R16380 CSoutput.n405 CSoutput.t131 2.82907
R16381 CSoutput.n403 CSoutput.t116 2.82907
R16382 CSoutput.n403 CSoutput.t160 2.82907
R16383 CSoutput.n401 CSoutput.t150 2.82907
R16384 CSoutput.n401 CSoutput.t140 2.82907
R16385 CSoutput.n399 CSoutput.t128 2.82907
R16386 CSoutput.n399 CSoutput.t219 2.82907
R16387 CSoutput.n397 CSoutput.t143 2.82907
R16388 CSoutput.n397 CSoutput.t147 2.82907
R16389 CSoutput.n395 CSoutput.t142 2.82907
R16390 CSoutput.n395 CSoutput.t235 2.82907
R16391 CSoutput.n393 CSoutput.t166 2.82907
R16392 CSoutput.n393 CSoutput.t133 2.82907
R16393 CSoutput.n391 CSoutput.t121 2.82907
R16394 CSoutput.n391 CSoutput.t205 2.82907
R16395 CSoutput.n389 CSoutput.t152 2.82907
R16396 CSoutput.n389 CSoutput.t158 2.82907
R16397 CSoutput.n388 CSoutput.t132 2.82907
R16398 CSoutput.n388 CSoutput.t223 2.82907
R16399 CSoutput.n385 CSoutput.t168 2.82907
R16400 CSoutput.n385 CSoutput.t181 2.82907
R16401 CSoutput.n383 CSoutput.t186 2.82907
R16402 CSoutput.n383 CSoutput.t190 2.82907
R16403 CSoutput.n381 CSoutput.t201 2.82907
R16404 CSoutput.n381 CSoutput.t176 2.82907
R16405 CSoutput.n379 CSoutput.t177 2.82907
R16406 CSoutput.n379 CSoutput.t185 2.82907
R16407 CSoutput.n377 CSoutput.t120 2.82907
R16408 CSoutput.n377 CSoutput.t202 2.82907
R16409 CSoutput.n375 CSoutput.t200 2.82907
R16410 CSoutput.n375 CSoutput.t174 2.82907
R16411 CSoutput.n373 CSoutput.t221 2.82907
R16412 CSoutput.n373 CSoutput.t118 2.82907
R16413 CSoutput.n371 CSoutput.t119 2.82907
R16414 CSoutput.n371 CSoutput.t210 2.82907
R16415 CSoutput.n369 CSoutput.t129 2.82907
R16416 CSoutput.n369 CSoutput.t220 2.82907
R16417 CSoutput.n368 CSoutput.t227 2.82907
R16418 CSoutput.n368 CSoutput.t117 2.82907
R16419 CSoutput.n366 CSoutput.t231 2.82907
R16420 CSoutput.n366 CSoutput.t175 2.82907
R16421 CSoutput.n364 CSoutput.t204 2.82907
R16422 CSoutput.n364 CSoutput.t215 2.82907
R16423 CSoutput.n362 CSoutput.t125 2.82907
R16424 CSoutput.n362 CSoutput.t151 2.82907
R16425 CSoutput.n360 CSoutput.t139 2.82907
R16426 CSoutput.n360 CSoutput.t171 2.82907
R16427 CSoutput.n358 CSoutput.t184 2.82907
R16428 CSoutput.n358 CSoutput.t198 2.82907
R16429 CSoutput.n356 CSoutput.t167 2.82907
R16430 CSoutput.n356 CSoutput.t222 2.82907
R16431 CSoutput.n354 CSoutput.t191 2.82907
R16432 CSoutput.n354 CSoutput.t157 2.82907
R16433 CSoutput.n352 CSoutput.t144 2.82907
R16434 CSoutput.n352 CSoutput.t170 2.82907
R16435 CSoutput.n350 CSoutput.t154 2.82907
R16436 CSoutput.n350 CSoutput.t163 2.82907
R16437 CSoutput.n349 CSoutput.t164 2.82907
R16438 CSoutput.n349 CSoutput.t232 2.82907
R16439 CSoutput.n448 CSoutput.t182 2.82907
R16440 CSoutput.n448 CSoutput.t214 2.82907
R16441 CSoutput.n449 CSoutput.t145 2.82907
R16442 CSoutput.n449 CSoutput.t162 2.82907
R16443 CSoutput.n451 CSoutput.t172 2.82907
R16444 CSoutput.n451 CSoutput.t193 2.82907
R16445 CSoutput.n453 CSoutput.t216 2.82907
R16446 CSoutput.n453 CSoutput.t178 2.82907
R16447 CSoutput.n455 CSoutput.t188 2.82907
R16448 CSoutput.n455 CSoutput.t228 2.82907
R16449 CSoutput.n457 CSoutput.t123 2.82907
R16450 CSoutput.n457 CSoutput.t148 2.82907
R16451 CSoutput.n459 CSoutput.t179 2.82907
R16452 CSoutput.n459 CSoutput.t208 2.82907
R16453 CSoutput.n461 CSoutput.t224 2.82907
R16454 CSoutput.n461 CSoutput.t134 2.82907
R16455 CSoutput.n463 CSoutput.t169 2.82907
R16456 CSoutput.n463 CSoutput.t189 2.82907
R16457 CSoutput.n465 CSoutput.t124 2.82907
R16458 CSoutput.n465 CSoutput.t159 2.82907
R16459 CSoutput.n428 CSoutput.t135 2.82907
R16460 CSoutput.n428 CSoutput.t126 2.82907
R16461 CSoutput.n429 CSoutput.t122 2.82907
R16462 CSoutput.n429 CSoutput.t233 2.82907
R16463 CSoutput.n431 CSoutput.t234 2.82907
R16464 CSoutput.n431 CSoutput.t136 2.82907
R16465 CSoutput.n433 CSoutput.t137 2.82907
R16466 CSoutput.n433 CSoutput.t194 2.82907
R16467 CSoutput.n435 CSoutput.t195 2.82907
R16468 CSoutput.n435 CSoutput.t226 2.82907
R16469 CSoutput.n437 CSoutput.t229 2.82907
R16470 CSoutput.n437 CSoutput.t218 2.82907
R16471 CSoutput.n439 CSoutput.t209 2.82907
R16472 CSoutput.n439 CSoutput.t196 2.82907
R16473 CSoutput.n441 CSoutput.t197 2.82907
R16474 CSoutput.n441 CSoutput.t230 2.82907
R16475 CSoutput.n443 CSoutput.t183 2.82907
R16476 CSoutput.n443 CSoutput.t211 2.82907
R16477 CSoutput.n445 CSoutput.t217 2.82907
R16478 CSoutput.n445 CSoutput.t192 2.82907
R16479 CSoutput.n409 CSoutput.t146 2.82907
R16480 CSoutput.n409 CSoutput.t203 2.82907
R16481 CSoutput.n410 CSoutput.t199 2.82907
R16482 CSoutput.n410 CSoutput.t173 2.82907
R16483 CSoutput.n412 CSoutput.t207 2.82907
R16484 CSoutput.n412 CSoutput.t161 2.82907
R16485 CSoutput.n414 CSoutput.t187 2.82907
R16486 CSoutput.n414 CSoutput.t225 2.82907
R16487 CSoutput.n416 CSoutput.t141 2.82907
R16488 CSoutput.n416 CSoutput.t206 2.82907
R16489 CSoutput.n418 CSoutput.t127 2.82907
R16490 CSoutput.n418 CSoutput.t213 2.82907
R16491 CSoutput.n420 CSoutput.t212 2.82907
R16492 CSoutput.n420 CSoutput.t153 2.82907
R16493 CSoutput.n422 CSoutput.t180 2.82907
R16494 CSoutput.n422 CSoutput.t149 2.82907
R16495 CSoutput.n424 CSoutput.t155 2.82907
R16496 CSoutput.n424 CSoutput.t130 2.82907
R16497 CSoutput.n426 CSoutput.t138 2.82907
R16498 CSoutput.n426 CSoutput.t156 2.82907
R16499 CSoutput.n348 CSoutput.n138 2.57547
R16500 CSoutput.n75 CSoutput.n1 2.45513
R16501 CSoutput.n229 CSoutput.n227 2.251
R16502 CSoutput.n229 CSoutput.n226 2.251
R16503 CSoutput.n229 CSoutput.n225 2.251
R16504 CSoutput.n229 CSoutput.n224 2.251
R16505 CSoutput.n198 CSoutput.n197 2.251
R16506 CSoutput.n198 CSoutput.n196 2.251
R16507 CSoutput.n198 CSoutput.n195 2.251
R16508 CSoutput.n198 CSoutput.n194 2.251
R16509 CSoutput.n271 CSoutput.n270 2.251
R16510 CSoutput.n236 CSoutput.n234 2.251
R16511 CSoutput.n236 CSoutput.n233 2.251
R16512 CSoutput.n236 CSoutput.n232 2.251
R16513 CSoutput.n254 CSoutput.n236 2.251
R16514 CSoutput.n242 CSoutput.n241 2.251
R16515 CSoutput.n242 CSoutput.n240 2.251
R16516 CSoutput.n242 CSoutput.n239 2.251
R16517 CSoutput.n242 CSoutput.n238 2.251
R16518 CSoutput.n268 CSoutput.n208 2.251
R16519 CSoutput.n263 CSoutput.n261 2.251
R16520 CSoutput.n263 CSoutput.n260 2.251
R16521 CSoutput.n263 CSoutput.n259 2.251
R16522 CSoutput.n263 CSoutput.n258 2.251
R16523 CSoutput.n164 CSoutput.n163 2.251
R16524 CSoutput.n164 CSoutput.n162 2.251
R16525 CSoutput.n164 CSoutput.n161 2.251
R16526 CSoutput.n164 CSoutput.n160 2.251
R16527 CSoutput.n281 CSoutput.n280 2.251
R16528 CSoutput.n198 CSoutput.n178 2.2505
R16529 CSoutput.n193 CSoutput.n178 2.2505
R16530 CSoutput.n191 CSoutput.n178 2.2505
R16531 CSoutput.n190 CSoutput.n178 2.2505
R16532 CSoutput.n275 CSoutput.n178 2.2505
R16533 CSoutput.n273 CSoutput.n178 2.2505
R16534 CSoutput.n271 CSoutput.n178 2.2505
R16535 CSoutput.n201 CSoutput.n178 2.2505
R16536 CSoutput.n200 CSoutput.n178 2.2505
R16537 CSoutput.n204 CSoutput.n178 2.2505
R16538 CSoutput.n203 CSoutput.n178 2.2505
R16539 CSoutput.n186 CSoutput.n178 2.2505
R16540 CSoutput.n278 CSoutput.n178 2.2505
R16541 CSoutput.n278 CSoutput.n277 2.2505
R16542 CSoutput.n242 CSoutput.n213 2.2505
R16543 CSoutput.n223 CSoutput.n213 2.2505
R16544 CSoutput.n244 CSoutput.n213 2.2505
R16545 CSoutput.n222 CSoutput.n213 2.2505
R16546 CSoutput.n246 CSoutput.n213 2.2505
R16547 CSoutput.n213 CSoutput.n207 2.2505
R16548 CSoutput.n268 CSoutput.n213 2.2505
R16549 CSoutput.n266 CSoutput.n213 2.2505
R16550 CSoutput.n248 CSoutput.n213 2.2505
R16551 CSoutput.n220 CSoutput.n213 2.2505
R16552 CSoutput.n250 CSoutput.n213 2.2505
R16553 CSoutput.n219 CSoutput.n213 2.2505
R16554 CSoutput.n264 CSoutput.n213 2.2505
R16555 CSoutput.n264 CSoutput.n217 2.2505
R16556 CSoutput.n164 CSoutput.n144 2.2505
R16557 CSoutput.n159 CSoutput.n144 2.2505
R16558 CSoutput.n157 CSoutput.n144 2.2505
R16559 CSoutput.n156 CSoutput.n144 2.2505
R16560 CSoutput.n285 CSoutput.n144 2.2505
R16561 CSoutput.n283 CSoutput.n144 2.2505
R16562 CSoutput.n281 CSoutput.n144 2.2505
R16563 CSoutput.n167 CSoutput.n144 2.2505
R16564 CSoutput.n166 CSoutput.n144 2.2505
R16565 CSoutput.n170 CSoutput.n144 2.2505
R16566 CSoutput.n169 CSoutput.n144 2.2505
R16567 CSoutput.n152 CSoutput.n144 2.2505
R16568 CSoutput.n288 CSoutput.n144 2.2505
R16569 CSoutput.n288 CSoutput.n287 2.2505
R16570 CSoutput.n206 CSoutput.n199 2.25024
R16571 CSoutput.n206 CSoutput.n192 2.25024
R16572 CSoutput.n274 CSoutput.n206 2.25024
R16573 CSoutput.n206 CSoutput.n202 2.25024
R16574 CSoutput.n206 CSoutput.n205 2.25024
R16575 CSoutput.n206 CSoutput.n173 2.25024
R16576 CSoutput.n256 CSoutput.n253 2.25024
R16577 CSoutput.n256 CSoutput.n252 2.25024
R16578 CSoutput.n256 CSoutput.n251 2.25024
R16579 CSoutput.n256 CSoutput.n218 2.25024
R16580 CSoutput.n256 CSoutput.n255 2.25024
R16581 CSoutput.n257 CSoutput.n256 2.25024
R16582 CSoutput.n172 CSoutput.n165 2.25024
R16583 CSoutput.n172 CSoutput.n158 2.25024
R16584 CSoutput.n284 CSoutput.n172 2.25024
R16585 CSoutput.n172 CSoutput.n168 2.25024
R16586 CSoutput.n172 CSoutput.n171 2.25024
R16587 CSoutput.n172 CSoutput.n139 2.25024
R16588 CSoutput.n273 CSoutput.n183 1.50111
R16589 CSoutput.n221 CSoutput.n207 1.50111
R16590 CSoutput.n283 CSoutput.n149 1.50111
R16591 CSoutput.n229 CSoutput.n228 1.501
R16592 CSoutput.n236 CSoutput.n235 1.501
R16593 CSoutput.n263 CSoutput.n262 1.501
R16594 CSoutput.n277 CSoutput.n188 1.12536
R16595 CSoutput.n277 CSoutput.n189 1.12536
R16596 CSoutput.n277 CSoutput.n276 1.12536
R16597 CSoutput.n237 CSoutput.n217 1.12536
R16598 CSoutput.n243 CSoutput.n217 1.12536
R16599 CSoutput.n245 CSoutput.n217 1.12536
R16600 CSoutput.n287 CSoutput.n154 1.12536
R16601 CSoutput.n287 CSoutput.n155 1.12536
R16602 CSoutput.n287 CSoutput.n286 1.12536
R16603 CSoutput.n277 CSoutput.n184 1.12536
R16604 CSoutput.n277 CSoutput.n185 1.12536
R16605 CSoutput.n277 CSoutput.n187 1.12536
R16606 CSoutput.n267 CSoutput.n217 1.12536
R16607 CSoutput.n247 CSoutput.n217 1.12536
R16608 CSoutput.n249 CSoutput.n217 1.12536
R16609 CSoutput.n287 CSoutput.n150 1.12536
R16610 CSoutput.n287 CSoutput.n151 1.12536
R16611 CSoutput.n287 CSoutput.n153 1.12536
R16612 CSoutput.n31 CSoutput.n30 0.669944
R16613 CSoutput.n62 CSoutput.n61 0.669944
R16614 CSoutput.n392 CSoutput.n390 0.573776
R16615 CSoutput.n394 CSoutput.n392 0.573776
R16616 CSoutput.n396 CSoutput.n394 0.573776
R16617 CSoutput.n398 CSoutput.n396 0.573776
R16618 CSoutput.n400 CSoutput.n398 0.573776
R16619 CSoutput.n402 CSoutput.n400 0.573776
R16620 CSoutput.n404 CSoutput.n402 0.573776
R16621 CSoutput.n406 CSoutput.n404 0.573776
R16622 CSoutput.n372 CSoutput.n370 0.573776
R16623 CSoutput.n374 CSoutput.n372 0.573776
R16624 CSoutput.n376 CSoutput.n374 0.573776
R16625 CSoutput.n378 CSoutput.n376 0.573776
R16626 CSoutput.n380 CSoutput.n378 0.573776
R16627 CSoutput.n382 CSoutput.n380 0.573776
R16628 CSoutput.n384 CSoutput.n382 0.573776
R16629 CSoutput.n386 CSoutput.n384 0.573776
R16630 CSoutput.n353 CSoutput.n351 0.573776
R16631 CSoutput.n355 CSoutput.n353 0.573776
R16632 CSoutput.n357 CSoutput.n355 0.573776
R16633 CSoutput.n359 CSoutput.n357 0.573776
R16634 CSoutput.n361 CSoutput.n359 0.573776
R16635 CSoutput.n363 CSoutput.n361 0.573776
R16636 CSoutput.n365 CSoutput.n363 0.573776
R16637 CSoutput.n367 CSoutput.n365 0.573776
R16638 CSoutput.n466 CSoutput.n464 0.573776
R16639 CSoutput.n464 CSoutput.n462 0.573776
R16640 CSoutput.n462 CSoutput.n460 0.573776
R16641 CSoutput.n460 CSoutput.n458 0.573776
R16642 CSoutput.n458 CSoutput.n456 0.573776
R16643 CSoutput.n456 CSoutput.n454 0.573776
R16644 CSoutput.n454 CSoutput.n452 0.573776
R16645 CSoutput.n452 CSoutput.n450 0.573776
R16646 CSoutput.n446 CSoutput.n444 0.573776
R16647 CSoutput.n444 CSoutput.n442 0.573776
R16648 CSoutput.n442 CSoutput.n440 0.573776
R16649 CSoutput.n440 CSoutput.n438 0.573776
R16650 CSoutput.n438 CSoutput.n436 0.573776
R16651 CSoutput.n436 CSoutput.n434 0.573776
R16652 CSoutput.n434 CSoutput.n432 0.573776
R16653 CSoutput.n432 CSoutput.n430 0.573776
R16654 CSoutput.n427 CSoutput.n425 0.573776
R16655 CSoutput.n425 CSoutput.n423 0.573776
R16656 CSoutput.n423 CSoutput.n421 0.573776
R16657 CSoutput.n421 CSoutput.n419 0.573776
R16658 CSoutput.n419 CSoutput.n417 0.573776
R16659 CSoutput.n417 CSoutput.n415 0.573776
R16660 CSoutput.n415 CSoutput.n413 0.573776
R16661 CSoutput.n413 CSoutput.n411 0.573776
R16662 CSoutput.n469 CSoutput.n288 0.53442
R16663 CSoutput.n332 CSoutput.n330 0.358259
R16664 CSoutput.n334 CSoutput.n332 0.358259
R16665 CSoutput.n336 CSoutput.n334 0.358259
R16666 CSoutput.n338 CSoutput.n336 0.358259
R16667 CSoutput.n340 CSoutput.n338 0.358259
R16668 CSoutput.n342 CSoutput.n340 0.358259
R16669 CSoutput.n344 CSoutput.n342 0.358259
R16670 CSoutput.n346 CSoutput.n344 0.358259
R16671 CSoutput.n312 CSoutput.n310 0.358259
R16672 CSoutput.n314 CSoutput.n312 0.358259
R16673 CSoutput.n316 CSoutput.n314 0.358259
R16674 CSoutput.n318 CSoutput.n316 0.358259
R16675 CSoutput.n320 CSoutput.n318 0.358259
R16676 CSoutput.n322 CSoutput.n320 0.358259
R16677 CSoutput.n324 CSoutput.n322 0.358259
R16678 CSoutput.n326 CSoutput.n324 0.358259
R16679 CSoutput.n293 CSoutput.n291 0.358259
R16680 CSoutput.n295 CSoutput.n293 0.358259
R16681 CSoutput.n297 CSoutput.n295 0.358259
R16682 CSoutput.n299 CSoutput.n297 0.358259
R16683 CSoutput.n301 CSoutput.n299 0.358259
R16684 CSoutput.n303 CSoutput.n301 0.358259
R16685 CSoutput.n305 CSoutput.n303 0.358259
R16686 CSoutput.n307 CSoutput.n305 0.358259
R16687 CSoutput.n136 CSoutput.n134 0.358259
R16688 CSoutput.n134 CSoutput.n132 0.358259
R16689 CSoutput.n132 CSoutput.n130 0.358259
R16690 CSoutput.n130 CSoutput.n128 0.358259
R16691 CSoutput.n128 CSoutput.n126 0.358259
R16692 CSoutput.n126 CSoutput.n124 0.358259
R16693 CSoutput.n124 CSoutput.n122 0.358259
R16694 CSoutput.n122 CSoutput.n120 0.358259
R16695 CSoutput.n116 CSoutput.n114 0.358259
R16696 CSoutput.n114 CSoutput.n112 0.358259
R16697 CSoutput.n112 CSoutput.n110 0.358259
R16698 CSoutput.n110 CSoutput.n108 0.358259
R16699 CSoutput.n108 CSoutput.n106 0.358259
R16700 CSoutput.n106 CSoutput.n104 0.358259
R16701 CSoutput.n104 CSoutput.n102 0.358259
R16702 CSoutput.n102 CSoutput.n100 0.358259
R16703 CSoutput.n97 CSoutput.n95 0.358259
R16704 CSoutput.n95 CSoutput.n93 0.358259
R16705 CSoutput.n93 CSoutput.n91 0.358259
R16706 CSoutput.n91 CSoutput.n89 0.358259
R16707 CSoutput.n89 CSoutput.n87 0.358259
R16708 CSoutput.n87 CSoutput.n85 0.358259
R16709 CSoutput.n85 CSoutput.n83 0.358259
R16710 CSoutput.n83 CSoutput.n81 0.358259
R16711 CSoutput.n21 CSoutput.n20 0.169105
R16712 CSoutput.n21 CSoutput.n16 0.169105
R16713 CSoutput.n26 CSoutput.n16 0.169105
R16714 CSoutput.n27 CSoutput.n26 0.169105
R16715 CSoutput.n27 CSoutput.n14 0.169105
R16716 CSoutput.n32 CSoutput.n14 0.169105
R16717 CSoutput.n33 CSoutput.n32 0.169105
R16718 CSoutput.n34 CSoutput.n33 0.169105
R16719 CSoutput.n34 CSoutput.n12 0.169105
R16720 CSoutput.n39 CSoutput.n12 0.169105
R16721 CSoutput.n40 CSoutput.n39 0.169105
R16722 CSoutput.n40 CSoutput.n10 0.169105
R16723 CSoutput.n45 CSoutput.n10 0.169105
R16724 CSoutput.n46 CSoutput.n45 0.169105
R16725 CSoutput.n47 CSoutput.n46 0.169105
R16726 CSoutput.n47 CSoutput.n8 0.169105
R16727 CSoutput.n52 CSoutput.n8 0.169105
R16728 CSoutput.n53 CSoutput.n52 0.169105
R16729 CSoutput.n53 CSoutput.n6 0.169105
R16730 CSoutput.n58 CSoutput.n6 0.169105
R16731 CSoutput.n59 CSoutput.n58 0.169105
R16732 CSoutput.n60 CSoutput.n59 0.169105
R16733 CSoutput.n60 CSoutput.n4 0.169105
R16734 CSoutput.n66 CSoutput.n4 0.169105
R16735 CSoutput.n67 CSoutput.n66 0.169105
R16736 CSoutput.n68 CSoutput.n67 0.169105
R16737 CSoutput.n68 CSoutput.n2 0.169105
R16738 CSoutput.n73 CSoutput.n2 0.169105
R16739 CSoutput.n74 CSoutput.n73 0.169105
R16740 CSoutput.n74 CSoutput.n0 0.169105
R16741 CSoutput.n78 CSoutput.n0 0.169105
R16742 CSoutput.n231 CSoutput.n230 0.0910737
R16743 CSoutput.n282 CSoutput.n279 0.0723685
R16744 CSoutput.n236 CSoutput.n231 0.0522944
R16745 CSoutput.n279 CSoutput.n278 0.0499135
R16746 CSoutput.n230 CSoutput.n229 0.0499135
R16747 CSoutput.n264 CSoutput.n263 0.0464294
R16748 CSoutput.n272 CSoutput.n269 0.0391444
R16749 CSoutput.n231 CSoutput.t240 0.023435
R16750 CSoutput.n279 CSoutput.t243 0.02262
R16751 CSoutput.n230 CSoutput.t246 0.02262
R16752 CSoutput CSoutput.n469 0.0052
R16753 CSoutput.n201 CSoutput.n184 0.00365111
R16754 CSoutput.n204 CSoutput.n185 0.00365111
R16755 CSoutput.n187 CSoutput.n186 0.00365111
R16756 CSoutput.n229 CSoutput.n188 0.00365111
R16757 CSoutput.n193 CSoutput.n189 0.00365111
R16758 CSoutput.n276 CSoutput.n190 0.00365111
R16759 CSoutput.n267 CSoutput.n266 0.00365111
R16760 CSoutput.n247 CSoutput.n220 0.00365111
R16761 CSoutput.n249 CSoutput.n219 0.00365111
R16762 CSoutput.n237 CSoutput.n236 0.00365111
R16763 CSoutput.n243 CSoutput.n223 0.00365111
R16764 CSoutput.n245 CSoutput.n222 0.00365111
R16765 CSoutput.n167 CSoutput.n150 0.00365111
R16766 CSoutput.n170 CSoutput.n151 0.00365111
R16767 CSoutput.n153 CSoutput.n152 0.00365111
R16768 CSoutput.n263 CSoutput.n154 0.00365111
R16769 CSoutput.n159 CSoutput.n155 0.00365111
R16770 CSoutput.n286 CSoutput.n156 0.00365111
R16771 CSoutput.n198 CSoutput.n188 0.00340054
R16772 CSoutput.n191 CSoutput.n189 0.00340054
R16773 CSoutput.n276 CSoutput.n275 0.00340054
R16774 CSoutput.n271 CSoutput.n184 0.00340054
R16775 CSoutput.n200 CSoutput.n185 0.00340054
R16776 CSoutput.n203 CSoutput.n187 0.00340054
R16777 CSoutput.n242 CSoutput.n237 0.00340054
R16778 CSoutput.n244 CSoutput.n243 0.00340054
R16779 CSoutput.n246 CSoutput.n245 0.00340054
R16780 CSoutput.n268 CSoutput.n267 0.00340054
R16781 CSoutput.n248 CSoutput.n247 0.00340054
R16782 CSoutput.n250 CSoutput.n249 0.00340054
R16783 CSoutput.n164 CSoutput.n154 0.00340054
R16784 CSoutput.n157 CSoutput.n155 0.00340054
R16785 CSoutput.n286 CSoutput.n285 0.00340054
R16786 CSoutput.n281 CSoutput.n150 0.00340054
R16787 CSoutput.n166 CSoutput.n151 0.00340054
R16788 CSoutput.n169 CSoutput.n153 0.00340054
R16789 CSoutput.n199 CSoutput.n193 0.00252698
R16790 CSoutput.n192 CSoutput.n190 0.00252698
R16791 CSoutput.n274 CSoutput.n273 0.00252698
R16792 CSoutput.n202 CSoutput.n200 0.00252698
R16793 CSoutput.n205 CSoutput.n203 0.00252698
R16794 CSoutput.n278 CSoutput.n173 0.00252698
R16795 CSoutput.n199 CSoutput.n198 0.00252698
R16796 CSoutput.n192 CSoutput.n191 0.00252698
R16797 CSoutput.n275 CSoutput.n274 0.00252698
R16798 CSoutput.n202 CSoutput.n201 0.00252698
R16799 CSoutput.n205 CSoutput.n204 0.00252698
R16800 CSoutput.n186 CSoutput.n173 0.00252698
R16801 CSoutput.n253 CSoutput.n223 0.00252698
R16802 CSoutput.n252 CSoutput.n222 0.00252698
R16803 CSoutput.n251 CSoutput.n207 0.00252698
R16804 CSoutput.n248 CSoutput.n218 0.00252698
R16805 CSoutput.n255 CSoutput.n250 0.00252698
R16806 CSoutput.n264 CSoutput.n257 0.00252698
R16807 CSoutput.n253 CSoutput.n242 0.00252698
R16808 CSoutput.n252 CSoutput.n244 0.00252698
R16809 CSoutput.n251 CSoutput.n246 0.00252698
R16810 CSoutput.n266 CSoutput.n218 0.00252698
R16811 CSoutput.n255 CSoutput.n220 0.00252698
R16812 CSoutput.n257 CSoutput.n219 0.00252698
R16813 CSoutput.n165 CSoutput.n159 0.00252698
R16814 CSoutput.n158 CSoutput.n156 0.00252698
R16815 CSoutput.n284 CSoutput.n283 0.00252698
R16816 CSoutput.n168 CSoutput.n166 0.00252698
R16817 CSoutput.n171 CSoutput.n169 0.00252698
R16818 CSoutput.n288 CSoutput.n139 0.00252698
R16819 CSoutput.n165 CSoutput.n164 0.00252698
R16820 CSoutput.n158 CSoutput.n157 0.00252698
R16821 CSoutput.n285 CSoutput.n284 0.00252698
R16822 CSoutput.n168 CSoutput.n167 0.00252698
R16823 CSoutput.n171 CSoutput.n170 0.00252698
R16824 CSoutput.n152 CSoutput.n139 0.00252698
R16825 CSoutput.n273 CSoutput.n272 0.0020275
R16826 CSoutput.n272 CSoutput.n271 0.0020275
R16827 CSoutput.n269 CSoutput.n207 0.0020275
R16828 CSoutput.n269 CSoutput.n268 0.0020275
R16829 CSoutput.n283 CSoutput.n282 0.0020275
R16830 CSoutput.n282 CSoutput.n281 0.0020275
R16831 CSoutput.n183 CSoutput.n182 0.00166668
R16832 CSoutput.n265 CSoutput.n221 0.00166668
R16833 CSoutput.n149 CSoutput.n148 0.00166668
R16834 CSoutput.n287 CSoutput.n149 0.00133328
R16835 CSoutput.n221 CSoutput.n217 0.00133328
R16836 CSoutput.n277 CSoutput.n183 0.00133328
R16837 CSoutput.n280 CSoutput.n172 0.001
R16838 CSoutput.n258 CSoutput.n172 0.001
R16839 CSoutput.n160 CSoutput.n140 0.001
R16840 CSoutput.n259 CSoutput.n140 0.001
R16841 CSoutput.n161 CSoutput.n141 0.001
R16842 CSoutput.n260 CSoutput.n141 0.001
R16843 CSoutput.n162 CSoutput.n142 0.001
R16844 CSoutput.n261 CSoutput.n142 0.001
R16845 CSoutput.n163 CSoutput.n143 0.001
R16846 CSoutput.n262 CSoutput.n143 0.001
R16847 CSoutput.n256 CSoutput.n208 0.001
R16848 CSoutput.n256 CSoutput.n254 0.001
R16849 CSoutput.n238 CSoutput.n209 0.001
R16850 CSoutput.n232 CSoutput.n209 0.001
R16851 CSoutput.n239 CSoutput.n210 0.001
R16852 CSoutput.n233 CSoutput.n210 0.001
R16853 CSoutput.n240 CSoutput.n211 0.001
R16854 CSoutput.n234 CSoutput.n211 0.001
R16855 CSoutput.n241 CSoutput.n212 0.001
R16856 CSoutput.n235 CSoutput.n212 0.001
R16857 CSoutput.n270 CSoutput.n206 0.001
R16858 CSoutput.n224 CSoutput.n206 0.001
R16859 CSoutput.n194 CSoutput.n174 0.001
R16860 CSoutput.n225 CSoutput.n174 0.001
R16861 CSoutput.n195 CSoutput.n175 0.001
R16862 CSoutput.n226 CSoutput.n175 0.001
R16863 CSoutput.n196 CSoutput.n176 0.001
R16864 CSoutput.n227 CSoutput.n176 0.001
R16865 CSoutput.n197 CSoutput.n177 0.001
R16866 CSoutput.n228 CSoutput.n177 0.001
R16867 CSoutput.n228 CSoutput.n178 0.001
R16868 CSoutput.n227 CSoutput.n179 0.001
R16869 CSoutput.n226 CSoutput.n180 0.001
R16870 CSoutput.n225 CSoutput.t260 0.001
R16871 CSoutput.n224 CSoutput.n181 0.001
R16872 CSoutput.n197 CSoutput.n179 0.001
R16873 CSoutput.n196 CSoutput.n180 0.001
R16874 CSoutput.n195 CSoutput.t260 0.001
R16875 CSoutput.n194 CSoutput.n181 0.001
R16876 CSoutput.n270 CSoutput.n182 0.001
R16877 CSoutput.n235 CSoutput.n213 0.001
R16878 CSoutput.n234 CSoutput.n214 0.001
R16879 CSoutput.n233 CSoutput.n215 0.001
R16880 CSoutput.n232 CSoutput.t256 0.001
R16881 CSoutput.n254 CSoutput.n216 0.001
R16882 CSoutput.n241 CSoutput.n214 0.001
R16883 CSoutput.n240 CSoutput.n215 0.001
R16884 CSoutput.n239 CSoutput.t256 0.001
R16885 CSoutput.n238 CSoutput.n216 0.001
R16886 CSoutput.n265 CSoutput.n208 0.001
R16887 CSoutput.n262 CSoutput.n144 0.001
R16888 CSoutput.n261 CSoutput.n145 0.001
R16889 CSoutput.n260 CSoutput.n146 0.001
R16890 CSoutput.n259 CSoutput.t255 0.001
R16891 CSoutput.n258 CSoutput.n147 0.001
R16892 CSoutput.n163 CSoutput.n145 0.001
R16893 CSoutput.n162 CSoutput.n146 0.001
R16894 CSoutput.n161 CSoutput.t255 0.001
R16895 CSoutput.n160 CSoutput.n147 0.001
R16896 CSoutput.n280 CSoutput.n148 0.001
R16897 a_n1986_13878.n3 a_n1986_13878.t11 539.01
R16898 a_n1986_13878.n90 a_n1986_13878.t13 512.366
R16899 a_n1986_13878.n89 a_n1986_13878.t33 512.366
R16900 a_n1986_13878.n51 a_n1986_13878.t17 512.366
R16901 a_n1986_13878.n88 a_n1986_13878.t29 512.366
R16902 a_n1986_13878.n7 a_n1986_13878.t67 539.01
R16903 a_n1986_13878.n79 a_n1986_13878.t50 512.366
R16904 a_n1986_13878.n78 a_n1986_13878.t54 512.366
R16905 a_n1986_13878.n52 a_n1986_13878.t44 512.366
R16906 a_n1986_13878.n77 a_n1986_13878.t59 512.366
R16907 a_n1986_13878.n20 a_n1986_13878.t27 539.01
R16908 a_n1986_13878.n60 a_n1986_13878.t21 512.366
R16909 a_n1986_13878.n61 a_n1986_13878.t23 512.366
R16910 a_n1986_13878.n55 a_n1986_13878.t15 512.366
R16911 a_n1986_13878.n62 a_n1986_13878.t25 512.366
R16912 a_n1986_13878.n24 a_n1986_13878.t62 539.01
R16913 a_n1986_13878.n57 a_n1986_13878.t63 512.366
R16914 a_n1986_13878.n58 a_n1986_13878.t42 512.366
R16915 a_n1986_13878.n56 a_n1986_13878.t48 512.366
R16916 a_n1986_13878.n59 a_n1986_13878.t57 512.366
R16917 a_n1986_13878.n74 a_n1986_13878.t56 512.366
R16918 a_n1986_13878.n64 a_n1986_13878.t47 512.366
R16919 a_n1986_13878.n75 a_n1986_13878.t41 512.366
R16920 a_n1986_13878.n72 a_n1986_13878.t64 512.366
R16921 a_n1986_13878.n65 a_n1986_13878.t53 512.366
R16922 a_n1986_13878.n73 a_n1986_13878.t52 512.366
R16923 a_n1986_13878.n70 a_n1986_13878.t60 512.366
R16924 a_n1986_13878.n66 a_n1986_13878.t45 512.366
R16925 a_n1986_13878.n71 a_n1986_13878.t46 512.366
R16926 a_n1986_13878.n68 a_n1986_13878.t49 512.366
R16927 a_n1986_13878.n67 a_n1986_13878.t58 512.366
R16928 a_n1986_13878.n69 a_n1986_13878.t40 512.366
R16929 a_n1986_13878.n50 a_n1986_13878.n0 70.3058
R16930 a_n1986_13878.n47 a_n1986_13878.n5 70.3058
R16931 a_n1986_13878.n17 a_n1986_13878.n36 70.3058
R16932 a_n1986_13878.n21 a_n1986_13878.n33 70.3058
R16933 a_n1986_13878.n32 a_n1986_13878.n22 70.1674
R16934 a_n1986_13878.n32 a_n1986_13878.n56 20.9683
R16935 a_n1986_13878.n22 a_n1986_13878.n31 75.0448
R16936 a_n1986_13878.n58 a_n1986_13878.n31 11.2134
R16937 a_n1986_13878.n23 a_n1986_13878.n24 44.8194
R16938 a_n1986_13878.n35 a_n1986_13878.n18 70.1674
R16939 a_n1986_13878.n35 a_n1986_13878.n55 20.9683
R16940 a_n1986_13878.n18 a_n1986_13878.n34 75.0448
R16941 a_n1986_13878.n61 a_n1986_13878.n34 11.2134
R16942 a_n1986_13878.n19 a_n1986_13878.n20 44.8194
R16943 a_n1986_13878.n8 a_n1986_13878.n44 70.1674
R16944 a_n1986_13878.n10 a_n1986_13878.n42 70.1674
R16945 a_n1986_13878.n12 a_n1986_13878.n40 70.1674
R16946 a_n1986_13878.n15 a_n1986_13878.n38 70.1674
R16947 a_n1986_13878.n69 a_n1986_13878.n38 20.9683
R16948 a_n1986_13878.n37 a_n1986_13878.n16 75.0448
R16949 a_n1986_13878.n37 a_n1986_13878.n67 11.2134
R16950 a_n1986_13878.n16 a_n1986_13878.n68 161.3
R16951 a_n1986_13878.n71 a_n1986_13878.n40 20.9683
R16952 a_n1986_13878.n39 a_n1986_13878.n13 75.0448
R16953 a_n1986_13878.n39 a_n1986_13878.n66 11.2134
R16954 a_n1986_13878.n13 a_n1986_13878.n70 161.3
R16955 a_n1986_13878.n73 a_n1986_13878.n42 20.9683
R16956 a_n1986_13878.n41 a_n1986_13878.n11 75.0448
R16957 a_n1986_13878.n41 a_n1986_13878.n65 11.2134
R16958 a_n1986_13878.n11 a_n1986_13878.n72 161.3
R16959 a_n1986_13878.n75 a_n1986_13878.n44 20.9683
R16960 a_n1986_13878.n43 a_n1986_13878.n9 75.0448
R16961 a_n1986_13878.n43 a_n1986_13878.n64 11.2134
R16962 a_n1986_13878.n9 a_n1986_13878.n74 161.3
R16963 a_n1986_13878.n6 a_n1986_13878.n46 70.1674
R16964 a_n1986_13878.n46 a_n1986_13878.n52 20.9683
R16965 a_n1986_13878.n45 a_n1986_13878.n6 75.0448
R16966 a_n1986_13878.n78 a_n1986_13878.n45 11.2134
R16967 a_n1986_13878.n4 a_n1986_13878.n7 44.8194
R16968 a_n1986_13878.n2 a_n1986_13878.n49 70.1674
R16969 a_n1986_13878.n49 a_n1986_13878.n51 20.9683
R16970 a_n1986_13878.n48 a_n1986_13878.n2 75.0448
R16971 a_n1986_13878.n89 a_n1986_13878.n48 11.2134
R16972 a_n1986_13878.n1 a_n1986_13878.n3 44.8194
R16973 a_n1986_13878.n29 a_n1986_13878.n86 81.2902
R16974 a_n1986_13878.n30 a_n1986_13878.n82 81.2902
R16975 a_n1986_13878.n30 a_n1986_13878.n80 81.2902
R16976 a_n1986_13878.n29 a_n1986_13878.n87 80.9324
R16977 a_n1986_13878.n29 a_n1986_13878.n85 80.9324
R16978 a_n1986_13878.n28 a_n1986_13878.n84 80.9324
R16979 a_n1986_13878.n30 a_n1986_13878.n83 80.9324
R16980 a_n1986_13878.n30 a_n1986_13878.n81 80.9324
R16981 a_n1986_13878.n27 a_n1986_13878.t20 74.6477
R16982 a_n1986_13878.n25 a_n1986_13878.t28 74.6477
R16983 a_n1986_13878.t12 a_n1986_13878.n94 74.2899
R16984 a_n1986_13878.n26 a_n1986_13878.t32 74.2897
R16985 a_n1986_13878.n27 a_n1986_13878.n92 70.6783
R16986 a_n1986_13878.n27 a_n1986_13878.n93 70.6783
R16987 a_n1986_13878.n26 a_n1986_13878.n54 70.6783
R16988 a_n1986_13878.n25 a_n1986_13878.n53 70.6783
R16989 a_n1986_13878.n90 a_n1986_13878.n89 48.2005
R16990 a_n1986_13878.n88 a_n1986_13878.n49 20.9683
R16991 a_n1986_13878.n79 a_n1986_13878.n78 48.2005
R16992 a_n1986_13878.n77 a_n1986_13878.n46 20.9683
R16993 a_n1986_13878.n61 a_n1986_13878.n60 48.2005
R16994 a_n1986_13878.n62 a_n1986_13878.n35 20.9683
R16995 a_n1986_13878.n58 a_n1986_13878.n57 48.2005
R16996 a_n1986_13878.n59 a_n1986_13878.n32 20.9683
R16997 a_n1986_13878.n74 a_n1986_13878.n64 48.2005
R16998 a_n1986_13878.t61 a_n1986_13878.n44 533.335
R16999 a_n1986_13878.n72 a_n1986_13878.n65 48.2005
R17000 a_n1986_13878.t66 a_n1986_13878.n42 533.335
R17001 a_n1986_13878.n70 a_n1986_13878.n66 48.2005
R17002 a_n1986_13878.t55 a_n1986_13878.n40 533.335
R17003 a_n1986_13878.n68 a_n1986_13878.n67 48.2005
R17004 a_n1986_13878.t51 a_n1986_13878.n38 533.335
R17005 a_n1986_13878.n50 a_n1986_13878.t19 533.058
R17006 a_n1986_13878.n47 a_n1986_13878.t65 533.058
R17007 a_n1986_13878.t31 a_n1986_13878.n36 533.058
R17008 a_n1986_13878.t43 a_n1986_13878.n33 533.058
R17009 a_n1986_13878.n48 a_n1986_13878.n51 35.3134
R17010 a_n1986_13878.n45 a_n1986_13878.n52 35.3134
R17011 a_n1986_13878.n55 a_n1986_13878.n34 35.3134
R17012 a_n1986_13878.n56 a_n1986_13878.n31 35.3134
R17013 a_n1986_13878.n75 a_n1986_13878.n43 35.3134
R17014 a_n1986_13878.n73 a_n1986_13878.n41 35.3134
R17015 a_n1986_13878.n71 a_n1986_13878.n39 35.3134
R17016 a_n1986_13878.n69 a_n1986_13878.n37 35.3134
R17017 a_n1986_13878.n28 a_n1986_13878.n30 31.0592
R17018 a_n1986_13878.n0 a_n1986_13878.n29 23.891
R17019 a_n1986_13878.n23 a_n1986_13878.n14 12.046
R17020 a_n1986_13878.n5 a_n1986_13878.n76 11.8414
R17021 a_n1986_13878.n91 a_n1986_13878.n1 10.5365
R17022 a_n1986_13878.n63 a_n1986_13878.n26 9.50122
R17023 a_n1986_13878.n16 a_n1986_13878.n14 7.47588
R17024 a_n1986_13878.n76 a_n1986_13878.n8 7.47588
R17025 a_n1986_13878.n63 a_n1986_13878.n17 6.70126
R17026 a_n1986_13878.n94 a_n1986_13878.n91 5.65783
R17027 a_n1986_13878.n76 a_n1986_13878.n63 5.3452
R17028 a_n1986_13878.n19 a_n1986_13878.n21 3.95126
R17029 a_n1986_13878.n92 a_n1986_13878.t18 3.61217
R17030 a_n1986_13878.n92 a_n1986_13878.t30 3.61217
R17031 a_n1986_13878.n93 a_n1986_13878.t14 3.61217
R17032 a_n1986_13878.n93 a_n1986_13878.t34 3.61217
R17033 a_n1986_13878.n54 a_n1986_13878.t16 3.61217
R17034 a_n1986_13878.n54 a_n1986_13878.t26 3.61217
R17035 a_n1986_13878.n53 a_n1986_13878.t22 3.61217
R17036 a_n1986_13878.n53 a_n1986_13878.t24 3.61217
R17037 a_n1986_13878.n0 a_n1986_13878.n4 3.42095
R17038 a_n1986_13878.n86 a_n1986_13878.t0 2.82907
R17039 a_n1986_13878.n86 a_n1986_13878.t39 2.82907
R17040 a_n1986_13878.n87 a_n1986_13878.t4 2.82907
R17041 a_n1986_13878.n87 a_n1986_13878.t6 2.82907
R17042 a_n1986_13878.n85 a_n1986_13878.t37 2.82907
R17043 a_n1986_13878.n85 a_n1986_13878.t7 2.82907
R17044 a_n1986_13878.n84 a_n1986_13878.t8 2.82907
R17045 a_n1986_13878.n84 a_n1986_13878.t38 2.82907
R17046 a_n1986_13878.n82 a_n1986_13878.t2 2.82907
R17047 a_n1986_13878.n82 a_n1986_13878.t36 2.82907
R17048 a_n1986_13878.n83 a_n1986_13878.t3 2.82907
R17049 a_n1986_13878.n83 a_n1986_13878.t10 2.82907
R17050 a_n1986_13878.n81 a_n1986_13878.t35 2.82907
R17051 a_n1986_13878.n81 a_n1986_13878.t1 2.82907
R17052 a_n1986_13878.n80 a_n1986_13878.t9 2.82907
R17053 a_n1986_13878.n80 a_n1986_13878.t5 2.82907
R17054 a_n1986_13878.n91 a_n1986_13878.n14 1.30542
R17055 a_n1986_13878.n11 a_n1986_13878.n12 1.04595
R17056 a_n1986_13878.n3 a_n1986_13878.n90 13.657
R17057 a_n1986_13878.n88 a_n1986_13878.n50 21.4216
R17058 a_n1986_13878.n7 a_n1986_13878.n79 13.657
R17059 a_n1986_13878.n77 a_n1986_13878.n47 21.4216
R17060 a_n1986_13878.n60 a_n1986_13878.n20 13.657
R17061 a_n1986_13878.n36 a_n1986_13878.n62 21.4216
R17062 a_n1986_13878.n57 a_n1986_13878.n24 13.657
R17063 a_n1986_13878.n33 a_n1986_13878.n59 21.4216
R17064 a_n1986_13878.n2 a_n1986_13878.n0 1.2505
R17065 a_n1986_13878.n23 a_n1986_13878.n22 0.758076
R17066 a_n1986_13878.n22 a_n1986_13878.n21 0.758076
R17067 a_n1986_13878.n19 a_n1986_13878.n18 0.758076
R17068 a_n1986_13878.n18 a_n1986_13878.n17 0.758076
R17069 a_n1986_13878.n16 a_n1986_13878.n15 0.758076
R17070 a_n1986_13878.n13 a_n1986_13878.n12 0.758076
R17071 a_n1986_13878.n11 a_n1986_13878.n10 0.758076
R17072 a_n1986_13878.n9 a_n1986_13878.n8 0.758076
R17073 a_n1986_13878.n6 a_n1986_13878.n4 0.758076
R17074 a_n1986_13878.n6 a_n1986_13878.n5 0.758076
R17075 a_n1986_13878.n2 a_n1986_13878.n1 0.758076
R17076 a_n1986_13878.n29 a_n1986_13878.n28 0.716017
R17077 a_n1986_13878.n94 a_n1986_13878.n27 0.716017
R17078 a_n1986_13878.n26 a_n1986_13878.n25 0.716017
R17079 a_n1986_13878.n13 a_n1986_13878.n15 0.67853
R17080 a_n1986_13878.n9 a_n1986_13878.n10 0.67853
R17081 vdd.n327 vdd.n291 756.745
R17082 vdd.n268 vdd.n232 756.745
R17083 vdd.n225 vdd.n189 756.745
R17084 vdd.n166 vdd.n130 756.745
R17085 vdd.n124 vdd.n88 756.745
R17086 vdd.n65 vdd.n29 756.745
R17087 vdd.n1746 vdd.n1710 756.745
R17088 vdd.n1805 vdd.n1769 756.745
R17089 vdd.n1644 vdd.n1608 756.745
R17090 vdd.n1703 vdd.n1667 756.745
R17091 vdd.n1543 vdd.n1507 756.745
R17092 vdd.n1602 vdd.n1566 756.745
R17093 vdd.n2177 vdd.t219 640.208
R17094 vdd.n965 vdd.t204 640.208
R17095 vdd.n2151 vdd.t242 640.208
R17096 vdd.n957 vdd.t230 640.208
R17097 vdd.n2922 vdd.t180 640.208
R17098 vdd.n2642 vdd.t227 640.208
R17099 vdd.n832 vdd.t208 640.208
R17100 vdd.n2639 vdd.t212 640.208
R17101 vdd.n799 vdd.t216 640.208
R17102 vdd.n1027 vdd.t223 640.208
R17103 vdd.n1317 vdd.t195 592.009
R17104 vdd.n1355 vdd.t184 592.009
R17105 vdd.n1251 vdd.t198 592.009
R17106 vdd.n2333 vdd.t176 592.009
R17107 vdd.n1970 vdd.t188 592.009
R17108 vdd.n1930 vdd.t201 592.009
R17109 vdd.n426 vdd.t191 592.009
R17110 vdd.n440 vdd.t233 592.009
R17111 vdd.n452 vdd.t239 592.009
R17112 vdd.n768 vdd.t169 592.009
R17113 vdd.n3184 vdd.t173 592.009
R17114 vdd.n688 vdd.t236 592.009
R17115 vdd.n328 vdd.n327 585
R17116 vdd.n326 vdd.n293 585
R17117 vdd.n325 vdd.n324 585
R17118 vdd.n296 vdd.n294 585
R17119 vdd.n319 vdd.n318 585
R17120 vdd.n317 vdd.n316 585
R17121 vdd.n300 vdd.n299 585
R17122 vdd.n311 vdd.n310 585
R17123 vdd.n309 vdd.n308 585
R17124 vdd.n304 vdd.n303 585
R17125 vdd.n269 vdd.n268 585
R17126 vdd.n267 vdd.n234 585
R17127 vdd.n266 vdd.n265 585
R17128 vdd.n237 vdd.n235 585
R17129 vdd.n260 vdd.n259 585
R17130 vdd.n258 vdd.n257 585
R17131 vdd.n241 vdd.n240 585
R17132 vdd.n252 vdd.n251 585
R17133 vdd.n250 vdd.n249 585
R17134 vdd.n245 vdd.n244 585
R17135 vdd.n226 vdd.n225 585
R17136 vdd.n224 vdd.n191 585
R17137 vdd.n223 vdd.n222 585
R17138 vdd.n194 vdd.n192 585
R17139 vdd.n217 vdd.n216 585
R17140 vdd.n215 vdd.n214 585
R17141 vdd.n198 vdd.n197 585
R17142 vdd.n209 vdd.n208 585
R17143 vdd.n207 vdd.n206 585
R17144 vdd.n202 vdd.n201 585
R17145 vdd.n167 vdd.n166 585
R17146 vdd.n165 vdd.n132 585
R17147 vdd.n164 vdd.n163 585
R17148 vdd.n135 vdd.n133 585
R17149 vdd.n158 vdd.n157 585
R17150 vdd.n156 vdd.n155 585
R17151 vdd.n139 vdd.n138 585
R17152 vdd.n150 vdd.n149 585
R17153 vdd.n148 vdd.n147 585
R17154 vdd.n143 vdd.n142 585
R17155 vdd.n125 vdd.n124 585
R17156 vdd.n123 vdd.n90 585
R17157 vdd.n122 vdd.n121 585
R17158 vdd.n93 vdd.n91 585
R17159 vdd.n116 vdd.n115 585
R17160 vdd.n114 vdd.n113 585
R17161 vdd.n97 vdd.n96 585
R17162 vdd.n108 vdd.n107 585
R17163 vdd.n106 vdd.n105 585
R17164 vdd.n101 vdd.n100 585
R17165 vdd.n66 vdd.n65 585
R17166 vdd.n64 vdd.n31 585
R17167 vdd.n63 vdd.n62 585
R17168 vdd.n34 vdd.n32 585
R17169 vdd.n57 vdd.n56 585
R17170 vdd.n55 vdd.n54 585
R17171 vdd.n38 vdd.n37 585
R17172 vdd.n49 vdd.n48 585
R17173 vdd.n47 vdd.n46 585
R17174 vdd.n42 vdd.n41 585
R17175 vdd.n1747 vdd.n1746 585
R17176 vdd.n1745 vdd.n1712 585
R17177 vdd.n1744 vdd.n1743 585
R17178 vdd.n1715 vdd.n1713 585
R17179 vdd.n1738 vdd.n1737 585
R17180 vdd.n1736 vdd.n1735 585
R17181 vdd.n1719 vdd.n1718 585
R17182 vdd.n1730 vdd.n1729 585
R17183 vdd.n1728 vdd.n1727 585
R17184 vdd.n1723 vdd.n1722 585
R17185 vdd.n1806 vdd.n1805 585
R17186 vdd.n1804 vdd.n1771 585
R17187 vdd.n1803 vdd.n1802 585
R17188 vdd.n1774 vdd.n1772 585
R17189 vdd.n1797 vdd.n1796 585
R17190 vdd.n1795 vdd.n1794 585
R17191 vdd.n1778 vdd.n1777 585
R17192 vdd.n1789 vdd.n1788 585
R17193 vdd.n1787 vdd.n1786 585
R17194 vdd.n1782 vdd.n1781 585
R17195 vdd.n1645 vdd.n1644 585
R17196 vdd.n1643 vdd.n1610 585
R17197 vdd.n1642 vdd.n1641 585
R17198 vdd.n1613 vdd.n1611 585
R17199 vdd.n1636 vdd.n1635 585
R17200 vdd.n1634 vdd.n1633 585
R17201 vdd.n1617 vdd.n1616 585
R17202 vdd.n1628 vdd.n1627 585
R17203 vdd.n1626 vdd.n1625 585
R17204 vdd.n1621 vdd.n1620 585
R17205 vdd.n1704 vdd.n1703 585
R17206 vdd.n1702 vdd.n1669 585
R17207 vdd.n1701 vdd.n1700 585
R17208 vdd.n1672 vdd.n1670 585
R17209 vdd.n1695 vdd.n1694 585
R17210 vdd.n1693 vdd.n1692 585
R17211 vdd.n1676 vdd.n1675 585
R17212 vdd.n1687 vdd.n1686 585
R17213 vdd.n1685 vdd.n1684 585
R17214 vdd.n1680 vdd.n1679 585
R17215 vdd.n1544 vdd.n1543 585
R17216 vdd.n1542 vdd.n1509 585
R17217 vdd.n1541 vdd.n1540 585
R17218 vdd.n1512 vdd.n1510 585
R17219 vdd.n1535 vdd.n1534 585
R17220 vdd.n1533 vdd.n1532 585
R17221 vdd.n1516 vdd.n1515 585
R17222 vdd.n1527 vdd.n1526 585
R17223 vdd.n1525 vdd.n1524 585
R17224 vdd.n1520 vdd.n1519 585
R17225 vdd.n1603 vdd.n1602 585
R17226 vdd.n1601 vdd.n1568 585
R17227 vdd.n1600 vdd.n1599 585
R17228 vdd.n1571 vdd.n1569 585
R17229 vdd.n1594 vdd.n1593 585
R17230 vdd.n1592 vdd.n1591 585
R17231 vdd.n1575 vdd.n1574 585
R17232 vdd.n1586 vdd.n1585 585
R17233 vdd.n1584 vdd.n1583 585
R17234 vdd.n1579 vdd.n1578 585
R17235 vdd.n3356 vdd.n392 509.269
R17236 vdd.n3352 vdd.n393 509.269
R17237 vdd.n3224 vdd.n685 509.269
R17238 vdd.n3221 vdd.n684 509.269
R17239 vdd.n2328 vdd.n1075 509.269
R17240 vdd.n2331 vdd.n2330 509.269
R17241 vdd.n1224 vdd.n1188 509.269
R17242 vdd.n1420 vdd.n1189 509.269
R17243 vdd.n305 vdd.t115 329.043
R17244 vdd.n246 vdd.t122 329.043
R17245 vdd.n203 vdd.t112 329.043
R17246 vdd.n144 vdd.t108 329.043
R17247 vdd.n102 vdd.t269 329.043
R17248 vdd.n43 vdd.t251 329.043
R17249 vdd.n1724 vdd.t56 329.043
R17250 vdd.n1783 vdd.t59 329.043
R17251 vdd.n1622 vdd.t247 329.043
R17252 vdd.n1681 vdd.t283 329.043
R17253 vdd.n1521 vdd.t44 329.043
R17254 vdd.n1580 vdd.t101 329.043
R17255 vdd.n1317 vdd.t197 319.788
R17256 vdd.n1355 vdd.t187 319.788
R17257 vdd.n1251 vdd.t200 319.788
R17258 vdd.n2333 vdd.t178 319.788
R17259 vdd.n1970 vdd.t189 319.788
R17260 vdd.n1930 vdd.t202 319.788
R17261 vdd.n426 vdd.t193 319.788
R17262 vdd.n440 vdd.t234 319.788
R17263 vdd.n452 vdd.t240 319.788
R17264 vdd.n768 vdd.t172 319.788
R17265 vdd.n3184 vdd.t175 319.788
R17266 vdd.n688 vdd.t238 319.788
R17267 vdd.n1318 vdd.t196 303.69
R17268 vdd.n1356 vdd.t186 303.69
R17269 vdd.n1252 vdd.t199 303.69
R17270 vdd.n2334 vdd.t179 303.69
R17271 vdd.n1971 vdd.t190 303.69
R17272 vdd.n1931 vdd.t203 303.69
R17273 vdd.n427 vdd.t194 303.69
R17274 vdd.n441 vdd.t235 303.69
R17275 vdd.n453 vdd.t241 303.69
R17276 vdd.n769 vdd.t171 303.69
R17277 vdd.n3185 vdd.t174 303.69
R17278 vdd.n689 vdd.t237 303.69
R17279 vdd.n2865 vdd.n913 297.074
R17280 vdd.n3058 vdd.n809 297.074
R17281 vdd.n2995 vdd.n806 297.074
R17282 vdd.n2788 vdd.n914 297.074
R17283 vdd.n2603 vdd.n954 297.074
R17284 vdd.n2534 vdd.n2533 297.074
R17285 vdd.n2280 vdd.n1050 297.074
R17286 vdd.n2376 vdd.n1048 297.074
R17287 vdd.n2974 vdd.n807 297.074
R17288 vdd.n3061 vdd.n3060 297.074
R17289 vdd.n2637 vdd.n915 297.074
R17290 vdd.n2863 vdd.n916 297.074
R17291 vdd.n2531 vdd.n963 297.074
R17292 vdd.n961 vdd.n936 297.074
R17293 vdd.n2217 vdd.n1051 297.074
R17294 vdd.n2374 vdd.n1052 297.074
R17295 vdd.n2976 vdd.n807 185
R17296 vdd.n3059 vdd.n807 185
R17297 vdd.n2978 vdd.n2977 185
R17298 vdd.n2977 vdd.n805 185
R17299 vdd.n2979 vdd.n839 185
R17300 vdd.n2989 vdd.n839 185
R17301 vdd.n2980 vdd.n848 185
R17302 vdd.n848 vdd.n846 185
R17303 vdd.n2982 vdd.n2981 185
R17304 vdd.n2983 vdd.n2982 185
R17305 vdd.n2935 vdd.n847 185
R17306 vdd.n847 vdd.n843 185
R17307 vdd.n2934 vdd.n2933 185
R17308 vdd.n2933 vdd.n2932 185
R17309 vdd.n850 vdd.n849 185
R17310 vdd.n851 vdd.n850 185
R17311 vdd.n2925 vdd.n2924 185
R17312 vdd.n2926 vdd.n2925 185
R17313 vdd.n2921 vdd.n860 185
R17314 vdd.n860 vdd.n857 185
R17315 vdd.n2920 vdd.n2919 185
R17316 vdd.n2919 vdd.n2918 185
R17317 vdd.n862 vdd.n861 185
R17318 vdd.n870 vdd.n862 185
R17319 vdd.n2911 vdd.n2910 185
R17320 vdd.n2912 vdd.n2911 185
R17321 vdd.n2909 vdd.n871 185
R17322 vdd.n2760 vdd.n871 185
R17323 vdd.n2908 vdd.n2907 185
R17324 vdd.n2907 vdd.n2906 185
R17325 vdd.n873 vdd.n872 185
R17326 vdd.n874 vdd.n873 185
R17327 vdd.n2899 vdd.n2898 185
R17328 vdd.n2900 vdd.n2899 185
R17329 vdd.n2897 vdd.n883 185
R17330 vdd.n883 vdd.n880 185
R17331 vdd.n2896 vdd.n2895 185
R17332 vdd.n2895 vdd.n2894 185
R17333 vdd.n885 vdd.n884 185
R17334 vdd.n893 vdd.n885 185
R17335 vdd.n2887 vdd.n2886 185
R17336 vdd.n2888 vdd.n2887 185
R17337 vdd.n2885 vdd.n894 185
R17338 vdd.n900 vdd.n894 185
R17339 vdd.n2884 vdd.n2883 185
R17340 vdd.n2883 vdd.n2882 185
R17341 vdd.n896 vdd.n895 185
R17342 vdd.n897 vdd.n896 185
R17343 vdd.n2875 vdd.n2874 185
R17344 vdd.n2876 vdd.n2875 185
R17345 vdd.n2873 vdd.n906 185
R17346 vdd.n2781 vdd.n906 185
R17347 vdd.n2872 vdd.n2871 185
R17348 vdd.n2871 vdd.n2870 185
R17349 vdd.n908 vdd.n907 185
R17350 vdd.t147 vdd.n908 185
R17351 vdd.n2863 vdd.n2862 185
R17352 vdd.n2864 vdd.n2863 185
R17353 vdd.n2861 vdd.n916 185
R17354 vdd.n2860 vdd.n2859 185
R17355 vdd.n918 vdd.n917 185
R17356 vdd.n2646 vdd.n2645 185
R17357 vdd.n2648 vdd.n2647 185
R17358 vdd.n2650 vdd.n2649 185
R17359 vdd.n2652 vdd.n2651 185
R17360 vdd.n2654 vdd.n2653 185
R17361 vdd.n2656 vdd.n2655 185
R17362 vdd.n2658 vdd.n2657 185
R17363 vdd.n2660 vdd.n2659 185
R17364 vdd.n2662 vdd.n2661 185
R17365 vdd.n2664 vdd.n2663 185
R17366 vdd.n2666 vdd.n2665 185
R17367 vdd.n2668 vdd.n2667 185
R17368 vdd.n2670 vdd.n2669 185
R17369 vdd.n2672 vdd.n2671 185
R17370 vdd.n2674 vdd.n2673 185
R17371 vdd.n2676 vdd.n2675 185
R17372 vdd.n2678 vdd.n2677 185
R17373 vdd.n2680 vdd.n2679 185
R17374 vdd.n2682 vdd.n2681 185
R17375 vdd.n2684 vdd.n2683 185
R17376 vdd.n2686 vdd.n2685 185
R17377 vdd.n2688 vdd.n2687 185
R17378 vdd.n2690 vdd.n2689 185
R17379 vdd.n2692 vdd.n2691 185
R17380 vdd.n2694 vdd.n2693 185
R17381 vdd.n2696 vdd.n2695 185
R17382 vdd.n2698 vdd.n2697 185
R17383 vdd.n2700 vdd.n2699 185
R17384 vdd.n2702 vdd.n2701 185
R17385 vdd.n2704 vdd.n2703 185
R17386 vdd.n2706 vdd.n2705 185
R17387 vdd.n2707 vdd.n2637 185
R17388 vdd.n2857 vdd.n2637 185
R17389 vdd.n3062 vdd.n3061 185
R17390 vdd.n3063 vdd.n798 185
R17391 vdd.n3065 vdd.n3064 185
R17392 vdd.n3067 vdd.n796 185
R17393 vdd.n3069 vdd.n3068 185
R17394 vdd.n3070 vdd.n795 185
R17395 vdd.n3072 vdd.n3071 185
R17396 vdd.n3074 vdd.n793 185
R17397 vdd.n3076 vdd.n3075 185
R17398 vdd.n3077 vdd.n792 185
R17399 vdd.n3079 vdd.n3078 185
R17400 vdd.n3081 vdd.n790 185
R17401 vdd.n3083 vdd.n3082 185
R17402 vdd.n3084 vdd.n789 185
R17403 vdd.n3086 vdd.n3085 185
R17404 vdd.n3088 vdd.n788 185
R17405 vdd.n3089 vdd.n786 185
R17406 vdd.n3092 vdd.n3091 185
R17407 vdd.n787 vdd.n785 185
R17408 vdd.n2948 vdd.n2947 185
R17409 vdd.n2950 vdd.n2949 185
R17410 vdd.n2952 vdd.n2944 185
R17411 vdd.n2954 vdd.n2953 185
R17412 vdd.n2955 vdd.n2943 185
R17413 vdd.n2957 vdd.n2956 185
R17414 vdd.n2959 vdd.n2941 185
R17415 vdd.n2961 vdd.n2960 185
R17416 vdd.n2962 vdd.n2940 185
R17417 vdd.n2964 vdd.n2963 185
R17418 vdd.n2966 vdd.n2938 185
R17419 vdd.n2968 vdd.n2967 185
R17420 vdd.n2969 vdd.n2937 185
R17421 vdd.n2971 vdd.n2970 185
R17422 vdd.n2973 vdd.n2936 185
R17423 vdd.n2975 vdd.n2974 185
R17424 vdd.n2974 vdd.n692 185
R17425 vdd.n3060 vdd.n802 185
R17426 vdd.n3060 vdd.n3059 185
R17427 vdd.n2712 vdd.n804 185
R17428 vdd.n805 vdd.n804 185
R17429 vdd.n2713 vdd.n838 185
R17430 vdd.n2989 vdd.n838 185
R17431 vdd.n2715 vdd.n2714 185
R17432 vdd.n2714 vdd.n846 185
R17433 vdd.n2716 vdd.n845 185
R17434 vdd.n2983 vdd.n845 185
R17435 vdd.n2718 vdd.n2717 185
R17436 vdd.n2717 vdd.n843 185
R17437 vdd.n2719 vdd.n853 185
R17438 vdd.n2932 vdd.n853 185
R17439 vdd.n2721 vdd.n2720 185
R17440 vdd.n2720 vdd.n851 185
R17441 vdd.n2722 vdd.n859 185
R17442 vdd.n2926 vdd.n859 185
R17443 vdd.n2724 vdd.n2723 185
R17444 vdd.n2723 vdd.n857 185
R17445 vdd.n2725 vdd.n864 185
R17446 vdd.n2918 vdd.n864 185
R17447 vdd.n2727 vdd.n2726 185
R17448 vdd.n2726 vdd.n870 185
R17449 vdd.n2728 vdd.n869 185
R17450 vdd.n2912 vdd.n869 185
R17451 vdd.n2762 vdd.n2761 185
R17452 vdd.n2761 vdd.n2760 185
R17453 vdd.n2763 vdd.n876 185
R17454 vdd.n2906 vdd.n876 185
R17455 vdd.n2765 vdd.n2764 185
R17456 vdd.n2764 vdd.n874 185
R17457 vdd.n2766 vdd.n882 185
R17458 vdd.n2900 vdd.n882 185
R17459 vdd.n2768 vdd.n2767 185
R17460 vdd.n2767 vdd.n880 185
R17461 vdd.n2769 vdd.n887 185
R17462 vdd.n2894 vdd.n887 185
R17463 vdd.n2771 vdd.n2770 185
R17464 vdd.n2770 vdd.n893 185
R17465 vdd.n2772 vdd.n892 185
R17466 vdd.n2888 vdd.n892 185
R17467 vdd.n2774 vdd.n2773 185
R17468 vdd.n2773 vdd.n900 185
R17469 vdd.n2775 vdd.n899 185
R17470 vdd.n2882 vdd.n899 185
R17471 vdd.n2777 vdd.n2776 185
R17472 vdd.n2776 vdd.n897 185
R17473 vdd.n2778 vdd.n905 185
R17474 vdd.n2876 vdd.n905 185
R17475 vdd.n2780 vdd.n2779 185
R17476 vdd.n2781 vdd.n2780 185
R17477 vdd.n2711 vdd.n910 185
R17478 vdd.n2870 vdd.n910 185
R17479 vdd.n2710 vdd.n2709 185
R17480 vdd.n2709 vdd.t147 185
R17481 vdd.n2708 vdd.n915 185
R17482 vdd.n2864 vdd.n915 185
R17483 vdd.n2328 vdd.n2327 185
R17484 vdd.n2329 vdd.n2328 185
R17485 vdd.n1076 vdd.n1074 185
R17486 vdd.n1894 vdd.n1074 185
R17487 vdd.n1897 vdd.n1896 185
R17488 vdd.n1896 vdd.n1895 185
R17489 vdd.n1079 vdd.n1078 185
R17490 vdd.n1080 vdd.n1079 185
R17491 vdd.n1883 vdd.n1882 185
R17492 vdd.n1884 vdd.n1883 185
R17493 vdd.n1088 vdd.n1087 185
R17494 vdd.n1875 vdd.n1087 185
R17495 vdd.n1878 vdd.n1877 185
R17496 vdd.n1877 vdd.n1876 185
R17497 vdd.n1091 vdd.n1090 185
R17498 vdd.n1098 vdd.n1091 185
R17499 vdd.n1866 vdd.n1865 185
R17500 vdd.n1867 vdd.n1866 185
R17501 vdd.n1100 vdd.n1099 185
R17502 vdd.n1099 vdd.n1097 185
R17503 vdd.n1861 vdd.n1860 185
R17504 vdd.n1860 vdd.n1859 185
R17505 vdd.n1103 vdd.n1102 185
R17506 vdd.n1104 vdd.n1103 185
R17507 vdd.n1850 vdd.n1849 185
R17508 vdd.n1851 vdd.n1850 185
R17509 vdd.n1111 vdd.n1110 185
R17510 vdd.n1842 vdd.n1110 185
R17511 vdd.n1845 vdd.n1844 185
R17512 vdd.n1844 vdd.n1843 185
R17513 vdd.n1114 vdd.n1113 185
R17514 vdd.n1120 vdd.n1114 185
R17515 vdd.n1833 vdd.n1832 185
R17516 vdd.n1834 vdd.n1833 185
R17517 vdd.n1122 vdd.n1121 185
R17518 vdd.n1825 vdd.n1121 185
R17519 vdd.n1828 vdd.n1827 185
R17520 vdd.n1827 vdd.n1826 185
R17521 vdd.n1125 vdd.n1124 185
R17522 vdd.n1126 vdd.n1125 185
R17523 vdd.n1816 vdd.n1815 185
R17524 vdd.n1817 vdd.n1816 185
R17525 vdd.n1134 vdd.n1133 185
R17526 vdd.n1133 vdd.n1132 185
R17527 vdd.n1504 vdd.n1503 185
R17528 vdd.n1503 vdd.n1502 185
R17529 vdd.n1137 vdd.n1136 185
R17530 vdd.n1143 vdd.n1137 185
R17531 vdd.n1493 vdd.n1492 185
R17532 vdd.n1494 vdd.n1493 185
R17533 vdd.n1145 vdd.n1144 185
R17534 vdd.n1485 vdd.n1144 185
R17535 vdd.n1488 vdd.n1487 185
R17536 vdd.n1487 vdd.n1486 185
R17537 vdd.n1148 vdd.n1147 185
R17538 vdd.n1155 vdd.n1148 185
R17539 vdd.n1476 vdd.n1475 185
R17540 vdd.n1477 vdd.n1476 185
R17541 vdd.n1157 vdd.n1156 185
R17542 vdd.n1156 vdd.n1154 185
R17543 vdd.n1471 vdd.n1470 185
R17544 vdd.n1470 vdd.n1469 185
R17545 vdd.n1160 vdd.n1159 185
R17546 vdd.n1161 vdd.n1160 185
R17547 vdd.n1460 vdd.n1459 185
R17548 vdd.n1461 vdd.n1460 185
R17549 vdd.n1168 vdd.n1167 185
R17550 vdd.n1452 vdd.n1167 185
R17551 vdd.n1455 vdd.n1454 185
R17552 vdd.n1454 vdd.n1453 185
R17553 vdd.n1171 vdd.n1170 185
R17554 vdd.n1177 vdd.n1171 185
R17555 vdd.n1443 vdd.n1442 185
R17556 vdd.n1444 vdd.n1443 185
R17557 vdd.n1179 vdd.n1178 185
R17558 vdd.n1435 vdd.n1178 185
R17559 vdd.n1438 vdd.n1437 185
R17560 vdd.n1437 vdd.n1436 185
R17561 vdd.n1182 vdd.n1181 185
R17562 vdd.n1183 vdd.n1182 185
R17563 vdd.n1426 vdd.n1425 185
R17564 vdd.n1427 vdd.n1426 185
R17565 vdd.n1190 vdd.n1189 185
R17566 vdd.n1225 vdd.n1189 185
R17567 vdd.n1421 vdd.n1420 185
R17568 vdd.n1193 vdd.n1192 185
R17569 vdd.n1417 vdd.n1416 185
R17570 vdd.n1418 vdd.n1417 185
R17571 vdd.n1227 vdd.n1226 185
R17572 vdd.n1412 vdd.n1229 185
R17573 vdd.n1411 vdd.n1230 185
R17574 vdd.n1410 vdd.n1231 185
R17575 vdd.n1233 vdd.n1232 185
R17576 vdd.n1406 vdd.n1235 185
R17577 vdd.n1405 vdd.n1236 185
R17578 vdd.n1404 vdd.n1237 185
R17579 vdd.n1239 vdd.n1238 185
R17580 vdd.n1400 vdd.n1241 185
R17581 vdd.n1399 vdd.n1242 185
R17582 vdd.n1398 vdd.n1243 185
R17583 vdd.n1245 vdd.n1244 185
R17584 vdd.n1394 vdd.n1247 185
R17585 vdd.n1393 vdd.n1248 185
R17586 vdd.n1392 vdd.n1249 185
R17587 vdd.n1253 vdd.n1250 185
R17588 vdd.n1388 vdd.n1255 185
R17589 vdd.n1387 vdd.n1256 185
R17590 vdd.n1386 vdd.n1257 185
R17591 vdd.n1259 vdd.n1258 185
R17592 vdd.n1382 vdd.n1261 185
R17593 vdd.n1381 vdd.n1262 185
R17594 vdd.n1380 vdd.n1263 185
R17595 vdd.n1265 vdd.n1264 185
R17596 vdd.n1376 vdd.n1267 185
R17597 vdd.n1375 vdd.n1268 185
R17598 vdd.n1374 vdd.n1269 185
R17599 vdd.n1271 vdd.n1270 185
R17600 vdd.n1370 vdd.n1273 185
R17601 vdd.n1369 vdd.n1274 185
R17602 vdd.n1368 vdd.n1275 185
R17603 vdd.n1277 vdd.n1276 185
R17604 vdd.n1364 vdd.n1279 185
R17605 vdd.n1363 vdd.n1280 185
R17606 vdd.n1362 vdd.n1281 185
R17607 vdd.n1283 vdd.n1282 185
R17608 vdd.n1358 vdd.n1285 185
R17609 vdd.n1357 vdd.n1354 185
R17610 vdd.n1353 vdd.n1286 185
R17611 vdd.n1288 vdd.n1287 185
R17612 vdd.n1349 vdd.n1290 185
R17613 vdd.n1348 vdd.n1291 185
R17614 vdd.n1347 vdd.n1292 185
R17615 vdd.n1294 vdd.n1293 185
R17616 vdd.n1343 vdd.n1296 185
R17617 vdd.n1342 vdd.n1297 185
R17618 vdd.n1341 vdd.n1298 185
R17619 vdd.n1300 vdd.n1299 185
R17620 vdd.n1337 vdd.n1302 185
R17621 vdd.n1336 vdd.n1303 185
R17622 vdd.n1335 vdd.n1304 185
R17623 vdd.n1306 vdd.n1305 185
R17624 vdd.n1331 vdd.n1308 185
R17625 vdd.n1330 vdd.n1309 185
R17626 vdd.n1329 vdd.n1310 185
R17627 vdd.n1312 vdd.n1311 185
R17628 vdd.n1325 vdd.n1314 185
R17629 vdd.n1324 vdd.n1315 185
R17630 vdd.n1323 vdd.n1316 185
R17631 vdd.n1320 vdd.n1224 185
R17632 vdd.n1418 vdd.n1224 185
R17633 vdd.n2332 vdd.n2331 185
R17634 vdd.n2336 vdd.n1069 185
R17635 vdd.n1999 vdd.n1068 185
R17636 vdd.n2002 vdd.n2001 185
R17637 vdd.n2004 vdd.n2003 185
R17638 vdd.n2007 vdd.n2006 185
R17639 vdd.n2009 vdd.n2008 185
R17640 vdd.n2011 vdd.n1997 185
R17641 vdd.n2013 vdd.n2012 185
R17642 vdd.n2014 vdd.n1991 185
R17643 vdd.n2016 vdd.n2015 185
R17644 vdd.n2018 vdd.n1989 185
R17645 vdd.n2020 vdd.n2019 185
R17646 vdd.n2021 vdd.n1984 185
R17647 vdd.n2023 vdd.n2022 185
R17648 vdd.n2025 vdd.n1982 185
R17649 vdd.n2027 vdd.n2026 185
R17650 vdd.n2028 vdd.n1978 185
R17651 vdd.n2030 vdd.n2029 185
R17652 vdd.n2032 vdd.n1975 185
R17653 vdd.n2034 vdd.n2033 185
R17654 vdd.n1976 vdd.n1969 185
R17655 vdd.n2038 vdd.n1973 185
R17656 vdd.n2039 vdd.n1965 185
R17657 vdd.n2041 vdd.n2040 185
R17658 vdd.n2043 vdd.n1963 185
R17659 vdd.n2045 vdd.n2044 185
R17660 vdd.n2046 vdd.n1958 185
R17661 vdd.n2048 vdd.n2047 185
R17662 vdd.n2050 vdd.n1956 185
R17663 vdd.n2052 vdd.n2051 185
R17664 vdd.n2053 vdd.n1951 185
R17665 vdd.n2055 vdd.n2054 185
R17666 vdd.n2057 vdd.n1949 185
R17667 vdd.n2059 vdd.n2058 185
R17668 vdd.n2060 vdd.n1944 185
R17669 vdd.n2062 vdd.n2061 185
R17670 vdd.n2064 vdd.n1942 185
R17671 vdd.n2066 vdd.n2065 185
R17672 vdd.n2067 vdd.n1938 185
R17673 vdd.n2069 vdd.n2068 185
R17674 vdd.n2071 vdd.n1935 185
R17675 vdd.n2073 vdd.n2072 185
R17676 vdd.n1936 vdd.n1929 185
R17677 vdd.n2077 vdd.n1933 185
R17678 vdd.n2078 vdd.n1925 185
R17679 vdd.n2080 vdd.n2079 185
R17680 vdd.n2082 vdd.n1923 185
R17681 vdd.n2084 vdd.n2083 185
R17682 vdd.n2085 vdd.n1918 185
R17683 vdd.n2087 vdd.n2086 185
R17684 vdd.n2089 vdd.n1916 185
R17685 vdd.n2091 vdd.n2090 185
R17686 vdd.n2092 vdd.n1911 185
R17687 vdd.n2094 vdd.n2093 185
R17688 vdd.n2096 vdd.n1910 185
R17689 vdd.n2097 vdd.n1907 185
R17690 vdd.n2100 vdd.n2099 185
R17691 vdd.n1909 vdd.n1905 185
R17692 vdd.n2317 vdd.n1903 185
R17693 vdd.n2319 vdd.n2318 185
R17694 vdd.n2321 vdd.n1901 185
R17695 vdd.n2323 vdd.n2322 185
R17696 vdd.n2324 vdd.n1075 185
R17697 vdd.n2330 vdd.n1072 185
R17698 vdd.n2330 vdd.n2329 185
R17699 vdd.n1083 vdd.n1071 185
R17700 vdd.n1894 vdd.n1071 185
R17701 vdd.n1893 vdd.n1892 185
R17702 vdd.n1895 vdd.n1893 185
R17703 vdd.n1082 vdd.n1081 185
R17704 vdd.n1081 vdd.n1080 185
R17705 vdd.n1886 vdd.n1885 185
R17706 vdd.n1885 vdd.n1884 185
R17707 vdd.n1086 vdd.n1085 185
R17708 vdd.n1875 vdd.n1086 185
R17709 vdd.n1874 vdd.n1873 185
R17710 vdd.n1876 vdd.n1874 185
R17711 vdd.n1093 vdd.n1092 185
R17712 vdd.n1098 vdd.n1092 185
R17713 vdd.n1869 vdd.n1868 185
R17714 vdd.n1868 vdd.n1867 185
R17715 vdd.n1096 vdd.n1095 185
R17716 vdd.n1097 vdd.n1096 185
R17717 vdd.n1858 vdd.n1857 185
R17718 vdd.n1859 vdd.n1858 185
R17719 vdd.n1106 vdd.n1105 185
R17720 vdd.n1105 vdd.n1104 185
R17721 vdd.n1853 vdd.n1852 185
R17722 vdd.n1852 vdd.n1851 185
R17723 vdd.n1109 vdd.n1108 185
R17724 vdd.n1842 vdd.n1109 185
R17725 vdd.n1841 vdd.n1840 185
R17726 vdd.n1843 vdd.n1841 185
R17727 vdd.n1116 vdd.n1115 185
R17728 vdd.n1120 vdd.n1115 185
R17729 vdd.n1836 vdd.n1835 185
R17730 vdd.n1835 vdd.n1834 185
R17731 vdd.n1119 vdd.n1118 185
R17732 vdd.n1825 vdd.n1119 185
R17733 vdd.n1824 vdd.n1823 185
R17734 vdd.n1826 vdd.n1824 185
R17735 vdd.n1128 vdd.n1127 185
R17736 vdd.n1127 vdd.n1126 185
R17737 vdd.n1819 vdd.n1818 185
R17738 vdd.n1818 vdd.n1817 185
R17739 vdd.n1131 vdd.n1130 185
R17740 vdd.n1132 vdd.n1131 185
R17741 vdd.n1501 vdd.n1500 185
R17742 vdd.n1502 vdd.n1501 185
R17743 vdd.n1139 vdd.n1138 185
R17744 vdd.n1143 vdd.n1138 185
R17745 vdd.n1496 vdd.n1495 185
R17746 vdd.n1495 vdd.n1494 185
R17747 vdd.n1142 vdd.n1141 185
R17748 vdd.n1485 vdd.n1142 185
R17749 vdd.n1484 vdd.n1483 185
R17750 vdd.n1486 vdd.n1484 185
R17751 vdd.n1150 vdd.n1149 185
R17752 vdd.n1155 vdd.n1149 185
R17753 vdd.n1479 vdd.n1478 185
R17754 vdd.n1478 vdd.n1477 185
R17755 vdd.n1153 vdd.n1152 185
R17756 vdd.n1154 vdd.n1153 185
R17757 vdd.n1468 vdd.n1467 185
R17758 vdd.n1469 vdd.n1468 185
R17759 vdd.n1163 vdd.n1162 185
R17760 vdd.n1162 vdd.n1161 185
R17761 vdd.n1463 vdd.n1462 185
R17762 vdd.n1462 vdd.n1461 185
R17763 vdd.n1166 vdd.n1165 185
R17764 vdd.n1452 vdd.n1166 185
R17765 vdd.n1451 vdd.n1450 185
R17766 vdd.n1453 vdd.n1451 185
R17767 vdd.n1173 vdd.n1172 185
R17768 vdd.n1177 vdd.n1172 185
R17769 vdd.n1446 vdd.n1445 185
R17770 vdd.n1445 vdd.n1444 185
R17771 vdd.n1176 vdd.n1175 185
R17772 vdd.n1435 vdd.n1176 185
R17773 vdd.n1434 vdd.n1433 185
R17774 vdd.n1436 vdd.n1434 185
R17775 vdd.n1185 vdd.n1184 185
R17776 vdd.n1184 vdd.n1183 185
R17777 vdd.n1429 vdd.n1428 185
R17778 vdd.n1428 vdd.n1427 185
R17779 vdd.n1188 vdd.n1187 185
R17780 vdd.n1225 vdd.n1188 185
R17781 vdd.n956 vdd.n954 185
R17782 vdd.n2532 vdd.n954 185
R17783 vdd.n2454 vdd.n973 185
R17784 vdd.n973 vdd.t159 185
R17785 vdd.n2456 vdd.n2455 185
R17786 vdd.n2457 vdd.n2456 185
R17787 vdd.n2453 vdd.n972 185
R17788 vdd.n2156 vdd.n972 185
R17789 vdd.n2452 vdd.n2451 185
R17790 vdd.n2451 vdd.n2450 185
R17791 vdd.n975 vdd.n974 185
R17792 vdd.n976 vdd.n975 185
R17793 vdd.n2441 vdd.n2440 185
R17794 vdd.n2442 vdd.n2441 185
R17795 vdd.n2439 vdd.n986 185
R17796 vdd.n986 vdd.n983 185
R17797 vdd.n2438 vdd.n2437 185
R17798 vdd.n2437 vdd.n2436 185
R17799 vdd.n988 vdd.n987 185
R17800 vdd.n989 vdd.n988 185
R17801 vdd.n2429 vdd.n2428 185
R17802 vdd.n2430 vdd.n2429 185
R17803 vdd.n2427 vdd.n997 185
R17804 vdd.n1002 vdd.n997 185
R17805 vdd.n2426 vdd.n2425 185
R17806 vdd.n2425 vdd.n2424 185
R17807 vdd.n999 vdd.n998 185
R17808 vdd.n1008 vdd.n999 185
R17809 vdd.n2417 vdd.n2416 185
R17810 vdd.n2418 vdd.n2417 185
R17811 vdd.n2415 vdd.n1009 185
R17812 vdd.n2257 vdd.n1009 185
R17813 vdd.n2414 vdd.n2413 185
R17814 vdd.n2413 vdd.n2412 185
R17815 vdd.n1011 vdd.n1010 185
R17816 vdd.n1012 vdd.n1011 185
R17817 vdd.n2405 vdd.n2404 185
R17818 vdd.n2406 vdd.n2405 185
R17819 vdd.n2403 vdd.n1021 185
R17820 vdd.n1021 vdd.n1018 185
R17821 vdd.n2402 vdd.n2401 185
R17822 vdd.n2401 vdd.n2400 185
R17823 vdd.n1023 vdd.n1022 185
R17824 vdd.n1033 vdd.n1023 185
R17825 vdd.n2392 vdd.n2391 185
R17826 vdd.n2393 vdd.n2392 185
R17827 vdd.n2390 vdd.n1034 185
R17828 vdd.n1034 vdd.n1030 185
R17829 vdd.n2389 vdd.n2388 185
R17830 vdd.n2388 vdd.n2387 185
R17831 vdd.n1036 vdd.n1035 185
R17832 vdd.n1037 vdd.n1036 185
R17833 vdd.n2380 vdd.n2379 185
R17834 vdd.n2381 vdd.n2380 185
R17835 vdd.n2378 vdd.n1046 185
R17836 vdd.n1046 vdd.n1043 185
R17837 vdd.n2377 vdd.n2376 185
R17838 vdd.n2376 vdd.n2375 185
R17839 vdd.n1048 vdd.n1047 185
R17840 vdd.n2112 vdd.n2111 185
R17841 vdd.n2113 vdd.n2109 185
R17842 vdd.n2109 vdd.n1049 185
R17843 vdd.n2115 vdd.n2114 185
R17844 vdd.n2117 vdd.n2108 185
R17845 vdd.n2120 vdd.n2119 185
R17846 vdd.n2121 vdd.n2107 185
R17847 vdd.n2123 vdd.n2122 185
R17848 vdd.n2125 vdd.n2106 185
R17849 vdd.n2128 vdd.n2127 185
R17850 vdd.n2129 vdd.n2105 185
R17851 vdd.n2131 vdd.n2130 185
R17852 vdd.n2133 vdd.n2104 185
R17853 vdd.n2136 vdd.n2135 185
R17854 vdd.n2137 vdd.n2103 185
R17855 vdd.n2139 vdd.n2138 185
R17856 vdd.n2141 vdd.n2102 185
R17857 vdd.n2314 vdd.n2142 185
R17858 vdd.n2313 vdd.n2312 185
R17859 vdd.n2310 vdd.n2143 185
R17860 vdd.n2308 vdd.n2307 185
R17861 vdd.n2306 vdd.n2144 185
R17862 vdd.n2305 vdd.n2304 185
R17863 vdd.n2302 vdd.n2145 185
R17864 vdd.n2300 vdd.n2299 185
R17865 vdd.n2298 vdd.n2146 185
R17866 vdd.n2297 vdd.n2296 185
R17867 vdd.n2294 vdd.n2147 185
R17868 vdd.n2292 vdd.n2291 185
R17869 vdd.n2290 vdd.n2148 185
R17870 vdd.n2289 vdd.n2288 185
R17871 vdd.n2286 vdd.n2149 185
R17872 vdd.n2284 vdd.n2283 185
R17873 vdd.n2282 vdd.n2150 185
R17874 vdd.n2281 vdd.n2280 185
R17875 vdd.n2535 vdd.n2534 185
R17876 vdd.n2537 vdd.n2536 185
R17877 vdd.n2539 vdd.n2538 185
R17878 vdd.n2542 vdd.n2541 185
R17879 vdd.n2544 vdd.n2543 185
R17880 vdd.n2546 vdd.n2545 185
R17881 vdd.n2548 vdd.n2547 185
R17882 vdd.n2550 vdd.n2549 185
R17883 vdd.n2552 vdd.n2551 185
R17884 vdd.n2554 vdd.n2553 185
R17885 vdd.n2556 vdd.n2555 185
R17886 vdd.n2558 vdd.n2557 185
R17887 vdd.n2560 vdd.n2559 185
R17888 vdd.n2562 vdd.n2561 185
R17889 vdd.n2564 vdd.n2563 185
R17890 vdd.n2566 vdd.n2565 185
R17891 vdd.n2568 vdd.n2567 185
R17892 vdd.n2570 vdd.n2569 185
R17893 vdd.n2572 vdd.n2571 185
R17894 vdd.n2574 vdd.n2573 185
R17895 vdd.n2576 vdd.n2575 185
R17896 vdd.n2578 vdd.n2577 185
R17897 vdd.n2580 vdd.n2579 185
R17898 vdd.n2582 vdd.n2581 185
R17899 vdd.n2584 vdd.n2583 185
R17900 vdd.n2586 vdd.n2585 185
R17901 vdd.n2588 vdd.n2587 185
R17902 vdd.n2590 vdd.n2589 185
R17903 vdd.n2592 vdd.n2591 185
R17904 vdd.n2594 vdd.n2593 185
R17905 vdd.n2596 vdd.n2595 185
R17906 vdd.n2598 vdd.n2597 185
R17907 vdd.n2600 vdd.n2599 185
R17908 vdd.n2601 vdd.n955 185
R17909 vdd.n2603 vdd.n2602 185
R17910 vdd.n2604 vdd.n2603 185
R17911 vdd.n2533 vdd.n959 185
R17912 vdd.n2533 vdd.n2532 185
R17913 vdd.n2154 vdd.n960 185
R17914 vdd.t159 vdd.n960 185
R17915 vdd.n2155 vdd.n970 185
R17916 vdd.n2457 vdd.n970 185
R17917 vdd.n2158 vdd.n2157 185
R17918 vdd.n2157 vdd.n2156 185
R17919 vdd.n2159 vdd.n977 185
R17920 vdd.n2450 vdd.n977 185
R17921 vdd.n2161 vdd.n2160 185
R17922 vdd.n2160 vdd.n976 185
R17923 vdd.n2162 vdd.n984 185
R17924 vdd.n2442 vdd.n984 185
R17925 vdd.n2164 vdd.n2163 185
R17926 vdd.n2163 vdd.n983 185
R17927 vdd.n2165 vdd.n990 185
R17928 vdd.n2436 vdd.n990 185
R17929 vdd.n2167 vdd.n2166 185
R17930 vdd.n2166 vdd.n989 185
R17931 vdd.n2168 vdd.n995 185
R17932 vdd.n2430 vdd.n995 185
R17933 vdd.n2170 vdd.n2169 185
R17934 vdd.n2169 vdd.n1002 185
R17935 vdd.n2171 vdd.n1000 185
R17936 vdd.n2424 vdd.n1000 185
R17937 vdd.n2173 vdd.n2172 185
R17938 vdd.n2172 vdd.n1008 185
R17939 vdd.n2174 vdd.n1006 185
R17940 vdd.n2418 vdd.n1006 185
R17941 vdd.n2259 vdd.n2258 185
R17942 vdd.n2258 vdd.n2257 185
R17943 vdd.n2260 vdd.n1013 185
R17944 vdd.n2412 vdd.n1013 185
R17945 vdd.n2262 vdd.n2261 185
R17946 vdd.n2261 vdd.n1012 185
R17947 vdd.n2263 vdd.n1019 185
R17948 vdd.n2406 vdd.n1019 185
R17949 vdd.n2265 vdd.n2264 185
R17950 vdd.n2264 vdd.n1018 185
R17951 vdd.n2266 vdd.n1024 185
R17952 vdd.n2400 vdd.n1024 185
R17953 vdd.n2268 vdd.n2267 185
R17954 vdd.n2267 vdd.n1033 185
R17955 vdd.n2269 vdd.n1031 185
R17956 vdd.n2393 vdd.n1031 185
R17957 vdd.n2271 vdd.n2270 185
R17958 vdd.n2270 vdd.n1030 185
R17959 vdd.n2272 vdd.n1038 185
R17960 vdd.n2387 vdd.n1038 185
R17961 vdd.n2274 vdd.n2273 185
R17962 vdd.n2273 vdd.n1037 185
R17963 vdd.n2275 vdd.n1044 185
R17964 vdd.n2381 vdd.n1044 185
R17965 vdd.n2277 vdd.n2276 185
R17966 vdd.n2276 vdd.n1043 185
R17967 vdd.n2278 vdd.n1050 185
R17968 vdd.n2375 vdd.n1050 185
R17969 vdd.n3357 vdd.n3356 185
R17970 vdd.n3356 vdd.n3355 185
R17971 vdd.n3358 vdd.n387 185
R17972 vdd.n387 vdd.n386 185
R17973 vdd.n3360 vdd.n3359 185
R17974 vdd.n3361 vdd.n3360 185
R17975 vdd.n382 vdd.n381 185
R17976 vdd.n3362 vdd.n382 185
R17977 vdd.n3365 vdd.n3364 185
R17978 vdd.n3364 vdd.n3363 185
R17979 vdd.n3366 vdd.n376 185
R17980 vdd.n376 vdd.n375 185
R17981 vdd.n3368 vdd.n3367 185
R17982 vdd.n3369 vdd.n3368 185
R17983 vdd.n371 vdd.n370 185
R17984 vdd.n3370 vdd.n371 185
R17985 vdd.n3373 vdd.n3372 185
R17986 vdd.n3372 vdd.n3371 185
R17987 vdd.n3374 vdd.n365 185
R17988 vdd.n3331 vdd.n365 185
R17989 vdd.n3376 vdd.n3375 185
R17990 vdd.n3377 vdd.n3376 185
R17991 vdd.n360 vdd.n359 185
R17992 vdd.n3378 vdd.n360 185
R17993 vdd.n3381 vdd.n3380 185
R17994 vdd.n3380 vdd.n3379 185
R17995 vdd.n3382 vdd.n354 185
R17996 vdd.n361 vdd.n354 185
R17997 vdd.n3384 vdd.n3383 185
R17998 vdd.n3385 vdd.n3384 185
R17999 vdd.n350 vdd.n349 185
R18000 vdd.n3386 vdd.n350 185
R18001 vdd.n3389 vdd.n3388 185
R18002 vdd.n3388 vdd.n3387 185
R18003 vdd.n3390 vdd.n345 185
R18004 vdd.n345 vdd.n344 185
R18005 vdd.n3392 vdd.n3391 185
R18006 vdd.n3393 vdd.n3392 185
R18007 vdd.n339 vdd.n337 185
R18008 vdd.n3394 vdd.n339 185
R18009 vdd.n3397 vdd.n3396 185
R18010 vdd.n3396 vdd.n3395 185
R18011 vdd.n338 vdd.n336 185
R18012 vdd.n340 vdd.n338 185
R18013 vdd.n3307 vdd.n3306 185
R18014 vdd.n3308 vdd.n3307 185
R18015 vdd.n635 vdd.n634 185
R18016 vdd.n634 vdd.n633 185
R18017 vdd.n3302 vdd.n3301 185
R18018 vdd.n3301 vdd.n3300 185
R18019 vdd.n638 vdd.n637 185
R18020 vdd.n644 vdd.n638 185
R18021 vdd.n3288 vdd.n3287 185
R18022 vdd.n3289 vdd.n3288 185
R18023 vdd.n646 vdd.n645 185
R18024 vdd.n3280 vdd.n645 185
R18025 vdd.n3283 vdd.n3282 185
R18026 vdd.n3282 vdd.n3281 185
R18027 vdd.n649 vdd.n648 185
R18028 vdd.n656 vdd.n649 185
R18029 vdd.n3271 vdd.n3270 185
R18030 vdd.n3272 vdd.n3271 185
R18031 vdd.n658 vdd.n657 185
R18032 vdd.n657 vdd.n655 185
R18033 vdd.n3266 vdd.n3265 185
R18034 vdd.n3265 vdd.n3264 185
R18035 vdd.n661 vdd.n660 185
R18036 vdd.n662 vdd.n661 185
R18037 vdd.n3255 vdd.n3254 185
R18038 vdd.n3256 vdd.n3255 185
R18039 vdd.n669 vdd.n668 185
R18040 vdd.n3247 vdd.n668 185
R18041 vdd.n3250 vdd.n3249 185
R18042 vdd.n3249 vdd.n3248 185
R18043 vdd.n672 vdd.n671 185
R18044 vdd.n679 vdd.n672 185
R18045 vdd.n3238 vdd.n3237 185
R18046 vdd.n3239 vdd.n3238 185
R18047 vdd.n681 vdd.n680 185
R18048 vdd.n680 vdd.n678 185
R18049 vdd.n3233 vdd.n3232 185
R18050 vdd.n3232 vdd.n3231 185
R18051 vdd.n684 vdd.n683 185
R18052 vdd.n723 vdd.n684 185
R18053 vdd.n3221 vdd.n3220 185
R18054 vdd.n3219 vdd.n725 185
R18055 vdd.n3218 vdd.n724 185
R18056 vdd.n3223 vdd.n724 185
R18057 vdd.n729 vdd.n728 185
R18058 vdd.n733 vdd.n732 185
R18059 vdd.n3214 vdd.n734 185
R18060 vdd.n3213 vdd.n3212 185
R18061 vdd.n3211 vdd.n3210 185
R18062 vdd.n3209 vdd.n3208 185
R18063 vdd.n3207 vdd.n3206 185
R18064 vdd.n3205 vdd.n3204 185
R18065 vdd.n3203 vdd.n3202 185
R18066 vdd.n3201 vdd.n3200 185
R18067 vdd.n3199 vdd.n3198 185
R18068 vdd.n3197 vdd.n3196 185
R18069 vdd.n3195 vdd.n3194 185
R18070 vdd.n3193 vdd.n3192 185
R18071 vdd.n3191 vdd.n3190 185
R18072 vdd.n3189 vdd.n3188 185
R18073 vdd.n3187 vdd.n3186 185
R18074 vdd.n3178 vdd.n747 185
R18075 vdd.n3180 vdd.n3179 185
R18076 vdd.n3177 vdd.n3176 185
R18077 vdd.n3175 vdd.n3174 185
R18078 vdd.n3173 vdd.n3172 185
R18079 vdd.n3171 vdd.n3170 185
R18080 vdd.n3169 vdd.n3168 185
R18081 vdd.n3167 vdd.n3166 185
R18082 vdd.n3165 vdd.n3164 185
R18083 vdd.n3163 vdd.n3162 185
R18084 vdd.n3161 vdd.n3160 185
R18085 vdd.n3159 vdd.n3158 185
R18086 vdd.n3157 vdd.n3156 185
R18087 vdd.n3155 vdd.n3154 185
R18088 vdd.n3153 vdd.n3152 185
R18089 vdd.n3151 vdd.n3150 185
R18090 vdd.n3149 vdd.n3148 185
R18091 vdd.n3147 vdd.n3146 185
R18092 vdd.n3145 vdd.n3144 185
R18093 vdd.n3143 vdd.n3142 185
R18094 vdd.n3141 vdd.n3140 185
R18095 vdd.n3139 vdd.n3138 185
R18096 vdd.n3132 vdd.n767 185
R18097 vdd.n3134 vdd.n3133 185
R18098 vdd.n3131 vdd.n3130 185
R18099 vdd.n3129 vdd.n3128 185
R18100 vdd.n3127 vdd.n3126 185
R18101 vdd.n3125 vdd.n3124 185
R18102 vdd.n3123 vdd.n3122 185
R18103 vdd.n3121 vdd.n3120 185
R18104 vdd.n3119 vdd.n3118 185
R18105 vdd.n3117 vdd.n3116 185
R18106 vdd.n3115 vdd.n3114 185
R18107 vdd.n3113 vdd.n3112 185
R18108 vdd.n3111 vdd.n3110 185
R18109 vdd.n3109 vdd.n3108 185
R18110 vdd.n3107 vdd.n3106 185
R18111 vdd.n3105 vdd.n3104 185
R18112 vdd.n3103 vdd.n3102 185
R18113 vdd.n3101 vdd.n3100 185
R18114 vdd.n3099 vdd.n3098 185
R18115 vdd.n3097 vdd.n3096 185
R18116 vdd.n3095 vdd.n691 185
R18117 vdd.n3225 vdd.n3224 185
R18118 vdd.n3224 vdd.n3223 185
R18119 vdd.n3352 vdd.n3351 185
R18120 vdd.n618 vdd.n425 185
R18121 vdd.n617 vdd.n616 185
R18122 vdd.n615 vdd.n614 185
R18123 vdd.n613 vdd.n430 185
R18124 vdd.n609 vdd.n608 185
R18125 vdd.n607 vdd.n606 185
R18126 vdd.n605 vdd.n604 185
R18127 vdd.n603 vdd.n432 185
R18128 vdd.n599 vdd.n598 185
R18129 vdd.n597 vdd.n596 185
R18130 vdd.n595 vdd.n594 185
R18131 vdd.n593 vdd.n434 185
R18132 vdd.n589 vdd.n588 185
R18133 vdd.n587 vdd.n586 185
R18134 vdd.n585 vdd.n584 185
R18135 vdd.n583 vdd.n436 185
R18136 vdd.n579 vdd.n578 185
R18137 vdd.n577 vdd.n576 185
R18138 vdd.n575 vdd.n574 185
R18139 vdd.n573 vdd.n438 185
R18140 vdd.n569 vdd.n568 185
R18141 vdd.n567 vdd.n566 185
R18142 vdd.n565 vdd.n564 185
R18143 vdd.n563 vdd.n442 185
R18144 vdd.n559 vdd.n558 185
R18145 vdd.n557 vdd.n556 185
R18146 vdd.n555 vdd.n554 185
R18147 vdd.n553 vdd.n444 185
R18148 vdd.n549 vdd.n548 185
R18149 vdd.n547 vdd.n546 185
R18150 vdd.n545 vdd.n544 185
R18151 vdd.n543 vdd.n446 185
R18152 vdd.n539 vdd.n538 185
R18153 vdd.n537 vdd.n536 185
R18154 vdd.n535 vdd.n534 185
R18155 vdd.n533 vdd.n448 185
R18156 vdd.n529 vdd.n528 185
R18157 vdd.n527 vdd.n526 185
R18158 vdd.n525 vdd.n524 185
R18159 vdd.n523 vdd.n450 185
R18160 vdd.n519 vdd.n518 185
R18161 vdd.n517 vdd.n516 185
R18162 vdd.n515 vdd.n514 185
R18163 vdd.n513 vdd.n454 185
R18164 vdd.n509 vdd.n508 185
R18165 vdd.n507 vdd.n506 185
R18166 vdd.n505 vdd.n504 185
R18167 vdd.n503 vdd.n456 185
R18168 vdd.n499 vdd.n498 185
R18169 vdd.n497 vdd.n496 185
R18170 vdd.n495 vdd.n494 185
R18171 vdd.n493 vdd.n458 185
R18172 vdd.n489 vdd.n488 185
R18173 vdd.n487 vdd.n486 185
R18174 vdd.n485 vdd.n484 185
R18175 vdd.n483 vdd.n460 185
R18176 vdd.n479 vdd.n478 185
R18177 vdd.n477 vdd.n476 185
R18178 vdd.n475 vdd.n474 185
R18179 vdd.n473 vdd.n462 185
R18180 vdd.n469 vdd.n468 185
R18181 vdd.n467 vdd.n466 185
R18182 vdd.n465 vdd.n392 185
R18183 vdd.n3348 vdd.n393 185
R18184 vdd.n3355 vdd.n393 185
R18185 vdd.n3347 vdd.n3346 185
R18186 vdd.n3346 vdd.n386 185
R18187 vdd.n3345 vdd.n385 185
R18188 vdd.n3361 vdd.n385 185
R18189 vdd.n621 vdd.n384 185
R18190 vdd.n3362 vdd.n384 185
R18191 vdd.n3341 vdd.n383 185
R18192 vdd.n3363 vdd.n383 185
R18193 vdd.n3340 vdd.n3339 185
R18194 vdd.n3339 vdd.n375 185
R18195 vdd.n3338 vdd.n374 185
R18196 vdd.n3369 vdd.n374 185
R18197 vdd.n623 vdd.n373 185
R18198 vdd.n3370 vdd.n373 185
R18199 vdd.n3334 vdd.n372 185
R18200 vdd.n3371 vdd.n372 185
R18201 vdd.n3333 vdd.n3332 185
R18202 vdd.n3332 vdd.n3331 185
R18203 vdd.n3330 vdd.n364 185
R18204 vdd.n3377 vdd.n364 185
R18205 vdd.n625 vdd.n363 185
R18206 vdd.n3378 vdd.n363 185
R18207 vdd.n3326 vdd.n362 185
R18208 vdd.n3379 vdd.n362 185
R18209 vdd.n3325 vdd.n3324 185
R18210 vdd.n3324 vdd.n361 185
R18211 vdd.n3323 vdd.n353 185
R18212 vdd.n3385 vdd.n353 185
R18213 vdd.n627 vdd.n352 185
R18214 vdd.n3386 vdd.n352 185
R18215 vdd.n3319 vdd.n351 185
R18216 vdd.n3387 vdd.n351 185
R18217 vdd.n3318 vdd.n3317 185
R18218 vdd.n3317 vdd.n344 185
R18219 vdd.n3316 vdd.n343 185
R18220 vdd.n3393 vdd.n343 185
R18221 vdd.n629 vdd.n342 185
R18222 vdd.n3394 vdd.n342 185
R18223 vdd.n3312 vdd.n341 185
R18224 vdd.n3395 vdd.n341 185
R18225 vdd.n3311 vdd.n3310 185
R18226 vdd.n3310 vdd.n340 185
R18227 vdd.n3309 vdd.n631 185
R18228 vdd.n3309 vdd.n3308 185
R18229 vdd.n3297 vdd.n632 185
R18230 vdd.n633 vdd.n632 185
R18231 vdd.n3299 vdd.n3298 185
R18232 vdd.n3300 vdd.n3299 185
R18233 vdd.n640 vdd.n639 185
R18234 vdd.n644 vdd.n639 185
R18235 vdd.n3291 vdd.n3290 185
R18236 vdd.n3290 vdd.n3289 185
R18237 vdd.n643 vdd.n642 185
R18238 vdd.n3280 vdd.n643 185
R18239 vdd.n3279 vdd.n3278 185
R18240 vdd.n3281 vdd.n3279 185
R18241 vdd.n651 vdd.n650 185
R18242 vdd.n656 vdd.n650 185
R18243 vdd.n3274 vdd.n3273 185
R18244 vdd.n3273 vdd.n3272 185
R18245 vdd.n654 vdd.n653 185
R18246 vdd.n655 vdd.n654 185
R18247 vdd.n3263 vdd.n3262 185
R18248 vdd.n3264 vdd.n3263 185
R18249 vdd.n664 vdd.n663 185
R18250 vdd.n663 vdd.n662 185
R18251 vdd.n3258 vdd.n3257 185
R18252 vdd.n3257 vdd.n3256 185
R18253 vdd.n667 vdd.n666 185
R18254 vdd.n3247 vdd.n667 185
R18255 vdd.n3246 vdd.n3245 185
R18256 vdd.n3248 vdd.n3246 185
R18257 vdd.n674 vdd.n673 185
R18258 vdd.n679 vdd.n673 185
R18259 vdd.n3241 vdd.n3240 185
R18260 vdd.n3240 vdd.n3239 185
R18261 vdd.n677 vdd.n676 185
R18262 vdd.n678 vdd.n677 185
R18263 vdd.n3230 vdd.n3229 185
R18264 vdd.n3231 vdd.n3230 185
R18265 vdd.n686 vdd.n685 185
R18266 vdd.n723 vdd.n685 185
R18267 vdd.n913 vdd.n912 185
R18268 vdd.n2855 vdd.n2854 185
R18269 vdd.n2853 vdd.n2638 185
R18270 vdd.n2857 vdd.n2638 185
R18271 vdd.n2852 vdd.n2851 185
R18272 vdd.n2850 vdd.n2849 185
R18273 vdd.n2848 vdd.n2847 185
R18274 vdd.n2846 vdd.n2845 185
R18275 vdd.n2844 vdd.n2843 185
R18276 vdd.n2842 vdd.n2841 185
R18277 vdd.n2840 vdd.n2839 185
R18278 vdd.n2838 vdd.n2837 185
R18279 vdd.n2836 vdd.n2835 185
R18280 vdd.n2834 vdd.n2833 185
R18281 vdd.n2832 vdd.n2831 185
R18282 vdd.n2830 vdd.n2829 185
R18283 vdd.n2828 vdd.n2827 185
R18284 vdd.n2826 vdd.n2825 185
R18285 vdd.n2824 vdd.n2823 185
R18286 vdd.n2822 vdd.n2821 185
R18287 vdd.n2820 vdd.n2819 185
R18288 vdd.n2818 vdd.n2817 185
R18289 vdd.n2816 vdd.n2815 185
R18290 vdd.n2814 vdd.n2813 185
R18291 vdd.n2812 vdd.n2811 185
R18292 vdd.n2810 vdd.n2809 185
R18293 vdd.n2808 vdd.n2807 185
R18294 vdd.n2806 vdd.n2805 185
R18295 vdd.n2804 vdd.n2803 185
R18296 vdd.n2802 vdd.n2801 185
R18297 vdd.n2800 vdd.n2799 185
R18298 vdd.n2798 vdd.n2797 185
R18299 vdd.n2796 vdd.n2795 185
R18300 vdd.n2793 vdd.n2792 185
R18301 vdd.n2791 vdd.n2790 185
R18302 vdd.n2789 vdd.n2788 185
R18303 vdd.n2995 vdd.n2994 185
R18304 vdd.n2997 vdd.n834 185
R18305 vdd.n2999 vdd.n2998 185
R18306 vdd.n3001 vdd.n831 185
R18307 vdd.n3003 vdd.n3002 185
R18308 vdd.n3005 vdd.n829 185
R18309 vdd.n3007 vdd.n3006 185
R18310 vdd.n3008 vdd.n828 185
R18311 vdd.n3010 vdd.n3009 185
R18312 vdd.n3012 vdd.n826 185
R18313 vdd.n3014 vdd.n3013 185
R18314 vdd.n3015 vdd.n825 185
R18315 vdd.n3017 vdd.n3016 185
R18316 vdd.n3019 vdd.n823 185
R18317 vdd.n3021 vdd.n3020 185
R18318 vdd.n3022 vdd.n822 185
R18319 vdd.n3024 vdd.n3023 185
R18320 vdd.n3026 vdd.n731 185
R18321 vdd.n3028 vdd.n3027 185
R18322 vdd.n3030 vdd.n820 185
R18323 vdd.n3032 vdd.n3031 185
R18324 vdd.n3033 vdd.n819 185
R18325 vdd.n3035 vdd.n3034 185
R18326 vdd.n3037 vdd.n817 185
R18327 vdd.n3039 vdd.n3038 185
R18328 vdd.n3040 vdd.n816 185
R18329 vdd.n3042 vdd.n3041 185
R18330 vdd.n3044 vdd.n814 185
R18331 vdd.n3046 vdd.n3045 185
R18332 vdd.n3047 vdd.n813 185
R18333 vdd.n3049 vdd.n3048 185
R18334 vdd.n3051 vdd.n812 185
R18335 vdd.n3052 vdd.n811 185
R18336 vdd.n3055 vdd.n3054 185
R18337 vdd.n3056 vdd.n809 185
R18338 vdd.n809 vdd.n692 185
R18339 vdd.n2993 vdd.n806 185
R18340 vdd.n3059 vdd.n806 185
R18341 vdd.n2992 vdd.n2991 185
R18342 vdd.n2991 vdd.n805 185
R18343 vdd.n2990 vdd.n836 185
R18344 vdd.n2990 vdd.n2989 185
R18345 vdd.n2744 vdd.n837 185
R18346 vdd.n846 vdd.n837 185
R18347 vdd.n2745 vdd.n844 185
R18348 vdd.n2983 vdd.n844 185
R18349 vdd.n2747 vdd.n2746 185
R18350 vdd.n2746 vdd.n843 185
R18351 vdd.n2748 vdd.n852 185
R18352 vdd.n2932 vdd.n852 185
R18353 vdd.n2750 vdd.n2749 185
R18354 vdd.n2749 vdd.n851 185
R18355 vdd.n2751 vdd.n858 185
R18356 vdd.n2926 vdd.n858 185
R18357 vdd.n2753 vdd.n2752 185
R18358 vdd.n2752 vdd.n857 185
R18359 vdd.n2754 vdd.n863 185
R18360 vdd.n2918 vdd.n863 185
R18361 vdd.n2756 vdd.n2755 185
R18362 vdd.n2755 vdd.n870 185
R18363 vdd.n2757 vdd.n868 185
R18364 vdd.n2912 vdd.n868 185
R18365 vdd.n2759 vdd.n2758 185
R18366 vdd.n2760 vdd.n2759 185
R18367 vdd.n2743 vdd.n875 185
R18368 vdd.n2906 vdd.n875 185
R18369 vdd.n2742 vdd.n2741 185
R18370 vdd.n2741 vdd.n874 185
R18371 vdd.n2740 vdd.n881 185
R18372 vdd.n2900 vdd.n881 185
R18373 vdd.n2739 vdd.n2738 185
R18374 vdd.n2738 vdd.n880 185
R18375 vdd.n2737 vdd.n886 185
R18376 vdd.n2894 vdd.n886 185
R18377 vdd.n2736 vdd.n2735 185
R18378 vdd.n2735 vdd.n893 185
R18379 vdd.n2734 vdd.n891 185
R18380 vdd.n2888 vdd.n891 185
R18381 vdd.n2733 vdd.n2732 185
R18382 vdd.n2732 vdd.n900 185
R18383 vdd.n2731 vdd.n898 185
R18384 vdd.n2882 vdd.n898 185
R18385 vdd.n2730 vdd.n2729 185
R18386 vdd.n2729 vdd.n897 185
R18387 vdd.n2641 vdd.n904 185
R18388 vdd.n2876 vdd.n904 185
R18389 vdd.n2783 vdd.n2782 185
R18390 vdd.n2782 vdd.n2781 185
R18391 vdd.n2784 vdd.n909 185
R18392 vdd.n2870 vdd.n909 185
R18393 vdd.n2786 vdd.n2785 185
R18394 vdd.n2785 vdd.t147 185
R18395 vdd.n2787 vdd.n914 185
R18396 vdd.n2864 vdd.n914 185
R18397 vdd.n2866 vdd.n2865 185
R18398 vdd.n2865 vdd.n2864 185
R18399 vdd.n2867 vdd.n911 185
R18400 vdd.n911 vdd.t147 185
R18401 vdd.n2869 vdd.n2868 185
R18402 vdd.n2870 vdd.n2869 185
R18403 vdd.n903 vdd.n902 185
R18404 vdd.n2781 vdd.n903 185
R18405 vdd.n2878 vdd.n2877 185
R18406 vdd.n2877 vdd.n2876 185
R18407 vdd.n2879 vdd.n901 185
R18408 vdd.n901 vdd.n897 185
R18409 vdd.n2881 vdd.n2880 185
R18410 vdd.n2882 vdd.n2881 185
R18411 vdd.n890 vdd.n889 185
R18412 vdd.n900 vdd.n890 185
R18413 vdd.n2890 vdd.n2889 185
R18414 vdd.n2889 vdd.n2888 185
R18415 vdd.n2891 vdd.n888 185
R18416 vdd.n893 vdd.n888 185
R18417 vdd.n2893 vdd.n2892 185
R18418 vdd.n2894 vdd.n2893 185
R18419 vdd.n879 vdd.n878 185
R18420 vdd.n880 vdd.n879 185
R18421 vdd.n2902 vdd.n2901 185
R18422 vdd.n2901 vdd.n2900 185
R18423 vdd.n2903 vdd.n877 185
R18424 vdd.n877 vdd.n874 185
R18425 vdd.n2905 vdd.n2904 185
R18426 vdd.n2906 vdd.n2905 185
R18427 vdd.n867 vdd.n866 185
R18428 vdd.n2760 vdd.n867 185
R18429 vdd.n2914 vdd.n2913 185
R18430 vdd.n2913 vdd.n2912 185
R18431 vdd.n2915 vdd.n865 185
R18432 vdd.n870 vdd.n865 185
R18433 vdd.n2917 vdd.n2916 185
R18434 vdd.n2918 vdd.n2917 185
R18435 vdd.n856 vdd.n855 185
R18436 vdd.n857 vdd.n856 185
R18437 vdd.n2928 vdd.n2927 185
R18438 vdd.n2927 vdd.n2926 185
R18439 vdd.n2929 vdd.n854 185
R18440 vdd.n854 vdd.n851 185
R18441 vdd.n2931 vdd.n2930 185
R18442 vdd.n2932 vdd.n2931 185
R18443 vdd.n842 vdd.n841 185
R18444 vdd.n843 vdd.n842 185
R18445 vdd.n2985 vdd.n2984 185
R18446 vdd.n2984 vdd.n2983 185
R18447 vdd.n2986 vdd.n840 185
R18448 vdd.n846 vdd.n840 185
R18449 vdd.n2988 vdd.n2987 185
R18450 vdd.n2989 vdd.n2988 185
R18451 vdd.n810 vdd.n808 185
R18452 vdd.n808 vdd.n805 185
R18453 vdd.n3058 vdd.n3057 185
R18454 vdd.n3059 vdd.n3058 185
R18455 vdd.n2531 vdd.n2530 185
R18456 vdd.n2532 vdd.n2531 185
R18457 vdd.n964 vdd.n962 185
R18458 vdd.n962 vdd.t159 185
R18459 vdd.n2446 vdd.n971 185
R18460 vdd.n2457 vdd.n971 185
R18461 vdd.n2447 vdd.n980 185
R18462 vdd.n2156 vdd.n980 185
R18463 vdd.n2449 vdd.n2448 185
R18464 vdd.n2450 vdd.n2449 185
R18465 vdd.n2445 vdd.n979 185
R18466 vdd.n979 vdd.n976 185
R18467 vdd.n2444 vdd.n2443 185
R18468 vdd.n2443 vdd.n2442 185
R18469 vdd.n982 vdd.n981 185
R18470 vdd.n983 vdd.n982 185
R18471 vdd.n2435 vdd.n2434 185
R18472 vdd.n2436 vdd.n2435 185
R18473 vdd.n2433 vdd.n992 185
R18474 vdd.n992 vdd.n989 185
R18475 vdd.n2432 vdd.n2431 185
R18476 vdd.n2431 vdd.n2430 185
R18477 vdd.n994 vdd.n993 185
R18478 vdd.n1002 vdd.n994 185
R18479 vdd.n2423 vdd.n2422 185
R18480 vdd.n2424 vdd.n2423 185
R18481 vdd.n2421 vdd.n1003 185
R18482 vdd.n1008 vdd.n1003 185
R18483 vdd.n2420 vdd.n2419 185
R18484 vdd.n2419 vdd.n2418 185
R18485 vdd.n1005 vdd.n1004 185
R18486 vdd.n2257 vdd.n1005 185
R18487 vdd.n2411 vdd.n2410 185
R18488 vdd.n2412 vdd.n2411 185
R18489 vdd.n2409 vdd.n1015 185
R18490 vdd.n1015 vdd.n1012 185
R18491 vdd.n2408 vdd.n2407 185
R18492 vdd.n2407 vdd.n2406 185
R18493 vdd.n1017 vdd.n1016 185
R18494 vdd.n1018 vdd.n1017 185
R18495 vdd.n2399 vdd.n2398 185
R18496 vdd.n2400 vdd.n2399 185
R18497 vdd.n2396 vdd.n1026 185
R18498 vdd.n1033 vdd.n1026 185
R18499 vdd.n2395 vdd.n2394 185
R18500 vdd.n2394 vdd.n2393 185
R18501 vdd.n1029 vdd.n1028 185
R18502 vdd.n1030 vdd.n1029 185
R18503 vdd.n2386 vdd.n2385 185
R18504 vdd.n2387 vdd.n2386 185
R18505 vdd.n2384 vdd.n1040 185
R18506 vdd.n1040 vdd.n1037 185
R18507 vdd.n2383 vdd.n2382 185
R18508 vdd.n2382 vdd.n2381 185
R18509 vdd.n1042 vdd.n1041 185
R18510 vdd.n1043 vdd.n1042 185
R18511 vdd.n2374 vdd.n2373 185
R18512 vdd.n2375 vdd.n2374 185
R18513 vdd.n2462 vdd.n936 185
R18514 vdd.n2604 vdd.n936 185
R18515 vdd.n2464 vdd.n2463 185
R18516 vdd.n2466 vdd.n2465 185
R18517 vdd.n2468 vdd.n2467 185
R18518 vdd.n2470 vdd.n2469 185
R18519 vdd.n2472 vdd.n2471 185
R18520 vdd.n2474 vdd.n2473 185
R18521 vdd.n2476 vdd.n2475 185
R18522 vdd.n2478 vdd.n2477 185
R18523 vdd.n2480 vdd.n2479 185
R18524 vdd.n2482 vdd.n2481 185
R18525 vdd.n2484 vdd.n2483 185
R18526 vdd.n2486 vdd.n2485 185
R18527 vdd.n2488 vdd.n2487 185
R18528 vdd.n2490 vdd.n2489 185
R18529 vdd.n2492 vdd.n2491 185
R18530 vdd.n2494 vdd.n2493 185
R18531 vdd.n2496 vdd.n2495 185
R18532 vdd.n2498 vdd.n2497 185
R18533 vdd.n2500 vdd.n2499 185
R18534 vdd.n2502 vdd.n2501 185
R18535 vdd.n2504 vdd.n2503 185
R18536 vdd.n2506 vdd.n2505 185
R18537 vdd.n2508 vdd.n2507 185
R18538 vdd.n2510 vdd.n2509 185
R18539 vdd.n2512 vdd.n2511 185
R18540 vdd.n2514 vdd.n2513 185
R18541 vdd.n2516 vdd.n2515 185
R18542 vdd.n2518 vdd.n2517 185
R18543 vdd.n2520 vdd.n2519 185
R18544 vdd.n2522 vdd.n2521 185
R18545 vdd.n2524 vdd.n2523 185
R18546 vdd.n2526 vdd.n2525 185
R18547 vdd.n2528 vdd.n2527 185
R18548 vdd.n2529 vdd.n963 185
R18549 vdd.n2461 vdd.n961 185
R18550 vdd.n2532 vdd.n961 185
R18551 vdd.n2460 vdd.n2459 185
R18552 vdd.n2459 vdd.t159 185
R18553 vdd.n2458 vdd.n968 185
R18554 vdd.n2458 vdd.n2457 185
R18555 vdd.n2238 vdd.n969 185
R18556 vdd.n2156 vdd.n969 185
R18557 vdd.n2239 vdd.n978 185
R18558 vdd.n2450 vdd.n978 185
R18559 vdd.n2241 vdd.n2240 185
R18560 vdd.n2240 vdd.n976 185
R18561 vdd.n2242 vdd.n985 185
R18562 vdd.n2442 vdd.n985 185
R18563 vdd.n2244 vdd.n2243 185
R18564 vdd.n2243 vdd.n983 185
R18565 vdd.n2245 vdd.n991 185
R18566 vdd.n2436 vdd.n991 185
R18567 vdd.n2247 vdd.n2246 185
R18568 vdd.n2246 vdd.n989 185
R18569 vdd.n2248 vdd.n996 185
R18570 vdd.n2430 vdd.n996 185
R18571 vdd.n2250 vdd.n2249 185
R18572 vdd.n2249 vdd.n1002 185
R18573 vdd.n2251 vdd.n1001 185
R18574 vdd.n2424 vdd.n1001 185
R18575 vdd.n2253 vdd.n2252 185
R18576 vdd.n2252 vdd.n1008 185
R18577 vdd.n2254 vdd.n1007 185
R18578 vdd.n2418 vdd.n1007 185
R18579 vdd.n2256 vdd.n2255 185
R18580 vdd.n2257 vdd.n2256 185
R18581 vdd.n2237 vdd.n1014 185
R18582 vdd.n2412 vdd.n1014 185
R18583 vdd.n2236 vdd.n2235 185
R18584 vdd.n2235 vdd.n1012 185
R18585 vdd.n2234 vdd.n1020 185
R18586 vdd.n2406 vdd.n1020 185
R18587 vdd.n2233 vdd.n2232 185
R18588 vdd.n2232 vdd.n1018 185
R18589 vdd.n2231 vdd.n1025 185
R18590 vdd.n2400 vdd.n1025 185
R18591 vdd.n2230 vdd.n2229 185
R18592 vdd.n2229 vdd.n1033 185
R18593 vdd.n2228 vdd.n1032 185
R18594 vdd.n2393 vdd.n1032 185
R18595 vdd.n2227 vdd.n2226 185
R18596 vdd.n2226 vdd.n1030 185
R18597 vdd.n2225 vdd.n1039 185
R18598 vdd.n2387 vdd.n1039 185
R18599 vdd.n2224 vdd.n2223 185
R18600 vdd.n2223 vdd.n1037 185
R18601 vdd.n2222 vdd.n1045 185
R18602 vdd.n2381 vdd.n1045 185
R18603 vdd.n2221 vdd.n2220 185
R18604 vdd.n2220 vdd.n1043 185
R18605 vdd.n2219 vdd.n1051 185
R18606 vdd.n2375 vdd.n1051 185
R18607 vdd.n2372 vdd.n1052 185
R18608 vdd.n2371 vdd.n2370 185
R18609 vdd.n2368 vdd.n1053 185
R18610 vdd.n2366 vdd.n2365 185
R18611 vdd.n2364 vdd.n1054 185
R18612 vdd.n2363 vdd.n2362 185
R18613 vdd.n2360 vdd.n1055 185
R18614 vdd.n2358 vdd.n2357 185
R18615 vdd.n2356 vdd.n1056 185
R18616 vdd.n2355 vdd.n2354 185
R18617 vdd.n2352 vdd.n1057 185
R18618 vdd.n2350 vdd.n2349 185
R18619 vdd.n2348 vdd.n1058 185
R18620 vdd.n2347 vdd.n2346 185
R18621 vdd.n2344 vdd.n1059 185
R18622 vdd.n2342 vdd.n2341 185
R18623 vdd.n2340 vdd.n1060 185
R18624 vdd.n2339 vdd.n1062 185
R18625 vdd.n2184 vdd.n1063 185
R18626 vdd.n2187 vdd.n2186 185
R18627 vdd.n2189 vdd.n2188 185
R18628 vdd.n2191 vdd.n2183 185
R18629 vdd.n2194 vdd.n2193 185
R18630 vdd.n2195 vdd.n2182 185
R18631 vdd.n2197 vdd.n2196 185
R18632 vdd.n2199 vdd.n2181 185
R18633 vdd.n2202 vdd.n2201 185
R18634 vdd.n2203 vdd.n2180 185
R18635 vdd.n2205 vdd.n2204 185
R18636 vdd.n2207 vdd.n2179 185
R18637 vdd.n2210 vdd.n2209 185
R18638 vdd.n2211 vdd.n2176 185
R18639 vdd.n2214 vdd.n2213 185
R18640 vdd.n2216 vdd.n2175 185
R18641 vdd.n2218 vdd.n2217 185
R18642 vdd.n2217 vdd.n1049 185
R18643 vdd.n327 vdd.n326 171.744
R18644 vdd.n326 vdd.n325 171.744
R18645 vdd.n325 vdd.n294 171.744
R18646 vdd.n318 vdd.n294 171.744
R18647 vdd.n318 vdd.n317 171.744
R18648 vdd.n317 vdd.n299 171.744
R18649 vdd.n310 vdd.n299 171.744
R18650 vdd.n310 vdd.n309 171.744
R18651 vdd.n309 vdd.n303 171.744
R18652 vdd.n268 vdd.n267 171.744
R18653 vdd.n267 vdd.n266 171.744
R18654 vdd.n266 vdd.n235 171.744
R18655 vdd.n259 vdd.n235 171.744
R18656 vdd.n259 vdd.n258 171.744
R18657 vdd.n258 vdd.n240 171.744
R18658 vdd.n251 vdd.n240 171.744
R18659 vdd.n251 vdd.n250 171.744
R18660 vdd.n250 vdd.n244 171.744
R18661 vdd.n225 vdd.n224 171.744
R18662 vdd.n224 vdd.n223 171.744
R18663 vdd.n223 vdd.n192 171.744
R18664 vdd.n216 vdd.n192 171.744
R18665 vdd.n216 vdd.n215 171.744
R18666 vdd.n215 vdd.n197 171.744
R18667 vdd.n208 vdd.n197 171.744
R18668 vdd.n208 vdd.n207 171.744
R18669 vdd.n207 vdd.n201 171.744
R18670 vdd.n166 vdd.n165 171.744
R18671 vdd.n165 vdd.n164 171.744
R18672 vdd.n164 vdd.n133 171.744
R18673 vdd.n157 vdd.n133 171.744
R18674 vdd.n157 vdd.n156 171.744
R18675 vdd.n156 vdd.n138 171.744
R18676 vdd.n149 vdd.n138 171.744
R18677 vdd.n149 vdd.n148 171.744
R18678 vdd.n148 vdd.n142 171.744
R18679 vdd.n124 vdd.n123 171.744
R18680 vdd.n123 vdd.n122 171.744
R18681 vdd.n122 vdd.n91 171.744
R18682 vdd.n115 vdd.n91 171.744
R18683 vdd.n115 vdd.n114 171.744
R18684 vdd.n114 vdd.n96 171.744
R18685 vdd.n107 vdd.n96 171.744
R18686 vdd.n107 vdd.n106 171.744
R18687 vdd.n106 vdd.n100 171.744
R18688 vdd.n65 vdd.n64 171.744
R18689 vdd.n64 vdd.n63 171.744
R18690 vdd.n63 vdd.n32 171.744
R18691 vdd.n56 vdd.n32 171.744
R18692 vdd.n56 vdd.n55 171.744
R18693 vdd.n55 vdd.n37 171.744
R18694 vdd.n48 vdd.n37 171.744
R18695 vdd.n48 vdd.n47 171.744
R18696 vdd.n47 vdd.n41 171.744
R18697 vdd.n1746 vdd.n1745 171.744
R18698 vdd.n1745 vdd.n1744 171.744
R18699 vdd.n1744 vdd.n1713 171.744
R18700 vdd.n1737 vdd.n1713 171.744
R18701 vdd.n1737 vdd.n1736 171.744
R18702 vdd.n1736 vdd.n1718 171.744
R18703 vdd.n1729 vdd.n1718 171.744
R18704 vdd.n1729 vdd.n1728 171.744
R18705 vdd.n1728 vdd.n1722 171.744
R18706 vdd.n1805 vdd.n1804 171.744
R18707 vdd.n1804 vdd.n1803 171.744
R18708 vdd.n1803 vdd.n1772 171.744
R18709 vdd.n1796 vdd.n1772 171.744
R18710 vdd.n1796 vdd.n1795 171.744
R18711 vdd.n1795 vdd.n1777 171.744
R18712 vdd.n1788 vdd.n1777 171.744
R18713 vdd.n1788 vdd.n1787 171.744
R18714 vdd.n1787 vdd.n1781 171.744
R18715 vdd.n1644 vdd.n1643 171.744
R18716 vdd.n1643 vdd.n1642 171.744
R18717 vdd.n1642 vdd.n1611 171.744
R18718 vdd.n1635 vdd.n1611 171.744
R18719 vdd.n1635 vdd.n1634 171.744
R18720 vdd.n1634 vdd.n1616 171.744
R18721 vdd.n1627 vdd.n1616 171.744
R18722 vdd.n1627 vdd.n1626 171.744
R18723 vdd.n1626 vdd.n1620 171.744
R18724 vdd.n1703 vdd.n1702 171.744
R18725 vdd.n1702 vdd.n1701 171.744
R18726 vdd.n1701 vdd.n1670 171.744
R18727 vdd.n1694 vdd.n1670 171.744
R18728 vdd.n1694 vdd.n1693 171.744
R18729 vdd.n1693 vdd.n1675 171.744
R18730 vdd.n1686 vdd.n1675 171.744
R18731 vdd.n1686 vdd.n1685 171.744
R18732 vdd.n1685 vdd.n1679 171.744
R18733 vdd.n1543 vdd.n1542 171.744
R18734 vdd.n1542 vdd.n1541 171.744
R18735 vdd.n1541 vdd.n1510 171.744
R18736 vdd.n1534 vdd.n1510 171.744
R18737 vdd.n1534 vdd.n1533 171.744
R18738 vdd.n1533 vdd.n1515 171.744
R18739 vdd.n1526 vdd.n1515 171.744
R18740 vdd.n1526 vdd.n1525 171.744
R18741 vdd.n1525 vdd.n1519 171.744
R18742 vdd.n1602 vdd.n1601 171.744
R18743 vdd.n1601 vdd.n1600 171.744
R18744 vdd.n1600 vdd.n1569 171.744
R18745 vdd.n1593 vdd.n1569 171.744
R18746 vdd.n1593 vdd.n1592 171.744
R18747 vdd.n1592 vdd.n1574 171.744
R18748 vdd.n1585 vdd.n1574 171.744
R18749 vdd.n1585 vdd.n1584 171.744
R18750 vdd.n1584 vdd.n1578 171.744
R18751 vdd.n468 vdd.n467 146.341
R18752 vdd.n474 vdd.n473 146.341
R18753 vdd.n478 vdd.n477 146.341
R18754 vdd.n484 vdd.n483 146.341
R18755 vdd.n488 vdd.n487 146.341
R18756 vdd.n494 vdd.n493 146.341
R18757 vdd.n498 vdd.n497 146.341
R18758 vdd.n504 vdd.n503 146.341
R18759 vdd.n508 vdd.n507 146.341
R18760 vdd.n514 vdd.n513 146.341
R18761 vdd.n518 vdd.n517 146.341
R18762 vdd.n524 vdd.n523 146.341
R18763 vdd.n528 vdd.n527 146.341
R18764 vdd.n534 vdd.n533 146.341
R18765 vdd.n538 vdd.n537 146.341
R18766 vdd.n544 vdd.n543 146.341
R18767 vdd.n548 vdd.n547 146.341
R18768 vdd.n554 vdd.n553 146.341
R18769 vdd.n558 vdd.n557 146.341
R18770 vdd.n564 vdd.n563 146.341
R18771 vdd.n568 vdd.n567 146.341
R18772 vdd.n574 vdd.n573 146.341
R18773 vdd.n578 vdd.n577 146.341
R18774 vdd.n584 vdd.n583 146.341
R18775 vdd.n588 vdd.n587 146.341
R18776 vdd.n594 vdd.n593 146.341
R18777 vdd.n598 vdd.n597 146.341
R18778 vdd.n604 vdd.n603 146.341
R18779 vdd.n608 vdd.n607 146.341
R18780 vdd.n614 vdd.n613 146.341
R18781 vdd.n616 vdd.n425 146.341
R18782 vdd.n3230 vdd.n685 146.341
R18783 vdd.n3230 vdd.n677 146.341
R18784 vdd.n3240 vdd.n677 146.341
R18785 vdd.n3240 vdd.n673 146.341
R18786 vdd.n3246 vdd.n673 146.341
R18787 vdd.n3246 vdd.n667 146.341
R18788 vdd.n3257 vdd.n667 146.341
R18789 vdd.n3257 vdd.n663 146.341
R18790 vdd.n3263 vdd.n663 146.341
R18791 vdd.n3263 vdd.n654 146.341
R18792 vdd.n3273 vdd.n654 146.341
R18793 vdd.n3273 vdd.n650 146.341
R18794 vdd.n3279 vdd.n650 146.341
R18795 vdd.n3279 vdd.n643 146.341
R18796 vdd.n3290 vdd.n643 146.341
R18797 vdd.n3290 vdd.n639 146.341
R18798 vdd.n3299 vdd.n639 146.341
R18799 vdd.n3299 vdd.n632 146.341
R18800 vdd.n3309 vdd.n632 146.341
R18801 vdd.n3310 vdd.n3309 146.341
R18802 vdd.n3310 vdd.n341 146.341
R18803 vdd.n342 vdd.n341 146.341
R18804 vdd.n343 vdd.n342 146.341
R18805 vdd.n3317 vdd.n343 146.341
R18806 vdd.n3317 vdd.n351 146.341
R18807 vdd.n352 vdd.n351 146.341
R18808 vdd.n353 vdd.n352 146.341
R18809 vdd.n3324 vdd.n353 146.341
R18810 vdd.n3324 vdd.n362 146.341
R18811 vdd.n363 vdd.n362 146.341
R18812 vdd.n364 vdd.n363 146.341
R18813 vdd.n3332 vdd.n364 146.341
R18814 vdd.n3332 vdd.n372 146.341
R18815 vdd.n373 vdd.n372 146.341
R18816 vdd.n374 vdd.n373 146.341
R18817 vdd.n3339 vdd.n374 146.341
R18818 vdd.n3339 vdd.n383 146.341
R18819 vdd.n384 vdd.n383 146.341
R18820 vdd.n385 vdd.n384 146.341
R18821 vdd.n3346 vdd.n385 146.341
R18822 vdd.n3346 vdd.n393 146.341
R18823 vdd.n725 vdd.n724 146.341
R18824 vdd.n728 vdd.n724 146.341
R18825 vdd.n734 vdd.n733 146.341
R18826 vdd.n3212 vdd.n3211 146.341
R18827 vdd.n3208 vdd.n3207 146.341
R18828 vdd.n3204 vdd.n3203 146.341
R18829 vdd.n3200 vdd.n3199 146.341
R18830 vdd.n3196 vdd.n3195 146.341
R18831 vdd.n3192 vdd.n3191 146.341
R18832 vdd.n3188 vdd.n3187 146.341
R18833 vdd.n3179 vdd.n3178 146.341
R18834 vdd.n3176 vdd.n3175 146.341
R18835 vdd.n3172 vdd.n3171 146.341
R18836 vdd.n3168 vdd.n3167 146.341
R18837 vdd.n3164 vdd.n3163 146.341
R18838 vdd.n3160 vdd.n3159 146.341
R18839 vdd.n3156 vdd.n3155 146.341
R18840 vdd.n3152 vdd.n3151 146.341
R18841 vdd.n3148 vdd.n3147 146.341
R18842 vdd.n3144 vdd.n3143 146.341
R18843 vdd.n3140 vdd.n3139 146.341
R18844 vdd.n3133 vdd.n3132 146.341
R18845 vdd.n3130 vdd.n3129 146.341
R18846 vdd.n3126 vdd.n3125 146.341
R18847 vdd.n3122 vdd.n3121 146.341
R18848 vdd.n3118 vdd.n3117 146.341
R18849 vdd.n3114 vdd.n3113 146.341
R18850 vdd.n3110 vdd.n3109 146.341
R18851 vdd.n3106 vdd.n3105 146.341
R18852 vdd.n3102 vdd.n3101 146.341
R18853 vdd.n3098 vdd.n3097 146.341
R18854 vdd.n3224 vdd.n691 146.341
R18855 vdd.n3232 vdd.n684 146.341
R18856 vdd.n3232 vdd.n680 146.341
R18857 vdd.n3238 vdd.n680 146.341
R18858 vdd.n3238 vdd.n672 146.341
R18859 vdd.n3249 vdd.n672 146.341
R18860 vdd.n3249 vdd.n668 146.341
R18861 vdd.n3255 vdd.n668 146.341
R18862 vdd.n3255 vdd.n661 146.341
R18863 vdd.n3265 vdd.n661 146.341
R18864 vdd.n3265 vdd.n657 146.341
R18865 vdd.n3271 vdd.n657 146.341
R18866 vdd.n3271 vdd.n649 146.341
R18867 vdd.n3282 vdd.n649 146.341
R18868 vdd.n3282 vdd.n645 146.341
R18869 vdd.n3288 vdd.n645 146.341
R18870 vdd.n3288 vdd.n638 146.341
R18871 vdd.n3301 vdd.n638 146.341
R18872 vdd.n3301 vdd.n634 146.341
R18873 vdd.n3307 vdd.n634 146.341
R18874 vdd.n3307 vdd.n338 146.341
R18875 vdd.n3396 vdd.n338 146.341
R18876 vdd.n3396 vdd.n339 146.341
R18877 vdd.n3392 vdd.n339 146.341
R18878 vdd.n3392 vdd.n345 146.341
R18879 vdd.n3388 vdd.n345 146.341
R18880 vdd.n3388 vdd.n350 146.341
R18881 vdd.n3384 vdd.n350 146.341
R18882 vdd.n3384 vdd.n354 146.341
R18883 vdd.n3380 vdd.n354 146.341
R18884 vdd.n3380 vdd.n360 146.341
R18885 vdd.n3376 vdd.n360 146.341
R18886 vdd.n3376 vdd.n365 146.341
R18887 vdd.n3372 vdd.n365 146.341
R18888 vdd.n3372 vdd.n371 146.341
R18889 vdd.n3368 vdd.n371 146.341
R18890 vdd.n3368 vdd.n376 146.341
R18891 vdd.n3364 vdd.n376 146.341
R18892 vdd.n3364 vdd.n382 146.341
R18893 vdd.n3360 vdd.n382 146.341
R18894 vdd.n3360 vdd.n387 146.341
R18895 vdd.n3356 vdd.n387 146.341
R18896 vdd.n2322 vdd.n2321 146.341
R18897 vdd.n2319 vdd.n1903 146.341
R18898 vdd.n2099 vdd.n1909 146.341
R18899 vdd.n2097 vdd.n2096 146.341
R18900 vdd.n2094 vdd.n1911 146.341
R18901 vdd.n2090 vdd.n2089 146.341
R18902 vdd.n2087 vdd.n1918 146.341
R18903 vdd.n2083 vdd.n2082 146.341
R18904 vdd.n2080 vdd.n1925 146.341
R18905 vdd.n1936 vdd.n1933 146.341
R18906 vdd.n2072 vdd.n2071 146.341
R18907 vdd.n2069 vdd.n1938 146.341
R18908 vdd.n2065 vdd.n2064 146.341
R18909 vdd.n2062 vdd.n1944 146.341
R18910 vdd.n2058 vdd.n2057 146.341
R18911 vdd.n2055 vdd.n1951 146.341
R18912 vdd.n2051 vdd.n2050 146.341
R18913 vdd.n2048 vdd.n1958 146.341
R18914 vdd.n2044 vdd.n2043 146.341
R18915 vdd.n2041 vdd.n1965 146.341
R18916 vdd.n1976 vdd.n1973 146.341
R18917 vdd.n2033 vdd.n2032 146.341
R18918 vdd.n2030 vdd.n1978 146.341
R18919 vdd.n2026 vdd.n2025 146.341
R18920 vdd.n2023 vdd.n1984 146.341
R18921 vdd.n2019 vdd.n2018 146.341
R18922 vdd.n2016 vdd.n1991 146.341
R18923 vdd.n2012 vdd.n2011 146.341
R18924 vdd.n2009 vdd.n2006 146.341
R18925 vdd.n2004 vdd.n2001 146.341
R18926 vdd.n1999 vdd.n1069 146.341
R18927 vdd.n1428 vdd.n1188 146.341
R18928 vdd.n1428 vdd.n1184 146.341
R18929 vdd.n1434 vdd.n1184 146.341
R18930 vdd.n1434 vdd.n1176 146.341
R18931 vdd.n1445 vdd.n1176 146.341
R18932 vdd.n1445 vdd.n1172 146.341
R18933 vdd.n1451 vdd.n1172 146.341
R18934 vdd.n1451 vdd.n1166 146.341
R18935 vdd.n1462 vdd.n1166 146.341
R18936 vdd.n1462 vdd.n1162 146.341
R18937 vdd.n1468 vdd.n1162 146.341
R18938 vdd.n1468 vdd.n1153 146.341
R18939 vdd.n1478 vdd.n1153 146.341
R18940 vdd.n1478 vdd.n1149 146.341
R18941 vdd.n1484 vdd.n1149 146.341
R18942 vdd.n1484 vdd.n1142 146.341
R18943 vdd.n1495 vdd.n1142 146.341
R18944 vdd.n1495 vdd.n1138 146.341
R18945 vdd.n1501 vdd.n1138 146.341
R18946 vdd.n1501 vdd.n1131 146.341
R18947 vdd.n1818 vdd.n1131 146.341
R18948 vdd.n1818 vdd.n1127 146.341
R18949 vdd.n1824 vdd.n1127 146.341
R18950 vdd.n1824 vdd.n1119 146.341
R18951 vdd.n1835 vdd.n1119 146.341
R18952 vdd.n1835 vdd.n1115 146.341
R18953 vdd.n1841 vdd.n1115 146.341
R18954 vdd.n1841 vdd.n1109 146.341
R18955 vdd.n1852 vdd.n1109 146.341
R18956 vdd.n1852 vdd.n1105 146.341
R18957 vdd.n1858 vdd.n1105 146.341
R18958 vdd.n1858 vdd.n1096 146.341
R18959 vdd.n1868 vdd.n1096 146.341
R18960 vdd.n1868 vdd.n1092 146.341
R18961 vdd.n1874 vdd.n1092 146.341
R18962 vdd.n1874 vdd.n1086 146.341
R18963 vdd.n1885 vdd.n1086 146.341
R18964 vdd.n1885 vdd.n1081 146.341
R18965 vdd.n1893 vdd.n1081 146.341
R18966 vdd.n1893 vdd.n1071 146.341
R18967 vdd.n2330 vdd.n1071 146.341
R18968 vdd.n1417 vdd.n1193 146.341
R18969 vdd.n1417 vdd.n1226 146.341
R18970 vdd.n1230 vdd.n1229 146.341
R18971 vdd.n1232 vdd.n1231 146.341
R18972 vdd.n1236 vdd.n1235 146.341
R18973 vdd.n1238 vdd.n1237 146.341
R18974 vdd.n1242 vdd.n1241 146.341
R18975 vdd.n1244 vdd.n1243 146.341
R18976 vdd.n1248 vdd.n1247 146.341
R18977 vdd.n1250 vdd.n1249 146.341
R18978 vdd.n1256 vdd.n1255 146.341
R18979 vdd.n1258 vdd.n1257 146.341
R18980 vdd.n1262 vdd.n1261 146.341
R18981 vdd.n1264 vdd.n1263 146.341
R18982 vdd.n1268 vdd.n1267 146.341
R18983 vdd.n1270 vdd.n1269 146.341
R18984 vdd.n1274 vdd.n1273 146.341
R18985 vdd.n1276 vdd.n1275 146.341
R18986 vdd.n1280 vdd.n1279 146.341
R18987 vdd.n1282 vdd.n1281 146.341
R18988 vdd.n1354 vdd.n1285 146.341
R18989 vdd.n1287 vdd.n1286 146.341
R18990 vdd.n1291 vdd.n1290 146.341
R18991 vdd.n1293 vdd.n1292 146.341
R18992 vdd.n1297 vdd.n1296 146.341
R18993 vdd.n1299 vdd.n1298 146.341
R18994 vdd.n1303 vdd.n1302 146.341
R18995 vdd.n1305 vdd.n1304 146.341
R18996 vdd.n1309 vdd.n1308 146.341
R18997 vdd.n1311 vdd.n1310 146.341
R18998 vdd.n1315 vdd.n1314 146.341
R18999 vdd.n1316 vdd.n1224 146.341
R19000 vdd.n1426 vdd.n1189 146.341
R19001 vdd.n1426 vdd.n1182 146.341
R19002 vdd.n1437 vdd.n1182 146.341
R19003 vdd.n1437 vdd.n1178 146.341
R19004 vdd.n1443 vdd.n1178 146.341
R19005 vdd.n1443 vdd.n1171 146.341
R19006 vdd.n1454 vdd.n1171 146.341
R19007 vdd.n1454 vdd.n1167 146.341
R19008 vdd.n1460 vdd.n1167 146.341
R19009 vdd.n1460 vdd.n1160 146.341
R19010 vdd.n1470 vdd.n1160 146.341
R19011 vdd.n1470 vdd.n1156 146.341
R19012 vdd.n1476 vdd.n1156 146.341
R19013 vdd.n1476 vdd.n1148 146.341
R19014 vdd.n1487 vdd.n1148 146.341
R19015 vdd.n1487 vdd.n1144 146.341
R19016 vdd.n1493 vdd.n1144 146.341
R19017 vdd.n1493 vdd.n1137 146.341
R19018 vdd.n1503 vdd.n1137 146.341
R19019 vdd.n1503 vdd.n1133 146.341
R19020 vdd.n1816 vdd.n1133 146.341
R19021 vdd.n1816 vdd.n1125 146.341
R19022 vdd.n1827 vdd.n1125 146.341
R19023 vdd.n1827 vdd.n1121 146.341
R19024 vdd.n1833 vdd.n1121 146.341
R19025 vdd.n1833 vdd.n1114 146.341
R19026 vdd.n1844 vdd.n1114 146.341
R19027 vdd.n1844 vdd.n1110 146.341
R19028 vdd.n1850 vdd.n1110 146.341
R19029 vdd.n1850 vdd.n1103 146.341
R19030 vdd.n1860 vdd.n1103 146.341
R19031 vdd.n1860 vdd.n1099 146.341
R19032 vdd.n1866 vdd.n1099 146.341
R19033 vdd.n1866 vdd.n1091 146.341
R19034 vdd.n1877 vdd.n1091 146.341
R19035 vdd.n1877 vdd.n1087 146.341
R19036 vdd.n1883 vdd.n1087 146.341
R19037 vdd.n1883 vdd.n1079 146.341
R19038 vdd.n1896 vdd.n1079 146.341
R19039 vdd.n1896 vdd.n1074 146.341
R19040 vdd.n2328 vdd.n1074 146.341
R19041 vdd.n1073 vdd.n1049 141.707
R19042 vdd.n3223 vdd.n692 141.707
R19043 vdd.n2177 vdd.t222 127.284
R19044 vdd.n965 vdd.t206 127.284
R19045 vdd.n2151 vdd.t244 127.284
R19046 vdd.n957 vdd.t231 127.284
R19047 vdd.n2922 vdd.t182 127.284
R19048 vdd.n2922 vdd.t183 127.284
R19049 vdd.n2642 vdd.t229 127.284
R19050 vdd.n832 vdd.t210 127.284
R19051 vdd.n2639 vdd.t215 127.284
R19052 vdd.n799 vdd.t217 127.284
R19053 vdd.n1027 vdd.t225 127.284
R19054 vdd.n1027 vdd.t226 127.284
R19055 vdd.n22 vdd.n20 117.314
R19056 vdd.n17 vdd.n15 117.314
R19057 vdd.n27 vdd.n26 116.927
R19058 vdd.n24 vdd.n23 116.927
R19059 vdd.n22 vdd.n21 116.927
R19060 vdd.n17 vdd.n16 116.927
R19061 vdd.n19 vdd.n18 116.927
R19062 vdd.n27 vdd.n25 116.927
R19063 vdd.n2178 vdd.t221 111.188
R19064 vdd.n966 vdd.t207 111.188
R19065 vdd.n2152 vdd.t243 111.188
R19066 vdd.n958 vdd.t232 111.188
R19067 vdd.n2643 vdd.t228 111.188
R19068 vdd.n833 vdd.t211 111.188
R19069 vdd.n2640 vdd.t214 111.188
R19070 vdd.n800 vdd.t218 111.188
R19071 vdd.n2865 vdd.n911 99.5127
R19072 vdd.n2869 vdd.n911 99.5127
R19073 vdd.n2869 vdd.n903 99.5127
R19074 vdd.n2877 vdd.n903 99.5127
R19075 vdd.n2877 vdd.n901 99.5127
R19076 vdd.n2881 vdd.n901 99.5127
R19077 vdd.n2881 vdd.n890 99.5127
R19078 vdd.n2889 vdd.n890 99.5127
R19079 vdd.n2889 vdd.n888 99.5127
R19080 vdd.n2893 vdd.n888 99.5127
R19081 vdd.n2893 vdd.n879 99.5127
R19082 vdd.n2901 vdd.n879 99.5127
R19083 vdd.n2901 vdd.n877 99.5127
R19084 vdd.n2905 vdd.n877 99.5127
R19085 vdd.n2905 vdd.n867 99.5127
R19086 vdd.n2913 vdd.n867 99.5127
R19087 vdd.n2913 vdd.n865 99.5127
R19088 vdd.n2917 vdd.n865 99.5127
R19089 vdd.n2917 vdd.n856 99.5127
R19090 vdd.n2927 vdd.n856 99.5127
R19091 vdd.n2927 vdd.n854 99.5127
R19092 vdd.n2931 vdd.n854 99.5127
R19093 vdd.n2931 vdd.n842 99.5127
R19094 vdd.n2984 vdd.n842 99.5127
R19095 vdd.n2984 vdd.n840 99.5127
R19096 vdd.n2988 vdd.n840 99.5127
R19097 vdd.n2988 vdd.n808 99.5127
R19098 vdd.n3058 vdd.n808 99.5127
R19099 vdd.n3054 vdd.n809 99.5127
R19100 vdd.n3052 vdd.n3051 99.5127
R19101 vdd.n3049 vdd.n813 99.5127
R19102 vdd.n3045 vdd.n3044 99.5127
R19103 vdd.n3042 vdd.n816 99.5127
R19104 vdd.n3038 vdd.n3037 99.5127
R19105 vdd.n3035 vdd.n819 99.5127
R19106 vdd.n3031 vdd.n3030 99.5127
R19107 vdd.n3028 vdd.n3026 99.5127
R19108 vdd.n3024 vdd.n822 99.5127
R19109 vdd.n3020 vdd.n3019 99.5127
R19110 vdd.n3017 vdd.n825 99.5127
R19111 vdd.n3013 vdd.n3012 99.5127
R19112 vdd.n3010 vdd.n828 99.5127
R19113 vdd.n3006 vdd.n3005 99.5127
R19114 vdd.n3003 vdd.n831 99.5127
R19115 vdd.n2998 vdd.n2997 99.5127
R19116 vdd.n2785 vdd.n914 99.5127
R19117 vdd.n2785 vdd.n909 99.5127
R19118 vdd.n2782 vdd.n909 99.5127
R19119 vdd.n2782 vdd.n904 99.5127
R19120 vdd.n2729 vdd.n904 99.5127
R19121 vdd.n2729 vdd.n898 99.5127
R19122 vdd.n2732 vdd.n898 99.5127
R19123 vdd.n2732 vdd.n891 99.5127
R19124 vdd.n2735 vdd.n891 99.5127
R19125 vdd.n2735 vdd.n886 99.5127
R19126 vdd.n2738 vdd.n886 99.5127
R19127 vdd.n2738 vdd.n881 99.5127
R19128 vdd.n2741 vdd.n881 99.5127
R19129 vdd.n2741 vdd.n875 99.5127
R19130 vdd.n2759 vdd.n875 99.5127
R19131 vdd.n2759 vdd.n868 99.5127
R19132 vdd.n2755 vdd.n868 99.5127
R19133 vdd.n2755 vdd.n863 99.5127
R19134 vdd.n2752 vdd.n863 99.5127
R19135 vdd.n2752 vdd.n858 99.5127
R19136 vdd.n2749 vdd.n858 99.5127
R19137 vdd.n2749 vdd.n852 99.5127
R19138 vdd.n2746 vdd.n852 99.5127
R19139 vdd.n2746 vdd.n844 99.5127
R19140 vdd.n844 vdd.n837 99.5127
R19141 vdd.n2990 vdd.n837 99.5127
R19142 vdd.n2991 vdd.n2990 99.5127
R19143 vdd.n2991 vdd.n806 99.5127
R19144 vdd.n2855 vdd.n2638 99.5127
R19145 vdd.n2851 vdd.n2638 99.5127
R19146 vdd.n2849 vdd.n2848 99.5127
R19147 vdd.n2845 vdd.n2844 99.5127
R19148 vdd.n2841 vdd.n2840 99.5127
R19149 vdd.n2837 vdd.n2836 99.5127
R19150 vdd.n2833 vdd.n2832 99.5127
R19151 vdd.n2829 vdd.n2828 99.5127
R19152 vdd.n2825 vdd.n2824 99.5127
R19153 vdd.n2821 vdd.n2820 99.5127
R19154 vdd.n2817 vdd.n2816 99.5127
R19155 vdd.n2813 vdd.n2812 99.5127
R19156 vdd.n2809 vdd.n2808 99.5127
R19157 vdd.n2805 vdd.n2804 99.5127
R19158 vdd.n2801 vdd.n2800 99.5127
R19159 vdd.n2797 vdd.n2796 99.5127
R19160 vdd.n2792 vdd.n2791 99.5127
R19161 vdd.n2603 vdd.n955 99.5127
R19162 vdd.n2599 vdd.n2598 99.5127
R19163 vdd.n2595 vdd.n2594 99.5127
R19164 vdd.n2591 vdd.n2590 99.5127
R19165 vdd.n2587 vdd.n2586 99.5127
R19166 vdd.n2583 vdd.n2582 99.5127
R19167 vdd.n2579 vdd.n2578 99.5127
R19168 vdd.n2575 vdd.n2574 99.5127
R19169 vdd.n2571 vdd.n2570 99.5127
R19170 vdd.n2567 vdd.n2566 99.5127
R19171 vdd.n2563 vdd.n2562 99.5127
R19172 vdd.n2559 vdd.n2558 99.5127
R19173 vdd.n2555 vdd.n2554 99.5127
R19174 vdd.n2551 vdd.n2550 99.5127
R19175 vdd.n2547 vdd.n2546 99.5127
R19176 vdd.n2543 vdd.n2542 99.5127
R19177 vdd.n2538 vdd.n2537 99.5127
R19178 vdd.n2276 vdd.n1050 99.5127
R19179 vdd.n2276 vdd.n1044 99.5127
R19180 vdd.n2273 vdd.n1044 99.5127
R19181 vdd.n2273 vdd.n1038 99.5127
R19182 vdd.n2270 vdd.n1038 99.5127
R19183 vdd.n2270 vdd.n1031 99.5127
R19184 vdd.n2267 vdd.n1031 99.5127
R19185 vdd.n2267 vdd.n1024 99.5127
R19186 vdd.n2264 vdd.n1024 99.5127
R19187 vdd.n2264 vdd.n1019 99.5127
R19188 vdd.n2261 vdd.n1019 99.5127
R19189 vdd.n2261 vdd.n1013 99.5127
R19190 vdd.n2258 vdd.n1013 99.5127
R19191 vdd.n2258 vdd.n1006 99.5127
R19192 vdd.n2172 vdd.n1006 99.5127
R19193 vdd.n2172 vdd.n1000 99.5127
R19194 vdd.n2169 vdd.n1000 99.5127
R19195 vdd.n2169 vdd.n995 99.5127
R19196 vdd.n2166 vdd.n995 99.5127
R19197 vdd.n2166 vdd.n990 99.5127
R19198 vdd.n2163 vdd.n990 99.5127
R19199 vdd.n2163 vdd.n984 99.5127
R19200 vdd.n2160 vdd.n984 99.5127
R19201 vdd.n2160 vdd.n977 99.5127
R19202 vdd.n2157 vdd.n977 99.5127
R19203 vdd.n2157 vdd.n970 99.5127
R19204 vdd.n970 vdd.n960 99.5127
R19205 vdd.n2533 vdd.n960 99.5127
R19206 vdd.n2111 vdd.n2109 99.5127
R19207 vdd.n2115 vdd.n2109 99.5127
R19208 vdd.n2119 vdd.n2117 99.5127
R19209 vdd.n2123 vdd.n2107 99.5127
R19210 vdd.n2127 vdd.n2125 99.5127
R19211 vdd.n2131 vdd.n2105 99.5127
R19212 vdd.n2135 vdd.n2133 99.5127
R19213 vdd.n2139 vdd.n2103 99.5127
R19214 vdd.n2142 vdd.n2141 99.5127
R19215 vdd.n2312 vdd.n2310 99.5127
R19216 vdd.n2308 vdd.n2144 99.5127
R19217 vdd.n2304 vdd.n2302 99.5127
R19218 vdd.n2300 vdd.n2146 99.5127
R19219 vdd.n2296 vdd.n2294 99.5127
R19220 vdd.n2292 vdd.n2148 99.5127
R19221 vdd.n2288 vdd.n2286 99.5127
R19222 vdd.n2284 vdd.n2150 99.5127
R19223 vdd.n2376 vdd.n1046 99.5127
R19224 vdd.n2380 vdd.n1046 99.5127
R19225 vdd.n2380 vdd.n1036 99.5127
R19226 vdd.n2388 vdd.n1036 99.5127
R19227 vdd.n2388 vdd.n1034 99.5127
R19228 vdd.n2392 vdd.n1034 99.5127
R19229 vdd.n2392 vdd.n1023 99.5127
R19230 vdd.n2401 vdd.n1023 99.5127
R19231 vdd.n2401 vdd.n1021 99.5127
R19232 vdd.n2405 vdd.n1021 99.5127
R19233 vdd.n2405 vdd.n1011 99.5127
R19234 vdd.n2413 vdd.n1011 99.5127
R19235 vdd.n2413 vdd.n1009 99.5127
R19236 vdd.n2417 vdd.n1009 99.5127
R19237 vdd.n2417 vdd.n999 99.5127
R19238 vdd.n2425 vdd.n999 99.5127
R19239 vdd.n2425 vdd.n997 99.5127
R19240 vdd.n2429 vdd.n997 99.5127
R19241 vdd.n2429 vdd.n988 99.5127
R19242 vdd.n2437 vdd.n988 99.5127
R19243 vdd.n2437 vdd.n986 99.5127
R19244 vdd.n2441 vdd.n986 99.5127
R19245 vdd.n2441 vdd.n975 99.5127
R19246 vdd.n2451 vdd.n975 99.5127
R19247 vdd.n2451 vdd.n972 99.5127
R19248 vdd.n2456 vdd.n972 99.5127
R19249 vdd.n2456 vdd.n973 99.5127
R19250 vdd.n973 vdd.n954 99.5127
R19251 vdd.n2974 vdd.n2973 99.5127
R19252 vdd.n2971 vdd.n2937 99.5127
R19253 vdd.n2967 vdd.n2966 99.5127
R19254 vdd.n2964 vdd.n2940 99.5127
R19255 vdd.n2960 vdd.n2959 99.5127
R19256 vdd.n2957 vdd.n2943 99.5127
R19257 vdd.n2953 vdd.n2952 99.5127
R19258 vdd.n2950 vdd.n2947 99.5127
R19259 vdd.n3091 vdd.n787 99.5127
R19260 vdd.n3089 vdd.n3088 99.5127
R19261 vdd.n3086 vdd.n789 99.5127
R19262 vdd.n3082 vdd.n3081 99.5127
R19263 vdd.n3079 vdd.n792 99.5127
R19264 vdd.n3075 vdd.n3074 99.5127
R19265 vdd.n3072 vdd.n795 99.5127
R19266 vdd.n3068 vdd.n3067 99.5127
R19267 vdd.n3065 vdd.n798 99.5127
R19268 vdd.n2709 vdd.n915 99.5127
R19269 vdd.n2709 vdd.n910 99.5127
R19270 vdd.n2780 vdd.n910 99.5127
R19271 vdd.n2780 vdd.n905 99.5127
R19272 vdd.n2776 vdd.n905 99.5127
R19273 vdd.n2776 vdd.n899 99.5127
R19274 vdd.n2773 vdd.n899 99.5127
R19275 vdd.n2773 vdd.n892 99.5127
R19276 vdd.n2770 vdd.n892 99.5127
R19277 vdd.n2770 vdd.n887 99.5127
R19278 vdd.n2767 vdd.n887 99.5127
R19279 vdd.n2767 vdd.n882 99.5127
R19280 vdd.n2764 vdd.n882 99.5127
R19281 vdd.n2764 vdd.n876 99.5127
R19282 vdd.n2761 vdd.n876 99.5127
R19283 vdd.n2761 vdd.n869 99.5127
R19284 vdd.n2726 vdd.n869 99.5127
R19285 vdd.n2726 vdd.n864 99.5127
R19286 vdd.n2723 vdd.n864 99.5127
R19287 vdd.n2723 vdd.n859 99.5127
R19288 vdd.n2720 vdd.n859 99.5127
R19289 vdd.n2720 vdd.n853 99.5127
R19290 vdd.n2717 vdd.n853 99.5127
R19291 vdd.n2717 vdd.n845 99.5127
R19292 vdd.n2714 vdd.n845 99.5127
R19293 vdd.n2714 vdd.n838 99.5127
R19294 vdd.n838 vdd.n804 99.5127
R19295 vdd.n3060 vdd.n804 99.5127
R19296 vdd.n2859 vdd.n918 99.5127
R19297 vdd.n2647 vdd.n2646 99.5127
R19298 vdd.n2651 vdd.n2650 99.5127
R19299 vdd.n2655 vdd.n2654 99.5127
R19300 vdd.n2659 vdd.n2658 99.5127
R19301 vdd.n2663 vdd.n2662 99.5127
R19302 vdd.n2667 vdd.n2666 99.5127
R19303 vdd.n2671 vdd.n2670 99.5127
R19304 vdd.n2675 vdd.n2674 99.5127
R19305 vdd.n2679 vdd.n2678 99.5127
R19306 vdd.n2683 vdd.n2682 99.5127
R19307 vdd.n2687 vdd.n2686 99.5127
R19308 vdd.n2691 vdd.n2690 99.5127
R19309 vdd.n2695 vdd.n2694 99.5127
R19310 vdd.n2699 vdd.n2698 99.5127
R19311 vdd.n2703 vdd.n2702 99.5127
R19312 vdd.n2705 vdd.n2637 99.5127
R19313 vdd.n2863 vdd.n908 99.5127
R19314 vdd.n2871 vdd.n908 99.5127
R19315 vdd.n2871 vdd.n906 99.5127
R19316 vdd.n2875 vdd.n906 99.5127
R19317 vdd.n2875 vdd.n896 99.5127
R19318 vdd.n2883 vdd.n896 99.5127
R19319 vdd.n2883 vdd.n894 99.5127
R19320 vdd.n2887 vdd.n894 99.5127
R19321 vdd.n2887 vdd.n885 99.5127
R19322 vdd.n2895 vdd.n885 99.5127
R19323 vdd.n2895 vdd.n883 99.5127
R19324 vdd.n2899 vdd.n883 99.5127
R19325 vdd.n2899 vdd.n873 99.5127
R19326 vdd.n2907 vdd.n873 99.5127
R19327 vdd.n2907 vdd.n871 99.5127
R19328 vdd.n2911 vdd.n871 99.5127
R19329 vdd.n2911 vdd.n862 99.5127
R19330 vdd.n2919 vdd.n862 99.5127
R19331 vdd.n2919 vdd.n860 99.5127
R19332 vdd.n2925 vdd.n860 99.5127
R19333 vdd.n2925 vdd.n850 99.5127
R19334 vdd.n2933 vdd.n850 99.5127
R19335 vdd.n2933 vdd.n847 99.5127
R19336 vdd.n2982 vdd.n847 99.5127
R19337 vdd.n2982 vdd.n848 99.5127
R19338 vdd.n848 vdd.n839 99.5127
R19339 vdd.n2977 vdd.n839 99.5127
R19340 vdd.n2977 vdd.n807 99.5127
R19341 vdd.n2527 vdd.n2526 99.5127
R19342 vdd.n2523 vdd.n2522 99.5127
R19343 vdd.n2519 vdd.n2518 99.5127
R19344 vdd.n2515 vdd.n2514 99.5127
R19345 vdd.n2511 vdd.n2510 99.5127
R19346 vdd.n2507 vdd.n2506 99.5127
R19347 vdd.n2503 vdd.n2502 99.5127
R19348 vdd.n2499 vdd.n2498 99.5127
R19349 vdd.n2495 vdd.n2494 99.5127
R19350 vdd.n2491 vdd.n2490 99.5127
R19351 vdd.n2487 vdd.n2486 99.5127
R19352 vdd.n2483 vdd.n2482 99.5127
R19353 vdd.n2479 vdd.n2478 99.5127
R19354 vdd.n2475 vdd.n2474 99.5127
R19355 vdd.n2471 vdd.n2470 99.5127
R19356 vdd.n2467 vdd.n2466 99.5127
R19357 vdd.n2463 vdd.n936 99.5127
R19358 vdd.n2220 vdd.n1051 99.5127
R19359 vdd.n2220 vdd.n1045 99.5127
R19360 vdd.n2223 vdd.n1045 99.5127
R19361 vdd.n2223 vdd.n1039 99.5127
R19362 vdd.n2226 vdd.n1039 99.5127
R19363 vdd.n2226 vdd.n1032 99.5127
R19364 vdd.n2229 vdd.n1032 99.5127
R19365 vdd.n2229 vdd.n1025 99.5127
R19366 vdd.n2232 vdd.n1025 99.5127
R19367 vdd.n2232 vdd.n1020 99.5127
R19368 vdd.n2235 vdd.n1020 99.5127
R19369 vdd.n2235 vdd.n1014 99.5127
R19370 vdd.n2256 vdd.n1014 99.5127
R19371 vdd.n2256 vdd.n1007 99.5127
R19372 vdd.n2252 vdd.n1007 99.5127
R19373 vdd.n2252 vdd.n1001 99.5127
R19374 vdd.n2249 vdd.n1001 99.5127
R19375 vdd.n2249 vdd.n996 99.5127
R19376 vdd.n2246 vdd.n996 99.5127
R19377 vdd.n2246 vdd.n991 99.5127
R19378 vdd.n2243 vdd.n991 99.5127
R19379 vdd.n2243 vdd.n985 99.5127
R19380 vdd.n2240 vdd.n985 99.5127
R19381 vdd.n2240 vdd.n978 99.5127
R19382 vdd.n978 vdd.n969 99.5127
R19383 vdd.n2458 vdd.n969 99.5127
R19384 vdd.n2459 vdd.n2458 99.5127
R19385 vdd.n2459 vdd.n961 99.5127
R19386 vdd.n2370 vdd.n2368 99.5127
R19387 vdd.n2366 vdd.n1054 99.5127
R19388 vdd.n2362 vdd.n2360 99.5127
R19389 vdd.n2358 vdd.n1056 99.5127
R19390 vdd.n2354 vdd.n2352 99.5127
R19391 vdd.n2350 vdd.n1058 99.5127
R19392 vdd.n2346 vdd.n2344 99.5127
R19393 vdd.n2342 vdd.n1060 99.5127
R19394 vdd.n2184 vdd.n1062 99.5127
R19395 vdd.n2189 vdd.n2186 99.5127
R19396 vdd.n2193 vdd.n2191 99.5127
R19397 vdd.n2197 vdd.n2182 99.5127
R19398 vdd.n2201 vdd.n2199 99.5127
R19399 vdd.n2205 vdd.n2180 99.5127
R19400 vdd.n2209 vdd.n2207 99.5127
R19401 vdd.n2214 vdd.n2176 99.5127
R19402 vdd.n2217 vdd.n2216 99.5127
R19403 vdd.n2374 vdd.n1042 99.5127
R19404 vdd.n2382 vdd.n1042 99.5127
R19405 vdd.n2382 vdd.n1040 99.5127
R19406 vdd.n2386 vdd.n1040 99.5127
R19407 vdd.n2386 vdd.n1029 99.5127
R19408 vdd.n2394 vdd.n1029 99.5127
R19409 vdd.n2394 vdd.n1026 99.5127
R19410 vdd.n2399 vdd.n1026 99.5127
R19411 vdd.n2399 vdd.n1017 99.5127
R19412 vdd.n2407 vdd.n1017 99.5127
R19413 vdd.n2407 vdd.n1015 99.5127
R19414 vdd.n2411 vdd.n1015 99.5127
R19415 vdd.n2411 vdd.n1005 99.5127
R19416 vdd.n2419 vdd.n1005 99.5127
R19417 vdd.n2419 vdd.n1003 99.5127
R19418 vdd.n2423 vdd.n1003 99.5127
R19419 vdd.n2423 vdd.n994 99.5127
R19420 vdd.n2431 vdd.n994 99.5127
R19421 vdd.n2431 vdd.n992 99.5127
R19422 vdd.n2435 vdd.n992 99.5127
R19423 vdd.n2435 vdd.n982 99.5127
R19424 vdd.n2443 vdd.n982 99.5127
R19425 vdd.n2443 vdd.n979 99.5127
R19426 vdd.n2449 vdd.n979 99.5127
R19427 vdd.n2449 vdd.n980 99.5127
R19428 vdd.n980 vdd.n971 99.5127
R19429 vdd.n971 vdd.n962 99.5127
R19430 vdd.n2531 vdd.n962 99.5127
R19431 vdd.n9 vdd.n7 98.9633
R19432 vdd.n2 vdd.n0 98.9633
R19433 vdd.n9 vdd.n8 98.6055
R19434 vdd.n11 vdd.n10 98.6055
R19435 vdd.n13 vdd.n12 98.6055
R19436 vdd.n6 vdd.n5 98.6055
R19437 vdd.n4 vdd.n3 98.6055
R19438 vdd.n2 vdd.n1 98.6055
R19439 vdd.t115 vdd.n303 85.8723
R19440 vdd.t122 vdd.n244 85.8723
R19441 vdd.t112 vdd.n201 85.8723
R19442 vdd.t108 vdd.n142 85.8723
R19443 vdd.t269 vdd.n100 85.8723
R19444 vdd.t251 vdd.n41 85.8723
R19445 vdd.t56 vdd.n1722 85.8723
R19446 vdd.t59 vdd.n1781 85.8723
R19447 vdd.t247 vdd.n1620 85.8723
R19448 vdd.t283 vdd.n1679 85.8723
R19449 vdd.t44 vdd.n1519 85.8723
R19450 vdd.t101 vdd.n1578 85.8723
R19451 vdd.n2923 vdd.n2922 78.546
R19452 vdd.n2397 vdd.n1027 78.546
R19453 vdd.n290 vdd.n289 75.1835
R19454 vdd.n288 vdd.n287 75.1835
R19455 vdd.n286 vdd.n285 75.1835
R19456 vdd.n284 vdd.n283 75.1835
R19457 vdd.n282 vdd.n281 75.1835
R19458 vdd.n280 vdd.n279 75.1835
R19459 vdd.n278 vdd.n277 75.1835
R19460 vdd.n276 vdd.n275 75.1835
R19461 vdd.n274 vdd.n273 75.1835
R19462 vdd.n188 vdd.n187 75.1835
R19463 vdd.n186 vdd.n185 75.1835
R19464 vdd.n184 vdd.n183 75.1835
R19465 vdd.n182 vdd.n181 75.1835
R19466 vdd.n180 vdd.n179 75.1835
R19467 vdd.n178 vdd.n177 75.1835
R19468 vdd.n176 vdd.n175 75.1835
R19469 vdd.n174 vdd.n173 75.1835
R19470 vdd.n172 vdd.n171 75.1835
R19471 vdd.n87 vdd.n86 75.1835
R19472 vdd.n85 vdd.n84 75.1835
R19473 vdd.n83 vdd.n82 75.1835
R19474 vdd.n81 vdd.n80 75.1835
R19475 vdd.n79 vdd.n78 75.1835
R19476 vdd.n77 vdd.n76 75.1835
R19477 vdd.n75 vdd.n74 75.1835
R19478 vdd.n73 vdd.n72 75.1835
R19479 vdd.n71 vdd.n70 75.1835
R19480 vdd.n1752 vdd.n1751 75.1835
R19481 vdd.n1754 vdd.n1753 75.1835
R19482 vdd.n1756 vdd.n1755 75.1835
R19483 vdd.n1758 vdd.n1757 75.1835
R19484 vdd.n1760 vdd.n1759 75.1835
R19485 vdd.n1762 vdd.n1761 75.1835
R19486 vdd.n1764 vdd.n1763 75.1835
R19487 vdd.n1766 vdd.n1765 75.1835
R19488 vdd.n1768 vdd.n1767 75.1835
R19489 vdd.n1650 vdd.n1649 75.1835
R19490 vdd.n1652 vdd.n1651 75.1835
R19491 vdd.n1654 vdd.n1653 75.1835
R19492 vdd.n1656 vdd.n1655 75.1835
R19493 vdd.n1658 vdd.n1657 75.1835
R19494 vdd.n1660 vdd.n1659 75.1835
R19495 vdd.n1662 vdd.n1661 75.1835
R19496 vdd.n1664 vdd.n1663 75.1835
R19497 vdd.n1666 vdd.n1665 75.1835
R19498 vdd.n1549 vdd.n1548 75.1835
R19499 vdd.n1551 vdd.n1550 75.1835
R19500 vdd.n1553 vdd.n1552 75.1835
R19501 vdd.n1555 vdd.n1554 75.1835
R19502 vdd.n1557 vdd.n1556 75.1835
R19503 vdd.n1559 vdd.n1558 75.1835
R19504 vdd.n1561 vdd.n1560 75.1835
R19505 vdd.n1563 vdd.n1562 75.1835
R19506 vdd.n1565 vdd.n1564 75.1835
R19507 vdd.n2858 vdd.n2857 72.8958
R19508 vdd.n2857 vdd.n2621 72.8958
R19509 vdd.n2857 vdd.n2622 72.8958
R19510 vdd.n2857 vdd.n2623 72.8958
R19511 vdd.n2857 vdd.n2624 72.8958
R19512 vdd.n2857 vdd.n2625 72.8958
R19513 vdd.n2857 vdd.n2626 72.8958
R19514 vdd.n2857 vdd.n2627 72.8958
R19515 vdd.n2857 vdd.n2628 72.8958
R19516 vdd.n2857 vdd.n2629 72.8958
R19517 vdd.n2857 vdd.n2630 72.8958
R19518 vdd.n2857 vdd.n2631 72.8958
R19519 vdd.n2857 vdd.n2632 72.8958
R19520 vdd.n2857 vdd.n2633 72.8958
R19521 vdd.n2857 vdd.n2634 72.8958
R19522 vdd.n2857 vdd.n2635 72.8958
R19523 vdd.n2857 vdd.n2636 72.8958
R19524 vdd.n803 vdd.n692 72.8958
R19525 vdd.n3066 vdd.n692 72.8958
R19526 vdd.n797 vdd.n692 72.8958
R19527 vdd.n3073 vdd.n692 72.8958
R19528 vdd.n794 vdd.n692 72.8958
R19529 vdd.n3080 vdd.n692 72.8958
R19530 vdd.n791 vdd.n692 72.8958
R19531 vdd.n3087 vdd.n692 72.8958
R19532 vdd.n3090 vdd.n692 72.8958
R19533 vdd.n2946 vdd.n692 72.8958
R19534 vdd.n2951 vdd.n692 72.8958
R19535 vdd.n2945 vdd.n692 72.8958
R19536 vdd.n2958 vdd.n692 72.8958
R19537 vdd.n2942 vdd.n692 72.8958
R19538 vdd.n2965 vdd.n692 72.8958
R19539 vdd.n2939 vdd.n692 72.8958
R19540 vdd.n2972 vdd.n692 72.8958
R19541 vdd.n2110 vdd.n1049 72.8958
R19542 vdd.n2116 vdd.n1049 72.8958
R19543 vdd.n2118 vdd.n1049 72.8958
R19544 vdd.n2124 vdd.n1049 72.8958
R19545 vdd.n2126 vdd.n1049 72.8958
R19546 vdd.n2132 vdd.n1049 72.8958
R19547 vdd.n2134 vdd.n1049 72.8958
R19548 vdd.n2140 vdd.n1049 72.8958
R19549 vdd.n2311 vdd.n1049 72.8958
R19550 vdd.n2309 vdd.n1049 72.8958
R19551 vdd.n2303 vdd.n1049 72.8958
R19552 vdd.n2301 vdd.n1049 72.8958
R19553 vdd.n2295 vdd.n1049 72.8958
R19554 vdd.n2293 vdd.n1049 72.8958
R19555 vdd.n2287 vdd.n1049 72.8958
R19556 vdd.n2285 vdd.n1049 72.8958
R19557 vdd.n2279 vdd.n1049 72.8958
R19558 vdd.n2604 vdd.n937 72.8958
R19559 vdd.n2604 vdd.n938 72.8958
R19560 vdd.n2604 vdd.n939 72.8958
R19561 vdd.n2604 vdd.n940 72.8958
R19562 vdd.n2604 vdd.n941 72.8958
R19563 vdd.n2604 vdd.n942 72.8958
R19564 vdd.n2604 vdd.n943 72.8958
R19565 vdd.n2604 vdd.n944 72.8958
R19566 vdd.n2604 vdd.n945 72.8958
R19567 vdd.n2604 vdd.n946 72.8958
R19568 vdd.n2604 vdd.n947 72.8958
R19569 vdd.n2604 vdd.n948 72.8958
R19570 vdd.n2604 vdd.n949 72.8958
R19571 vdd.n2604 vdd.n950 72.8958
R19572 vdd.n2604 vdd.n951 72.8958
R19573 vdd.n2604 vdd.n952 72.8958
R19574 vdd.n2604 vdd.n953 72.8958
R19575 vdd.n2857 vdd.n2856 72.8958
R19576 vdd.n2857 vdd.n2605 72.8958
R19577 vdd.n2857 vdd.n2606 72.8958
R19578 vdd.n2857 vdd.n2607 72.8958
R19579 vdd.n2857 vdd.n2608 72.8958
R19580 vdd.n2857 vdd.n2609 72.8958
R19581 vdd.n2857 vdd.n2610 72.8958
R19582 vdd.n2857 vdd.n2611 72.8958
R19583 vdd.n2857 vdd.n2612 72.8958
R19584 vdd.n2857 vdd.n2613 72.8958
R19585 vdd.n2857 vdd.n2614 72.8958
R19586 vdd.n2857 vdd.n2615 72.8958
R19587 vdd.n2857 vdd.n2616 72.8958
R19588 vdd.n2857 vdd.n2617 72.8958
R19589 vdd.n2857 vdd.n2618 72.8958
R19590 vdd.n2857 vdd.n2619 72.8958
R19591 vdd.n2857 vdd.n2620 72.8958
R19592 vdd.n2996 vdd.n692 72.8958
R19593 vdd.n835 vdd.n692 72.8958
R19594 vdd.n3004 vdd.n692 72.8958
R19595 vdd.n830 vdd.n692 72.8958
R19596 vdd.n3011 vdd.n692 72.8958
R19597 vdd.n827 vdd.n692 72.8958
R19598 vdd.n3018 vdd.n692 72.8958
R19599 vdd.n824 vdd.n692 72.8958
R19600 vdd.n3025 vdd.n692 72.8958
R19601 vdd.n3029 vdd.n692 72.8958
R19602 vdd.n821 vdd.n692 72.8958
R19603 vdd.n3036 vdd.n692 72.8958
R19604 vdd.n818 vdd.n692 72.8958
R19605 vdd.n3043 vdd.n692 72.8958
R19606 vdd.n815 vdd.n692 72.8958
R19607 vdd.n3050 vdd.n692 72.8958
R19608 vdd.n3053 vdd.n692 72.8958
R19609 vdd.n2604 vdd.n935 72.8958
R19610 vdd.n2604 vdd.n934 72.8958
R19611 vdd.n2604 vdd.n933 72.8958
R19612 vdd.n2604 vdd.n932 72.8958
R19613 vdd.n2604 vdd.n931 72.8958
R19614 vdd.n2604 vdd.n930 72.8958
R19615 vdd.n2604 vdd.n929 72.8958
R19616 vdd.n2604 vdd.n928 72.8958
R19617 vdd.n2604 vdd.n927 72.8958
R19618 vdd.n2604 vdd.n926 72.8958
R19619 vdd.n2604 vdd.n925 72.8958
R19620 vdd.n2604 vdd.n924 72.8958
R19621 vdd.n2604 vdd.n923 72.8958
R19622 vdd.n2604 vdd.n922 72.8958
R19623 vdd.n2604 vdd.n921 72.8958
R19624 vdd.n2604 vdd.n920 72.8958
R19625 vdd.n2604 vdd.n919 72.8958
R19626 vdd.n2369 vdd.n1049 72.8958
R19627 vdd.n2367 vdd.n1049 72.8958
R19628 vdd.n2361 vdd.n1049 72.8958
R19629 vdd.n2359 vdd.n1049 72.8958
R19630 vdd.n2353 vdd.n1049 72.8958
R19631 vdd.n2351 vdd.n1049 72.8958
R19632 vdd.n2345 vdd.n1049 72.8958
R19633 vdd.n2343 vdd.n1049 72.8958
R19634 vdd.n1061 vdd.n1049 72.8958
R19635 vdd.n2185 vdd.n1049 72.8958
R19636 vdd.n2190 vdd.n1049 72.8958
R19637 vdd.n2192 vdd.n1049 72.8958
R19638 vdd.n2198 vdd.n1049 72.8958
R19639 vdd.n2200 vdd.n1049 72.8958
R19640 vdd.n2206 vdd.n1049 72.8958
R19641 vdd.n2208 vdd.n1049 72.8958
R19642 vdd.n2215 vdd.n1049 72.8958
R19643 vdd.n1419 vdd.n1418 66.2847
R19644 vdd.n1418 vdd.n1194 66.2847
R19645 vdd.n1418 vdd.n1195 66.2847
R19646 vdd.n1418 vdd.n1196 66.2847
R19647 vdd.n1418 vdd.n1197 66.2847
R19648 vdd.n1418 vdd.n1198 66.2847
R19649 vdd.n1418 vdd.n1199 66.2847
R19650 vdd.n1418 vdd.n1200 66.2847
R19651 vdd.n1418 vdd.n1201 66.2847
R19652 vdd.n1418 vdd.n1202 66.2847
R19653 vdd.n1418 vdd.n1203 66.2847
R19654 vdd.n1418 vdd.n1204 66.2847
R19655 vdd.n1418 vdd.n1205 66.2847
R19656 vdd.n1418 vdd.n1206 66.2847
R19657 vdd.n1418 vdd.n1207 66.2847
R19658 vdd.n1418 vdd.n1208 66.2847
R19659 vdd.n1418 vdd.n1209 66.2847
R19660 vdd.n1418 vdd.n1210 66.2847
R19661 vdd.n1418 vdd.n1211 66.2847
R19662 vdd.n1418 vdd.n1212 66.2847
R19663 vdd.n1418 vdd.n1213 66.2847
R19664 vdd.n1418 vdd.n1214 66.2847
R19665 vdd.n1418 vdd.n1215 66.2847
R19666 vdd.n1418 vdd.n1216 66.2847
R19667 vdd.n1418 vdd.n1217 66.2847
R19668 vdd.n1418 vdd.n1218 66.2847
R19669 vdd.n1418 vdd.n1219 66.2847
R19670 vdd.n1418 vdd.n1220 66.2847
R19671 vdd.n1418 vdd.n1221 66.2847
R19672 vdd.n1418 vdd.n1222 66.2847
R19673 vdd.n1418 vdd.n1223 66.2847
R19674 vdd.n1073 vdd.n1070 66.2847
R19675 vdd.n2000 vdd.n1073 66.2847
R19676 vdd.n2005 vdd.n1073 66.2847
R19677 vdd.n2010 vdd.n1073 66.2847
R19678 vdd.n1998 vdd.n1073 66.2847
R19679 vdd.n2017 vdd.n1073 66.2847
R19680 vdd.n1990 vdd.n1073 66.2847
R19681 vdd.n2024 vdd.n1073 66.2847
R19682 vdd.n1983 vdd.n1073 66.2847
R19683 vdd.n2031 vdd.n1073 66.2847
R19684 vdd.n1977 vdd.n1073 66.2847
R19685 vdd.n1972 vdd.n1073 66.2847
R19686 vdd.n2042 vdd.n1073 66.2847
R19687 vdd.n1964 vdd.n1073 66.2847
R19688 vdd.n2049 vdd.n1073 66.2847
R19689 vdd.n1957 vdd.n1073 66.2847
R19690 vdd.n2056 vdd.n1073 66.2847
R19691 vdd.n1950 vdd.n1073 66.2847
R19692 vdd.n2063 vdd.n1073 66.2847
R19693 vdd.n1943 vdd.n1073 66.2847
R19694 vdd.n2070 vdd.n1073 66.2847
R19695 vdd.n1937 vdd.n1073 66.2847
R19696 vdd.n1932 vdd.n1073 66.2847
R19697 vdd.n2081 vdd.n1073 66.2847
R19698 vdd.n1924 vdd.n1073 66.2847
R19699 vdd.n2088 vdd.n1073 66.2847
R19700 vdd.n1917 vdd.n1073 66.2847
R19701 vdd.n2095 vdd.n1073 66.2847
R19702 vdd.n2098 vdd.n1073 66.2847
R19703 vdd.n1908 vdd.n1073 66.2847
R19704 vdd.n2320 vdd.n1073 66.2847
R19705 vdd.n1902 vdd.n1073 66.2847
R19706 vdd.n3223 vdd.n3222 66.2847
R19707 vdd.n3223 vdd.n693 66.2847
R19708 vdd.n3223 vdd.n694 66.2847
R19709 vdd.n3223 vdd.n695 66.2847
R19710 vdd.n3223 vdd.n696 66.2847
R19711 vdd.n3223 vdd.n697 66.2847
R19712 vdd.n3223 vdd.n698 66.2847
R19713 vdd.n3223 vdd.n699 66.2847
R19714 vdd.n3223 vdd.n700 66.2847
R19715 vdd.n3223 vdd.n701 66.2847
R19716 vdd.n3223 vdd.n702 66.2847
R19717 vdd.n3223 vdd.n703 66.2847
R19718 vdd.n3223 vdd.n704 66.2847
R19719 vdd.n3223 vdd.n705 66.2847
R19720 vdd.n3223 vdd.n706 66.2847
R19721 vdd.n3223 vdd.n707 66.2847
R19722 vdd.n3223 vdd.n708 66.2847
R19723 vdd.n3223 vdd.n709 66.2847
R19724 vdd.n3223 vdd.n710 66.2847
R19725 vdd.n3223 vdd.n711 66.2847
R19726 vdd.n3223 vdd.n712 66.2847
R19727 vdd.n3223 vdd.n713 66.2847
R19728 vdd.n3223 vdd.n714 66.2847
R19729 vdd.n3223 vdd.n715 66.2847
R19730 vdd.n3223 vdd.n716 66.2847
R19731 vdd.n3223 vdd.n717 66.2847
R19732 vdd.n3223 vdd.n718 66.2847
R19733 vdd.n3223 vdd.n719 66.2847
R19734 vdd.n3223 vdd.n720 66.2847
R19735 vdd.n3223 vdd.n721 66.2847
R19736 vdd.n3223 vdd.n722 66.2847
R19737 vdd.n3354 vdd.n3353 66.2847
R19738 vdd.n3354 vdd.n424 66.2847
R19739 vdd.n3354 vdd.n423 66.2847
R19740 vdd.n3354 vdd.n422 66.2847
R19741 vdd.n3354 vdd.n421 66.2847
R19742 vdd.n3354 vdd.n420 66.2847
R19743 vdd.n3354 vdd.n419 66.2847
R19744 vdd.n3354 vdd.n418 66.2847
R19745 vdd.n3354 vdd.n417 66.2847
R19746 vdd.n3354 vdd.n416 66.2847
R19747 vdd.n3354 vdd.n415 66.2847
R19748 vdd.n3354 vdd.n414 66.2847
R19749 vdd.n3354 vdd.n413 66.2847
R19750 vdd.n3354 vdd.n412 66.2847
R19751 vdd.n3354 vdd.n411 66.2847
R19752 vdd.n3354 vdd.n410 66.2847
R19753 vdd.n3354 vdd.n409 66.2847
R19754 vdd.n3354 vdd.n408 66.2847
R19755 vdd.n3354 vdd.n407 66.2847
R19756 vdd.n3354 vdd.n406 66.2847
R19757 vdd.n3354 vdd.n405 66.2847
R19758 vdd.n3354 vdd.n404 66.2847
R19759 vdd.n3354 vdd.n403 66.2847
R19760 vdd.n3354 vdd.n402 66.2847
R19761 vdd.n3354 vdd.n401 66.2847
R19762 vdd.n3354 vdd.n400 66.2847
R19763 vdd.n3354 vdd.n399 66.2847
R19764 vdd.n3354 vdd.n398 66.2847
R19765 vdd.n3354 vdd.n397 66.2847
R19766 vdd.n3354 vdd.n396 66.2847
R19767 vdd.n3354 vdd.n395 66.2847
R19768 vdd.n3354 vdd.n394 66.2847
R19769 vdd.n467 vdd.n394 52.4337
R19770 vdd.n473 vdd.n395 52.4337
R19771 vdd.n477 vdd.n396 52.4337
R19772 vdd.n483 vdd.n397 52.4337
R19773 vdd.n487 vdd.n398 52.4337
R19774 vdd.n493 vdd.n399 52.4337
R19775 vdd.n497 vdd.n400 52.4337
R19776 vdd.n503 vdd.n401 52.4337
R19777 vdd.n507 vdd.n402 52.4337
R19778 vdd.n513 vdd.n403 52.4337
R19779 vdd.n517 vdd.n404 52.4337
R19780 vdd.n523 vdd.n405 52.4337
R19781 vdd.n527 vdd.n406 52.4337
R19782 vdd.n533 vdd.n407 52.4337
R19783 vdd.n537 vdd.n408 52.4337
R19784 vdd.n543 vdd.n409 52.4337
R19785 vdd.n547 vdd.n410 52.4337
R19786 vdd.n553 vdd.n411 52.4337
R19787 vdd.n557 vdd.n412 52.4337
R19788 vdd.n563 vdd.n413 52.4337
R19789 vdd.n567 vdd.n414 52.4337
R19790 vdd.n573 vdd.n415 52.4337
R19791 vdd.n577 vdd.n416 52.4337
R19792 vdd.n583 vdd.n417 52.4337
R19793 vdd.n587 vdd.n418 52.4337
R19794 vdd.n593 vdd.n419 52.4337
R19795 vdd.n597 vdd.n420 52.4337
R19796 vdd.n603 vdd.n421 52.4337
R19797 vdd.n607 vdd.n422 52.4337
R19798 vdd.n613 vdd.n423 52.4337
R19799 vdd.n616 vdd.n424 52.4337
R19800 vdd.n3353 vdd.n3352 52.4337
R19801 vdd.n3222 vdd.n3221 52.4337
R19802 vdd.n728 vdd.n693 52.4337
R19803 vdd.n734 vdd.n694 52.4337
R19804 vdd.n3211 vdd.n695 52.4337
R19805 vdd.n3207 vdd.n696 52.4337
R19806 vdd.n3203 vdd.n697 52.4337
R19807 vdd.n3199 vdd.n698 52.4337
R19808 vdd.n3195 vdd.n699 52.4337
R19809 vdd.n3191 vdd.n700 52.4337
R19810 vdd.n3187 vdd.n701 52.4337
R19811 vdd.n3179 vdd.n702 52.4337
R19812 vdd.n3175 vdd.n703 52.4337
R19813 vdd.n3171 vdd.n704 52.4337
R19814 vdd.n3167 vdd.n705 52.4337
R19815 vdd.n3163 vdd.n706 52.4337
R19816 vdd.n3159 vdd.n707 52.4337
R19817 vdd.n3155 vdd.n708 52.4337
R19818 vdd.n3151 vdd.n709 52.4337
R19819 vdd.n3147 vdd.n710 52.4337
R19820 vdd.n3143 vdd.n711 52.4337
R19821 vdd.n3139 vdd.n712 52.4337
R19822 vdd.n3133 vdd.n713 52.4337
R19823 vdd.n3129 vdd.n714 52.4337
R19824 vdd.n3125 vdd.n715 52.4337
R19825 vdd.n3121 vdd.n716 52.4337
R19826 vdd.n3117 vdd.n717 52.4337
R19827 vdd.n3113 vdd.n718 52.4337
R19828 vdd.n3109 vdd.n719 52.4337
R19829 vdd.n3105 vdd.n720 52.4337
R19830 vdd.n3101 vdd.n721 52.4337
R19831 vdd.n3097 vdd.n722 52.4337
R19832 vdd.n2322 vdd.n1902 52.4337
R19833 vdd.n2320 vdd.n2319 52.4337
R19834 vdd.n1909 vdd.n1908 52.4337
R19835 vdd.n2098 vdd.n2097 52.4337
R19836 vdd.n2095 vdd.n2094 52.4337
R19837 vdd.n2090 vdd.n1917 52.4337
R19838 vdd.n2088 vdd.n2087 52.4337
R19839 vdd.n2083 vdd.n1924 52.4337
R19840 vdd.n2081 vdd.n2080 52.4337
R19841 vdd.n1933 vdd.n1932 52.4337
R19842 vdd.n2072 vdd.n1937 52.4337
R19843 vdd.n2070 vdd.n2069 52.4337
R19844 vdd.n2065 vdd.n1943 52.4337
R19845 vdd.n2063 vdd.n2062 52.4337
R19846 vdd.n2058 vdd.n1950 52.4337
R19847 vdd.n2056 vdd.n2055 52.4337
R19848 vdd.n2051 vdd.n1957 52.4337
R19849 vdd.n2049 vdd.n2048 52.4337
R19850 vdd.n2044 vdd.n1964 52.4337
R19851 vdd.n2042 vdd.n2041 52.4337
R19852 vdd.n1973 vdd.n1972 52.4337
R19853 vdd.n2033 vdd.n1977 52.4337
R19854 vdd.n2031 vdd.n2030 52.4337
R19855 vdd.n2026 vdd.n1983 52.4337
R19856 vdd.n2024 vdd.n2023 52.4337
R19857 vdd.n2019 vdd.n1990 52.4337
R19858 vdd.n2017 vdd.n2016 52.4337
R19859 vdd.n2012 vdd.n1998 52.4337
R19860 vdd.n2010 vdd.n2009 52.4337
R19861 vdd.n2005 vdd.n2004 52.4337
R19862 vdd.n2000 vdd.n1999 52.4337
R19863 vdd.n2331 vdd.n1070 52.4337
R19864 vdd.n1420 vdd.n1419 52.4337
R19865 vdd.n1226 vdd.n1194 52.4337
R19866 vdd.n1230 vdd.n1195 52.4337
R19867 vdd.n1232 vdd.n1196 52.4337
R19868 vdd.n1236 vdd.n1197 52.4337
R19869 vdd.n1238 vdd.n1198 52.4337
R19870 vdd.n1242 vdd.n1199 52.4337
R19871 vdd.n1244 vdd.n1200 52.4337
R19872 vdd.n1248 vdd.n1201 52.4337
R19873 vdd.n1250 vdd.n1202 52.4337
R19874 vdd.n1256 vdd.n1203 52.4337
R19875 vdd.n1258 vdd.n1204 52.4337
R19876 vdd.n1262 vdd.n1205 52.4337
R19877 vdd.n1264 vdd.n1206 52.4337
R19878 vdd.n1268 vdd.n1207 52.4337
R19879 vdd.n1270 vdd.n1208 52.4337
R19880 vdd.n1274 vdd.n1209 52.4337
R19881 vdd.n1276 vdd.n1210 52.4337
R19882 vdd.n1280 vdd.n1211 52.4337
R19883 vdd.n1282 vdd.n1212 52.4337
R19884 vdd.n1354 vdd.n1213 52.4337
R19885 vdd.n1287 vdd.n1214 52.4337
R19886 vdd.n1291 vdd.n1215 52.4337
R19887 vdd.n1293 vdd.n1216 52.4337
R19888 vdd.n1297 vdd.n1217 52.4337
R19889 vdd.n1299 vdd.n1218 52.4337
R19890 vdd.n1303 vdd.n1219 52.4337
R19891 vdd.n1305 vdd.n1220 52.4337
R19892 vdd.n1309 vdd.n1221 52.4337
R19893 vdd.n1311 vdd.n1222 52.4337
R19894 vdd.n1315 vdd.n1223 52.4337
R19895 vdd.n1419 vdd.n1193 52.4337
R19896 vdd.n1229 vdd.n1194 52.4337
R19897 vdd.n1231 vdd.n1195 52.4337
R19898 vdd.n1235 vdd.n1196 52.4337
R19899 vdd.n1237 vdd.n1197 52.4337
R19900 vdd.n1241 vdd.n1198 52.4337
R19901 vdd.n1243 vdd.n1199 52.4337
R19902 vdd.n1247 vdd.n1200 52.4337
R19903 vdd.n1249 vdd.n1201 52.4337
R19904 vdd.n1255 vdd.n1202 52.4337
R19905 vdd.n1257 vdd.n1203 52.4337
R19906 vdd.n1261 vdd.n1204 52.4337
R19907 vdd.n1263 vdd.n1205 52.4337
R19908 vdd.n1267 vdd.n1206 52.4337
R19909 vdd.n1269 vdd.n1207 52.4337
R19910 vdd.n1273 vdd.n1208 52.4337
R19911 vdd.n1275 vdd.n1209 52.4337
R19912 vdd.n1279 vdd.n1210 52.4337
R19913 vdd.n1281 vdd.n1211 52.4337
R19914 vdd.n1285 vdd.n1212 52.4337
R19915 vdd.n1286 vdd.n1213 52.4337
R19916 vdd.n1290 vdd.n1214 52.4337
R19917 vdd.n1292 vdd.n1215 52.4337
R19918 vdd.n1296 vdd.n1216 52.4337
R19919 vdd.n1298 vdd.n1217 52.4337
R19920 vdd.n1302 vdd.n1218 52.4337
R19921 vdd.n1304 vdd.n1219 52.4337
R19922 vdd.n1308 vdd.n1220 52.4337
R19923 vdd.n1310 vdd.n1221 52.4337
R19924 vdd.n1314 vdd.n1222 52.4337
R19925 vdd.n1316 vdd.n1223 52.4337
R19926 vdd.n1070 vdd.n1069 52.4337
R19927 vdd.n2001 vdd.n2000 52.4337
R19928 vdd.n2006 vdd.n2005 52.4337
R19929 vdd.n2011 vdd.n2010 52.4337
R19930 vdd.n1998 vdd.n1991 52.4337
R19931 vdd.n2018 vdd.n2017 52.4337
R19932 vdd.n1990 vdd.n1984 52.4337
R19933 vdd.n2025 vdd.n2024 52.4337
R19934 vdd.n1983 vdd.n1978 52.4337
R19935 vdd.n2032 vdd.n2031 52.4337
R19936 vdd.n1977 vdd.n1976 52.4337
R19937 vdd.n1972 vdd.n1965 52.4337
R19938 vdd.n2043 vdd.n2042 52.4337
R19939 vdd.n1964 vdd.n1958 52.4337
R19940 vdd.n2050 vdd.n2049 52.4337
R19941 vdd.n1957 vdd.n1951 52.4337
R19942 vdd.n2057 vdd.n2056 52.4337
R19943 vdd.n1950 vdd.n1944 52.4337
R19944 vdd.n2064 vdd.n2063 52.4337
R19945 vdd.n1943 vdd.n1938 52.4337
R19946 vdd.n2071 vdd.n2070 52.4337
R19947 vdd.n1937 vdd.n1936 52.4337
R19948 vdd.n1932 vdd.n1925 52.4337
R19949 vdd.n2082 vdd.n2081 52.4337
R19950 vdd.n1924 vdd.n1918 52.4337
R19951 vdd.n2089 vdd.n2088 52.4337
R19952 vdd.n1917 vdd.n1911 52.4337
R19953 vdd.n2096 vdd.n2095 52.4337
R19954 vdd.n2099 vdd.n2098 52.4337
R19955 vdd.n1908 vdd.n1903 52.4337
R19956 vdd.n2321 vdd.n2320 52.4337
R19957 vdd.n1902 vdd.n1075 52.4337
R19958 vdd.n3222 vdd.n725 52.4337
R19959 vdd.n733 vdd.n693 52.4337
R19960 vdd.n3212 vdd.n694 52.4337
R19961 vdd.n3208 vdd.n695 52.4337
R19962 vdd.n3204 vdd.n696 52.4337
R19963 vdd.n3200 vdd.n697 52.4337
R19964 vdd.n3196 vdd.n698 52.4337
R19965 vdd.n3192 vdd.n699 52.4337
R19966 vdd.n3188 vdd.n700 52.4337
R19967 vdd.n3178 vdd.n701 52.4337
R19968 vdd.n3176 vdd.n702 52.4337
R19969 vdd.n3172 vdd.n703 52.4337
R19970 vdd.n3168 vdd.n704 52.4337
R19971 vdd.n3164 vdd.n705 52.4337
R19972 vdd.n3160 vdd.n706 52.4337
R19973 vdd.n3156 vdd.n707 52.4337
R19974 vdd.n3152 vdd.n708 52.4337
R19975 vdd.n3148 vdd.n709 52.4337
R19976 vdd.n3144 vdd.n710 52.4337
R19977 vdd.n3140 vdd.n711 52.4337
R19978 vdd.n3132 vdd.n712 52.4337
R19979 vdd.n3130 vdd.n713 52.4337
R19980 vdd.n3126 vdd.n714 52.4337
R19981 vdd.n3122 vdd.n715 52.4337
R19982 vdd.n3118 vdd.n716 52.4337
R19983 vdd.n3114 vdd.n717 52.4337
R19984 vdd.n3110 vdd.n718 52.4337
R19985 vdd.n3106 vdd.n719 52.4337
R19986 vdd.n3102 vdd.n720 52.4337
R19987 vdd.n3098 vdd.n721 52.4337
R19988 vdd.n722 vdd.n691 52.4337
R19989 vdd.n3353 vdd.n425 52.4337
R19990 vdd.n614 vdd.n424 52.4337
R19991 vdd.n608 vdd.n423 52.4337
R19992 vdd.n604 vdd.n422 52.4337
R19993 vdd.n598 vdd.n421 52.4337
R19994 vdd.n594 vdd.n420 52.4337
R19995 vdd.n588 vdd.n419 52.4337
R19996 vdd.n584 vdd.n418 52.4337
R19997 vdd.n578 vdd.n417 52.4337
R19998 vdd.n574 vdd.n416 52.4337
R19999 vdd.n568 vdd.n415 52.4337
R20000 vdd.n564 vdd.n414 52.4337
R20001 vdd.n558 vdd.n413 52.4337
R20002 vdd.n554 vdd.n412 52.4337
R20003 vdd.n548 vdd.n411 52.4337
R20004 vdd.n544 vdd.n410 52.4337
R20005 vdd.n538 vdd.n409 52.4337
R20006 vdd.n534 vdd.n408 52.4337
R20007 vdd.n528 vdd.n407 52.4337
R20008 vdd.n524 vdd.n406 52.4337
R20009 vdd.n518 vdd.n405 52.4337
R20010 vdd.n514 vdd.n404 52.4337
R20011 vdd.n508 vdd.n403 52.4337
R20012 vdd.n504 vdd.n402 52.4337
R20013 vdd.n498 vdd.n401 52.4337
R20014 vdd.n494 vdd.n400 52.4337
R20015 vdd.n488 vdd.n399 52.4337
R20016 vdd.n484 vdd.n398 52.4337
R20017 vdd.n478 vdd.n397 52.4337
R20018 vdd.n474 vdd.n396 52.4337
R20019 vdd.n468 vdd.n395 52.4337
R20020 vdd.n394 vdd.n392 52.4337
R20021 vdd.t129 vdd.t142 51.4683
R20022 vdd.n274 vdd.n272 42.0461
R20023 vdd.n172 vdd.n170 42.0461
R20024 vdd.n71 vdd.n69 42.0461
R20025 vdd.n1752 vdd.n1750 42.0461
R20026 vdd.n1650 vdd.n1648 42.0461
R20027 vdd.n1549 vdd.n1547 42.0461
R20028 vdd.n332 vdd.n331 41.6884
R20029 vdd.n230 vdd.n229 41.6884
R20030 vdd.n129 vdd.n128 41.6884
R20031 vdd.n1810 vdd.n1809 41.6884
R20032 vdd.n1708 vdd.n1707 41.6884
R20033 vdd.n1607 vdd.n1606 41.6884
R20034 vdd.n1319 vdd.n1318 41.1157
R20035 vdd.n1357 vdd.n1356 41.1157
R20036 vdd.n1253 vdd.n1252 41.1157
R20037 vdd.n428 vdd.n427 41.1157
R20038 vdd.n566 vdd.n441 41.1157
R20039 vdd.n454 vdd.n453 41.1157
R20040 vdd.n3053 vdd.n3052 39.2114
R20041 vdd.n3050 vdd.n3049 39.2114
R20042 vdd.n3045 vdd.n815 39.2114
R20043 vdd.n3043 vdd.n3042 39.2114
R20044 vdd.n3038 vdd.n818 39.2114
R20045 vdd.n3036 vdd.n3035 39.2114
R20046 vdd.n3031 vdd.n821 39.2114
R20047 vdd.n3029 vdd.n3028 39.2114
R20048 vdd.n3025 vdd.n3024 39.2114
R20049 vdd.n3020 vdd.n824 39.2114
R20050 vdd.n3018 vdd.n3017 39.2114
R20051 vdd.n3013 vdd.n827 39.2114
R20052 vdd.n3011 vdd.n3010 39.2114
R20053 vdd.n3006 vdd.n830 39.2114
R20054 vdd.n3004 vdd.n3003 39.2114
R20055 vdd.n2998 vdd.n835 39.2114
R20056 vdd.n2996 vdd.n2995 39.2114
R20057 vdd.n2856 vdd.n913 39.2114
R20058 vdd.n2851 vdd.n2605 39.2114
R20059 vdd.n2848 vdd.n2606 39.2114
R20060 vdd.n2844 vdd.n2607 39.2114
R20061 vdd.n2840 vdd.n2608 39.2114
R20062 vdd.n2836 vdd.n2609 39.2114
R20063 vdd.n2832 vdd.n2610 39.2114
R20064 vdd.n2828 vdd.n2611 39.2114
R20065 vdd.n2824 vdd.n2612 39.2114
R20066 vdd.n2820 vdd.n2613 39.2114
R20067 vdd.n2816 vdd.n2614 39.2114
R20068 vdd.n2812 vdd.n2615 39.2114
R20069 vdd.n2808 vdd.n2616 39.2114
R20070 vdd.n2804 vdd.n2617 39.2114
R20071 vdd.n2800 vdd.n2618 39.2114
R20072 vdd.n2796 vdd.n2619 39.2114
R20073 vdd.n2791 vdd.n2620 39.2114
R20074 vdd.n2599 vdd.n953 39.2114
R20075 vdd.n2595 vdd.n952 39.2114
R20076 vdd.n2591 vdd.n951 39.2114
R20077 vdd.n2587 vdd.n950 39.2114
R20078 vdd.n2583 vdd.n949 39.2114
R20079 vdd.n2579 vdd.n948 39.2114
R20080 vdd.n2575 vdd.n947 39.2114
R20081 vdd.n2571 vdd.n946 39.2114
R20082 vdd.n2567 vdd.n945 39.2114
R20083 vdd.n2563 vdd.n944 39.2114
R20084 vdd.n2559 vdd.n943 39.2114
R20085 vdd.n2555 vdd.n942 39.2114
R20086 vdd.n2551 vdd.n941 39.2114
R20087 vdd.n2547 vdd.n940 39.2114
R20088 vdd.n2543 vdd.n939 39.2114
R20089 vdd.n2538 vdd.n938 39.2114
R20090 vdd.n2534 vdd.n937 39.2114
R20091 vdd.n2110 vdd.n1048 39.2114
R20092 vdd.n2116 vdd.n2115 39.2114
R20093 vdd.n2119 vdd.n2118 39.2114
R20094 vdd.n2124 vdd.n2123 39.2114
R20095 vdd.n2127 vdd.n2126 39.2114
R20096 vdd.n2132 vdd.n2131 39.2114
R20097 vdd.n2135 vdd.n2134 39.2114
R20098 vdd.n2140 vdd.n2139 39.2114
R20099 vdd.n2311 vdd.n2142 39.2114
R20100 vdd.n2310 vdd.n2309 39.2114
R20101 vdd.n2303 vdd.n2144 39.2114
R20102 vdd.n2302 vdd.n2301 39.2114
R20103 vdd.n2295 vdd.n2146 39.2114
R20104 vdd.n2294 vdd.n2293 39.2114
R20105 vdd.n2287 vdd.n2148 39.2114
R20106 vdd.n2286 vdd.n2285 39.2114
R20107 vdd.n2279 vdd.n2150 39.2114
R20108 vdd.n2972 vdd.n2971 39.2114
R20109 vdd.n2967 vdd.n2939 39.2114
R20110 vdd.n2965 vdd.n2964 39.2114
R20111 vdd.n2960 vdd.n2942 39.2114
R20112 vdd.n2958 vdd.n2957 39.2114
R20113 vdd.n2953 vdd.n2945 39.2114
R20114 vdd.n2951 vdd.n2950 39.2114
R20115 vdd.n2946 vdd.n787 39.2114
R20116 vdd.n3090 vdd.n3089 39.2114
R20117 vdd.n3087 vdd.n3086 39.2114
R20118 vdd.n3082 vdd.n791 39.2114
R20119 vdd.n3080 vdd.n3079 39.2114
R20120 vdd.n3075 vdd.n794 39.2114
R20121 vdd.n3073 vdd.n3072 39.2114
R20122 vdd.n3068 vdd.n797 39.2114
R20123 vdd.n3066 vdd.n3065 39.2114
R20124 vdd.n3061 vdd.n803 39.2114
R20125 vdd.n2858 vdd.n916 39.2114
R20126 vdd.n2621 vdd.n918 39.2114
R20127 vdd.n2647 vdd.n2622 39.2114
R20128 vdd.n2651 vdd.n2623 39.2114
R20129 vdd.n2655 vdd.n2624 39.2114
R20130 vdd.n2659 vdd.n2625 39.2114
R20131 vdd.n2663 vdd.n2626 39.2114
R20132 vdd.n2667 vdd.n2627 39.2114
R20133 vdd.n2671 vdd.n2628 39.2114
R20134 vdd.n2675 vdd.n2629 39.2114
R20135 vdd.n2679 vdd.n2630 39.2114
R20136 vdd.n2683 vdd.n2631 39.2114
R20137 vdd.n2687 vdd.n2632 39.2114
R20138 vdd.n2691 vdd.n2633 39.2114
R20139 vdd.n2695 vdd.n2634 39.2114
R20140 vdd.n2699 vdd.n2635 39.2114
R20141 vdd.n2703 vdd.n2636 39.2114
R20142 vdd.n2859 vdd.n2858 39.2114
R20143 vdd.n2646 vdd.n2621 39.2114
R20144 vdd.n2650 vdd.n2622 39.2114
R20145 vdd.n2654 vdd.n2623 39.2114
R20146 vdd.n2658 vdd.n2624 39.2114
R20147 vdd.n2662 vdd.n2625 39.2114
R20148 vdd.n2666 vdd.n2626 39.2114
R20149 vdd.n2670 vdd.n2627 39.2114
R20150 vdd.n2674 vdd.n2628 39.2114
R20151 vdd.n2678 vdd.n2629 39.2114
R20152 vdd.n2682 vdd.n2630 39.2114
R20153 vdd.n2686 vdd.n2631 39.2114
R20154 vdd.n2690 vdd.n2632 39.2114
R20155 vdd.n2694 vdd.n2633 39.2114
R20156 vdd.n2698 vdd.n2634 39.2114
R20157 vdd.n2702 vdd.n2635 39.2114
R20158 vdd.n2705 vdd.n2636 39.2114
R20159 vdd.n803 vdd.n798 39.2114
R20160 vdd.n3067 vdd.n3066 39.2114
R20161 vdd.n797 vdd.n795 39.2114
R20162 vdd.n3074 vdd.n3073 39.2114
R20163 vdd.n794 vdd.n792 39.2114
R20164 vdd.n3081 vdd.n3080 39.2114
R20165 vdd.n791 vdd.n789 39.2114
R20166 vdd.n3088 vdd.n3087 39.2114
R20167 vdd.n3091 vdd.n3090 39.2114
R20168 vdd.n2947 vdd.n2946 39.2114
R20169 vdd.n2952 vdd.n2951 39.2114
R20170 vdd.n2945 vdd.n2943 39.2114
R20171 vdd.n2959 vdd.n2958 39.2114
R20172 vdd.n2942 vdd.n2940 39.2114
R20173 vdd.n2966 vdd.n2965 39.2114
R20174 vdd.n2939 vdd.n2937 39.2114
R20175 vdd.n2973 vdd.n2972 39.2114
R20176 vdd.n2111 vdd.n2110 39.2114
R20177 vdd.n2117 vdd.n2116 39.2114
R20178 vdd.n2118 vdd.n2107 39.2114
R20179 vdd.n2125 vdd.n2124 39.2114
R20180 vdd.n2126 vdd.n2105 39.2114
R20181 vdd.n2133 vdd.n2132 39.2114
R20182 vdd.n2134 vdd.n2103 39.2114
R20183 vdd.n2141 vdd.n2140 39.2114
R20184 vdd.n2312 vdd.n2311 39.2114
R20185 vdd.n2309 vdd.n2308 39.2114
R20186 vdd.n2304 vdd.n2303 39.2114
R20187 vdd.n2301 vdd.n2300 39.2114
R20188 vdd.n2296 vdd.n2295 39.2114
R20189 vdd.n2293 vdd.n2292 39.2114
R20190 vdd.n2288 vdd.n2287 39.2114
R20191 vdd.n2285 vdd.n2284 39.2114
R20192 vdd.n2280 vdd.n2279 39.2114
R20193 vdd.n2537 vdd.n937 39.2114
R20194 vdd.n2542 vdd.n938 39.2114
R20195 vdd.n2546 vdd.n939 39.2114
R20196 vdd.n2550 vdd.n940 39.2114
R20197 vdd.n2554 vdd.n941 39.2114
R20198 vdd.n2558 vdd.n942 39.2114
R20199 vdd.n2562 vdd.n943 39.2114
R20200 vdd.n2566 vdd.n944 39.2114
R20201 vdd.n2570 vdd.n945 39.2114
R20202 vdd.n2574 vdd.n946 39.2114
R20203 vdd.n2578 vdd.n947 39.2114
R20204 vdd.n2582 vdd.n948 39.2114
R20205 vdd.n2586 vdd.n949 39.2114
R20206 vdd.n2590 vdd.n950 39.2114
R20207 vdd.n2594 vdd.n951 39.2114
R20208 vdd.n2598 vdd.n952 39.2114
R20209 vdd.n955 vdd.n953 39.2114
R20210 vdd.n2856 vdd.n2855 39.2114
R20211 vdd.n2849 vdd.n2605 39.2114
R20212 vdd.n2845 vdd.n2606 39.2114
R20213 vdd.n2841 vdd.n2607 39.2114
R20214 vdd.n2837 vdd.n2608 39.2114
R20215 vdd.n2833 vdd.n2609 39.2114
R20216 vdd.n2829 vdd.n2610 39.2114
R20217 vdd.n2825 vdd.n2611 39.2114
R20218 vdd.n2821 vdd.n2612 39.2114
R20219 vdd.n2817 vdd.n2613 39.2114
R20220 vdd.n2813 vdd.n2614 39.2114
R20221 vdd.n2809 vdd.n2615 39.2114
R20222 vdd.n2805 vdd.n2616 39.2114
R20223 vdd.n2801 vdd.n2617 39.2114
R20224 vdd.n2797 vdd.n2618 39.2114
R20225 vdd.n2792 vdd.n2619 39.2114
R20226 vdd.n2788 vdd.n2620 39.2114
R20227 vdd.n2997 vdd.n2996 39.2114
R20228 vdd.n835 vdd.n831 39.2114
R20229 vdd.n3005 vdd.n3004 39.2114
R20230 vdd.n830 vdd.n828 39.2114
R20231 vdd.n3012 vdd.n3011 39.2114
R20232 vdd.n827 vdd.n825 39.2114
R20233 vdd.n3019 vdd.n3018 39.2114
R20234 vdd.n824 vdd.n822 39.2114
R20235 vdd.n3026 vdd.n3025 39.2114
R20236 vdd.n3030 vdd.n3029 39.2114
R20237 vdd.n821 vdd.n819 39.2114
R20238 vdd.n3037 vdd.n3036 39.2114
R20239 vdd.n818 vdd.n816 39.2114
R20240 vdd.n3044 vdd.n3043 39.2114
R20241 vdd.n815 vdd.n813 39.2114
R20242 vdd.n3051 vdd.n3050 39.2114
R20243 vdd.n3054 vdd.n3053 39.2114
R20244 vdd.n963 vdd.n919 39.2114
R20245 vdd.n2526 vdd.n920 39.2114
R20246 vdd.n2522 vdd.n921 39.2114
R20247 vdd.n2518 vdd.n922 39.2114
R20248 vdd.n2514 vdd.n923 39.2114
R20249 vdd.n2510 vdd.n924 39.2114
R20250 vdd.n2506 vdd.n925 39.2114
R20251 vdd.n2502 vdd.n926 39.2114
R20252 vdd.n2498 vdd.n927 39.2114
R20253 vdd.n2494 vdd.n928 39.2114
R20254 vdd.n2490 vdd.n929 39.2114
R20255 vdd.n2486 vdd.n930 39.2114
R20256 vdd.n2482 vdd.n931 39.2114
R20257 vdd.n2478 vdd.n932 39.2114
R20258 vdd.n2474 vdd.n933 39.2114
R20259 vdd.n2470 vdd.n934 39.2114
R20260 vdd.n2466 vdd.n935 39.2114
R20261 vdd.n2369 vdd.n1052 39.2114
R20262 vdd.n2368 vdd.n2367 39.2114
R20263 vdd.n2361 vdd.n1054 39.2114
R20264 vdd.n2360 vdd.n2359 39.2114
R20265 vdd.n2353 vdd.n1056 39.2114
R20266 vdd.n2352 vdd.n2351 39.2114
R20267 vdd.n2345 vdd.n1058 39.2114
R20268 vdd.n2344 vdd.n2343 39.2114
R20269 vdd.n1061 vdd.n1060 39.2114
R20270 vdd.n2185 vdd.n2184 39.2114
R20271 vdd.n2190 vdd.n2189 39.2114
R20272 vdd.n2193 vdd.n2192 39.2114
R20273 vdd.n2198 vdd.n2197 39.2114
R20274 vdd.n2201 vdd.n2200 39.2114
R20275 vdd.n2206 vdd.n2205 39.2114
R20276 vdd.n2209 vdd.n2208 39.2114
R20277 vdd.n2215 vdd.n2214 39.2114
R20278 vdd.n2463 vdd.n935 39.2114
R20279 vdd.n2467 vdd.n934 39.2114
R20280 vdd.n2471 vdd.n933 39.2114
R20281 vdd.n2475 vdd.n932 39.2114
R20282 vdd.n2479 vdd.n931 39.2114
R20283 vdd.n2483 vdd.n930 39.2114
R20284 vdd.n2487 vdd.n929 39.2114
R20285 vdd.n2491 vdd.n928 39.2114
R20286 vdd.n2495 vdd.n927 39.2114
R20287 vdd.n2499 vdd.n926 39.2114
R20288 vdd.n2503 vdd.n925 39.2114
R20289 vdd.n2507 vdd.n924 39.2114
R20290 vdd.n2511 vdd.n923 39.2114
R20291 vdd.n2515 vdd.n922 39.2114
R20292 vdd.n2519 vdd.n921 39.2114
R20293 vdd.n2523 vdd.n920 39.2114
R20294 vdd.n2527 vdd.n919 39.2114
R20295 vdd.n2370 vdd.n2369 39.2114
R20296 vdd.n2367 vdd.n2366 39.2114
R20297 vdd.n2362 vdd.n2361 39.2114
R20298 vdd.n2359 vdd.n2358 39.2114
R20299 vdd.n2354 vdd.n2353 39.2114
R20300 vdd.n2351 vdd.n2350 39.2114
R20301 vdd.n2346 vdd.n2345 39.2114
R20302 vdd.n2343 vdd.n2342 39.2114
R20303 vdd.n1062 vdd.n1061 39.2114
R20304 vdd.n2186 vdd.n2185 39.2114
R20305 vdd.n2191 vdd.n2190 39.2114
R20306 vdd.n2192 vdd.n2182 39.2114
R20307 vdd.n2199 vdd.n2198 39.2114
R20308 vdd.n2200 vdd.n2180 39.2114
R20309 vdd.n2207 vdd.n2206 39.2114
R20310 vdd.n2208 vdd.n2176 39.2114
R20311 vdd.n2216 vdd.n2215 39.2114
R20312 vdd.n2335 vdd.n2334 37.2369
R20313 vdd.n2038 vdd.n1971 37.2369
R20314 vdd.n2077 vdd.n1931 37.2369
R20315 vdd.n3138 vdd.n769 37.2369
R20316 vdd.n3186 vdd.n3185 37.2369
R20317 vdd.n690 vdd.n689 37.2369
R20318 vdd.n2377 vdd.n1047 31.6883
R20319 vdd.n2602 vdd.n956 31.6883
R20320 vdd.n2535 vdd.n959 31.6883
R20321 vdd.n2281 vdd.n2278 31.6883
R20322 vdd.n2789 vdd.n2787 31.6883
R20323 vdd.n2994 vdd.n2993 31.6883
R20324 vdd.n2866 vdd.n912 31.6883
R20325 vdd.n3057 vdd.n3056 31.6883
R20326 vdd.n2976 vdd.n2975 31.6883
R20327 vdd.n3062 vdd.n802 31.6883
R20328 vdd.n2708 vdd.n2707 31.6883
R20329 vdd.n2862 vdd.n2861 31.6883
R20330 vdd.n2373 vdd.n2372 31.6883
R20331 vdd.n2530 vdd.n2529 31.6883
R20332 vdd.n2462 vdd.n2461 31.6883
R20333 vdd.n2219 vdd.n2218 31.6883
R20334 vdd.n2212 vdd.n2178 30.449
R20335 vdd.n967 vdd.n966 30.449
R20336 vdd.n2153 vdd.n2152 30.449
R20337 vdd.n2540 vdd.n958 30.449
R20338 vdd.n2644 vdd.n2643 30.449
R20339 vdd.n3000 vdd.n833 30.449
R20340 vdd.n2794 vdd.n2640 30.449
R20341 vdd.n801 vdd.n800 30.449
R20342 vdd.n1418 vdd.n1225 22.2201
R20343 vdd.n2329 vdd.n1073 22.2201
R20344 vdd.n3223 vdd.n723 22.2201
R20345 vdd.n3355 vdd.n3354 22.2201
R20346 vdd.n1429 vdd.n1187 19.3944
R20347 vdd.n1429 vdd.n1185 19.3944
R20348 vdd.n1433 vdd.n1185 19.3944
R20349 vdd.n1433 vdd.n1175 19.3944
R20350 vdd.n1446 vdd.n1175 19.3944
R20351 vdd.n1446 vdd.n1173 19.3944
R20352 vdd.n1450 vdd.n1173 19.3944
R20353 vdd.n1450 vdd.n1165 19.3944
R20354 vdd.n1463 vdd.n1165 19.3944
R20355 vdd.n1463 vdd.n1163 19.3944
R20356 vdd.n1467 vdd.n1163 19.3944
R20357 vdd.n1467 vdd.n1152 19.3944
R20358 vdd.n1479 vdd.n1152 19.3944
R20359 vdd.n1479 vdd.n1150 19.3944
R20360 vdd.n1483 vdd.n1150 19.3944
R20361 vdd.n1483 vdd.n1141 19.3944
R20362 vdd.n1496 vdd.n1141 19.3944
R20363 vdd.n1496 vdd.n1139 19.3944
R20364 vdd.n1500 vdd.n1139 19.3944
R20365 vdd.n1500 vdd.n1130 19.3944
R20366 vdd.n1819 vdd.n1130 19.3944
R20367 vdd.n1819 vdd.n1128 19.3944
R20368 vdd.n1823 vdd.n1128 19.3944
R20369 vdd.n1823 vdd.n1118 19.3944
R20370 vdd.n1836 vdd.n1118 19.3944
R20371 vdd.n1836 vdd.n1116 19.3944
R20372 vdd.n1840 vdd.n1116 19.3944
R20373 vdd.n1840 vdd.n1108 19.3944
R20374 vdd.n1853 vdd.n1108 19.3944
R20375 vdd.n1853 vdd.n1106 19.3944
R20376 vdd.n1857 vdd.n1106 19.3944
R20377 vdd.n1857 vdd.n1095 19.3944
R20378 vdd.n1869 vdd.n1095 19.3944
R20379 vdd.n1869 vdd.n1093 19.3944
R20380 vdd.n1873 vdd.n1093 19.3944
R20381 vdd.n1873 vdd.n1085 19.3944
R20382 vdd.n1886 vdd.n1085 19.3944
R20383 vdd.n1886 vdd.n1082 19.3944
R20384 vdd.n1892 vdd.n1082 19.3944
R20385 vdd.n1892 vdd.n1083 19.3944
R20386 vdd.n1083 vdd.n1072 19.3944
R20387 vdd.n1353 vdd.n1288 19.3944
R20388 vdd.n1349 vdd.n1288 19.3944
R20389 vdd.n1349 vdd.n1348 19.3944
R20390 vdd.n1348 vdd.n1347 19.3944
R20391 vdd.n1347 vdd.n1294 19.3944
R20392 vdd.n1343 vdd.n1294 19.3944
R20393 vdd.n1343 vdd.n1342 19.3944
R20394 vdd.n1342 vdd.n1341 19.3944
R20395 vdd.n1341 vdd.n1300 19.3944
R20396 vdd.n1337 vdd.n1300 19.3944
R20397 vdd.n1337 vdd.n1336 19.3944
R20398 vdd.n1336 vdd.n1335 19.3944
R20399 vdd.n1335 vdd.n1306 19.3944
R20400 vdd.n1331 vdd.n1306 19.3944
R20401 vdd.n1331 vdd.n1330 19.3944
R20402 vdd.n1330 vdd.n1329 19.3944
R20403 vdd.n1329 vdd.n1312 19.3944
R20404 vdd.n1325 vdd.n1312 19.3944
R20405 vdd.n1325 vdd.n1324 19.3944
R20406 vdd.n1324 vdd.n1323 19.3944
R20407 vdd.n1388 vdd.n1387 19.3944
R20408 vdd.n1387 vdd.n1386 19.3944
R20409 vdd.n1386 vdd.n1259 19.3944
R20410 vdd.n1382 vdd.n1259 19.3944
R20411 vdd.n1382 vdd.n1381 19.3944
R20412 vdd.n1381 vdd.n1380 19.3944
R20413 vdd.n1380 vdd.n1265 19.3944
R20414 vdd.n1376 vdd.n1265 19.3944
R20415 vdd.n1376 vdd.n1375 19.3944
R20416 vdd.n1375 vdd.n1374 19.3944
R20417 vdd.n1374 vdd.n1271 19.3944
R20418 vdd.n1370 vdd.n1271 19.3944
R20419 vdd.n1370 vdd.n1369 19.3944
R20420 vdd.n1369 vdd.n1368 19.3944
R20421 vdd.n1368 vdd.n1277 19.3944
R20422 vdd.n1364 vdd.n1277 19.3944
R20423 vdd.n1364 vdd.n1363 19.3944
R20424 vdd.n1363 vdd.n1362 19.3944
R20425 vdd.n1362 vdd.n1283 19.3944
R20426 vdd.n1358 vdd.n1283 19.3944
R20427 vdd.n1421 vdd.n1192 19.3944
R20428 vdd.n1416 vdd.n1192 19.3944
R20429 vdd.n1416 vdd.n1227 19.3944
R20430 vdd.n1412 vdd.n1227 19.3944
R20431 vdd.n1412 vdd.n1411 19.3944
R20432 vdd.n1411 vdd.n1410 19.3944
R20433 vdd.n1410 vdd.n1233 19.3944
R20434 vdd.n1406 vdd.n1233 19.3944
R20435 vdd.n1406 vdd.n1405 19.3944
R20436 vdd.n1405 vdd.n1404 19.3944
R20437 vdd.n1404 vdd.n1239 19.3944
R20438 vdd.n1400 vdd.n1239 19.3944
R20439 vdd.n1400 vdd.n1399 19.3944
R20440 vdd.n1399 vdd.n1398 19.3944
R20441 vdd.n1398 vdd.n1245 19.3944
R20442 vdd.n1394 vdd.n1245 19.3944
R20443 vdd.n1394 vdd.n1393 19.3944
R20444 vdd.n1393 vdd.n1392 19.3944
R20445 vdd.n2034 vdd.n1969 19.3944
R20446 vdd.n2034 vdd.n1975 19.3944
R20447 vdd.n2029 vdd.n1975 19.3944
R20448 vdd.n2029 vdd.n2028 19.3944
R20449 vdd.n2028 vdd.n2027 19.3944
R20450 vdd.n2027 vdd.n1982 19.3944
R20451 vdd.n2022 vdd.n1982 19.3944
R20452 vdd.n2022 vdd.n2021 19.3944
R20453 vdd.n2021 vdd.n2020 19.3944
R20454 vdd.n2020 vdd.n1989 19.3944
R20455 vdd.n2015 vdd.n1989 19.3944
R20456 vdd.n2015 vdd.n2014 19.3944
R20457 vdd.n2014 vdd.n2013 19.3944
R20458 vdd.n2013 vdd.n1997 19.3944
R20459 vdd.n2008 vdd.n1997 19.3944
R20460 vdd.n2008 vdd.n2007 19.3944
R20461 vdd.n2003 vdd.n2002 19.3944
R20462 vdd.n2336 vdd.n1068 19.3944
R20463 vdd.n2073 vdd.n1929 19.3944
R20464 vdd.n2073 vdd.n1935 19.3944
R20465 vdd.n2068 vdd.n1935 19.3944
R20466 vdd.n2068 vdd.n2067 19.3944
R20467 vdd.n2067 vdd.n2066 19.3944
R20468 vdd.n2066 vdd.n1942 19.3944
R20469 vdd.n2061 vdd.n1942 19.3944
R20470 vdd.n2061 vdd.n2060 19.3944
R20471 vdd.n2060 vdd.n2059 19.3944
R20472 vdd.n2059 vdd.n1949 19.3944
R20473 vdd.n2054 vdd.n1949 19.3944
R20474 vdd.n2054 vdd.n2053 19.3944
R20475 vdd.n2053 vdd.n2052 19.3944
R20476 vdd.n2052 vdd.n1956 19.3944
R20477 vdd.n2047 vdd.n1956 19.3944
R20478 vdd.n2047 vdd.n2046 19.3944
R20479 vdd.n2046 vdd.n2045 19.3944
R20480 vdd.n2045 vdd.n1963 19.3944
R20481 vdd.n2040 vdd.n1963 19.3944
R20482 vdd.n2040 vdd.n2039 19.3944
R20483 vdd.n2324 vdd.n2323 19.3944
R20484 vdd.n2323 vdd.n1901 19.3944
R20485 vdd.n2318 vdd.n2317 19.3944
R20486 vdd.n2100 vdd.n1905 19.3944
R20487 vdd.n2100 vdd.n1907 19.3944
R20488 vdd.n1910 vdd.n1907 19.3944
R20489 vdd.n2093 vdd.n1910 19.3944
R20490 vdd.n2093 vdd.n2092 19.3944
R20491 vdd.n2092 vdd.n2091 19.3944
R20492 vdd.n2091 vdd.n1916 19.3944
R20493 vdd.n2086 vdd.n1916 19.3944
R20494 vdd.n2086 vdd.n2085 19.3944
R20495 vdd.n2085 vdd.n2084 19.3944
R20496 vdd.n2084 vdd.n1923 19.3944
R20497 vdd.n2079 vdd.n1923 19.3944
R20498 vdd.n2079 vdd.n2078 19.3944
R20499 vdd.n1425 vdd.n1190 19.3944
R20500 vdd.n1425 vdd.n1181 19.3944
R20501 vdd.n1438 vdd.n1181 19.3944
R20502 vdd.n1438 vdd.n1179 19.3944
R20503 vdd.n1442 vdd.n1179 19.3944
R20504 vdd.n1442 vdd.n1170 19.3944
R20505 vdd.n1455 vdd.n1170 19.3944
R20506 vdd.n1455 vdd.n1168 19.3944
R20507 vdd.n1459 vdd.n1168 19.3944
R20508 vdd.n1459 vdd.n1159 19.3944
R20509 vdd.n1471 vdd.n1159 19.3944
R20510 vdd.n1471 vdd.n1157 19.3944
R20511 vdd.n1475 vdd.n1157 19.3944
R20512 vdd.n1475 vdd.n1147 19.3944
R20513 vdd.n1488 vdd.n1147 19.3944
R20514 vdd.n1488 vdd.n1145 19.3944
R20515 vdd.n1492 vdd.n1145 19.3944
R20516 vdd.n1492 vdd.n1136 19.3944
R20517 vdd.n1504 vdd.n1136 19.3944
R20518 vdd.n1504 vdd.n1134 19.3944
R20519 vdd.n1815 vdd.n1134 19.3944
R20520 vdd.n1815 vdd.n1124 19.3944
R20521 vdd.n1828 vdd.n1124 19.3944
R20522 vdd.n1828 vdd.n1122 19.3944
R20523 vdd.n1832 vdd.n1122 19.3944
R20524 vdd.n1832 vdd.n1113 19.3944
R20525 vdd.n1845 vdd.n1113 19.3944
R20526 vdd.n1845 vdd.n1111 19.3944
R20527 vdd.n1849 vdd.n1111 19.3944
R20528 vdd.n1849 vdd.n1102 19.3944
R20529 vdd.n1861 vdd.n1102 19.3944
R20530 vdd.n1861 vdd.n1100 19.3944
R20531 vdd.n1865 vdd.n1100 19.3944
R20532 vdd.n1865 vdd.n1090 19.3944
R20533 vdd.n1878 vdd.n1090 19.3944
R20534 vdd.n1878 vdd.n1088 19.3944
R20535 vdd.n1882 vdd.n1088 19.3944
R20536 vdd.n1882 vdd.n1078 19.3944
R20537 vdd.n1897 vdd.n1078 19.3944
R20538 vdd.n1897 vdd.n1076 19.3944
R20539 vdd.n2327 vdd.n1076 19.3944
R20540 vdd.n3229 vdd.n686 19.3944
R20541 vdd.n3229 vdd.n676 19.3944
R20542 vdd.n3241 vdd.n676 19.3944
R20543 vdd.n3241 vdd.n674 19.3944
R20544 vdd.n3245 vdd.n674 19.3944
R20545 vdd.n3245 vdd.n666 19.3944
R20546 vdd.n3258 vdd.n666 19.3944
R20547 vdd.n3258 vdd.n664 19.3944
R20548 vdd.n3262 vdd.n664 19.3944
R20549 vdd.n3262 vdd.n653 19.3944
R20550 vdd.n3274 vdd.n653 19.3944
R20551 vdd.n3274 vdd.n651 19.3944
R20552 vdd.n3278 vdd.n651 19.3944
R20553 vdd.n3278 vdd.n642 19.3944
R20554 vdd.n3291 vdd.n642 19.3944
R20555 vdd.n3291 vdd.n640 19.3944
R20556 vdd.n3298 vdd.n640 19.3944
R20557 vdd.n3298 vdd.n3297 19.3944
R20558 vdd.n3297 vdd.n631 19.3944
R20559 vdd.n3311 vdd.n631 19.3944
R20560 vdd.n3312 vdd.n3311 19.3944
R20561 vdd.n3312 vdd.n629 19.3944
R20562 vdd.n3316 vdd.n629 19.3944
R20563 vdd.n3318 vdd.n3316 19.3944
R20564 vdd.n3319 vdd.n3318 19.3944
R20565 vdd.n3319 vdd.n627 19.3944
R20566 vdd.n3323 vdd.n627 19.3944
R20567 vdd.n3325 vdd.n3323 19.3944
R20568 vdd.n3326 vdd.n3325 19.3944
R20569 vdd.n3326 vdd.n625 19.3944
R20570 vdd.n3330 vdd.n625 19.3944
R20571 vdd.n3333 vdd.n3330 19.3944
R20572 vdd.n3334 vdd.n3333 19.3944
R20573 vdd.n3334 vdd.n623 19.3944
R20574 vdd.n3338 vdd.n623 19.3944
R20575 vdd.n3340 vdd.n3338 19.3944
R20576 vdd.n3341 vdd.n3340 19.3944
R20577 vdd.n3341 vdd.n621 19.3944
R20578 vdd.n3345 vdd.n621 19.3944
R20579 vdd.n3347 vdd.n3345 19.3944
R20580 vdd.n3348 vdd.n3347 19.3944
R20581 vdd.n569 vdd.n438 19.3944
R20582 vdd.n575 vdd.n438 19.3944
R20583 vdd.n576 vdd.n575 19.3944
R20584 vdd.n579 vdd.n576 19.3944
R20585 vdd.n579 vdd.n436 19.3944
R20586 vdd.n585 vdd.n436 19.3944
R20587 vdd.n586 vdd.n585 19.3944
R20588 vdd.n589 vdd.n586 19.3944
R20589 vdd.n589 vdd.n434 19.3944
R20590 vdd.n595 vdd.n434 19.3944
R20591 vdd.n596 vdd.n595 19.3944
R20592 vdd.n599 vdd.n596 19.3944
R20593 vdd.n599 vdd.n432 19.3944
R20594 vdd.n605 vdd.n432 19.3944
R20595 vdd.n606 vdd.n605 19.3944
R20596 vdd.n609 vdd.n606 19.3944
R20597 vdd.n609 vdd.n430 19.3944
R20598 vdd.n615 vdd.n430 19.3944
R20599 vdd.n617 vdd.n615 19.3944
R20600 vdd.n618 vdd.n617 19.3944
R20601 vdd.n516 vdd.n515 19.3944
R20602 vdd.n519 vdd.n516 19.3944
R20603 vdd.n519 vdd.n450 19.3944
R20604 vdd.n525 vdd.n450 19.3944
R20605 vdd.n526 vdd.n525 19.3944
R20606 vdd.n529 vdd.n526 19.3944
R20607 vdd.n529 vdd.n448 19.3944
R20608 vdd.n535 vdd.n448 19.3944
R20609 vdd.n536 vdd.n535 19.3944
R20610 vdd.n539 vdd.n536 19.3944
R20611 vdd.n539 vdd.n446 19.3944
R20612 vdd.n545 vdd.n446 19.3944
R20613 vdd.n546 vdd.n545 19.3944
R20614 vdd.n549 vdd.n546 19.3944
R20615 vdd.n549 vdd.n444 19.3944
R20616 vdd.n555 vdd.n444 19.3944
R20617 vdd.n556 vdd.n555 19.3944
R20618 vdd.n559 vdd.n556 19.3944
R20619 vdd.n559 vdd.n442 19.3944
R20620 vdd.n565 vdd.n442 19.3944
R20621 vdd.n466 vdd.n465 19.3944
R20622 vdd.n469 vdd.n466 19.3944
R20623 vdd.n469 vdd.n462 19.3944
R20624 vdd.n475 vdd.n462 19.3944
R20625 vdd.n476 vdd.n475 19.3944
R20626 vdd.n479 vdd.n476 19.3944
R20627 vdd.n479 vdd.n460 19.3944
R20628 vdd.n485 vdd.n460 19.3944
R20629 vdd.n486 vdd.n485 19.3944
R20630 vdd.n489 vdd.n486 19.3944
R20631 vdd.n489 vdd.n458 19.3944
R20632 vdd.n495 vdd.n458 19.3944
R20633 vdd.n496 vdd.n495 19.3944
R20634 vdd.n499 vdd.n496 19.3944
R20635 vdd.n499 vdd.n456 19.3944
R20636 vdd.n505 vdd.n456 19.3944
R20637 vdd.n506 vdd.n505 19.3944
R20638 vdd.n509 vdd.n506 19.3944
R20639 vdd.n3233 vdd.n683 19.3944
R20640 vdd.n3233 vdd.n681 19.3944
R20641 vdd.n3237 vdd.n681 19.3944
R20642 vdd.n3237 vdd.n671 19.3944
R20643 vdd.n3250 vdd.n671 19.3944
R20644 vdd.n3250 vdd.n669 19.3944
R20645 vdd.n3254 vdd.n669 19.3944
R20646 vdd.n3254 vdd.n660 19.3944
R20647 vdd.n3266 vdd.n660 19.3944
R20648 vdd.n3266 vdd.n658 19.3944
R20649 vdd.n3270 vdd.n658 19.3944
R20650 vdd.n3270 vdd.n648 19.3944
R20651 vdd.n3283 vdd.n648 19.3944
R20652 vdd.n3283 vdd.n646 19.3944
R20653 vdd.n3287 vdd.n646 19.3944
R20654 vdd.n3287 vdd.n637 19.3944
R20655 vdd.n3302 vdd.n637 19.3944
R20656 vdd.n3302 vdd.n635 19.3944
R20657 vdd.n3306 vdd.n635 19.3944
R20658 vdd.n3306 vdd.n336 19.3944
R20659 vdd.n3397 vdd.n336 19.3944
R20660 vdd.n3397 vdd.n337 19.3944
R20661 vdd.n3391 vdd.n337 19.3944
R20662 vdd.n3391 vdd.n3390 19.3944
R20663 vdd.n3390 vdd.n3389 19.3944
R20664 vdd.n3389 vdd.n349 19.3944
R20665 vdd.n3383 vdd.n349 19.3944
R20666 vdd.n3383 vdd.n3382 19.3944
R20667 vdd.n3382 vdd.n3381 19.3944
R20668 vdd.n3381 vdd.n359 19.3944
R20669 vdd.n3375 vdd.n359 19.3944
R20670 vdd.n3375 vdd.n3374 19.3944
R20671 vdd.n3374 vdd.n3373 19.3944
R20672 vdd.n3373 vdd.n370 19.3944
R20673 vdd.n3367 vdd.n370 19.3944
R20674 vdd.n3367 vdd.n3366 19.3944
R20675 vdd.n3366 vdd.n3365 19.3944
R20676 vdd.n3365 vdd.n381 19.3944
R20677 vdd.n3359 vdd.n381 19.3944
R20678 vdd.n3359 vdd.n3358 19.3944
R20679 vdd.n3358 vdd.n3357 19.3944
R20680 vdd.n3180 vdd.n747 19.3944
R20681 vdd.n3180 vdd.n3177 19.3944
R20682 vdd.n3177 vdd.n3174 19.3944
R20683 vdd.n3174 vdd.n3173 19.3944
R20684 vdd.n3173 vdd.n3170 19.3944
R20685 vdd.n3170 vdd.n3169 19.3944
R20686 vdd.n3169 vdd.n3166 19.3944
R20687 vdd.n3166 vdd.n3165 19.3944
R20688 vdd.n3165 vdd.n3162 19.3944
R20689 vdd.n3162 vdd.n3161 19.3944
R20690 vdd.n3161 vdd.n3158 19.3944
R20691 vdd.n3158 vdd.n3157 19.3944
R20692 vdd.n3157 vdd.n3154 19.3944
R20693 vdd.n3154 vdd.n3153 19.3944
R20694 vdd.n3153 vdd.n3150 19.3944
R20695 vdd.n3150 vdd.n3149 19.3944
R20696 vdd.n3149 vdd.n3146 19.3944
R20697 vdd.n3146 vdd.n3145 19.3944
R20698 vdd.n3145 vdd.n3142 19.3944
R20699 vdd.n3142 vdd.n3141 19.3944
R20700 vdd.n3220 vdd.n3219 19.3944
R20701 vdd.n3219 vdd.n3218 19.3944
R20702 vdd.n732 vdd.n729 19.3944
R20703 vdd.n3214 vdd.n3213 19.3944
R20704 vdd.n3213 vdd.n3210 19.3944
R20705 vdd.n3210 vdd.n3209 19.3944
R20706 vdd.n3209 vdd.n3206 19.3944
R20707 vdd.n3206 vdd.n3205 19.3944
R20708 vdd.n3205 vdd.n3202 19.3944
R20709 vdd.n3202 vdd.n3201 19.3944
R20710 vdd.n3201 vdd.n3198 19.3944
R20711 vdd.n3198 vdd.n3197 19.3944
R20712 vdd.n3197 vdd.n3194 19.3944
R20713 vdd.n3194 vdd.n3193 19.3944
R20714 vdd.n3193 vdd.n3190 19.3944
R20715 vdd.n3190 vdd.n3189 19.3944
R20716 vdd.n3134 vdd.n767 19.3944
R20717 vdd.n3134 vdd.n3131 19.3944
R20718 vdd.n3131 vdd.n3128 19.3944
R20719 vdd.n3128 vdd.n3127 19.3944
R20720 vdd.n3127 vdd.n3124 19.3944
R20721 vdd.n3124 vdd.n3123 19.3944
R20722 vdd.n3123 vdd.n3120 19.3944
R20723 vdd.n3120 vdd.n3119 19.3944
R20724 vdd.n3119 vdd.n3116 19.3944
R20725 vdd.n3116 vdd.n3115 19.3944
R20726 vdd.n3115 vdd.n3112 19.3944
R20727 vdd.n3112 vdd.n3111 19.3944
R20728 vdd.n3111 vdd.n3108 19.3944
R20729 vdd.n3108 vdd.n3107 19.3944
R20730 vdd.n3107 vdd.n3104 19.3944
R20731 vdd.n3104 vdd.n3103 19.3944
R20732 vdd.n3100 vdd.n3099 19.3944
R20733 vdd.n3096 vdd.n3095 19.3944
R20734 vdd.n1357 vdd.n1353 19.0066
R20735 vdd.n2038 vdd.n1969 19.0066
R20736 vdd.n569 vdd.n566 19.0066
R20737 vdd.n3138 vdd.n767 19.0066
R20738 vdd.n2178 vdd.n2177 16.0975
R20739 vdd.n966 vdd.n965 16.0975
R20740 vdd.n1318 vdd.n1317 16.0975
R20741 vdd.n1356 vdd.n1355 16.0975
R20742 vdd.n1252 vdd.n1251 16.0975
R20743 vdd.n2334 vdd.n2333 16.0975
R20744 vdd.n1971 vdd.n1970 16.0975
R20745 vdd.n1931 vdd.n1930 16.0975
R20746 vdd.n2152 vdd.n2151 16.0975
R20747 vdd.n958 vdd.n957 16.0975
R20748 vdd.n2643 vdd.n2642 16.0975
R20749 vdd.n427 vdd.n426 16.0975
R20750 vdd.n441 vdd.n440 16.0975
R20751 vdd.n453 vdd.n452 16.0975
R20752 vdd.n769 vdd.n768 16.0975
R20753 vdd.n3185 vdd.n3184 16.0975
R20754 vdd.n833 vdd.n832 16.0975
R20755 vdd.n2640 vdd.n2639 16.0975
R20756 vdd.n689 vdd.n688 16.0975
R20757 vdd.n800 vdd.n799 16.0975
R20758 vdd.t142 vdd.n2604 15.4182
R20759 vdd.n2857 vdd.t129 15.4182
R20760 vdd.n28 vdd.n27 14.7341
R20761 vdd.n2375 vdd.n1049 14.5112
R20762 vdd.n3059 vdd.n692 14.5112
R20763 vdd.n328 vdd.n293 13.1884
R20764 vdd.n269 vdd.n234 13.1884
R20765 vdd.n226 vdd.n191 13.1884
R20766 vdd.n167 vdd.n132 13.1884
R20767 vdd.n125 vdd.n90 13.1884
R20768 vdd.n66 vdd.n31 13.1884
R20769 vdd.n1747 vdd.n1712 13.1884
R20770 vdd.n1806 vdd.n1771 13.1884
R20771 vdd.n1645 vdd.n1610 13.1884
R20772 vdd.n1704 vdd.n1669 13.1884
R20773 vdd.n1544 vdd.n1509 13.1884
R20774 vdd.n1603 vdd.n1568 13.1884
R20775 vdd.n1388 vdd.n1253 12.9944
R20776 vdd.n1392 vdd.n1253 12.9944
R20777 vdd.n2077 vdd.n1929 12.9944
R20778 vdd.n2078 vdd.n2077 12.9944
R20779 vdd.n515 vdd.n454 12.9944
R20780 vdd.n509 vdd.n454 12.9944
R20781 vdd.n3186 vdd.n747 12.9944
R20782 vdd.n3189 vdd.n3186 12.9944
R20783 vdd.n329 vdd.n291 12.8005
R20784 vdd.n324 vdd.n295 12.8005
R20785 vdd.n270 vdd.n232 12.8005
R20786 vdd.n265 vdd.n236 12.8005
R20787 vdd.n227 vdd.n189 12.8005
R20788 vdd.n222 vdd.n193 12.8005
R20789 vdd.n168 vdd.n130 12.8005
R20790 vdd.n163 vdd.n134 12.8005
R20791 vdd.n126 vdd.n88 12.8005
R20792 vdd.n121 vdd.n92 12.8005
R20793 vdd.n67 vdd.n29 12.8005
R20794 vdd.n62 vdd.n33 12.8005
R20795 vdd.n1748 vdd.n1710 12.8005
R20796 vdd.n1743 vdd.n1714 12.8005
R20797 vdd.n1807 vdd.n1769 12.8005
R20798 vdd.n1802 vdd.n1773 12.8005
R20799 vdd.n1646 vdd.n1608 12.8005
R20800 vdd.n1641 vdd.n1612 12.8005
R20801 vdd.n1705 vdd.n1667 12.8005
R20802 vdd.n1700 vdd.n1671 12.8005
R20803 vdd.n1545 vdd.n1507 12.8005
R20804 vdd.n1540 vdd.n1511 12.8005
R20805 vdd.n1604 vdd.n1566 12.8005
R20806 vdd.n1599 vdd.n1570 12.8005
R20807 vdd.n323 vdd.n296 12.0247
R20808 vdd.n264 vdd.n237 12.0247
R20809 vdd.n221 vdd.n194 12.0247
R20810 vdd.n162 vdd.n135 12.0247
R20811 vdd.n120 vdd.n93 12.0247
R20812 vdd.n61 vdd.n34 12.0247
R20813 vdd.n1742 vdd.n1715 12.0247
R20814 vdd.n1801 vdd.n1774 12.0247
R20815 vdd.n1640 vdd.n1613 12.0247
R20816 vdd.n1699 vdd.n1672 12.0247
R20817 vdd.n1539 vdd.n1512 12.0247
R20818 vdd.n1598 vdd.n1571 12.0247
R20819 vdd.n1427 vdd.n1183 11.337
R20820 vdd.n1436 vdd.n1183 11.337
R20821 vdd.n1436 vdd.n1435 11.337
R20822 vdd.n1444 vdd.n1177 11.337
R20823 vdd.n1453 vdd.n1452 11.337
R20824 vdd.n1469 vdd.n1161 11.337
R20825 vdd.n1477 vdd.n1154 11.337
R20826 vdd.n1486 vdd.n1485 11.337
R20827 vdd.n1494 vdd.n1143 11.337
R20828 vdd.n1817 vdd.n1132 11.337
R20829 vdd.n1826 vdd.n1126 11.337
R20830 vdd.n1834 vdd.n1120 11.337
R20831 vdd.n1843 vdd.n1842 11.337
R20832 vdd.n1859 vdd.n1104 11.337
R20833 vdd.n1867 vdd.n1097 11.337
R20834 vdd.n1876 vdd.n1875 11.337
R20835 vdd.n1884 vdd.n1080 11.337
R20836 vdd.n1895 vdd.n1080 11.337
R20837 vdd.n1895 vdd.n1894 11.337
R20838 vdd.n3231 vdd.n678 11.337
R20839 vdd.n3239 vdd.n678 11.337
R20840 vdd.n3239 vdd.n679 11.337
R20841 vdd.n3248 vdd.n3247 11.337
R20842 vdd.n3264 vdd.n662 11.337
R20843 vdd.n3272 vdd.n655 11.337
R20844 vdd.n3281 vdd.n3280 11.337
R20845 vdd.n3289 vdd.n644 11.337
R20846 vdd.n3308 vdd.n633 11.337
R20847 vdd.n3395 vdd.n340 11.337
R20848 vdd.n3393 vdd.n344 11.337
R20849 vdd.n3387 vdd.n3386 11.337
R20850 vdd.n3379 vdd.n361 11.337
R20851 vdd.n3378 vdd.n3377 11.337
R20852 vdd.n3371 vdd.n3370 11.337
R20853 vdd.n3369 vdd.n375 11.337
R20854 vdd.n3363 vdd.n3362 11.337
R20855 vdd.n3362 vdd.n3361 11.337
R20856 vdd.n3361 vdd.n386 11.337
R20857 vdd.n320 vdd.n319 11.249
R20858 vdd.n261 vdd.n260 11.249
R20859 vdd.n218 vdd.n217 11.249
R20860 vdd.n159 vdd.n158 11.249
R20861 vdd.n117 vdd.n116 11.249
R20862 vdd.n58 vdd.n57 11.249
R20863 vdd.n1739 vdd.n1738 11.249
R20864 vdd.n1798 vdd.n1797 11.249
R20865 vdd.n1637 vdd.n1636 11.249
R20866 vdd.n1696 vdd.n1695 11.249
R20867 vdd.n1536 vdd.n1535 11.249
R20868 vdd.n1595 vdd.n1594 11.249
R20869 vdd.n1225 vdd.t185 11.2237
R20870 vdd.n3355 vdd.t192 11.2237
R20871 vdd.n2532 vdd.t157 11.1103
R20872 vdd.n2864 vdd.t145 11.1103
R20873 vdd.t45 vdd.n1098 10.7702
R20874 vdd.n3256 vdd.t271 10.7702
R20875 vdd.n305 vdd.n304 10.7238
R20876 vdd.n246 vdd.n245 10.7238
R20877 vdd.n203 vdd.n202 10.7238
R20878 vdd.n144 vdd.n143 10.7238
R20879 vdd.n102 vdd.n101 10.7238
R20880 vdd.n43 vdd.n42 10.7238
R20881 vdd.n1724 vdd.n1723 10.7238
R20882 vdd.n1783 vdd.n1782 10.7238
R20883 vdd.n1622 vdd.n1621 10.7238
R20884 vdd.n1681 vdd.n1680 10.7238
R20885 vdd.n1521 vdd.n1520 10.7238
R20886 vdd.n1580 vdd.n1579 10.7238
R20887 vdd.n2378 vdd.n2377 10.6151
R20888 vdd.n2379 vdd.n2378 10.6151
R20889 vdd.n2379 vdd.n1035 10.6151
R20890 vdd.n2389 vdd.n1035 10.6151
R20891 vdd.n2390 vdd.n2389 10.6151
R20892 vdd.n2391 vdd.n2390 10.6151
R20893 vdd.n2391 vdd.n1022 10.6151
R20894 vdd.n2402 vdd.n1022 10.6151
R20895 vdd.n2403 vdd.n2402 10.6151
R20896 vdd.n2404 vdd.n2403 10.6151
R20897 vdd.n2404 vdd.n1010 10.6151
R20898 vdd.n2414 vdd.n1010 10.6151
R20899 vdd.n2415 vdd.n2414 10.6151
R20900 vdd.n2416 vdd.n2415 10.6151
R20901 vdd.n2416 vdd.n998 10.6151
R20902 vdd.n2426 vdd.n998 10.6151
R20903 vdd.n2427 vdd.n2426 10.6151
R20904 vdd.n2428 vdd.n2427 10.6151
R20905 vdd.n2428 vdd.n987 10.6151
R20906 vdd.n2438 vdd.n987 10.6151
R20907 vdd.n2439 vdd.n2438 10.6151
R20908 vdd.n2440 vdd.n2439 10.6151
R20909 vdd.n2440 vdd.n974 10.6151
R20910 vdd.n2452 vdd.n974 10.6151
R20911 vdd.n2453 vdd.n2452 10.6151
R20912 vdd.n2455 vdd.n2453 10.6151
R20913 vdd.n2455 vdd.n2454 10.6151
R20914 vdd.n2454 vdd.n956 10.6151
R20915 vdd.n2602 vdd.n2601 10.6151
R20916 vdd.n2601 vdd.n2600 10.6151
R20917 vdd.n2600 vdd.n2597 10.6151
R20918 vdd.n2597 vdd.n2596 10.6151
R20919 vdd.n2596 vdd.n2593 10.6151
R20920 vdd.n2593 vdd.n2592 10.6151
R20921 vdd.n2592 vdd.n2589 10.6151
R20922 vdd.n2589 vdd.n2588 10.6151
R20923 vdd.n2588 vdd.n2585 10.6151
R20924 vdd.n2585 vdd.n2584 10.6151
R20925 vdd.n2584 vdd.n2581 10.6151
R20926 vdd.n2581 vdd.n2580 10.6151
R20927 vdd.n2580 vdd.n2577 10.6151
R20928 vdd.n2577 vdd.n2576 10.6151
R20929 vdd.n2576 vdd.n2573 10.6151
R20930 vdd.n2573 vdd.n2572 10.6151
R20931 vdd.n2572 vdd.n2569 10.6151
R20932 vdd.n2569 vdd.n2568 10.6151
R20933 vdd.n2568 vdd.n2565 10.6151
R20934 vdd.n2565 vdd.n2564 10.6151
R20935 vdd.n2564 vdd.n2561 10.6151
R20936 vdd.n2561 vdd.n2560 10.6151
R20937 vdd.n2560 vdd.n2557 10.6151
R20938 vdd.n2557 vdd.n2556 10.6151
R20939 vdd.n2556 vdd.n2553 10.6151
R20940 vdd.n2553 vdd.n2552 10.6151
R20941 vdd.n2552 vdd.n2549 10.6151
R20942 vdd.n2549 vdd.n2548 10.6151
R20943 vdd.n2548 vdd.n2545 10.6151
R20944 vdd.n2545 vdd.n2544 10.6151
R20945 vdd.n2544 vdd.n2541 10.6151
R20946 vdd.n2539 vdd.n2536 10.6151
R20947 vdd.n2536 vdd.n2535 10.6151
R20948 vdd.n2278 vdd.n2277 10.6151
R20949 vdd.n2277 vdd.n2275 10.6151
R20950 vdd.n2275 vdd.n2274 10.6151
R20951 vdd.n2274 vdd.n2272 10.6151
R20952 vdd.n2272 vdd.n2271 10.6151
R20953 vdd.n2271 vdd.n2269 10.6151
R20954 vdd.n2269 vdd.n2268 10.6151
R20955 vdd.n2268 vdd.n2266 10.6151
R20956 vdd.n2266 vdd.n2265 10.6151
R20957 vdd.n2265 vdd.n2263 10.6151
R20958 vdd.n2263 vdd.n2262 10.6151
R20959 vdd.n2262 vdd.n2260 10.6151
R20960 vdd.n2260 vdd.n2259 10.6151
R20961 vdd.n2259 vdd.n2174 10.6151
R20962 vdd.n2174 vdd.n2173 10.6151
R20963 vdd.n2173 vdd.n2171 10.6151
R20964 vdd.n2171 vdd.n2170 10.6151
R20965 vdd.n2170 vdd.n2168 10.6151
R20966 vdd.n2168 vdd.n2167 10.6151
R20967 vdd.n2167 vdd.n2165 10.6151
R20968 vdd.n2165 vdd.n2164 10.6151
R20969 vdd.n2164 vdd.n2162 10.6151
R20970 vdd.n2162 vdd.n2161 10.6151
R20971 vdd.n2161 vdd.n2159 10.6151
R20972 vdd.n2159 vdd.n2158 10.6151
R20973 vdd.n2158 vdd.n2155 10.6151
R20974 vdd.n2155 vdd.n2154 10.6151
R20975 vdd.n2154 vdd.n959 10.6151
R20976 vdd.n2112 vdd.n1047 10.6151
R20977 vdd.n2113 vdd.n2112 10.6151
R20978 vdd.n2114 vdd.n2113 10.6151
R20979 vdd.n2114 vdd.n2108 10.6151
R20980 vdd.n2120 vdd.n2108 10.6151
R20981 vdd.n2121 vdd.n2120 10.6151
R20982 vdd.n2122 vdd.n2121 10.6151
R20983 vdd.n2122 vdd.n2106 10.6151
R20984 vdd.n2128 vdd.n2106 10.6151
R20985 vdd.n2129 vdd.n2128 10.6151
R20986 vdd.n2130 vdd.n2129 10.6151
R20987 vdd.n2130 vdd.n2104 10.6151
R20988 vdd.n2136 vdd.n2104 10.6151
R20989 vdd.n2137 vdd.n2136 10.6151
R20990 vdd.n2138 vdd.n2137 10.6151
R20991 vdd.n2138 vdd.n2102 10.6151
R20992 vdd.n2314 vdd.n2102 10.6151
R20993 vdd.n2314 vdd.n2313 10.6151
R20994 vdd.n2313 vdd.n2143 10.6151
R20995 vdd.n2307 vdd.n2143 10.6151
R20996 vdd.n2307 vdd.n2306 10.6151
R20997 vdd.n2306 vdd.n2305 10.6151
R20998 vdd.n2305 vdd.n2145 10.6151
R20999 vdd.n2299 vdd.n2145 10.6151
R21000 vdd.n2299 vdd.n2298 10.6151
R21001 vdd.n2298 vdd.n2297 10.6151
R21002 vdd.n2297 vdd.n2147 10.6151
R21003 vdd.n2291 vdd.n2147 10.6151
R21004 vdd.n2291 vdd.n2290 10.6151
R21005 vdd.n2290 vdd.n2289 10.6151
R21006 vdd.n2289 vdd.n2149 10.6151
R21007 vdd.n2283 vdd.n2282 10.6151
R21008 vdd.n2282 vdd.n2281 10.6151
R21009 vdd.n2787 vdd.n2786 10.6151
R21010 vdd.n2786 vdd.n2784 10.6151
R21011 vdd.n2784 vdd.n2783 10.6151
R21012 vdd.n2783 vdd.n2641 10.6151
R21013 vdd.n2730 vdd.n2641 10.6151
R21014 vdd.n2731 vdd.n2730 10.6151
R21015 vdd.n2733 vdd.n2731 10.6151
R21016 vdd.n2734 vdd.n2733 10.6151
R21017 vdd.n2736 vdd.n2734 10.6151
R21018 vdd.n2737 vdd.n2736 10.6151
R21019 vdd.n2739 vdd.n2737 10.6151
R21020 vdd.n2740 vdd.n2739 10.6151
R21021 vdd.n2742 vdd.n2740 10.6151
R21022 vdd.n2743 vdd.n2742 10.6151
R21023 vdd.n2758 vdd.n2743 10.6151
R21024 vdd.n2758 vdd.n2757 10.6151
R21025 vdd.n2757 vdd.n2756 10.6151
R21026 vdd.n2756 vdd.n2754 10.6151
R21027 vdd.n2754 vdd.n2753 10.6151
R21028 vdd.n2753 vdd.n2751 10.6151
R21029 vdd.n2751 vdd.n2750 10.6151
R21030 vdd.n2750 vdd.n2748 10.6151
R21031 vdd.n2748 vdd.n2747 10.6151
R21032 vdd.n2747 vdd.n2745 10.6151
R21033 vdd.n2745 vdd.n2744 10.6151
R21034 vdd.n2744 vdd.n836 10.6151
R21035 vdd.n2992 vdd.n836 10.6151
R21036 vdd.n2993 vdd.n2992 10.6151
R21037 vdd.n2854 vdd.n912 10.6151
R21038 vdd.n2854 vdd.n2853 10.6151
R21039 vdd.n2853 vdd.n2852 10.6151
R21040 vdd.n2852 vdd.n2850 10.6151
R21041 vdd.n2850 vdd.n2847 10.6151
R21042 vdd.n2847 vdd.n2846 10.6151
R21043 vdd.n2846 vdd.n2843 10.6151
R21044 vdd.n2843 vdd.n2842 10.6151
R21045 vdd.n2842 vdd.n2839 10.6151
R21046 vdd.n2839 vdd.n2838 10.6151
R21047 vdd.n2838 vdd.n2835 10.6151
R21048 vdd.n2835 vdd.n2834 10.6151
R21049 vdd.n2834 vdd.n2831 10.6151
R21050 vdd.n2831 vdd.n2830 10.6151
R21051 vdd.n2830 vdd.n2827 10.6151
R21052 vdd.n2827 vdd.n2826 10.6151
R21053 vdd.n2826 vdd.n2823 10.6151
R21054 vdd.n2823 vdd.n2822 10.6151
R21055 vdd.n2822 vdd.n2819 10.6151
R21056 vdd.n2819 vdd.n2818 10.6151
R21057 vdd.n2818 vdd.n2815 10.6151
R21058 vdd.n2815 vdd.n2814 10.6151
R21059 vdd.n2814 vdd.n2811 10.6151
R21060 vdd.n2811 vdd.n2810 10.6151
R21061 vdd.n2810 vdd.n2807 10.6151
R21062 vdd.n2807 vdd.n2806 10.6151
R21063 vdd.n2806 vdd.n2803 10.6151
R21064 vdd.n2803 vdd.n2802 10.6151
R21065 vdd.n2802 vdd.n2799 10.6151
R21066 vdd.n2799 vdd.n2798 10.6151
R21067 vdd.n2798 vdd.n2795 10.6151
R21068 vdd.n2793 vdd.n2790 10.6151
R21069 vdd.n2790 vdd.n2789 10.6151
R21070 vdd.n2867 vdd.n2866 10.6151
R21071 vdd.n2868 vdd.n2867 10.6151
R21072 vdd.n2868 vdd.n902 10.6151
R21073 vdd.n2878 vdd.n902 10.6151
R21074 vdd.n2879 vdd.n2878 10.6151
R21075 vdd.n2880 vdd.n2879 10.6151
R21076 vdd.n2880 vdd.n889 10.6151
R21077 vdd.n2890 vdd.n889 10.6151
R21078 vdd.n2891 vdd.n2890 10.6151
R21079 vdd.n2892 vdd.n2891 10.6151
R21080 vdd.n2892 vdd.n878 10.6151
R21081 vdd.n2902 vdd.n878 10.6151
R21082 vdd.n2903 vdd.n2902 10.6151
R21083 vdd.n2904 vdd.n2903 10.6151
R21084 vdd.n2904 vdd.n866 10.6151
R21085 vdd.n2914 vdd.n866 10.6151
R21086 vdd.n2915 vdd.n2914 10.6151
R21087 vdd.n2916 vdd.n2915 10.6151
R21088 vdd.n2916 vdd.n855 10.6151
R21089 vdd.n2928 vdd.n855 10.6151
R21090 vdd.n2929 vdd.n2928 10.6151
R21091 vdd.n2930 vdd.n2929 10.6151
R21092 vdd.n2930 vdd.n841 10.6151
R21093 vdd.n2985 vdd.n841 10.6151
R21094 vdd.n2986 vdd.n2985 10.6151
R21095 vdd.n2987 vdd.n2986 10.6151
R21096 vdd.n2987 vdd.n810 10.6151
R21097 vdd.n3057 vdd.n810 10.6151
R21098 vdd.n3056 vdd.n3055 10.6151
R21099 vdd.n3055 vdd.n811 10.6151
R21100 vdd.n812 vdd.n811 10.6151
R21101 vdd.n3048 vdd.n812 10.6151
R21102 vdd.n3048 vdd.n3047 10.6151
R21103 vdd.n3047 vdd.n3046 10.6151
R21104 vdd.n3046 vdd.n814 10.6151
R21105 vdd.n3041 vdd.n814 10.6151
R21106 vdd.n3041 vdd.n3040 10.6151
R21107 vdd.n3040 vdd.n3039 10.6151
R21108 vdd.n3039 vdd.n817 10.6151
R21109 vdd.n3034 vdd.n817 10.6151
R21110 vdd.n3034 vdd.n3033 10.6151
R21111 vdd.n3033 vdd.n3032 10.6151
R21112 vdd.n3032 vdd.n820 10.6151
R21113 vdd.n3027 vdd.n820 10.6151
R21114 vdd.n3027 vdd.n731 10.6151
R21115 vdd.n3023 vdd.n731 10.6151
R21116 vdd.n3023 vdd.n3022 10.6151
R21117 vdd.n3022 vdd.n3021 10.6151
R21118 vdd.n3021 vdd.n823 10.6151
R21119 vdd.n3016 vdd.n823 10.6151
R21120 vdd.n3016 vdd.n3015 10.6151
R21121 vdd.n3015 vdd.n3014 10.6151
R21122 vdd.n3014 vdd.n826 10.6151
R21123 vdd.n3009 vdd.n826 10.6151
R21124 vdd.n3009 vdd.n3008 10.6151
R21125 vdd.n3008 vdd.n3007 10.6151
R21126 vdd.n3007 vdd.n829 10.6151
R21127 vdd.n3002 vdd.n829 10.6151
R21128 vdd.n3002 vdd.n3001 10.6151
R21129 vdd.n2999 vdd.n834 10.6151
R21130 vdd.n2994 vdd.n834 10.6151
R21131 vdd.n2975 vdd.n2936 10.6151
R21132 vdd.n2970 vdd.n2936 10.6151
R21133 vdd.n2970 vdd.n2969 10.6151
R21134 vdd.n2969 vdd.n2968 10.6151
R21135 vdd.n2968 vdd.n2938 10.6151
R21136 vdd.n2963 vdd.n2938 10.6151
R21137 vdd.n2963 vdd.n2962 10.6151
R21138 vdd.n2962 vdd.n2961 10.6151
R21139 vdd.n2961 vdd.n2941 10.6151
R21140 vdd.n2956 vdd.n2941 10.6151
R21141 vdd.n2956 vdd.n2955 10.6151
R21142 vdd.n2955 vdd.n2954 10.6151
R21143 vdd.n2954 vdd.n2944 10.6151
R21144 vdd.n2949 vdd.n2944 10.6151
R21145 vdd.n2949 vdd.n2948 10.6151
R21146 vdd.n2948 vdd.n785 10.6151
R21147 vdd.n3092 vdd.n785 10.6151
R21148 vdd.n3092 vdd.n786 10.6151
R21149 vdd.n788 vdd.n786 10.6151
R21150 vdd.n3085 vdd.n788 10.6151
R21151 vdd.n3085 vdd.n3084 10.6151
R21152 vdd.n3084 vdd.n3083 10.6151
R21153 vdd.n3083 vdd.n790 10.6151
R21154 vdd.n3078 vdd.n790 10.6151
R21155 vdd.n3078 vdd.n3077 10.6151
R21156 vdd.n3077 vdd.n3076 10.6151
R21157 vdd.n3076 vdd.n793 10.6151
R21158 vdd.n3071 vdd.n793 10.6151
R21159 vdd.n3071 vdd.n3070 10.6151
R21160 vdd.n3070 vdd.n3069 10.6151
R21161 vdd.n3069 vdd.n796 10.6151
R21162 vdd.n3064 vdd.n3063 10.6151
R21163 vdd.n3063 vdd.n3062 10.6151
R21164 vdd.n2710 vdd.n2708 10.6151
R21165 vdd.n2711 vdd.n2710 10.6151
R21166 vdd.n2779 vdd.n2711 10.6151
R21167 vdd.n2779 vdd.n2778 10.6151
R21168 vdd.n2778 vdd.n2777 10.6151
R21169 vdd.n2777 vdd.n2775 10.6151
R21170 vdd.n2775 vdd.n2774 10.6151
R21171 vdd.n2774 vdd.n2772 10.6151
R21172 vdd.n2772 vdd.n2771 10.6151
R21173 vdd.n2771 vdd.n2769 10.6151
R21174 vdd.n2769 vdd.n2768 10.6151
R21175 vdd.n2768 vdd.n2766 10.6151
R21176 vdd.n2766 vdd.n2765 10.6151
R21177 vdd.n2765 vdd.n2763 10.6151
R21178 vdd.n2763 vdd.n2762 10.6151
R21179 vdd.n2762 vdd.n2728 10.6151
R21180 vdd.n2728 vdd.n2727 10.6151
R21181 vdd.n2727 vdd.n2725 10.6151
R21182 vdd.n2725 vdd.n2724 10.6151
R21183 vdd.n2724 vdd.n2722 10.6151
R21184 vdd.n2722 vdd.n2721 10.6151
R21185 vdd.n2721 vdd.n2719 10.6151
R21186 vdd.n2719 vdd.n2718 10.6151
R21187 vdd.n2718 vdd.n2716 10.6151
R21188 vdd.n2716 vdd.n2715 10.6151
R21189 vdd.n2715 vdd.n2713 10.6151
R21190 vdd.n2713 vdd.n2712 10.6151
R21191 vdd.n2712 vdd.n802 10.6151
R21192 vdd.n2861 vdd.n2860 10.6151
R21193 vdd.n2860 vdd.n917 10.6151
R21194 vdd.n2645 vdd.n917 10.6151
R21195 vdd.n2648 vdd.n2645 10.6151
R21196 vdd.n2649 vdd.n2648 10.6151
R21197 vdd.n2652 vdd.n2649 10.6151
R21198 vdd.n2653 vdd.n2652 10.6151
R21199 vdd.n2656 vdd.n2653 10.6151
R21200 vdd.n2657 vdd.n2656 10.6151
R21201 vdd.n2660 vdd.n2657 10.6151
R21202 vdd.n2661 vdd.n2660 10.6151
R21203 vdd.n2664 vdd.n2661 10.6151
R21204 vdd.n2665 vdd.n2664 10.6151
R21205 vdd.n2668 vdd.n2665 10.6151
R21206 vdd.n2669 vdd.n2668 10.6151
R21207 vdd.n2672 vdd.n2669 10.6151
R21208 vdd.n2673 vdd.n2672 10.6151
R21209 vdd.n2676 vdd.n2673 10.6151
R21210 vdd.n2677 vdd.n2676 10.6151
R21211 vdd.n2680 vdd.n2677 10.6151
R21212 vdd.n2681 vdd.n2680 10.6151
R21213 vdd.n2684 vdd.n2681 10.6151
R21214 vdd.n2685 vdd.n2684 10.6151
R21215 vdd.n2688 vdd.n2685 10.6151
R21216 vdd.n2689 vdd.n2688 10.6151
R21217 vdd.n2692 vdd.n2689 10.6151
R21218 vdd.n2693 vdd.n2692 10.6151
R21219 vdd.n2696 vdd.n2693 10.6151
R21220 vdd.n2697 vdd.n2696 10.6151
R21221 vdd.n2700 vdd.n2697 10.6151
R21222 vdd.n2701 vdd.n2700 10.6151
R21223 vdd.n2706 vdd.n2704 10.6151
R21224 vdd.n2707 vdd.n2706 10.6151
R21225 vdd.n2862 vdd.n907 10.6151
R21226 vdd.n2872 vdd.n907 10.6151
R21227 vdd.n2873 vdd.n2872 10.6151
R21228 vdd.n2874 vdd.n2873 10.6151
R21229 vdd.n2874 vdd.n895 10.6151
R21230 vdd.n2884 vdd.n895 10.6151
R21231 vdd.n2885 vdd.n2884 10.6151
R21232 vdd.n2886 vdd.n2885 10.6151
R21233 vdd.n2886 vdd.n884 10.6151
R21234 vdd.n2896 vdd.n884 10.6151
R21235 vdd.n2897 vdd.n2896 10.6151
R21236 vdd.n2898 vdd.n2897 10.6151
R21237 vdd.n2898 vdd.n872 10.6151
R21238 vdd.n2908 vdd.n872 10.6151
R21239 vdd.n2909 vdd.n2908 10.6151
R21240 vdd.n2910 vdd.n2909 10.6151
R21241 vdd.n2910 vdd.n861 10.6151
R21242 vdd.n2920 vdd.n861 10.6151
R21243 vdd.n2921 vdd.n2920 10.6151
R21244 vdd.n2924 vdd.n2921 10.6151
R21245 vdd.n2934 vdd.n849 10.6151
R21246 vdd.n2935 vdd.n2934 10.6151
R21247 vdd.n2981 vdd.n2935 10.6151
R21248 vdd.n2981 vdd.n2980 10.6151
R21249 vdd.n2980 vdd.n2979 10.6151
R21250 vdd.n2979 vdd.n2978 10.6151
R21251 vdd.n2978 vdd.n2976 10.6151
R21252 vdd.n2373 vdd.n1041 10.6151
R21253 vdd.n2383 vdd.n1041 10.6151
R21254 vdd.n2384 vdd.n2383 10.6151
R21255 vdd.n2385 vdd.n2384 10.6151
R21256 vdd.n2385 vdd.n1028 10.6151
R21257 vdd.n2395 vdd.n1028 10.6151
R21258 vdd.n2396 vdd.n2395 10.6151
R21259 vdd.n2398 vdd.n1016 10.6151
R21260 vdd.n2408 vdd.n1016 10.6151
R21261 vdd.n2409 vdd.n2408 10.6151
R21262 vdd.n2410 vdd.n2409 10.6151
R21263 vdd.n2410 vdd.n1004 10.6151
R21264 vdd.n2420 vdd.n1004 10.6151
R21265 vdd.n2421 vdd.n2420 10.6151
R21266 vdd.n2422 vdd.n2421 10.6151
R21267 vdd.n2422 vdd.n993 10.6151
R21268 vdd.n2432 vdd.n993 10.6151
R21269 vdd.n2433 vdd.n2432 10.6151
R21270 vdd.n2434 vdd.n2433 10.6151
R21271 vdd.n2434 vdd.n981 10.6151
R21272 vdd.n2444 vdd.n981 10.6151
R21273 vdd.n2445 vdd.n2444 10.6151
R21274 vdd.n2448 vdd.n2445 10.6151
R21275 vdd.n2448 vdd.n2447 10.6151
R21276 vdd.n2447 vdd.n2446 10.6151
R21277 vdd.n2446 vdd.n964 10.6151
R21278 vdd.n2530 vdd.n964 10.6151
R21279 vdd.n2529 vdd.n2528 10.6151
R21280 vdd.n2528 vdd.n2525 10.6151
R21281 vdd.n2525 vdd.n2524 10.6151
R21282 vdd.n2524 vdd.n2521 10.6151
R21283 vdd.n2521 vdd.n2520 10.6151
R21284 vdd.n2520 vdd.n2517 10.6151
R21285 vdd.n2517 vdd.n2516 10.6151
R21286 vdd.n2516 vdd.n2513 10.6151
R21287 vdd.n2513 vdd.n2512 10.6151
R21288 vdd.n2512 vdd.n2509 10.6151
R21289 vdd.n2509 vdd.n2508 10.6151
R21290 vdd.n2508 vdd.n2505 10.6151
R21291 vdd.n2505 vdd.n2504 10.6151
R21292 vdd.n2504 vdd.n2501 10.6151
R21293 vdd.n2501 vdd.n2500 10.6151
R21294 vdd.n2500 vdd.n2497 10.6151
R21295 vdd.n2497 vdd.n2496 10.6151
R21296 vdd.n2496 vdd.n2493 10.6151
R21297 vdd.n2493 vdd.n2492 10.6151
R21298 vdd.n2492 vdd.n2489 10.6151
R21299 vdd.n2489 vdd.n2488 10.6151
R21300 vdd.n2488 vdd.n2485 10.6151
R21301 vdd.n2485 vdd.n2484 10.6151
R21302 vdd.n2484 vdd.n2481 10.6151
R21303 vdd.n2481 vdd.n2480 10.6151
R21304 vdd.n2480 vdd.n2477 10.6151
R21305 vdd.n2477 vdd.n2476 10.6151
R21306 vdd.n2476 vdd.n2473 10.6151
R21307 vdd.n2473 vdd.n2472 10.6151
R21308 vdd.n2472 vdd.n2469 10.6151
R21309 vdd.n2469 vdd.n2468 10.6151
R21310 vdd.n2465 vdd.n2464 10.6151
R21311 vdd.n2464 vdd.n2462 10.6151
R21312 vdd.n2221 vdd.n2219 10.6151
R21313 vdd.n2222 vdd.n2221 10.6151
R21314 vdd.n2224 vdd.n2222 10.6151
R21315 vdd.n2225 vdd.n2224 10.6151
R21316 vdd.n2227 vdd.n2225 10.6151
R21317 vdd.n2228 vdd.n2227 10.6151
R21318 vdd.n2230 vdd.n2228 10.6151
R21319 vdd.n2231 vdd.n2230 10.6151
R21320 vdd.n2233 vdd.n2231 10.6151
R21321 vdd.n2234 vdd.n2233 10.6151
R21322 vdd.n2236 vdd.n2234 10.6151
R21323 vdd.n2237 vdd.n2236 10.6151
R21324 vdd.n2255 vdd.n2237 10.6151
R21325 vdd.n2255 vdd.n2254 10.6151
R21326 vdd.n2254 vdd.n2253 10.6151
R21327 vdd.n2253 vdd.n2251 10.6151
R21328 vdd.n2251 vdd.n2250 10.6151
R21329 vdd.n2250 vdd.n2248 10.6151
R21330 vdd.n2248 vdd.n2247 10.6151
R21331 vdd.n2247 vdd.n2245 10.6151
R21332 vdd.n2245 vdd.n2244 10.6151
R21333 vdd.n2244 vdd.n2242 10.6151
R21334 vdd.n2242 vdd.n2241 10.6151
R21335 vdd.n2241 vdd.n2239 10.6151
R21336 vdd.n2239 vdd.n2238 10.6151
R21337 vdd.n2238 vdd.n968 10.6151
R21338 vdd.n2460 vdd.n968 10.6151
R21339 vdd.n2461 vdd.n2460 10.6151
R21340 vdd.n2372 vdd.n2371 10.6151
R21341 vdd.n2371 vdd.n1053 10.6151
R21342 vdd.n2365 vdd.n1053 10.6151
R21343 vdd.n2365 vdd.n2364 10.6151
R21344 vdd.n2364 vdd.n2363 10.6151
R21345 vdd.n2363 vdd.n1055 10.6151
R21346 vdd.n2357 vdd.n1055 10.6151
R21347 vdd.n2357 vdd.n2356 10.6151
R21348 vdd.n2356 vdd.n2355 10.6151
R21349 vdd.n2355 vdd.n1057 10.6151
R21350 vdd.n2349 vdd.n1057 10.6151
R21351 vdd.n2349 vdd.n2348 10.6151
R21352 vdd.n2348 vdd.n2347 10.6151
R21353 vdd.n2347 vdd.n1059 10.6151
R21354 vdd.n2341 vdd.n1059 10.6151
R21355 vdd.n2341 vdd.n2340 10.6151
R21356 vdd.n2340 vdd.n2339 10.6151
R21357 vdd.n2339 vdd.n1063 10.6151
R21358 vdd.n2187 vdd.n1063 10.6151
R21359 vdd.n2188 vdd.n2187 10.6151
R21360 vdd.n2188 vdd.n2183 10.6151
R21361 vdd.n2194 vdd.n2183 10.6151
R21362 vdd.n2195 vdd.n2194 10.6151
R21363 vdd.n2196 vdd.n2195 10.6151
R21364 vdd.n2196 vdd.n2181 10.6151
R21365 vdd.n2202 vdd.n2181 10.6151
R21366 vdd.n2203 vdd.n2202 10.6151
R21367 vdd.n2204 vdd.n2203 10.6151
R21368 vdd.n2204 vdd.n2179 10.6151
R21369 vdd.n2210 vdd.n2179 10.6151
R21370 vdd.n2211 vdd.n2210 10.6151
R21371 vdd.n2213 vdd.n2175 10.6151
R21372 vdd.n2218 vdd.n2175 10.6151
R21373 vdd.n1851 vdd.t41 10.5435
R21374 vdd.n656 vdd.t85 10.5435
R21375 vdd.n316 vdd.n298 10.4732
R21376 vdd.n257 vdd.n239 10.4732
R21377 vdd.n214 vdd.n196 10.4732
R21378 vdd.n155 vdd.n137 10.4732
R21379 vdd.n113 vdd.n95 10.4732
R21380 vdd.n54 vdd.n36 10.4732
R21381 vdd.n1735 vdd.n1717 10.4732
R21382 vdd.n1794 vdd.n1776 10.4732
R21383 vdd.n1633 vdd.n1615 10.4732
R21384 vdd.n1692 vdd.n1674 10.4732
R21385 vdd.n1532 vdd.n1514 10.4732
R21386 vdd.n1591 vdd.n1573 10.4732
R21387 vdd.t10 vdd.n1825 10.3167
R21388 vdd.n3300 vdd.t67 10.3167
R21389 vdd.n1502 vdd.t4 10.09
R21390 vdd.n3394 vdd.t0 10.09
R21391 vdd.t52 vdd.n1155 9.86327
R21392 vdd.n3385 vdd.t265 9.86327
R21393 vdd.n315 vdd.n300 9.69747
R21394 vdd.n256 vdd.n241 9.69747
R21395 vdd.n213 vdd.n198 9.69747
R21396 vdd.n154 vdd.n139 9.69747
R21397 vdd.n112 vdd.n97 9.69747
R21398 vdd.n53 vdd.n38 9.69747
R21399 vdd.n1734 vdd.n1719 9.69747
R21400 vdd.n1793 vdd.n1778 9.69747
R21401 vdd.n1632 vdd.n1617 9.69747
R21402 vdd.n1691 vdd.n1676 9.69747
R21403 vdd.n1531 vdd.n1516 9.69747
R21404 vdd.n1590 vdd.n1575 9.69747
R21405 vdd.n2315 vdd.n2314 9.67831
R21406 vdd.n3216 vdd.n731 9.67831
R21407 vdd.n3093 vdd.n3092 9.67831
R21408 vdd.n2339 vdd.n2338 9.67831
R21409 vdd.n1461 vdd.t28 9.63654
R21410 vdd.n3331 vdd.t60 9.63654
R21411 vdd.n331 vdd.n330 9.45567
R21412 vdd.n272 vdd.n271 9.45567
R21413 vdd.n229 vdd.n228 9.45567
R21414 vdd.n170 vdd.n169 9.45567
R21415 vdd.n128 vdd.n127 9.45567
R21416 vdd.n69 vdd.n68 9.45567
R21417 vdd.n1750 vdd.n1749 9.45567
R21418 vdd.n1809 vdd.n1808 9.45567
R21419 vdd.n1648 vdd.n1647 9.45567
R21420 vdd.n1707 vdd.n1706 9.45567
R21421 vdd.n1547 vdd.n1546 9.45567
R21422 vdd.n1606 vdd.n1605 9.45567
R21423 vdd.n1435 vdd.t58 9.40981
R21424 vdd.n3363 vdd.t111 9.40981
R21425 vdd.n2075 vdd.n1929 9.3005
R21426 vdd.n2074 vdd.n2073 9.3005
R21427 vdd.n1935 vdd.n1934 9.3005
R21428 vdd.n2068 vdd.n1939 9.3005
R21429 vdd.n2067 vdd.n1940 9.3005
R21430 vdd.n2066 vdd.n1941 9.3005
R21431 vdd.n1945 vdd.n1942 9.3005
R21432 vdd.n2061 vdd.n1946 9.3005
R21433 vdd.n2060 vdd.n1947 9.3005
R21434 vdd.n2059 vdd.n1948 9.3005
R21435 vdd.n1952 vdd.n1949 9.3005
R21436 vdd.n2054 vdd.n1953 9.3005
R21437 vdd.n2053 vdd.n1954 9.3005
R21438 vdd.n2052 vdd.n1955 9.3005
R21439 vdd.n1959 vdd.n1956 9.3005
R21440 vdd.n2047 vdd.n1960 9.3005
R21441 vdd.n2046 vdd.n1961 9.3005
R21442 vdd.n2045 vdd.n1962 9.3005
R21443 vdd.n1966 vdd.n1963 9.3005
R21444 vdd.n2040 vdd.n1967 9.3005
R21445 vdd.n2039 vdd.n1968 9.3005
R21446 vdd.n2038 vdd.n2037 9.3005
R21447 vdd.n2036 vdd.n1969 9.3005
R21448 vdd.n2035 vdd.n2034 9.3005
R21449 vdd.n1975 vdd.n1974 9.3005
R21450 vdd.n2029 vdd.n1979 9.3005
R21451 vdd.n2028 vdd.n1980 9.3005
R21452 vdd.n2027 vdd.n1981 9.3005
R21453 vdd.n1985 vdd.n1982 9.3005
R21454 vdd.n2022 vdd.n1986 9.3005
R21455 vdd.n2021 vdd.n1987 9.3005
R21456 vdd.n2020 vdd.n1988 9.3005
R21457 vdd.n1992 vdd.n1989 9.3005
R21458 vdd.n2015 vdd.n1993 9.3005
R21459 vdd.n2014 vdd.n1994 9.3005
R21460 vdd.n2013 vdd.n1995 9.3005
R21461 vdd.n1997 vdd.n1996 9.3005
R21462 vdd.n2008 vdd.n1064 9.3005
R21463 vdd.n2077 vdd.n2076 9.3005
R21464 vdd.n2101 vdd.n2100 9.3005
R21465 vdd.n1907 vdd.n1906 9.3005
R21466 vdd.n1912 vdd.n1910 9.3005
R21467 vdd.n2093 vdd.n1913 9.3005
R21468 vdd.n2092 vdd.n1914 9.3005
R21469 vdd.n2091 vdd.n1915 9.3005
R21470 vdd.n1919 vdd.n1916 9.3005
R21471 vdd.n2086 vdd.n1920 9.3005
R21472 vdd.n2085 vdd.n1921 9.3005
R21473 vdd.n2084 vdd.n1922 9.3005
R21474 vdd.n1926 vdd.n1923 9.3005
R21475 vdd.n2079 vdd.n1927 9.3005
R21476 vdd.n2078 vdd.n1928 9.3005
R21477 vdd.n2323 vdd.n1900 9.3005
R21478 vdd.n2325 vdd.n2324 9.3005
R21479 vdd.n1815 vdd.n1814 9.3005
R21480 vdd.n1124 vdd.n1123 9.3005
R21481 vdd.n1829 vdd.n1828 9.3005
R21482 vdd.n1830 vdd.n1122 9.3005
R21483 vdd.n1832 vdd.n1831 9.3005
R21484 vdd.n1113 vdd.n1112 9.3005
R21485 vdd.n1846 vdd.n1845 9.3005
R21486 vdd.n1847 vdd.n1111 9.3005
R21487 vdd.n1849 vdd.n1848 9.3005
R21488 vdd.n1102 vdd.n1101 9.3005
R21489 vdd.n1862 vdd.n1861 9.3005
R21490 vdd.n1863 vdd.n1100 9.3005
R21491 vdd.n1865 vdd.n1864 9.3005
R21492 vdd.n1090 vdd.n1089 9.3005
R21493 vdd.n1879 vdd.n1878 9.3005
R21494 vdd.n1880 vdd.n1088 9.3005
R21495 vdd.n1882 vdd.n1881 9.3005
R21496 vdd.n1078 vdd.n1077 9.3005
R21497 vdd.n1898 vdd.n1897 9.3005
R21498 vdd.n1899 vdd.n1076 9.3005
R21499 vdd.n2327 vdd.n2326 9.3005
R21500 vdd.n307 vdd.n306 9.3005
R21501 vdd.n302 vdd.n301 9.3005
R21502 vdd.n313 vdd.n312 9.3005
R21503 vdd.n315 vdd.n314 9.3005
R21504 vdd.n298 vdd.n297 9.3005
R21505 vdd.n321 vdd.n320 9.3005
R21506 vdd.n323 vdd.n322 9.3005
R21507 vdd.n295 vdd.n292 9.3005
R21508 vdd.n330 vdd.n329 9.3005
R21509 vdd.n248 vdd.n247 9.3005
R21510 vdd.n243 vdd.n242 9.3005
R21511 vdd.n254 vdd.n253 9.3005
R21512 vdd.n256 vdd.n255 9.3005
R21513 vdd.n239 vdd.n238 9.3005
R21514 vdd.n262 vdd.n261 9.3005
R21515 vdd.n264 vdd.n263 9.3005
R21516 vdd.n236 vdd.n233 9.3005
R21517 vdd.n271 vdd.n270 9.3005
R21518 vdd.n205 vdd.n204 9.3005
R21519 vdd.n200 vdd.n199 9.3005
R21520 vdd.n211 vdd.n210 9.3005
R21521 vdd.n213 vdd.n212 9.3005
R21522 vdd.n196 vdd.n195 9.3005
R21523 vdd.n219 vdd.n218 9.3005
R21524 vdd.n221 vdd.n220 9.3005
R21525 vdd.n193 vdd.n190 9.3005
R21526 vdd.n228 vdd.n227 9.3005
R21527 vdd.n146 vdd.n145 9.3005
R21528 vdd.n141 vdd.n140 9.3005
R21529 vdd.n152 vdd.n151 9.3005
R21530 vdd.n154 vdd.n153 9.3005
R21531 vdd.n137 vdd.n136 9.3005
R21532 vdd.n160 vdd.n159 9.3005
R21533 vdd.n162 vdd.n161 9.3005
R21534 vdd.n134 vdd.n131 9.3005
R21535 vdd.n169 vdd.n168 9.3005
R21536 vdd.n104 vdd.n103 9.3005
R21537 vdd.n99 vdd.n98 9.3005
R21538 vdd.n110 vdd.n109 9.3005
R21539 vdd.n112 vdd.n111 9.3005
R21540 vdd.n95 vdd.n94 9.3005
R21541 vdd.n118 vdd.n117 9.3005
R21542 vdd.n120 vdd.n119 9.3005
R21543 vdd.n92 vdd.n89 9.3005
R21544 vdd.n127 vdd.n126 9.3005
R21545 vdd.n45 vdd.n44 9.3005
R21546 vdd.n40 vdd.n39 9.3005
R21547 vdd.n51 vdd.n50 9.3005
R21548 vdd.n53 vdd.n52 9.3005
R21549 vdd.n36 vdd.n35 9.3005
R21550 vdd.n59 vdd.n58 9.3005
R21551 vdd.n61 vdd.n60 9.3005
R21552 vdd.n33 vdd.n30 9.3005
R21553 vdd.n68 vdd.n67 9.3005
R21554 vdd.n3138 vdd.n3137 9.3005
R21555 vdd.n3141 vdd.n766 9.3005
R21556 vdd.n3142 vdd.n765 9.3005
R21557 vdd.n3145 vdd.n764 9.3005
R21558 vdd.n3146 vdd.n763 9.3005
R21559 vdd.n3149 vdd.n762 9.3005
R21560 vdd.n3150 vdd.n761 9.3005
R21561 vdd.n3153 vdd.n760 9.3005
R21562 vdd.n3154 vdd.n759 9.3005
R21563 vdd.n3157 vdd.n758 9.3005
R21564 vdd.n3158 vdd.n757 9.3005
R21565 vdd.n3161 vdd.n756 9.3005
R21566 vdd.n3162 vdd.n755 9.3005
R21567 vdd.n3165 vdd.n754 9.3005
R21568 vdd.n3166 vdd.n753 9.3005
R21569 vdd.n3169 vdd.n752 9.3005
R21570 vdd.n3170 vdd.n751 9.3005
R21571 vdd.n3173 vdd.n750 9.3005
R21572 vdd.n3174 vdd.n749 9.3005
R21573 vdd.n3177 vdd.n748 9.3005
R21574 vdd.n3181 vdd.n3180 9.3005
R21575 vdd.n3182 vdd.n747 9.3005
R21576 vdd.n3186 vdd.n3183 9.3005
R21577 vdd.n3189 vdd.n746 9.3005
R21578 vdd.n3190 vdd.n745 9.3005
R21579 vdd.n3193 vdd.n744 9.3005
R21580 vdd.n3194 vdd.n743 9.3005
R21581 vdd.n3197 vdd.n742 9.3005
R21582 vdd.n3198 vdd.n741 9.3005
R21583 vdd.n3201 vdd.n740 9.3005
R21584 vdd.n3202 vdd.n739 9.3005
R21585 vdd.n3205 vdd.n738 9.3005
R21586 vdd.n3206 vdd.n737 9.3005
R21587 vdd.n3209 vdd.n736 9.3005
R21588 vdd.n3210 vdd.n735 9.3005
R21589 vdd.n3213 vdd.n730 9.3005
R21590 vdd.n3219 vdd.n727 9.3005
R21591 vdd.n3220 vdd.n726 9.3005
R21592 vdd.n3234 vdd.n3233 9.3005
R21593 vdd.n3235 vdd.n681 9.3005
R21594 vdd.n3237 vdd.n3236 9.3005
R21595 vdd.n671 vdd.n670 9.3005
R21596 vdd.n3251 vdd.n3250 9.3005
R21597 vdd.n3252 vdd.n669 9.3005
R21598 vdd.n3254 vdd.n3253 9.3005
R21599 vdd.n660 vdd.n659 9.3005
R21600 vdd.n3267 vdd.n3266 9.3005
R21601 vdd.n3268 vdd.n658 9.3005
R21602 vdd.n3270 vdd.n3269 9.3005
R21603 vdd.n648 vdd.n647 9.3005
R21604 vdd.n3284 vdd.n3283 9.3005
R21605 vdd.n3285 vdd.n646 9.3005
R21606 vdd.n3287 vdd.n3286 9.3005
R21607 vdd.n637 vdd.n636 9.3005
R21608 vdd.n3303 vdd.n3302 9.3005
R21609 vdd.n3304 vdd.n635 9.3005
R21610 vdd.n3306 vdd.n3305 9.3005
R21611 vdd.n336 vdd.n334 9.3005
R21612 vdd.n683 vdd.n682 9.3005
R21613 vdd.n3398 vdd.n3397 9.3005
R21614 vdd.n337 vdd.n335 9.3005
R21615 vdd.n3391 vdd.n346 9.3005
R21616 vdd.n3390 vdd.n347 9.3005
R21617 vdd.n3389 vdd.n348 9.3005
R21618 vdd.n355 vdd.n349 9.3005
R21619 vdd.n3383 vdd.n356 9.3005
R21620 vdd.n3382 vdd.n357 9.3005
R21621 vdd.n3381 vdd.n358 9.3005
R21622 vdd.n366 vdd.n359 9.3005
R21623 vdd.n3375 vdd.n367 9.3005
R21624 vdd.n3374 vdd.n368 9.3005
R21625 vdd.n3373 vdd.n369 9.3005
R21626 vdd.n377 vdd.n370 9.3005
R21627 vdd.n3367 vdd.n378 9.3005
R21628 vdd.n3366 vdd.n379 9.3005
R21629 vdd.n3365 vdd.n380 9.3005
R21630 vdd.n388 vdd.n381 9.3005
R21631 vdd.n3359 vdd.n389 9.3005
R21632 vdd.n3358 vdd.n390 9.3005
R21633 vdd.n3357 vdd.n391 9.3005
R21634 vdd.n466 vdd.n463 9.3005
R21635 vdd.n470 vdd.n469 9.3005
R21636 vdd.n471 vdd.n462 9.3005
R21637 vdd.n475 vdd.n472 9.3005
R21638 vdd.n476 vdd.n461 9.3005
R21639 vdd.n480 vdd.n479 9.3005
R21640 vdd.n481 vdd.n460 9.3005
R21641 vdd.n485 vdd.n482 9.3005
R21642 vdd.n486 vdd.n459 9.3005
R21643 vdd.n490 vdd.n489 9.3005
R21644 vdd.n491 vdd.n458 9.3005
R21645 vdd.n495 vdd.n492 9.3005
R21646 vdd.n496 vdd.n457 9.3005
R21647 vdd.n500 vdd.n499 9.3005
R21648 vdd.n501 vdd.n456 9.3005
R21649 vdd.n505 vdd.n502 9.3005
R21650 vdd.n506 vdd.n455 9.3005
R21651 vdd.n510 vdd.n509 9.3005
R21652 vdd.n511 vdd.n454 9.3005
R21653 vdd.n515 vdd.n512 9.3005
R21654 vdd.n516 vdd.n451 9.3005
R21655 vdd.n520 vdd.n519 9.3005
R21656 vdd.n521 vdd.n450 9.3005
R21657 vdd.n525 vdd.n522 9.3005
R21658 vdd.n526 vdd.n449 9.3005
R21659 vdd.n530 vdd.n529 9.3005
R21660 vdd.n531 vdd.n448 9.3005
R21661 vdd.n535 vdd.n532 9.3005
R21662 vdd.n536 vdd.n447 9.3005
R21663 vdd.n540 vdd.n539 9.3005
R21664 vdd.n541 vdd.n446 9.3005
R21665 vdd.n545 vdd.n542 9.3005
R21666 vdd.n546 vdd.n445 9.3005
R21667 vdd.n550 vdd.n549 9.3005
R21668 vdd.n551 vdd.n444 9.3005
R21669 vdd.n555 vdd.n552 9.3005
R21670 vdd.n556 vdd.n443 9.3005
R21671 vdd.n560 vdd.n559 9.3005
R21672 vdd.n561 vdd.n442 9.3005
R21673 vdd.n565 vdd.n562 9.3005
R21674 vdd.n566 vdd.n439 9.3005
R21675 vdd.n570 vdd.n569 9.3005
R21676 vdd.n571 vdd.n438 9.3005
R21677 vdd.n575 vdd.n572 9.3005
R21678 vdd.n576 vdd.n437 9.3005
R21679 vdd.n580 vdd.n579 9.3005
R21680 vdd.n581 vdd.n436 9.3005
R21681 vdd.n585 vdd.n582 9.3005
R21682 vdd.n586 vdd.n435 9.3005
R21683 vdd.n590 vdd.n589 9.3005
R21684 vdd.n591 vdd.n434 9.3005
R21685 vdd.n595 vdd.n592 9.3005
R21686 vdd.n596 vdd.n433 9.3005
R21687 vdd.n600 vdd.n599 9.3005
R21688 vdd.n601 vdd.n432 9.3005
R21689 vdd.n605 vdd.n602 9.3005
R21690 vdd.n606 vdd.n431 9.3005
R21691 vdd.n610 vdd.n609 9.3005
R21692 vdd.n611 vdd.n430 9.3005
R21693 vdd.n615 vdd.n612 9.3005
R21694 vdd.n617 vdd.n429 9.3005
R21695 vdd.n619 vdd.n618 9.3005
R21696 vdd.n3351 vdd.n3350 9.3005
R21697 vdd.n465 vdd.n464 9.3005
R21698 vdd.n3229 vdd.n3228 9.3005
R21699 vdd.n676 vdd.n675 9.3005
R21700 vdd.n3242 vdd.n3241 9.3005
R21701 vdd.n3243 vdd.n674 9.3005
R21702 vdd.n3245 vdd.n3244 9.3005
R21703 vdd.n666 vdd.n665 9.3005
R21704 vdd.n3259 vdd.n3258 9.3005
R21705 vdd.n3260 vdd.n664 9.3005
R21706 vdd.n3262 vdd.n3261 9.3005
R21707 vdd.n653 vdd.n652 9.3005
R21708 vdd.n3275 vdd.n3274 9.3005
R21709 vdd.n3276 vdd.n651 9.3005
R21710 vdd.n3278 vdd.n3277 9.3005
R21711 vdd.n642 vdd.n641 9.3005
R21712 vdd.n3292 vdd.n3291 9.3005
R21713 vdd.n3293 vdd.n640 9.3005
R21714 vdd.n3298 vdd.n3294 9.3005
R21715 vdd.n3297 vdd.n3296 9.3005
R21716 vdd.n3295 vdd.n631 9.3005
R21717 vdd.n3311 vdd.n630 9.3005
R21718 vdd.n3313 vdd.n3312 9.3005
R21719 vdd.n3314 vdd.n629 9.3005
R21720 vdd.n3316 vdd.n3315 9.3005
R21721 vdd.n3318 vdd.n628 9.3005
R21722 vdd.n3320 vdd.n3319 9.3005
R21723 vdd.n3321 vdd.n627 9.3005
R21724 vdd.n3323 vdd.n3322 9.3005
R21725 vdd.n3325 vdd.n626 9.3005
R21726 vdd.n3327 vdd.n3326 9.3005
R21727 vdd.n3328 vdd.n625 9.3005
R21728 vdd.n3330 vdd.n3329 9.3005
R21729 vdd.n3333 vdd.n624 9.3005
R21730 vdd.n3335 vdd.n3334 9.3005
R21731 vdd.n3336 vdd.n623 9.3005
R21732 vdd.n3338 vdd.n3337 9.3005
R21733 vdd.n3340 vdd.n622 9.3005
R21734 vdd.n3342 vdd.n3341 9.3005
R21735 vdd.n3343 vdd.n621 9.3005
R21736 vdd.n3345 vdd.n3344 9.3005
R21737 vdd.n3347 vdd.n620 9.3005
R21738 vdd.n3349 vdd.n3348 9.3005
R21739 vdd.n3227 vdd.n686 9.3005
R21740 vdd.n3226 vdd.n3225 9.3005
R21741 vdd.n3095 vdd.n687 9.3005
R21742 vdd.n3104 vdd.n783 9.3005
R21743 vdd.n3107 vdd.n782 9.3005
R21744 vdd.n3108 vdd.n781 9.3005
R21745 vdd.n3111 vdd.n780 9.3005
R21746 vdd.n3112 vdd.n779 9.3005
R21747 vdd.n3115 vdd.n778 9.3005
R21748 vdd.n3116 vdd.n777 9.3005
R21749 vdd.n3119 vdd.n776 9.3005
R21750 vdd.n3120 vdd.n775 9.3005
R21751 vdd.n3123 vdd.n774 9.3005
R21752 vdd.n3124 vdd.n773 9.3005
R21753 vdd.n3127 vdd.n772 9.3005
R21754 vdd.n3128 vdd.n771 9.3005
R21755 vdd.n3131 vdd.n770 9.3005
R21756 vdd.n3135 vdd.n3134 9.3005
R21757 vdd.n3136 vdd.n767 9.3005
R21758 vdd.n2337 vdd.n2336 9.3005
R21759 vdd.n2332 vdd.n1067 9.3005
R21760 vdd.n1430 vdd.n1429 9.3005
R21761 vdd.n1431 vdd.n1185 9.3005
R21762 vdd.n1433 vdd.n1432 9.3005
R21763 vdd.n1175 vdd.n1174 9.3005
R21764 vdd.n1447 vdd.n1446 9.3005
R21765 vdd.n1448 vdd.n1173 9.3005
R21766 vdd.n1450 vdd.n1449 9.3005
R21767 vdd.n1165 vdd.n1164 9.3005
R21768 vdd.n1464 vdd.n1463 9.3005
R21769 vdd.n1465 vdd.n1163 9.3005
R21770 vdd.n1467 vdd.n1466 9.3005
R21771 vdd.n1152 vdd.n1151 9.3005
R21772 vdd.n1480 vdd.n1479 9.3005
R21773 vdd.n1481 vdd.n1150 9.3005
R21774 vdd.n1483 vdd.n1482 9.3005
R21775 vdd.n1141 vdd.n1140 9.3005
R21776 vdd.n1497 vdd.n1496 9.3005
R21777 vdd.n1498 vdd.n1139 9.3005
R21778 vdd.n1500 vdd.n1499 9.3005
R21779 vdd.n1130 vdd.n1129 9.3005
R21780 vdd.n1820 vdd.n1819 9.3005
R21781 vdd.n1821 vdd.n1128 9.3005
R21782 vdd.n1823 vdd.n1822 9.3005
R21783 vdd.n1118 vdd.n1117 9.3005
R21784 vdd.n1837 vdd.n1836 9.3005
R21785 vdd.n1838 vdd.n1116 9.3005
R21786 vdd.n1840 vdd.n1839 9.3005
R21787 vdd.n1108 vdd.n1107 9.3005
R21788 vdd.n1854 vdd.n1853 9.3005
R21789 vdd.n1855 vdd.n1106 9.3005
R21790 vdd.n1857 vdd.n1856 9.3005
R21791 vdd.n1095 vdd.n1094 9.3005
R21792 vdd.n1870 vdd.n1869 9.3005
R21793 vdd.n1871 vdd.n1093 9.3005
R21794 vdd.n1873 vdd.n1872 9.3005
R21795 vdd.n1085 vdd.n1084 9.3005
R21796 vdd.n1887 vdd.n1886 9.3005
R21797 vdd.n1888 vdd.n1082 9.3005
R21798 vdd.n1892 vdd.n1891 9.3005
R21799 vdd.n1890 vdd.n1083 9.3005
R21800 vdd.n1889 vdd.n1072 9.3005
R21801 vdd.n1187 vdd.n1186 9.3005
R21802 vdd.n1323 vdd.n1322 9.3005
R21803 vdd.n1324 vdd.n1313 9.3005
R21804 vdd.n1326 vdd.n1325 9.3005
R21805 vdd.n1327 vdd.n1312 9.3005
R21806 vdd.n1329 vdd.n1328 9.3005
R21807 vdd.n1330 vdd.n1307 9.3005
R21808 vdd.n1332 vdd.n1331 9.3005
R21809 vdd.n1333 vdd.n1306 9.3005
R21810 vdd.n1335 vdd.n1334 9.3005
R21811 vdd.n1336 vdd.n1301 9.3005
R21812 vdd.n1338 vdd.n1337 9.3005
R21813 vdd.n1339 vdd.n1300 9.3005
R21814 vdd.n1341 vdd.n1340 9.3005
R21815 vdd.n1342 vdd.n1295 9.3005
R21816 vdd.n1344 vdd.n1343 9.3005
R21817 vdd.n1345 vdd.n1294 9.3005
R21818 vdd.n1347 vdd.n1346 9.3005
R21819 vdd.n1348 vdd.n1289 9.3005
R21820 vdd.n1350 vdd.n1349 9.3005
R21821 vdd.n1351 vdd.n1288 9.3005
R21822 vdd.n1353 vdd.n1352 9.3005
R21823 vdd.n1357 vdd.n1284 9.3005
R21824 vdd.n1359 vdd.n1358 9.3005
R21825 vdd.n1360 vdd.n1283 9.3005
R21826 vdd.n1362 vdd.n1361 9.3005
R21827 vdd.n1363 vdd.n1278 9.3005
R21828 vdd.n1365 vdd.n1364 9.3005
R21829 vdd.n1366 vdd.n1277 9.3005
R21830 vdd.n1368 vdd.n1367 9.3005
R21831 vdd.n1369 vdd.n1272 9.3005
R21832 vdd.n1371 vdd.n1370 9.3005
R21833 vdd.n1372 vdd.n1271 9.3005
R21834 vdd.n1374 vdd.n1373 9.3005
R21835 vdd.n1375 vdd.n1266 9.3005
R21836 vdd.n1377 vdd.n1376 9.3005
R21837 vdd.n1378 vdd.n1265 9.3005
R21838 vdd.n1380 vdd.n1379 9.3005
R21839 vdd.n1381 vdd.n1260 9.3005
R21840 vdd.n1383 vdd.n1382 9.3005
R21841 vdd.n1384 vdd.n1259 9.3005
R21842 vdd.n1386 vdd.n1385 9.3005
R21843 vdd.n1387 vdd.n1254 9.3005
R21844 vdd.n1389 vdd.n1388 9.3005
R21845 vdd.n1390 vdd.n1253 9.3005
R21846 vdd.n1392 vdd.n1391 9.3005
R21847 vdd.n1393 vdd.n1246 9.3005
R21848 vdd.n1395 vdd.n1394 9.3005
R21849 vdd.n1396 vdd.n1245 9.3005
R21850 vdd.n1398 vdd.n1397 9.3005
R21851 vdd.n1399 vdd.n1240 9.3005
R21852 vdd.n1401 vdd.n1400 9.3005
R21853 vdd.n1402 vdd.n1239 9.3005
R21854 vdd.n1404 vdd.n1403 9.3005
R21855 vdd.n1405 vdd.n1234 9.3005
R21856 vdd.n1407 vdd.n1406 9.3005
R21857 vdd.n1408 vdd.n1233 9.3005
R21858 vdd.n1410 vdd.n1409 9.3005
R21859 vdd.n1411 vdd.n1228 9.3005
R21860 vdd.n1413 vdd.n1412 9.3005
R21861 vdd.n1414 vdd.n1227 9.3005
R21862 vdd.n1416 vdd.n1415 9.3005
R21863 vdd.n1192 vdd.n1191 9.3005
R21864 vdd.n1422 vdd.n1421 9.3005
R21865 vdd.n1321 vdd.n1320 9.3005
R21866 vdd.n1425 vdd.n1424 9.3005
R21867 vdd.n1181 vdd.n1180 9.3005
R21868 vdd.n1439 vdd.n1438 9.3005
R21869 vdd.n1440 vdd.n1179 9.3005
R21870 vdd.n1442 vdd.n1441 9.3005
R21871 vdd.n1170 vdd.n1169 9.3005
R21872 vdd.n1456 vdd.n1455 9.3005
R21873 vdd.n1457 vdd.n1168 9.3005
R21874 vdd.n1459 vdd.n1458 9.3005
R21875 vdd.n1159 vdd.n1158 9.3005
R21876 vdd.n1472 vdd.n1471 9.3005
R21877 vdd.n1473 vdd.n1157 9.3005
R21878 vdd.n1475 vdd.n1474 9.3005
R21879 vdd.n1147 vdd.n1146 9.3005
R21880 vdd.n1489 vdd.n1488 9.3005
R21881 vdd.n1490 vdd.n1145 9.3005
R21882 vdd.n1492 vdd.n1491 9.3005
R21883 vdd.n1136 vdd.n1135 9.3005
R21884 vdd.n1505 vdd.n1504 9.3005
R21885 vdd.n1506 vdd.n1134 9.3005
R21886 vdd.n1423 vdd.n1190 9.3005
R21887 vdd.n1726 vdd.n1725 9.3005
R21888 vdd.n1721 vdd.n1720 9.3005
R21889 vdd.n1732 vdd.n1731 9.3005
R21890 vdd.n1734 vdd.n1733 9.3005
R21891 vdd.n1717 vdd.n1716 9.3005
R21892 vdd.n1740 vdd.n1739 9.3005
R21893 vdd.n1742 vdd.n1741 9.3005
R21894 vdd.n1714 vdd.n1711 9.3005
R21895 vdd.n1749 vdd.n1748 9.3005
R21896 vdd.n1785 vdd.n1784 9.3005
R21897 vdd.n1780 vdd.n1779 9.3005
R21898 vdd.n1791 vdd.n1790 9.3005
R21899 vdd.n1793 vdd.n1792 9.3005
R21900 vdd.n1776 vdd.n1775 9.3005
R21901 vdd.n1799 vdd.n1798 9.3005
R21902 vdd.n1801 vdd.n1800 9.3005
R21903 vdd.n1773 vdd.n1770 9.3005
R21904 vdd.n1808 vdd.n1807 9.3005
R21905 vdd.n1624 vdd.n1623 9.3005
R21906 vdd.n1619 vdd.n1618 9.3005
R21907 vdd.n1630 vdd.n1629 9.3005
R21908 vdd.n1632 vdd.n1631 9.3005
R21909 vdd.n1615 vdd.n1614 9.3005
R21910 vdd.n1638 vdd.n1637 9.3005
R21911 vdd.n1640 vdd.n1639 9.3005
R21912 vdd.n1612 vdd.n1609 9.3005
R21913 vdd.n1647 vdd.n1646 9.3005
R21914 vdd.n1683 vdd.n1682 9.3005
R21915 vdd.n1678 vdd.n1677 9.3005
R21916 vdd.n1689 vdd.n1688 9.3005
R21917 vdd.n1691 vdd.n1690 9.3005
R21918 vdd.n1674 vdd.n1673 9.3005
R21919 vdd.n1697 vdd.n1696 9.3005
R21920 vdd.n1699 vdd.n1698 9.3005
R21921 vdd.n1671 vdd.n1668 9.3005
R21922 vdd.n1706 vdd.n1705 9.3005
R21923 vdd.n1523 vdd.n1522 9.3005
R21924 vdd.n1518 vdd.n1517 9.3005
R21925 vdd.n1529 vdd.n1528 9.3005
R21926 vdd.n1531 vdd.n1530 9.3005
R21927 vdd.n1514 vdd.n1513 9.3005
R21928 vdd.n1537 vdd.n1536 9.3005
R21929 vdd.n1539 vdd.n1538 9.3005
R21930 vdd.n1511 vdd.n1508 9.3005
R21931 vdd.n1546 vdd.n1545 9.3005
R21932 vdd.n1582 vdd.n1581 9.3005
R21933 vdd.n1577 vdd.n1576 9.3005
R21934 vdd.n1588 vdd.n1587 9.3005
R21935 vdd.n1590 vdd.n1589 9.3005
R21936 vdd.n1573 vdd.n1572 9.3005
R21937 vdd.n1596 vdd.n1595 9.3005
R21938 vdd.n1598 vdd.n1597 9.3005
R21939 vdd.n1570 vdd.n1567 9.3005
R21940 vdd.n1605 vdd.n1604 9.3005
R21941 vdd.n1461 vdd.t78 9.18308
R21942 vdd.n3331 vdd.t80 9.18308
R21943 vdd.n1155 vdd.t119 8.95635
R21944 vdd.n2329 vdd.t177 8.95635
R21945 vdd.n723 vdd.t170 8.95635
R21946 vdd.t90 vdd.n3385 8.95635
R21947 vdd.n312 vdd.n311 8.92171
R21948 vdd.n253 vdd.n252 8.92171
R21949 vdd.n210 vdd.n209 8.92171
R21950 vdd.n151 vdd.n150 8.92171
R21951 vdd.n109 vdd.n108 8.92171
R21952 vdd.n50 vdd.n49 8.92171
R21953 vdd.n1731 vdd.n1730 8.92171
R21954 vdd.n1790 vdd.n1789 8.92171
R21955 vdd.n1629 vdd.n1628 8.92171
R21956 vdd.n1688 vdd.n1687 8.92171
R21957 vdd.n1528 vdd.n1527 8.92171
R21958 vdd.n1587 vdd.n1586 8.92171
R21959 vdd.n231 vdd.n129 8.81535
R21960 vdd.n1709 vdd.n1607 8.81535
R21961 vdd.n1502 vdd.t6 8.72962
R21962 vdd.t2 vdd.n3394 8.72962
R21963 vdd.n1825 vdd.t34 8.50289
R21964 vdd.n3300 vdd.t73 8.50289
R21965 vdd.n28 vdd.n14 8.42249
R21966 vdd.n1851 vdd.t64 8.27616
R21967 vdd.t102 vdd.n656 8.27616
R21968 vdd.n3400 vdd.n3399 8.16225
R21969 vdd.n1813 vdd.n1812 8.16225
R21970 vdd.n308 vdd.n302 8.14595
R21971 vdd.n249 vdd.n243 8.14595
R21972 vdd.n206 vdd.n200 8.14595
R21973 vdd.n147 vdd.n141 8.14595
R21974 vdd.n105 vdd.n99 8.14595
R21975 vdd.n46 vdd.n40 8.14595
R21976 vdd.n1727 vdd.n1721 8.14595
R21977 vdd.n1786 vdd.n1780 8.14595
R21978 vdd.n1625 vdd.n1619 8.14595
R21979 vdd.n1684 vdd.n1678 8.14595
R21980 vdd.n1524 vdd.n1518 8.14595
R21981 vdd.n1583 vdd.n1577 8.14595
R21982 vdd.n2923 vdd.n849 8.11757
R21983 vdd.n2397 vdd.n2396 8.11757
R21984 vdd.n1098 vdd.t54 8.04943
R21985 vdd.n3256 vdd.t105 8.04943
R21986 vdd.n2375 vdd.n1043 7.70933
R21987 vdd.n2381 vdd.n1043 7.70933
R21988 vdd.n2387 vdd.n1037 7.70933
R21989 vdd.n2387 vdd.n1030 7.70933
R21990 vdd.n2393 vdd.n1030 7.70933
R21991 vdd.n2393 vdd.n1033 7.70933
R21992 vdd.n2400 vdd.n1018 7.70933
R21993 vdd.n2406 vdd.n1018 7.70933
R21994 vdd.n2412 vdd.n1012 7.70933
R21995 vdd.n2418 vdd.n1008 7.70933
R21996 vdd.n2424 vdd.n1002 7.70933
R21997 vdd.n2436 vdd.n989 7.70933
R21998 vdd.n2442 vdd.n983 7.70933
R21999 vdd.n2442 vdd.n976 7.70933
R22000 vdd.n2450 vdd.n976 7.70933
R22001 vdd.n2457 vdd.t159 7.70933
R22002 vdd.n2532 vdd.t159 7.70933
R22003 vdd.n2864 vdd.t147 7.70933
R22004 vdd.n2870 vdd.t147 7.70933
R22005 vdd.n2876 vdd.n897 7.70933
R22006 vdd.n2882 vdd.n897 7.70933
R22007 vdd.n2882 vdd.n900 7.70933
R22008 vdd.n2888 vdd.n893 7.70933
R22009 vdd.n2900 vdd.n880 7.70933
R22010 vdd.n2906 vdd.n874 7.70933
R22011 vdd.n2912 vdd.n870 7.70933
R22012 vdd.n2918 vdd.n857 7.70933
R22013 vdd.n2926 vdd.n857 7.70933
R22014 vdd.n2932 vdd.n851 7.70933
R22015 vdd.n2932 vdd.n843 7.70933
R22016 vdd.n2983 vdd.n843 7.70933
R22017 vdd.n2983 vdd.n846 7.70933
R22018 vdd.n2989 vdd.n805 7.70933
R22019 vdd.n3059 vdd.n805 7.70933
R22020 vdd.n307 vdd.n304 7.3702
R22021 vdd.n248 vdd.n245 7.3702
R22022 vdd.n205 vdd.n202 7.3702
R22023 vdd.n146 vdd.n143 7.3702
R22024 vdd.n104 vdd.n101 7.3702
R22025 vdd.n45 vdd.n42 7.3702
R22026 vdd.n1726 vdd.n1723 7.3702
R22027 vdd.n1785 vdd.n1782 7.3702
R22028 vdd.n1624 vdd.n1621 7.3702
R22029 vdd.n1683 vdd.n1680 7.3702
R22030 vdd.n1523 vdd.n1520 7.3702
R22031 vdd.n1582 vdd.n1579 7.3702
R22032 vdd.n1884 vdd.t43 7.1425
R22033 vdd.n679 vdd.t107 7.1425
R22034 vdd.n1358 vdd.n1357 6.98232
R22035 vdd.n2039 vdd.n2038 6.98232
R22036 vdd.n566 vdd.n565 6.98232
R22037 vdd.n3141 vdd.n3138 6.98232
R22038 vdd.t82 vdd.n1097 6.91577
R22039 vdd.n3264 vdd.t94 6.91577
R22040 vdd.n1843 vdd.t69 6.68904
R22041 vdd.n3280 vdd.t8 6.68904
R22042 vdd.t47 vdd.n1126 6.46231
R22043 vdd.n3308 vdd.t88 6.46231
R22044 vdd.n3400 vdd.n333 6.38151
R22045 vdd.n1812 vdd.n1811 6.38151
R22046 vdd.n1494 vdd.t76 6.23558
R22047 vdd.t32 vdd.n344 6.23558
R22048 vdd.t92 vdd.n1154 6.00885
R22049 vdd.n2412 vdd.t161 6.00885
R22050 vdd.n2912 vdd.t151 6.00885
R22051 vdd.n3379 vdd.t36 6.00885
R22052 vdd.n1033 vdd.t224 5.89549
R22053 vdd.t181 vdd.n851 5.89549
R22054 vdd.n308 vdd.n307 5.81868
R22055 vdd.n249 vdd.n248 5.81868
R22056 vdd.n206 vdd.n205 5.81868
R22057 vdd.n147 vdd.n146 5.81868
R22058 vdd.n105 vdd.n104 5.81868
R22059 vdd.n46 vdd.n45 5.81868
R22060 vdd.n1727 vdd.n1726 5.81868
R22061 vdd.n1786 vdd.n1785 5.81868
R22062 vdd.n1625 vdd.n1624 5.81868
R22063 vdd.n1684 vdd.n1683 5.81868
R22064 vdd.n1524 vdd.n1523 5.81868
R22065 vdd.n1583 vdd.n1582 5.81868
R22066 vdd.n1453 vdd.t252 5.78212
R22067 vdd.t220 vdd.n1037 5.78212
R22068 vdd.n2156 vdd.t205 5.78212
R22069 vdd.n2781 vdd.t213 5.78212
R22070 vdd.n846 vdd.t209 5.78212
R22071 vdd.n3370 vdd.t30 5.78212
R22072 vdd.n2540 vdd.n2539 5.77611
R22073 vdd.n2283 vdd.n2153 5.77611
R22074 vdd.n2794 vdd.n2793 5.77611
R22075 vdd.n3000 vdd.n2999 5.77611
R22076 vdd.n3064 vdd.n801 5.77611
R22077 vdd.n2704 vdd.n2644 5.77611
R22078 vdd.n2465 vdd.n967 5.77611
R22079 vdd.n2213 vdd.n2212 5.77611
R22080 vdd.n1320 vdd.n1319 5.62474
R22081 vdd.n2335 vdd.n2332 5.62474
R22082 vdd.n3351 vdd.n428 5.62474
R22083 vdd.n3225 vdd.n690 5.62474
R22084 vdd.n1177 vdd.t252 5.55539
R22085 vdd.t30 vdd.n3369 5.55539
R22086 vdd.t165 vdd.n989 5.44203
R22087 vdd.n893 vdd.t155 5.44203
R22088 vdd.n1469 vdd.t92 5.32866
R22089 vdd.t36 vdd.n3378 5.32866
R22090 vdd.n1485 vdd.t76 5.10193
R22091 vdd.t131 vdd.n1012 5.10193
R22092 vdd.n1002 vdd.t139 5.10193
R22093 vdd.t152 vdd.n880 5.10193
R22094 vdd.n870 vdd.t136 5.10193
R22095 vdd.n3387 vdd.t32 5.10193
R22096 vdd.n311 vdd.n302 5.04292
R22097 vdd.n252 vdd.n243 5.04292
R22098 vdd.n209 vdd.n200 5.04292
R22099 vdd.n150 vdd.n141 5.04292
R22100 vdd.n108 vdd.n99 5.04292
R22101 vdd.n49 vdd.n40 5.04292
R22102 vdd.n1730 vdd.n1721 5.04292
R22103 vdd.n1789 vdd.n1780 5.04292
R22104 vdd.n1628 vdd.n1619 5.04292
R22105 vdd.n1687 vdd.n1678 5.04292
R22106 vdd.n1527 vdd.n1518 5.04292
R22107 vdd.n1586 vdd.n1577 5.04292
R22108 vdd.n1817 vdd.t47 4.8752
R22109 vdd.t128 vdd.t137 4.8752
R22110 vdd.t162 vdd.t149 4.8752
R22111 vdd.t140 vdd.t123 4.8752
R22112 vdd.t163 vdd.t144 4.8752
R22113 vdd.t88 vdd.n340 4.8752
R22114 vdd.n2541 vdd.n2540 4.83952
R22115 vdd.n2153 vdd.n2149 4.83952
R22116 vdd.n2795 vdd.n2794 4.83952
R22117 vdd.n3001 vdd.n3000 4.83952
R22118 vdd.n801 vdd.n796 4.83952
R22119 vdd.n2701 vdd.n2644 4.83952
R22120 vdd.n2468 vdd.n967 4.83952
R22121 vdd.n2212 vdd.n2211 4.83952
R22122 vdd.n2007 vdd.n1065 4.74817
R22123 vdd.n2002 vdd.n1066 4.74817
R22124 vdd.n1904 vdd.n1901 4.74817
R22125 vdd.n2316 vdd.n1905 4.74817
R22126 vdd.n2318 vdd.n1904 4.74817
R22127 vdd.n2317 vdd.n2316 4.74817
R22128 vdd.n3218 vdd.n3217 4.74817
R22129 vdd.n3215 vdd.n3214 4.74817
R22130 vdd.n3215 vdd.n732 4.74817
R22131 vdd.n3217 vdd.n729 4.74817
R22132 vdd.n3100 vdd.n784 4.74817
R22133 vdd.n3096 vdd.n3094 4.74817
R22134 vdd.n3099 vdd.n3094 4.74817
R22135 vdd.n3103 vdd.n784 4.74817
R22136 vdd.n2003 vdd.n1065 4.74817
R22137 vdd.n1068 vdd.n1066 4.74817
R22138 vdd.n333 vdd.n332 4.7074
R22139 vdd.n231 vdd.n230 4.7074
R22140 vdd.n1811 vdd.n1810 4.7074
R22141 vdd.n1709 vdd.n1708 4.7074
R22142 vdd.n1120 vdd.t69 4.64847
R22143 vdd.n3289 vdd.t8 4.64847
R22144 vdd.n2418 vdd.t153 4.53511
R22145 vdd.n2906 vdd.t132 4.53511
R22146 vdd.n1859 vdd.t82 4.42174
R22147 vdd.t94 vdd.n655 4.42174
R22148 vdd.n2450 vdd.t134 4.30838
R22149 vdd.n2876 vdd.t124 4.30838
R22150 vdd.n312 vdd.n300 4.26717
R22151 vdd.n253 vdd.n241 4.26717
R22152 vdd.n210 vdd.n198 4.26717
R22153 vdd.n151 vdd.n139 4.26717
R22154 vdd.n109 vdd.n97 4.26717
R22155 vdd.n50 vdd.n38 4.26717
R22156 vdd.n1731 vdd.n1719 4.26717
R22157 vdd.n1790 vdd.n1778 4.26717
R22158 vdd.n1629 vdd.n1617 4.26717
R22159 vdd.n1688 vdd.n1676 4.26717
R22160 vdd.n1528 vdd.n1516 4.26717
R22161 vdd.n1587 vdd.n1575 4.26717
R22162 vdd.n1875 vdd.t43 4.19501
R22163 vdd.n3248 vdd.t107 4.19501
R22164 vdd.n333 vdd.n231 4.10845
R22165 vdd.n1811 vdd.n1709 4.10845
R22166 vdd.n289 vdd.t97 4.06363
R22167 vdd.n289 vdd.t31 4.06363
R22168 vdd.n287 vdd.t248 4.06363
R22169 vdd.n287 vdd.t290 4.06363
R22170 vdd.n285 vdd.t91 4.06363
R22171 vdd.n285 vdd.t266 4.06363
R22172 vdd.n283 vdd.t1 4.06363
R22173 vdd.n283 vdd.t33 4.06363
R22174 vdd.n281 vdd.t89 4.06363
R22175 vdd.n281 vdd.t3 4.06363
R22176 vdd.n279 vdd.t74 4.06363
R22177 vdd.n279 vdd.t104 4.06363
R22178 vdd.n277 vdd.t86 4.06363
R22179 vdd.n277 vdd.t38 4.06363
R22180 vdd.n275 vdd.t95 4.06363
R22181 vdd.n275 vdd.t288 4.06363
R22182 vdd.n273 vdd.t121 4.06363
R22183 vdd.n273 vdd.t295 4.06363
R22184 vdd.n187 vdd.t285 4.06363
R22185 vdd.n187 vdd.t273 4.06363
R22186 vdd.n185 vdd.t279 4.06363
R22187 vdd.n185 vdd.t292 4.06363
R22188 vdd.n183 vdd.t287 4.06363
R22189 vdd.n183 vdd.t284 4.06363
R22190 vdd.n181 vdd.t39 4.06363
R22191 vdd.n181 vdd.t51 4.06363
R22192 vdd.n179 vdd.t256 4.06363
R22193 vdd.n179 vdd.t40 4.06363
R22194 vdd.n177 vdd.t267 4.06363
R22195 vdd.n177 vdd.t68 4.06363
R22196 vdd.n175 vdd.t113 4.06363
R22197 vdd.n175 vdd.t9 4.06363
R22198 vdd.n173 vdd.t282 4.06363
R22199 vdd.n173 vdd.t103 4.06363
R22200 vdd.n171 vdd.t106 4.06363
R22201 vdd.n171 vdd.t278 4.06363
R22202 vdd.n86 vdd.t61 4.06363
R22203 vdd.n86 vdd.t167 4.06363
R22204 vdd.n84 vdd.t37 4.06363
R22205 vdd.n84 vdd.t81 4.06363
R22206 vdd.n82 vdd.t268 4.06363
R22207 vdd.n82 vdd.t293 4.06363
R22208 vdd.n80 vdd.t50 4.06363
R22209 vdd.n80 vdd.t274 4.06363
R22210 vdd.n78 vdd.t255 4.06363
R22211 vdd.n78 vdd.t66 4.06363
R22212 vdd.n76 vdd.t291 4.06363
R22213 vdd.n76 vdd.t168 4.06363
R22214 vdd.n74 vdd.t117 4.06363
R22215 vdd.n74 vdd.t71 4.06363
R22216 vdd.n72 vdd.t250 4.06363
R22217 vdd.n72 vdd.t264 4.06363
R22218 vdd.n70 vdd.t286 4.06363
R22219 vdd.n70 vdd.t272 4.06363
R22220 vdd.n1751 vdd.t62 4.06363
R22221 vdd.n1751 vdd.t55 4.06363
R22222 vdd.n1753 vdd.t259 4.06363
R22223 vdd.n1753 vdd.t87 4.06363
R22224 vdd.n1755 vdd.t110 4.06363
R22225 vdd.n1755 vdd.t57 4.06363
R22226 vdd.n1757 vdd.t11 4.06363
R22227 vdd.n1757 vdd.t245 4.06363
R22228 vdd.n1759 vdd.t281 4.06363
R22229 vdd.n1759 vdd.t100 4.06363
R22230 vdd.n1761 vdd.t270 4.06363
R22231 vdd.n1761 vdd.t280 4.06363
R22232 vdd.n1763 vdd.t118 4.06363
R22233 vdd.n1763 vdd.t120 4.06363
R22234 vdd.n1765 vdd.t99 4.06363
R22235 vdd.n1765 vdd.t93 4.06363
R22236 vdd.n1767 vdd.t260 4.06363
R22237 vdd.n1767 vdd.t29 4.06363
R22238 vdd.n1649 vdd.t46 4.06363
R22239 vdd.n1649 vdd.t294 4.06363
R22240 vdd.n1651 vdd.t114 4.06363
R22241 vdd.n1651 vdd.t83 4.06363
R22242 vdd.n1653 vdd.t72 4.06363
R22243 vdd.n1653 vdd.t42 4.06363
R22244 vdd.n1655 vdd.t258 4.06363
R22245 vdd.n1655 vdd.t84 4.06363
R22246 vdd.n1657 vdd.t7 4.06363
R22247 vdd.n1657 vdd.t63 4.06363
R22248 vdd.n1659 vdd.t262 4.06363
R22249 vdd.n1659 vdd.t5 4.06363
R22250 vdd.n1661 vdd.t276 4.06363
R22251 vdd.n1661 vdd.t277 4.06363
R22252 vdd.n1663 vdd.t96 4.06363
R22253 vdd.n1663 vdd.t254 4.06363
R22254 vdd.n1665 vdd.t253 4.06363
R22255 vdd.n1665 vdd.t75 4.06363
R22256 vdd.n1548 vdd.t275 4.06363
R22257 vdd.n1548 vdd.t257 4.06363
R22258 vdd.n1550 vdd.t65 4.06363
R22259 vdd.n1550 vdd.t246 4.06363
R22260 vdd.n1552 vdd.t70 4.06363
R22261 vdd.n1552 vdd.t116 4.06363
R22262 vdd.n1554 vdd.t109 4.06363
R22263 vdd.n1554 vdd.t35 4.06363
R22264 vdd.n1556 vdd.t98 4.06363
R22265 vdd.n1556 vdd.t48 4.06363
R22266 vdd.n1558 vdd.t77 4.06363
R22267 vdd.n1558 vdd.t49 4.06363
R22268 vdd.n1560 vdd.t53 4.06363
R22269 vdd.n1560 vdd.t249 4.06363
R22270 vdd.n1562 vdd.t79 4.06363
R22271 vdd.n1562 vdd.t261 4.06363
R22272 vdd.n1564 vdd.t289 4.06363
R22273 vdd.n1564 vdd.t263 4.06363
R22274 vdd.n26 vdd.t13 3.9605
R22275 vdd.n26 vdd.t14 3.9605
R22276 vdd.n23 vdd.t12 3.9605
R22277 vdd.n23 vdd.t20 3.9605
R22278 vdd.n21 vdd.t19 3.9605
R22279 vdd.n21 vdd.t16 3.9605
R22280 vdd.n20 vdd.t17 3.9605
R22281 vdd.n20 vdd.t18 3.9605
R22282 vdd.n15 vdd.t27 3.9605
R22283 vdd.n15 vdd.t15 3.9605
R22284 vdd.n16 vdd.t22 3.9605
R22285 vdd.n16 vdd.t23 3.9605
R22286 vdd.n18 vdd.t26 3.9605
R22287 vdd.n18 vdd.t25 3.9605
R22288 vdd.n25 vdd.t24 3.9605
R22289 vdd.n25 vdd.t21 3.9605
R22290 vdd.n7 vdd.t164 3.61217
R22291 vdd.n7 vdd.t133 3.61217
R22292 vdd.n8 vdd.t141 3.61217
R22293 vdd.n8 vdd.t156 3.61217
R22294 vdd.n10 vdd.t148 3.61217
R22295 vdd.n10 vdd.t125 3.61217
R22296 vdd.n12 vdd.t130 3.61217
R22297 vdd.n12 vdd.t146 3.61217
R22298 vdd.n5 vdd.t158 3.61217
R22299 vdd.n5 vdd.t143 3.61217
R22300 vdd.n3 vdd.t135 3.61217
R22301 vdd.n3 vdd.t160 3.61217
R22302 vdd.n1 vdd.t166 3.61217
R22303 vdd.n1 vdd.t150 3.61217
R22304 vdd.n0 vdd.t154 3.61217
R22305 vdd.n0 vdd.t138 3.61217
R22306 vdd.n316 vdd.n315 3.49141
R22307 vdd.n257 vdd.n256 3.49141
R22308 vdd.n214 vdd.n213 3.49141
R22309 vdd.n155 vdd.n154 3.49141
R22310 vdd.n113 vdd.n112 3.49141
R22311 vdd.n54 vdd.n53 3.49141
R22312 vdd.n1735 vdd.n1734 3.49141
R22313 vdd.n1794 vdd.n1793 3.49141
R22314 vdd.n1633 vdd.n1632 3.49141
R22315 vdd.n1692 vdd.n1691 3.49141
R22316 vdd.n1532 vdd.n1531 3.49141
R22317 vdd.n1591 vdd.n1590 3.49141
R22318 vdd.n2156 vdd.t134 3.40145
R22319 vdd.n2604 vdd.t157 3.40145
R22320 vdd.n2857 vdd.t145 3.40145
R22321 vdd.n2781 vdd.t124 3.40145
R22322 vdd.n1876 vdd.t54 3.28809
R22323 vdd.n3247 vdd.t105 3.28809
R22324 vdd.n2257 vdd.t153 3.17472
R22325 vdd.n2760 vdd.t132 3.17472
R22326 vdd.t64 vdd.n1104 3.06136
R22327 vdd.n3272 vdd.t102 3.06136
R22328 vdd.n1834 vdd.t34 2.83463
R22329 vdd.n644 vdd.t73 2.83463
R22330 vdd.n319 vdd.n298 2.71565
R22331 vdd.n260 vdd.n239 2.71565
R22332 vdd.n217 vdd.n196 2.71565
R22333 vdd.n158 vdd.n137 2.71565
R22334 vdd.n116 vdd.n95 2.71565
R22335 vdd.n57 vdd.n36 2.71565
R22336 vdd.n1738 vdd.n1717 2.71565
R22337 vdd.n1797 vdd.n1776 2.71565
R22338 vdd.n1636 vdd.n1615 2.71565
R22339 vdd.n1695 vdd.n1674 2.71565
R22340 vdd.n1535 vdd.n1514 2.71565
R22341 vdd.n1594 vdd.n1573 2.71565
R22342 vdd.t6 vdd.n1132 2.6079
R22343 vdd.n2406 vdd.t131 2.6079
R22344 vdd.n2430 vdd.t139 2.6079
R22345 vdd.n2894 vdd.t152 2.6079
R22346 vdd.n2918 vdd.t136 2.6079
R22347 vdd.n3395 vdd.t2 2.6079
R22348 vdd.n2924 vdd.n2923 2.49806
R22349 vdd.n2398 vdd.n2397 2.49806
R22350 vdd.n306 vdd.n305 2.4129
R22351 vdd.n247 vdd.n246 2.4129
R22352 vdd.n204 vdd.n203 2.4129
R22353 vdd.n145 vdd.n144 2.4129
R22354 vdd.n103 vdd.n102 2.4129
R22355 vdd.n44 vdd.n43 2.4129
R22356 vdd.n1725 vdd.n1724 2.4129
R22357 vdd.n1784 vdd.n1783 2.4129
R22358 vdd.n1623 vdd.n1622 2.4129
R22359 vdd.n1682 vdd.n1681 2.4129
R22360 vdd.n1522 vdd.n1521 2.4129
R22361 vdd.n1581 vdd.n1580 2.4129
R22362 vdd.n1486 vdd.t119 2.38117
R22363 vdd.n1894 vdd.t177 2.38117
R22364 vdd.n3231 vdd.t170 2.38117
R22365 vdd.n3386 vdd.t90 2.38117
R22366 vdd.n2315 vdd.n1904 2.27742
R22367 vdd.n2316 vdd.n2315 2.27742
R22368 vdd.n3216 vdd.n3215 2.27742
R22369 vdd.n3217 vdd.n3216 2.27742
R22370 vdd.n3094 vdd.n3093 2.27742
R22371 vdd.n3093 vdd.n784 2.27742
R22372 vdd.n2338 vdd.n1065 2.27742
R22373 vdd.n2338 vdd.n1066 2.27742
R22374 vdd.n2430 vdd.t165 2.2678
R22375 vdd.n2894 vdd.t155 2.2678
R22376 vdd.t78 vdd.n1161 2.15444
R22377 vdd.n3377 vdd.t80 2.15444
R22378 vdd.t149 vdd.n983 2.04107
R22379 vdd.n900 vdd.t140 2.04107
R22380 vdd.n320 vdd.n296 1.93989
R22381 vdd.n261 vdd.n237 1.93989
R22382 vdd.n218 vdd.n194 1.93989
R22383 vdd.n159 vdd.n135 1.93989
R22384 vdd.n117 vdd.n93 1.93989
R22385 vdd.n58 vdd.n34 1.93989
R22386 vdd.n1739 vdd.n1715 1.93989
R22387 vdd.n1798 vdd.n1774 1.93989
R22388 vdd.n1637 vdd.n1613 1.93989
R22389 vdd.n1696 vdd.n1672 1.93989
R22390 vdd.n1536 vdd.n1512 1.93989
R22391 vdd.n1595 vdd.n1571 1.93989
R22392 vdd.n1444 vdd.t58 1.92771
R22393 vdd.n2381 vdd.t220 1.92771
R22394 vdd.n2457 vdd.t205 1.92771
R22395 vdd.n2870 vdd.t213 1.92771
R22396 vdd.n2989 vdd.t209 1.92771
R22397 vdd.t111 vdd.n375 1.92771
R22398 vdd.n1452 vdd.t28 1.70098
R22399 vdd.n2257 vdd.t161 1.70098
R22400 vdd.n1008 vdd.t128 1.70098
R22401 vdd.t144 vdd.n874 1.70098
R22402 vdd.n2760 vdd.t151 1.70098
R22403 vdd.n3371 vdd.t60 1.70098
R22404 vdd.n1477 vdd.t52 1.47425
R22405 vdd.n361 vdd.t265 1.47425
R22406 vdd.n1143 vdd.t4 1.24752
R22407 vdd.t0 vdd.n3393 1.24752
R22408 vdd.n331 vdd.n291 1.16414
R22409 vdd.n324 vdd.n323 1.16414
R22410 vdd.n272 vdd.n232 1.16414
R22411 vdd.n265 vdd.n264 1.16414
R22412 vdd.n229 vdd.n189 1.16414
R22413 vdd.n222 vdd.n221 1.16414
R22414 vdd.n170 vdd.n130 1.16414
R22415 vdd.n163 vdd.n162 1.16414
R22416 vdd.n128 vdd.n88 1.16414
R22417 vdd.n121 vdd.n120 1.16414
R22418 vdd.n69 vdd.n29 1.16414
R22419 vdd.n62 vdd.n61 1.16414
R22420 vdd.n1750 vdd.n1710 1.16414
R22421 vdd.n1743 vdd.n1742 1.16414
R22422 vdd.n1809 vdd.n1769 1.16414
R22423 vdd.n1802 vdd.n1801 1.16414
R22424 vdd.n1648 vdd.n1608 1.16414
R22425 vdd.n1641 vdd.n1640 1.16414
R22426 vdd.n1707 vdd.n1667 1.16414
R22427 vdd.n1700 vdd.n1699 1.16414
R22428 vdd.n1547 vdd.n1507 1.16414
R22429 vdd.n1540 vdd.n1539 1.16414
R22430 vdd.n1606 vdd.n1566 1.16414
R22431 vdd.n1599 vdd.n1598 1.16414
R22432 vdd.n2424 vdd.t137 1.13415
R22433 vdd.n2900 vdd.t163 1.13415
R22434 vdd.n1826 vdd.t10 1.02079
R22435 vdd.t224 vdd.t127 1.02079
R22436 vdd.t126 vdd.t181 1.02079
R22437 vdd.t67 vdd.n633 1.02079
R22438 vdd.n1323 vdd.n1319 0.970197
R22439 vdd.n2336 vdd.n2335 0.970197
R22440 vdd.n618 vdd.n428 0.970197
R22441 vdd.n3095 vdd.n690 0.970197
R22442 vdd.n1812 vdd.n28 0.90431
R22443 vdd vdd.n3400 0.896477
R22444 vdd.n1842 vdd.t41 0.794056
R22445 vdd.n2400 vdd.t127 0.794056
R22446 vdd.n2436 vdd.t162 0.794056
R22447 vdd.n2888 vdd.t123 0.794056
R22448 vdd.n2926 vdd.t126 0.794056
R22449 vdd.n3281 vdd.t85 0.794056
R22450 vdd.n1867 vdd.t45 0.567326
R22451 vdd.t271 vdd.n662 0.567326
R22452 vdd.n2326 vdd.n2325 0.530988
R22453 vdd.n726 vdd.n682 0.530988
R22454 vdd.n464 vdd.n391 0.530988
R22455 vdd.n3350 vdd.n3349 0.530988
R22456 vdd.n3227 vdd.n3226 0.530988
R22457 vdd.n1889 vdd.n1067 0.530988
R22458 vdd.n1321 vdd.n1186 0.530988
R22459 vdd.n1423 vdd.n1422 0.530988
R22460 vdd.n4 vdd.n2 0.459552
R22461 vdd.n11 vdd.n9 0.459552
R22462 vdd.n329 vdd.n328 0.388379
R22463 vdd.n295 vdd.n293 0.388379
R22464 vdd.n270 vdd.n269 0.388379
R22465 vdd.n236 vdd.n234 0.388379
R22466 vdd.n227 vdd.n226 0.388379
R22467 vdd.n193 vdd.n191 0.388379
R22468 vdd.n168 vdd.n167 0.388379
R22469 vdd.n134 vdd.n132 0.388379
R22470 vdd.n126 vdd.n125 0.388379
R22471 vdd.n92 vdd.n90 0.388379
R22472 vdd.n67 vdd.n66 0.388379
R22473 vdd.n33 vdd.n31 0.388379
R22474 vdd.n1748 vdd.n1747 0.388379
R22475 vdd.n1714 vdd.n1712 0.388379
R22476 vdd.n1807 vdd.n1806 0.388379
R22477 vdd.n1773 vdd.n1771 0.388379
R22478 vdd.n1646 vdd.n1645 0.388379
R22479 vdd.n1612 vdd.n1610 0.388379
R22480 vdd.n1705 vdd.n1704 0.388379
R22481 vdd.n1671 vdd.n1669 0.388379
R22482 vdd.n1545 vdd.n1544 0.388379
R22483 vdd.n1511 vdd.n1509 0.388379
R22484 vdd.n1604 vdd.n1603 0.388379
R22485 vdd.n1570 vdd.n1568 0.388379
R22486 vdd.n19 vdd.n17 0.387128
R22487 vdd.n24 vdd.n22 0.387128
R22488 vdd.n6 vdd.n4 0.358259
R22489 vdd.n13 vdd.n11 0.358259
R22490 vdd.n276 vdd.n274 0.358259
R22491 vdd.n278 vdd.n276 0.358259
R22492 vdd.n280 vdd.n278 0.358259
R22493 vdd.n282 vdd.n280 0.358259
R22494 vdd.n284 vdd.n282 0.358259
R22495 vdd.n286 vdd.n284 0.358259
R22496 vdd.n288 vdd.n286 0.358259
R22497 vdd.n290 vdd.n288 0.358259
R22498 vdd.n332 vdd.n290 0.358259
R22499 vdd.n174 vdd.n172 0.358259
R22500 vdd.n176 vdd.n174 0.358259
R22501 vdd.n178 vdd.n176 0.358259
R22502 vdd.n180 vdd.n178 0.358259
R22503 vdd.n182 vdd.n180 0.358259
R22504 vdd.n184 vdd.n182 0.358259
R22505 vdd.n186 vdd.n184 0.358259
R22506 vdd.n188 vdd.n186 0.358259
R22507 vdd.n230 vdd.n188 0.358259
R22508 vdd.n73 vdd.n71 0.358259
R22509 vdd.n75 vdd.n73 0.358259
R22510 vdd.n77 vdd.n75 0.358259
R22511 vdd.n79 vdd.n77 0.358259
R22512 vdd.n81 vdd.n79 0.358259
R22513 vdd.n83 vdd.n81 0.358259
R22514 vdd.n85 vdd.n83 0.358259
R22515 vdd.n87 vdd.n85 0.358259
R22516 vdd.n129 vdd.n87 0.358259
R22517 vdd.n1810 vdd.n1768 0.358259
R22518 vdd.n1768 vdd.n1766 0.358259
R22519 vdd.n1766 vdd.n1764 0.358259
R22520 vdd.n1764 vdd.n1762 0.358259
R22521 vdd.n1762 vdd.n1760 0.358259
R22522 vdd.n1760 vdd.n1758 0.358259
R22523 vdd.n1758 vdd.n1756 0.358259
R22524 vdd.n1756 vdd.n1754 0.358259
R22525 vdd.n1754 vdd.n1752 0.358259
R22526 vdd.n1708 vdd.n1666 0.358259
R22527 vdd.n1666 vdd.n1664 0.358259
R22528 vdd.n1664 vdd.n1662 0.358259
R22529 vdd.n1662 vdd.n1660 0.358259
R22530 vdd.n1660 vdd.n1658 0.358259
R22531 vdd.n1658 vdd.n1656 0.358259
R22532 vdd.n1656 vdd.n1654 0.358259
R22533 vdd.n1654 vdd.n1652 0.358259
R22534 vdd.n1652 vdd.n1650 0.358259
R22535 vdd.n1607 vdd.n1565 0.358259
R22536 vdd.n1565 vdd.n1563 0.358259
R22537 vdd.n1563 vdd.n1561 0.358259
R22538 vdd.n1561 vdd.n1559 0.358259
R22539 vdd.n1559 vdd.n1557 0.358259
R22540 vdd.n1557 vdd.n1555 0.358259
R22541 vdd.n1555 vdd.n1553 0.358259
R22542 vdd.n1553 vdd.n1551 0.358259
R22543 vdd.n1551 vdd.n1549 0.358259
R22544 vdd.n14 vdd.n6 0.334552
R22545 vdd.n14 vdd.n13 0.334552
R22546 vdd.n27 vdd.n19 0.21707
R22547 vdd.n27 vdd.n24 0.21707
R22548 vdd.n330 vdd.n292 0.155672
R22549 vdd.n322 vdd.n292 0.155672
R22550 vdd.n322 vdd.n321 0.155672
R22551 vdd.n321 vdd.n297 0.155672
R22552 vdd.n314 vdd.n297 0.155672
R22553 vdd.n314 vdd.n313 0.155672
R22554 vdd.n313 vdd.n301 0.155672
R22555 vdd.n306 vdd.n301 0.155672
R22556 vdd.n271 vdd.n233 0.155672
R22557 vdd.n263 vdd.n233 0.155672
R22558 vdd.n263 vdd.n262 0.155672
R22559 vdd.n262 vdd.n238 0.155672
R22560 vdd.n255 vdd.n238 0.155672
R22561 vdd.n255 vdd.n254 0.155672
R22562 vdd.n254 vdd.n242 0.155672
R22563 vdd.n247 vdd.n242 0.155672
R22564 vdd.n228 vdd.n190 0.155672
R22565 vdd.n220 vdd.n190 0.155672
R22566 vdd.n220 vdd.n219 0.155672
R22567 vdd.n219 vdd.n195 0.155672
R22568 vdd.n212 vdd.n195 0.155672
R22569 vdd.n212 vdd.n211 0.155672
R22570 vdd.n211 vdd.n199 0.155672
R22571 vdd.n204 vdd.n199 0.155672
R22572 vdd.n169 vdd.n131 0.155672
R22573 vdd.n161 vdd.n131 0.155672
R22574 vdd.n161 vdd.n160 0.155672
R22575 vdd.n160 vdd.n136 0.155672
R22576 vdd.n153 vdd.n136 0.155672
R22577 vdd.n153 vdd.n152 0.155672
R22578 vdd.n152 vdd.n140 0.155672
R22579 vdd.n145 vdd.n140 0.155672
R22580 vdd.n127 vdd.n89 0.155672
R22581 vdd.n119 vdd.n89 0.155672
R22582 vdd.n119 vdd.n118 0.155672
R22583 vdd.n118 vdd.n94 0.155672
R22584 vdd.n111 vdd.n94 0.155672
R22585 vdd.n111 vdd.n110 0.155672
R22586 vdd.n110 vdd.n98 0.155672
R22587 vdd.n103 vdd.n98 0.155672
R22588 vdd.n68 vdd.n30 0.155672
R22589 vdd.n60 vdd.n30 0.155672
R22590 vdd.n60 vdd.n59 0.155672
R22591 vdd.n59 vdd.n35 0.155672
R22592 vdd.n52 vdd.n35 0.155672
R22593 vdd.n52 vdd.n51 0.155672
R22594 vdd.n51 vdd.n39 0.155672
R22595 vdd.n44 vdd.n39 0.155672
R22596 vdd.n1749 vdd.n1711 0.155672
R22597 vdd.n1741 vdd.n1711 0.155672
R22598 vdd.n1741 vdd.n1740 0.155672
R22599 vdd.n1740 vdd.n1716 0.155672
R22600 vdd.n1733 vdd.n1716 0.155672
R22601 vdd.n1733 vdd.n1732 0.155672
R22602 vdd.n1732 vdd.n1720 0.155672
R22603 vdd.n1725 vdd.n1720 0.155672
R22604 vdd.n1808 vdd.n1770 0.155672
R22605 vdd.n1800 vdd.n1770 0.155672
R22606 vdd.n1800 vdd.n1799 0.155672
R22607 vdd.n1799 vdd.n1775 0.155672
R22608 vdd.n1792 vdd.n1775 0.155672
R22609 vdd.n1792 vdd.n1791 0.155672
R22610 vdd.n1791 vdd.n1779 0.155672
R22611 vdd.n1784 vdd.n1779 0.155672
R22612 vdd.n1647 vdd.n1609 0.155672
R22613 vdd.n1639 vdd.n1609 0.155672
R22614 vdd.n1639 vdd.n1638 0.155672
R22615 vdd.n1638 vdd.n1614 0.155672
R22616 vdd.n1631 vdd.n1614 0.155672
R22617 vdd.n1631 vdd.n1630 0.155672
R22618 vdd.n1630 vdd.n1618 0.155672
R22619 vdd.n1623 vdd.n1618 0.155672
R22620 vdd.n1706 vdd.n1668 0.155672
R22621 vdd.n1698 vdd.n1668 0.155672
R22622 vdd.n1698 vdd.n1697 0.155672
R22623 vdd.n1697 vdd.n1673 0.155672
R22624 vdd.n1690 vdd.n1673 0.155672
R22625 vdd.n1690 vdd.n1689 0.155672
R22626 vdd.n1689 vdd.n1677 0.155672
R22627 vdd.n1682 vdd.n1677 0.155672
R22628 vdd.n1546 vdd.n1508 0.155672
R22629 vdd.n1538 vdd.n1508 0.155672
R22630 vdd.n1538 vdd.n1537 0.155672
R22631 vdd.n1537 vdd.n1513 0.155672
R22632 vdd.n1530 vdd.n1513 0.155672
R22633 vdd.n1530 vdd.n1529 0.155672
R22634 vdd.n1529 vdd.n1517 0.155672
R22635 vdd.n1522 vdd.n1517 0.155672
R22636 vdd.n1605 vdd.n1567 0.155672
R22637 vdd.n1597 vdd.n1567 0.155672
R22638 vdd.n1597 vdd.n1596 0.155672
R22639 vdd.n1596 vdd.n1572 0.155672
R22640 vdd.n1589 vdd.n1572 0.155672
R22641 vdd.n1589 vdd.n1588 0.155672
R22642 vdd.n1588 vdd.n1576 0.155672
R22643 vdd.n1581 vdd.n1576 0.155672
R22644 vdd.n2101 vdd.n1906 0.152939
R22645 vdd.n1912 vdd.n1906 0.152939
R22646 vdd.n1913 vdd.n1912 0.152939
R22647 vdd.n1914 vdd.n1913 0.152939
R22648 vdd.n1915 vdd.n1914 0.152939
R22649 vdd.n1919 vdd.n1915 0.152939
R22650 vdd.n1920 vdd.n1919 0.152939
R22651 vdd.n1921 vdd.n1920 0.152939
R22652 vdd.n1922 vdd.n1921 0.152939
R22653 vdd.n1926 vdd.n1922 0.152939
R22654 vdd.n1927 vdd.n1926 0.152939
R22655 vdd.n1928 vdd.n1927 0.152939
R22656 vdd.n2076 vdd.n1928 0.152939
R22657 vdd.n2076 vdd.n2075 0.152939
R22658 vdd.n2075 vdd.n2074 0.152939
R22659 vdd.n2074 vdd.n1934 0.152939
R22660 vdd.n1939 vdd.n1934 0.152939
R22661 vdd.n1940 vdd.n1939 0.152939
R22662 vdd.n1941 vdd.n1940 0.152939
R22663 vdd.n1945 vdd.n1941 0.152939
R22664 vdd.n1946 vdd.n1945 0.152939
R22665 vdd.n1947 vdd.n1946 0.152939
R22666 vdd.n1948 vdd.n1947 0.152939
R22667 vdd.n1952 vdd.n1948 0.152939
R22668 vdd.n1953 vdd.n1952 0.152939
R22669 vdd.n1954 vdd.n1953 0.152939
R22670 vdd.n1955 vdd.n1954 0.152939
R22671 vdd.n1959 vdd.n1955 0.152939
R22672 vdd.n1960 vdd.n1959 0.152939
R22673 vdd.n1961 vdd.n1960 0.152939
R22674 vdd.n1962 vdd.n1961 0.152939
R22675 vdd.n1966 vdd.n1962 0.152939
R22676 vdd.n1967 vdd.n1966 0.152939
R22677 vdd.n1968 vdd.n1967 0.152939
R22678 vdd.n2037 vdd.n1968 0.152939
R22679 vdd.n2037 vdd.n2036 0.152939
R22680 vdd.n2036 vdd.n2035 0.152939
R22681 vdd.n2035 vdd.n1974 0.152939
R22682 vdd.n1979 vdd.n1974 0.152939
R22683 vdd.n1980 vdd.n1979 0.152939
R22684 vdd.n1981 vdd.n1980 0.152939
R22685 vdd.n1985 vdd.n1981 0.152939
R22686 vdd.n1986 vdd.n1985 0.152939
R22687 vdd.n1987 vdd.n1986 0.152939
R22688 vdd.n1988 vdd.n1987 0.152939
R22689 vdd.n1992 vdd.n1988 0.152939
R22690 vdd.n1993 vdd.n1992 0.152939
R22691 vdd.n1994 vdd.n1993 0.152939
R22692 vdd.n1995 vdd.n1994 0.152939
R22693 vdd.n1996 vdd.n1995 0.152939
R22694 vdd.n1996 vdd.n1064 0.152939
R22695 vdd.n2325 vdd.n1900 0.152939
R22696 vdd.n1814 vdd.n1123 0.152939
R22697 vdd.n1829 vdd.n1123 0.152939
R22698 vdd.n1830 vdd.n1829 0.152939
R22699 vdd.n1831 vdd.n1830 0.152939
R22700 vdd.n1831 vdd.n1112 0.152939
R22701 vdd.n1846 vdd.n1112 0.152939
R22702 vdd.n1847 vdd.n1846 0.152939
R22703 vdd.n1848 vdd.n1847 0.152939
R22704 vdd.n1848 vdd.n1101 0.152939
R22705 vdd.n1862 vdd.n1101 0.152939
R22706 vdd.n1863 vdd.n1862 0.152939
R22707 vdd.n1864 vdd.n1863 0.152939
R22708 vdd.n1864 vdd.n1089 0.152939
R22709 vdd.n1879 vdd.n1089 0.152939
R22710 vdd.n1880 vdd.n1879 0.152939
R22711 vdd.n1881 vdd.n1880 0.152939
R22712 vdd.n1881 vdd.n1077 0.152939
R22713 vdd.n1898 vdd.n1077 0.152939
R22714 vdd.n1899 vdd.n1898 0.152939
R22715 vdd.n2326 vdd.n1899 0.152939
R22716 vdd.n735 vdd.n730 0.152939
R22717 vdd.n736 vdd.n735 0.152939
R22718 vdd.n737 vdd.n736 0.152939
R22719 vdd.n738 vdd.n737 0.152939
R22720 vdd.n739 vdd.n738 0.152939
R22721 vdd.n740 vdd.n739 0.152939
R22722 vdd.n741 vdd.n740 0.152939
R22723 vdd.n742 vdd.n741 0.152939
R22724 vdd.n743 vdd.n742 0.152939
R22725 vdd.n744 vdd.n743 0.152939
R22726 vdd.n745 vdd.n744 0.152939
R22727 vdd.n746 vdd.n745 0.152939
R22728 vdd.n3183 vdd.n746 0.152939
R22729 vdd.n3183 vdd.n3182 0.152939
R22730 vdd.n3182 vdd.n3181 0.152939
R22731 vdd.n3181 vdd.n748 0.152939
R22732 vdd.n749 vdd.n748 0.152939
R22733 vdd.n750 vdd.n749 0.152939
R22734 vdd.n751 vdd.n750 0.152939
R22735 vdd.n752 vdd.n751 0.152939
R22736 vdd.n753 vdd.n752 0.152939
R22737 vdd.n754 vdd.n753 0.152939
R22738 vdd.n755 vdd.n754 0.152939
R22739 vdd.n756 vdd.n755 0.152939
R22740 vdd.n757 vdd.n756 0.152939
R22741 vdd.n758 vdd.n757 0.152939
R22742 vdd.n759 vdd.n758 0.152939
R22743 vdd.n760 vdd.n759 0.152939
R22744 vdd.n761 vdd.n760 0.152939
R22745 vdd.n762 vdd.n761 0.152939
R22746 vdd.n763 vdd.n762 0.152939
R22747 vdd.n764 vdd.n763 0.152939
R22748 vdd.n765 vdd.n764 0.152939
R22749 vdd.n766 vdd.n765 0.152939
R22750 vdd.n3137 vdd.n766 0.152939
R22751 vdd.n3137 vdd.n3136 0.152939
R22752 vdd.n3136 vdd.n3135 0.152939
R22753 vdd.n3135 vdd.n770 0.152939
R22754 vdd.n771 vdd.n770 0.152939
R22755 vdd.n772 vdd.n771 0.152939
R22756 vdd.n773 vdd.n772 0.152939
R22757 vdd.n774 vdd.n773 0.152939
R22758 vdd.n775 vdd.n774 0.152939
R22759 vdd.n776 vdd.n775 0.152939
R22760 vdd.n777 vdd.n776 0.152939
R22761 vdd.n778 vdd.n777 0.152939
R22762 vdd.n779 vdd.n778 0.152939
R22763 vdd.n780 vdd.n779 0.152939
R22764 vdd.n781 vdd.n780 0.152939
R22765 vdd.n782 vdd.n781 0.152939
R22766 vdd.n783 vdd.n782 0.152939
R22767 vdd.n727 vdd.n726 0.152939
R22768 vdd.n3234 vdd.n682 0.152939
R22769 vdd.n3235 vdd.n3234 0.152939
R22770 vdd.n3236 vdd.n3235 0.152939
R22771 vdd.n3236 vdd.n670 0.152939
R22772 vdd.n3251 vdd.n670 0.152939
R22773 vdd.n3252 vdd.n3251 0.152939
R22774 vdd.n3253 vdd.n3252 0.152939
R22775 vdd.n3253 vdd.n659 0.152939
R22776 vdd.n3267 vdd.n659 0.152939
R22777 vdd.n3268 vdd.n3267 0.152939
R22778 vdd.n3269 vdd.n3268 0.152939
R22779 vdd.n3269 vdd.n647 0.152939
R22780 vdd.n3284 vdd.n647 0.152939
R22781 vdd.n3285 vdd.n3284 0.152939
R22782 vdd.n3286 vdd.n3285 0.152939
R22783 vdd.n3286 vdd.n636 0.152939
R22784 vdd.n3303 vdd.n636 0.152939
R22785 vdd.n3304 vdd.n3303 0.152939
R22786 vdd.n3305 vdd.n3304 0.152939
R22787 vdd.n3305 vdd.n334 0.152939
R22788 vdd.n3398 vdd.n335 0.152939
R22789 vdd.n346 vdd.n335 0.152939
R22790 vdd.n347 vdd.n346 0.152939
R22791 vdd.n348 vdd.n347 0.152939
R22792 vdd.n355 vdd.n348 0.152939
R22793 vdd.n356 vdd.n355 0.152939
R22794 vdd.n357 vdd.n356 0.152939
R22795 vdd.n358 vdd.n357 0.152939
R22796 vdd.n366 vdd.n358 0.152939
R22797 vdd.n367 vdd.n366 0.152939
R22798 vdd.n368 vdd.n367 0.152939
R22799 vdd.n369 vdd.n368 0.152939
R22800 vdd.n377 vdd.n369 0.152939
R22801 vdd.n378 vdd.n377 0.152939
R22802 vdd.n379 vdd.n378 0.152939
R22803 vdd.n380 vdd.n379 0.152939
R22804 vdd.n388 vdd.n380 0.152939
R22805 vdd.n389 vdd.n388 0.152939
R22806 vdd.n390 vdd.n389 0.152939
R22807 vdd.n391 vdd.n390 0.152939
R22808 vdd.n464 vdd.n463 0.152939
R22809 vdd.n470 vdd.n463 0.152939
R22810 vdd.n471 vdd.n470 0.152939
R22811 vdd.n472 vdd.n471 0.152939
R22812 vdd.n472 vdd.n461 0.152939
R22813 vdd.n480 vdd.n461 0.152939
R22814 vdd.n481 vdd.n480 0.152939
R22815 vdd.n482 vdd.n481 0.152939
R22816 vdd.n482 vdd.n459 0.152939
R22817 vdd.n490 vdd.n459 0.152939
R22818 vdd.n491 vdd.n490 0.152939
R22819 vdd.n492 vdd.n491 0.152939
R22820 vdd.n492 vdd.n457 0.152939
R22821 vdd.n500 vdd.n457 0.152939
R22822 vdd.n501 vdd.n500 0.152939
R22823 vdd.n502 vdd.n501 0.152939
R22824 vdd.n502 vdd.n455 0.152939
R22825 vdd.n510 vdd.n455 0.152939
R22826 vdd.n511 vdd.n510 0.152939
R22827 vdd.n512 vdd.n511 0.152939
R22828 vdd.n512 vdd.n451 0.152939
R22829 vdd.n520 vdd.n451 0.152939
R22830 vdd.n521 vdd.n520 0.152939
R22831 vdd.n522 vdd.n521 0.152939
R22832 vdd.n522 vdd.n449 0.152939
R22833 vdd.n530 vdd.n449 0.152939
R22834 vdd.n531 vdd.n530 0.152939
R22835 vdd.n532 vdd.n531 0.152939
R22836 vdd.n532 vdd.n447 0.152939
R22837 vdd.n540 vdd.n447 0.152939
R22838 vdd.n541 vdd.n540 0.152939
R22839 vdd.n542 vdd.n541 0.152939
R22840 vdd.n542 vdd.n445 0.152939
R22841 vdd.n550 vdd.n445 0.152939
R22842 vdd.n551 vdd.n550 0.152939
R22843 vdd.n552 vdd.n551 0.152939
R22844 vdd.n552 vdd.n443 0.152939
R22845 vdd.n560 vdd.n443 0.152939
R22846 vdd.n561 vdd.n560 0.152939
R22847 vdd.n562 vdd.n561 0.152939
R22848 vdd.n562 vdd.n439 0.152939
R22849 vdd.n570 vdd.n439 0.152939
R22850 vdd.n571 vdd.n570 0.152939
R22851 vdd.n572 vdd.n571 0.152939
R22852 vdd.n572 vdd.n437 0.152939
R22853 vdd.n580 vdd.n437 0.152939
R22854 vdd.n581 vdd.n580 0.152939
R22855 vdd.n582 vdd.n581 0.152939
R22856 vdd.n582 vdd.n435 0.152939
R22857 vdd.n590 vdd.n435 0.152939
R22858 vdd.n591 vdd.n590 0.152939
R22859 vdd.n592 vdd.n591 0.152939
R22860 vdd.n592 vdd.n433 0.152939
R22861 vdd.n600 vdd.n433 0.152939
R22862 vdd.n601 vdd.n600 0.152939
R22863 vdd.n602 vdd.n601 0.152939
R22864 vdd.n602 vdd.n431 0.152939
R22865 vdd.n610 vdd.n431 0.152939
R22866 vdd.n611 vdd.n610 0.152939
R22867 vdd.n612 vdd.n611 0.152939
R22868 vdd.n612 vdd.n429 0.152939
R22869 vdd.n619 vdd.n429 0.152939
R22870 vdd.n3350 vdd.n619 0.152939
R22871 vdd.n3228 vdd.n3227 0.152939
R22872 vdd.n3228 vdd.n675 0.152939
R22873 vdd.n3242 vdd.n675 0.152939
R22874 vdd.n3243 vdd.n3242 0.152939
R22875 vdd.n3244 vdd.n3243 0.152939
R22876 vdd.n3244 vdd.n665 0.152939
R22877 vdd.n3259 vdd.n665 0.152939
R22878 vdd.n3260 vdd.n3259 0.152939
R22879 vdd.n3261 vdd.n3260 0.152939
R22880 vdd.n3261 vdd.n652 0.152939
R22881 vdd.n3275 vdd.n652 0.152939
R22882 vdd.n3276 vdd.n3275 0.152939
R22883 vdd.n3277 vdd.n3276 0.152939
R22884 vdd.n3277 vdd.n641 0.152939
R22885 vdd.n3292 vdd.n641 0.152939
R22886 vdd.n3293 vdd.n3292 0.152939
R22887 vdd.n3294 vdd.n3293 0.152939
R22888 vdd.n3296 vdd.n3294 0.152939
R22889 vdd.n3296 vdd.n3295 0.152939
R22890 vdd.n3295 vdd.n630 0.152939
R22891 vdd.n3313 vdd.n630 0.152939
R22892 vdd.n3314 vdd.n3313 0.152939
R22893 vdd.n3315 vdd.n3314 0.152939
R22894 vdd.n3315 vdd.n628 0.152939
R22895 vdd.n3320 vdd.n628 0.152939
R22896 vdd.n3321 vdd.n3320 0.152939
R22897 vdd.n3322 vdd.n3321 0.152939
R22898 vdd.n3322 vdd.n626 0.152939
R22899 vdd.n3327 vdd.n626 0.152939
R22900 vdd.n3328 vdd.n3327 0.152939
R22901 vdd.n3329 vdd.n3328 0.152939
R22902 vdd.n3329 vdd.n624 0.152939
R22903 vdd.n3335 vdd.n624 0.152939
R22904 vdd.n3336 vdd.n3335 0.152939
R22905 vdd.n3337 vdd.n3336 0.152939
R22906 vdd.n3337 vdd.n622 0.152939
R22907 vdd.n3342 vdd.n622 0.152939
R22908 vdd.n3343 vdd.n3342 0.152939
R22909 vdd.n3344 vdd.n3343 0.152939
R22910 vdd.n3344 vdd.n620 0.152939
R22911 vdd.n3349 vdd.n620 0.152939
R22912 vdd.n3226 vdd.n687 0.152939
R22913 vdd.n2337 vdd.n1067 0.152939
R22914 vdd.n1430 vdd.n1186 0.152939
R22915 vdd.n1431 vdd.n1430 0.152939
R22916 vdd.n1432 vdd.n1431 0.152939
R22917 vdd.n1432 vdd.n1174 0.152939
R22918 vdd.n1447 vdd.n1174 0.152939
R22919 vdd.n1448 vdd.n1447 0.152939
R22920 vdd.n1449 vdd.n1448 0.152939
R22921 vdd.n1449 vdd.n1164 0.152939
R22922 vdd.n1464 vdd.n1164 0.152939
R22923 vdd.n1465 vdd.n1464 0.152939
R22924 vdd.n1466 vdd.n1465 0.152939
R22925 vdd.n1466 vdd.n1151 0.152939
R22926 vdd.n1480 vdd.n1151 0.152939
R22927 vdd.n1481 vdd.n1480 0.152939
R22928 vdd.n1482 vdd.n1481 0.152939
R22929 vdd.n1482 vdd.n1140 0.152939
R22930 vdd.n1497 vdd.n1140 0.152939
R22931 vdd.n1498 vdd.n1497 0.152939
R22932 vdd.n1499 vdd.n1498 0.152939
R22933 vdd.n1499 vdd.n1129 0.152939
R22934 vdd.n1820 vdd.n1129 0.152939
R22935 vdd.n1821 vdd.n1820 0.152939
R22936 vdd.n1822 vdd.n1821 0.152939
R22937 vdd.n1822 vdd.n1117 0.152939
R22938 vdd.n1837 vdd.n1117 0.152939
R22939 vdd.n1838 vdd.n1837 0.152939
R22940 vdd.n1839 vdd.n1838 0.152939
R22941 vdd.n1839 vdd.n1107 0.152939
R22942 vdd.n1854 vdd.n1107 0.152939
R22943 vdd.n1855 vdd.n1854 0.152939
R22944 vdd.n1856 vdd.n1855 0.152939
R22945 vdd.n1856 vdd.n1094 0.152939
R22946 vdd.n1870 vdd.n1094 0.152939
R22947 vdd.n1871 vdd.n1870 0.152939
R22948 vdd.n1872 vdd.n1871 0.152939
R22949 vdd.n1872 vdd.n1084 0.152939
R22950 vdd.n1887 vdd.n1084 0.152939
R22951 vdd.n1888 vdd.n1887 0.152939
R22952 vdd.n1891 vdd.n1888 0.152939
R22953 vdd.n1891 vdd.n1890 0.152939
R22954 vdd.n1890 vdd.n1889 0.152939
R22955 vdd.n1422 vdd.n1191 0.152939
R22956 vdd.n1415 vdd.n1191 0.152939
R22957 vdd.n1415 vdd.n1414 0.152939
R22958 vdd.n1414 vdd.n1413 0.152939
R22959 vdd.n1413 vdd.n1228 0.152939
R22960 vdd.n1409 vdd.n1228 0.152939
R22961 vdd.n1409 vdd.n1408 0.152939
R22962 vdd.n1408 vdd.n1407 0.152939
R22963 vdd.n1407 vdd.n1234 0.152939
R22964 vdd.n1403 vdd.n1234 0.152939
R22965 vdd.n1403 vdd.n1402 0.152939
R22966 vdd.n1402 vdd.n1401 0.152939
R22967 vdd.n1401 vdd.n1240 0.152939
R22968 vdd.n1397 vdd.n1240 0.152939
R22969 vdd.n1397 vdd.n1396 0.152939
R22970 vdd.n1396 vdd.n1395 0.152939
R22971 vdd.n1395 vdd.n1246 0.152939
R22972 vdd.n1391 vdd.n1246 0.152939
R22973 vdd.n1391 vdd.n1390 0.152939
R22974 vdd.n1390 vdd.n1389 0.152939
R22975 vdd.n1389 vdd.n1254 0.152939
R22976 vdd.n1385 vdd.n1254 0.152939
R22977 vdd.n1385 vdd.n1384 0.152939
R22978 vdd.n1384 vdd.n1383 0.152939
R22979 vdd.n1383 vdd.n1260 0.152939
R22980 vdd.n1379 vdd.n1260 0.152939
R22981 vdd.n1379 vdd.n1378 0.152939
R22982 vdd.n1378 vdd.n1377 0.152939
R22983 vdd.n1377 vdd.n1266 0.152939
R22984 vdd.n1373 vdd.n1266 0.152939
R22985 vdd.n1373 vdd.n1372 0.152939
R22986 vdd.n1372 vdd.n1371 0.152939
R22987 vdd.n1371 vdd.n1272 0.152939
R22988 vdd.n1367 vdd.n1272 0.152939
R22989 vdd.n1367 vdd.n1366 0.152939
R22990 vdd.n1366 vdd.n1365 0.152939
R22991 vdd.n1365 vdd.n1278 0.152939
R22992 vdd.n1361 vdd.n1278 0.152939
R22993 vdd.n1361 vdd.n1360 0.152939
R22994 vdd.n1360 vdd.n1359 0.152939
R22995 vdd.n1359 vdd.n1284 0.152939
R22996 vdd.n1352 vdd.n1284 0.152939
R22997 vdd.n1352 vdd.n1351 0.152939
R22998 vdd.n1351 vdd.n1350 0.152939
R22999 vdd.n1350 vdd.n1289 0.152939
R23000 vdd.n1346 vdd.n1289 0.152939
R23001 vdd.n1346 vdd.n1345 0.152939
R23002 vdd.n1345 vdd.n1344 0.152939
R23003 vdd.n1344 vdd.n1295 0.152939
R23004 vdd.n1340 vdd.n1295 0.152939
R23005 vdd.n1340 vdd.n1339 0.152939
R23006 vdd.n1339 vdd.n1338 0.152939
R23007 vdd.n1338 vdd.n1301 0.152939
R23008 vdd.n1334 vdd.n1301 0.152939
R23009 vdd.n1334 vdd.n1333 0.152939
R23010 vdd.n1333 vdd.n1332 0.152939
R23011 vdd.n1332 vdd.n1307 0.152939
R23012 vdd.n1328 vdd.n1307 0.152939
R23013 vdd.n1328 vdd.n1327 0.152939
R23014 vdd.n1327 vdd.n1326 0.152939
R23015 vdd.n1326 vdd.n1313 0.152939
R23016 vdd.n1322 vdd.n1313 0.152939
R23017 vdd.n1322 vdd.n1321 0.152939
R23018 vdd.n1424 vdd.n1423 0.152939
R23019 vdd.n1424 vdd.n1180 0.152939
R23020 vdd.n1439 vdd.n1180 0.152939
R23021 vdd.n1440 vdd.n1439 0.152939
R23022 vdd.n1441 vdd.n1440 0.152939
R23023 vdd.n1441 vdd.n1169 0.152939
R23024 vdd.n1456 vdd.n1169 0.152939
R23025 vdd.n1457 vdd.n1456 0.152939
R23026 vdd.n1458 vdd.n1457 0.152939
R23027 vdd.n1458 vdd.n1158 0.152939
R23028 vdd.n1472 vdd.n1158 0.152939
R23029 vdd.n1473 vdd.n1472 0.152939
R23030 vdd.n1474 vdd.n1473 0.152939
R23031 vdd.n1474 vdd.n1146 0.152939
R23032 vdd.n1489 vdd.n1146 0.152939
R23033 vdd.n1490 vdd.n1489 0.152939
R23034 vdd.n1491 vdd.n1490 0.152939
R23035 vdd.n1491 vdd.n1135 0.152939
R23036 vdd.n1505 vdd.n1135 0.152939
R23037 vdd.n1506 vdd.n1505 0.152939
R23038 vdd.n1427 vdd.t185 0.113865
R23039 vdd.t192 vdd.n386 0.113865
R23040 vdd.n2315 vdd.n1900 0.110256
R23041 vdd.n3216 vdd.n727 0.110256
R23042 vdd.n3093 vdd.n687 0.110256
R23043 vdd.n2338 vdd.n2337 0.110256
R23044 vdd.n1814 vdd.n1813 0.0695946
R23045 vdd.n3399 vdd.n334 0.0695946
R23046 vdd.n3399 vdd.n3398 0.0695946
R23047 vdd.n1813 vdd.n1506 0.0695946
R23048 vdd.n2315 vdd.n2101 0.0431829
R23049 vdd.n2338 vdd.n1064 0.0431829
R23050 vdd.n3216 vdd.n730 0.0431829
R23051 vdd.n3093 vdd.n783 0.0431829
R23052 vdd vdd.n28 0.00833333
R23053 a_n1986_8322.n14 a_n1986_8322.t12 74.6477
R23054 a_n1986_8322.n7 a_n1986_8322.t6 74.6477
R23055 a_n1986_8322.n1 a_n1986_8322.t3 74.6474
R23056 a_n1986_8322.n15 a_n1986_8322.t10 74.2899
R23057 a_n1986_8322.n16 a_n1986_8322.t13 74.2899
R23058 a_n1986_8322.n12 a_n1986_8322.t14 74.2899
R23059 a_n1986_8322.n4 a_n1986_8322.t19 74.2899
R23060 a_n1986_8322.n10 a_n1986_8322.t18 74.2899
R23061 a_n1986_8322.n14 a_n1986_8322.n13 70.6783
R23062 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R23063 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R23064 a_n1986_8322.n7 a_n1986_8322.n6 70.6783
R23065 a_n1986_8322.n9 a_n1986_8322.n8 70.6783
R23066 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R23067 a_n1986_8322.n11 a_n1986_8322.n10 22.7556
R23068 a_n1986_8322.n5 a_n1986_8322.t0 10.1306
R23069 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R23070 a_n1986_8322.n5 a_n1986_8322.n4 5.83671
R23071 a_n1986_8322.n11 a_n1986_8322.n5 5.3452
R23072 a_n1986_8322.n13 a_n1986_8322.t16 3.61217
R23073 a_n1986_8322.n13 a_n1986_8322.t15 3.61217
R23074 a_n1986_8322.n0 a_n1986_8322.t5 3.61217
R23075 a_n1986_8322.n0 a_n1986_8322.t8 3.61217
R23076 a_n1986_8322.n2 a_n1986_8322.t7 3.61217
R23077 a_n1986_8322.n2 a_n1986_8322.t1 3.61217
R23078 a_n1986_8322.n6 a_n1986_8322.t2 3.61217
R23079 a_n1986_8322.n6 a_n1986_8322.t20 3.61217
R23080 a_n1986_8322.n8 a_n1986_8322.t4 3.61217
R23081 a_n1986_8322.n8 a_n1986_8322.t9 3.61217
R23082 a_n1986_8322.n18 a_n1986_8322.t11 3.61217
R23083 a_n1986_8322.t17 a_n1986_8322.n18 3.61217
R23084 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R23085 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R23086 a_n1986_8322.n10 a_n1986_8322.n9 0.358259
R23087 a_n1986_8322.n9 a_n1986_8322.n7 0.358259
R23088 a_n1986_8322.n17 a_n1986_8322.n12 0.358259
R23089 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R23090 a_n1986_8322.n15 a_n1986_8322.n14 0.358259
R23091 a_n1986_8322.n16 a_n1986_8322.n15 0.101793
R23092 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R23093 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R23094 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R23095 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R23096 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R23097 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R23098 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R23099 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R23100 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R23101 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R23102 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R23103 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R23104 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R23105 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R23106 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R23107 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R23108 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R23109 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R23110 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R23111 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R23112 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R23113 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R23114 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R23115 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R23116 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R23117 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R23118 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R23119 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R23120 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R23121 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R23122 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R23123 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R23124 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R23125 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R23126 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R23127 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R23128 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R23129 a_n7636_8799.n225 a_n7636_8799.t57 485.149
R23130 a_n7636_8799.n287 a_n7636_8799.t68 485.149
R23131 a_n7636_8799.n350 a_n7636_8799.t106 485.149
R23132 a_n7636_8799.n35 a_n7636_8799.t129 485.149
R23133 a_n7636_8799.n97 a_n7636_8799.t143 485.149
R23134 a_n7636_8799.n160 a_n7636_8799.t105 485.149
R23135 a_n7636_8799.n268 a_n7636_8799.t79 464.166
R23136 a_n7636_8799.n267 a_n7636_8799.t78 464.166
R23137 a_n7636_8799.n209 a_n7636_8799.t51 464.166
R23138 a_n7636_8799.n261 a_n7636_8799.t127 464.166
R23139 a_n7636_8799.n260 a_n7636_8799.t82 464.166
R23140 a_n7636_8799.n212 a_n7636_8799.t58 464.166
R23141 a_n7636_8799.n254 a_n7636_8799.t133 464.166
R23142 a_n7636_8799.n253 a_n7636_8799.t99 464.166
R23143 a_n7636_8799.n215 a_n7636_8799.t97 464.166
R23144 a_n7636_8799.n247 a_n7636_8799.t32 464.166
R23145 a_n7636_8799.n246 a_n7636_8799.t103 464.166
R23146 a_n7636_8799.n218 a_n7636_8799.t102 464.166
R23147 a_n7636_8799.n240 a_n7636_8799.t34 464.166
R23148 a_n7636_8799.n239 a_n7636_8799.t33 464.166
R23149 a_n7636_8799.n221 a_n7636_8799.t119 464.166
R23150 a_n7636_8799.n233 a_n7636_8799.t53 464.166
R23151 a_n7636_8799.n232 a_n7636_8799.t36 464.166
R23152 a_n7636_8799.n224 a_n7636_8799.t123 464.166
R23153 a_n7636_8799.n226 a_n7636_8799.t81 464.166
R23154 a_n7636_8799.n330 a_n7636_8799.t89 464.166
R23155 a_n7636_8799.n329 a_n7636_8799.t88 464.166
R23156 a_n7636_8799.n271 a_n7636_8799.t66 464.166
R23157 a_n7636_8799.n323 a_n7636_8799.t142 464.166
R23158 a_n7636_8799.n322 a_n7636_8799.t96 464.166
R23159 a_n7636_8799.n274 a_n7636_8799.t69 464.166
R23160 a_n7636_8799.n316 a_n7636_8799.t28 464.166
R23161 a_n7636_8799.n315 a_n7636_8799.t112 464.166
R23162 a_n7636_8799.n277 a_n7636_8799.t111 464.166
R23163 a_n7636_8799.n309 a_n7636_8799.t42 464.166
R23164 a_n7636_8799.n308 a_n7636_8799.t115 464.166
R23165 a_n7636_8799.n280 a_n7636_8799.t114 464.166
R23166 a_n7636_8799.n302 a_n7636_8799.t46 464.166
R23167 a_n7636_8799.n301 a_n7636_8799.t45 464.166
R23168 a_n7636_8799.n283 a_n7636_8799.t136 464.166
R23169 a_n7636_8799.n295 a_n7636_8799.t67 464.166
R23170 a_n7636_8799.n294 a_n7636_8799.t48 464.166
R23171 a_n7636_8799.n286 a_n7636_8799.t137 464.166
R23172 a_n7636_8799.n288 a_n7636_8799.t95 464.166
R23173 a_n7636_8799.n393 a_n7636_8799.t146 464.166
R23174 a_n7636_8799.n392 a_n7636_8799.t44 464.166
R23175 a_n7636_8799.n334 a_n7636_8799.t94 464.166
R23176 a_n7636_8799.n386 a_n7636_8799.t31 464.166
R23177 a_n7636_8799.n385 a_n7636_8799.t118 464.166
R23178 a_n7636_8799.n337 a_n7636_8799.t55 464.166
R23179 a_n7636_8799.n379 a_n7636_8799.t101 464.166
R23180 a_n7636_8799.n378 a_n7636_8799.t37 464.166
R23181 a_n7636_8799.n340 a_n7636_8799.t61 464.166
R23182 a_n7636_8799.n372 a_n7636_8799.t141 464.166
R23183 a_n7636_8799.n371 a_n7636_8799.t110 464.166
R23184 a_n7636_8799.n343 a_n7636_8799.t135 464.166
R23185 a_n7636_8799.n365 a_n7636_8799.t92 464.166
R23186 a_n7636_8799.n364 a_n7636_8799.t113 464.166
R23187 a_n7636_8799.n346 a_n7636_8799.t49 464.166
R23188 a_n7636_8799.n358 a_n7636_8799.t132 464.166
R23189 a_n7636_8799.n357 a_n7636_8799.t73 464.166
R23190 a_n7636_8799.n349 a_n7636_8799.t124 464.166
R23191 a_n7636_8799.n351 a_n7636_8799.t60 464.166
R23192 a_n7636_8799.n36 a_n7636_8799.t130 464.166
R23193 a_n7636_8799.n38 a_n7636_8799.t80 464.166
R23194 a_n7636_8799.n42 a_n7636_8799.t109 464.166
R23195 a_n7636_8799.n43 a_n7636_8799.t126 464.166
R23196 a_n7636_8799.n31 a_n7636_8799.t76 464.166
R23197 a_n7636_8799.n49 a_n7636_8799.t77 464.166
R23198 a_n7636_8799.n50 a_n7636_8799.t107 464.166
R23199 a_n7636_8799.n54 a_n7636_8799.t64 464.166
R23200 a_n7636_8799.n56 a_n7636_8799.t65 464.166
R23201 a_n7636_8799.n27 a_n7636_8799.t104 464.166
R23202 a_n7636_8799.n61 a_n7636_8799.t29 464.166
R23203 a_n7636_8799.n25 a_n7636_8799.t62 464.166
R23204 a_n7636_8799.n66 a_n7636_8799.t85 464.166
R23205 a_n7636_8799.n68 a_n7636_8799.t128 464.166
R23206 a_n7636_8799.n72 a_n7636_8799.t41 464.166
R23207 a_n7636_8799.n73 a_n7636_8799.t59 464.166
R23208 a_n7636_8799.n21 a_n7636_8799.t125 464.166
R23209 a_n7636_8799.n79 a_n7636_8799.t38 464.166
R23210 a_n7636_8799.n80 a_n7636_8799.t39 464.166
R23211 a_n7636_8799.n98 a_n7636_8799.t147 464.166
R23212 a_n7636_8799.n100 a_n7636_8799.t90 464.166
R23213 a_n7636_8799.n104 a_n7636_8799.t122 464.166
R23214 a_n7636_8799.n105 a_n7636_8799.t140 464.166
R23215 a_n7636_8799.n93 a_n7636_8799.t86 464.166
R23216 a_n7636_8799.n111 a_n7636_8799.t87 464.166
R23217 a_n7636_8799.n112 a_n7636_8799.t120 464.166
R23218 a_n7636_8799.n116 a_n7636_8799.t74 464.166
R23219 a_n7636_8799.n118 a_n7636_8799.t75 464.166
R23220 a_n7636_8799.n89 a_n7636_8799.t116 464.166
R23221 a_n7636_8799.n123 a_n7636_8799.t40 464.166
R23222 a_n7636_8799.n87 a_n7636_8799.t71 464.166
R23223 a_n7636_8799.n128 a_n7636_8799.t98 464.166
R23224 a_n7636_8799.n130 a_n7636_8799.t144 464.166
R23225 a_n7636_8799.n134 a_n7636_8799.t56 464.166
R23226 a_n7636_8799.n135 a_n7636_8799.t70 464.166
R23227 a_n7636_8799.n83 a_n7636_8799.t138 464.166
R23228 a_n7636_8799.n141 a_n7636_8799.t50 464.166
R23229 a_n7636_8799.n142 a_n7636_8799.t52 464.166
R23230 a_n7636_8799.n161 a_n7636_8799.t83 464.166
R23231 a_n7636_8799.n163 a_n7636_8799.t121 464.166
R23232 a_n7636_8799.n167 a_n7636_8799.t72 464.166
R23233 a_n7636_8799.n168 a_n7636_8799.t131 464.166
R23234 a_n7636_8799.n156 a_n7636_8799.t47 464.166
R23235 a_n7636_8799.n174 a_n7636_8799.t30 464.166
R23236 a_n7636_8799.n175 a_n7636_8799.t91 464.166
R23237 a_n7636_8799.n179 a_n7636_8799.t134 464.166
R23238 a_n7636_8799.n181 a_n7636_8799.t108 464.166
R23239 a_n7636_8799.n152 a_n7636_8799.t139 464.166
R23240 a_n7636_8799.n186 a_n7636_8799.t84 464.166
R23241 a_n7636_8799.n150 a_n7636_8799.t35 464.166
R23242 a_n7636_8799.n191 a_n7636_8799.t100 464.166
R23243 a_n7636_8799.n193 a_n7636_8799.t54 464.166
R23244 a_n7636_8799.n197 a_n7636_8799.t117 464.166
R23245 a_n7636_8799.n198 a_n7636_8799.t63 464.166
R23246 a_n7636_8799.n146 a_n7636_8799.t93 464.166
R23247 a_n7636_8799.n204 a_n7636_8799.t43 464.166
R23248 a_n7636_8799.n205 a_n7636_8799.t145 464.166
R23249 a_n7636_8799.n228 a_n7636_8799.n227 161.3
R23250 a_n7636_8799.n229 a_n7636_8799.n224 161.3
R23251 a_n7636_8799.n231 a_n7636_8799.n230 161.3
R23252 a_n7636_8799.n232 a_n7636_8799.n223 161.3
R23253 a_n7636_8799.n233 a_n7636_8799.n222 161.3
R23254 a_n7636_8799.n235 a_n7636_8799.n234 161.3
R23255 a_n7636_8799.n236 a_n7636_8799.n221 161.3
R23256 a_n7636_8799.n238 a_n7636_8799.n237 161.3
R23257 a_n7636_8799.n239 a_n7636_8799.n220 161.3
R23258 a_n7636_8799.n240 a_n7636_8799.n219 161.3
R23259 a_n7636_8799.n242 a_n7636_8799.n241 161.3
R23260 a_n7636_8799.n243 a_n7636_8799.n218 161.3
R23261 a_n7636_8799.n245 a_n7636_8799.n244 161.3
R23262 a_n7636_8799.n246 a_n7636_8799.n217 161.3
R23263 a_n7636_8799.n247 a_n7636_8799.n216 161.3
R23264 a_n7636_8799.n249 a_n7636_8799.n248 161.3
R23265 a_n7636_8799.n250 a_n7636_8799.n215 161.3
R23266 a_n7636_8799.n252 a_n7636_8799.n251 161.3
R23267 a_n7636_8799.n253 a_n7636_8799.n214 161.3
R23268 a_n7636_8799.n254 a_n7636_8799.n213 161.3
R23269 a_n7636_8799.n256 a_n7636_8799.n255 161.3
R23270 a_n7636_8799.n257 a_n7636_8799.n212 161.3
R23271 a_n7636_8799.n259 a_n7636_8799.n258 161.3
R23272 a_n7636_8799.n260 a_n7636_8799.n211 161.3
R23273 a_n7636_8799.n261 a_n7636_8799.n210 161.3
R23274 a_n7636_8799.n263 a_n7636_8799.n262 161.3
R23275 a_n7636_8799.n264 a_n7636_8799.n209 161.3
R23276 a_n7636_8799.n266 a_n7636_8799.n265 161.3
R23277 a_n7636_8799.n267 a_n7636_8799.n208 161.3
R23278 a_n7636_8799.n269 a_n7636_8799.n268 161.3
R23279 a_n7636_8799.n290 a_n7636_8799.n289 161.3
R23280 a_n7636_8799.n291 a_n7636_8799.n286 161.3
R23281 a_n7636_8799.n293 a_n7636_8799.n292 161.3
R23282 a_n7636_8799.n294 a_n7636_8799.n285 161.3
R23283 a_n7636_8799.n295 a_n7636_8799.n284 161.3
R23284 a_n7636_8799.n297 a_n7636_8799.n296 161.3
R23285 a_n7636_8799.n298 a_n7636_8799.n283 161.3
R23286 a_n7636_8799.n300 a_n7636_8799.n299 161.3
R23287 a_n7636_8799.n301 a_n7636_8799.n282 161.3
R23288 a_n7636_8799.n302 a_n7636_8799.n281 161.3
R23289 a_n7636_8799.n304 a_n7636_8799.n303 161.3
R23290 a_n7636_8799.n305 a_n7636_8799.n280 161.3
R23291 a_n7636_8799.n307 a_n7636_8799.n306 161.3
R23292 a_n7636_8799.n308 a_n7636_8799.n279 161.3
R23293 a_n7636_8799.n309 a_n7636_8799.n278 161.3
R23294 a_n7636_8799.n311 a_n7636_8799.n310 161.3
R23295 a_n7636_8799.n312 a_n7636_8799.n277 161.3
R23296 a_n7636_8799.n314 a_n7636_8799.n313 161.3
R23297 a_n7636_8799.n315 a_n7636_8799.n276 161.3
R23298 a_n7636_8799.n316 a_n7636_8799.n275 161.3
R23299 a_n7636_8799.n318 a_n7636_8799.n317 161.3
R23300 a_n7636_8799.n319 a_n7636_8799.n274 161.3
R23301 a_n7636_8799.n321 a_n7636_8799.n320 161.3
R23302 a_n7636_8799.n322 a_n7636_8799.n273 161.3
R23303 a_n7636_8799.n323 a_n7636_8799.n272 161.3
R23304 a_n7636_8799.n325 a_n7636_8799.n324 161.3
R23305 a_n7636_8799.n326 a_n7636_8799.n271 161.3
R23306 a_n7636_8799.n328 a_n7636_8799.n327 161.3
R23307 a_n7636_8799.n329 a_n7636_8799.n270 161.3
R23308 a_n7636_8799.n331 a_n7636_8799.n330 161.3
R23309 a_n7636_8799.n353 a_n7636_8799.n352 161.3
R23310 a_n7636_8799.n354 a_n7636_8799.n349 161.3
R23311 a_n7636_8799.n356 a_n7636_8799.n355 161.3
R23312 a_n7636_8799.n357 a_n7636_8799.n348 161.3
R23313 a_n7636_8799.n358 a_n7636_8799.n347 161.3
R23314 a_n7636_8799.n360 a_n7636_8799.n359 161.3
R23315 a_n7636_8799.n361 a_n7636_8799.n346 161.3
R23316 a_n7636_8799.n363 a_n7636_8799.n362 161.3
R23317 a_n7636_8799.n364 a_n7636_8799.n345 161.3
R23318 a_n7636_8799.n365 a_n7636_8799.n344 161.3
R23319 a_n7636_8799.n367 a_n7636_8799.n366 161.3
R23320 a_n7636_8799.n368 a_n7636_8799.n343 161.3
R23321 a_n7636_8799.n370 a_n7636_8799.n369 161.3
R23322 a_n7636_8799.n371 a_n7636_8799.n342 161.3
R23323 a_n7636_8799.n372 a_n7636_8799.n341 161.3
R23324 a_n7636_8799.n374 a_n7636_8799.n373 161.3
R23325 a_n7636_8799.n375 a_n7636_8799.n340 161.3
R23326 a_n7636_8799.n377 a_n7636_8799.n376 161.3
R23327 a_n7636_8799.n378 a_n7636_8799.n339 161.3
R23328 a_n7636_8799.n379 a_n7636_8799.n338 161.3
R23329 a_n7636_8799.n381 a_n7636_8799.n380 161.3
R23330 a_n7636_8799.n382 a_n7636_8799.n337 161.3
R23331 a_n7636_8799.n384 a_n7636_8799.n383 161.3
R23332 a_n7636_8799.n385 a_n7636_8799.n336 161.3
R23333 a_n7636_8799.n386 a_n7636_8799.n335 161.3
R23334 a_n7636_8799.n388 a_n7636_8799.n387 161.3
R23335 a_n7636_8799.n389 a_n7636_8799.n334 161.3
R23336 a_n7636_8799.n391 a_n7636_8799.n390 161.3
R23337 a_n7636_8799.n392 a_n7636_8799.n333 161.3
R23338 a_n7636_8799.n394 a_n7636_8799.n393 161.3
R23339 a_n7636_8799.n81 a_n7636_8799.n80 161.3
R23340 a_n7636_8799.n79 a_n7636_8799.n20 161.3
R23341 a_n7636_8799.n78 a_n7636_8799.n77 161.3
R23342 a_n7636_8799.n76 a_n7636_8799.n21 161.3
R23343 a_n7636_8799.n75 a_n7636_8799.n74 161.3
R23344 a_n7636_8799.n73 a_n7636_8799.n22 161.3
R23345 a_n7636_8799.n72 a_n7636_8799.n71 161.3
R23346 a_n7636_8799.n70 a_n7636_8799.n23 161.3
R23347 a_n7636_8799.n69 a_n7636_8799.n68 161.3
R23348 a_n7636_8799.n67 a_n7636_8799.n24 161.3
R23349 a_n7636_8799.n66 a_n7636_8799.n65 161.3
R23350 a_n7636_8799.n64 a_n7636_8799.n25 161.3
R23351 a_n7636_8799.n63 a_n7636_8799.n62 161.3
R23352 a_n7636_8799.n61 a_n7636_8799.n26 161.3
R23353 a_n7636_8799.n60 a_n7636_8799.n59 161.3
R23354 a_n7636_8799.n58 a_n7636_8799.n27 161.3
R23355 a_n7636_8799.n57 a_n7636_8799.n56 161.3
R23356 a_n7636_8799.n55 a_n7636_8799.n28 161.3
R23357 a_n7636_8799.n54 a_n7636_8799.n53 161.3
R23358 a_n7636_8799.n52 a_n7636_8799.n29 161.3
R23359 a_n7636_8799.n51 a_n7636_8799.n50 161.3
R23360 a_n7636_8799.n49 a_n7636_8799.n30 161.3
R23361 a_n7636_8799.n48 a_n7636_8799.n47 161.3
R23362 a_n7636_8799.n46 a_n7636_8799.n31 161.3
R23363 a_n7636_8799.n45 a_n7636_8799.n44 161.3
R23364 a_n7636_8799.n43 a_n7636_8799.n32 161.3
R23365 a_n7636_8799.n42 a_n7636_8799.n41 161.3
R23366 a_n7636_8799.n40 a_n7636_8799.n33 161.3
R23367 a_n7636_8799.n39 a_n7636_8799.n38 161.3
R23368 a_n7636_8799.n37 a_n7636_8799.n34 161.3
R23369 a_n7636_8799.n143 a_n7636_8799.n142 161.3
R23370 a_n7636_8799.n141 a_n7636_8799.n82 161.3
R23371 a_n7636_8799.n140 a_n7636_8799.n139 161.3
R23372 a_n7636_8799.n138 a_n7636_8799.n83 161.3
R23373 a_n7636_8799.n137 a_n7636_8799.n136 161.3
R23374 a_n7636_8799.n135 a_n7636_8799.n84 161.3
R23375 a_n7636_8799.n134 a_n7636_8799.n133 161.3
R23376 a_n7636_8799.n132 a_n7636_8799.n85 161.3
R23377 a_n7636_8799.n131 a_n7636_8799.n130 161.3
R23378 a_n7636_8799.n129 a_n7636_8799.n86 161.3
R23379 a_n7636_8799.n128 a_n7636_8799.n127 161.3
R23380 a_n7636_8799.n126 a_n7636_8799.n87 161.3
R23381 a_n7636_8799.n125 a_n7636_8799.n124 161.3
R23382 a_n7636_8799.n123 a_n7636_8799.n88 161.3
R23383 a_n7636_8799.n122 a_n7636_8799.n121 161.3
R23384 a_n7636_8799.n120 a_n7636_8799.n89 161.3
R23385 a_n7636_8799.n119 a_n7636_8799.n118 161.3
R23386 a_n7636_8799.n117 a_n7636_8799.n90 161.3
R23387 a_n7636_8799.n116 a_n7636_8799.n115 161.3
R23388 a_n7636_8799.n114 a_n7636_8799.n91 161.3
R23389 a_n7636_8799.n113 a_n7636_8799.n112 161.3
R23390 a_n7636_8799.n111 a_n7636_8799.n92 161.3
R23391 a_n7636_8799.n110 a_n7636_8799.n109 161.3
R23392 a_n7636_8799.n108 a_n7636_8799.n93 161.3
R23393 a_n7636_8799.n107 a_n7636_8799.n106 161.3
R23394 a_n7636_8799.n105 a_n7636_8799.n94 161.3
R23395 a_n7636_8799.n104 a_n7636_8799.n103 161.3
R23396 a_n7636_8799.n102 a_n7636_8799.n95 161.3
R23397 a_n7636_8799.n101 a_n7636_8799.n100 161.3
R23398 a_n7636_8799.n99 a_n7636_8799.n96 161.3
R23399 a_n7636_8799.n206 a_n7636_8799.n205 161.3
R23400 a_n7636_8799.n204 a_n7636_8799.n145 161.3
R23401 a_n7636_8799.n203 a_n7636_8799.n202 161.3
R23402 a_n7636_8799.n201 a_n7636_8799.n146 161.3
R23403 a_n7636_8799.n200 a_n7636_8799.n199 161.3
R23404 a_n7636_8799.n198 a_n7636_8799.n147 161.3
R23405 a_n7636_8799.n197 a_n7636_8799.n196 161.3
R23406 a_n7636_8799.n195 a_n7636_8799.n148 161.3
R23407 a_n7636_8799.n194 a_n7636_8799.n193 161.3
R23408 a_n7636_8799.n192 a_n7636_8799.n149 161.3
R23409 a_n7636_8799.n191 a_n7636_8799.n190 161.3
R23410 a_n7636_8799.n189 a_n7636_8799.n150 161.3
R23411 a_n7636_8799.n188 a_n7636_8799.n187 161.3
R23412 a_n7636_8799.n186 a_n7636_8799.n151 161.3
R23413 a_n7636_8799.n185 a_n7636_8799.n184 161.3
R23414 a_n7636_8799.n183 a_n7636_8799.n152 161.3
R23415 a_n7636_8799.n182 a_n7636_8799.n181 161.3
R23416 a_n7636_8799.n180 a_n7636_8799.n153 161.3
R23417 a_n7636_8799.n179 a_n7636_8799.n178 161.3
R23418 a_n7636_8799.n177 a_n7636_8799.n154 161.3
R23419 a_n7636_8799.n176 a_n7636_8799.n175 161.3
R23420 a_n7636_8799.n174 a_n7636_8799.n155 161.3
R23421 a_n7636_8799.n173 a_n7636_8799.n172 161.3
R23422 a_n7636_8799.n171 a_n7636_8799.n156 161.3
R23423 a_n7636_8799.n170 a_n7636_8799.n169 161.3
R23424 a_n7636_8799.n168 a_n7636_8799.n157 161.3
R23425 a_n7636_8799.n167 a_n7636_8799.n166 161.3
R23426 a_n7636_8799.n165 a_n7636_8799.n158 161.3
R23427 a_n7636_8799.n164 a_n7636_8799.n163 161.3
R23428 a_n7636_8799.n162 a_n7636_8799.n159 161.3
R23429 a_n7636_8799.n2 a_n7636_8799.n0 98.9633
R23430 a_n7636_8799.n402 a_n7636_8799.n401 98.9631
R23431 a_n7636_8799.n400 a_n7636_8799.n399 98.6055
R23432 a_n7636_8799.n4 a_n7636_8799.n3 98.6055
R23433 a_n7636_8799.n2 a_n7636_8799.n1 98.6055
R23434 a_n7636_8799.n403 a_n7636_8799.n402 98.6054
R23435 a_n7636_8799.n7 a_n7636_8799.n5 81.2902
R23436 a_n7636_8799.n13 a_n7636_8799.n11 81.2902
R23437 a_n7636_8799.n10 a_n7636_8799.n8 81.2902
R23438 a_n7636_8799.n16 a_n7636_8799.n15 80.9324
R23439 a_n7636_8799.n18 a_n7636_8799.n17 80.9324
R23440 a_n7636_8799.n7 a_n7636_8799.n6 80.9324
R23441 a_n7636_8799.n13 a_n7636_8799.n12 80.9324
R23442 a_n7636_8799.n10 a_n7636_8799.n9 80.9324
R23443 a_n7636_8799.n228 a_n7636_8799.n225 70.4033
R23444 a_n7636_8799.n290 a_n7636_8799.n287 70.4033
R23445 a_n7636_8799.n353 a_n7636_8799.n350 70.4033
R23446 a_n7636_8799.n35 a_n7636_8799.n34 70.4033
R23447 a_n7636_8799.n97 a_n7636_8799.n96 70.4033
R23448 a_n7636_8799.n160 a_n7636_8799.n159 70.4033
R23449 a_n7636_8799.n268 a_n7636_8799.n267 48.2005
R23450 a_n7636_8799.n261 a_n7636_8799.n260 48.2005
R23451 a_n7636_8799.n254 a_n7636_8799.n253 48.2005
R23452 a_n7636_8799.n247 a_n7636_8799.n246 48.2005
R23453 a_n7636_8799.n240 a_n7636_8799.n239 48.2005
R23454 a_n7636_8799.n233 a_n7636_8799.n232 48.2005
R23455 a_n7636_8799.n330 a_n7636_8799.n329 48.2005
R23456 a_n7636_8799.n323 a_n7636_8799.n322 48.2005
R23457 a_n7636_8799.n316 a_n7636_8799.n315 48.2005
R23458 a_n7636_8799.n309 a_n7636_8799.n308 48.2005
R23459 a_n7636_8799.n302 a_n7636_8799.n301 48.2005
R23460 a_n7636_8799.n295 a_n7636_8799.n294 48.2005
R23461 a_n7636_8799.n393 a_n7636_8799.n392 48.2005
R23462 a_n7636_8799.n386 a_n7636_8799.n385 48.2005
R23463 a_n7636_8799.n379 a_n7636_8799.n378 48.2005
R23464 a_n7636_8799.n372 a_n7636_8799.n371 48.2005
R23465 a_n7636_8799.n365 a_n7636_8799.n364 48.2005
R23466 a_n7636_8799.n358 a_n7636_8799.n357 48.2005
R23467 a_n7636_8799.n43 a_n7636_8799.n42 48.2005
R23468 a_n7636_8799.n50 a_n7636_8799.n49 48.2005
R23469 a_n7636_8799.n56 a_n7636_8799.n27 48.2005
R23470 a_n7636_8799.n66 a_n7636_8799.n25 48.2005
R23471 a_n7636_8799.n73 a_n7636_8799.n72 48.2005
R23472 a_n7636_8799.n80 a_n7636_8799.n79 48.2005
R23473 a_n7636_8799.n105 a_n7636_8799.n104 48.2005
R23474 a_n7636_8799.n112 a_n7636_8799.n111 48.2005
R23475 a_n7636_8799.n118 a_n7636_8799.n89 48.2005
R23476 a_n7636_8799.n128 a_n7636_8799.n87 48.2005
R23477 a_n7636_8799.n135 a_n7636_8799.n134 48.2005
R23478 a_n7636_8799.n142 a_n7636_8799.n141 48.2005
R23479 a_n7636_8799.n168 a_n7636_8799.n167 48.2005
R23480 a_n7636_8799.n175 a_n7636_8799.n174 48.2005
R23481 a_n7636_8799.n181 a_n7636_8799.n152 48.2005
R23482 a_n7636_8799.n191 a_n7636_8799.n150 48.2005
R23483 a_n7636_8799.n198 a_n7636_8799.n197 48.2005
R23484 a_n7636_8799.n205 a_n7636_8799.n204 48.2005
R23485 a_n7636_8799.n266 a_n7636_8799.n209 40.1672
R23486 a_n7636_8799.n227 a_n7636_8799.n224 40.1672
R23487 a_n7636_8799.n328 a_n7636_8799.n271 40.1672
R23488 a_n7636_8799.n289 a_n7636_8799.n286 40.1672
R23489 a_n7636_8799.n391 a_n7636_8799.n334 40.1672
R23490 a_n7636_8799.n352 a_n7636_8799.n349 40.1672
R23491 a_n7636_8799.n38 a_n7636_8799.n37 40.1672
R23492 a_n7636_8799.n78 a_n7636_8799.n21 40.1672
R23493 a_n7636_8799.n100 a_n7636_8799.n99 40.1672
R23494 a_n7636_8799.n140 a_n7636_8799.n83 40.1672
R23495 a_n7636_8799.n163 a_n7636_8799.n162 40.1672
R23496 a_n7636_8799.n203 a_n7636_8799.n146 40.1672
R23497 a_n7636_8799.n259 a_n7636_8799.n212 38.7066
R23498 a_n7636_8799.n234 a_n7636_8799.n221 38.7066
R23499 a_n7636_8799.n321 a_n7636_8799.n274 38.7066
R23500 a_n7636_8799.n296 a_n7636_8799.n283 38.7066
R23501 a_n7636_8799.n384 a_n7636_8799.n337 38.7066
R23502 a_n7636_8799.n359 a_n7636_8799.n346 38.7066
R23503 a_n7636_8799.n44 a_n7636_8799.n31 38.7066
R23504 a_n7636_8799.n68 a_n7636_8799.n23 38.7066
R23505 a_n7636_8799.n106 a_n7636_8799.n93 38.7066
R23506 a_n7636_8799.n130 a_n7636_8799.n85 38.7066
R23507 a_n7636_8799.n169 a_n7636_8799.n156 38.7066
R23508 a_n7636_8799.n193 a_n7636_8799.n148 38.7066
R23509 a_n7636_8799.n252 a_n7636_8799.n215 37.246
R23510 a_n7636_8799.n241 a_n7636_8799.n218 37.246
R23511 a_n7636_8799.n314 a_n7636_8799.n277 37.246
R23512 a_n7636_8799.n303 a_n7636_8799.n280 37.246
R23513 a_n7636_8799.n377 a_n7636_8799.n340 37.246
R23514 a_n7636_8799.n366 a_n7636_8799.n343 37.246
R23515 a_n7636_8799.n54 a_n7636_8799.n29 37.246
R23516 a_n7636_8799.n62 a_n7636_8799.n61 37.246
R23517 a_n7636_8799.n116 a_n7636_8799.n91 37.246
R23518 a_n7636_8799.n124 a_n7636_8799.n123 37.246
R23519 a_n7636_8799.n179 a_n7636_8799.n154 37.246
R23520 a_n7636_8799.n187 a_n7636_8799.n186 37.246
R23521 a_n7636_8799.n248 a_n7636_8799.n215 35.7853
R23522 a_n7636_8799.n245 a_n7636_8799.n218 35.7853
R23523 a_n7636_8799.n310 a_n7636_8799.n277 35.7853
R23524 a_n7636_8799.n307 a_n7636_8799.n280 35.7853
R23525 a_n7636_8799.n373 a_n7636_8799.n340 35.7853
R23526 a_n7636_8799.n370 a_n7636_8799.n343 35.7853
R23527 a_n7636_8799.n55 a_n7636_8799.n54 35.7853
R23528 a_n7636_8799.n61 a_n7636_8799.n60 35.7853
R23529 a_n7636_8799.n117 a_n7636_8799.n116 35.7853
R23530 a_n7636_8799.n123 a_n7636_8799.n122 35.7853
R23531 a_n7636_8799.n180 a_n7636_8799.n179 35.7853
R23532 a_n7636_8799.n186 a_n7636_8799.n185 35.7853
R23533 a_n7636_8799.n255 a_n7636_8799.n212 34.3247
R23534 a_n7636_8799.n238 a_n7636_8799.n221 34.3247
R23535 a_n7636_8799.n317 a_n7636_8799.n274 34.3247
R23536 a_n7636_8799.n300 a_n7636_8799.n283 34.3247
R23537 a_n7636_8799.n380 a_n7636_8799.n337 34.3247
R23538 a_n7636_8799.n363 a_n7636_8799.n346 34.3247
R23539 a_n7636_8799.n48 a_n7636_8799.n31 34.3247
R23540 a_n7636_8799.n68 a_n7636_8799.n67 34.3247
R23541 a_n7636_8799.n110 a_n7636_8799.n93 34.3247
R23542 a_n7636_8799.n130 a_n7636_8799.n129 34.3247
R23543 a_n7636_8799.n173 a_n7636_8799.n156 34.3247
R23544 a_n7636_8799.n193 a_n7636_8799.n192 34.3247
R23545 a_n7636_8799.n262 a_n7636_8799.n209 32.8641
R23546 a_n7636_8799.n231 a_n7636_8799.n224 32.8641
R23547 a_n7636_8799.n324 a_n7636_8799.n271 32.8641
R23548 a_n7636_8799.n293 a_n7636_8799.n286 32.8641
R23549 a_n7636_8799.n387 a_n7636_8799.n334 32.8641
R23550 a_n7636_8799.n356 a_n7636_8799.n349 32.8641
R23551 a_n7636_8799.n38 a_n7636_8799.n33 32.8641
R23552 a_n7636_8799.n74 a_n7636_8799.n21 32.8641
R23553 a_n7636_8799.n100 a_n7636_8799.n95 32.8641
R23554 a_n7636_8799.n136 a_n7636_8799.n83 32.8641
R23555 a_n7636_8799.n163 a_n7636_8799.n158 32.8641
R23556 a_n7636_8799.n199 a_n7636_8799.n146 32.8641
R23557 a_n7636_8799.n16 a_n7636_8799.n14 31.4401
R23558 a_n7636_8799.n400 a_n7636_8799.n398 30.3191
R23559 a_n7636_8799.n226 a_n7636_8799.n225 20.9576
R23560 a_n7636_8799.n288 a_n7636_8799.n287 20.9576
R23561 a_n7636_8799.n351 a_n7636_8799.n350 20.9576
R23562 a_n7636_8799.n36 a_n7636_8799.n35 20.9576
R23563 a_n7636_8799.n98 a_n7636_8799.n97 20.9576
R23564 a_n7636_8799.n161 a_n7636_8799.n160 20.9576
R23565 a_n7636_8799.n398 a_n7636_8799.n4 18.1305
R23566 a_n7636_8799.n262 a_n7636_8799.n261 15.3369
R23567 a_n7636_8799.n232 a_n7636_8799.n231 15.3369
R23568 a_n7636_8799.n324 a_n7636_8799.n323 15.3369
R23569 a_n7636_8799.n294 a_n7636_8799.n293 15.3369
R23570 a_n7636_8799.n387 a_n7636_8799.n386 15.3369
R23571 a_n7636_8799.n357 a_n7636_8799.n356 15.3369
R23572 a_n7636_8799.n42 a_n7636_8799.n33 15.3369
R23573 a_n7636_8799.n74 a_n7636_8799.n73 15.3369
R23574 a_n7636_8799.n104 a_n7636_8799.n95 15.3369
R23575 a_n7636_8799.n136 a_n7636_8799.n135 15.3369
R23576 a_n7636_8799.n167 a_n7636_8799.n158 15.3369
R23577 a_n7636_8799.n199 a_n7636_8799.n198 15.3369
R23578 a_n7636_8799.n255 a_n7636_8799.n254 13.8763
R23579 a_n7636_8799.n239 a_n7636_8799.n238 13.8763
R23580 a_n7636_8799.n317 a_n7636_8799.n316 13.8763
R23581 a_n7636_8799.n301 a_n7636_8799.n300 13.8763
R23582 a_n7636_8799.n380 a_n7636_8799.n379 13.8763
R23583 a_n7636_8799.n364 a_n7636_8799.n363 13.8763
R23584 a_n7636_8799.n49 a_n7636_8799.n48 13.8763
R23585 a_n7636_8799.n67 a_n7636_8799.n66 13.8763
R23586 a_n7636_8799.n111 a_n7636_8799.n110 13.8763
R23587 a_n7636_8799.n129 a_n7636_8799.n128 13.8763
R23588 a_n7636_8799.n174 a_n7636_8799.n173 13.8763
R23589 a_n7636_8799.n192 a_n7636_8799.n191 13.8763
R23590 a_n7636_8799.n248 a_n7636_8799.n247 12.4157
R23591 a_n7636_8799.n246 a_n7636_8799.n245 12.4157
R23592 a_n7636_8799.n310 a_n7636_8799.n309 12.4157
R23593 a_n7636_8799.n308 a_n7636_8799.n307 12.4157
R23594 a_n7636_8799.n373 a_n7636_8799.n372 12.4157
R23595 a_n7636_8799.n371 a_n7636_8799.n370 12.4157
R23596 a_n7636_8799.n56 a_n7636_8799.n55 12.4157
R23597 a_n7636_8799.n60 a_n7636_8799.n27 12.4157
R23598 a_n7636_8799.n118 a_n7636_8799.n117 12.4157
R23599 a_n7636_8799.n122 a_n7636_8799.n89 12.4157
R23600 a_n7636_8799.n181 a_n7636_8799.n180 12.4157
R23601 a_n7636_8799.n185 a_n7636_8799.n152 12.4157
R23602 a_n7636_8799.n397 a_n7636_8799.n19 12.3339
R23603 a_n7636_8799.n398 a_n7636_8799.n397 11.4887
R23604 a_n7636_8799.n253 a_n7636_8799.n252 10.955
R23605 a_n7636_8799.n241 a_n7636_8799.n240 10.955
R23606 a_n7636_8799.n315 a_n7636_8799.n314 10.955
R23607 a_n7636_8799.n303 a_n7636_8799.n302 10.955
R23608 a_n7636_8799.n378 a_n7636_8799.n377 10.955
R23609 a_n7636_8799.n366 a_n7636_8799.n365 10.955
R23610 a_n7636_8799.n50 a_n7636_8799.n29 10.955
R23611 a_n7636_8799.n62 a_n7636_8799.n25 10.955
R23612 a_n7636_8799.n112 a_n7636_8799.n91 10.955
R23613 a_n7636_8799.n124 a_n7636_8799.n87 10.955
R23614 a_n7636_8799.n175 a_n7636_8799.n154 10.955
R23615 a_n7636_8799.n187 a_n7636_8799.n150 10.955
R23616 a_n7636_8799.n260 a_n7636_8799.n259 9.49444
R23617 a_n7636_8799.n234 a_n7636_8799.n233 9.49444
R23618 a_n7636_8799.n322 a_n7636_8799.n321 9.49444
R23619 a_n7636_8799.n296 a_n7636_8799.n295 9.49444
R23620 a_n7636_8799.n385 a_n7636_8799.n384 9.49444
R23621 a_n7636_8799.n359 a_n7636_8799.n358 9.49444
R23622 a_n7636_8799.n44 a_n7636_8799.n43 9.49444
R23623 a_n7636_8799.n72 a_n7636_8799.n23 9.49444
R23624 a_n7636_8799.n106 a_n7636_8799.n105 9.49444
R23625 a_n7636_8799.n134 a_n7636_8799.n85 9.49444
R23626 a_n7636_8799.n169 a_n7636_8799.n168 9.49444
R23627 a_n7636_8799.n197 a_n7636_8799.n148 9.49444
R23628 a_n7636_8799.n332 a_n7636_8799.n269 9.04406
R23629 a_n7636_8799.n144 a_n7636_8799.n81 9.04406
R23630 a_n7636_8799.n267 a_n7636_8799.n266 8.03383
R23631 a_n7636_8799.n227 a_n7636_8799.n226 8.03383
R23632 a_n7636_8799.n329 a_n7636_8799.n328 8.03383
R23633 a_n7636_8799.n289 a_n7636_8799.n288 8.03383
R23634 a_n7636_8799.n392 a_n7636_8799.n391 8.03383
R23635 a_n7636_8799.n352 a_n7636_8799.n351 8.03383
R23636 a_n7636_8799.n37 a_n7636_8799.n36 8.03383
R23637 a_n7636_8799.n79 a_n7636_8799.n78 8.03383
R23638 a_n7636_8799.n99 a_n7636_8799.n98 8.03383
R23639 a_n7636_8799.n141 a_n7636_8799.n140 8.03383
R23640 a_n7636_8799.n162 a_n7636_8799.n161 8.03383
R23641 a_n7636_8799.n204 a_n7636_8799.n203 8.03383
R23642 a_n7636_8799.n396 a_n7636_8799.n207 6.81251
R23643 a_n7636_8799.n396 a_n7636_8799.n395 6.5703
R23644 a_n7636_8799.n332 a_n7636_8799.n331 4.93611
R23645 a_n7636_8799.n395 a_n7636_8799.n394 4.93611
R23646 a_n7636_8799.n144 a_n7636_8799.n143 4.93611
R23647 a_n7636_8799.n207 a_n7636_8799.n206 4.93611
R23648 a_n7636_8799.n395 a_n7636_8799.n332 4.10845
R23649 a_n7636_8799.n207 a_n7636_8799.n144 4.10845
R23650 a_n7636_8799.n401 a_n7636_8799.t12 3.61217
R23651 a_n7636_8799.n401 a_n7636_8799.t17 3.61217
R23652 a_n7636_8799.n399 a_n7636_8799.t10 3.61217
R23653 a_n7636_8799.n399 a_n7636_8799.t9 3.61217
R23654 a_n7636_8799.n3 a_n7636_8799.t11 3.61217
R23655 a_n7636_8799.n3 a_n7636_8799.t8 3.61217
R23656 a_n7636_8799.n1 a_n7636_8799.t13 3.61217
R23657 a_n7636_8799.n1 a_n7636_8799.t16 3.61217
R23658 a_n7636_8799.n0 a_n7636_8799.t7 3.61217
R23659 a_n7636_8799.n0 a_n7636_8799.t14 3.61217
R23660 a_n7636_8799.t18 a_n7636_8799.n403 3.61217
R23661 a_n7636_8799.n403 a_n7636_8799.t15 3.61217
R23662 a_n7636_8799.n397 a_n7636_8799.n396 3.4105
R23663 a_n7636_8799.n15 a_n7636_8799.t6 2.82907
R23664 a_n7636_8799.n15 a_n7636_8799.t2 2.82907
R23665 a_n7636_8799.n17 a_n7636_8799.t4 2.82907
R23666 a_n7636_8799.n17 a_n7636_8799.t5 2.82907
R23667 a_n7636_8799.n6 a_n7636_8799.t26 2.82907
R23668 a_n7636_8799.n6 a_n7636_8799.t1 2.82907
R23669 a_n7636_8799.n5 a_n7636_8799.t25 2.82907
R23670 a_n7636_8799.n5 a_n7636_8799.t22 2.82907
R23671 a_n7636_8799.n11 a_n7636_8799.t3 2.82907
R23672 a_n7636_8799.n11 a_n7636_8799.t23 2.82907
R23673 a_n7636_8799.n12 a_n7636_8799.t20 2.82907
R23674 a_n7636_8799.n12 a_n7636_8799.t19 2.82907
R23675 a_n7636_8799.n9 a_n7636_8799.t0 2.82907
R23676 a_n7636_8799.n9 a_n7636_8799.t24 2.82907
R23677 a_n7636_8799.n8 a_n7636_8799.t21 2.82907
R23678 a_n7636_8799.n8 a_n7636_8799.t27 2.82907
R23679 a_n7636_8799.n18 a_n7636_8799.n16 0.358259
R23680 a_n7636_8799.n4 a_n7636_8799.n2 0.358259
R23681 a_n7636_8799.n402 a_n7636_8799.n400 0.358259
R23682 a_n7636_8799.n269 a_n7636_8799.n208 0.189894
R23683 a_n7636_8799.n265 a_n7636_8799.n208 0.189894
R23684 a_n7636_8799.n265 a_n7636_8799.n264 0.189894
R23685 a_n7636_8799.n264 a_n7636_8799.n263 0.189894
R23686 a_n7636_8799.n263 a_n7636_8799.n210 0.189894
R23687 a_n7636_8799.n211 a_n7636_8799.n210 0.189894
R23688 a_n7636_8799.n258 a_n7636_8799.n211 0.189894
R23689 a_n7636_8799.n258 a_n7636_8799.n257 0.189894
R23690 a_n7636_8799.n257 a_n7636_8799.n256 0.189894
R23691 a_n7636_8799.n256 a_n7636_8799.n213 0.189894
R23692 a_n7636_8799.n214 a_n7636_8799.n213 0.189894
R23693 a_n7636_8799.n251 a_n7636_8799.n214 0.189894
R23694 a_n7636_8799.n251 a_n7636_8799.n250 0.189894
R23695 a_n7636_8799.n250 a_n7636_8799.n249 0.189894
R23696 a_n7636_8799.n249 a_n7636_8799.n216 0.189894
R23697 a_n7636_8799.n217 a_n7636_8799.n216 0.189894
R23698 a_n7636_8799.n244 a_n7636_8799.n217 0.189894
R23699 a_n7636_8799.n244 a_n7636_8799.n243 0.189894
R23700 a_n7636_8799.n243 a_n7636_8799.n242 0.189894
R23701 a_n7636_8799.n242 a_n7636_8799.n219 0.189894
R23702 a_n7636_8799.n220 a_n7636_8799.n219 0.189894
R23703 a_n7636_8799.n237 a_n7636_8799.n220 0.189894
R23704 a_n7636_8799.n237 a_n7636_8799.n236 0.189894
R23705 a_n7636_8799.n236 a_n7636_8799.n235 0.189894
R23706 a_n7636_8799.n235 a_n7636_8799.n222 0.189894
R23707 a_n7636_8799.n223 a_n7636_8799.n222 0.189894
R23708 a_n7636_8799.n230 a_n7636_8799.n223 0.189894
R23709 a_n7636_8799.n230 a_n7636_8799.n229 0.189894
R23710 a_n7636_8799.n229 a_n7636_8799.n228 0.189894
R23711 a_n7636_8799.n331 a_n7636_8799.n270 0.189894
R23712 a_n7636_8799.n327 a_n7636_8799.n270 0.189894
R23713 a_n7636_8799.n327 a_n7636_8799.n326 0.189894
R23714 a_n7636_8799.n326 a_n7636_8799.n325 0.189894
R23715 a_n7636_8799.n325 a_n7636_8799.n272 0.189894
R23716 a_n7636_8799.n273 a_n7636_8799.n272 0.189894
R23717 a_n7636_8799.n320 a_n7636_8799.n273 0.189894
R23718 a_n7636_8799.n320 a_n7636_8799.n319 0.189894
R23719 a_n7636_8799.n319 a_n7636_8799.n318 0.189894
R23720 a_n7636_8799.n318 a_n7636_8799.n275 0.189894
R23721 a_n7636_8799.n276 a_n7636_8799.n275 0.189894
R23722 a_n7636_8799.n313 a_n7636_8799.n276 0.189894
R23723 a_n7636_8799.n313 a_n7636_8799.n312 0.189894
R23724 a_n7636_8799.n312 a_n7636_8799.n311 0.189894
R23725 a_n7636_8799.n311 a_n7636_8799.n278 0.189894
R23726 a_n7636_8799.n279 a_n7636_8799.n278 0.189894
R23727 a_n7636_8799.n306 a_n7636_8799.n279 0.189894
R23728 a_n7636_8799.n306 a_n7636_8799.n305 0.189894
R23729 a_n7636_8799.n305 a_n7636_8799.n304 0.189894
R23730 a_n7636_8799.n304 a_n7636_8799.n281 0.189894
R23731 a_n7636_8799.n282 a_n7636_8799.n281 0.189894
R23732 a_n7636_8799.n299 a_n7636_8799.n282 0.189894
R23733 a_n7636_8799.n299 a_n7636_8799.n298 0.189894
R23734 a_n7636_8799.n298 a_n7636_8799.n297 0.189894
R23735 a_n7636_8799.n297 a_n7636_8799.n284 0.189894
R23736 a_n7636_8799.n285 a_n7636_8799.n284 0.189894
R23737 a_n7636_8799.n292 a_n7636_8799.n285 0.189894
R23738 a_n7636_8799.n292 a_n7636_8799.n291 0.189894
R23739 a_n7636_8799.n291 a_n7636_8799.n290 0.189894
R23740 a_n7636_8799.n394 a_n7636_8799.n333 0.189894
R23741 a_n7636_8799.n390 a_n7636_8799.n333 0.189894
R23742 a_n7636_8799.n390 a_n7636_8799.n389 0.189894
R23743 a_n7636_8799.n389 a_n7636_8799.n388 0.189894
R23744 a_n7636_8799.n388 a_n7636_8799.n335 0.189894
R23745 a_n7636_8799.n336 a_n7636_8799.n335 0.189894
R23746 a_n7636_8799.n383 a_n7636_8799.n336 0.189894
R23747 a_n7636_8799.n383 a_n7636_8799.n382 0.189894
R23748 a_n7636_8799.n382 a_n7636_8799.n381 0.189894
R23749 a_n7636_8799.n381 a_n7636_8799.n338 0.189894
R23750 a_n7636_8799.n339 a_n7636_8799.n338 0.189894
R23751 a_n7636_8799.n376 a_n7636_8799.n339 0.189894
R23752 a_n7636_8799.n376 a_n7636_8799.n375 0.189894
R23753 a_n7636_8799.n375 a_n7636_8799.n374 0.189894
R23754 a_n7636_8799.n374 a_n7636_8799.n341 0.189894
R23755 a_n7636_8799.n342 a_n7636_8799.n341 0.189894
R23756 a_n7636_8799.n369 a_n7636_8799.n342 0.189894
R23757 a_n7636_8799.n369 a_n7636_8799.n368 0.189894
R23758 a_n7636_8799.n368 a_n7636_8799.n367 0.189894
R23759 a_n7636_8799.n367 a_n7636_8799.n344 0.189894
R23760 a_n7636_8799.n345 a_n7636_8799.n344 0.189894
R23761 a_n7636_8799.n362 a_n7636_8799.n345 0.189894
R23762 a_n7636_8799.n362 a_n7636_8799.n361 0.189894
R23763 a_n7636_8799.n361 a_n7636_8799.n360 0.189894
R23764 a_n7636_8799.n360 a_n7636_8799.n347 0.189894
R23765 a_n7636_8799.n348 a_n7636_8799.n347 0.189894
R23766 a_n7636_8799.n355 a_n7636_8799.n348 0.189894
R23767 a_n7636_8799.n355 a_n7636_8799.n354 0.189894
R23768 a_n7636_8799.n354 a_n7636_8799.n353 0.189894
R23769 a_n7636_8799.n39 a_n7636_8799.n34 0.189894
R23770 a_n7636_8799.n40 a_n7636_8799.n39 0.189894
R23771 a_n7636_8799.n41 a_n7636_8799.n40 0.189894
R23772 a_n7636_8799.n41 a_n7636_8799.n32 0.189894
R23773 a_n7636_8799.n45 a_n7636_8799.n32 0.189894
R23774 a_n7636_8799.n46 a_n7636_8799.n45 0.189894
R23775 a_n7636_8799.n47 a_n7636_8799.n46 0.189894
R23776 a_n7636_8799.n47 a_n7636_8799.n30 0.189894
R23777 a_n7636_8799.n51 a_n7636_8799.n30 0.189894
R23778 a_n7636_8799.n52 a_n7636_8799.n51 0.189894
R23779 a_n7636_8799.n53 a_n7636_8799.n52 0.189894
R23780 a_n7636_8799.n53 a_n7636_8799.n28 0.189894
R23781 a_n7636_8799.n57 a_n7636_8799.n28 0.189894
R23782 a_n7636_8799.n58 a_n7636_8799.n57 0.189894
R23783 a_n7636_8799.n59 a_n7636_8799.n58 0.189894
R23784 a_n7636_8799.n59 a_n7636_8799.n26 0.189894
R23785 a_n7636_8799.n63 a_n7636_8799.n26 0.189894
R23786 a_n7636_8799.n64 a_n7636_8799.n63 0.189894
R23787 a_n7636_8799.n65 a_n7636_8799.n64 0.189894
R23788 a_n7636_8799.n65 a_n7636_8799.n24 0.189894
R23789 a_n7636_8799.n69 a_n7636_8799.n24 0.189894
R23790 a_n7636_8799.n70 a_n7636_8799.n69 0.189894
R23791 a_n7636_8799.n71 a_n7636_8799.n70 0.189894
R23792 a_n7636_8799.n71 a_n7636_8799.n22 0.189894
R23793 a_n7636_8799.n75 a_n7636_8799.n22 0.189894
R23794 a_n7636_8799.n76 a_n7636_8799.n75 0.189894
R23795 a_n7636_8799.n77 a_n7636_8799.n76 0.189894
R23796 a_n7636_8799.n77 a_n7636_8799.n20 0.189894
R23797 a_n7636_8799.n81 a_n7636_8799.n20 0.189894
R23798 a_n7636_8799.n101 a_n7636_8799.n96 0.189894
R23799 a_n7636_8799.n102 a_n7636_8799.n101 0.189894
R23800 a_n7636_8799.n103 a_n7636_8799.n102 0.189894
R23801 a_n7636_8799.n103 a_n7636_8799.n94 0.189894
R23802 a_n7636_8799.n107 a_n7636_8799.n94 0.189894
R23803 a_n7636_8799.n108 a_n7636_8799.n107 0.189894
R23804 a_n7636_8799.n109 a_n7636_8799.n108 0.189894
R23805 a_n7636_8799.n109 a_n7636_8799.n92 0.189894
R23806 a_n7636_8799.n113 a_n7636_8799.n92 0.189894
R23807 a_n7636_8799.n114 a_n7636_8799.n113 0.189894
R23808 a_n7636_8799.n115 a_n7636_8799.n114 0.189894
R23809 a_n7636_8799.n115 a_n7636_8799.n90 0.189894
R23810 a_n7636_8799.n119 a_n7636_8799.n90 0.189894
R23811 a_n7636_8799.n120 a_n7636_8799.n119 0.189894
R23812 a_n7636_8799.n121 a_n7636_8799.n120 0.189894
R23813 a_n7636_8799.n121 a_n7636_8799.n88 0.189894
R23814 a_n7636_8799.n125 a_n7636_8799.n88 0.189894
R23815 a_n7636_8799.n126 a_n7636_8799.n125 0.189894
R23816 a_n7636_8799.n127 a_n7636_8799.n126 0.189894
R23817 a_n7636_8799.n127 a_n7636_8799.n86 0.189894
R23818 a_n7636_8799.n131 a_n7636_8799.n86 0.189894
R23819 a_n7636_8799.n132 a_n7636_8799.n131 0.189894
R23820 a_n7636_8799.n133 a_n7636_8799.n132 0.189894
R23821 a_n7636_8799.n133 a_n7636_8799.n84 0.189894
R23822 a_n7636_8799.n137 a_n7636_8799.n84 0.189894
R23823 a_n7636_8799.n138 a_n7636_8799.n137 0.189894
R23824 a_n7636_8799.n139 a_n7636_8799.n138 0.189894
R23825 a_n7636_8799.n139 a_n7636_8799.n82 0.189894
R23826 a_n7636_8799.n143 a_n7636_8799.n82 0.189894
R23827 a_n7636_8799.n164 a_n7636_8799.n159 0.189894
R23828 a_n7636_8799.n165 a_n7636_8799.n164 0.189894
R23829 a_n7636_8799.n166 a_n7636_8799.n165 0.189894
R23830 a_n7636_8799.n166 a_n7636_8799.n157 0.189894
R23831 a_n7636_8799.n170 a_n7636_8799.n157 0.189894
R23832 a_n7636_8799.n171 a_n7636_8799.n170 0.189894
R23833 a_n7636_8799.n172 a_n7636_8799.n171 0.189894
R23834 a_n7636_8799.n172 a_n7636_8799.n155 0.189894
R23835 a_n7636_8799.n176 a_n7636_8799.n155 0.189894
R23836 a_n7636_8799.n177 a_n7636_8799.n176 0.189894
R23837 a_n7636_8799.n178 a_n7636_8799.n177 0.189894
R23838 a_n7636_8799.n178 a_n7636_8799.n153 0.189894
R23839 a_n7636_8799.n182 a_n7636_8799.n153 0.189894
R23840 a_n7636_8799.n183 a_n7636_8799.n182 0.189894
R23841 a_n7636_8799.n184 a_n7636_8799.n183 0.189894
R23842 a_n7636_8799.n184 a_n7636_8799.n151 0.189894
R23843 a_n7636_8799.n188 a_n7636_8799.n151 0.189894
R23844 a_n7636_8799.n189 a_n7636_8799.n188 0.189894
R23845 a_n7636_8799.n190 a_n7636_8799.n189 0.189894
R23846 a_n7636_8799.n190 a_n7636_8799.n149 0.189894
R23847 a_n7636_8799.n194 a_n7636_8799.n149 0.189894
R23848 a_n7636_8799.n195 a_n7636_8799.n194 0.189894
R23849 a_n7636_8799.n196 a_n7636_8799.n195 0.189894
R23850 a_n7636_8799.n196 a_n7636_8799.n147 0.189894
R23851 a_n7636_8799.n200 a_n7636_8799.n147 0.189894
R23852 a_n7636_8799.n201 a_n7636_8799.n200 0.189894
R23853 a_n7636_8799.n202 a_n7636_8799.n201 0.189894
R23854 a_n7636_8799.n202 a_n7636_8799.n145 0.189894
R23855 a_n7636_8799.n206 a_n7636_8799.n145 0.189894
R23856 a_n7636_8799.n14 a_n7636_8799.n10 0.179379
R23857 a_n7636_8799.n14 a_n7636_8799.n13 0.179379
R23858 a_n7636_8799.n19 a_n7636_8799.n7 0.179379
R23859 a_n7636_8799.n19 a_n7636_8799.n18 0.179379
R23860 plus.n27 plus.t19 436.949
R23861 plus.n5 plus.t11 436.949
R23862 plus.n28 plus.t5 415.966
R23863 plus.n30 plus.t17 415.966
R23864 plus.n34 plus.t20 415.966
R23865 plus.n35 plus.t10 415.966
R23866 plus.n23 plus.t6 415.966
R23867 plus.n41 plus.t9 415.966
R23868 plus.n42 plus.t16 415.966
R23869 plus.n20 plus.t7 415.966
R23870 plus.n19 plus.t15 415.966
R23871 plus.n1 plus.t12 415.966
R23872 plus.n13 plus.t18 415.966
R23873 plus.n12 plus.t14 415.966
R23874 plus.n4 plus.t8 415.966
R23875 plus.n6 plus.t13 415.966
R23876 plus.n46 plus.t4 243.97
R23877 plus.n46 plus.n45 223.454
R23878 plus.n48 plus.n47 223.454
R23879 plus.n43 plus.n42 161.3
R23880 plus.n41 plus.n22 161.3
R23881 plus.n40 plus.n39 161.3
R23882 plus.n38 plus.n23 161.3
R23883 plus.n37 plus.n36 161.3
R23884 plus.n35 plus.n24 161.3
R23885 plus.n34 plus.n33 161.3
R23886 plus.n32 plus.n25 161.3
R23887 plus.n31 plus.n30 161.3
R23888 plus.n29 plus.n26 161.3
R23889 plus.n8 plus.n7 161.3
R23890 plus.n9 plus.n4 161.3
R23891 plus.n11 plus.n10 161.3
R23892 plus.n12 plus.n3 161.3
R23893 plus.n13 plus.n2 161.3
R23894 plus.n15 plus.n14 161.3
R23895 plus.n16 plus.n1 161.3
R23896 plus.n18 plus.n17 161.3
R23897 plus.n19 plus.n0 161.3
R23898 plus.n21 plus.n20 161.3
R23899 plus.n27 plus.n26 70.4033
R23900 plus.n8 plus.n5 70.4033
R23901 plus.n35 plus.n34 48.2005
R23902 plus.n42 plus.n41 48.2005
R23903 plus.n20 plus.n19 48.2005
R23904 plus.n13 plus.n12 48.2005
R23905 plus.n30 plus.n29 37.246
R23906 plus.n40 plus.n23 37.246
R23907 plus.n18 plus.n1 37.246
R23908 plus.n7 plus.n4 37.246
R23909 plus.n30 plus.n25 35.7853
R23910 plus.n36 plus.n23 35.7853
R23911 plus.n14 plus.n1 35.7853
R23912 plus.n11 plus.n4 35.7853
R23913 plus.n44 plus.n43 28.5744
R23914 plus.n28 plus.n27 20.9576
R23915 plus.n6 plus.n5 20.9576
R23916 plus.n45 plus.t0 19.8005
R23917 plus.n45 plus.t1 19.8005
R23918 plus.n47 plus.t3 19.8005
R23919 plus.n47 plus.t2 19.8005
R23920 plus plus.n49 14.5359
R23921 plus.n34 plus.n25 12.4157
R23922 plus.n36 plus.n35 12.4157
R23923 plus.n14 plus.n13 12.4157
R23924 plus.n12 plus.n11 12.4157
R23925 plus.n44 plus.n21 11.76
R23926 plus.n29 plus.n28 10.955
R23927 plus.n41 plus.n40 10.955
R23928 plus.n19 plus.n18 10.955
R23929 plus.n7 plus.n6 10.955
R23930 plus.n49 plus.n48 5.40567
R23931 plus.n49 plus.n44 1.188
R23932 plus.n48 plus.n46 0.716017
R23933 plus.n31 plus.n26 0.189894
R23934 plus.n32 plus.n31 0.189894
R23935 plus.n33 plus.n32 0.189894
R23936 plus.n33 plus.n24 0.189894
R23937 plus.n37 plus.n24 0.189894
R23938 plus.n38 plus.n37 0.189894
R23939 plus.n39 plus.n38 0.189894
R23940 plus.n39 plus.n22 0.189894
R23941 plus.n43 plus.n22 0.189894
R23942 plus.n21 plus.n0 0.189894
R23943 plus.n17 plus.n0 0.189894
R23944 plus.n17 plus.n16 0.189894
R23945 plus.n16 plus.n15 0.189894
R23946 plus.n15 plus.n2 0.189894
R23947 plus.n3 plus.n2 0.189894
R23948 plus.n10 plus.n3 0.189894
R23949 plus.n10 plus.n9 0.189894
R23950 plus.n9 plus.n8 0.189894
R23951 a_n2903_n3924.n10 a_n2903_n3924.t35 214.994
R23952 a_n2903_n3924.n0 a_n2903_n3924.t39 214.975
R23953 a_n2903_n3924.n0 a_n2903_n3924.t36 214.321
R23954 a_n2903_n3924.n11 a_n2903_n3924.t11 214.321
R23955 a_n2903_n3924.n12 a_n2903_n3924.t38 214.321
R23956 a_n2903_n3924.n13 a_n2903_n3924.t12 214.321
R23957 a_n2903_n3924.n14 a_n2903_n3924.t8 214.321
R23958 a_n2903_n3924.n10 a_n2903_n3924.t5 214.321
R23959 a_n2903_n3924.n1 a_n2903_n3924.t14 55.8337
R23960 a_n2903_n3924.n2 a_n2903_n3924.t37 55.8337
R23961 a_n2903_n3924.n9 a_n2903_n3924.t10 55.8337
R23962 a_n2903_n3924.n34 a_n2903_n3924.t17 55.8335
R23963 a_n2903_n3924.n32 a_n2903_n3924.t32 55.8335
R23964 a_n2903_n3924.n25 a_n2903_n3924.t29 55.8335
R23965 a_n2903_n3924.n24 a_n2903_n3924.t22 55.8335
R23966 a_n2903_n3924.n17 a_n2903_n3924.t26 55.8335
R23967 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R23968 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R23969 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R23970 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R23971 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R23972 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R23973 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R23974 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R23975 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R23976 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R23977 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R23978 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R23979 a_n2903_n3924.n16 a_n2903_n3924.n9 12.1555
R23980 a_n2903_n3924.n34 a_n2903_n3924.n33 12.1555
R23981 a_n2903_n3924.n17 a_n2903_n3924.n16 5.07593
R23982 a_n2903_n3924.n33 a_n2903_n3924.n32 5.07593
R23983 a_n2903_n3924.n35 a_n2903_n3924.t27 2.82907
R23984 a_n2903_n3924.n35 a_n2903_n3924.t24 2.82907
R23985 a_n2903_n3924.n37 a_n2903_n3924.t13 2.82907
R23986 a_n2903_n3924.n37 a_n2903_n3924.t23 2.82907
R23987 a_n2903_n3924.n3 a_n2903_n3924.t7 2.82907
R23988 a_n2903_n3924.n3 a_n2903_n3924.t0 2.82907
R23989 a_n2903_n3924.n5 a_n2903_n3924.t9 2.82907
R23990 a_n2903_n3924.n5 a_n2903_n3924.t4 2.82907
R23991 a_n2903_n3924.n7 a_n2903_n3924.t34 2.82907
R23992 a_n2903_n3924.n7 a_n2903_n3924.t33 2.82907
R23993 a_n2903_n3924.n30 a_n2903_n3924.t30 2.82907
R23994 a_n2903_n3924.n30 a_n2903_n3924.t2 2.82907
R23995 a_n2903_n3924.n28 a_n2903_n3924.t1 2.82907
R23996 a_n2903_n3924.n28 a_n2903_n3924.t3 2.82907
R23997 a_n2903_n3924.n26 a_n2903_n3924.t6 2.82907
R23998 a_n2903_n3924.n26 a_n2903_n3924.t31 2.82907
R23999 a_n2903_n3924.n22 a_n2903_n3924.t25 2.82907
R24000 a_n2903_n3924.n22 a_n2903_n3924.t20 2.82907
R24001 a_n2903_n3924.n20 a_n2903_n3924.t15 2.82907
R24002 a_n2903_n3924.n20 a_n2903_n3924.t19 2.82907
R24003 a_n2903_n3924.n18 a_n2903_n3924.t18 2.82907
R24004 a_n2903_n3924.n18 a_n2903_n3924.t21 2.82907
R24005 a_n2903_n3924.t28 a_n2903_n3924.n40 2.82907
R24006 a_n2903_n3924.n40 a_n2903_n3924.t16 2.82907
R24007 a_n2903_n3924.n33 a_n2903_n3924.n0 1.95694
R24008 a_n2903_n3924.n16 a_n2903_n3924.n15 1.95694
R24009 a_n2903_n3924.n11 a_n2903_n3924.n0 0.69018
R24010 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R24011 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R24012 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R24013 a_n2903_n3924.n15 a_n2903_n3924.n10 0.511401
R24014 a_n2903_n3924.n19 a_n2903_n3924.n17 0.358259
R24015 a_n2903_n3924.n21 a_n2903_n3924.n19 0.358259
R24016 a_n2903_n3924.n23 a_n2903_n3924.n21 0.358259
R24017 a_n2903_n3924.n24 a_n2903_n3924.n23 0.358259
R24018 a_n2903_n3924.n27 a_n2903_n3924.n25 0.358259
R24019 a_n2903_n3924.n29 a_n2903_n3924.n27 0.358259
R24020 a_n2903_n3924.n31 a_n2903_n3924.n29 0.358259
R24021 a_n2903_n3924.n32 a_n2903_n3924.n31 0.358259
R24022 a_n2903_n3924.n9 a_n2903_n3924.n8 0.358259
R24023 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R24024 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R24025 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R24026 a_n2903_n3924.n39 a_n2903_n3924.n1 0.358259
R24027 a_n2903_n3924.n39 a_n2903_n3924.n38 0.358259
R24028 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R24029 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R24030 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R24031 a_n2903_n3924.n2 a_n2903_n3924.n1 0.235414
R24032 a_n2903_n3924.n15 a_n2903_n3924.n14 0.16111
R24033 output.n41 output.n15 289.615
R24034 output.n72 output.n46 289.615
R24035 output.n104 output.n78 289.615
R24036 output.n136 output.n110 289.615
R24037 output.n77 output.n45 197.26
R24038 output.n77 output.n76 196.298
R24039 output.n109 output.n108 196.298
R24040 output.n141 output.n140 196.298
R24041 output.n42 output.n41 185
R24042 output.n40 output.n39 185
R24043 output.n19 output.n18 185
R24044 output.n34 output.n33 185
R24045 output.n32 output.n31 185
R24046 output.n23 output.n22 185
R24047 output.n26 output.n25 185
R24048 output.n73 output.n72 185
R24049 output.n71 output.n70 185
R24050 output.n50 output.n49 185
R24051 output.n65 output.n64 185
R24052 output.n63 output.n62 185
R24053 output.n54 output.n53 185
R24054 output.n57 output.n56 185
R24055 output.n105 output.n104 185
R24056 output.n103 output.n102 185
R24057 output.n82 output.n81 185
R24058 output.n97 output.n96 185
R24059 output.n95 output.n94 185
R24060 output.n86 output.n85 185
R24061 output.n89 output.n88 185
R24062 output.n137 output.n136 185
R24063 output.n135 output.n134 185
R24064 output.n114 output.n113 185
R24065 output.n129 output.n128 185
R24066 output.n127 output.n126 185
R24067 output.n118 output.n117 185
R24068 output.n121 output.n120 185
R24069 output.t16 output.n24 147.661
R24070 output.t18 output.n55 147.661
R24071 output.t19 output.n87 147.661
R24072 output.t17 output.n119 147.661
R24073 output.n41 output.n40 104.615
R24074 output.n40 output.n18 104.615
R24075 output.n33 output.n18 104.615
R24076 output.n33 output.n32 104.615
R24077 output.n32 output.n22 104.615
R24078 output.n25 output.n22 104.615
R24079 output.n72 output.n71 104.615
R24080 output.n71 output.n49 104.615
R24081 output.n64 output.n49 104.615
R24082 output.n64 output.n63 104.615
R24083 output.n63 output.n53 104.615
R24084 output.n56 output.n53 104.615
R24085 output.n104 output.n103 104.615
R24086 output.n103 output.n81 104.615
R24087 output.n96 output.n81 104.615
R24088 output.n96 output.n95 104.615
R24089 output.n95 output.n85 104.615
R24090 output.n88 output.n85 104.615
R24091 output.n136 output.n135 104.615
R24092 output.n135 output.n113 104.615
R24093 output.n128 output.n113 104.615
R24094 output.n128 output.n127 104.615
R24095 output.n127 output.n117 104.615
R24096 output.n120 output.n117 104.615
R24097 output.n1 output.t1 77.056
R24098 output.n14 output.t2 76.6694
R24099 output.n1 output.n0 72.7095
R24100 output.n3 output.n2 72.7095
R24101 output.n5 output.n4 72.7095
R24102 output.n7 output.n6 72.7095
R24103 output.n9 output.n8 72.7095
R24104 output.n11 output.n10 72.7095
R24105 output.n13 output.n12 72.7095
R24106 output.n25 output.t16 52.3082
R24107 output.n56 output.t18 52.3082
R24108 output.n88 output.t19 52.3082
R24109 output.n120 output.t17 52.3082
R24110 output.n26 output.n24 15.6674
R24111 output.n57 output.n55 15.6674
R24112 output.n89 output.n87 15.6674
R24113 output.n121 output.n119 15.6674
R24114 output.n27 output.n23 12.8005
R24115 output.n58 output.n54 12.8005
R24116 output.n90 output.n86 12.8005
R24117 output.n122 output.n118 12.8005
R24118 output.n31 output.n30 12.0247
R24119 output.n62 output.n61 12.0247
R24120 output.n94 output.n93 12.0247
R24121 output.n126 output.n125 12.0247
R24122 output.n34 output.n21 11.249
R24123 output.n65 output.n52 11.249
R24124 output.n97 output.n84 11.249
R24125 output.n129 output.n116 11.249
R24126 output.n35 output.n19 10.4732
R24127 output.n66 output.n50 10.4732
R24128 output.n98 output.n82 10.4732
R24129 output.n130 output.n114 10.4732
R24130 output.n39 output.n38 9.69747
R24131 output.n70 output.n69 9.69747
R24132 output.n102 output.n101 9.69747
R24133 output.n134 output.n133 9.69747
R24134 output.n45 output.n44 9.45567
R24135 output.n76 output.n75 9.45567
R24136 output.n108 output.n107 9.45567
R24137 output.n140 output.n139 9.45567
R24138 output.n44 output.n43 9.3005
R24139 output.n17 output.n16 9.3005
R24140 output.n38 output.n37 9.3005
R24141 output.n36 output.n35 9.3005
R24142 output.n21 output.n20 9.3005
R24143 output.n30 output.n29 9.3005
R24144 output.n28 output.n27 9.3005
R24145 output.n75 output.n74 9.3005
R24146 output.n48 output.n47 9.3005
R24147 output.n69 output.n68 9.3005
R24148 output.n67 output.n66 9.3005
R24149 output.n52 output.n51 9.3005
R24150 output.n61 output.n60 9.3005
R24151 output.n59 output.n58 9.3005
R24152 output.n107 output.n106 9.3005
R24153 output.n80 output.n79 9.3005
R24154 output.n101 output.n100 9.3005
R24155 output.n99 output.n98 9.3005
R24156 output.n84 output.n83 9.3005
R24157 output.n93 output.n92 9.3005
R24158 output.n91 output.n90 9.3005
R24159 output.n139 output.n138 9.3005
R24160 output.n112 output.n111 9.3005
R24161 output.n133 output.n132 9.3005
R24162 output.n131 output.n130 9.3005
R24163 output.n116 output.n115 9.3005
R24164 output.n125 output.n124 9.3005
R24165 output.n123 output.n122 9.3005
R24166 output.n42 output.n17 8.92171
R24167 output.n73 output.n48 8.92171
R24168 output.n105 output.n80 8.92171
R24169 output.n137 output.n112 8.92171
R24170 output output.n141 8.15037
R24171 output.n43 output.n15 8.14595
R24172 output.n74 output.n46 8.14595
R24173 output.n106 output.n78 8.14595
R24174 output.n138 output.n110 8.14595
R24175 output.n45 output.n15 5.81868
R24176 output.n76 output.n46 5.81868
R24177 output.n108 output.n78 5.81868
R24178 output.n140 output.n110 5.81868
R24179 output.n43 output.n42 5.04292
R24180 output.n74 output.n73 5.04292
R24181 output.n106 output.n105 5.04292
R24182 output.n138 output.n137 5.04292
R24183 output.n28 output.n24 4.38594
R24184 output.n59 output.n55 4.38594
R24185 output.n91 output.n87 4.38594
R24186 output.n123 output.n119 4.38594
R24187 output.n39 output.n17 4.26717
R24188 output.n70 output.n48 4.26717
R24189 output.n102 output.n80 4.26717
R24190 output.n134 output.n112 4.26717
R24191 output.n0 output.t11 3.9605
R24192 output.n0 output.t9 3.9605
R24193 output.n2 output.t0 3.9605
R24194 output.n2 output.t3 3.9605
R24195 output.n4 output.t5 3.9605
R24196 output.n4 output.t13 3.9605
R24197 output.n6 output.t15 3.9605
R24198 output.n6 output.t6 3.9605
R24199 output.n8 output.t7 3.9605
R24200 output.n8 output.t12 3.9605
R24201 output.n10 output.t14 3.9605
R24202 output.n10 output.t4 3.9605
R24203 output.n12 output.t10 3.9605
R24204 output.n12 output.t8 3.9605
R24205 output.n38 output.n19 3.49141
R24206 output.n69 output.n50 3.49141
R24207 output.n101 output.n82 3.49141
R24208 output.n133 output.n114 3.49141
R24209 output.n35 output.n34 2.71565
R24210 output.n66 output.n65 2.71565
R24211 output.n98 output.n97 2.71565
R24212 output.n130 output.n129 2.71565
R24213 output.n31 output.n21 1.93989
R24214 output.n62 output.n52 1.93989
R24215 output.n94 output.n84 1.93989
R24216 output.n126 output.n116 1.93989
R24217 output.n30 output.n23 1.16414
R24218 output.n61 output.n54 1.16414
R24219 output.n93 output.n86 1.16414
R24220 output.n125 output.n118 1.16414
R24221 output.n141 output.n109 0.962709
R24222 output.n109 output.n77 0.962709
R24223 output.n27 output.n26 0.388379
R24224 output.n58 output.n57 0.388379
R24225 output.n90 output.n89 0.388379
R24226 output.n122 output.n121 0.388379
R24227 output.n14 output.n13 0.387128
R24228 output.n13 output.n11 0.387128
R24229 output.n11 output.n9 0.387128
R24230 output.n9 output.n7 0.387128
R24231 output.n7 output.n5 0.387128
R24232 output.n5 output.n3 0.387128
R24233 output.n3 output.n1 0.387128
R24234 output.n44 output.n16 0.155672
R24235 output.n37 output.n16 0.155672
R24236 output.n37 output.n36 0.155672
R24237 output.n36 output.n20 0.155672
R24238 output.n29 output.n20 0.155672
R24239 output.n29 output.n28 0.155672
R24240 output.n75 output.n47 0.155672
R24241 output.n68 output.n47 0.155672
R24242 output.n68 output.n67 0.155672
R24243 output.n67 output.n51 0.155672
R24244 output.n60 output.n51 0.155672
R24245 output.n60 output.n59 0.155672
R24246 output.n107 output.n79 0.155672
R24247 output.n100 output.n79 0.155672
R24248 output.n100 output.n99 0.155672
R24249 output.n99 output.n83 0.155672
R24250 output.n92 output.n83 0.155672
R24251 output.n92 output.n91 0.155672
R24252 output.n139 output.n111 0.155672
R24253 output.n132 output.n111 0.155672
R24254 output.n132 output.n131 0.155672
R24255 output.n131 output.n115 0.155672
R24256 output.n124 output.n115 0.155672
R24257 output.n124 output.n123 0.155672
R24258 output output.n14 0.126227
R24259 diffpairibias.n0 diffpairibias.t18 436.822
R24260 diffpairibias.n21 diffpairibias.t19 435.479
R24261 diffpairibias.n20 diffpairibias.t16 435.479
R24262 diffpairibias.n19 diffpairibias.t17 435.479
R24263 diffpairibias.n18 diffpairibias.t21 435.479
R24264 diffpairibias.n0 diffpairibias.t22 435.479
R24265 diffpairibias.n1 diffpairibias.t20 435.479
R24266 diffpairibias.n2 diffpairibias.t23 435.479
R24267 diffpairibias.n10 diffpairibias.t0 377.536
R24268 diffpairibias.n10 diffpairibias.t8 376.193
R24269 diffpairibias.n11 diffpairibias.t10 376.193
R24270 diffpairibias.n12 diffpairibias.t6 376.193
R24271 diffpairibias.n13 diffpairibias.t2 376.193
R24272 diffpairibias.n14 diffpairibias.t12 376.193
R24273 diffpairibias.n15 diffpairibias.t4 376.193
R24274 diffpairibias.n16 diffpairibias.t14 376.193
R24275 diffpairibias.n3 diffpairibias.t1 113.368
R24276 diffpairibias.n3 diffpairibias.t9 112.698
R24277 diffpairibias.n4 diffpairibias.t11 112.698
R24278 diffpairibias.n5 diffpairibias.t7 112.698
R24279 diffpairibias.n6 diffpairibias.t3 112.698
R24280 diffpairibias.n7 diffpairibias.t13 112.698
R24281 diffpairibias.n8 diffpairibias.t5 112.698
R24282 diffpairibias.n9 diffpairibias.t15 112.698
R24283 diffpairibias.n17 diffpairibias.n16 4.77242
R24284 diffpairibias.n17 diffpairibias.n9 4.30807
R24285 diffpairibias.n18 diffpairibias.n17 4.13945
R24286 diffpairibias.n16 diffpairibias.n15 1.34352
R24287 diffpairibias.n15 diffpairibias.n14 1.34352
R24288 diffpairibias.n14 diffpairibias.n13 1.34352
R24289 diffpairibias.n13 diffpairibias.n12 1.34352
R24290 diffpairibias.n12 diffpairibias.n11 1.34352
R24291 diffpairibias.n11 diffpairibias.n10 1.34352
R24292 diffpairibias.n2 diffpairibias.n1 1.34352
R24293 diffpairibias.n1 diffpairibias.n0 1.34352
R24294 diffpairibias.n19 diffpairibias.n18 1.34352
R24295 diffpairibias.n20 diffpairibias.n19 1.34352
R24296 diffpairibias.n21 diffpairibias.n20 1.34352
R24297 diffpairibias.n22 diffpairibias.n21 0.862419
R24298 diffpairibias diffpairibias.n22 0.684875
R24299 diffpairibias.n9 diffpairibias.n8 0.672012
R24300 diffpairibias.n8 diffpairibias.n7 0.672012
R24301 diffpairibias.n7 diffpairibias.n6 0.672012
R24302 diffpairibias.n6 diffpairibias.n5 0.672012
R24303 diffpairibias.n5 diffpairibias.n4 0.672012
R24304 diffpairibias.n4 diffpairibias.n3 0.672012
R24305 diffpairibias.n22 diffpairibias.n2 0.190907
R24306 minus.n27 minus.t20 436.949
R24307 minus.n5 minus.t11 436.949
R24308 minus.n42 minus.t17 415.966
R24309 minus.n41 minus.t10 415.966
R24310 minus.n23 minus.t5 415.966
R24311 minus.n35 minus.t13 415.966
R24312 minus.n34 minus.t9 415.966
R24313 minus.n26 minus.t19 415.966
R24314 minus.n28 minus.t7 415.966
R24315 minus.n6 minus.t14 415.966
R24316 minus.n8 minus.t8 415.966
R24317 minus.n12 minus.t12 415.966
R24318 minus.n13 minus.t18 415.966
R24319 minus.n1 minus.t15 415.966
R24320 minus.n19 minus.t16 415.966
R24321 minus.n20 minus.t6 415.966
R24322 minus.n48 minus.t1 243.255
R24323 minus.n47 minus.n45 224.169
R24324 minus.n47 minus.n46 223.454
R24325 minus.n30 minus.n29 161.3
R24326 minus.n31 minus.n26 161.3
R24327 minus.n33 minus.n32 161.3
R24328 minus.n34 minus.n25 161.3
R24329 minus.n35 minus.n24 161.3
R24330 minus.n37 minus.n36 161.3
R24331 minus.n38 minus.n23 161.3
R24332 minus.n40 minus.n39 161.3
R24333 minus.n41 minus.n22 161.3
R24334 minus.n43 minus.n42 161.3
R24335 minus.n21 minus.n20 161.3
R24336 minus.n19 minus.n0 161.3
R24337 minus.n18 minus.n17 161.3
R24338 minus.n16 minus.n1 161.3
R24339 minus.n15 minus.n14 161.3
R24340 minus.n13 minus.n2 161.3
R24341 minus.n12 minus.n11 161.3
R24342 minus.n10 minus.n3 161.3
R24343 minus.n9 minus.n8 161.3
R24344 minus.n7 minus.n4 161.3
R24345 minus.n30 minus.n27 70.4033
R24346 minus.n5 minus.n4 70.4033
R24347 minus.n42 minus.n41 48.2005
R24348 minus.n35 minus.n34 48.2005
R24349 minus.n13 minus.n12 48.2005
R24350 minus.n20 minus.n19 48.2005
R24351 minus.n40 minus.n23 37.246
R24352 minus.n29 minus.n26 37.246
R24353 minus.n8 minus.n7 37.246
R24354 minus.n18 minus.n1 37.246
R24355 minus.n36 minus.n23 35.7853
R24356 minus.n33 minus.n26 35.7853
R24357 minus.n8 minus.n3 35.7853
R24358 minus.n14 minus.n1 35.7853
R24359 minus.n44 minus.n43 28.7903
R24360 minus.n28 minus.n27 20.9576
R24361 minus.n6 minus.n5 20.9576
R24362 minus.n46 minus.t3 19.8005
R24363 minus.n46 minus.t4 19.8005
R24364 minus.n45 minus.t2 19.8005
R24365 minus.n45 minus.t0 19.8005
R24366 minus.n36 minus.n35 12.4157
R24367 minus.n34 minus.n33 12.4157
R24368 minus.n12 minus.n3 12.4157
R24369 minus.n14 minus.n13 12.4157
R24370 minus minus.n49 12.1137
R24371 minus.n44 minus.n21 11.9759
R24372 minus.n41 minus.n40 10.955
R24373 minus.n29 minus.n28 10.955
R24374 minus.n7 minus.n6 10.955
R24375 minus.n19 minus.n18 10.955
R24376 minus.n49 minus.n48 4.80222
R24377 minus.n49 minus.n44 0.972091
R24378 minus.n48 minus.n47 0.716017
R24379 minus.n43 minus.n22 0.189894
R24380 minus.n39 minus.n22 0.189894
R24381 minus.n39 minus.n38 0.189894
R24382 minus.n38 minus.n37 0.189894
R24383 minus.n37 minus.n24 0.189894
R24384 minus.n25 minus.n24 0.189894
R24385 minus.n32 minus.n25 0.189894
R24386 minus.n32 minus.n31 0.189894
R24387 minus.n31 minus.n30 0.189894
R24388 minus.n9 minus.n4 0.189894
R24389 minus.n10 minus.n9 0.189894
R24390 minus.n11 minus.n10 0.189894
R24391 minus.n11 minus.n2 0.189894
R24392 minus.n15 minus.n2 0.189894
R24393 minus.n16 minus.n15 0.189894
R24394 minus.n17 minus.n16 0.189894
R24395 minus.n17 minus.n0 0.189894
R24396 minus.n21 minus.n0 0.189894
R24397 outputibias.n27 outputibias.n1 289.615
R24398 outputibias.n58 outputibias.n32 289.615
R24399 outputibias.n90 outputibias.n64 289.615
R24400 outputibias.n122 outputibias.n96 289.615
R24401 outputibias.n28 outputibias.n27 185
R24402 outputibias.n26 outputibias.n25 185
R24403 outputibias.n5 outputibias.n4 185
R24404 outputibias.n20 outputibias.n19 185
R24405 outputibias.n18 outputibias.n17 185
R24406 outputibias.n9 outputibias.n8 185
R24407 outputibias.n12 outputibias.n11 185
R24408 outputibias.n59 outputibias.n58 185
R24409 outputibias.n57 outputibias.n56 185
R24410 outputibias.n36 outputibias.n35 185
R24411 outputibias.n51 outputibias.n50 185
R24412 outputibias.n49 outputibias.n48 185
R24413 outputibias.n40 outputibias.n39 185
R24414 outputibias.n43 outputibias.n42 185
R24415 outputibias.n91 outputibias.n90 185
R24416 outputibias.n89 outputibias.n88 185
R24417 outputibias.n68 outputibias.n67 185
R24418 outputibias.n83 outputibias.n82 185
R24419 outputibias.n81 outputibias.n80 185
R24420 outputibias.n72 outputibias.n71 185
R24421 outputibias.n75 outputibias.n74 185
R24422 outputibias.n123 outputibias.n122 185
R24423 outputibias.n121 outputibias.n120 185
R24424 outputibias.n100 outputibias.n99 185
R24425 outputibias.n115 outputibias.n114 185
R24426 outputibias.n113 outputibias.n112 185
R24427 outputibias.n104 outputibias.n103 185
R24428 outputibias.n107 outputibias.n106 185
R24429 outputibias.n0 outputibias.t8 178.945
R24430 outputibias.n133 outputibias.t11 177.018
R24431 outputibias.n132 outputibias.t9 177.018
R24432 outputibias.n0 outputibias.t10 177.018
R24433 outputibias.t7 outputibias.n10 147.661
R24434 outputibias.t1 outputibias.n41 147.661
R24435 outputibias.t3 outputibias.n73 147.661
R24436 outputibias.t5 outputibias.n105 147.661
R24437 outputibias.n128 outputibias.t6 132.363
R24438 outputibias.n128 outputibias.t0 130.436
R24439 outputibias.n129 outputibias.t2 130.436
R24440 outputibias.n130 outputibias.t4 130.436
R24441 outputibias.n27 outputibias.n26 104.615
R24442 outputibias.n26 outputibias.n4 104.615
R24443 outputibias.n19 outputibias.n4 104.615
R24444 outputibias.n19 outputibias.n18 104.615
R24445 outputibias.n18 outputibias.n8 104.615
R24446 outputibias.n11 outputibias.n8 104.615
R24447 outputibias.n58 outputibias.n57 104.615
R24448 outputibias.n57 outputibias.n35 104.615
R24449 outputibias.n50 outputibias.n35 104.615
R24450 outputibias.n50 outputibias.n49 104.615
R24451 outputibias.n49 outputibias.n39 104.615
R24452 outputibias.n42 outputibias.n39 104.615
R24453 outputibias.n90 outputibias.n89 104.615
R24454 outputibias.n89 outputibias.n67 104.615
R24455 outputibias.n82 outputibias.n67 104.615
R24456 outputibias.n82 outputibias.n81 104.615
R24457 outputibias.n81 outputibias.n71 104.615
R24458 outputibias.n74 outputibias.n71 104.615
R24459 outputibias.n122 outputibias.n121 104.615
R24460 outputibias.n121 outputibias.n99 104.615
R24461 outputibias.n114 outputibias.n99 104.615
R24462 outputibias.n114 outputibias.n113 104.615
R24463 outputibias.n113 outputibias.n103 104.615
R24464 outputibias.n106 outputibias.n103 104.615
R24465 outputibias.n63 outputibias.n31 95.6354
R24466 outputibias.n63 outputibias.n62 94.6732
R24467 outputibias.n95 outputibias.n94 94.6732
R24468 outputibias.n127 outputibias.n126 94.6732
R24469 outputibias.n11 outputibias.t7 52.3082
R24470 outputibias.n42 outputibias.t1 52.3082
R24471 outputibias.n74 outputibias.t3 52.3082
R24472 outputibias.n106 outputibias.t5 52.3082
R24473 outputibias.n12 outputibias.n10 15.6674
R24474 outputibias.n43 outputibias.n41 15.6674
R24475 outputibias.n75 outputibias.n73 15.6674
R24476 outputibias.n107 outputibias.n105 15.6674
R24477 outputibias.n13 outputibias.n9 12.8005
R24478 outputibias.n44 outputibias.n40 12.8005
R24479 outputibias.n76 outputibias.n72 12.8005
R24480 outputibias.n108 outputibias.n104 12.8005
R24481 outputibias.n17 outputibias.n16 12.0247
R24482 outputibias.n48 outputibias.n47 12.0247
R24483 outputibias.n80 outputibias.n79 12.0247
R24484 outputibias.n112 outputibias.n111 12.0247
R24485 outputibias.n20 outputibias.n7 11.249
R24486 outputibias.n51 outputibias.n38 11.249
R24487 outputibias.n83 outputibias.n70 11.249
R24488 outputibias.n115 outputibias.n102 11.249
R24489 outputibias.n21 outputibias.n5 10.4732
R24490 outputibias.n52 outputibias.n36 10.4732
R24491 outputibias.n84 outputibias.n68 10.4732
R24492 outputibias.n116 outputibias.n100 10.4732
R24493 outputibias.n25 outputibias.n24 9.69747
R24494 outputibias.n56 outputibias.n55 9.69747
R24495 outputibias.n88 outputibias.n87 9.69747
R24496 outputibias.n120 outputibias.n119 9.69747
R24497 outputibias.n31 outputibias.n30 9.45567
R24498 outputibias.n62 outputibias.n61 9.45567
R24499 outputibias.n94 outputibias.n93 9.45567
R24500 outputibias.n126 outputibias.n125 9.45567
R24501 outputibias.n30 outputibias.n29 9.3005
R24502 outputibias.n3 outputibias.n2 9.3005
R24503 outputibias.n24 outputibias.n23 9.3005
R24504 outputibias.n22 outputibias.n21 9.3005
R24505 outputibias.n7 outputibias.n6 9.3005
R24506 outputibias.n16 outputibias.n15 9.3005
R24507 outputibias.n14 outputibias.n13 9.3005
R24508 outputibias.n61 outputibias.n60 9.3005
R24509 outputibias.n34 outputibias.n33 9.3005
R24510 outputibias.n55 outputibias.n54 9.3005
R24511 outputibias.n53 outputibias.n52 9.3005
R24512 outputibias.n38 outputibias.n37 9.3005
R24513 outputibias.n47 outputibias.n46 9.3005
R24514 outputibias.n45 outputibias.n44 9.3005
R24515 outputibias.n93 outputibias.n92 9.3005
R24516 outputibias.n66 outputibias.n65 9.3005
R24517 outputibias.n87 outputibias.n86 9.3005
R24518 outputibias.n85 outputibias.n84 9.3005
R24519 outputibias.n70 outputibias.n69 9.3005
R24520 outputibias.n79 outputibias.n78 9.3005
R24521 outputibias.n77 outputibias.n76 9.3005
R24522 outputibias.n125 outputibias.n124 9.3005
R24523 outputibias.n98 outputibias.n97 9.3005
R24524 outputibias.n119 outputibias.n118 9.3005
R24525 outputibias.n117 outputibias.n116 9.3005
R24526 outputibias.n102 outputibias.n101 9.3005
R24527 outputibias.n111 outputibias.n110 9.3005
R24528 outputibias.n109 outputibias.n108 9.3005
R24529 outputibias.n28 outputibias.n3 8.92171
R24530 outputibias.n59 outputibias.n34 8.92171
R24531 outputibias.n91 outputibias.n66 8.92171
R24532 outputibias.n123 outputibias.n98 8.92171
R24533 outputibias.n29 outputibias.n1 8.14595
R24534 outputibias.n60 outputibias.n32 8.14595
R24535 outputibias.n92 outputibias.n64 8.14595
R24536 outputibias.n124 outputibias.n96 8.14595
R24537 outputibias.n31 outputibias.n1 5.81868
R24538 outputibias.n62 outputibias.n32 5.81868
R24539 outputibias.n94 outputibias.n64 5.81868
R24540 outputibias.n126 outputibias.n96 5.81868
R24541 outputibias.n131 outputibias.n130 5.20947
R24542 outputibias.n29 outputibias.n28 5.04292
R24543 outputibias.n60 outputibias.n59 5.04292
R24544 outputibias.n92 outputibias.n91 5.04292
R24545 outputibias.n124 outputibias.n123 5.04292
R24546 outputibias.n131 outputibias.n127 4.42209
R24547 outputibias.n14 outputibias.n10 4.38594
R24548 outputibias.n45 outputibias.n41 4.38594
R24549 outputibias.n77 outputibias.n73 4.38594
R24550 outputibias.n109 outputibias.n105 4.38594
R24551 outputibias.n132 outputibias.n131 4.28454
R24552 outputibias.n25 outputibias.n3 4.26717
R24553 outputibias.n56 outputibias.n34 4.26717
R24554 outputibias.n88 outputibias.n66 4.26717
R24555 outputibias.n120 outputibias.n98 4.26717
R24556 outputibias.n24 outputibias.n5 3.49141
R24557 outputibias.n55 outputibias.n36 3.49141
R24558 outputibias.n87 outputibias.n68 3.49141
R24559 outputibias.n119 outputibias.n100 3.49141
R24560 outputibias.n21 outputibias.n20 2.71565
R24561 outputibias.n52 outputibias.n51 2.71565
R24562 outputibias.n84 outputibias.n83 2.71565
R24563 outputibias.n116 outputibias.n115 2.71565
R24564 outputibias.n17 outputibias.n7 1.93989
R24565 outputibias.n48 outputibias.n38 1.93989
R24566 outputibias.n80 outputibias.n70 1.93989
R24567 outputibias.n112 outputibias.n102 1.93989
R24568 outputibias.n130 outputibias.n129 1.9266
R24569 outputibias.n129 outputibias.n128 1.9266
R24570 outputibias.n133 outputibias.n132 1.92658
R24571 outputibias.n134 outputibias.n133 1.29913
R24572 outputibias.n16 outputibias.n9 1.16414
R24573 outputibias.n47 outputibias.n40 1.16414
R24574 outputibias.n79 outputibias.n72 1.16414
R24575 outputibias.n111 outputibias.n104 1.16414
R24576 outputibias.n127 outputibias.n95 0.962709
R24577 outputibias.n95 outputibias.n63 0.962709
R24578 outputibias.n13 outputibias.n12 0.388379
R24579 outputibias.n44 outputibias.n43 0.388379
R24580 outputibias.n76 outputibias.n75 0.388379
R24581 outputibias.n108 outputibias.n107 0.388379
R24582 outputibias.n134 outputibias.n0 0.337251
R24583 outputibias outputibias.n134 0.302375
R24584 outputibias.n30 outputibias.n2 0.155672
R24585 outputibias.n23 outputibias.n2 0.155672
R24586 outputibias.n23 outputibias.n22 0.155672
R24587 outputibias.n22 outputibias.n6 0.155672
R24588 outputibias.n15 outputibias.n6 0.155672
R24589 outputibias.n15 outputibias.n14 0.155672
R24590 outputibias.n61 outputibias.n33 0.155672
R24591 outputibias.n54 outputibias.n33 0.155672
R24592 outputibias.n54 outputibias.n53 0.155672
R24593 outputibias.n53 outputibias.n37 0.155672
R24594 outputibias.n46 outputibias.n37 0.155672
R24595 outputibias.n46 outputibias.n45 0.155672
R24596 outputibias.n93 outputibias.n65 0.155672
R24597 outputibias.n86 outputibias.n65 0.155672
R24598 outputibias.n86 outputibias.n85 0.155672
R24599 outputibias.n85 outputibias.n69 0.155672
R24600 outputibias.n78 outputibias.n69 0.155672
R24601 outputibias.n78 outputibias.n77 0.155672
R24602 outputibias.n125 outputibias.n97 0.155672
R24603 outputibias.n118 outputibias.n97 0.155672
R24604 outputibias.n118 outputibias.n117 0.155672
R24605 outputibias.n117 outputibias.n101 0.155672
R24606 outputibias.n110 outputibias.n101 0.155672
R24607 outputibias.n110 outputibias.n109 0.155672
C0 plus commonsourceibias 0.268404f
C1 output outputibias 2.34152f
C2 vdd output 7.23429f
C3 CSoutput output 6.13881f
C4 CSoutput outputibias 0.032386f
C5 vdd CSoutput 0.140616p
C6 minus diffpairibias 1.62e-19
C7 commonsourceibias output 0.006808f
C8 vdd plus 0.0849f
C9 CSoutput minus 3.23017f
C10 plus diffpairibias 2.39e-19
C11 commonsourceibias outputibias 0.003832f
C12 CSoutput plus 0.849039f
C13 vdd commonsourceibias 0.004218f
C14 commonsourceibias diffpairibias 0.06482f
C15 minus plus 8.922501f
C16 CSoutput commonsourceibias 66.33679f
C17 minus commonsourceibias 0.314643f
C18 diffpairibias gnd 48.979836f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.222623p
C22 plus gnd 29.663897f
C23 minus gnd 26.37718f
C24 CSoutput gnd 0.143502p
C25 vdd gnd 0.439059p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t1 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t3 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t2 gnd 0.108319f
C162 outputibias.t0 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 minus.n0 gnd 0.030236f
C174 minus.t15 gnd 0.305475f
C175 minus.n1 gnd 0.141231f
C176 minus.n2 gnd 0.030236f
C177 minus.n3 gnd 0.006861f
C178 minus.n4 gnd 0.096268f
C179 minus.t11 gnd 0.312107f
C180 minus.n5 gnd 0.13165f
C181 minus.t14 gnd 0.305475f
C182 minus.n6 gnd 0.13946f
C183 minus.n7 gnd 0.006861f
C184 minus.t8 gnd 0.305475f
C185 minus.n8 gnd 0.141231f
C186 minus.n9 gnd 0.030236f
C187 minus.n10 gnd 0.030236f
C188 minus.n11 gnd 0.030236f
C189 minus.t12 gnd 0.305475f
C190 minus.n12 gnd 0.139646f
C191 minus.t18 gnd 0.305475f
C192 minus.n13 gnd 0.139646f
C193 minus.n14 gnd 0.006861f
C194 minus.n15 gnd 0.030236f
C195 minus.n16 gnd 0.030236f
C196 minus.n17 gnd 0.030236f
C197 minus.n18 gnd 0.006861f
C198 minus.t16 gnd 0.305475f
C199 minus.n19 gnd 0.13946f
C200 minus.t6 gnd 0.305475f
C201 minus.n20 gnd 0.138062f
C202 minus.n21 gnd 0.341781f
C203 minus.n22 gnd 0.030236f
C204 minus.t17 gnd 0.305475f
C205 minus.t10 gnd 0.305475f
C206 minus.t5 gnd 0.305475f
C207 minus.n23 gnd 0.141231f
C208 minus.n24 gnd 0.030236f
C209 minus.t13 gnd 0.305475f
C210 minus.t9 gnd 0.305475f
C211 minus.n25 gnd 0.030236f
C212 minus.t19 gnd 0.305475f
C213 minus.n26 gnd 0.141231f
C214 minus.t20 gnd 0.312107f
C215 minus.n27 gnd 0.13165f
C216 minus.t7 gnd 0.305475f
C217 minus.n28 gnd 0.13946f
C218 minus.n29 gnd 0.006861f
C219 minus.n30 gnd 0.096268f
C220 minus.n31 gnd 0.030236f
C221 minus.n32 gnd 0.030236f
C222 minus.n33 gnd 0.006861f
C223 minus.n34 gnd 0.139646f
C224 minus.n35 gnd 0.139646f
C225 minus.n36 gnd 0.006861f
C226 minus.n37 gnd 0.030236f
C227 minus.n38 gnd 0.030236f
C228 minus.n39 gnd 0.030236f
C229 minus.n40 gnd 0.006861f
C230 minus.n41 gnd 0.13946f
C231 minus.n42 gnd 0.138062f
C232 minus.n43 gnd 0.813811f
C233 minus.n44 gnd 1.25224f
C234 minus.t2 gnd 0.009321f
C235 minus.t0 gnd 0.009321f
C236 minus.n45 gnd 0.030649f
C237 minus.t3 gnd 0.009321f
C238 minus.t4 gnd 0.009321f
C239 minus.n46 gnd 0.03023f
C240 minus.n47 gnd 0.257996f
C241 minus.t1 gnd 0.051879f
C242 minus.n48 gnd 0.140786f
C243 minus.n49 gnd 2.30203f
C244 diffpairibias.t18 gnd 0.087401f
C245 diffpairibias.t22 gnd 0.087239f
C246 diffpairibias.n0 gnd 0.102784f
C247 diffpairibias.t20 gnd 0.087239f
C248 diffpairibias.n1 gnd 0.050171f
C249 diffpairibias.t23 gnd 0.087239f
C250 diffpairibias.n2 gnd 0.039841f
C251 diffpairibias.t1 gnd 0.083757f
C252 diffpairibias.t9 gnd 0.083392f
C253 diffpairibias.n3 gnd 0.131682f
C254 diffpairibias.t11 gnd 0.083392f
C255 diffpairibias.n4 gnd 0.07027f
C256 diffpairibias.t7 gnd 0.083392f
C257 diffpairibias.n5 gnd 0.07027f
C258 diffpairibias.t3 gnd 0.083392f
C259 diffpairibias.n6 gnd 0.07027f
C260 diffpairibias.t13 gnd 0.083392f
C261 diffpairibias.n7 gnd 0.07027f
C262 diffpairibias.t5 gnd 0.083392f
C263 diffpairibias.n8 gnd 0.07027f
C264 diffpairibias.t15 gnd 0.083392f
C265 diffpairibias.n9 gnd 0.099771f
C266 diffpairibias.t0 gnd 0.08427f
C267 diffpairibias.t8 gnd 0.084123f
C268 diffpairibias.n10 gnd 0.091784f
C269 diffpairibias.t10 gnd 0.084123f
C270 diffpairibias.n11 gnd 0.050681f
C271 diffpairibias.t6 gnd 0.084123f
C272 diffpairibias.n12 gnd 0.050681f
C273 diffpairibias.t2 gnd 0.084123f
C274 diffpairibias.n13 gnd 0.050681f
C275 diffpairibias.t12 gnd 0.084123f
C276 diffpairibias.n14 gnd 0.050681f
C277 diffpairibias.t4 gnd 0.084123f
C278 diffpairibias.n15 gnd 0.050681f
C279 diffpairibias.t14 gnd 0.084123f
C280 diffpairibias.n16 gnd 0.059977f
C281 diffpairibias.n17 gnd 0.226448f
C282 diffpairibias.t21 gnd 0.087239f
C283 diffpairibias.n18 gnd 0.050181f
C284 diffpairibias.t17 gnd 0.087239f
C285 diffpairibias.n19 gnd 0.050171f
C286 diffpairibias.t16 gnd 0.087239f
C287 diffpairibias.n20 gnd 0.050171f
C288 diffpairibias.t19 gnd 0.087239f
C289 diffpairibias.n21 gnd 0.045859f
C290 diffpairibias.n22 gnd 0.046268f
C291 output.t1 gnd 0.464308f
C292 output.t11 gnd 0.044422f
C293 output.t9 gnd 0.044422f
C294 output.n0 gnd 0.364624f
C295 output.n1 gnd 0.614102f
C296 output.t0 gnd 0.044422f
C297 output.t3 gnd 0.044422f
C298 output.n2 gnd 0.364624f
C299 output.n3 gnd 0.350265f
C300 output.t5 gnd 0.044422f
C301 output.t13 gnd 0.044422f
C302 output.n4 gnd 0.364624f
C303 output.n5 gnd 0.350265f
C304 output.t15 gnd 0.044422f
C305 output.t6 gnd 0.044422f
C306 output.n6 gnd 0.364624f
C307 output.n7 gnd 0.350265f
C308 output.t7 gnd 0.044422f
C309 output.t12 gnd 0.044422f
C310 output.n8 gnd 0.364624f
C311 output.n9 gnd 0.350265f
C312 output.t14 gnd 0.044422f
C313 output.t4 gnd 0.044422f
C314 output.n10 gnd 0.364624f
C315 output.n11 gnd 0.350265f
C316 output.t10 gnd 0.044422f
C317 output.t8 gnd 0.044422f
C318 output.n12 gnd 0.364624f
C319 output.n13 gnd 0.350265f
C320 output.t2 gnd 0.462979f
C321 output.n14 gnd 0.28994f
C322 output.n15 gnd 0.015803f
C323 output.n16 gnd 0.011243f
C324 output.n17 gnd 0.006041f
C325 output.n18 gnd 0.01428f
C326 output.n19 gnd 0.006397f
C327 output.n20 gnd 0.011243f
C328 output.n21 gnd 0.006041f
C329 output.n22 gnd 0.01428f
C330 output.n23 gnd 0.006397f
C331 output.n24 gnd 0.048111f
C332 output.t16 gnd 0.023274f
C333 output.n25 gnd 0.01071f
C334 output.n26 gnd 0.008435f
C335 output.n27 gnd 0.006041f
C336 output.n28 gnd 0.267512f
C337 output.n29 gnd 0.011243f
C338 output.n30 gnd 0.006041f
C339 output.n31 gnd 0.006397f
C340 output.n32 gnd 0.01428f
C341 output.n33 gnd 0.01428f
C342 output.n34 gnd 0.006397f
C343 output.n35 gnd 0.006041f
C344 output.n36 gnd 0.011243f
C345 output.n37 gnd 0.011243f
C346 output.n38 gnd 0.006041f
C347 output.n39 gnd 0.006397f
C348 output.n40 gnd 0.01428f
C349 output.n41 gnd 0.030913f
C350 output.n42 gnd 0.006397f
C351 output.n43 gnd 0.006041f
C352 output.n44 gnd 0.025987f
C353 output.n45 gnd 0.097665f
C354 output.n46 gnd 0.015803f
C355 output.n47 gnd 0.011243f
C356 output.n48 gnd 0.006041f
C357 output.n49 gnd 0.01428f
C358 output.n50 gnd 0.006397f
C359 output.n51 gnd 0.011243f
C360 output.n52 gnd 0.006041f
C361 output.n53 gnd 0.01428f
C362 output.n54 gnd 0.006397f
C363 output.n55 gnd 0.048111f
C364 output.t18 gnd 0.023274f
C365 output.n56 gnd 0.01071f
C366 output.n57 gnd 0.008435f
C367 output.n58 gnd 0.006041f
C368 output.n59 gnd 0.267512f
C369 output.n60 gnd 0.011243f
C370 output.n61 gnd 0.006041f
C371 output.n62 gnd 0.006397f
C372 output.n63 gnd 0.01428f
C373 output.n64 gnd 0.01428f
C374 output.n65 gnd 0.006397f
C375 output.n66 gnd 0.006041f
C376 output.n67 gnd 0.011243f
C377 output.n68 gnd 0.011243f
C378 output.n69 gnd 0.006041f
C379 output.n70 gnd 0.006397f
C380 output.n71 gnd 0.01428f
C381 output.n72 gnd 0.030913f
C382 output.n73 gnd 0.006397f
C383 output.n74 gnd 0.006041f
C384 output.n75 gnd 0.025987f
C385 output.n76 gnd 0.09306f
C386 output.n77 gnd 1.65264f
C387 output.n78 gnd 0.015803f
C388 output.n79 gnd 0.011243f
C389 output.n80 gnd 0.006041f
C390 output.n81 gnd 0.01428f
C391 output.n82 gnd 0.006397f
C392 output.n83 gnd 0.011243f
C393 output.n84 gnd 0.006041f
C394 output.n85 gnd 0.01428f
C395 output.n86 gnd 0.006397f
C396 output.n87 gnd 0.048111f
C397 output.t19 gnd 0.023274f
C398 output.n88 gnd 0.01071f
C399 output.n89 gnd 0.008435f
C400 output.n90 gnd 0.006041f
C401 output.n91 gnd 0.267512f
C402 output.n92 gnd 0.011243f
C403 output.n93 gnd 0.006041f
C404 output.n94 gnd 0.006397f
C405 output.n95 gnd 0.01428f
C406 output.n96 gnd 0.01428f
C407 output.n97 gnd 0.006397f
C408 output.n98 gnd 0.006041f
C409 output.n99 gnd 0.011243f
C410 output.n100 gnd 0.011243f
C411 output.n101 gnd 0.006041f
C412 output.n102 gnd 0.006397f
C413 output.n103 gnd 0.01428f
C414 output.n104 gnd 0.030913f
C415 output.n105 gnd 0.006397f
C416 output.n106 gnd 0.006041f
C417 output.n107 gnd 0.025987f
C418 output.n108 gnd 0.09306f
C419 output.n109 gnd 0.713089f
C420 output.n110 gnd 0.015803f
C421 output.n111 gnd 0.011243f
C422 output.n112 gnd 0.006041f
C423 output.n113 gnd 0.01428f
C424 output.n114 gnd 0.006397f
C425 output.n115 gnd 0.011243f
C426 output.n116 gnd 0.006041f
C427 output.n117 gnd 0.01428f
C428 output.n118 gnd 0.006397f
C429 output.n119 gnd 0.048111f
C430 output.t17 gnd 0.023274f
C431 output.n120 gnd 0.01071f
C432 output.n121 gnd 0.008435f
C433 output.n122 gnd 0.006041f
C434 output.n123 gnd 0.267512f
C435 output.n124 gnd 0.011243f
C436 output.n125 gnd 0.006041f
C437 output.n126 gnd 0.006397f
C438 output.n127 gnd 0.01428f
C439 output.n128 gnd 0.01428f
C440 output.n129 gnd 0.006397f
C441 output.n130 gnd 0.006041f
C442 output.n131 gnd 0.011243f
C443 output.n132 gnd 0.011243f
C444 output.n133 gnd 0.006041f
C445 output.n134 gnd 0.006397f
C446 output.n135 gnd 0.01428f
C447 output.n136 gnd 0.030913f
C448 output.n137 gnd 0.006397f
C449 output.n138 gnd 0.006041f
C450 output.n139 gnd 0.025987f
C451 output.n140 gnd 0.09306f
C452 output.n141 gnd 1.67353f
C453 a_n2903_n3924.n0 gnd 2.07284f
C454 a_n2903_n3924.t16 gnd 0.094832f
C455 a_n2903_n3924.t14 gnd 0.985605f
C456 a_n2903_n3924.n1 gnd 0.334506f
C457 a_n2903_n3924.t39 gnd 1.22783f
C458 a_n2903_n3924.t37 gnd 0.985605f
C459 a_n2903_n3924.n2 gnd 0.334506f
C460 a_n2903_n3924.t7 gnd 0.094832f
C461 a_n2903_n3924.t0 gnd 0.094832f
C462 a_n2903_n3924.n3 gnd 0.774508f
C463 a_n2903_n3924.n4 gnd 0.314114f
C464 a_n2903_n3924.t9 gnd 0.094832f
C465 a_n2903_n3924.t4 gnd 0.094832f
C466 a_n2903_n3924.n5 gnd 0.774508f
C467 a_n2903_n3924.n6 gnd 0.314114f
C468 a_n2903_n3924.t34 gnd 0.094832f
C469 a_n2903_n3924.t33 gnd 0.094832f
C470 a_n2903_n3924.n7 gnd 0.774508f
C471 a_n2903_n3924.n8 gnd 0.314114f
C472 a_n2903_n3924.t10 gnd 0.985605f
C473 a_n2903_n3924.n9 gnd 0.850542f
C474 a_n2903_n3924.t35 gnd 1.22634f
C475 a_n2903_n3924.t5 gnd 1.22459f
C476 a_n2903_n3924.n10 gnd 1.34231f
C477 a_n2903_n3924.t36 gnd 1.22459f
C478 a_n2903_n3924.t11 gnd 1.22459f
C479 a_n2903_n3924.n11 gnd 0.8625f
C480 a_n2903_n3924.t38 gnd 1.22459f
C481 a_n2903_n3924.n12 gnd 0.8625f
C482 a_n2903_n3924.t12 gnd 1.22459f
C483 a_n2903_n3924.n13 gnd 0.8625f
C484 a_n2903_n3924.t8 gnd 1.22459f
C485 a_n2903_n3924.n14 gnd 0.614303f
C486 a_n2903_n3924.n15 gnd 0.466167f
C487 a_n2903_n3924.n16 gnd 0.885261f
C488 a_n2903_n3924.t26 gnd 0.985601f
C489 a_n2903_n3924.n17 gnd 0.54064f
C490 a_n2903_n3924.t18 gnd 0.094832f
C491 a_n2903_n3924.t21 gnd 0.094832f
C492 a_n2903_n3924.n18 gnd 0.774507f
C493 a_n2903_n3924.n19 gnd 0.314115f
C494 a_n2903_n3924.t15 gnd 0.094832f
C495 a_n2903_n3924.t19 gnd 0.094832f
C496 a_n2903_n3924.n20 gnd 0.774507f
C497 a_n2903_n3924.n21 gnd 0.314115f
C498 a_n2903_n3924.t25 gnd 0.094832f
C499 a_n2903_n3924.t20 gnd 0.094832f
C500 a_n2903_n3924.n22 gnd 0.774507f
C501 a_n2903_n3924.n23 gnd 0.314115f
C502 a_n2903_n3924.t22 gnd 0.985601f
C503 a_n2903_n3924.n24 gnd 0.334509f
C504 a_n2903_n3924.t29 gnd 0.985601f
C505 a_n2903_n3924.n25 gnd 0.334509f
C506 a_n2903_n3924.t6 gnd 0.094832f
C507 a_n2903_n3924.t31 gnd 0.094832f
C508 a_n2903_n3924.n26 gnd 0.774507f
C509 a_n2903_n3924.n27 gnd 0.314115f
C510 a_n2903_n3924.t1 gnd 0.094832f
C511 a_n2903_n3924.t3 gnd 0.094832f
C512 a_n2903_n3924.n28 gnd 0.774507f
C513 a_n2903_n3924.n29 gnd 0.314115f
C514 a_n2903_n3924.t30 gnd 0.094832f
C515 a_n2903_n3924.t2 gnd 0.094832f
C516 a_n2903_n3924.n30 gnd 0.774507f
C517 a_n2903_n3924.n31 gnd 0.314115f
C518 a_n2903_n3924.t32 gnd 0.985601f
C519 a_n2903_n3924.n32 gnd 0.54064f
C520 a_n2903_n3924.n33 gnd 0.885261f
C521 a_n2903_n3924.t17 gnd 0.985601f
C522 a_n2903_n3924.n34 gnd 0.850545f
C523 a_n2903_n3924.t27 gnd 0.094832f
C524 a_n2903_n3924.t24 gnd 0.094832f
C525 a_n2903_n3924.n35 gnd 0.774508f
C526 a_n2903_n3924.n36 gnd 0.314114f
C527 a_n2903_n3924.t13 gnd 0.094832f
C528 a_n2903_n3924.t23 gnd 0.094832f
C529 a_n2903_n3924.n37 gnd 0.774508f
C530 a_n2903_n3924.n38 gnd 0.314114f
C531 a_n2903_n3924.n39 gnd 0.314113f
C532 a_n2903_n3924.n40 gnd 0.774509f
C533 a_n2903_n3924.t28 gnd 0.094832f
C534 plus.n0 gnd 0.021615f
C535 plus.t7 gnd 0.21837f
C536 plus.t15 gnd 0.21837f
C537 plus.t12 gnd 0.21837f
C538 plus.n1 gnd 0.100959f
C539 plus.n2 gnd 0.021615f
C540 plus.t18 gnd 0.21837f
C541 plus.n3 gnd 0.021615f
C542 plus.t14 gnd 0.21837f
C543 plus.t8 gnd 0.21837f
C544 plus.n4 gnd 0.100959f
C545 plus.t11 gnd 0.223111f
C546 plus.n5 gnd 0.094111f
C547 plus.t13 gnd 0.21837f
C548 plus.n6 gnd 0.099693f
C549 plus.n7 gnd 0.004905f
C550 plus.n8 gnd 0.068817f
C551 plus.n9 gnd 0.021615f
C552 plus.n10 gnd 0.021615f
C553 plus.n11 gnd 0.004905f
C554 plus.n12 gnd 0.099827f
C555 plus.n13 gnd 0.099827f
C556 plus.n14 gnd 0.004905f
C557 plus.n15 gnd 0.021615f
C558 plus.n16 gnd 0.021615f
C559 plus.n17 gnd 0.021615f
C560 plus.n18 gnd 0.004905f
C561 plus.n19 gnd 0.099693f
C562 plus.n20 gnd 0.098694f
C563 plus.n21 gnd 0.238743f
C564 plus.n22 gnd 0.021615f
C565 plus.t6 gnd 0.21837f
C566 plus.n23 gnd 0.100959f
C567 plus.n24 gnd 0.021615f
C568 plus.n25 gnd 0.004905f
C569 plus.t20 gnd 0.21837f
C570 plus.n26 gnd 0.068817f
C571 plus.t5 gnd 0.21837f
C572 plus.t19 gnd 0.223111f
C573 plus.n27 gnd 0.094111f
C574 plus.n28 gnd 0.099693f
C575 plus.n29 gnd 0.004905f
C576 plus.t17 gnd 0.21837f
C577 plus.n30 gnd 0.100959f
C578 plus.n31 gnd 0.021615f
C579 plus.n32 gnd 0.021615f
C580 plus.n33 gnd 0.021615f
C581 plus.n34 gnd 0.099827f
C582 plus.t10 gnd 0.21837f
C583 plus.n35 gnd 0.099827f
C584 plus.n36 gnd 0.004905f
C585 plus.n37 gnd 0.021615f
C586 plus.n38 gnd 0.021615f
C587 plus.n39 gnd 0.021615f
C588 plus.n40 gnd 0.004905f
C589 plus.t9 gnd 0.21837f
C590 plus.n41 gnd 0.099693f
C591 plus.t16 gnd 0.21837f
C592 plus.n42 gnd 0.098694f
C593 plus.n43 gnd 0.57307f
C594 plus.n44 gnd 0.886647f
C595 plus.t4 gnd 0.037313f
C596 plus.t0 gnd 0.006663f
C597 plus.t1 gnd 0.006663f
C598 plus.n45 gnd 0.02161f
C599 plus.n46 gnd 0.167758f
C600 plus.t3 gnd 0.006663f
C601 plus.t2 gnd 0.006663f
C602 plus.n47 gnd 0.02161f
C603 plus.n48 gnd 0.125923f
C604 plus.n49 gnd 2.50274f
C605 a_n7636_8799.t15 gnd 0.144643f
C606 a_n7636_8799.t7 gnd 0.144643f
C607 a_n7636_8799.t14 gnd 0.144643f
C608 a_n7636_8799.n0 gnd 1.14082f
C609 a_n7636_8799.t13 gnd 0.144643f
C610 a_n7636_8799.t16 gnd 0.144643f
C611 a_n7636_8799.n1 gnd 1.13894f
C612 a_n7636_8799.n2 gnd 1.02377f
C613 a_n7636_8799.t11 gnd 0.144643f
C614 a_n7636_8799.t8 gnd 0.144643f
C615 a_n7636_8799.n3 gnd 1.13894f
C616 a_n7636_8799.n4 gnd 1.85609f
C617 a_n7636_8799.t25 gnd 0.1125f
C618 a_n7636_8799.t22 gnd 0.1125f
C619 a_n7636_8799.n5 gnd 0.995675f
C620 a_n7636_8799.t26 gnd 0.1125f
C621 a_n7636_8799.t1 gnd 0.1125f
C622 a_n7636_8799.n6 gnd 0.994091f
C623 a_n7636_8799.n7 gnd 0.655186f
C624 a_n7636_8799.t21 gnd 0.1125f
C625 a_n7636_8799.t27 gnd 0.1125f
C626 a_n7636_8799.n8 gnd 0.995675f
C627 a_n7636_8799.t0 gnd 0.1125f
C628 a_n7636_8799.t24 gnd 0.1125f
C629 a_n7636_8799.n9 gnd 0.99409f
C630 a_n7636_8799.n10 gnd 0.655188f
C631 a_n7636_8799.t3 gnd 0.1125f
C632 a_n7636_8799.t23 gnd 0.1125f
C633 a_n7636_8799.n11 gnd 0.995675f
C634 a_n7636_8799.t20 gnd 0.1125f
C635 a_n7636_8799.t19 gnd 0.1125f
C636 a_n7636_8799.n12 gnd 0.99409f
C637 a_n7636_8799.n13 gnd 0.655188f
C638 a_n7636_8799.n14 gnd 1.79181f
C639 a_n7636_8799.t6 gnd 0.1125f
C640 a_n7636_8799.t2 gnd 0.1125f
C641 a_n7636_8799.n15 gnd 0.994091f
C642 a_n7636_8799.n16 gnd 2.39774f
C643 a_n7636_8799.t4 gnd 0.1125f
C644 a_n7636_8799.t5 gnd 0.1125f
C645 a_n7636_8799.n17 gnd 0.994091f
C646 a_n7636_8799.n18 gnd 0.296749f
C647 a_n7636_8799.n19 gnd 0.449457f
C648 a_n7636_8799.n20 gnd 0.052134f
C649 a_n7636_8799.t125 gnd 0.599757f
C650 a_n7636_8799.n21 gnd 0.267863f
C651 a_n7636_8799.n22 gnd 0.052134f
C652 a_n7636_8799.n23 gnd 0.01183f
C653 a_n7636_8799.t41 gnd 0.599757f
C654 a_n7636_8799.n24 gnd 0.052134f
C655 a_n7636_8799.t62 gnd 0.599757f
C656 a_n7636_8799.n25 gnd 0.26481f
C657 a_n7636_8799.t85 gnd 0.599757f
C658 a_n7636_8799.n26 gnd 0.052134f
C659 a_n7636_8799.t104 gnd 0.599757f
C660 a_n7636_8799.n27 gnd 0.265131f
C661 a_n7636_8799.n28 gnd 0.052134f
C662 a_n7636_8799.n29 gnd 0.01183f
C663 a_n7636_8799.t64 gnd 0.599757f
C664 a_n7636_8799.n30 gnd 0.052134f
C665 a_n7636_8799.t76 gnd 0.599757f
C666 a_n7636_8799.n31 gnd 0.267863f
C667 a_n7636_8799.n32 gnd 0.052134f
C668 a_n7636_8799.n33 gnd 0.01183f
C669 a_n7636_8799.t109 gnd 0.599757f
C670 a_n7636_8799.n34 gnd 0.164706f
C671 a_n7636_8799.t130 gnd 0.599757f
C672 a_n7636_8799.t129 gnd 0.611109f
C673 a_n7636_8799.n35 gnd 0.251423f
C674 a_n7636_8799.n36 gnd 0.264167f
C675 a_n7636_8799.n37 gnd 0.01183f
C676 a_n7636_8799.t80 gnd 0.599757f
C677 a_n7636_8799.n38 gnd 0.267863f
C678 a_n7636_8799.n39 gnd 0.052134f
C679 a_n7636_8799.n40 gnd 0.052134f
C680 a_n7636_8799.n41 gnd 0.052134f
C681 a_n7636_8799.n42 gnd 0.265774f
C682 a_n7636_8799.t126 gnd 0.599757f
C683 a_n7636_8799.n43 gnd 0.264488f
C684 a_n7636_8799.n44 gnd 0.01183f
C685 a_n7636_8799.n45 gnd 0.052134f
C686 a_n7636_8799.n46 gnd 0.052134f
C687 a_n7636_8799.n47 gnd 0.052134f
C688 a_n7636_8799.n48 gnd 0.01183f
C689 a_n7636_8799.t77 gnd 0.599757f
C690 a_n7636_8799.n49 gnd 0.265452f
C691 a_n7636_8799.t107 gnd 0.599757f
C692 a_n7636_8799.n50 gnd 0.26481f
C693 a_n7636_8799.n51 gnd 0.052134f
C694 a_n7636_8799.n52 gnd 0.052134f
C695 a_n7636_8799.n53 gnd 0.052134f
C696 a_n7636_8799.n54 gnd 0.267863f
C697 a_n7636_8799.n55 gnd 0.01183f
C698 a_n7636_8799.t65 gnd 0.599757f
C699 a_n7636_8799.n56 gnd 0.265131f
C700 a_n7636_8799.n57 gnd 0.052134f
C701 a_n7636_8799.n58 gnd 0.052134f
C702 a_n7636_8799.n59 gnd 0.052134f
C703 a_n7636_8799.n60 gnd 0.01183f
C704 a_n7636_8799.t29 gnd 0.599757f
C705 a_n7636_8799.n61 gnd 0.267863f
C706 a_n7636_8799.n62 gnd 0.01183f
C707 a_n7636_8799.n63 gnd 0.052134f
C708 a_n7636_8799.n64 gnd 0.052134f
C709 a_n7636_8799.n65 gnd 0.052134f
C710 a_n7636_8799.n66 gnd 0.265452f
C711 a_n7636_8799.n67 gnd 0.01183f
C712 a_n7636_8799.t128 gnd 0.599757f
C713 a_n7636_8799.n68 gnd 0.267863f
C714 a_n7636_8799.n69 gnd 0.052134f
C715 a_n7636_8799.n70 gnd 0.052134f
C716 a_n7636_8799.n71 gnd 0.052134f
C717 a_n7636_8799.n72 gnd 0.264488f
C718 a_n7636_8799.t59 gnd 0.599757f
C719 a_n7636_8799.n73 gnd 0.265774f
C720 a_n7636_8799.n74 gnd 0.01183f
C721 a_n7636_8799.n75 gnd 0.052134f
C722 a_n7636_8799.n76 gnd 0.052134f
C723 a_n7636_8799.n77 gnd 0.052134f
C724 a_n7636_8799.n78 gnd 0.01183f
C725 a_n7636_8799.t38 gnd 0.599757f
C726 a_n7636_8799.n79 gnd 0.264167f
C727 a_n7636_8799.t39 gnd 0.599757f
C728 a_n7636_8799.n80 gnd 0.262399f
C729 a_n7636_8799.n81 gnd 0.295587f
C730 a_n7636_8799.n82 gnd 0.052134f
C731 a_n7636_8799.t138 gnd 0.599757f
C732 a_n7636_8799.n83 gnd 0.267863f
C733 a_n7636_8799.n84 gnd 0.052134f
C734 a_n7636_8799.n85 gnd 0.01183f
C735 a_n7636_8799.t56 gnd 0.599757f
C736 a_n7636_8799.n86 gnd 0.052134f
C737 a_n7636_8799.t71 gnd 0.599757f
C738 a_n7636_8799.n87 gnd 0.26481f
C739 a_n7636_8799.t98 gnd 0.599757f
C740 a_n7636_8799.n88 gnd 0.052134f
C741 a_n7636_8799.t116 gnd 0.599757f
C742 a_n7636_8799.n89 gnd 0.265131f
C743 a_n7636_8799.n90 gnd 0.052134f
C744 a_n7636_8799.n91 gnd 0.01183f
C745 a_n7636_8799.t74 gnd 0.599757f
C746 a_n7636_8799.n92 gnd 0.052134f
C747 a_n7636_8799.t86 gnd 0.599757f
C748 a_n7636_8799.n93 gnd 0.267863f
C749 a_n7636_8799.n94 gnd 0.052134f
C750 a_n7636_8799.n95 gnd 0.01183f
C751 a_n7636_8799.t122 gnd 0.599757f
C752 a_n7636_8799.n96 gnd 0.164706f
C753 a_n7636_8799.t147 gnd 0.599757f
C754 a_n7636_8799.t143 gnd 0.611109f
C755 a_n7636_8799.n97 gnd 0.251423f
C756 a_n7636_8799.n98 gnd 0.264167f
C757 a_n7636_8799.n99 gnd 0.01183f
C758 a_n7636_8799.t90 gnd 0.599757f
C759 a_n7636_8799.n100 gnd 0.267863f
C760 a_n7636_8799.n101 gnd 0.052134f
C761 a_n7636_8799.n102 gnd 0.052134f
C762 a_n7636_8799.n103 gnd 0.052134f
C763 a_n7636_8799.n104 gnd 0.265774f
C764 a_n7636_8799.t140 gnd 0.599757f
C765 a_n7636_8799.n105 gnd 0.264488f
C766 a_n7636_8799.n106 gnd 0.01183f
C767 a_n7636_8799.n107 gnd 0.052134f
C768 a_n7636_8799.n108 gnd 0.052134f
C769 a_n7636_8799.n109 gnd 0.052134f
C770 a_n7636_8799.n110 gnd 0.01183f
C771 a_n7636_8799.t87 gnd 0.599757f
C772 a_n7636_8799.n111 gnd 0.265452f
C773 a_n7636_8799.t120 gnd 0.599757f
C774 a_n7636_8799.n112 gnd 0.26481f
C775 a_n7636_8799.n113 gnd 0.052134f
C776 a_n7636_8799.n114 gnd 0.052134f
C777 a_n7636_8799.n115 gnd 0.052134f
C778 a_n7636_8799.n116 gnd 0.267863f
C779 a_n7636_8799.n117 gnd 0.01183f
C780 a_n7636_8799.t75 gnd 0.599757f
C781 a_n7636_8799.n118 gnd 0.265131f
C782 a_n7636_8799.n119 gnd 0.052134f
C783 a_n7636_8799.n120 gnd 0.052134f
C784 a_n7636_8799.n121 gnd 0.052134f
C785 a_n7636_8799.n122 gnd 0.01183f
C786 a_n7636_8799.t40 gnd 0.599757f
C787 a_n7636_8799.n123 gnd 0.267863f
C788 a_n7636_8799.n124 gnd 0.01183f
C789 a_n7636_8799.n125 gnd 0.052134f
C790 a_n7636_8799.n126 gnd 0.052134f
C791 a_n7636_8799.n127 gnd 0.052134f
C792 a_n7636_8799.n128 gnd 0.265452f
C793 a_n7636_8799.n129 gnd 0.01183f
C794 a_n7636_8799.t144 gnd 0.599757f
C795 a_n7636_8799.n130 gnd 0.267863f
C796 a_n7636_8799.n131 gnd 0.052134f
C797 a_n7636_8799.n132 gnd 0.052134f
C798 a_n7636_8799.n133 gnd 0.052134f
C799 a_n7636_8799.n134 gnd 0.264488f
C800 a_n7636_8799.t70 gnd 0.599757f
C801 a_n7636_8799.n135 gnd 0.265774f
C802 a_n7636_8799.n136 gnd 0.01183f
C803 a_n7636_8799.n137 gnd 0.052134f
C804 a_n7636_8799.n138 gnd 0.052134f
C805 a_n7636_8799.n139 gnd 0.052134f
C806 a_n7636_8799.n140 gnd 0.01183f
C807 a_n7636_8799.t50 gnd 0.599757f
C808 a_n7636_8799.n141 gnd 0.264167f
C809 a_n7636_8799.t52 gnd 0.599757f
C810 a_n7636_8799.n142 gnd 0.262399f
C811 a_n7636_8799.n143 gnd 0.129945f
C812 a_n7636_8799.n144 gnd 0.901652f
C813 a_n7636_8799.n145 gnd 0.052134f
C814 a_n7636_8799.t93 gnd 0.599757f
C815 a_n7636_8799.n146 gnd 0.267863f
C816 a_n7636_8799.n147 gnd 0.052134f
C817 a_n7636_8799.n148 gnd 0.01183f
C818 a_n7636_8799.t117 gnd 0.599757f
C819 a_n7636_8799.n149 gnd 0.052134f
C820 a_n7636_8799.t35 gnd 0.599757f
C821 a_n7636_8799.n150 gnd 0.26481f
C822 a_n7636_8799.t100 gnd 0.599757f
C823 a_n7636_8799.n151 gnd 0.052134f
C824 a_n7636_8799.t139 gnd 0.599757f
C825 a_n7636_8799.n152 gnd 0.265131f
C826 a_n7636_8799.n153 gnd 0.052134f
C827 a_n7636_8799.n154 gnd 0.01183f
C828 a_n7636_8799.t134 gnd 0.599757f
C829 a_n7636_8799.n155 gnd 0.052134f
C830 a_n7636_8799.t47 gnd 0.599757f
C831 a_n7636_8799.n156 gnd 0.267863f
C832 a_n7636_8799.n157 gnd 0.052134f
C833 a_n7636_8799.n158 gnd 0.01183f
C834 a_n7636_8799.t72 gnd 0.599757f
C835 a_n7636_8799.n159 gnd 0.164706f
C836 a_n7636_8799.t83 gnd 0.599757f
C837 a_n7636_8799.t105 gnd 0.611109f
C838 a_n7636_8799.n160 gnd 0.251423f
C839 a_n7636_8799.n161 gnd 0.264167f
C840 a_n7636_8799.n162 gnd 0.01183f
C841 a_n7636_8799.t121 gnd 0.599757f
C842 a_n7636_8799.n163 gnd 0.267863f
C843 a_n7636_8799.n164 gnd 0.052134f
C844 a_n7636_8799.n165 gnd 0.052134f
C845 a_n7636_8799.n166 gnd 0.052134f
C846 a_n7636_8799.n167 gnd 0.265774f
C847 a_n7636_8799.t131 gnd 0.599757f
C848 a_n7636_8799.n168 gnd 0.264488f
C849 a_n7636_8799.n169 gnd 0.01183f
C850 a_n7636_8799.n170 gnd 0.052134f
C851 a_n7636_8799.n171 gnd 0.052134f
C852 a_n7636_8799.n172 gnd 0.052134f
C853 a_n7636_8799.n173 gnd 0.01183f
C854 a_n7636_8799.t30 gnd 0.599757f
C855 a_n7636_8799.n174 gnd 0.265452f
C856 a_n7636_8799.t91 gnd 0.599757f
C857 a_n7636_8799.n175 gnd 0.26481f
C858 a_n7636_8799.n176 gnd 0.052134f
C859 a_n7636_8799.n177 gnd 0.052134f
C860 a_n7636_8799.n178 gnd 0.052134f
C861 a_n7636_8799.n179 gnd 0.267863f
C862 a_n7636_8799.n180 gnd 0.01183f
C863 a_n7636_8799.t108 gnd 0.599757f
C864 a_n7636_8799.n181 gnd 0.265131f
C865 a_n7636_8799.n182 gnd 0.052134f
C866 a_n7636_8799.n183 gnd 0.052134f
C867 a_n7636_8799.n184 gnd 0.052134f
C868 a_n7636_8799.n185 gnd 0.01183f
C869 a_n7636_8799.t84 gnd 0.599757f
C870 a_n7636_8799.n186 gnd 0.267863f
C871 a_n7636_8799.n187 gnd 0.01183f
C872 a_n7636_8799.n188 gnd 0.052134f
C873 a_n7636_8799.n189 gnd 0.052134f
C874 a_n7636_8799.n190 gnd 0.052134f
C875 a_n7636_8799.n191 gnd 0.265452f
C876 a_n7636_8799.n192 gnd 0.01183f
C877 a_n7636_8799.t54 gnd 0.599757f
C878 a_n7636_8799.n193 gnd 0.267863f
C879 a_n7636_8799.n194 gnd 0.052134f
C880 a_n7636_8799.n195 gnd 0.052134f
C881 a_n7636_8799.n196 gnd 0.052134f
C882 a_n7636_8799.n197 gnd 0.264488f
C883 a_n7636_8799.t63 gnd 0.599757f
C884 a_n7636_8799.n198 gnd 0.265774f
C885 a_n7636_8799.n199 gnd 0.01183f
C886 a_n7636_8799.n200 gnd 0.052134f
C887 a_n7636_8799.n201 gnd 0.052134f
C888 a_n7636_8799.n202 gnd 0.052134f
C889 a_n7636_8799.n203 gnd 0.01183f
C890 a_n7636_8799.t43 gnd 0.599757f
C891 a_n7636_8799.n204 gnd 0.264167f
C892 a_n7636_8799.t145 gnd 0.599757f
C893 a_n7636_8799.n205 gnd 0.262399f
C894 a_n7636_8799.n206 gnd 0.129945f
C895 a_n7636_8799.n207 gnd 1.40196f
C896 a_n7636_8799.n208 gnd 0.052134f
C897 a_n7636_8799.t79 gnd 0.599757f
C898 a_n7636_8799.t78 gnd 0.599757f
C899 a_n7636_8799.t51 gnd 0.599757f
C900 a_n7636_8799.n209 gnd 0.267863f
C901 a_n7636_8799.n210 gnd 0.052134f
C902 a_n7636_8799.t127 gnd 0.599757f
C903 a_n7636_8799.t82 gnd 0.599757f
C904 a_n7636_8799.n211 gnd 0.052134f
C905 a_n7636_8799.t58 gnd 0.599757f
C906 a_n7636_8799.n212 gnd 0.267863f
C907 a_n7636_8799.n213 gnd 0.052134f
C908 a_n7636_8799.t133 gnd 0.599757f
C909 a_n7636_8799.t99 gnd 0.599757f
C910 a_n7636_8799.n214 gnd 0.052134f
C911 a_n7636_8799.t97 gnd 0.599757f
C912 a_n7636_8799.n215 gnd 0.267863f
C913 a_n7636_8799.n216 gnd 0.052134f
C914 a_n7636_8799.t32 gnd 0.599757f
C915 a_n7636_8799.t103 gnd 0.599757f
C916 a_n7636_8799.n217 gnd 0.052134f
C917 a_n7636_8799.t102 gnd 0.599757f
C918 a_n7636_8799.n218 gnd 0.267863f
C919 a_n7636_8799.n219 gnd 0.052134f
C920 a_n7636_8799.t34 gnd 0.599757f
C921 a_n7636_8799.t33 gnd 0.599757f
C922 a_n7636_8799.n220 gnd 0.052134f
C923 a_n7636_8799.t119 gnd 0.599757f
C924 a_n7636_8799.n221 gnd 0.267863f
C925 a_n7636_8799.n222 gnd 0.052134f
C926 a_n7636_8799.t53 gnd 0.599757f
C927 a_n7636_8799.t36 gnd 0.599757f
C928 a_n7636_8799.n223 gnd 0.052134f
C929 a_n7636_8799.t123 gnd 0.599757f
C930 a_n7636_8799.n224 gnd 0.267863f
C931 a_n7636_8799.t57 gnd 0.611109f
C932 a_n7636_8799.n225 gnd 0.251423f
C933 a_n7636_8799.t81 gnd 0.599757f
C934 a_n7636_8799.n226 gnd 0.264167f
C935 a_n7636_8799.n227 gnd 0.01183f
C936 a_n7636_8799.n228 gnd 0.164706f
C937 a_n7636_8799.n229 gnd 0.052134f
C938 a_n7636_8799.n230 gnd 0.052134f
C939 a_n7636_8799.n231 gnd 0.01183f
C940 a_n7636_8799.n232 gnd 0.265774f
C941 a_n7636_8799.n233 gnd 0.264488f
C942 a_n7636_8799.n234 gnd 0.01183f
C943 a_n7636_8799.n235 gnd 0.052134f
C944 a_n7636_8799.n236 gnd 0.052134f
C945 a_n7636_8799.n237 gnd 0.052134f
C946 a_n7636_8799.n238 gnd 0.01183f
C947 a_n7636_8799.n239 gnd 0.265452f
C948 a_n7636_8799.n240 gnd 0.26481f
C949 a_n7636_8799.n241 gnd 0.01183f
C950 a_n7636_8799.n242 gnd 0.052134f
C951 a_n7636_8799.n243 gnd 0.052134f
C952 a_n7636_8799.n244 gnd 0.052134f
C953 a_n7636_8799.n245 gnd 0.01183f
C954 a_n7636_8799.n246 gnd 0.265131f
C955 a_n7636_8799.n247 gnd 0.265131f
C956 a_n7636_8799.n248 gnd 0.01183f
C957 a_n7636_8799.n249 gnd 0.052134f
C958 a_n7636_8799.n250 gnd 0.052134f
C959 a_n7636_8799.n251 gnd 0.052134f
C960 a_n7636_8799.n252 gnd 0.01183f
C961 a_n7636_8799.n253 gnd 0.26481f
C962 a_n7636_8799.n254 gnd 0.265452f
C963 a_n7636_8799.n255 gnd 0.01183f
C964 a_n7636_8799.n256 gnd 0.052134f
C965 a_n7636_8799.n257 gnd 0.052134f
C966 a_n7636_8799.n258 gnd 0.052134f
C967 a_n7636_8799.n259 gnd 0.01183f
C968 a_n7636_8799.n260 gnd 0.264488f
C969 a_n7636_8799.n261 gnd 0.265774f
C970 a_n7636_8799.n262 gnd 0.01183f
C971 a_n7636_8799.n263 gnd 0.052134f
C972 a_n7636_8799.n264 gnd 0.052134f
C973 a_n7636_8799.n265 gnd 0.052134f
C974 a_n7636_8799.n266 gnd 0.01183f
C975 a_n7636_8799.n267 gnd 0.264167f
C976 a_n7636_8799.n268 gnd 0.262399f
C977 a_n7636_8799.n269 gnd 0.295587f
C978 a_n7636_8799.n270 gnd 0.052134f
C979 a_n7636_8799.t89 gnd 0.599757f
C980 a_n7636_8799.t88 gnd 0.599757f
C981 a_n7636_8799.t66 gnd 0.599757f
C982 a_n7636_8799.n271 gnd 0.267863f
C983 a_n7636_8799.n272 gnd 0.052134f
C984 a_n7636_8799.t142 gnd 0.599757f
C985 a_n7636_8799.t96 gnd 0.599757f
C986 a_n7636_8799.n273 gnd 0.052134f
C987 a_n7636_8799.t69 gnd 0.599757f
C988 a_n7636_8799.n274 gnd 0.267863f
C989 a_n7636_8799.n275 gnd 0.052134f
C990 a_n7636_8799.t28 gnd 0.599757f
C991 a_n7636_8799.t112 gnd 0.599757f
C992 a_n7636_8799.n276 gnd 0.052134f
C993 a_n7636_8799.t111 gnd 0.599757f
C994 a_n7636_8799.n277 gnd 0.267863f
C995 a_n7636_8799.n278 gnd 0.052134f
C996 a_n7636_8799.t42 gnd 0.599757f
C997 a_n7636_8799.t115 gnd 0.599757f
C998 a_n7636_8799.n279 gnd 0.052134f
C999 a_n7636_8799.t114 gnd 0.599757f
C1000 a_n7636_8799.n280 gnd 0.267863f
C1001 a_n7636_8799.n281 gnd 0.052134f
C1002 a_n7636_8799.t46 gnd 0.599757f
C1003 a_n7636_8799.t45 gnd 0.599757f
C1004 a_n7636_8799.n282 gnd 0.052134f
C1005 a_n7636_8799.t136 gnd 0.599757f
C1006 a_n7636_8799.n283 gnd 0.267863f
C1007 a_n7636_8799.n284 gnd 0.052134f
C1008 a_n7636_8799.t67 gnd 0.599757f
C1009 a_n7636_8799.t48 gnd 0.599757f
C1010 a_n7636_8799.n285 gnd 0.052134f
C1011 a_n7636_8799.t137 gnd 0.599757f
C1012 a_n7636_8799.n286 gnd 0.267863f
C1013 a_n7636_8799.t68 gnd 0.611109f
C1014 a_n7636_8799.n287 gnd 0.251423f
C1015 a_n7636_8799.t95 gnd 0.599757f
C1016 a_n7636_8799.n288 gnd 0.264167f
C1017 a_n7636_8799.n289 gnd 0.01183f
C1018 a_n7636_8799.n290 gnd 0.164706f
C1019 a_n7636_8799.n291 gnd 0.052134f
C1020 a_n7636_8799.n292 gnd 0.052134f
C1021 a_n7636_8799.n293 gnd 0.01183f
C1022 a_n7636_8799.n294 gnd 0.265774f
C1023 a_n7636_8799.n295 gnd 0.264488f
C1024 a_n7636_8799.n296 gnd 0.01183f
C1025 a_n7636_8799.n297 gnd 0.052134f
C1026 a_n7636_8799.n298 gnd 0.052134f
C1027 a_n7636_8799.n299 gnd 0.052134f
C1028 a_n7636_8799.n300 gnd 0.01183f
C1029 a_n7636_8799.n301 gnd 0.265452f
C1030 a_n7636_8799.n302 gnd 0.26481f
C1031 a_n7636_8799.n303 gnd 0.01183f
C1032 a_n7636_8799.n304 gnd 0.052134f
C1033 a_n7636_8799.n305 gnd 0.052134f
C1034 a_n7636_8799.n306 gnd 0.052134f
C1035 a_n7636_8799.n307 gnd 0.01183f
C1036 a_n7636_8799.n308 gnd 0.265131f
C1037 a_n7636_8799.n309 gnd 0.265131f
C1038 a_n7636_8799.n310 gnd 0.01183f
C1039 a_n7636_8799.n311 gnd 0.052134f
C1040 a_n7636_8799.n312 gnd 0.052134f
C1041 a_n7636_8799.n313 gnd 0.052134f
C1042 a_n7636_8799.n314 gnd 0.01183f
C1043 a_n7636_8799.n315 gnd 0.26481f
C1044 a_n7636_8799.n316 gnd 0.265452f
C1045 a_n7636_8799.n317 gnd 0.01183f
C1046 a_n7636_8799.n318 gnd 0.052134f
C1047 a_n7636_8799.n319 gnd 0.052134f
C1048 a_n7636_8799.n320 gnd 0.052134f
C1049 a_n7636_8799.n321 gnd 0.01183f
C1050 a_n7636_8799.n322 gnd 0.264488f
C1051 a_n7636_8799.n323 gnd 0.265774f
C1052 a_n7636_8799.n324 gnd 0.01183f
C1053 a_n7636_8799.n325 gnd 0.052134f
C1054 a_n7636_8799.n326 gnd 0.052134f
C1055 a_n7636_8799.n327 gnd 0.052134f
C1056 a_n7636_8799.n328 gnd 0.01183f
C1057 a_n7636_8799.n329 gnd 0.264167f
C1058 a_n7636_8799.n330 gnd 0.262399f
C1059 a_n7636_8799.n331 gnd 0.129945f
C1060 a_n7636_8799.n332 gnd 0.901652f
C1061 a_n7636_8799.n333 gnd 0.052134f
C1062 a_n7636_8799.t146 gnd 0.599757f
C1063 a_n7636_8799.t44 gnd 0.599757f
C1064 a_n7636_8799.t94 gnd 0.599757f
C1065 a_n7636_8799.n334 gnd 0.267863f
C1066 a_n7636_8799.n335 gnd 0.052134f
C1067 a_n7636_8799.t31 gnd 0.599757f
C1068 a_n7636_8799.t118 gnd 0.599757f
C1069 a_n7636_8799.n336 gnd 0.052134f
C1070 a_n7636_8799.t55 gnd 0.599757f
C1071 a_n7636_8799.n337 gnd 0.267863f
C1072 a_n7636_8799.n338 gnd 0.052134f
C1073 a_n7636_8799.t101 gnd 0.599757f
C1074 a_n7636_8799.t37 gnd 0.599757f
C1075 a_n7636_8799.n339 gnd 0.052134f
C1076 a_n7636_8799.t61 gnd 0.599757f
C1077 a_n7636_8799.n340 gnd 0.267863f
C1078 a_n7636_8799.n341 gnd 0.052134f
C1079 a_n7636_8799.t141 gnd 0.599757f
C1080 a_n7636_8799.t110 gnd 0.599757f
C1081 a_n7636_8799.n342 gnd 0.052134f
C1082 a_n7636_8799.t135 gnd 0.599757f
C1083 a_n7636_8799.n343 gnd 0.267863f
C1084 a_n7636_8799.n344 gnd 0.052134f
C1085 a_n7636_8799.t92 gnd 0.599757f
C1086 a_n7636_8799.t113 gnd 0.599757f
C1087 a_n7636_8799.n345 gnd 0.052134f
C1088 a_n7636_8799.t49 gnd 0.599757f
C1089 a_n7636_8799.n346 gnd 0.267863f
C1090 a_n7636_8799.n347 gnd 0.052134f
C1091 a_n7636_8799.t132 gnd 0.599757f
C1092 a_n7636_8799.t73 gnd 0.599757f
C1093 a_n7636_8799.n348 gnd 0.052134f
C1094 a_n7636_8799.t124 gnd 0.599757f
C1095 a_n7636_8799.n349 gnd 0.267863f
C1096 a_n7636_8799.t106 gnd 0.611109f
C1097 a_n7636_8799.n350 gnd 0.251423f
C1098 a_n7636_8799.t60 gnd 0.599757f
C1099 a_n7636_8799.n351 gnd 0.264167f
C1100 a_n7636_8799.n352 gnd 0.01183f
C1101 a_n7636_8799.n353 gnd 0.164706f
C1102 a_n7636_8799.n354 gnd 0.052134f
C1103 a_n7636_8799.n355 gnd 0.052134f
C1104 a_n7636_8799.n356 gnd 0.01183f
C1105 a_n7636_8799.n357 gnd 0.265774f
C1106 a_n7636_8799.n358 gnd 0.264488f
C1107 a_n7636_8799.n359 gnd 0.01183f
C1108 a_n7636_8799.n360 gnd 0.052134f
C1109 a_n7636_8799.n361 gnd 0.052134f
C1110 a_n7636_8799.n362 gnd 0.052134f
C1111 a_n7636_8799.n363 gnd 0.01183f
C1112 a_n7636_8799.n364 gnd 0.265452f
C1113 a_n7636_8799.n365 gnd 0.26481f
C1114 a_n7636_8799.n366 gnd 0.01183f
C1115 a_n7636_8799.n367 gnd 0.052134f
C1116 a_n7636_8799.n368 gnd 0.052134f
C1117 a_n7636_8799.n369 gnd 0.052134f
C1118 a_n7636_8799.n370 gnd 0.01183f
C1119 a_n7636_8799.n371 gnd 0.265131f
C1120 a_n7636_8799.n372 gnd 0.265131f
C1121 a_n7636_8799.n373 gnd 0.01183f
C1122 a_n7636_8799.n374 gnd 0.052134f
C1123 a_n7636_8799.n375 gnd 0.052134f
C1124 a_n7636_8799.n376 gnd 0.052134f
C1125 a_n7636_8799.n377 gnd 0.01183f
C1126 a_n7636_8799.n378 gnd 0.26481f
C1127 a_n7636_8799.n379 gnd 0.265452f
C1128 a_n7636_8799.n380 gnd 0.01183f
C1129 a_n7636_8799.n381 gnd 0.052134f
C1130 a_n7636_8799.n382 gnd 0.052134f
C1131 a_n7636_8799.n383 gnd 0.052134f
C1132 a_n7636_8799.n384 gnd 0.01183f
C1133 a_n7636_8799.n385 gnd 0.264488f
C1134 a_n7636_8799.n386 gnd 0.265774f
C1135 a_n7636_8799.n387 gnd 0.01183f
C1136 a_n7636_8799.n388 gnd 0.052134f
C1137 a_n7636_8799.n389 gnd 0.052134f
C1138 a_n7636_8799.n390 gnd 0.052134f
C1139 a_n7636_8799.n391 gnd 0.01183f
C1140 a_n7636_8799.n392 gnd 0.264167f
C1141 a_n7636_8799.n393 gnd 0.262399f
C1142 a_n7636_8799.n394 gnd 0.129945f
C1143 a_n7636_8799.n395 gnd 1.17929f
C1144 a_n7636_8799.n396 gnd 12.302401f
C1145 a_n7636_8799.n397 gnd 4.38935f
C1146 a_n7636_8799.n398 gnd 5.71736f
C1147 a_n7636_8799.t10 gnd 0.144643f
C1148 a_n7636_8799.t9 gnd 0.144643f
C1149 a_n7636_8799.n399 gnd 1.13894f
C1150 a_n7636_8799.n400 gnd 2.91857f
C1151 a_n7636_8799.t12 gnd 0.144643f
C1152 a_n7636_8799.t17 gnd 0.144643f
C1153 a_n7636_8799.n401 gnd 1.14082f
C1154 a_n7636_8799.n402 gnd 1.02377f
C1155 a_n7636_8799.n403 gnd 1.13894f
C1156 a_n7636_8799.t18 gnd 0.144643f
C1157 a_n1808_13878.t4 gnd 0.185195f
C1158 a_n1808_13878.t0 gnd 0.185195f
C1159 a_n1808_13878.t2 gnd 0.185195f
C1160 a_n1808_13878.n0 gnd 1.4598f
C1161 a_n1808_13878.t6 gnd 0.185195f
C1162 a_n1808_13878.t1 gnd 0.185195f
C1163 a_n1808_13878.n1 gnd 1.45825f
C1164 a_n1808_13878.n2 gnd 2.03762f
C1165 a_n1808_13878.t5 gnd 0.185195f
C1166 a_n1808_13878.t9 gnd 0.185195f
C1167 a_n1808_13878.n3 gnd 1.46067f
C1168 a_n1808_13878.t10 gnd 0.185195f
C1169 a_n1808_13878.t3 gnd 0.185195f
C1170 a_n1808_13878.n4 gnd 1.45825f
C1171 a_n1808_13878.n5 gnd 1.31079f
C1172 a_n1808_13878.t7 gnd 0.185195f
C1173 a_n1808_13878.t8 gnd 0.185195f
C1174 a_n1808_13878.n6 gnd 1.45825f
C1175 a_n1808_13878.n7 gnd 1.80025f
C1176 a_n1808_13878.t13 gnd 1.73408f
C1177 a_n1808_13878.t16 gnd 0.185195f
C1178 a_n1808_13878.t17 gnd 0.185195f
C1179 a_n1808_13878.n8 gnd 1.30452f
C1180 a_n1808_13878.n9 gnd 1.4576f
C1181 a_n1808_13878.t12 gnd 1.73062f
C1182 a_n1808_13878.n10 gnd 0.733487f
C1183 a_n1808_13878.t15 gnd 1.73062f
C1184 a_n1808_13878.n11 gnd 0.733487f
C1185 a_n1808_13878.t18 gnd 0.185195f
C1186 a_n1808_13878.t19 gnd 0.185195f
C1187 a_n1808_13878.n12 gnd 1.30452f
C1188 a_n1808_13878.n13 gnd 0.74059f
C1189 a_n1808_13878.t14 gnd 1.73062f
C1190 a_n1808_13878.n14 gnd 1.7272f
C1191 a_n1808_13878.n15 gnd 2.51438f
C1192 a_n1808_13878.n16 gnd 3.69301f
C1193 a_n1808_13878.n17 gnd 1.45826f
C1194 a_n1808_13878.t11 gnd 0.185195f
C1195 a_n1986_8322.t0 gnd 0.125549p
C1196 a_n1986_8322.t11 gnd 0.093526f
C1197 a_n1986_8322.t3 gnd 0.875728f
C1198 a_n1986_8322.t5 gnd 0.093526f
C1199 a_n1986_8322.t8 gnd 0.093526f
C1200 a_n1986_8322.n0 gnd 0.658798f
C1201 a_n1986_8322.n1 gnd 0.736111f
C1202 a_n1986_8322.t7 gnd 0.093526f
C1203 a_n1986_8322.t1 gnd 0.093526f
C1204 a_n1986_8322.n2 gnd 0.658798f
C1205 a_n1986_8322.n3 gnd 0.374008f
C1206 a_n1986_8322.t19 gnd 0.873987f
C1207 a_n1986_8322.n4 gnd 0.766467f
C1208 a_n1986_8322.n5 gnd 3.77945f
C1209 a_n1986_8322.t6 gnd 0.875731f
C1210 a_n1986_8322.t2 gnd 0.093526f
C1211 a_n1986_8322.t20 gnd 0.093526f
C1212 a_n1986_8322.n6 gnd 0.658798f
C1213 a_n1986_8322.n7 gnd 0.736109f
C1214 a_n1986_8322.t4 gnd 0.093526f
C1215 a_n1986_8322.t9 gnd 0.093526f
C1216 a_n1986_8322.n8 gnd 0.658798f
C1217 a_n1986_8322.n9 gnd 0.374008f
C1218 a_n1986_8322.t18 gnd 0.873987f
C1219 a_n1986_8322.n10 gnd 1.39886f
C1220 a_n1986_8322.n11 gnd 1.5906f
C1221 a_n1986_8322.t14 gnd 0.873987f
C1222 a_n1986_8322.n12 gnd 0.872256f
C1223 a_n1986_8322.t12 gnd 0.875731f
C1224 a_n1986_8322.t16 gnd 0.093526f
C1225 a_n1986_8322.t15 gnd 0.093526f
C1226 a_n1986_8322.n13 gnd 0.658798f
C1227 a_n1986_8322.n14 gnd 0.736109f
C1228 a_n1986_8322.t10 gnd 0.873987f
C1229 a_n1986_8322.n15 gnd 0.37042f
C1230 a_n1986_8322.t13 gnd 0.873987f
C1231 a_n1986_8322.n16 gnd 0.37042f
C1232 a_n1986_8322.n17 gnd 0.374006f
C1233 a_n1986_8322.n18 gnd 0.658799f
C1234 a_n1986_8322.t17 gnd 0.093526f
C1235 vdd.t154 gnd 0.040782f
C1236 vdd.t138 gnd 0.040782f
C1237 vdd.n0 gnd 0.321655f
C1238 vdd.t166 gnd 0.040782f
C1239 vdd.t150 gnd 0.040782f
C1240 vdd.n1 gnd 0.321124f
C1241 vdd.n2 gnd 0.296137f
C1242 vdd.t135 gnd 0.040782f
C1243 vdd.t160 gnd 0.040782f
C1244 vdd.n3 gnd 0.321124f
C1245 vdd.n4 gnd 0.149768f
C1246 vdd.t158 gnd 0.040782f
C1247 vdd.t143 gnd 0.040782f
C1248 vdd.n5 gnd 0.321124f
C1249 vdd.n6 gnd 0.140529f
C1250 vdd.t164 gnd 0.040782f
C1251 vdd.t133 gnd 0.040782f
C1252 vdd.n7 gnd 0.321655f
C1253 vdd.t141 gnd 0.040782f
C1254 vdd.t156 gnd 0.040782f
C1255 vdd.n8 gnd 0.321124f
C1256 vdd.n9 gnd 0.296137f
C1257 vdd.t148 gnd 0.040782f
C1258 vdd.t125 gnd 0.040782f
C1259 vdd.n10 gnd 0.321124f
C1260 vdd.n11 gnd 0.149768f
C1261 vdd.t130 gnd 0.040782f
C1262 vdd.t146 gnd 0.040782f
C1263 vdd.n12 gnd 0.321124f
C1264 vdd.n13 gnd 0.140529f
C1265 vdd.n14 gnd 0.099352f
C1266 vdd.t27 gnd 0.022657f
C1267 vdd.t15 gnd 0.022657f
C1268 vdd.n15 gnd 0.208545f
C1269 vdd.t22 gnd 0.022657f
C1270 vdd.t23 gnd 0.022657f
C1271 vdd.n16 gnd 0.207935f
C1272 vdd.n17 gnd 0.361872f
C1273 vdd.t26 gnd 0.022657f
C1274 vdd.t25 gnd 0.022657f
C1275 vdd.n18 gnd 0.207935f
C1276 vdd.n19 gnd 0.149711f
C1277 vdd.t17 gnd 0.022657f
C1278 vdd.t18 gnd 0.022657f
C1279 vdd.n20 gnd 0.208545f
C1280 vdd.t19 gnd 0.022657f
C1281 vdd.t16 gnd 0.022657f
C1282 vdd.n21 gnd 0.207935f
C1283 vdd.n22 gnd 0.361872f
C1284 vdd.t12 gnd 0.022657f
C1285 vdd.t20 gnd 0.022657f
C1286 vdd.n23 gnd 0.207935f
C1287 vdd.n24 gnd 0.149711f
C1288 vdd.t24 gnd 0.022657f
C1289 vdd.t21 gnd 0.022657f
C1290 vdd.n25 gnd 0.207935f
C1291 vdd.t13 gnd 0.022657f
C1292 vdd.t14 gnd 0.022657f
C1293 vdd.n26 gnd 0.207935f
C1294 vdd.n27 gnd 23.0465f
C1295 vdd.n28 gnd 8.9102f
C1296 vdd.n29 gnd 0.006179f
C1297 vdd.n30 gnd 0.005734f
C1298 vdd.n31 gnd 0.003172f
C1299 vdd.n32 gnd 0.007283f
C1300 vdd.n33 gnd 0.003081f
C1301 vdd.n34 gnd 0.003263f
C1302 vdd.n35 gnd 0.005734f
C1303 vdd.n36 gnd 0.003081f
C1304 vdd.n37 gnd 0.007283f
C1305 vdd.n38 gnd 0.003263f
C1306 vdd.n39 gnd 0.005734f
C1307 vdd.n40 gnd 0.003081f
C1308 vdd.n41 gnd 0.005462f
C1309 vdd.n42 gnd 0.005479f
C1310 vdd.t251 gnd 0.015647f
C1311 vdd.n43 gnd 0.034815f
C1312 vdd.n44 gnd 0.181183f
C1313 vdd.n45 gnd 0.003081f
C1314 vdd.n46 gnd 0.003263f
C1315 vdd.n47 gnd 0.007283f
C1316 vdd.n48 gnd 0.007283f
C1317 vdd.n49 gnd 0.003263f
C1318 vdd.n50 gnd 0.003081f
C1319 vdd.n51 gnd 0.005734f
C1320 vdd.n52 gnd 0.005734f
C1321 vdd.n53 gnd 0.003081f
C1322 vdd.n54 gnd 0.003263f
C1323 vdd.n55 gnd 0.007283f
C1324 vdd.n56 gnd 0.007283f
C1325 vdd.n57 gnd 0.003263f
C1326 vdd.n58 gnd 0.003081f
C1327 vdd.n59 gnd 0.005734f
C1328 vdd.n60 gnd 0.005734f
C1329 vdd.n61 gnd 0.003081f
C1330 vdd.n62 gnd 0.003263f
C1331 vdd.n63 gnd 0.007283f
C1332 vdd.n64 gnd 0.007283f
C1333 vdd.n65 gnd 0.017219f
C1334 vdd.n66 gnd 0.003172f
C1335 vdd.n67 gnd 0.003081f
C1336 vdd.n68 gnd 0.014821f
C1337 vdd.n69 gnd 0.010347f
C1338 vdd.t286 gnd 0.036251f
C1339 vdd.t272 gnd 0.036251f
C1340 vdd.n70 gnd 0.24914f
C1341 vdd.n71 gnd 0.195911f
C1342 vdd.t250 gnd 0.036251f
C1343 vdd.t264 gnd 0.036251f
C1344 vdd.n72 gnd 0.24914f
C1345 vdd.n73 gnd 0.158099f
C1346 vdd.t117 gnd 0.036251f
C1347 vdd.t71 gnd 0.036251f
C1348 vdd.n74 gnd 0.24914f
C1349 vdd.n75 gnd 0.158099f
C1350 vdd.t291 gnd 0.036251f
C1351 vdd.t168 gnd 0.036251f
C1352 vdd.n76 gnd 0.24914f
C1353 vdd.n77 gnd 0.158099f
C1354 vdd.t255 gnd 0.036251f
C1355 vdd.t66 gnd 0.036251f
C1356 vdd.n78 gnd 0.24914f
C1357 vdd.n79 gnd 0.158099f
C1358 vdd.t50 gnd 0.036251f
C1359 vdd.t274 gnd 0.036251f
C1360 vdd.n80 gnd 0.24914f
C1361 vdd.n81 gnd 0.158099f
C1362 vdd.t268 gnd 0.036251f
C1363 vdd.t293 gnd 0.036251f
C1364 vdd.n82 gnd 0.24914f
C1365 vdd.n83 gnd 0.158099f
C1366 vdd.t37 gnd 0.036251f
C1367 vdd.t81 gnd 0.036251f
C1368 vdd.n84 gnd 0.24914f
C1369 vdd.n85 gnd 0.158099f
C1370 vdd.t61 gnd 0.036251f
C1371 vdd.t167 gnd 0.036251f
C1372 vdd.n86 gnd 0.24914f
C1373 vdd.n87 gnd 0.158099f
C1374 vdd.n88 gnd 0.006179f
C1375 vdd.n89 gnd 0.005734f
C1376 vdd.n90 gnd 0.003172f
C1377 vdd.n91 gnd 0.007283f
C1378 vdd.n92 gnd 0.003081f
C1379 vdd.n93 gnd 0.003263f
C1380 vdd.n94 gnd 0.005734f
C1381 vdd.n95 gnd 0.003081f
C1382 vdd.n96 gnd 0.007283f
C1383 vdd.n97 gnd 0.003263f
C1384 vdd.n98 gnd 0.005734f
C1385 vdd.n99 gnd 0.003081f
C1386 vdd.n100 gnd 0.005462f
C1387 vdd.n101 gnd 0.005479f
C1388 vdd.t269 gnd 0.015647f
C1389 vdd.n102 gnd 0.034815f
C1390 vdd.n103 gnd 0.181183f
C1391 vdd.n104 gnd 0.003081f
C1392 vdd.n105 gnd 0.003263f
C1393 vdd.n106 gnd 0.007283f
C1394 vdd.n107 gnd 0.007283f
C1395 vdd.n108 gnd 0.003263f
C1396 vdd.n109 gnd 0.003081f
C1397 vdd.n110 gnd 0.005734f
C1398 vdd.n111 gnd 0.005734f
C1399 vdd.n112 gnd 0.003081f
C1400 vdd.n113 gnd 0.003263f
C1401 vdd.n114 gnd 0.007283f
C1402 vdd.n115 gnd 0.007283f
C1403 vdd.n116 gnd 0.003263f
C1404 vdd.n117 gnd 0.003081f
C1405 vdd.n118 gnd 0.005734f
C1406 vdd.n119 gnd 0.005734f
C1407 vdd.n120 gnd 0.003081f
C1408 vdd.n121 gnd 0.003263f
C1409 vdd.n122 gnd 0.007283f
C1410 vdd.n123 gnd 0.007283f
C1411 vdd.n124 gnd 0.017219f
C1412 vdd.n125 gnd 0.003172f
C1413 vdd.n126 gnd 0.003081f
C1414 vdd.n127 gnd 0.014821f
C1415 vdd.n128 gnd 0.010023f
C1416 vdd.n129 gnd 0.117626f
C1417 vdd.n130 gnd 0.006179f
C1418 vdd.n131 gnd 0.005734f
C1419 vdd.n132 gnd 0.003172f
C1420 vdd.n133 gnd 0.007283f
C1421 vdd.n134 gnd 0.003081f
C1422 vdd.n135 gnd 0.003263f
C1423 vdd.n136 gnd 0.005734f
C1424 vdd.n137 gnd 0.003081f
C1425 vdd.n138 gnd 0.007283f
C1426 vdd.n139 gnd 0.003263f
C1427 vdd.n140 gnd 0.005734f
C1428 vdd.n141 gnd 0.003081f
C1429 vdd.n142 gnd 0.005462f
C1430 vdd.n143 gnd 0.005479f
C1431 vdd.t108 gnd 0.015647f
C1432 vdd.n144 gnd 0.034815f
C1433 vdd.n145 gnd 0.181183f
C1434 vdd.n146 gnd 0.003081f
C1435 vdd.n147 gnd 0.003263f
C1436 vdd.n148 gnd 0.007283f
C1437 vdd.n149 gnd 0.007283f
C1438 vdd.n150 gnd 0.003263f
C1439 vdd.n151 gnd 0.003081f
C1440 vdd.n152 gnd 0.005734f
C1441 vdd.n153 gnd 0.005734f
C1442 vdd.n154 gnd 0.003081f
C1443 vdd.n155 gnd 0.003263f
C1444 vdd.n156 gnd 0.007283f
C1445 vdd.n157 gnd 0.007283f
C1446 vdd.n158 gnd 0.003263f
C1447 vdd.n159 gnd 0.003081f
C1448 vdd.n160 gnd 0.005734f
C1449 vdd.n161 gnd 0.005734f
C1450 vdd.n162 gnd 0.003081f
C1451 vdd.n163 gnd 0.003263f
C1452 vdd.n164 gnd 0.007283f
C1453 vdd.n165 gnd 0.007283f
C1454 vdd.n166 gnd 0.017219f
C1455 vdd.n167 gnd 0.003172f
C1456 vdd.n168 gnd 0.003081f
C1457 vdd.n169 gnd 0.014821f
C1458 vdd.n170 gnd 0.010347f
C1459 vdd.t106 gnd 0.036251f
C1460 vdd.t278 gnd 0.036251f
C1461 vdd.n171 gnd 0.24914f
C1462 vdd.n172 gnd 0.195911f
C1463 vdd.t282 gnd 0.036251f
C1464 vdd.t103 gnd 0.036251f
C1465 vdd.n173 gnd 0.24914f
C1466 vdd.n174 gnd 0.158099f
C1467 vdd.t113 gnd 0.036251f
C1468 vdd.t9 gnd 0.036251f
C1469 vdd.n175 gnd 0.24914f
C1470 vdd.n176 gnd 0.158099f
C1471 vdd.t267 gnd 0.036251f
C1472 vdd.t68 gnd 0.036251f
C1473 vdd.n177 gnd 0.24914f
C1474 vdd.n178 gnd 0.158099f
C1475 vdd.t256 gnd 0.036251f
C1476 vdd.t40 gnd 0.036251f
C1477 vdd.n179 gnd 0.24914f
C1478 vdd.n180 gnd 0.158099f
C1479 vdd.t39 gnd 0.036251f
C1480 vdd.t51 gnd 0.036251f
C1481 vdd.n181 gnd 0.24914f
C1482 vdd.n182 gnd 0.158099f
C1483 vdd.t287 gnd 0.036251f
C1484 vdd.t284 gnd 0.036251f
C1485 vdd.n183 gnd 0.24914f
C1486 vdd.n184 gnd 0.158099f
C1487 vdd.t279 gnd 0.036251f
C1488 vdd.t292 gnd 0.036251f
C1489 vdd.n185 gnd 0.24914f
C1490 vdd.n186 gnd 0.158099f
C1491 vdd.t285 gnd 0.036251f
C1492 vdd.t273 gnd 0.036251f
C1493 vdd.n187 gnd 0.24914f
C1494 vdd.n188 gnd 0.158099f
C1495 vdd.n189 gnd 0.006179f
C1496 vdd.n190 gnd 0.005734f
C1497 vdd.n191 gnd 0.003172f
C1498 vdd.n192 gnd 0.007283f
C1499 vdd.n193 gnd 0.003081f
C1500 vdd.n194 gnd 0.003263f
C1501 vdd.n195 gnd 0.005734f
C1502 vdd.n196 gnd 0.003081f
C1503 vdd.n197 gnd 0.007283f
C1504 vdd.n198 gnd 0.003263f
C1505 vdd.n199 gnd 0.005734f
C1506 vdd.n200 gnd 0.003081f
C1507 vdd.n201 gnd 0.005462f
C1508 vdd.n202 gnd 0.005479f
C1509 vdd.t112 gnd 0.015647f
C1510 vdd.n203 gnd 0.034815f
C1511 vdd.n204 gnd 0.181183f
C1512 vdd.n205 gnd 0.003081f
C1513 vdd.n206 gnd 0.003263f
C1514 vdd.n207 gnd 0.007283f
C1515 vdd.n208 gnd 0.007283f
C1516 vdd.n209 gnd 0.003263f
C1517 vdd.n210 gnd 0.003081f
C1518 vdd.n211 gnd 0.005734f
C1519 vdd.n212 gnd 0.005734f
C1520 vdd.n213 gnd 0.003081f
C1521 vdd.n214 gnd 0.003263f
C1522 vdd.n215 gnd 0.007283f
C1523 vdd.n216 gnd 0.007283f
C1524 vdd.n217 gnd 0.003263f
C1525 vdd.n218 gnd 0.003081f
C1526 vdd.n219 gnd 0.005734f
C1527 vdd.n220 gnd 0.005734f
C1528 vdd.n221 gnd 0.003081f
C1529 vdd.n222 gnd 0.003263f
C1530 vdd.n223 gnd 0.007283f
C1531 vdd.n224 gnd 0.007283f
C1532 vdd.n225 gnd 0.017219f
C1533 vdd.n226 gnd 0.003172f
C1534 vdd.n227 gnd 0.003081f
C1535 vdd.n228 gnd 0.014821f
C1536 vdd.n229 gnd 0.010023f
C1537 vdd.n230 gnd 0.069976f
C1538 vdd.n231 gnd 0.252141f
C1539 vdd.n232 gnd 0.006179f
C1540 vdd.n233 gnd 0.005734f
C1541 vdd.n234 gnd 0.003172f
C1542 vdd.n235 gnd 0.007283f
C1543 vdd.n236 gnd 0.003081f
C1544 vdd.n237 gnd 0.003263f
C1545 vdd.n238 gnd 0.005734f
C1546 vdd.n239 gnd 0.003081f
C1547 vdd.n240 gnd 0.007283f
C1548 vdd.n241 gnd 0.003263f
C1549 vdd.n242 gnd 0.005734f
C1550 vdd.n243 gnd 0.003081f
C1551 vdd.n244 gnd 0.005462f
C1552 vdd.n245 gnd 0.005479f
C1553 vdd.t122 gnd 0.015647f
C1554 vdd.n246 gnd 0.034815f
C1555 vdd.n247 gnd 0.181183f
C1556 vdd.n248 gnd 0.003081f
C1557 vdd.n249 gnd 0.003263f
C1558 vdd.n250 gnd 0.007283f
C1559 vdd.n251 gnd 0.007283f
C1560 vdd.n252 gnd 0.003263f
C1561 vdd.n253 gnd 0.003081f
C1562 vdd.n254 gnd 0.005734f
C1563 vdd.n255 gnd 0.005734f
C1564 vdd.n256 gnd 0.003081f
C1565 vdd.n257 gnd 0.003263f
C1566 vdd.n258 gnd 0.007283f
C1567 vdd.n259 gnd 0.007283f
C1568 vdd.n260 gnd 0.003263f
C1569 vdd.n261 gnd 0.003081f
C1570 vdd.n262 gnd 0.005734f
C1571 vdd.n263 gnd 0.005734f
C1572 vdd.n264 gnd 0.003081f
C1573 vdd.n265 gnd 0.003263f
C1574 vdd.n266 gnd 0.007283f
C1575 vdd.n267 gnd 0.007283f
C1576 vdd.n268 gnd 0.017219f
C1577 vdd.n269 gnd 0.003172f
C1578 vdd.n270 gnd 0.003081f
C1579 vdd.n271 gnd 0.014821f
C1580 vdd.n272 gnd 0.010347f
C1581 vdd.t121 gnd 0.036251f
C1582 vdd.t295 gnd 0.036251f
C1583 vdd.n273 gnd 0.24914f
C1584 vdd.n274 gnd 0.195911f
C1585 vdd.t95 gnd 0.036251f
C1586 vdd.t288 gnd 0.036251f
C1587 vdd.n275 gnd 0.24914f
C1588 vdd.n276 gnd 0.158099f
C1589 vdd.t86 gnd 0.036251f
C1590 vdd.t38 gnd 0.036251f
C1591 vdd.n277 gnd 0.24914f
C1592 vdd.n278 gnd 0.158099f
C1593 vdd.t74 gnd 0.036251f
C1594 vdd.t104 gnd 0.036251f
C1595 vdd.n279 gnd 0.24914f
C1596 vdd.n280 gnd 0.158099f
C1597 vdd.t89 gnd 0.036251f
C1598 vdd.t3 gnd 0.036251f
C1599 vdd.n281 gnd 0.24914f
C1600 vdd.n282 gnd 0.158099f
C1601 vdd.t1 gnd 0.036251f
C1602 vdd.t33 gnd 0.036251f
C1603 vdd.n283 gnd 0.24914f
C1604 vdd.n284 gnd 0.158099f
C1605 vdd.t91 gnd 0.036251f
C1606 vdd.t266 gnd 0.036251f
C1607 vdd.n285 gnd 0.24914f
C1608 vdd.n286 gnd 0.158099f
C1609 vdd.t248 gnd 0.036251f
C1610 vdd.t290 gnd 0.036251f
C1611 vdd.n287 gnd 0.24914f
C1612 vdd.n288 gnd 0.158099f
C1613 vdd.t97 gnd 0.036251f
C1614 vdd.t31 gnd 0.036251f
C1615 vdd.n289 gnd 0.24914f
C1616 vdd.n290 gnd 0.158099f
C1617 vdd.n291 gnd 0.006179f
C1618 vdd.n292 gnd 0.005734f
C1619 vdd.n293 gnd 0.003172f
C1620 vdd.n294 gnd 0.007283f
C1621 vdd.n295 gnd 0.003081f
C1622 vdd.n296 gnd 0.003263f
C1623 vdd.n297 gnd 0.005734f
C1624 vdd.n298 gnd 0.003081f
C1625 vdd.n299 gnd 0.007283f
C1626 vdd.n300 gnd 0.003263f
C1627 vdd.n301 gnd 0.005734f
C1628 vdd.n302 gnd 0.003081f
C1629 vdd.n303 gnd 0.005462f
C1630 vdd.n304 gnd 0.005479f
C1631 vdd.t115 gnd 0.015647f
C1632 vdd.n305 gnd 0.034815f
C1633 vdd.n306 gnd 0.181183f
C1634 vdd.n307 gnd 0.003081f
C1635 vdd.n308 gnd 0.003263f
C1636 vdd.n309 gnd 0.007283f
C1637 vdd.n310 gnd 0.007283f
C1638 vdd.n311 gnd 0.003263f
C1639 vdd.n312 gnd 0.003081f
C1640 vdd.n313 gnd 0.005734f
C1641 vdd.n314 gnd 0.005734f
C1642 vdd.n315 gnd 0.003081f
C1643 vdd.n316 gnd 0.003263f
C1644 vdd.n317 gnd 0.007283f
C1645 vdd.n318 gnd 0.007283f
C1646 vdd.n319 gnd 0.003263f
C1647 vdd.n320 gnd 0.003081f
C1648 vdd.n321 gnd 0.005734f
C1649 vdd.n322 gnd 0.005734f
C1650 vdd.n323 gnd 0.003081f
C1651 vdd.n324 gnd 0.003263f
C1652 vdd.n325 gnd 0.007283f
C1653 vdd.n326 gnd 0.007283f
C1654 vdd.n327 gnd 0.017219f
C1655 vdd.n328 gnd 0.003172f
C1656 vdd.n329 gnd 0.003081f
C1657 vdd.n330 gnd 0.014821f
C1658 vdd.n331 gnd 0.010023f
C1659 vdd.n332 gnd 0.069976f
C1660 vdd.n333 gnd 0.288647f
C1661 vdd.n334 gnd 0.008654f
C1662 vdd.n335 gnd 0.01126f
C1663 vdd.n336 gnd 0.009063f
C1664 vdd.n337 gnd 0.009063f
C1665 vdd.n338 gnd 0.01126f
C1666 vdd.n339 gnd 0.01126f
C1667 vdd.n340 gnd 0.822741f
C1668 vdd.n341 gnd 0.01126f
C1669 vdd.n342 gnd 0.01126f
C1670 vdd.n343 gnd 0.01126f
C1671 vdd.n344 gnd 0.891782f
C1672 vdd.n345 gnd 0.01126f
C1673 vdd.n346 gnd 0.01126f
C1674 vdd.n347 gnd 0.01126f
C1675 vdd.n348 gnd 0.01126f
C1676 vdd.n349 gnd 0.009063f
C1677 vdd.n350 gnd 0.01126f
C1678 vdd.t32 gnd 0.575343f
C1679 vdd.n351 gnd 0.01126f
C1680 vdd.n352 gnd 0.01126f
C1681 vdd.n353 gnd 0.01126f
C1682 vdd.t265 gnd 0.575343f
C1683 vdd.n354 gnd 0.01126f
C1684 vdd.n355 gnd 0.01126f
C1685 vdd.n356 gnd 0.01126f
C1686 vdd.n357 gnd 0.01126f
C1687 vdd.n358 gnd 0.01126f
C1688 vdd.n359 gnd 0.009063f
C1689 vdd.n360 gnd 0.01126f
C1690 vdd.n361 gnd 0.650138f
C1691 vdd.n362 gnd 0.01126f
C1692 vdd.n363 gnd 0.01126f
C1693 vdd.n364 gnd 0.01126f
C1694 vdd.t80 gnd 0.575343f
C1695 vdd.n365 gnd 0.01126f
C1696 vdd.n366 gnd 0.01126f
C1697 vdd.n367 gnd 0.01126f
C1698 vdd.n368 gnd 0.01126f
C1699 vdd.n369 gnd 0.01126f
C1700 vdd.n370 gnd 0.009063f
C1701 vdd.n371 gnd 0.01126f
C1702 vdd.t60 gnd 0.575343f
C1703 vdd.n372 gnd 0.01126f
C1704 vdd.n373 gnd 0.01126f
C1705 vdd.n374 gnd 0.01126f
C1706 vdd.n375 gnd 0.673151f
C1707 vdd.n376 gnd 0.01126f
C1708 vdd.n377 gnd 0.01126f
C1709 vdd.n378 gnd 0.01126f
C1710 vdd.n379 gnd 0.01126f
C1711 vdd.n380 gnd 0.01126f
C1712 vdd.n381 gnd 0.009063f
C1713 vdd.n382 gnd 0.01126f
C1714 vdd.t111 gnd 0.575343f
C1715 vdd.n383 gnd 0.01126f
C1716 vdd.n384 gnd 0.01126f
C1717 vdd.n385 gnd 0.01126f
C1718 vdd.n386 gnd 0.581097f
C1719 vdd.n387 gnd 0.01126f
C1720 vdd.n388 gnd 0.01126f
C1721 vdd.n389 gnd 0.01126f
C1722 vdd.n390 gnd 0.01126f
C1723 vdd.n391 gnd 0.027238f
C1724 vdd.n392 gnd 0.027822f
C1725 vdd.t192 gnd 0.575343f
C1726 vdd.n393 gnd 0.027238f
C1727 vdd.n425 gnd 0.01126f
C1728 vdd.t194 gnd 0.138524f
C1729 vdd.t193 gnd 0.148044f
C1730 vdd.t191 gnd 0.18091f
C1731 vdd.n426 gnd 0.231901f
C1732 vdd.n427 gnd 0.195745f
C1733 vdd.n428 gnd 0.014863f
C1734 vdd.n429 gnd 0.01126f
C1735 vdd.n430 gnd 0.009063f
C1736 vdd.n431 gnd 0.01126f
C1737 vdd.n432 gnd 0.009063f
C1738 vdd.n433 gnd 0.01126f
C1739 vdd.n434 gnd 0.009063f
C1740 vdd.n435 gnd 0.01126f
C1741 vdd.n436 gnd 0.009063f
C1742 vdd.n437 gnd 0.01126f
C1743 vdd.n438 gnd 0.009063f
C1744 vdd.n439 gnd 0.01126f
C1745 vdd.t235 gnd 0.138524f
C1746 vdd.t234 gnd 0.148044f
C1747 vdd.t233 gnd 0.18091f
C1748 vdd.n440 gnd 0.231901f
C1749 vdd.n441 gnd 0.195745f
C1750 vdd.n442 gnd 0.009063f
C1751 vdd.n443 gnd 0.01126f
C1752 vdd.n444 gnd 0.009063f
C1753 vdd.n445 gnd 0.01126f
C1754 vdd.n446 gnd 0.009063f
C1755 vdd.n447 gnd 0.01126f
C1756 vdd.n448 gnd 0.009063f
C1757 vdd.n449 gnd 0.01126f
C1758 vdd.n450 gnd 0.009063f
C1759 vdd.n451 gnd 0.01126f
C1760 vdd.t241 gnd 0.138524f
C1761 vdd.t240 gnd 0.148044f
C1762 vdd.t239 gnd 0.18091f
C1763 vdd.n452 gnd 0.231901f
C1764 vdd.n453 gnd 0.195745f
C1765 vdd.n454 gnd 0.019394f
C1766 vdd.n455 gnd 0.01126f
C1767 vdd.n456 gnd 0.009063f
C1768 vdd.n457 gnd 0.01126f
C1769 vdd.n458 gnd 0.009063f
C1770 vdd.n459 gnd 0.01126f
C1771 vdd.n460 gnd 0.009063f
C1772 vdd.n461 gnd 0.01126f
C1773 vdd.n462 gnd 0.009063f
C1774 vdd.n463 gnd 0.01126f
C1775 vdd.n464 gnd 0.027822f
C1776 vdd.n465 gnd 0.007522f
C1777 vdd.n466 gnd 0.009063f
C1778 vdd.n467 gnd 0.01126f
C1779 vdd.n468 gnd 0.01126f
C1780 vdd.n469 gnd 0.009063f
C1781 vdd.n470 gnd 0.01126f
C1782 vdd.n471 gnd 0.01126f
C1783 vdd.n472 gnd 0.01126f
C1784 vdd.n473 gnd 0.01126f
C1785 vdd.n474 gnd 0.01126f
C1786 vdd.n475 gnd 0.009063f
C1787 vdd.n476 gnd 0.009063f
C1788 vdd.n477 gnd 0.01126f
C1789 vdd.n478 gnd 0.01126f
C1790 vdd.n479 gnd 0.009063f
C1791 vdd.n480 gnd 0.01126f
C1792 vdd.n481 gnd 0.01126f
C1793 vdd.n482 gnd 0.01126f
C1794 vdd.n483 gnd 0.01126f
C1795 vdd.n484 gnd 0.01126f
C1796 vdd.n485 gnd 0.009063f
C1797 vdd.n486 gnd 0.009063f
C1798 vdd.n487 gnd 0.01126f
C1799 vdd.n488 gnd 0.01126f
C1800 vdd.n489 gnd 0.009063f
C1801 vdd.n490 gnd 0.01126f
C1802 vdd.n491 gnd 0.01126f
C1803 vdd.n492 gnd 0.01126f
C1804 vdd.n493 gnd 0.01126f
C1805 vdd.n494 gnd 0.01126f
C1806 vdd.n495 gnd 0.009063f
C1807 vdd.n496 gnd 0.009063f
C1808 vdd.n497 gnd 0.01126f
C1809 vdd.n498 gnd 0.01126f
C1810 vdd.n499 gnd 0.009063f
C1811 vdd.n500 gnd 0.01126f
C1812 vdd.n501 gnd 0.01126f
C1813 vdd.n502 gnd 0.01126f
C1814 vdd.n503 gnd 0.01126f
C1815 vdd.n504 gnd 0.01126f
C1816 vdd.n505 gnd 0.009063f
C1817 vdd.n506 gnd 0.009063f
C1818 vdd.n507 gnd 0.01126f
C1819 vdd.n508 gnd 0.01126f
C1820 vdd.n509 gnd 0.007567f
C1821 vdd.n510 gnd 0.01126f
C1822 vdd.n511 gnd 0.01126f
C1823 vdd.n512 gnd 0.01126f
C1824 vdd.n513 gnd 0.01126f
C1825 vdd.n514 gnd 0.01126f
C1826 vdd.n515 gnd 0.007567f
C1827 vdd.n516 gnd 0.009063f
C1828 vdd.n517 gnd 0.01126f
C1829 vdd.n518 gnd 0.01126f
C1830 vdd.n519 gnd 0.009063f
C1831 vdd.n520 gnd 0.01126f
C1832 vdd.n521 gnd 0.01126f
C1833 vdd.n522 gnd 0.01126f
C1834 vdd.n523 gnd 0.01126f
C1835 vdd.n524 gnd 0.01126f
C1836 vdd.n525 gnd 0.009063f
C1837 vdd.n526 gnd 0.009063f
C1838 vdd.n527 gnd 0.01126f
C1839 vdd.n528 gnd 0.01126f
C1840 vdd.n529 gnd 0.009063f
C1841 vdd.n530 gnd 0.01126f
C1842 vdd.n531 gnd 0.01126f
C1843 vdd.n532 gnd 0.01126f
C1844 vdd.n533 gnd 0.01126f
C1845 vdd.n534 gnd 0.01126f
C1846 vdd.n535 gnd 0.009063f
C1847 vdd.n536 gnd 0.009063f
C1848 vdd.n537 gnd 0.01126f
C1849 vdd.n538 gnd 0.01126f
C1850 vdd.n539 gnd 0.009063f
C1851 vdd.n540 gnd 0.01126f
C1852 vdd.n541 gnd 0.01126f
C1853 vdd.n542 gnd 0.01126f
C1854 vdd.n543 gnd 0.01126f
C1855 vdd.n544 gnd 0.01126f
C1856 vdd.n545 gnd 0.009063f
C1857 vdd.n546 gnd 0.009063f
C1858 vdd.n547 gnd 0.01126f
C1859 vdd.n548 gnd 0.01126f
C1860 vdd.n549 gnd 0.009063f
C1861 vdd.n550 gnd 0.01126f
C1862 vdd.n551 gnd 0.01126f
C1863 vdd.n552 gnd 0.01126f
C1864 vdd.n553 gnd 0.01126f
C1865 vdd.n554 gnd 0.01126f
C1866 vdd.n555 gnd 0.009063f
C1867 vdd.n556 gnd 0.009063f
C1868 vdd.n557 gnd 0.01126f
C1869 vdd.n558 gnd 0.01126f
C1870 vdd.n559 gnd 0.009063f
C1871 vdd.n560 gnd 0.01126f
C1872 vdd.n561 gnd 0.01126f
C1873 vdd.n562 gnd 0.01126f
C1874 vdd.n563 gnd 0.01126f
C1875 vdd.n564 gnd 0.01126f
C1876 vdd.n565 gnd 0.006163f
C1877 vdd.n566 gnd 0.019394f
C1878 vdd.n567 gnd 0.01126f
C1879 vdd.n568 gnd 0.01126f
C1880 vdd.n569 gnd 0.008972f
C1881 vdd.n570 gnd 0.01126f
C1882 vdd.n571 gnd 0.01126f
C1883 vdd.n572 gnd 0.01126f
C1884 vdd.n573 gnd 0.01126f
C1885 vdd.n574 gnd 0.01126f
C1886 vdd.n575 gnd 0.009063f
C1887 vdd.n576 gnd 0.009063f
C1888 vdd.n577 gnd 0.01126f
C1889 vdd.n578 gnd 0.01126f
C1890 vdd.n579 gnd 0.009063f
C1891 vdd.n580 gnd 0.01126f
C1892 vdd.n581 gnd 0.01126f
C1893 vdd.n582 gnd 0.01126f
C1894 vdd.n583 gnd 0.01126f
C1895 vdd.n584 gnd 0.01126f
C1896 vdd.n585 gnd 0.009063f
C1897 vdd.n586 gnd 0.009063f
C1898 vdd.n587 gnd 0.01126f
C1899 vdd.n588 gnd 0.01126f
C1900 vdd.n589 gnd 0.009063f
C1901 vdd.n590 gnd 0.01126f
C1902 vdd.n591 gnd 0.01126f
C1903 vdd.n592 gnd 0.01126f
C1904 vdd.n593 gnd 0.01126f
C1905 vdd.n594 gnd 0.01126f
C1906 vdd.n595 gnd 0.009063f
C1907 vdd.n596 gnd 0.009063f
C1908 vdd.n597 gnd 0.01126f
C1909 vdd.n598 gnd 0.01126f
C1910 vdd.n599 gnd 0.009063f
C1911 vdd.n600 gnd 0.01126f
C1912 vdd.n601 gnd 0.01126f
C1913 vdd.n602 gnd 0.01126f
C1914 vdd.n603 gnd 0.01126f
C1915 vdd.n604 gnd 0.01126f
C1916 vdd.n605 gnd 0.009063f
C1917 vdd.n606 gnd 0.009063f
C1918 vdd.n607 gnd 0.01126f
C1919 vdd.n608 gnd 0.01126f
C1920 vdd.n609 gnd 0.009063f
C1921 vdd.n610 gnd 0.01126f
C1922 vdd.n611 gnd 0.01126f
C1923 vdd.n612 gnd 0.01126f
C1924 vdd.n613 gnd 0.01126f
C1925 vdd.n614 gnd 0.01126f
C1926 vdd.n615 gnd 0.009063f
C1927 vdd.n616 gnd 0.01126f
C1928 vdd.n617 gnd 0.009063f
C1929 vdd.n618 gnd 0.004758f
C1930 vdd.n619 gnd 0.01126f
C1931 vdd.n620 gnd 0.01126f
C1932 vdd.n621 gnd 0.009063f
C1933 vdd.n622 gnd 0.01126f
C1934 vdd.n623 gnd 0.009063f
C1935 vdd.n624 gnd 0.01126f
C1936 vdd.n625 gnd 0.009063f
C1937 vdd.n626 gnd 0.01126f
C1938 vdd.n627 gnd 0.009063f
C1939 vdd.n628 gnd 0.01126f
C1940 vdd.n629 gnd 0.009063f
C1941 vdd.n630 gnd 0.01126f
C1942 vdd.n631 gnd 0.009063f
C1943 vdd.n632 gnd 0.01126f
C1944 vdd.n633 gnd 0.627124f
C1945 vdd.t88 gnd 0.575343f
C1946 vdd.n634 gnd 0.01126f
C1947 vdd.n635 gnd 0.009063f
C1948 vdd.n636 gnd 0.01126f
C1949 vdd.n637 gnd 0.009063f
C1950 vdd.n638 gnd 0.01126f
C1951 vdd.t73 gnd 0.575343f
C1952 vdd.n639 gnd 0.01126f
C1953 vdd.n640 gnd 0.009063f
C1954 vdd.n641 gnd 0.01126f
C1955 vdd.n642 gnd 0.009063f
C1956 vdd.n643 gnd 0.01126f
C1957 vdd.t8 gnd 0.575343f
C1958 vdd.n644 gnd 0.719179f
C1959 vdd.n645 gnd 0.01126f
C1960 vdd.n646 gnd 0.009063f
C1961 vdd.n647 gnd 0.01126f
C1962 vdd.n648 gnd 0.009063f
C1963 vdd.n649 gnd 0.01126f
C1964 vdd.t85 gnd 0.575343f
C1965 vdd.n650 gnd 0.01126f
C1966 vdd.n651 gnd 0.009063f
C1967 vdd.n652 gnd 0.01126f
C1968 vdd.n653 gnd 0.009063f
C1969 vdd.n654 gnd 0.01126f
C1970 vdd.n655 gnd 0.799727f
C1971 vdd.n656 gnd 0.95507f
C1972 vdd.t102 gnd 0.575343f
C1973 vdd.n657 gnd 0.01126f
C1974 vdd.n658 gnd 0.009063f
C1975 vdd.n659 gnd 0.01126f
C1976 vdd.n660 gnd 0.009063f
C1977 vdd.n661 gnd 0.01126f
C1978 vdd.n662 gnd 0.60411f
C1979 vdd.n663 gnd 0.01126f
C1980 vdd.n664 gnd 0.009063f
C1981 vdd.n665 gnd 0.01126f
C1982 vdd.n666 gnd 0.009063f
C1983 vdd.n667 gnd 0.01126f
C1984 vdd.t105 gnd 0.575343f
C1985 vdd.t271 gnd 0.575343f
C1986 vdd.n668 gnd 0.01126f
C1987 vdd.n669 gnd 0.009063f
C1988 vdd.n670 gnd 0.01126f
C1989 vdd.n671 gnd 0.009063f
C1990 vdd.n672 gnd 0.01126f
C1991 vdd.t107 gnd 0.575343f
C1992 vdd.n673 gnd 0.01126f
C1993 vdd.n674 gnd 0.009063f
C1994 vdd.n675 gnd 0.01126f
C1995 vdd.n676 gnd 0.009063f
C1996 vdd.n677 gnd 0.01126f
C1997 vdd.n678 gnd 1.15069f
C1998 vdd.n679 gnd 0.937809f
C1999 vdd.n680 gnd 0.01126f
C2000 vdd.n681 gnd 0.009063f
C2001 vdd.n682 gnd 0.027238f
C2002 vdd.n683 gnd 0.007522f
C2003 vdd.n684 gnd 0.027238f
C2004 vdd.t170 gnd 0.575343f
C2005 vdd.n685 gnd 0.027238f
C2006 vdd.n686 gnd 0.007522f
C2007 vdd.n687 gnd 0.009683f
C2008 vdd.t237 gnd 0.138524f
C2009 vdd.t238 gnd 0.148044f
C2010 vdd.t236 gnd 0.18091f
C2011 vdd.n688 gnd 0.231901f
C2012 vdd.n689 gnd 0.194839f
C2013 vdd.n690 gnd 0.013957f
C2014 vdd.n691 gnd 0.01126f
C2015 vdd.n692 gnd 7.92823f
C2016 vdd.n723 gnd 1.58219f
C2017 vdd.n724 gnd 0.01126f
C2018 vdd.n725 gnd 0.01126f
C2019 vdd.n726 gnd 0.027822f
C2020 vdd.n727 gnd 0.009683f
C2021 vdd.n728 gnd 0.01126f
C2022 vdd.n729 gnd 0.009063f
C2023 vdd.n730 gnd 0.007206f
C2024 vdd.n731 gnd 0.018399f
C2025 vdd.n732 gnd 0.009063f
C2026 vdd.n733 gnd 0.01126f
C2027 vdd.n734 gnd 0.01126f
C2028 vdd.n735 gnd 0.01126f
C2029 vdd.n736 gnd 0.01126f
C2030 vdd.n737 gnd 0.01126f
C2031 vdd.n738 gnd 0.01126f
C2032 vdd.n739 gnd 0.01126f
C2033 vdd.n740 gnd 0.01126f
C2034 vdd.n741 gnd 0.01126f
C2035 vdd.n742 gnd 0.01126f
C2036 vdd.n743 gnd 0.01126f
C2037 vdd.n744 gnd 0.01126f
C2038 vdd.n745 gnd 0.01126f
C2039 vdd.n746 gnd 0.01126f
C2040 vdd.n747 gnd 0.007567f
C2041 vdd.n748 gnd 0.01126f
C2042 vdd.n749 gnd 0.01126f
C2043 vdd.n750 gnd 0.01126f
C2044 vdd.n751 gnd 0.01126f
C2045 vdd.n752 gnd 0.01126f
C2046 vdd.n753 gnd 0.01126f
C2047 vdd.n754 gnd 0.01126f
C2048 vdd.n755 gnd 0.01126f
C2049 vdd.n756 gnd 0.01126f
C2050 vdd.n757 gnd 0.01126f
C2051 vdd.n758 gnd 0.01126f
C2052 vdd.n759 gnd 0.01126f
C2053 vdd.n760 gnd 0.01126f
C2054 vdd.n761 gnd 0.01126f
C2055 vdd.n762 gnd 0.01126f
C2056 vdd.n763 gnd 0.01126f
C2057 vdd.n764 gnd 0.01126f
C2058 vdd.n765 gnd 0.01126f
C2059 vdd.n766 gnd 0.01126f
C2060 vdd.n767 gnd 0.008972f
C2061 vdd.t171 gnd 0.138524f
C2062 vdd.t172 gnd 0.148044f
C2063 vdd.t169 gnd 0.18091f
C2064 vdd.n768 gnd 0.231901f
C2065 vdd.n769 gnd 0.194839f
C2066 vdd.n770 gnd 0.01126f
C2067 vdd.n771 gnd 0.01126f
C2068 vdd.n772 gnd 0.01126f
C2069 vdd.n773 gnd 0.01126f
C2070 vdd.n774 gnd 0.01126f
C2071 vdd.n775 gnd 0.01126f
C2072 vdd.n776 gnd 0.01126f
C2073 vdd.n777 gnd 0.01126f
C2074 vdd.n778 gnd 0.01126f
C2075 vdd.n779 gnd 0.01126f
C2076 vdd.n780 gnd 0.01126f
C2077 vdd.n781 gnd 0.01126f
C2078 vdd.n782 gnd 0.01126f
C2079 vdd.n783 gnd 0.007206f
C2080 vdd.n785 gnd 0.007657f
C2081 vdd.n786 gnd 0.007657f
C2082 vdd.n787 gnd 0.007657f
C2083 vdd.n788 gnd 0.007657f
C2084 vdd.n789 gnd 0.007657f
C2085 vdd.n790 gnd 0.007657f
C2086 vdd.n792 gnd 0.007657f
C2087 vdd.n793 gnd 0.007657f
C2088 vdd.n795 gnd 0.007657f
C2089 vdd.n796 gnd 0.005574f
C2090 vdd.n798 gnd 0.007657f
C2091 vdd.t218 gnd 0.309402f
C2092 vdd.t217 gnd 0.316711f
C2093 vdd.t216 gnd 0.201989f
C2094 vdd.n799 gnd 0.109164f
C2095 vdd.n800 gnd 0.061921f
C2096 vdd.n801 gnd 0.010943f
C2097 vdd.n802 gnd 0.017895f
C2098 vdd.n804 gnd 0.007657f
C2099 vdd.n805 gnd 0.782467f
C2100 vdd.n806 gnd 0.016963f
C2101 vdd.n807 gnd 0.016963f
C2102 vdd.n808 gnd 0.007657f
C2103 vdd.n809 gnd 0.018168f
C2104 vdd.n810 gnd 0.007657f
C2105 vdd.n811 gnd 0.007657f
C2106 vdd.n812 gnd 0.007657f
C2107 vdd.n813 gnd 0.007657f
C2108 vdd.n814 gnd 0.007657f
C2109 vdd.n816 gnd 0.007657f
C2110 vdd.n817 gnd 0.007657f
C2111 vdd.n819 gnd 0.007657f
C2112 vdd.n820 gnd 0.007657f
C2113 vdd.n822 gnd 0.007657f
C2114 vdd.n823 gnd 0.007657f
C2115 vdd.n825 gnd 0.007657f
C2116 vdd.n826 gnd 0.007657f
C2117 vdd.n828 gnd 0.007657f
C2118 vdd.n829 gnd 0.007657f
C2119 vdd.n831 gnd 0.007657f
C2120 vdd.t211 gnd 0.309402f
C2121 vdd.t210 gnd 0.316711f
C2122 vdd.t208 gnd 0.201989f
C2123 vdd.n832 gnd 0.109164f
C2124 vdd.n833 gnd 0.061921f
C2125 vdd.n834 gnd 0.007657f
C2126 vdd.n836 gnd 0.007657f
C2127 vdd.n837 gnd 0.007657f
C2128 vdd.t209 gnd 0.391233f
C2129 vdd.n838 gnd 0.007657f
C2130 vdd.n839 gnd 0.007657f
C2131 vdd.n840 gnd 0.007657f
C2132 vdd.n841 gnd 0.007657f
C2133 vdd.n842 gnd 0.007657f
C2134 vdd.n843 gnd 0.782467f
C2135 vdd.n844 gnd 0.007657f
C2136 vdd.n845 gnd 0.007657f
C2137 vdd.n846 gnd 0.684658f
C2138 vdd.n847 gnd 0.007657f
C2139 vdd.n848 gnd 0.007657f
C2140 vdd.n849 gnd 0.006756f
C2141 vdd.n850 gnd 0.007657f
C2142 vdd.n851 gnd 0.690412f
C2143 vdd.n852 gnd 0.007657f
C2144 vdd.n853 gnd 0.007657f
C2145 vdd.n854 gnd 0.007657f
C2146 vdd.n855 gnd 0.007657f
C2147 vdd.n856 gnd 0.007657f
C2148 vdd.n857 gnd 0.782467f
C2149 vdd.n858 gnd 0.007657f
C2150 vdd.n859 gnd 0.007657f
C2151 vdd.t181 gnd 0.350959f
C2152 vdd.t126 gnd 0.092055f
C2153 vdd.n860 gnd 0.007657f
C2154 vdd.n861 gnd 0.007657f
C2155 vdd.n862 gnd 0.007657f
C2156 vdd.t136 gnd 0.391233f
C2157 vdd.n863 gnd 0.007657f
C2158 vdd.n864 gnd 0.007657f
C2159 vdd.n865 gnd 0.007657f
C2160 vdd.n866 gnd 0.007657f
C2161 vdd.n867 gnd 0.007657f
C2162 vdd.t151 gnd 0.391233f
C2163 vdd.n868 gnd 0.007657f
C2164 vdd.n869 gnd 0.007657f
C2165 vdd.n870 gnd 0.650138f
C2166 vdd.n871 gnd 0.007657f
C2167 vdd.n872 gnd 0.007657f
C2168 vdd.n873 gnd 0.007657f
C2169 vdd.n874 gnd 0.477535f
C2170 vdd.n875 gnd 0.007657f
C2171 vdd.n876 gnd 0.007657f
C2172 vdd.t132 gnd 0.391233f
C2173 vdd.n877 gnd 0.007657f
C2174 vdd.n878 gnd 0.007657f
C2175 vdd.n879 gnd 0.007657f
C2176 vdd.n880 gnd 0.650138f
C2177 vdd.n881 gnd 0.007657f
C2178 vdd.n882 gnd 0.007657f
C2179 vdd.t144 gnd 0.333699f
C2180 vdd.t163 gnd 0.304932f
C2181 vdd.n883 gnd 0.007657f
C2182 vdd.n884 gnd 0.007657f
C2183 vdd.n885 gnd 0.007657f
C2184 vdd.t155 gnd 0.391233f
C2185 vdd.n886 gnd 0.007657f
C2186 vdd.n887 gnd 0.007657f
C2187 vdd.t152 gnd 0.391233f
C2188 vdd.n888 gnd 0.007657f
C2189 vdd.n889 gnd 0.007657f
C2190 vdd.n890 gnd 0.007657f
C2191 vdd.t123 gnd 0.287672f
C2192 vdd.n891 gnd 0.007657f
C2193 vdd.n892 gnd 0.007657f
C2194 vdd.n893 gnd 0.667398f
C2195 vdd.n894 gnd 0.007657f
C2196 vdd.n895 gnd 0.007657f
C2197 vdd.n896 gnd 0.007657f
C2198 vdd.n897 gnd 0.782467f
C2199 vdd.n898 gnd 0.007657f
C2200 vdd.n899 gnd 0.007657f
C2201 vdd.t140 gnd 0.350959f
C2202 vdd.n900 gnd 0.494795f
C2203 vdd.n901 gnd 0.007657f
C2204 vdd.n902 gnd 0.007657f
C2205 vdd.n903 gnd 0.007657f
C2206 vdd.t124 gnd 0.391233f
C2207 vdd.n904 gnd 0.007657f
C2208 vdd.n905 gnd 0.007657f
C2209 vdd.n906 gnd 0.007657f
C2210 vdd.n907 gnd 0.007657f
C2211 vdd.n908 gnd 0.007657f
C2212 vdd.t147 gnd 0.782467f
C2213 vdd.n909 gnd 0.007657f
C2214 vdd.n910 gnd 0.007657f
C2215 vdd.t213 gnd 0.391233f
C2216 vdd.n911 gnd 0.007657f
C2217 vdd.n912 gnd 0.018168f
C2218 vdd.n913 gnd 0.018168f
C2219 vdd.t145 gnd 0.736439f
C2220 vdd.n914 gnd 0.016963f
C2221 vdd.n915 gnd 0.016963f
C2222 vdd.n916 gnd 0.018168f
C2223 vdd.n917 gnd 0.007657f
C2224 vdd.n918 gnd 0.007657f
C2225 vdd.t157 gnd 0.736439f
C2226 vdd.n936 gnd 0.018168f
C2227 vdd.n954 gnd 0.016963f
C2228 vdd.n955 gnd 0.007657f
C2229 vdd.n956 gnd 0.016963f
C2230 vdd.t232 gnd 0.309402f
C2231 vdd.t231 gnd 0.316711f
C2232 vdd.t230 gnd 0.201989f
C2233 vdd.n957 gnd 0.109164f
C2234 vdd.n958 gnd 0.061921f
C2235 vdd.n959 gnd 0.017895f
C2236 vdd.n960 gnd 0.007657f
C2237 vdd.t159 gnd 0.782467f
C2238 vdd.n961 gnd 0.016963f
C2239 vdd.n962 gnd 0.007657f
C2240 vdd.n963 gnd 0.018168f
C2241 vdd.n964 gnd 0.007657f
C2242 vdd.t207 gnd 0.309402f
C2243 vdd.t206 gnd 0.316711f
C2244 vdd.t204 gnd 0.201989f
C2245 vdd.n965 gnd 0.109164f
C2246 vdd.n966 gnd 0.061921f
C2247 vdd.n967 gnd 0.010943f
C2248 vdd.n968 gnd 0.007657f
C2249 vdd.n969 gnd 0.007657f
C2250 vdd.t205 gnd 0.391233f
C2251 vdd.n970 gnd 0.007657f
C2252 vdd.n971 gnd 0.007657f
C2253 vdd.n972 gnd 0.007657f
C2254 vdd.n973 gnd 0.007657f
C2255 vdd.n974 gnd 0.007657f
C2256 vdd.n975 gnd 0.007657f
C2257 vdd.n976 gnd 0.782467f
C2258 vdd.n977 gnd 0.007657f
C2259 vdd.n978 gnd 0.007657f
C2260 vdd.t134 gnd 0.391233f
C2261 vdd.n979 gnd 0.007657f
C2262 vdd.n980 gnd 0.007657f
C2263 vdd.n981 gnd 0.007657f
C2264 vdd.n982 gnd 0.007657f
C2265 vdd.n983 gnd 0.494795f
C2266 vdd.n984 gnd 0.007657f
C2267 vdd.n985 gnd 0.007657f
C2268 vdd.n986 gnd 0.007657f
C2269 vdd.n987 gnd 0.007657f
C2270 vdd.n988 gnd 0.007657f
C2271 vdd.n989 gnd 0.667398f
C2272 vdd.n990 gnd 0.007657f
C2273 vdd.n991 gnd 0.007657f
C2274 vdd.t149 gnd 0.350959f
C2275 vdd.t162 gnd 0.287672f
C2276 vdd.n992 gnd 0.007657f
C2277 vdd.n993 gnd 0.007657f
C2278 vdd.n994 gnd 0.007657f
C2279 vdd.t139 gnd 0.391233f
C2280 vdd.n995 gnd 0.007657f
C2281 vdd.n996 gnd 0.007657f
C2282 vdd.t165 gnd 0.391233f
C2283 vdd.n997 gnd 0.007657f
C2284 vdd.n998 gnd 0.007657f
C2285 vdd.n999 gnd 0.007657f
C2286 vdd.t137 gnd 0.304932f
C2287 vdd.n1000 gnd 0.007657f
C2288 vdd.n1001 gnd 0.007657f
C2289 vdd.n1002 gnd 0.650138f
C2290 vdd.n1003 gnd 0.007657f
C2291 vdd.n1004 gnd 0.007657f
C2292 vdd.n1005 gnd 0.007657f
C2293 vdd.t153 gnd 0.391233f
C2294 vdd.n1006 gnd 0.007657f
C2295 vdd.n1007 gnd 0.007657f
C2296 vdd.t128 gnd 0.333699f
C2297 vdd.n1008 gnd 0.477535f
C2298 vdd.n1009 gnd 0.007657f
C2299 vdd.n1010 gnd 0.007657f
C2300 vdd.n1011 gnd 0.007657f
C2301 vdd.n1012 gnd 0.650138f
C2302 vdd.n1013 gnd 0.007657f
C2303 vdd.n1014 gnd 0.007657f
C2304 vdd.t161 gnd 0.391233f
C2305 vdd.n1015 gnd 0.007657f
C2306 vdd.n1016 gnd 0.007657f
C2307 vdd.n1017 gnd 0.007657f
C2308 vdd.n1018 gnd 0.782467f
C2309 vdd.n1019 gnd 0.007657f
C2310 vdd.n1020 gnd 0.007657f
C2311 vdd.t131 gnd 0.391233f
C2312 vdd.n1021 gnd 0.007657f
C2313 vdd.n1022 gnd 0.007657f
C2314 vdd.n1023 gnd 0.007657f
C2315 vdd.t127 gnd 0.092055f
C2316 vdd.n1024 gnd 0.007657f
C2317 vdd.n1025 gnd 0.007657f
C2318 vdd.n1026 gnd 0.007657f
C2319 vdd.t225 gnd 0.316711f
C2320 vdd.t223 gnd 0.201989f
C2321 vdd.t226 gnd 0.316711f
C2322 vdd.n1027 gnd 0.178004f
C2323 vdd.n1028 gnd 0.007657f
C2324 vdd.n1029 gnd 0.007657f
C2325 vdd.n1030 gnd 0.782467f
C2326 vdd.n1031 gnd 0.007657f
C2327 vdd.n1032 gnd 0.007657f
C2328 vdd.t224 gnd 0.350959f
C2329 vdd.n1033 gnd 0.690412f
C2330 vdd.n1034 gnd 0.007657f
C2331 vdd.n1035 gnd 0.007657f
C2332 vdd.n1036 gnd 0.007657f
C2333 vdd.n1037 gnd 0.684658f
C2334 vdd.n1038 gnd 0.007657f
C2335 vdd.n1039 gnd 0.007657f
C2336 vdd.n1040 gnd 0.007657f
C2337 vdd.n1041 gnd 0.007657f
C2338 vdd.n1042 gnd 0.007657f
C2339 vdd.n1043 gnd 0.782467f
C2340 vdd.n1044 gnd 0.007657f
C2341 vdd.n1045 gnd 0.007657f
C2342 vdd.t220 gnd 0.391233f
C2343 vdd.n1046 gnd 0.007657f
C2344 vdd.n1047 gnd 0.018168f
C2345 vdd.n1048 gnd 0.018168f
C2346 vdd.n1049 gnd 7.92823f
C2347 vdd.n1050 gnd 0.016963f
C2348 vdd.n1051 gnd 0.016963f
C2349 vdd.n1052 gnd 0.018168f
C2350 vdd.n1053 gnd 0.007657f
C2351 vdd.n1054 gnd 0.007657f
C2352 vdd.n1055 gnd 0.007657f
C2353 vdd.n1056 gnd 0.007657f
C2354 vdd.n1057 gnd 0.007657f
C2355 vdd.n1058 gnd 0.007657f
C2356 vdd.n1059 gnd 0.007657f
C2357 vdd.n1060 gnd 0.007657f
C2358 vdd.n1062 gnd 0.007657f
C2359 vdd.n1063 gnd 0.007657f
C2360 vdd.n1064 gnd 0.007206f
C2361 vdd.n1067 gnd 0.027822f
C2362 vdd.n1068 gnd 0.009063f
C2363 vdd.n1069 gnd 0.01126f
C2364 vdd.n1071 gnd 0.01126f
C2365 vdd.n1072 gnd 0.007522f
C2366 vdd.t177 gnd 0.575343f
C2367 vdd.n1073 gnd 8.31946f
C2368 vdd.n1074 gnd 0.01126f
C2369 vdd.n1075 gnd 0.027822f
C2370 vdd.n1076 gnd 0.009063f
C2371 vdd.n1077 gnd 0.01126f
C2372 vdd.n1078 gnd 0.009063f
C2373 vdd.n1079 gnd 0.01126f
C2374 vdd.n1080 gnd 1.15069f
C2375 vdd.n1081 gnd 0.01126f
C2376 vdd.n1082 gnd 0.009063f
C2377 vdd.n1083 gnd 0.009063f
C2378 vdd.n1084 gnd 0.01126f
C2379 vdd.n1085 gnd 0.009063f
C2380 vdd.n1086 gnd 0.01126f
C2381 vdd.t43 gnd 0.575343f
C2382 vdd.n1087 gnd 0.01126f
C2383 vdd.n1088 gnd 0.009063f
C2384 vdd.n1089 gnd 0.01126f
C2385 vdd.n1090 gnd 0.009063f
C2386 vdd.n1091 gnd 0.01126f
C2387 vdd.t54 gnd 0.575343f
C2388 vdd.n1092 gnd 0.01126f
C2389 vdd.n1093 gnd 0.009063f
C2390 vdd.n1094 gnd 0.01126f
C2391 vdd.n1095 gnd 0.009063f
C2392 vdd.n1096 gnd 0.01126f
C2393 vdd.n1097 gnd 0.926302f
C2394 vdd.n1098 gnd 0.95507f
C2395 vdd.t45 gnd 0.575343f
C2396 vdd.n1099 gnd 0.01126f
C2397 vdd.n1100 gnd 0.009063f
C2398 vdd.n1101 gnd 0.01126f
C2399 vdd.n1102 gnd 0.009063f
C2400 vdd.n1103 gnd 0.01126f
C2401 vdd.n1104 gnd 0.730686f
C2402 vdd.n1105 gnd 0.01126f
C2403 vdd.n1106 gnd 0.009063f
C2404 vdd.n1107 gnd 0.01126f
C2405 vdd.n1108 gnd 0.009063f
C2406 vdd.n1109 gnd 0.01126f
C2407 vdd.t41 gnd 0.575343f
C2408 vdd.t64 gnd 0.575343f
C2409 vdd.n1110 gnd 0.01126f
C2410 vdd.n1111 gnd 0.009063f
C2411 vdd.n1112 gnd 0.01126f
C2412 vdd.n1113 gnd 0.009063f
C2413 vdd.n1114 gnd 0.01126f
C2414 vdd.t69 gnd 0.575343f
C2415 vdd.n1115 gnd 0.01126f
C2416 vdd.n1116 gnd 0.009063f
C2417 vdd.n1117 gnd 0.01126f
C2418 vdd.n1118 gnd 0.009063f
C2419 vdd.n1119 gnd 0.01126f
C2420 vdd.t34 gnd 0.575343f
C2421 vdd.n1120 gnd 0.811234f
C2422 vdd.n1121 gnd 0.01126f
C2423 vdd.n1122 gnd 0.009063f
C2424 vdd.n1123 gnd 0.01126f
C2425 vdd.n1124 gnd 0.009063f
C2426 vdd.n1125 gnd 0.01126f
C2427 vdd.n1126 gnd 0.903289f
C2428 vdd.n1127 gnd 0.01126f
C2429 vdd.n1128 gnd 0.009063f
C2430 vdd.n1129 gnd 0.01126f
C2431 vdd.n1130 gnd 0.009063f
C2432 vdd.n1131 gnd 0.01126f
C2433 vdd.n1132 gnd 0.707672f
C2434 vdd.t47 gnd 0.575343f
C2435 vdd.n1133 gnd 0.01126f
C2436 vdd.n1134 gnd 0.009063f
C2437 vdd.n1135 gnd 0.01126f
C2438 vdd.n1136 gnd 0.009063f
C2439 vdd.n1137 gnd 0.01126f
C2440 vdd.t4 gnd 0.575343f
C2441 vdd.n1138 gnd 0.01126f
C2442 vdd.n1139 gnd 0.009063f
C2443 vdd.n1140 gnd 0.01126f
C2444 vdd.n1141 gnd 0.009063f
C2445 vdd.n1142 gnd 0.01126f
C2446 vdd.t76 gnd 0.575343f
C2447 vdd.n1143 gnd 0.638631f
C2448 vdd.n1144 gnd 0.01126f
C2449 vdd.n1145 gnd 0.009063f
C2450 vdd.n1146 gnd 0.01126f
C2451 vdd.n1147 gnd 0.009063f
C2452 vdd.n1148 gnd 0.01126f
C2453 vdd.t119 gnd 0.575343f
C2454 vdd.n1149 gnd 0.01126f
C2455 vdd.n1150 gnd 0.009063f
C2456 vdd.n1151 gnd 0.01126f
C2457 vdd.n1152 gnd 0.009063f
C2458 vdd.n1153 gnd 0.01126f
C2459 vdd.n1154 gnd 0.880275f
C2460 vdd.n1155 gnd 0.95507f
C2461 vdd.t52 gnd 0.575343f
C2462 vdd.n1156 gnd 0.01126f
C2463 vdd.n1157 gnd 0.009063f
C2464 vdd.n1158 gnd 0.01126f
C2465 vdd.n1159 gnd 0.009063f
C2466 vdd.n1160 gnd 0.01126f
C2467 vdd.n1161 gnd 0.684658f
C2468 vdd.n1162 gnd 0.01126f
C2469 vdd.n1163 gnd 0.009063f
C2470 vdd.n1164 gnd 0.01126f
C2471 vdd.n1165 gnd 0.009063f
C2472 vdd.n1166 gnd 0.01126f
C2473 vdd.t28 gnd 0.575343f
C2474 vdd.t78 gnd 0.575343f
C2475 vdd.n1167 gnd 0.01126f
C2476 vdd.n1168 gnd 0.009063f
C2477 vdd.n1169 gnd 0.01126f
C2478 vdd.n1170 gnd 0.009063f
C2479 vdd.n1171 gnd 0.01126f
C2480 vdd.t252 gnd 0.575343f
C2481 vdd.n1172 gnd 0.01126f
C2482 vdd.n1173 gnd 0.009063f
C2483 vdd.n1174 gnd 0.01126f
C2484 vdd.n1175 gnd 0.009063f
C2485 vdd.n1176 gnd 0.01126f
C2486 vdd.t58 gnd 0.575343f
C2487 vdd.n1177 gnd 0.857261f
C2488 vdd.n1178 gnd 0.01126f
C2489 vdd.n1179 gnd 0.009063f
C2490 vdd.n1180 gnd 0.01126f
C2491 vdd.n1181 gnd 0.009063f
C2492 vdd.n1182 gnd 0.01126f
C2493 vdd.n1183 gnd 1.15069f
C2494 vdd.n1184 gnd 0.01126f
C2495 vdd.n1185 gnd 0.009063f
C2496 vdd.n1186 gnd 0.027238f
C2497 vdd.n1187 gnd 0.007522f
C2498 vdd.n1188 gnd 0.027238f
C2499 vdd.t185 gnd 0.575343f
C2500 vdd.n1189 gnd 0.027238f
C2501 vdd.n1190 gnd 0.007522f
C2502 vdd.n1191 gnd 0.01126f
C2503 vdd.n1192 gnd 0.009063f
C2504 vdd.n1193 gnd 0.01126f
C2505 vdd.n1224 gnd 0.027822f
C2506 vdd.n1225 gnd 1.69726f
C2507 vdd.n1226 gnd 0.01126f
C2508 vdd.n1227 gnd 0.009063f
C2509 vdd.n1228 gnd 0.01126f
C2510 vdd.n1229 gnd 0.01126f
C2511 vdd.n1230 gnd 0.01126f
C2512 vdd.n1231 gnd 0.01126f
C2513 vdd.n1232 gnd 0.01126f
C2514 vdd.n1233 gnd 0.009063f
C2515 vdd.n1234 gnd 0.01126f
C2516 vdd.n1235 gnd 0.01126f
C2517 vdd.n1236 gnd 0.01126f
C2518 vdd.n1237 gnd 0.01126f
C2519 vdd.n1238 gnd 0.01126f
C2520 vdd.n1239 gnd 0.009063f
C2521 vdd.n1240 gnd 0.01126f
C2522 vdd.n1241 gnd 0.01126f
C2523 vdd.n1242 gnd 0.01126f
C2524 vdd.n1243 gnd 0.01126f
C2525 vdd.n1244 gnd 0.01126f
C2526 vdd.n1245 gnd 0.009063f
C2527 vdd.n1246 gnd 0.01126f
C2528 vdd.n1247 gnd 0.01126f
C2529 vdd.n1248 gnd 0.01126f
C2530 vdd.n1249 gnd 0.01126f
C2531 vdd.n1250 gnd 0.01126f
C2532 vdd.t199 gnd 0.138524f
C2533 vdd.t200 gnd 0.148044f
C2534 vdd.t198 gnd 0.18091f
C2535 vdd.n1251 gnd 0.231901f
C2536 vdd.n1252 gnd 0.195745f
C2537 vdd.n1253 gnd 0.019394f
C2538 vdd.n1254 gnd 0.01126f
C2539 vdd.n1255 gnd 0.01126f
C2540 vdd.n1256 gnd 0.01126f
C2541 vdd.n1257 gnd 0.01126f
C2542 vdd.n1258 gnd 0.01126f
C2543 vdd.n1259 gnd 0.009063f
C2544 vdd.n1260 gnd 0.01126f
C2545 vdd.n1261 gnd 0.01126f
C2546 vdd.n1262 gnd 0.01126f
C2547 vdd.n1263 gnd 0.01126f
C2548 vdd.n1264 gnd 0.01126f
C2549 vdd.n1265 gnd 0.009063f
C2550 vdd.n1266 gnd 0.01126f
C2551 vdd.n1267 gnd 0.01126f
C2552 vdd.n1268 gnd 0.01126f
C2553 vdd.n1269 gnd 0.01126f
C2554 vdd.n1270 gnd 0.01126f
C2555 vdd.n1271 gnd 0.009063f
C2556 vdd.n1272 gnd 0.01126f
C2557 vdd.n1273 gnd 0.01126f
C2558 vdd.n1274 gnd 0.01126f
C2559 vdd.n1275 gnd 0.01126f
C2560 vdd.n1276 gnd 0.01126f
C2561 vdd.n1277 gnd 0.009063f
C2562 vdd.n1278 gnd 0.01126f
C2563 vdd.n1279 gnd 0.01126f
C2564 vdd.n1280 gnd 0.01126f
C2565 vdd.n1281 gnd 0.01126f
C2566 vdd.n1282 gnd 0.01126f
C2567 vdd.n1283 gnd 0.009063f
C2568 vdd.n1284 gnd 0.01126f
C2569 vdd.n1285 gnd 0.01126f
C2570 vdd.n1286 gnd 0.01126f
C2571 vdd.n1287 gnd 0.01126f
C2572 vdd.n1288 gnd 0.009063f
C2573 vdd.n1289 gnd 0.01126f
C2574 vdd.n1290 gnd 0.01126f
C2575 vdd.n1291 gnd 0.01126f
C2576 vdd.n1292 gnd 0.01126f
C2577 vdd.n1293 gnd 0.01126f
C2578 vdd.n1294 gnd 0.009063f
C2579 vdd.n1295 gnd 0.01126f
C2580 vdd.n1296 gnd 0.01126f
C2581 vdd.n1297 gnd 0.01126f
C2582 vdd.n1298 gnd 0.01126f
C2583 vdd.n1299 gnd 0.01126f
C2584 vdd.n1300 gnd 0.009063f
C2585 vdd.n1301 gnd 0.01126f
C2586 vdd.n1302 gnd 0.01126f
C2587 vdd.n1303 gnd 0.01126f
C2588 vdd.n1304 gnd 0.01126f
C2589 vdd.n1305 gnd 0.01126f
C2590 vdd.n1306 gnd 0.009063f
C2591 vdd.n1307 gnd 0.01126f
C2592 vdd.n1308 gnd 0.01126f
C2593 vdd.n1309 gnd 0.01126f
C2594 vdd.n1310 gnd 0.01126f
C2595 vdd.n1311 gnd 0.01126f
C2596 vdd.n1312 gnd 0.009063f
C2597 vdd.n1313 gnd 0.01126f
C2598 vdd.n1314 gnd 0.01126f
C2599 vdd.n1315 gnd 0.01126f
C2600 vdd.n1316 gnd 0.01126f
C2601 vdd.t196 gnd 0.138524f
C2602 vdd.t197 gnd 0.148044f
C2603 vdd.t195 gnd 0.18091f
C2604 vdd.n1317 gnd 0.231901f
C2605 vdd.n1318 gnd 0.195745f
C2606 vdd.n1319 gnd 0.014863f
C2607 vdd.n1320 gnd 0.004305f
C2608 vdd.n1321 gnd 0.027822f
C2609 vdd.n1322 gnd 0.01126f
C2610 vdd.n1323 gnd 0.004758f
C2611 vdd.n1324 gnd 0.009063f
C2612 vdd.n1325 gnd 0.009063f
C2613 vdd.n1326 gnd 0.01126f
C2614 vdd.n1327 gnd 0.01126f
C2615 vdd.n1328 gnd 0.01126f
C2616 vdd.n1329 gnd 0.009063f
C2617 vdd.n1330 gnd 0.009063f
C2618 vdd.n1331 gnd 0.009063f
C2619 vdd.n1332 gnd 0.01126f
C2620 vdd.n1333 gnd 0.01126f
C2621 vdd.n1334 gnd 0.01126f
C2622 vdd.n1335 gnd 0.009063f
C2623 vdd.n1336 gnd 0.009063f
C2624 vdd.n1337 gnd 0.009063f
C2625 vdd.n1338 gnd 0.01126f
C2626 vdd.n1339 gnd 0.01126f
C2627 vdd.n1340 gnd 0.01126f
C2628 vdd.n1341 gnd 0.009063f
C2629 vdd.n1342 gnd 0.009063f
C2630 vdd.n1343 gnd 0.009063f
C2631 vdd.n1344 gnd 0.01126f
C2632 vdd.n1345 gnd 0.01126f
C2633 vdd.n1346 gnd 0.01126f
C2634 vdd.n1347 gnd 0.009063f
C2635 vdd.n1348 gnd 0.009063f
C2636 vdd.n1349 gnd 0.009063f
C2637 vdd.n1350 gnd 0.01126f
C2638 vdd.n1351 gnd 0.01126f
C2639 vdd.n1352 gnd 0.01126f
C2640 vdd.n1353 gnd 0.008972f
C2641 vdd.n1354 gnd 0.01126f
C2642 vdd.t186 gnd 0.138524f
C2643 vdd.t187 gnd 0.148044f
C2644 vdd.t184 gnd 0.18091f
C2645 vdd.n1355 gnd 0.231901f
C2646 vdd.n1356 gnd 0.195745f
C2647 vdd.n1357 gnd 0.019394f
C2648 vdd.n1358 gnd 0.006163f
C2649 vdd.n1359 gnd 0.01126f
C2650 vdd.n1360 gnd 0.01126f
C2651 vdd.n1361 gnd 0.01126f
C2652 vdd.n1362 gnd 0.009063f
C2653 vdd.n1363 gnd 0.009063f
C2654 vdd.n1364 gnd 0.009063f
C2655 vdd.n1365 gnd 0.01126f
C2656 vdd.n1366 gnd 0.01126f
C2657 vdd.n1367 gnd 0.01126f
C2658 vdd.n1368 gnd 0.009063f
C2659 vdd.n1369 gnd 0.009063f
C2660 vdd.n1370 gnd 0.009063f
C2661 vdd.n1371 gnd 0.01126f
C2662 vdd.n1372 gnd 0.01126f
C2663 vdd.n1373 gnd 0.01126f
C2664 vdd.n1374 gnd 0.009063f
C2665 vdd.n1375 gnd 0.009063f
C2666 vdd.n1376 gnd 0.009063f
C2667 vdd.n1377 gnd 0.01126f
C2668 vdd.n1378 gnd 0.01126f
C2669 vdd.n1379 gnd 0.01126f
C2670 vdd.n1380 gnd 0.009063f
C2671 vdd.n1381 gnd 0.009063f
C2672 vdd.n1382 gnd 0.009063f
C2673 vdd.n1383 gnd 0.01126f
C2674 vdd.n1384 gnd 0.01126f
C2675 vdd.n1385 gnd 0.01126f
C2676 vdd.n1386 gnd 0.009063f
C2677 vdd.n1387 gnd 0.009063f
C2678 vdd.n1388 gnd 0.007567f
C2679 vdd.n1389 gnd 0.01126f
C2680 vdd.n1390 gnd 0.01126f
C2681 vdd.n1391 gnd 0.01126f
C2682 vdd.n1392 gnd 0.007567f
C2683 vdd.n1393 gnd 0.009063f
C2684 vdd.n1394 gnd 0.009063f
C2685 vdd.n1395 gnd 0.01126f
C2686 vdd.n1396 gnd 0.01126f
C2687 vdd.n1397 gnd 0.01126f
C2688 vdd.n1398 gnd 0.009063f
C2689 vdd.n1399 gnd 0.009063f
C2690 vdd.n1400 gnd 0.009063f
C2691 vdd.n1401 gnd 0.01126f
C2692 vdd.n1402 gnd 0.01126f
C2693 vdd.n1403 gnd 0.01126f
C2694 vdd.n1404 gnd 0.009063f
C2695 vdd.n1405 gnd 0.009063f
C2696 vdd.n1406 gnd 0.009063f
C2697 vdd.n1407 gnd 0.01126f
C2698 vdd.n1408 gnd 0.01126f
C2699 vdd.n1409 gnd 0.01126f
C2700 vdd.n1410 gnd 0.009063f
C2701 vdd.n1411 gnd 0.009063f
C2702 vdd.n1412 gnd 0.009063f
C2703 vdd.n1413 gnd 0.01126f
C2704 vdd.n1414 gnd 0.01126f
C2705 vdd.n1415 gnd 0.01126f
C2706 vdd.n1416 gnd 0.009063f
C2707 vdd.n1417 gnd 0.01126f
C2708 vdd.n1418 gnd 2.72713f
C2709 vdd.n1420 gnd 0.027822f
C2710 vdd.n1421 gnd 0.007522f
C2711 vdd.n1422 gnd 0.027822f
C2712 vdd.n1423 gnd 0.027238f
C2713 vdd.n1424 gnd 0.01126f
C2714 vdd.n1425 gnd 0.009063f
C2715 vdd.n1426 gnd 0.01126f
C2716 vdd.n1427 gnd 0.581097f
C2717 vdd.n1428 gnd 0.01126f
C2718 vdd.n1429 gnd 0.009063f
C2719 vdd.n1430 gnd 0.01126f
C2720 vdd.n1431 gnd 0.01126f
C2721 vdd.n1432 gnd 0.01126f
C2722 vdd.n1433 gnd 0.009063f
C2723 vdd.n1434 gnd 0.01126f
C2724 vdd.n1435 gnd 1.05288f
C2725 vdd.n1436 gnd 1.15069f
C2726 vdd.n1437 gnd 0.01126f
C2727 vdd.n1438 gnd 0.009063f
C2728 vdd.n1439 gnd 0.01126f
C2729 vdd.n1440 gnd 0.01126f
C2730 vdd.n1441 gnd 0.01126f
C2731 vdd.n1442 gnd 0.009063f
C2732 vdd.n1443 gnd 0.01126f
C2733 vdd.n1444 gnd 0.673151f
C2734 vdd.n1445 gnd 0.01126f
C2735 vdd.n1446 gnd 0.009063f
C2736 vdd.n1447 gnd 0.01126f
C2737 vdd.n1448 gnd 0.01126f
C2738 vdd.n1449 gnd 0.01126f
C2739 vdd.n1450 gnd 0.009063f
C2740 vdd.n1451 gnd 0.01126f
C2741 vdd.n1452 gnd 0.661645f
C2742 vdd.n1453 gnd 0.868768f
C2743 vdd.n1454 gnd 0.01126f
C2744 vdd.n1455 gnd 0.009063f
C2745 vdd.n1456 gnd 0.01126f
C2746 vdd.n1457 gnd 0.01126f
C2747 vdd.n1458 gnd 0.01126f
C2748 vdd.n1459 gnd 0.009063f
C2749 vdd.n1460 gnd 0.01126f
C2750 vdd.n1461 gnd 0.95507f
C2751 vdd.n1462 gnd 0.01126f
C2752 vdd.n1463 gnd 0.009063f
C2753 vdd.n1464 gnd 0.01126f
C2754 vdd.n1465 gnd 0.01126f
C2755 vdd.n1466 gnd 0.01126f
C2756 vdd.n1467 gnd 0.009063f
C2757 vdd.n1468 gnd 0.01126f
C2758 vdd.t92 gnd 0.575343f
C2759 vdd.n1469 gnd 0.845754f
C2760 vdd.n1470 gnd 0.01126f
C2761 vdd.n1471 gnd 0.009063f
C2762 vdd.n1472 gnd 0.01126f
C2763 vdd.n1473 gnd 0.01126f
C2764 vdd.n1474 gnd 0.01126f
C2765 vdd.n1475 gnd 0.009063f
C2766 vdd.n1476 gnd 0.01126f
C2767 vdd.n1477 gnd 0.650138f
C2768 vdd.n1478 gnd 0.01126f
C2769 vdd.n1479 gnd 0.009063f
C2770 vdd.n1480 gnd 0.01126f
C2771 vdd.n1481 gnd 0.01126f
C2772 vdd.n1482 gnd 0.01126f
C2773 vdd.n1483 gnd 0.009063f
C2774 vdd.n1484 gnd 0.01126f
C2775 vdd.n1485 gnd 0.834248f
C2776 vdd.n1486 gnd 0.696165f
C2777 vdd.n1487 gnd 0.01126f
C2778 vdd.n1488 gnd 0.009063f
C2779 vdd.n1489 gnd 0.01126f
C2780 vdd.n1490 gnd 0.01126f
C2781 vdd.n1491 gnd 0.01126f
C2782 vdd.n1492 gnd 0.009063f
C2783 vdd.n1493 gnd 0.01126f
C2784 vdd.n1494 gnd 0.891782f
C2785 vdd.n1495 gnd 0.01126f
C2786 vdd.n1496 gnd 0.009063f
C2787 vdd.n1497 gnd 0.01126f
C2788 vdd.n1498 gnd 0.01126f
C2789 vdd.n1499 gnd 0.01126f
C2790 vdd.n1500 gnd 0.009063f
C2791 vdd.n1501 gnd 0.01126f
C2792 vdd.t6 gnd 0.575343f
C2793 vdd.n1502 gnd 0.95507f
C2794 vdd.n1503 gnd 0.01126f
C2795 vdd.n1504 gnd 0.009063f
C2796 vdd.n1505 gnd 0.01126f
C2797 vdd.n1506 gnd 0.008654f
C2798 vdd.n1507 gnd 0.006179f
C2799 vdd.n1508 gnd 0.005734f
C2800 vdd.n1509 gnd 0.003172f
C2801 vdd.n1510 gnd 0.007283f
C2802 vdd.n1511 gnd 0.003081f
C2803 vdd.n1512 gnd 0.003263f
C2804 vdd.n1513 gnd 0.005734f
C2805 vdd.n1514 gnd 0.003081f
C2806 vdd.n1515 gnd 0.007283f
C2807 vdd.n1516 gnd 0.003263f
C2808 vdd.n1517 gnd 0.005734f
C2809 vdd.n1518 gnd 0.003081f
C2810 vdd.n1519 gnd 0.005462f
C2811 vdd.n1520 gnd 0.005479f
C2812 vdd.t44 gnd 0.015647f
C2813 vdd.n1521 gnd 0.034815f
C2814 vdd.n1522 gnd 0.181183f
C2815 vdd.n1523 gnd 0.003081f
C2816 vdd.n1524 gnd 0.003263f
C2817 vdd.n1525 gnd 0.007283f
C2818 vdd.n1526 gnd 0.007283f
C2819 vdd.n1527 gnd 0.003263f
C2820 vdd.n1528 gnd 0.003081f
C2821 vdd.n1529 gnd 0.005734f
C2822 vdd.n1530 gnd 0.005734f
C2823 vdd.n1531 gnd 0.003081f
C2824 vdd.n1532 gnd 0.003263f
C2825 vdd.n1533 gnd 0.007283f
C2826 vdd.n1534 gnd 0.007283f
C2827 vdd.n1535 gnd 0.003263f
C2828 vdd.n1536 gnd 0.003081f
C2829 vdd.n1537 gnd 0.005734f
C2830 vdd.n1538 gnd 0.005734f
C2831 vdd.n1539 gnd 0.003081f
C2832 vdd.n1540 gnd 0.003263f
C2833 vdd.n1541 gnd 0.007283f
C2834 vdd.n1542 gnd 0.007283f
C2835 vdd.n1543 gnd 0.017219f
C2836 vdd.n1544 gnd 0.003172f
C2837 vdd.n1545 gnd 0.003081f
C2838 vdd.n1546 gnd 0.014821f
C2839 vdd.n1547 gnd 0.010347f
C2840 vdd.t275 gnd 0.036251f
C2841 vdd.t257 gnd 0.036251f
C2842 vdd.n1548 gnd 0.24914f
C2843 vdd.n1549 gnd 0.195911f
C2844 vdd.t65 gnd 0.036251f
C2845 vdd.t246 gnd 0.036251f
C2846 vdd.n1550 gnd 0.24914f
C2847 vdd.n1551 gnd 0.158099f
C2848 vdd.t70 gnd 0.036251f
C2849 vdd.t116 gnd 0.036251f
C2850 vdd.n1552 gnd 0.24914f
C2851 vdd.n1553 gnd 0.158099f
C2852 vdd.t109 gnd 0.036251f
C2853 vdd.t35 gnd 0.036251f
C2854 vdd.n1554 gnd 0.24914f
C2855 vdd.n1555 gnd 0.158099f
C2856 vdd.t98 gnd 0.036251f
C2857 vdd.t48 gnd 0.036251f
C2858 vdd.n1556 gnd 0.24914f
C2859 vdd.n1557 gnd 0.158099f
C2860 vdd.t77 gnd 0.036251f
C2861 vdd.t49 gnd 0.036251f
C2862 vdd.n1558 gnd 0.24914f
C2863 vdd.n1559 gnd 0.158099f
C2864 vdd.t53 gnd 0.036251f
C2865 vdd.t249 gnd 0.036251f
C2866 vdd.n1560 gnd 0.24914f
C2867 vdd.n1561 gnd 0.158099f
C2868 vdd.t79 gnd 0.036251f
C2869 vdd.t261 gnd 0.036251f
C2870 vdd.n1562 gnd 0.24914f
C2871 vdd.n1563 gnd 0.158099f
C2872 vdd.t289 gnd 0.036251f
C2873 vdd.t263 gnd 0.036251f
C2874 vdd.n1564 gnd 0.24914f
C2875 vdd.n1565 gnd 0.158099f
C2876 vdd.n1566 gnd 0.006179f
C2877 vdd.n1567 gnd 0.005734f
C2878 vdd.n1568 gnd 0.003172f
C2879 vdd.n1569 gnd 0.007283f
C2880 vdd.n1570 gnd 0.003081f
C2881 vdd.n1571 gnd 0.003263f
C2882 vdd.n1572 gnd 0.005734f
C2883 vdd.n1573 gnd 0.003081f
C2884 vdd.n1574 gnd 0.007283f
C2885 vdd.n1575 gnd 0.003263f
C2886 vdd.n1576 gnd 0.005734f
C2887 vdd.n1577 gnd 0.003081f
C2888 vdd.n1578 gnd 0.005462f
C2889 vdd.n1579 gnd 0.005479f
C2890 vdd.t101 gnd 0.015647f
C2891 vdd.n1580 gnd 0.034815f
C2892 vdd.n1581 gnd 0.181183f
C2893 vdd.n1582 gnd 0.003081f
C2894 vdd.n1583 gnd 0.003263f
C2895 vdd.n1584 gnd 0.007283f
C2896 vdd.n1585 gnd 0.007283f
C2897 vdd.n1586 gnd 0.003263f
C2898 vdd.n1587 gnd 0.003081f
C2899 vdd.n1588 gnd 0.005734f
C2900 vdd.n1589 gnd 0.005734f
C2901 vdd.n1590 gnd 0.003081f
C2902 vdd.n1591 gnd 0.003263f
C2903 vdd.n1592 gnd 0.007283f
C2904 vdd.n1593 gnd 0.007283f
C2905 vdd.n1594 gnd 0.003263f
C2906 vdd.n1595 gnd 0.003081f
C2907 vdd.n1596 gnd 0.005734f
C2908 vdd.n1597 gnd 0.005734f
C2909 vdd.n1598 gnd 0.003081f
C2910 vdd.n1599 gnd 0.003263f
C2911 vdd.n1600 gnd 0.007283f
C2912 vdd.n1601 gnd 0.007283f
C2913 vdd.n1602 gnd 0.017219f
C2914 vdd.n1603 gnd 0.003172f
C2915 vdd.n1604 gnd 0.003081f
C2916 vdd.n1605 gnd 0.014821f
C2917 vdd.n1606 gnd 0.010023f
C2918 vdd.n1607 gnd 0.117626f
C2919 vdd.n1608 gnd 0.006179f
C2920 vdd.n1609 gnd 0.005734f
C2921 vdd.n1610 gnd 0.003172f
C2922 vdd.n1611 gnd 0.007283f
C2923 vdd.n1612 gnd 0.003081f
C2924 vdd.n1613 gnd 0.003263f
C2925 vdd.n1614 gnd 0.005734f
C2926 vdd.n1615 gnd 0.003081f
C2927 vdd.n1616 gnd 0.007283f
C2928 vdd.n1617 gnd 0.003263f
C2929 vdd.n1618 gnd 0.005734f
C2930 vdd.n1619 gnd 0.003081f
C2931 vdd.n1620 gnd 0.005462f
C2932 vdd.n1621 gnd 0.005479f
C2933 vdd.t247 gnd 0.015647f
C2934 vdd.n1622 gnd 0.034815f
C2935 vdd.n1623 gnd 0.181183f
C2936 vdd.n1624 gnd 0.003081f
C2937 vdd.n1625 gnd 0.003263f
C2938 vdd.n1626 gnd 0.007283f
C2939 vdd.n1627 gnd 0.007283f
C2940 vdd.n1628 gnd 0.003263f
C2941 vdd.n1629 gnd 0.003081f
C2942 vdd.n1630 gnd 0.005734f
C2943 vdd.n1631 gnd 0.005734f
C2944 vdd.n1632 gnd 0.003081f
C2945 vdd.n1633 gnd 0.003263f
C2946 vdd.n1634 gnd 0.007283f
C2947 vdd.n1635 gnd 0.007283f
C2948 vdd.n1636 gnd 0.003263f
C2949 vdd.n1637 gnd 0.003081f
C2950 vdd.n1638 gnd 0.005734f
C2951 vdd.n1639 gnd 0.005734f
C2952 vdd.n1640 gnd 0.003081f
C2953 vdd.n1641 gnd 0.003263f
C2954 vdd.n1642 gnd 0.007283f
C2955 vdd.n1643 gnd 0.007283f
C2956 vdd.n1644 gnd 0.017219f
C2957 vdd.n1645 gnd 0.003172f
C2958 vdd.n1646 gnd 0.003081f
C2959 vdd.n1647 gnd 0.014821f
C2960 vdd.n1648 gnd 0.010347f
C2961 vdd.t46 gnd 0.036251f
C2962 vdd.t294 gnd 0.036251f
C2963 vdd.n1649 gnd 0.24914f
C2964 vdd.n1650 gnd 0.195911f
C2965 vdd.t114 gnd 0.036251f
C2966 vdd.t83 gnd 0.036251f
C2967 vdd.n1651 gnd 0.24914f
C2968 vdd.n1652 gnd 0.158099f
C2969 vdd.t72 gnd 0.036251f
C2970 vdd.t42 gnd 0.036251f
C2971 vdd.n1653 gnd 0.24914f
C2972 vdd.n1654 gnd 0.158099f
C2973 vdd.t258 gnd 0.036251f
C2974 vdd.t84 gnd 0.036251f
C2975 vdd.n1655 gnd 0.24914f
C2976 vdd.n1656 gnd 0.158099f
C2977 vdd.t7 gnd 0.036251f
C2978 vdd.t63 gnd 0.036251f
C2979 vdd.n1657 gnd 0.24914f
C2980 vdd.n1658 gnd 0.158099f
C2981 vdd.t262 gnd 0.036251f
C2982 vdd.t5 gnd 0.036251f
C2983 vdd.n1659 gnd 0.24914f
C2984 vdd.n1660 gnd 0.158099f
C2985 vdd.t276 gnd 0.036251f
C2986 vdd.t277 gnd 0.036251f
C2987 vdd.n1661 gnd 0.24914f
C2988 vdd.n1662 gnd 0.158099f
C2989 vdd.t96 gnd 0.036251f
C2990 vdd.t254 gnd 0.036251f
C2991 vdd.n1663 gnd 0.24914f
C2992 vdd.n1664 gnd 0.158099f
C2993 vdd.t253 gnd 0.036251f
C2994 vdd.t75 gnd 0.036251f
C2995 vdd.n1665 gnd 0.24914f
C2996 vdd.n1666 gnd 0.158099f
C2997 vdd.n1667 gnd 0.006179f
C2998 vdd.n1668 gnd 0.005734f
C2999 vdd.n1669 gnd 0.003172f
C3000 vdd.n1670 gnd 0.007283f
C3001 vdd.n1671 gnd 0.003081f
C3002 vdd.n1672 gnd 0.003263f
C3003 vdd.n1673 gnd 0.005734f
C3004 vdd.n1674 gnd 0.003081f
C3005 vdd.n1675 gnd 0.007283f
C3006 vdd.n1676 gnd 0.003263f
C3007 vdd.n1677 gnd 0.005734f
C3008 vdd.n1678 gnd 0.003081f
C3009 vdd.n1679 gnd 0.005462f
C3010 vdd.n1680 gnd 0.005479f
C3011 vdd.t283 gnd 0.015647f
C3012 vdd.n1681 gnd 0.034815f
C3013 vdd.n1682 gnd 0.181183f
C3014 vdd.n1683 gnd 0.003081f
C3015 vdd.n1684 gnd 0.003263f
C3016 vdd.n1685 gnd 0.007283f
C3017 vdd.n1686 gnd 0.007283f
C3018 vdd.n1687 gnd 0.003263f
C3019 vdd.n1688 gnd 0.003081f
C3020 vdd.n1689 gnd 0.005734f
C3021 vdd.n1690 gnd 0.005734f
C3022 vdd.n1691 gnd 0.003081f
C3023 vdd.n1692 gnd 0.003263f
C3024 vdd.n1693 gnd 0.007283f
C3025 vdd.n1694 gnd 0.007283f
C3026 vdd.n1695 gnd 0.003263f
C3027 vdd.n1696 gnd 0.003081f
C3028 vdd.n1697 gnd 0.005734f
C3029 vdd.n1698 gnd 0.005734f
C3030 vdd.n1699 gnd 0.003081f
C3031 vdd.n1700 gnd 0.003263f
C3032 vdd.n1701 gnd 0.007283f
C3033 vdd.n1702 gnd 0.007283f
C3034 vdd.n1703 gnd 0.017219f
C3035 vdd.n1704 gnd 0.003172f
C3036 vdd.n1705 gnd 0.003081f
C3037 vdd.n1706 gnd 0.014821f
C3038 vdd.n1707 gnd 0.010023f
C3039 vdd.n1708 gnd 0.069976f
C3040 vdd.n1709 gnd 0.252141f
C3041 vdd.n1710 gnd 0.006179f
C3042 vdd.n1711 gnd 0.005734f
C3043 vdd.n1712 gnd 0.003172f
C3044 vdd.n1713 gnd 0.007283f
C3045 vdd.n1714 gnd 0.003081f
C3046 vdd.n1715 gnd 0.003263f
C3047 vdd.n1716 gnd 0.005734f
C3048 vdd.n1717 gnd 0.003081f
C3049 vdd.n1718 gnd 0.007283f
C3050 vdd.n1719 gnd 0.003263f
C3051 vdd.n1720 gnd 0.005734f
C3052 vdd.n1721 gnd 0.003081f
C3053 vdd.n1722 gnd 0.005462f
C3054 vdd.n1723 gnd 0.005479f
C3055 vdd.t56 gnd 0.015647f
C3056 vdd.n1724 gnd 0.034815f
C3057 vdd.n1725 gnd 0.181183f
C3058 vdd.n1726 gnd 0.003081f
C3059 vdd.n1727 gnd 0.003263f
C3060 vdd.n1728 gnd 0.007283f
C3061 vdd.n1729 gnd 0.007283f
C3062 vdd.n1730 gnd 0.003263f
C3063 vdd.n1731 gnd 0.003081f
C3064 vdd.n1732 gnd 0.005734f
C3065 vdd.n1733 gnd 0.005734f
C3066 vdd.n1734 gnd 0.003081f
C3067 vdd.n1735 gnd 0.003263f
C3068 vdd.n1736 gnd 0.007283f
C3069 vdd.n1737 gnd 0.007283f
C3070 vdd.n1738 gnd 0.003263f
C3071 vdd.n1739 gnd 0.003081f
C3072 vdd.n1740 gnd 0.005734f
C3073 vdd.n1741 gnd 0.005734f
C3074 vdd.n1742 gnd 0.003081f
C3075 vdd.n1743 gnd 0.003263f
C3076 vdd.n1744 gnd 0.007283f
C3077 vdd.n1745 gnd 0.007283f
C3078 vdd.n1746 gnd 0.017219f
C3079 vdd.n1747 gnd 0.003172f
C3080 vdd.n1748 gnd 0.003081f
C3081 vdd.n1749 gnd 0.014821f
C3082 vdd.n1750 gnd 0.010347f
C3083 vdd.t62 gnd 0.036251f
C3084 vdd.t55 gnd 0.036251f
C3085 vdd.n1751 gnd 0.24914f
C3086 vdd.n1752 gnd 0.195911f
C3087 vdd.t259 gnd 0.036251f
C3088 vdd.t87 gnd 0.036251f
C3089 vdd.n1753 gnd 0.24914f
C3090 vdd.n1754 gnd 0.158099f
C3091 vdd.t110 gnd 0.036251f
C3092 vdd.t57 gnd 0.036251f
C3093 vdd.n1755 gnd 0.24914f
C3094 vdd.n1756 gnd 0.158099f
C3095 vdd.t11 gnd 0.036251f
C3096 vdd.t245 gnd 0.036251f
C3097 vdd.n1757 gnd 0.24914f
C3098 vdd.n1758 gnd 0.158099f
C3099 vdd.t281 gnd 0.036251f
C3100 vdd.t100 gnd 0.036251f
C3101 vdd.n1759 gnd 0.24914f
C3102 vdd.n1760 gnd 0.158099f
C3103 vdd.t270 gnd 0.036251f
C3104 vdd.t280 gnd 0.036251f
C3105 vdd.n1761 gnd 0.24914f
C3106 vdd.n1762 gnd 0.158099f
C3107 vdd.t118 gnd 0.036251f
C3108 vdd.t120 gnd 0.036251f
C3109 vdd.n1763 gnd 0.24914f
C3110 vdd.n1764 gnd 0.158099f
C3111 vdd.t99 gnd 0.036251f
C3112 vdd.t93 gnd 0.036251f
C3113 vdd.n1765 gnd 0.24914f
C3114 vdd.n1766 gnd 0.158099f
C3115 vdd.t260 gnd 0.036251f
C3116 vdd.t29 gnd 0.036251f
C3117 vdd.n1767 gnd 0.24914f
C3118 vdd.n1768 gnd 0.158099f
C3119 vdd.n1769 gnd 0.006179f
C3120 vdd.n1770 gnd 0.005734f
C3121 vdd.n1771 gnd 0.003172f
C3122 vdd.n1772 gnd 0.007283f
C3123 vdd.n1773 gnd 0.003081f
C3124 vdd.n1774 gnd 0.003263f
C3125 vdd.n1775 gnd 0.005734f
C3126 vdd.n1776 gnd 0.003081f
C3127 vdd.n1777 gnd 0.007283f
C3128 vdd.n1778 gnd 0.003263f
C3129 vdd.n1779 gnd 0.005734f
C3130 vdd.n1780 gnd 0.003081f
C3131 vdd.n1781 gnd 0.005462f
C3132 vdd.n1782 gnd 0.005479f
C3133 vdd.t59 gnd 0.015647f
C3134 vdd.n1783 gnd 0.034815f
C3135 vdd.n1784 gnd 0.181183f
C3136 vdd.n1785 gnd 0.003081f
C3137 vdd.n1786 gnd 0.003263f
C3138 vdd.n1787 gnd 0.007283f
C3139 vdd.n1788 gnd 0.007283f
C3140 vdd.n1789 gnd 0.003263f
C3141 vdd.n1790 gnd 0.003081f
C3142 vdd.n1791 gnd 0.005734f
C3143 vdd.n1792 gnd 0.005734f
C3144 vdd.n1793 gnd 0.003081f
C3145 vdd.n1794 gnd 0.003263f
C3146 vdd.n1795 gnd 0.007283f
C3147 vdd.n1796 gnd 0.007283f
C3148 vdd.n1797 gnd 0.003263f
C3149 vdd.n1798 gnd 0.003081f
C3150 vdd.n1799 gnd 0.005734f
C3151 vdd.n1800 gnd 0.005734f
C3152 vdd.n1801 gnd 0.003081f
C3153 vdd.n1802 gnd 0.003263f
C3154 vdd.n1803 gnd 0.007283f
C3155 vdd.n1804 gnd 0.007283f
C3156 vdd.n1805 gnd 0.017219f
C3157 vdd.n1806 gnd 0.003172f
C3158 vdd.n1807 gnd 0.003081f
C3159 vdd.n1808 gnd 0.014821f
C3160 vdd.n1809 gnd 0.010023f
C3161 vdd.n1810 gnd 0.069976f
C3162 vdd.n1811 gnd 0.288647f
C3163 vdd.n1812 gnd 2.89194f
C3164 vdd.n1813 gnd 0.664139f
C3165 vdd.n1814 gnd 0.008654f
C3166 vdd.n1815 gnd 0.009063f
C3167 vdd.n1816 gnd 0.01126f
C3168 vdd.n1817 gnd 0.822741f
C3169 vdd.n1818 gnd 0.01126f
C3170 vdd.n1819 gnd 0.009063f
C3171 vdd.n1820 gnd 0.01126f
C3172 vdd.n1821 gnd 0.01126f
C3173 vdd.n1822 gnd 0.01126f
C3174 vdd.n1823 gnd 0.009063f
C3175 vdd.n1824 gnd 0.01126f
C3176 vdd.n1825 gnd 0.95507f
C3177 vdd.t10 gnd 0.575343f
C3178 vdd.n1826 gnd 0.627124f
C3179 vdd.n1827 gnd 0.01126f
C3180 vdd.n1828 gnd 0.009063f
C3181 vdd.n1829 gnd 0.01126f
C3182 vdd.n1830 gnd 0.01126f
C3183 vdd.n1831 gnd 0.01126f
C3184 vdd.n1832 gnd 0.009063f
C3185 vdd.n1833 gnd 0.01126f
C3186 vdd.n1834 gnd 0.719179f
C3187 vdd.n1835 gnd 0.01126f
C3188 vdd.n1836 gnd 0.009063f
C3189 vdd.n1837 gnd 0.01126f
C3190 vdd.n1838 gnd 0.01126f
C3191 vdd.n1839 gnd 0.01126f
C3192 vdd.n1840 gnd 0.009063f
C3193 vdd.n1841 gnd 0.01126f
C3194 vdd.n1842 gnd 0.615617f
C3195 vdd.n1843 gnd 0.914796f
C3196 vdd.n1844 gnd 0.01126f
C3197 vdd.n1845 gnd 0.009063f
C3198 vdd.n1846 gnd 0.01126f
C3199 vdd.n1847 gnd 0.01126f
C3200 vdd.n1848 gnd 0.01126f
C3201 vdd.n1849 gnd 0.009063f
C3202 vdd.n1850 gnd 0.01126f
C3203 vdd.n1851 gnd 0.95507f
C3204 vdd.n1852 gnd 0.01126f
C3205 vdd.n1853 gnd 0.009063f
C3206 vdd.n1854 gnd 0.01126f
C3207 vdd.n1855 gnd 0.01126f
C3208 vdd.n1856 gnd 0.01126f
C3209 vdd.n1857 gnd 0.009063f
C3210 vdd.n1858 gnd 0.01126f
C3211 vdd.t82 gnd 0.575343f
C3212 vdd.n1859 gnd 0.799727f
C3213 vdd.n1860 gnd 0.01126f
C3214 vdd.n1861 gnd 0.009063f
C3215 vdd.n1862 gnd 0.01126f
C3216 vdd.n1863 gnd 0.01126f
C3217 vdd.n1864 gnd 0.01126f
C3218 vdd.n1865 gnd 0.009063f
C3219 vdd.n1866 gnd 0.01126f
C3220 vdd.n1867 gnd 0.60411f
C3221 vdd.n1868 gnd 0.01126f
C3222 vdd.n1869 gnd 0.009063f
C3223 vdd.n1870 gnd 0.01126f
C3224 vdd.n1871 gnd 0.01126f
C3225 vdd.n1872 gnd 0.01126f
C3226 vdd.n1873 gnd 0.009063f
C3227 vdd.n1874 gnd 0.01126f
C3228 vdd.n1875 gnd 0.78822f
C3229 vdd.n1876 gnd 0.742193f
C3230 vdd.n1877 gnd 0.01126f
C3231 vdd.n1878 gnd 0.009063f
C3232 vdd.n1879 gnd 0.01126f
C3233 vdd.n1880 gnd 0.01126f
C3234 vdd.n1881 gnd 0.01126f
C3235 vdd.n1882 gnd 0.009063f
C3236 vdd.n1883 gnd 0.01126f
C3237 vdd.n1884 gnd 0.937809f
C3238 vdd.n1885 gnd 0.01126f
C3239 vdd.n1886 gnd 0.009063f
C3240 vdd.n1887 gnd 0.01126f
C3241 vdd.n1888 gnd 0.01126f
C3242 vdd.n1889 gnd 0.027238f
C3243 vdd.n1890 gnd 0.01126f
C3244 vdd.n1891 gnd 0.01126f
C3245 vdd.n1892 gnd 0.009063f
C3246 vdd.n1893 gnd 0.01126f
C3247 vdd.n1894 gnd 0.696165f
C3248 vdd.n1895 gnd 1.15069f
C3249 vdd.n1896 gnd 0.01126f
C3250 vdd.n1897 gnd 0.009063f
C3251 vdd.n1898 gnd 0.01126f
C3252 vdd.n1899 gnd 0.01126f
C3253 vdd.n1900 gnd 0.009683f
C3254 vdd.n1901 gnd 0.009063f
C3255 vdd.n1903 gnd 0.01126f
C3256 vdd.n1905 gnd 0.009063f
C3257 vdd.n1906 gnd 0.01126f
C3258 vdd.n1907 gnd 0.009063f
C3259 vdd.n1909 gnd 0.01126f
C3260 vdd.n1910 gnd 0.009063f
C3261 vdd.n1911 gnd 0.01126f
C3262 vdd.n1912 gnd 0.01126f
C3263 vdd.n1913 gnd 0.01126f
C3264 vdd.n1914 gnd 0.01126f
C3265 vdd.n1915 gnd 0.01126f
C3266 vdd.n1916 gnd 0.009063f
C3267 vdd.n1918 gnd 0.01126f
C3268 vdd.n1919 gnd 0.01126f
C3269 vdd.n1920 gnd 0.01126f
C3270 vdd.n1921 gnd 0.01126f
C3271 vdd.n1922 gnd 0.01126f
C3272 vdd.n1923 gnd 0.009063f
C3273 vdd.n1925 gnd 0.01126f
C3274 vdd.n1926 gnd 0.01126f
C3275 vdd.n1927 gnd 0.01126f
C3276 vdd.n1928 gnd 0.01126f
C3277 vdd.n1929 gnd 0.007567f
C3278 vdd.t203 gnd 0.138524f
C3279 vdd.t202 gnd 0.148044f
C3280 vdd.t201 gnd 0.18091f
C3281 vdd.n1930 gnd 0.231901f
C3282 vdd.n1931 gnd 0.194839f
C3283 vdd.n1933 gnd 0.01126f
C3284 vdd.n1934 gnd 0.01126f
C3285 vdd.n1935 gnd 0.009063f
C3286 vdd.n1936 gnd 0.01126f
C3287 vdd.n1938 gnd 0.01126f
C3288 vdd.n1939 gnd 0.01126f
C3289 vdd.n1940 gnd 0.01126f
C3290 vdd.n1941 gnd 0.01126f
C3291 vdd.n1942 gnd 0.009063f
C3292 vdd.n1944 gnd 0.01126f
C3293 vdd.n1945 gnd 0.01126f
C3294 vdd.n1946 gnd 0.01126f
C3295 vdd.n1947 gnd 0.01126f
C3296 vdd.n1948 gnd 0.01126f
C3297 vdd.n1949 gnd 0.009063f
C3298 vdd.n1951 gnd 0.01126f
C3299 vdd.n1952 gnd 0.01126f
C3300 vdd.n1953 gnd 0.01126f
C3301 vdd.n1954 gnd 0.01126f
C3302 vdd.n1955 gnd 0.01126f
C3303 vdd.n1956 gnd 0.009063f
C3304 vdd.n1958 gnd 0.01126f
C3305 vdd.n1959 gnd 0.01126f
C3306 vdd.n1960 gnd 0.01126f
C3307 vdd.n1961 gnd 0.01126f
C3308 vdd.n1962 gnd 0.01126f
C3309 vdd.n1963 gnd 0.009063f
C3310 vdd.n1965 gnd 0.01126f
C3311 vdd.n1966 gnd 0.01126f
C3312 vdd.n1967 gnd 0.01126f
C3313 vdd.n1968 gnd 0.01126f
C3314 vdd.n1969 gnd 0.008972f
C3315 vdd.t190 gnd 0.138524f
C3316 vdd.t189 gnd 0.148044f
C3317 vdd.t188 gnd 0.18091f
C3318 vdd.n1970 gnd 0.231901f
C3319 vdd.n1971 gnd 0.194839f
C3320 vdd.n1973 gnd 0.01126f
C3321 vdd.n1974 gnd 0.01126f
C3322 vdd.n1975 gnd 0.009063f
C3323 vdd.n1976 gnd 0.01126f
C3324 vdd.n1978 gnd 0.01126f
C3325 vdd.n1979 gnd 0.01126f
C3326 vdd.n1980 gnd 0.01126f
C3327 vdd.n1981 gnd 0.01126f
C3328 vdd.n1982 gnd 0.009063f
C3329 vdd.n1984 gnd 0.01126f
C3330 vdd.n1985 gnd 0.01126f
C3331 vdd.n1986 gnd 0.01126f
C3332 vdd.n1987 gnd 0.01126f
C3333 vdd.n1988 gnd 0.01126f
C3334 vdd.n1989 gnd 0.009063f
C3335 vdd.n1991 gnd 0.01126f
C3336 vdd.n1992 gnd 0.01126f
C3337 vdd.n1993 gnd 0.01126f
C3338 vdd.n1994 gnd 0.01126f
C3339 vdd.n1995 gnd 0.01126f
C3340 vdd.n1996 gnd 0.01126f
C3341 vdd.n1997 gnd 0.009063f
C3342 vdd.n1999 gnd 0.01126f
C3343 vdd.n2001 gnd 0.01126f
C3344 vdd.n2002 gnd 0.009063f
C3345 vdd.n2003 gnd 0.009063f
C3346 vdd.n2004 gnd 0.01126f
C3347 vdd.n2006 gnd 0.01126f
C3348 vdd.n2007 gnd 0.009063f
C3349 vdd.n2008 gnd 0.009063f
C3350 vdd.n2009 gnd 0.01126f
C3351 vdd.n2011 gnd 0.01126f
C3352 vdd.n2012 gnd 0.01126f
C3353 vdd.n2013 gnd 0.009063f
C3354 vdd.n2014 gnd 0.009063f
C3355 vdd.n2015 gnd 0.009063f
C3356 vdd.n2016 gnd 0.01126f
C3357 vdd.n2018 gnd 0.01126f
C3358 vdd.n2019 gnd 0.01126f
C3359 vdd.n2020 gnd 0.009063f
C3360 vdd.n2021 gnd 0.009063f
C3361 vdd.n2022 gnd 0.009063f
C3362 vdd.n2023 gnd 0.01126f
C3363 vdd.n2025 gnd 0.01126f
C3364 vdd.n2026 gnd 0.01126f
C3365 vdd.n2027 gnd 0.009063f
C3366 vdd.n2028 gnd 0.009063f
C3367 vdd.n2029 gnd 0.009063f
C3368 vdd.n2030 gnd 0.01126f
C3369 vdd.n2032 gnd 0.01126f
C3370 vdd.n2033 gnd 0.01126f
C3371 vdd.n2034 gnd 0.009063f
C3372 vdd.n2035 gnd 0.01126f
C3373 vdd.n2036 gnd 0.01126f
C3374 vdd.n2037 gnd 0.01126f
C3375 vdd.n2038 gnd 0.018488f
C3376 vdd.n2039 gnd 0.006163f
C3377 vdd.n2040 gnd 0.009063f
C3378 vdd.n2041 gnd 0.01126f
C3379 vdd.n2043 gnd 0.01126f
C3380 vdd.n2044 gnd 0.01126f
C3381 vdd.n2045 gnd 0.009063f
C3382 vdd.n2046 gnd 0.009063f
C3383 vdd.n2047 gnd 0.009063f
C3384 vdd.n2048 gnd 0.01126f
C3385 vdd.n2050 gnd 0.01126f
C3386 vdd.n2051 gnd 0.01126f
C3387 vdd.n2052 gnd 0.009063f
C3388 vdd.n2053 gnd 0.009063f
C3389 vdd.n2054 gnd 0.009063f
C3390 vdd.n2055 gnd 0.01126f
C3391 vdd.n2057 gnd 0.01126f
C3392 vdd.n2058 gnd 0.01126f
C3393 vdd.n2059 gnd 0.009063f
C3394 vdd.n2060 gnd 0.009063f
C3395 vdd.n2061 gnd 0.009063f
C3396 vdd.n2062 gnd 0.01126f
C3397 vdd.n2064 gnd 0.01126f
C3398 vdd.n2065 gnd 0.01126f
C3399 vdd.n2066 gnd 0.009063f
C3400 vdd.n2067 gnd 0.009063f
C3401 vdd.n2068 gnd 0.009063f
C3402 vdd.n2069 gnd 0.01126f
C3403 vdd.n2071 gnd 0.01126f
C3404 vdd.n2072 gnd 0.01126f
C3405 vdd.n2073 gnd 0.009063f
C3406 vdd.n2074 gnd 0.01126f
C3407 vdd.n2075 gnd 0.01126f
C3408 vdd.n2076 gnd 0.01126f
C3409 vdd.n2077 gnd 0.018488f
C3410 vdd.n2078 gnd 0.007567f
C3411 vdd.n2079 gnd 0.009063f
C3412 vdd.n2080 gnd 0.01126f
C3413 vdd.n2082 gnd 0.01126f
C3414 vdd.n2083 gnd 0.01126f
C3415 vdd.n2084 gnd 0.009063f
C3416 vdd.n2085 gnd 0.009063f
C3417 vdd.n2086 gnd 0.009063f
C3418 vdd.n2087 gnd 0.01126f
C3419 vdd.n2089 gnd 0.01126f
C3420 vdd.n2090 gnd 0.01126f
C3421 vdd.n2091 gnd 0.009063f
C3422 vdd.n2092 gnd 0.009063f
C3423 vdd.n2093 gnd 0.009063f
C3424 vdd.n2094 gnd 0.01126f
C3425 vdd.n2096 gnd 0.01126f
C3426 vdd.n2097 gnd 0.01126f
C3427 vdd.n2099 gnd 0.01126f
C3428 vdd.n2100 gnd 0.009063f
C3429 vdd.n2101 gnd 0.007206f
C3430 vdd.n2102 gnd 0.007657f
C3431 vdd.n2103 gnd 0.007657f
C3432 vdd.n2104 gnd 0.007657f
C3433 vdd.n2105 gnd 0.007657f
C3434 vdd.n2106 gnd 0.007657f
C3435 vdd.n2107 gnd 0.007657f
C3436 vdd.n2108 gnd 0.007657f
C3437 vdd.n2109 gnd 0.007657f
C3438 vdd.n2111 gnd 0.007657f
C3439 vdd.n2112 gnd 0.007657f
C3440 vdd.n2113 gnd 0.007657f
C3441 vdd.n2114 gnd 0.007657f
C3442 vdd.n2115 gnd 0.007657f
C3443 vdd.n2117 gnd 0.007657f
C3444 vdd.n2119 gnd 0.007657f
C3445 vdd.n2120 gnd 0.007657f
C3446 vdd.n2121 gnd 0.007657f
C3447 vdd.n2122 gnd 0.007657f
C3448 vdd.n2123 gnd 0.007657f
C3449 vdd.n2125 gnd 0.007657f
C3450 vdd.n2127 gnd 0.007657f
C3451 vdd.n2128 gnd 0.007657f
C3452 vdd.n2129 gnd 0.007657f
C3453 vdd.n2130 gnd 0.007657f
C3454 vdd.n2131 gnd 0.007657f
C3455 vdd.n2133 gnd 0.007657f
C3456 vdd.n2135 gnd 0.007657f
C3457 vdd.n2136 gnd 0.007657f
C3458 vdd.n2137 gnd 0.007657f
C3459 vdd.n2138 gnd 0.007657f
C3460 vdd.n2139 gnd 0.007657f
C3461 vdd.n2141 gnd 0.007657f
C3462 vdd.n2142 gnd 0.007657f
C3463 vdd.n2143 gnd 0.007657f
C3464 vdd.n2144 gnd 0.007657f
C3465 vdd.n2145 gnd 0.007657f
C3466 vdd.n2146 gnd 0.007657f
C3467 vdd.n2147 gnd 0.007657f
C3468 vdd.n2148 gnd 0.007657f
C3469 vdd.n2149 gnd 0.005574f
C3470 vdd.n2150 gnd 0.007657f
C3471 vdd.t243 gnd 0.309402f
C3472 vdd.t244 gnd 0.316711f
C3473 vdd.t242 gnd 0.201989f
C3474 vdd.n2151 gnd 0.109164f
C3475 vdd.n2152 gnd 0.061921f
C3476 vdd.n2153 gnd 0.010943f
C3477 vdd.n2154 gnd 0.007657f
C3478 vdd.n2155 gnd 0.007657f
C3479 vdd.n2156 gnd 0.466028f
C3480 vdd.n2157 gnd 0.007657f
C3481 vdd.n2158 gnd 0.007657f
C3482 vdd.n2159 gnd 0.007657f
C3483 vdd.n2160 gnd 0.007657f
C3484 vdd.n2161 gnd 0.007657f
C3485 vdd.n2162 gnd 0.007657f
C3486 vdd.n2163 gnd 0.007657f
C3487 vdd.n2164 gnd 0.007657f
C3488 vdd.n2165 gnd 0.007657f
C3489 vdd.n2166 gnd 0.007657f
C3490 vdd.n2167 gnd 0.007657f
C3491 vdd.n2168 gnd 0.007657f
C3492 vdd.n2169 gnd 0.007657f
C3493 vdd.n2170 gnd 0.007657f
C3494 vdd.n2171 gnd 0.007657f
C3495 vdd.n2172 gnd 0.007657f
C3496 vdd.n2173 gnd 0.007657f
C3497 vdd.n2174 gnd 0.007657f
C3498 vdd.n2175 gnd 0.007657f
C3499 vdd.n2176 gnd 0.007657f
C3500 vdd.t221 gnd 0.309402f
C3501 vdd.t222 gnd 0.316711f
C3502 vdd.t219 gnd 0.201989f
C3503 vdd.n2177 gnd 0.109164f
C3504 vdd.n2178 gnd 0.061921f
C3505 vdd.n2179 gnd 0.007657f
C3506 vdd.n2180 gnd 0.007657f
C3507 vdd.n2181 gnd 0.007657f
C3508 vdd.n2182 gnd 0.007657f
C3509 vdd.n2183 gnd 0.007657f
C3510 vdd.n2184 gnd 0.007657f
C3511 vdd.n2186 gnd 0.007657f
C3512 vdd.n2187 gnd 0.007657f
C3513 vdd.n2188 gnd 0.007657f
C3514 vdd.n2189 gnd 0.007657f
C3515 vdd.n2191 gnd 0.007657f
C3516 vdd.n2193 gnd 0.007657f
C3517 vdd.n2194 gnd 0.007657f
C3518 vdd.n2195 gnd 0.007657f
C3519 vdd.n2196 gnd 0.007657f
C3520 vdd.n2197 gnd 0.007657f
C3521 vdd.n2199 gnd 0.007657f
C3522 vdd.n2201 gnd 0.007657f
C3523 vdd.n2202 gnd 0.007657f
C3524 vdd.n2203 gnd 0.007657f
C3525 vdd.n2204 gnd 0.007657f
C3526 vdd.n2205 gnd 0.007657f
C3527 vdd.n2207 gnd 0.007657f
C3528 vdd.n2209 gnd 0.007657f
C3529 vdd.n2210 gnd 0.007657f
C3530 vdd.n2211 gnd 0.005574f
C3531 vdd.n2212 gnd 0.010943f
C3532 vdd.n2213 gnd 0.005911f
C3533 vdd.n2214 gnd 0.007657f
C3534 vdd.n2216 gnd 0.007657f
C3535 vdd.n2217 gnd 0.018168f
C3536 vdd.n2218 gnd 0.018168f
C3537 vdd.n2219 gnd 0.016963f
C3538 vdd.n2220 gnd 0.007657f
C3539 vdd.n2221 gnd 0.007657f
C3540 vdd.n2222 gnd 0.007657f
C3541 vdd.n2223 gnd 0.007657f
C3542 vdd.n2224 gnd 0.007657f
C3543 vdd.n2225 gnd 0.007657f
C3544 vdd.n2226 gnd 0.007657f
C3545 vdd.n2227 gnd 0.007657f
C3546 vdd.n2228 gnd 0.007657f
C3547 vdd.n2229 gnd 0.007657f
C3548 vdd.n2230 gnd 0.007657f
C3549 vdd.n2231 gnd 0.007657f
C3550 vdd.n2232 gnd 0.007657f
C3551 vdd.n2233 gnd 0.007657f
C3552 vdd.n2234 gnd 0.007657f
C3553 vdd.n2235 gnd 0.007657f
C3554 vdd.n2236 gnd 0.007657f
C3555 vdd.n2237 gnd 0.007657f
C3556 vdd.n2238 gnd 0.007657f
C3557 vdd.n2239 gnd 0.007657f
C3558 vdd.n2240 gnd 0.007657f
C3559 vdd.n2241 gnd 0.007657f
C3560 vdd.n2242 gnd 0.007657f
C3561 vdd.n2243 gnd 0.007657f
C3562 vdd.n2244 gnd 0.007657f
C3563 vdd.n2245 gnd 0.007657f
C3564 vdd.n2246 gnd 0.007657f
C3565 vdd.n2247 gnd 0.007657f
C3566 vdd.n2248 gnd 0.007657f
C3567 vdd.n2249 gnd 0.007657f
C3568 vdd.n2250 gnd 0.007657f
C3569 vdd.n2251 gnd 0.007657f
C3570 vdd.n2252 gnd 0.007657f
C3571 vdd.n2253 gnd 0.007657f
C3572 vdd.n2254 gnd 0.007657f
C3573 vdd.n2255 gnd 0.007657f
C3574 vdd.n2256 gnd 0.007657f
C3575 vdd.n2257 gnd 0.247398f
C3576 vdd.n2258 gnd 0.007657f
C3577 vdd.n2259 gnd 0.007657f
C3578 vdd.n2260 gnd 0.007657f
C3579 vdd.n2261 gnd 0.007657f
C3580 vdd.n2262 gnd 0.007657f
C3581 vdd.n2263 gnd 0.007657f
C3582 vdd.n2264 gnd 0.007657f
C3583 vdd.n2265 gnd 0.007657f
C3584 vdd.n2266 gnd 0.007657f
C3585 vdd.n2267 gnd 0.007657f
C3586 vdd.n2268 gnd 0.007657f
C3587 vdd.n2269 gnd 0.007657f
C3588 vdd.n2270 gnd 0.007657f
C3589 vdd.n2271 gnd 0.007657f
C3590 vdd.n2272 gnd 0.007657f
C3591 vdd.n2273 gnd 0.007657f
C3592 vdd.n2274 gnd 0.007657f
C3593 vdd.n2275 gnd 0.007657f
C3594 vdd.n2276 gnd 0.007657f
C3595 vdd.n2277 gnd 0.007657f
C3596 vdd.n2278 gnd 0.016963f
C3597 vdd.n2280 gnd 0.018168f
C3598 vdd.n2281 gnd 0.018168f
C3599 vdd.n2282 gnd 0.007657f
C3600 vdd.n2283 gnd 0.005911f
C3601 vdd.n2284 gnd 0.007657f
C3602 vdd.n2286 gnd 0.007657f
C3603 vdd.n2288 gnd 0.007657f
C3604 vdd.n2289 gnd 0.007657f
C3605 vdd.n2290 gnd 0.007657f
C3606 vdd.n2291 gnd 0.007657f
C3607 vdd.n2292 gnd 0.007657f
C3608 vdd.n2294 gnd 0.007657f
C3609 vdd.n2296 gnd 0.007657f
C3610 vdd.n2297 gnd 0.007657f
C3611 vdd.n2298 gnd 0.007657f
C3612 vdd.n2299 gnd 0.007657f
C3613 vdd.n2300 gnd 0.007657f
C3614 vdd.n2302 gnd 0.007657f
C3615 vdd.n2304 gnd 0.007657f
C3616 vdd.n2305 gnd 0.007657f
C3617 vdd.n2306 gnd 0.007657f
C3618 vdd.n2307 gnd 0.007657f
C3619 vdd.n2308 gnd 0.007657f
C3620 vdd.n2310 gnd 0.007657f
C3621 vdd.n2312 gnd 0.007657f
C3622 vdd.n2313 gnd 0.007657f
C3623 vdd.n2314 gnd 0.022838f
C3624 vdd.n2315 gnd 0.677016f
C3625 vdd.n2317 gnd 0.009063f
C3626 vdd.n2318 gnd 0.009063f
C3627 vdd.n2319 gnd 0.01126f
C3628 vdd.n2321 gnd 0.01126f
C3629 vdd.n2322 gnd 0.01126f
C3630 vdd.n2323 gnd 0.009063f
C3631 vdd.n2324 gnd 0.007522f
C3632 vdd.n2325 gnd 0.027822f
C3633 vdd.n2326 gnd 0.027238f
C3634 vdd.n2327 gnd 0.007522f
C3635 vdd.n2328 gnd 0.027238f
C3636 vdd.n2329 gnd 1.58219f
C3637 vdd.n2330 gnd 0.027238f
C3638 vdd.n2331 gnd 0.027822f
C3639 vdd.n2332 gnd 0.004305f
C3640 vdd.t179 gnd 0.138524f
C3641 vdd.t178 gnd 0.148044f
C3642 vdd.t176 gnd 0.18091f
C3643 vdd.n2333 gnd 0.231901f
C3644 vdd.n2334 gnd 0.194839f
C3645 vdd.n2335 gnd 0.013957f
C3646 vdd.n2336 gnd 0.004758f
C3647 vdd.n2337 gnd 0.009683f
C3648 vdd.n2338 gnd 0.677016f
C3649 vdd.n2339 gnd 0.022838f
C3650 vdd.n2340 gnd 0.007657f
C3651 vdd.n2341 gnd 0.007657f
C3652 vdd.n2342 gnd 0.007657f
C3653 vdd.n2344 gnd 0.007657f
C3654 vdd.n2346 gnd 0.007657f
C3655 vdd.n2347 gnd 0.007657f
C3656 vdd.n2348 gnd 0.007657f
C3657 vdd.n2349 gnd 0.007657f
C3658 vdd.n2350 gnd 0.007657f
C3659 vdd.n2352 gnd 0.007657f
C3660 vdd.n2354 gnd 0.007657f
C3661 vdd.n2355 gnd 0.007657f
C3662 vdd.n2356 gnd 0.007657f
C3663 vdd.n2357 gnd 0.007657f
C3664 vdd.n2358 gnd 0.007657f
C3665 vdd.n2360 gnd 0.007657f
C3666 vdd.n2362 gnd 0.007657f
C3667 vdd.n2363 gnd 0.007657f
C3668 vdd.n2364 gnd 0.007657f
C3669 vdd.n2365 gnd 0.007657f
C3670 vdd.n2366 gnd 0.007657f
C3671 vdd.n2368 gnd 0.007657f
C3672 vdd.n2370 gnd 0.007657f
C3673 vdd.n2371 gnd 0.007657f
C3674 vdd.n2372 gnd 0.018168f
C3675 vdd.n2373 gnd 0.016963f
C3676 vdd.n2374 gnd 0.016963f
C3677 vdd.n2375 gnd 1.12767f
C3678 vdd.n2376 gnd 0.016963f
C3679 vdd.n2377 gnd 0.016963f
C3680 vdd.n2378 gnd 0.007657f
C3681 vdd.n2379 gnd 0.007657f
C3682 vdd.n2380 gnd 0.007657f
C3683 vdd.n2381 gnd 0.489042f
C3684 vdd.n2382 gnd 0.007657f
C3685 vdd.n2383 gnd 0.007657f
C3686 vdd.n2384 gnd 0.007657f
C3687 vdd.n2385 gnd 0.007657f
C3688 vdd.n2386 gnd 0.007657f
C3689 vdd.n2387 gnd 0.782467f
C3690 vdd.n2388 gnd 0.007657f
C3691 vdd.n2389 gnd 0.007657f
C3692 vdd.n2390 gnd 0.007657f
C3693 vdd.n2391 gnd 0.007657f
C3694 vdd.n2392 gnd 0.007657f
C3695 vdd.n2393 gnd 0.782467f
C3696 vdd.n2394 gnd 0.007657f
C3697 vdd.n2395 gnd 0.007657f
C3698 vdd.n2396 gnd 0.006756f
C3699 vdd.n2397 gnd 0.02218f
C3700 vdd.n2398 gnd 0.004729f
C3701 vdd.n2399 gnd 0.007657f
C3702 vdd.n2400 gnd 0.431507f
C3703 vdd.n2401 gnd 0.007657f
C3704 vdd.n2402 gnd 0.007657f
C3705 vdd.n2403 gnd 0.007657f
C3706 vdd.n2404 gnd 0.007657f
C3707 vdd.n2405 gnd 0.007657f
C3708 vdd.n2406 gnd 0.523562f
C3709 vdd.n2407 gnd 0.007657f
C3710 vdd.n2408 gnd 0.007657f
C3711 vdd.n2409 gnd 0.007657f
C3712 vdd.n2410 gnd 0.007657f
C3713 vdd.n2411 gnd 0.007657f
C3714 vdd.n2412 gnd 0.696165f
C3715 vdd.n2413 gnd 0.007657f
C3716 vdd.n2414 gnd 0.007657f
C3717 vdd.n2415 gnd 0.007657f
C3718 vdd.n2416 gnd 0.007657f
C3719 vdd.n2417 gnd 0.007657f
C3720 vdd.n2418 gnd 0.621371f
C3721 vdd.n2419 gnd 0.007657f
C3722 vdd.n2420 gnd 0.007657f
C3723 vdd.n2421 gnd 0.007657f
C3724 vdd.n2422 gnd 0.007657f
C3725 vdd.n2423 gnd 0.007657f
C3726 vdd.n2424 gnd 0.448768f
C3727 vdd.n2425 gnd 0.007657f
C3728 vdd.n2426 gnd 0.007657f
C3729 vdd.n2427 gnd 0.007657f
C3730 vdd.n2428 gnd 0.007657f
C3731 vdd.n2429 gnd 0.007657f
C3732 vdd.n2430 gnd 0.247398f
C3733 vdd.n2431 gnd 0.007657f
C3734 vdd.n2432 gnd 0.007657f
C3735 vdd.n2433 gnd 0.007657f
C3736 vdd.n2434 gnd 0.007657f
C3737 vdd.n2435 gnd 0.007657f
C3738 vdd.n2436 gnd 0.431507f
C3739 vdd.n2437 gnd 0.007657f
C3740 vdd.n2438 gnd 0.007657f
C3741 vdd.n2439 gnd 0.007657f
C3742 vdd.n2440 gnd 0.007657f
C3743 vdd.n2441 gnd 0.007657f
C3744 vdd.n2442 gnd 0.782467f
C3745 vdd.n2443 gnd 0.007657f
C3746 vdd.n2444 gnd 0.007657f
C3747 vdd.n2445 gnd 0.007657f
C3748 vdd.n2446 gnd 0.007657f
C3749 vdd.n2447 gnd 0.007657f
C3750 vdd.n2448 gnd 0.007657f
C3751 vdd.n2449 gnd 0.007657f
C3752 vdd.n2450 gnd 0.609864f
C3753 vdd.n2451 gnd 0.007657f
C3754 vdd.n2452 gnd 0.007657f
C3755 vdd.n2453 gnd 0.007657f
C3756 vdd.n2454 gnd 0.007657f
C3757 vdd.n2455 gnd 0.007657f
C3758 vdd.n2456 gnd 0.007657f
C3759 vdd.n2457 gnd 0.489042f
C3760 vdd.n2458 gnd 0.007657f
C3761 vdd.n2459 gnd 0.007657f
C3762 vdd.n2460 gnd 0.007657f
C3763 vdd.n2461 gnd 0.017895f
C3764 vdd.n2462 gnd 0.017235f
C3765 vdd.n2463 gnd 0.007657f
C3766 vdd.n2464 gnd 0.007657f
C3767 vdd.n2465 gnd 0.005911f
C3768 vdd.n2466 gnd 0.007657f
C3769 vdd.n2467 gnd 0.007657f
C3770 vdd.n2468 gnd 0.005574f
C3771 vdd.n2469 gnd 0.007657f
C3772 vdd.n2470 gnd 0.007657f
C3773 vdd.n2471 gnd 0.007657f
C3774 vdd.n2472 gnd 0.007657f
C3775 vdd.n2473 gnd 0.007657f
C3776 vdd.n2474 gnd 0.007657f
C3777 vdd.n2475 gnd 0.007657f
C3778 vdd.n2476 gnd 0.007657f
C3779 vdd.n2477 gnd 0.007657f
C3780 vdd.n2478 gnd 0.007657f
C3781 vdd.n2479 gnd 0.007657f
C3782 vdd.n2480 gnd 0.007657f
C3783 vdd.n2481 gnd 0.007657f
C3784 vdd.n2482 gnd 0.007657f
C3785 vdd.n2483 gnd 0.007657f
C3786 vdd.n2484 gnd 0.007657f
C3787 vdd.n2485 gnd 0.007657f
C3788 vdd.n2486 gnd 0.007657f
C3789 vdd.n2487 gnd 0.007657f
C3790 vdd.n2488 gnd 0.007657f
C3791 vdd.n2489 gnd 0.007657f
C3792 vdd.n2490 gnd 0.007657f
C3793 vdd.n2491 gnd 0.007657f
C3794 vdd.n2492 gnd 0.007657f
C3795 vdd.n2493 gnd 0.007657f
C3796 vdd.n2494 gnd 0.007657f
C3797 vdd.n2495 gnd 0.007657f
C3798 vdd.n2496 gnd 0.007657f
C3799 vdd.n2497 gnd 0.007657f
C3800 vdd.n2498 gnd 0.007657f
C3801 vdd.n2499 gnd 0.007657f
C3802 vdd.n2500 gnd 0.007657f
C3803 vdd.n2501 gnd 0.007657f
C3804 vdd.n2502 gnd 0.007657f
C3805 vdd.n2503 gnd 0.007657f
C3806 vdd.n2504 gnd 0.007657f
C3807 vdd.n2505 gnd 0.007657f
C3808 vdd.n2506 gnd 0.007657f
C3809 vdd.n2507 gnd 0.007657f
C3810 vdd.n2508 gnd 0.007657f
C3811 vdd.n2509 gnd 0.007657f
C3812 vdd.n2510 gnd 0.007657f
C3813 vdd.n2511 gnd 0.007657f
C3814 vdd.n2512 gnd 0.007657f
C3815 vdd.n2513 gnd 0.007657f
C3816 vdd.n2514 gnd 0.007657f
C3817 vdd.n2515 gnd 0.007657f
C3818 vdd.n2516 gnd 0.007657f
C3819 vdd.n2517 gnd 0.007657f
C3820 vdd.n2518 gnd 0.007657f
C3821 vdd.n2519 gnd 0.007657f
C3822 vdd.n2520 gnd 0.007657f
C3823 vdd.n2521 gnd 0.007657f
C3824 vdd.n2522 gnd 0.007657f
C3825 vdd.n2523 gnd 0.007657f
C3826 vdd.n2524 gnd 0.007657f
C3827 vdd.n2525 gnd 0.007657f
C3828 vdd.n2526 gnd 0.007657f
C3829 vdd.n2527 gnd 0.007657f
C3830 vdd.n2528 gnd 0.007657f
C3831 vdd.n2529 gnd 0.018168f
C3832 vdd.n2530 gnd 0.016963f
C3833 vdd.n2531 gnd 0.016963f
C3834 vdd.n2532 gnd 0.95507f
C3835 vdd.n2533 gnd 0.016963f
C3836 vdd.n2534 gnd 0.018168f
C3837 vdd.n2535 gnd 0.017235f
C3838 vdd.n2536 gnd 0.007657f
C3839 vdd.n2537 gnd 0.007657f
C3840 vdd.n2538 gnd 0.007657f
C3841 vdd.n2539 gnd 0.005911f
C3842 vdd.n2540 gnd 0.010943f
C3843 vdd.n2541 gnd 0.005574f
C3844 vdd.n2542 gnd 0.007657f
C3845 vdd.n2543 gnd 0.007657f
C3846 vdd.n2544 gnd 0.007657f
C3847 vdd.n2545 gnd 0.007657f
C3848 vdd.n2546 gnd 0.007657f
C3849 vdd.n2547 gnd 0.007657f
C3850 vdd.n2548 gnd 0.007657f
C3851 vdd.n2549 gnd 0.007657f
C3852 vdd.n2550 gnd 0.007657f
C3853 vdd.n2551 gnd 0.007657f
C3854 vdd.n2552 gnd 0.007657f
C3855 vdd.n2553 gnd 0.007657f
C3856 vdd.n2554 gnd 0.007657f
C3857 vdd.n2555 gnd 0.007657f
C3858 vdd.n2556 gnd 0.007657f
C3859 vdd.n2557 gnd 0.007657f
C3860 vdd.n2558 gnd 0.007657f
C3861 vdd.n2559 gnd 0.007657f
C3862 vdd.n2560 gnd 0.007657f
C3863 vdd.n2561 gnd 0.007657f
C3864 vdd.n2562 gnd 0.007657f
C3865 vdd.n2563 gnd 0.007657f
C3866 vdd.n2564 gnd 0.007657f
C3867 vdd.n2565 gnd 0.007657f
C3868 vdd.n2566 gnd 0.007657f
C3869 vdd.n2567 gnd 0.007657f
C3870 vdd.n2568 gnd 0.007657f
C3871 vdd.n2569 gnd 0.007657f
C3872 vdd.n2570 gnd 0.007657f
C3873 vdd.n2571 gnd 0.007657f
C3874 vdd.n2572 gnd 0.007657f
C3875 vdd.n2573 gnd 0.007657f
C3876 vdd.n2574 gnd 0.007657f
C3877 vdd.n2575 gnd 0.007657f
C3878 vdd.n2576 gnd 0.007657f
C3879 vdd.n2577 gnd 0.007657f
C3880 vdd.n2578 gnd 0.007657f
C3881 vdd.n2579 gnd 0.007657f
C3882 vdd.n2580 gnd 0.007657f
C3883 vdd.n2581 gnd 0.007657f
C3884 vdd.n2582 gnd 0.007657f
C3885 vdd.n2583 gnd 0.007657f
C3886 vdd.n2584 gnd 0.007657f
C3887 vdd.n2585 gnd 0.007657f
C3888 vdd.n2586 gnd 0.007657f
C3889 vdd.n2587 gnd 0.007657f
C3890 vdd.n2588 gnd 0.007657f
C3891 vdd.n2589 gnd 0.007657f
C3892 vdd.n2590 gnd 0.007657f
C3893 vdd.n2591 gnd 0.007657f
C3894 vdd.n2592 gnd 0.007657f
C3895 vdd.n2593 gnd 0.007657f
C3896 vdd.n2594 gnd 0.007657f
C3897 vdd.n2595 gnd 0.007657f
C3898 vdd.n2596 gnd 0.007657f
C3899 vdd.n2597 gnd 0.007657f
C3900 vdd.n2598 gnd 0.007657f
C3901 vdd.n2599 gnd 0.007657f
C3902 vdd.n2600 gnd 0.007657f
C3903 vdd.n2601 gnd 0.007657f
C3904 vdd.n2602 gnd 0.018168f
C3905 vdd.n2603 gnd 0.018168f
C3906 vdd.n2604 gnd 0.95507f
C3907 vdd.t142 gnd 3.39452f
C3908 vdd.t129 gnd 3.39452f
C3909 vdd.n2637 gnd 0.018168f
C3910 vdd.n2638 gnd 0.007657f
C3911 vdd.t214 gnd 0.309402f
C3912 vdd.t215 gnd 0.316711f
C3913 vdd.t212 gnd 0.201989f
C3914 vdd.n2639 gnd 0.109164f
C3915 vdd.n2640 gnd 0.061921f
C3916 vdd.n2641 gnd 0.007657f
C3917 vdd.t228 gnd 0.309402f
C3918 vdd.t229 gnd 0.316711f
C3919 vdd.t227 gnd 0.201989f
C3920 vdd.n2642 gnd 0.109164f
C3921 vdd.n2643 gnd 0.061921f
C3922 vdd.n2644 gnd 0.010943f
C3923 vdd.n2645 gnd 0.007657f
C3924 vdd.n2646 gnd 0.007657f
C3925 vdd.n2647 gnd 0.007657f
C3926 vdd.n2648 gnd 0.007657f
C3927 vdd.n2649 gnd 0.007657f
C3928 vdd.n2650 gnd 0.007657f
C3929 vdd.n2651 gnd 0.007657f
C3930 vdd.n2652 gnd 0.007657f
C3931 vdd.n2653 gnd 0.007657f
C3932 vdd.n2654 gnd 0.007657f
C3933 vdd.n2655 gnd 0.007657f
C3934 vdd.n2656 gnd 0.007657f
C3935 vdd.n2657 gnd 0.007657f
C3936 vdd.n2658 gnd 0.007657f
C3937 vdd.n2659 gnd 0.007657f
C3938 vdd.n2660 gnd 0.007657f
C3939 vdd.n2661 gnd 0.007657f
C3940 vdd.n2662 gnd 0.007657f
C3941 vdd.n2663 gnd 0.007657f
C3942 vdd.n2664 gnd 0.007657f
C3943 vdd.n2665 gnd 0.007657f
C3944 vdd.n2666 gnd 0.007657f
C3945 vdd.n2667 gnd 0.007657f
C3946 vdd.n2668 gnd 0.007657f
C3947 vdd.n2669 gnd 0.007657f
C3948 vdd.n2670 gnd 0.007657f
C3949 vdd.n2671 gnd 0.007657f
C3950 vdd.n2672 gnd 0.007657f
C3951 vdd.n2673 gnd 0.007657f
C3952 vdd.n2674 gnd 0.007657f
C3953 vdd.n2675 gnd 0.007657f
C3954 vdd.n2676 gnd 0.007657f
C3955 vdd.n2677 gnd 0.007657f
C3956 vdd.n2678 gnd 0.007657f
C3957 vdd.n2679 gnd 0.007657f
C3958 vdd.n2680 gnd 0.007657f
C3959 vdd.n2681 gnd 0.007657f
C3960 vdd.n2682 gnd 0.007657f
C3961 vdd.n2683 gnd 0.007657f
C3962 vdd.n2684 gnd 0.007657f
C3963 vdd.n2685 gnd 0.007657f
C3964 vdd.n2686 gnd 0.007657f
C3965 vdd.n2687 gnd 0.007657f
C3966 vdd.n2688 gnd 0.007657f
C3967 vdd.n2689 gnd 0.007657f
C3968 vdd.n2690 gnd 0.007657f
C3969 vdd.n2691 gnd 0.007657f
C3970 vdd.n2692 gnd 0.007657f
C3971 vdd.n2693 gnd 0.007657f
C3972 vdd.n2694 gnd 0.007657f
C3973 vdd.n2695 gnd 0.007657f
C3974 vdd.n2696 gnd 0.007657f
C3975 vdd.n2697 gnd 0.007657f
C3976 vdd.n2698 gnd 0.007657f
C3977 vdd.n2699 gnd 0.007657f
C3978 vdd.n2700 gnd 0.007657f
C3979 vdd.n2701 gnd 0.005574f
C3980 vdd.n2702 gnd 0.007657f
C3981 vdd.n2703 gnd 0.007657f
C3982 vdd.n2704 gnd 0.005911f
C3983 vdd.n2705 gnd 0.007657f
C3984 vdd.n2706 gnd 0.007657f
C3985 vdd.n2707 gnd 0.018168f
C3986 vdd.n2708 gnd 0.016963f
C3987 vdd.n2709 gnd 0.007657f
C3988 vdd.n2710 gnd 0.007657f
C3989 vdd.n2711 gnd 0.007657f
C3990 vdd.n2712 gnd 0.007657f
C3991 vdd.n2713 gnd 0.007657f
C3992 vdd.n2714 gnd 0.007657f
C3993 vdd.n2715 gnd 0.007657f
C3994 vdd.n2716 gnd 0.007657f
C3995 vdd.n2717 gnd 0.007657f
C3996 vdd.n2718 gnd 0.007657f
C3997 vdd.n2719 gnd 0.007657f
C3998 vdd.n2720 gnd 0.007657f
C3999 vdd.n2721 gnd 0.007657f
C4000 vdd.n2722 gnd 0.007657f
C4001 vdd.n2723 gnd 0.007657f
C4002 vdd.n2724 gnd 0.007657f
C4003 vdd.n2725 gnd 0.007657f
C4004 vdd.n2726 gnd 0.007657f
C4005 vdd.n2727 gnd 0.007657f
C4006 vdd.n2728 gnd 0.007657f
C4007 vdd.n2729 gnd 0.007657f
C4008 vdd.n2730 gnd 0.007657f
C4009 vdd.n2731 gnd 0.007657f
C4010 vdd.n2732 gnd 0.007657f
C4011 vdd.n2733 gnd 0.007657f
C4012 vdd.n2734 gnd 0.007657f
C4013 vdd.n2735 gnd 0.007657f
C4014 vdd.n2736 gnd 0.007657f
C4015 vdd.n2737 gnd 0.007657f
C4016 vdd.n2738 gnd 0.007657f
C4017 vdd.n2739 gnd 0.007657f
C4018 vdd.n2740 gnd 0.007657f
C4019 vdd.n2741 gnd 0.007657f
C4020 vdd.n2742 gnd 0.007657f
C4021 vdd.n2743 gnd 0.007657f
C4022 vdd.n2744 gnd 0.007657f
C4023 vdd.n2745 gnd 0.007657f
C4024 vdd.n2746 gnd 0.007657f
C4025 vdd.n2747 gnd 0.007657f
C4026 vdd.n2748 gnd 0.007657f
C4027 vdd.n2749 gnd 0.007657f
C4028 vdd.n2750 gnd 0.007657f
C4029 vdd.n2751 gnd 0.007657f
C4030 vdd.n2752 gnd 0.007657f
C4031 vdd.n2753 gnd 0.007657f
C4032 vdd.n2754 gnd 0.007657f
C4033 vdd.n2755 gnd 0.007657f
C4034 vdd.n2756 gnd 0.007657f
C4035 vdd.n2757 gnd 0.007657f
C4036 vdd.n2758 gnd 0.007657f
C4037 vdd.n2759 gnd 0.007657f
C4038 vdd.n2760 gnd 0.247398f
C4039 vdd.n2761 gnd 0.007657f
C4040 vdd.n2762 gnd 0.007657f
C4041 vdd.n2763 gnd 0.007657f
C4042 vdd.n2764 gnd 0.007657f
C4043 vdd.n2765 gnd 0.007657f
C4044 vdd.n2766 gnd 0.007657f
C4045 vdd.n2767 gnd 0.007657f
C4046 vdd.n2768 gnd 0.007657f
C4047 vdd.n2769 gnd 0.007657f
C4048 vdd.n2770 gnd 0.007657f
C4049 vdd.n2771 gnd 0.007657f
C4050 vdd.n2772 gnd 0.007657f
C4051 vdd.n2773 gnd 0.007657f
C4052 vdd.n2774 gnd 0.007657f
C4053 vdd.n2775 gnd 0.007657f
C4054 vdd.n2776 gnd 0.007657f
C4055 vdd.n2777 gnd 0.007657f
C4056 vdd.n2778 gnd 0.007657f
C4057 vdd.n2779 gnd 0.007657f
C4058 vdd.n2780 gnd 0.007657f
C4059 vdd.n2781 gnd 0.466028f
C4060 vdd.n2782 gnd 0.007657f
C4061 vdd.n2783 gnd 0.007657f
C4062 vdd.n2784 gnd 0.007657f
C4063 vdd.n2785 gnd 0.007657f
C4064 vdd.n2786 gnd 0.007657f
C4065 vdd.n2787 gnd 0.016963f
C4066 vdd.n2788 gnd 0.018168f
C4067 vdd.n2789 gnd 0.018168f
C4068 vdd.n2790 gnd 0.007657f
C4069 vdd.n2791 gnd 0.007657f
C4070 vdd.n2792 gnd 0.007657f
C4071 vdd.n2793 gnd 0.005911f
C4072 vdd.n2794 gnd 0.010943f
C4073 vdd.n2795 gnd 0.005574f
C4074 vdd.n2796 gnd 0.007657f
C4075 vdd.n2797 gnd 0.007657f
C4076 vdd.n2798 gnd 0.007657f
C4077 vdd.n2799 gnd 0.007657f
C4078 vdd.n2800 gnd 0.007657f
C4079 vdd.n2801 gnd 0.007657f
C4080 vdd.n2802 gnd 0.007657f
C4081 vdd.n2803 gnd 0.007657f
C4082 vdd.n2804 gnd 0.007657f
C4083 vdd.n2805 gnd 0.007657f
C4084 vdd.n2806 gnd 0.007657f
C4085 vdd.n2807 gnd 0.007657f
C4086 vdd.n2808 gnd 0.007657f
C4087 vdd.n2809 gnd 0.007657f
C4088 vdd.n2810 gnd 0.007657f
C4089 vdd.n2811 gnd 0.007657f
C4090 vdd.n2812 gnd 0.007657f
C4091 vdd.n2813 gnd 0.007657f
C4092 vdd.n2814 gnd 0.007657f
C4093 vdd.n2815 gnd 0.007657f
C4094 vdd.n2816 gnd 0.007657f
C4095 vdd.n2817 gnd 0.007657f
C4096 vdd.n2818 gnd 0.007657f
C4097 vdd.n2819 gnd 0.007657f
C4098 vdd.n2820 gnd 0.007657f
C4099 vdd.n2821 gnd 0.007657f
C4100 vdd.n2822 gnd 0.007657f
C4101 vdd.n2823 gnd 0.007657f
C4102 vdd.n2824 gnd 0.007657f
C4103 vdd.n2825 gnd 0.007657f
C4104 vdd.n2826 gnd 0.007657f
C4105 vdd.n2827 gnd 0.007657f
C4106 vdd.n2828 gnd 0.007657f
C4107 vdd.n2829 gnd 0.007657f
C4108 vdd.n2830 gnd 0.007657f
C4109 vdd.n2831 gnd 0.007657f
C4110 vdd.n2832 gnd 0.007657f
C4111 vdd.n2833 gnd 0.007657f
C4112 vdd.n2834 gnd 0.007657f
C4113 vdd.n2835 gnd 0.007657f
C4114 vdd.n2836 gnd 0.007657f
C4115 vdd.n2837 gnd 0.007657f
C4116 vdd.n2838 gnd 0.007657f
C4117 vdd.n2839 gnd 0.007657f
C4118 vdd.n2840 gnd 0.007657f
C4119 vdd.n2841 gnd 0.007657f
C4120 vdd.n2842 gnd 0.007657f
C4121 vdd.n2843 gnd 0.007657f
C4122 vdd.n2844 gnd 0.007657f
C4123 vdd.n2845 gnd 0.007657f
C4124 vdd.n2846 gnd 0.007657f
C4125 vdd.n2847 gnd 0.007657f
C4126 vdd.n2848 gnd 0.007657f
C4127 vdd.n2849 gnd 0.007657f
C4128 vdd.n2850 gnd 0.007657f
C4129 vdd.n2851 gnd 0.007657f
C4130 vdd.n2852 gnd 0.007657f
C4131 vdd.n2853 gnd 0.007657f
C4132 vdd.n2854 gnd 0.007657f
C4133 vdd.n2855 gnd 0.007657f
C4134 vdd.n2857 gnd 0.95507f
C4135 vdd.n2859 gnd 0.007657f
C4136 vdd.n2860 gnd 0.007657f
C4137 vdd.n2861 gnd 0.018168f
C4138 vdd.n2862 gnd 0.016963f
C4139 vdd.n2863 gnd 0.016963f
C4140 vdd.n2864 gnd 0.95507f
C4141 vdd.n2865 gnd 0.016963f
C4142 vdd.n2866 gnd 0.016963f
C4143 vdd.n2867 gnd 0.007657f
C4144 vdd.n2868 gnd 0.007657f
C4145 vdd.n2869 gnd 0.007657f
C4146 vdd.n2870 gnd 0.489042f
C4147 vdd.n2871 gnd 0.007657f
C4148 vdd.n2872 gnd 0.007657f
C4149 vdd.n2873 gnd 0.007657f
C4150 vdd.n2874 gnd 0.007657f
C4151 vdd.n2875 gnd 0.007657f
C4152 vdd.n2876 gnd 0.609864f
C4153 vdd.n2877 gnd 0.007657f
C4154 vdd.n2878 gnd 0.007657f
C4155 vdd.n2879 gnd 0.007657f
C4156 vdd.n2880 gnd 0.007657f
C4157 vdd.n2881 gnd 0.007657f
C4158 vdd.n2882 gnd 0.782467f
C4159 vdd.n2883 gnd 0.007657f
C4160 vdd.n2884 gnd 0.007657f
C4161 vdd.n2885 gnd 0.007657f
C4162 vdd.n2886 gnd 0.007657f
C4163 vdd.n2887 gnd 0.007657f
C4164 vdd.n2888 gnd 0.431507f
C4165 vdd.n2889 gnd 0.007657f
C4166 vdd.n2890 gnd 0.007657f
C4167 vdd.n2891 gnd 0.007657f
C4168 vdd.n2892 gnd 0.007657f
C4169 vdd.n2893 gnd 0.007657f
C4170 vdd.n2894 gnd 0.247398f
C4171 vdd.n2895 gnd 0.007657f
C4172 vdd.n2896 gnd 0.007657f
C4173 vdd.n2897 gnd 0.007657f
C4174 vdd.n2898 gnd 0.007657f
C4175 vdd.n2899 gnd 0.007657f
C4176 vdd.n2900 gnd 0.448768f
C4177 vdd.n2901 gnd 0.007657f
C4178 vdd.n2902 gnd 0.007657f
C4179 vdd.n2903 gnd 0.007657f
C4180 vdd.n2904 gnd 0.007657f
C4181 vdd.n2905 gnd 0.007657f
C4182 vdd.n2906 gnd 0.621371f
C4183 vdd.n2907 gnd 0.007657f
C4184 vdd.n2908 gnd 0.007657f
C4185 vdd.n2909 gnd 0.007657f
C4186 vdd.n2910 gnd 0.007657f
C4187 vdd.n2911 gnd 0.007657f
C4188 vdd.n2912 gnd 0.696165f
C4189 vdd.n2913 gnd 0.007657f
C4190 vdd.n2914 gnd 0.007657f
C4191 vdd.n2915 gnd 0.007657f
C4192 vdd.n2916 gnd 0.007657f
C4193 vdd.n2917 gnd 0.007657f
C4194 vdd.n2918 gnd 0.523562f
C4195 vdd.n2919 gnd 0.007657f
C4196 vdd.n2920 gnd 0.007657f
C4197 vdd.n2921 gnd 0.007657f
C4198 vdd.t182 gnd 0.316711f
C4199 vdd.t180 gnd 0.201989f
C4200 vdd.t183 gnd 0.316711f
C4201 vdd.n2922 gnd 0.178004f
C4202 vdd.n2923 gnd 0.02218f
C4203 vdd.n2924 gnd 0.004729f
C4204 vdd.n2925 gnd 0.007657f
C4205 vdd.n2926 gnd 0.431507f
C4206 vdd.n2927 gnd 0.007657f
C4207 vdd.n2928 gnd 0.007657f
C4208 vdd.n2929 gnd 0.007657f
C4209 vdd.n2930 gnd 0.007657f
C4210 vdd.n2931 gnd 0.007657f
C4211 vdd.n2932 gnd 0.782467f
C4212 vdd.n2933 gnd 0.007657f
C4213 vdd.n2934 gnd 0.007657f
C4214 vdd.n2935 gnd 0.007657f
C4215 vdd.n2936 gnd 0.007657f
C4216 vdd.n2937 gnd 0.007657f
C4217 vdd.n2938 gnd 0.007657f
C4218 vdd.n2940 gnd 0.007657f
C4219 vdd.n2941 gnd 0.007657f
C4220 vdd.n2943 gnd 0.007657f
C4221 vdd.n2944 gnd 0.007657f
C4222 vdd.n2947 gnd 0.007657f
C4223 vdd.n2948 gnd 0.007657f
C4224 vdd.n2949 gnd 0.007657f
C4225 vdd.n2950 gnd 0.007657f
C4226 vdd.n2952 gnd 0.007657f
C4227 vdd.n2953 gnd 0.007657f
C4228 vdd.n2954 gnd 0.007657f
C4229 vdd.n2955 gnd 0.007657f
C4230 vdd.n2956 gnd 0.007657f
C4231 vdd.n2957 gnd 0.007657f
C4232 vdd.n2959 gnd 0.007657f
C4233 vdd.n2960 gnd 0.007657f
C4234 vdd.n2961 gnd 0.007657f
C4235 vdd.n2962 gnd 0.007657f
C4236 vdd.n2963 gnd 0.007657f
C4237 vdd.n2964 gnd 0.007657f
C4238 vdd.n2966 gnd 0.007657f
C4239 vdd.n2967 gnd 0.007657f
C4240 vdd.n2968 gnd 0.007657f
C4241 vdd.n2969 gnd 0.007657f
C4242 vdd.n2970 gnd 0.007657f
C4243 vdd.n2971 gnd 0.007657f
C4244 vdd.n2973 gnd 0.007657f
C4245 vdd.n2974 gnd 0.018168f
C4246 vdd.n2975 gnd 0.018168f
C4247 vdd.n2976 gnd 0.016963f
C4248 vdd.n2977 gnd 0.007657f
C4249 vdd.n2978 gnd 0.007657f
C4250 vdd.n2979 gnd 0.007657f
C4251 vdd.n2980 gnd 0.007657f
C4252 vdd.n2981 gnd 0.007657f
C4253 vdd.n2982 gnd 0.007657f
C4254 vdd.n2983 gnd 0.782467f
C4255 vdd.n2984 gnd 0.007657f
C4256 vdd.n2985 gnd 0.007657f
C4257 vdd.n2986 gnd 0.007657f
C4258 vdd.n2987 gnd 0.007657f
C4259 vdd.n2988 gnd 0.007657f
C4260 vdd.n2989 gnd 0.489042f
C4261 vdd.n2990 gnd 0.007657f
C4262 vdd.n2991 gnd 0.007657f
C4263 vdd.n2992 gnd 0.007657f
C4264 vdd.n2993 gnd 0.017895f
C4265 vdd.n2994 gnd 0.017235f
C4266 vdd.n2995 gnd 0.018168f
C4267 vdd.n2997 gnd 0.007657f
C4268 vdd.n2998 gnd 0.007657f
C4269 vdd.n2999 gnd 0.005911f
C4270 vdd.n3000 gnd 0.010943f
C4271 vdd.n3001 gnd 0.005574f
C4272 vdd.n3002 gnd 0.007657f
C4273 vdd.n3003 gnd 0.007657f
C4274 vdd.n3005 gnd 0.007657f
C4275 vdd.n3006 gnd 0.007657f
C4276 vdd.n3007 gnd 0.007657f
C4277 vdd.n3008 gnd 0.007657f
C4278 vdd.n3009 gnd 0.007657f
C4279 vdd.n3010 gnd 0.007657f
C4280 vdd.n3012 gnd 0.007657f
C4281 vdd.n3013 gnd 0.007657f
C4282 vdd.n3014 gnd 0.007657f
C4283 vdd.n3015 gnd 0.007657f
C4284 vdd.n3016 gnd 0.007657f
C4285 vdd.n3017 gnd 0.007657f
C4286 vdd.n3019 gnd 0.007657f
C4287 vdd.n3020 gnd 0.007657f
C4288 vdd.n3021 gnd 0.007657f
C4289 vdd.n3022 gnd 0.007657f
C4290 vdd.n3023 gnd 0.007657f
C4291 vdd.n3024 gnd 0.007657f
C4292 vdd.n3026 gnd 0.007657f
C4293 vdd.n3027 gnd 0.007657f
C4294 vdd.n3028 gnd 0.007657f
C4295 vdd.n3030 gnd 0.007657f
C4296 vdd.n3031 gnd 0.007657f
C4297 vdd.n3032 gnd 0.007657f
C4298 vdd.n3033 gnd 0.007657f
C4299 vdd.n3034 gnd 0.007657f
C4300 vdd.n3035 gnd 0.007657f
C4301 vdd.n3037 gnd 0.007657f
C4302 vdd.n3038 gnd 0.007657f
C4303 vdd.n3039 gnd 0.007657f
C4304 vdd.n3040 gnd 0.007657f
C4305 vdd.n3041 gnd 0.007657f
C4306 vdd.n3042 gnd 0.007657f
C4307 vdd.n3044 gnd 0.007657f
C4308 vdd.n3045 gnd 0.007657f
C4309 vdd.n3046 gnd 0.007657f
C4310 vdd.n3047 gnd 0.007657f
C4311 vdd.n3048 gnd 0.007657f
C4312 vdd.n3049 gnd 0.007657f
C4313 vdd.n3051 gnd 0.007657f
C4314 vdd.n3052 gnd 0.007657f
C4315 vdd.n3054 gnd 0.007657f
C4316 vdd.n3055 gnd 0.007657f
C4317 vdd.n3056 gnd 0.018168f
C4318 vdd.n3057 gnd 0.016963f
C4319 vdd.n3058 gnd 0.016963f
C4320 vdd.n3059 gnd 1.12767f
C4321 vdd.n3060 gnd 0.016963f
C4322 vdd.n3061 gnd 0.018168f
C4323 vdd.n3062 gnd 0.017235f
C4324 vdd.n3063 gnd 0.007657f
C4325 vdd.n3064 gnd 0.005911f
C4326 vdd.n3065 gnd 0.007657f
C4327 vdd.n3067 gnd 0.007657f
C4328 vdd.n3068 gnd 0.007657f
C4329 vdd.n3069 gnd 0.007657f
C4330 vdd.n3070 gnd 0.007657f
C4331 vdd.n3071 gnd 0.007657f
C4332 vdd.n3072 gnd 0.007657f
C4333 vdd.n3074 gnd 0.007657f
C4334 vdd.n3075 gnd 0.007657f
C4335 vdd.n3076 gnd 0.007657f
C4336 vdd.n3077 gnd 0.007657f
C4337 vdd.n3078 gnd 0.007657f
C4338 vdd.n3079 gnd 0.007657f
C4339 vdd.n3081 gnd 0.007657f
C4340 vdd.n3082 gnd 0.007657f
C4341 vdd.n3083 gnd 0.007657f
C4342 vdd.n3084 gnd 0.007657f
C4343 vdd.n3085 gnd 0.007657f
C4344 vdd.n3086 gnd 0.007657f
C4345 vdd.n3088 gnd 0.007657f
C4346 vdd.n3089 gnd 0.007657f
C4347 vdd.n3091 gnd 0.007657f
C4348 vdd.n3092 gnd 0.018399f
C4349 vdd.n3093 gnd 0.681454f
C4350 vdd.n3095 gnd 0.004758f
C4351 vdd.n3096 gnd 0.009063f
C4352 vdd.n3097 gnd 0.01126f
C4353 vdd.n3098 gnd 0.01126f
C4354 vdd.n3099 gnd 0.009063f
C4355 vdd.n3100 gnd 0.009063f
C4356 vdd.n3101 gnd 0.01126f
C4357 vdd.n3102 gnd 0.01126f
C4358 vdd.n3103 gnd 0.009063f
C4359 vdd.n3104 gnd 0.009063f
C4360 vdd.n3105 gnd 0.01126f
C4361 vdd.n3106 gnd 0.01126f
C4362 vdd.n3107 gnd 0.009063f
C4363 vdd.n3108 gnd 0.009063f
C4364 vdd.n3109 gnd 0.01126f
C4365 vdd.n3110 gnd 0.01126f
C4366 vdd.n3111 gnd 0.009063f
C4367 vdd.n3112 gnd 0.009063f
C4368 vdd.n3113 gnd 0.01126f
C4369 vdd.n3114 gnd 0.01126f
C4370 vdd.n3115 gnd 0.009063f
C4371 vdd.n3116 gnd 0.009063f
C4372 vdd.n3117 gnd 0.01126f
C4373 vdd.n3118 gnd 0.01126f
C4374 vdd.n3119 gnd 0.009063f
C4375 vdd.n3120 gnd 0.009063f
C4376 vdd.n3121 gnd 0.01126f
C4377 vdd.n3122 gnd 0.01126f
C4378 vdd.n3123 gnd 0.009063f
C4379 vdd.n3124 gnd 0.009063f
C4380 vdd.n3125 gnd 0.01126f
C4381 vdd.n3126 gnd 0.01126f
C4382 vdd.n3127 gnd 0.009063f
C4383 vdd.n3128 gnd 0.009063f
C4384 vdd.n3129 gnd 0.01126f
C4385 vdd.n3130 gnd 0.01126f
C4386 vdd.n3131 gnd 0.009063f
C4387 vdd.n3132 gnd 0.01126f
C4388 vdd.n3133 gnd 0.01126f
C4389 vdd.n3134 gnd 0.009063f
C4390 vdd.n3135 gnd 0.01126f
C4391 vdd.n3136 gnd 0.01126f
C4392 vdd.n3137 gnd 0.01126f
C4393 vdd.n3138 gnd 0.018488f
C4394 vdd.n3139 gnd 0.01126f
C4395 vdd.n3140 gnd 0.01126f
C4396 vdd.n3141 gnd 0.006163f
C4397 vdd.n3142 gnd 0.009063f
C4398 vdd.n3143 gnd 0.01126f
C4399 vdd.n3144 gnd 0.01126f
C4400 vdd.n3145 gnd 0.009063f
C4401 vdd.n3146 gnd 0.009063f
C4402 vdd.n3147 gnd 0.01126f
C4403 vdd.n3148 gnd 0.01126f
C4404 vdd.n3149 gnd 0.009063f
C4405 vdd.n3150 gnd 0.009063f
C4406 vdd.n3151 gnd 0.01126f
C4407 vdd.n3152 gnd 0.01126f
C4408 vdd.n3153 gnd 0.009063f
C4409 vdd.n3154 gnd 0.009063f
C4410 vdd.n3155 gnd 0.01126f
C4411 vdd.n3156 gnd 0.01126f
C4412 vdd.n3157 gnd 0.009063f
C4413 vdd.n3158 gnd 0.009063f
C4414 vdd.n3159 gnd 0.01126f
C4415 vdd.n3160 gnd 0.01126f
C4416 vdd.n3161 gnd 0.009063f
C4417 vdd.n3162 gnd 0.009063f
C4418 vdd.n3163 gnd 0.01126f
C4419 vdd.n3164 gnd 0.01126f
C4420 vdd.n3165 gnd 0.009063f
C4421 vdd.n3166 gnd 0.009063f
C4422 vdd.n3167 gnd 0.01126f
C4423 vdd.n3168 gnd 0.01126f
C4424 vdd.n3169 gnd 0.009063f
C4425 vdd.n3170 gnd 0.009063f
C4426 vdd.n3171 gnd 0.01126f
C4427 vdd.n3172 gnd 0.01126f
C4428 vdd.n3173 gnd 0.009063f
C4429 vdd.n3174 gnd 0.009063f
C4430 vdd.n3175 gnd 0.01126f
C4431 vdd.n3176 gnd 0.01126f
C4432 vdd.n3177 gnd 0.009063f
C4433 vdd.n3178 gnd 0.01126f
C4434 vdd.n3179 gnd 0.01126f
C4435 vdd.n3180 gnd 0.009063f
C4436 vdd.n3181 gnd 0.01126f
C4437 vdd.n3182 gnd 0.01126f
C4438 vdd.n3183 gnd 0.01126f
C4439 vdd.t174 gnd 0.138524f
C4440 vdd.t175 gnd 0.148044f
C4441 vdd.t173 gnd 0.18091f
C4442 vdd.n3184 gnd 0.231901f
C4443 vdd.n3185 gnd 0.194839f
C4444 vdd.n3186 gnd 0.018488f
C4445 vdd.n3187 gnd 0.01126f
C4446 vdd.n3188 gnd 0.01126f
C4447 vdd.n3189 gnd 0.007567f
C4448 vdd.n3190 gnd 0.009063f
C4449 vdd.n3191 gnd 0.01126f
C4450 vdd.n3192 gnd 0.01126f
C4451 vdd.n3193 gnd 0.009063f
C4452 vdd.n3194 gnd 0.009063f
C4453 vdd.n3195 gnd 0.01126f
C4454 vdd.n3196 gnd 0.01126f
C4455 vdd.n3197 gnd 0.009063f
C4456 vdd.n3198 gnd 0.009063f
C4457 vdd.n3199 gnd 0.01126f
C4458 vdd.n3200 gnd 0.01126f
C4459 vdd.n3201 gnd 0.009063f
C4460 vdd.n3202 gnd 0.009063f
C4461 vdd.n3203 gnd 0.01126f
C4462 vdd.n3204 gnd 0.01126f
C4463 vdd.n3205 gnd 0.009063f
C4464 vdd.n3206 gnd 0.009063f
C4465 vdd.n3207 gnd 0.01126f
C4466 vdd.n3208 gnd 0.01126f
C4467 vdd.n3209 gnd 0.009063f
C4468 vdd.n3210 gnd 0.009063f
C4469 vdd.n3211 gnd 0.01126f
C4470 vdd.n3212 gnd 0.01126f
C4471 vdd.n3213 gnd 0.009063f
C4472 vdd.n3214 gnd 0.009063f
C4473 vdd.n3216 gnd 0.681454f
C4474 vdd.n3218 gnd 0.009063f
C4475 vdd.n3219 gnd 0.009063f
C4476 vdd.n3220 gnd 0.007522f
C4477 vdd.n3221 gnd 0.027822f
C4478 vdd.n3223 gnd 8.31946f
C4479 vdd.n3224 gnd 0.027822f
C4480 vdd.n3225 gnd 0.004305f
C4481 vdd.n3226 gnd 0.027822f
C4482 vdd.n3227 gnd 0.027238f
C4483 vdd.n3228 gnd 0.01126f
C4484 vdd.n3229 gnd 0.009063f
C4485 vdd.n3230 gnd 0.01126f
C4486 vdd.n3231 gnd 0.696165f
C4487 vdd.n3232 gnd 0.01126f
C4488 vdd.n3233 gnd 0.009063f
C4489 vdd.n3234 gnd 0.01126f
C4490 vdd.n3235 gnd 0.01126f
C4491 vdd.n3236 gnd 0.01126f
C4492 vdd.n3237 gnd 0.009063f
C4493 vdd.n3238 gnd 0.01126f
C4494 vdd.n3239 gnd 1.15069f
C4495 vdd.n3240 gnd 0.01126f
C4496 vdd.n3241 gnd 0.009063f
C4497 vdd.n3242 gnd 0.01126f
C4498 vdd.n3243 gnd 0.01126f
C4499 vdd.n3244 gnd 0.01126f
C4500 vdd.n3245 gnd 0.009063f
C4501 vdd.n3246 gnd 0.01126f
C4502 vdd.n3247 gnd 0.742193f
C4503 vdd.n3248 gnd 0.78822f
C4504 vdd.n3249 gnd 0.01126f
C4505 vdd.n3250 gnd 0.009063f
C4506 vdd.n3251 gnd 0.01126f
C4507 vdd.n3252 gnd 0.01126f
C4508 vdd.n3253 gnd 0.01126f
C4509 vdd.n3254 gnd 0.009063f
C4510 vdd.n3255 gnd 0.01126f
C4511 vdd.n3256 gnd 0.95507f
C4512 vdd.n3257 gnd 0.01126f
C4513 vdd.n3258 gnd 0.009063f
C4514 vdd.n3259 gnd 0.01126f
C4515 vdd.n3260 gnd 0.01126f
C4516 vdd.n3261 gnd 0.01126f
C4517 vdd.n3262 gnd 0.009063f
C4518 vdd.n3263 gnd 0.01126f
C4519 vdd.t94 gnd 0.575343f
C4520 vdd.n3264 gnd 0.926302f
C4521 vdd.n3265 gnd 0.01126f
C4522 vdd.n3266 gnd 0.009063f
C4523 vdd.n3267 gnd 0.01126f
C4524 vdd.n3268 gnd 0.01126f
C4525 vdd.n3269 gnd 0.01126f
C4526 vdd.n3270 gnd 0.009063f
C4527 vdd.n3271 gnd 0.01126f
C4528 vdd.n3272 gnd 0.730686f
C4529 vdd.n3273 gnd 0.01126f
C4530 vdd.n3274 gnd 0.009063f
C4531 vdd.n3275 gnd 0.01126f
C4532 vdd.n3276 gnd 0.01126f
C4533 vdd.n3277 gnd 0.01126f
C4534 vdd.n3278 gnd 0.009063f
C4535 vdd.n3279 gnd 0.01126f
C4536 vdd.n3280 gnd 0.914796f
C4537 vdd.n3281 gnd 0.615617f
C4538 vdd.n3282 gnd 0.01126f
C4539 vdd.n3283 gnd 0.009063f
C4540 vdd.n3284 gnd 0.01126f
C4541 vdd.n3285 gnd 0.01126f
C4542 vdd.n3286 gnd 0.01126f
C4543 vdd.n3287 gnd 0.009063f
C4544 vdd.n3288 gnd 0.01126f
C4545 vdd.n3289 gnd 0.811234f
C4546 vdd.n3290 gnd 0.01126f
C4547 vdd.n3291 gnd 0.009063f
C4548 vdd.n3292 gnd 0.01126f
C4549 vdd.n3293 gnd 0.01126f
C4550 vdd.n3294 gnd 0.01126f
C4551 vdd.n3295 gnd 0.01126f
C4552 vdd.n3296 gnd 0.01126f
C4553 vdd.n3297 gnd 0.009063f
C4554 vdd.n3298 gnd 0.009063f
C4555 vdd.n3299 gnd 0.01126f
C4556 vdd.t67 gnd 0.575343f
C4557 vdd.n3300 gnd 0.95507f
C4558 vdd.n3301 gnd 0.01126f
C4559 vdd.n3302 gnd 0.009063f
C4560 vdd.n3303 gnd 0.01126f
C4561 vdd.n3304 gnd 0.01126f
C4562 vdd.n3305 gnd 0.01126f
C4563 vdd.n3306 gnd 0.009063f
C4564 vdd.n3307 gnd 0.01126f
C4565 vdd.n3308 gnd 0.903289f
C4566 vdd.n3309 gnd 0.01126f
C4567 vdd.n3310 gnd 0.01126f
C4568 vdd.n3311 gnd 0.009063f
C4569 vdd.n3312 gnd 0.009063f
C4570 vdd.n3313 gnd 0.01126f
C4571 vdd.n3314 gnd 0.01126f
C4572 vdd.n3315 gnd 0.01126f
C4573 vdd.n3316 gnd 0.009063f
C4574 vdd.n3317 gnd 0.01126f
C4575 vdd.n3318 gnd 0.009063f
C4576 vdd.n3319 gnd 0.009063f
C4577 vdd.n3320 gnd 0.01126f
C4578 vdd.n3321 gnd 0.01126f
C4579 vdd.n3322 gnd 0.01126f
C4580 vdd.n3323 gnd 0.009063f
C4581 vdd.n3324 gnd 0.01126f
C4582 vdd.n3325 gnd 0.009063f
C4583 vdd.n3326 gnd 0.009063f
C4584 vdd.n3327 gnd 0.01126f
C4585 vdd.n3328 gnd 0.01126f
C4586 vdd.n3329 gnd 0.01126f
C4587 vdd.n3330 gnd 0.009063f
C4588 vdd.n3331 gnd 0.95507f
C4589 vdd.n3332 gnd 0.01126f
C4590 vdd.n3333 gnd 0.009063f
C4591 vdd.n3334 gnd 0.009063f
C4592 vdd.n3335 gnd 0.01126f
C4593 vdd.n3336 gnd 0.01126f
C4594 vdd.n3337 gnd 0.01126f
C4595 vdd.n3338 gnd 0.009063f
C4596 vdd.n3339 gnd 0.01126f
C4597 vdd.n3340 gnd 0.009063f
C4598 vdd.n3341 gnd 0.009063f
C4599 vdd.n3342 gnd 0.01126f
C4600 vdd.n3343 gnd 0.01126f
C4601 vdd.n3344 gnd 0.01126f
C4602 vdd.n3345 gnd 0.009063f
C4603 vdd.n3346 gnd 0.01126f
C4604 vdd.n3347 gnd 0.009063f
C4605 vdd.n3348 gnd 0.007522f
C4606 vdd.n3349 gnd 0.027238f
C4607 vdd.n3350 gnd 0.027822f
C4608 vdd.n3351 gnd 0.004305f
C4609 vdd.n3352 gnd 0.027822f
C4610 vdd.n3354 gnd 2.72713f
C4611 vdd.n3355 gnd 1.69726f
C4612 vdd.n3356 gnd 0.027238f
C4613 vdd.n3357 gnd 0.007522f
C4614 vdd.n3358 gnd 0.009063f
C4615 vdd.n3359 gnd 0.009063f
C4616 vdd.n3360 gnd 0.01126f
C4617 vdd.n3361 gnd 1.15069f
C4618 vdd.n3362 gnd 1.15069f
C4619 vdd.n3363 gnd 1.05288f
C4620 vdd.n3364 gnd 0.01126f
C4621 vdd.n3365 gnd 0.009063f
C4622 vdd.n3366 gnd 0.009063f
C4623 vdd.n3367 gnd 0.009063f
C4624 vdd.n3368 gnd 0.01126f
C4625 vdd.n3369 gnd 0.857261f
C4626 vdd.t30 gnd 0.575343f
C4627 vdd.n3370 gnd 0.868768f
C4628 vdd.n3371 gnd 0.661645f
C4629 vdd.n3372 gnd 0.01126f
C4630 vdd.n3373 gnd 0.009063f
C4631 vdd.n3374 gnd 0.009063f
C4632 vdd.n3375 gnd 0.009063f
C4633 vdd.n3376 gnd 0.01126f
C4634 vdd.n3377 gnd 0.684658f
C4635 vdd.n3378 gnd 0.845754f
C4636 vdd.t36 gnd 0.575343f
C4637 vdd.n3379 gnd 0.880275f
C4638 vdd.n3380 gnd 0.01126f
C4639 vdd.n3381 gnd 0.009063f
C4640 vdd.n3382 gnd 0.009063f
C4641 vdd.n3383 gnd 0.009063f
C4642 vdd.n3384 gnd 0.01126f
C4643 vdd.n3385 gnd 0.95507f
C4644 vdd.t90 gnd 0.575343f
C4645 vdd.n3386 gnd 0.696165f
C4646 vdd.n3387 gnd 0.834248f
C4647 vdd.n3388 gnd 0.01126f
C4648 vdd.n3389 gnd 0.009063f
C4649 vdd.n3390 gnd 0.009063f
C4650 vdd.n3391 gnd 0.009063f
C4651 vdd.n3392 gnd 0.01126f
C4652 vdd.n3393 gnd 0.638631f
C4653 vdd.t0 gnd 0.575343f
C4654 vdd.n3394 gnd 0.95507f
C4655 vdd.t2 gnd 0.575343f
C4656 vdd.n3395 gnd 0.707672f
C4657 vdd.n3396 gnd 0.01126f
C4658 vdd.n3397 gnd 0.009063f
C4659 vdd.n3398 gnd 0.008654f
C4660 vdd.n3399 gnd 0.664139f
C4661 vdd.n3400 gnd 2.87926f
C4662 a_n1986_13878.n0 gnd 3.20192f
C4663 a_n1986_13878.n1 gnd 0.64915f
C4664 a_n1986_13878.n2 gnd 0.219304f
C4665 a_n1986_13878.n3 gnd 0.286909f
C4666 a_n1986_13878.n4 gnd 0.452885f
C4667 a_n1986_13878.n5 gnd 0.674778f
C4668 a_n1986_13878.n6 gnd 0.219304f
C4669 a_n1986_13878.n7 gnd 0.286909f
C4670 a_n1986_13878.n8 gnd 0.534226f
C4671 a_n1986_13878.n9 gnd 0.208083f
C4672 a_n1986_13878.n10 gnd 0.153257f
C4673 a_n1986_13878.n11 gnd 0.240872f
C4674 a_n1986_13878.n12 gnd 0.186046f
C4675 a_n1986_13878.n13 gnd 0.208083f
C4676 a_n1986_13878.n14 gnd 1.02197f
C4677 a_n1986_13878.n15 gnd 0.153257f
C4678 a_n1986_13878.n16 gnd 0.589052f
C4679 a_n1986_13878.n17 gnd 0.439018f
C4680 a_n1986_13878.n18 gnd 0.219304f
C4681 a_n1986_13878.n19 gnd 0.500138f
C4682 a_n1986_13878.n20 gnd 0.286909f
C4683 a_n1986_13878.n21 gnd 0.445312f
C4684 a_n1986_13878.n22 gnd 0.219304f
C4685 a_n1986_13878.n23 gnd 0.742922f
C4686 a_n1986_13878.n24 gnd 0.286909f
C4687 a_n1986_13878.n25 gnd 1.19721f
C4688 a_n1986_13878.n26 gnd 1.9455f
C4689 a_n1986_13878.n27 gnd 1.8055f
C4690 a_n1986_13878.n28 gnd 2.46475f
C4691 a_n1986_13878.n29 gnd 3.82161f
C4692 a_n1986_13878.n30 gnd 3.20861f
C4693 a_n1986_13878.n31 gnd 0.008491f
C4694 a_n1986_13878.n33 gnd 0.290112f
C4695 a_n1986_13878.n34 gnd 0.008491f
C4696 a_n1986_13878.n36 gnd 0.290112f
C4697 a_n1986_13878.n37 gnd 0.008491f
C4698 a_n1986_13878.n38 gnd 0.2897f
C4699 a_n1986_13878.n39 gnd 0.008491f
C4700 a_n1986_13878.n40 gnd 0.2897f
C4701 a_n1986_13878.n41 gnd 0.008491f
C4702 a_n1986_13878.n42 gnd 0.2897f
C4703 a_n1986_13878.n43 gnd 0.008491f
C4704 a_n1986_13878.n44 gnd 0.2897f
C4705 a_n1986_13878.n45 gnd 0.008491f
C4706 a_n1986_13878.n47 gnd 0.290112f
C4707 a_n1986_13878.n48 gnd 0.008491f
C4708 a_n1986_13878.n50 gnd 0.290112f
C4709 a_n1986_13878.t11 gnd 0.722451f
C4710 a_n1986_13878.t13 gnd 0.707549f
C4711 a_n1986_13878.t33 gnd 0.707549f
C4712 a_n1986_13878.t17 gnd 0.707549f
C4713 a_n1986_13878.n51 gnd 0.311083f
C4714 a_n1986_13878.t29 gnd 0.707549f
C4715 a_n1986_13878.t19 gnd 0.719248f
C4716 a_n1986_13878.t67 gnd 0.722451f
C4717 a_n1986_13878.t50 gnd 0.707549f
C4718 a_n1986_13878.t54 gnd 0.707549f
C4719 a_n1986_13878.t44 gnd 0.707549f
C4720 a_n1986_13878.n52 gnd 0.311083f
C4721 a_n1986_13878.t59 gnd 0.707549f
C4722 a_n1986_13878.t65 gnd 0.719248f
C4723 a_n1986_13878.t28 gnd 1.4243f
C4724 a_n1986_13878.t22 gnd 0.152112f
C4725 a_n1986_13878.t24 gnd 0.152112f
C4726 a_n1986_13878.n53 gnd 1.07147f
C4727 a_n1986_13878.t16 gnd 0.152112f
C4728 a_n1986_13878.t26 gnd 0.152112f
C4729 a_n1986_13878.n54 gnd 1.07147f
C4730 a_n1986_13878.t32 gnd 1.42146f
C4731 a_n1986_13878.t15 gnd 0.707549f
C4732 a_n1986_13878.n55 gnd 0.311083f
C4733 a_n1986_13878.t25 gnd 0.707549f
C4734 a_n1986_13878.t21 gnd 0.707549f
C4735 a_n1986_13878.t48 gnd 0.707549f
C4736 a_n1986_13878.n56 gnd 0.311083f
C4737 a_n1986_13878.t57 gnd 0.707549f
C4738 a_n1986_13878.t63 gnd 0.707549f
C4739 a_n1986_13878.t62 gnd 0.722451f
C4740 a_n1986_13878.n57 gnd 0.313741f
C4741 a_n1986_13878.t42 gnd 0.707549f
C4742 a_n1986_13878.n58 gnd 0.307133f
C4743 a_n1986_13878.n59 gnd 0.313742f
C4744 a_n1986_13878.t43 gnd 0.719248f
C4745 a_n1986_13878.t27 gnd 0.722451f
C4746 a_n1986_13878.n60 gnd 0.313741f
C4747 a_n1986_13878.t23 gnd 0.707549f
C4748 a_n1986_13878.n61 gnd 0.307133f
C4749 a_n1986_13878.n62 gnd 0.313742f
C4750 a_n1986_13878.t31 gnd 0.719248f
C4751 a_n1986_13878.n63 gnd 1.14966f
C4752 a_n1986_13878.t47 gnd 0.707549f
C4753 a_n1986_13878.n64 gnd 0.307133f
C4754 a_n1986_13878.t53 gnd 0.707549f
C4755 a_n1986_13878.n65 gnd 0.307133f
C4756 a_n1986_13878.t45 gnd 0.707549f
C4757 a_n1986_13878.n66 gnd 0.307133f
C4758 a_n1986_13878.t58 gnd 0.707549f
C4759 a_n1986_13878.n67 gnd 0.307133f
C4760 a_n1986_13878.t49 gnd 0.707549f
C4761 a_n1986_13878.n68 gnd 0.301556f
C4762 a_n1986_13878.t40 gnd 0.707549f
C4763 a_n1986_13878.n69 gnd 0.311083f
C4764 a_n1986_13878.t51 gnd 0.719405f
C4765 a_n1986_13878.t60 gnd 0.707549f
C4766 a_n1986_13878.n70 gnd 0.301556f
C4767 a_n1986_13878.t46 gnd 0.707549f
C4768 a_n1986_13878.n71 gnd 0.311083f
C4769 a_n1986_13878.t55 gnd 0.719405f
C4770 a_n1986_13878.t64 gnd 0.707549f
C4771 a_n1986_13878.n72 gnd 0.301556f
C4772 a_n1986_13878.t52 gnd 0.707549f
C4773 a_n1986_13878.n73 gnd 0.311083f
C4774 a_n1986_13878.t66 gnd 0.719405f
C4775 a_n1986_13878.t56 gnd 0.707549f
C4776 a_n1986_13878.n74 gnd 0.301556f
C4777 a_n1986_13878.t41 gnd 0.707549f
C4778 a_n1986_13878.n75 gnd 0.311083f
C4779 a_n1986_13878.t61 gnd 0.719405f
C4780 a_n1986_13878.n76 gnd 1.35928f
C4781 a_n1986_13878.n77 gnd 0.313742f
C4782 a_n1986_13878.n78 gnd 0.307133f
C4783 a_n1986_13878.n79 gnd 0.313741f
C4784 a_n1986_13878.t9 gnd 0.118309f
C4785 a_n1986_13878.t5 gnd 0.118309f
C4786 a_n1986_13878.n80 gnd 1.04709f
C4787 a_n1986_13878.t35 gnd 0.118309f
C4788 a_n1986_13878.t1 gnd 0.118309f
C4789 a_n1986_13878.n81 gnd 1.04542f
C4790 a_n1986_13878.t2 gnd 0.118309f
C4791 a_n1986_13878.t36 gnd 0.118309f
C4792 a_n1986_13878.n82 gnd 1.04709f
C4793 a_n1986_13878.t3 gnd 0.118309f
C4794 a_n1986_13878.t10 gnd 0.118309f
C4795 a_n1986_13878.n83 gnd 1.04542f
C4796 a_n1986_13878.t8 gnd 0.118309f
C4797 a_n1986_13878.t38 gnd 0.118309f
C4798 a_n1986_13878.n84 gnd 1.04542f
C4799 a_n1986_13878.t37 gnd 0.118309f
C4800 a_n1986_13878.t7 gnd 0.118309f
C4801 a_n1986_13878.n85 gnd 1.04542f
C4802 a_n1986_13878.t0 gnd 0.118309f
C4803 a_n1986_13878.t39 gnd 0.118309f
C4804 a_n1986_13878.n86 gnd 1.04709f
C4805 a_n1986_13878.t4 gnd 0.118309f
C4806 a_n1986_13878.t6 gnd 0.118309f
C4807 a_n1986_13878.n87 gnd 1.04542f
C4808 a_n1986_13878.n88 gnd 0.313742f
C4809 a_n1986_13878.n89 gnd 0.307133f
C4810 a_n1986_13878.n90 gnd 0.313741f
C4811 a_n1986_13878.n91 gnd 0.799185f
C4812 a_n1986_13878.t20 gnd 1.4243f
C4813 a_n1986_13878.t18 gnd 0.152112f
C4814 a_n1986_13878.t30 gnd 0.152112f
C4815 a_n1986_13878.n92 gnd 1.07147f
C4816 a_n1986_13878.t14 gnd 0.152112f
C4817 a_n1986_13878.t34 gnd 0.152112f
C4818 a_n1986_13878.n93 gnd 1.07147f
C4819 a_n1986_13878.n94 gnd 1.1624f
C4820 a_n1986_13878.t12 gnd 1.42146f
C4821 CSoutput.n0 gnd 0.049279f
C4822 CSoutput.t249 gnd 0.325971f
C4823 CSoutput.n1 gnd 0.147192f
C4824 CSoutput.n2 gnd 0.049279f
C4825 CSoutput.t247 gnd 0.325971f
C4826 CSoutput.n3 gnd 0.039058f
C4827 CSoutput.n4 gnd 0.049279f
C4828 CSoutput.t261 gnd 0.325971f
C4829 CSoutput.n5 gnd 0.03368f
C4830 CSoutput.n6 gnd 0.049279f
C4831 CSoutput.t244 gnd 0.325971f
C4832 CSoutput.t253 gnd 0.325971f
C4833 CSoutput.n7 gnd 0.145588f
C4834 CSoutput.n8 gnd 0.049279f
C4835 CSoutput.t252 gnd 0.325971f
C4836 CSoutput.n9 gnd 0.032112f
C4837 CSoutput.n10 gnd 0.049279f
C4838 CSoutput.t241 gnd 0.325971f
C4839 CSoutput.t245 gnd 0.325971f
C4840 CSoutput.n11 gnd 0.145588f
C4841 CSoutput.n12 gnd 0.049279f
C4842 CSoutput.t251 gnd 0.325971f
C4843 CSoutput.n13 gnd 0.03368f
C4844 CSoutput.n14 gnd 0.049279f
C4845 CSoutput.t254 gnd 0.325971f
C4846 CSoutput.t242 gnd 0.325971f
C4847 CSoutput.n15 gnd 0.145588f
C4848 CSoutput.n16 gnd 0.049279f
C4849 CSoutput.t250 gnd 0.325971f
C4850 CSoutput.n17 gnd 0.035972f
C4851 CSoutput.t258 gnd 0.389544f
C4852 CSoutput.t248 gnd 0.325971f
C4853 CSoutput.n18 gnd 0.185859f
C4854 CSoutput.n19 gnd 0.180348f
C4855 CSoutput.n20 gnd 0.209225f
C4856 CSoutput.n21 gnd 0.049279f
C4857 CSoutput.n22 gnd 0.041129f
C4858 CSoutput.n23 gnd 0.145588f
C4859 CSoutput.n24 gnd 0.039647f
C4860 CSoutput.n25 gnd 0.039058f
C4861 CSoutput.n26 gnd 0.049279f
C4862 CSoutput.n27 gnd 0.049279f
C4863 CSoutput.n28 gnd 0.040813f
C4864 CSoutput.n29 gnd 0.034651f
C4865 CSoutput.n30 gnd 0.148829f
C4866 CSoutput.n31 gnd 0.035128f
C4867 CSoutput.n32 gnd 0.049279f
C4868 CSoutput.n33 gnd 0.049279f
C4869 CSoutput.n34 gnd 0.049279f
C4870 CSoutput.n35 gnd 0.040378f
C4871 CSoutput.n36 gnd 0.145588f
C4872 CSoutput.n37 gnd 0.038616f
C4873 CSoutput.n38 gnd 0.040089f
C4874 CSoutput.n39 gnd 0.049279f
C4875 CSoutput.n40 gnd 0.049279f
C4876 CSoutput.n41 gnd 0.04112f
C4877 CSoutput.n42 gnd 0.037584f
C4878 CSoutput.n43 gnd 0.145588f
C4879 CSoutput.n44 gnd 0.038537f
C4880 CSoutput.n45 gnd 0.049279f
C4881 CSoutput.n46 gnd 0.049279f
C4882 CSoutput.n47 gnd 0.049279f
C4883 CSoutput.n48 gnd 0.038537f
C4884 CSoutput.n49 gnd 0.145588f
C4885 CSoutput.n50 gnd 0.037584f
C4886 CSoutput.n51 gnd 0.04112f
C4887 CSoutput.n52 gnd 0.049279f
C4888 CSoutput.n53 gnd 0.049279f
C4889 CSoutput.n54 gnd 0.040089f
C4890 CSoutput.n55 gnd 0.038616f
C4891 CSoutput.n56 gnd 0.145588f
C4892 CSoutput.n57 gnd 0.040378f
C4893 CSoutput.n58 gnd 0.049279f
C4894 CSoutput.n59 gnd 0.049279f
C4895 CSoutput.n60 gnd 0.049279f
C4896 CSoutput.n61 gnd 0.035128f
C4897 CSoutput.n62 gnd 0.148829f
C4898 CSoutput.n63 gnd 0.034651f
C4899 CSoutput.t257 gnd 0.325971f
C4900 CSoutput.n64 gnd 0.145588f
C4901 CSoutput.n65 gnd 0.040813f
C4902 CSoutput.n66 gnd 0.049279f
C4903 CSoutput.n67 gnd 0.049279f
C4904 CSoutput.n68 gnd 0.049279f
C4905 CSoutput.n69 gnd 0.039647f
C4906 CSoutput.n70 gnd 0.145588f
C4907 CSoutput.n71 gnd 0.041129f
C4908 CSoutput.n72 gnd 0.035972f
C4909 CSoutput.n73 gnd 0.049279f
C4910 CSoutput.n74 gnd 0.049279f
C4911 CSoutput.n75 gnd 0.037305f
C4912 CSoutput.n76 gnd 0.022156f
C4913 CSoutput.t259 gnd 0.366251f
C4914 CSoutput.n77 gnd 0.181939f
C4915 CSoutput.n78 gnd 0.744303f
C4916 CSoutput.t83 gnd 0.061469f
C4917 CSoutput.t15 gnd 0.061469f
C4918 CSoutput.n79 gnd 0.475912f
C4919 CSoutput.t73 gnd 0.061469f
C4920 CSoutput.t99 gnd 0.061469f
C4921 CSoutput.n80 gnd 0.475063f
C4922 CSoutput.n81 gnd 0.482188f
C4923 CSoutput.t64 gnd 0.061469f
C4924 CSoutput.t29 gnd 0.061469f
C4925 CSoutput.n82 gnd 0.475063f
C4926 CSoutput.n83 gnd 0.237602f
C4927 CSoutput.t9 gnd 0.061469f
C4928 CSoutput.t32 gnd 0.061469f
C4929 CSoutput.n84 gnd 0.475063f
C4930 CSoutput.n85 gnd 0.237602f
C4931 CSoutput.t17 gnd 0.061469f
C4932 CSoutput.t58 gnd 0.061469f
C4933 CSoutput.n86 gnd 0.475063f
C4934 CSoutput.n87 gnd 0.237602f
C4935 CSoutput.t18 gnd 0.061469f
C4936 CSoutput.t50 gnd 0.061469f
C4937 CSoutput.n88 gnd 0.475063f
C4938 CSoutput.n89 gnd 0.237602f
C4939 CSoutput.t76 gnd 0.061469f
C4940 CSoutput.t37 gnd 0.061469f
C4941 CSoutput.n90 gnd 0.475063f
C4942 CSoutput.n91 gnd 0.237602f
C4943 CSoutput.t87 gnd 0.061469f
C4944 CSoutput.t21 gnd 0.061469f
C4945 CSoutput.n92 gnd 0.475063f
C4946 CSoutput.n93 gnd 0.237602f
C4947 CSoutput.t89 gnd 0.061469f
C4948 CSoutput.t38 gnd 0.061469f
C4949 CSoutput.n94 gnd 0.475063f
C4950 CSoutput.n95 gnd 0.237602f
C4951 CSoutput.t53 gnd 0.061469f
C4952 CSoutput.t113 gnd 0.061469f
C4953 CSoutput.n96 gnd 0.475063f
C4954 CSoutput.n97 gnd 0.435707f
C4955 CSoutput.t238 gnd 0.061469f
C4956 CSoutput.t74 gnd 0.061469f
C4957 CSoutput.n98 gnd 0.475912f
C4958 CSoutput.t40 gnd 0.061469f
C4959 CSoutput.t16 gnd 0.061469f
C4960 CSoutput.n99 gnd 0.475063f
C4961 CSoutput.n100 gnd 0.482188f
C4962 CSoutput.t14 gnd 0.061469f
C4963 CSoutput.t62 gnd 0.061469f
C4964 CSoutput.n101 gnd 0.475063f
C4965 CSoutput.n102 gnd 0.237602f
C4966 CSoutput.t41 gnd 0.061469f
C4967 CSoutput.t34 gnd 0.061469f
C4968 CSoutput.n103 gnd 0.475063f
C4969 CSoutput.n104 gnd 0.237602f
C4970 CSoutput.t28 gnd 0.061469f
C4971 CSoutput.t84 gnd 0.061469f
C4972 CSoutput.n105 gnd 0.475063f
C4973 CSoutput.n106 gnd 0.237602f
C4974 CSoutput.t2 gnd 0.061469f
C4975 CSoutput.t3 gnd 0.061469f
C4976 CSoutput.n107 gnd 0.475063f
C4977 CSoutput.n108 gnd 0.237602f
C4978 CSoutput.t101 gnd 0.061469f
C4979 CSoutput.t88 gnd 0.061469f
C4980 CSoutput.n109 gnd 0.475063f
C4981 CSoutput.n110 gnd 0.237602f
C4982 CSoutput.t80 gnd 0.061469f
C4983 CSoutput.t100 gnd 0.061469f
C4984 CSoutput.n111 gnd 0.475063f
C4985 CSoutput.n112 gnd 0.237602f
C4986 CSoutput.t36 gnd 0.061469f
C4987 CSoutput.t48 gnd 0.061469f
C4988 CSoutput.n113 gnd 0.475063f
C4989 CSoutput.n114 gnd 0.237602f
C4990 CSoutput.t107 gnd 0.061469f
C4991 CSoutput.t79 gnd 0.061469f
C4992 CSoutput.n115 gnd 0.475063f
C4993 CSoutput.n116 gnd 0.354324f
C4994 CSoutput.n117 gnd 0.446801f
C4995 CSoutput.t22 gnd 0.061469f
C4996 CSoutput.t23 gnd 0.061469f
C4997 CSoutput.n118 gnd 0.475912f
C4998 CSoutput.t43 gnd 0.061469f
C4999 CSoutput.t27 gnd 0.061469f
C5000 CSoutput.n119 gnd 0.475063f
C5001 CSoutput.n120 gnd 0.482188f
C5002 CSoutput.t24 gnd 0.061469f
C5003 CSoutput.t85 gnd 0.061469f
C5004 CSoutput.n121 gnd 0.475063f
C5005 CSoutput.n122 gnd 0.237602f
C5006 CSoutput.t72 gnd 0.061469f
C5007 CSoutput.t59 gnd 0.061469f
C5008 CSoutput.n123 gnd 0.475063f
C5009 CSoutput.n124 gnd 0.237602f
C5010 CSoutput.t52 gnd 0.061469f
C5011 CSoutput.t5 gnd 0.061469f
C5012 CSoutput.n125 gnd 0.475063f
C5013 CSoutput.n126 gnd 0.237602f
C5014 CSoutput.t104 gnd 0.061469f
C5015 CSoutput.t105 gnd 0.061469f
C5016 CSoutput.n127 gnd 0.475063f
C5017 CSoutput.n128 gnd 0.237602f
C5018 CSoutput.t67 gnd 0.061469f
C5019 CSoutput.t95 gnd 0.061469f
C5020 CSoutput.n129 gnd 0.475063f
C5021 CSoutput.n130 gnd 0.237602f
C5022 CSoutput.t46 gnd 0.061469f
C5023 CSoutput.t66 gnd 0.061469f
C5024 CSoutput.n131 gnd 0.475063f
C5025 CSoutput.n132 gnd 0.237602f
C5026 CSoutput.t6 gnd 0.061469f
C5027 CSoutput.t51 gnd 0.061469f
C5028 CSoutput.n133 gnd 0.475063f
C5029 CSoutput.n134 gnd 0.237602f
C5030 CSoutput.t25 gnd 0.061469f
C5031 CSoutput.t86 gnd 0.061469f
C5032 CSoutput.n135 gnd 0.475063f
C5033 CSoutput.n136 gnd 0.354324f
C5034 CSoutput.n137 gnd 0.499409f
C5035 CSoutput.n138 gnd 9.86747f
C5036 CSoutput.n140 gnd 0.871739f
C5037 CSoutput.n141 gnd 0.653804f
C5038 CSoutput.n142 gnd 0.871739f
C5039 CSoutput.n143 gnd 0.871739f
C5040 CSoutput.n144 gnd 2.34699f
C5041 CSoutput.n145 gnd 0.871739f
C5042 CSoutput.n146 gnd 0.871739f
C5043 CSoutput.t255 gnd 1.08967f
C5044 CSoutput.n147 gnd 0.871739f
C5045 CSoutput.n148 gnd 0.871739f
C5046 CSoutput.n152 gnd 0.871739f
C5047 CSoutput.n156 gnd 0.871739f
C5048 CSoutput.n157 gnd 0.871739f
C5049 CSoutput.n159 gnd 0.871739f
C5050 CSoutput.n164 gnd 0.871739f
C5051 CSoutput.n166 gnd 0.871739f
C5052 CSoutput.n167 gnd 0.871739f
C5053 CSoutput.n169 gnd 0.871739f
C5054 CSoutput.n170 gnd 0.871739f
C5055 CSoutput.n172 gnd 0.871739f
C5056 CSoutput.t243 gnd 14.5667f
C5057 CSoutput.n174 gnd 0.871739f
C5058 CSoutput.n175 gnd 0.653804f
C5059 CSoutput.n176 gnd 0.871739f
C5060 CSoutput.n177 gnd 0.871739f
C5061 CSoutput.n178 gnd 2.34699f
C5062 CSoutput.n179 gnd 0.871739f
C5063 CSoutput.n180 gnd 0.871739f
C5064 CSoutput.t260 gnd 1.08967f
C5065 CSoutput.n181 gnd 0.871739f
C5066 CSoutput.n182 gnd 0.871739f
C5067 CSoutput.n186 gnd 0.871739f
C5068 CSoutput.n190 gnd 0.871739f
C5069 CSoutput.n191 gnd 0.871739f
C5070 CSoutput.n193 gnd 0.871739f
C5071 CSoutput.n198 gnd 0.871739f
C5072 CSoutput.n200 gnd 0.871739f
C5073 CSoutput.n201 gnd 0.871739f
C5074 CSoutput.n203 gnd 0.871739f
C5075 CSoutput.n204 gnd 0.871739f
C5076 CSoutput.n206 gnd 0.871739f
C5077 CSoutput.n207 gnd 0.653804f
C5078 CSoutput.n209 gnd 0.871739f
C5079 CSoutput.n210 gnd 0.653804f
C5080 CSoutput.n211 gnd 0.871739f
C5081 CSoutput.n212 gnd 0.871739f
C5082 CSoutput.n213 gnd 2.34699f
C5083 CSoutput.n214 gnd 0.871739f
C5084 CSoutput.n215 gnd 0.871739f
C5085 CSoutput.t256 gnd 1.08967f
C5086 CSoutput.n216 gnd 0.871739f
C5087 CSoutput.n217 gnd 2.34699f
C5088 CSoutput.n219 gnd 0.871739f
C5089 CSoutput.n220 gnd 0.871739f
C5090 CSoutput.n222 gnd 0.871739f
C5091 CSoutput.n223 gnd 0.871739f
C5092 CSoutput.t240 gnd 14.329301f
C5093 CSoutput.t246 gnd 14.5667f
C5094 CSoutput.n229 gnd 2.73477f
C5095 CSoutput.n230 gnd 11.1405f
C5096 CSoutput.n231 gnd 11.6066f
C5097 CSoutput.n236 gnd 2.9625f
C5098 CSoutput.n242 gnd 0.871739f
C5099 CSoutput.n244 gnd 0.871739f
C5100 CSoutput.n246 gnd 0.871739f
C5101 CSoutput.n248 gnd 0.871739f
C5102 CSoutput.n250 gnd 0.871739f
C5103 CSoutput.n256 gnd 0.871739f
C5104 CSoutput.n263 gnd 1.59931f
C5105 CSoutput.n264 gnd 1.59931f
C5106 CSoutput.n265 gnd 0.871739f
C5107 CSoutput.n266 gnd 0.871739f
C5108 CSoutput.n268 gnd 0.653804f
C5109 CSoutput.n269 gnd 0.559925f
C5110 CSoutput.n271 gnd 0.653804f
C5111 CSoutput.n272 gnd 0.559925f
C5112 CSoutput.n273 gnd 0.653804f
C5113 CSoutput.n275 gnd 0.871739f
C5114 CSoutput.n277 gnd 2.34699f
C5115 CSoutput.n278 gnd 2.73477f
C5116 CSoutput.n279 gnd 10.2464f
C5117 CSoutput.n281 gnd 0.653804f
C5118 CSoutput.n282 gnd 1.68228f
C5119 CSoutput.n283 gnd 0.653804f
C5120 CSoutput.n285 gnd 0.871739f
C5121 CSoutput.n287 gnd 2.34699f
C5122 CSoutput.n288 gnd 5.11212f
C5123 CSoutput.t78 gnd 0.061469f
C5124 CSoutput.t110 gnd 0.061469f
C5125 CSoutput.n289 gnd 0.475912f
C5126 CSoutput.t96 gnd 0.061469f
C5127 CSoutput.t77 gnd 0.061469f
C5128 CSoutput.n290 gnd 0.475063f
C5129 CSoutput.n291 gnd 0.482188f
C5130 CSoutput.t90 gnd 0.061469f
C5131 CSoutput.t65 gnd 0.061469f
C5132 CSoutput.n292 gnd 0.475063f
C5133 CSoutput.n293 gnd 0.237602f
C5134 CSoutput.t33 gnd 0.061469f
C5135 CSoutput.t115 gnd 0.061469f
C5136 CSoutput.n294 gnd 0.475063f
C5137 CSoutput.n295 gnd 0.237602f
C5138 CSoutput.t71 gnd 0.061469f
C5139 CSoutput.t81 gnd 0.061469f
C5140 CSoutput.n296 gnd 0.475063f
C5141 CSoutput.n297 gnd 0.237602f
C5142 CSoutput.t30 gnd 0.061469f
C5143 CSoutput.t19 gnd 0.061469f
C5144 CSoutput.n298 gnd 0.475063f
C5145 CSoutput.n299 gnd 0.237602f
C5146 CSoutput.t98 gnd 0.061469f
C5147 CSoutput.t93 gnd 0.061469f
C5148 CSoutput.n300 gnd 0.475063f
C5149 CSoutput.n301 gnd 0.237602f
C5150 CSoutput.t237 gnd 0.061469f
C5151 CSoutput.t10 gnd 0.061469f
C5152 CSoutput.n302 gnd 0.475063f
C5153 CSoutput.n303 gnd 0.237602f
C5154 CSoutput.t39 gnd 0.061469f
C5155 CSoutput.t26 gnd 0.061469f
C5156 CSoutput.n304 gnd 0.475063f
C5157 CSoutput.n305 gnd 0.237602f
C5158 CSoutput.t70 gnd 0.061469f
C5159 CSoutput.t94 gnd 0.061469f
C5160 CSoutput.n306 gnd 0.475063f
C5161 CSoutput.n307 gnd 0.435707f
C5162 CSoutput.t57 gnd 0.061469f
C5163 CSoutput.t56 gnd 0.061469f
C5164 CSoutput.n308 gnd 0.475912f
C5165 CSoutput.t102 gnd 0.061469f
C5166 CSoutput.t106 gnd 0.061469f
C5167 CSoutput.n309 gnd 0.475063f
C5168 CSoutput.n310 gnd 0.482188f
C5169 CSoutput.t54 gnd 0.061469f
C5170 CSoutput.t61 gnd 0.061469f
C5171 CSoutput.n311 gnd 0.475063f
C5172 CSoutput.n312 gnd 0.237602f
C5173 CSoutput.t4 gnd 0.061469f
C5174 CSoutput.t92 gnd 0.061469f
C5175 CSoutput.n313 gnd 0.475063f
C5176 CSoutput.n314 gnd 0.237602f
C5177 CSoutput.t31 gnd 0.061469f
C5178 CSoutput.t82 gnd 0.061469f
C5179 CSoutput.n315 gnd 0.475063f
C5180 CSoutput.n316 gnd 0.237602f
C5181 CSoutput.t13 gnd 0.061469f
C5182 CSoutput.t12 gnd 0.061469f
C5183 CSoutput.n317 gnd 0.475063f
C5184 CSoutput.n318 gnd 0.237602f
C5185 CSoutput.t20 gnd 0.061469f
C5186 CSoutput.t111 gnd 0.061469f
C5187 CSoutput.n319 gnd 0.475063f
C5188 CSoutput.n320 gnd 0.237602f
C5189 CSoutput.t108 gnd 0.061469f
C5190 CSoutput.t103 gnd 0.061469f
C5191 CSoutput.n321 gnd 0.475063f
C5192 CSoutput.n322 gnd 0.237602f
C5193 CSoutput.t236 gnd 0.061469f
C5194 CSoutput.t109 gnd 0.061469f
C5195 CSoutput.n323 gnd 0.475063f
C5196 CSoutput.n324 gnd 0.237602f
C5197 CSoutput.t97 gnd 0.061469f
C5198 CSoutput.t60 gnd 0.061469f
C5199 CSoutput.n325 gnd 0.475063f
C5200 CSoutput.n326 gnd 0.354324f
C5201 CSoutput.n327 gnd 0.446801f
C5202 CSoutput.t69 gnd 0.061469f
C5203 CSoutput.t68 gnd 0.061469f
C5204 CSoutput.n328 gnd 0.475912f
C5205 CSoutput.t239 gnd 0.061469f
C5206 CSoutput.t47 gnd 0.061469f
C5207 CSoutput.n329 gnd 0.475063f
C5208 CSoutput.n330 gnd 0.482188f
C5209 CSoutput.t112 gnd 0.061469f
C5210 CSoutput.t42 gnd 0.061469f
C5211 CSoutput.n331 gnd 0.475063f
C5212 CSoutput.n332 gnd 0.237602f
C5213 CSoutput.t11 gnd 0.061469f
C5214 CSoutput.t35 gnd 0.061469f
C5215 CSoutput.n333 gnd 0.475063f
C5216 CSoutput.n334 gnd 0.237602f
C5217 CSoutput.t55 gnd 0.061469f
C5218 CSoutput.t44 gnd 0.061469f
C5219 CSoutput.n335 gnd 0.475063f
C5220 CSoutput.n336 gnd 0.237602f
C5221 CSoutput.t1 gnd 0.061469f
C5222 CSoutput.t0 gnd 0.061469f
C5223 CSoutput.n337 gnd 0.475063f
C5224 CSoutput.n338 gnd 0.237602f
C5225 CSoutput.t8 gnd 0.061469f
C5226 CSoutput.t45 gnd 0.061469f
C5227 CSoutput.n339 gnd 0.475063f
C5228 CSoutput.n340 gnd 0.237602f
C5229 CSoutput.t91 gnd 0.061469f
C5230 CSoutput.t75 gnd 0.061469f
C5231 CSoutput.n341 gnd 0.475063f
C5232 CSoutput.n342 gnd 0.237602f
C5233 CSoutput.t114 gnd 0.061469f
C5234 CSoutput.t49 gnd 0.061469f
C5235 CSoutput.n343 gnd 0.475063f
C5236 CSoutput.n344 gnd 0.237602f
C5237 CSoutput.t7 gnd 0.061469f
C5238 CSoutput.t63 gnd 0.061469f
C5239 CSoutput.n345 gnd 0.475061f
C5240 CSoutput.n346 gnd 0.354326f
C5241 CSoutput.n347 gnd 0.499409f
C5242 CSoutput.n348 gnd 13.799999f
C5243 CSoutput.t164 gnd 0.053785f
C5244 CSoutput.t232 gnd 0.053785f
C5245 CSoutput.n349 gnd 0.476855f
C5246 CSoutput.t154 gnd 0.053785f
C5247 CSoutput.t163 gnd 0.053785f
C5248 CSoutput.n350 gnd 0.475265f
C5249 CSoutput.n351 gnd 0.442858f
C5250 CSoutput.t144 gnd 0.053785f
C5251 CSoutput.t170 gnd 0.053785f
C5252 CSoutput.n352 gnd 0.475265f
C5253 CSoutput.n353 gnd 0.218308f
C5254 CSoutput.t191 gnd 0.053785f
C5255 CSoutput.t157 gnd 0.053785f
C5256 CSoutput.n354 gnd 0.475265f
C5257 CSoutput.n355 gnd 0.218308f
C5258 CSoutput.t167 gnd 0.053785f
C5259 CSoutput.t222 gnd 0.053785f
C5260 CSoutput.n356 gnd 0.475265f
C5261 CSoutput.n357 gnd 0.218308f
C5262 CSoutput.t184 gnd 0.053785f
C5263 CSoutput.t198 gnd 0.053785f
C5264 CSoutput.n358 gnd 0.475265f
C5265 CSoutput.n359 gnd 0.218308f
C5266 CSoutput.t139 gnd 0.053785f
C5267 CSoutput.t171 gnd 0.053785f
C5268 CSoutput.n360 gnd 0.475265f
C5269 CSoutput.n361 gnd 0.218308f
C5270 CSoutput.t125 gnd 0.053785f
C5271 CSoutput.t151 gnd 0.053785f
C5272 CSoutput.n362 gnd 0.475265f
C5273 CSoutput.n363 gnd 0.218308f
C5274 CSoutput.t204 gnd 0.053785f
C5275 CSoutput.t215 gnd 0.053785f
C5276 CSoutput.n364 gnd 0.475265f
C5277 CSoutput.n365 gnd 0.218308f
C5278 CSoutput.t231 gnd 0.053785f
C5279 CSoutput.t175 gnd 0.053785f
C5280 CSoutput.n366 gnd 0.475265f
C5281 CSoutput.n367 gnd 0.402657f
C5282 CSoutput.t227 gnd 0.053785f
C5283 CSoutput.t117 gnd 0.053785f
C5284 CSoutput.n368 gnd 0.476855f
C5285 CSoutput.t129 gnd 0.053785f
C5286 CSoutput.t220 gnd 0.053785f
C5287 CSoutput.n369 gnd 0.475265f
C5288 CSoutput.n370 gnd 0.442858f
C5289 CSoutput.t119 gnd 0.053785f
C5290 CSoutput.t210 gnd 0.053785f
C5291 CSoutput.n371 gnd 0.475265f
C5292 CSoutput.n372 gnd 0.218308f
C5293 CSoutput.t221 gnd 0.053785f
C5294 CSoutput.t118 gnd 0.053785f
C5295 CSoutput.n373 gnd 0.475265f
C5296 CSoutput.n374 gnd 0.218308f
C5297 CSoutput.t200 gnd 0.053785f
C5298 CSoutput.t174 gnd 0.053785f
C5299 CSoutput.n375 gnd 0.475265f
C5300 CSoutput.n376 gnd 0.218308f
C5301 CSoutput.t120 gnd 0.053785f
C5302 CSoutput.t202 gnd 0.053785f
C5303 CSoutput.n377 gnd 0.475265f
C5304 CSoutput.n378 gnd 0.218308f
C5305 CSoutput.t177 gnd 0.053785f
C5306 CSoutput.t185 gnd 0.053785f
C5307 CSoutput.n379 gnd 0.475265f
C5308 CSoutput.n380 gnd 0.218308f
C5309 CSoutput.t201 gnd 0.053785f
C5310 CSoutput.t176 gnd 0.053785f
C5311 CSoutput.n381 gnd 0.475265f
C5312 CSoutput.n382 gnd 0.218308f
C5313 CSoutput.t186 gnd 0.053785f
C5314 CSoutput.t190 gnd 0.053785f
C5315 CSoutput.n383 gnd 0.475265f
C5316 CSoutput.n384 gnd 0.218308f
C5317 CSoutput.t168 gnd 0.053785f
C5318 CSoutput.t181 gnd 0.053785f
C5319 CSoutput.n385 gnd 0.475265f
C5320 CSoutput.n386 gnd 0.331438f
C5321 CSoutput.n387 gnd 0.418047f
C5322 CSoutput.t132 gnd 0.053785f
C5323 CSoutput.t223 gnd 0.053785f
C5324 CSoutput.n388 gnd 0.476855f
C5325 CSoutput.t152 gnd 0.053785f
C5326 CSoutput.t158 gnd 0.053785f
C5327 CSoutput.n389 gnd 0.475265f
C5328 CSoutput.n390 gnd 0.442858f
C5329 CSoutput.t121 gnd 0.053785f
C5330 CSoutput.t205 gnd 0.053785f
C5331 CSoutput.n391 gnd 0.475265f
C5332 CSoutput.n392 gnd 0.218308f
C5333 CSoutput.t166 gnd 0.053785f
C5334 CSoutput.t133 gnd 0.053785f
C5335 CSoutput.n393 gnd 0.475265f
C5336 CSoutput.n394 gnd 0.218308f
C5337 CSoutput.t142 gnd 0.053785f
C5338 CSoutput.t235 gnd 0.053785f
C5339 CSoutput.n395 gnd 0.475265f
C5340 CSoutput.n396 gnd 0.218308f
C5341 CSoutput.t143 gnd 0.053785f
C5342 CSoutput.t147 gnd 0.053785f
C5343 CSoutput.n397 gnd 0.475265f
C5344 CSoutput.n398 gnd 0.218308f
C5345 CSoutput.t128 gnd 0.053785f
C5346 CSoutput.t219 gnd 0.053785f
C5347 CSoutput.n399 gnd 0.475265f
C5348 CSoutput.n400 gnd 0.218308f
C5349 CSoutput.t150 gnd 0.053785f
C5350 CSoutput.t140 gnd 0.053785f
C5351 CSoutput.n401 gnd 0.475265f
C5352 CSoutput.n402 gnd 0.218308f
C5353 CSoutput.t116 gnd 0.053785f
C5354 CSoutput.t160 gnd 0.053785f
C5355 CSoutput.n403 gnd 0.475265f
C5356 CSoutput.n404 gnd 0.218308f
C5357 CSoutput.t165 gnd 0.053785f
C5358 CSoutput.t131 gnd 0.053785f
C5359 CSoutput.n405 gnd 0.475265f
C5360 CSoutput.n406 gnd 0.331438f
C5361 CSoutput.n407 gnd 0.448917f
C5362 CSoutput.n408 gnd 14.4386f
C5363 CSoutput.t146 gnd 0.053785f
C5364 CSoutput.t203 gnd 0.053785f
C5365 CSoutput.n409 gnd 0.476855f
C5366 CSoutput.t199 gnd 0.053785f
C5367 CSoutput.t173 gnd 0.053785f
C5368 CSoutput.n410 gnd 0.475265f
C5369 CSoutput.n411 gnd 0.442858f
C5370 CSoutput.t207 gnd 0.053785f
C5371 CSoutput.t161 gnd 0.053785f
C5372 CSoutput.n412 gnd 0.475265f
C5373 CSoutput.n413 gnd 0.218308f
C5374 CSoutput.t187 gnd 0.053785f
C5375 CSoutput.t225 gnd 0.053785f
C5376 CSoutput.n414 gnd 0.475265f
C5377 CSoutput.n415 gnd 0.218308f
C5378 CSoutput.t141 gnd 0.053785f
C5379 CSoutput.t206 gnd 0.053785f
C5380 CSoutput.n416 gnd 0.475265f
C5381 CSoutput.n417 gnd 0.218308f
C5382 CSoutput.t127 gnd 0.053785f
C5383 CSoutput.t213 gnd 0.053785f
C5384 CSoutput.n418 gnd 0.475265f
C5385 CSoutput.n419 gnd 0.218308f
C5386 CSoutput.t212 gnd 0.053785f
C5387 CSoutput.t153 gnd 0.053785f
C5388 CSoutput.n420 gnd 0.475265f
C5389 CSoutput.n421 gnd 0.218308f
C5390 CSoutput.t180 gnd 0.053785f
C5391 CSoutput.t149 gnd 0.053785f
C5392 CSoutput.n422 gnd 0.475265f
C5393 CSoutput.n423 gnd 0.218308f
C5394 CSoutput.t155 gnd 0.053785f
C5395 CSoutput.t130 gnd 0.053785f
C5396 CSoutput.n424 gnd 0.475265f
C5397 CSoutput.n425 gnd 0.218308f
C5398 CSoutput.t138 gnd 0.053785f
C5399 CSoutput.t156 gnd 0.053785f
C5400 CSoutput.n426 gnd 0.475265f
C5401 CSoutput.n427 gnd 0.402657f
C5402 CSoutput.t135 gnd 0.053785f
C5403 CSoutput.t126 gnd 0.053785f
C5404 CSoutput.n428 gnd 0.476855f
C5405 CSoutput.t122 gnd 0.053785f
C5406 CSoutput.t233 gnd 0.053785f
C5407 CSoutput.n429 gnd 0.475265f
C5408 CSoutput.n430 gnd 0.442858f
C5409 CSoutput.t234 gnd 0.053785f
C5410 CSoutput.t136 gnd 0.053785f
C5411 CSoutput.n431 gnd 0.475265f
C5412 CSoutput.n432 gnd 0.218308f
C5413 CSoutput.t137 gnd 0.053785f
C5414 CSoutput.t194 gnd 0.053785f
C5415 CSoutput.n433 gnd 0.475265f
C5416 CSoutput.n434 gnd 0.218308f
C5417 CSoutput.t195 gnd 0.053785f
C5418 CSoutput.t226 gnd 0.053785f
C5419 CSoutput.n435 gnd 0.475265f
C5420 CSoutput.n436 gnd 0.218308f
C5421 CSoutput.t229 gnd 0.053785f
C5422 CSoutput.t218 gnd 0.053785f
C5423 CSoutput.n437 gnd 0.475265f
C5424 CSoutput.n438 gnd 0.218308f
C5425 CSoutput.t209 gnd 0.053785f
C5426 CSoutput.t196 gnd 0.053785f
C5427 CSoutput.n439 gnd 0.475265f
C5428 CSoutput.n440 gnd 0.218308f
C5429 CSoutput.t197 gnd 0.053785f
C5430 CSoutput.t230 gnd 0.053785f
C5431 CSoutput.n441 gnd 0.475265f
C5432 CSoutput.n442 gnd 0.218308f
C5433 CSoutput.t183 gnd 0.053785f
C5434 CSoutput.t211 gnd 0.053785f
C5435 CSoutput.n443 gnd 0.475265f
C5436 CSoutput.n444 gnd 0.218308f
C5437 CSoutput.t217 gnd 0.053785f
C5438 CSoutput.t192 gnd 0.053785f
C5439 CSoutput.n445 gnd 0.475265f
C5440 CSoutput.n446 gnd 0.331438f
C5441 CSoutput.n447 gnd 0.418047f
C5442 CSoutput.t182 gnd 0.053785f
C5443 CSoutput.t214 gnd 0.053785f
C5444 CSoutput.n448 gnd 0.476855f
C5445 CSoutput.t145 gnd 0.053785f
C5446 CSoutput.t162 gnd 0.053785f
C5447 CSoutput.n449 gnd 0.475265f
C5448 CSoutput.n450 gnd 0.442858f
C5449 CSoutput.t172 gnd 0.053785f
C5450 CSoutput.t193 gnd 0.053785f
C5451 CSoutput.n451 gnd 0.475265f
C5452 CSoutput.n452 gnd 0.218308f
C5453 CSoutput.t216 gnd 0.053785f
C5454 CSoutput.t178 gnd 0.053785f
C5455 CSoutput.n453 gnd 0.475265f
C5456 CSoutput.n454 gnd 0.218308f
C5457 CSoutput.t188 gnd 0.053785f
C5458 CSoutput.t228 gnd 0.053785f
C5459 CSoutput.n455 gnd 0.475265f
C5460 CSoutput.n456 gnd 0.218308f
C5461 CSoutput.t123 gnd 0.053785f
C5462 CSoutput.t148 gnd 0.053785f
C5463 CSoutput.n457 gnd 0.475265f
C5464 CSoutput.n458 gnd 0.218308f
C5465 CSoutput.t179 gnd 0.053785f
C5466 CSoutput.t208 gnd 0.053785f
C5467 CSoutput.n459 gnd 0.475265f
C5468 CSoutput.n460 gnd 0.218308f
C5469 CSoutput.t224 gnd 0.053785f
C5470 CSoutput.t134 gnd 0.053785f
C5471 CSoutput.n461 gnd 0.475265f
C5472 CSoutput.n462 gnd 0.218308f
C5473 CSoutput.t169 gnd 0.053785f
C5474 CSoutput.t189 gnd 0.053785f
C5475 CSoutput.n463 gnd 0.475265f
C5476 CSoutput.n464 gnd 0.218308f
C5477 CSoutput.t124 gnd 0.053785f
C5478 CSoutput.t159 gnd 0.053785f
C5479 CSoutput.n465 gnd 0.475265f
C5480 CSoutput.n466 gnd 0.331438f
C5481 CSoutput.n467 gnd 0.448917f
C5482 CSoutput.n468 gnd 8.57409f
C5483 CSoutput.n469 gnd 15.068401f
C5484 commonsourceibias.n0 gnd 0.012817f
C5485 commonsourceibias.t151 gnd 0.194086f
C5486 commonsourceibias.t83 gnd 0.17946f
C5487 commonsourceibias.n1 gnd 0.009349f
C5488 commonsourceibias.n2 gnd 0.009605f
C5489 commonsourceibias.t161 gnd 0.17946f
C5490 commonsourceibias.n3 gnd 0.012358f
C5491 commonsourceibias.n4 gnd 0.009605f
C5492 commonsourceibias.t152 gnd 0.17946f
C5493 commonsourceibias.n5 gnd 0.071604f
C5494 commonsourceibias.t171 gnd 0.17946f
C5495 commonsourceibias.n6 gnd 0.009057f
C5496 commonsourceibias.n7 gnd 0.009605f
C5497 commonsourceibias.t145 gnd 0.17946f
C5498 commonsourceibias.n8 gnd 0.012174f
C5499 commonsourceibias.n9 gnd 0.009605f
C5500 commonsourceibias.t124 gnd 0.17946f
C5501 commonsourceibias.n10 gnd 0.071604f
C5502 commonsourceibias.t158 gnd 0.17946f
C5503 commonsourceibias.n11 gnd 0.008798f
C5504 commonsourceibias.n12 gnd 0.009605f
C5505 commonsourceibias.t148 gnd 0.17946f
C5506 commonsourceibias.n13 gnd 0.01197f
C5507 commonsourceibias.n14 gnd 0.012817f
C5508 commonsourceibias.t52 gnd 0.194086f
C5509 commonsourceibias.t20 gnd 0.17946f
C5510 commonsourceibias.n15 gnd 0.009349f
C5511 commonsourceibias.n16 gnd 0.009605f
C5512 commonsourceibias.t66 gnd 0.17946f
C5513 commonsourceibias.n17 gnd 0.012358f
C5514 commonsourceibias.n18 gnd 0.009605f
C5515 commonsourceibias.t50 gnd 0.17946f
C5516 commonsourceibias.n19 gnd 0.071604f
C5517 commonsourceibias.t0 gnd 0.17946f
C5518 commonsourceibias.n20 gnd 0.009057f
C5519 commonsourceibias.n21 gnd 0.009605f
C5520 commonsourceibias.t56 gnd 0.17946f
C5521 commonsourceibias.n22 gnd 0.012174f
C5522 commonsourceibias.n23 gnd 0.009605f
C5523 commonsourceibias.t42 gnd 0.17946f
C5524 commonsourceibias.n24 gnd 0.071604f
C5525 commonsourceibias.t72 gnd 0.17946f
C5526 commonsourceibias.n25 gnd 0.008798f
C5527 commonsourceibias.n26 gnd 0.009605f
C5528 commonsourceibias.t54 gnd 0.17946f
C5529 commonsourceibias.n27 gnd 0.01197f
C5530 commonsourceibias.n28 gnd 0.009605f
C5531 commonsourceibias.t34 gnd 0.17946f
C5532 commonsourceibias.n29 gnd 0.071604f
C5533 commonsourceibias.t38 gnd 0.17946f
C5534 commonsourceibias.n30 gnd 0.008571f
C5535 commonsourceibias.n31 gnd 0.009605f
C5536 commonsourceibias.t44 gnd 0.17946f
C5537 commonsourceibias.n32 gnd 0.011742f
C5538 commonsourceibias.n33 gnd 0.009605f
C5539 commonsourceibias.t6 gnd 0.17946f
C5540 commonsourceibias.n34 gnd 0.071604f
C5541 commonsourceibias.t58 gnd 0.17946f
C5542 commonsourceibias.n35 gnd 0.008375f
C5543 commonsourceibias.n36 gnd 0.009605f
C5544 commonsourceibias.t10 gnd 0.17946f
C5545 commonsourceibias.n37 gnd 0.011489f
C5546 commonsourceibias.n38 gnd 0.009605f
C5547 commonsourceibias.t76 gnd 0.17946f
C5548 commonsourceibias.n39 gnd 0.071604f
C5549 commonsourceibias.t22 gnd 0.17946f
C5550 commonsourceibias.n40 gnd 0.008208f
C5551 commonsourceibias.n41 gnd 0.009605f
C5552 commonsourceibias.t32 gnd 0.17946f
C5553 commonsourceibias.n42 gnd 0.011208f
C5554 commonsourceibias.t62 gnd 0.199526f
C5555 commonsourceibias.t18 gnd 0.17946f
C5556 commonsourceibias.n43 gnd 0.078221f
C5557 commonsourceibias.n44 gnd 0.085838f
C5558 commonsourceibias.n45 gnd 0.03983f
C5559 commonsourceibias.n46 gnd 0.009605f
C5560 commonsourceibias.n47 gnd 0.009349f
C5561 commonsourceibias.n48 gnd 0.013398f
C5562 commonsourceibias.n49 gnd 0.071604f
C5563 commonsourceibias.n50 gnd 0.013389f
C5564 commonsourceibias.n51 gnd 0.009605f
C5565 commonsourceibias.n52 gnd 0.009605f
C5566 commonsourceibias.n53 gnd 0.009605f
C5567 commonsourceibias.n54 gnd 0.012358f
C5568 commonsourceibias.n55 gnd 0.071604f
C5569 commonsourceibias.n56 gnd 0.012648f
C5570 commonsourceibias.n57 gnd 0.012288f
C5571 commonsourceibias.n58 gnd 0.009605f
C5572 commonsourceibias.n59 gnd 0.009605f
C5573 commonsourceibias.n60 gnd 0.009605f
C5574 commonsourceibias.n61 gnd 0.009057f
C5575 commonsourceibias.n62 gnd 0.01341f
C5576 commonsourceibias.n63 gnd 0.071604f
C5577 commonsourceibias.n64 gnd 0.013406f
C5578 commonsourceibias.n65 gnd 0.009605f
C5579 commonsourceibias.n66 gnd 0.009605f
C5580 commonsourceibias.n67 gnd 0.009605f
C5581 commonsourceibias.n68 gnd 0.012174f
C5582 commonsourceibias.n69 gnd 0.071604f
C5583 commonsourceibias.n70 gnd 0.012558f
C5584 commonsourceibias.n71 gnd 0.012378f
C5585 commonsourceibias.n72 gnd 0.009605f
C5586 commonsourceibias.n73 gnd 0.009605f
C5587 commonsourceibias.n74 gnd 0.009605f
C5588 commonsourceibias.n75 gnd 0.008798f
C5589 commonsourceibias.n76 gnd 0.013415f
C5590 commonsourceibias.n77 gnd 0.071604f
C5591 commonsourceibias.n78 gnd 0.013414f
C5592 commonsourceibias.n79 gnd 0.009605f
C5593 commonsourceibias.n80 gnd 0.009605f
C5594 commonsourceibias.n81 gnd 0.009605f
C5595 commonsourceibias.n82 gnd 0.01197f
C5596 commonsourceibias.n83 gnd 0.071604f
C5597 commonsourceibias.n84 gnd 0.012468f
C5598 commonsourceibias.n85 gnd 0.012468f
C5599 commonsourceibias.n86 gnd 0.009605f
C5600 commonsourceibias.n87 gnd 0.009605f
C5601 commonsourceibias.n88 gnd 0.009605f
C5602 commonsourceibias.n89 gnd 0.008571f
C5603 commonsourceibias.n90 gnd 0.013414f
C5604 commonsourceibias.n91 gnd 0.071604f
C5605 commonsourceibias.n92 gnd 0.013415f
C5606 commonsourceibias.n93 gnd 0.009605f
C5607 commonsourceibias.n94 gnd 0.009605f
C5608 commonsourceibias.n95 gnd 0.009605f
C5609 commonsourceibias.n96 gnd 0.011742f
C5610 commonsourceibias.n97 gnd 0.071604f
C5611 commonsourceibias.n98 gnd 0.012378f
C5612 commonsourceibias.n99 gnd 0.012558f
C5613 commonsourceibias.n100 gnd 0.009605f
C5614 commonsourceibias.n101 gnd 0.009605f
C5615 commonsourceibias.n102 gnd 0.009605f
C5616 commonsourceibias.n103 gnd 0.008375f
C5617 commonsourceibias.n104 gnd 0.013406f
C5618 commonsourceibias.n105 gnd 0.071604f
C5619 commonsourceibias.n106 gnd 0.01341f
C5620 commonsourceibias.n107 gnd 0.009605f
C5621 commonsourceibias.n108 gnd 0.009605f
C5622 commonsourceibias.n109 gnd 0.009605f
C5623 commonsourceibias.n110 gnd 0.011489f
C5624 commonsourceibias.n111 gnd 0.071604f
C5625 commonsourceibias.n112 gnd 0.012288f
C5626 commonsourceibias.n113 gnd 0.012648f
C5627 commonsourceibias.n114 gnd 0.009605f
C5628 commonsourceibias.n115 gnd 0.009605f
C5629 commonsourceibias.n116 gnd 0.009605f
C5630 commonsourceibias.n117 gnd 0.008208f
C5631 commonsourceibias.n118 gnd 0.013389f
C5632 commonsourceibias.n119 gnd 0.071604f
C5633 commonsourceibias.n120 gnd 0.013398f
C5634 commonsourceibias.n121 gnd 0.009605f
C5635 commonsourceibias.n122 gnd 0.009605f
C5636 commonsourceibias.n123 gnd 0.009605f
C5637 commonsourceibias.n124 gnd 0.011208f
C5638 commonsourceibias.n125 gnd 0.071604f
C5639 commonsourceibias.n126 gnd 0.011785f
C5640 commonsourceibias.n127 gnd 0.085919f
C5641 commonsourceibias.n128 gnd 0.095702f
C5642 commonsourceibias.t53 gnd 0.020728f
C5643 commonsourceibias.t21 gnd 0.020728f
C5644 commonsourceibias.n129 gnd 0.183157f
C5645 commonsourceibias.n130 gnd 0.158432f
C5646 commonsourceibias.t67 gnd 0.020728f
C5647 commonsourceibias.t51 gnd 0.020728f
C5648 commonsourceibias.n131 gnd 0.183157f
C5649 commonsourceibias.n132 gnd 0.084131f
C5650 commonsourceibias.t1 gnd 0.020728f
C5651 commonsourceibias.t57 gnd 0.020728f
C5652 commonsourceibias.n133 gnd 0.183157f
C5653 commonsourceibias.n134 gnd 0.084131f
C5654 commonsourceibias.t43 gnd 0.020728f
C5655 commonsourceibias.t73 gnd 0.020728f
C5656 commonsourceibias.n135 gnd 0.183157f
C5657 commonsourceibias.n136 gnd 0.084131f
C5658 commonsourceibias.t55 gnd 0.020728f
C5659 commonsourceibias.t35 gnd 0.020728f
C5660 commonsourceibias.n137 gnd 0.183157f
C5661 commonsourceibias.n138 gnd 0.070287f
C5662 commonsourceibias.t19 gnd 0.020728f
C5663 commonsourceibias.t63 gnd 0.020728f
C5664 commonsourceibias.n139 gnd 0.18377f
C5665 commonsourceibias.t23 gnd 0.020728f
C5666 commonsourceibias.t33 gnd 0.020728f
C5667 commonsourceibias.n140 gnd 0.183157f
C5668 commonsourceibias.n141 gnd 0.170668f
C5669 commonsourceibias.t11 gnd 0.020728f
C5670 commonsourceibias.t77 gnd 0.020728f
C5671 commonsourceibias.n142 gnd 0.183157f
C5672 commonsourceibias.n143 gnd 0.084131f
C5673 commonsourceibias.t7 gnd 0.020728f
C5674 commonsourceibias.t59 gnd 0.020728f
C5675 commonsourceibias.n144 gnd 0.183157f
C5676 commonsourceibias.n145 gnd 0.084131f
C5677 commonsourceibias.t39 gnd 0.020728f
C5678 commonsourceibias.t45 gnd 0.020728f
C5679 commonsourceibias.n146 gnd 0.183157f
C5680 commonsourceibias.n147 gnd 0.070287f
C5681 commonsourceibias.n148 gnd 0.085111f
C5682 commonsourceibias.n149 gnd 0.062167f
C5683 commonsourceibias.t93 gnd 0.17946f
C5684 commonsourceibias.n150 gnd 0.071604f
C5685 commonsourceibias.t131 gnd 0.17946f
C5686 commonsourceibias.n151 gnd 0.071604f
C5687 commonsourceibias.n152 gnd 0.009605f
C5688 commonsourceibias.t117 gnd 0.17946f
C5689 commonsourceibias.n153 gnd 0.071604f
C5690 commonsourceibias.n154 gnd 0.009605f
C5691 commonsourceibias.t176 gnd 0.17946f
C5692 commonsourceibias.n155 gnd 0.071604f
C5693 commonsourceibias.n156 gnd 0.009605f
C5694 commonsourceibias.t144 gnd 0.17946f
C5695 commonsourceibias.n157 gnd 0.008375f
C5696 commonsourceibias.n158 gnd 0.009605f
C5697 commonsourceibias.t190 gnd 0.17946f
C5698 commonsourceibias.n159 gnd 0.011489f
C5699 commonsourceibias.n160 gnd 0.009605f
C5700 commonsourceibias.t164 gnd 0.17946f
C5701 commonsourceibias.n161 gnd 0.071604f
C5702 commonsourceibias.t111 gnd 0.17946f
C5703 commonsourceibias.n162 gnd 0.008208f
C5704 commonsourceibias.n163 gnd 0.009605f
C5705 commonsourceibias.t100 gnd 0.17946f
C5706 commonsourceibias.n164 gnd 0.011208f
C5707 commonsourceibias.t140 gnd 0.199526f
C5708 commonsourceibias.t84 gnd 0.17946f
C5709 commonsourceibias.n165 gnd 0.078221f
C5710 commonsourceibias.n166 gnd 0.085838f
C5711 commonsourceibias.n167 gnd 0.03983f
C5712 commonsourceibias.n168 gnd 0.009605f
C5713 commonsourceibias.n169 gnd 0.009349f
C5714 commonsourceibias.n170 gnd 0.013398f
C5715 commonsourceibias.n171 gnd 0.071604f
C5716 commonsourceibias.n172 gnd 0.013389f
C5717 commonsourceibias.n173 gnd 0.009605f
C5718 commonsourceibias.n174 gnd 0.009605f
C5719 commonsourceibias.n175 gnd 0.009605f
C5720 commonsourceibias.n176 gnd 0.012358f
C5721 commonsourceibias.n177 gnd 0.071604f
C5722 commonsourceibias.n178 gnd 0.012648f
C5723 commonsourceibias.n179 gnd 0.012288f
C5724 commonsourceibias.n180 gnd 0.009605f
C5725 commonsourceibias.n181 gnd 0.009605f
C5726 commonsourceibias.n182 gnd 0.009605f
C5727 commonsourceibias.n183 gnd 0.009057f
C5728 commonsourceibias.n184 gnd 0.01341f
C5729 commonsourceibias.n185 gnd 0.071604f
C5730 commonsourceibias.n186 gnd 0.013406f
C5731 commonsourceibias.n187 gnd 0.009605f
C5732 commonsourceibias.n188 gnd 0.009605f
C5733 commonsourceibias.n189 gnd 0.009605f
C5734 commonsourceibias.n190 gnd 0.012174f
C5735 commonsourceibias.n191 gnd 0.071604f
C5736 commonsourceibias.n192 gnd 0.012558f
C5737 commonsourceibias.n193 gnd 0.012378f
C5738 commonsourceibias.n194 gnd 0.009605f
C5739 commonsourceibias.n195 gnd 0.009605f
C5740 commonsourceibias.n196 gnd 0.011742f
C5741 commonsourceibias.n197 gnd 0.008798f
C5742 commonsourceibias.n198 gnd 0.013415f
C5743 commonsourceibias.n199 gnd 0.009605f
C5744 commonsourceibias.n200 gnd 0.009605f
C5745 commonsourceibias.n201 gnd 0.013414f
C5746 commonsourceibias.n202 gnd 0.008571f
C5747 commonsourceibias.n203 gnd 0.01197f
C5748 commonsourceibias.n204 gnd 0.009605f
C5749 commonsourceibias.n205 gnd 0.008391f
C5750 commonsourceibias.n206 gnd 0.012468f
C5751 commonsourceibias.n207 gnd 0.012468f
C5752 commonsourceibias.n208 gnd 0.008391f
C5753 commonsourceibias.n209 gnd 0.009605f
C5754 commonsourceibias.n210 gnd 0.009605f
C5755 commonsourceibias.n211 gnd 0.008571f
C5756 commonsourceibias.n212 gnd 0.013414f
C5757 commonsourceibias.n213 gnd 0.071604f
C5758 commonsourceibias.n214 gnd 0.013415f
C5759 commonsourceibias.n215 gnd 0.009605f
C5760 commonsourceibias.n216 gnd 0.009605f
C5761 commonsourceibias.n217 gnd 0.009605f
C5762 commonsourceibias.n218 gnd 0.011742f
C5763 commonsourceibias.n219 gnd 0.071604f
C5764 commonsourceibias.n220 gnd 0.012378f
C5765 commonsourceibias.n221 gnd 0.012558f
C5766 commonsourceibias.n222 gnd 0.009605f
C5767 commonsourceibias.n223 gnd 0.009605f
C5768 commonsourceibias.n224 gnd 0.009605f
C5769 commonsourceibias.n225 gnd 0.008375f
C5770 commonsourceibias.n226 gnd 0.013406f
C5771 commonsourceibias.n227 gnd 0.071604f
C5772 commonsourceibias.n228 gnd 0.01341f
C5773 commonsourceibias.n229 gnd 0.009605f
C5774 commonsourceibias.n230 gnd 0.009605f
C5775 commonsourceibias.n231 gnd 0.009605f
C5776 commonsourceibias.n232 gnd 0.011489f
C5777 commonsourceibias.n233 gnd 0.071604f
C5778 commonsourceibias.n234 gnd 0.012288f
C5779 commonsourceibias.n235 gnd 0.012648f
C5780 commonsourceibias.n236 gnd 0.009605f
C5781 commonsourceibias.n237 gnd 0.009605f
C5782 commonsourceibias.n238 gnd 0.009605f
C5783 commonsourceibias.n239 gnd 0.008208f
C5784 commonsourceibias.n240 gnd 0.013389f
C5785 commonsourceibias.n241 gnd 0.071604f
C5786 commonsourceibias.n242 gnd 0.013398f
C5787 commonsourceibias.n243 gnd 0.009605f
C5788 commonsourceibias.n244 gnd 0.009605f
C5789 commonsourceibias.n245 gnd 0.009605f
C5790 commonsourceibias.n246 gnd 0.011208f
C5791 commonsourceibias.n247 gnd 0.071604f
C5792 commonsourceibias.n248 gnd 0.011785f
C5793 commonsourceibias.n249 gnd 0.085919f
C5794 commonsourceibias.n250 gnd 0.056156f
C5795 commonsourceibias.n251 gnd 0.012817f
C5796 commonsourceibias.t88 gnd 0.194086f
C5797 commonsourceibias.t198 gnd 0.17946f
C5798 commonsourceibias.n252 gnd 0.009349f
C5799 commonsourceibias.n253 gnd 0.009605f
C5800 commonsourceibias.t186 gnd 0.17946f
C5801 commonsourceibias.n254 gnd 0.012358f
C5802 commonsourceibias.n255 gnd 0.009605f
C5803 commonsourceibias.t95 gnd 0.17946f
C5804 commonsourceibias.n256 gnd 0.071604f
C5805 commonsourceibias.t196 gnd 0.17946f
C5806 commonsourceibias.n257 gnd 0.009057f
C5807 commonsourceibias.n258 gnd 0.009605f
C5808 commonsourceibias.t105 gnd 0.17946f
C5809 commonsourceibias.n259 gnd 0.012174f
C5810 commonsourceibias.n260 gnd 0.009605f
C5811 commonsourceibias.t94 gnd 0.17946f
C5812 commonsourceibias.n261 gnd 0.071604f
C5813 commonsourceibias.t197 gnd 0.17946f
C5814 commonsourceibias.n262 gnd 0.008798f
C5815 commonsourceibias.n263 gnd 0.009605f
C5816 commonsourceibias.t115 gnd 0.17946f
C5817 commonsourceibias.n264 gnd 0.01197f
C5818 commonsourceibias.n265 gnd 0.009605f
C5819 commonsourceibias.t141 gnd 0.17946f
C5820 commonsourceibias.n266 gnd 0.071604f
C5821 commonsourceibias.t195 gnd 0.17946f
C5822 commonsourceibias.n267 gnd 0.008571f
C5823 commonsourceibias.n268 gnd 0.009605f
C5824 commonsourceibias.t113 gnd 0.17946f
C5825 commonsourceibias.n269 gnd 0.011742f
C5826 commonsourceibias.n270 gnd 0.009605f
C5827 commonsourceibias.t138 gnd 0.17946f
C5828 commonsourceibias.n271 gnd 0.071604f
C5829 commonsourceibias.t130 gnd 0.17946f
C5830 commonsourceibias.n272 gnd 0.008375f
C5831 commonsourceibias.n273 gnd 0.009605f
C5832 commonsourceibias.t114 gnd 0.17946f
C5833 commonsourceibias.n274 gnd 0.011489f
C5834 commonsourceibias.n275 gnd 0.009605f
C5835 commonsourceibias.t139 gnd 0.17946f
C5836 commonsourceibias.n276 gnd 0.071604f
C5837 commonsourceibias.t129 gnd 0.17946f
C5838 commonsourceibias.n277 gnd 0.008208f
C5839 commonsourceibias.n278 gnd 0.009605f
C5840 commonsourceibias.t125 gnd 0.17946f
C5841 commonsourceibias.n279 gnd 0.011208f
C5842 commonsourceibias.t134 gnd 0.199526f
C5843 commonsourceibias.t147 gnd 0.17946f
C5844 commonsourceibias.n280 gnd 0.078221f
C5845 commonsourceibias.n281 gnd 0.085838f
C5846 commonsourceibias.n282 gnd 0.03983f
C5847 commonsourceibias.n283 gnd 0.009605f
C5848 commonsourceibias.n284 gnd 0.009349f
C5849 commonsourceibias.n285 gnd 0.013398f
C5850 commonsourceibias.n286 gnd 0.071604f
C5851 commonsourceibias.n287 gnd 0.013389f
C5852 commonsourceibias.n288 gnd 0.009605f
C5853 commonsourceibias.n289 gnd 0.009605f
C5854 commonsourceibias.n290 gnd 0.009605f
C5855 commonsourceibias.n291 gnd 0.012358f
C5856 commonsourceibias.n292 gnd 0.071604f
C5857 commonsourceibias.n293 gnd 0.012648f
C5858 commonsourceibias.n294 gnd 0.012288f
C5859 commonsourceibias.n295 gnd 0.009605f
C5860 commonsourceibias.n296 gnd 0.009605f
C5861 commonsourceibias.n297 gnd 0.009605f
C5862 commonsourceibias.n298 gnd 0.009057f
C5863 commonsourceibias.n299 gnd 0.01341f
C5864 commonsourceibias.n300 gnd 0.071604f
C5865 commonsourceibias.n301 gnd 0.013406f
C5866 commonsourceibias.n302 gnd 0.009605f
C5867 commonsourceibias.n303 gnd 0.009605f
C5868 commonsourceibias.n304 gnd 0.009605f
C5869 commonsourceibias.n305 gnd 0.012174f
C5870 commonsourceibias.n306 gnd 0.071604f
C5871 commonsourceibias.n307 gnd 0.012558f
C5872 commonsourceibias.n308 gnd 0.012378f
C5873 commonsourceibias.n309 gnd 0.009605f
C5874 commonsourceibias.n310 gnd 0.009605f
C5875 commonsourceibias.n311 gnd 0.009605f
C5876 commonsourceibias.n312 gnd 0.008798f
C5877 commonsourceibias.n313 gnd 0.013415f
C5878 commonsourceibias.n314 gnd 0.071604f
C5879 commonsourceibias.n315 gnd 0.013414f
C5880 commonsourceibias.n316 gnd 0.009605f
C5881 commonsourceibias.n317 gnd 0.009605f
C5882 commonsourceibias.n318 gnd 0.009605f
C5883 commonsourceibias.n319 gnd 0.01197f
C5884 commonsourceibias.n320 gnd 0.071604f
C5885 commonsourceibias.n321 gnd 0.012468f
C5886 commonsourceibias.n322 gnd 0.012468f
C5887 commonsourceibias.n323 gnd 0.009605f
C5888 commonsourceibias.n324 gnd 0.009605f
C5889 commonsourceibias.n325 gnd 0.009605f
C5890 commonsourceibias.n326 gnd 0.008571f
C5891 commonsourceibias.n327 gnd 0.013414f
C5892 commonsourceibias.n328 gnd 0.071604f
C5893 commonsourceibias.n329 gnd 0.013415f
C5894 commonsourceibias.n330 gnd 0.009605f
C5895 commonsourceibias.n331 gnd 0.009605f
C5896 commonsourceibias.n332 gnd 0.009605f
C5897 commonsourceibias.n333 gnd 0.011742f
C5898 commonsourceibias.n334 gnd 0.071604f
C5899 commonsourceibias.n335 gnd 0.012378f
C5900 commonsourceibias.n336 gnd 0.012558f
C5901 commonsourceibias.n337 gnd 0.009605f
C5902 commonsourceibias.n338 gnd 0.009605f
C5903 commonsourceibias.n339 gnd 0.009605f
C5904 commonsourceibias.n340 gnd 0.008375f
C5905 commonsourceibias.n341 gnd 0.013406f
C5906 commonsourceibias.n342 gnd 0.071604f
C5907 commonsourceibias.n343 gnd 0.01341f
C5908 commonsourceibias.n344 gnd 0.009605f
C5909 commonsourceibias.n345 gnd 0.009605f
C5910 commonsourceibias.n346 gnd 0.009605f
C5911 commonsourceibias.n347 gnd 0.011489f
C5912 commonsourceibias.n348 gnd 0.071604f
C5913 commonsourceibias.n349 gnd 0.012288f
C5914 commonsourceibias.n350 gnd 0.012648f
C5915 commonsourceibias.n351 gnd 0.009605f
C5916 commonsourceibias.n352 gnd 0.009605f
C5917 commonsourceibias.n353 gnd 0.009605f
C5918 commonsourceibias.n354 gnd 0.008208f
C5919 commonsourceibias.n355 gnd 0.013389f
C5920 commonsourceibias.n356 gnd 0.071604f
C5921 commonsourceibias.n357 gnd 0.013398f
C5922 commonsourceibias.n358 gnd 0.009605f
C5923 commonsourceibias.n359 gnd 0.009605f
C5924 commonsourceibias.n360 gnd 0.009605f
C5925 commonsourceibias.n361 gnd 0.011208f
C5926 commonsourceibias.n362 gnd 0.071604f
C5927 commonsourceibias.n363 gnd 0.011785f
C5928 commonsourceibias.n364 gnd 0.085919f
C5929 commonsourceibias.n365 gnd 0.029883f
C5930 commonsourceibias.n366 gnd 0.153509f
C5931 commonsourceibias.n367 gnd 0.012817f
C5932 commonsourceibias.t92 gnd 0.17946f
C5933 commonsourceibias.n368 gnd 0.009349f
C5934 commonsourceibias.n369 gnd 0.009605f
C5935 commonsourceibias.t163 gnd 0.17946f
C5936 commonsourceibias.n370 gnd 0.012358f
C5937 commonsourceibias.n371 gnd 0.009605f
C5938 commonsourceibias.t157 gnd 0.17946f
C5939 commonsourceibias.n372 gnd 0.071604f
C5940 commonsourceibias.t194 gnd 0.17946f
C5941 commonsourceibias.n373 gnd 0.009057f
C5942 commonsourceibias.n374 gnd 0.009605f
C5943 commonsourceibias.t110 gnd 0.17946f
C5944 commonsourceibias.n375 gnd 0.012174f
C5945 commonsourceibias.n376 gnd 0.009605f
C5946 commonsourceibias.t149 gnd 0.17946f
C5947 commonsourceibias.n377 gnd 0.071604f
C5948 commonsourceibias.t182 gnd 0.17946f
C5949 commonsourceibias.n378 gnd 0.008798f
C5950 commonsourceibias.n379 gnd 0.009605f
C5951 commonsourceibias.t173 gnd 0.17946f
C5952 commonsourceibias.n380 gnd 0.01197f
C5953 commonsourceibias.n381 gnd 0.009605f
C5954 commonsourceibias.t80 gnd 0.17946f
C5955 commonsourceibias.n382 gnd 0.071604f
C5956 commonsourceibias.t172 gnd 0.17946f
C5957 commonsourceibias.n383 gnd 0.008571f
C5958 commonsourceibias.n384 gnd 0.009605f
C5959 commonsourceibias.t168 gnd 0.17946f
C5960 commonsourceibias.n385 gnd 0.011742f
C5961 commonsourceibias.n386 gnd 0.009605f
C5962 commonsourceibias.t187 gnd 0.17946f
C5963 commonsourceibias.n387 gnd 0.071604f
C5964 commonsourceibias.t96 gnd 0.17946f
C5965 commonsourceibias.n388 gnd 0.008375f
C5966 commonsourceibias.n389 gnd 0.009605f
C5967 commonsourceibias.t165 gnd 0.17946f
C5968 commonsourceibias.n390 gnd 0.011489f
C5969 commonsourceibias.n391 gnd 0.009605f
C5970 commonsourceibias.t175 gnd 0.17946f
C5971 commonsourceibias.n392 gnd 0.071604f
C5972 commonsourceibias.t199 gnd 0.17946f
C5973 commonsourceibias.n393 gnd 0.008208f
C5974 commonsourceibias.n394 gnd 0.009605f
C5975 commonsourceibias.t155 gnd 0.17946f
C5976 commonsourceibias.n395 gnd 0.011208f
C5977 commonsourceibias.t184 gnd 0.199526f
C5978 commonsourceibias.t150 gnd 0.17946f
C5979 commonsourceibias.n396 gnd 0.078221f
C5980 commonsourceibias.n397 gnd 0.085838f
C5981 commonsourceibias.n398 gnd 0.03983f
C5982 commonsourceibias.n399 gnd 0.009605f
C5983 commonsourceibias.n400 gnd 0.009349f
C5984 commonsourceibias.n401 gnd 0.013398f
C5985 commonsourceibias.n402 gnd 0.071604f
C5986 commonsourceibias.n403 gnd 0.013389f
C5987 commonsourceibias.n404 gnd 0.009605f
C5988 commonsourceibias.n405 gnd 0.009605f
C5989 commonsourceibias.n406 gnd 0.009605f
C5990 commonsourceibias.n407 gnd 0.012358f
C5991 commonsourceibias.n408 gnd 0.071604f
C5992 commonsourceibias.n409 gnd 0.012648f
C5993 commonsourceibias.n410 gnd 0.012288f
C5994 commonsourceibias.n411 gnd 0.009605f
C5995 commonsourceibias.n412 gnd 0.009605f
C5996 commonsourceibias.n413 gnd 0.009605f
C5997 commonsourceibias.n414 gnd 0.009057f
C5998 commonsourceibias.n415 gnd 0.01341f
C5999 commonsourceibias.n416 gnd 0.071604f
C6000 commonsourceibias.n417 gnd 0.013406f
C6001 commonsourceibias.n418 gnd 0.009605f
C6002 commonsourceibias.n419 gnd 0.009605f
C6003 commonsourceibias.n420 gnd 0.009605f
C6004 commonsourceibias.n421 gnd 0.012174f
C6005 commonsourceibias.n422 gnd 0.071604f
C6006 commonsourceibias.n423 gnd 0.012558f
C6007 commonsourceibias.n424 gnd 0.012378f
C6008 commonsourceibias.n425 gnd 0.009605f
C6009 commonsourceibias.n426 gnd 0.009605f
C6010 commonsourceibias.n427 gnd 0.009605f
C6011 commonsourceibias.n428 gnd 0.008798f
C6012 commonsourceibias.n429 gnd 0.013415f
C6013 commonsourceibias.n430 gnd 0.071604f
C6014 commonsourceibias.n431 gnd 0.013414f
C6015 commonsourceibias.n432 gnd 0.009605f
C6016 commonsourceibias.n433 gnd 0.009605f
C6017 commonsourceibias.n434 gnd 0.009605f
C6018 commonsourceibias.n435 gnd 0.01197f
C6019 commonsourceibias.n436 gnd 0.071604f
C6020 commonsourceibias.n437 gnd 0.012468f
C6021 commonsourceibias.n438 gnd 0.012468f
C6022 commonsourceibias.n439 gnd 0.009605f
C6023 commonsourceibias.n440 gnd 0.009605f
C6024 commonsourceibias.n441 gnd 0.009605f
C6025 commonsourceibias.n442 gnd 0.008571f
C6026 commonsourceibias.n443 gnd 0.013414f
C6027 commonsourceibias.n444 gnd 0.071604f
C6028 commonsourceibias.n445 gnd 0.013415f
C6029 commonsourceibias.n446 gnd 0.009605f
C6030 commonsourceibias.n447 gnd 0.009605f
C6031 commonsourceibias.n448 gnd 0.009605f
C6032 commonsourceibias.n449 gnd 0.011742f
C6033 commonsourceibias.n450 gnd 0.071604f
C6034 commonsourceibias.n451 gnd 0.012378f
C6035 commonsourceibias.n452 gnd 0.012558f
C6036 commonsourceibias.n453 gnd 0.009605f
C6037 commonsourceibias.n454 gnd 0.009605f
C6038 commonsourceibias.n455 gnd 0.009605f
C6039 commonsourceibias.n456 gnd 0.008375f
C6040 commonsourceibias.n457 gnd 0.013406f
C6041 commonsourceibias.n458 gnd 0.071604f
C6042 commonsourceibias.n459 gnd 0.01341f
C6043 commonsourceibias.n460 gnd 0.009605f
C6044 commonsourceibias.n461 gnd 0.009605f
C6045 commonsourceibias.n462 gnd 0.009605f
C6046 commonsourceibias.n463 gnd 0.011489f
C6047 commonsourceibias.n464 gnd 0.071604f
C6048 commonsourceibias.n465 gnd 0.012288f
C6049 commonsourceibias.n466 gnd 0.012648f
C6050 commonsourceibias.n467 gnd 0.009605f
C6051 commonsourceibias.n468 gnd 0.009605f
C6052 commonsourceibias.n469 gnd 0.009605f
C6053 commonsourceibias.n470 gnd 0.008208f
C6054 commonsourceibias.n471 gnd 0.013389f
C6055 commonsourceibias.n472 gnd 0.071604f
C6056 commonsourceibias.n473 gnd 0.013398f
C6057 commonsourceibias.n474 gnd 0.009605f
C6058 commonsourceibias.n475 gnd 0.009605f
C6059 commonsourceibias.n476 gnd 0.009605f
C6060 commonsourceibias.n477 gnd 0.011208f
C6061 commonsourceibias.n478 gnd 0.071604f
C6062 commonsourceibias.n479 gnd 0.011785f
C6063 commonsourceibias.t183 gnd 0.194086f
C6064 commonsourceibias.n480 gnd 0.085919f
C6065 commonsourceibias.n481 gnd 0.029883f
C6066 commonsourceibias.n482 gnd 0.456424f
C6067 commonsourceibias.n483 gnd 0.012817f
C6068 commonsourceibias.t112 gnd 0.194086f
C6069 commonsourceibias.t169 gnd 0.17946f
C6070 commonsourceibias.n484 gnd 0.009349f
C6071 commonsourceibias.n485 gnd 0.009605f
C6072 commonsourceibias.t142 gnd 0.17946f
C6073 commonsourceibias.n486 gnd 0.012358f
C6074 commonsourceibias.n487 gnd 0.009605f
C6075 commonsourceibias.t154 gnd 0.17946f
C6076 commonsourceibias.n488 gnd 0.009057f
C6077 commonsourceibias.n489 gnd 0.009605f
C6078 commonsourceibias.t108 gnd 0.17946f
C6079 commonsourceibias.n490 gnd 0.012174f
C6080 commonsourceibias.n491 gnd 0.009605f
C6081 commonsourceibias.t128 gnd 0.17946f
C6082 commonsourceibias.n492 gnd 0.008798f
C6083 commonsourceibias.n493 gnd 0.009605f
C6084 commonsourceibias.t109 gnd 0.17946f
C6085 commonsourceibias.n494 gnd 0.01197f
C6086 commonsourceibias.t5 gnd 0.020728f
C6087 commonsourceibias.t71 gnd 0.020728f
C6088 commonsourceibias.n495 gnd 0.18377f
C6089 commonsourceibias.t69 gnd 0.020728f
C6090 commonsourceibias.t15 gnd 0.020728f
C6091 commonsourceibias.n496 gnd 0.183157f
C6092 commonsourceibias.n497 gnd 0.170668f
C6093 commonsourceibias.t37 gnd 0.020728f
C6094 commonsourceibias.t79 gnd 0.020728f
C6095 commonsourceibias.n498 gnd 0.183157f
C6096 commonsourceibias.n499 gnd 0.084131f
C6097 commonsourceibias.t29 gnd 0.020728f
C6098 commonsourceibias.t65 gnd 0.020728f
C6099 commonsourceibias.n500 gnd 0.183157f
C6100 commonsourceibias.n501 gnd 0.084131f
C6101 commonsourceibias.t13 gnd 0.020728f
C6102 commonsourceibias.t31 gnd 0.020728f
C6103 commonsourceibias.n502 gnd 0.183157f
C6104 commonsourceibias.n503 gnd 0.070287f
C6105 commonsourceibias.n504 gnd 0.012817f
C6106 commonsourceibias.t2 gnd 0.17946f
C6107 commonsourceibias.n505 gnd 0.009349f
C6108 commonsourceibias.n506 gnd 0.009605f
C6109 commonsourceibias.t60 gnd 0.17946f
C6110 commonsourceibias.n507 gnd 0.012358f
C6111 commonsourceibias.n508 gnd 0.009605f
C6112 commonsourceibias.t74 gnd 0.17946f
C6113 commonsourceibias.n509 gnd 0.009057f
C6114 commonsourceibias.n510 gnd 0.009605f
C6115 commonsourceibias.t26 gnd 0.17946f
C6116 commonsourceibias.n511 gnd 0.012174f
C6117 commonsourceibias.n512 gnd 0.009605f
C6118 commonsourceibias.t40 gnd 0.17946f
C6119 commonsourceibias.n513 gnd 0.008798f
C6120 commonsourceibias.n514 gnd 0.009605f
C6121 commonsourceibias.t24 gnd 0.17946f
C6122 commonsourceibias.n515 gnd 0.01197f
C6123 commonsourceibias.n516 gnd 0.009605f
C6124 commonsourceibias.t30 gnd 0.17946f
C6125 commonsourceibias.n517 gnd 0.008571f
C6126 commonsourceibias.n518 gnd 0.009605f
C6127 commonsourceibias.t12 gnd 0.17946f
C6128 commonsourceibias.n519 gnd 0.011742f
C6129 commonsourceibias.n520 gnd 0.009605f
C6130 commonsourceibias.t28 gnd 0.17946f
C6131 commonsourceibias.n521 gnd 0.008375f
C6132 commonsourceibias.n522 gnd 0.009605f
C6133 commonsourceibias.t78 gnd 0.17946f
C6134 commonsourceibias.n523 gnd 0.011489f
C6135 commonsourceibias.n524 gnd 0.009605f
C6136 commonsourceibias.t14 gnd 0.17946f
C6137 commonsourceibias.n525 gnd 0.008208f
C6138 commonsourceibias.n526 gnd 0.009605f
C6139 commonsourceibias.t68 gnd 0.17946f
C6140 commonsourceibias.n527 gnd 0.011208f
C6141 commonsourceibias.t4 gnd 0.199526f
C6142 commonsourceibias.t70 gnd 0.17946f
C6143 commonsourceibias.n528 gnd 0.078221f
C6144 commonsourceibias.n529 gnd 0.085838f
C6145 commonsourceibias.n530 gnd 0.03983f
C6146 commonsourceibias.n531 gnd 0.009605f
C6147 commonsourceibias.n532 gnd 0.009349f
C6148 commonsourceibias.n533 gnd 0.013398f
C6149 commonsourceibias.n534 gnd 0.071604f
C6150 commonsourceibias.n535 gnd 0.013389f
C6151 commonsourceibias.n536 gnd 0.009605f
C6152 commonsourceibias.n537 gnd 0.009605f
C6153 commonsourceibias.n538 gnd 0.009605f
C6154 commonsourceibias.n539 gnd 0.012358f
C6155 commonsourceibias.n540 gnd 0.071604f
C6156 commonsourceibias.n541 gnd 0.012648f
C6157 commonsourceibias.t36 gnd 0.17946f
C6158 commonsourceibias.n542 gnd 0.071604f
C6159 commonsourceibias.n543 gnd 0.012288f
C6160 commonsourceibias.n544 gnd 0.009605f
C6161 commonsourceibias.n545 gnd 0.009605f
C6162 commonsourceibias.n546 gnd 0.009605f
C6163 commonsourceibias.n547 gnd 0.009057f
C6164 commonsourceibias.n548 gnd 0.01341f
C6165 commonsourceibias.n549 gnd 0.071604f
C6166 commonsourceibias.n550 gnd 0.013406f
C6167 commonsourceibias.n551 gnd 0.009605f
C6168 commonsourceibias.n552 gnd 0.009605f
C6169 commonsourceibias.n553 gnd 0.009605f
C6170 commonsourceibias.n554 gnd 0.012174f
C6171 commonsourceibias.n555 gnd 0.071604f
C6172 commonsourceibias.n556 gnd 0.012558f
C6173 commonsourceibias.t64 gnd 0.17946f
C6174 commonsourceibias.n557 gnd 0.071604f
C6175 commonsourceibias.n558 gnd 0.012378f
C6176 commonsourceibias.n559 gnd 0.009605f
C6177 commonsourceibias.n560 gnd 0.009605f
C6178 commonsourceibias.n561 gnd 0.009605f
C6179 commonsourceibias.n562 gnd 0.008798f
C6180 commonsourceibias.n563 gnd 0.013415f
C6181 commonsourceibias.n564 gnd 0.071604f
C6182 commonsourceibias.n565 gnd 0.013414f
C6183 commonsourceibias.n566 gnd 0.009605f
C6184 commonsourceibias.n567 gnd 0.009605f
C6185 commonsourceibias.n568 gnd 0.009605f
C6186 commonsourceibias.n569 gnd 0.01197f
C6187 commonsourceibias.n570 gnd 0.071604f
C6188 commonsourceibias.n571 gnd 0.012468f
C6189 commonsourceibias.t8 gnd 0.17946f
C6190 commonsourceibias.n572 gnd 0.071604f
C6191 commonsourceibias.n573 gnd 0.012468f
C6192 commonsourceibias.n574 gnd 0.009605f
C6193 commonsourceibias.n575 gnd 0.009605f
C6194 commonsourceibias.n576 gnd 0.009605f
C6195 commonsourceibias.n577 gnd 0.008571f
C6196 commonsourceibias.n578 gnd 0.013414f
C6197 commonsourceibias.n579 gnd 0.071604f
C6198 commonsourceibias.n580 gnd 0.013415f
C6199 commonsourceibias.n581 gnd 0.009605f
C6200 commonsourceibias.n582 gnd 0.009605f
C6201 commonsourceibias.n583 gnd 0.009605f
C6202 commonsourceibias.n584 gnd 0.011742f
C6203 commonsourceibias.n585 gnd 0.071604f
C6204 commonsourceibias.n586 gnd 0.012378f
C6205 commonsourceibias.t16 gnd 0.17946f
C6206 commonsourceibias.n587 gnd 0.071604f
C6207 commonsourceibias.n588 gnd 0.012558f
C6208 commonsourceibias.n589 gnd 0.009605f
C6209 commonsourceibias.n590 gnd 0.009605f
C6210 commonsourceibias.n591 gnd 0.009605f
C6211 commonsourceibias.n592 gnd 0.008375f
C6212 commonsourceibias.n593 gnd 0.013406f
C6213 commonsourceibias.n594 gnd 0.071604f
C6214 commonsourceibias.n595 gnd 0.01341f
C6215 commonsourceibias.n596 gnd 0.009605f
C6216 commonsourceibias.n597 gnd 0.009605f
C6217 commonsourceibias.n598 gnd 0.009605f
C6218 commonsourceibias.n599 gnd 0.011489f
C6219 commonsourceibias.n600 gnd 0.071604f
C6220 commonsourceibias.n601 gnd 0.012288f
C6221 commonsourceibias.t46 gnd 0.17946f
C6222 commonsourceibias.n602 gnd 0.071604f
C6223 commonsourceibias.n603 gnd 0.012648f
C6224 commonsourceibias.n604 gnd 0.009605f
C6225 commonsourceibias.n605 gnd 0.009605f
C6226 commonsourceibias.n606 gnd 0.009605f
C6227 commonsourceibias.n607 gnd 0.008208f
C6228 commonsourceibias.n608 gnd 0.013389f
C6229 commonsourceibias.n609 gnd 0.071604f
C6230 commonsourceibias.n610 gnd 0.013398f
C6231 commonsourceibias.n611 gnd 0.009605f
C6232 commonsourceibias.n612 gnd 0.009605f
C6233 commonsourceibias.n613 gnd 0.009605f
C6234 commonsourceibias.n614 gnd 0.011208f
C6235 commonsourceibias.n615 gnd 0.071604f
C6236 commonsourceibias.n616 gnd 0.011785f
C6237 commonsourceibias.t48 gnd 0.194086f
C6238 commonsourceibias.n617 gnd 0.085919f
C6239 commonsourceibias.n618 gnd 0.095702f
C6240 commonsourceibias.t3 gnd 0.020728f
C6241 commonsourceibias.t49 gnd 0.020728f
C6242 commonsourceibias.n619 gnd 0.183157f
C6243 commonsourceibias.n620 gnd 0.158432f
C6244 commonsourceibias.t47 gnd 0.020728f
C6245 commonsourceibias.t61 gnd 0.020728f
C6246 commonsourceibias.n621 gnd 0.183157f
C6247 commonsourceibias.n622 gnd 0.084131f
C6248 commonsourceibias.t27 gnd 0.020728f
C6249 commonsourceibias.t75 gnd 0.020728f
C6250 commonsourceibias.n623 gnd 0.183157f
C6251 commonsourceibias.n624 gnd 0.084131f
C6252 commonsourceibias.t41 gnd 0.020728f
C6253 commonsourceibias.t17 gnd 0.020728f
C6254 commonsourceibias.n625 gnd 0.183157f
C6255 commonsourceibias.n626 gnd 0.084131f
C6256 commonsourceibias.t9 gnd 0.020728f
C6257 commonsourceibias.t25 gnd 0.020728f
C6258 commonsourceibias.n627 gnd 0.183157f
C6259 commonsourceibias.n628 gnd 0.070287f
C6260 commonsourceibias.n629 gnd 0.085111f
C6261 commonsourceibias.n630 gnd 0.062167f
C6262 commonsourceibias.t102 gnd 0.17946f
C6263 commonsourceibias.n631 gnd 0.071604f
C6264 commonsourceibias.n632 gnd 0.009605f
C6265 commonsourceibias.t188 gnd 0.17946f
C6266 commonsourceibias.n633 gnd 0.071604f
C6267 commonsourceibias.n634 gnd 0.009605f
C6268 commonsourceibias.t162 gnd 0.17946f
C6269 commonsourceibias.n635 gnd 0.071604f
C6270 commonsourceibias.n636 gnd 0.009605f
C6271 commonsourceibias.t103 gnd 0.17946f
C6272 commonsourceibias.n637 gnd 0.008375f
C6273 commonsourceibias.n638 gnd 0.009605f
C6274 commonsourceibias.t166 gnd 0.17946f
C6275 commonsourceibias.n639 gnd 0.011489f
C6276 commonsourceibias.n640 gnd 0.009605f
C6277 commonsourceibias.t185 gnd 0.17946f
C6278 commonsourceibias.n641 gnd 0.008208f
C6279 commonsourceibias.n642 gnd 0.009605f
C6280 commonsourceibias.t160 gnd 0.17946f
C6281 commonsourceibias.n643 gnd 0.011208f
C6282 commonsourceibias.t177 gnd 0.199526f
C6283 commonsourceibias.t159 gnd 0.17946f
C6284 commonsourceibias.n644 gnd 0.078221f
C6285 commonsourceibias.n645 gnd 0.085838f
C6286 commonsourceibias.n646 gnd 0.03983f
C6287 commonsourceibias.n647 gnd 0.009605f
C6288 commonsourceibias.n648 gnd 0.009349f
C6289 commonsourceibias.n649 gnd 0.013398f
C6290 commonsourceibias.n650 gnd 0.071604f
C6291 commonsourceibias.n651 gnd 0.013389f
C6292 commonsourceibias.n652 gnd 0.009605f
C6293 commonsourceibias.n653 gnd 0.009605f
C6294 commonsourceibias.n654 gnd 0.009605f
C6295 commonsourceibias.n655 gnd 0.012358f
C6296 commonsourceibias.n656 gnd 0.071604f
C6297 commonsourceibias.n657 gnd 0.012648f
C6298 commonsourceibias.t135 gnd 0.17946f
C6299 commonsourceibias.n658 gnd 0.071604f
C6300 commonsourceibias.n659 gnd 0.012288f
C6301 commonsourceibias.n660 gnd 0.009605f
C6302 commonsourceibias.n661 gnd 0.009605f
C6303 commonsourceibias.n662 gnd 0.009605f
C6304 commonsourceibias.n663 gnd 0.009057f
C6305 commonsourceibias.n664 gnd 0.01341f
C6306 commonsourceibias.n665 gnd 0.071604f
C6307 commonsourceibias.n666 gnd 0.013406f
C6308 commonsourceibias.n667 gnd 0.009605f
C6309 commonsourceibias.n668 gnd 0.009605f
C6310 commonsourceibias.n669 gnd 0.009605f
C6311 commonsourceibias.n670 gnd 0.012174f
C6312 commonsourceibias.n671 gnd 0.071604f
C6313 commonsourceibias.n672 gnd 0.012558f
C6314 commonsourceibias.n673 gnd 0.012378f
C6315 commonsourceibias.n674 gnd 0.009605f
C6316 commonsourceibias.n675 gnd 0.009605f
C6317 commonsourceibias.n676 gnd 0.011742f
C6318 commonsourceibias.n677 gnd 0.008798f
C6319 commonsourceibias.n678 gnd 0.013415f
C6320 commonsourceibias.n679 gnd 0.009605f
C6321 commonsourceibias.n680 gnd 0.009605f
C6322 commonsourceibias.n681 gnd 0.013414f
C6323 commonsourceibias.n682 gnd 0.008571f
C6324 commonsourceibias.n683 gnd 0.01197f
C6325 commonsourceibias.n684 gnd 0.009605f
C6326 commonsourceibias.n685 gnd 0.008391f
C6327 commonsourceibias.n686 gnd 0.012468f
C6328 commonsourceibias.t174 gnd 0.17946f
C6329 commonsourceibias.n687 gnd 0.071604f
C6330 commonsourceibias.n688 gnd 0.012468f
C6331 commonsourceibias.n689 gnd 0.008391f
C6332 commonsourceibias.n690 gnd 0.009605f
C6333 commonsourceibias.n691 gnd 0.009605f
C6334 commonsourceibias.n692 gnd 0.008571f
C6335 commonsourceibias.n693 gnd 0.013414f
C6336 commonsourceibias.n694 gnd 0.071604f
C6337 commonsourceibias.n695 gnd 0.013415f
C6338 commonsourceibias.n696 gnd 0.009605f
C6339 commonsourceibias.n697 gnd 0.009605f
C6340 commonsourceibias.n698 gnd 0.009605f
C6341 commonsourceibias.n699 gnd 0.011742f
C6342 commonsourceibias.n700 gnd 0.071604f
C6343 commonsourceibias.n701 gnd 0.012378f
C6344 commonsourceibias.t90 gnd 0.17946f
C6345 commonsourceibias.n702 gnd 0.071604f
C6346 commonsourceibias.n703 gnd 0.012558f
C6347 commonsourceibias.n704 gnd 0.009605f
C6348 commonsourceibias.n705 gnd 0.009605f
C6349 commonsourceibias.n706 gnd 0.009605f
C6350 commonsourceibias.n707 gnd 0.008375f
C6351 commonsourceibias.n708 gnd 0.013406f
C6352 commonsourceibias.n709 gnd 0.071604f
C6353 commonsourceibias.n710 gnd 0.01341f
C6354 commonsourceibias.n711 gnd 0.009605f
C6355 commonsourceibias.n712 gnd 0.009605f
C6356 commonsourceibias.n713 gnd 0.009605f
C6357 commonsourceibias.n714 gnd 0.011489f
C6358 commonsourceibias.n715 gnd 0.071604f
C6359 commonsourceibias.n716 gnd 0.012288f
C6360 commonsourceibias.t116 gnd 0.17946f
C6361 commonsourceibias.n717 gnd 0.071604f
C6362 commonsourceibias.n718 gnd 0.012648f
C6363 commonsourceibias.n719 gnd 0.009605f
C6364 commonsourceibias.n720 gnd 0.009605f
C6365 commonsourceibias.n721 gnd 0.009605f
C6366 commonsourceibias.n722 gnd 0.008208f
C6367 commonsourceibias.n723 gnd 0.013389f
C6368 commonsourceibias.n724 gnd 0.071604f
C6369 commonsourceibias.n725 gnd 0.013398f
C6370 commonsourceibias.n726 gnd 0.009605f
C6371 commonsourceibias.n727 gnd 0.009605f
C6372 commonsourceibias.n728 gnd 0.009605f
C6373 commonsourceibias.n729 gnd 0.011208f
C6374 commonsourceibias.n730 gnd 0.071604f
C6375 commonsourceibias.n731 gnd 0.011785f
C6376 commonsourceibias.n732 gnd 0.085919f
C6377 commonsourceibias.n733 gnd 0.056156f
C6378 commonsourceibias.n734 gnd 0.012817f
C6379 commonsourceibias.t180 gnd 0.17946f
C6380 commonsourceibias.n735 gnd 0.009349f
C6381 commonsourceibias.n736 gnd 0.009605f
C6382 commonsourceibias.t82 gnd 0.17946f
C6383 commonsourceibias.n737 gnd 0.012358f
C6384 commonsourceibias.n738 gnd 0.009605f
C6385 commonsourceibias.t179 gnd 0.17946f
C6386 commonsourceibias.n739 gnd 0.009057f
C6387 commonsourceibias.n740 gnd 0.009605f
C6388 commonsourceibias.t81 gnd 0.17946f
C6389 commonsourceibias.n741 gnd 0.012174f
C6390 commonsourceibias.n742 gnd 0.009605f
C6391 commonsourceibias.t178 gnd 0.17946f
C6392 commonsourceibias.n743 gnd 0.008798f
C6393 commonsourceibias.n744 gnd 0.009605f
C6394 commonsourceibias.t89 gnd 0.17946f
C6395 commonsourceibias.n745 gnd 0.01197f
C6396 commonsourceibias.n746 gnd 0.009605f
C6397 commonsourceibias.t97 gnd 0.17946f
C6398 commonsourceibias.n747 gnd 0.008571f
C6399 commonsourceibias.n748 gnd 0.009605f
C6400 commonsourceibias.t86 gnd 0.17946f
C6401 commonsourceibias.n749 gnd 0.011742f
C6402 commonsourceibias.n750 gnd 0.009605f
C6403 commonsourceibias.t106 gnd 0.17946f
C6404 commonsourceibias.n751 gnd 0.008375f
C6405 commonsourceibias.n752 gnd 0.009605f
C6406 commonsourceibias.t85 gnd 0.17946f
C6407 commonsourceibias.n753 gnd 0.011489f
C6408 commonsourceibias.n754 gnd 0.009605f
C6409 commonsourceibias.t104 gnd 0.17946f
C6410 commonsourceibias.n755 gnd 0.008208f
C6411 commonsourceibias.n756 gnd 0.009605f
C6412 commonsourceibias.t132 gnd 0.17946f
C6413 commonsourceibias.n757 gnd 0.011208f
C6414 commonsourceibias.t98 gnd 0.199526f
C6415 commonsourceibias.t123 gnd 0.17946f
C6416 commonsourceibias.n758 gnd 0.078221f
C6417 commonsourceibias.n759 gnd 0.085838f
C6418 commonsourceibias.n760 gnd 0.03983f
C6419 commonsourceibias.n761 gnd 0.009605f
C6420 commonsourceibias.n762 gnd 0.009349f
C6421 commonsourceibias.n763 gnd 0.013398f
C6422 commonsourceibias.n764 gnd 0.071604f
C6423 commonsourceibias.n765 gnd 0.013389f
C6424 commonsourceibias.n766 gnd 0.009605f
C6425 commonsourceibias.n767 gnd 0.009605f
C6426 commonsourceibias.n768 gnd 0.009605f
C6427 commonsourceibias.n769 gnd 0.012358f
C6428 commonsourceibias.n770 gnd 0.071604f
C6429 commonsourceibias.n771 gnd 0.012648f
C6430 commonsourceibias.t118 gnd 0.17946f
C6431 commonsourceibias.n772 gnd 0.071604f
C6432 commonsourceibias.n773 gnd 0.012288f
C6433 commonsourceibias.n774 gnd 0.009605f
C6434 commonsourceibias.n775 gnd 0.009605f
C6435 commonsourceibias.n776 gnd 0.009605f
C6436 commonsourceibias.n777 gnd 0.009057f
C6437 commonsourceibias.n778 gnd 0.01341f
C6438 commonsourceibias.n779 gnd 0.071604f
C6439 commonsourceibias.n780 gnd 0.013406f
C6440 commonsourceibias.n781 gnd 0.009605f
C6441 commonsourceibias.n782 gnd 0.009605f
C6442 commonsourceibias.n783 gnd 0.009605f
C6443 commonsourceibias.n784 gnd 0.012174f
C6444 commonsourceibias.n785 gnd 0.071604f
C6445 commonsourceibias.n786 gnd 0.012558f
C6446 commonsourceibias.t119 gnd 0.17946f
C6447 commonsourceibias.n787 gnd 0.071604f
C6448 commonsourceibias.n788 gnd 0.012378f
C6449 commonsourceibias.n789 gnd 0.009605f
C6450 commonsourceibias.n790 gnd 0.009605f
C6451 commonsourceibias.n791 gnd 0.009605f
C6452 commonsourceibias.n792 gnd 0.008798f
C6453 commonsourceibias.n793 gnd 0.013415f
C6454 commonsourceibias.n794 gnd 0.071604f
C6455 commonsourceibias.n795 gnd 0.013414f
C6456 commonsourceibias.n796 gnd 0.009605f
C6457 commonsourceibias.n797 gnd 0.009605f
C6458 commonsourceibias.n798 gnd 0.009605f
C6459 commonsourceibias.n799 gnd 0.01197f
C6460 commonsourceibias.n800 gnd 0.071604f
C6461 commonsourceibias.n801 gnd 0.012468f
C6462 commonsourceibias.t120 gnd 0.17946f
C6463 commonsourceibias.n802 gnd 0.071604f
C6464 commonsourceibias.n803 gnd 0.012468f
C6465 commonsourceibias.n804 gnd 0.009605f
C6466 commonsourceibias.n805 gnd 0.009605f
C6467 commonsourceibias.n806 gnd 0.009605f
C6468 commonsourceibias.n807 gnd 0.008571f
C6469 commonsourceibias.n808 gnd 0.013414f
C6470 commonsourceibias.n809 gnd 0.071604f
C6471 commonsourceibias.n810 gnd 0.013415f
C6472 commonsourceibias.n811 gnd 0.009605f
C6473 commonsourceibias.n812 gnd 0.009605f
C6474 commonsourceibias.n813 gnd 0.009605f
C6475 commonsourceibias.n814 gnd 0.011742f
C6476 commonsourceibias.n815 gnd 0.071604f
C6477 commonsourceibias.n816 gnd 0.012378f
C6478 commonsourceibias.t121 gnd 0.17946f
C6479 commonsourceibias.n817 gnd 0.071604f
C6480 commonsourceibias.n818 gnd 0.012558f
C6481 commonsourceibias.n819 gnd 0.009605f
C6482 commonsourceibias.n820 gnd 0.009605f
C6483 commonsourceibias.n821 gnd 0.009605f
C6484 commonsourceibias.n822 gnd 0.008375f
C6485 commonsourceibias.n823 gnd 0.013406f
C6486 commonsourceibias.n824 gnd 0.071604f
C6487 commonsourceibias.n825 gnd 0.01341f
C6488 commonsourceibias.n826 gnd 0.009605f
C6489 commonsourceibias.n827 gnd 0.009605f
C6490 commonsourceibias.n828 gnd 0.009605f
C6491 commonsourceibias.n829 gnd 0.011489f
C6492 commonsourceibias.n830 gnd 0.071604f
C6493 commonsourceibias.n831 gnd 0.012288f
C6494 commonsourceibias.t193 gnd 0.17946f
C6495 commonsourceibias.n832 gnd 0.071604f
C6496 commonsourceibias.n833 gnd 0.012648f
C6497 commonsourceibias.n834 gnd 0.009605f
C6498 commonsourceibias.n835 gnd 0.009605f
C6499 commonsourceibias.n836 gnd 0.009605f
C6500 commonsourceibias.n837 gnd 0.008208f
C6501 commonsourceibias.n838 gnd 0.013389f
C6502 commonsourceibias.n839 gnd 0.071604f
C6503 commonsourceibias.n840 gnd 0.013398f
C6504 commonsourceibias.n841 gnd 0.009605f
C6505 commonsourceibias.n842 gnd 0.009605f
C6506 commonsourceibias.n843 gnd 0.009605f
C6507 commonsourceibias.n844 gnd 0.011208f
C6508 commonsourceibias.n845 gnd 0.071604f
C6509 commonsourceibias.n846 gnd 0.011785f
C6510 commonsourceibias.t189 gnd 0.194086f
C6511 commonsourceibias.n847 gnd 0.085919f
C6512 commonsourceibias.n848 gnd 0.029883f
C6513 commonsourceibias.n849 gnd 0.153509f
C6514 commonsourceibias.n850 gnd 0.012817f
C6515 commonsourceibias.t133 gnd 0.17946f
C6516 commonsourceibias.n851 gnd 0.009349f
C6517 commonsourceibias.n852 gnd 0.009605f
C6518 commonsourceibias.t153 gnd 0.17946f
C6519 commonsourceibias.n853 gnd 0.012358f
C6520 commonsourceibias.n854 gnd 0.009605f
C6521 commonsourceibias.t122 gnd 0.17946f
C6522 commonsourceibias.n855 gnd 0.009057f
C6523 commonsourceibias.n856 gnd 0.009605f
C6524 commonsourceibias.t143 gnd 0.17946f
C6525 commonsourceibias.n857 gnd 0.012174f
C6526 commonsourceibias.n858 gnd 0.009605f
C6527 commonsourceibias.t99 gnd 0.17946f
C6528 commonsourceibias.n859 gnd 0.008798f
C6529 commonsourceibias.n860 gnd 0.009605f
C6530 commonsourceibias.t87 gnd 0.17946f
C6531 commonsourceibias.n861 gnd 0.01197f
C6532 commonsourceibias.n862 gnd 0.009605f
C6533 commonsourceibias.t167 gnd 0.17946f
C6534 commonsourceibias.n863 gnd 0.008571f
C6535 commonsourceibias.n864 gnd 0.009605f
C6536 commonsourceibias.t192 gnd 0.17946f
C6537 commonsourceibias.n865 gnd 0.011742f
C6538 commonsourceibias.n866 gnd 0.009605f
C6539 commonsourceibias.t136 gnd 0.17946f
C6540 commonsourceibias.n867 gnd 0.008375f
C6541 commonsourceibias.n868 gnd 0.009605f
C6542 commonsourceibias.t181 gnd 0.17946f
C6543 commonsourceibias.n869 gnd 0.011489f
C6544 commonsourceibias.n870 gnd 0.009605f
C6545 commonsourceibias.t126 gnd 0.17946f
C6546 commonsourceibias.n871 gnd 0.008208f
C6547 commonsourceibias.n872 gnd 0.009605f
C6548 commonsourceibias.t146 gnd 0.17946f
C6549 commonsourceibias.n873 gnd 0.011208f
C6550 commonsourceibias.t191 gnd 0.199526f
C6551 commonsourceibias.t156 gnd 0.17946f
C6552 commonsourceibias.n874 gnd 0.078221f
C6553 commonsourceibias.n875 gnd 0.085838f
C6554 commonsourceibias.n876 gnd 0.03983f
C6555 commonsourceibias.n877 gnd 0.009605f
C6556 commonsourceibias.n878 gnd 0.009349f
C6557 commonsourceibias.n879 gnd 0.013398f
C6558 commonsourceibias.n880 gnd 0.071604f
C6559 commonsourceibias.n881 gnd 0.013389f
C6560 commonsourceibias.n882 gnd 0.009605f
C6561 commonsourceibias.n883 gnd 0.009605f
C6562 commonsourceibias.n884 gnd 0.009605f
C6563 commonsourceibias.n885 gnd 0.012358f
C6564 commonsourceibias.n886 gnd 0.071604f
C6565 commonsourceibias.n887 gnd 0.012648f
C6566 commonsourceibias.t91 gnd 0.17946f
C6567 commonsourceibias.n888 gnd 0.071604f
C6568 commonsourceibias.n889 gnd 0.012288f
C6569 commonsourceibias.n890 gnd 0.009605f
C6570 commonsourceibias.n891 gnd 0.009605f
C6571 commonsourceibias.n892 gnd 0.009605f
C6572 commonsourceibias.n893 gnd 0.009057f
C6573 commonsourceibias.n894 gnd 0.01341f
C6574 commonsourceibias.n895 gnd 0.071604f
C6575 commonsourceibias.n896 gnd 0.013406f
C6576 commonsourceibias.n897 gnd 0.009605f
C6577 commonsourceibias.n898 gnd 0.009605f
C6578 commonsourceibias.n899 gnd 0.009605f
C6579 commonsourceibias.n900 gnd 0.012174f
C6580 commonsourceibias.n901 gnd 0.071604f
C6581 commonsourceibias.n902 gnd 0.012558f
C6582 commonsourceibias.t107 gnd 0.17946f
C6583 commonsourceibias.n903 gnd 0.071604f
C6584 commonsourceibias.n904 gnd 0.012378f
C6585 commonsourceibias.n905 gnd 0.009605f
C6586 commonsourceibias.n906 gnd 0.009605f
C6587 commonsourceibias.n907 gnd 0.009605f
C6588 commonsourceibias.n908 gnd 0.008798f
C6589 commonsourceibias.n909 gnd 0.013415f
C6590 commonsourceibias.n910 gnd 0.071604f
C6591 commonsourceibias.n911 gnd 0.013414f
C6592 commonsourceibias.n912 gnd 0.009605f
C6593 commonsourceibias.n913 gnd 0.009605f
C6594 commonsourceibias.n914 gnd 0.009605f
C6595 commonsourceibias.n915 gnd 0.01197f
C6596 commonsourceibias.n916 gnd 0.071604f
C6597 commonsourceibias.n917 gnd 0.012468f
C6598 commonsourceibias.t127 gnd 0.17946f
C6599 commonsourceibias.n918 gnd 0.071604f
C6600 commonsourceibias.n919 gnd 0.012468f
C6601 commonsourceibias.n920 gnd 0.009605f
C6602 commonsourceibias.n921 gnd 0.009605f
C6603 commonsourceibias.n922 gnd 0.009605f
C6604 commonsourceibias.n923 gnd 0.008571f
C6605 commonsourceibias.n924 gnd 0.013414f
C6606 commonsourceibias.n925 gnd 0.071604f
C6607 commonsourceibias.n926 gnd 0.013415f
C6608 commonsourceibias.n927 gnd 0.009605f
C6609 commonsourceibias.n928 gnd 0.009605f
C6610 commonsourceibias.n929 gnd 0.009605f
C6611 commonsourceibias.n930 gnd 0.011742f
C6612 commonsourceibias.n931 gnd 0.071604f
C6613 commonsourceibias.n932 gnd 0.012378f
C6614 commonsourceibias.t137 gnd 0.17946f
C6615 commonsourceibias.n933 gnd 0.071604f
C6616 commonsourceibias.n934 gnd 0.012558f
C6617 commonsourceibias.n935 gnd 0.009605f
C6618 commonsourceibias.n936 gnd 0.009605f
C6619 commonsourceibias.n937 gnd 0.009605f
C6620 commonsourceibias.n938 gnd 0.008375f
C6621 commonsourceibias.n939 gnd 0.013406f
C6622 commonsourceibias.n940 gnd 0.071604f
C6623 commonsourceibias.n941 gnd 0.01341f
C6624 commonsourceibias.n942 gnd 0.009605f
C6625 commonsourceibias.n943 gnd 0.009605f
C6626 commonsourceibias.n944 gnd 0.009605f
C6627 commonsourceibias.n945 gnd 0.011489f
C6628 commonsourceibias.n946 gnd 0.071604f
C6629 commonsourceibias.n947 gnd 0.012288f
C6630 commonsourceibias.t170 gnd 0.17946f
C6631 commonsourceibias.n948 gnd 0.071604f
C6632 commonsourceibias.n949 gnd 0.012648f
C6633 commonsourceibias.n950 gnd 0.009605f
C6634 commonsourceibias.n951 gnd 0.009605f
C6635 commonsourceibias.n952 gnd 0.009605f
C6636 commonsourceibias.n953 gnd 0.008208f
C6637 commonsourceibias.n954 gnd 0.013389f
C6638 commonsourceibias.n955 gnd 0.071604f
C6639 commonsourceibias.n956 gnd 0.013398f
C6640 commonsourceibias.n957 gnd 0.009605f
C6641 commonsourceibias.n958 gnd 0.009605f
C6642 commonsourceibias.n959 gnd 0.009605f
C6643 commonsourceibias.n960 gnd 0.011208f
C6644 commonsourceibias.n961 gnd 0.071604f
C6645 commonsourceibias.n962 gnd 0.011785f
C6646 commonsourceibias.t101 gnd 0.194086f
C6647 commonsourceibias.n963 gnd 0.085919f
C6648 commonsourceibias.n964 gnd 0.029883f
C6649 commonsourceibias.n965 gnd 0.202572f
C6650 commonsourceibias.n966 gnd 5.28148f
.ends

