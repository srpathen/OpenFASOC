* NGSPICE file created from opamp625.ext - technology: sky130A

.subckt opamp625 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2804_13878.t29 a_n2982_13878.t52 a_n2982_13878.t53 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t113 commonsourceibias.t64 gnd.t296 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2804_13878.t0 a_n2982_13878.t72 vdd.t196 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t216 a_n9628_8799.t48 CSoutput.t200 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 gnd.t295 commonsourceibias.t65 CSoutput.t112 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 CSoutput.t111 commonsourceibias.t66 gnd.t294 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 CSoutput.t110 commonsourceibias.t67 gnd.t293 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 CSoutput.t201 a_n9628_8799.t49 vdd.t217 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X8 vdd.t230 a_n9628_8799.t50 CSoutput.t214 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 a_n2982_8322.t29 a_n2982_13878.t73 a_n9628_8799.t24 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X10 CSoutput.t215 a_n9628_8799.t51 vdd.t231 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 vdd.t118 a_n9628_8799.t52 CSoutput.t162 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 gnd.t123 gnd.t121 gnd.t122 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X13 output.t15 CSoutput.t216 vdd.t6 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X14 CSoutput.t163 a_n9628_8799.t53 vdd.t119 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 CSoutput.t109 commonsourceibias.t68 gnd.t292 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 gnd.t120 gnd.t118 gnd.t119 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X17 gnd.t117 gnd.t116 plus.t4 gnd.t53 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X18 gnd.t291 commonsourceibias.t69 CSoutput.t108 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 vdd.t7 CSoutput.t217 output.t14 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t107 commonsourceibias.t70 gnd.t290 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X21 a_n9628_8799.t47 plus.t5 a_n2903_n3924.t33 gnd.t345 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X22 gnd.t289 commonsourceibias.t71 CSoutput.t106 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t70 a_n9628_8799.t54 CSoutput.t128 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 vdd.t71 a_n9628_8799.t55 CSoutput.t129 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X25 CSoutput.t105 commonsourceibias.t72 gnd.t288 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 minus.t4 gnd.t113 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X27 CSoutput.t104 commonsourceibias.t73 gnd.t287 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 gnd.t286 commonsourceibias.t74 CSoutput.t103 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X29 commonsourceibias.t51 commonsourceibias.t50 gnd.t283 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 CSoutput.t136 a_n9628_8799.t56 vdd.t81 vdd.t67 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 CSoutput.t102 commonsourceibias.t75 gnd.t285 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 a_n9628_8799.t23 a_n2982_13878.t74 a_n2982_8322.t28 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X33 vdd.t82 a_n9628_8799.t57 CSoutput.t137 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X34 vdd.t36 a_n9628_8799.t58 CSoutput.t16 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 CSoutput.t17 a_n9628_8799.t59 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X36 a_n9628_8799.t30 a_n2982_13878.t75 a_n2982_8322.t27 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X37 CSoutput.t101 commonsourceibias.t76 gnd.t284 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 gnd.t282 commonsourceibias.t77 CSoutput.t100 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 gnd.t112 gnd.t110 gnd.t111 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X40 a_n9628_8799.t6 plus.t6 a_n2903_n3924.t32 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X41 CSoutput.t99 commonsourceibias.t78 gnd.t281 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 CSoutput.t98 commonsourceibias.t79 gnd.t280 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 gnd.t109 gnd.t107 gnd.t108 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X44 CSoutput.t97 commonsourceibias.t80 gnd.t279 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X45 vdd.t8 CSoutput.t218 output.t13 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X46 CSoutput.t198 a_n9628_8799.t60 vdd.t214 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 a_n2903_n3924.t50 diffpairibias.t16 gnd.t352 gnd.t351 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X48 a_n2903_n3924.t2 minus.t5 a_n2982_13878.t1 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X49 CSoutput.t199 a_n9628_8799.t61 vdd.t215 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 vdd.t26 a_n9628_8799.t62 CSoutput.t10 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X51 gnd.t278 commonsourceibias.t81 CSoutput.t96 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 a_n2903_n3924.t31 plus.t7 a_n9628_8799.t11 gnd.t320 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X53 vdd.t28 a_n9628_8799.t63 CSoutput.t11 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 CSoutput.t95 commonsourceibias.t82 gnd.t277 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X55 a_n2982_13878.t13 minus.t6 a_n2903_n3924.t42 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X56 output.t16 outputibias.t8 gnd.t318 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X57 gnd.t276 commonsourceibias.t48 commonsourceibias.t49 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 CSoutput.t94 commonsourceibias.t83 gnd.t275 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 CSoutput.t219 a_n2982_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X60 a_n2903_n3924.t30 plus.t8 a_n9628_8799.t13 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X61 vdd.t307 vdd.t305 vdd.t306 vdd.t296 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X62 a_n2903_n3924.t49 minus.t7 a_n2982_13878.t19 gnd.t321 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X63 gnd.t274 commonsourceibias.t84 CSoutput.t93 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 vdd.t115 a_n9628_8799.t64 CSoutput.t160 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 vdd.t39 CSoutput.t220 output.t12 gnd.t130 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X66 a_n2804_13878.t28 a_n2982_13878.t54 a_n2982_13878.t55 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X67 CSoutput.t92 commonsourceibias.t85 gnd.t273 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 gnd.t272 commonsourceibias.t86 CSoutput.t91 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 output.t11 CSoutput.t221 vdd.t40 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X70 a_n2982_13878.t57 a_n2982_13878.t56 a_n2804_13878.t27 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X71 CSoutput.t90 commonsourceibias.t87 gnd.t271 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 vdd.t304 vdd.t302 vdd.t303 vdd.t296 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X73 gnd.t270 commonsourceibias.t88 CSoutput.t89 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 CSoutput.t161 a_n9628_8799.t65 vdd.t117 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd.t301 vdd.t299 vdd.t300 vdd.t278 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X76 gnd.t269 commonsourceibias.t60 commonsourceibias.t61 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 a_n2903_n3924.t9 minus.t8 a_n2982_13878.t5 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X78 vdd.t137 a_n9628_8799.t66 CSoutput.t178 vdd.t69 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 CSoutput.t88 commonsourceibias.t89 gnd.t268 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 vdd.t138 a_n9628_8799.t67 CSoutput.t179 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X81 gnd.t106 gnd.t103 gnd.t105 gnd.t104 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X82 gnd.t102 gnd.t100 gnd.t101 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X83 CSoutput.t87 commonsourceibias.t90 gnd.t267 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 diffpairibias.t15 diffpairibias.t14 gnd.t358 gnd.t357 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X85 CSoutput.t172 a_n9628_8799.t68 vdd.t130 vdd.t67 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 a_n2982_13878.t59 a_n2982_13878.t58 a_n2804_13878.t26 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X87 CSoutput.t86 commonsourceibias.t91 gnd.t266 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X88 CSoutput.t173 a_n9628_8799.t69 vdd.t132 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 CSoutput.t85 commonsourceibias.t92 gnd.t265 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 gnd.t264 commonsourceibias.t93 CSoutput.t84 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n9628_8799.t29 a_n2982_13878.t76 a_n2982_8322.t26 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 gnd.t263 commonsourceibias.t94 CSoutput.t83 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 vdd.t212 a_n9628_8799.t70 CSoutput.t196 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X94 CSoutput.t197 a_n9628_8799.t71 vdd.t213 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X95 gnd.t262 commonsourceibias.t95 CSoutput.t82 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X96 CSoutput.t222 a_n2982_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X97 a_n2982_13878.t0 minus.t9 a_n2903_n3924.t1 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X98 a_n2982_13878.t61 a_n2982_13878.t60 a_n2804_13878.t25 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X99 gnd.t99 gnd.t97 plus.t3 gnd.t98 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X100 vdd.t228 a_n9628_8799.t72 CSoutput.t212 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 vdd.t229 a_n9628_8799.t73 CSoutput.t213 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n9628_8799.t26 a_n2982_13878.t77 a_n2982_8322.t25 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X103 CSoutput.t158 a_n9628_8799.t74 vdd.t112 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 CSoutput.t81 commonsourceibias.t96 gnd.t261 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 diffpairibias.t13 diffpairibias.t12 gnd.t366 gnd.t365 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X106 CSoutput.t159 a_n9628_8799.t75 vdd.t113 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 gnd.t253 commonsourceibias.t2 commonsourceibias.t3 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t254 commonsourceibias.t97 CSoutput.t80 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X109 a_n9628_8799.t25 a_n2982_13878.t78 a_n2982_8322.t24 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X110 CSoutput.t79 commonsourceibias.t98 gnd.t260 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 gnd.t259 commonsourceibias.t99 CSoutput.t78 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X112 gnd.t96 gnd.t94 gnd.t95 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X113 CSoutput.t77 commonsourceibias.t100 gnd.t258 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 CSoutput.t76 commonsourceibias.t101 gnd.t255 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 a_n2982_8322.t23 a_n2982_13878.t79 a_n9628_8799.t22 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X116 gnd.t257 commonsourceibias.t102 CSoutput.t75 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 CSoutput.t126 a_n9628_8799.t76 vdd.t66 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X118 plus.t2 gnd.t91 gnd.t93 gnd.t92 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X119 gnd.t256 commonsourceibias.t62 commonsourceibias.t63 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 output.t10 CSoutput.t223 vdd.t41 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X121 vdd.t47 CSoutput.t224 output.t9 gnd.t301 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X122 a_n9628_8799.t0 plus.t9 a_n2903_n3924.t29 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X123 vdd.t298 vdd.t295 vdd.t297 vdd.t296 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X124 gnd.t252 commonsourceibias.t103 CSoutput.t74 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X125 a_n2903_n3924.t0 diffpairibias.t17 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X126 CSoutput.t127 a_n9628_8799.t77 vdd.t68 vdd.t67 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X127 vdd.t79 a_n9628_8799.t78 CSoutput.t134 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X128 gnd.t90 gnd.t88 gnd.t89 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X129 a_n2903_n3924.t48 minus.t10 a_n2982_13878.t18 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X130 vdd.t80 a_n9628_8799.t79 CSoutput.t135 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 a_n2982_13878.t63 a_n2982_13878.t62 a_n2804_13878.t24 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X132 vdd.t210 a_n9628_8799.t80 CSoutput.t194 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 gnd.t251 commonsourceibias.t104 CSoutput.t73 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 a_n9628_8799.t21 a_n2982_13878.t80 a_n2982_8322.t22 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X135 a_n2982_13878.t51 a_n2982_13878.t50 a_n2804_13878.t23 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X136 a_n2982_13878.t11 minus.t11 a_n2903_n3924.t40 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X137 gnd.t87 gnd.t85 gnd.t86 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X138 vdd.t48 CSoutput.t225 output.t8 gnd.t302 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X139 a_n2903_n3924.t28 plus.t10 a_n9628_8799.t7 gnd.t310 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X140 CSoutput.t72 commonsourceibias.t105 gnd.t250 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 CSoutput.t195 a_n9628_8799.t81 vdd.t211 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 vdd.t22 a_n9628_8799.t82 CSoutput.t8 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X143 gnd.t249 commonsourceibias.t106 CSoutput.t71 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 CSoutput.t9 a_n9628_8799.t83 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X145 a_n2903_n3924.t53 minus.t12 a_n2982_13878.t69 gnd.t350 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X146 vdd.t294 vdd.t292 vdd.t293 vdd.t285 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X147 gnd.t248 commonsourceibias.t0 commonsourceibias.t1 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 output.t7 CSoutput.t226 vdd.t49 gnd.t303 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X149 gnd.t247 commonsourceibias.t107 CSoutput.t70 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X150 CSoutput.t156 a_n9628_8799.t84 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 vdd.t291 vdd.t288 vdd.t290 vdd.t289 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X152 a_n2804_13878.t22 a_n2982_13878.t46 a_n2982_13878.t47 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X153 CSoutput.t157 a_n9628_8799.t85 vdd.t111 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X154 vdd.t135 a_n9628_8799.t86 CSoutput.t176 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 vdd.t192 a_n2982_13878.t81 a_n2982_8322.t37 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 a_n2982_13878.t23 a_n2982_13878.t22 a_n2804_13878.t21 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X157 a_n2982_8322.t36 a_n2982_13878.t82 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X158 gnd.t246 commonsourceibias.t108 CSoutput.t69 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X159 a_n2903_n3924.t51 diffpairibias.t18 gnd.t356 gnd.t355 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X160 CSoutput.t177 a_n9628_8799.t87 vdd.t136 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 output.t6 CSoutput.t227 vdd.t50 gnd.t304 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X162 gnd.t245 commonsourceibias.t109 CSoutput.t68 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n2982_13878.t4 minus.t13 a_n2903_n3924.t8 gnd.t324 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X164 gnd.t244 commonsourceibias.t16 commonsourceibias.t17 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 CSoutput.t67 commonsourceibias.t110 gnd.t243 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 gnd.t242 commonsourceibias.t111 CSoutput.t66 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 CSoutput.t65 commonsourceibias.t112 gnd.t241 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X168 CSoutput.t64 commonsourceibias.t113 gnd.t240 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 a_n2903_n3924.t27 plus.t11 a_n9628_8799.t4 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X170 vdd.t188 a_n2982_13878.t83 a_n2804_13878.t2 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X171 gnd.t84 gnd.t82 minus.t3 gnd.t83 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X172 vdd.t287 vdd.t284 vdd.t286 vdd.t285 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X173 gnd.t81 gnd.t79 gnd.t80 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X174 a_n2804_13878.t20 a_n2982_13878.t32 a_n2982_13878.t33 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 vdd.t30 a_n9628_8799.t88 CSoutput.t12 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X176 vdd.t31 a_n9628_8799.t89 CSoutput.t13 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X177 a_n2982_8322.t21 a_n2982_13878.t84 a_n9628_8799.t32 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X178 a_n9628_8799.t17 plus.t12 a_n2903_n3924.t26 gnd.t335 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X179 vdd.t283 vdd.t281 vdd.t282 vdd.t258 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X180 vdd.t280 vdd.t277 vdd.t279 vdd.t278 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X181 a_n2982_8322.t35 a_n2982_13878.t85 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X182 a_n9628_8799.t31 a_n2982_13878.t86 a_n2982_8322.t20 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X183 a_n2982_13878.t6 minus.t14 a_n2903_n3924.t34 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X184 CSoutput.t0 a_n9628_8799.t90 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X185 diffpairibias.t11 diffpairibias.t10 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 vdd.t3 a_n9628_8799.t91 CSoutput.t1 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X187 a_n2982_13878.t27 a_n2982_13878.t26 a_n2804_13878.t19 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X188 CSoutput.t63 commonsourceibias.t114 gnd.t239 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n9628_8799.t34 a_n2982_13878.t87 a_n2982_8322.t19 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X190 CSoutput.t192 a_n9628_8799.t92 vdd.t208 vdd.t131 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X191 CSoutput.t193 a_n9628_8799.t93 vdd.t209 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 commonsourceibias.t15 commonsourceibias.t14 gnd.t238 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 gnd.t237 commonsourceibias.t115 CSoutput.t62 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 a_n2804_13878.t18 a_n2982_13878.t24 a_n2982_13878.t25 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X195 gnd.t78 gnd.t75 gnd.t77 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X196 CSoutput.t61 commonsourceibias.t116 gnd.t236 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 a_n9628_8799.t10 plus.t13 a_n2903_n3924.t25 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X198 a_n2903_n3924.t35 minus.t15 a_n2982_13878.t7 gnd.t328 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X199 a_n2903_n3924.t38 minus.t16 a_n2982_13878.t9 gnd.t336 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X200 vdd.t276 vdd.t274 vdd.t275 vdd.t237 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X201 CSoutput.t210 a_n9628_8799.t94 vdd.t226 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 outputibias.t7 outputibias.t6 gnd.t342 gnd.t341 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X203 vdd.t83 CSoutput.t228 output.t5 gnd.t325 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X204 a_n2982_13878.t68 minus.t17 a_n2903_n3924.t52 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X205 CSoutput.t60 commonsourceibias.t117 gnd.t235 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 gnd.t74 gnd.t72 gnd.t73 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X207 vdd.t181 a_n2982_13878.t88 a_n2982_8322.t34 vdd.t180 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X208 a_n2804_13878.t17 a_n2982_13878.t48 a_n2982_13878.t49 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 vdd.t227 a_n9628_8799.t95 CSoutput.t211 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 vdd.t107 a_n9628_8799.t96 CSoutput.t154 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 a_n2982_13878.t21 a_n2982_13878.t20 a_n2804_13878.t16 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X212 gnd.t234 commonsourceibias.t118 CSoutput.t59 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 gnd.t233 commonsourceibias.t119 CSoutput.t58 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 commonsourceibias.t41 commonsourceibias.t40 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 outputibias.t5 outputibias.t4 gnd.t347 gnd.t346 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X216 gnd.t230 commonsourceibias.t120 CSoutput.t57 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X217 vdd.t108 a_n9628_8799.t97 CSoutput.t155 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 vdd.t206 a_n9628_8799.t98 CSoutput.t190 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X219 CSoutput.t191 a_n9628_8799.t99 vdd.t207 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 CSoutput.t56 commonsourceibias.t121 gnd.t229 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 a_n2903_n3924.t43 diffpairibias.t19 gnd.t344 gnd.t343 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X222 gnd.t71 gnd.t68 gnd.t70 gnd.t69 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X223 vdd.t273 vdd.t271 vdd.t272 vdd.t245 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X224 a_n2903_n3924.t36 diffpairibias.t20 gnd.t332 gnd.t331 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X225 commonsourceibias.t39 commonsourceibias.t38 gnd.t228 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 a_n2982_13878.t15 minus.t18 a_n2903_n3924.t45 gnd.t345 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X227 vdd.t224 a_n9628_8799.t100 CSoutput.t208 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X228 vdd.t225 a_n9628_8799.t101 CSoutput.t209 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 CSoutput.t152 a_n9628_8799.t102 vdd.t103 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 gnd.t67 gnd.t65 gnd.t66 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X231 gnd.t64 gnd.t62 gnd.t63 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X232 gnd.t61 gnd.t59 minus.t2 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X233 vdd.t270 vdd.t268 vdd.t269 vdd.t258 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X234 CSoutput.t55 commonsourceibias.t122 gnd.t226 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 CSoutput.t54 commonsourceibias.t123 gnd.t225 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 a_n2804_13878.t15 a_n2982_13878.t40 a_n2982_13878.t41 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X237 CSoutput.t153 a_n9628_8799.t103 vdd.t105 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 a_n2982_8322.t18 a_n2982_13878.t89 a_n9628_8799.t33 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X239 CSoutput.t142 a_n9628_8799.t104 vdd.t90 vdd.t59 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X240 commonsourceibias.t35 commonsourceibias.t34 gnd.t222 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 a_n2982_13878.t3 minus.t19 a_n2903_n3924.t6 gnd.t309 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X242 CSoutput.t229 a_n2982_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X243 gnd.t224 commonsourceibias.t36 commonsourceibias.t37 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 diffpairibias.t9 diffpairibias.t8 gnd.t334 gnd.t333 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X245 a_n2804_13878.t4 a_n2982_13878.t90 vdd.t177 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 vdd.t175 a_n2982_13878.t91 a_n2804_13878.t3 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X247 CSoutput.t53 commonsourceibias.t124 gnd.t221 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 CSoutput.t52 commonsourceibias.t125 gnd.t220 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t143 a_n9628_8799.t105 vdd.t92 vdd.t91 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 CSoutput.t230 a_n2982_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X251 a_n2903_n3924.t24 plus.t14 a_n9628_8799.t45 gnd.t136 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X252 gnd.t219 commonsourceibias.t32 commonsourceibias.t33 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 vdd.t203 a_n9628_8799.t106 CSoutput.t188 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X254 vdd.t205 a_n9628_8799.t107 CSoutput.t189 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X255 vdd.t18 a_n9628_8799.t108 CSoutput.t6 vdd.t17 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 commonsourceibias.t31 commonsourceibias.t30 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 CSoutput.t7 a_n9628_8799.t109 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 a_n2903_n3924.t55 minus.t20 a_n2982_13878.t71 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X259 a_n2804_13878.t14 a_n2982_13878.t30 a_n2982_13878.t31 vdd.t173 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X260 a_n2903_n3924.t23 plus.t15 a_n9628_8799.t12 gnd.t321 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X261 gnd.t215 commonsourceibias.t126 CSoutput.t51 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 a_n2903_n3924.t4 minus.t21 a_n2982_13878.t2 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X263 commonsourceibias.t29 commonsourceibias.t28 gnd.t214 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X264 a_n9628_8799.t14 plus.t16 a_n2903_n3924.t22 gnd.t330 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X265 vdd.t101 a_n9628_8799.t110 CSoutput.t150 vdd.t21 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X266 vdd.t102 a_n9628_8799.t111 CSoutput.t151 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 output.t18 outputibias.t9 gnd.t360 gnd.t359 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X268 CSoutput.t14 a_n9628_8799.t112 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 gnd.t213 commonsourceibias.t26 commonsourceibias.t27 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 a_n2982_8322.t17 a_n2982_13878.t92 a_n9628_8799.t28 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X271 a_n2982_13878.t65 a_n2982_13878.t64 a_n2804_13878.t13 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X272 CSoutput.t50 commonsourceibias.t127 gnd.t212 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 CSoutput.t15 a_n9628_8799.t113 vdd.t35 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X274 diffpairibias.t7 diffpairibias.t6 gnd.t362 gnd.t361 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X275 vdd.t14 a_n9628_8799.t114 CSoutput.t4 vdd.t13 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X276 a_n2804_13878.t12 a_n2982_13878.t36 a_n2982_13878.t37 vdd.t171 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X277 commonsourceibias.t47 commonsourceibias.t46 gnd.t198 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 vdd.t170 a_n2982_13878.t93 a_n2982_8322.t33 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X279 vdd.t84 CSoutput.t231 output.t4 gnd.t326 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X280 vdd.t16 a_n9628_8799.t115 CSoutput.t5 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X281 gnd.t211 commonsourceibias.t128 CSoutput.t49 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X282 CSoutput.t170 a_n9628_8799.t116 vdd.t128 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X283 gnd.t210 commonsourceibias.t12 commonsourceibias.t13 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X284 CSoutput.t48 commonsourceibias.t129 gnd.t199 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X285 a_n2804_13878.t1 a_n2982_13878.t94 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X286 plus.t1 gnd.t56 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X287 vdd.t129 a_n9628_8799.t117 CSoutput.t171 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 CSoutput.t202 a_n9628_8799.t118 vdd.t218 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X289 CSoutput.t203 a_n9628_8799.t119 vdd.t219 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 gnd.t55 gnd.t52 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X291 gnd.t208 commonsourceibias.t130 CSoutput.t47 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 gnd.t51 gnd.t49 minus.t1 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X293 gnd.t48 gnd.t45 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X294 vdd.t63 a_n9628_8799.t120 CSoutput.t124 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 gnd.t44 gnd.t41 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X296 vdd.t267 vdd.t265 vdd.t266 vdd.t241 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X297 a_n2903_n3924.t3 diffpairibias.t21 gnd.t298 gnd.t297 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X298 a_n2982_8322.t16 a_n2982_13878.t95 a_n9628_8799.t27 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X299 vdd.t165 a_n2982_13878.t96 a_n2982_8322.t32 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X300 gnd.t207 commonsourceibias.t10 commonsourceibias.t11 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 vdd.t65 a_n9628_8799.t121 CSoutput.t125 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 gnd.t40 gnd.t38 gnd.t39 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X303 gnd.t206 commonsourceibias.t8 commonsourceibias.t9 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 a_n2903_n3924.t21 plus.t17 a_n9628_8799.t1 gnd.t129 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X305 vdd.t264 vdd.t261 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X306 gnd.t37 gnd.t35 gnd.t36 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X307 CSoutput.t46 commonsourceibias.t131 gnd.t205 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 vdd.t86 a_n9628_8799.t122 CSoutput.t138 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 vdd.t87 a_n9628_8799.t123 CSoutput.t139 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 output.t3 CSoutput.t232 vdd.t45 gnd.t299 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X311 vdd.t88 a_n9628_8799.t124 CSoutput.t140 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 CSoutput.t141 a_n9628_8799.t125 vdd.t89 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X313 a_n9628_8799.t2 plus.t18 a_n2903_n3924.t20 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X314 CSoutput.t118 a_n9628_8799.t126 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 CSoutput.t45 commonsourceibias.t132 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 CSoutput.t119 a_n9628_8799.t127 vdd.t57 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X317 CSoutput.t116 a_n9628_8799.t128 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 a_n2903_n3924.t47 minus.t22 a_n2982_13878.t17 gnd.t310 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X319 a_n2804_13878.t11 a_n2982_13878.t42 a_n2982_13878.t43 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X320 a_n2982_8322.t15 a_n2982_13878.t97 a_n9628_8799.t36 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X321 diffpairibias.t5 diffpairibias.t4 gnd.t316 gnd.t315 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X322 a_n2903_n3924.t46 minus.t23 a_n2982_13878.t16 gnd.t320 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X323 a_n9628_8799.t8 plus.t19 a_n2903_n3924.t19 gnd.t311 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X324 gnd.t34 gnd.t31 gnd.t33 gnd.t32 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X325 CSoutput.t117 a_n9628_8799.t129 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X326 CSoutput.t168 a_n9628_8799.t130 vdd.t126 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 gnd.t202 commonsourceibias.t6 commonsourceibias.t7 gnd.t201 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X328 vdd.t260 vdd.t257 vdd.t259 vdd.t258 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X329 vdd.t127 a_n9628_8799.t131 CSoutput.t169 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 CSoutput.t44 commonsourceibias.t133 gnd.t200 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 CSoutput.t233 a_n2982_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X332 a_n2982_8322.t31 a_n2982_13878.t98 vdd.t162 vdd.t161 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X333 CSoutput.t114 a_n9628_8799.t132 vdd.t42 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 outputibias.t3 outputibias.t2 gnd.t349 gnd.t348 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X335 a_n2903_n3924.t18 plus.t20 a_n9628_8799.t5 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X336 vdd.t44 a_n9628_8799.t133 CSoutput.t115 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 gnd.t196 commonsourceibias.t134 CSoutput.t43 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 CSoutput.t164 a_n9628_8799.t134 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 output.t19 outputibias.t10 gnd.t364 gnd.t363 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X340 vdd.t160 a_n2982_13878.t99 a_n2804_13878.t31 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X341 vdd.t122 a_n9628_8799.t135 CSoutput.t165 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput.t180 a_n9628_8799.t136 vdd.t139 vdd.t116 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 vdd.t140 a_n9628_8799.t137 CSoutput.t181 vdd.t64 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 a_n9628_8799.t18 plus.t21 a_n2903_n3924.t17 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X345 gnd.t195 commonsourceibias.t135 CSoutput.t42 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 a_n2903_n3924.t41 minus.t24 a_n2982_13878.t12 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X347 output.t17 outputibias.t11 gnd.t338 gnd.t337 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X348 gnd.t194 commonsourceibias.t136 CSoutput.t41 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 a_n2982_8322.t14 a_n2982_13878.t100 a_n9628_8799.t35 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X350 commonsourceibias.t45 commonsourceibias.t44 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 a_n9628_8799.t38 a_n2982_13878.t101 a_n2982_8322.t13 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X352 a_n2804_13878.t30 a_n2982_13878.t102 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X353 gnd.t191 commonsourceibias.t137 CSoutput.t40 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 vdd.t201 a_n9628_8799.t138 CSoutput.t186 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 vdd.t256 vdd.t254 vdd.t255 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X356 vdd.t253 vdd.t251 vdd.t252 vdd.t245 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X357 vdd.t202 a_n9628_8799.t139 CSoutput.t187 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 CSoutput.t206 a_n9628_8799.t140 vdd.t222 vdd.t51 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 CSoutput.t207 a_n9628_8799.t141 vdd.t223 vdd.t34 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X360 CSoutput.t148 a_n9628_8799.t142 vdd.t98 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 commonsourceibias.t43 commonsourceibias.t42 gnd.t190 gnd.t189 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 a_n2982_13878.t45 a_n2982_13878.t44 a_n2804_13878.t10 vdd.t146 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X363 a_n9628_8799.t37 a_n2982_13878.t103 a_n2982_8322.t12 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X364 a_n9628_8799.t46 plus.t22 a_n2903_n3924.t16 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X365 gnd.t30 gnd.t27 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X366 a_n9628_8799.t40 a_n2982_13878.t104 a_n2982_8322.t11 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X367 gnd.t188 commonsourceibias.t138 CSoutput.t39 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X368 a_n2982_8322.t10 a_n2982_13878.t105 a_n9628_8799.t39 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X369 commonsourceibias.t25 commonsourceibias.t24 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 gnd.t185 commonsourceibias.t139 CSoutput.t38 gnd.t184 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 a_n2982_13878.t10 minus.t25 a_n2903_n3924.t39 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X372 CSoutput.t37 commonsourceibias.t140 gnd.t183 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X373 vdd.t100 a_n9628_8799.t143 CSoutput.t149 vdd.t99 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 gnd.t182 commonsourceibias.t22 commonsourceibias.t23 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X375 CSoutput.t122 a_n9628_8799.t144 vdd.t61 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t123 a_n9628_8799.t145 vdd.t62 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X377 CSoutput.t132 a_n9628_8799.t146 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 CSoutput.t133 a_n9628_8799.t147 vdd.t78 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 gnd.t26 gnd.t23 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X380 a_n2804_13878.t9 a_n2982_13878.t34 a_n2982_13878.t35 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X381 vdd.t199 a_n9628_8799.t148 CSoutput.t184 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 vdd.t200 a_n9628_8799.t149 CSoutput.t185 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 vdd.t10 a_n9628_8799.t150 CSoutput.t2 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 gnd.t180 commonsourceibias.t20 commonsourceibias.t21 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X385 a_n2903_n3924.t15 plus.t23 a_n9628_8799.t20 gnd.t336 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X386 commonsourceibias.t19 commonsourceibias.t18 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 gnd.t177 commonsourceibias.t141 CSoutput.t36 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X388 a_n9628_8799.t9 plus.t24 a_n2903_n3924.t14 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X389 a_n2903_n3924.t7 diffpairibias.t22 gnd.t323 gnd.t322 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X390 gnd.t176 commonsourceibias.t142 CSoutput.t35 gnd.t175 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X391 vdd.t12 a_n9628_8799.t151 CSoutput.t3 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X392 CSoutput.t34 commonsourceibias.t143 gnd.t174 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X393 output.t2 CSoutput.t234 vdd.t46 gnd.t300 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X394 gnd.t173 commonsourceibias.t144 CSoutput.t33 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X395 CSoutput.t146 a_n9628_8799.t152 vdd.t95 vdd.t59 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 CSoutput.t32 commonsourceibias.t145 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 a_n2982_13878.t67 a_n2982_13878.t66 a_n2804_13878.t8 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X398 gnd.t22 gnd.t19 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X399 a_n9628_8799.t44 a_n2982_13878.t106 a_n2982_8322.t9 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X400 vdd.t96 a_n9628_8799.t153 CSoutput.t147 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 CSoutput.t235 a_n2982_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X402 CSoutput.t174 a_n9628_8799.t154 vdd.t133 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 vdd.t250 vdd.t248 vdd.t249 vdd.t241 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X404 a_n2903_n3924.t13 plus.t25 a_n9628_8799.t19 gnd.t350 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X405 CSoutput.t31 commonsourceibias.t146 gnd.t169 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 gnd.t168 commonsourceibias.t147 CSoutput.t30 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X407 commonsourceibias.t5 commonsourceibias.t4 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X408 CSoutput.t175 a_n9628_8799.t155 vdd.t134 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X409 diffpairibias.t3 diffpairibias.t2 gnd.t125 gnd.t124 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X410 outputibias.t1 outputibias.t0 gnd.t340 gnd.t339 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X411 a_n2982_8322.t8 a_n2982_13878.t107 a_n9628_8799.t43 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X412 gnd.t164 commonsourceibias.t148 CSoutput.t29 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 vdd.t247 vdd.t244 vdd.t246 vdd.t245 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X414 vdd.t124 a_n9628_8799.t156 CSoutput.t166 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 CSoutput.t167 a_n9628_8799.t157 vdd.t125 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X416 gnd.t15 gnd.t12 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X417 CSoutput.t182 a_n9628_8799.t158 vdd.t197 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X418 diffpairibias.t1 diffpairibias.t0 gnd.t354 gnd.t353 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X419 gnd.t163 commonsourceibias.t149 CSoutput.t28 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X420 gnd.t18 gnd.t16 plus.t0 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X421 a_n9628_8799.t15 plus.t26 a_n2903_n3924.t12 gnd.t324 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X422 commonsourceibias.t55 commonsourceibias.t54 gnd.t161 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 gnd.t160 commonsourceibias.t150 CSoutput.t27 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 CSoutput.t26 commonsourceibias.t151 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X425 minus.t0 gnd.t9 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X426 vdd.t148 a_n2982_13878.t108 a_n2804_13878.t5 vdd.t147 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X427 CSoutput.t183 a_n9628_8799.t159 vdd.t198 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X428 CSoutput.t204 a_n9628_8799.t160 vdd.t220 vdd.t76 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X429 vdd.t221 a_n9628_8799.t161 CSoutput.t205 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X430 vdd.t93 a_n9628_8799.t162 CSoutput.t144 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X431 gnd.t142 commonsourceibias.t58 commonsourceibias.t59 gnd.t141 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X432 a_n2982_8322.t7 a_n2982_13878.t109 a_n9628_8799.t42 vdd.t146 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X433 vdd.t4 CSoutput.t236 output.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X434 gnd.t144 commonsourceibias.t152 CSoutput.t25 gnd.t143 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X435 a_n2982_13878.t8 minus.t26 a_n2903_n3924.t37 gnd.t335 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X436 commonsourceibias.t53 commonsourceibias.t52 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X437 output.t0 CSoutput.t237 vdd.t5 gnd.t1 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X438 gnd.t155 commonsourceibias.t153 CSoutput.t24 gnd.t154 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X439 gnd.t8 gnd.t5 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X440 gnd.t153 commonsourceibias.t154 CSoutput.t23 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X441 a_n2982_8322.t6 a_n2982_13878.t110 a_n9628_8799.t41 vdd.t145 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X442 vdd.t94 a_n9628_8799.t163 CSoutput.t145 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X443 vdd.t58 a_n9628_8799.t164 CSoutput.t120 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X444 CSoutput.t121 a_n9628_8799.t165 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X445 gnd.t151 commonsourceibias.t155 CSoutput.t22 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X446 a_n2903_n3924.t11 plus.t27 a_n9628_8799.t3 gnd.t134 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X447 vdd.t243 vdd.t240 vdd.t242 vdd.t241 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X448 a_n2982_8322.t30 a_n2982_13878.t111 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X449 a_n2982_13878.t14 minus.t27 a_n2903_n3924.t44 gnd.t330 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X450 gnd.t150 commonsourceibias.t156 CSoutput.t21 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X451 a_n2804_13878.t7 a_n2982_13878.t38 a_n2982_13878.t39 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X452 gnd.t148 commonsourceibias.t157 CSoutput.t20 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X453 CSoutput.t19 commonsourceibias.t158 gnd.t146 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X454 commonsourceibias.t57 commonsourceibias.t56 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X455 CSoutput.t18 commonsourceibias.t159 gnd.t138 gnd.t137 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X456 vdd.t239 vdd.t236 vdd.t238 vdd.t237 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X457 a_n2903_n3924.t5 diffpairibias.t23 gnd.t313 gnd.t312 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X458 a_n2982_13878.t70 minus.t28 a_n2903_n3924.t54 gnd.t319 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X459 vdd.t235 vdd.t232 vdd.t234 vdd.t233 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X460 vdd.t73 a_n9628_8799.t166 CSoutput.t130 vdd.t72 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X461 CSoutput.t131 a_n9628_8799.t167 vdd.t75 vdd.t74 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X462 a_n2982_13878.t29 a_n2982_13878.t28 a_n2804_13878.t6 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X463 a_n2903_n3924.t10 plus.t28 a_n9628_8799.t16 gnd.t328 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
R0 a_n2982_13878.n137 a_n2982_13878.t94 512.366
R1 a_n2982_13878.n136 a_n2982_13878.t83 512.366
R2 a_n2982_13878.n135 a_n2982_13878.t72 512.366
R3 a_n2982_13878.n139 a_n2982_13878.t102 512.366
R4 a_n2982_13878.n138 a_n2982_13878.t91 512.366
R5 a_n2982_13878.n134 a_n2982_13878.t90 512.366
R6 a_n2982_13878.n141 a_n2982_13878.t98 512.366
R7 a_n2982_13878.n140 a_n2982_13878.t81 512.366
R8 a_n2982_13878.n133 a_n2982_13878.t82 512.366
R9 a_n2982_13878.n143 a_n2982_13878.t85 512.366
R10 a_n2982_13878.n142 a_n2982_13878.t96 512.366
R11 a_n2982_13878.n132 a_n2982_13878.t111 512.366
R12 a_n2982_13878.n31 a_n2982_13878.t110 538.698
R13 a_n2982_13878.n118 a_n2982_13878.t87 512.366
R14 a_n2982_13878.n117 a_n2982_13878.t92 512.366
R15 a_n2982_13878.n109 a_n2982_13878.t80 512.366
R16 a_n2982_13878.n116 a_n2982_13878.t97 512.366
R17 a_n2982_13878.n115 a_n2982_13878.t106 512.366
R18 a_n2982_13878.n110 a_n2982_13878.t107 512.366
R19 a_n2982_13878.n114 a_n2982_13878.t74 512.366
R20 a_n2982_13878.n113 a_n2982_13878.t89 512.366
R21 a_n2982_13878.n111 a_n2982_13878.t77 512.366
R22 a_n2982_13878.n112 a_n2982_13878.t84 512.366
R23 a_n2982_13878.n25 a_n2982_13878.t44 538.698
R24 a_n2982_13878.n125 a_n2982_13878.t32 512.366
R25 a_n2982_13878.n124 a_n2982_13878.t60 512.366
R26 a_n2982_13878.n94 a_n2982_13878.t40 512.366
R27 a_n2982_13878.n123 a_n2982_13878.t22 512.366
R28 a_n2982_13878.n122 a_n2982_13878.t30 512.366
R29 a_n2982_13878.n95 a_n2982_13878.t66 512.366
R30 a_n2982_13878.n121 a_n2982_13878.t42 512.366
R31 a_n2982_13878.n120 a_n2982_13878.t62 512.366
R32 a_n2982_13878.n96 a_n2982_13878.t34 512.366
R33 a_n2982_13878.n119 a_n2982_13878.t26 512.366
R34 a_n2982_13878.n13 a_n2982_13878.t50 538.698
R35 a_n2982_13878.n151 a_n2982_13878.t52 512.366
R36 a_n2982_13878.n89 a_n2982_13878.t28 512.366
R37 a_n2982_13878.n152 a_n2982_13878.t24 512.366
R38 a_n2982_13878.n88 a_n2982_13878.t56 512.366
R39 a_n2982_13878.n153 a_n2982_13878.t54 512.366
R40 a_n2982_13878.n154 a_n2982_13878.t20 512.366
R41 a_n2982_13878.n87 a_n2982_13878.t48 512.366
R42 a_n2982_13878.n155 a_n2982_13878.t58 512.366
R43 a_n2982_13878.n86 a_n2982_13878.t36 512.366
R44 a_n2982_13878.n156 a_n2982_13878.t64 512.366
R45 a_n2982_13878.n19 a_n2982_13878.t109 538.698
R46 a_n2982_13878.n145 a_n2982_13878.t78 512.366
R47 a_n2982_13878.n93 a_n2982_13878.t79 512.366
R48 a_n2982_13878.n146 a_n2982_13878.t104 512.366
R49 a_n2982_13878.n92 a_n2982_13878.t105 512.366
R50 a_n2982_13878.n147 a_n2982_13878.t76 512.366
R51 a_n2982_13878.n148 a_n2982_13878.t100 512.366
R52 a_n2982_13878.n91 a_n2982_13878.t101 512.366
R53 a_n2982_13878.n149 a_n2982_13878.t73 512.366
R54 a_n2982_13878.n90 a_n2982_13878.t86 512.366
R55 a_n2982_13878.n150 a_n2982_13878.t95 512.366
R56 a_n2982_13878.n0 a_n2982_13878.n82 70.1674
R57 a_n2982_13878.n2 a_n2982_13878.n80 70.1674
R58 a_n2982_13878.n4 a_n2982_13878.n78 70.1674
R59 a_n2982_13878.n6 a_n2982_13878.n76 70.1674
R60 a_n2982_13878.n51 a_n2982_13878.n26 70.5844
R61 a_n2982_13878.n83 a_n2982_13878.n20 70.5844
R62 a_n2982_13878.n26 a_n2982_13878.n49 70.1674
R63 a_n2982_13878.n49 a_n2982_13878.n111 20.9683
R64 a_n2982_13878.n48 a_n2982_13878.n27 74.73
R65 a_n2982_13878.n113 a_n2982_13878.n48 11.843
R66 a_n2982_13878.n47 a_n2982_13878.n27 80.4688
R67 a_n2982_13878.n47 a_n2982_13878.n114 0.365327
R68 a_n2982_13878.n28 a_n2982_13878.n46 75.0448
R69 a_n2982_13878.n45 a_n2982_13878.n28 70.1674
R70 a_n2982_13878.n116 a_n2982_13878.n45 20.9683
R71 a_n2982_13878.n30 a_n2982_13878.n44 70.3058
R72 a_n2982_13878.n44 a_n2982_13878.n109 20.6913
R73 a_n2982_13878.n43 a_n2982_13878.n30 75.3623
R74 a_n2982_13878.n117 a_n2982_13878.n43 10.5784
R75 a_n2982_13878.n29 a_n2982_13878.n31 44.7878
R76 a_n2982_13878.n20 a_n2982_13878.n58 70.1674
R77 a_n2982_13878.n58 a_n2982_13878.n96 20.9683
R78 a_n2982_13878.n57 a_n2982_13878.n21 74.73
R79 a_n2982_13878.n120 a_n2982_13878.n57 11.843
R80 a_n2982_13878.n56 a_n2982_13878.n21 80.4688
R81 a_n2982_13878.n56 a_n2982_13878.n121 0.365327
R82 a_n2982_13878.n22 a_n2982_13878.n55 75.0448
R83 a_n2982_13878.n54 a_n2982_13878.n22 70.1674
R84 a_n2982_13878.n123 a_n2982_13878.n54 20.9683
R85 a_n2982_13878.n24 a_n2982_13878.n53 70.3058
R86 a_n2982_13878.n53 a_n2982_13878.n94 20.6913
R87 a_n2982_13878.n52 a_n2982_13878.n24 75.3623
R88 a_n2982_13878.n124 a_n2982_13878.n52 10.5784
R89 a_n2982_13878.n23 a_n2982_13878.n25 44.7878
R90 a_n2982_13878.n9 a_n2982_13878.n74 70.5844
R91 a_n2982_13878.n15 a_n2982_13878.n66 70.5844
R92 a_n2982_13878.n65 a_n2982_13878.n15 70.1674
R93 a_n2982_13878.n65 a_n2982_13878.n90 20.9683
R94 a_n2982_13878.n14 a_n2982_13878.n64 74.73
R95 a_n2982_13878.n149 a_n2982_13878.n64 11.843
R96 a_n2982_13878.n63 a_n2982_13878.n14 80.4688
R97 a_n2982_13878.n63 a_n2982_13878.n91 0.365327
R98 a_n2982_13878.n16 a_n2982_13878.n62 75.0448
R99 a_n2982_13878.n61 a_n2982_13878.n16 70.1674
R100 a_n2982_13878.n61 a_n2982_13878.n92 20.9683
R101 a_n2982_13878.n17 a_n2982_13878.n60 70.3058
R102 a_n2982_13878.n146 a_n2982_13878.n60 20.6913
R103 a_n2982_13878.n59 a_n2982_13878.n17 75.3623
R104 a_n2982_13878.n59 a_n2982_13878.n93 10.5784
R105 a_n2982_13878.n19 a_n2982_13878.n18 44.7878
R106 a_n2982_13878.n73 a_n2982_13878.n9 70.1674
R107 a_n2982_13878.n73 a_n2982_13878.n86 20.9683
R108 a_n2982_13878.n8 a_n2982_13878.n72 74.73
R109 a_n2982_13878.n155 a_n2982_13878.n72 11.843
R110 a_n2982_13878.n71 a_n2982_13878.n8 80.4688
R111 a_n2982_13878.n71 a_n2982_13878.n87 0.365327
R112 a_n2982_13878.n10 a_n2982_13878.n70 75.0448
R113 a_n2982_13878.n69 a_n2982_13878.n10 70.1674
R114 a_n2982_13878.n69 a_n2982_13878.n88 20.9683
R115 a_n2982_13878.n11 a_n2982_13878.n68 70.3058
R116 a_n2982_13878.n152 a_n2982_13878.n68 20.6913
R117 a_n2982_13878.n67 a_n2982_13878.n11 75.3623
R118 a_n2982_13878.n67 a_n2982_13878.n89 10.5784
R119 a_n2982_13878.n13 a_n2982_13878.n12 44.7878
R120 a_n2982_13878.n76 a_n2982_13878.n132 20.9683
R121 a_n2982_13878.n75 a_n2982_13878.n7 75.0448
R122 a_n2982_13878.n142 a_n2982_13878.n75 11.2134
R123 a_n2982_13878.n7 a_n2982_13878.n143 161.3
R124 a_n2982_13878.n78 a_n2982_13878.n133 20.9683
R125 a_n2982_13878.n77 a_n2982_13878.n5 75.0448
R126 a_n2982_13878.n140 a_n2982_13878.n77 11.2134
R127 a_n2982_13878.n5 a_n2982_13878.n141 161.3
R128 a_n2982_13878.n80 a_n2982_13878.n134 20.9683
R129 a_n2982_13878.n79 a_n2982_13878.n3 75.0448
R130 a_n2982_13878.n138 a_n2982_13878.n79 11.2134
R131 a_n2982_13878.n3 a_n2982_13878.n139 161.3
R132 a_n2982_13878.n82 a_n2982_13878.n135 20.9683
R133 a_n2982_13878.n81 a_n2982_13878.n1 75.0448
R134 a_n2982_13878.n136 a_n2982_13878.n81 11.2134
R135 a_n2982_13878.n1 a_n2982_13878.n137 161.3
R136 a_n2982_13878.n41 a_n2982_13878.n106 81.2902
R137 a_n2982_13878.n42 a_n2982_13878.n100 81.2902
R138 a_n2982_13878.n32 a_n2982_13878.n97 81.2902
R139 a_n2982_13878.n41 a_n2982_13878.n107 80.9324
R140 a_n2982_13878.n34 a_n2982_13878.n108 80.9324
R141 a_n2982_13878.n34 a_n2982_13878.n105 80.9324
R142 a_n2982_13878.n34 a_n2982_13878.n104 80.9324
R143 a_n2982_13878.n33 a_n2982_13878.n103 80.9324
R144 a_n2982_13878.n42 a_n2982_13878.n101 80.9324
R145 a_n2982_13878.n32 a_n2982_13878.n102 80.9324
R146 a_n2982_13878.n32 a_n2982_13878.n99 80.9324
R147 a_n2982_13878.n32 a_n2982_13878.n98 80.9324
R148 a_n2982_13878.n38 a_n2982_13878.t51 74.6477
R149 a_n2982_13878.n37 a_n2982_13878.t39 74.6477
R150 a_n2982_13878.n36 a_n2982_13878.t45 74.2899
R151 a_n2982_13878.n39 a_n2982_13878.t47 74.2897
R152 a_n2982_13878.n39 a_n2982_13878.n158 70.6783
R153 a_n2982_13878.n40 a_n2982_13878.n159 70.6783
R154 a_n2982_13878.n38 a_n2982_13878.n85 70.6783
R155 a_n2982_13878.n38 a_n2982_13878.n84 70.6783
R156 a_n2982_13878.n37 a_n2982_13878.n126 70.6783
R157 a_n2982_13878.n37 a_n2982_13878.n127 70.6783
R158 a_n2982_13878.n35 a_n2982_13878.n128 70.6783
R159 a_n2982_13878.n35 a_n2982_13878.n129 70.6783
R160 a_n2982_13878.n36 a_n2982_13878.n130 70.6783
R161 a_n2982_13878.n160 a_n2982_13878.n40 70.6782
R162 a_n2982_13878.n137 a_n2982_13878.n136 48.2005
R163 a_n2982_13878.t99 a_n2982_13878.n82 533.335
R164 a_n2982_13878.n139 a_n2982_13878.n138 48.2005
R165 a_n2982_13878.t108 a_n2982_13878.n80 533.335
R166 a_n2982_13878.n141 a_n2982_13878.n140 48.2005
R167 a_n2982_13878.t93 a_n2982_13878.n78 533.335
R168 a_n2982_13878.n143 a_n2982_13878.n142 48.2005
R169 a_n2982_13878.t88 a_n2982_13878.n76 533.335
R170 a_n2982_13878.n118 a_n2982_13878.n117 48.2005
R171 a_n2982_13878.n45 a_n2982_13878.n115 20.9683
R172 a_n2982_13878.n114 a_n2982_13878.n110 48.2005
R173 a_n2982_13878.n112 a_n2982_13878.n49 20.9683
R174 a_n2982_13878.n125 a_n2982_13878.n124 48.2005
R175 a_n2982_13878.n54 a_n2982_13878.n122 20.9683
R176 a_n2982_13878.n121 a_n2982_13878.n95 48.2005
R177 a_n2982_13878.n119 a_n2982_13878.n58 20.9683
R178 a_n2982_13878.n151 a_n2982_13878.n89 48.2005
R179 a_n2982_13878.n153 a_n2982_13878.n69 20.9683
R180 a_n2982_13878.n154 a_n2982_13878.n87 48.2005
R181 a_n2982_13878.n156 a_n2982_13878.n73 20.9683
R182 a_n2982_13878.n145 a_n2982_13878.n93 48.2005
R183 a_n2982_13878.n147 a_n2982_13878.n61 20.9683
R184 a_n2982_13878.n148 a_n2982_13878.n91 48.2005
R185 a_n2982_13878.n150 a_n2982_13878.n65 20.9683
R186 a_n2982_13878.n116 a_n2982_13878.n44 21.4216
R187 a_n2982_13878.n123 a_n2982_13878.n53 21.4216
R188 a_n2982_13878.n88 a_n2982_13878.n68 21.4216
R189 a_n2982_13878.n92 a_n2982_13878.n60 21.4216
R190 a_n2982_13878.n51 a_n2982_13878.t103 532.5
R191 a_n2982_13878.n83 a_n2982_13878.t38 532.5
R192 a_n2982_13878.t46 a_n2982_13878.n74 532.5
R193 a_n2982_13878.t75 a_n2982_13878.n66 532.5
R194 a_n2982_13878.n33 a_n2982_13878.n32 31.7747
R195 a_n2982_13878.n48 a_n2982_13878.n111 34.4824
R196 a_n2982_13878.n57 a_n2982_13878.n96 34.4824
R197 a_n2982_13878.n86 a_n2982_13878.n72 34.4824
R198 a_n2982_13878.n90 a_n2982_13878.n64 34.4824
R199 a_n2982_13878.n81 a_n2982_13878.n135 35.3134
R200 a_n2982_13878.n79 a_n2982_13878.n134 35.3134
R201 a_n2982_13878.n77 a_n2982_13878.n133 35.3134
R202 a_n2982_13878.n75 a_n2982_13878.n132 35.3134
R203 a_n2982_13878.n115 a_n2982_13878.n46 35.3134
R204 a_n2982_13878.n46 a_n2982_13878.n110 11.2134
R205 a_n2982_13878.n122 a_n2982_13878.n55 35.3134
R206 a_n2982_13878.n55 a_n2982_13878.n95 11.2134
R207 a_n2982_13878.n70 a_n2982_13878.n153 35.3134
R208 a_n2982_13878.n154 a_n2982_13878.n70 11.2134
R209 a_n2982_13878.n62 a_n2982_13878.n147 35.3134
R210 a_n2982_13878.n148 a_n2982_13878.n62 11.2134
R211 a_n2982_13878.n20 a_n2982_13878.n34 23.891
R212 a_n2982_13878.n43 a_n2982_13878.n109 36.139
R213 a_n2982_13878.n52 a_n2982_13878.n94 36.139
R214 a_n2982_13878.n152 a_n2982_13878.n67 36.139
R215 a_n2982_13878.n146 a_n2982_13878.n59 36.139
R216 a_n2982_13878.n18 a_n2982_13878.n144 13.9285
R217 a_n2982_13878.n26 a_n2982_13878.n50 13.724
R218 a_n2982_13878.n131 a_n2982_13878.n23 12.4191
R219 a_n2982_13878.n144 a_n2982_13878.n7 11.2486
R220 a_n2982_13878.n0 a_n2982_13878.n50 11.2486
R221 a_n2982_13878.n39 a_n2982_13878.n157 10.5745
R222 a_n2982_13878.n157 a_n2982_13878.n9 8.58383
R223 a_n2982_13878.n131 a_n2982_13878.n36 6.7311
R224 a_n2982_13878.n157 a_n2982_13878.n50 5.3452
R225 a_n2982_13878.n20 a_n2982_13878.n29 3.94368
R226 a_n2982_13878.n12 a_n2982_13878.n15 3.94368
R227 a_n2982_13878.n158 a_n2982_13878.t37 3.61217
R228 a_n2982_13878.n158 a_n2982_13878.t65 3.61217
R229 a_n2982_13878.n159 a_n2982_13878.t49 3.61217
R230 a_n2982_13878.n159 a_n2982_13878.t59 3.61217
R231 a_n2982_13878.n85 a_n2982_13878.t25 3.61217
R232 a_n2982_13878.n85 a_n2982_13878.t57 3.61217
R233 a_n2982_13878.n84 a_n2982_13878.t53 3.61217
R234 a_n2982_13878.n84 a_n2982_13878.t29 3.61217
R235 a_n2982_13878.n126 a_n2982_13878.t35 3.61217
R236 a_n2982_13878.n126 a_n2982_13878.t27 3.61217
R237 a_n2982_13878.n127 a_n2982_13878.t43 3.61217
R238 a_n2982_13878.n127 a_n2982_13878.t63 3.61217
R239 a_n2982_13878.n128 a_n2982_13878.t31 3.61217
R240 a_n2982_13878.n128 a_n2982_13878.t67 3.61217
R241 a_n2982_13878.n129 a_n2982_13878.t41 3.61217
R242 a_n2982_13878.n129 a_n2982_13878.t23 3.61217
R243 a_n2982_13878.n130 a_n2982_13878.t33 3.61217
R244 a_n2982_13878.n130 a_n2982_13878.t61 3.61217
R245 a_n2982_13878.n160 a_n2982_13878.t55 3.61217
R246 a_n2982_13878.t21 a_n2982_13878.n160 3.61217
R247 a_n2982_13878.n106 a_n2982_13878.t19 2.82907
R248 a_n2982_13878.n106 a_n2982_13878.t8 2.82907
R249 a_n2982_13878.n107 a_n2982_13878.t18 2.82907
R250 a_n2982_13878.n107 a_n2982_13878.t10 2.82907
R251 a_n2982_13878.n108 a_n2982_13878.t1 2.82907
R252 a_n2982_13878.n108 a_n2982_13878.t68 2.82907
R253 a_n2982_13878.n105 a_n2982_13878.t16 2.82907
R254 a_n2982_13878.n105 a_n2982_13878.t11 2.82907
R255 a_n2982_13878.n104 a_n2982_13878.t2 2.82907
R256 a_n2982_13878.n104 a_n2982_13878.t6 2.82907
R257 a_n2982_13878.n103 a_n2982_13878.t9 2.82907
R258 a_n2982_13878.n103 a_n2982_13878.t70 2.82907
R259 a_n2982_13878.n100 a_n2982_13878.t7 2.82907
R260 a_n2982_13878.n100 a_n2982_13878.t0 2.82907
R261 a_n2982_13878.n101 a_n2982_13878.t71 2.82907
R262 a_n2982_13878.n101 a_n2982_13878.t14 2.82907
R263 a_n2982_13878.n102 a_n2982_13878.t17 2.82907
R264 a_n2982_13878.n102 a_n2982_13878.t13 2.82907
R265 a_n2982_13878.n99 a_n2982_13878.t12 2.82907
R266 a_n2982_13878.n99 a_n2982_13878.t3 2.82907
R267 a_n2982_13878.n98 a_n2982_13878.t5 2.82907
R268 a_n2982_13878.n98 a_n2982_13878.t4 2.82907
R269 a_n2982_13878.n97 a_n2982_13878.t69 2.82907
R270 a_n2982_13878.n97 a_n2982_13878.t15 2.82907
R271 a_n2982_13878.n31 a_n2982_13878.n118 14.1668
R272 a_n2982_13878.n112 a_n2982_13878.n51 22.3251
R273 a_n2982_13878.n25 a_n2982_13878.n125 14.1668
R274 a_n2982_13878.n119 a_n2982_13878.n83 22.3251
R275 a_n2982_13878.n151 a_n2982_13878.n13 14.1668
R276 a_n2982_13878.n74 a_n2982_13878.n156 22.3251
R277 a_n2982_13878.n145 a_n2982_13878.n19 14.1668
R278 a_n2982_13878.n66 a_n2982_13878.n150 22.3251
R279 a_n2982_13878.n144 a_n2982_13878.n131 1.30542
R280 a_n2982_13878.n4 a_n2982_13878.n3 1.04595
R281 a_n2982_13878.n47 a_n2982_13878.n113 47.835
R282 a_n2982_13878.n56 a_n2982_13878.n120 47.835
R283 a_n2982_13878.n155 a_n2982_13878.n71 47.835
R284 a_n2982_13878.n149 a_n2982_13878.n63 47.835
R285 a_n2982_13878.n27 a_n2982_13878.n26 1.13686
R286 a_n2982_13878.n15 a_n2982_13878.n14 1.13686
R287 a_n2982_13878.n9 a_n2982_13878.n8 1.13686
R288 a_n2982_13878.n21 a_n2982_13878.n20 1.09898
R289 a_n2982_13878.n40 a_n2982_13878.n38 1.07378
R290 a_n2982_13878.n36 a_n2982_13878.n35 1.07378
R291 a_n2982_13878.n32 a_n2982_13878.n42 1.07378
R292 a_n2982_13878.n30 a_n2982_13878.n29 0.758076
R293 a_n2982_13878.n30 a_n2982_13878.n28 0.758076
R294 a_n2982_13878.n28 a_n2982_13878.n27 0.758076
R295 a_n2982_13878.n24 a_n2982_13878.n23 0.758076
R296 a_n2982_13878.n24 a_n2982_13878.n22 0.758076
R297 a_n2982_13878.n22 a_n2982_13878.n21 0.758076
R298 a_n2982_13878.n17 a_n2982_13878.n18 0.758076
R299 a_n2982_13878.n16 a_n2982_13878.n17 0.758076
R300 a_n2982_13878.n14 a_n2982_13878.n16 0.758076
R301 a_n2982_13878.n11 a_n2982_13878.n12 0.758076
R302 a_n2982_13878.n10 a_n2982_13878.n11 0.758076
R303 a_n2982_13878.n8 a_n2982_13878.n10 0.758076
R304 a_n2982_13878.n7 a_n2982_13878.n6 0.758076
R305 a_n2982_13878.n5 a_n2982_13878.n4 0.758076
R306 a_n2982_13878.n3 a_n2982_13878.n2 0.758076
R307 a_n2982_13878.n1 a_n2982_13878.n0 0.758076
R308 a_n2982_13878.n34 a_n2982_13878.n41 0.716017
R309 a_n2982_13878.n40 a_n2982_13878.n39 0.716017
R310 a_n2982_13878.n35 a_n2982_13878.n37 0.716017
R311 a_n2982_13878.n34 a_n2982_13878.n33 0.716017
R312 a_n2982_13878.n6 a_n2982_13878.n5 0.67853
R313 a_n2982_13878.n2 a_n2982_13878.n1 0.67853
R314 a_n2804_13878.n29 a_n2804_13878.n28 98.9632
R315 a_n2804_13878.n2 a_n2804_13878.n0 98.7517
R316 a_n2804_13878.n22 a_n2804_13878.n21 98.6055
R317 a_n2804_13878.n24 a_n2804_13878.n23 98.6055
R318 a_n2804_13878.n26 a_n2804_13878.n25 98.6055
R319 a_n2804_13878.n28 a_n2804_13878.n27 98.6055
R320 a_n2804_13878.n10 a_n2804_13878.n9 98.6055
R321 a_n2804_13878.n8 a_n2804_13878.n7 98.6055
R322 a_n2804_13878.n6 a_n2804_13878.n5 98.6055
R323 a_n2804_13878.n4 a_n2804_13878.n3 98.6055
R324 a_n2804_13878.n2 a_n2804_13878.n1 98.6055
R325 a_n2804_13878.n20 a_n2804_13878.n19 98.6054
R326 a_n2804_13878.n12 a_n2804_13878.t30 74.6477
R327 a_n2804_13878.n17 a_n2804_13878.t31 74.2899
R328 a_n2804_13878.n14 a_n2804_13878.t1 74.2899
R329 a_n2804_13878.n13 a_n2804_13878.t5 74.2899
R330 a_n2804_13878.n16 a_n2804_13878.n15 70.6783
R331 a_n2804_13878.n12 a_n2804_13878.n11 70.6783
R332 a_n2804_13878.n18 a_n2804_13878.n10 15.7159
R333 a_n2804_13878.n20 a_n2804_13878.n18 12.6495
R334 a_n2804_13878.n18 a_n2804_13878.n17 8.38735
R335 a_n2804_13878.n19 a_n2804_13878.t13 3.61217
R336 a_n2804_13878.n19 a_n2804_13878.t22 3.61217
R337 a_n2804_13878.n21 a_n2804_13878.t26 3.61217
R338 a_n2804_13878.n21 a_n2804_13878.t12 3.61217
R339 a_n2804_13878.n23 a_n2804_13878.t16 3.61217
R340 a_n2804_13878.n23 a_n2804_13878.t17 3.61217
R341 a_n2804_13878.n25 a_n2804_13878.t27 3.61217
R342 a_n2804_13878.n25 a_n2804_13878.t28 3.61217
R343 a_n2804_13878.n27 a_n2804_13878.t6 3.61217
R344 a_n2804_13878.n27 a_n2804_13878.t18 3.61217
R345 a_n2804_13878.n15 a_n2804_13878.t2 3.61217
R346 a_n2804_13878.n15 a_n2804_13878.t0 3.61217
R347 a_n2804_13878.n11 a_n2804_13878.t3 3.61217
R348 a_n2804_13878.n11 a_n2804_13878.t4 3.61217
R349 a_n2804_13878.n9 a_n2804_13878.t19 3.61217
R350 a_n2804_13878.n9 a_n2804_13878.t7 3.61217
R351 a_n2804_13878.n7 a_n2804_13878.t24 3.61217
R352 a_n2804_13878.n7 a_n2804_13878.t9 3.61217
R353 a_n2804_13878.n5 a_n2804_13878.t8 3.61217
R354 a_n2804_13878.n5 a_n2804_13878.t11 3.61217
R355 a_n2804_13878.n3 a_n2804_13878.t21 3.61217
R356 a_n2804_13878.n3 a_n2804_13878.t14 3.61217
R357 a_n2804_13878.n1 a_n2804_13878.t25 3.61217
R358 a_n2804_13878.n1 a_n2804_13878.t15 3.61217
R359 a_n2804_13878.n0 a_n2804_13878.t10 3.61217
R360 a_n2804_13878.n0 a_n2804_13878.t20 3.61217
R361 a_n2804_13878.n29 a_n2804_13878.t23 3.61217
R362 a_n2804_13878.t29 a_n2804_13878.n29 3.61217
R363 a_n2804_13878.n13 a_n2804_13878.n12 0.358259
R364 a_n2804_13878.n16 a_n2804_13878.n14 0.358259
R365 a_n2804_13878.n17 a_n2804_13878.n16 0.358259
R366 a_n2804_13878.n28 a_n2804_13878.n26 0.358259
R367 a_n2804_13878.n26 a_n2804_13878.n24 0.358259
R368 a_n2804_13878.n24 a_n2804_13878.n22 0.358259
R369 a_n2804_13878.n22 a_n2804_13878.n20 0.358259
R370 a_n2804_13878.n4 a_n2804_13878.n2 0.146627
R371 a_n2804_13878.n6 a_n2804_13878.n4 0.146627
R372 a_n2804_13878.n8 a_n2804_13878.n6 0.146627
R373 a_n2804_13878.n10 a_n2804_13878.n8 0.146627
R374 a_n2804_13878.n14 a_n2804_13878.n13 0.101793
R375 vdd.n327 vdd.n291 756.745
R376 vdd.n268 vdd.n232 756.745
R377 vdd.n225 vdd.n189 756.745
R378 vdd.n166 vdd.n130 756.745
R379 vdd.n124 vdd.n88 756.745
R380 vdd.n65 vdd.n29 756.745
R381 vdd.n2201 vdd.n2165 756.745
R382 vdd.n2260 vdd.n2224 756.745
R383 vdd.n2099 vdd.n2063 756.745
R384 vdd.n2158 vdd.n2122 756.745
R385 vdd.n1998 vdd.n1962 756.745
R386 vdd.n2057 vdd.n2021 756.745
R387 vdd.n1315 vdd.t236 640.208
R388 vdd.n1010 vdd.t277 640.208
R389 vdd.n1319 vdd.t274 640.208
R390 vdd.n1001 vdd.t299 640.208
R391 vdd.n896 vdd.t261 640.208
R392 vdd.n2823 vdd.t292 640.208
R393 vdd.n832 vdd.t254 640.208
R394 vdd.n2820 vdd.t284 640.208
R395 vdd.n799 vdd.t232 640.208
R396 vdd.n1071 vdd.t288 640.208
R397 vdd.n1772 vdd.t302 592.009
R398 vdd.n1810 vdd.t295 592.009
R399 vdd.n1706 vdd.t305 592.009
R400 vdd.n2362 vdd.t265 592.009
R401 vdd.n1248 vdd.t240 592.009
R402 vdd.n1208 vdd.t248 592.009
R403 vdd.n426 vdd.t271 592.009
R404 vdd.n440 vdd.t244 592.009
R405 vdd.n452 vdd.t251 592.009
R406 vdd.n768 vdd.t268 592.009
R407 vdd.n3456 vdd.t281 592.009
R408 vdd.n688 vdd.t257 592.009
R409 vdd.n328 vdd.n327 585
R410 vdd.n326 vdd.n293 585
R411 vdd.n325 vdd.n324 585
R412 vdd.n296 vdd.n294 585
R413 vdd.n319 vdd.n318 585
R414 vdd.n317 vdd.n316 585
R415 vdd.n300 vdd.n299 585
R416 vdd.n311 vdd.n310 585
R417 vdd.n309 vdd.n308 585
R418 vdd.n304 vdd.n303 585
R419 vdd.n269 vdd.n268 585
R420 vdd.n267 vdd.n234 585
R421 vdd.n266 vdd.n265 585
R422 vdd.n237 vdd.n235 585
R423 vdd.n260 vdd.n259 585
R424 vdd.n258 vdd.n257 585
R425 vdd.n241 vdd.n240 585
R426 vdd.n252 vdd.n251 585
R427 vdd.n250 vdd.n249 585
R428 vdd.n245 vdd.n244 585
R429 vdd.n226 vdd.n225 585
R430 vdd.n224 vdd.n191 585
R431 vdd.n223 vdd.n222 585
R432 vdd.n194 vdd.n192 585
R433 vdd.n217 vdd.n216 585
R434 vdd.n215 vdd.n214 585
R435 vdd.n198 vdd.n197 585
R436 vdd.n209 vdd.n208 585
R437 vdd.n207 vdd.n206 585
R438 vdd.n202 vdd.n201 585
R439 vdd.n167 vdd.n166 585
R440 vdd.n165 vdd.n132 585
R441 vdd.n164 vdd.n163 585
R442 vdd.n135 vdd.n133 585
R443 vdd.n158 vdd.n157 585
R444 vdd.n156 vdd.n155 585
R445 vdd.n139 vdd.n138 585
R446 vdd.n150 vdd.n149 585
R447 vdd.n148 vdd.n147 585
R448 vdd.n143 vdd.n142 585
R449 vdd.n125 vdd.n124 585
R450 vdd.n123 vdd.n90 585
R451 vdd.n122 vdd.n121 585
R452 vdd.n93 vdd.n91 585
R453 vdd.n116 vdd.n115 585
R454 vdd.n114 vdd.n113 585
R455 vdd.n97 vdd.n96 585
R456 vdd.n108 vdd.n107 585
R457 vdd.n106 vdd.n105 585
R458 vdd.n101 vdd.n100 585
R459 vdd.n66 vdd.n65 585
R460 vdd.n64 vdd.n31 585
R461 vdd.n63 vdd.n62 585
R462 vdd.n34 vdd.n32 585
R463 vdd.n57 vdd.n56 585
R464 vdd.n55 vdd.n54 585
R465 vdd.n38 vdd.n37 585
R466 vdd.n49 vdd.n48 585
R467 vdd.n47 vdd.n46 585
R468 vdd.n42 vdd.n41 585
R469 vdd.n2202 vdd.n2201 585
R470 vdd.n2200 vdd.n2167 585
R471 vdd.n2199 vdd.n2198 585
R472 vdd.n2170 vdd.n2168 585
R473 vdd.n2193 vdd.n2192 585
R474 vdd.n2191 vdd.n2190 585
R475 vdd.n2174 vdd.n2173 585
R476 vdd.n2185 vdd.n2184 585
R477 vdd.n2183 vdd.n2182 585
R478 vdd.n2178 vdd.n2177 585
R479 vdd.n2261 vdd.n2260 585
R480 vdd.n2259 vdd.n2226 585
R481 vdd.n2258 vdd.n2257 585
R482 vdd.n2229 vdd.n2227 585
R483 vdd.n2252 vdd.n2251 585
R484 vdd.n2250 vdd.n2249 585
R485 vdd.n2233 vdd.n2232 585
R486 vdd.n2244 vdd.n2243 585
R487 vdd.n2242 vdd.n2241 585
R488 vdd.n2237 vdd.n2236 585
R489 vdd.n2100 vdd.n2099 585
R490 vdd.n2098 vdd.n2065 585
R491 vdd.n2097 vdd.n2096 585
R492 vdd.n2068 vdd.n2066 585
R493 vdd.n2091 vdd.n2090 585
R494 vdd.n2089 vdd.n2088 585
R495 vdd.n2072 vdd.n2071 585
R496 vdd.n2083 vdd.n2082 585
R497 vdd.n2081 vdd.n2080 585
R498 vdd.n2076 vdd.n2075 585
R499 vdd.n2159 vdd.n2158 585
R500 vdd.n2157 vdd.n2124 585
R501 vdd.n2156 vdd.n2155 585
R502 vdd.n2127 vdd.n2125 585
R503 vdd.n2150 vdd.n2149 585
R504 vdd.n2148 vdd.n2147 585
R505 vdd.n2131 vdd.n2130 585
R506 vdd.n2142 vdd.n2141 585
R507 vdd.n2140 vdd.n2139 585
R508 vdd.n2135 vdd.n2134 585
R509 vdd.n1999 vdd.n1998 585
R510 vdd.n1997 vdd.n1964 585
R511 vdd.n1996 vdd.n1995 585
R512 vdd.n1967 vdd.n1965 585
R513 vdd.n1990 vdd.n1989 585
R514 vdd.n1988 vdd.n1987 585
R515 vdd.n1971 vdd.n1970 585
R516 vdd.n1982 vdd.n1981 585
R517 vdd.n1980 vdd.n1979 585
R518 vdd.n1975 vdd.n1974 585
R519 vdd.n2058 vdd.n2057 585
R520 vdd.n2056 vdd.n2023 585
R521 vdd.n2055 vdd.n2054 585
R522 vdd.n2026 vdd.n2024 585
R523 vdd.n2049 vdd.n2048 585
R524 vdd.n2047 vdd.n2046 585
R525 vdd.n2030 vdd.n2029 585
R526 vdd.n2041 vdd.n2040 585
R527 vdd.n2039 vdd.n2038 585
R528 vdd.n2034 vdd.n2033 585
R529 vdd.n3628 vdd.n392 509.269
R530 vdd.n3624 vdd.n393 509.269
R531 vdd.n3496 vdd.n685 509.269
R532 vdd.n3493 vdd.n684 509.269
R533 vdd.n2357 vdd.n1530 509.269
R534 vdd.n2360 vdd.n2359 509.269
R535 vdd.n1679 vdd.n1643 509.269
R536 vdd.n1875 vdd.n1644 509.269
R537 vdd.n305 vdd.t62 329.043
R538 vdd.n246 vdd.t71 329.043
R539 vdd.n203 vdd.t198 329.043
R540 vdd.n144 vdd.t138 329.043
R541 vdd.n102 vdd.t24 329.043
R542 vdd.n43 vdd.t14 329.043
R543 vdd.n2179 vdd.t57 329.043
R544 vdd.n2238 vdd.t206 329.043
R545 vdd.n2077 vdd.t223 329.043
R546 vdd.n2136 vdd.t101 329.043
R547 vdd.n1976 vdd.t35 329.043
R548 vdd.n2035 vdd.t22 329.043
R549 vdd.n1772 vdd.t304 319.788
R550 vdd.n1810 vdd.t298 319.788
R551 vdd.n1706 vdd.t307 319.788
R552 vdd.n2362 vdd.t266 319.788
R553 vdd.n1248 vdd.t242 319.788
R554 vdd.n1208 vdd.t249 319.788
R555 vdd.n426 vdd.t272 319.788
R556 vdd.n440 vdd.t246 319.788
R557 vdd.n452 vdd.t252 319.788
R558 vdd.n768 vdd.t270 319.788
R559 vdd.n3456 vdd.t283 319.788
R560 vdd.n688 vdd.t260 319.788
R561 vdd.n1773 vdd.t303 303.69
R562 vdd.n1811 vdd.t297 303.69
R563 vdd.n1707 vdd.t306 303.69
R564 vdd.n2363 vdd.t267 303.69
R565 vdd.n1249 vdd.t243 303.69
R566 vdd.n1209 vdd.t250 303.69
R567 vdd.n427 vdd.t273 303.69
R568 vdd.n441 vdd.t247 303.69
R569 vdd.n453 vdd.t253 303.69
R570 vdd.n769 vdd.t269 303.69
R571 vdd.n3457 vdd.t282 303.69
R572 vdd.n689 vdd.t259 303.69
R573 vdd.n3090 vdd.n960 279.512
R574 vdd.n3330 vdd.n809 279.512
R575 vdd.n3267 vdd.n806 279.512
R576 vdd.n3022 vdd.n3021 279.512
R577 vdd.n2783 vdd.n998 279.512
R578 vdd.n2714 vdd.n2713 279.512
R579 vdd.n1355 vdd.n1354 279.512
R580 vdd.n2508 vdd.n1138 279.512
R581 vdd.n3246 vdd.n807 279.512
R582 vdd.n3333 vdd.n3332 279.512
R583 vdd.n2895 vdd.n2818 279.512
R584 vdd.n2826 vdd.n956 279.512
R585 vdd.n2711 vdd.n1008 279.512
R586 vdd.n1006 vdd.n980 279.512
R587 vdd.n1480 vdd.n1175 279.512
R588 vdd.n1280 vdd.n1133 279.512
R589 vdd.n2506 vdd.n1141 254.619
R590 vdd.n3495 vdd.n692 254.619
R591 vdd.n3248 vdd.n807 185
R592 vdd.n3331 vdd.n807 185
R593 vdd.n3250 vdd.n3249 185
R594 vdd.n3249 vdd.n805 185
R595 vdd.n3251 vdd.n839 185
R596 vdd.n3261 vdd.n839 185
R597 vdd.n3252 vdd.n848 185
R598 vdd.n848 vdd.n846 185
R599 vdd.n3254 vdd.n3253 185
R600 vdd.n3255 vdd.n3254 185
R601 vdd.n3207 vdd.n847 185
R602 vdd.n847 vdd.n843 185
R603 vdd.n3206 vdd.n3205 185
R604 vdd.n3205 vdd.n3204 185
R605 vdd.n850 vdd.n849 185
R606 vdd.n851 vdd.n850 185
R607 vdd.n3197 vdd.n3196 185
R608 vdd.n3198 vdd.n3197 185
R609 vdd.n3195 vdd.n859 185
R610 vdd.n864 vdd.n859 185
R611 vdd.n3194 vdd.n3193 185
R612 vdd.n3193 vdd.n3192 185
R613 vdd.n861 vdd.n860 185
R614 vdd.n870 vdd.n861 185
R615 vdd.n3185 vdd.n3184 185
R616 vdd.n3186 vdd.n3185 185
R617 vdd.n3183 vdd.n871 185
R618 vdd.n877 vdd.n871 185
R619 vdd.n3182 vdd.n3181 185
R620 vdd.n3181 vdd.n3180 185
R621 vdd.n873 vdd.n872 185
R622 vdd.n874 vdd.n873 185
R623 vdd.n3173 vdd.n3172 185
R624 vdd.n3174 vdd.n3173 185
R625 vdd.n3171 vdd.n884 185
R626 vdd.n884 vdd.n881 185
R627 vdd.n3170 vdd.n3169 185
R628 vdd.n3169 vdd.n3168 185
R629 vdd.n886 vdd.n885 185
R630 vdd.n887 vdd.n886 185
R631 vdd.n3161 vdd.n3160 185
R632 vdd.n3162 vdd.n3161 185
R633 vdd.n3159 vdd.n895 185
R634 vdd.n901 vdd.n895 185
R635 vdd.n3158 vdd.n3157 185
R636 vdd.n3157 vdd.n3156 185
R637 vdd.n3147 vdd.n898 185
R638 vdd.n908 vdd.n898 185
R639 vdd.n3149 vdd.n3148 185
R640 vdd.n3150 vdd.n3149 185
R641 vdd.n3146 vdd.n909 185
R642 vdd.n909 vdd.n905 185
R643 vdd.n3145 vdd.n3144 185
R644 vdd.n3144 vdd.n3143 185
R645 vdd.n911 vdd.n910 185
R646 vdd.n912 vdd.n911 185
R647 vdd.n3136 vdd.n3135 185
R648 vdd.n3137 vdd.n3136 185
R649 vdd.n3134 vdd.n920 185
R650 vdd.n925 vdd.n920 185
R651 vdd.n3133 vdd.n3132 185
R652 vdd.n3132 vdd.n3131 185
R653 vdd.n922 vdd.n921 185
R654 vdd.n931 vdd.n922 185
R655 vdd.n3124 vdd.n3123 185
R656 vdd.n3125 vdd.n3124 185
R657 vdd.n3122 vdd.n932 185
R658 vdd.n2998 vdd.n932 185
R659 vdd.n3121 vdd.n3120 185
R660 vdd.n3120 vdd.n3119 185
R661 vdd.n934 vdd.n933 185
R662 vdd.n3004 vdd.n934 185
R663 vdd.n3112 vdd.n3111 185
R664 vdd.n3113 vdd.n3112 185
R665 vdd.n3110 vdd.n943 185
R666 vdd.n943 vdd.n940 185
R667 vdd.n3109 vdd.n3108 185
R668 vdd.n3108 vdd.n3107 185
R669 vdd.n945 vdd.n944 185
R670 vdd.n946 vdd.n945 185
R671 vdd.n3100 vdd.n3099 185
R672 vdd.n3101 vdd.n3100 185
R673 vdd.n3098 vdd.n954 185
R674 vdd.n3016 vdd.n954 185
R675 vdd.n3097 vdd.n3096 185
R676 vdd.n3096 vdd.n3095 185
R677 vdd.n956 vdd.n955 185
R678 vdd.n957 vdd.n956 185
R679 vdd.n2827 vdd.n2826 185
R680 vdd.n2829 vdd.n2828 185
R681 vdd.n2831 vdd.n2830 185
R682 vdd.n2833 vdd.n2832 185
R683 vdd.n2835 vdd.n2834 185
R684 vdd.n2837 vdd.n2836 185
R685 vdd.n2839 vdd.n2838 185
R686 vdd.n2841 vdd.n2840 185
R687 vdd.n2843 vdd.n2842 185
R688 vdd.n2845 vdd.n2844 185
R689 vdd.n2847 vdd.n2846 185
R690 vdd.n2849 vdd.n2848 185
R691 vdd.n2851 vdd.n2850 185
R692 vdd.n2853 vdd.n2852 185
R693 vdd.n2855 vdd.n2854 185
R694 vdd.n2857 vdd.n2856 185
R695 vdd.n2859 vdd.n2858 185
R696 vdd.n2861 vdd.n2860 185
R697 vdd.n2863 vdd.n2862 185
R698 vdd.n2865 vdd.n2864 185
R699 vdd.n2867 vdd.n2866 185
R700 vdd.n2869 vdd.n2868 185
R701 vdd.n2871 vdd.n2870 185
R702 vdd.n2873 vdd.n2872 185
R703 vdd.n2875 vdd.n2874 185
R704 vdd.n2877 vdd.n2876 185
R705 vdd.n2879 vdd.n2878 185
R706 vdd.n2881 vdd.n2880 185
R707 vdd.n2883 vdd.n2882 185
R708 vdd.n2885 vdd.n2884 185
R709 vdd.n2887 vdd.n2886 185
R710 vdd.n2889 vdd.n2888 185
R711 vdd.n2891 vdd.n2890 185
R712 vdd.n2893 vdd.n2892 185
R713 vdd.n2894 vdd.n2818 185
R714 vdd.n3088 vdd.n2818 185
R715 vdd.n3334 vdd.n3333 185
R716 vdd.n3335 vdd.n798 185
R717 vdd.n3337 vdd.n3336 185
R718 vdd.n3339 vdd.n796 185
R719 vdd.n3341 vdd.n3340 185
R720 vdd.n3342 vdd.n795 185
R721 vdd.n3344 vdd.n3343 185
R722 vdd.n3346 vdd.n793 185
R723 vdd.n3348 vdd.n3347 185
R724 vdd.n3349 vdd.n792 185
R725 vdd.n3351 vdd.n3350 185
R726 vdd.n3353 vdd.n790 185
R727 vdd.n3355 vdd.n3354 185
R728 vdd.n3356 vdd.n789 185
R729 vdd.n3358 vdd.n3357 185
R730 vdd.n3360 vdd.n788 185
R731 vdd.n3361 vdd.n786 185
R732 vdd.n3364 vdd.n3363 185
R733 vdd.n787 vdd.n785 185
R734 vdd.n3220 vdd.n3219 185
R735 vdd.n3222 vdd.n3221 185
R736 vdd.n3224 vdd.n3216 185
R737 vdd.n3226 vdd.n3225 185
R738 vdd.n3227 vdd.n3215 185
R739 vdd.n3229 vdd.n3228 185
R740 vdd.n3231 vdd.n3213 185
R741 vdd.n3233 vdd.n3232 185
R742 vdd.n3234 vdd.n3212 185
R743 vdd.n3236 vdd.n3235 185
R744 vdd.n3238 vdd.n3210 185
R745 vdd.n3240 vdd.n3239 185
R746 vdd.n3241 vdd.n3209 185
R747 vdd.n3243 vdd.n3242 185
R748 vdd.n3245 vdd.n3208 185
R749 vdd.n3247 vdd.n3246 185
R750 vdd.n3246 vdd.n692 185
R751 vdd.n3332 vdd.n802 185
R752 vdd.n3332 vdd.n3331 185
R753 vdd.n2949 vdd.n804 185
R754 vdd.n805 vdd.n804 185
R755 vdd.n2950 vdd.n838 185
R756 vdd.n3261 vdd.n838 185
R757 vdd.n2952 vdd.n2951 185
R758 vdd.n2951 vdd.n846 185
R759 vdd.n2953 vdd.n845 185
R760 vdd.n3255 vdd.n845 185
R761 vdd.n2955 vdd.n2954 185
R762 vdd.n2954 vdd.n843 185
R763 vdd.n2956 vdd.n853 185
R764 vdd.n3204 vdd.n853 185
R765 vdd.n2958 vdd.n2957 185
R766 vdd.n2957 vdd.n851 185
R767 vdd.n2959 vdd.n858 185
R768 vdd.n3198 vdd.n858 185
R769 vdd.n2961 vdd.n2960 185
R770 vdd.n2960 vdd.n864 185
R771 vdd.n2962 vdd.n863 185
R772 vdd.n3192 vdd.n863 185
R773 vdd.n2964 vdd.n2963 185
R774 vdd.n2963 vdd.n870 185
R775 vdd.n2965 vdd.n869 185
R776 vdd.n3186 vdd.n869 185
R777 vdd.n2967 vdd.n2966 185
R778 vdd.n2966 vdd.n877 185
R779 vdd.n2968 vdd.n876 185
R780 vdd.n3180 vdd.n876 185
R781 vdd.n2970 vdd.n2969 185
R782 vdd.n2969 vdd.n874 185
R783 vdd.n2971 vdd.n883 185
R784 vdd.n3174 vdd.n883 185
R785 vdd.n2973 vdd.n2972 185
R786 vdd.n2972 vdd.n881 185
R787 vdd.n2974 vdd.n889 185
R788 vdd.n3168 vdd.n889 185
R789 vdd.n2976 vdd.n2975 185
R790 vdd.n2975 vdd.n887 185
R791 vdd.n2977 vdd.n894 185
R792 vdd.n3162 vdd.n894 185
R793 vdd.n2979 vdd.n2978 185
R794 vdd.n2978 vdd.n901 185
R795 vdd.n2980 vdd.n900 185
R796 vdd.n3156 vdd.n900 185
R797 vdd.n2982 vdd.n2981 185
R798 vdd.n2981 vdd.n908 185
R799 vdd.n2983 vdd.n907 185
R800 vdd.n3150 vdd.n907 185
R801 vdd.n2985 vdd.n2984 185
R802 vdd.n2984 vdd.n905 185
R803 vdd.n2986 vdd.n914 185
R804 vdd.n3143 vdd.n914 185
R805 vdd.n2988 vdd.n2987 185
R806 vdd.n2987 vdd.n912 185
R807 vdd.n2989 vdd.n919 185
R808 vdd.n3137 vdd.n919 185
R809 vdd.n2991 vdd.n2990 185
R810 vdd.n2990 vdd.n925 185
R811 vdd.n2992 vdd.n924 185
R812 vdd.n3131 vdd.n924 185
R813 vdd.n2994 vdd.n2993 185
R814 vdd.n2993 vdd.n931 185
R815 vdd.n2995 vdd.n930 185
R816 vdd.n3125 vdd.n930 185
R817 vdd.n2997 vdd.n2996 185
R818 vdd.n2998 vdd.n2997 185
R819 vdd.n2898 vdd.n936 185
R820 vdd.n3119 vdd.n936 185
R821 vdd.n3006 vdd.n3005 185
R822 vdd.n3005 vdd.n3004 185
R823 vdd.n3007 vdd.n942 185
R824 vdd.n3113 vdd.n942 185
R825 vdd.n3009 vdd.n3008 185
R826 vdd.n3008 vdd.n940 185
R827 vdd.n3010 vdd.n948 185
R828 vdd.n3107 vdd.n948 185
R829 vdd.n3012 vdd.n3011 185
R830 vdd.n3011 vdd.n946 185
R831 vdd.n3013 vdd.n953 185
R832 vdd.n3101 vdd.n953 185
R833 vdd.n3015 vdd.n3014 185
R834 vdd.n3016 vdd.n3015 185
R835 vdd.n2897 vdd.n959 185
R836 vdd.n3095 vdd.n959 185
R837 vdd.n2896 vdd.n2895 185
R838 vdd.n2895 vdd.n957 185
R839 vdd.n2357 vdd.n2356 185
R840 vdd.n2358 vdd.n2357 185
R841 vdd.n1531 vdd.n1529 185
R842 vdd.n2349 vdd.n1529 185
R843 vdd.n2352 vdd.n2351 185
R844 vdd.n2351 vdd.n2350 185
R845 vdd.n1534 vdd.n1533 185
R846 vdd.n1535 vdd.n1534 185
R847 vdd.n2338 vdd.n2337 185
R848 vdd.n2339 vdd.n2338 185
R849 vdd.n1543 vdd.n1542 185
R850 vdd.n2330 vdd.n1542 185
R851 vdd.n2333 vdd.n2332 185
R852 vdd.n2332 vdd.n2331 185
R853 vdd.n1546 vdd.n1545 185
R854 vdd.n1553 vdd.n1546 185
R855 vdd.n2321 vdd.n2320 185
R856 vdd.n2322 vdd.n2321 185
R857 vdd.n1555 vdd.n1554 185
R858 vdd.n1554 vdd.n1552 185
R859 vdd.n2316 vdd.n2315 185
R860 vdd.n2315 vdd.n2314 185
R861 vdd.n1558 vdd.n1557 185
R862 vdd.n1559 vdd.n1558 185
R863 vdd.n2305 vdd.n2304 185
R864 vdd.n2306 vdd.n2305 185
R865 vdd.n1566 vdd.n1565 185
R866 vdd.n2297 vdd.n1565 185
R867 vdd.n2300 vdd.n2299 185
R868 vdd.n2299 vdd.n2298 185
R869 vdd.n1569 vdd.n1568 185
R870 vdd.n1575 vdd.n1569 185
R871 vdd.n2288 vdd.n2287 185
R872 vdd.n2289 vdd.n2288 185
R873 vdd.n1577 vdd.n1576 185
R874 vdd.n2280 vdd.n1576 185
R875 vdd.n2283 vdd.n2282 185
R876 vdd.n2282 vdd.n2281 185
R877 vdd.n1580 vdd.n1579 185
R878 vdd.n1581 vdd.n1580 185
R879 vdd.n2271 vdd.n2270 185
R880 vdd.n2272 vdd.n2271 185
R881 vdd.n1589 vdd.n1588 185
R882 vdd.n1588 vdd.n1587 185
R883 vdd.n1959 vdd.n1958 185
R884 vdd.n1958 vdd.n1957 185
R885 vdd.n1592 vdd.n1591 185
R886 vdd.n1598 vdd.n1592 185
R887 vdd.n1948 vdd.n1947 185
R888 vdd.n1949 vdd.n1948 185
R889 vdd.n1600 vdd.n1599 185
R890 vdd.n1940 vdd.n1599 185
R891 vdd.n1943 vdd.n1942 185
R892 vdd.n1942 vdd.n1941 185
R893 vdd.n1603 vdd.n1602 185
R894 vdd.n1610 vdd.n1603 185
R895 vdd.n1931 vdd.n1930 185
R896 vdd.n1932 vdd.n1931 185
R897 vdd.n1612 vdd.n1611 185
R898 vdd.n1611 vdd.n1609 185
R899 vdd.n1926 vdd.n1925 185
R900 vdd.n1925 vdd.n1924 185
R901 vdd.n1615 vdd.n1614 185
R902 vdd.n1616 vdd.n1615 185
R903 vdd.n1915 vdd.n1914 185
R904 vdd.n1916 vdd.n1915 185
R905 vdd.n1623 vdd.n1622 185
R906 vdd.n1907 vdd.n1622 185
R907 vdd.n1910 vdd.n1909 185
R908 vdd.n1909 vdd.n1908 185
R909 vdd.n1626 vdd.n1625 185
R910 vdd.n1632 vdd.n1626 185
R911 vdd.n1898 vdd.n1897 185
R912 vdd.n1899 vdd.n1898 185
R913 vdd.n1634 vdd.n1633 185
R914 vdd.n1890 vdd.n1633 185
R915 vdd.n1893 vdd.n1892 185
R916 vdd.n1892 vdd.n1891 185
R917 vdd.n1637 vdd.n1636 185
R918 vdd.n1638 vdd.n1637 185
R919 vdd.n1881 vdd.n1880 185
R920 vdd.n1882 vdd.n1881 185
R921 vdd.n1645 vdd.n1644 185
R922 vdd.n1680 vdd.n1644 185
R923 vdd.n1876 vdd.n1875 185
R924 vdd.n1648 vdd.n1647 185
R925 vdd.n1872 vdd.n1871 185
R926 vdd.n1873 vdd.n1872 185
R927 vdd.n1682 vdd.n1681 185
R928 vdd.n1867 vdd.n1684 185
R929 vdd.n1866 vdd.n1685 185
R930 vdd.n1865 vdd.n1686 185
R931 vdd.n1688 vdd.n1687 185
R932 vdd.n1861 vdd.n1690 185
R933 vdd.n1860 vdd.n1691 185
R934 vdd.n1859 vdd.n1692 185
R935 vdd.n1694 vdd.n1693 185
R936 vdd.n1855 vdd.n1696 185
R937 vdd.n1854 vdd.n1697 185
R938 vdd.n1853 vdd.n1698 185
R939 vdd.n1700 vdd.n1699 185
R940 vdd.n1849 vdd.n1702 185
R941 vdd.n1848 vdd.n1703 185
R942 vdd.n1847 vdd.n1704 185
R943 vdd.n1708 vdd.n1705 185
R944 vdd.n1843 vdd.n1710 185
R945 vdd.n1842 vdd.n1711 185
R946 vdd.n1841 vdd.n1712 185
R947 vdd.n1714 vdd.n1713 185
R948 vdd.n1837 vdd.n1716 185
R949 vdd.n1836 vdd.n1717 185
R950 vdd.n1835 vdd.n1718 185
R951 vdd.n1720 vdd.n1719 185
R952 vdd.n1831 vdd.n1722 185
R953 vdd.n1830 vdd.n1723 185
R954 vdd.n1829 vdd.n1724 185
R955 vdd.n1726 vdd.n1725 185
R956 vdd.n1825 vdd.n1728 185
R957 vdd.n1824 vdd.n1729 185
R958 vdd.n1823 vdd.n1730 185
R959 vdd.n1732 vdd.n1731 185
R960 vdd.n1819 vdd.n1734 185
R961 vdd.n1818 vdd.n1735 185
R962 vdd.n1817 vdd.n1736 185
R963 vdd.n1738 vdd.n1737 185
R964 vdd.n1813 vdd.n1740 185
R965 vdd.n1812 vdd.n1809 185
R966 vdd.n1808 vdd.n1741 185
R967 vdd.n1743 vdd.n1742 185
R968 vdd.n1804 vdd.n1745 185
R969 vdd.n1803 vdd.n1746 185
R970 vdd.n1802 vdd.n1747 185
R971 vdd.n1749 vdd.n1748 185
R972 vdd.n1798 vdd.n1751 185
R973 vdd.n1797 vdd.n1752 185
R974 vdd.n1796 vdd.n1753 185
R975 vdd.n1755 vdd.n1754 185
R976 vdd.n1792 vdd.n1757 185
R977 vdd.n1791 vdd.n1758 185
R978 vdd.n1790 vdd.n1759 185
R979 vdd.n1761 vdd.n1760 185
R980 vdd.n1786 vdd.n1763 185
R981 vdd.n1785 vdd.n1764 185
R982 vdd.n1784 vdd.n1765 185
R983 vdd.n1767 vdd.n1766 185
R984 vdd.n1780 vdd.n1769 185
R985 vdd.n1779 vdd.n1770 185
R986 vdd.n1778 vdd.n1771 185
R987 vdd.n1775 vdd.n1679 185
R988 vdd.n1873 vdd.n1679 185
R989 vdd.n2361 vdd.n2360 185
R990 vdd.n2365 vdd.n1525 185
R991 vdd.n1524 vdd.n1518 185
R992 vdd.n1522 vdd.n1521 185
R993 vdd.n1520 vdd.n1279 185
R994 vdd.n2369 vdd.n1276 185
R995 vdd.n2371 vdd.n2370 185
R996 vdd.n2373 vdd.n1274 185
R997 vdd.n2375 vdd.n2374 185
R998 vdd.n2376 vdd.n1269 185
R999 vdd.n2378 vdd.n2377 185
R1000 vdd.n2380 vdd.n1267 185
R1001 vdd.n2382 vdd.n2381 185
R1002 vdd.n2383 vdd.n1262 185
R1003 vdd.n2385 vdd.n2384 185
R1004 vdd.n2387 vdd.n1260 185
R1005 vdd.n2389 vdd.n2388 185
R1006 vdd.n2390 vdd.n1256 185
R1007 vdd.n2392 vdd.n2391 185
R1008 vdd.n2394 vdd.n1253 185
R1009 vdd.n2396 vdd.n2395 185
R1010 vdd.n1254 vdd.n1247 185
R1011 vdd.n2400 vdd.n1251 185
R1012 vdd.n2401 vdd.n1243 185
R1013 vdd.n2403 vdd.n2402 185
R1014 vdd.n2405 vdd.n1241 185
R1015 vdd.n2407 vdd.n2406 185
R1016 vdd.n2408 vdd.n1236 185
R1017 vdd.n2410 vdd.n2409 185
R1018 vdd.n2412 vdd.n1234 185
R1019 vdd.n2414 vdd.n2413 185
R1020 vdd.n2415 vdd.n1229 185
R1021 vdd.n2417 vdd.n2416 185
R1022 vdd.n2419 vdd.n1227 185
R1023 vdd.n2421 vdd.n2420 185
R1024 vdd.n2422 vdd.n1222 185
R1025 vdd.n2424 vdd.n2423 185
R1026 vdd.n2426 vdd.n1220 185
R1027 vdd.n2428 vdd.n2427 185
R1028 vdd.n2429 vdd.n1216 185
R1029 vdd.n2431 vdd.n2430 185
R1030 vdd.n2433 vdd.n1213 185
R1031 vdd.n2435 vdd.n2434 185
R1032 vdd.n1214 vdd.n1207 185
R1033 vdd.n2439 vdd.n1211 185
R1034 vdd.n2440 vdd.n1203 185
R1035 vdd.n2442 vdd.n2441 185
R1036 vdd.n2444 vdd.n1201 185
R1037 vdd.n2446 vdd.n2445 185
R1038 vdd.n2447 vdd.n1196 185
R1039 vdd.n2449 vdd.n2448 185
R1040 vdd.n2451 vdd.n1194 185
R1041 vdd.n2453 vdd.n2452 185
R1042 vdd.n2454 vdd.n1189 185
R1043 vdd.n2456 vdd.n2455 185
R1044 vdd.n2458 vdd.n1187 185
R1045 vdd.n2460 vdd.n2459 185
R1046 vdd.n2461 vdd.n1185 185
R1047 vdd.n2463 vdd.n2462 185
R1048 vdd.n2466 vdd.n2465 185
R1049 vdd.n2468 vdd.n2467 185
R1050 vdd.n2470 vdd.n1183 185
R1051 vdd.n2472 vdd.n2471 185
R1052 vdd.n1530 vdd.n1182 185
R1053 vdd.n2359 vdd.n1528 185
R1054 vdd.n2359 vdd.n2358 185
R1055 vdd.n1538 vdd.n1527 185
R1056 vdd.n2349 vdd.n1527 185
R1057 vdd.n2348 vdd.n2347 185
R1058 vdd.n2350 vdd.n2348 185
R1059 vdd.n1537 vdd.n1536 185
R1060 vdd.n1536 vdd.n1535 185
R1061 vdd.n2341 vdd.n2340 185
R1062 vdd.n2340 vdd.n2339 185
R1063 vdd.n1541 vdd.n1540 185
R1064 vdd.n2330 vdd.n1541 185
R1065 vdd.n2329 vdd.n2328 185
R1066 vdd.n2331 vdd.n2329 185
R1067 vdd.n1548 vdd.n1547 185
R1068 vdd.n1553 vdd.n1547 185
R1069 vdd.n2324 vdd.n2323 185
R1070 vdd.n2323 vdd.n2322 185
R1071 vdd.n1551 vdd.n1550 185
R1072 vdd.n1552 vdd.n1551 185
R1073 vdd.n2313 vdd.n2312 185
R1074 vdd.n2314 vdd.n2313 185
R1075 vdd.n1561 vdd.n1560 185
R1076 vdd.n1560 vdd.n1559 185
R1077 vdd.n2308 vdd.n2307 185
R1078 vdd.n2307 vdd.n2306 185
R1079 vdd.n1564 vdd.n1563 185
R1080 vdd.n2297 vdd.n1564 185
R1081 vdd.n2296 vdd.n2295 185
R1082 vdd.n2298 vdd.n2296 185
R1083 vdd.n1571 vdd.n1570 185
R1084 vdd.n1575 vdd.n1570 185
R1085 vdd.n2291 vdd.n2290 185
R1086 vdd.n2290 vdd.n2289 185
R1087 vdd.n1574 vdd.n1573 185
R1088 vdd.n2280 vdd.n1574 185
R1089 vdd.n2279 vdd.n2278 185
R1090 vdd.n2281 vdd.n2279 185
R1091 vdd.n1583 vdd.n1582 185
R1092 vdd.n1582 vdd.n1581 185
R1093 vdd.n2274 vdd.n2273 185
R1094 vdd.n2273 vdd.n2272 185
R1095 vdd.n1586 vdd.n1585 185
R1096 vdd.n1587 vdd.n1586 185
R1097 vdd.n1956 vdd.n1955 185
R1098 vdd.n1957 vdd.n1956 185
R1099 vdd.n1594 vdd.n1593 185
R1100 vdd.n1598 vdd.n1593 185
R1101 vdd.n1951 vdd.n1950 185
R1102 vdd.n1950 vdd.n1949 185
R1103 vdd.n1597 vdd.n1596 185
R1104 vdd.n1940 vdd.n1597 185
R1105 vdd.n1939 vdd.n1938 185
R1106 vdd.n1941 vdd.n1939 185
R1107 vdd.n1605 vdd.n1604 185
R1108 vdd.n1610 vdd.n1604 185
R1109 vdd.n1934 vdd.n1933 185
R1110 vdd.n1933 vdd.n1932 185
R1111 vdd.n1608 vdd.n1607 185
R1112 vdd.n1609 vdd.n1608 185
R1113 vdd.n1923 vdd.n1922 185
R1114 vdd.n1924 vdd.n1923 185
R1115 vdd.n1618 vdd.n1617 185
R1116 vdd.n1617 vdd.n1616 185
R1117 vdd.n1918 vdd.n1917 185
R1118 vdd.n1917 vdd.n1916 185
R1119 vdd.n1621 vdd.n1620 185
R1120 vdd.n1907 vdd.n1621 185
R1121 vdd.n1906 vdd.n1905 185
R1122 vdd.n1908 vdd.n1906 185
R1123 vdd.n1628 vdd.n1627 185
R1124 vdd.n1632 vdd.n1627 185
R1125 vdd.n1901 vdd.n1900 185
R1126 vdd.n1900 vdd.n1899 185
R1127 vdd.n1631 vdd.n1630 185
R1128 vdd.n1890 vdd.n1631 185
R1129 vdd.n1889 vdd.n1888 185
R1130 vdd.n1891 vdd.n1889 185
R1131 vdd.n1640 vdd.n1639 185
R1132 vdd.n1639 vdd.n1638 185
R1133 vdd.n1884 vdd.n1883 185
R1134 vdd.n1883 vdd.n1882 185
R1135 vdd.n1643 vdd.n1642 185
R1136 vdd.n1680 vdd.n1643 185
R1137 vdd.n1000 vdd.n998 185
R1138 vdd.n2712 vdd.n998 185
R1139 vdd.n2634 vdd.n1018 185
R1140 vdd.n1018 vdd.n1005 185
R1141 vdd.n2636 vdd.n2635 185
R1142 vdd.n2637 vdd.n2636 185
R1143 vdd.n2633 vdd.n1017 185
R1144 vdd.n1399 vdd.n1017 185
R1145 vdd.n2632 vdd.n2631 185
R1146 vdd.n2631 vdd.n2630 185
R1147 vdd.n1020 vdd.n1019 185
R1148 vdd.n1021 vdd.n1020 185
R1149 vdd.n2621 vdd.n2620 185
R1150 vdd.n2622 vdd.n2621 185
R1151 vdd.n2619 vdd.n1031 185
R1152 vdd.n1031 vdd.n1028 185
R1153 vdd.n2618 vdd.n2617 185
R1154 vdd.n2617 vdd.n2616 185
R1155 vdd.n1033 vdd.n1032 185
R1156 vdd.n1425 vdd.n1033 185
R1157 vdd.n2609 vdd.n2608 185
R1158 vdd.n2610 vdd.n2609 185
R1159 vdd.n2607 vdd.n1041 185
R1160 vdd.n1046 vdd.n1041 185
R1161 vdd.n2606 vdd.n2605 185
R1162 vdd.n2605 vdd.n2604 185
R1163 vdd.n1043 vdd.n1042 185
R1164 vdd.n1052 vdd.n1043 185
R1165 vdd.n2597 vdd.n2596 185
R1166 vdd.n2598 vdd.n2597 185
R1167 vdd.n2595 vdd.n1053 185
R1168 vdd.n1437 vdd.n1053 185
R1169 vdd.n2594 vdd.n2593 185
R1170 vdd.n2593 vdd.n2592 185
R1171 vdd.n1055 vdd.n1054 185
R1172 vdd.n1056 vdd.n1055 185
R1173 vdd.n2585 vdd.n2584 185
R1174 vdd.n2586 vdd.n2585 185
R1175 vdd.n2583 vdd.n1065 185
R1176 vdd.n1065 vdd.n1062 185
R1177 vdd.n2582 vdd.n2581 185
R1178 vdd.n2581 vdd.n2580 185
R1179 vdd.n1067 vdd.n1066 185
R1180 vdd.n1076 vdd.n1067 185
R1181 vdd.n2572 vdd.n2571 185
R1182 vdd.n2573 vdd.n2572 185
R1183 vdd.n2570 vdd.n1077 185
R1184 vdd.n1083 vdd.n1077 185
R1185 vdd.n2569 vdd.n2568 185
R1186 vdd.n2568 vdd.n2567 185
R1187 vdd.n1079 vdd.n1078 185
R1188 vdd.n1080 vdd.n1079 185
R1189 vdd.n2560 vdd.n2559 185
R1190 vdd.n2561 vdd.n2560 185
R1191 vdd.n2558 vdd.n1090 185
R1192 vdd.n1090 vdd.n1087 185
R1193 vdd.n2557 vdd.n2556 185
R1194 vdd.n2556 vdd.n2555 185
R1195 vdd.n1092 vdd.n1091 185
R1196 vdd.n1093 vdd.n1092 185
R1197 vdd.n2548 vdd.n2547 185
R1198 vdd.n2549 vdd.n2548 185
R1199 vdd.n2546 vdd.n1101 185
R1200 vdd.n1106 vdd.n1101 185
R1201 vdd.n2545 vdd.n2544 185
R1202 vdd.n2544 vdd.n2543 185
R1203 vdd.n1103 vdd.n1102 185
R1204 vdd.n1112 vdd.n1103 185
R1205 vdd.n2536 vdd.n2535 185
R1206 vdd.n2537 vdd.n2536 185
R1207 vdd.n2534 vdd.n1113 185
R1208 vdd.n1119 vdd.n1113 185
R1209 vdd.n2533 vdd.n2532 185
R1210 vdd.n2532 vdd.n2531 185
R1211 vdd.n1115 vdd.n1114 185
R1212 vdd.n1116 vdd.n1115 185
R1213 vdd.n2524 vdd.n2523 185
R1214 vdd.n2525 vdd.n2524 185
R1215 vdd.n2522 vdd.n1126 185
R1216 vdd.n1126 vdd.n1123 185
R1217 vdd.n2521 vdd.n2520 185
R1218 vdd.n2520 vdd.n2519 185
R1219 vdd.n1128 vdd.n1127 185
R1220 vdd.n1137 vdd.n1128 185
R1221 vdd.n2512 vdd.n2511 185
R1222 vdd.n2513 vdd.n2512 185
R1223 vdd.n2510 vdd.n1138 185
R1224 vdd.n1138 vdd.n1134 185
R1225 vdd.n2509 vdd.n2508 185
R1226 vdd.n1140 vdd.n1139 185
R1227 vdd.n2505 vdd.n2504 185
R1228 vdd.n2506 vdd.n2505 185
R1229 vdd.n2503 vdd.n1176 185
R1230 vdd.n2502 vdd.n2501 185
R1231 vdd.n2500 vdd.n2499 185
R1232 vdd.n2498 vdd.n2497 185
R1233 vdd.n2496 vdd.n2495 185
R1234 vdd.n2494 vdd.n2493 185
R1235 vdd.n2492 vdd.n2491 185
R1236 vdd.n2490 vdd.n2489 185
R1237 vdd.n2488 vdd.n2487 185
R1238 vdd.n2486 vdd.n2485 185
R1239 vdd.n2484 vdd.n2483 185
R1240 vdd.n2482 vdd.n2481 185
R1241 vdd.n2480 vdd.n2479 185
R1242 vdd.n2478 vdd.n2477 185
R1243 vdd.n2476 vdd.n2475 185
R1244 vdd.n1321 vdd.n1177 185
R1245 vdd.n1323 vdd.n1322 185
R1246 vdd.n1325 vdd.n1324 185
R1247 vdd.n1327 vdd.n1326 185
R1248 vdd.n1329 vdd.n1328 185
R1249 vdd.n1331 vdd.n1330 185
R1250 vdd.n1333 vdd.n1332 185
R1251 vdd.n1335 vdd.n1334 185
R1252 vdd.n1337 vdd.n1336 185
R1253 vdd.n1339 vdd.n1338 185
R1254 vdd.n1341 vdd.n1340 185
R1255 vdd.n1343 vdd.n1342 185
R1256 vdd.n1345 vdd.n1344 185
R1257 vdd.n1347 vdd.n1346 185
R1258 vdd.n1350 vdd.n1349 185
R1259 vdd.n1352 vdd.n1351 185
R1260 vdd.n1354 vdd.n1353 185
R1261 vdd.n2715 vdd.n2714 185
R1262 vdd.n2717 vdd.n2716 185
R1263 vdd.n2719 vdd.n2718 185
R1264 vdd.n2722 vdd.n2721 185
R1265 vdd.n2724 vdd.n2723 185
R1266 vdd.n2726 vdd.n2725 185
R1267 vdd.n2728 vdd.n2727 185
R1268 vdd.n2730 vdd.n2729 185
R1269 vdd.n2732 vdd.n2731 185
R1270 vdd.n2734 vdd.n2733 185
R1271 vdd.n2736 vdd.n2735 185
R1272 vdd.n2738 vdd.n2737 185
R1273 vdd.n2740 vdd.n2739 185
R1274 vdd.n2742 vdd.n2741 185
R1275 vdd.n2744 vdd.n2743 185
R1276 vdd.n2746 vdd.n2745 185
R1277 vdd.n2748 vdd.n2747 185
R1278 vdd.n2750 vdd.n2749 185
R1279 vdd.n2752 vdd.n2751 185
R1280 vdd.n2754 vdd.n2753 185
R1281 vdd.n2756 vdd.n2755 185
R1282 vdd.n2758 vdd.n2757 185
R1283 vdd.n2760 vdd.n2759 185
R1284 vdd.n2762 vdd.n2761 185
R1285 vdd.n2764 vdd.n2763 185
R1286 vdd.n2766 vdd.n2765 185
R1287 vdd.n2768 vdd.n2767 185
R1288 vdd.n2770 vdd.n2769 185
R1289 vdd.n2772 vdd.n2771 185
R1290 vdd.n2774 vdd.n2773 185
R1291 vdd.n2776 vdd.n2775 185
R1292 vdd.n2778 vdd.n2777 185
R1293 vdd.n2780 vdd.n2779 185
R1294 vdd.n2781 vdd.n999 185
R1295 vdd.n2783 vdd.n2782 185
R1296 vdd.n2784 vdd.n2783 185
R1297 vdd.n2713 vdd.n1003 185
R1298 vdd.n2713 vdd.n2712 185
R1299 vdd.n1397 vdd.n1004 185
R1300 vdd.n1005 vdd.n1004 185
R1301 vdd.n1398 vdd.n1015 185
R1302 vdd.n2637 vdd.n1015 185
R1303 vdd.n1401 vdd.n1400 185
R1304 vdd.n1400 vdd.n1399 185
R1305 vdd.n1402 vdd.n1022 185
R1306 vdd.n2630 vdd.n1022 185
R1307 vdd.n1404 vdd.n1403 185
R1308 vdd.n1403 vdd.n1021 185
R1309 vdd.n1405 vdd.n1029 185
R1310 vdd.n2622 vdd.n1029 185
R1311 vdd.n1407 vdd.n1406 185
R1312 vdd.n1406 vdd.n1028 185
R1313 vdd.n1408 vdd.n1034 185
R1314 vdd.n2616 vdd.n1034 185
R1315 vdd.n1427 vdd.n1426 185
R1316 vdd.n1426 vdd.n1425 185
R1317 vdd.n1428 vdd.n1039 185
R1318 vdd.n2610 vdd.n1039 185
R1319 vdd.n1430 vdd.n1429 185
R1320 vdd.n1429 vdd.n1046 185
R1321 vdd.n1431 vdd.n1044 185
R1322 vdd.n2604 vdd.n1044 185
R1323 vdd.n1433 vdd.n1432 185
R1324 vdd.n1432 vdd.n1052 185
R1325 vdd.n1434 vdd.n1050 185
R1326 vdd.n2598 vdd.n1050 185
R1327 vdd.n1436 vdd.n1435 185
R1328 vdd.n1437 vdd.n1436 185
R1329 vdd.n1396 vdd.n1057 185
R1330 vdd.n2592 vdd.n1057 185
R1331 vdd.n1395 vdd.n1394 185
R1332 vdd.n1394 vdd.n1056 185
R1333 vdd.n1393 vdd.n1063 185
R1334 vdd.n2586 vdd.n1063 185
R1335 vdd.n1392 vdd.n1391 185
R1336 vdd.n1391 vdd.n1062 185
R1337 vdd.n1390 vdd.n1068 185
R1338 vdd.n2580 vdd.n1068 185
R1339 vdd.n1389 vdd.n1388 185
R1340 vdd.n1388 vdd.n1076 185
R1341 vdd.n1387 vdd.n1074 185
R1342 vdd.n2573 vdd.n1074 185
R1343 vdd.n1386 vdd.n1385 185
R1344 vdd.n1385 vdd.n1083 185
R1345 vdd.n1384 vdd.n1081 185
R1346 vdd.n2567 vdd.n1081 185
R1347 vdd.n1383 vdd.n1382 185
R1348 vdd.n1382 vdd.n1080 185
R1349 vdd.n1381 vdd.n1088 185
R1350 vdd.n2561 vdd.n1088 185
R1351 vdd.n1380 vdd.n1379 185
R1352 vdd.n1379 vdd.n1087 185
R1353 vdd.n1378 vdd.n1094 185
R1354 vdd.n2555 vdd.n1094 185
R1355 vdd.n1377 vdd.n1376 185
R1356 vdd.n1376 vdd.n1093 185
R1357 vdd.n1375 vdd.n1099 185
R1358 vdd.n2549 vdd.n1099 185
R1359 vdd.n1374 vdd.n1373 185
R1360 vdd.n1373 vdd.n1106 185
R1361 vdd.n1372 vdd.n1104 185
R1362 vdd.n2543 vdd.n1104 185
R1363 vdd.n1371 vdd.n1370 185
R1364 vdd.n1370 vdd.n1112 185
R1365 vdd.n1369 vdd.n1110 185
R1366 vdd.n2537 vdd.n1110 185
R1367 vdd.n1368 vdd.n1367 185
R1368 vdd.n1367 vdd.n1119 185
R1369 vdd.n1366 vdd.n1117 185
R1370 vdd.n2531 vdd.n1117 185
R1371 vdd.n1365 vdd.n1364 185
R1372 vdd.n1364 vdd.n1116 185
R1373 vdd.n1363 vdd.n1124 185
R1374 vdd.n2525 vdd.n1124 185
R1375 vdd.n1362 vdd.n1361 185
R1376 vdd.n1361 vdd.n1123 185
R1377 vdd.n1360 vdd.n1129 185
R1378 vdd.n2519 vdd.n1129 185
R1379 vdd.n1359 vdd.n1358 185
R1380 vdd.n1358 vdd.n1137 185
R1381 vdd.n1357 vdd.n1135 185
R1382 vdd.n2513 vdd.n1135 185
R1383 vdd.n1356 vdd.n1355 185
R1384 vdd.n1355 vdd.n1134 185
R1385 vdd.n3629 vdd.n3628 185
R1386 vdd.n3628 vdd.n3627 185
R1387 vdd.n3630 vdd.n387 185
R1388 vdd.n387 vdd.n386 185
R1389 vdd.n3632 vdd.n3631 185
R1390 vdd.n3633 vdd.n3632 185
R1391 vdd.n382 vdd.n381 185
R1392 vdd.n3634 vdd.n382 185
R1393 vdd.n3637 vdd.n3636 185
R1394 vdd.n3636 vdd.n3635 185
R1395 vdd.n3638 vdd.n376 185
R1396 vdd.n376 vdd.n375 185
R1397 vdd.n3640 vdd.n3639 185
R1398 vdd.n3641 vdd.n3640 185
R1399 vdd.n371 vdd.n370 185
R1400 vdd.n3642 vdd.n371 185
R1401 vdd.n3645 vdd.n3644 185
R1402 vdd.n3644 vdd.n3643 185
R1403 vdd.n3646 vdd.n365 185
R1404 vdd.n3603 vdd.n365 185
R1405 vdd.n3648 vdd.n3647 185
R1406 vdd.n3649 vdd.n3648 185
R1407 vdd.n360 vdd.n359 185
R1408 vdd.n3650 vdd.n360 185
R1409 vdd.n3653 vdd.n3652 185
R1410 vdd.n3652 vdd.n3651 185
R1411 vdd.n3654 vdd.n354 185
R1412 vdd.n361 vdd.n354 185
R1413 vdd.n3656 vdd.n3655 185
R1414 vdd.n3657 vdd.n3656 185
R1415 vdd.n350 vdd.n349 185
R1416 vdd.n3658 vdd.n350 185
R1417 vdd.n3661 vdd.n3660 185
R1418 vdd.n3660 vdd.n3659 185
R1419 vdd.n3662 vdd.n345 185
R1420 vdd.n345 vdd.n344 185
R1421 vdd.n3664 vdd.n3663 185
R1422 vdd.n3665 vdd.n3664 185
R1423 vdd.n339 vdd.n337 185
R1424 vdd.n3666 vdd.n339 185
R1425 vdd.n3669 vdd.n3668 185
R1426 vdd.n3668 vdd.n3667 185
R1427 vdd.n338 vdd.n336 185
R1428 vdd.n340 vdd.n338 185
R1429 vdd.n3579 vdd.n3578 185
R1430 vdd.n3580 vdd.n3579 185
R1431 vdd.n635 vdd.n634 185
R1432 vdd.n634 vdd.n633 185
R1433 vdd.n3574 vdd.n3573 185
R1434 vdd.n3573 vdd.n3572 185
R1435 vdd.n638 vdd.n637 185
R1436 vdd.n644 vdd.n638 185
R1437 vdd.n3560 vdd.n3559 185
R1438 vdd.n3561 vdd.n3560 185
R1439 vdd.n646 vdd.n645 185
R1440 vdd.n3552 vdd.n645 185
R1441 vdd.n3555 vdd.n3554 185
R1442 vdd.n3554 vdd.n3553 185
R1443 vdd.n649 vdd.n648 185
R1444 vdd.n656 vdd.n649 185
R1445 vdd.n3543 vdd.n3542 185
R1446 vdd.n3544 vdd.n3543 185
R1447 vdd.n658 vdd.n657 185
R1448 vdd.n657 vdd.n655 185
R1449 vdd.n3538 vdd.n3537 185
R1450 vdd.n3537 vdd.n3536 185
R1451 vdd.n661 vdd.n660 185
R1452 vdd.n662 vdd.n661 185
R1453 vdd.n3527 vdd.n3526 185
R1454 vdd.n3528 vdd.n3527 185
R1455 vdd.n669 vdd.n668 185
R1456 vdd.n3519 vdd.n668 185
R1457 vdd.n3522 vdd.n3521 185
R1458 vdd.n3521 vdd.n3520 185
R1459 vdd.n672 vdd.n671 185
R1460 vdd.n679 vdd.n672 185
R1461 vdd.n3510 vdd.n3509 185
R1462 vdd.n3511 vdd.n3510 185
R1463 vdd.n681 vdd.n680 185
R1464 vdd.n680 vdd.n678 185
R1465 vdd.n3505 vdd.n3504 185
R1466 vdd.n3504 vdd.n3503 185
R1467 vdd.n684 vdd.n683 185
R1468 vdd.n723 vdd.n684 185
R1469 vdd.n3493 vdd.n3492 185
R1470 vdd.n3491 vdd.n725 185
R1471 vdd.n3490 vdd.n724 185
R1472 vdd.n3495 vdd.n724 185
R1473 vdd.n729 vdd.n728 185
R1474 vdd.n733 vdd.n732 185
R1475 vdd.n3486 vdd.n734 185
R1476 vdd.n3485 vdd.n3484 185
R1477 vdd.n3483 vdd.n3482 185
R1478 vdd.n3481 vdd.n3480 185
R1479 vdd.n3479 vdd.n3478 185
R1480 vdd.n3477 vdd.n3476 185
R1481 vdd.n3475 vdd.n3474 185
R1482 vdd.n3473 vdd.n3472 185
R1483 vdd.n3471 vdd.n3470 185
R1484 vdd.n3469 vdd.n3468 185
R1485 vdd.n3467 vdd.n3466 185
R1486 vdd.n3465 vdd.n3464 185
R1487 vdd.n3463 vdd.n3462 185
R1488 vdd.n3461 vdd.n3460 185
R1489 vdd.n3459 vdd.n3458 185
R1490 vdd.n3450 vdd.n747 185
R1491 vdd.n3452 vdd.n3451 185
R1492 vdd.n3449 vdd.n3448 185
R1493 vdd.n3447 vdd.n3446 185
R1494 vdd.n3445 vdd.n3444 185
R1495 vdd.n3443 vdd.n3442 185
R1496 vdd.n3441 vdd.n3440 185
R1497 vdd.n3439 vdd.n3438 185
R1498 vdd.n3437 vdd.n3436 185
R1499 vdd.n3435 vdd.n3434 185
R1500 vdd.n3433 vdd.n3432 185
R1501 vdd.n3431 vdd.n3430 185
R1502 vdd.n3429 vdd.n3428 185
R1503 vdd.n3427 vdd.n3426 185
R1504 vdd.n3425 vdd.n3424 185
R1505 vdd.n3423 vdd.n3422 185
R1506 vdd.n3421 vdd.n3420 185
R1507 vdd.n3419 vdd.n3418 185
R1508 vdd.n3417 vdd.n3416 185
R1509 vdd.n3415 vdd.n3414 185
R1510 vdd.n3413 vdd.n3412 185
R1511 vdd.n3411 vdd.n3410 185
R1512 vdd.n3404 vdd.n767 185
R1513 vdd.n3406 vdd.n3405 185
R1514 vdd.n3403 vdd.n3402 185
R1515 vdd.n3401 vdd.n3400 185
R1516 vdd.n3399 vdd.n3398 185
R1517 vdd.n3397 vdd.n3396 185
R1518 vdd.n3395 vdd.n3394 185
R1519 vdd.n3393 vdd.n3392 185
R1520 vdd.n3391 vdd.n3390 185
R1521 vdd.n3389 vdd.n3388 185
R1522 vdd.n3387 vdd.n3386 185
R1523 vdd.n3385 vdd.n3384 185
R1524 vdd.n3383 vdd.n3382 185
R1525 vdd.n3381 vdd.n3380 185
R1526 vdd.n3379 vdd.n3378 185
R1527 vdd.n3377 vdd.n3376 185
R1528 vdd.n3375 vdd.n3374 185
R1529 vdd.n3373 vdd.n3372 185
R1530 vdd.n3371 vdd.n3370 185
R1531 vdd.n3369 vdd.n3368 185
R1532 vdd.n3367 vdd.n691 185
R1533 vdd.n3497 vdd.n3496 185
R1534 vdd.n3496 vdd.n3495 185
R1535 vdd.n3624 vdd.n3623 185
R1536 vdd.n618 vdd.n425 185
R1537 vdd.n617 vdd.n616 185
R1538 vdd.n615 vdd.n614 185
R1539 vdd.n613 vdd.n430 185
R1540 vdd.n609 vdd.n608 185
R1541 vdd.n607 vdd.n606 185
R1542 vdd.n605 vdd.n604 185
R1543 vdd.n603 vdd.n432 185
R1544 vdd.n599 vdd.n598 185
R1545 vdd.n597 vdd.n596 185
R1546 vdd.n595 vdd.n594 185
R1547 vdd.n593 vdd.n434 185
R1548 vdd.n589 vdd.n588 185
R1549 vdd.n587 vdd.n586 185
R1550 vdd.n585 vdd.n584 185
R1551 vdd.n583 vdd.n436 185
R1552 vdd.n579 vdd.n578 185
R1553 vdd.n577 vdd.n576 185
R1554 vdd.n575 vdd.n574 185
R1555 vdd.n573 vdd.n438 185
R1556 vdd.n569 vdd.n568 185
R1557 vdd.n567 vdd.n566 185
R1558 vdd.n565 vdd.n564 185
R1559 vdd.n563 vdd.n442 185
R1560 vdd.n559 vdd.n558 185
R1561 vdd.n557 vdd.n556 185
R1562 vdd.n555 vdd.n554 185
R1563 vdd.n553 vdd.n444 185
R1564 vdd.n549 vdd.n548 185
R1565 vdd.n547 vdd.n546 185
R1566 vdd.n545 vdd.n544 185
R1567 vdd.n543 vdd.n446 185
R1568 vdd.n539 vdd.n538 185
R1569 vdd.n537 vdd.n536 185
R1570 vdd.n535 vdd.n534 185
R1571 vdd.n533 vdd.n448 185
R1572 vdd.n529 vdd.n528 185
R1573 vdd.n527 vdd.n526 185
R1574 vdd.n525 vdd.n524 185
R1575 vdd.n523 vdd.n450 185
R1576 vdd.n519 vdd.n518 185
R1577 vdd.n517 vdd.n516 185
R1578 vdd.n515 vdd.n514 185
R1579 vdd.n513 vdd.n454 185
R1580 vdd.n509 vdd.n508 185
R1581 vdd.n507 vdd.n506 185
R1582 vdd.n505 vdd.n504 185
R1583 vdd.n503 vdd.n456 185
R1584 vdd.n499 vdd.n498 185
R1585 vdd.n497 vdd.n496 185
R1586 vdd.n495 vdd.n494 185
R1587 vdd.n493 vdd.n458 185
R1588 vdd.n489 vdd.n488 185
R1589 vdd.n487 vdd.n486 185
R1590 vdd.n485 vdd.n484 185
R1591 vdd.n483 vdd.n460 185
R1592 vdd.n479 vdd.n478 185
R1593 vdd.n477 vdd.n476 185
R1594 vdd.n475 vdd.n474 185
R1595 vdd.n473 vdd.n462 185
R1596 vdd.n469 vdd.n468 185
R1597 vdd.n467 vdd.n466 185
R1598 vdd.n465 vdd.n392 185
R1599 vdd.n3620 vdd.n393 185
R1600 vdd.n3627 vdd.n393 185
R1601 vdd.n3619 vdd.n3618 185
R1602 vdd.n3618 vdd.n386 185
R1603 vdd.n3617 vdd.n385 185
R1604 vdd.n3633 vdd.n385 185
R1605 vdd.n621 vdd.n384 185
R1606 vdd.n3634 vdd.n384 185
R1607 vdd.n3613 vdd.n383 185
R1608 vdd.n3635 vdd.n383 185
R1609 vdd.n3612 vdd.n3611 185
R1610 vdd.n3611 vdd.n375 185
R1611 vdd.n3610 vdd.n374 185
R1612 vdd.n3641 vdd.n374 185
R1613 vdd.n623 vdd.n373 185
R1614 vdd.n3642 vdd.n373 185
R1615 vdd.n3606 vdd.n372 185
R1616 vdd.n3643 vdd.n372 185
R1617 vdd.n3605 vdd.n3604 185
R1618 vdd.n3604 vdd.n3603 185
R1619 vdd.n3602 vdd.n364 185
R1620 vdd.n3649 vdd.n364 185
R1621 vdd.n625 vdd.n363 185
R1622 vdd.n3650 vdd.n363 185
R1623 vdd.n3598 vdd.n362 185
R1624 vdd.n3651 vdd.n362 185
R1625 vdd.n3597 vdd.n3596 185
R1626 vdd.n3596 vdd.n361 185
R1627 vdd.n3595 vdd.n353 185
R1628 vdd.n3657 vdd.n353 185
R1629 vdd.n627 vdd.n352 185
R1630 vdd.n3658 vdd.n352 185
R1631 vdd.n3591 vdd.n351 185
R1632 vdd.n3659 vdd.n351 185
R1633 vdd.n3590 vdd.n3589 185
R1634 vdd.n3589 vdd.n344 185
R1635 vdd.n3588 vdd.n343 185
R1636 vdd.n3665 vdd.n343 185
R1637 vdd.n629 vdd.n342 185
R1638 vdd.n3666 vdd.n342 185
R1639 vdd.n3584 vdd.n341 185
R1640 vdd.n3667 vdd.n341 185
R1641 vdd.n3583 vdd.n3582 185
R1642 vdd.n3582 vdd.n340 185
R1643 vdd.n3581 vdd.n631 185
R1644 vdd.n3581 vdd.n3580 185
R1645 vdd.n3569 vdd.n632 185
R1646 vdd.n633 vdd.n632 185
R1647 vdd.n3571 vdd.n3570 185
R1648 vdd.n3572 vdd.n3571 185
R1649 vdd.n640 vdd.n639 185
R1650 vdd.n644 vdd.n639 185
R1651 vdd.n3563 vdd.n3562 185
R1652 vdd.n3562 vdd.n3561 185
R1653 vdd.n643 vdd.n642 185
R1654 vdd.n3552 vdd.n643 185
R1655 vdd.n3551 vdd.n3550 185
R1656 vdd.n3553 vdd.n3551 185
R1657 vdd.n651 vdd.n650 185
R1658 vdd.n656 vdd.n650 185
R1659 vdd.n3546 vdd.n3545 185
R1660 vdd.n3545 vdd.n3544 185
R1661 vdd.n654 vdd.n653 185
R1662 vdd.n655 vdd.n654 185
R1663 vdd.n3535 vdd.n3534 185
R1664 vdd.n3536 vdd.n3535 185
R1665 vdd.n664 vdd.n663 185
R1666 vdd.n663 vdd.n662 185
R1667 vdd.n3530 vdd.n3529 185
R1668 vdd.n3529 vdd.n3528 185
R1669 vdd.n667 vdd.n666 185
R1670 vdd.n3519 vdd.n667 185
R1671 vdd.n3518 vdd.n3517 185
R1672 vdd.n3520 vdd.n3518 185
R1673 vdd.n674 vdd.n673 185
R1674 vdd.n679 vdd.n673 185
R1675 vdd.n3513 vdd.n3512 185
R1676 vdd.n3512 vdd.n3511 185
R1677 vdd.n677 vdd.n676 185
R1678 vdd.n678 vdd.n677 185
R1679 vdd.n3502 vdd.n3501 185
R1680 vdd.n3503 vdd.n3502 185
R1681 vdd.n686 vdd.n685 185
R1682 vdd.n723 vdd.n685 185
R1683 vdd.n3091 vdd.n3090 185
R1684 vdd.n962 vdd.n961 185
R1685 vdd.n3087 vdd.n3086 185
R1686 vdd.n3088 vdd.n3087 185
R1687 vdd.n3085 vdd.n2819 185
R1688 vdd.n3084 vdd.n3083 185
R1689 vdd.n3082 vdd.n3081 185
R1690 vdd.n3080 vdd.n3079 185
R1691 vdd.n3078 vdd.n3077 185
R1692 vdd.n3076 vdd.n3075 185
R1693 vdd.n3074 vdd.n3073 185
R1694 vdd.n3072 vdd.n3071 185
R1695 vdd.n3070 vdd.n3069 185
R1696 vdd.n3068 vdd.n3067 185
R1697 vdd.n3066 vdd.n3065 185
R1698 vdd.n3064 vdd.n3063 185
R1699 vdd.n3062 vdd.n3061 185
R1700 vdd.n3060 vdd.n3059 185
R1701 vdd.n3058 vdd.n3057 185
R1702 vdd.n3056 vdd.n3055 185
R1703 vdd.n3054 vdd.n3053 185
R1704 vdd.n3052 vdd.n3051 185
R1705 vdd.n3050 vdd.n3049 185
R1706 vdd.n3048 vdd.n3047 185
R1707 vdd.n3046 vdd.n3045 185
R1708 vdd.n3044 vdd.n3043 185
R1709 vdd.n3042 vdd.n3041 185
R1710 vdd.n3040 vdd.n3039 185
R1711 vdd.n3038 vdd.n3037 185
R1712 vdd.n3036 vdd.n3035 185
R1713 vdd.n3034 vdd.n3033 185
R1714 vdd.n3032 vdd.n3031 185
R1715 vdd.n3030 vdd.n3029 185
R1716 vdd.n3027 vdd.n3026 185
R1717 vdd.n3025 vdd.n3024 185
R1718 vdd.n3023 vdd.n3022 185
R1719 vdd.n3267 vdd.n3266 185
R1720 vdd.n3269 vdd.n834 185
R1721 vdd.n3271 vdd.n3270 185
R1722 vdd.n3273 vdd.n831 185
R1723 vdd.n3275 vdd.n3274 185
R1724 vdd.n3277 vdd.n829 185
R1725 vdd.n3279 vdd.n3278 185
R1726 vdd.n3280 vdd.n828 185
R1727 vdd.n3282 vdd.n3281 185
R1728 vdd.n3284 vdd.n826 185
R1729 vdd.n3286 vdd.n3285 185
R1730 vdd.n3287 vdd.n825 185
R1731 vdd.n3289 vdd.n3288 185
R1732 vdd.n3291 vdd.n823 185
R1733 vdd.n3293 vdd.n3292 185
R1734 vdd.n3294 vdd.n822 185
R1735 vdd.n3296 vdd.n3295 185
R1736 vdd.n3298 vdd.n731 185
R1737 vdd.n3300 vdd.n3299 185
R1738 vdd.n3302 vdd.n820 185
R1739 vdd.n3304 vdd.n3303 185
R1740 vdd.n3305 vdd.n819 185
R1741 vdd.n3307 vdd.n3306 185
R1742 vdd.n3309 vdd.n817 185
R1743 vdd.n3311 vdd.n3310 185
R1744 vdd.n3312 vdd.n816 185
R1745 vdd.n3314 vdd.n3313 185
R1746 vdd.n3316 vdd.n814 185
R1747 vdd.n3318 vdd.n3317 185
R1748 vdd.n3319 vdd.n813 185
R1749 vdd.n3321 vdd.n3320 185
R1750 vdd.n3323 vdd.n812 185
R1751 vdd.n3324 vdd.n811 185
R1752 vdd.n3327 vdd.n3326 185
R1753 vdd.n3328 vdd.n809 185
R1754 vdd.n809 vdd.n692 185
R1755 vdd.n3265 vdd.n806 185
R1756 vdd.n3331 vdd.n806 185
R1757 vdd.n3264 vdd.n3263 185
R1758 vdd.n3263 vdd.n805 185
R1759 vdd.n3262 vdd.n836 185
R1760 vdd.n3262 vdd.n3261 185
R1761 vdd.n2905 vdd.n837 185
R1762 vdd.n846 vdd.n837 185
R1763 vdd.n2906 vdd.n844 185
R1764 vdd.n3255 vdd.n844 185
R1765 vdd.n2908 vdd.n2907 185
R1766 vdd.n2907 vdd.n843 185
R1767 vdd.n2909 vdd.n852 185
R1768 vdd.n3204 vdd.n852 185
R1769 vdd.n2911 vdd.n2910 185
R1770 vdd.n2910 vdd.n851 185
R1771 vdd.n2912 vdd.n857 185
R1772 vdd.n3198 vdd.n857 185
R1773 vdd.n2914 vdd.n2913 185
R1774 vdd.n2913 vdd.n864 185
R1775 vdd.n2915 vdd.n862 185
R1776 vdd.n3192 vdd.n862 185
R1777 vdd.n2917 vdd.n2916 185
R1778 vdd.n2916 vdd.n870 185
R1779 vdd.n2918 vdd.n868 185
R1780 vdd.n3186 vdd.n868 185
R1781 vdd.n2920 vdd.n2919 185
R1782 vdd.n2919 vdd.n877 185
R1783 vdd.n2921 vdd.n875 185
R1784 vdd.n3180 vdd.n875 185
R1785 vdd.n2923 vdd.n2922 185
R1786 vdd.n2922 vdd.n874 185
R1787 vdd.n2924 vdd.n882 185
R1788 vdd.n3174 vdd.n882 185
R1789 vdd.n2926 vdd.n2925 185
R1790 vdd.n2925 vdd.n881 185
R1791 vdd.n2927 vdd.n888 185
R1792 vdd.n3168 vdd.n888 185
R1793 vdd.n2929 vdd.n2928 185
R1794 vdd.n2928 vdd.n887 185
R1795 vdd.n2930 vdd.n893 185
R1796 vdd.n3162 vdd.n893 185
R1797 vdd.n2932 vdd.n2931 185
R1798 vdd.n2931 vdd.n901 185
R1799 vdd.n2933 vdd.n899 185
R1800 vdd.n3156 vdd.n899 185
R1801 vdd.n2935 vdd.n2934 185
R1802 vdd.n2934 vdd.n908 185
R1803 vdd.n2936 vdd.n906 185
R1804 vdd.n3150 vdd.n906 185
R1805 vdd.n2938 vdd.n2937 185
R1806 vdd.n2937 vdd.n905 185
R1807 vdd.n2939 vdd.n913 185
R1808 vdd.n3143 vdd.n913 185
R1809 vdd.n2941 vdd.n2940 185
R1810 vdd.n2940 vdd.n912 185
R1811 vdd.n2942 vdd.n918 185
R1812 vdd.n3137 vdd.n918 185
R1813 vdd.n2944 vdd.n2943 185
R1814 vdd.n2943 vdd.n925 185
R1815 vdd.n2945 vdd.n923 185
R1816 vdd.n3131 vdd.n923 185
R1817 vdd.n2947 vdd.n2946 185
R1818 vdd.n2946 vdd.n931 185
R1819 vdd.n2948 vdd.n929 185
R1820 vdd.n3125 vdd.n929 185
R1821 vdd.n3000 vdd.n2999 185
R1822 vdd.n2999 vdd.n2998 185
R1823 vdd.n3001 vdd.n935 185
R1824 vdd.n3119 vdd.n935 185
R1825 vdd.n3003 vdd.n3002 185
R1826 vdd.n3004 vdd.n3003 185
R1827 vdd.n2904 vdd.n941 185
R1828 vdd.n3113 vdd.n941 185
R1829 vdd.n2903 vdd.n2902 185
R1830 vdd.n2902 vdd.n940 185
R1831 vdd.n2901 vdd.n947 185
R1832 vdd.n3107 vdd.n947 185
R1833 vdd.n2900 vdd.n2899 185
R1834 vdd.n2899 vdd.n946 185
R1835 vdd.n2822 vdd.n952 185
R1836 vdd.n3101 vdd.n952 185
R1837 vdd.n3018 vdd.n3017 185
R1838 vdd.n3017 vdd.n3016 185
R1839 vdd.n3019 vdd.n958 185
R1840 vdd.n3095 vdd.n958 185
R1841 vdd.n3021 vdd.n3020 185
R1842 vdd.n3021 vdd.n957 185
R1843 vdd.n3092 vdd.n960 185
R1844 vdd.n960 vdd.n957 185
R1845 vdd.n3094 vdd.n3093 185
R1846 vdd.n3095 vdd.n3094 185
R1847 vdd.n951 vdd.n950 185
R1848 vdd.n3016 vdd.n951 185
R1849 vdd.n3103 vdd.n3102 185
R1850 vdd.n3102 vdd.n3101 185
R1851 vdd.n3104 vdd.n949 185
R1852 vdd.n949 vdd.n946 185
R1853 vdd.n3106 vdd.n3105 185
R1854 vdd.n3107 vdd.n3106 185
R1855 vdd.n939 vdd.n938 185
R1856 vdd.n940 vdd.n939 185
R1857 vdd.n3115 vdd.n3114 185
R1858 vdd.n3114 vdd.n3113 185
R1859 vdd.n3116 vdd.n937 185
R1860 vdd.n3004 vdd.n937 185
R1861 vdd.n3118 vdd.n3117 185
R1862 vdd.n3119 vdd.n3118 185
R1863 vdd.n928 vdd.n927 185
R1864 vdd.n2998 vdd.n928 185
R1865 vdd.n3127 vdd.n3126 185
R1866 vdd.n3126 vdd.n3125 185
R1867 vdd.n3128 vdd.n926 185
R1868 vdd.n931 vdd.n926 185
R1869 vdd.n3130 vdd.n3129 185
R1870 vdd.n3131 vdd.n3130 185
R1871 vdd.n917 vdd.n916 185
R1872 vdd.n925 vdd.n917 185
R1873 vdd.n3139 vdd.n3138 185
R1874 vdd.n3138 vdd.n3137 185
R1875 vdd.n3140 vdd.n915 185
R1876 vdd.n915 vdd.n912 185
R1877 vdd.n3142 vdd.n3141 185
R1878 vdd.n3143 vdd.n3142 185
R1879 vdd.n904 vdd.n903 185
R1880 vdd.n905 vdd.n904 185
R1881 vdd.n3152 vdd.n3151 185
R1882 vdd.n3151 vdd.n3150 185
R1883 vdd.n3153 vdd.n902 185
R1884 vdd.n908 vdd.n902 185
R1885 vdd.n3155 vdd.n3154 185
R1886 vdd.n3156 vdd.n3155 185
R1887 vdd.n892 vdd.n891 185
R1888 vdd.n901 vdd.n892 185
R1889 vdd.n3164 vdd.n3163 185
R1890 vdd.n3163 vdd.n3162 185
R1891 vdd.n3165 vdd.n890 185
R1892 vdd.n890 vdd.n887 185
R1893 vdd.n3167 vdd.n3166 185
R1894 vdd.n3168 vdd.n3167 185
R1895 vdd.n880 vdd.n879 185
R1896 vdd.n881 vdd.n880 185
R1897 vdd.n3176 vdd.n3175 185
R1898 vdd.n3175 vdd.n3174 185
R1899 vdd.n3177 vdd.n878 185
R1900 vdd.n878 vdd.n874 185
R1901 vdd.n3179 vdd.n3178 185
R1902 vdd.n3180 vdd.n3179 185
R1903 vdd.n867 vdd.n866 185
R1904 vdd.n877 vdd.n867 185
R1905 vdd.n3188 vdd.n3187 185
R1906 vdd.n3187 vdd.n3186 185
R1907 vdd.n3189 vdd.n865 185
R1908 vdd.n870 vdd.n865 185
R1909 vdd.n3191 vdd.n3190 185
R1910 vdd.n3192 vdd.n3191 185
R1911 vdd.n856 vdd.n855 185
R1912 vdd.n864 vdd.n856 185
R1913 vdd.n3200 vdd.n3199 185
R1914 vdd.n3199 vdd.n3198 185
R1915 vdd.n3201 vdd.n854 185
R1916 vdd.n854 vdd.n851 185
R1917 vdd.n3203 vdd.n3202 185
R1918 vdd.n3204 vdd.n3203 185
R1919 vdd.n842 vdd.n841 185
R1920 vdd.n843 vdd.n842 185
R1921 vdd.n3257 vdd.n3256 185
R1922 vdd.n3256 vdd.n3255 185
R1923 vdd.n3258 vdd.n840 185
R1924 vdd.n846 vdd.n840 185
R1925 vdd.n3260 vdd.n3259 185
R1926 vdd.n3261 vdd.n3260 185
R1927 vdd.n810 vdd.n808 185
R1928 vdd.n808 vdd.n805 185
R1929 vdd.n3330 vdd.n3329 185
R1930 vdd.n3331 vdd.n3330 185
R1931 vdd.n2711 vdd.n2710 185
R1932 vdd.n2712 vdd.n2711 185
R1933 vdd.n1009 vdd.n1007 185
R1934 vdd.n1007 vdd.n1005 185
R1935 vdd.n2626 vdd.n1016 185
R1936 vdd.n2637 vdd.n1016 185
R1937 vdd.n2627 vdd.n1025 185
R1938 vdd.n1399 vdd.n1025 185
R1939 vdd.n2629 vdd.n2628 185
R1940 vdd.n2630 vdd.n2629 185
R1941 vdd.n2625 vdd.n1024 185
R1942 vdd.n1024 vdd.n1021 185
R1943 vdd.n2624 vdd.n2623 185
R1944 vdd.n2623 vdd.n2622 185
R1945 vdd.n1027 vdd.n1026 185
R1946 vdd.n1028 vdd.n1027 185
R1947 vdd.n2615 vdd.n2614 185
R1948 vdd.n2616 vdd.n2615 185
R1949 vdd.n2613 vdd.n1036 185
R1950 vdd.n1425 vdd.n1036 185
R1951 vdd.n2612 vdd.n2611 185
R1952 vdd.n2611 vdd.n2610 185
R1953 vdd.n1038 vdd.n1037 185
R1954 vdd.n1046 vdd.n1038 185
R1955 vdd.n2603 vdd.n2602 185
R1956 vdd.n2604 vdd.n2603 185
R1957 vdd.n2601 vdd.n1047 185
R1958 vdd.n1052 vdd.n1047 185
R1959 vdd.n2600 vdd.n2599 185
R1960 vdd.n2599 vdd.n2598 185
R1961 vdd.n1049 vdd.n1048 185
R1962 vdd.n1437 vdd.n1049 185
R1963 vdd.n2591 vdd.n2590 185
R1964 vdd.n2592 vdd.n2591 185
R1965 vdd.n2589 vdd.n1059 185
R1966 vdd.n1059 vdd.n1056 185
R1967 vdd.n2588 vdd.n2587 185
R1968 vdd.n2587 vdd.n2586 185
R1969 vdd.n1061 vdd.n1060 185
R1970 vdd.n1062 vdd.n1061 185
R1971 vdd.n2579 vdd.n2578 185
R1972 vdd.n2580 vdd.n2579 185
R1973 vdd.n2576 vdd.n1070 185
R1974 vdd.n1076 vdd.n1070 185
R1975 vdd.n2575 vdd.n2574 185
R1976 vdd.n2574 vdd.n2573 185
R1977 vdd.n1073 vdd.n1072 185
R1978 vdd.n1083 vdd.n1073 185
R1979 vdd.n2566 vdd.n2565 185
R1980 vdd.n2567 vdd.n2566 185
R1981 vdd.n2564 vdd.n1084 185
R1982 vdd.n1084 vdd.n1080 185
R1983 vdd.n2563 vdd.n2562 185
R1984 vdd.n2562 vdd.n2561 185
R1985 vdd.n1086 vdd.n1085 185
R1986 vdd.n1087 vdd.n1086 185
R1987 vdd.n2554 vdd.n2553 185
R1988 vdd.n2555 vdd.n2554 185
R1989 vdd.n2552 vdd.n1096 185
R1990 vdd.n1096 vdd.n1093 185
R1991 vdd.n2551 vdd.n2550 185
R1992 vdd.n2550 vdd.n2549 185
R1993 vdd.n1098 vdd.n1097 185
R1994 vdd.n1106 vdd.n1098 185
R1995 vdd.n2542 vdd.n2541 185
R1996 vdd.n2543 vdd.n2542 185
R1997 vdd.n2540 vdd.n1107 185
R1998 vdd.n1112 vdd.n1107 185
R1999 vdd.n2539 vdd.n2538 185
R2000 vdd.n2538 vdd.n2537 185
R2001 vdd.n1109 vdd.n1108 185
R2002 vdd.n1119 vdd.n1109 185
R2003 vdd.n2530 vdd.n2529 185
R2004 vdd.n2531 vdd.n2530 185
R2005 vdd.n2528 vdd.n1120 185
R2006 vdd.n1120 vdd.n1116 185
R2007 vdd.n2527 vdd.n2526 185
R2008 vdd.n2526 vdd.n2525 185
R2009 vdd.n1122 vdd.n1121 185
R2010 vdd.n1123 vdd.n1122 185
R2011 vdd.n2518 vdd.n2517 185
R2012 vdd.n2519 vdd.n2518 185
R2013 vdd.n2516 vdd.n1131 185
R2014 vdd.n1137 vdd.n1131 185
R2015 vdd.n2515 vdd.n2514 185
R2016 vdd.n2514 vdd.n2513 185
R2017 vdd.n1133 vdd.n1132 185
R2018 vdd.n1134 vdd.n1133 185
R2019 vdd.n2642 vdd.n980 185
R2020 vdd.n2784 vdd.n980 185
R2021 vdd.n2644 vdd.n2643 185
R2022 vdd.n2646 vdd.n2645 185
R2023 vdd.n2648 vdd.n2647 185
R2024 vdd.n2650 vdd.n2649 185
R2025 vdd.n2652 vdd.n2651 185
R2026 vdd.n2654 vdd.n2653 185
R2027 vdd.n2656 vdd.n2655 185
R2028 vdd.n2658 vdd.n2657 185
R2029 vdd.n2660 vdd.n2659 185
R2030 vdd.n2662 vdd.n2661 185
R2031 vdd.n2664 vdd.n2663 185
R2032 vdd.n2666 vdd.n2665 185
R2033 vdd.n2668 vdd.n2667 185
R2034 vdd.n2670 vdd.n2669 185
R2035 vdd.n2672 vdd.n2671 185
R2036 vdd.n2674 vdd.n2673 185
R2037 vdd.n2676 vdd.n2675 185
R2038 vdd.n2678 vdd.n2677 185
R2039 vdd.n2680 vdd.n2679 185
R2040 vdd.n2682 vdd.n2681 185
R2041 vdd.n2684 vdd.n2683 185
R2042 vdd.n2686 vdd.n2685 185
R2043 vdd.n2688 vdd.n2687 185
R2044 vdd.n2690 vdd.n2689 185
R2045 vdd.n2692 vdd.n2691 185
R2046 vdd.n2694 vdd.n2693 185
R2047 vdd.n2696 vdd.n2695 185
R2048 vdd.n2698 vdd.n2697 185
R2049 vdd.n2700 vdd.n2699 185
R2050 vdd.n2702 vdd.n2701 185
R2051 vdd.n2704 vdd.n2703 185
R2052 vdd.n2706 vdd.n2705 185
R2053 vdd.n2708 vdd.n2707 185
R2054 vdd.n2709 vdd.n1008 185
R2055 vdd.n2641 vdd.n1006 185
R2056 vdd.n2712 vdd.n1006 185
R2057 vdd.n2640 vdd.n2639 185
R2058 vdd.n2639 vdd.n1005 185
R2059 vdd.n2638 vdd.n1013 185
R2060 vdd.n2638 vdd.n2637 185
R2061 vdd.n1415 vdd.n1014 185
R2062 vdd.n1399 vdd.n1014 185
R2063 vdd.n1416 vdd.n1023 185
R2064 vdd.n2630 vdd.n1023 185
R2065 vdd.n1418 vdd.n1417 185
R2066 vdd.n1417 vdd.n1021 185
R2067 vdd.n1419 vdd.n1030 185
R2068 vdd.n2622 vdd.n1030 185
R2069 vdd.n1421 vdd.n1420 185
R2070 vdd.n1420 vdd.n1028 185
R2071 vdd.n1422 vdd.n1035 185
R2072 vdd.n2616 vdd.n1035 185
R2073 vdd.n1424 vdd.n1423 185
R2074 vdd.n1425 vdd.n1424 185
R2075 vdd.n1414 vdd.n1040 185
R2076 vdd.n2610 vdd.n1040 185
R2077 vdd.n1413 vdd.n1412 185
R2078 vdd.n1412 vdd.n1046 185
R2079 vdd.n1411 vdd.n1045 185
R2080 vdd.n2604 vdd.n1045 185
R2081 vdd.n1410 vdd.n1409 185
R2082 vdd.n1409 vdd.n1052 185
R2083 vdd.n1318 vdd.n1051 185
R2084 vdd.n2598 vdd.n1051 185
R2085 vdd.n1439 vdd.n1438 185
R2086 vdd.n1438 vdd.n1437 185
R2087 vdd.n1440 vdd.n1058 185
R2088 vdd.n2592 vdd.n1058 185
R2089 vdd.n1442 vdd.n1441 185
R2090 vdd.n1441 vdd.n1056 185
R2091 vdd.n1443 vdd.n1064 185
R2092 vdd.n2586 vdd.n1064 185
R2093 vdd.n1445 vdd.n1444 185
R2094 vdd.n1444 vdd.n1062 185
R2095 vdd.n1446 vdd.n1069 185
R2096 vdd.n2580 vdd.n1069 185
R2097 vdd.n1448 vdd.n1447 185
R2098 vdd.n1447 vdd.n1076 185
R2099 vdd.n1449 vdd.n1075 185
R2100 vdd.n2573 vdd.n1075 185
R2101 vdd.n1451 vdd.n1450 185
R2102 vdd.n1450 vdd.n1083 185
R2103 vdd.n1452 vdd.n1082 185
R2104 vdd.n2567 vdd.n1082 185
R2105 vdd.n1454 vdd.n1453 185
R2106 vdd.n1453 vdd.n1080 185
R2107 vdd.n1455 vdd.n1089 185
R2108 vdd.n2561 vdd.n1089 185
R2109 vdd.n1457 vdd.n1456 185
R2110 vdd.n1456 vdd.n1087 185
R2111 vdd.n1458 vdd.n1095 185
R2112 vdd.n2555 vdd.n1095 185
R2113 vdd.n1460 vdd.n1459 185
R2114 vdd.n1459 vdd.n1093 185
R2115 vdd.n1461 vdd.n1100 185
R2116 vdd.n2549 vdd.n1100 185
R2117 vdd.n1463 vdd.n1462 185
R2118 vdd.n1462 vdd.n1106 185
R2119 vdd.n1464 vdd.n1105 185
R2120 vdd.n2543 vdd.n1105 185
R2121 vdd.n1466 vdd.n1465 185
R2122 vdd.n1465 vdd.n1112 185
R2123 vdd.n1467 vdd.n1111 185
R2124 vdd.n2537 vdd.n1111 185
R2125 vdd.n1469 vdd.n1468 185
R2126 vdd.n1468 vdd.n1119 185
R2127 vdd.n1470 vdd.n1118 185
R2128 vdd.n2531 vdd.n1118 185
R2129 vdd.n1472 vdd.n1471 185
R2130 vdd.n1471 vdd.n1116 185
R2131 vdd.n1473 vdd.n1125 185
R2132 vdd.n2525 vdd.n1125 185
R2133 vdd.n1475 vdd.n1474 185
R2134 vdd.n1474 vdd.n1123 185
R2135 vdd.n1476 vdd.n1130 185
R2136 vdd.n2519 vdd.n1130 185
R2137 vdd.n1478 vdd.n1477 185
R2138 vdd.n1477 vdd.n1137 185
R2139 vdd.n1479 vdd.n1136 185
R2140 vdd.n2513 vdd.n1136 185
R2141 vdd.n1481 vdd.n1480 185
R2142 vdd.n1480 vdd.n1134 185
R2143 vdd.n1281 vdd.n1280 185
R2144 vdd.n1283 vdd.n1282 185
R2145 vdd.n1285 vdd.n1284 185
R2146 vdd.n1287 vdd.n1286 185
R2147 vdd.n1289 vdd.n1288 185
R2148 vdd.n1291 vdd.n1290 185
R2149 vdd.n1293 vdd.n1292 185
R2150 vdd.n1295 vdd.n1294 185
R2151 vdd.n1297 vdd.n1296 185
R2152 vdd.n1299 vdd.n1298 185
R2153 vdd.n1301 vdd.n1300 185
R2154 vdd.n1303 vdd.n1302 185
R2155 vdd.n1305 vdd.n1304 185
R2156 vdd.n1307 vdd.n1306 185
R2157 vdd.n1309 vdd.n1308 185
R2158 vdd.n1311 vdd.n1310 185
R2159 vdd.n1313 vdd.n1312 185
R2160 vdd.n1515 vdd.n1314 185
R2161 vdd.n1514 vdd.n1513 185
R2162 vdd.n1512 vdd.n1511 185
R2163 vdd.n1510 vdd.n1509 185
R2164 vdd.n1508 vdd.n1507 185
R2165 vdd.n1506 vdd.n1505 185
R2166 vdd.n1504 vdd.n1503 185
R2167 vdd.n1502 vdd.n1501 185
R2168 vdd.n1500 vdd.n1499 185
R2169 vdd.n1498 vdd.n1497 185
R2170 vdd.n1496 vdd.n1495 185
R2171 vdd.n1494 vdd.n1493 185
R2172 vdd.n1492 vdd.n1491 185
R2173 vdd.n1490 vdd.n1489 185
R2174 vdd.n1488 vdd.n1487 185
R2175 vdd.n1486 vdd.n1485 185
R2176 vdd.n1484 vdd.n1483 185
R2177 vdd.n1482 vdd.n1175 185
R2178 vdd.n2506 vdd.n1175 185
R2179 vdd.n327 vdd.n326 171.744
R2180 vdd.n326 vdd.n325 171.744
R2181 vdd.n325 vdd.n294 171.744
R2182 vdd.n318 vdd.n294 171.744
R2183 vdd.n318 vdd.n317 171.744
R2184 vdd.n317 vdd.n299 171.744
R2185 vdd.n310 vdd.n299 171.744
R2186 vdd.n310 vdd.n309 171.744
R2187 vdd.n309 vdd.n303 171.744
R2188 vdd.n268 vdd.n267 171.744
R2189 vdd.n267 vdd.n266 171.744
R2190 vdd.n266 vdd.n235 171.744
R2191 vdd.n259 vdd.n235 171.744
R2192 vdd.n259 vdd.n258 171.744
R2193 vdd.n258 vdd.n240 171.744
R2194 vdd.n251 vdd.n240 171.744
R2195 vdd.n251 vdd.n250 171.744
R2196 vdd.n250 vdd.n244 171.744
R2197 vdd.n225 vdd.n224 171.744
R2198 vdd.n224 vdd.n223 171.744
R2199 vdd.n223 vdd.n192 171.744
R2200 vdd.n216 vdd.n192 171.744
R2201 vdd.n216 vdd.n215 171.744
R2202 vdd.n215 vdd.n197 171.744
R2203 vdd.n208 vdd.n197 171.744
R2204 vdd.n208 vdd.n207 171.744
R2205 vdd.n207 vdd.n201 171.744
R2206 vdd.n166 vdd.n165 171.744
R2207 vdd.n165 vdd.n164 171.744
R2208 vdd.n164 vdd.n133 171.744
R2209 vdd.n157 vdd.n133 171.744
R2210 vdd.n157 vdd.n156 171.744
R2211 vdd.n156 vdd.n138 171.744
R2212 vdd.n149 vdd.n138 171.744
R2213 vdd.n149 vdd.n148 171.744
R2214 vdd.n148 vdd.n142 171.744
R2215 vdd.n124 vdd.n123 171.744
R2216 vdd.n123 vdd.n122 171.744
R2217 vdd.n122 vdd.n91 171.744
R2218 vdd.n115 vdd.n91 171.744
R2219 vdd.n115 vdd.n114 171.744
R2220 vdd.n114 vdd.n96 171.744
R2221 vdd.n107 vdd.n96 171.744
R2222 vdd.n107 vdd.n106 171.744
R2223 vdd.n106 vdd.n100 171.744
R2224 vdd.n65 vdd.n64 171.744
R2225 vdd.n64 vdd.n63 171.744
R2226 vdd.n63 vdd.n32 171.744
R2227 vdd.n56 vdd.n32 171.744
R2228 vdd.n56 vdd.n55 171.744
R2229 vdd.n55 vdd.n37 171.744
R2230 vdd.n48 vdd.n37 171.744
R2231 vdd.n48 vdd.n47 171.744
R2232 vdd.n47 vdd.n41 171.744
R2233 vdd.n2201 vdd.n2200 171.744
R2234 vdd.n2200 vdd.n2199 171.744
R2235 vdd.n2199 vdd.n2168 171.744
R2236 vdd.n2192 vdd.n2168 171.744
R2237 vdd.n2192 vdd.n2191 171.744
R2238 vdd.n2191 vdd.n2173 171.744
R2239 vdd.n2184 vdd.n2173 171.744
R2240 vdd.n2184 vdd.n2183 171.744
R2241 vdd.n2183 vdd.n2177 171.744
R2242 vdd.n2260 vdd.n2259 171.744
R2243 vdd.n2259 vdd.n2258 171.744
R2244 vdd.n2258 vdd.n2227 171.744
R2245 vdd.n2251 vdd.n2227 171.744
R2246 vdd.n2251 vdd.n2250 171.744
R2247 vdd.n2250 vdd.n2232 171.744
R2248 vdd.n2243 vdd.n2232 171.744
R2249 vdd.n2243 vdd.n2242 171.744
R2250 vdd.n2242 vdd.n2236 171.744
R2251 vdd.n2099 vdd.n2098 171.744
R2252 vdd.n2098 vdd.n2097 171.744
R2253 vdd.n2097 vdd.n2066 171.744
R2254 vdd.n2090 vdd.n2066 171.744
R2255 vdd.n2090 vdd.n2089 171.744
R2256 vdd.n2089 vdd.n2071 171.744
R2257 vdd.n2082 vdd.n2071 171.744
R2258 vdd.n2082 vdd.n2081 171.744
R2259 vdd.n2081 vdd.n2075 171.744
R2260 vdd.n2158 vdd.n2157 171.744
R2261 vdd.n2157 vdd.n2156 171.744
R2262 vdd.n2156 vdd.n2125 171.744
R2263 vdd.n2149 vdd.n2125 171.744
R2264 vdd.n2149 vdd.n2148 171.744
R2265 vdd.n2148 vdd.n2130 171.744
R2266 vdd.n2141 vdd.n2130 171.744
R2267 vdd.n2141 vdd.n2140 171.744
R2268 vdd.n2140 vdd.n2134 171.744
R2269 vdd.n1998 vdd.n1997 171.744
R2270 vdd.n1997 vdd.n1996 171.744
R2271 vdd.n1996 vdd.n1965 171.744
R2272 vdd.n1989 vdd.n1965 171.744
R2273 vdd.n1989 vdd.n1988 171.744
R2274 vdd.n1988 vdd.n1970 171.744
R2275 vdd.n1981 vdd.n1970 171.744
R2276 vdd.n1981 vdd.n1980 171.744
R2277 vdd.n1980 vdd.n1974 171.744
R2278 vdd.n2057 vdd.n2056 171.744
R2279 vdd.n2056 vdd.n2055 171.744
R2280 vdd.n2055 vdd.n2024 171.744
R2281 vdd.n2048 vdd.n2024 171.744
R2282 vdd.n2048 vdd.n2047 171.744
R2283 vdd.n2047 vdd.n2029 171.744
R2284 vdd.n2040 vdd.n2029 171.744
R2285 vdd.n2040 vdd.n2039 171.744
R2286 vdd.n2039 vdd.n2033 171.744
R2287 vdd.n468 vdd.n467 146.341
R2288 vdd.n474 vdd.n473 146.341
R2289 vdd.n478 vdd.n477 146.341
R2290 vdd.n484 vdd.n483 146.341
R2291 vdd.n488 vdd.n487 146.341
R2292 vdd.n494 vdd.n493 146.341
R2293 vdd.n498 vdd.n497 146.341
R2294 vdd.n504 vdd.n503 146.341
R2295 vdd.n508 vdd.n507 146.341
R2296 vdd.n514 vdd.n513 146.341
R2297 vdd.n518 vdd.n517 146.341
R2298 vdd.n524 vdd.n523 146.341
R2299 vdd.n528 vdd.n527 146.341
R2300 vdd.n534 vdd.n533 146.341
R2301 vdd.n538 vdd.n537 146.341
R2302 vdd.n544 vdd.n543 146.341
R2303 vdd.n548 vdd.n547 146.341
R2304 vdd.n554 vdd.n553 146.341
R2305 vdd.n558 vdd.n557 146.341
R2306 vdd.n564 vdd.n563 146.341
R2307 vdd.n568 vdd.n567 146.341
R2308 vdd.n574 vdd.n573 146.341
R2309 vdd.n578 vdd.n577 146.341
R2310 vdd.n584 vdd.n583 146.341
R2311 vdd.n588 vdd.n587 146.341
R2312 vdd.n594 vdd.n593 146.341
R2313 vdd.n598 vdd.n597 146.341
R2314 vdd.n604 vdd.n603 146.341
R2315 vdd.n608 vdd.n607 146.341
R2316 vdd.n614 vdd.n613 146.341
R2317 vdd.n616 vdd.n425 146.341
R2318 vdd.n3502 vdd.n685 146.341
R2319 vdd.n3502 vdd.n677 146.341
R2320 vdd.n3512 vdd.n677 146.341
R2321 vdd.n3512 vdd.n673 146.341
R2322 vdd.n3518 vdd.n673 146.341
R2323 vdd.n3518 vdd.n667 146.341
R2324 vdd.n3529 vdd.n667 146.341
R2325 vdd.n3529 vdd.n663 146.341
R2326 vdd.n3535 vdd.n663 146.341
R2327 vdd.n3535 vdd.n654 146.341
R2328 vdd.n3545 vdd.n654 146.341
R2329 vdd.n3545 vdd.n650 146.341
R2330 vdd.n3551 vdd.n650 146.341
R2331 vdd.n3551 vdd.n643 146.341
R2332 vdd.n3562 vdd.n643 146.341
R2333 vdd.n3562 vdd.n639 146.341
R2334 vdd.n3571 vdd.n639 146.341
R2335 vdd.n3571 vdd.n632 146.341
R2336 vdd.n3581 vdd.n632 146.341
R2337 vdd.n3582 vdd.n3581 146.341
R2338 vdd.n3582 vdd.n341 146.341
R2339 vdd.n342 vdd.n341 146.341
R2340 vdd.n343 vdd.n342 146.341
R2341 vdd.n3589 vdd.n343 146.341
R2342 vdd.n3589 vdd.n351 146.341
R2343 vdd.n352 vdd.n351 146.341
R2344 vdd.n353 vdd.n352 146.341
R2345 vdd.n3596 vdd.n353 146.341
R2346 vdd.n3596 vdd.n362 146.341
R2347 vdd.n363 vdd.n362 146.341
R2348 vdd.n364 vdd.n363 146.341
R2349 vdd.n3604 vdd.n364 146.341
R2350 vdd.n3604 vdd.n372 146.341
R2351 vdd.n373 vdd.n372 146.341
R2352 vdd.n374 vdd.n373 146.341
R2353 vdd.n3611 vdd.n374 146.341
R2354 vdd.n3611 vdd.n383 146.341
R2355 vdd.n384 vdd.n383 146.341
R2356 vdd.n385 vdd.n384 146.341
R2357 vdd.n3618 vdd.n385 146.341
R2358 vdd.n3618 vdd.n393 146.341
R2359 vdd.n725 vdd.n724 146.341
R2360 vdd.n728 vdd.n724 146.341
R2361 vdd.n734 vdd.n733 146.341
R2362 vdd.n3484 vdd.n3483 146.341
R2363 vdd.n3480 vdd.n3479 146.341
R2364 vdd.n3476 vdd.n3475 146.341
R2365 vdd.n3472 vdd.n3471 146.341
R2366 vdd.n3468 vdd.n3467 146.341
R2367 vdd.n3464 vdd.n3463 146.341
R2368 vdd.n3460 vdd.n3459 146.341
R2369 vdd.n3451 vdd.n3450 146.341
R2370 vdd.n3448 vdd.n3447 146.341
R2371 vdd.n3444 vdd.n3443 146.341
R2372 vdd.n3440 vdd.n3439 146.341
R2373 vdd.n3436 vdd.n3435 146.341
R2374 vdd.n3432 vdd.n3431 146.341
R2375 vdd.n3428 vdd.n3427 146.341
R2376 vdd.n3424 vdd.n3423 146.341
R2377 vdd.n3420 vdd.n3419 146.341
R2378 vdd.n3416 vdd.n3415 146.341
R2379 vdd.n3412 vdd.n3411 146.341
R2380 vdd.n3405 vdd.n3404 146.341
R2381 vdd.n3402 vdd.n3401 146.341
R2382 vdd.n3398 vdd.n3397 146.341
R2383 vdd.n3394 vdd.n3393 146.341
R2384 vdd.n3390 vdd.n3389 146.341
R2385 vdd.n3386 vdd.n3385 146.341
R2386 vdd.n3382 vdd.n3381 146.341
R2387 vdd.n3378 vdd.n3377 146.341
R2388 vdd.n3374 vdd.n3373 146.341
R2389 vdd.n3370 vdd.n3369 146.341
R2390 vdd.n3496 vdd.n691 146.341
R2391 vdd.n3504 vdd.n684 146.341
R2392 vdd.n3504 vdd.n680 146.341
R2393 vdd.n3510 vdd.n680 146.341
R2394 vdd.n3510 vdd.n672 146.341
R2395 vdd.n3521 vdd.n672 146.341
R2396 vdd.n3521 vdd.n668 146.341
R2397 vdd.n3527 vdd.n668 146.341
R2398 vdd.n3527 vdd.n661 146.341
R2399 vdd.n3537 vdd.n661 146.341
R2400 vdd.n3537 vdd.n657 146.341
R2401 vdd.n3543 vdd.n657 146.341
R2402 vdd.n3543 vdd.n649 146.341
R2403 vdd.n3554 vdd.n649 146.341
R2404 vdd.n3554 vdd.n645 146.341
R2405 vdd.n3560 vdd.n645 146.341
R2406 vdd.n3560 vdd.n638 146.341
R2407 vdd.n3573 vdd.n638 146.341
R2408 vdd.n3573 vdd.n634 146.341
R2409 vdd.n3579 vdd.n634 146.341
R2410 vdd.n3579 vdd.n338 146.341
R2411 vdd.n3668 vdd.n338 146.341
R2412 vdd.n3668 vdd.n339 146.341
R2413 vdd.n3664 vdd.n339 146.341
R2414 vdd.n3664 vdd.n345 146.341
R2415 vdd.n3660 vdd.n345 146.341
R2416 vdd.n3660 vdd.n350 146.341
R2417 vdd.n3656 vdd.n350 146.341
R2418 vdd.n3656 vdd.n354 146.341
R2419 vdd.n3652 vdd.n354 146.341
R2420 vdd.n3652 vdd.n360 146.341
R2421 vdd.n3648 vdd.n360 146.341
R2422 vdd.n3648 vdd.n365 146.341
R2423 vdd.n3644 vdd.n365 146.341
R2424 vdd.n3644 vdd.n371 146.341
R2425 vdd.n3640 vdd.n371 146.341
R2426 vdd.n3640 vdd.n376 146.341
R2427 vdd.n3636 vdd.n376 146.341
R2428 vdd.n3636 vdd.n382 146.341
R2429 vdd.n3632 vdd.n382 146.341
R2430 vdd.n3632 vdd.n387 146.341
R2431 vdd.n3628 vdd.n387 146.341
R2432 vdd.n2471 vdd.n2470 146.341
R2433 vdd.n2468 vdd.n2465 146.341
R2434 vdd.n2463 vdd.n1185 146.341
R2435 vdd.n2459 vdd.n2458 146.341
R2436 vdd.n2456 vdd.n1189 146.341
R2437 vdd.n2452 vdd.n2451 146.341
R2438 vdd.n2449 vdd.n1196 146.341
R2439 vdd.n2445 vdd.n2444 146.341
R2440 vdd.n2442 vdd.n1203 146.341
R2441 vdd.n1214 vdd.n1211 146.341
R2442 vdd.n2434 vdd.n2433 146.341
R2443 vdd.n2431 vdd.n1216 146.341
R2444 vdd.n2427 vdd.n2426 146.341
R2445 vdd.n2424 vdd.n1222 146.341
R2446 vdd.n2420 vdd.n2419 146.341
R2447 vdd.n2417 vdd.n1229 146.341
R2448 vdd.n2413 vdd.n2412 146.341
R2449 vdd.n2410 vdd.n1236 146.341
R2450 vdd.n2406 vdd.n2405 146.341
R2451 vdd.n2403 vdd.n1243 146.341
R2452 vdd.n1254 vdd.n1251 146.341
R2453 vdd.n2395 vdd.n2394 146.341
R2454 vdd.n2392 vdd.n1256 146.341
R2455 vdd.n2388 vdd.n2387 146.341
R2456 vdd.n2385 vdd.n1262 146.341
R2457 vdd.n2381 vdd.n2380 146.341
R2458 vdd.n2378 vdd.n1269 146.341
R2459 vdd.n2374 vdd.n2373 146.341
R2460 vdd.n2371 vdd.n1276 146.341
R2461 vdd.n1522 vdd.n1520 146.341
R2462 vdd.n1525 vdd.n1524 146.341
R2463 vdd.n1883 vdd.n1643 146.341
R2464 vdd.n1883 vdd.n1639 146.341
R2465 vdd.n1889 vdd.n1639 146.341
R2466 vdd.n1889 vdd.n1631 146.341
R2467 vdd.n1900 vdd.n1631 146.341
R2468 vdd.n1900 vdd.n1627 146.341
R2469 vdd.n1906 vdd.n1627 146.341
R2470 vdd.n1906 vdd.n1621 146.341
R2471 vdd.n1917 vdd.n1621 146.341
R2472 vdd.n1917 vdd.n1617 146.341
R2473 vdd.n1923 vdd.n1617 146.341
R2474 vdd.n1923 vdd.n1608 146.341
R2475 vdd.n1933 vdd.n1608 146.341
R2476 vdd.n1933 vdd.n1604 146.341
R2477 vdd.n1939 vdd.n1604 146.341
R2478 vdd.n1939 vdd.n1597 146.341
R2479 vdd.n1950 vdd.n1597 146.341
R2480 vdd.n1950 vdd.n1593 146.341
R2481 vdd.n1956 vdd.n1593 146.341
R2482 vdd.n1956 vdd.n1586 146.341
R2483 vdd.n2273 vdd.n1586 146.341
R2484 vdd.n2273 vdd.n1582 146.341
R2485 vdd.n2279 vdd.n1582 146.341
R2486 vdd.n2279 vdd.n1574 146.341
R2487 vdd.n2290 vdd.n1574 146.341
R2488 vdd.n2290 vdd.n1570 146.341
R2489 vdd.n2296 vdd.n1570 146.341
R2490 vdd.n2296 vdd.n1564 146.341
R2491 vdd.n2307 vdd.n1564 146.341
R2492 vdd.n2307 vdd.n1560 146.341
R2493 vdd.n2313 vdd.n1560 146.341
R2494 vdd.n2313 vdd.n1551 146.341
R2495 vdd.n2323 vdd.n1551 146.341
R2496 vdd.n2323 vdd.n1547 146.341
R2497 vdd.n2329 vdd.n1547 146.341
R2498 vdd.n2329 vdd.n1541 146.341
R2499 vdd.n2340 vdd.n1541 146.341
R2500 vdd.n2340 vdd.n1536 146.341
R2501 vdd.n2348 vdd.n1536 146.341
R2502 vdd.n2348 vdd.n1527 146.341
R2503 vdd.n2359 vdd.n1527 146.341
R2504 vdd.n1872 vdd.n1648 146.341
R2505 vdd.n1872 vdd.n1681 146.341
R2506 vdd.n1685 vdd.n1684 146.341
R2507 vdd.n1687 vdd.n1686 146.341
R2508 vdd.n1691 vdd.n1690 146.341
R2509 vdd.n1693 vdd.n1692 146.341
R2510 vdd.n1697 vdd.n1696 146.341
R2511 vdd.n1699 vdd.n1698 146.341
R2512 vdd.n1703 vdd.n1702 146.341
R2513 vdd.n1705 vdd.n1704 146.341
R2514 vdd.n1711 vdd.n1710 146.341
R2515 vdd.n1713 vdd.n1712 146.341
R2516 vdd.n1717 vdd.n1716 146.341
R2517 vdd.n1719 vdd.n1718 146.341
R2518 vdd.n1723 vdd.n1722 146.341
R2519 vdd.n1725 vdd.n1724 146.341
R2520 vdd.n1729 vdd.n1728 146.341
R2521 vdd.n1731 vdd.n1730 146.341
R2522 vdd.n1735 vdd.n1734 146.341
R2523 vdd.n1737 vdd.n1736 146.341
R2524 vdd.n1809 vdd.n1740 146.341
R2525 vdd.n1742 vdd.n1741 146.341
R2526 vdd.n1746 vdd.n1745 146.341
R2527 vdd.n1748 vdd.n1747 146.341
R2528 vdd.n1752 vdd.n1751 146.341
R2529 vdd.n1754 vdd.n1753 146.341
R2530 vdd.n1758 vdd.n1757 146.341
R2531 vdd.n1760 vdd.n1759 146.341
R2532 vdd.n1764 vdd.n1763 146.341
R2533 vdd.n1766 vdd.n1765 146.341
R2534 vdd.n1770 vdd.n1769 146.341
R2535 vdd.n1771 vdd.n1679 146.341
R2536 vdd.n1881 vdd.n1644 146.341
R2537 vdd.n1881 vdd.n1637 146.341
R2538 vdd.n1892 vdd.n1637 146.341
R2539 vdd.n1892 vdd.n1633 146.341
R2540 vdd.n1898 vdd.n1633 146.341
R2541 vdd.n1898 vdd.n1626 146.341
R2542 vdd.n1909 vdd.n1626 146.341
R2543 vdd.n1909 vdd.n1622 146.341
R2544 vdd.n1915 vdd.n1622 146.341
R2545 vdd.n1915 vdd.n1615 146.341
R2546 vdd.n1925 vdd.n1615 146.341
R2547 vdd.n1925 vdd.n1611 146.341
R2548 vdd.n1931 vdd.n1611 146.341
R2549 vdd.n1931 vdd.n1603 146.341
R2550 vdd.n1942 vdd.n1603 146.341
R2551 vdd.n1942 vdd.n1599 146.341
R2552 vdd.n1948 vdd.n1599 146.341
R2553 vdd.n1948 vdd.n1592 146.341
R2554 vdd.n1958 vdd.n1592 146.341
R2555 vdd.n1958 vdd.n1588 146.341
R2556 vdd.n2271 vdd.n1588 146.341
R2557 vdd.n2271 vdd.n1580 146.341
R2558 vdd.n2282 vdd.n1580 146.341
R2559 vdd.n2282 vdd.n1576 146.341
R2560 vdd.n2288 vdd.n1576 146.341
R2561 vdd.n2288 vdd.n1569 146.341
R2562 vdd.n2299 vdd.n1569 146.341
R2563 vdd.n2299 vdd.n1565 146.341
R2564 vdd.n2305 vdd.n1565 146.341
R2565 vdd.n2305 vdd.n1558 146.341
R2566 vdd.n2315 vdd.n1558 146.341
R2567 vdd.n2315 vdd.n1554 146.341
R2568 vdd.n2321 vdd.n1554 146.341
R2569 vdd.n2321 vdd.n1546 146.341
R2570 vdd.n2332 vdd.n1546 146.341
R2571 vdd.n2332 vdd.n1542 146.341
R2572 vdd.n2338 vdd.n1542 146.341
R2573 vdd.n2338 vdd.n1534 146.341
R2574 vdd.n2351 vdd.n1534 146.341
R2575 vdd.n2351 vdd.n1529 146.341
R2576 vdd.n2357 vdd.n1529 146.341
R2577 vdd.n1315 vdd.t239 127.284
R2578 vdd.n1010 vdd.t279 127.284
R2579 vdd.n1319 vdd.t276 127.284
R2580 vdd.n1001 vdd.t300 127.284
R2581 vdd.n896 vdd.t263 127.284
R2582 vdd.n896 vdd.t264 127.284
R2583 vdd.n2823 vdd.t294 127.284
R2584 vdd.n832 vdd.t255 127.284
R2585 vdd.n2820 vdd.t287 127.284
R2586 vdd.n799 vdd.t234 127.284
R2587 vdd.n1071 vdd.t290 127.284
R2588 vdd.n1071 vdd.t291 127.284
R2589 vdd.n22 vdd.n20 117.314
R2590 vdd.n17 vdd.n15 117.314
R2591 vdd.n27 vdd.n26 116.927
R2592 vdd.n24 vdd.n23 116.927
R2593 vdd.n22 vdd.n21 116.927
R2594 vdd.n17 vdd.n16 116.927
R2595 vdd.n19 vdd.n18 116.927
R2596 vdd.n27 vdd.n25 116.927
R2597 vdd.n1316 vdd.t238 111.188
R2598 vdd.n1011 vdd.t280 111.188
R2599 vdd.n1320 vdd.t275 111.188
R2600 vdd.n1002 vdd.t301 111.188
R2601 vdd.n2824 vdd.t293 111.188
R2602 vdd.n833 vdd.t256 111.188
R2603 vdd.n2821 vdd.t286 111.188
R2604 vdd.n800 vdd.t235 111.188
R2605 vdd.n3094 vdd.n960 99.5127
R2606 vdd.n3094 vdd.n951 99.5127
R2607 vdd.n3102 vdd.n951 99.5127
R2608 vdd.n3102 vdd.n949 99.5127
R2609 vdd.n3106 vdd.n949 99.5127
R2610 vdd.n3106 vdd.n939 99.5127
R2611 vdd.n3114 vdd.n939 99.5127
R2612 vdd.n3114 vdd.n937 99.5127
R2613 vdd.n3118 vdd.n937 99.5127
R2614 vdd.n3118 vdd.n928 99.5127
R2615 vdd.n3126 vdd.n928 99.5127
R2616 vdd.n3126 vdd.n926 99.5127
R2617 vdd.n3130 vdd.n926 99.5127
R2618 vdd.n3130 vdd.n917 99.5127
R2619 vdd.n3138 vdd.n917 99.5127
R2620 vdd.n3138 vdd.n915 99.5127
R2621 vdd.n3142 vdd.n915 99.5127
R2622 vdd.n3142 vdd.n904 99.5127
R2623 vdd.n3151 vdd.n904 99.5127
R2624 vdd.n3151 vdd.n902 99.5127
R2625 vdd.n3155 vdd.n902 99.5127
R2626 vdd.n3155 vdd.n892 99.5127
R2627 vdd.n3163 vdd.n892 99.5127
R2628 vdd.n3163 vdd.n890 99.5127
R2629 vdd.n3167 vdd.n890 99.5127
R2630 vdd.n3167 vdd.n880 99.5127
R2631 vdd.n3175 vdd.n880 99.5127
R2632 vdd.n3175 vdd.n878 99.5127
R2633 vdd.n3179 vdd.n878 99.5127
R2634 vdd.n3179 vdd.n867 99.5127
R2635 vdd.n3187 vdd.n867 99.5127
R2636 vdd.n3187 vdd.n865 99.5127
R2637 vdd.n3191 vdd.n865 99.5127
R2638 vdd.n3191 vdd.n856 99.5127
R2639 vdd.n3199 vdd.n856 99.5127
R2640 vdd.n3199 vdd.n854 99.5127
R2641 vdd.n3203 vdd.n854 99.5127
R2642 vdd.n3203 vdd.n842 99.5127
R2643 vdd.n3256 vdd.n842 99.5127
R2644 vdd.n3256 vdd.n840 99.5127
R2645 vdd.n3260 vdd.n840 99.5127
R2646 vdd.n3260 vdd.n808 99.5127
R2647 vdd.n3330 vdd.n808 99.5127
R2648 vdd.n3326 vdd.n809 99.5127
R2649 vdd.n3324 vdd.n3323 99.5127
R2650 vdd.n3321 vdd.n813 99.5127
R2651 vdd.n3317 vdd.n3316 99.5127
R2652 vdd.n3314 vdd.n816 99.5127
R2653 vdd.n3310 vdd.n3309 99.5127
R2654 vdd.n3307 vdd.n819 99.5127
R2655 vdd.n3303 vdd.n3302 99.5127
R2656 vdd.n3300 vdd.n3298 99.5127
R2657 vdd.n3296 vdd.n822 99.5127
R2658 vdd.n3292 vdd.n3291 99.5127
R2659 vdd.n3289 vdd.n825 99.5127
R2660 vdd.n3285 vdd.n3284 99.5127
R2661 vdd.n3282 vdd.n828 99.5127
R2662 vdd.n3278 vdd.n3277 99.5127
R2663 vdd.n3275 vdd.n831 99.5127
R2664 vdd.n3270 vdd.n3269 99.5127
R2665 vdd.n3021 vdd.n958 99.5127
R2666 vdd.n3017 vdd.n958 99.5127
R2667 vdd.n3017 vdd.n952 99.5127
R2668 vdd.n2899 vdd.n952 99.5127
R2669 vdd.n2899 vdd.n947 99.5127
R2670 vdd.n2902 vdd.n947 99.5127
R2671 vdd.n2902 vdd.n941 99.5127
R2672 vdd.n3003 vdd.n941 99.5127
R2673 vdd.n3003 vdd.n935 99.5127
R2674 vdd.n2999 vdd.n935 99.5127
R2675 vdd.n2999 vdd.n929 99.5127
R2676 vdd.n2946 vdd.n929 99.5127
R2677 vdd.n2946 vdd.n923 99.5127
R2678 vdd.n2943 vdd.n923 99.5127
R2679 vdd.n2943 vdd.n918 99.5127
R2680 vdd.n2940 vdd.n918 99.5127
R2681 vdd.n2940 vdd.n913 99.5127
R2682 vdd.n2937 vdd.n913 99.5127
R2683 vdd.n2937 vdd.n906 99.5127
R2684 vdd.n2934 vdd.n906 99.5127
R2685 vdd.n2934 vdd.n899 99.5127
R2686 vdd.n2931 vdd.n899 99.5127
R2687 vdd.n2931 vdd.n893 99.5127
R2688 vdd.n2928 vdd.n893 99.5127
R2689 vdd.n2928 vdd.n888 99.5127
R2690 vdd.n2925 vdd.n888 99.5127
R2691 vdd.n2925 vdd.n882 99.5127
R2692 vdd.n2922 vdd.n882 99.5127
R2693 vdd.n2922 vdd.n875 99.5127
R2694 vdd.n2919 vdd.n875 99.5127
R2695 vdd.n2919 vdd.n868 99.5127
R2696 vdd.n2916 vdd.n868 99.5127
R2697 vdd.n2916 vdd.n862 99.5127
R2698 vdd.n2913 vdd.n862 99.5127
R2699 vdd.n2913 vdd.n857 99.5127
R2700 vdd.n2910 vdd.n857 99.5127
R2701 vdd.n2910 vdd.n852 99.5127
R2702 vdd.n2907 vdd.n852 99.5127
R2703 vdd.n2907 vdd.n844 99.5127
R2704 vdd.n844 vdd.n837 99.5127
R2705 vdd.n3262 vdd.n837 99.5127
R2706 vdd.n3263 vdd.n3262 99.5127
R2707 vdd.n3263 vdd.n806 99.5127
R2708 vdd.n3087 vdd.n962 99.5127
R2709 vdd.n3087 vdd.n2819 99.5127
R2710 vdd.n3083 vdd.n3082 99.5127
R2711 vdd.n3079 vdd.n3078 99.5127
R2712 vdd.n3075 vdd.n3074 99.5127
R2713 vdd.n3071 vdd.n3070 99.5127
R2714 vdd.n3067 vdd.n3066 99.5127
R2715 vdd.n3063 vdd.n3062 99.5127
R2716 vdd.n3059 vdd.n3058 99.5127
R2717 vdd.n3055 vdd.n3054 99.5127
R2718 vdd.n3051 vdd.n3050 99.5127
R2719 vdd.n3047 vdd.n3046 99.5127
R2720 vdd.n3043 vdd.n3042 99.5127
R2721 vdd.n3039 vdd.n3038 99.5127
R2722 vdd.n3035 vdd.n3034 99.5127
R2723 vdd.n3031 vdd.n3030 99.5127
R2724 vdd.n3026 vdd.n3025 99.5127
R2725 vdd.n2783 vdd.n999 99.5127
R2726 vdd.n2779 vdd.n2778 99.5127
R2727 vdd.n2775 vdd.n2774 99.5127
R2728 vdd.n2771 vdd.n2770 99.5127
R2729 vdd.n2767 vdd.n2766 99.5127
R2730 vdd.n2763 vdd.n2762 99.5127
R2731 vdd.n2759 vdd.n2758 99.5127
R2732 vdd.n2755 vdd.n2754 99.5127
R2733 vdd.n2751 vdd.n2750 99.5127
R2734 vdd.n2747 vdd.n2746 99.5127
R2735 vdd.n2743 vdd.n2742 99.5127
R2736 vdd.n2739 vdd.n2738 99.5127
R2737 vdd.n2735 vdd.n2734 99.5127
R2738 vdd.n2731 vdd.n2730 99.5127
R2739 vdd.n2727 vdd.n2726 99.5127
R2740 vdd.n2723 vdd.n2722 99.5127
R2741 vdd.n2718 vdd.n2717 99.5127
R2742 vdd.n1355 vdd.n1135 99.5127
R2743 vdd.n1358 vdd.n1135 99.5127
R2744 vdd.n1358 vdd.n1129 99.5127
R2745 vdd.n1361 vdd.n1129 99.5127
R2746 vdd.n1361 vdd.n1124 99.5127
R2747 vdd.n1364 vdd.n1124 99.5127
R2748 vdd.n1364 vdd.n1117 99.5127
R2749 vdd.n1367 vdd.n1117 99.5127
R2750 vdd.n1367 vdd.n1110 99.5127
R2751 vdd.n1370 vdd.n1110 99.5127
R2752 vdd.n1370 vdd.n1104 99.5127
R2753 vdd.n1373 vdd.n1104 99.5127
R2754 vdd.n1373 vdd.n1099 99.5127
R2755 vdd.n1376 vdd.n1099 99.5127
R2756 vdd.n1376 vdd.n1094 99.5127
R2757 vdd.n1379 vdd.n1094 99.5127
R2758 vdd.n1379 vdd.n1088 99.5127
R2759 vdd.n1382 vdd.n1088 99.5127
R2760 vdd.n1382 vdd.n1081 99.5127
R2761 vdd.n1385 vdd.n1081 99.5127
R2762 vdd.n1385 vdd.n1074 99.5127
R2763 vdd.n1388 vdd.n1074 99.5127
R2764 vdd.n1388 vdd.n1068 99.5127
R2765 vdd.n1391 vdd.n1068 99.5127
R2766 vdd.n1391 vdd.n1063 99.5127
R2767 vdd.n1394 vdd.n1063 99.5127
R2768 vdd.n1394 vdd.n1057 99.5127
R2769 vdd.n1436 vdd.n1057 99.5127
R2770 vdd.n1436 vdd.n1050 99.5127
R2771 vdd.n1432 vdd.n1050 99.5127
R2772 vdd.n1432 vdd.n1044 99.5127
R2773 vdd.n1429 vdd.n1044 99.5127
R2774 vdd.n1429 vdd.n1039 99.5127
R2775 vdd.n1426 vdd.n1039 99.5127
R2776 vdd.n1426 vdd.n1034 99.5127
R2777 vdd.n1406 vdd.n1034 99.5127
R2778 vdd.n1406 vdd.n1029 99.5127
R2779 vdd.n1403 vdd.n1029 99.5127
R2780 vdd.n1403 vdd.n1022 99.5127
R2781 vdd.n1400 vdd.n1022 99.5127
R2782 vdd.n1400 vdd.n1015 99.5127
R2783 vdd.n1015 vdd.n1004 99.5127
R2784 vdd.n2713 vdd.n1004 99.5127
R2785 vdd.n2505 vdd.n1140 99.5127
R2786 vdd.n2505 vdd.n1176 99.5127
R2787 vdd.n2501 vdd.n2500 99.5127
R2788 vdd.n2497 vdd.n2496 99.5127
R2789 vdd.n2493 vdd.n2492 99.5127
R2790 vdd.n2489 vdd.n2488 99.5127
R2791 vdd.n2485 vdd.n2484 99.5127
R2792 vdd.n2481 vdd.n2480 99.5127
R2793 vdd.n2477 vdd.n2476 99.5127
R2794 vdd.n1322 vdd.n1321 99.5127
R2795 vdd.n1326 vdd.n1325 99.5127
R2796 vdd.n1330 vdd.n1329 99.5127
R2797 vdd.n1334 vdd.n1333 99.5127
R2798 vdd.n1338 vdd.n1337 99.5127
R2799 vdd.n1342 vdd.n1341 99.5127
R2800 vdd.n1346 vdd.n1345 99.5127
R2801 vdd.n1351 vdd.n1350 99.5127
R2802 vdd.n2512 vdd.n1138 99.5127
R2803 vdd.n2512 vdd.n1128 99.5127
R2804 vdd.n2520 vdd.n1128 99.5127
R2805 vdd.n2520 vdd.n1126 99.5127
R2806 vdd.n2524 vdd.n1126 99.5127
R2807 vdd.n2524 vdd.n1115 99.5127
R2808 vdd.n2532 vdd.n1115 99.5127
R2809 vdd.n2532 vdd.n1113 99.5127
R2810 vdd.n2536 vdd.n1113 99.5127
R2811 vdd.n2536 vdd.n1103 99.5127
R2812 vdd.n2544 vdd.n1103 99.5127
R2813 vdd.n2544 vdd.n1101 99.5127
R2814 vdd.n2548 vdd.n1101 99.5127
R2815 vdd.n2548 vdd.n1092 99.5127
R2816 vdd.n2556 vdd.n1092 99.5127
R2817 vdd.n2556 vdd.n1090 99.5127
R2818 vdd.n2560 vdd.n1090 99.5127
R2819 vdd.n2560 vdd.n1079 99.5127
R2820 vdd.n2568 vdd.n1079 99.5127
R2821 vdd.n2568 vdd.n1077 99.5127
R2822 vdd.n2572 vdd.n1077 99.5127
R2823 vdd.n2572 vdd.n1067 99.5127
R2824 vdd.n2581 vdd.n1067 99.5127
R2825 vdd.n2581 vdd.n1065 99.5127
R2826 vdd.n2585 vdd.n1065 99.5127
R2827 vdd.n2585 vdd.n1055 99.5127
R2828 vdd.n2593 vdd.n1055 99.5127
R2829 vdd.n2593 vdd.n1053 99.5127
R2830 vdd.n2597 vdd.n1053 99.5127
R2831 vdd.n2597 vdd.n1043 99.5127
R2832 vdd.n2605 vdd.n1043 99.5127
R2833 vdd.n2605 vdd.n1041 99.5127
R2834 vdd.n2609 vdd.n1041 99.5127
R2835 vdd.n2609 vdd.n1033 99.5127
R2836 vdd.n2617 vdd.n1033 99.5127
R2837 vdd.n2617 vdd.n1031 99.5127
R2838 vdd.n2621 vdd.n1031 99.5127
R2839 vdd.n2621 vdd.n1020 99.5127
R2840 vdd.n2631 vdd.n1020 99.5127
R2841 vdd.n2631 vdd.n1017 99.5127
R2842 vdd.n2636 vdd.n1017 99.5127
R2843 vdd.n2636 vdd.n1018 99.5127
R2844 vdd.n1018 vdd.n998 99.5127
R2845 vdd.n3246 vdd.n3245 99.5127
R2846 vdd.n3243 vdd.n3209 99.5127
R2847 vdd.n3239 vdd.n3238 99.5127
R2848 vdd.n3236 vdd.n3212 99.5127
R2849 vdd.n3232 vdd.n3231 99.5127
R2850 vdd.n3229 vdd.n3215 99.5127
R2851 vdd.n3225 vdd.n3224 99.5127
R2852 vdd.n3222 vdd.n3219 99.5127
R2853 vdd.n3363 vdd.n787 99.5127
R2854 vdd.n3361 vdd.n3360 99.5127
R2855 vdd.n3358 vdd.n789 99.5127
R2856 vdd.n3354 vdd.n3353 99.5127
R2857 vdd.n3351 vdd.n792 99.5127
R2858 vdd.n3347 vdd.n3346 99.5127
R2859 vdd.n3344 vdd.n795 99.5127
R2860 vdd.n3340 vdd.n3339 99.5127
R2861 vdd.n3337 vdd.n798 99.5127
R2862 vdd.n2895 vdd.n959 99.5127
R2863 vdd.n3015 vdd.n959 99.5127
R2864 vdd.n3015 vdd.n953 99.5127
R2865 vdd.n3011 vdd.n953 99.5127
R2866 vdd.n3011 vdd.n948 99.5127
R2867 vdd.n3008 vdd.n948 99.5127
R2868 vdd.n3008 vdd.n942 99.5127
R2869 vdd.n3005 vdd.n942 99.5127
R2870 vdd.n3005 vdd.n936 99.5127
R2871 vdd.n2997 vdd.n936 99.5127
R2872 vdd.n2997 vdd.n930 99.5127
R2873 vdd.n2993 vdd.n930 99.5127
R2874 vdd.n2993 vdd.n924 99.5127
R2875 vdd.n2990 vdd.n924 99.5127
R2876 vdd.n2990 vdd.n919 99.5127
R2877 vdd.n2987 vdd.n919 99.5127
R2878 vdd.n2987 vdd.n914 99.5127
R2879 vdd.n2984 vdd.n914 99.5127
R2880 vdd.n2984 vdd.n907 99.5127
R2881 vdd.n2981 vdd.n907 99.5127
R2882 vdd.n2981 vdd.n900 99.5127
R2883 vdd.n2978 vdd.n900 99.5127
R2884 vdd.n2978 vdd.n894 99.5127
R2885 vdd.n2975 vdd.n894 99.5127
R2886 vdd.n2975 vdd.n889 99.5127
R2887 vdd.n2972 vdd.n889 99.5127
R2888 vdd.n2972 vdd.n883 99.5127
R2889 vdd.n2969 vdd.n883 99.5127
R2890 vdd.n2969 vdd.n876 99.5127
R2891 vdd.n2966 vdd.n876 99.5127
R2892 vdd.n2966 vdd.n869 99.5127
R2893 vdd.n2963 vdd.n869 99.5127
R2894 vdd.n2963 vdd.n863 99.5127
R2895 vdd.n2960 vdd.n863 99.5127
R2896 vdd.n2960 vdd.n858 99.5127
R2897 vdd.n2957 vdd.n858 99.5127
R2898 vdd.n2957 vdd.n853 99.5127
R2899 vdd.n2954 vdd.n853 99.5127
R2900 vdd.n2954 vdd.n845 99.5127
R2901 vdd.n2951 vdd.n845 99.5127
R2902 vdd.n2951 vdd.n838 99.5127
R2903 vdd.n838 vdd.n804 99.5127
R2904 vdd.n3332 vdd.n804 99.5127
R2905 vdd.n2830 vdd.n2829 99.5127
R2906 vdd.n2834 vdd.n2833 99.5127
R2907 vdd.n2838 vdd.n2837 99.5127
R2908 vdd.n2842 vdd.n2841 99.5127
R2909 vdd.n2846 vdd.n2845 99.5127
R2910 vdd.n2850 vdd.n2849 99.5127
R2911 vdd.n2854 vdd.n2853 99.5127
R2912 vdd.n2858 vdd.n2857 99.5127
R2913 vdd.n2862 vdd.n2861 99.5127
R2914 vdd.n2866 vdd.n2865 99.5127
R2915 vdd.n2870 vdd.n2869 99.5127
R2916 vdd.n2874 vdd.n2873 99.5127
R2917 vdd.n2878 vdd.n2877 99.5127
R2918 vdd.n2882 vdd.n2881 99.5127
R2919 vdd.n2886 vdd.n2885 99.5127
R2920 vdd.n2890 vdd.n2889 99.5127
R2921 vdd.n2892 vdd.n2818 99.5127
R2922 vdd.n3096 vdd.n956 99.5127
R2923 vdd.n3096 vdd.n954 99.5127
R2924 vdd.n3100 vdd.n954 99.5127
R2925 vdd.n3100 vdd.n945 99.5127
R2926 vdd.n3108 vdd.n945 99.5127
R2927 vdd.n3108 vdd.n943 99.5127
R2928 vdd.n3112 vdd.n943 99.5127
R2929 vdd.n3112 vdd.n934 99.5127
R2930 vdd.n3120 vdd.n934 99.5127
R2931 vdd.n3120 vdd.n932 99.5127
R2932 vdd.n3124 vdd.n932 99.5127
R2933 vdd.n3124 vdd.n922 99.5127
R2934 vdd.n3132 vdd.n922 99.5127
R2935 vdd.n3132 vdd.n920 99.5127
R2936 vdd.n3136 vdd.n920 99.5127
R2937 vdd.n3136 vdd.n911 99.5127
R2938 vdd.n3144 vdd.n911 99.5127
R2939 vdd.n3144 vdd.n909 99.5127
R2940 vdd.n3149 vdd.n909 99.5127
R2941 vdd.n3149 vdd.n898 99.5127
R2942 vdd.n3157 vdd.n898 99.5127
R2943 vdd.n3157 vdd.n895 99.5127
R2944 vdd.n3161 vdd.n895 99.5127
R2945 vdd.n3161 vdd.n886 99.5127
R2946 vdd.n3169 vdd.n886 99.5127
R2947 vdd.n3169 vdd.n884 99.5127
R2948 vdd.n3173 vdd.n884 99.5127
R2949 vdd.n3173 vdd.n873 99.5127
R2950 vdd.n3181 vdd.n873 99.5127
R2951 vdd.n3181 vdd.n871 99.5127
R2952 vdd.n3185 vdd.n871 99.5127
R2953 vdd.n3185 vdd.n861 99.5127
R2954 vdd.n3193 vdd.n861 99.5127
R2955 vdd.n3193 vdd.n859 99.5127
R2956 vdd.n3197 vdd.n859 99.5127
R2957 vdd.n3197 vdd.n850 99.5127
R2958 vdd.n3205 vdd.n850 99.5127
R2959 vdd.n3205 vdd.n847 99.5127
R2960 vdd.n3254 vdd.n847 99.5127
R2961 vdd.n3254 vdd.n848 99.5127
R2962 vdd.n848 vdd.n839 99.5127
R2963 vdd.n3249 vdd.n839 99.5127
R2964 vdd.n3249 vdd.n807 99.5127
R2965 vdd.n2707 vdd.n2706 99.5127
R2966 vdd.n2703 vdd.n2702 99.5127
R2967 vdd.n2699 vdd.n2698 99.5127
R2968 vdd.n2695 vdd.n2694 99.5127
R2969 vdd.n2691 vdd.n2690 99.5127
R2970 vdd.n2687 vdd.n2686 99.5127
R2971 vdd.n2683 vdd.n2682 99.5127
R2972 vdd.n2679 vdd.n2678 99.5127
R2973 vdd.n2675 vdd.n2674 99.5127
R2974 vdd.n2671 vdd.n2670 99.5127
R2975 vdd.n2667 vdd.n2666 99.5127
R2976 vdd.n2663 vdd.n2662 99.5127
R2977 vdd.n2659 vdd.n2658 99.5127
R2978 vdd.n2655 vdd.n2654 99.5127
R2979 vdd.n2651 vdd.n2650 99.5127
R2980 vdd.n2647 vdd.n2646 99.5127
R2981 vdd.n2643 vdd.n980 99.5127
R2982 vdd.n1480 vdd.n1136 99.5127
R2983 vdd.n1477 vdd.n1136 99.5127
R2984 vdd.n1477 vdd.n1130 99.5127
R2985 vdd.n1474 vdd.n1130 99.5127
R2986 vdd.n1474 vdd.n1125 99.5127
R2987 vdd.n1471 vdd.n1125 99.5127
R2988 vdd.n1471 vdd.n1118 99.5127
R2989 vdd.n1468 vdd.n1118 99.5127
R2990 vdd.n1468 vdd.n1111 99.5127
R2991 vdd.n1465 vdd.n1111 99.5127
R2992 vdd.n1465 vdd.n1105 99.5127
R2993 vdd.n1462 vdd.n1105 99.5127
R2994 vdd.n1462 vdd.n1100 99.5127
R2995 vdd.n1459 vdd.n1100 99.5127
R2996 vdd.n1459 vdd.n1095 99.5127
R2997 vdd.n1456 vdd.n1095 99.5127
R2998 vdd.n1456 vdd.n1089 99.5127
R2999 vdd.n1453 vdd.n1089 99.5127
R3000 vdd.n1453 vdd.n1082 99.5127
R3001 vdd.n1450 vdd.n1082 99.5127
R3002 vdd.n1450 vdd.n1075 99.5127
R3003 vdd.n1447 vdd.n1075 99.5127
R3004 vdd.n1447 vdd.n1069 99.5127
R3005 vdd.n1444 vdd.n1069 99.5127
R3006 vdd.n1444 vdd.n1064 99.5127
R3007 vdd.n1441 vdd.n1064 99.5127
R3008 vdd.n1441 vdd.n1058 99.5127
R3009 vdd.n1438 vdd.n1058 99.5127
R3010 vdd.n1438 vdd.n1051 99.5127
R3011 vdd.n1409 vdd.n1051 99.5127
R3012 vdd.n1409 vdd.n1045 99.5127
R3013 vdd.n1412 vdd.n1045 99.5127
R3014 vdd.n1412 vdd.n1040 99.5127
R3015 vdd.n1424 vdd.n1040 99.5127
R3016 vdd.n1424 vdd.n1035 99.5127
R3017 vdd.n1420 vdd.n1035 99.5127
R3018 vdd.n1420 vdd.n1030 99.5127
R3019 vdd.n1417 vdd.n1030 99.5127
R3020 vdd.n1417 vdd.n1023 99.5127
R3021 vdd.n1023 vdd.n1014 99.5127
R3022 vdd.n2638 vdd.n1014 99.5127
R3023 vdd.n2639 vdd.n2638 99.5127
R3024 vdd.n2639 vdd.n1006 99.5127
R3025 vdd.n1284 vdd.n1283 99.5127
R3026 vdd.n1288 vdd.n1287 99.5127
R3027 vdd.n1292 vdd.n1291 99.5127
R3028 vdd.n1296 vdd.n1295 99.5127
R3029 vdd.n1300 vdd.n1299 99.5127
R3030 vdd.n1304 vdd.n1303 99.5127
R3031 vdd.n1308 vdd.n1307 99.5127
R3032 vdd.n1312 vdd.n1311 99.5127
R3033 vdd.n1513 vdd.n1314 99.5127
R3034 vdd.n1511 vdd.n1510 99.5127
R3035 vdd.n1507 vdd.n1506 99.5127
R3036 vdd.n1503 vdd.n1502 99.5127
R3037 vdd.n1499 vdd.n1498 99.5127
R3038 vdd.n1495 vdd.n1494 99.5127
R3039 vdd.n1491 vdd.n1490 99.5127
R3040 vdd.n1487 vdd.n1486 99.5127
R3041 vdd.n1483 vdd.n1175 99.5127
R3042 vdd.n2514 vdd.n1133 99.5127
R3043 vdd.n2514 vdd.n1131 99.5127
R3044 vdd.n2518 vdd.n1131 99.5127
R3045 vdd.n2518 vdd.n1122 99.5127
R3046 vdd.n2526 vdd.n1122 99.5127
R3047 vdd.n2526 vdd.n1120 99.5127
R3048 vdd.n2530 vdd.n1120 99.5127
R3049 vdd.n2530 vdd.n1109 99.5127
R3050 vdd.n2538 vdd.n1109 99.5127
R3051 vdd.n2538 vdd.n1107 99.5127
R3052 vdd.n2542 vdd.n1107 99.5127
R3053 vdd.n2542 vdd.n1098 99.5127
R3054 vdd.n2550 vdd.n1098 99.5127
R3055 vdd.n2550 vdd.n1096 99.5127
R3056 vdd.n2554 vdd.n1096 99.5127
R3057 vdd.n2554 vdd.n1086 99.5127
R3058 vdd.n2562 vdd.n1086 99.5127
R3059 vdd.n2562 vdd.n1084 99.5127
R3060 vdd.n2566 vdd.n1084 99.5127
R3061 vdd.n2566 vdd.n1073 99.5127
R3062 vdd.n2574 vdd.n1073 99.5127
R3063 vdd.n2574 vdd.n1070 99.5127
R3064 vdd.n2579 vdd.n1070 99.5127
R3065 vdd.n2579 vdd.n1061 99.5127
R3066 vdd.n2587 vdd.n1061 99.5127
R3067 vdd.n2587 vdd.n1059 99.5127
R3068 vdd.n2591 vdd.n1059 99.5127
R3069 vdd.n2591 vdd.n1049 99.5127
R3070 vdd.n2599 vdd.n1049 99.5127
R3071 vdd.n2599 vdd.n1047 99.5127
R3072 vdd.n2603 vdd.n1047 99.5127
R3073 vdd.n2603 vdd.n1038 99.5127
R3074 vdd.n2611 vdd.n1038 99.5127
R3075 vdd.n2611 vdd.n1036 99.5127
R3076 vdd.n2615 vdd.n1036 99.5127
R3077 vdd.n2615 vdd.n1027 99.5127
R3078 vdd.n2623 vdd.n1027 99.5127
R3079 vdd.n2623 vdd.n1024 99.5127
R3080 vdd.n2629 vdd.n1024 99.5127
R3081 vdd.n2629 vdd.n1025 99.5127
R3082 vdd.n1025 vdd.n1016 99.5127
R3083 vdd.n1016 vdd.n1007 99.5127
R3084 vdd.n2711 vdd.n1007 99.5127
R3085 vdd.n9 vdd.n7 98.9633
R3086 vdd.n2 vdd.n0 98.9633
R3087 vdd.n9 vdd.n8 98.6055
R3088 vdd.n11 vdd.n10 98.6055
R3089 vdd.n13 vdd.n12 98.6055
R3090 vdd.n6 vdd.n5 98.6055
R3091 vdd.n4 vdd.n3 98.6055
R3092 vdd.n2 vdd.n1 98.6055
R3093 vdd.t62 vdd.n303 85.8723
R3094 vdd.t71 vdd.n244 85.8723
R3095 vdd.t198 vdd.n201 85.8723
R3096 vdd.t138 vdd.n142 85.8723
R3097 vdd.t24 vdd.n100 85.8723
R3098 vdd.t14 vdd.n41 85.8723
R3099 vdd.t57 vdd.n2177 85.8723
R3100 vdd.t206 vdd.n2236 85.8723
R3101 vdd.t223 vdd.n2075 85.8723
R3102 vdd.t101 vdd.n2134 85.8723
R3103 vdd.t35 vdd.n1974 85.8723
R3104 vdd.t22 vdd.n2033 85.8723
R3105 vdd.n897 vdd.n896 78.546
R3106 vdd.n2577 vdd.n1071 78.546
R3107 vdd.n290 vdd.n289 75.1835
R3108 vdd.n288 vdd.n287 75.1835
R3109 vdd.n286 vdd.n285 75.1835
R3110 vdd.n284 vdd.n283 75.1835
R3111 vdd.n282 vdd.n281 75.1835
R3112 vdd.n280 vdd.n279 75.1835
R3113 vdd.n278 vdd.n277 75.1835
R3114 vdd.n276 vdd.n275 75.1835
R3115 vdd.n274 vdd.n273 75.1835
R3116 vdd.n188 vdd.n187 75.1835
R3117 vdd.n186 vdd.n185 75.1835
R3118 vdd.n184 vdd.n183 75.1835
R3119 vdd.n182 vdd.n181 75.1835
R3120 vdd.n180 vdd.n179 75.1835
R3121 vdd.n178 vdd.n177 75.1835
R3122 vdd.n176 vdd.n175 75.1835
R3123 vdd.n174 vdd.n173 75.1835
R3124 vdd.n172 vdd.n171 75.1835
R3125 vdd.n87 vdd.n86 75.1835
R3126 vdd.n85 vdd.n84 75.1835
R3127 vdd.n83 vdd.n82 75.1835
R3128 vdd.n81 vdd.n80 75.1835
R3129 vdd.n79 vdd.n78 75.1835
R3130 vdd.n77 vdd.n76 75.1835
R3131 vdd.n75 vdd.n74 75.1835
R3132 vdd.n73 vdd.n72 75.1835
R3133 vdd.n71 vdd.n70 75.1835
R3134 vdd.n2207 vdd.n2206 75.1835
R3135 vdd.n2209 vdd.n2208 75.1835
R3136 vdd.n2211 vdd.n2210 75.1835
R3137 vdd.n2213 vdd.n2212 75.1835
R3138 vdd.n2215 vdd.n2214 75.1835
R3139 vdd.n2217 vdd.n2216 75.1835
R3140 vdd.n2219 vdd.n2218 75.1835
R3141 vdd.n2221 vdd.n2220 75.1835
R3142 vdd.n2223 vdd.n2222 75.1835
R3143 vdd.n2105 vdd.n2104 75.1835
R3144 vdd.n2107 vdd.n2106 75.1835
R3145 vdd.n2109 vdd.n2108 75.1835
R3146 vdd.n2111 vdd.n2110 75.1835
R3147 vdd.n2113 vdd.n2112 75.1835
R3148 vdd.n2115 vdd.n2114 75.1835
R3149 vdd.n2117 vdd.n2116 75.1835
R3150 vdd.n2119 vdd.n2118 75.1835
R3151 vdd.n2121 vdd.n2120 75.1835
R3152 vdd.n2004 vdd.n2003 75.1835
R3153 vdd.n2006 vdd.n2005 75.1835
R3154 vdd.n2008 vdd.n2007 75.1835
R3155 vdd.n2010 vdd.n2009 75.1835
R3156 vdd.n2012 vdd.n2011 75.1835
R3157 vdd.n2014 vdd.n2013 75.1835
R3158 vdd.n2016 vdd.n2015 75.1835
R3159 vdd.n2018 vdd.n2017 75.1835
R3160 vdd.n2020 vdd.n2019 75.1835
R3161 vdd.n3088 vdd.n2801 72.8958
R3162 vdd.n3088 vdd.n2802 72.8958
R3163 vdd.n3088 vdd.n2803 72.8958
R3164 vdd.n3088 vdd.n2804 72.8958
R3165 vdd.n3088 vdd.n2805 72.8958
R3166 vdd.n3088 vdd.n2806 72.8958
R3167 vdd.n3088 vdd.n2807 72.8958
R3168 vdd.n3088 vdd.n2808 72.8958
R3169 vdd.n3088 vdd.n2809 72.8958
R3170 vdd.n3088 vdd.n2810 72.8958
R3171 vdd.n3088 vdd.n2811 72.8958
R3172 vdd.n3088 vdd.n2812 72.8958
R3173 vdd.n3088 vdd.n2813 72.8958
R3174 vdd.n3088 vdd.n2814 72.8958
R3175 vdd.n3088 vdd.n2815 72.8958
R3176 vdd.n3088 vdd.n2816 72.8958
R3177 vdd.n3088 vdd.n2817 72.8958
R3178 vdd.n803 vdd.n692 72.8958
R3179 vdd.n3338 vdd.n692 72.8958
R3180 vdd.n797 vdd.n692 72.8958
R3181 vdd.n3345 vdd.n692 72.8958
R3182 vdd.n794 vdd.n692 72.8958
R3183 vdd.n3352 vdd.n692 72.8958
R3184 vdd.n791 vdd.n692 72.8958
R3185 vdd.n3359 vdd.n692 72.8958
R3186 vdd.n3362 vdd.n692 72.8958
R3187 vdd.n3218 vdd.n692 72.8958
R3188 vdd.n3223 vdd.n692 72.8958
R3189 vdd.n3217 vdd.n692 72.8958
R3190 vdd.n3230 vdd.n692 72.8958
R3191 vdd.n3214 vdd.n692 72.8958
R3192 vdd.n3237 vdd.n692 72.8958
R3193 vdd.n3211 vdd.n692 72.8958
R3194 vdd.n3244 vdd.n692 72.8958
R3195 vdd.n2507 vdd.n2506 72.8958
R3196 vdd.n2506 vdd.n1142 72.8958
R3197 vdd.n2506 vdd.n1143 72.8958
R3198 vdd.n2506 vdd.n1144 72.8958
R3199 vdd.n2506 vdd.n1145 72.8958
R3200 vdd.n2506 vdd.n1146 72.8958
R3201 vdd.n2506 vdd.n1147 72.8958
R3202 vdd.n2506 vdd.n1148 72.8958
R3203 vdd.n2506 vdd.n1149 72.8958
R3204 vdd.n2506 vdd.n1150 72.8958
R3205 vdd.n2506 vdd.n1151 72.8958
R3206 vdd.n2506 vdd.n1152 72.8958
R3207 vdd.n2506 vdd.n1153 72.8958
R3208 vdd.n2506 vdd.n1154 72.8958
R3209 vdd.n2506 vdd.n1155 72.8958
R3210 vdd.n2506 vdd.n1156 72.8958
R3211 vdd.n2506 vdd.n1157 72.8958
R3212 vdd.n2784 vdd.n981 72.8958
R3213 vdd.n2784 vdd.n982 72.8958
R3214 vdd.n2784 vdd.n983 72.8958
R3215 vdd.n2784 vdd.n984 72.8958
R3216 vdd.n2784 vdd.n985 72.8958
R3217 vdd.n2784 vdd.n986 72.8958
R3218 vdd.n2784 vdd.n987 72.8958
R3219 vdd.n2784 vdd.n988 72.8958
R3220 vdd.n2784 vdd.n989 72.8958
R3221 vdd.n2784 vdd.n990 72.8958
R3222 vdd.n2784 vdd.n991 72.8958
R3223 vdd.n2784 vdd.n992 72.8958
R3224 vdd.n2784 vdd.n993 72.8958
R3225 vdd.n2784 vdd.n994 72.8958
R3226 vdd.n2784 vdd.n995 72.8958
R3227 vdd.n2784 vdd.n996 72.8958
R3228 vdd.n2784 vdd.n997 72.8958
R3229 vdd.n3089 vdd.n3088 72.8958
R3230 vdd.n3088 vdd.n2785 72.8958
R3231 vdd.n3088 vdd.n2786 72.8958
R3232 vdd.n3088 vdd.n2787 72.8958
R3233 vdd.n3088 vdd.n2788 72.8958
R3234 vdd.n3088 vdd.n2789 72.8958
R3235 vdd.n3088 vdd.n2790 72.8958
R3236 vdd.n3088 vdd.n2791 72.8958
R3237 vdd.n3088 vdd.n2792 72.8958
R3238 vdd.n3088 vdd.n2793 72.8958
R3239 vdd.n3088 vdd.n2794 72.8958
R3240 vdd.n3088 vdd.n2795 72.8958
R3241 vdd.n3088 vdd.n2796 72.8958
R3242 vdd.n3088 vdd.n2797 72.8958
R3243 vdd.n3088 vdd.n2798 72.8958
R3244 vdd.n3088 vdd.n2799 72.8958
R3245 vdd.n3088 vdd.n2800 72.8958
R3246 vdd.n3268 vdd.n692 72.8958
R3247 vdd.n835 vdd.n692 72.8958
R3248 vdd.n3276 vdd.n692 72.8958
R3249 vdd.n830 vdd.n692 72.8958
R3250 vdd.n3283 vdd.n692 72.8958
R3251 vdd.n827 vdd.n692 72.8958
R3252 vdd.n3290 vdd.n692 72.8958
R3253 vdd.n824 vdd.n692 72.8958
R3254 vdd.n3297 vdd.n692 72.8958
R3255 vdd.n3301 vdd.n692 72.8958
R3256 vdd.n821 vdd.n692 72.8958
R3257 vdd.n3308 vdd.n692 72.8958
R3258 vdd.n818 vdd.n692 72.8958
R3259 vdd.n3315 vdd.n692 72.8958
R3260 vdd.n815 vdd.n692 72.8958
R3261 vdd.n3322 vdd.n692 72.8958
R3262 vdd.n3325 vdd.n692 72.8958
R3263 vdd.n2784 vdd.n979 72.8958
R3264 vdd.n2784 vdd.n978 72.8958
R3265 vdd.n2784 vdd.n977 72.8958
R3266 vdd.n2784 vdd.n976 72.8958
R3267 vdd.n2784 vdd.n975 72.8958
R3268 vdd.n2784 vdd.n974 72.8958
R3269 vdd.n2784 vdd.n973 72.8958
R3270 vdd.n2784 vdd.n972 72.8958
R3271 vdd.n2784 vdd.n971 72.8958
R3272 vdd.n2784 vdd.n970 72.8958
R3273 vdd.n2784 vdd.n969 72.8958
R3274 vdd.n2784 vdd.n968 72.8958
R3275 vdd.n2784 vdd.n967 72.8958
R3276 vdd.n2784 vdd.n966 72.8958
R3277 vdd.n2784 vdd.n965 72.8958
R3278 vdd.n2784 vdd.n964 72.8958
R3279 vdd.n2784 vdd.n963 72.8958
R3280 vdd.n2506 vdd.n1158 72.8958
R3281 vdd.n2506 vdd.n1159 72.8958
R3282 vdd.n2506 vdd.n1160 72.8958
R3283 vdd.n2506 vdd.n1161 72.8958
R3284 vdd.n2506 vdd.n1162 72.8958
R3285 vdd.n2506 vdd.n1163 72.8958
R3286 vdd.n2506 vdd.n1164 72.8958
R3287 vdd.n2506 vdd.n1165 72.8958
R3288 vdd.n2506 vdd.n1166 72.8958
R3289 vdd.n2506 vdd.n1167 72.8958
R3290 vdd.n2506 vdd.n1168 72.8958
R3291 vdd.n2506 vdd.n1169 72.8958
R3292 vdd.n2506 vdd.n1170 72.8958
R3293 vdd.n2506 vdd.n1171 72.8958
R3294 vdd.n2506 vdd.n1172 72.8958
R3295 vdd.n2506 vdd.n1173 72.8958
R3296 vdd.n2506 vdd.n1174 72.8958
R3297 vdd.n1874 vdd.n1873 66.2847
R3298 vdd.n1873 vdd.n1649 66.2847
R3299 vdd.n1873 vdd.n1650 66.2847
R3300 vdd.n1873 vdd.n1651 66.2847
R3301 vdd.n1873 vdd.n1652 66.2847
R3302 vdd.n1873 vdd.n1653 66.2847
R3303 vdd.n1873 vdd.n1654 66.2847
R3304 vdd.n1873 vdd.n1655 66.2847
R3305 vdd.n1873 vdd.n1656 66.2847
R3306 vdd.n1873 vdd.n1657 66.2847
R3307 vdd.n1873 vdd.n1658 66.2847
R3308 vdd.n1873 vdd.n1659 66.2847
R3309 vdd.n1873 vdd.n1660 66.2847
R3310 vdd.n1873 vdd.n1661 66.2847
R3311 vdd.n1873 vdd.n1662 66.2847
R3312 vdd.n1873 vdd.n1663 66.2847
R3313 vdd.n1873 vdd.n1664 66.2847
R3314 vdd.n1873 vdd.n1665 66.2847
R3315 vdd.n1873 vdd.n1666 66.2847
R3316 vdd.n1873 vdd.n1667 66.2847
R3317 vdd.n1873 vdd.n1668 66.2847
R3318 vdd.n1873 vdd.n1669 66.2847
R3319 vdd.n1873 vdd.n1670 66.2847
R3320 vdd.n1873 vdd.n1671 66.2847
R3321 vdd.n1873 vdd.n1672 66.2847
R3322 vdd.n1873 vdd.n1673 66.2847
R3323 vdd.n1873 vdd.n1674 66.2847
R3324 vdd.n1873 vdd.n1675 66.2847
R3325 vdd.n1873 vdd.n1676 66.2847
R3326 vdd.n1873 vdd.n1677 66.2847
R3327 vdd.n1873 vdd.n1678 66.2847
R3328 vdd.n1526 vdd.n1141 66.2847
R3329 vdd.n1523 vdd.n1141 66.2847
R3330 vdd.n1519 vdd.n1141 66.2847
R3331 vdd.n2372 vdd.n1141 66.2847
R3332 vdd.n1275 vdd.n1141 66.2847
R3333 vdd.n2379 vdd.n1141 66.2847
R3334 vdd.n1268 vdd.n1141 66.2847
R3335 vdd.n2386 vdd.n1141 66.2847
R3336 vdd.n1261 vdd.n1141 66.2847
R3337 vdd.n2393 vdd.n1141 66.2847
R3338 vdd.n1255 vdd.n1141 66.2847
R3339 vdd.n1250 vdd.n1141 66.2847
R3340 vdd.n2404 vdd.n1141 66.2847
R3341 vdd.n1242 vdd.n1141 66.2847
R3342 vdd.n2411 vdd.n1141 66.2847
R3343 vdd.n1235 vdd.n1141 66.2847
R3344 vdd.n2418 vdd.n1141 66.2847
R3345 vdd.n1228 vdd.n1141 66.2847
R3346 vdd.n2425 vdd.n1141 66.2847
R3347 vdd.n1221 vdd.n1141 66.2847
R3348 vdd.n2432 vdd.n1141 66.2847
R3349 vdd.n1215 vdd.n1141 66.2847
R3350 vdd.n1210 vdd.n1141 66.2847
R3351 vdd.n2443 vdd.n1141 66.2847
R3352 vdd.n1202 vdd.n1141 66.2847
R3353 vdd.n2450 vdd.n1141 66.2847
R3354 vdd.n1195 vdd.n1141 66.2847
R3355 vdd.n2457 vdd.n1141 66.2847
R3356 vdd.n1188 vdd.n1141 66.2847
R3357 vdd.n2464 vdd.n1141 66.2847
R3358 vdd.n2469 vdd.n1141 66.2847
R3359 vdd.n1184 vdd.n1141 66.2847
R3360 vdd.n3495 vdd.n3494 66.2847
R3361 vdd.n3495 vdd.n693 66.2847
R3362 vdd.n3495 vdd.n694 66.2847
R3363 vdd.n3495 vdd.n695 66.2847
R3364 vdd.n3495 vdd.n696 66.2847
R3365 vdd.n3495 vdd.n697 66.2847
R3366 vdd.n3495 vdd.n698 66.2847
R3367 vdd.n3495 vdd.n699 66.2847
R3368 vdd.n3495 vdd.n700 66.2847
R3369 vdd.n3495 vdd.n701 66.2847
R3370 vdd.n3495 vdd.n702 66.2847
R3371 vdd.n3495 vdd.n703 66.2847
R3372 vdd.n3495 vdd.n704 66.2847
R3373 vdd.n3495 vdd.n705 66.2847
R3374 vdd.n3495 vdd.n706 66.2847
R3375 vdd.n3495 vdd.n707 66.2847
R3376 vdd.n3495 vdd.n708 66.2847
R3377 vdd.n3495 vdd.n709 66.2847
R3378 vdd.n3495 vdd.n710 66.2847
R3379 vdd.n3495 vdd.n711 66.2847
R3380 vdd.n3495 vdd.n712 66.2847
R3381 vdd.n3495 vdd.n713 66.2847
R3382 vdd.n3495 vdd.n714 66.2847
R3383 vdd.n3495 vdd.n715 66.2847
R3384 vdd.n3495 vdd.n716 66.2847
R3385 vdd.n3495 vdd.n717 66.2847
R3386 vdd.n3495 vdd.n718 66.2847
R3387 vdd.n3495 vdd.n719 66.2847
R3388 vdd.n3495 vdd.n720 66.2847
R3389 vdd.n3495 vdd.n721 66.2847
R3390 vdd.n3495 vdd.n722 66.2847
R3391 vdd.n3626 vdd.n3625 66.2847
R3392 vdd.n3626 vdd.n424 66.2847
R3393 vdd.n3626 vdd.n423 66.2847
R3394 vdd.n3626 vdd.n422 66.2847
R3395 vdd.n3626 vdd.n421 66.2847
R3396 vdd.n3626 vdd.n420 66.2847
R3397 vdd.n3626 vdd.n419 66.2847
R3398 vdd.n3626 vdd.n418 66.2847
R3399 vdd.n3626 vdd.n417 66.2847
R3400 vdd.n3626 vdd.n416 66.2847
R3401 vdd.n3626 vdd.n415 66.2847
R3402 vdd.n3626 vdd.n414 66.2847
R3403 vdd.n3626 vdd.n413 66.2847
R3404 vdd.n3626 vdd.n412 66.2847
R3405 vdd.n3626 vdd.n411 66.2847
R3406 vdd.n3626 vdd.n410 66.2847
R3407 vdd.n3626 vdd.n409 66.2847
R3408 vdd.n3626 vdd.n408 66.2847
R3409 vdd.n3626 vdd.n407 66.2847
R3410 vdd.n3626 vdd.n406 66.2847
R3411 vdd.n3626 vdd.n405 66.2847
R3412 vdd.n3626 vdd.n404 66.2847
R3413 vdd.n3626 vdd.n403 66.2847
R3414 vdd.n3626 vdd.n402 66.2847
R3415 vdd.n3626 vdd.n401 66.2847
R3416 vdd.n3626 vdd.n400 66.2847
R3417 vdd.n3626 vdd.n399 66.2847
R3418 vdd.n3626 vdd.n398 66.2847
R3419 vdd.n3626 vdd.n397 66.2847
R3420 vdd.n3626 vdd.n396 66.2847
R3421 vdd.n3626 vdd.n395 66.2847
R3422 vdd.n3626 vdd.n394 66.2847
R3423 vdd.n467 vdd.n394 52.4337
R3424 vdd.n473 vdd.n395 52.4337
R3425 vdd.n477 vdd.n396 52.4337
R3426 vdd.n483 vdd.n397 52.4337
R3427 vdd.n487 vdd.n398 52.4337
R3428 vdd.n493 vdd.n399 52.4337
R3429 vdd.n497 vdd.n400 52.4337
R3430 vdd.n503 vdd.n401 52.4337
R3431 vdd.n507 vdd.n402 52.4337
R3432 vdd.n513 vdd.n403 52.4337
R3433 vdd.n517 vdd.n404 52.4337
R3434 vdd.n523 vdd.n405 52.4337
R3435 vdd.n527 vdd.n406 52.4337
R3436 vdd.n533 vdd.n407 52.4337
R3437 vdd.n537 vdd.n408 52.4337
R3438 vdd.n543 vdd.n409 52.4337
R3439 vdd.n547 vdd.n410 52.4337
R3440 vdd.n553 vdd.n411 52.4337
R3441 vdd.n557 vdd.n412 52.4337
R3442 vdd.n563 vdd.n413 52.4337
R3443 vdd.n567 vdd.n414 52.4337
R3444 vdd.n573 vdd.n415 52.4337
R3445 vdd.n577 vdd.n416 52.4337
R3446 vdd.n583 vdd.n417 52.4337
R3447 vdd.n587 vdd.n418 52.4337
R3448 vdd.n593 vdd.n419 52.4337
R3449 vdd.n597 vdd.n420 52.4337
R3450 vdd.n603 vdd.n421 52.4337
R3451 vdd.n607 vdd.n422 52.4337
R3452 vdd.n613 vdd.n423 52.4337
R3453 vdd.n616 vdd.n424 52.4337
R3454 vdd.n3625 vdd.n3624 52.4337
R3455 vdd.n3494 vdd.n3493 52.4337
R3456 vdd.n728 vdd.n693 52.4337
R3457 vdd.n734 vdd.n694 52.4337
R3458 vdd.n3483 vdd.n695 52.4337
R3459 vdd.n3479 vdd.n696 52.4337
R3460 vdd.n3475 vdd.n697 52.4337
R3461 vdd.n3471 vdd.n698 52.4337
R3462 vdd.n3467 vdd.n699 52.4337
R3463 vdd.n3463 vdd.n700 52.4337
R3464 vdd.n3459 vdd.n701 52.4337
R3465 vdd.n3451 vdd.n702 52.4337
R3466 vdd.n3447 vdd.n703 52.4337
R3467 vdd.n3443 vdd.n704 52.4337
R3468 vdd.n3439 vdd.n705 52.4337
R3469 vdd.n3435 vdd.n706 52.4337
R3470 vdd.n3431 vdd.n707 52.4337
R3471 vdd.n3427 vdd.n708 52.4337
R3472 vdd.n3423 vdd.n709 52.4337
R3473 vdd.n3419 vdd.n710 52.4337
R3474 vdd.n3415 vdd.n711 52.4337
R3475 vdd.n3411 vdd.n712 52.4337
R3476 vdd.n3405 vdd.n713 52.4337
R3477 vdd.n3401 vdd.n714 52.4337
R3478 vdd.n3397 vdd.n715 52.4337
R3479 vdd.n3393 vdd.n716 52.4337
R3480 vdd.n3389 vdd.n717 52.4337
R3481 vdd.n3385 vdd.n718 52.4337
R3482 vdd.n3381 vdd.n719 52.4337
R3483 vdd.n3377 vdd.n720 52.4337
R3484 vdd.n3373 vdd.n721 52.4337
R3485 vdd.n3369 vdd.n722 52.4337
R3486 vdd.n2471 vdd.n1184 52.4337
R3487 vdd.n2469 vdd.n2468 52.4337
R3488 vdd.n2464 vdd.n2463 52.4337
R3489 vdd.n2459 vdd.n1188 52.4337
R3490 vdd.n2457 vdd.n2456 52.4337
R3491 vdd.n2452 vdd.n1195 52.4337
R3492 vdd.n2450 vdd.n2449 52.4337
R3493 vdd.n2445 vdd.n1202 52.4337
R3494 vdd.n2443 vdd.n2442 52.4337
R3495 vdd.n1211 vdd.n1210 52.4337
R3496 vdd.n2434 vdd.n1215 52.4337
R3497 vdd.n2432 vdd.n2431 52.4337
R3498 vdd.n2427 vdd.n1221 52.4337
R3499 vdd.n2425 vdd.n2424 52.4337
R3500 vdd.n2420 vdd.n1228 52.4337
R3501 vdd.n2418 vdd.n2417 52.4337
R3502 vdd.n2413 vdd.n1235 52.4337
R3503 vdd.n2411 vdd.n2410 52.4337
R3504 vdd.n2406 vdd.n1242 52.4337
R3505 vdd.n2404 vdd.n2403 52.4337
R3506 vdd.n1251 vdd.n1250 52.4337
R3507 vdd.n2395 vdd.n1255 52.4337
R3508 vdd.n2393 vdd.n2392 52.4337
R3509 vdd.n2388 vdd.n1261 52.4337
R3510 vdd.n2386 vdd.n2385 52.4337
R3511 vdd.n2381 vdd.n1268 52.4337
R3512 vdd.n2379 vdd.n2378 52.4337
R3513 vdd.n2374 vdd.n1275 52.4337
R3514 vdd.n2372 vdd.n2371 52.4337
R3515 vdd.n1520 vdd.n1519 52.4337
R3516 vdd.n1524 vdd.n1523 52.4337
R3517 vdd.n2360 vdd.n1526 52.4337
R3518 vdd.n1875 vdd.n1874 52.4337
R3519 vdd.n1681 vdd.n1649 52.4337
R3520 vdd.n1685 vdd.n1650 52.4337
R3521 vdd.n1687 vdd.n1651 52.4337
R3522 vdd.n1691 vdd.n1652 52.4337
R3523 vdd.n1693 vdd.n1653 52.4337
R3524 vdd.n1697 vdd.n1654 52.4337
R3525 vdd.n1699 vdd.n1655 52.4337
R3526 vdd.n1703 vdd.n1656 52.4337
R3527 vdd.n1705 vdd.n1657 52.4337
R3528 vdd.n1711 vdd.n1658 52.4337
R3529 vdd.n1713 vdd.n1659 52.4337
R3530 vdd.n1717 vdd.n1660 52.4337
R3531 vdd.n1719 vdd.n1661 52.4337
R3532 vdd.n1723 vdd.n1662 52.4337
R3533 vdd.n1725 vdd.n1663 52.4337
R3534 vdd.n1729 vdd.n1664 52.4337
R3535 vdd.n1731 vdd.n1665 52.4337
R3536 vdd.n1735 vdd.n1666 52.4337
R3537 vdd.n1737 vdd.n1667 52.4337
R3538 vdd.n1809 vdd.n1668 52.4337
R3539 vdd.n1742 vdd.n1669 52.4337
R3540 vdd.n1746 vdd.n1670 52.4337
R3541 vdd.n1748 vdd.n1671 52.4337
R3542 vdd.n1752 vdd.n1672 52.4337
R3543 vdd.n1754 vdd.n1673 52.4337
R3544 vdd.n1758 vdd.n1674 52.4337
R3545 vdd.n1760 vdd.n1675 52.4337
R3546 vdd.n1764 vdd.n1676 52.4337
R3547 vdd.n1766 vdd.n1677 52.4337
R3548 vdd.n1770 vdd.n1678 52.4337
R3549 vdd.n1874 vdd.n1648 52.4337
R3550 vdd.n1684 vdd.n1649 52.4337
R3551 vdd.n1686 vdd.n1650 52.4337
R3552 vdd.n1690 vdd.n1651 52.4337
R3553 vdd.n1692 vdd.n1652 52.4337
R3554 vdd.n1696 vdd.n1653 52.4337
R3555 vdd.n1698 vdd.n1654 52.4337
R3556 vdd.n1702 vdd.n1655 52.4337
R3557 vdd.n1704 vdd.n1656 52.4337
R3558 vdd.n1710 vdd.n1657 52.4337
R3559 vdd.n1712 vdd.n1658 52.4337
R3560 vdd.n1716 vdd.n1659 52.4337
R3561 vdd.n1718 vdd.n1660 52.4337
R3562 vdd.n1722 vdd.n1661 52.4337
R3563 vdd.n1724 vdd.n1662 52.4337
R3564 vdd.n1728 vdd.n1663 52.4337
R3565 vdd.n1730 vdd.n1664 52.4337
R3566 vdd.n1734 vdd.n1665 52.4337
R3567 vdd.n1736 vdd.n1666 52.4337
R3568 vdd.n1740 vdd.n1667 52.4337
R3569 vdd.n1741 vdd.n1668 52.4337
R3570 vdd.n1745 vdd.n1669 52.4337
R3571 vdd.n1747 vdd.n1670 52.4337
R3572 vdd.n1751 vdd.n1671 52.4337
R3573 vdd.n1753 vdd.n1672 52.4337
R3574 vdd.n1757 vdd.n1673 52.4337
R3575 vdd.n1759 vdd.n1674 52.4337
R3576 vdd.n1763 vdd.n1675 52.4337
R3577 vdd.n1765 vdd.n1676 52.4337
R3578 vdd.n1769 vdd.n1677 52.4337
R3579 vdd.n1771 vdd.n1678 52.4337
R3580 vdd.n1526 vdd.n1525 52.4337
R3581 vdd.n1523 vdd.n1522 52.4337
R3582 vdd.n1519 vdd.n1276 52.4337
R3583 vdd.n2373 vdd.n2372 52.4337
R3584 vdd.n1275 vdd.n1269 52.4337
R3585 vdd.n2380 vdd.n2379 52.4337
R3586 vdd.n1268 vdd.n1262 52.4337
R3587 vdd.n2387 vdd.n2386 52.4337
R3588 vdd.n1261 vdd.n1256 52.4337
R3589 vdd.n2394 vdd.n2393 52.4337
R3590 vdd.n1255 vdd.n1254 52.4337
R3591 vdd.n1250 vdd.n1243 52.4337
R3592 vdd.n2405 vdd.n2404 52.4337
R3593 vdd.n1242 vdd.n1236 52.4337
R3594 vdd.n2412 vdd.n2411 52.4337
R3595 vdd.n1235 vdd.n1229 52.4337
R3596 vdd.n2419 vdd.n2418 52.4337
R3597 vdd.n1228 vdd.n1222 52.4337
R3598 vdd.n2426 vdd.n2425 52.4337
R3599 vdd.n1221 vdd.n1216 52.4337
R3600 vdd.n2433 vdd.n2432 52.4337
R3601 vdd.n1215 vdd.n1214 52.4337
R3602 vdd.n1210 vdd.n1203 52.4337
R3603 vdd.n2444 vdd.n2443 52.4337
R3604 vdd.n1202 vdd.n1196 52.4337
R3605 vdd.n2451 vdd.n2450 52.4337
R3606 vdd.n1195 vdd.n1189 52.4337
R3607 vdd.n2458 vdd.n2457 52.4337
R3608 vdd.n1188 vdd.n1185 52.4337
R3609 vdd.n2465 vdd.n2464 52.4337
R3610 vdd.n2470 vdd.n2469 52.4337
R3611 vdd.n1530 vdd.n1184 52.4337
R3612 vdd.n3494 vdd.n725 52.4337
R3613 vdd.n733 vdd.n693 52.4337
R3614 vdd.n3484 vdd.n694 52.4337
R3615 vdd.n3480 vdd.n695 52.4337
R3616 vdd.n3476 vdd.n696 52.4337
R3617 vdd.n3472 vdd.n697 52.4337
R3618 vdd.n3468 vdd.n698 52.4337
R3619 vdd.n3464 vdd.n699 52.4337
R3620 vdd.n3460 vdd.n700 52.4337
R3621 vdd.n3450 vdd.n701 52.4337
R3622 vdd.n3448 vdd.n702 52.4337
R3623 vdd.n3444 vdd.n703 52.4337
R3624 vdd.n3440 vdd.n704 52.4337
R3625 vdd.n3436 vdd.n705 52.4337
R3626 vdd.n3432 vdd.n706 52.4337
R3627 vdd.n3428 vdd.n707 52.4337
R3628 vdd.n3424 vdd.n708 52.4337
R3629 vdd.n3420 vdd.n709 52.4337
R3630 vdd.n3416 vdd.n710 52.4337
R3631 vdd.n3412 vdd.n711 52.4337
R3632 vdd.n3404 vdd.n712 52.4337
R3633 vdd.n3402 vdd.n713 52.4337
R3634 vdd.n3398 vdd.n714 52.4337
R3635 vdd.n3394 vdd.n715 52.4337
R3636 vdd.n3390 vdd.n716 52.4337
R3637 vdd.n3386 vdd.n717 52.4337
R3638 vdd.n3382 vdd.n718 52.4337
R3639 vdd.n3378 vdd.n719 52.4337
R3640 vdd.n3374 vdd.n720 52.4337
R3641 vdd.n3370 vdd.n721 52.4337
R3642 vdd.n722 vdd.n691 52.4337
R3643 vdd.n3625 vdd.n425 52.4337
R3644 vdd.n614 vdd.n424 52.4337
R3645 vdd.n608 vdd.n423 52.4337
R3646 vdd.n604 vdd.n422 52.4337
R3647 vdd.n598 vdd.n421 52.4337
R3648 vdd.n594 vdd.n420 52.4337
R3649 vdd.n588 vdd.n419 52.4337
R3650 vdd.n584 vdd.n418 52.4337
R3651 vdd.n578 vdd.n417 52.4337
R3652 vdd.n574 vdd.n416 52.4337
R3653 vdd.n568 vdd.n415 52.4337
R3654 vdd.n564 vdd.n414 52.4337
R3655 vdd.n558 vdd.n413 52.4337
R3656 vdd.n554 vdd.n412 52.4337
R3657 vdd.n548 vdd.n411 52.4337
R3658 vdd.n544 vdd.n410 52.4337
R3659 vdd.n538 vdd.n409 52.4337
R3660 vdd.n534 vdd.n408 52.4337
R3661 vdd.n528 vdd.n407 52.4337
R3662 vdd.n524 vdd.n406 52.4337
R3663 vdd.n518 vdd.n405 52.4337
R3664 vdd.n514 vdd.n404 52.4337
R3665 vdd.n508 vdd.n403 52.4337
R3666 vdd.n504 vdd.n402 52.4337
R3667 vdd.n498 vdd.n401 52.4337
R3668 vdd.n494 vdd.n400 52.4337
R3669 vdd.n488 vdd.n399 52.4337
R3670 vdd.n484 vdd.n398 52.4337
R3671 vdd.n478 vdd.n397 52.4337
R3672 vdd.n474 vdd.n396 52.4337
R3673 vdd.n468 vdd.n395 52.4337
R3674 vdd.n394 vdd.n392 52.4337
R3675 vdd.t156 vdd.t169 51.4683
R3676 vdd.n274 vdd.n272 42.0461
R3677 vdd.n172 vdd.n170 42.0461
R3678 vdd.n71 vdd.n69 42.0461
R3679 vdd.n2207 vdd.n2205 42.0461
R3680 vdd.n2105 vdd.n2103 42.0461
R3681 vdd.n2004 vdd.n2002 42.0461
R3682 vdd.n332 vdd.n331 41.6884
R3683 vdd.n230 vdd.n229 41.6884
R3684 vdd.n129 vdd.n128 41.6884
R3685 vdd.n2265 vdd.n2264 41.6884
R3686 vdd.n2163 vdd.n2162 41.6884
R3687 vdd.n2062 vdd.n2061 41.6884
R3688 vdd.n1774 vdd.n1773 41.1157
R3689 vdd.n1812 vdd.n1811 41.1157
R3690 vdd.n1708 vdd.n1707 41.1157
R3691 vdd.n428 vdd.n427 41.1157
R3692 vdd.n566 vdd.n441 41.1157
R3693 vdd.n454 vdd.n453 41.1157
R3694 vdd.n3325 vdd.n3324 39.2114
R3695 vdd.n3322 vdd.n3321 39.2114
R3696 vdd.n3317 vdd.n815 39.2114
R3697 vdd.n3315 vdd.n3314 39.2114
R3698 vdd.n3310 vdd.n818 39.2114
R3699 vdd.n3308 vdd.n3307 39.2114
R3700 vdd.n3303 vdd.n821 39.2114
R3701 vdd.n3301 vdd.n3300 39.2114
R3702 vdd.n3297 vdd.n3296 39.2114
R3703 vdd.n3292 vdd.n824 39.2114
R3704 vdd.n3290 vdd.n3289 39.2114
R3705 vdd.n3285 vdd.n827 39.2114
R3706 vdd.n3283 vdd.n3282 39.2114
R3707 vdd.n3278 vdd.n830 39.2114
R3708 vdd.n3276 vdd.n3275 39.2114
R3709 vdd.n3270 vdd.n835 39.2114
R3710 vdd.n3268 vdd.n3267 39.2114
R3711 vdd.n3090 vdd.n3089 39.2114
R3712 vdd.n2819 vdd.n2785 39.2114
R3713 vdd.n3082 vdd.n2786 39.2114
R3714 vdd.n3078 vdd.n2787 39.2114
R3715 vdd.n3074 vdd.n2788 39.2114
R3716 vdd.n3070 vdd.n2789 39.2114
R3717 vdd.n3066 vdd.n2790 39.2114
R3718 vdd.n3062 vdd.n2791 39.2114
R3719 vdd.n3058 vdd.n2792 39.2114
R3720 vdd.n3054 vdd.n2793 39.2114
R3721 vdd.n3050 vdd.n2794 39.2114
R3722 vdd.n3046 vdd.n2795 39.2114
R3723 vdd.n3042 vdd.n2796 39.2114
R3724 vdd.n3038 vdd.n2797 39.2114
R3725 vdd.n3034 vdd.n2798 39.2114
R3726 vdd.n3030 vdd.n2799 39.2114
R3727 vdd.n3025 vdd.n2800 39.2114
R3728 vdd.n2779 vdd.n997 39.2114
R3729 vdd.n2775 vdd.n996 39.2114
R3730 vdd.n2771 vdd.n995 39.2114
R3731 vdd.n2767 vdd.n994 39.2114
R3732 vdd.n2763 vdd.n993 39.2114
R3733 vdd.n2759 vdd.n992 39.2114
R3734 vdd.n2755 vdd.n991 39.2114
R3735 vdd.n2751 vdd.n990 39.2114
R3736 vdd.n2747 vdd.n989 39.2114
R3737 vdd.n2743 vdd.n988 39.2114
R3738 vdd.n2739 vdd.n987 39.2114
R3739 vdd.n2735 vdd.n986 39.2114
R3740 vdd.n2731 vdd.n985 39.2114
R3741 vdd.n2727 vdd.n984 39.2114
R3742 vdd.n2723 vdd.n983 39.2114
R3743 vdd.n2718 vdd.n982 39.2114
R3744 vdd.n2714 vdd.n981 39.2114
R3745 vdd.n2508 vdd.n2507 39.2114
R3746 vdd.n1176 vdd.n1142 39.2114
R3747 vdd.n2500 vdd.n1143 39.2114
R3748 vdd.n2496 vdd.n1144 39.2114
R3749 vdd.n2492 vdd.n1145 39.2114
R3750 vdd.n2488 vdd.n1146 39.2114
R3751 vdd.n2484 vdd.n1147 39.2114
R3752 vdd.n2480 vdd.n1148 39.2114
R3753 vdd.n2476 vdd.n1149 39.2114
R3754 vdd.n1322 vdd.n1150 39.2114
R3755 vdd.n1326 vdd.n1151 39.2114
R3756 vdd.n1330 vdd.n1152 39.2114
R3757 vdd.n1334 vdd.n1153 39.2114
R3758 vdd.n1338 vdd.n1154 39.2114
R3759 vdd.n1342 vdd.n1155 39.2114
R3760 vdd.n1346 vdd.n1156 39.2114
R3761 vdd.n1351 vdd.n1157 39.2114
R3762 vdd.n3244 vdd.n3243 39.2114
R3763 vdd.n3239 vdd.n3211 39.2114
R3764 vdd.n3237 vdd.n3236 39.2114
R3765 vdd.n3232 vdd.n3214 39.2114
R3766 vdd.n3230 vdd.n3229 39.2114
R3767 vdd.n3225 vdd.n3217 39.2114
R3768 vdd.n3223 vdd.n3222 39.2114
R3769 vdd.n3218 vdd.n787 39.2114
R3770 vdd.n3362 vdd.n3361 39.2114
R3771 vdd.n3359 vdd.n3358 39.2114
R3772 vdd.n3354 vdd.n791 39.2114
R3773 vdd.n3352 vdd.n3351 39.2114
R3774 vdd.n3347 vdd.n794 39.2114
R3775 vdd.n3345 vdd.n3344 39.2114
R3776 vdd.n3340 vdd.n797 39.2114
R3777 vdd.n3338 vdd.n3337 39.2114
R3778 vdd.n3333 vdd.n803 39.2114
R3779 vdd.n2826 vdd.n2801 39.2114
R3780 vdd.n2830 vdd.n2802 39.2114
R3781 vdd.n2834 vdd.n2803 39.2114
R3782 vdd.n2838 vdd.n2804 39.2114
R3783 vdd.n2842 vdd.n2805 39.2114
R3784 vdd.n2846 vdd.n2806 39.2114
R3785 vdd.n2850 vdd.n2807 39.2114
R3786 vdd.n2854 vdd.n2808 39.2114
R3787 vdd.n2858 vdd.n2809 39.2114
R3788 vdd.n2862 vdd.n2810 39.2114
R3789 vdd.n2866 vdd.n2811 39.2114
R3790 vdd.n2870 vdd.n2812 39.2114
R3791 vdd.n2874 vdd.n2813 39.2114
R3792 vdd.n2878 vdd.n2814 39.2114
R3793 vdd.n2882 vdd.n2815 39.2114
R3794 vdd.n2886 vdd.n2816 39.2114
R3795 vdd.n2890 vdd.n2817 39.2114
R3796 vdd.n2829 vdd.n2801 39.2114
R3797 vdd.n2833 vdd.n2802 39.2114
R3798 vdd.n2837 vdd.n2803 39.2114
R3799 vdd.n2841 vdd.n2804 39.2114
R3800 vdd.n2845 vdd.n2805 39.2114
R3801 vdd.n2849 vdd.n2806 39.2114
R3802 vdd.n2853 vdd.n2807 39.2114
R3803 vdd.n2857 vdd.n2808 39.2114
R3804 vdd.n2861 vdd.n2809 39.2114
R3805 vdd.n2865 vdd.n2810 39.2114
R3806 vdd.n2869 vdd.n2811 39.2114
R3807 vdd.n2873 vdd.n2812 39.2114
R3808 vdd.n2877 vdd.n2813 39.2114
R3809 vdd.n2881 vdd.n2814 39.2114
R3810 vdd.n2885 vdd.n2815 39.2114
R3811 vdd.n2889 vdd.n2816 39.2114
R3812 vdd.n2892 vdd.n2817 39.2114
R3813 vdd.n803 vdd.n798 39.2114
R3814 vdd.n3339 vdd.n3338 39.2114
R3815 vdd.n797 vdd.n795 39.2114
R3816 vdd.n3346 vdd.n3345 39.2114
R3817 vdd.n794 vdd.n792 39.2114
R3818 vdd.n3353 vdd.n3352 39.2114
R3819 vdd.n791 vdd.n789 39.2114
R3820 vdd.n3360 vdd.n3359 39.2114
R3821 vdd.n3363 vdd.n3362 39.2114
R3822 vdd.n3219 vdd.n3218 39.2114
R3823 vdd.n3224 vdd.n3223 39.2114
R3824 vdd.n3217 vdd.n3215 39.2114
R3825 vdd.n3231 vdd.n3230 39.2114
R3826 vdd.n3214 vdd.n3212 39.2114
R3827 vdd.n3238 vdd.n3237 39.2114
R3828 vdd.n3211 vdd.n3209 39.2114
R3829 vdd.n3245 vdd.n3244 39.2114
R3830 vdd.n2507 vdd.n1140 39.2114
R3831 vdd.n2501 vdd.n1142 39.2114
R3832 vdd.n2497 vdd.n1143 39.2114
R3833 vdd.n2493 vdd.n1144 39.2114
R3834 vdd.n2489 vdd.n1145 39.2114
R3835 vdd.n2485 vdd.n1146 39.2114
R3836 vdd.n2481 vdd.n1147 39.2114
R3837 vdd.n2477 vdd.n1148 39.2114
R3838 vdd.n1321 vdd.n1149 39.2114
R3839 vdd.n1325 vdd.n1150 39.2114
R3840 vdd.n1329 vdd.n1151 39.2114
R3841 vdd.n1333 vdd.n1152 39.2114
R3842 vdd.n1337 vdd.n1153 39.2114
R3843 vdd.n1341 vdd.n1154 39.2114
R3844 vdd.n1345 vdd.n1155 39.2114
R3845 vdd.n1350 vdd.n1156 39.2114
R3846 vdd.n1354 vdd.n1157 39.2114
R3847 vdd.n2717 vdd.n981 39.2114
R3848 vdd.n2722 vdd.n982 39.2114
R3849 vdd.n2726 vdd.n983 39.2114
R3850 vdd.n2730 vdd.n984 39.2114
R3851 vdd.n2734 vdd.n985 39.2114
R3852 vdd.n2738 vdd.n986 39.2114
R3853 vdd.n2742 vdd.n987 39.2114
R3854 vdd.n2746 vdd.n988 39.2114
R3855 vdd.n2750 vdd.n989 39.2114
R3856 vdd.n2754 vdd.n990 39.2114
R3857 vdd.n2758 vdd.n991 39.2114
R3858 vdd.n2762 vdd.n992 39.2114
R3859 vdd.n2766 vdd.n993 39.2114
R3860 vdd.n2770 vdd.n994 39.2114
R3861 vdd.n2774 vdd.n995 39.2114
R3862 vdd.n2778 vdd.n996 39.2114
R3863 vdd.n999 vdd.n997 39.2114
R3864 vdd.n3089 vdd.n962 39.2114
R3865 vdd.n3083 vdd.n2785 39.2114
R3866 vdd.n3079 vdd.n2786 39.2114
R3867 vdd.n3075 vdd.n2787 39.2114
R3868 vdd.n3071 vdd.n2788 39.2114
R3869 vdd.n3067 vdd.n2789 39.2114
R3870 vdd.n3063 vdd.n2790 39.2114
R3871 vdd.n3059 vdd.n2791 39.2114
R3872 vdd.n3055 vdd.n2792 39.2114
R3873 vdd.n3051 vdd.n2793 39.2114
R3874 vdd.n3047 vdd.n2794 39.2114
R3875 vdd.n3043 vdd.n2795 39.2114
R3876 vdd.n3039 vdd.n2796 39.2114
R3877 vdd.n3035 vdd.n2797 39.2114
R3878 vdd.n3031 vdd.n2798 39.2114
R3879 vdd.n3026 vdd.n2799 39.2114
R3880 vdd.n3022 vdd.n2800 39.2114
R3881 vdd.n3269 vdd.n3268 39.2114
R3882 vdd.n835 vdd.n831 39.2114
R3883 vdd.n3277 vdd.n3276 39.2114
R3884 vdd.n830 vdd.n828 39.2114
R3885 vdd.n3284 vdd.n3283 39.2114
R3886 vdd.n827 vdd.n825 39.2114
R3887 vdd.n3291 vdd.n3290 39.2114
R3888 vdd.n824 vdd.n822 39.2114
R3889 vdd.n3298 vdd.n3297 39.2114
R3890 vdd.n3302 vdd.n3301 39.2114
R3891 vdd.n821 vdd.n819 39.2114
R3892 vdd.n3309 vdd.n3308 39.2114
R3893 vdd.n818 vdd.n816 39.2114
R3894 vdd.n3316 vdd.n3315 39.2114
R3895 vdd.n815 vdd.n813 39.2114
R3896 vdd.n3323 vdd.n3322 39.2114
R3897 vdd.n3326 vdd.n3325 39.2114
R3898 vdd.n1008 vdd.n963 39.2114
R3899 vdd.n2706 vdd.n964 39.2114
R3900 vdd.n2702 vdd.n965 39.2114
R3901 vdd.n2698 vdd.n966 39.2114
R3902 vdd.n2694 vdd.n967 39.2114
R3903 vdd.n2690 vdd.n968 39.2114
R3904 vdd.n2686 vdd.n969 39.2114
R3905 vdd.n2682 vdd.n970 39.2114
R3906 vdd.n2678 vdd.n971 39.2114
R3907 vdd.n2674 vdd.n972 39.2114
R3908 vdd.n2670 vdd.n973 39.2114
R3909 vdd.n2666 vdd.n974 39.2114
R3910 vdd.n2662 vdd.n975 39.2114
R3911 vdd.n2658 vdd.n976 39.2114
R3912 vdd.n2654 vdd.n977 39.2114
R3913 vdd.n2650 vdd.n978 39.2114
R3914 vdd.n2646 vdd.n979 39.2114
R3915 vdd.n1280 vdd.n1158 39.2114
R3916 vdd.n1284 vdd.n1159 39.2114
R3917 vdd.n1288 vdd.n1160 39.2114
R3918 vdd.n1292 vdd.n1161 39.2114
R3919 vdd.n1296 vdd.n1162 39.2114
R3920 vdd.n1300 vdd.n1163 39.2114
R3921 vdd.n1304 vdd.n1164 39.2114
R3922 vdd.n1308 vdd.n1165 39.2114
R3923 vdd.n1312 vdd.n1166 39.2114
R3924 vdd.n1513 vdd.n1167 39.2114
R3925 vdd.n1510 vdd.n1168 39.2114
R3926 vdd.n1506 vdd.n1169 39.2114
R3927 vdd.n1502 vdd.n1170 39.2114
R3928 vdd.n1498 vdd.n1171 39.2114
R3929 vdd.n1494 vdd.n1172 39.2114
R3930 vdd.n1490 vdd.n1173 39.2114
R3931 vdd.n1486 vdd.n1174 39.2114
R3932 vdd.n2643 vdd.n979 39.2114
R3933 vdd.n2647 vdd.n978 39.2114
R3934 vdd.n2651 vdd.n977 39.2114
R3935 vdd.n2655 vdd.n976 39.2114
R3936 vdd.n2659 vdd.n975 39.2114
R3937 vdd.n2663 vdd.n974 39.2114
R3938 vdd.n2667 vdd.n973 39.2114
R3939 vdd.n2671 vdd.n972 39.2114
R3940 vdd.n2675 vdd.n971 39.2114
R3941 vdd.n2679 vdd.n970 39.2114
R3942 vdd.n2683 vdd.n969 39.2114
R3943 vdd.n2687 vdd.n968 39.2114
R3944 vdd.n2691 vdd.n967 39.2114
R3945 vdd.n2695 vdd.n966 39.2114
R3946 vdd.n2699 vdd.n965 39.2114
R3947 vdd.n2703 vdd.n964 39.2114
R3948 vdd.n2707 vdd.n963 39.2114
R3949 vdd.n1283 vdd.n1158 39.2114
R3950 vdd.n1287 vdd.n1159 39.2114
R3951 vdd.n1291 vdd.n1160 39.2114
R3952 vdd.n1295 vdd.n1161 39.2114
R3953 vdd.n1299 vdd.n1162 39.2114
R3954 vdd.n1303 vdd.n1163 39.2114
R3955 vdd.n1307 vdd.n1164 39.2114
R3956 vdd.n1311 vdd.n1165 39.2114
R3957 vdd.n1314 vdd.n1166 39.2114
R3958 vdd.n1511 vdd.n1167 39.2114
R3959 vdd.n1507 vdd.n1168 39.2114
R3960 vdd.n1503 vdd.n1169 39.2114
R3961 vdd.n1499 vdd.n1170 39.2114
R3962 vdd.n1495 vdd.n1171 39.2114
R3963 vdd.n1491 vdd.n1172 39.2114
R3964 vdd.n1487 vdd.n1173 39.2114
R3965 vdd.n1483 vdd.n1174 39.2114
R3966 vdd.n2364 vdd.n2363 37.2369
R3967 vdd.n2400 vdd.n1249 37.2369
R3968 vdd.n2439 vdd.n1209 37.2369
R3969 vdd.n3410 vdd.n769 37.2369
R3970 vdd.n3458 vdd.n3457 37.2369
R3971 vdd.n690 vdd.n689 37.2369
R3972 vdd.n1317 vdd.n1316 30.449
R3973 vdd.n1012 vdd.n1011 30.449
R3974 vdd.n1348 vdd.n1320 30.449
R3975 vdd.n2720 vdd.n1002 30.449
R3976 vdd.n2825 vdd.n2824 30.449
R3977 vdd.n3272 vdd.n833 30.449
R3978 vdd.n3028 vdd.n2821 30.449
R3979 vdd.n801 vdd.n800 30.449
R3980 vdd.n2510 vdd.n2509 29.8151
R3981 vdd.n2782 vdd.n1000 29.8151
R3982 vdd.n2715 vdd.n1003 29.8151
R3983 vdd.n1356 vdd.n1353 29.8151
R3984 vdd.n3023 vdd.n3020 29.8151
R3985 vdd.n3266 vdd.n3265 29.8151
R3986 vdd.n3092 vdd.n3091 29.8151
R3987 vdd.n3329 vdd.n3328 29.8151
R3988 vdd.n3248 vdd.n3247 29.8151
R3989 vdd.n3334 vdd.n802 29.8151
R3990 vdd.n2896 vdd.n2894 29.8151
R3991 vdd.n2827 vdd.n955 29.8151
R3992 vdd.n1281 vdd.n1132 29.8151
R3993 vdd.n2710 vdd.n2709 29.8151
R3994 vdd.n2642 vdd.n2641 29.8151
R3995 vdd.n1482 vdd.n1481 29.8151
R3996 vdd.n1873 vdd.n1680 22.2201
R3997 vdd.n2358 vdd.n1141 22.2201
R3998 vdd.n3495 vdd.n723 22.2201
R3999 vdd.n3627 vdd.n3626 22.2201
R4000 vdd.n1884 vdd.n1642 19.3944
R4001 vdd.n1884 vdd.n1640 19.3944
R4002 vdd.n1888 vdd.n1640 19.3944
R4003 vdd.n1888 vdd.n1630 19.3944
R4004 vdd.n1901 vdd.n1630 19.3944
R4005 vdd.n1901 vdd.n1628 19.3944
R4006 vdd.n1905 vdd.n1628 19.3944
R4007 vdd.n1905 vdd.n1620 19.3944
R4008 vdd.n1918 vdd.n1620 19.3944
R4009 vdd.n1918 vdd.n1618 19.3944
R4010 vdd.n1922 vdd.n1618 19.3944
R4011 vdd.n1922 vdd.n1607 19.3944
R4012 vdd.n1934 vdd.n1607 19.3944
R4013 vdd.n1934 vdd.n1605 19.3944
R4014 vdd.n1938 vdd.n1605 19.3944
R4015 vdd.n1938 vdd.n1596 19.3944
R4016 vdd.n1951 vdd.n1596 19.3944
R4017 vdd.n1951 vdd.n1594 19.3944
R4018 vdd.n1955 vdd.n1594 19.3944
R4019 vdd.n1955 vdd.n1585 19.3944
R4020 vdd.n2274 vdd.n1585 19.3944
R4021 vdd.n2274 vdd.n1583 19.3944
R4022 vdd.n2278 vdd.n1583 19.3944
R4023 vdd.n2278 vdd.n1573 19.3944
R4024 vdd.n2291 vdd.n1573 19.3944
R4025 vdd.n2291 vdd.n1571 19.3944
R4026 vdd.n2295 vdd.n1571 19.3944
R4027 vdd.n2295 vdd.n1563 19.3944
R4028 vdd.n2308 vdd.n1563 19.3944
R4029 vdd.n2308 vdd.n1561 19.3944
R4030 vdd.n2312 vdd.n1561 19.3944
R4031 vdd.n2312 vdd.n1550 19.3944
R4032 vdd.n2324 vdd.n1550 19.3944
R4033 vdd.n2324 vdd.n1548 19.3944
R4034 vdd.n2328 vdd.n1548 19.3944
R4035 vdd.n2328 vdd.n1540 19.3944
R4036 vdd.n2341 vdd.n1540 19.3944
R4037 vdd.n2341 vdd.n1537 19.3944
R4038 vdd.n2347 vdd.n1537 19.3944
R4039 vdd.n2347 vdd.n1538 19.3944
R4040 vdd.n1538 vdd.n1528 19.3944
R4041 vdd.n1808 vdd.n1743 19.3944
R4042 vdd.n1804 vdd.n1743 19.3944
R4043 vdd.n1804 vdd.n1803 19.3944
R4044 vdd.n1803 vdd.n1802 19.3944
R4045 vdd.n1802 vdd.n1749 19.3944
R4046 vdd.n1798 vdd.n1749 19.3944
R4047 vdd.n1798 vdd.n1797 19.3944
R4048 vdd.n1797 vdd.n1796 19.3944
R4049 vdd.n1796 vdd.n1755 19.3944
R4050 vdd.n1792 vdd.n1755 19.3944
R4051 vdd.n1792 vdd.n1791 19.3944
R4052 vdd.n1791 vdd.n1790 19.3944
R4053 vdd.n1790 vdd.n1761 19.3944
R4054 vdd.n1786 vdd.n1761 19.3944
R4055 vdd.n1786 vdd.n1785 19.3944
R4056 vdd.n1785 vdd.n1784 19.3944
R4057 vdd.n1784 vdd.n1767 19.3944
R4058 vdd.n1780 vdd.n1767 19.3944
R4059 vdd.n1780 vdd.n1779 19.3944
R4060 vdd.n1779 vdd.n1778 19.3944
R4061 vdd.n1843 vdd.n1842 19.3944
R4062 vdd.n1842 vdd.n1841 19.3944
R4063 vdd.n1841 vdd.n1714 19.3944
R4064 vdd.n1837 vdd.n1714 19.3944
R4065 vdd.n1837 vdd.n1836 19.3944
R4066 vdd.n1836 vdd.n1835 19.3944
R4067 vdd.n1835 vdd.n1720 19.3944
R4068 vdd.n1831 vdd.n1720 19.3944
R4069 vdd.n1831 vdd.n1830 19.3944
R4070 vdd.n1830 vdd.n1829 19.3944
R4071 vdd.n1829 vdd.n1726 19.3944
R4072 vdd.n1825 vdd.n1726 19.3944
R4073 vdd.n1825 vdd.n1824 19.3944
R4074 vdd.n1824 vdd.n1823 19.3944
R4075 vdd.n1823 vdd.n1732 19.3944
R4076 vdd.n1819 vdd.n1732 19.3944
R4077 vdd.n1819 vdd.n1818 19.3944
R4078 vdd.n1818 vdd.n1817 19.3944
R4079 vdd.n1817 vdd.n1738 19.3944
R4080 vdd.n1813 vdd.n1738 19.3944
R4081 vdd.n1876 vdd.n1647 19.3944
R4082 vdd.n1871 vdd.n1647 19.3944
R4083 vdd.n1871 vdd.n1682 19.3944
R4084 vdd.n1867 vdd.n1682 19.3944
R4085 vdd.n1867 vdd.n1866 19.3944
R4086 vdd.n1866 vdd.n1865 19.3944
R4087 vdd.n1865 vdd.n1688 19.3944
R4088 vdd.n1861 vdd.n1688 19.3944
R4089 vdd.n1861 vdd.n1860 19.3944
R4090 vdd.n1860 vdd.n1859 19.3944
R4091 vdd.n1859 vdd.n1694 19.3944
R4092 vdd.n1855 vdd.n1694 19.3944
R4093 vdd.n1855 vdd.n1854 19.3944
R4094 vdd.n1854 vdd.n1853 19.3944
R4095 vdd.n1853 vdd.n1700 19.3944
R4096 vdd.n1849 vdd.n1700 19.3944
R4097 vdd.n1849 vdd.n1848 19.3944
R4098 vdd.n1848 vdd.n1847 19.3944
R4099 vdd.n2396 vdd.n1247 19.3944
R4100 vdd.n2396 vdd.n1253 19.3944
R4101 vdd.n2391 vdd.n1253 19.3944
R4102 vdd.n2391 vdd.n2390 19.3944
R4103 vdd.n2390 vdd.n2389 19.3944
R4104 vdd.n2389 vdd.n1260 19.3944
R4105 vdd.n2384 vdd.n1260 19.3944
R4106 vdd.n2384 vdd.n2383 19.3944
R4107 vdd.n2383 vdd.n2382 19.3944
R4108 vdd.n2382 vdd.n1267 19.3944
R4109 vdd.n2377 vdd.n1267 19.3944
R4110 vdd.n2377 vdd.n2376 19.3944
R4111 vdd.n2376 vdd.n2375 19.3944
R4112 vdd.n2375 vdd.n1274 19.3944
R4113 vdd.n2370 vdd.n1274 19.3944
R4114 vdd.n2370 vdd.n2369 19.3944
R4115 vdd.n1521 vdd.n1279 19.3944
R4116 vdd.n2365 vdd.n1518 19.3944
R4117 vdd.n2435 vdd.n1207 19.3944
R4118 vdd.n2435 vdd.n1213 19.3944
R4119 vdd.n2430 vdd.n1213 19.3944
R4120 vdd.n2430 vdd.n2429 19.3944
R4121 vdd.n2429 vdd.n2428 19.3944
R4122 vdd.n2428 vdd.n1220 19.3944
R4123 vdd.n2423 vdd.n1220 19.3944
R4124 vdd.n2423 vdd.n2422 19.3944
R4125 vdd.n2422 vdd.n2421 19.3944
R4126 vdd.n2421 vdd.n1227 19.3944
R4127 vdd.n2416 vdd.n1227 19.3944
R4128 vdd.n2416 vdd.n2415 19.3944
R4129 vdd.n2415 vdd.n2414 19.3944
R4130 vdd.n2414 vdd.n1234 19.3944
R4131 vdd.n2409 vdd.n1234 19.3944
R4132 vdd.n2409 vdd.n2408 19.3944
R4133 vdd.n2408 vdd.n2407 19.3944
R4134 vdd.n2407 vdd.n1241 19.3944
R4135 vdd.n2402 vdd.n1241 19.3944
R4136 vdd.n2402 vdd.n2401 19.3944
R4137 vdd.n2472 vdd.n1182 19.3944
R4138 vdd.n2472 vdd.n1183 19.3944
R4139 vdd.n2467 vdd.n2466 19.3944
R4140 vdd.n2462 vdd.n2461 19.3944
R4141 vdd.n2461 vdd.n2460 19.3944
R4142 vdd.n2460 vdd.n1187 19.3944
R4143 vdd.n2455 vdd.n1187 19.3944
R4144 vdd.n2455 vdd.n2454 19.3944
R4145 vdd.n2454 vdd.n2453 19.3944
R4146 vdd.n2453 vdd.n1194 19.3944
R4147 vdd.n2448 vdd.n1194 19.3944
R4148 vdd.n2448 vdd.n2447 19.3944
R4149 vdd.n2447 vdd.n2446 19.3944
R4150 vdd.n2446 vdd.n1201 19.3944
R4151 vdd.n2441 vdd.n1201 19.3944
R4152 vdd.n2441 vdd.n2440 19.3944
R4153 vdd.n1880 vdd.n1645 19.3944
R4154 vdd.n1880 vdd.n1636 19.3944
R4155 vdd.n1893 vdd.n1636 19.3944
R4156 vdd.n1893 vdd.n1634 19.3944
R4157 vdd.n1897 vdd.n1634 19.3944
R4158 vdd.n1897 vdd.n1625 19.3944
R4159 vdd.n1910 vdd.n1625 19.3944
R4160 vdd.n1910 vdd.n1623 19.3944
R4161 vdd.n1914 vdd.n1623 19.3944
R4162 vdd.n1914 vdd.n1614 19.3944
R4163 vdd.n1926 vdd.n1614 19.3944
R4164 vdd.n1926 vdd.n1612 19.3944
R4165 vdd.n1930 vdd.n1612 19.3944
R4166 vdd.n1930 vdd.n1602 19.3944
R4167 vdd.n1943 vdd.n1602 19.3944
R4168 vdd.n1943 vdd.n1600 19.3944
R4169 vdd.n1947 vdd.n1600 19.3944
R4170 vdd.n1947 vdd.n1591 19.3944
R4171 vdd.n1959 vdd.n1591 19.3944
R4172 vdd.n1959 vdd.n1589 19.3944
R4173 vdd.n2270 vdd.n1589 19.3944
R4174 vdd.n2270 vdd.n1579 19.3944
R4175 vdd.n2283 vdd.n1579 19.3944
R4176 vdd.n2283 vdd.n1577 19.3944
R4177 vdd.n2287 vdd.n1577 19.3944
R4178 vdd.n2287 vdd.n1568 19.3944
R4179 vdd.n2300 vdd.n1568 19.3944
R4180 vdd.n2300 vdd.n1566 19.3944
R4181 vdd.n2304 vdd.n1566 19.3944
R4182 vdd.n2304 vdd.n1557 19.3944
R4183 vdd.n2316 vdd.n1557 19.3944
R4184 vdd.n2316 vdd.n1555 19.3944
R4185 vdd.n2320 vdd.n1555 19.3944
R4186 vdd.n2320 vdd.n1545 19.3944
R4187 vdd.n2333 vdd.n1545 19.3944
R4188 vdd.n2333 vdd.n1543 19.3944
R4189 vdd.n2337 vdd.n1543 19.3944
R4190 vdd.n2337 vdd.n1533 19.3944
R4191 vdd.n2352 vdd.n1533 19.3944
R4192 vdd.n2352 vdd.n1531 19.3944
R4193 vdd.n2356 vdd.n1531 19.3944
R4194 vdd.n3501 vdd.n686 19.3944
R4195 vdd.n3501 vdd.n676 19.3944
R4196 vdd.n3513 vdd.n676 19.3944
R4197 vdd.n3513 vdd.n674 19.3944
R4198 vdd.n3517 vdd.n674 19.3944
R4199 vdd.n3517 vdd.n666 19.3944
R4200 vdd.n3530 vdd.n666 19.3944
R4201 vdd.n3530 vdd.n664 19.3944
R4202 vdd.n3534 vdd.n664 19.3944
R4203 vdd.n3534 vdd.n653 19.3944
R4204 vdd.n3546 vdd.n653 19.3944
R4205 vdd.n3546 vdd.n651 19.3944
R4206 vdd.n3550 vdd.n651 19.3944
R4207 vdd.n3550 vdd.n642 19.3944
R4208 vdd.n3563 vdd.n642 19.3944
R4209 vdd.n3563 vdd.n640 19.3944
R4210 vdd.n3570 vdd.n640 19.3944
R4211 vdd.n3570 vdd.n3569 19.3944
R4212 vdd.n3569 vdd.n631 19.3944
R4213 vdd.n3583 vdd.n631 19.3944
R4214 vdd.n3584 vdd.n3583 19.3944
R4215 vdd.n3584 vdd.n629 19.3944
R4216 vdd.n3588 vdd.n629 19.3944
R4217 vdd.n3590 vdd.n3588 19.3944
R4218 vdd.n3591 vdd.n3590 19.3944
R4219 vdd.n3591 vdd.n627 19.3944
R4220 vdd.n3595 vdd.n627 19.3944
R4221 vdd.n3597 vdd.n3595 19.3944
R4222 vdd.n3598 vdd.n3597 19.3944
R4223 vdd.n3598 vdd.n625 19.3944
R4224 vdd.n3602 vdd.n625 19.3944
R4225 vdd.n3605 vdd.n3602 19.3944
R4226 vdd.n3606 vdd.n3605 19.3944
R4227 vdd.n3606 vdd.n623 19.3944
R4228 vdd.n3610 vdd.n623 19.3944
R4229 vdd.n3612 vdd.n3610 19.3944
R4230 vdd.n3613 vdd.n3612 19.3944
R4231 vdd.n3613 vdd.n621 19.3944
R4232 vdd.n3617 vdd.n621 19.3944
R4233 vdd.n3619 vdd.n3617 19.3944
R4234 vdd.n3620 vdd.n3619 19.3944
R4235 vdd.n569 vdd.n438 19.3944
R4236 vdd.n575 vdd.n438 19.3944
R4237 vdd.n576 vdd.n575 19.3944
R4238 vdd.n579 vdd.n576 19.3944
R4239 vdd.n579 vdd.n436 19.3944
R4240 vdd.n585 vdd.n436 19.3944
R4241 vdd.n586 vdd.n585 19.3944
R4242 vdd.n589 vdd.n586 19.3944
R4243 vdd.n589 vdd.n434 19.3944
R4244 vdd.n595 vdd.n434 19.3944
R4245 vdd.n596 vdd.n595 19.3944
R4246 vdd.n599 vdd.n596 19.3944
R4247 vdd.n599 vdd.n432 19.3944
R4248 vdd.n605 vdd.n432 19.3944
R4249 vdd.n606 vdd.n605 19.3944
R4250 vdd.n609 vdd.n606 19.3944
R4251 vdd.n609 vdd.n430 19.3944
R4252 vdd.n615 vdd.n430 19.3944
R4253 vdd.n617 vdd.n615 19.3944
R4254 vdd.n618 vdd.n617 19.3944
R4255 vdd.n516 vdd.n515 19.3944
R4256 vdd.n519 vdd.n516 19.3944
R4257 vdd.n519 vdd.n450 19.3944
R4258 vdd.n525 vdd.n450 19.3944
R4259 vdd.n526 vdd.n525 19.3944
R4260 vdd.n529 vdd.n526 19.3944
R4261 vdd.n529 vdd.n448 19.3944
R4262 vdd.n535 vdd.n448 19.3944
R4263 vdd.n536 vdd.n535 19.3944
R4264 vdd.n539 vdd.n536 19.3944
R4265 vdd.n539 vdd.n446 19.3944
R4266 vdd.n545 vdd.n446 19.3944
R4267 vdd.n546 vdd.n545 19.3944
R4268 vdd.n549 vdd.n546 19.3944
R4269 vdd.n549 vdd.n444 19.3944
R4270 vdd.n555 vdd.n444 19.3944
R4271 vdd.n556 vdd.n555 19.3944
R4272 vdd.n559 vdd.n556 19.3944
R4273 vdd.n559 vdd.n442 19.3944
R4274 vdd.n565 vdd.n442 19.3944
R4275 vdd.n466 vdd.n465 19.3944
R4276 vdd.n469 vdd.n466 19.3944
R4277 vdd.n469 vdd.n462 19.3944
R4278 vdd.n475 vdd.n462 19.3944
R4279 vdd.n476 vdd.n475 19.3944
R4280 vdd.n479 vdd.n476 19.3944
R4281 vdd.n479 vdd.n460 19.3944
R4282 vdd.n485 vdd.n460 19.3944
R4283 vdd.n486 vdd.n485 19.3944
R4284 vdd.n489 vdd.n486 19.3944
R4285 vdd.n489 vdd.n458 19.3944
R4286 vdd.n495 vdd.n458 19.3944
R4287 vdd.n496 vdd.n495 19.3944
R4288 vdd.n499 vdd.n496 19.3944
R4289 vdd.n499 vdd.n456 19.3944
R4290 vdd.n505 vdd.n456 19.3944
R4291 vdd.n506 vdd.n505 19.3944
R4292 vdd.n509 vdd.n506 19.3944
R4293 vdd.n3505 vdd.n683 19.3944
R4294 vdd.n3505 vdd.n681 19.3944
R4295 vdd.n3509 vdd.n681 19.3944
R4296 vdd.n3509 vdd.n671 19.3944
R4297 vdd.n3522 vdd.n671 19.3944
R4298 vdd.n3522 vdd.n669 19.3944
R4299 vdd.n3526 vdd.n669 19.3944
R4300 vdd.n3526 vdd.n660 19.3944
R4301 vdd.n3538 vdd.n660 19.3944
R4302 vdd.n3538 vdd.n658 19.3944
R4303 vdd.n3542 vdd.n658 19.3944
R4304 vdd.n3542 vdd.n648 19.3944
R4305 vdd.n3555 vdd.n648 19.3944
R4306 vdd.n3555 vdd.n646 19.3944
R4307 vdd.n3559 vdd.n646 19.3944
R4308 vdd.n3559 vdd.n637 19.3944
R4309 vdd.n3574 vdd.n637 19.3944
R4310 vdd.n3574 vdd.n635 19.3944
R4311 vdd.n3578 vdd.n635 19.3944
R4312 vdd.n3578 vdd.n336 19.3944
R4313 vdd.n3669 vdd.n336 19.3944
R4314 vdd.n3669 vdd.n337 19.3944
R4315 vdd.n3663 vdd.n337 19.3944
R4316 vdd.n3663 vdd.n3662 19.3944
R4317 vdd.n3662 vdd.n3661 19.3944
R4318 vdd.n3661 vdd.n349 19.3944
R4319 vdd.n3655 vdd.n349 19.3944
R4320 vdd.n3655 vdd.n3654 19.3944
R4321 vdd.n3654 vdd.n3653 19.3944
R4322 vdd.n3653 vdd.n359 19.3944
R4323 vdd.n3647 vdd.n359 19.3944
R4324 vdd.n3647 vdd.n3646 19.3944
R4325 vdd.n3646 vdd.n3645 19.3944
R4326 vdd.n3645 vdd.n370 19.3944
R4327 vdd.n3639 vdd.n370 19.3944
R4328 vdd.n3639 vdd.n3638 19.3944
R4329 vdd.n3638 vdd.n3637 19.3944
R4330 vdd.n3637 vdd.n381 19.3944
R4331 vdd.n3631 vdd.n381 19.3944
R4332 vdd.n3631 vdd.n3630 19.3944
R4333 vdd.n3630 vdd.n3629 19.3944
R4334 vdd.n3452 vdd.n747 19.3944
R4335 vdd.n3452 vdd.n3449 19.3944
R4336 vdd.n3449 vdd.n3446 19.3944
R4337 vdd.n3446 vdd.n3445 19.3944
R4338 vdd.n3445 vdd.n3442 19.3944
R4339 vdd.n3442 vdd.n3441 19.3944
R4340 vdd.n3441 vdd.n3438 19.3944
R4341 vdd.n3438 vdd.n3437 19.3944
R4342 vdd.n3437 vdd.n3434 19.3944
R4343 vdd.n3434 vdd.n3433 19.3944
R4344 vdd.n3433 vdd.n3430 19.3944
R4345 vdd.n3430 vdd.n3429 19.3944
R4346 vdd.n3429 vdd.n3426 19.3944
R4347 vdd.n3426 vdd.n3425 19.3944
R4348 vdd.n3425 vdd.n3422 19.3944
R4349 vdd.n3422 vdd.n3421 19.3944
R4350 vdd.n3421 vdd.n3418 19.3944
R4351 vdd.n3418 vdd.n3417 19.3944
R4352 vdd.n3417 vdd.n3414 19.3944
R4353 vdd.n3414 vdd.n3413 19.3944
R4354 vdd.n3492 vdd.n3491 19.3944
R4355 vdd.n3491 vdd.n3490 19.3944
R4356 vdd.n732 vdd.n729 19.3944
R4357 vdd.n3486 vdd.n3485 19.3944
R4358 vdd.n3485 vdd.n3482 19.3944
R4359 vdd.n3482 vdd.n3481 19.3944
R4360 vdd.n3481 vdd.n3478 19.3944
R4361 vdd.n3478 vdd.n3477 19.3944
R4362 vdd.n3477 vdd.n3474 19.3944
R4363 vdd.n3474 vdd.n3473 19.3944
R4364 vdd.n3473 vdd.n3470 19.3944
R4365 vdd.n3470 vdd.n3469 19.3944
R4366 vdd.n3469 vdd.n3466 19.3944
R4367 vdd.n3466 vdd.n3465 19.3944
R4368 vdd.n3465 vdd.n3462 19.3944
R4369 vdd.n3462 vdd.n3461 19.3944
R4370 vdd.n3406 vdd.n767 19.3944
R4371 vdd.n3406 vdd.n3403 19.3944
R4372 vdd.n3403 vdd.n3400 19.3944
R4373 vdd.n3400 vdd.n3399 19.3944
R4374 vdd.n3399 vdd.n3396 19.3944
R4375 vdd.n3396 vdd.n3395 19.3944
R4376 vdd.n3395 vdd.n3392 19.3944
R4377 vdd.n3392 vdd.n3391 19.3944
R4378 vdd.n3391 vdd.n3388 19.3944
R4379 vdd.n3388 vdd.n3387 19.3944
R4380 vdd.n3387 vdd.n3384 19.3944
R4381 vdd.n3384 vdd.n3383 19.3944
R4382 vdd.n3383 vdd.n3380 19.3944
R4383 vdd.n3380 vdd.n3379 19.3944
R4384 vdd.n3379 vdd.n3376 19.3944
R4385 vdd.n3376 vdd.n3375 19.3944
R4386 vdd.n3372 vdd.n3371 19.3944
R4387 vdd.n3368 vdd.n3367 19.3944
R4388 vdd.n1812 vdd.n1808 19.0066
R4389 vdd.n2400 vdd.n1247 19.0066
R4390 vdd.n569 vdd.n566 19.0066
R4391 vdd.n3410 vdd.n767 19.0066
R4392 vdd.n1316 vdd.n1315 16.0975
R4393 vdd.n1011 vdd.n1010 16.0975
R4394 vdd.n1773 vdd.n1772 16.0975
R4395 vdd.n1811 vdd.n1810 16.0975
R4396 vdd.n1707 vdd.n1706 16.0975
R4397 vdd.n2363 vdd.n2362 16.0975
R4398 vdd.n1249 vdd.n1248 16.0975
R4399 vdd.n1209 vdd.n1208 16.0975
R4400 vdd.n1320 vdd.n1319 16.0975
R4401 vdd.n1002 vdd.n1001 16.0975
R4402 vdd.n2824 vdd.n2823 16.0975
R4403 vdd.n427 vdd.n426 16.0975
R4404 vdd.n441 vdd.n440 16.0975
R4405 vdd.n453 vdd.n452 16.0975
R4406 vdd.n769 vdd.n768 16.0975
R4407 vdd.n3457 vdd.n3456 16.0975
R4408 vdd.n833 vdd.n832 16.0975
R4409 vdd.n2821 vdd.n2820 16.0975
R4410 vdd.n689 vdd.n688 16.0975
R4411 vdd.n800 vdd.n799 16.0975
R4412 vdd.t169 vdd.n2784 15.4182
R4413 vdd.n3088 vdd.t156 15.4182
R4414 vdd.n28 vdd.n27 14.6072
R4415 vdd.n328 vdd.n293 13.1884
R4416 vdd.n269 vdd.n234 13.1884
R4417 vdd.n226 vdd.n191 13.1884
R4418 vdd.n167 vdd.n132 13.1884
R4419 vdd.n125 vdd.n90 13.1884
R4420 vdd.n66 vdd.n31 13.1884
R4421 vdd.n2202 vdd.n2167 13.1884
R4422 vdd.n2261 vdd.n2226 13.1884
R4423 vdd.n2100 vdd.n2065 13.1884
R4424 vdd.n2159 vdd.n2124 13.1884
R4425 vdd.n1999 vdd.n1964 13.1884
R4426 vdd.n2058 vdd.n2023 13.1884
R4427 vdd.n2506 vdd.n1134 13.1509
R4428 vdd.n3331 vdd.n692 13.1509
R4429 vdd.n1843 vdd.n1708 12.9944
R4430 vdd.n1847 vdd.n1708 12.9944
R4431 vdd.n2439 vdd.n1207 12.9944
R4432 vdd.n2440 vdd.n2439 12.9944
R4433 vdd.n515 vdd.n454 12.9944
R4434 vdd.n509 vdd.n454 12.9944
R4435 vdd.n3458 vdd.n747 12.9944
R4436 vdd.n3461 vdd.n3458 12.9944
R4437 vdd.n329 vdd.n291 12.8005
R4438 vdd.n324 vdd.n295 12.8005
R4439 vdd.n270 vdd.n232 12.8005
R4440 vdd.n265 vdd.n236 12.8005
R4441 vdd.n227 vdd.n189 12.8005
R4442 vdd.n222 vdd.n193 12.8005
R4443 vdd.n168 vdd.n130 12.8005
R4444 vdd.n163 vdd.n134 12.8005
R4445 vdd.n126 vdd.n88 12.8005
R4446 vdd.n121 vdd.n92 12.8005
R4447 vdd.n67 vdd.n29 12.8005
R4448 vdd.n62 vdd.n33 12.8005
R4449 vdd.n2203 vdd.n2165 12.8005
R4450 vdd.n2198 vdd.n2169 12.8005
R4451 vdd.n2262 vdd.n2224 12.8005
R4452 vdd.n2257 vdd.n2228 12.8005
R4453 vdd.n2101 vdd.n2063 12.8005
R4454 vdd.n2096 vdd.n2067 12.8005
R4455 vdd.n2160 vdd.n2122 12.8005
R4456 vdd.n2155 vdd.n2126 12.8005
R4457 vdd.n2000 vdd.n1962 12.8005
R4458 vdd.n1995 vdd.n1966 12.8005
R4459 vdd.n2059 vdd.n2021 12.8005
R4460 vdd.n2054 vdd.n2025 12.8005
R4461 vdd.n323 vdd.n296 12.0247
R4462 vdd.n264 vdd.n237 12.0247
R4463 vdd.n221 vdd.n194 12.0247
R4464 vdd.n162 vdd.n135 12.0247
R4465 vdd.n120 vdd.n93 12.0247
R4466 vdd.n61 vdd.n34 12.0247
R4467 vdd.n2197 vdd.n2170 12.0247
R4468 vdd.n2256 vdd.n2229 12.0247
R4469 vdd.n2095 vdd.n2068 12.0247
R4470 vdd.n2154 vdd.n2127 12.0247
R4471 vdd.n1994 vdd.n1967 12.0247
R4472 vdd.n2053 vdd.n2026 12.0247
R4473 vdd.n1882 vdd.n1638 11.337
R4474 vdd.n1891 vdd.n1638 11.337
R4475 vdd.n1891 vdd.n1890 11.337
R4476 vdd.n1899 vdd.n1632 11.337
R4477 vdd.n1908 vdd.n1907 11.337
R4478 vdd.n1924 vdd.n1616 11.337
R4479 vdd.n1932 vdd.n1609 11.337
R4480 vdd.n1941 vdd.n1940 11.337
R4481 vdd.n1949 vdd.n1598 11.337
R4482 vdd.n2272 vdd.n1587 11.337
R4483 vdd.n2281 vdd.n1581 11.337
R4484 vdd.n2289 vdd.n1575 11.337
R4485 vdd.n2298 vdd.n2297 11.337
R4486 vdd.n2314 vdd.n1559 11.337
R4487 vdd.n2322 vdd.n1552 11.337
R4488 vdd.n2331 vdd.n2330 11.337
R4489 vdd.n2339 vdd.n1535 11.337
R4490 vdd.n2350 vdd.n1535 11.337
R4491 vdd.n2350 vdd.n2349 11.337
R4492 vdd.n3503 vdd.n678 11.337
R4493 vdd.n3511 vdd.n678 11.337
R4494 vdd.n3511 vdd.n679 11.337
R4495 vdd.n3520 vdd.n3519 11.337
R4496 vdd.n3536 vdd.n662 11.337
R4497 vdd.n3544 vdd.n655 11.337
R4498 vdd.n3553 vdd.n3552 11.337
R4499 vdd.n3561 vdd.n644 11.337
R4500 vdd.n3580 vdd.n633 11.337
R4501 vdd.n3667 vdd.n340 11.337
R4502 vdd.n3665 vdd.n344 11.337
R4503 vdd.n3659 vdd.n3658 11.337
R4504 vdd.n3651 vdd.n361 11.337
R4505 vdd.n3650 vdd.n3649 11.337
R4506 vdd.n3643 vdd.n3642 11.337
R4507 vdd.n3641 vdd.n375 11.337
R4508 vdd.n3635 vdd.n3634 11.337
R4509 vdd.n3634 vdd.n3633 11.337
R4510 vdd.n3633 vdd.n386 11.337
R4511 vdd.n320 vdd.n319 11.249
R4512 vdd.n261 vdd.n260 11.249
R4513 vdd.n218 vdd.n217 11.249
R4514 vdd.n159 vdd.n158 11.249
R4515 vdd.n117 vdd.n116 11.249
R4516 vdd.n58 vdd.n57 11.249
R4517 vdd.n2194 vdd.n2193 11.249
R4518 vdd.n2253 vdd.n2252 11.249
R4519 vdd.n2092 vdd.n2091 11.249
R4520 vdd.n2151 vdd.n2150 11.249
R4521 vdd.n1991 vdd.n1990 11.249
R4522 vdd.n2050 vdd.n2049 11.249
R4523 vdd.n1680 vdd.t296 11.2237
R4524 vdd.n3627 vdd.t245 11.2237
R4525 vdd.t91 vdd.n1553 10.7702
R4526 vdd.n3528 vdd.t123 10.7702
R4527 vdd.n305 vdd.n304 10.7238
R4528 vdd.n246 vdd.n245 10.7238
R4529 vdd.n203 vdd.n202 10.7238
R4530 vdd.n144 vdd.n143 10.7238
R4531 vdd.n102 vdd.n101 10.7238
R4532 vdd.n43 vdd.n42 10.7238
R4533 vdd.n2179 vdd.n2178 10.7238
R4534 vdd.n2238 vdd.n2237 10.7238
R4535 vdd.n2077 vdd.n2076 10.7238
R4536 vdd.n2136 vdd.n2135 10.7238
R4537 vdd.n1976 vdd.n1975 10.7238
R4538 vdd.n2035 vdd.n2034 10.7238
R4539 vdd.n2511 vdd.n2510 10.6151
R4540 vdd.n2511 vdd.n1127 10.6151
R4541 vdd.n2521 vdd.n1127 10.6151
R4542 vdd.n2522 vdd.n2521 10.6151
R4543 vdd.n2523 vdd.n2522 10.6151
R4544 vdd.n2523 vdd.n1114 10.6151
R4545 vdd.n2533 vdd.n1114 10.6151
R4546 vdd.n2534 vdd.n2533 10.6151
R4547 vdd.n2535 vdd.n2534 10.6151
R4548 vdd.n2535 vdd.n1102 10.6151
R4549 vdd.n2545 vdd.n1102 10.6151
R4550 vdd.n2546 vdd.n2545 10.6151
R4551 vdd.n2547 vdd.n2546 10.6151
R4552 vdd.n2547 vdd.n1091 10.6151
R4553 vdd.n2557 vdd.n1091 10.6151
R4554 vdd.n2558 vdd.n2557 10.6151
R4555 vdd.n2559 vdd.n2558 10.6151
R4556 vdd.n2559 vdd.n1078 10.6151
R4557 vdd.n2569 vdd.n1078 10.6151
R4558 vdd.n2570 vdd.n2569 10.6151
R4559 vdd.n2571 vdd.n2570 10.6151
R4560 vdd.n2571 vdd.n1066 10.6151
R4561 vdd.n2582 vdd.n1066 10.6151
R4562 vdd.n2583 vdd.n2582 10.6151
R4563 vdd.n2584 vdd.n2583 10.6151
R4564 vdd.n2584 vdd.n1054 10.6151
R4565 vdd.n2594 vdd.n1054 10.6151
R4566 vdd.n2595 vdd.n2594 10.6151
R4567 vdd.n2596 vdd.n2595 10.6151
R4568 vdd.n2596 vdd.n1042 10.6151
R4569 vdd.n2606 vdd.n1042 10.6151
R4570 vdd.n2607 vdd.n2606 10.6151
R4571 vdd.n2608 vdd.n2607 10.6151
R4572 vdd.n2608 vdd.n1032 10.6151
R4573 vdd.n2618 vdd.n1032 10.6151
R4574 vdd.n2619 vdd.n2618 10.6151
R4575 vdd.n2620 vdd.n2619 10.6151
R4576 vdd.n2620 vdd.n1019 10.6151
R4577 vdd.n2632 vdd.n1019 10.6151
R4578 vdd.n2633 vdd.n2632 10.6151
R4579 vdd.n2635 vdd.n2633 10.6151
R4580 vdd.n2635 vdd.n2634 10.6151
R4581 vdd.n2634 vdd.n1000 10.6151
R4582 vdd.n2782 vdd.n2781 10.6151
R4583 vdd.n2781 vdd.n2780 10.6151
R4584 vdd.n2780 vdd.n2777 10.6151
R4585 vdd.n2777 vdd.n2776 10.6151
R4586 vdd.n2776 vdd.n2773 10.6151
R4587 vdd.n2773 vdd.n2772 10.6151
R4588 vdd.n2772 vdd.n2769 10.6151
R4589 vdd.n2769 vdd.n2768 10.6151
R4590 vdd.n2768 vdd.n2765 10.6151
R4591 vdd.n2765 vdd.n2764 10.6151
R4592 vdd.n2764 vdd.n2761 10.6151
R4593 vdd.n2761 vdd.n2760 10.6151
R4594 vdd.n2760 vdd.n2757 10.6151
R4595 vdd.n2757 vdd.n2756 10.6151
R4596 vdd.n2756 vdd.n2753 10.6151
R4597 vdd.n2753 vdd.n2752 10.6151
R4598 vdd.n2752 vdd.n2749 10.6151
R4599 vdd.n2749 vdd.n2748 10.6151
R4600 vdd.n2748 vdd.n2745 10.6151
R4601 vdd.n2745 vdd.n2744 10.6151
R4602 vdd.n2744 vdd.n2741 10.6151
R4603 vdd.n2741 vdd.n2740 10.6151
R4604 vdd.n2740 vdd.n2737 10.6151
R4605 vdd.n2737 vdd.n2736 10.6151
R4606 vdd.n2736 vdd.n2733 10.6151
R4607 vdd.n2733 vdd.n2732 10.6151
R4608 vdd.n2732 vdd.n2729 10.6151
R4609 vdd.n2729 vdd.n2728 10.6151
R4610 vdd.n2728 vdd.n2725 10.6151
R4611 vdd.n2725 vdd.n2724 10.6151
R4612 vdd.n2724 vdd.n2721 10.6151
R4613 vdd.n2719 vdd.n2716 10.6151
R4614 vdd.n2716 vdd.n2715 10.6151
R4615 vdd.n1357 vdd.n1356 10.6151
R4616 vdd.n1359 vdd.n1357 10.6151
R4617 vdd.n1360 vdd.n1359 10.6151
R4618 vdd.n1362 vdd.n1360 10.6151
R4619 vdd.n1363 vdd.n1362 10.6151
R4620 vdd.n1365 vdd.n1363 10.6151
R4621 vdd.n1366 vdd.n1365 10.6151
R4622 vdd.n1368 vdd.n1366 10.6151
R4623 vdd.n1369 vdd.n1368 10.6151
R4624 vdd.n1371 vdd.n1369 10.6151
R4625 vdd.n1372 vdd.n1371 10.6151
R4626 vdd.n1374 vdd.n1372 10.6151
R4627 vdd.n1375 vdd.n1374 10.6151
R4628 vdd.n1377 vdd.n1375 10.6151
R4629 vdd.n1378 vdd.n1377 10.6151
R4630 vdd.n1380 vdd.n1378 10.6151
R4631 vdd.n1381 vdd.n1380 10.6151
R4632 vdd.n1383 vdd.n1381 10.6151
R4633 vdd.n1384 vdd.n1383 10.6151
R4634 vdd.n1386 vdd.n1384 10.6151
R4635 vdd.n1387 vdd.n1386 10.6151
R4636 vdd.n1389 vdd.n1387 10.6151
R4637 vdd.n1390 vdd.n1389 10.6151
R4638 vdd.n1392 vdd.n1390 10.6151
R4639 vdd.n1393 vdd.n1392 10.6151
R4640 vdd.n1395 vdd.n1393 10.6151
R4641 vdd.n1396 vdd.n1395 10.6151
R4642 vdd.n1435 vdd.n1396 10.6151
R4643 vdd.n1435 vdd.n1434 10.6151
R4644 vdd.n1434 vdd.n1433 10.6151
R4645 vdd.n1433 vdd.n1431 10.6151
R4646 vdd.n1431 vdd.n1430 10.6151
R4647 vdd.n1430 vdd.n1428 10.6151
R4648 vdd.n1428 vdd.n1427 10.6151
R4649 vdd.n1427 vdd.n1408 10.6151
R4650 vdd.n1408 vdd.n1407 10.6151
R4651 vdd.n1407 vdd.n1405 10.6151
R4652 vdd.n1405 vdd.n1404 10.6151
R4653 vdd.n1404 vdd.n1402 10.6151
R4654 vdd.n1402 vdd.n1401 10.6151
R4655 vdd.n1401 vdd.n1398 10.6151
R4656 vdd.n1398 vdd.n1397 10.6151
R4657 vdd.n1397 vdd.n1003 10.6151
R4658 vdd.n2509 vdd.n1139 10.6151
R4659 vdd.n2504 vdd.n1139 10.6151
R4660 vdd.n2504 vdd.n2503 10.6151
R4661 vdd.n2503 vdd.n2502 10.6151
R4662 vdd.n2502 vdd.n2499 10.6151
R4663 vdd.n2499 vdd.n2498 10.6151
R4664 vdd.n2498 vdd.n2495 10.6151
R4665 vdd.n2495 vdd.n2494 10.6151
R4666 vdd.n2494 vdd.n2491 10.6151
R4667 vdd.n2491 vdd.n2490 10.6151
R4668 vdd.n2490 vdd.n2487 10.6151
R4669 vdd.n2487 vdd.n2486 10.6151
R4670 vdd.n2486 vdd.n2483 10.6151
R4671 vdd.n2483 vdd.n2482 10.6151
R4672 vdd.n2482 vdd.n2479 10.6151
R4673 vdd.n2479 vdd.n2478 10.6151
R4674 vdd.n2478 vdd.n2475 10.6151
R4675 vdd.n2475 vdd.n1177 10.6151
R4676 vdd.n1323 vdd.n1177 10.6151
R4677 vdd.n1324 vdd.n1323 10.6151
R4678 vdd.n1327 vdd.n1324 10.6151
R4679 vdd.n1328 vdd.n1327 10.6151
R4680 vdd.n1331 vdd.n1328 10.6151
R4681 vdd.n1332 vdd.n1331 10.6151
R4682 vdd.n1335 vdd.n1332 10.6151
R4683 vdd.n1336 vdd.n1335 10.6151
R4684 vdd.n1339 vdd.n1336 10.6151
R4685 vdd.n1340 vdd.n1339 10.6151
R4686 vdd.n1343 vdd.n1340 10.6151
R4687 vdd.n1344 vdd.n1343 10.6151
R4688 vdd.n1347 vdd.n1344 10.6151
R4689 vdd.n1352 vdd.n1349 10.6151
R4690 vdd.n1353 vdd.n1352 10.6151
R4691 vdd.n3020 vdd.n3019 10.6151
R4692 vdd.n3019 vdd.n3018 10.6151
R4693 vdd.n3018 vdd.n2822 10.6151
R4694 vdd.n2900 vdd.n2822 10.6151
R4695 vdd.n2901 vdd.n2900 10.6151
R4696 vdd.n2903 vdd.n2901 10.6151
R4697 vdd.n2904 vdd.n2903 10.6151
R4698 vdd.n3002 vdd.n2904 10.6151
R4699 vdd.n3002 vdd.n3001 10.6151
R4700 vdd.n3001 vdd.n3000 10.6151
R4701 vdd.n3000 vdd.n2948 10.6151
R4702 vdd.n2948 vdd.n2947 10.6151
R4703 vdd.n2947 vdd.n2945 10.6151
R4704 vdd.n2945 vdd.n2944 10.6151
R4705 vdd.n2944 vdd.n2942 10.6151
R4706 vdd.n2942 vdd.n2941 10.6151
R4707 vdd.n2941 vdd.n2939 10.6151
R4708 vdd.n2939 vdd.n2938 10.6151
R4709 vdd.n2938 vdd.n2936 10.6151
R4710 vdd.n2936 vdd.n2935 10.6151
R4711 vdd.n2935 vdd.n2933 10.6151
R4712 vdd.n2933 vdd.n2932 10.6151
R4713 vdd.n2932 vdd.n2930 10.6151
R4714 vdd.n2930 vdd.n2929 10.6151
R4715 vdd.n2929 vdd.n2927 10.6151
R4716 vdd.n2927 vdd.n2926 10.6151
R4717 vdd.n2926 vdd.n2924 10.6151
R4718 vdd.n2924 vdd.n2923 10.6151
R4719 vdd.n2923 vdd.n2921 10.6151
R4720 vdd.n2921 vdd.n2920 10.6151
R4721 vdd.n2920 vdd.n2918 10.6151
R4722 vdd.n2918 vdd.n2917 10.6151
R4723 vdd.n2917 vdd.n2915 10.6151
R4724 vdd.n2915 vdd.n2914 10.6151
R4725 vdd.n2914 vdd.n2912 10.6151
R4726 vdd.n2912 vdd.n2911 10.6151
R4727 vdd.n2911 vdd.n2909 10.6151
R4728 vdd.n2909 vdd.n2908 10.6151
R4729 vdd.n2908 vdd.n2906 10.6151
R4730 vdd.n2906 vdd.n2905 10.6151
R4731 vdd.n2905 vdd.n836 10.6151
R4732 vdd.n3264 vdd.n836 10.6151
R4733 vdd.n3265 vdd.n3264 10.6151
R4734 vdd.n3091 vdd.n961 10.6151
R4735 vdd.n3086 vdd.n961 10.6151
R4736 vdd.n3086 vdd.n3085 10.6151
R4737 vdd.n3085 vdd.n3084 10.6151
R4738 vdd.n3084 vdd.n3081 10.6151
R4739 vdd.n3081 vdd.n3080 10.6151
R4740 vdd.n3080 vdd.n3077 10.6151
R4741 vdd.n3077 vdd.n3076 10.6151
R4742 vdd.n3076 vdd.n3073 10.6151
R4743 vdd.n3073 vdd.n3072 10.6151
R4744 vdd.n3072 vdd.n3069 10.6151
R4745 vdd.n3069 vdd.n3068 10.6151
R4746 vdd.n3068 vdd.n3065 10.6151
R4747 vdd.n3065 vdd.n3064 10.6151
R4748 vdd.n3064 vdd.n3061 10.6151
R4749 vdd.n3061 vdd.n3060 10.6151
R4750 vdd.n3060 vdd.n3057 10.6151
R4751 vdd.n3057 vdd.n3056 10.6151
R4752 vdd.n3056 vdd.n3053 10.6151
R4753 vdd.n3053 vdd.n3052 10.6151
R4754 vdd.n3052 vdd.n3049 10.6151
R4755 vdd.n3049 vdd.n3048 10.6151
R4756 vdd.n3048 vdd.n3045 10.6151
R4757 vdd.n3045 vdd.n3044 10.6151
R4758 vdd.n3044 vdd.n3041 10.6151
R4759 vdd.n3041 vdd.n3040 10.6151
R4760 vdd.n3040 vdd.n3037 10.6151
R4761 vdd.n3037 vdd.n3036 10.6151
R4762 vdd.n3036 vdd.n3033 10.6151
R4763 vdd.n3033 vdd.n3032 10.6151
R4764 vdd.n3032 vdd.n3029 10.6151
R4765 vdd.n3027 vdd.n3024 10.6151
R4766 vdd.n3024 vdd.n3023 10.6151
R4767 vdd.n3093 vdd.n3092 10.6151
R4768 vdd.n3093 vdd.n950 10.6151
R4769 vdd.n3103 vdd.n950 10.6151
R4770 vdd.n3104 vdd.n3103 10.6151
R4771 vdd.n3105 vdd.n3104 10.6151
R4772 vdd.n3105 vdd.n938 10.6151
R4773 vdd.n3115 vdd.n938 10.6151
R4774 vdd.n3116 vdd.n3115 10.6151
R4775 vdd.n3117 vdd.n3116 10.6151
R4776 vdd.n3117 vdd.n927 10.6151
R4777 vdd.n3127 vdd.n927 10.6151
R4778 vdd.n3128 vdd.n3127 10.6151
R4779 vdd.n3129 vdd.n3128 10.6151
R4780 vdd.n3129 vdd.n916 10.6151
R4781 vdd.n3139 vdd.n916 10.6151
R4782 vdd.n3140 vdd.n3139 10.6151
R4783 vdd.n3141 vdd.n3140 10.6151
R4784 vdd.n3141 vdd.n903 10.6151
R4785 vdd.n3152 vdd.n903 10.6151
R4786 vdd.n3153 vdd.n3152 10.6151
R4787 vdd.n3154 vdd.n3153 10.6151
R4788 vdd.n3154 vdd.n891 10.6151
R4789 vdd.n3164 vdd.n891 10.6151
R4790 vdd.n3165 vdd.n3164 10.6151
R4791 vdd.n3166 vdd.n3165 10.6151
R4792 vdd.n3166 vdd.n879 10.6151
R4793 vdd.n3176 vdd.n879 10.6151
R4794 vdd.n3177 vdd.n3176 10.6151
R4795 vdd.n3178 vdd.n3177 10.6151
R4796 vdd.n3178 vdd.n866 10.6151
R4797 vdd.n3188 vdd.n866 10.6151
R4798 vdd.n3189 vdd.n3188 10.6151
R4799 vdd.n3190 vdd.n3189 10.6151
R4800 vdd.n3190 vdd.n855 10.6151
R4801 vdd.n3200 vdd.n855 10.6151
R4802 vdd.n3201 vdd.n3200 10.6151
R4803 vdd.n3202 vdd.n3201 10.6151
R4804 vdd.n3202 vdd.n841 10.6151
R4805 vdd.n3257 vdd.n841 10.6151
R4806 vdd.n3258 vdd.n3257 10.6151
R4807 vdd.n3259 vdd.n3258 10.6151
R4808 vdd.n3259 vdd.n810 10.6151
R4809 vdd.n3329 vdd.n810 10.6151
R4810 vdd.n3328 vdd.n3327 10.6151
R4811 vdd.n3327 vdd.n811 10.6151
R4812 vdd.n812 vdd.n811 10.6151
R4813 vdd.n3320 vdd.n812 10.6151
R4814 vdd.n3320 vdd.n3319 10.6151
R4815 vdd.n3319 vdd.n3318 10.6151
R4816 vdd.n3318 vdd.n814 10.6151
R4817 vdd.n3313 vdd.n814 10.6151
R4818 vdd.n3313 vdd.n3312 10.6151
R4819 vdd.n3312 vdd.n3311 10.6151
R4820 vdd.n3311 vdd.n817 10.6151
R4821 vdd.n3306 vdd.n817 10.6151
R4822 vdd.n3306 vdd.n3305 10.6151
R4823 vdd.n3305 vdd.n3304 10.6151
R4824 vdd.n3304 vdd.n820 10.6151
R4825 vdd.n3299 vdd.n820 10.6151
R4826 vdd.n3299 vdd.n731 10.6151
R4827 vdd.n3295 vdd.n731 10.6151
R4828 vdd.n3295 vdd.n3294 10.6151
R4829 vdd.n3294 vdd.n3293 10.6151
R4830 vdd.n3293 vdd.n823 10.6151
R4831 vdd.n3288 vdd.n823 10.6151
R4832 vdd.n3288 vdd.n3287 10.6151
R4833 vdd.n3287 vdd.n3286 10.6151
R4834 vdd.n3286 vdd.n826 10.6151
R4835 vdd.n3281 vdd.n826 10.6151
R4836 vdd.n3281 vdd.n3280 10.6151
R4837 vdd.n3280 vdd.n3279 10.6151
R4838 vdd.n3279 vdd.n829 10.6151
R4839 vdd.n3274 vdd.n829 10.6151
R4840 vdd.n3274 vdd.n3273 10.6151
R4841 vdd.n3271 vdd.n834 10.6151
R4842 vdd.n3266 vdd.n834 10.6151
R4843 vdd.n3247 vdd.n3208 10.6151
R4844 vdd.n3242 vdd.n3208 10.6151
R4845 vdd.n3242 vdd.n3241 10.6151
R4846 vdd.n3241 vdd.n3240 10.6151
R4847 vdd.n3240 vdd.n3210 10.6151
R4848 vdd.n3235 vdd.n3210 10.6151
R4849 vdd.n3235 vdd.n3234 10.6151
R4850 vdd.n3234 vdd.n3233 10.6151
R4851 vdd.n3233 vdd.n3213 10.6151
R4852 vdd.n3228 vdd.n3213 10.6151
R4853 vdd.n3228 vdd.n3227 10.6151
R4854 vdd.n3227 vdd.n3226 10.6151
R4855 vdd.n3226 vdd.n3216 10.6151
R4856 vdd.n3221 vdd.n3216 10.6151
R4857 vdd.n3221 vdd.n3220 10.6151
R4858 vdd.n3220 vdd.n785 10.6151
R4859 vdd.n3364 vdd.n785 10.6151
R4860 vdd.n3364 vdd.n786 10.6151
R4861 vdd.n788 vdd.n786 10.6151
R4862 vdd.n3357 vdd.n788 10.6151
R4863 vdd.n3357 vdd.n3356 10.6151
R4864 vdd.n3356 vdd.n3355 10.6151
R4865 vdd.n3355 vdd.n790 10.6151
R4866 vdd.n3350 vdd.n790 10.6151
R4867 vdd.n3350 vdd.n3349 10.6151
R4868 vdd.n3349 vdd.n3348 10.6151
R4869 vdd.n3348 vdd.n793 10.6151
R4870 vdd.n3343 vdd.n793 10.6151
R4871 vdd.n3343 vdd.n3342 10.6151
R4872 vdd.n3342 vdd.n3341 10.6151
R4873 vdd.n3341 vdd.n796 10.6151
R4874 vdd.n3336 vdd.n3335 10.6151
R4875 vdd.n3335 vdd.n3334 10.6151
R4876 vdd.n2897 vdd.n2896 10.6151
R4877 vdd.n3014 vdd.n2897 10.6151
R4878 vdd.n3014 vdd.n3013 10.6151
R4879 vdd.n3013 vdd.n3012 10.6151
R4880 vdd.n3012 vdd.n3010 10.6151
R4881 vdd.n3010 vdd.n3009 10.6151
R4882 vdd.n3009 vdd.n3007 10.6151
R4883 vdd.n3007 vdd.n3006 10.6151
R4884 vdd.n3006 vdd.n2898 10.6151
R4885 vdd.n2996 vdd.n2898 10.6151
R4886 vdd.n2996 vdd.n2995 10.6151
R4887 vdd.n2995 vdd.n2994 10.6151
R4888 vdd.n2994 vdd.n2992 10.6151
R4889 vdd.n2992 vdd.n2991 10.6151
R4890 vdd.n2991 vdd.n2989 10.6151
R4891 vdd.n2989 vdd.n2988 10.6151
R4892 vdd.n2988 vdd.n2986 10.6151
R4893 vdd.n2986 vdd.n2985 10.6151
R4894 vdd.n2985 vdd.n2983 10.6151
R4895 vdd.n2983 vdd.n2982 10.6151
R4896 vdd.n2982 vdd.n2980 10.6151
R4897 vdd.n2980 vdd.n2979 10.6151
R4898 vdd.n2979 vdd.n2977 10.6151
R4899 vdd.n2977 vdd.n2976 10.6151
R4900 vdd.n2976 vdd.n2974 10.6151
R4901 vdd.n2974 vdd.n2973 10.6151
R4902 vdd.n2973 vdd.n2971 10.6151
R4903 vdd.n2971 vdd.n2970 10.6151
R4904 vdd.n2970 vdd.n2968 10.6151
R4905 vdd.n2968 vdd.n2967 10.6151
R4906 vdd.n2967 vdd.n2965 10.6151
R4907 vdd.n2965 vdd.n2964 10.6151
R4908 vdd.n2964 vdd.n2962 10.6151
R4909 vdd.n2962 vdd.n2961 10.6151
R4910 vdd.n2961 vdd.n2959 10.6151
R4911 vdd.n2959 vdd.n2958 10.6151
R4912 vdd.n2958 vdd.n2956 10.6151
R4913 vdd.n2956 vdd.n2955 10.6151
R4914 vdd.n2955 vdd.n2953 10.6151
R4915 vdd.n2953 vdd.n2952 10.6151
R4916 vdd.n2952 vdd.n2950 10.6151
R4917 vdd.n2950 vdd.n2949 10.6151
R4918 vdd.n2949 vdd.n802 10.6151
R4919 vdd.n2828 vdd.n2827 10.6151
R4920 vdd.n2831 vdd.n2828 10.6151
R4921 vdd.n2832 vdd.n2831 10.6151
R4922 vdd.n2835 vdd.n2832 10.6151
R4923 vdd.n2836 vdd.n2835 10.6151
R4924 vdd.n2839 vdd.n2836 10.6151
R4925 vdd.n2840 vdd.n2839 10.6151
R4926 vdd.n2843 vdd.n2840 10.6151
R4927 vdd.n2844 vdd.n2843 10.6151
R4928 vdd.n2847 vdd.n2844 10.6151
R4929 vdd.n2848 vdd.n2847 10.6151
R4930 vdd.n2851 vdd.n2848 10.6151
R4931 vdd.n2852 vdd.n2851 10.6151
R4932 vdd.n2855 vdd.n2852 10.6151
R4933 vdd.n2856 vdd.n2855 10.6151
R4934 vdd.n2859 vdd.n2856 10.6151
R4935 vdd.n2860 vdd.n2859 10.6151
R4936 vdd.n2863 vdd.n2860 10.6151
R4937 vdd.n2864 vdd.n2863 10.6151
R4938 vdd.n2867 vdd.n2864 10.6151
R4939 vdd.n2868 vdd.n2867 10.6151
R4940 vdd.n2871 vdd.n2868 10.6151
R4941 vdd.n2872 vdd.n2871 10.6151
R4942 vdd.n2875 vdd.n2872 10.6151
R4943 vdd.n2876 vdd.n2875 10.6151
R4944 vdd.n2879 vdd.n2876 10.6151
R4945 vdd.n2880 vdd.n2879 10.6151
R4946 vdd.n2883 vdd.n2880 10.6151
R4947 vdd.n2884 vdd.n2883 10.6151
R4948 vdd.n2887 vdd.n2884 10.6151
R4949 vdd.n2888 vdd.n2887 10.6151
R4950 vdd.n2893 vdd.n2891 10.6151
R4951 vdd.n2894 vdd.n2893 10.6151
R4952 vdd.n3097 vdd.n955 10.6151
R4953 vdd.n3098 vdd.n3097 10.6151
R4954 vdd.n3099 vdd.n3098 10.6151
R4955 vdd.n3099 vdd.n944 10.6151
R4956 vdd.n3109 vdd.n944 10.6151
R4957 vdd.n3110 vdd.n3109 10.6151
R4958 vdd.n3111 vdd.n3110 10.6151
R4959 vdd.n3111 vdd.n933 10.6151
R4960 vdd.n3121 vdd.n933 10.6151
R4961 vdd.n3122 vdd.n3121 10.6151
R4962 vdd.n3123 vdd.n3122 10.6151
R4963 vdd.n3123 vdd.n921 10.6151
R4964 vdd.n3133 vdd.n921 10.6151
R4965 vdd.n3134 vdd.n3133 10.6151
R4966 vdd.n3135 vdd.n3134 10.6151
R4967 vdd.n3135 vdd.n910 10.6151
R4968 vdd.n3145 vdd.n910 10.6151
R4969 vdd.n3146 vdd.n3145 10.6151
R4970 vdd.n3148 vdd.n3146 10.6151
R4971 vdd.n3148 vdd.n3147 10.6151
R4972 vdd.n3159 vdd.n3158 10.6151
R4973 vdd.n3160 vdd.n3159 10.6151
R4974 vdd.n3160 vdd.n885 10.6151
R4975 vdd.n3170 vdd.n885 10.6151
R4976 vdd.n3171 vdd.n3170 10.6151
R4977 vdd.n3172 vdd.n3171 10.6151
R4978 vdd.n3172 vdd.n872 10.6151
R4979 vdd.n3182 vdd.n872 10.6151
R4980 vdd.n3183 vdd.n3182 10.6151
R4981 vdd.n3184 vdd.n3183 10.6151
R4982 vdd.n3184 vdd.n860 10.6151
R4983 vdd.n3194 vdd.n860 10.6151
R4984 vdd.n3195 vdd.n3194 10.6151
R4985 vdd.n3196 vdd.n3195 10.6151
R4986 vdd.n3196 vdd.n849 10.6151
R4987 vdd.n3206 vdd.n849 10.6151
R4988 vdd.n3207 vdd.n3206 10.6151
R4989 vdd.n3253 vdd.n3207 10.6151
R4990 vdd.n3253 vdd.n3252 10.6151
R4991 vdd.n3252 vdd.n3251 10.6151
R4992 vdd.n3251 vdd.n3250 10.6151
R4993 vdd.n3250 vdd.n3248 10.6151
R4994 vdd.n2515 vdd.n1132 10.6151
R4995 vdd.n2516 vdd.n2515 10.6151
R4996 vdd.n2517 vdd.n2516 10.6151
R4997 vdd.n2517 vdd.n1121 10.6151
R4998 vdd.n2527 vdd.n1121 10.6151
R4999 vdd.n2528 vdd.n2527 10.6151
R5000 vdd.n2529 vdd.n2528 10.6151
R5001 vdd.n2529 vdd.n1108 10.6151
R5002 vdd.n2539 vdd.n1108 10.6151
R5003 vdd.n2540 vdd.n2539 10.6151
R5004 vdd.n2541 vdd.n2540 10.6151
R5005 vdd.n2541 vdd.n1097 10.6151
R5006 vdd.n2551 vdd.n1097 10.6151
R5007 vdd.n2552 vdd.n2551 10.6151
R5008 vdd.n2553 vdd.n2552 10.6151
R5009 vdd.n2553 vdd.n1085 10.6151
R5010 vdd.n2563 vdd.n1085 10.6151
R5011 vdd.n2564 vdd.n2563 10.6151
R5012 vdd.n2565 vdd.n2564 10.6151
R5013 vdd.n2565 vdd.n1072 10.6151
R5014 vdd.n2575 vdd.n1072 10.6151
R5015 vdd.n2576 vdd.n2575 10.6151
R5016 vdd.n2578 vdd.n1060 10.6151
R5017 vdd.n2588 vdd.n1060 10.6151
R5018 vdd.n2589 vdd.n2588 10.6151
R5019 vdd.n2590 vdd.n2589 10.6151
R5020 vdd.n2590 vdd.n1048 10.6151
R5021 vdd.n2600 vdd.n1048 10.6151
R5022 vdd.n2601 vdd.n2600 10.6151
R5023 vdd.n2602 vdd.n2601 10.6151
R5024 vdd.n2602 vdd.n1037 10.6151
R5025 vdd.n2612 vdd.n1037 10.6151
R5026 vdd.n2613 vdd.n2612 10.6151
R5027 vdd.n2614 vdd.n2613 10.6151
R5028 vdd.n2614 vdd.n1026 10.6151
R5029 vdd.n2624 vdd.n1026 10.6151
R5030 vdd.n2625 vdd.n2624 10.6151
R5031 vdd.n2628 vdd.n2625 10.6151
R5032 vdd.n2628 vdd.n2627 10.6151
R5033 vdd.n2627 vdd.n2626 10.6151
R5034 vdd.n2626 vdd.n1009 10.6151
R5035 vdd.n2710 vdd.n1009 10.6151
R5036 vdd.n2709 vdd.n2708 10.6151
R5037 vdd.n2708 vdd.n2705 10.6151
R5038 vdd.n2705 vdd.n2704 10.6151
R5039 vdd.n2704 vdd.n2701 10.6151
R5040 vdd.n2701 vdd.n2700 10.6151
R5041 vdd.n2700 vdd.n2697 10.6151
R5042 vdd.n2697 vdd.n2696 10.6151
R5043 vdd.n2696 vdd.n2693 10.6151
R5044 vdd.n2693 vdd.n2692 10.6151
R5045 vdd.n2692 vdd.n2689 10.6151
R5046 vdd.n2689 vdd.n2688 10.6151
R5047 vdd.n2688 vdd.n2685 10.6151
R5048 vdd.n2685 vdd.n2684 10.6151
R5049 vdd.n2684 vdd.n2681 10.6151
R5050 vdd.n2681 vdd.n2680 10.6151
R5051 vdd.n2680 vdd.n2677 10.6151
R5052 vdd.n2677 vdd.n2676 10.6151
R5053 vdd.n2676 vdd.n2673 10.6151
R5054 vdd.n2673 vdd.n2672 10.6151
R5055 vdd.n2672 vdd.n2669 10.6151
R5056 vdd.n2669 vdd.n2668 10.6151
R5057 vdd.n2668 vdd.n2665 10.6151
R5058 vdd.n2665 vdd.n2664 10.6151
R5059 vdd.n2664 vdd.n2661 10.6151
R5060 vdd.n2661 vdd.n2660 10.6151
R5061 vdd.n2660 vdd.n2657 10.6151
R5062 vdd.n2657 vdd.n2656 10.6151
R5063 vdd.n2656 vdd.n2653 10.6151
R5064 vdd.n2653 vdd.n2652 10.6151
R5065 vdd.n2652 vdd.n2649 10.6151
R5066 vdd.n2649 vdd.n2648 10.6151
R5067 vdd.n2645 vdd.n2644 10.6151
R5068 vdd.n2644 vdd.n2642 10.6151
R5069 vdd.n1481 vdd.n1479 10.6151
R5070 vdd.n1479 vdd.n1478 10.6151
R5071 vdd.n1478 vdd.n1476 10.6151
R5072 vdd.n1476 vdd.n1475 10.6151
R5073 vdd.n1475 vdd.n1473 10.6151
R5074 vdd.n1473 vdd.n1472 10.6151
R5075 vdd.n1472 vdd.n1470 10.6151
R5076 vdd.n1470 vdd.n1469 10.6151
R5077 vdd.n1469 vdd.n1467 10.6151
R5078 vdd.n1467 vdd.n1466 10.6151
R5079 vdd.n1466 vdd.n1464 10.6151
R5080 vdd.n1464 vdd.n1463 10.6151
R5081 vdd.n1463 vdd.n1461 10.6151
R5082 vdd.n1461 vdd.n1460 10.6151
R5083 vdd.n1460 vdd.n1458 10.6151
R5084 vdd.n1458 vdd.n1457 10.6151
R5085 vdd.n1457 vdd.n1455 10.6151
R5086 vdd.n1455 vdd.n1454 10.6151
R5087 vdd.n1454 vdd.n1452 10.6151
R5088 vdd.n1452 vdd.n1451 10.6151
R5089 vdd.n1451 vdd.n1449 10.6151
R5090 vdd.n1449 vdd.n1448 10.6151
R5091 vdd.n1448 vdd.n1446 10.6151
R5092 vdd.n1446 vdd.n1445 10.6151
R5093 vdd.n1445 vdd.n1443 10.6151
R5094 vdd.n1443 vdd.n1442 10.6151
R5095 vdd.n1442 vdd.n1440 10.6151
R5096 vdd.n1440 vdd.n1439 10.6151
R5097 vdd.n1439 vdd.n1318 10.6151
R5098 vdd.n1410 vdd.n1318 10.6151
R5099 vdd.n1411 vdd.n1410 10.6151
R5100 vdd.n1413 vdd.n1411 10.6151
R5101 vdd.n1414 vdd.n1413 10.6151
R5102 vdd.n1423 vdd.n1414 10.6151
R5103 vdd.n1423 vdd.n1422 10.6151
R5104 vdd.n1422 vdd.n1421 10.6151
R5105 vdd.n1421 vdd.n1419 10.6151
R5106 vdd.n1419 vdd.n1418 10.6151
R5107 vdd.n1418 vdd.n1416 10.6151
R5108 vdd.n1416 vdd.n1415 10.6151
R5109 vdd.n1415 vdd.n1013 10.6151
R5110 vdd.n2640 vdd.n1013 10.6151
R5111 vdd.n2641 vdd.n2640 10.6151
R5112 vdd.n1282 vdd.n1281 10.6151
R5113 vdd.n1285 vdd.n1282 10.6151
R5114 vdd.n1286 vdd.n1285 10.6151
R5115 vdd.n1289 vdd.n1286 10.6151
R5116 vdd.n1290 vdd.n1289 10.6151
R5117 vdd.n1293 vdd.n1290 10.6151
R5118 vdd.n1294 vdd.n1293 10.6151
R5119 vdd.n1297 vdd.n1294 10.6151
R5120 vdd.n1298 vdd.n1297 10.6151
R5121 vdd.n1301 vdd.n1298 10.6151
R5122 vdd.n1302 vdd.n1301 10.6151
R5123 vdd.n1305 vdd.n1302 10.6151
R5124 vdd.n1306 vdd.n1305 10.6151
R5125 vdd.n1309 vdd.n1306 10.6151
R5126 vdd.n1310 vdd.n1309 10.6151
R5127 vdd.n1313 vdd.n1310 10.6151
R5128 vdd.n1515 vdd.n1313 10.6151
R5129 vdd.n1515 vdd.n1514 10.6151
R5130 vdd.n1514 vdd.n1512 10.6151
R5131 vdd.n1512 vdd.n1509 10.6151
R5132 vdd.n1509 vdd.n1508 10.6151
R5133 vdd.n1508 vdd.n1505 10.6151
R5134 vdd.n1505 vdd.n1504 10.6151
R5135 vdd.n1504 vdd.n1501 10.6151
R5136 vdd.n1501 vdd.n1500 10.6151
R5137 vdd.n1500 vdd.n1497 10.6151
R5138 vdd.n1497 vdd.n1496 10.6151
R5139 vdd.n1496 vdd.n1493 10.6151
R5140 vdd.n1493 vdd.n1492 10.6151
R5141 vdd.n1492 vdd.n1489 10.6151
R5142 vdd.n1489 vdd.n1488 10.6151
R5143 vdd.n1485 vdd.n1484 10.6151
R5144 vdd.n1484 vdd.n1482 10.6151
R5145 vdd.n2306 vdd.t99 10.5435
R5146 vdd.n656 vdd.t76 10.5435
R5147 vdd.n316 vdd.n298 10.4732
R5148 vdd.n257 vdd.n239 10.4732
R5149 vdd.n214 vdd.n196 10.4732
R5150 vdd.n155 vdd.n137 10.4732
R5151 vdd.n113 vdd.n95 10.4732
R5152 vdd.n54 vdd.n36 10.4732
R5153 vdd.n2190 vdd.n2172 10.4732
R5154 vdd.n2249 vdd.n2231 10.4732
R5155 vdd.n2088 vdd.n2070 10.4732
R5156 vdd.n2147 vdd.n2129 10.4732
R5157 vdd.n1987 vdd.n1969 10.4732
R5158 vdd.n2046 vdd.n2028 10.4732
R5159 vdd.t53 vdd.n2280 10.3167
R5160 vdd.n3572 vdd.t27 10.3167
R5161 vdd.n1957 vdd.t43 10.09
R5162 vdd.n3666 vdd.t120 10.09
R5163 vdd.n2475 vdd.n2474 9.98956
R5164 vdd.n3488 vdd.n731 9.98956
R5165 vdd.n3365 vdd.n3364 9.98956
R5166 vdd.n2367 vdd.n1515 9.98956
R5167 vdd.t51 vdd.n1610 9.86327
R5168 vdd.n3657 vdd.t69 9.86327
R5169 vdd.n2712 vdd.t189 9.7499
R5170 vdd.t174 vdd.n957 9.7499
R5171 vdd.n315 vdd.n300 9.69747
R5172 vdd.n256 vdd.n241 9.69747
R5173 vdd.n213 vdd.n198 9.69747
R5174 vdd.n154 vdd.n139 9.69747
R5175 vdd.n112 vdd.n97 9.69747
R5176 vdd.n53 vdd.n38 9.69747
R5177 vdd.n2189 vdd.n2174 9.69747
R5178 vdd.n2248 vdd.n2233 9.69747
R5179 vdd.n2087 vdd.n2072 9.69747
R5180 vdd.n2146 vdd.n2131 9.69747
R5181 vdd.n1986 vdd.n1971 9.69747
R5182 vdd.n2045 vdd.n2030 9.69747
R5183 vdd.n1916 vdd.t85 9.63654
R5184 vdd.n3603 vdd.t37 9.63654
R5185 vdd.n331 vdd.n330 9.45567
R5186 vdd.n272 vdd.n271 9.45567
R5187 vdd.n229 vdd.n228 9.45567
R5188 vdd.n170 vdd.n169 9.45567
R5189 vdd.n128 vdd.n127 9.45567
R5190 vdd.n69 vdd.n68 9.45567
R5191 vdd.n2205 vdd.n2204 9.45567
R5192 vdd.n2264 vdd.n2263 9.45567
R5193 vdd.n2103 vdd.n2102 9.45567
R5194 vdd.n2162 vdd.n2161 9.45567
R5195 vdd.n2002 vdd.n2001 9.45567
R5196 vdd.n2061 vdd.n2060 9.45567
R5197 vdd.n1890 vdd.t21 9.40981
R5198 vdd.n3635 vdd.t23 9.40981
R5199 vdd.n2437 vdd.n1207 9.3005
R5200 vdd.n2436 vdd.n2435 9.3005
R5201 vdd.n1213 vdd.n1212 9.3005
R5202 vdd.n2430 vdd.n1217 9.3005
R5203 vdd.n2429 vdd.n1218 9.3005
R5204 vdd.n2428 vdd.n1219 9.3005
R5205 vdd.n1223 vdd.n1220 9.3005
R5206 vdd.n2423 vdd.n1224 9.3005
R5207 vdd.n2422 vdd.n1225 9.3005
R5208 vdd.n2421 vdd.n1226 9.3005
R5209 vdd.n1230 vdd.n1227 9.3005
R5210 vdd.n2416 vdd.n1231 9.3005
R5211 vdd.n2415 vdd.n1232 9.3005
R5212 vdd.n2414 vdd.n1233 9.3005
R5213 vdd.n1237 vdd.n1234 9.3005
R5214 vdd.n2409 vdd.n1238 9.3005
R5215 vdd.n2408 vdd.n1239 9.3005
R5216 vdd.n2407 vdd.n1240 9.3005
R5217 vdd.n1244 vdd.n1241 9.3005
R5218 vdd.n2402 vdd.n1245 9.3005
R5219 vdd.n2401 vdd.n1246 9.3005
R5220 vdd.n2400 vdd.n2399 9.3005
R5221 vdd.n2398 vdd.n1247 9.3005
R5222 vdd.n2397 vdd.n2396 9.3005
R5223 vdd.n1253 vdd.n1252 9.3005
R5224 vdd.n2391 vdd.n1257 9.3005
R5225 vdd.n2390 vdd.n1258 9.3005
R5226 vdd.n2389 vdd.n1259 9.3005
R5227 vdd.n1263 vdd.n1260 9.3005
R5228 vdd.n2384 vdd.n1264 9.3005
R5229 vdd.n2383 vdd.n1265 9.3005
R5230 vdd.n2382 vdd.n1266 9.3005
R5231 vdd.n1270 vdd.n1267 9.3005
R5232 vdd.n2377 vdd.n1271 9.3005
R5233 vdd.n2376 vdd.n1272 9.3005
R5234 vdd.n2375 vdd.n1273 9.3005
R5235 vdd.n1277 vdd.n1274 9.3005
R5236 vdd.n2370 vdd.n1278 9.3005
R5237 vdd.n2439 vdd.n2438 9.3005
R5238 vdd.n2461 vdd.n1178 9.3005
R5239 vdd.n2460 vdd.n1186 9.3005
R5240 vdd.n1190 vdd.n1187 9.3005
R5241 vdd.n2455 vdd.n1191 9.3005
R5242 vdd.n2454 vdd.n1192 9.3005
R5243 vdd.n2453 vdd.n1193 9.3005
R5244 vdd.n1197 vdd.n1194 9.3005
R5245 vdd.n2448 vdd.n1198 9.3005
R5246 vdd.n2447 vdd.n1199 9.3005
R5247 vdd.n2446 vdd.n1200 9.3005
R5248 vdd.n1204 vdd.n1201 9.3005
R5249 vdd.n2441 vdd.n1205 9.3005
R5250 vdd.n2440 vdd.n1206 9.3005
R5251 vdd.n2473 vdd.n2472 9.3005
R5252 vdd.n1182 vdd.n1181 9.3005
R5253 vdd.n2270 vdd.n2269 9.3005
R5254 vdd.n1579 vdd.n1578 9.3005
R5255 vdd.n2284 vdd.n2283 9.3005
R5256 vdd.n2285 vdd.n1577 9.3005
R5257 vdd.n2287 vdd.n2286 9.3005
R5258 vdd.n1568 vdd.n1567 9.3005
R5259 vdd.n2301 vdd.n2300 9.3005
R5260 vdd.n2302 vdd.n1566 9.3005
R5261 vdd.n2304 vdd.n2303 9.3005
R5262 vdd.n1557 vdd.n1556 9.3005
R5263 vdd.n2317 vdd.n2316 9.3005
R5264 vdd.n2318 vdd.n1555 9.3005
R5265 vdd.n2320 vdd.n2319 9.3005
R5266 vdd.n1545 vdd.n1544 9.3005
R5267 vdd.n2334 vdd.n2333 9.3005
R5268 vdd.n2335 vdd.n1543 9.3005
R5269 vdd.n2337 vdd.n2336 9.3005
R5270 vdd.n1533 vdd.n1532 9.3005
R5271 vdd.n2353 vdd.n2352 9.3005
R5272 vdd.n2354 vdd.n1531 9.3005
R5273 vdd.n2356 vdd.n2355 9.3005
R5274 vdd.n307 vdd.n306 9.3005
R5275 vdd.n302 vdd.n301 9.3005
R5276 vdd.n313 vdd.n312 9.3005
R5277 vdd.n315 vdd.n314 9.3005
R5278 vdd.n298 vdd.n297 9.3005
R5279 vdd.n321 vdd.n320 9.3005
R5280 vdd.n323 vdd.n322 9.3005
R5281 vdd.n295 vdd.n292 9.3005
R5282 vdd.n330 vdd.n329 9.3005
R5283 vdd.n248 vdd.n247 9.3005
R5284 vdd.n243 vdd.n242 9.3005
R5285 vdd.n254 vdd.n253 9.3005
R5286 vdd.n256 vdd.n255 9.3005
R5287 vdd.n239 vdd.n238 9.3005
R5288 vdd.n262 vdd.n261 9.3005
R5289 vdd.n264 vdd.n263 9.3005
R5290 vdd.n236 vdd.n233 9.3005
R5291 vdd.n271 vdd.n270 9.3005
R5292 vdd.n205 vdd.n204 9.3005
R5293 vdd.n200 vdd.n199 9.3005
R5294 vdd.n211 vdd.n210 9.3005
R5295 vdd.n213 vdd.n212 9.3005
R5296 vdd.n196 vdd.n195 9.3005
R5297 vdd.n219 vdd.n218 9.3005
R5298 vdd.n221 vdd.n220 9.3005
R5299 vdd.n193 vdd.n190 9.3005
R5300 vdd.n228 vdd.n227 9.3005
R5301 vdd.n146 vdd.n145 9.3005
R5302 vdd.n141 vdd.n140 9.3005
R5303 vdd.n152 vdd.n151 9.3005
R5304 vdd.n154 vdd.n153 9.3005
R5305 vdd.n137 vdd.n136 9.3005
R5306 vdd.n160 vdd.n159 9.3005
R5307 vdd.n162 vdd.n161 9.3005
R5308 vdd.n134 vdd.n131 9.3005
R5309 vdd.n169 vdd.n168 9.3005
R5310 vdd.n104 vdd.n103 9.3005
R5311 vdd.n99 vdd.n98 9.3005
R5312 vdd.n110 vdd.n109 9.3005
R5313 vdd.n112 vdd.n111 9.3005
R5314 vdd.n95 vdd.n94 9.3005
R5315 vdd.n118 vdd.n117 9.3005
R5316 vdd.n120 vdd.n119 9.3005
R5317 vdd.n92 vdd.n89 9.3005
R5318 vdd.n127 vdd.n126 9.3005
R5319 vdd.n45 vdd.n44 9.3005
R5320 vdd.n40 vdd.n39 9.3005
R5321 vdd.n51 vdd.n50 9.3005
R5322 vdd.n53 vdd.n52 9.3005
R5323 vdd.n36 vdd.n35 9.3005
R5324 vdd.n59 vdd.n58 9.3005
R5325 vdd.n61 vdd.n60 9.3005
R5326 vdd.n33 vdd.n30 9.3005
R5327 vdd.n68 vdd.n67 9.3005
R5328 vdd.n3410 vdd.n3409 9.3005
R5329 vdd.n3413 vdd.n766 9.3005
R5330 vdd.n3414 vdd.n765 9.3005
R5331 vdd.n3417 vdd.n764 9.3005
R5332 vdd.n3418 vdd.n763 9.3005
R5333 vdd.n3421 vdd.n762 9.3005
R5334 vdd.n3422 vdd.n761 9.3005
R5335 vdd.n3425 vdd.n760 9.3005
R5336 vdd.n3426 vdd.n759 9.3005
R5337 vdd.n3429 vdd.n758 9.3005
R5338 vdd.n3430 vdd.n757 9.3005
R5339 vdd.n3433 vdd.n756 9.3005
R5340 vdd.n3434 vdd.n755 9.3005
R5341 vdd.n3437 vdd.n754 9.3005
R5342 vdd.n3438 vdd.n753 9.3005
R5343 vdd.n3441 vdd.n752 9.3005
R5344 vdd.n3442 vdd.n751 9.3005
R5345 vdd.n3445 vdd.n750 9.3005
R5346 vdd.n3446 vdd.n749 9.3005
R5347 vdd.n3449 vdd.n748 9.3005
R5348 vdd.n3453 vdd.n3452 9.3005
R5349 vdd.n3454 vdd.n747 9.3005
R5350 vdd.n3458 vdd.n3455 9.3005
R5351 vdd.n3461 vdd.n746 9.3005
R5352 vdd.n3462 vdd.n745 9.3005
R5353 vdd.n3465 vdd.n744 9.3005
R5354 vdd.n3466 vdd.n743 9.3005
R5355 vdd.n3469 vdd.n742 9.3005
R5356 vdd.n3470 vdd.n741 9.3005
R5357 vdd.n3473 vdd.n740 9.3005
R5358 vdd.n3474 vdd.n739 9.3005
R5359 vdd.n3477 vdd.n738 9.3005
R5360 vdd.n3478 vdd.n737 9.3005
R5361 vdd.n3481 vdd.n736 9.3005
R5362 vdd.n3482 vdd.n735 9.3005
R5363 vdd.n3485 vdd.n730 9.3005
R5364 vdd.n3491 vdd.n727 9.3005
R5365 vdd.n3492 vdd.n726 9.3005
R5366 vdd.n3506 vdd.n3505 9.3005
R5367 vdd.n3507 vdd.n681 9.3005
R5368 vdd.n3509 vdd.n3508 9.3005
R5369 vdd.n671 vdd.n670 9.3005
R5370 vdd.n3523 vdd.n3522 9.3005
R5371 vdd.n3524 vdd.n669 9.3005
R5372 vdd.n3526 vdd.n3525 9.3005
R5373 vdd.n660 vdd.n659 9.3005
R5374 vdd.n3539 vdd.n3538 9.3005
R5375 vdd.n3540 vdd.n658 9.3005
R5376 vdd.n3542 vdd.n3541 9.3005
R5377 vdd.n648 vdd.n647 9.3005
R5378 vdd.n3556 vdd.n3555 9.3005
R5379 vdd.n3557 vdd.n646 9.3005
R5380 vdd.n3559 vdd.n3558 9.3005
R5381 vdd.n637 vdd.n636 9.3005
R5382 vdd.n3575 vdd.n3574 9.3005
R5383 vdd.n3576 vdd.n635 9.3005
R5384 vdd.n3578 vdd.n3577 9.3005
R5385 vdd.n336 vdd.n334 9.3005
R5386 vdd.n683 vdd.n682 9.3005
R5387 vdd.n3670 vdd.n3669 9.3005
R5388 vdd.n337 vdd.n335 9.3005
R5389 vdd.n3663 vdd.n346 9.3005
R5390 vdd.n3662 vdd.n347 9.3005
R5391 vdd.n3661 vdd.n348 9.3005
R5392 vdd.n355 vdd.n349 9.3005
R5393 vdd.n3655 vdd.n356 9.3005
R5394 vdd.n3654 vdd.n357 9.3005
R5395 vdd.n3653 vdd.n358 9.3005
R5396 vdd.n366 vdd.n359 9.3005
R5397 vdd.n3647 vdd.n367 9.3005
R5398 vdd.n3646 vdd.n368 9.3005
R5399 vdd.n3645 vdd.n369 9.3005
R5400 vdd.n377 vdd.n370 9.3005
R5401 vdd.n3639 vdd.n378 9.3005
R5402 vdd.n3638 vdd.n379 9.3005
R5403 vdd.n3637 vdd.n380 9.3005
R5404 vdd.n388 vdd.n381 9.3005
R5405 vdd.n3631 vdd.n389 9.3005
R5406 vdd.n3630 vdd.n390 9.3005
R5407 vdd.n3629 vdd.n391 9.3005
R5408 vdd.n466 vdd.n463 9.3005
R5409 vdd.n470 vdd.n469 9.3005
R5410 vdd.n471 vdd.n462 9.3005
R5411 vdd.n475 vdd.n472 9.3005
R5412 vdd.n476 vdd.n461 9.3005
R5413 vdd.n480 vdd.n479 9.3005
R5414 vdd.n481 vdd.n460 9.3005
R5415 vdd.n485 vdd.n482 9.3005
R5416 vdd.n486 vdd.n459 9.3005
R5417 vdd.n490 vdd.n489 9.3005
R5418 vdd.n491 vdd.n458 9.3005
R5419 vdd.n495 vdd.n492 9.3005
R5420 vdd.n496 vdd.n457 9.3005
R5421 vdd.n500 vdd.n499 9.3005
R5422 vdd.n501 vdd.n456 9.3005
R5423 vdd.n505 vdd.n502 9.3005
R5424 vdd.n506 vdd.n455 9.3005
R5425 vdd.n510 vdd.n509 9.3005
R5426 vdd.n511 vdd.n454 9.3005
R5427 vdd.n515 vdd.n512 9.3005
R5428 vdd.n516 vdd.n451 9.3005
R5429 vdd.n520 vdd.n519 9.3005
R5430 vdd.n521 vdd.n450 9.3005
R5431 vdd.n525 vdd.n522 9.3005
R5432 vdd.n526 vdd.n449 9.3005
R5433 vdd.n530 vdd.n529 9.3005
R5434 vdd.n531 vdd.n448 9.3005
R5435 vdd.n535 vdd.n532 9.3005
R5436 vdd.n536 vdd.n447 9.3005
R5437 vdd.n540 vdd.n539 9.3005
R5438 vdd.n541 vdd.n446 9.3005
R5439 vdd.n545 vdd.n542 9.3005
R5440 vdd.n546 vdd.n445 9.3005
R5441 vdd.n550 vdd.n549 9.3005
R5442 vdd.n551 vdd.n444 9.3005
R5443 vdd.n555 vdd.n552 9.3005
R5444 vdd.n556 vdd.n443 9.3005
R5445 vdd.n560 vdd.n559 9.3005
R5446 vdd.n561 vdd.n442 9.3005
R5447 vdd.n565 vdd.n562 9.3005
R5448 vdd.n566 vdd.n439 9.3005
R5449 vdd.n570 vdd.n569 9.3005
R5450 vdd.n571 vdd.n438 9.3005
R5451 vdd.n575 vdd.n572 9.3005
R5452 vdd.n576 vdd.n437 9.3005
R5453 vdd.n580 vdd.n579 9.3005
R5454 vdd.n581 vdd.n436 9.3005
R5455 vdd.n585 vdd.n582 9.3005
R5456 vdd.n586 vdd.n435 9.3005
R5457 vdd.n590 vdd.n589 9.3005
R5458 vdd.n591 vdd.n434 9.3005
R5459 vdd.n595 vdd.n592 9.3005
R5460 vdd.n596 vdd.n433 9.3005
R5461 vdd.n600 vdd.n599 9.3005
R5462 vdd.n601 vdd.n432 9.3005
R5463 vdd.n605 vdd.n602 9.3005
R5464 vdd.n606 vdd.n431 9.3005
R5465 vdd.n610 vdd.n609 9.3005
R5466 vdd.n611 vdd.n430 9.3005
R5467 vdd.n615 vdd.n612 9.3005
R5468 vdd.n617 vdd.n429 9.3005
R5469 vdd.n619 vdd.n618 9.3005
R5470 vdd.n3623 vdd.n3622 9.3005
R5471 vdd.n465 vdd.n464 9.3005
R5472 vdd.n3501 vdd.n3500 9.3005
R5473 vdd.n676 vdd.n675 9.3005
R5474 vdd.n3514 vdd.n3513 9.3005
R5475 vdd.n3515 vdd.n674 9.3005
R5476 vdd.n3517 vdd.n3516 9.3005
R5477 vdd.n666 vdd.n665 9.3005
R5478 vdd.n3531 vdd.n3530 9.3005
R5479 vdd.n3532 vdd.n664 9.3005
R5480 vdd.n3534 vdd.n3533 9.3005
R5481 vdd.n653 vdd.n652 9.3005
R5482 vdd.n3547 vdd.n3546 9.3005
R5483 vdd.n3548 vdd.n651 9.3005
R5484 vdd.n3550 vdd.n3549 9.3005
R5485 vdd.n642 vdd.n641 9.3005
R5486 vdd.n3564 vdd.n3563 9.3005
R5487 vdd.n3565 vdd.n640 9.3005
R5488 vdd.n3570 vdd.n3566 9.3005
R5489 vdd.n3569 vdd.n3568 9.3005
R5490 vdd.n3567 vdd.n631 9.3005
R5491 vdd.n3583 vdd.n630 9.3005
R5492 vdd.n3585 vdd.n3584 9.3005
R5493 vdd.n3586 vdd.n629 9.3005
R5494 vdd.n3588 vdd.n3587 9.3005
R5495 vdd.n3590 vdd.n628 9.3005
R5496 vdd.n3592 vdd.n3591 9.3005
R5497 vdd.n3593 vdd.n627 9.3005
R5498 vdd.n3595 vdd.n3594 9.3005
R5499 vdd.n3597 vdd.n626 9.3005
R5500 vdd.n3599 vdd.n3598 9.3005
R5501 vdd.n3600 vdd.n625 9.3005
R5502 vdd.n3602 vdd.n3601 9.3005
R5503 vdd.n3605 vdd.n624 9.3005
R5504 vdd.n3607 vdd.n3606 9.3005
R5505 vdd.n3608 vdd.n623 9.3005
R5506 vdd.n3610 vdd.n3609 9.3005
R5507 vdd.n3612 vdd.n622 9.3005
R5508 vdd.n3614 vdd.n3613 9.3005
R5509 vdd.n3615 vdd.n621 9.3005
R5510 vdd.n3617 vdd.n3616 9.3005
R5511 vdd.n3619 vdd.n620 9.3005
R5512 vdd.n3621 vdd.n3620 9.3005
R5513 vdd.n3499 vdd.n686 9.3005
R5514 vdd.n3498 vdd.n3497 9.3005
R5515 vdd.n3367 vdd.n687 9.3005
R5516 vdd.n3376 vdd.n783 9.3005
R5517 vdd.n3379 vdd.n782 9.3005
R5518 vdd.n3380 vdd.n781 9.3005
R5519 vdd.n3383 vdd.n780 9.3005
R5520 vdd.n3384 vdd.n779 9.3005
R5521 vdd.n3387 vdd.n778 9.3005
R5522 vdd.n3388 vdd.n777 9.3005
R5523 vdd.n3391 vdd.n776 9.3005
R5524 vdd.n3392 vdd.n775 9.3005
R5525 vdd.n3395 vdd.n774 9.3005
R5526 vdd.n3396 vdd.n773 9.3005
R5527 vdd.n3399 vdd.n772 9.3005
R5528 vdd.n3400 vdd.n771 9.3005
R5529 vdd.n3403 vdd.n770 9.3005
R5530 vdd.n3407 vdd.n3406 9.3005
R5531 vdd.n3408 vdd.n767 9.3005
R5532 vdd.n2366 vdd.n2365 9.3005
R5533 vdd.n2361 vdd.n1517 9.3005
R5534 vdd.n1885 vdd.n1884 9.3005
R5535 vdd.n1886 vdd.n1640 9.3005
R5536 vdd.n1888 vdd.n1887 9.3005
R5537 vdd.n1630 vdd.n1629 9.3005
R5538 vdd.n1902 vdd.n1901 9.3005
R5539 vdd.n1903 vdd.n1628 9.3005
R5540 vdd.n1905 vdd.n1904 9.3005
R5541 vdd.n1620 vdd.n1619 9.3005
R5542 vdd.n1919 vdd.n1918 9.3005
R5543 vdd.n1920 vdd.n1618 9.3005
R5544 vdd.n1922 vdd.n1921 9.3005
R5545 vdd.n1607 vdd.n1606 9.3005
R5546 vdd.n1935 vdd.n1934 9.3005
R5547 vdd.n1936 vdd.n1605 9.3005
R5548 vdd.n1938 vdd.n1937 9.3005
R5549 vdd.n1596 vdd.n1595 9.3005
R5550 vdd.n1952 vdd.n1951 9.3005
R5551 vdd.n1953 vdd.n1594 9.3005
R5552 vdd.n1955 vdd.n1954 9.3005
R5553 vdd.n1585 vdd.n1584 9.3005
R5554 vdd.n2275 vdd.n2274 9.3005
R5555 vdd.n2276 vdd.n1583 9.3005
R5556 vdd.n2278 vdd.n2277 9.3005
R5557 vdd.n1573 vdd.n1572 9.3005
R5558 vdd.n2292 vdd.n2291 9.3005
R5559 vdd.n2293 vdd.n1571 9.3005
R5560 vdd.n2295 vdd.n2294 9.3005
R5561 vdd.n1563 vdd.n1562 9.3005
R5562 vdd.n2309 vdd.n2308 9.3005
R5563 vdd.n2310 vdd.n1561 9.3005
R5564 vdd.n2312 vdd.n2311 9.3005
R5565 vdd.n1550 vdd.n1549 9.3005
R5566 vdd.n2325 vdd.n2324 9.3005
R5567 vdd.n2326 vdd.n1548 9.3005
R5568 vdd.n2328 vdd.n2327 9.3005
R5569 vdd.n1540 vdd.n1539 9.3005
R5570 vdd.n2342 vdd.n2341 9.3005
R5571 vdd.n2343 vdd.n1537 9.3005
R5572 vdd.n2347 vdd.n2346 9.3005
R5573 vdd.n2345 vdd.n1538 9.3005
R5574 vdd.n2344 vdd.n1528 9.3005
R5575 vdd.n1642 vdd.n1641 9.3005
R5576 vdd.n1778 vdd.n1777 9.3005
R5577 vdd.n1779 vdd.n1768 9.3005
R5578 vdd.n1781 vdd.n1780 9.3005
R5579 vdd.n1782 vdd.n1767 9.3005
R5580 vdd.n1784 vdd.n1783 9.3005
R5581 vdd.n1785 vdd.n1762 9.3005
R5582 vdd.n1787 vdd.n1786 9.3005
R5583 vdd.n1788 vdd.n1761 9.3005
R5584 vdd.n1790 vdd.n1789 9.3005
R5585 vdd.n1791 vdd.n1756 9.3005
R5586 vdd.n1793 vdd.n1792 9.3005
R5587 vdd.n1794 vdd.n1755 9.3005
R5588 vdd.n1796 vdd.n1795 9.3005
R5589 vdd.n1797 vdd.n1750 9.3005
R5590 vdd.n1799 vdd.n1798 9.3005
R5591 vdd.n1800 vdd.n1749 9.3005
R5592 vdd.n1802 vdd.n1801 9.3005
R5593 vdd.n1803 vdd.n1744 9.3005
R5594 vdd.n1805 vdd.n1804 9.3005
R5595 vdd.n1806 vdd.n1743 9.3005
R5596 vdd.n1808 vdd.n1807 9.3005
R5597 vdd.n1812 vdd.n1739 9.3005
R5598 vdd.n1814 vdd.n1813 9.3005
R5599 vdd.n1815 vdd.n1738 9.3005
R5600 vdd.n1817 vdd.n1816 9.3005
R5601 vdd.n1818 vdd.n1733 9.3005
R5602 vdd.n1820 vdd.n1819 9.3005
R5603 vdd.n1821 vdd.n1732 9.3005
R5604 vdd.n1823 vdd.n1822 9.3005
R5605 vdd.n1824 vdd.n1727 9.3005
R5606 vdd.n1826 vdd.n1825 9.3005
R5607 vdd.n1827 vdd.n1726 9.3005
R5608 vdd.n1829 vdd.n1828 9.3005
R5609 vdd.n1830 vdd.n1721 9.3005
R5610 vdd.n1832 vdd.n1831 9.3005
R5611 vdd.n1833 vdd.n1720 9.3005
R5612 vdd.n1835 vdd.n1834 9.3005
R5613 vdd.n1836 vdd.n1715 9.3005
R5614 vdd.n1838 vdd.n1837 9.3005
R5615 vdd.n1839 vdd.n1714 9.3005
R5616 vdd.n1841 vdd.n1840 9.3005
R5617 vdd.n1842 vdd.n1709 9.3005
R5618 vdd.n1844 vdd.n1843 9.3005
R5619 vdd.n1845 vdd.n1708 9.3005
R5620 vdd.n1847 vdd.n1846 9.3005
R5621 vdd.n1848 vdd.n1701 9.3005
R5622 vdd.n1850 vdd.n1849 9.3005
R5623 vdd.n1851 vdd.n1700 9.3005
R5624 vdd.n1853 vdd.n1852 9.3005
R5625 vdd.n1854 vdd.n1695 9.3005
R5626 vdd.n1856 vdd.n1855 9.3005
R5627 vdd.n1857 vdd.n1694 9.3005
R5628 vdd.n1859 vdd.n1858 9.3005
R5629 vdd.n1860 vdd.n1689 9.3005
R5630 vdd.n1862 vdd.n1861 9.3005
R5631 vdd.n1863 vdd.n1688 9.3005
R5632 vdd.n1865 vdd.n1864 9.3005
R5633 vdd.n1866 vdd.n1683 9.3005
R5634 vdd.n1868 vdd.n1867 9.3005
R5635 vdd.n1869 vdd.n1682 9.3005
R5636 vdd.n1871 vdd.n1870 9.3005
R5637 vdd.n1647 vdd.n1646 9.3005
R5638 vdd.n1877 vdd.n1876 9.3005
R5639 vdd.n1776 vdd.n1775 9.3005
R5640 vdd.n1880 vdd.n1879 9.3005
R5641 vdd.n1636 vdd.n1635 9.3005
R5642 vdd.n1894 vdd.n1893 9.3005
R5643 vdd.n1895 vdd.n1634 9.3005
R5644 vdd.n1897 vdd.n1896 9.3005
R5645 vdd.n1625 vdd.n1624 9.3005
R5646 vdd.n1911 vdd.n1910 9.3005
R5647 vdd.n1912 vdd.n1623 9.3005
R5648 vdd.n1914 vdd.n1913 9.3005
R5649 vdd.n1614 vdd.n1613 9.3005
R5650 vdd.n1927 vdd.n1926 9.3005
R5651 vdd.n1928 vdd.n1612 9.3005
R5652 vdd.n1930 vdd.n1929 9.3005
R5653 vdd.n1602 vdd.n1601 9.3005
R5654 vdd.n1944 vdd.n1943 9.3005
R5655 vdd.n1945 vdd.n1600 9.3005
R5656 vdd.n1947 vdd.n1946 9.3005
R5657 vdd.n1591 vdd.n1590 9.3005
R5658 vdd.n1960 vdd.n1959 9.3005
R5659 vdd.n1961 vdd.n1589 9.3005
R5660 vdd.n1878 vdd.n1645 9.3005
R5661 vdd.n2181 vdd.n2180 9.3005
R5662 vdd.n2176 vdd.n2175 9.3005
R5663 vdd.n2187 vdd.n2186 9.3005
R5664 vdd.n2189 vdd.n2188 9.3005
R5665 vdd.n2172 vdd.n2171 9.3005
R5666 vdd.n2195 vdd.n2194 9.3005
R5667 vdd.n2197 vdd.n2196 9.3005
R5668 vdd.n2169 vdd.n2166 9.3005
R5669 vdd.n2204 vdd.n2203 9.3005
R5670 vdd.n2240 vdd.n2239 9.3005
R5671 vdd.n2235 vdd.n2234 9.3005
R5672 vdd.n2246 vdd.n2245 9.3005
R5673 vdd.n2248 vdd.n2247 9.3005
R5674 vdd.n2231 vdd.n2230 9.3005
R5675 vdd.n2254 vdd.n2253 9.3005
R5676 vdd.n2256 vdd.n2255 9.3005
R5677 vdd.n2228 vdd.n2225 9.3005
R5678 vdd.n2263 vdd.n2262 9.3005
R5679 vdd.n2079 vdd.n2078 9.3005
R5680 vdd.n2074 vdd.n2073 9.3005
R5681 vdd.n2085 vdd.n2084 9.3005
R5682 vdd.n2087 vdd.n2086 9.3005
R5683 vdd.n2070 vdd.n2069 9.3005
R5684 vdd.n2093 vdd.n2092 9.3005
R5685 vdd.n2095 vdd.n2094 9.3005
R5686 vdd.n2067 vdd.n2064 9.3005
R5687 vdd.n2102 vdd.n2101 9.3005
R5688 vdd.n2138 vdd.n2137 9.3005
R5689 vdd.n2133 vdd.n2132 9.3005
R5690 vdd.n2144 vdd.n2143 9.3005
R5691 vdd.n2146 vdd.n2145 9.3005
R5692 vdd.n2129 vdd.n2128 9.3005
R5693 vdd.n2152 vdd.n2151 9.3005
R5694 vdd.n2154 vdd.n2153 9.3005
R5695 vdd.n2126 vdd.n2123 9.3005
R5696 vdd.n2161 vdd.n2160 9.3005
R5697 vdd.n1978 vdd.n1977 9.3005
R5698 vdd.n1973 vdd.n1972 9.3005
R5699 vdd.n1984 vdd.n1983 9.3005
R5700 vdd.n1986 vdd.n1985 9.3005
R5701 vdd.n1969 vdd.n1968 9.3005
R5702 vdd.n1992 vdd.n1991 9.3005
R5703 vdd.n1994 vdd.n1993 9.3005
R5704 vdd.n1966 vdd.n1963 9.3005
R5705 vdd.n2001 vdd.n2000 9.3005
R5706 vdd.n2037 vdd.n2036 9.3005
R5707 vdd.n2032 vdd.n2031 9.3005
R5708 vdd.n2043 vdd.n2042 9.3005
R5709 vdd.n2045 vdd.n2044 9.3005
R5710 vdd.n2028 vdd.n2027 9.3005
R5711 vdd.n2051 vdd.n2050 9.3005
R5712 vdd.n2053 vdd.n2052 9.3005
R5713 vdd.n2025 vdd.n2022 9.3005
R5714 vdd.n2060 vdd.n2059 9.3005
R5715 vdd.n1916 vdd.t67 9.18308
R5716 vdd.n3603 vdd.t72 9.18308
R5717 vdd.n1610 vdd.t114 8.95635
R5718 vdd.n2358 vdd.t241 8.95635
R5719 vdd.n723 vdd.t258 8.95635
R5720 vdd.t104 vdd.n3657 8.95635
R5721 vdd.n312 vdd.n311 8.92171
R5722 vdd.n253 vdd.n252 8.92171
R5723 vdd.n210 vdd.n209 8.92171
R5724 vdd.n151 vdd.n150 8.92171
R5725 vdd.n109 vdd.n108 8.92171
R5726 vdd.n50 vdd.n49 8.92171
R5727 vdd.n2186 vdd.n2185 8.92171
R5728 vdd.n2245 vdd.n2244 8.92171
R5729 vdd.n2084 vdd.n2083 8.92171
R5730 vdd.n2143 vdd.n2142 8.92171
R5731 vdd.n1983 vdd.n1982 8.92171
R5732 vdd.n2042 vdd.n2041 8.92171
R5733 vdd.n231 vdd.n129 8.81535
R5734 vdd.n2164 vdd.n2062 8.81535
R5735 vdd.n1957 vdd.t74 8.72962
R5736 vdd.t29 vdd.n3666 8.72962
R5737 vdd.n2280 vdd.t11 8.50289
R5738 vdd.n3572 vdd.t55 8.50289
R5739 vdd.n28 vdd.n14 8.42249
R5740 vdd.n2306 vdd.t0 8.27616
R5741 vdd.t2 vdd.n656 8.27616
R5742 vdd.n3672 vdd.n3671 8.16225
R5743 vdd.n2268 vdd.n2267 8.16225
R5744 vdd.n308 vdd.n302 8.14595
R5745 vdd.n249 vdd.n243 8.14595
R5746 vdd.n206 vdd.n200 8.14595
R5747 vdd.n147 vdd.n141 8.14595
R5748 vdd.n105 vdd.n99 8.14595
R5749 vdd.n46 vdd.n40 8.14595
R5750 vdd.n2182 vdd.n2176 8.14595
R5751 vdd.n2241 vdd.n2235 8.14595
R5752 vdd.n2080 vdd.n2074 8.14595
R5753 vdd.n2139 vdd.n2133 8.14595
R5754 vdd.n1979 vdd.n1973 8.14595
R5755 vdd.n2038 vdd.n2032 8.14595
R5756 vdd.n1553 vdd.t204 8.04943
R5757 vdd.n3528 vdd.t116 8.04943
R5758 vdd.n2513 vdd.n1134 7.70933
R5759 vdd.n2513 vdd.n1137 7.70933
R5760 vdd.n2519 vdd.n1123 7.70933
R5761 vdd.n2525 vdd.n1123 7.70933
R5762 vdd.n2525 vdd.n1116 7.70933
R5763 vdd.n2531 vdd.n1116 7.70933
R5764 vdd.n2531 vdd.n1119 7.70933
R5765 vdd.n2537 vdd.n1112 7.70933
R5766 vdd.n2543 vdd.n1106 7.70933
R5767 vdd.n2549 vdd.n1093 7.70933
R5768 vdd.n2555 vdd.n1093 7.70933
R5769 vdd.n2561 vdd.n1087 7.70933
R5770 vdd.n2567 vdd.n1080 7.70933
R5771 vdd.n2567 vdd.n1083 7.70933
R5772 vdd.n2573 vdd.n1076 7.70933
R5773 vdd.n2580 vdd.n1062 7.70933
R5774 vdd.n2586 vdd.n1062 7.70933
R5775 vdd.n2592 vdd.n1056 7.70933
R5776 vdd.n2598 vdd.n1052 7.70933
R5777 vdd.n2604 vdd.n1046 7.70933
R5778 vdd.n2622 vdd.n1028 7.70933
R5779 vdd.n2622 vdd.n1021 7.70933
R5780 vdd.n2630 vdd.n1021 7.70933
R5781 vdd.n2712 vdd.n1005 7.70933
R5782 vdd.n3095 vdd.n957 7.70933
R5783 vdd.n3107 vdd.n946 7.70933
R5784 vdd.n3107 vdd.n940 7.70933
R5785 vdd.n3113 vdd.n940 7.70933
R5786 vdd.n3125 vdd.n931 7.70933
R5787 vdd.n3131 vdd.n925 7.70933
R5788 vdd.n3143 vdd.n912 7.70933
R5789 vdd.n3150 vdd.n905 7.70933
R5790 vdd.n3150 vdd.n908 7.70933
R5791 vdd.n3156 vdd.n901 7.70933
R5792 vdd.n3162 vdd.n887 7.70933
R5793 vdd.n3168 vdd.n887 7.70933
R5794 vdd.n3174 vdd.n881 7.70933
R5795 vdd.n3180 vdd.n874 7.70933
R5796 vdd.n3180 vdd.n877 7.70933
R5797 vdd.n3186 vdd.n870 7.70933
R5798 vdd.n3192 vdd.n864 7.70933
R5799 vdd.n3198 vdd.n851 7.70933
R5800 vdd.n3204 vdd.n851 7.70933
R5801 vdd.n3204 vdd.n843 7.70933
R5802 vdd.n3255 vdd.n843 7.70933
R5803 vdd.n3255 vdd.n846 7.70933
R5804 vdd.n3261 vdd.n805 7.70933
R5805 vdd.n3331 vdd.n805 7.70933
R5806 vdd.n307 vdd.n304 7.3702
R5807 vdd.n248 vdd.n245 7.3702
R5808 vdd.n205 vdd.n202 7.3702
R5809 vdd.n146 vdd.n143 7.3702
R5810 vdd.n104 vdd.n101 7.3702
R5811 vdd.n45 vdd.n42 7.3702
R5812 vdd.n2181 vdd.n2178 7.3702
R5813 vdd.n2240 vdd.n2237 7.3702
R5814 vdd.n2079 vdd.n2076 7.3702
R5815 vdd.n2138 vdd.n2135 7.3702
R5816 vdd.n1978 vdd.n1975 7.3702
R5817 vdd.n2037 vdd.n2034 7.3702
R5818 vdd.n1106 vdd.t194 7.36923
R5819 vdd.n3186 vdd.t171 7.36923
R5820 vdd.n2339 vdd.t34 7.1425
R5821 vdd.n2537 vdd.t146 7.1425
R5822 vdd.n1425 vdd.t142 7.1425
R5823 vdd.n3119 vdd.t145 7.1425
R5824 vdd.n864 vdd.t155 7.1425
R5825 vdd.n679 vdd.t13 7.1425
R5826 vdd.n1813 vdd.n1812 6.98232
R5827 vdd.n2401 vdd.n2400 6.98232
R5828 vdd.n566 vdd.n565 6.98232
R5829 vdd.n3413 vdd.n3410 6.98232
R5830 vdd.t9 vdd.n1552 6.91577
R5831 vdd.n3536 vdd.t109 6.91577
R5832 vdd.n1425 vdd.t143 6.80241
R5833 vdd.n3119 vdd.t187 6.80241
R5834 vdd.n2298 vdd.t59 6.68904
R5835 vdd.n3552 vdd.t15 6.68904
R5836 vdd.t17 vdd.n1581 6.46231
R5837 vdd.n2561 vdd.t153 6.46231
R5838 vdd.t158 vdd.n1056 6.46231
R5839 vdd.n3143 vdd.t163 6.46231
R5840 vdd.t179 vdd.n881 6.46231
R5841 vdd.n3580 vdd.t19 6.46231
R5842 vdd.n3672 vdd.n333 6.38151
R5843 vdd.n2267 vdd.n2266 6.38151
R5844 vdd.n2637 vdd.t191 6.34895
R5845 vdd.n3016 vdd.t176 6.34895
R5846 vdd.n3158 vdd.n897 6.2444
R5847 vdd.n2577 vdd.n2576 6.2444
R5848 vdd.n1949 vdd.t131 6.23558
R5849 vdd.t64 vdd.n344 6.23558
R5850 vdd.t106 vdd.n1609 6.00885
R5851 vdd.n3651 vdd.t97 6.00885
R5852 vdd.n2598 vdd.t184 5.89549
R5853 vdd.n925 vdd.t159 5.89549
R5854 vdd.n308 vdd.n307 5.81868
R5855 vdd.n249 vdd.n248 5.81868
R5856 vdd.n206 vdd.n205 5.81868
R5857 vdd.n147 vdd.n146 5.81868
R5858 vdd.n105 vdd.n104 5.81868
R5859 vdd.n46 vdd.n45 5.81868
R5860 vdd.n2182 vdd.n2181 5.81868
R5861 vdd.n2241 vdd.n2240 5.81868
R5862 vdd.n2080 vdd.n2079 5.81868
R5863 vdd.n2139 vdd.n2138 5.81868
R5864 vdd.n1979 vdd.n1978 5.81868
R5865 vdd.n2038 vdd.n2037 5.81868
R5866 vdd.n1908 vdd.t32 5.78212
R5867 vdd.n3642 vdd.t25 5.78212
R5868 vdd.n2720 vdd.n2719 5.77611
R5869 vdd.n1349 vdd.n1348 5.77611
R5870 vdd.n3028 vdd.n3027 5.77611
R5871 vdd.n3272 vdd.n3271 5.77611
R5872 vdd.n3336 vdd.n801 5.77611
R5873 vdd.n2891 vdd.n2825 5.77611
R5874 vdd.n2645 vdd.n1012 5.77611
R5875 vdd.n1485 vdd.n1317 5.77611
R5876 vdd.n1775 vdd.n1774 5.62474
R5877 vdd.n2364 vdd.n2361 5.62474
R5878 vdd.n3623 vdd.n428 5.62474
R5879 vdd.n3497 vdd.n690 5.62474
R5880 vdd.n1632 vdd.t32 5.55539
R5881 vdd.n2573 vdd.t173 5.55539
R5882 vdd.n901 vdd.t149 5.55539
R5883 vdd.t25 vdd.n3641 5.55539
R5884 vdd.n1924 vdd.t106 5.32866
R5885 vdd.t97 vdd.n3650 5.32866
R5886 vdd.n1940 vdd.t131 5.10193
R5887 vdd.n3659 vdd.t64 5.10193
R5888 vdd.n311 vdd.n302 5.04292
R5889 vdd.n252 vdd.n243 5.04292
R5890 vdd.n209 vdd.n200 5.04292
R5891 vdd.n150 vdd.n141 5.04292
R5892 vdd.n108 vdd.n99 5.04292
R5893 vdd.n49 vdd.n40 5.04292
R5894 vdd.n2185 vdd.n2176 5.04292
R5895 vdd.n2244 vdd.n2235 5.04292
R5896 vdd.n2083 vdd.n2074 5.04292
R5897 vdd.n2142 vdd.n2133 5.04292
R5898 vdd.n1982 vdd.n1973 5.04292
R5899 vdd.n2041 vdd.n2032 5.04292
R5900 vdd.n2272 vdd.t17 4.8752
R5901 vdd.t152 vdd.t164 4.8752
R5902 vdd.t195 vdd.t141 4.8752
R5903 vdd.t19 vdd.n340 4.8752
R5904 vdd.n2721 vdd.n2720 4.83952
R5905 vdd.n1348 vdd.n1347 4.83952
R5906 vdd.n3029 vdd.n3028 4.83952
R5907 vdd.n3273 vdd.n3272 4.83952
R5908 vdd.n801 vdd.n796 4.83952
R5909 vdd.n2888 vdd.n2825 4.83952
R5910 vdd.n2648 vdd.n1012 4.83952
R5911 vdd.n1488 vdd.n1317 4.83952
R5912 vdd.n1399 vdd.t161 4.76184
R5913 vdd.n3101 vdd.t147 4.76184
R5914 vdd.n2369 vdd.n2368 4.74817
R5915 vdd.n1521 vdd.n1516 4.74817
R5916 vdd.n1183 vdd.n1180 4.74817
R5917 vdd.n2462 vdd.n1179 4.74817
R5918 vdd.n2467 vdd.n1180 4.74817
R5919 vdd.n2466 vdd.n1179 4.74817
R5920 vdd.n3490 vdd.n3489 4.74817
R5921 vdd.n3487 vdd.n3486 4.74817
R5922 vdd.n3487 vdd.n732 4.74817
R5923 vdd.n3489 vdd.n729 4.74817
R5924 vdd.n3372 vdd.n784 4.74817
R5925 vdd.n3368 vdd.n3366 4.74817
R5926 vdd.n3371 vdd.n3366 4.74817
R5927 vdd.n3375 vdd.n784 4.74817
R5928 vdd.n2368 vdd.n1279 4.74817
R5929 vdd.n1518 vdd.n1516 4.74817
R5930 vdd.n333 vdd.n332 4.7074
R5931 vdd.n231 vdd.n230 4.7074
R5932 vdd.n2266 vdd.n2265 4.7074
R5933 vdd.n2164 vdd.n2163 4.7074
R5934 vdd.n1575 vdd.t59 4.64847
R5935 vdd.t154 vdd.n1087 4.64847
R5936 vdd.n2592 vdd.t193 4.64847
R5937 vdd.t182 vdd.n912 4.64847
R5938 vdd.n3174 vdd.t178 4.64847
R5939 vdd.n3561 vdd.t15 4.64847
R5940 vdd.n1076 vdd.t289 4.53511
R5941 vdd.n3156 vdd.t262 4.53511
R5942 vdd.n2314 vdd.t9 4.42174
R5943 vdd.n2519 vdd.t237 4.42174
R5944 vdd.n1399 vdd.t278 4.42174
R5945 vdd.n3101 vdd.t285 4.42174
R5946 vdd.n846 vdd.t233 4.42174
R5947 vdd.t109 vdd.n655 4.42174
R5948 vdd.n3147 vdd.n897 4.37123
R5949 vdd.n2578 vdd.n2577 4.37123
R5950 vdd.n2616 vdd.t180 4.30838
R5951 vdd.n3004 vdd.t167 4.30838
R5952 vdd.n312 vdd.n300 4.26717
R5953 vdd.n253 vdd.n241 4.26717
R5954 vdd.n210 vdd.n198 4.26717
R5955 vdd.n151 vdd.n139 4.26717
R5956 vdd.n109 vdd.n97 4.26717
R5957 vdd.n50 vdd.n38 4.26717
R5958 vdd.n2186 vdd.n2174 4.26717
R5959 vdd.n2245 vdd.n2233 4.26717
R5960 vdd.n2084 vdd.n2072 4.26717
R5961 vdd.n2143 vdd.n2131 4.26717
R5962 vdd.n1983 vdd.n1971 4.26717
R5963 vdd.n2042 vdd.n2030 4.26717
R5964 vdd.n2330 vdd.t34 4.19501
R5965 vdd.n3520 vdd.t13 4.19501
R5966 vdd.n333 vdd.n231 4.10845
R5967 vdd.n2266 vdd.n2164 4.10845
R5968 vdd.n289 vdd.t38 4.06363
R5969 vdd.n289 vdd.t200 4.06363
R5970 vdd.n287 vdd.t98 4.06363
R5971 vdd.n287 vdd.t87 4.06363
R5972 vdd.n285 vdd.t209 4.06363
R5973 vdd.n285 vdd.t70 4.06363
R5974 vdd.n283 vdd.t197 4.06363
R5975 vdd.n283 vdd.t65 4.06363
R5976 vdd.n281 vdd.t219 4.06363
R5977 vdd.n281 vdd.t80 4.06363
R5978 vdd.n279 vdd.t66 4.06363
R5979 vdd.n279 vdd.t58 4.06363
R5980 vdd.n277 vdd.t77 4.06363
R5981 vdd.n277 vdd.t225 4.06363
R5982 vdd.n275 vdd.t113 4.06363
R5983 vdd.n275 vdd.t36 4.06363
R5984 vdd.n273 vdd.t119 4.06363
R5985 vdd.n273 vdd.t202 4.06363
R5986 vdd.n187 vdd.t112 4.06363
R5987 vdd.n187 vdd.t221 4.06363
R5988 vdd.n185 vdd.t125 4.06363
R5989 vdd.n185 vdd.t201 4.06363
R5990 vdd.n183 vdd.t105 4.06363
R5991 vdd.n183 vdd.t137 4.06363
R5992 vdd.n181 vdd.t217 4.06363
R5993 vdd.n181 vdd.t140 4.06363
R5994 vdd.n179 vdd.t42 4.06363
R5995 vdd.n179 vdd.t30 4.06363
R5996 vdd.n177 vdd.t136 4.06363
R5997 vdd.n177 vdd.t82 4.06363
R5998 vdd.n175 vdd.t220 4.06363
R5999 vdd.n175 vdd.t16 4.06363
R6000 vdd.n173 vdd.t110 4.06363
R6001 vdd.n173 vdd.t229 4.06363
R6002 vdd.n171 vdd.t117 4.06363
R6003 vdd.n171 vdd.t124 4.06363
R6004 vdd.n86 vdd.t89 4.06363
R6005 vdd.n86 vdd.t26 4.06363
R6006 vdd.n84 vdd.t103 4.06363
R6007 vdd.n84 vdd.t73 4.06363
R6008 vdd.n82 vdd.t218 4.06363
R6009 vdd.n82 vdd.t118 4.06363
R6010 vdd.n80 vdd.t121 4.06363
R6011 vdd.n80 vdd.t212 4.06363
R6012 vdd.n78 vdd.t20 4.06363
R6013 vdd.n78 vdd.t135 4.06363
R6014 vdd.n76 vdd.t56 4.06363
R6015 vdd.n76 vdd.t28 4.06363
R6016 vdd.n74 vdd.t78 4.06363
R6017 vdd.n74 vdd.t79 4.06363
R6018 vdd.n72 vdd.t133 4.06363
R6019 vdd.n72 vdd.t3 4.06363
R6020 vdd.n70 vdd.t139 4.06363
R6021 vdd.n70 vdd.t228 4.06363
R6022 vdd.n2206 vdd.t226 4.06363
R6023 vdd.n2206 vdd.t227 4.06363
R6024 vdd.n2208 vdd.t126 4.06363
R6025 vdd.n2208 vdd.t10 4.06363
R6026 vdd.n2210 vdd.t95 4.06363
R6027 vdd.n2210 vdd.t108 4.06363
R6028 vdd.n2212 vdd.t128 4.06363
R6029 vdd.n2212 vdd.t12 4.06363
R6030 vdd.n2214 vdd.t134 4.06363
R6031 vdd.n2214 vdd.t210 4.06363
R6032 vdd.n2216 vdd.t211 4.06363
R6033 vdd.n2216 vdd.t63 4.06363
R6034 vdd.n2218 vdd.t52 4.06363
R6035 vdd.n2218 vdd.t230 4.06363
R6036 vdd.n2220 vdd.t81 4.06363
R6037 vdd.n2220 vdd.t107 4.06363
R6038 vdd.n2222 vdd.t207 4.06363
R6039 vdd.n2222 vdd.t127 4.06363
R6040 vdd.n2104 vdd.t92 4.06363
R6041 vdd.n2104 vdd.t205 4.06363
R6042 vdd.n2106 vdd.t61 4.06363
R6043 vdd.n2106 vdd.t93 4.06363
R6044 vdd.n2108 vdd.t60 4.06363
R6045 vdd.n2108 vdd.t102 4.06363
R6046 vdd.n2110 vdd.t54 4.06363
R6047 vdd.n2110 vdd.t94 4.06363
R6048 vdd.n2112 vdd.t75 4.06363
R6049 vdd.n2112 vdd.t31 4.06363
R6050 vdd.n2114 vdd.t208 4.06363
R6051 vdd.n2114 vdd.t44 4.06363
R6052 vdd.n2116 vdd.t222 4.06363
R6053 vdd.n2116 vdd.t115 4.06363
R6054 vdd.n2118 vdd.t130 4.06363
R6055 vdd.n2118 vdd.t203 4.06363
R6056 vdd.n2120 vdd.t33 4.06363
R6057 vdd.n2120 vdd.t199 4.06363
R6058 vdd.n2003 vdd.t213 4.06363
R6059 vdd.n2003 vdd.t216 4.06363
R6060 vdd.n2005 vdd.t1 4.06363
R6061 vdd.n2005 vdd.t96 4.06363
R6062 vdd.n2007 vdd.t90 4.06363
R6063 vdd.n2007 vdd.t100 4.06363
R6064 vdd.n2009 vdd.t215 4.06363
R6065 vdd.n2009 vdd.t88 4.06363
R6066 vdd.n2011 vdd.t111 4.06363
R6067 vdd.n2011 vdd.t18 4.06363
R6068 vdd.n2013 vdd.t132 4.06363
R6069 vdd.n2013 vdd.t122 4.06363
R6070 vdd.n2015 vdd.t231 4.06363
R6071 vdd.n2015 vdd.t129 4.06363
R6072 vdd.n2017 vdd.t68 4.06363
R6073 vdd.n2017 vdd.t224 4.06363
R6074 vdd.n2019 vdd.t214 4.06363
R6075 vdd.n2019 vdd.t86 4.06363
R6076 vdd.n1112 vdd.t186 3.96828
R6077 vdd.n2610 vdd.t166 3.96828
R6078 vdd.n2998 vdd.t183 3.96828
R6079 vdd.n3192 vdd.t172 3.96828
R6080 vdd.n26 vdd.t46 3.9605
R6081 vdd.n26 vdd.t84 3.9605
R6082 vdd.n23 vdd.t5 3.9605
R6083 vdd.n23 vdd.t83 3.9605
R6084 vdd.n21 vdd.t50 3.9605
R6085 vdd.n21 vdd.t39 3.9605
R6086 vdd.n20 vdd.t6 3.9605
R6087 vdd.n20 vdd.t48 3.9605
R6088 vdd.n15 vdd.t49 3.9605
R6089 vdd.n15 vdd.t8 3.9605
R6090 vdd.n16 vdd.t45 3.9605
R6091 vdd.n16 vdd.t47 3.9605
R6092 vdd.n18 vdd.t40 3.9605
R6093 vdd.n18 vdd.t4 3.9605
R6094 vdd.n25 vdd.t41 3.9605
R6095 vdd.n25 vdd.t7 3.9605
R6096 vdd.n2543 vdd.t186 3.74155
R6097 vdd.n1046 vdd.t166 3.74155
R6098 vdd.n3125 vdd.t183 3.74155
R6099 vdd.n870 vdd.t172 3.74155
R6100 vdd.n7 vdd.t196 3.61217
R6101 vdd.n7 vdd.t160 3.61217
R6102 vdd.n8 vdd.t168 3.61217
R6103 vdd.n8 vdd.t188 3.61217
R6104 vdd.n10 vdd.t177 3.61217
R6105 vdd.n10 vdd.t148 3.61217
R6106 vdd.n12 vdd.t157 3.61217
R6107 vdd.n12 vdd.t175 3.61217
R6108 vdd.n5 vdd.t190 3.61217
R6109 vdd.n5 vdd.t170 3.61217
R6110 vdd.n3 vdd.t162 3.61217
R6111 vdd.n3 vdd.t192 3.61217
R6112 vdd.n1 vdd.t144 3.61217
R6113 vdd.n1 vdd.t181 3.61217
R6114 vdd.n0 vdd.t185 3.61217
R6115 vdd.n0 vdd.t165 3.61217
R6116 vdd.n316 vdd.n315 3.49141
R6117 vdd.n257 vdd.n256 3.49141
R6118 vdd.n214 vdd.n213 3.49141
R6119 vdd.n155 vdd.n154 3.49141
R6120 vdd.n113 vdd.n112 3.49141
R6121 vdd.n54 vdd.n53 3.49141
R6122 vdd.n2190 vdd.n2189 3.49141
R6123 vdd.n2249 vdd.n2248 3.49141
R6124 vdd.n2088 vdd.n2087 3.49141
R6125 vdd.n2147 vdd.n2146 3.49141
R6126 vdd.n1987 vdd.n1986 3.49141
R6127 vdd.n2046 vdd.n2045 3.49141
R6128 vdd.t180 vdd.n1028 3.40145
R6129 vdd.n2784 vdd.t189 3.40145
R6130 vdd.n3088 vdd.t174 3.40145
R6131 vdd.n3113 vdd.t167 3.40145
R6132 vdd.n2331 vdd.t204 3.28809
R6133 vdd.n1137 vdd.t237 3.28809
R6134 vdd.n2637 vdd.t278 3.28809
R6135 vdd.n3016 vdd.t285 3.28809
R6136 vdd.n3261 vdd.t233 3.28809
R6137 vdd.n3519 vdd.t116 3.28809
R6138 vdd.t0 vdd.n1559 3.06136
R6139 vdd.n2555 vdd.t154 3.06136
R6140 vdd.n1437 vdd.t193 3.06136
R6141 vdd.n3137 vdd.t182 3.06136
R6142 vdd.t178 vdd.n874 3.06136
R6143 vdd.n3544 vdd.t2 3.06136
R6144 vdd.n2630 vdd.t161 2.94799
R6145 vdd.t147 vdd.n946 2.94799
R6146 vdd.n2289 vdd.t11 2.83463
R6147 vdd.n644 vdd.t55 2.83463
R6148 vdd.n319 vdd.n298 2.71565
R6149 vdd.n260 vdd.n239 2.71565
R6150 vdd.n217 vdd.n196 2.71565
R6151 vdd.n158 vdd.n137 2.71565
R6152 vdd.n116 vdd.n95 2.71565
R6153 vdd.n57 vdd.n36 2.71565
R6154 vdd.n2193 vdd.n2172 2.71565
R6155 vdd.n2252 vdd.n2231 2.71565
R6156 vdd.n2091 vdd.n2070 2.71565
R6157 vdd.n2150 vdd.n2129 2.71565
R6158 vdd.n1990 vdd.n1969 2.71565
R6159 vdd.n2049 vdd.n2028 2.71565
R6160 vdd.t74 vdd.n1587 2.6079
R6161 vdd.n3667 vdd.t29 2.6079
R6162 vdd.n2604 vdd.t164 2.49453
R6163 vdd.n931 vdd.t195 2.49453
R6164 vdd.n306 vdd.n305 2.4129
R6165 vdd.n247 vdd.n246 2.4129
R6166 vdd.n204 vdd.n203 2.4129
R6167 vdd.n145 vdd.n144 2.4129
R6168 vdd.n103 vdd.n102 2.4129
R6169 vdd.n44 vdd.n43 2.4129
R6170 vdd.n2180 vdd.n2179 2.4129
R6171 vdd.n2239 vdd.n2238 2.4129
R6172 vdd.n2078 vdd.n2077 2.4129
R6173 vdd.n2137 vdd.n2136 2.4129
R6174 vdd.n1977 vdd.n1976 2.4129
R6175 vdd.n2036 vdd.n2035 2.4129
R6176 vdd.n1941 vdd.t114 2.38117
R6177 vdd.n2349 vdd.t241 2.38117
R6178 vdd.n3503 vdd.t258 2.38117
R6179 vdd.n3658 vdd.t104 2.38117
R6180 vdd.n2474 vdd.n1180 2.27742
R6181 vdd.n2474 vdd.n1179 2.27742
R6182 vdd.n3488 vdd.n3487 2.27742
R6183 vdd.n3489 vdd.n3488 2.27742
R6184 vdd.n3366 vdd.n3365 2.27742
R6185 vdd.n3365 vdd.n784 2.27742
R6186 vdd.n2368 vdd.n2367 2.27742
R6187 vdd.n2367 vdd.n1516 2.27742
R6188 vdd.t67 vdd.n1616 2.15444
R6189 vdd.n1083 vdd.t173 2.15444
R6190 vdd.n2580 vdd.t151 2.15444
R6191 vdd.n908 vdd.t150 2.15444
R6192 vdd.n3162 vdd.t149 2.15444
R6193 vdd.n3649 vdd.t72 2.15444
R6194 vdd.n320 vdd.n296 1.93989
R6195 vdd.n261 vdd.n237 1.93989
R6196 vdd.n218 vdd.n194 1.93989
R6197 vdd.n159 vdd.n135 1.93989
R6198 vdd.n117 vdd.n93 1.93989
R6199 vdd.n58 vdd.n34 1.93989
R6200 vdd.n2194 vdd.n2170 1.93989
R6201 vdd.n2253 vdd.n2229 1.93989
R6202 vdd.n2092 vdd.n2068 1.93989
R6203 vdd.n2151 vdd.n2127 1.93989
R6204 vdd.n1991 vdd.n1967 1.93989
R6205 vdd.n2050 vdd.n2026 1.93989
R6206 vdd.n1899 vdd.t21 1.92771
R6207 vdd.t23 vdd.n375 1.92771
R6208 vdd.n1437 vdd.t184 1.81434
R6209 vdd.n3137 vdd.t159 1.81434
R6210 vdd.n1907 vdd.t85 1.70098
R6211 vdd.n3643 vdd.t37 1.70098
R6212 vdd.n1932 vdd.t51 1.47425
R6213 vdd.n361 vdd.t69 1.47425
R6214 vdd.t191 vdd.n1005 1.36088
R6215 vdd.n3095 vdd.t176 1.36088
R6216 vdd.n1598 vdd.t43 1.24752
R6217 vdd.t153 vdd.n1080 1.24752
R6218 vdd.n2586 vdd.t158 1.24752
R6219 vdd.t163 vdd.n905 1.24752
R6220 vdd.n3168 vdd.t179 1.24752
R6221 vdd.t120 vdd.n3665 1.24752
R6222 vdd.n2267 vdd.n28 1.21639
R6223 vdd vdd.n3672 1.20856
R6224 vdd.n331 vdd.n291 1.16414
R6225 vdd.n324 vdd.n323 1.16414
R6226 vdd.n272 vdd.n232 1.16414
R6227 vdd.n265 vdd.n264 1.16414
R6228 vdd.n229 vdd.n189 1.16414
R6229 vdd.n222 vdd.n221 1.16414
R6230 vdd.n170 vdd.n130 1.16414
R6231 vdd.n163 vdd.n162 1.16414
R6232 vdd.n128 vdd.n88 1.16414
R6233 vdd.n121 vdd.n120 1.16414
R6234 vdd.n69 vdd.n29 1.16414
R6235 vdd.n62 vdd.n61 1.16414
R6236 vdd.n2205 vdd.n2165 1.16414
R6237 vdd.n2198 vdd.n2197 1.16414
R6238 vdd.n2264 vdd.n2224 1.16414
R6239 vdd.n2257 vdd.n2256 1.16414
R6240 vdd.n2103 vdd.n2063 1.16414
R6241 vdd.n2096 vdd.n2095 1.16414
R6242 vdd.n2162 vdd.n2122 1.16414
R6243 vdd.n2155 vdd.n2154 1.16414
R6244 vdd.n2002 vdd.n1962 1.16414
R6245 vdd.n1995 vdd.n1994 1.16414
R6246 vdd.n2061 vdd.n2021 1.16414
R6247 vdd.n2054 vdd.n2053 1.16414
R6248 vdd.n2281 vdd.t53 1.02079
R6249 vdd.t289 vdd.t151 1.02079
R6250 vdd.t150 vdd.t262 1.02079
R6251 vdd.t27 vdd.n633 1.02079
R6252 vdd.n1778 vdd.n1774 0.970197
R6253 vdd.n2365 vdd.n2364 0.970197
R6254 vdd.n618 vdd.n428 0.970197
R6255 vdd.n3367 vdd.n690 0.970197
R6256 vdd.n2610 vdd.t143 0.907421
R6257 vdd.n2998 vdd.t187 0.907421
R6258 vdd.n2297 vdd.t99 0.794056
R6259 vdd.n3553 vdd.t76 0.794056
R6260 vdd.n2322 vdd.t91 0.567326
R6261 vdd.n1119 vdd.t146 0.567326
R6262 vdd.n2616 vdd.t142 0.567326
R6263 vdd.n3004 vdd.t145 0.567326
R6264 vdd.n3198 vdd.t155 0.567326
R6265 vdd.t123 vdd.n662 0.567326
R6266 vdd.n2355 vdd.n1181 0.530988
R6267 vdd.n726 vdd.n682 0.530988
R6268 vdd.n464 vdd.n391 0.530988
R6269 vdd.n3622 vdd.n3621 0.530988
R6270 vdd.n3499 vdd.n3498 0.530988
R6271 vdd.n2344 vdd.n1517 0.530988
R6272 vdd.n1776 vdd.n1641 0.530988
R6273 vdd.n1878 vdd.n1877 0.530988
R6274 vdd.n4 vdd.n2 0.459552
R6275 vdd.n11 vdd.n9 0.459552
R6276 vdd.n329 vdd.n328 0.388379
R6277 vdd.n295 vdd.n293 0.388379
R6278 vdd.n270 vdd.n269 0.388379
R6279 vdd.n236 vdd.n234 0.388379
R6280 vdd.n227 vdd.n226 0.388379
R6281 vdd.n193 vdd.n191 0.388379
R6282 vdd.n168 vdd.n167 0.388379
R6283 vdd.n134 vdd.n132 0.388379
R6284 vdd.n126 vdd.n125 0.388379
R6285 vdd.n92 vdd.n90 0.388379
R6286 vdd.n67 vdd.n66 0.388379
R6287 vdd.n33 vdd.n31 0.388379
R6288 vdd.n2203 vdd.n2202 0.388379
R6289 vdd.n2169 vdd.n2167 0.388379
R6290 vdd.n2262 vdd.n2261 0.388379
R6291 vdd.n2228 vdd.n2226 0.388379
R6292 vdd.n2101 vdd.n2100 0.388379
R6293 vdd.n2067 vdd.n2065 0.388379
R6294 vdd.n2160 vdd.n2159 0.388379
R6295 vdd.n2126 vdd.n2124 0.388379
R6296 vdd.n2000 vdd.n1999 0.388379
R6297 vdd.n1966 vdd.n1964 0.388379
R6298 vdd.n2059 vdd.n2058 0.388379
R6299 vdd.n2025 vdd.n2023 0.388379
R6300 vdd.n19 vdd.n17 0.387128
R6301 vdd.n24 vdd.n22 0.387128
R6302 vdd.n6 vdd.n4 0.358259
R6303 vdd.n13 vdd.n11 0.358259
R6304 vdd.n276 vdd.n274 0.358259
R6305 vdd.n278 vdd.n276 0.358259
R6306 vdd.n280 vdd.n278 0.358259
R6307 vdd.n282 vdd.n280 0.358259
R6308 vdd.n284 vdd.n282 0.358259
R6309 vdd.n286 vdd.n284 0.358259
R6310 vdd.n288 vdd.n286 0.358259
R6311 vdd.n290 vdd.n288 0.358259
R6312 vdd.n332 vdd.n290 0.358259
R6313 vdd.n174 vdd.n172 0.358259
R6314 vdd.n176 vdd.n174 0.358259
R6315 vdd.n178 vdd.n176 0.358259
R6316 vdd.n180 vdd.n178 0.358259
R6317 vdd.n182 vdd.n180 0.358259
R6318 vdd.n184 vdd.n182 0.358259
R6319 vdd.n186 vdd.n184 0.358259
R6320 vdd.n188 vdd.n186 0.358259
R6321 vdd.n230 vdd.n188 0.358259
R6322 vdd.n73 vdd.n71 0.358259
R6323 vdd.n75 vdd.n73 0.358259
R6324 vdd.n77 vdd.n75 0.358259
R6325 vdd.n79 vdd.n77 0.358259
R6326 vdd.n81 vdd.n79 0.358259
R6327 vdd.n83 vdd.n81 0.358259
R6328 vdd.n85 vdd.n83 0.358259
R6329 vdd.n87 vdd.n85 0.358259
R6330 vdd.n129 vdd.n87 0.358259
R6331 vdd.n2265 vdd.n2223 0.358259
R6332 vdd.n2223 vdd.n2221 0.358259
R6333 vdd.n2221 vdd.n2219 0.358259
R6334 vdd.n2219 vdd.n2217 0.358259
R6335 vdd.n2217 vdd.n2215 0.358259
R6336 vdd.n2215 vdd.n2213 0.358259
R6337 vdd.n2213 vdd.n2211 0.358259
R6338 vdd.n2211 vdd.n2209 0.358259
R6339 vdd.n2209 vdd.n2207 0.358259
R6340 vdd.n2163 vdd.n2121 0.358259
R6341 vdd.n2121 vdd.n2119 0.358259
R6342 vdd.n2119 vdd.n2117 0.358259
R6343 vdd.n2117 vdd.n2115 0.358259
R6344 vdd.n2115 vdd.n2113 0.358259
R6345 vdd.n2113 vdd.n2111 0.358259
R6346 vdd.n2111 vdd.n2109 0.358259
R6347 vdd.n2109 vdd.n2107 0.358259
R6348 vdd.n2107 vdd.n2105 0.358259
R6349 vdd.n2062 vdd.n2020 0.358259
R6350 vdd.n2020 vdd.n2018 0.358259
R6351 vdd.n2018 vdd.n2016 0.358259
R6352 vdd.n2016 vdd.n2014 0.358259
R6353 vdd.n2014 vdd.n2012 0.358259
R6354 vdd.n2012 vdd.n2010 0.358259
R6355 vdd.n2010 vdd.n2008 0.358259
R6356 vdd.n2008 vdd.n2006 0.358259
R6357 vdd.n2006 vdd.n2004 0.358259
R6358 vdd.n2549 vdd.t194 0.340595
R6359 vdd.n1052 vdd.t152 0.340595
R6360 vdd.n3131 vdd.t141 0.340595
R6361 vdd.n877 vdd.t171 0.340595
R6362 vdd.n14 vdd.n6 0.334552
R6363 vdd.n14 vdd.n13 0.334552
R6364 vdd.n27 vdd.n19 0.21707
R6365 vdd.n27 vdd.n24 0.21707
R6366 vdd.n330 vdd.n292 0.155672
R6367 vdd.n322 vdd.n292 0.155672
R6368 vdd.n322 vdd.n321 0.155672
R6369 vdd.n321 vdd.n297 0.155672
R6370 vdd.n314 vdd.n297 0.155672
R6371 vdd.n314 vdd.n313 0.155672
R6372 vdd.n313 vdd.n301 0.155672
R6373 vdd.n306 vdd.n301 0.155672
R6374 vdd.n271 vdd.n233 0.155672
R6375 vdd.n263 vdd.n233 0.155672
R6376 vdd.n263 vdd.n262 0.155672
R6377 vdd.n262 vdd.n238 0.155672
R6378 vdd.n255 vdd.n238 0.155672
R6379 vdd.n255 vdd.n254 0.155672
R6380 vdd.n254 vdd.n242 0.155672
R6381 vdd.n247 vdd.n242 0.155672
R6382 vdd.n228 vdd.n190 0.155672
R6383 vdd.n220 vdd.n190 0.155672
R6384 vdd.n220 vdd.n219 0.155672
R6385 vdd.n219 vdd.n195 0.155672
R6386 vdd.n212 vdd.n195 0.155672
R6387 vdd.n212 vdd.n211 0.155672
R6388 vdd.n211 vdd.n199 0.155672
R6389 vdd.n204 vdd.n199 0.155672
R6390 vdd.n169 vdd.n131 0.155672
R6391 vdd.n161 vdd.n131 0.155672
R6392 vdd.n161 vdd.n160 0.155672
R6393 vdd.n160 vdd.n136 0.155672
R6394 vdd.n153 vdd.n136 0.155672
R6395 vdd.n153 vdd.n152 0.155672
R6396 vdd.n152 vdd.n140 0.155672
R6397 vdd.n145 vdd.n140 0.155672
R6398 vdd.n127 vdd.n89 0.155672
R6399 vdd.n119 vdd.n89 0.155672
R6400 vdd.n119 vdd.n118 0.155672
R6401 vdd.n118 vdd.n94 0.155672
R6402 vdd.n111 vdd.n94 0.155672
R6403 vdd.n111 vdd.n110 0.155672
R6404 vdd.n110 vdd.n98 0.155672
R6405 vdd.n103 vdd.n98 0.155672
R6406 vdd.n68 vdd.n30 0.155672
R6407 vdd.n60 vdd.n30 0.155672
R6408 vdd.n60 vdd.n59 0.155672
R6409 vdd.n59 vdd.n35 0.155672
R6410 vdd.n52 vdd.n35 0.155672
R6411 vdd.n52 vdd.n51 0.155672
R6412 vdd.n51 vdd.n39 0.155672
R6413 vdd.n44 vdd.n39 0.155672
R6414 vdd.n2204 vdd.n2166 0.155672
R6415 vdd.n2196 vdd.n2166 0.155672
R6416 vdd.n2196 vdd.n2195 0.155672
R6417 vdd.n2195 vdd.n2171 0.155672
R6418 vdd.n2188 vdd.n2171 0.155672
R6419 vdd.n2188 vdd.n2187 0.155672
R6420 vdd.n2187 vdd.n2175 0.155672
R6421 vdd.n2180 vdd.n2175 0.155672
R6422 vdd.n2263 vdd.n2225 0.155672
R6423 vdd.n2255 vdd.n2225 0.155672
R6424 vdd.n2255 vdd.n2254 0.155672
R6425 vdd.n2254 vdd.n2230 0.155672
R6426 vdd.n2247 vdd.n2230 0.155672
R6427 vdd.n2247 vdd.n2246 0.155672
R6428 vdd.n2246 vdd.n2234 0.155672
R6429 vdd.n2239 vdd.n2234 0.155672
R6430 vdd.n2102 vdd.n2064 0.155672
R6431 vdd.n2094 vdd.n2064 0.155672
R6432 vdd.n2094 vdd.n2093 0.155672
R6433 vdd.n2093 vdd.n2069 0.155672
R6434 vdd.n2086 vdd.n2069 0.155672
R6435 vdd.n2086 vdd.n2085 0.155672
R6436 vdd.n2085 vdd.n2073 0.155672
R6437 vdd.n2078 vdd.n2073 0.155672
R6438 vdd.n2161 vdd.n2123 0.155672
R6439 vdd.n2153 vdd.n2123 0.155672
R6440 vdd.n2153 vdd.n2152 0.155672
R6441 vdd.n2152 vdd.n2128 0.155672
R6442 vdd.n2145 vdd.n2128 0.155672
R6443 vdd.n2145 vdd.n2144 0.155672
R6444 vdd.n2144 vdd.n2132 0.155672
R6445 vdd.n2137 vdd.n2132 0.155672
R6446 vdd.n2001 vdd.n1963 0.155672
R6447 vdd.n1993 vdd.n1963 0.155672
R6448 vdd.n1993 vdd.n1992 0.155672
R6449 vdd.n1992 vdd.n1968 0.155672
R6450 vdd.n1985 vdd.n1968 0.155672
R6451 vdd.n1985 vdd.n1984 0.155672
R6452 vdd.n1984 vdd.n1972 0.155672
R6453 vdd.n1977 vdd.n1972 0.155672
R6454 vdd.n2060 vdd.n2022 0.155672
R6455 vdd.n2052 vdd.n2022 0.155672
R6456 vdd.n2052 vdd.n2051 0.155672
R6457 vdd.n2051 vdd.n2027 0.155672
R6458 vdd.n2044 vdd.n2027 0.155672
R6459 vdd.n2044 vdd.n2043 0.155672
R6460 vdd.n2043 vdd.n2031 0.155672
R6461 vdd.n2036 vdd.n2031 0.155672
R6462 vdd.n1186 vdd.n1178 0.152939
R6463 vdd.n1190 vdd.n1186 0.152939
R6464 vdd.n1191 vdd.n1190 0.152939
R6465 vdd.n1192 vdd.n1191 0.152939
R6466 vdd.n1193 vdd.n1192 0.152939
R6467 vdd.n1197 vdd.n1193 0.152939
R6468 vdd.n1198 vdd.n1197 0.152939
R6469 vdd.n1199 vdd.n1198 0.152939
R6470 vdd.n1200 vdd.n1199 0.152939
R6471 vdd.n1204 vdd.n1200 0.152939
R6472 vdd.n1205 vdd.n1204 0.152939
R6473 vdd.n1206 vdd.n1205 0.152939
R6474 vdd.n2438 vdd.n1206 0.152939
R6475 vdd.n2438 vdd.n2437 0.152939
R6476 vdd.n2437 vdd.n2436 0.152939
R6477 vdd.n2436 vdd.n1212 0.152939
R6478 vdd.n1217 vdd.n1212 0.152939
R6479 vdd.n1218 vdd.n1217 0.152939
R6480 vdd.n1219 vdd.n1218 0.152939
R6481 vdd.n1223 vdd.n1219 0.152939
R6482 vdd.n1224 vdd.n1223 0.152939
R6483 vdd.n1225 vdd.n1224 0.152939
R6484 vdd.n1226 vdd.n1225 0.152939
R6485 vdd.n1230 vdd.n1226 0.152939
R6486 vdd.n1231 vdd.n1230 0.152939
R6487 vdd.n1232 vdd.n1231 0.152939
R6488 vdd.n1233 vdd.n1232 0.152939
R6489 vdd.n1237 vdd.n1233 0.152939
R6490 vdd.n1238 vdd.n1237 0.152939
R6491 vdd.n1239 vdd.n1238 0.152939
R6492 vdd.n1240 vdd.n1239 0.152939
R6493 vdd.n1244 vdd.n1240 0.152939
R6494 vdd.n1245 vdd.n1244 0.152939
R6495 vdd.n1246 vdd.n1245 0.152939
R6496 vdd.n2399 vdd.n1246 0.152939
R6497 vdd.n2399 vdd.n2398 0.152939
R6498 vdd.n2398 vdd.n2397 0.152939
R6499 vdd.n2397 vdd.n1252 0.152939
R6500 vdd.n1257 vdd.n1252 0.152939
R6501 vdd.n1258 vdd.n1257 0.152939
R6502 vdd.n1259 vdd.n1258 0.152939
R6503 vdd.n1263 vdd.n1259 0.152939
R6504 vdd.n1264 vdd.n1263 0.152939
R6505 vdd.n1265 vdd.n1264 0.152939
R6506 vdd.n1266 vdd.n1265 0.152939
R6507 vdd.n1270 vdd.n1266 0.152939
R6508 vdd.n1271 vdd.n1270 0.152939
R6509 vdd.n1272 vdd.n1271 0.152939
R6510 vdd.n1273 vdd.n1272 0.152939
R6511 vdd.n1277 vdd.n1273 0.152939
R6512 vdd.n1278 vdd.n1277 0.152939
R6513 vdd.n2473 vdd.n1181 0.152939
R6514 vdd.n2269 vdd.n1578 0.152939
R6515 vdd.n2284 vdd.n1578 0.152939
R6516 vdd.n2285 vdd.n2284 0.152939
R6517 vdd.n2286 vdd.n2285 0.152939
R6518 vdd.n2286 vdd.n1567 0.152939
R6519 vdd.n2301 vdd.n1567 0.152939
R6520 vdd.n2302 vdd.n2301 0.152939
R6521 vdd.n2303 vdd.n2302 0.152939
R6522 vdd.n2303 vdd.n1556 0.152939
R6523 vdd.n2317 vdd.n1556 0.152939
R6524 vdd.n2318 vdd.n2317 0.152939
R6525 vdd.n2319 vdd.n2318 0.152939
R6526 vdd.n2319 vdd.n1544 0.152939
R6527 vdd.n2334 vdd.n1544 0.152939
R6528 vdd.n2335 vdd.n2334 0.152939
R6529 vdd.n2336 vdd.n2335 0.152939
R6530 vdd.n2336 vdd.n1532 0.152939
R6531 vdd.n2353 vdd.n1532 0.152939
R6532 vdd.n2354 vdd.n2353 0.152939
R6533 vdd.n2355 vdd.n2354 0.152939
R6534 vdd.n735 vdd.n730 0.152939
R6535 vdd.n736 vdd.n735 0.152939
R6536 vdd.n737 vdd.n736 0.152939
R6537 vdd.n738 vdd.n737 0.152939
R6538 vdd.n739 vdd.n738 0.152939
R6539 vdd.n740 vdd.n739 0.152939
R6540 vdd.n741 vdd.n740 0.152939
R6541 vdd.n742 vdd.n741 0.152939
R6542 vdd.n743 vdd.n742 0.152939
R6543 vdd.n744 vdd.n743 0.152939
R6544 vdd.n745 vdd.n744 0.152939
R6545 vdd.n746 vdd.n745 0.152939
R6546 vdd.n3455 vdd.n746 0.152939
R6547 vdd.n3455 vdd.n3454 0.152939
R6548 vdd.n3454 vdd.n3453 0.152939
R6549 vdd.n3453 vdd.n748 0.152939
R6550 vdd.n749 vdd.n748 0.152939
R6551 vdd.n750 vdd.n749 0.152939
R6552 vdd.n751 vdd.n750 0.152939
R6553 vdd.n752 vdd.n751 0.152939
R6554 vdd.n753 vdd.n752 0.152939
R6555 vdd.n754 vdd.n753 0.152939
R6556 vdd.n755 vdd.n754 0.152939
R6557 vdd.n756 vdd.n755 0.152939
R6558 vdd.n757 vdd.n756 0.152939
R6559 vdd.n758 vdd.n757 0.152939
R6560 vdd.n759 vdd.n758 0.152939
R6561 vdd.n760 vdd.n759 0.152939
R6562 vdd.n761 vdd.n760 0.152939
R6563 vdd.n762 vdd.n761 0.152939
R6564 vdd.n763 vdd.n762 0.152939
R6565 vdd.n764 vdd.n763 0.152939
R6566 vdd.n765 vdd.n764 0.152939
R6567 vdd.n766 vdd.n765 0.152939
R6568 vdd.n3409 vdd.n766 0.152939
R6569 vdd.n3409 vdd.n3408 0.152939
R6570 vdd.n3408 vdd.n3407 0.152939
R6571 vdd.n3407 vdd.n770 0.152939
R6572 vdd.n771 vdd.n770 0.152939
R6573 vdd.n772 vdd.n771 0.152939
R6574 vdd.n773 vdd.n772 0.152939
R6575 vdd.n774 vdd.n773 0.152939
R6576 vdd.n775 vdd.n774 0.152939
R6577 vdd.n776 vdd.n775 0.152939
R6578 vdd.n777 vdd.n776 0.152939
R6579 vdd.n778 vdd.n777 0.152939
R6580 vdd.n779 vdd.n778 0.152939
R6581 vdd.n780 vdd.n779 0.152939
R6582 vdd.n781 vdd.n780 0.152939
R6583 vdd.n782 vdd.n781 0.152939
R6584 vdd.n783 vdd.n782 0.152939
R6585 vdd.n727 vdd.n726 0.152939
R6586 vdd.n3506 vdd.n682 0.152939
R6587 vdd.n3507 vdd.n3506 0.152939
R6588 vdd.n3508 vdd.n3507 0.152939
R6589 vdd.n3508 vdd.n670 0.152939
R6590 vdd.n3523 vdd.n670 0.152939
R6591 vdd.n3524 vdd.n3523 0.152939
R6592 vdd.n3525 vdd.n3524 0.152939
R6593 vdd.n3525 vdd.n659 0.152939
R6594 vdd.n3539 vdd.n659 0.152939
R6595 vdd.n3540 vdd.n3539 0.152939
R6596 vdd.n3541 vdd.n3540 0.152939
R6597 vdd.n3541 vdd.n647 0.152939
R6598 vdd.n3556 vdd.n647 0.152939
R6599 vdd.n3557 vdd.n3556 0.152939
R6600 vdd.n3558 vdd.n3557 0.152939
R6601 vdd.n3558 vdd.n636 0.152939
R6602 vdd.n3575 vdd.n636 0.152939
R6603 vdd.n3576 vdd.n3575 0.152939
R6604 vdd.n3577 vdd.n3576 0.152939
R6605 vdd.n3577 vdd.n334 0.152939
R6606 vdd.n3670 vdd.n335 0.152939
R6607 vdd.n346 vdd.n335 0.152939
R6608 vdd.n347 vdd.n346 0.152939
R6609 vdd.n348 vdd.n347 0.152939
R6610 vdd.n355 vdd.n348 0.152939
R6611 vdd.n356 vdd.n355 0.152939
R6612 vdd.n357 vdd.n356 0.152939
R6613 vdd.n358 vdd.n357 0.152939
R6614 vdd.n366 vdd.n358 0.152939
R6615 vdd.n367 vdd.n366 0.152939
R6616 vdd.n368 vdd.n367 0.152939
R6617 vdd.n369 vdd.n368 0.152939
R6618 vdd.n377 vdd.n369 0.152939
R6619 vdd.n378 vdd.n377 0.152939
R6620 vdd.n379 vdd.n378 0.152939
R6621 vdd.n380 vdd.n379 0.152939
R6622 vdd.n388 vdd.n380 0.152939
R6623 vdd.n389 vdd.n388 0.152939
R6624 vdd.n390 vdd.n389 0.152939
R6625 vdd.n391 vdd.n390 0.152939
R6626 vdd.n464 vdd.n463 0.152939
R6627 vdd.n470 vdd.n463 0.152939
R6628 vdd.n471 vdd.n470 0.152939
R6629 vdd.n472 vdd.n471 0.152939
R6630 vdd.n472 vdd.n461 0.152939
R6631 vdd.n480 vdd.n461 0.152939
R6632 vdd.n481 vdd.n480 0.152939
R6633 vdd.n482 vdd.n481 0.152939
R6634 vdd.n482 vdd.n459 0.152939
R6635 vdd.n490 vdd.n459 0.152939
R6636 vdd.n491 vdd.n490 0.152939
R6637 vdd.n492 vdd.n491 0.152939
R6638 vdd.n492 vdd.n457 0.152939
R6639 vdd.n500 vdd.n457 0.152939
R6640 vdd.n501 vdd.n500 0.152939
R6641 vdd.n502 vdd.n501 0.152939
R6642 vdd.n502 vdd.n455 0.152939
R6643 vdd.n510 vdd.n455 0.152939
R6644 vdd.n511 vdd.n510 0.152939
R6645 vdd.n512 vdd.n511 0.152939
R6646 vdd.n512 vdd.n451 0.152939
R6647 vdd.n520 vdd.n451 0.152939
R6648 vdd.n521 vdd.n520 0.152939
R6649 vdd.n522 vdd.n521 0.152939
R6650 vdd.n522 vdd.n449 0.152939
R6651 vdd.n530 vdd.n449 0.152939
R6652 vdd.n531 vdd.n530 0.152939
R6653 vdd.n532 vdd.n531 0.152939
R6654 vdd.n532 vdd.n447 0.152939
R6655 vdd.n540 vdd.n447 0.152939
R6656 vdd.n541 vdd.n540 0.152939
R6657 vdd.n542 vdd.n541 0.152939
R6658 vdd.n542 vdd.n445 0.152939
R6659 vdd.n550 vdd.n445 0.152939
R6660 vdd.n551 vdd.n550 0.152939
R6661 vdd.n552 vdd.n551 0.152939
R6662 vdd.n552 vdd.n443 0.152939
R6663 vdd.n560 vdd.n443 0.152939
R6664 vdd.n561 vdd.n560 0.152939
R6665 vdd.n562 vdd.n561 0.152939
R6666 vdd.n562 vdd.n439 0.152939
R6667 vdd.n570 vdd.n439 0.152939
R6668 vdd.n571 vdd.n570 0.152939
R6669 vdd.n572 vdd.n571 0.152939
R6670 vdd.n572 vdd.n437 0.152939
R6671 vdd.n580 vdd.n437 0.152939
R6672 vdd.n581 vdd.n580 0.152939
R6673 vdd.n582 vdd.n581 0.152939
R6674 vdd.n582 vdd.n435 0.152939
R6675 vdd.n590 vdd.n435 0.152939
R6676 vdd.n591 vdd.n590 0.152939
R6677 vdd.n592 vdd.n591 0.152939
R6678 vdd.n592 vdd.n433 0.152939
R6679 vdd.n600 vdd.n433 0.152939
R6680 vdd.n601 vdd.n600 0.152939
R6681 vdd.n602 vdd.n601 0.152939
R6682 vdd.n602 vdd.n431 0.152939
R6683 vdd.n610 vdd.n431 0.152939
R6684 vdd.n611 vdd.n610 0.152939
R6685 vdd.n612 vdd.n611 0.152939
R6686 vdd.n612 vdd.n429 0.152939
R6687 vdd.n619 vdd.n429 0.152939
R6688 vdd.n3622 vdd.n619 0.152939
R6689 vdd.n3500 vdd.n3499 0.152939
R6690 vdd.n3500 vdd.n675 0.152939
R6691 vdd.n3514 vdd.n675 0.152939
R6692 vdd.n3515 vdd.n3514 0.152939
R6693 vdd.n3516 vdd.n3515 0.152939
R6694 vdd.n3516 vdd.n665 0.152939
R6695 vdd.n3531 vdd.n665 0.152939
R6696 vdd.n3532 vdd.n3531 0.152939
R6697 vdd.n3533 vdd.n3532 0.152939
R6698 vdd.n3533 vdd.n652 0.152939
R6699 vdd.n3547 vdd.n652 0.152939
R6700 vdd.n3548 vdd.n3547 0.152939
R6701 vdd.n3549 vdd.n3548 0.152939
R6702 vdd.n3549 vdd.n641 0.152939
R6703 vdd.n3564 vdd.n641 0.152939
R6704 vdd.n3565 vdd.n3564 0.152939
R6705 vdd.n3566 vdd.n3565 0.152939
R6706 vdd.n3568 vdd.n3566 0.152939
R6707 vdd.n3568 vdd.n3567 0.152939
R6708 vdd.n3567 vdd.n630 0.152939
R6709 vdd.n3585 vdd.n630 0.152939
R6710 vdd.n3586 vdd.n3585 0.152939
R6711 vdd.n3587 vdd.n3586 0.152939
R6712 vdd.n3587 vdd.n628 0.152939
R6713 vdd.n3592 vdd.n628 0.152939
R6714 vdd.n3593 vdd.n3592 0.152939
R6715 vdd.n3594 vdd.n3593 0.152939
R6716 vdd.n3594 vdd.n626 0.152939
R6717 vdd.n3599 vdd.n626 0.152939
R6718 vdd.n3600 vdd.n3599 0.152939
R6719 vdd.n3601 vdd.n3600 0.152939
R6720 vdd.n3601 vdd.n624 0.152939
R6721 vdd.n3607 vdd.n624 0.152939
R6722 vdd.n3608 vdd.n3607 0.152939
R6723 vdd.n3609 vdd.n3608 0.152939
R6724 vdd.n3609 vdd.n622 0.152939
R6725 vdd.n3614 vdd.n622 0.152939
R6726 vdd.n3615 vdd.n3614 0.152939
R6727 vdd.n3616 vdd.n3615 0.152939
R6728 vdd.n3616 vdd.n620 0.152939
R6729 vdd.n3621 vdd.n620 0.152939
R6730 vdd.n3498 vdd.n687 0.152939
R6731 vdd.n2366 vdd.n1517 0.152939
R6732 vdd.n1885 vdd.n1641 0.152939
R6733 vdd.n1886 vdd.n1885 0.152939
R6734 vdd.n1887 vdd.n1886 0.152939
R6735 vdd.n1887 vdd.n1629 0.152939
R6736 vdd.n1902 vdd.n1629 0.152939
R6737 vdd.n1903 vdd.n1902 0.152939
R6738 vdd.n1904 vdd.n1903 0.152939
R6739 vdd.n1904 vdd.n1619 0.152939
R6740 vdd.n1919 vdd.n1619 0.152939
R6741 vdd.n1920 vdd.n1919 0.152939
R6742 vdd.n1921 vdd.n1920 0.152939
R6743 vdd.n1921 vdd.n1606 0.152939
R6744 vdd.n1935 vdd.n1606 0.152939
R6745 vdd.n1936 vdd.n1935 0.152939
R6746 vdd.n1937 vdd.n1936 0.152939
R6747 vdd.n1937 vdd.n1595 0.152939
R6748 vdd.n1952 vdd.n1595 0.152939
R6749 vdd.n1953 vdd.n1952 0.152939
R6750 vdd.n1954 vdd.n1953 0.152939
R6751 vdd.n1954 vdd.n1584 0.152939
R6752 vdd.n2275 vdd.n1584 0.152939
R6753 vdd.n2276 vdd.n2275 0.152939
R6754 vdd.n2277 vdd.n2276 0.152939
R6755 vdd.n2277 vdd.n1572 0.152939
R6756 vdd.n2292 vdd.n1572 0.152939
R6757 vdd.n2293 vdd.n2292 0.152939
R6758 vdd.n2294 vdd.n2293 0.152939
R6759 vdd.n2294 vdd.n1562 0.152939
R6760 vdd.n2309 vdd.n1562 0.152939
R6761 vdd.n2310 vdd.n2309 0.152939
R6762 vdd.n2311 vdd.n2310 0.152939
R6763 vdd.n2311 vdd.n1549 0.152939
R6764 vdd.n2325 vdd.n1549 0.152939
R6765 vdd.n2326 vdd.n2325 0.152939
R6766 vdd.n2327 vdd.n2326 0.152939
R6767 vdd.n2327 vdd.n1539 0.152939
R6768 vdd.n2342 vdd.n1539 0.152939
R6769 vdd.n2343 vdd.n2342 0.152939
R6770 vdd.n2346 vdd.n2343 0.152939
R6771 vdd.n2346 vdd.n2345 0.152939
R6772 vdd.n2345 vdd.n2344 0.152939
R6773 vdd.n1877 vdd.n1646 0.152939
R6774 vdd.n1870 vdd.n1646 0.152939
R6775 vdd.n1870 vdd.n1869 0.152939
R6776 vdd.n1869 vdd.n1868 0.152939
R6777 vdd.n1868 vdd.n1683 0.152939
R6778 vdd.n1864 vdd.n1683 0.152939
R6779 vdd.n1864 vdd.n1863 0.152939
R6780 vdd.n1863 vdd.n1862 0.152939
R6781 vdd.n1862 vdd.n1689 0.152939
R6782 vdd.n1858 vdd.n1689 0.152939
R6783 vdd.n1858 vdd.n1857 0.152939
R6784 vdd.n1857 vdd.n1856 0.152939
R6785 vdd.n1856 vdd.n1695 0.152939
R6786 vdd.n1852 vdd.n1695 0.152939
R6787 vdd.n1852 vdd.n1851 0.152939
R6788 vdd.n1851 vdd.n1850 0.152939
R6789 vdd.n1850 vdd.n1701 0.152939
R6790 vdd.n1846 vdd.n1701 0.152939
R6791 vdd.n1846 vdd.n1845 0.152939
R6792 vdd.n1845 vdd.n1844 0.152939
R6793 vdd.n1844 vdd.n1709 0.152939
R6794 vdd.n1840 vdd.n1709 0.152939
R6795 vdd.n1840 vdd.n1839 0.152939
R6796 vdd.n1839 vdd.n1838 0.152939
R6797 vdd.n1838 vdd.n1715 0.152939
R6798 vdd.n1834 vdd.n1715 0.152939
R6799 vdd.n1834 vdd.n1833 0.152939
R6800 vdd.n1833 vdd.n1832 0.152939
R6801 vdd.n1832 vdd.n1721 0.152939
R6802 vdd.n1828 vdd.n1721 0.152939
R6803 vdd.n1828 vdd.n1827 0.152939
R6804 vdd.n1827 vdd.n1826 0.152939
R6805 vdd.n1826 vdd.n1727 0.152939
R6806 vdd.n1822 vdd.n1727 0.152939
R6807 vdd.n1822 vdd.n1821 0.152939
R6808 vdd.n1821 vdd.n1820 0.152939
R6809 vdd.n1820 vdd.n1733 0.152939
R6810 vdd.n1816 vdd.n1733 0.152939
R6811 vdd.n1816 vdd.n1815 0.152939
R6812 vdd.n1815 vdd.n1814 0.152939
R6813 vdd.n1814 vdd.n1739 0.152939
R6814 vdd.n1807 vdd.n1739 0.152939
R6815 vdd.n1807 vdd.n1806 0.152939
R6816 vdd.n1806 vdd.n1805 0.152939
R6817 vdd.n1805 vdd.n1744 0.152939
R6818 vdd.n1801 vdd.n1744 0.152939
R6819 vdd.n1801 vdd.n1800 0.152939
R6820 vdd.n1800 vdd.n1799 0.152939
R6821 vdd.n1799 vdd.n1750 0.152939
R6822 vdd.n1795 vdd.n1750 0.152939
R6823 vdd.n1795 vdd.n1794 0.152939
R6824 vdd.n1794 vdd.n1793 0.152939
R6825 vdd.n1793 vdd.n1756 0.152939
R6826 vdd.n1789 vdd.n1756 0.152939
R6827 vdd.n1789 vdd.n1788 0.152939
R6828 vdd.n1788 vdd.n1787 0.152939
R6829 vdd.n1787 vdd.n1762 0.152939
R6830 vdd.n1783 vdd.n1762 0.152939
R6831 vdd.n1783 vdd.n1782 0.152939
R6832 vdd.n1782 vdd.n1781 0.152939
R6833 vdd.n1781 vdd.n1768 0.152939
R6834 vdd.n1777 vdd.n1768 0.152939
R6835 vdd.n1777 vdd.n1776 0.152939
R6836 vdd.n1879 vdd.n1878 0.152939
R6837 vdd.n1879 vdd.n1635 0.152939
R6838 vdd.n1894 vdd.n1635 0.152939
R6839 vdd.n1895 vdd.n1894 0.152939
R6840 vdd.n1896 vdd.n1895 0.152939
R6841 vdd.n1896 vdd.n1624 0.152939
R6842 vdd.n1911 vdd.n1624 0.152939
R6843 vdd.n1912 vdd.n1911 0.152939
R6844 vdd.n1913 vdd.n1912 0.152939
R6845 vdd.n1913 vdd.n1613 0.152939
R6846 vdd.n1927 vdd.n1613 0.152939
R6847 vdd.n1928 vdd.n1927 0.152939
R6848 vdd.n1929 vdd.n1928 0.152939
R6849 vdd.n1929 vdd.n1601 0.152939
R6850 vdd.n1944 vdd.n1601 0.152939
R6851 vdd.n1945 vdd.n1944 0.152939
R6852 vdd.n1946 vdd.n1945 0.152939
R6853 vdd.n1946 vdd.n1590 0.152939
R6854 vdd.n1960 vdd.n1590 0.152939
R6855 vdd.n1961 vdd.n1960 0.152939
R6856 vdd.n1882 vdd.t296 0.113865
R6857 vdd.t245 vdd.n386 0.113865
R6858 vdd.n2474 vdd.n2473 0.110256
R6859 vdd.n3488 vdd.n727 0.110256
R6860 vdd.n3365 vdd.n687 0.110256
R6861 vdd.n2367 vdd.n2366 0.110256
R6862 vdd.n2269 vdd.n2268 0.0695946
R6863 vdd.n3671 vdd.n334 0.0695946
R6864 vdd.n3671 vdd.n3670 0.0695946
R6865 vdd.n2268 vdd.n1961 0.0695946
R6866 vdd.n2474 vdd.n1178 0.0431829
R6867 vdd.n2367 vdd.n1278 0.0431829
R6868 vdd.n3488 vdd.n730 0.0431829
R6869 vdd.n3365 vdd.n783 0.0431829
R6870 vdd vdd.n28 0.00833333
R6871 commonsourceibias.n35 commonsourceibias.t56 223.028
R6872 commonsourceibias.n128 commonsourceibias.t129 223.028
R6873 commonsourceibias.n307 commonsourceibias.t140 223.028
R6874 commonsourceibias.n217 commonsourceibias.t112 223.028
R6875 commonsourceibias.n454 commonsourceibias.t6 223.028
R6876 commonsourceibias.n395 commonsourceibias.t108 223.028
R6877 commonsourceibias.n679 commonsourceibias.t74 223.028
R6878 commonsourceibias.n589 commonsourceibias.t97 223.028
R6879 commonsourceibias.n99 commonsourceibias.t20 207.983
R6880 commonsourceibias.n192 commonsourceibias.t120 207.983
R6881 commonsourceibias.n371 commonsourceibias.t147 207.983
R6882 commonsourceibias.n281 commonsourceibias.t71 207.983
R6883 commonsourceibias.n520 commonsourceibias.t28 207.983
R6884 commonsourceibias.n566 commonsourceibias.t91 207.983
R6885 commonsourceibias.n745 commonsourceibias.t82 207.983
R6886 commonsourceibias.n655 commonsourceibias.t151 207.983
R6887 commonsourceibias.n97 commonsourceibias.t14 168.701
R6888 commonsourceibias.n91 commonsourceibias.t58 168.701
R6889 commonsourceibias.n17 commonsourceibias.t18 168.701
R6890 commonsourceibias.n83 commonsourceibias.t60 168.701
R6891 commonsourceibias.n77 commonsourceibias.t24 168.701
R6892 commonsourceibias.n22 commonsourceibias.t12 168.701
R6893 commonsourceibias.n69 commonsourceibias.t54 168.701
R6894 commonsourceibias.n63 commonsourceibias.t22 168.701
R6895 commonsourceibias.n25 commonsourceibias.t38 168.701
R6896 commonsourceibias.n27 commonsourceibias.t8 168.701
R6897 commonsourceibias.n29 commonsourceibias.t46 168.701
R6898 commonsourceibias.n46 commonsourceibias.t62 168.701
R6899 commonsourceibias.n40 commonsourceibias.t42 168.701
R6900 commonsourceibias.n34 commonsourceibias.t16 168.701
R6901 commonsourceibias.n190 commonsourceibias.t67 168.701
R6902 commonsourceibias.n184 commonsourceibias.t126 168.701
R6903 commonsourceibias.n5 commonsourceibias.t121 168.701
R6904 commonsourceibias.n176 commonsourceibias.t136 168.701
R6905 commonsourceibias.n170 commonsourceibias.t117 168.701
R6906 commonsourceibias.n10 commonsourceibias.t102 168.701
R6907 commonsourceibias.n162 commonsourceibias.t125 168.701
R6908 commonsourceibias.n156 commonsourceibias.t118 168.701
R6909 commonsourceibias.n118 commonsourceibias.t76 168.701
R6910 commonsourceibias.n120 commonsourceibias.t106 168.701
R6911 commonsourceibias.n122 commonsourceibias.t96 168.701
R6912 commonsourceibias.n139 commonsourceibias.t141 168.701
R6913 commonsourceibias.n133 commonsourceibias.t116 168.701
R6914 commonsourceibias.n127 commonsourceibias.t152 168.701
R6915 commonsourceibias.n306 commonsourceibias.t130 168.701
R6916 commonsourceibias.n312 commonsourceibias.t79 168.701
R6917 commonsourceibias.n318 commonsourceibias.t149 168.701
R6918 commonsourceibias.n301 commonsourceibias.t133 168.701
R6919 commonsourceibias.n299 commonsourceibias.t137 168.701
R6920 commonsourceibias.n297 commonsourceibias.t64 168.701
R6921 commonsourceibias.n335 commonsourceibias.t138 168.701
R6922 commonsourceibias.n341 commonsourceibias.t146 168.701
R6923 commonsourceibias.n294 commonsourceibias.t119 168.701
R6924 commonsourceibias.n349 commonsourceibias.t90 168.701
R6925 commonsourceibias.n355 commonsourceibias.t155 168.701
R6926 commonsourceibias.n289 commonsourceibias.t124 168.701
R6927 commonsourceibias.n363 commonsourceibias.t128 168.701
R6928 commonsourceibias.n369 commonsourceibias.t75 168.701
R6929 commonsourceibias.n279 commonsourceibias.t159 168.701
R6930 commonsourceibias.n273 commonsourceibias.t148 168.701
R6931 commonsourceibias.n199 commonsourceibias.t78 168.701
R6932 commonsourceibias.n265 commonsourceibias.t157 168.701
R6933 commonsourceibias.n259 commonsourceibias.t85 168.701
R6934 commonsourceibias.n204 commonsourceibias.t77 168.701
R6935 commonsourceibias.n251 commonsourceibias.t158 168.701
R6936 commonsourceibias.n245 commonsourceibias.t94 168.701
R6937 commonsourceibias.n207 commonsourceibias.t113 168.701
R6938 commonsourceibias.n209 commonsourceibias.t156 168.701
R6939 commonsourceibias.n211 commonsourceibias.t92 168.701
R6940 commonsourceibias.n228 commonsourceibias.t111 168.701
R6941 commonsourceibias.n222 commonsourceibias.t105 168.701
R6942 commonsourceibias.n216 commonsourceibias.t93 168.701
R6943 commonsourceibias.n453 commonsourceibias.t50 168.701
R6944 commonsourceibias.n459 commonsourceibias.t36 168.701
R6945 commonsourceibias.n465 commonsourceibias.t52 168.701
R6946 commonsourceibias.n448 commonsourceibias.t0 168.701
R6947 commonsourceibias.n446 commonsourceibias.t34 168.701
R6948 commonsourceibias.n444 commonsourceibias.t2 168.701
R6949 commonsourceibias.n482 commonsourceibias.t30 168.701
R6950 commonsourceibias.n488 commonsourceibias.t10 168.701
R6951 commonsourceibias.n490 commonsourceibias.t40 168.701
R6952 commonsourceibias.n497 commonsourceibias.t32 168.701
R6953 commonsourceibias.n503 commonsourceibias.t4 168.701
R6954 commonsourceibias.n505 commonsourceibias.t26 168.701
R6955 commonsourceibias.n512 commonsourceibias.t44 168.701
R6956 commonsourceibias.n518 commonsourceibias.t48 168.701
R6957 commonsourceibias.n564 commonsourceibias.t134 168.701
R6958 commonsourceibias.n558 commonsourceibias.t114 168.701
R6959 commonsourceibias.n551 commonsourceibias.t95 168.701
R6960 commonsourceibias.n549 commonsourceibias.t123 168.701
R6961 commonsourceibias.n543 commonsourceibias.t88 168.701
R6962 commonsourceibias.n536 commonsourceibias.t73 168.701
R6963 commonsourceibias.n534 commonsourceibias.t104 168.701
R6964 commonsourceibias.n394 commonsourceibias.t131 168.701
R6965 commonsourceibias.n400 commonsourceibias.t84 168.701
R6966 commonsourceibias.n406 commonsourceibias.t127 168.701
R6967 commonsourceibias.n389 commonsourceibias.t150 168.701
R6968 commonsourceibias.n387 commonsourceibias.t83 168.701
R6969 commonsourceibias.n385 commonsourceibias.t139 168.701
R6970 commonsourceibias.n423 commonsourceibias.t89 168.701
R6971 commonsourceibias.n678 commonsourceibias.t145 168.701
R6972 commonsourceibias.n684 commonsourceibias.t109 168.701
R6973 commonsourceibias.n690 commonsourceibias.t87 168.701
R6974 commonsourceibias.n673 commonsourceibias.t153 168.701
R6975 commonsourceibias.n671 commonsourceibias.t132 168.701
R6976 commonsourceibias.n669 commonsourceibias.t103 168.701
R6977 commonsourceibias.n707 commonsourceibias.t70 168.701
R6978 commonsourceibias.n713 commonsourceibias.t81 168.701
R6979 commonsourceibias.n715 commonsourceibias.t110 168.701
R6980 commonsourceibias.n722 commonsourceibias.t115 168.701
R6981 commonsourceibias.n728 commonsourceibias.t101 168.701
R6982 commonsourceibias.n730 commonsourceibias.t135 168.701
R6983 commonsourceibias.n737 commonsourceibias.t122 168.701
R6984 commonsourceibias.n743 commonsourceibias.t107 168.701
R6985 commonsourceibias.n588 commonsourceibias.t68 168.701
R6986 commonsourceibias.n594 commonsourceibias.t86 168.701
R6987 commonsourceibias.n600 commonsourceibias.t98 168.701
R6988 commonsourceibias.n583 commonsourceibias.t69 168.701
R6989 commonsourceibias.n581 commonsourceibias.t80 168.701
R6990 commonsourceibias.n579 commonsourceibias.t99 168.701
R6991 commonsourceibias.n617 commonsourceibias.t72 168.701
R6992 commonsourceibias.n623 commonsourceibias.t142 168.701
R6993 commonsourceibias.n625 commonsourceibias.t100 168.701
R6994 commonsourceibias.n632 commonsourceibias.t65 168.701
R6995 commonsourceibias.n638 commonsourceibias.t143 168.701
R6996 commonsourceibias.n640 commonsourceibias.t154 168.701
R6997 commonsourceibias.n647 commonsourceibias.t66 168.701
R6998 commonsourceibias.n653 commonsourceibias.t144 168.701
R6999 commonsourceibias.n36 commonsourceibias.n33 161.3
R7000 commonsourceibias.n38 commonsourceibias.n37 161.3
R7001 commonsourceibias.n39 commonsourceibias.n32 161.3
R7002 commonsourceibias.n42 commonsourceibias.n41 161.3
R7003 commonsourceibias.n43 commonsourceibias.n31 161.3
R7004 commonsourceibias.n45 commonsourceibias.n44 161.3
R7005 commonsourceibias.n47 commonsourceibias.n30 161.3
R7006 commonsourceibias.n49 commonsourceibias.n48 161.3
R7007 commonsourceibias.n51 commonsourceibias.n50 161.3
R7008 commonsourceibias.n52 commonsourceibias.n28 161.3
R7009 commonsourceibias.n54 commonsourceibias.n53 161.3
R7010 commonsourceibias.n56 commonsourceibias.n55 161.3
R7011 commonsourceibias.n57 commonsourceibias.n26 161.3
R7012 commonsourceibias.n59 commonsourceibias.n58 161.3
R7013 commonsourceibias.n61 commonsourceibias.n60 161.3
R7014 commonsourceibias.n62 commonsourceibias.n24 161.3
R7015 commonsourceibias.n65 commonsourceibias.n64 161.3
R7016 commonsourceibias.n66 commonsourceibias.n23 161.3
R7017 commonsourceibias.n68 commonsourceibias.n67 161.3
R7018 commonsourceibias.n70 commonsourceibias.n21 161.3
R7019 commonsourceibias.n72 commonsourceibias.n71 161.3
R7020 commonsourceibias.n73 commonsourceibias.n20 161.3
R7021 commonsourceibias.n75 commonsourceibias.n74 161.3
R7022 commonsourceibias.n76 commonsourceibias.n19 161.3
R7023 commonsourceibias.n79 commonsourceibias.n78 161.3
R7024 commonsourceibias.n80 commonsourceibias.n18 161.3
R7025 commonsourceibias.n82 commonsourceibias.n81 161.3
R7026 commonsourceibias.n84 commonsourceibias.n16 161.3
R7027 commonsourceibias.n86 commonsourceibias.n85 161.3
R7028 commonsourceibias.n87 commonsourceibias.n15 161.3
R7029 commonsourceibias.n89 commonsourceibias.n88 161.3
R7030 commonsourceibias.n90 commonsourceibias.n14 161.3
R7031 commonsourceibias.n93 commonsourceibias.n92 161.3
R7032 commonsourceibias.n94 commonsourceibias.n13 161.3
R7033 commonsourceibias.n96 commonsourceibias.n95 161.3
R7034 commonsourceibias.n98 commonsourceibias.n12 161.3
R7035 commonsourceibias.n129 commonsourceibias.n126 161.3
R7036 commonsourceibias.n131 commonsourceibias.n130 161.3
R7037 commonsourceibias.n132 commonsourceibias.n125 161.3
R7038 commonsourceibias.n135 commonsourceibias.n134 161.3
R7039 commonsourceibias.n136 commonsourceibias.n124 161.3
R7040 commonsourceibias.n138 commonsourceibias.n137 161.3
R7041 commonsourceibias.n140 commonsourceibias.n123 161.3
R7042 commonsourceibias.n142 commonsourceibias.n141 161.3
R7043 commonsourceibias.n144 commonsourceibias.n143 161.3
R7044 commonsourceibias.n145 commonsourceibias.n121 161.3
R7045 commonsourceibias.n147 commonsourceibias.n146 161.3
R7046 commonsourceibias.n149 commonsourceibias.n148 161.3
R7047 commonsourceibias.n150 commonsourceibias.n119 161.3
R7048 commonsourceibias.n152 commonsourceibias.n151 161.3
R7049 commonsourceibias.n154 commonsourceibias.n153 161.3
R7050 commonsourceibias.n155 commonsourceibias.n117 161.3
R7051 commonsourceibias.n158 commonsourceibias.n157 161.3
R7052 commonsourceibias.n159 commonsourceibias.n11 161.3
R7053 commonsourceibias.n161 commonsourceibias.n160 161.3
R7054 commonsourceibias.n163 commonsourceibias.n9 161.3
R7055 commonsourceibias.n165 commonsourceibias.n164 161.3
R7056 commonsourceibias.n166 commonsourceibias.n8 161.3
R7057 commonsourceibias.n168 commonsourceibias.n167 161.3
R7058 commonsourceibias.n169 commonsourceibias.n7 161.3
R7059 commonsourceibias.n172 commonsourceibias.n171 161.3
R7060 commonsourceibias.n173 commonsourceibias.n6 161.3
R7061 commonsourceibias.n175 commonsourceibias.n174 161.3
R7062 commonsourceibias.n177 commonsourceibias.n4 161.3
R7063 commonsourceibias.n179 commonsourceibias.n178 161.3
R7064 commonsourceibias.n180 commonsourceibias.n3 161.3
R7065 commonsourceibias.n182 commonsourceibias.n181 161.3
R7066 commonsourceibias.n183 commonsourceibias.n2 161.3
R7067 commonsourceibias.n186 commonsourceibias.n185 161.3
R7068 commonsourceibias.n187 commonsourceibias.n1 161.3
R7069 commonsourceibias.n189 commonsourceibias.n188 161.3
R7070 commonsourceibias.n191 commonsourceibias.n0 161.3
R7071 commonsourceibias.n370 commonsourceibias.n284 161.3
R7072 commonsourceibias.n368 commonsourceibias.n367 161.3
R7073 commonsourceibias.n366 commonsourceibias.n285 161.3
R7074 commonsourceibias.n365 commonsourceibias.n364 161.3
R7075 commonsourceibias.n362 commonsourceibias.n286 161.3
R7076 commonsourceibias.n361 commonsourceibias.n360 161.3
R7077 commonsourceibias.n359 commonsourceibias.n287 161.3
R7078 commonsourceibias.n358 commonsourceibias.n357 161.3
R7079 commonsourceibias.n356 commonsourceibias.n288 161.3
R7080 commonsourceibias.n354 commonsourceibias.n353 161.3
R7081 commonsourceibias.n352 commonsourceibias.n290 161.3
R7082 commonsourceibias.n351 commonsourceibias.n350 161.3
R7083 commonsourceibias.n348 commonsourceibias.n291 161.3
R7084 commonsourceibias.n347 commonsourceibias.n346 161.3
R7085 commonsourceibias.n345 commonsourceibias.n292 161.3
R7086 commonsourceibias.n344 commonsourceibias.n343 161.3
R7087 commonsourceibias.n342 commonsourceibias.n293 161.3
R7088 commonsourceibias.n340 commonsourceibias.n339 161.3
R7089 commonsourceibias.n338 commonsourceibias.n295 161.3
R7090 commonsourceibias.n337 commonsourceibias.n336 161.3
R7091 commonsourceibias.n334 commonsourceibias.n296 161.3
R7092 commonsourceibias.n333 commonsourceibias.n332 161.3
R7093 commonsourceibias.n331 commonsourceibias.n330 161.3
R7094 commonsourceibias.n329 commonsourceibias.n298 161.3
R7095 commonsourceibias.n328 commonsourceibias.n327 161.3
R7096 commonsourceibias.n326 commonsourceibias.n325 161.3
R7097 commonsourceibias.n324 commonsourceibias.n300 161.3
R7098 commonsourceibias.n323 commonsourceibias.n322 161.3
R7099 commonsourceibias.n321 commonsourceibias.n320 161.3
R7100 commonsourceibias.n319 commonsourceibias.n302 161.3
R7101 commonsourceibias.n317 commonsourceibias.n316 161.3
R7102 commonsourceibias.n315 commonsourceibias.n303 161.3
R7103 commonsourceibias.n314 commonsourceibias.n313 161.3
R7104 commonsourceibias.n311 commonsourceibias.n304 161.3
R7105 commonsourceibias.n310 commonsourceibias.n309 161.3
R7106 commonsourceibias.n308 commonsourceibias.n305 161.3
R7107 commonsourceibias.n218 commonsourceibias.n215 161.3
R7108 commonsourceibias.n220 commonsourceibias.n219 161.3
R7109 commonsourceibias.n221 commonsourceibias.n214 161.3
R7110 commonsourceibias.n224 commonsourceibias.n223 161.3
R7111 commonsourceibias.n225 commonsourceibias.n213 161.3
R7112 commonsourceibias.n227 commonsourceibias.n226 161.3
R7113 commonsourceibias.n229 commonsourceibias.n212 161.3
R7114 commonsourceibias.n231 commonsourceibias.n230 161.3
R7115 commonsourceibias.n233 commonsourceibias.n232 161.3
R7116 commonsourceibias.n234 commonsourceibias.n210 161.3
R7117 commonsourceibias.n236 commonsourceibias.n235 161.3
R7118 commonsourceibias.n238 commonsourceibias.n237 161.3
R7119 commonsourceibias.n239 commonsourceibias.n208 161.3
R7120 commonsourceibias.n241 commonsourceibias.n240 161.3
R7121 commonsourceibias.n243 commonsourceibias.n242 161.3
R7122 commonsourceibias.n244 commonsourceibias.n206 161.3
R7123 commonsourceibias.n247 commonsourceibias.n246 161.3
R7124 commonsourceibias.n248 commonsourceibias.n205 161.3
R7125 commonsourceibias.n250 commonsourceibias.n249 161.3
R7126 commonsourceibias.n252 commonsourceibias.n203 161.3
R7127 commonsourceibias.n254 commonsourceibias.n253 161.3
R7128 commonsourceibias.n255 commonsourceibias.n202 161.3
R7129 commonsourceibias.n257 commonsourceibias.n256 161.3
R7130 commonsourceibias.n258 commonsourceibias.n201 161.3
R7131 commonsourceibias.n261 commonsourceibias.n260 161.3
R7132 commonsourceibias.n262 commonsourceibias.n200 161.3
R7133 commonsourceibias.n264 commonsourceibias.n263 161.3
R7134 commonsourceibias.n266 commonsourceibias.n198 161.3
R7135 commonsourceibias.n268 commonsourceibias.n267 161.3
R7136 commonsourceibias.n269 commonsourceibias.n197 161.3
R7137 commonsourceibias.n271 commonsourceibias.n270 161.3
R7138 commonsourceibias.n272 commonsourceibias.n196 161.3
R7139 commonsourceibias.n275 commonsourceibias.n274 161.3
R7140 commonsourceibias.n276 commonsourceibias.n195 161.3
R7141 commonsourceibias.n278 commonsourceibias.n277 161.3
R7142 commonsourceibias.n280 commonsourceibias.n194 161.3
R7143 commonsourceibias.n519 commonsourceibias.n433 161.3
R7144 commonsourceibias.n517 commonsourceibias.n516 161.3
R7145 commonsourceibias.n515 commonsourceibias.n434 161.3
R7146 commonsourceibias.n514 commonsourceibias.n513 161.3
R7147 commonsourceibias.n511 commonsourceibias.n435 161.3
R7148 commonsourceibias.n510 commonsourceibias.n509 161.3
R7149 commonsourceibias.n508 commonsourceibias.n436 161.3
R7150 commonsourceibias.n507 commonsourceibias.n506 161.3
R7151 commonsourceibias.n504 commonsourceibias.n437 161.3
R7152 commonsourceibias.n502 commonsourceibias.n501 161.3
R7153 commonsourceibias.n500 commonsourceibias.n438 161.3
R7154 commonsourceibias.n499 commonsourceibias.n498 161.3
R7155 commonsourceibias.n496 commonsourceibias.n439 161.3
R7156 commonsourceibias.n495 commonsourceibias.n494 161.3
R7157 commonsourceibias.n493 commonsourceibias.n440 161.3
R7158 commonsourceibias.n492 commonsourceibias.n491 161.3
R7159 commonsourceibias.n489 commonsourceibias.n441 161.3
R7160 commonsourceibias.n487 commonsourceibias.n486 161.3
R7161 commonsourceibias.n485 commonsourceibias.n442 161.3
R7162 commonsourceibias.n484 commonsourceibias.n483 161.3
R7163 commonsourceibias.n481 commonsourceibias.n443 161.3
R7164 commonsourceibias.n480 commonsourceibias.n479 161.3
R7165 commonsourceibias.n478 commonsourceibias.n477 161.3
R7166 commonsourceibias.n476 commonsourceibias.n445 161.3
R7167 commonsourceibias.n475 commonsourceibias.n474 161.3
R7168 commonsourceibias.n473 commonsourceibias.n472 161.3
R7169 commonsourceibias.n471 commonsourceibias.n447 161.3
R7170 commonsourceibias.n470 commonsourceibias.n469 161.3
R7171 commonsourceibias.n468 commonsourceibias.n467 161.3
R7172 commonsourceibias.n466 commonsourceibias.n449 161.3
R7173 commonsourceibias.n464 commonsourceibias.n463 161.3
R7174 commonsourceibias.n462 commonsourceibias.n450 161.3
R7175 commonsourceibias.n461 commonsourceibias.n460 161.3
R7176 commonsourceibias.n458 commonsourceibias.n451 161.3
R7177 commonsourceibias.n457 commonsourceibias.n456 161.3
R7178 commonsourceibias.n455 commonsourceibias.n452 161.3
R7179 commonsourceibias.n425 commonsourceibias.n424 161.3
R7180 commonsourceibias.n422 commonsourceibias.n384 161.3
R7181 commonsourceibias.n421 commonsourceibias.n420 161.3
R7182 commonsourceibias.n419 commonsourceibias.n418 161.3
R7183 commonsourceibias.n417 commonsourceibias.n386 161.3
R7184 commonsourceibias.n416 commonsourceibias.n415 161.3
R7185 commonsourceibias.n414 commonsourceibias.n413 161.3
R7186 commonsourceibias.n412 commonsourceibias.n388 161.3
R7187 commonsourceibias.n411 commonsourceibias.n410 161.3
R7188 commonsourceibias.n409 commonsourceibias.n408 161.3
R7189 commonsourceibias.n407 commonsourceibias.n390 161.3
R7190 commonsourceibias.n405 commonsourceibias.n404 161.3
R7191 commonsourceibias.n403 commonsourceibias.n391 161.3
R7192 commonsourceibias.n402 commonsourceibias.n401 161.3
R7193 commonsourceibias.n399 commonsourceibias.n392 161.3
R7194 commonsourceibias.n398 commonsourceibias.n397 161.3
R7195 commonsourceibias.n396 commonsourceibias.n393 161.3
R7196 commonsourceibias.n531 commonsourceibias.n383 161.3
R7197 commonsourceibias.n565 commonsourceibias.n374 161.3
R7198 commonsourceibias.n563 commonsourceibias.n562 161.3
R7199 commonsourceibias.n561 commonsourceibias.n375 161.3
R7200 commonsourceibias.n560 commonsourceibias.n559 161.3
R7201 commonsourceibias.n557 commonsourceibias.n376 161.3
R7202 commonsourceibias.n556 commonsourceibias.n555 161.3
R7203 commonsourceibias.n554 commonsourceibias.n377 161.3
R7204 commonsourceibias.n553 commonsourceibias.n552 161.3
R7205 commonsourceibias.n550 commonsourceibias.n378 161.3
R7206 commonsourceibias.n548 commonsourceibias.n547 161.3
R7207 commonsourceibias.n546 commonsourceibias.n379 161.3
R7208 commonsourceibias.n545 commonsourceibias.n544 161.3
R7209 commonsourceibias.n542 commonsourceibias.n380 161.3
R7210 commonsourceibias.n541 commonsourceibias.n540 161.3
R7211 commonsourceibias.n539 commonsourceibias.n381 161.3
R7212 commonsourceibias.n538 commonsourceibias.n537 161.3
R7213 commonsourceibias.n535 commonsourceibias.n382 161.3
R7214 commonsourceibias.n533 commonsourceibias.n532 161.3
R7215 commonsourceibias.n744 commonsourceibias.n658 161.3
R7216 commonsourceibias.n742 commonsourceibias.n741 161.3
R7217 commonsourceibias.n740 commonsourceibias.n659 161.3
R7218 commonsourceibias.n739 commonsourceibias.n738 161.3
R7219 commonsourceibias.n736 commonsourceibias.n660 161.3
R7220 commonsourceibias.n735 commonsourceibias.n734 161.3
R7221 commonsourceibias.n733 commonsourceibias.n661 161.3
R7222 commonsourceibias.n732 commonsourceibias.n731 161.3
R7223 commonsourceibias.n729 commonsourceibias.n662 161.3
R7224 commonsourceibias.n727 commonsourceibias.n726 161.3
R7225 commonsourceibias.n725 commonsourceibias.n663 161.3
R7226 commonsourceibias.n724 commonsourceibias.n723 161.3
R7227 commonsourceibias.n721 commonsourceibias.n664 161.3
R7228 commonsourceibias.n720 commonsourceibias.n719 161.3
R7229 commonsourceibias.n718 commonsourceibias.n665 161.3
R7230 commonsourceibias.n717 commonsourceibias.n716 161.3
R7231 commonsourceibias.n714 commonsourceibias.n666 161.3
R7232 commonsourceibias.n712 commonsourceibias.n711 161.3
R7233 commonsourceibias.n710 commonsourceibias.n667 161.3
R7234 commonsourceibias.n709 commonsourceibias.n708 161.3
R7235 commonsourceibias.n706 commonsourceibias.n668 161.3
R7236 commonsourceibias.n705 commonsourceibias.n704 161.3
R7237 commonsourceibias.n703 commonsourceibias.n702 161.3
R7238 commonsourceibias.n701 commonsourceibias.n670 161.3
R7239 commonsourceibias.n700 commonsourceibias.n699 161.3
R7240 commonsourceibias.n698 commonsourceibias.n697 161.3
R7241 commonsourceibias.n696 commonsourceibias.n672 161.3
R7242 commonsourceibias.n695 commonsourceibias.n694 161.3
R7243 commonsourceibias.n693 commonsourceibias.n692 161.3
R7244 commonsourceibias.n691 commonsourceibias.n674 161.3
R7245 commonsourceibias.n689 commonsourceibias.n688 161.3
R7246 commonsourceibias.n687 commonsourceibias.n675 161.3
R7247 commonsourceibias.n686 commonsourceibias.n685 161.3
R7248 commonsourceibias.n683 commonsourceibias.n676 161.3
R7249 commonsourceibias.n682 commonsourceibias.n681 161.3
R7250 commonsourceibias.n680 commonsourceibias.n677 161.3
R7251 commonsourceibias.n654 commonsourceibias.n568 161.3
R7252 commonsourceibias.n652 commonsourceibias.n651 161.3
R7253 commonsourceibias.n650 commonsourceibias.n569 161.3
R7254 commonsourceibias.n649 commonsourceibias.n648 161.3
R7255 commonsourceibias.n646 commonsourceibias.n570 161.3
R7256 commonsourceibias.n645 commonsourceibias.n644 161.3
R7257 commonsourceibias.n643 commonsourceibias.n571 161.3
R7258 commonsourceibias.n642 commonsourceibias.n641 161.3
R7259 commonsourceibias.n639 commonsourceibias.n572 161.3
R7260 commonsourceibias.n637 commonsourceibias.n636 161.3
R7261 commonsourceibias.n635 commonsourceibias.n573 161.3
R7262 commonsourceibias.n634 commonsourceibias.n633 161.3
R7263 commonsourceibias.n631 commonsourceibias.n574 161.3
R7264 commonsourceibias.n630 commonsourceibias.n629 161.3
R7265 commonsourceibias.n628 commonsourceibias.n575 161.3
R7266 commonsourceibias.n627 commonsourceibias.n626 161.3
R7267 commonsourceibias.n624 commonsourceibias.n576 161.3
R7268 commonsourceibias.n622 commonsourceibias.n621 161.3
R7269 commonsourceibias.n620 commonsourceibias.n577 161.3
R7270 commonsourceibias.n619 commonsourceibias.n618 161.3
R7271 commonsourceibias.n616 commonsourceibias.n578 161.3
R7272 commonsourceibias.n615 commonsourceibias.n614 161.3
R7273 commonsourceibias.n613 commonsourceibias.n612 161.3
R7274 commonsourceibias.n611 commonsourceibias.n580 161.3
R7275 commonsourceibias.n610 commonsourceibias.n609 161.3
R7276 commonsourceibias.n608 commonsourceibias.n607 161.3
R7277 commonsourceibias.n606 commonsourceibias.n582 161.3
R7278 commonsourceibias.n605 commonsourceibias.n604 161.3
R7279 commonsourceibias.n603 commonsourceibias.n602 161.3
R7280 commonsourceibias.n601 commonsourceibias.n584 161.3
R7281 commonsourceibias.n599 commonsourceibias.n598 161.3
R7282 commonsourceibias.n597 commonsourceibias.n585 161.3
R7283 commonsourceibias.n596 commonsourceibias.n595 161.3
R7284 commonsourceibias.n593 commonsourceibias.n586 161.3
R7285 commonsourceibias.n592 commonsourceibias.n591 161.3
R7286 commonsourceibias.n590 commonsourceibias.n587 161.3
R7287 commonsourceibias.n111 commonsourceibias.n109 81.5057
R7288 commonsourceibias.n428 commonsourceibias.n426 81.5057
R7289 commonsourceibias.n111 commonsourceibias.n110 80.9324
R7290 commonsourceibias.n113 commonsourceibias.n112 80.9324
R7291 commonsourceibias.n115 commonsourceibias.n114 80.9324
R7292 commonsourceibias.n108 commonsourceibias.n107 80.9324
R7293 commonsourceibias.n106 commonsourceibias.n105 80.9324
R7294 commonsourceibias.n104 commonsourceibias.n103 80.9324
R7295 commonsourceibias.n102 commonsourceibias.n101 80.9324
R7296 commonsourceibias.n523 commonsourceibias.n522 80.9324
R7297 commonsourceibias.n525 commonsourceibias.n524 80.9324
R7298 commonsourceibias.n527 commonsourceibias.n526 80.9324
R7299 commonsourceibias.n529 commonsourceibias.n528 80.9324
R7300 commonsourceibias.n432 commonsourceibias.n431 80.9324
R7301 commonsourceibias.n430 commonsourceibias.n429 80.9324
R7302 commonsourceibias.n428 commonsourceibias.n427 80.9324
R7303 commonsourceibias.n100 commonsourceibias.n99 80.6037
R7304 commonsourceibias.n193 commonsourceibias.n192 80.6037
R7305 commonsourceibias.n372 commonsourceibias.n371 80.6037
R7306 commonsourceibias.n282 commonsourceibias.n281 80.6037
R7307 commonsourceibias.n521 commonsourceibias.n520 80.6037
R7308 commonsourceibias.n567 commonsourceibias.n566 80.6037
R7309 commonsourceibias.n746 commonsourceibias.n745 80.6037
R7310 commonsourceibias.n656 commonsourceibias.n655 80.6037
R7311 commonsourceibias.n85 commonsourceibias.n84 56.5617
R7312 commonsourceibias.n71 commonsourceibias.n70 56.5617
R7313 commonsourceibias.n62 commonsourceibias.n61 56.5617
R7314 commonsourceibias.n48 commonsourceibias.n47 56.5617
R7315 commonsourceibias.n178 commonsourceibias.n177 56.5617
R7316 commonsourceibias.n164 commonsourceibias.n163 56.5617
R7317 commonsourceibias.n155 commonsourceibias.n154 56.5617
R7318 commonsourceibias.n141 commonsourceibias.n140 56.5617
R7319 commonsourceibias.n320 commonsourceibias.n319 56.5617
R7320 commonsourceibias.n334 commonsourceibias.n333 56.5617
R7321 commonsourceibias.n343 commonsourceibias.n342 56.5617
R7322 commonsourceibias.n357 commonsourceibias.n356 56.5617
R7323 commonsourceibias.n267 commonsourceibias.n266 56.5617
R7324 commonsourceibias.n253 commonsourceibias.n252 56.5617
R7325 commonsourceibias.n244 commonsourceibias.n243 56.5617
R7326 commonsourceibias.n230 commonsourceibias.n229 56.5617
R7327 commonsourceibias.n467 commonsourceibias.n466 56.5617
R7328 commonsourceibias.n481 commonsourceibias.n480 56.5617
R7329 commonsourceibias.n491 commonsourceibias.n489 56.5617
R7330 commonsourceibias.n506 commonsourceibias.n504 56.5617
R7331 commonsourceibias.n552 commonsourceibias.n550 56.5617
R7332 commonsourceibias.n537 commonsourceibias.n535 56.5617
R7333 commonsourceibias.n408 commonsourceibias.n407 56.5617
R7334 commonsourceibias.n422 commonsourceibias.n421 56.5617
R7335 commonsourceibias.n692 commonsourceibias.n691 56.5617
R7336 commonsourceibias.n706 commonsourceibias.n705 56.5617
R7337 commonsourceibias.n716 commonsourceibias.n714 56.5617
R7338 commonsourceibias.n731 commonsourceibias.n729 56.5617
R7339 commonsourceibias.n602 commonsourceibias.n601 56.5617
R7340 commonsourceibias.n616 commonsourceibias.n615 56.5617
R7341 commonsourceibias.n626 commonsourceibias.n624 56.5617
R7342 commonsourceibias.n641 commonsourceibias.n639 56.5617
R7343 commonsourceibias.n76 commonsourceibias.n75 56.0773
R7344 commonsourceibias.n57 commonsourceibias.n56 56.0773
R7345 commonsourceibias.n169 commonsourceibias.n168 56.0773
R7346 commonsourceibias.n150 commonsourceibias.n149 56.0773
R7347 commonsourceibias.n329 commonsourceibias.n328 56.0773
R7348 commonsourceibias.n348 commonsourceibias.n347 56.0773
R7349 commonsourceibias.n258 commonsourceibias.n257 56.0773
R7350 commonsourceibias.n239 commonsourceibias.n238 56.0773
R7351 commonsourceibias.n476 commonsourceibias.n475 56.0773
R7352 commonsourceibias.n496 commonsourceibias.n495 56.0773
R7353 commonsourceibias.n542 commonsourceibias.n541 56.0773
R7354 commonsourceibias.n417 commonsourceibias.n416 56.0773
R7355 commonsourceibias.n701 commonsourceibias.n700 56.0773
R7356 commonsourceibias.n721 commonsourceibias.n720 56.0773
R7357 commonsourceibias.n611 commonsourceibias.n610 56.0773
R7358 commonsourceibias.n631 commonsourceibias.n630 56.0773
R7359 commonsourceibias.n99 commonsourceibias.n98 55.3321
R7360 commonsourceibias.n192 commonsourceibias.n191 55.3321
R7361 commonsourceibias.n371 commonsourceibias.n370 55.3321
R7362 commonsourceibias.n281 commonsourceibias.n280 55.3321
R7363 commonsourceibias.n520 commonsourceibias.n519 55.3321
R7364 commonsourceibias.n566 commonsourceibias.n565 55.3321
R7365 commonsourceibias.n745 commonsourceibias.n744 55.3321
R7366 commonsourceibias.n655 commonsourceibias.n654 55.3321
R7367 commonsourceibias.n90 commonsourceibias.n89 55.1086
R7368 commonsourceibias.n41 commonsourceibias.n31 55.1086
R7369 commonsourceibias.n183 commonsourceibias.n182 55.1086
R7370 commonsourceibias.n134 commonsourceibias.n124 55.1086
R7371 commonsourceibias.n313 commonsourceibias.n303 55.1086
R7372 commonsourceibias.n362 commonsourceibias.n361 55.1086
R7373 commonsourceibias.n272 commonsourceibias.n271 55.1086
R7374 commonsourceibias.n223 commonsourceibias.n213 55.1086
R7375 commonsourceibias.n460 commonsourceibias.n450 55.1086
R7376 commonsourceibias.n511 commonsourceibias.n510 55.1086
R7377 commonsourceibias.n557 commonsourceibias.n556 55.1086
R7378 commonsourceibias.n401 commonsourceibias.n391 55.1086
R7379 commonsourceibias.n685 commonsourceibias.n675 55.1086
R7380 commonsourceibias.n736 commonsourceibias.n735 55.1086
R7381 commonsourceibias.n595 commonsourceibias.n585 55.1086
R7382 commonsourceibias.n646 commonsourceibias.n645 55.1086
R7383 commonsourceibias.n35 commonsourceibias.n34 47.4592
R7384 commonsourceibias.n128 commonsourceibias.n127 47.4592
R7385 commonsourceibias.n307 commonsourceibias.n306 47.4592
R7386 commonsourceibias.n217 commonsourceibias.n216 47.4592
R7387 commonsourceibias.n454 commonsourceibias.n453 47.4592
R7388 commonsourceibias.n395 commonsourceibias.n394 47.4592
R7389 commonsourceibias.n679 commonsourceibias.n678 47.4592
R7390 commonsourceibias.n589 commonsourceibias.n588 47.4592
R7391 commonsourceibias.n308 commonsourceibias.n307 44.0436
R7392 commonsourceibias.n455 commonsourceibias.n454 44.0436
R7393 commonsourceibias.n396 commonsourceibias.n395 44.0436
R7394 commonsourceibias.n680 commonsourceibias.n679 44.0436
R7395 commonsourceibias.n590 commonsourceibias.n589 44.0436
R7396 commonsourceibias.n36 commonsourceibias.n35 44.0436
R7397 commonsourceibias.n129 commonsourceibias.n128 44.0436
R7398 commonsourceibias.n218 commonsourceibias.n217 44.0436
R7399 commonsourceibias.n92 commonsourceibias.n13 42.5146
R7400 commonsourceibias.n39 commonsourceibias.n38 42.5146
R7401 commonsourceibias.n185 commonsourceibias.n1 42.5146
R7402 commonsourceibias.n132 commonsourceibias.n131 42.5146
R7403 commonsourceibias.n311 commonsourceibias.n310 42.5146
R7404 commonsourceibias.n364 commonsourceibias.n285 42.5146
R7405 commonsourceibias.n274 commonsourceibias.n195 42.5146
R7406 commonsourceibias.n221 commonsourceibias.n220 42.5146
R7407 commonsourceibias.n458 commonsourceibias.n457 42.5146
R7408 commonsourceibias.n513 commonsourceibias.n434 42.5146
R7409 commonsourceibias.n559 commonsourceibias.n375 42.5146
R7410 commonsourceibias.n399 commonsourceibias.n398 42.5146
R7411 commonsourceibias.n683 commonsourceibias.n682 42.5146
R7412 commonsourceibias.n738 commonsourceibias.n659 42.5146
R7413 commonsourceibias.n593 commonsourceibias.n592 42.5146
R7414 commonsourceibias.n648 commonsourceibias.n569 42.5146
R7415 commonsourceibias.n78 commonsourceibias.n18 41.5458
R7416 commonsourceibias.n53 commonsourceibias.n52 41.5458
R7417 commonsourceibias.n171 commonsourceibias.n6 41.5458
R7418 commonsourceibias.n146 commonsourceibias.n145 41.5458
R7419 commonsourceibias.n325 commonsourceibias.n324 41.5458
R7420 commonsourceibias.n350 commonsourceibias.n290 41.5458
R7421 commonsourceibias.n260 commonsourceibias.n200 41.5458
R7422 commonsourceibias.n235 commonsourceibias.n234 41.5458
R7423 commonsourceibias.n472 commonsourceibias.n471 41.5458
R7424 commonsourceibias.n498 commonsourceibias.n438 41.5458
R7425 commonsourceibias.n544 commonsourceibias.n379 41.5458
R7426 commonsourceibias.n413 commonsourceibias.n412 41.5458
R7427 commonsourceibias.n697 commonsourceibias.n696 41.5458
R7428 commonsourceibias.n723 commonsourceibias.n663 41.5458
R7429 commonsourceibias.n607 commonsourceibias.n606 41.5458
R7430 commonsourceibias.n633 commonsourceibias.n573 41.5458
R7431 commonsourceibias.n68 commonsourceibias.n23 40.577
R7432 commonsourceibias.n64 commonsourceibias.n23 40.577
R7433 commonsourceibias.n161 commonsourceibias.n11 40.577
R7434 commonsourceibias.n157 commonsourceibias.n11 40.577
R7435 commonsourceibias.n336 commonsourceibias.n295 40.577
R7436 commonsourceibias.n340 commonsourceibias.n295 40.577
R7437 commonsourceibias.n250 commonsourceibias.n205 40.577
R7438 commonsourceibias.n246 commonsourceibias.n205 40.577
R7439 commonsourceibias.n483 commonsourceibias.n442 40.577
R7440 commonsourceibias.n487 commonsourceibias.n442 40.577
R7441 commonsourceibias.n533 commonsourceibias.n383 40.577
R7442 commonsourceibias.n424 commonsourceibias.n383 40.577
R7443 commonsourceibias.n708 commonsourceibias.n667 40.577
R7444 commonsourceibias.n712 commonsourceibias.n667 40.577
R7445 commonsourceibias.n618 commonsourceibias.n577 40.577
R7446 commonsourceibias.n622 commonsourceibias.n577 40.577
R7447 commonsourceibias.n82 commonsourceibias.n18 39.6083
R7448 commonsourceibias.n52 commonsourceibias.n51 39.6083
R7449 commonsourceibias.n175 commonsourceibias.n6 39.6083
R7450 commonsourceibias.n145 commonsourceibias.n144 39.6083
R7451 commonsourceibias.n324 commonsourceibias.n323 39.6083
R7452 commonsourceibias.n354 commonsourceibias.n290 39.6083
R7453 commonsourceibias.n264 commonsourceibias.n200 39.6083
R7454 commonsourceibias.n234 commonsourceibias.n233 39.6083
R7455 commonsourceibias.n471 commonsourceibias.n470 39.6083
R7456 commonsourceibias.n502 commonsourceibias.n438 39.6083
R7457 commonsourceibias.n548 commonsourceibias.n379 39.6083
R7458 commonsourceibias.n412 commonsourceibias.n411 39.6083
R7459 commonsourceibias.n696 commonsourceibias.n695 39.6083
R7460 commonsourceibias.n727 commonsourceibias.n663 39.6083
R7461 commonsourceibias.n606 commonsourceibias.n605 39.6083
R7462 commonsourceibias.n637 commonsourceibias.n573 39.6083
R7463 commonsourceibias.n96 commonsourceibias.n13 38.6395
R7464 commonsourceibias.n38 commonsourceibias.n33 38.6395
R7465 commonsourceibias.n189 commonsourceibias.n1 38.6395
R7466 commonsourceibias.n131 commonsourceibias.n126 38.6395
R7467 commonsourceibias.n310 commonsourceibias.n305 38.6395
R7468 commonsourceibias.n368 commonsourceibias.n285 38.6395
R7469 commonsourceibias.n278 commonsourceibias.n195 38.6395
R7470 commonsourceibias.n220 commonsourceibias.n215 38.6395
R7471 commonsourceibias.n457 commonsourceibias.n452 38.6395
R7472 commonsourceibias.n517 commonsourceibias.n434 38.6395
R7473 commonsourceibias.n563 commonsourceibias.n375 38.6395
R7474 commonsourceibias.n398 commonsourceibias.n393 38.6395
R7475 commonsourceibias.n682 commonsourceibias.n677 38.6395
R7476 commonsourceibias.n742 commonsourceibias.n659 38.6395
R7477 commonsourceibias.n592 commonsourceibias.n587 38.6395
R7478 commonsourceibias.n652 commonsourceibias.n569 38.6395
R7479 commonsourceibias.n89 commonsourceibias.n15 26.0455
R7480 commonsourceibias.n45 commonsourceibias.n31 26.0455
R7481 commonsourceibias.n182 commonsourceibias.n3 26.0455
R7482 commonsourceibias.n138 commonsourceibias.n124 26.0455
R7483 commonsourceibias.n317 commonsourceibias.n303 26.0455
R7484 commonsourceibias.n361 commonsourceibias.n287 26.0455
R7485 commonsourceibias.n271 commonsourceibias.n197 26.0455
R7486 commonsourceibias.n227 commonsourceibias.n213 26.0455
R7487 commonsourceibias.n464 commonsourceibias.n450 26.0455
R7488 commonsourceibias.n510 commonsourceibias.n436 26.0455
R7489 commonsourceibias.n556 commonsourceibias.n377 26.0455
R7490 commonsourceibias.n405 commonsourceibias.n391 26.0455
R7491 commonsourceibias.n689 commonsourceibias.n675 26.0455
R7492 commonsourceibias.n735 commonsourceibias.n661 26.0455
R7493 commonsourceibias.n599 commonsourceibias.n585 26.0455
R7494 commonsourceibias.n645 commonsourceibias.n571 26.0455
R7495 commonsourceibias.n75 commonsourceibias.n20 25.0767
R7496 commonsourceibias.n58 commonsourceibias.n57 25.0767
R7497 commonsourceibias.n168 commonsourceibias.n8 25.0767
R7498 commonsourceibias.n151 commonsourceibias.n150 25.0767
R7499 commonsourceibias.n330 commonsourceibias.n329 25.0767
R7500 commonsourceibias.n347 commonsourceibias.n292 25.0767
R7501 commonsourceibias.n257 commonsourceibias.n202 25.0767
R7502 commonsourceibias.n240 commonsourceibias.n239 25.0767
R7503 commonsourceibias.n477 commonsourceibias.n476 25.0767
R7504 commonsourceibias.n495 commonsourceibias.n440 25.0767
R7505 commonsourceibias.n541 commonsourceibias.n381 25.0767
R7506 commonsourceibias.n418 commonsourceibias.n417 25.0767
R7507 commonsourceibias.n702 commonsourceibias.n701 25.0767
R7508 commonsourceibias.n720 commonsourceibias.n665 25.0767
R7509 commonsourceibias.n612 commonsourceibias.n611 25.0767
R7510 commonsourceibias.n630 commonsourceibias.n575 25.0767
R7511 commonsourceibias.n71 commonsourceibias.n22 24.3464
R7512 commonsourceibias.n61 commonsourceibias.n25 24.3464
R7513 commonsourceibias.n164 commonsourceibias.n10 24.3464
R7514 commonsourceibias.n154 commonsourceibias.n118 24.3464
R7515 commonsourceibias.n333 commonsourceibias.n297 24.3464
R7516 commonsourceibias.n343 commonsourceibias.n294 24.3464
R7517 commonsourceibias.n253 commonsourceibias.n204 24.3464
R7518 commonsourceibias.n243 commonsourceibias.n207 24.3464
R7519 commonsourceibias.n480 commonsourceibias.n444 24.3464
R7520 commonsourceibias.n491 commonsourceibias.n490 24.3464
R7521 commonsourceibias.n537 commonsourceibias.n536 24.3464
R7522 commonsourceibias.n421 commonsourceibias.n385 24.3464
R7523 commonsourceibias.n705 commonsourceibias.n669 24.3464
R7524 commonsourceibias.n716 commonsourceibias.n715 24.3464
R7525 commonsourceibias.n615 commonsourceibias.n579 24.3464
R7526 commonsourceibias.n626 commonsourceibias.n625 24.3464
R7527 commonsourceibias.n85 commonsourceibias.n17 23.8546
R7528 commonsourceibias.n47 commonsourceibias.n46 23.8546
R7529 commonsourceibias.n178 commonsourceibias.n5 23.8546
R7530 commonsourceibias.n140 commonsourceibias.n139 23.8546
R7531 commonsourceibias.n319 commonsourceibias.n318 23.8546
R7532 commonsourceibias.n357 commonsourceibias.n289 23.8546
R7533 commonsourceibias.n267 commonsourceibias.n199 23.8546
R7534 commonsourceibias.n229 commonsourceibias.n228 23.8546
R7535 commonsourceibias.n466 commonsourceibias.n465 23.8546
R7536 commonsourceibias.n506 commonsourceibias.n505 23.8546
R7537 commonsourceibias.n552 commonsourceibias.n551 23.8546
R7538 commonsourceibias.n407 commonsourceibias.n406 23.8546
R7539 commonsourceibias.n691 commonsourceibias.n690 23.8546
R7540 commonsourceibias.n731 commonsourceibias.n730 23.8546
R7541 commonsourceibias.n601 commonsourceibias.n600 23.8546
R7542 commonsourceibias.n641 commonsourceibias.n640 23.8546
R7543 commonsourceibias.n98 commonsourceibias.n97 17.4607
R7544 commonsourceibias.n191 commonsourceibias.n190 17.4607
R7545 commonsourceibias.n370 commonsourceibias.n369 17.4607
R7546 commonsourceibias.n280 commonsourceibias.n279 17.4607
R7547 commonsourceibias.n519 commonsourceibias.n518 17.4607
R7548 commonsourceibias.n565 commonsourceibias.n564 17.4607
R7549 commonsourceibias.n744 commonsourceibias.n743 17.4607
R7550 commonsourceibias.n654 commonsourceibias.n653 17.4607
R7551 commonsourceibias.n84 commonsourceibias.n83 16.9689
R7552 commonsourceibias.n48 commonsourceibias.n29 16.9689
R7553 commonsourceibias.n177 commonsourceibias.n176 16.9689
R7554 commonsourceibias.n141 commonsourceibias.n122 16.9689
R7555 commonsourceibias.n320 commonsourceibias.n301 16.9689
R7556 commonsourceibias.n356 commonsourceibias.n355 16.9689
R7557 commonsourceibias.n266 commonsourceibias.n265 16.9689
R7558 commonsourceibias.n230 commonsourceibias.n211 16.9689
R7559 commonsourceibias.n467 commonsourceibias.n448 16.9689
R7560 commonsourceibias.n504 commonsourceibias.n503 16.9689
R7561 commonsourceibias.n550 commonsourceibias.n549 16.9689
R7562 commonsourceibias.n408 commonsourceibias.n389 16.9689
R7563 commonsourceibias.n692 commonsourceibias.n673 16.9689
R7564 commonsourceibias.n729 commonsourceibias.n728 16.9689
R7565 commonsourceibias.n602 commonsourceibias.n583 16.9689
R7566 commonsourceibias.n639 commonsourceibias.n638 16.9689
R7567 commonsourceibias.n70 commonsourceibias.n69 16.477
R7568 commonsourceibias.n63 commonsourceibias.n62 16.477
R7569 commonsourceibias.n163 commonsourceibias.n162 16.477
R7570 commonsourceibias.n156 commonsourceibias.n155 16.477
R7571 commonsourceibias.n335 commonsourceibias.n334 16.477
R7572 commonsourceibias.n342 commonsourceibias.n341 16.477
R7573 commonsourceibias.n252 commonsourceibias.n251 16.477
R7574 commonsourceibias.n245 commonsourceibias.n244 16.477
R7575 commonsourceibias.n482 commonsourceibias.n481 16.477
R7576 commonsourceibias.n489 commonsourceibias.n488 16.477
R7577 commonsourceibias.n535 commonsourceibias.n534 16.477
R7578 commonsourceibias.n423 commonsourceibias.n422 16.477
R7579 commonsourceibias.n707 commonsourceibias.n706 16.477
R7580 commonsourceibias.n714 commonsourceibias.n713 16.477
R7581 commonsourceibias.n617 commonsourceibias.n616 16.477
R7582 commonsourceibias.n624 commonsourceibias.n623 16.477
R7583 commonsourceibias.n77 commonsourceibias.n76 15.9852
R7584 commonsourceibias.n56 commonsourceibias.n27 15.9852
R7585 commonsourceibias.n170 commonsourceibias.n169 15.9852
R7586 commonsourceibias.n149 commonsourceibias.n120 15.9852
R7587 commonsourceibias.n328 commonsourceibias.n299 15.9852
R7588 commonsourceibias.n349 commonsourceibias.n348 15.9852
R7589 commonsourceibias.n259 commonsourceibias.n258 15.9852
R7590 commonsourceibias.n238 commonsourceibias.n209 15.9852
R7591 commonsourceibias.n475 commonsourceibias.n446 15.9852
R7592 commonsourceibias.n497 commonsourceibias.n496 15.9852
R7593 commonsourceibias.n543 commonsourceibias.n542 15.9852
R7594 commonsourceibias.n416 commonsourceibias.n387 15.9852
R7595 commonsourceibias.n700 commonsourceibias.n671 15.9852
R7596 commonsourceibias.n722 commonsourceibias.n721 15.9852
R7597 commonsourceibias.n610 commonsourceibias.n581 15.9852
R7598 commonsourceibias.n632 commonsourceibias.n631 15.9852
R7599 commonsourceibias.n91 commonsourceibias.n90 15.4934
R7600 commonsourceibias.n41 commonsourceibias.n40 15.4934
R7601 commonsourceibias.n184 commonsourceibias.n183 15.4934
R7602 commonsourceibias.n134 commonsourceibias.n133 15.4934
R7603 commonsourceibias.n313 commonsourceibias.n312 15.4934
R7604 commonsourceibias.n363 commonsourceibias.n362 15.4934
R7605 commonsourceibias.n273 commonsourceibias.n272 15.4934
R7606 commonsourceibias.n223 commonsourceibias.n222 15.4934
R7607 commonsourceibias.n460 commonsourceibias.n459 15.4934
R7608 commonsourceibias.n512 commonsourceibias.n511 15.4934
R7609 commonsourceibias.n558 commonsourceibias.n557 15.4934
R7610 commonsourceibias.n401 commonsourceibias.n400 15.4934
R7611 commonsourceibias.n685 commonsourceibias.n684 15.4934
R7612 commonsourceibias.n737 commonsourceibias.n736 15.4934
R7613 commonsourceibias.n595 commonsourceibias.n594 15.4934
R7614 commonsourceibias.n647 commonsourceibias.n646 15.4934
R7615 commonsourceibias.n102 commonsourceibias.n100 13.2663
R7616 commonsourceibias.n523 commonsourceibias.n521 13.2663
R7617 commonsourceibias.n748 commonsourceibias.n373 10.122
R7618 commonsourceibias.n159 commonsourceibias.n116 9.50363
R7619 commonsourceibias.n531 commonsourceibias.n530 9.50363
R7620 commonsourceibias.n92 commonsourceibias.n91 9.09948
R7621 commonsourceibias.n40 commonsourceibias.n39 9.09948
R7622 commonsourceibias.n185 commonsourceibias.n184 9.09948
R7623 commonsourceibias.n133 commonsourceibias.n132 9.09948
R7624 commonsourceibias.n312 commonsourceibias.n311 9.09948
R7625 commonsourceibias.n364 commonsourceibias.n363 9.09948
R7626 commonsourceibias.n274 commonsourceibias.n273 9.09948
R7627 commonsourceibias.n222 commonsourceibias.n221 9.09948
R7628 commonsourceibias.n459 commonsourceibias.n458 9.09948
R7629 commonsourceibias.n513 commonsourceibias.n512 9.09948
R7630 commonsourceibias.n559 commonsourceibias.n558 9.09948
R7631 commonsourceibias.n400 commonsourceibias.n399 9.09948
R7632 commonsourceibias.n684 commonsourceibias.n683 9.09948
R7633 commonsourceibias.n738 commonsourceibias.n737 9.09948
R7634 commonsourceibias.n594 commonsourceibias.n593 9.09948
R7635 commonsourceibias.n648 commonsourceibias.n647 9.09948
R7636 commonsourceibias.n283 commonsourceibias.n193 8.79451
R7637 commonsourceibias.n657 commonsourceibias.n567 8.79451
R7638 commonsourceibias.n78 commonsourceibias.n77 8.60764
R7639 commonsourceibias.n53 commonsourceibias.n27 8.60764
R7640 commonsourceibias.n171 commonsourceibias.n170 8.60764
R7641 commonsourceibias.n146 commonsourceibias.n120 8.60764
R7642 commonsourceibias.n325 commonsourceibias.n299 8.60764
R7643 commonsourceibias.n350 commonsourceibias.n349 8.60764
R7644 commonsourceibias.n260 commonsourceibias.n259 8.60764
R7645 commonsourceibias.n235 commonsourceibias.n209 8.60764
R7646 commonsourceibias.n472 commonsourceibias.n446 8.60764
R7647 commonsourceibias.n498 commonsourceibias.n497 8.60764
R7648 commonsourceibias.n544 commonsourceibias.n543 8.60764
R7649 commonsourceibias.n413 commonsourceibias.n387 8.60764
R7650 commonsourceibias.n697 commonsourceibias.n671 8.60764
R7651 commonsourceibias.n723 commonsourceibias.n722 8.60764
R7652 commonsourceibias.n607 commonsourceibias.n581 8.60764
R7653 commonsourceibias.n633 commonsourceibias.n632 8.60764
R7654 commonsourceibias.n748 commonsourceibias.n747 8.46921
R7655 commonsourceibias.n69 commonsourceibias.n68 8.11581
R7656 commonsourceibias.n64 commonsourceibias.n63 8.11581
R7657 commonsourceibias.n162 commonsourceibias.n161 8.11581
R7658 commonsourceibias.n157 commonsourceibias.n156 8.11581
R7659 commonsourceibias.n336 commonsourceibias.n335 8.11581
R7660 commonsourceibias.n341 commonsourceibias.n340 8.11581
R7661 commonsourceibias.n251 commonsourceibias.n250 8.11581
R7662 commonsourceibias.n246 commonsourceibias.n245 8.11581
R7663 commonsourceibias.n483 commonsourceibias.n482 8.11581
R7664 commonsourceibias.n488 commonsourceibias.n487 8.11581
R7665 commonsourceibias.n534 commonsourceibias.n533 8.11581
R7666 commonsourceibias.n424 commonsourceibias.n423 8.11581
R7667 commonsourceibias.n708 commonsourceibias.n707 8.11581
R7668 commonsourceibias.n713 commonsourceibias.n712 8.11581
R7669 commonsourceibias.n618 commonsourceibias.n617 8.11581
R7670 commonsourceibias.n623 commonsourceibias.n622 8.11581
R7671 commonsourceibias.n83 commonsourceibias.n82 7.62397
R7672 commonsourceibias.n51 commonsourceibias.n29 7.62397
R7673 commonsourceibias.n176 commonsourceibias.n175 7.62397
R7674 commonsourceibias.n144 commonsourceibias.n122 7.62397
R7675 commonsourceibias.n323 commonsourceibias.n301 7.62397
R7676 commonsourceibias.n355 commonsourceibias.n354 7.62397
R7677 commonsourceibias.n265 commonsourceibias.n264 7.62397
R7678 commonsourceibias.n233 commonsourceibias.n211 7.62397
R7679 commonsourceibias.n470 commonsourceibias.n448 7.62397
R7680 commonsourceibias.n503 commonsourceibias.n502 7.62397
R7681 commonsourceibias.n549 commonsourceibias.n548 7.62397
R7682 commonsourceibias.n411 commonsourceibias.n389 7.62397
R7683 commonsourceibias.n695 commonsourceibias.n673 7.62397
R7684 commonsourceibias.n728 commonsourceibias.n727 7.62397
R7685 commonsourceibias.n605 commonsourceibias.n583 7.62397
R7686 commonsourceibias.n638 commonsourceibias.n637 7.62397
R7687 commonsourceibias.n97 commonsourceibias.n96 7.13213
R7688 commonsourceibias.n34 commonsourceibias.n33 7.13213
R7689 commonsourceibias.n190 commonsourceibias.n189 7.13213
R7690 commonsourceibias.n127 commonsourceibias.n126 7.13213
R7691 commonsourceibias.n306 commonsourceibias.n305 7.13213
R7692 commonsourceibias.n369 commonsourceibias.n368 7.13213
R7693 commonsourceibias.n279 commonsourceibias.n278 7.13213
R7694 commonsourceibias.n216 commonsourceibias.n215 7.13213
R7695 commonsourceibias.n453 commonsourceibias.n452 7.13213
R7696 commonsourceibias.n518 commonsourceibias.n517 7.13213
R7697 commonsourceibias.n564 commonsourceibias.n563 7.13213
R7698 commonsourceibias.n394 commonsourceibias.n393 7.13213
R7699 commonsourceibias.n678 commonsourceibias.n677 7.13213
R7700 commonsourceibias.n743 commonsourceibias.n742 7.13213
R7701 commonsourceibias.n588 commonsourceibias.n587 7.13213
R7702 commonsourceibias.n653 commonsourceibias.n652 7.13213
R7703 commonsourceibias.n373 commonsourceibias.n372 5.06534
R7704 commonsourceibias.n283 commonsourceibias.n282 5.06534
R7705 commonsourceibias.n747 commonsourceibias.n746 5.06534
R7706 commonsourceibias.n657 commonsourceibias.n656 5.06534
R7707 commonsourceibias commonsourceibias.n748 4.08303
R7708 commonsourceibias.n373 commonsourceibias.n283 3.72967
R7709 commonsourceibias.n747 commonsourceibias.n657 3.72967
R7710 commonsourceibias.n109 commonsourceibias.t17 2.82907
R7711 commonsourceibias.n109 commonsourceibias.t57 2.82907
R7712 commonsourceibias.n110 commonsourceibias.t63 2.82907
R7713 commonsourceibias.n110 commonsourceibias.t43 2.82907
R7714 commonsourceibias.n112 commonsourceibias.t9 2.82907
R7715 commonsourceibias.n112 commonsourceibias.t47 2.82907
R7716 commonsourceibias.n114 commonsourceibias.t23 2.82907
R7717 commonsourceibias.n114 commonsourceibias.t39 2.82907
R7718 commonsourceibias.n107 commonsourceibias.t13 2.82907
R7719 commonsourceibias.n107 commonsourceibias.t55 2.82907
R7720 commonsourceibias.n105 commonsourceibias.t61 2.82907
R7721 commonsourceibias.n105 commonsourceibias.t25 2.82907
R7722 commonsourceibias.n103 commonsourceibias.t59 2.82907
R7723 commonsourceibias.n103 commonsourceibias.t19 2.82907
R7724 commonsourceibias.n101 commonsourceibias.t21 2.82907
R7725 commonsourceibias.n101 commonsourceibias.t15 2.82907
R7726 commonsourceibias.n522 commonsourceibias.t49 2.82907
R7727 commonsourceibias.n522 commonsourceibias.t29 2.82907
R7728 commonsourceibias.n524 commonsourceibias.t27 2.82907
R7729 commonsourceibias.n524 commonsourceibias.t45 2.82907
R7730 commonsourceibias.n526 commonsourceibias.t33 2.82907
R7731 commonsourceibias.n526 commonsourceibias.t5 2.82907
R7732 commonsourceibias.n528 commonsourceibias.t11 2.82907
R7733 commonsourceibias.n528 commonsourceibias.t41 2.82907
R7734 commonsourceibias.n431 commonsourceibias.t3 2.82907
R7735 commonsourceibias.n431 commonsourceibias.t31 2.82907
R7736 commonsourceibias.n429 commonsourceibias.t1 2.82907
R7737 commonsourceibias.n429 commonsourceibias.t35 2.82907
R7738 commonsourceibias.n427 commonsourceibias.t37 2.82907
R7739 commonsourceibias.n427 commonsourceibias.t53 2.82907
R7740 commonsourceibias.n426 commonsourceibias.t7 2.82907
R7741 commonsourceibias.n426 commonsourceibias.t51 2.82907
R7742 commonsourceibias.n17 commonsourceibias.n15 0.738255
R7743 commonsourceibias.n46 commonsourceibias.n45 0.738255
R7744 commonsourceibias.n5 commonsourceibias.n3 0.738255
R7745 commonsourceibias.n139 commonsourceibias.n138 0.738255
R7746 commonsourceibias.n318 commonsourceibias.n317 0.738255
R7747 commonsourceibias.n289 commonsourceibias.n287 0.738255
R7748 commonsourceibias.n199 commonsourceibias.n197 0.738255
R7749 commonsourceibias.n228 commonsourceibias.n227 0.738255
R7750 commonsourceibias.n465 commonsourceibias.n464 0.738255
R7751 commonsourceibias.n505 commonsourceibias.n436 0.738255
R7752 commonsourceibias.n551 commonsourceibias.n377 0.738255
R7753 commonsourceibias.n406 commonsourceibias.n405 0.738255
R7754 commonsourceibias.n690 commonsourceibias.n689 0.738255
R7755 commonsourceibias.n730 commonsourceibias.n661 0.738255
R7756 commonsourceibias.n600 commonsourceibias.n599 0.738255
R7757 commonsourceibias.n640 commonsourceibias.n571 0.738255
R7758 commonsourceibias.n104 commonsourceibias.n102 0.573776
R7759 commonsourceibias.n106 commonsourceibias.n104 0.573776
R7760 commonsourceibias.n108 commonsourceibias.n106 0.573776
R7761 commonsourceibias.n115 commonsourceibias.n113 0.573776
R7762 commonsourceibias.n113 commonsourceibias.n111 0.573776
R7763 commonsourceibias.n430 commonsourceibias.n428 0.573776
R7764 commonsourceibias.n432 commonsourceibias.n430 0.573776
R7765 commonsourceibias.n529 commonsourceibias.n527 0.573776
R7766 commonsourceibias.n527 commonsourceibias.n525 0.573776
R7767 commonsourceibias.n525 commonsourceibias.n523 0.573776
R7768 commonsourceibias.n116 commonsourceibias.n108 0.287138
R7769 commonsourceibias.n116 commonsourceibias.n115 0.287138
R7770 commonsourceibias.n530 commonsourceibias.n432 0.287138
R7771 commonsourceibias.n530 commonsourceibias.n529 0.287138
R7772 commonsourceibias.n100 commonsourceibias.n12 0.285035
R7773 commonsourceibias.n193 commonsourceibias.n0 0.285035
R7774 commonsourceibias.n372 commonsourceibias.n284 0.285035
R7775 commonsourceibias.n282 commonsourceibias.n194 0.285035
R7776 commonsourceibias.n521 commonsourceibias.n433 0.285035
R7777 commonsourceibias.n567 commonsourceibias.n374 0.285035
R7778 commonsourceibias.n746 commonsourceibias.n658 0.285035
R7779 commonsourceibias.n656 commonsourceibias.n568 0.285035
R7780 commonsourceibias.n22 commonsourceibias.n20 0.246418
R7781 commonsourceibias.n58 commonsourceibias.n25 0.246418
R7782 commonsourceibias.n10 commonsourceibias.n8 0.246418
R7783 commonsourceibias.n151 commonsourceibias.n118 0.246418
R7784 commonsourceibias.n330 commonsourceibias.n297 0.246418
R7785 commonsourceibias.n294 commonsourceibias.n292 0.246418
R7786 commonsourceibias.n204 commonsourceibias.n202 0.246418
R7787 commonsourceibias.n240 commonsourceibias.n207 0.246418
R7788 commonsourceibias.n477 commonsourceibias.n444 0.246418
R7789 commonsourceibias.n490 commonsourceibias.n440 0.246418
R7790 commonsourceibias.n536 commonsourceibias.n381 0.246418
R7791 commonsourceibias.n418 commonsourceibias.n385 0.246418
R7792 commonsourceibias.n702 commonsourceibias.n669 0.246418
R7793 commonsourceibias.n715 commonsourceibias.n665 0.246418
R7794 commonsourceibias.n612 commonsourceibias.n579 0.246418
R7795 commonsourceibias.n625 commonsourceibias.n575 0.246418
R7796 commonsourceibias.n95 commonsourceibias.n12 0.189894
R7797 commonsourceibias.n95 commonsourceibias.n94 0.189894
R7798 commonsourceibias.n94 commonsourceibias.n93 0.189894
R7799 commonsourceibias.n93 commonsourceibias.n14 0.189894
R7800 commonsourceibias.n88 commonsourceibias.n14 0.189894
R7801 commonsourceibias.n88 commonsourceibias.n87 0.189894
R7802 commonsourceibias.n87 commonsourceibias.n86 0.189894
R7803 commonsourceibias.n86 commonsourceibias.n16 0.189894
R7804 commonsourceibias.n81 commonsourceibias.n16 0.189894
R7805 commonsourceibias.n81 commonsourceibias.n80 0.189894
R7806 commonsourceibias.n80 commonsourceibias.n79 0.189894
R7807 commonsourceibias.n79 commonsourceibias.n19 0.189894
R7808 commonsourceibias.n74 commonsourceibias.n19 0.189894
R7809 commonsourceibias.n74 commonsourceibias.n73 0.189894
R7810 commonsourceibias.n73 commonsourceibias.n72 0.189894
R7811 commonsourceibias.n72 commonsourceibias.n21 0.189894
R7812 commonsourceibias.n67 commonsourceibias.n21 0.189894
R7813 commonsourceibias.n67 commonsourceibias.n66 0.189894
R7814 commonsourceibias.n66 commonsourceibias.n65 0.189894
R7815 commonsourceibias.n65 commonsourceibias.n24 0.189894
R7816 commonsourceibias.n60 commonsourceibias.n24 0.189894
R7817 commonsourceibias.n60 commonsourceibias.n59 0.189894
R7818 commonsourceibias.n59 commonsourceibias.n26 0.189894
R7819 commonsourceibias.n55 commonsourceibias.n26 0.189894
R7820 commonsourceibias.n55 commonsourceibias.n54 0.189894
R7821 commonsourceibias.n54 commonsourceibias.n28 0.189894
R7822 commonsourceibias.n50 commonsourceibias.n28 0.189894
R7823 commonsourceibias.n50 commonsourceibias.n49 0.189894
R7824 commonsourceibias.n49 commonsourceibias.n30 0.189894
R7825 commonsourceibias.n44 commonsourceibias.n30 0.189894
R7826 commonsourceibias.n44 commonsourceibias.n43 0.189894
R7827 commonsourceibias.n43 commonsourceibias.n42 0.189894
R7828 commonsourceibias.n42 commonsourceibias.n32 0.189894
R7829 commonsourceibias.n37 commonsourceibias.n32 0.189894
R7830 commonsourceibias.n37 commonsourceibias.n36 0.189894
R7831 commonsourceibias.n158 commonsourceibias.n117 0.189894
R7832 commonsourceibias.n153 commonsourceibias.n117 0.189894
R7833 commonsourceibias.n153 commonsourceibias.n152 0.189894
R7834 commonsourceibias.n152 commonsourceibias.n119 0.189894
R7835 commonsourceibias.n148 commonsourceibias.n119 0.189894
R7836 commonsourceibias.n148 commonsourceibias.n147 0.189894
R7837 commonsourceibias.n147 commonsourceibias.n121 0.189894
R7838 commonsourceibias.n143 commonsourceibias.n121 0.189894
R7839 commonsourceibias.n143 commonsourceibias.n142 0.189894
R7840 commonsourceibias.n142 commonsourceibias.n123 0.189894
R7841 commonsourceibias.n137 commonsourceibias.n123 0.189894
R7842 commonsourceibias.n137 commonsourceibias.n136 0.189894
R7843 commonsourceibias.n136 commonsourceibias.n135 0.189894
R7844 commonsourceibias.n135 commonsourceibias.n125 0.189894
R7845 commonsourceibias.n130 commonsourceibias.n125 0.189894
R7846 commonsourceibias.n130 commonsourceibias.n129 0.189894
R7847 commonsourceibias.n188 commonsourceibias.n0 0.189894
R7848 commonsourceibias.n188 commonsourceibias.n187 0.189894
R7849 commonsourceibias.n187 commonsourceibias.n186 0.189894
R7850 commonsourceibias.n186 commonsourceibias.n2 0.189894
R7851 commonsourceibias.n181 commonsourceibias.n2 0.189894
R7852 commonsourceibias.n181 commonsourceibias.n180 0.189894
R7853 commonsourceibias.n180 commonsourceibias.n179 0.189894
R7854 commonsourceibias.n179 commonsourceibias.n4 0.189894
R7855 commonsourceibias.n174 commonsourceibias.n4 0.189894
R7856 commonsourceibias.n174 commonsourceibias.n173 0.189894
R7857 commonsourceibias.n173 commonsourceibias.n172 0.189894
R7858 commonsourceibias.n172 commonsourceibias.n7 0.189894
R7859 commonsourceibias.n167 commonsourceibias.n7 0.189894
R7860 commonsourceibias.n167 commonsourceibias.n166 0.189894
R7861 commonsourceibias.n166 commonsourceibias.n165 0.189894
R7862 commonsourceibias.n165 commonsourceibias.n9 0.189894
R7863 commonsourceibias.n160 commonsourceibias.n9 0.189894
R7864 commonsourceibias.n367 commonsourceibias.n284 0.189894
R7865 commonsourceibias.n367 commonsourceibias.n366 0.189894
R7866 commonsourceibias.n366 commonsourceibias.n365 0.189894
R7867 commonsourceibias.n365 commonsourceibias.n286 0.189894
R7868 commonsourceibias.n360 commonsourceibias.n286 0.189894
R7869 commonsourceibias.n360 commonsourceibias.n359 0.189894
R7870 commonsourceibias.n359 commonsourceibias.n358 0.189894
R7871 commonsourceibias.n358 commonsourceibias.n288 0.189894
R7872 commonsourceibias.n353 commonsourceibias.n288 0.189894
R7873 commonsourceibias.n353 commonsourceibias.n352 0.189894
R7874 commonsourceibias.n352 commonsourceibias.n351 0.189894
R7875 commonsourceibias.n351 commonsourceibias.n291 0.189894
R7876 commonsourceibias.n346 commonsourceibias.n291 0.189894
R7877 commonsourceibias.n346 commonsourceibias.n345 0.189894
R7878 commonsourceibias.n345 commonsourceibias.n344 0.189894
R7879 commonsourceibias.n344 commonsourceibias.n293 0.189894
R7880 commonsourceibias.n339 commonsourceibias.n293 0.189894
R7881 commonsourceibias.n339 commonsourceibias.n338 0.189894
R7882 commonsourceibias.n338 commonsourceibias.n337 0.189894
R7883 commonsourceibias.n337 commonsourceibias.n296 0.189894
R7884 commonsourceibias.n332 commonsourceibias.n296 0.189894
R7885 commonsourceibias.n332 commonsourceibias.n331 0.189894
R7886 commonsourceibias.n331 commonsourceibias.n298 0.189894
R7887 commonsourceibias.n327 commonsourceibias.n298 0.189894
R7888 commonsourceibias.n327 commonsourceibias.n326 0.189894
R7889 commonsourceibias.n326 commonsourceibias.n300 0.189894
R7890 commonsourceibias.n322 commonsourceibias.n300 0.189894
R7891 commonsourceibias.n322 commonsourceibias.n321 0.189894
R7892 commonsourceibias.n321 commonsourceibias.n302 0.189894
R7893 commonsourceibias.n316 commonsourceibias.n302 0.189894
R7894 commonsourceibias.n316 commonsourceibias.n315 0.189894
R7895 commonsourceibias.n315 commonsourceibias.n314 0.189894
R7896 commonsourceibias.n314 commonsourceibias.n304 0.189894
R7897 commonsourceibias.n309 commonsourceibias.n304 0.189894
R7898 commonsourceibias.n309 commonsourceibias.n308 0.189894
R7899 commonsourceibias.n277 commonsourceibias.n194 0.189894
R7900 commonsourceibias.n277 commonsourceibias.n276 0.189894
R7901 commonsourceibias.n276 commonsourceibias.n275 0.189894
R7902 commonsourceibias.n275 commonsourceibias.n196 0.189894
R7903 commonsourceibias.n270 commonsourceibias.n196 0.189894
R7904 commonsourceibias.n270 commonsourceibias.n269 0.189894
R7905 commonsourceibias.n269 commonsourceibias.n268 0.189894
R7906 commonsourceibias.n268 commonsourceibias.n198 0.189894
R7907 commonsourceibias.n263 commonsourceibias.n198 0.189894
R7908 commonsourceibias.n263 commonsourceibias.n262 0.189894
R7909 commonsourceibias.n262 commonsourceibias.n261 0.189894
R7910 commonsourceibias.n261 commonsourceibias.n201 0.189894
R7911 commonsourceibias.n256 commonsourceibias.n201 0.189894
R7912 commonsourceibias.n256 commonsourceibias.n255 0.189894
R7913 commonsourceibias.n255 commonsourceibias.n254 0.189894
R7914 commonsourceibias.n254 commonsourceibias.n203 0.189894
R7915 commonsourceibias.n249 commonsourceibias.n203 0.189894
R7916 commonsourceibias.n249 commonsourceibias.n248 0.189894
R7917 commonsourceibias.n248 commonsourceibias.n247 0.189894
R7918 commonsourceibias.n247 commonsourceibias.n206 0.189894
R7919 commonsourceibias.n242 commonsourceibias.n206 0.189894
R7920 commonsourceibias.n242 commonsourceibias.n241 0.189894
R7921 commonsourceibias.n241 commonsourceibias.n208 0.189894
R7922 commonsourceibias.n237 commonsourceibias.n208 0.189894
R7923 commonsourceibias.n237 commonsourceibias.n236 0.189894
R7924 commonsourceibias.n236 commonsourceibias.n210 0.189894
R7925 commonsourceibias.n232 commonsourceibias.n210 0.189894
R7926 commonsourceibias.n232 commonsourceibias.n231 0.189894
R7927 commonsourceibias.n231 commonsourceibias.n212 0.189894
R7928 commonsourceibias.n226 commonsourceibias.n212 0.189894
R7929 commonsourceibias.n226 commonsourceibias.n225 0.189894
R7930 commonsourceibias.n225 commonsourceibias.n224 0.189894
R7931 commonsourceibias.n224 commonsourceibias.n214 0.189894
R7932 commonsourceibias.n219 commonsourceibias.n214 0.189894
R7933 commonsourceibias.n219 commonsourceibias.n218 0.189894
R7934 commonsourceibias.n456 commonsourceibias.n455 0.189894
R7935 commonsourceibias.n456 commonsourceibias.n451 0.189894
R7936 commonsourceibias.n461 commonsourceibias.n451 0.189894
R7937 commonsourceibias.n462 commonsourceibias.n461 0.189894
R7938 commonsourceibias.n463 commonsourceibias.n462 0.189894
R7939 commonsourceibias.n463 commonsourceibias.n449 0.189894
R7940 commonsourceibias.n468 commonsourceibias.n449 0.189894
R7941 commonsourceibias.n469 commonsourceibias.n468 0.189894
R7942 commonsourceibias.n469 commonsourceibias.n447 0.189894
R7943 commonsourceibias.n473 commonsourceibias.n447 0.189894
R7944 commonsourceibias.n474 commonsourceibias.n473 0.189894
R7945 commonsourceibias.n474 commonsourceibias.n445 0.189894
R7946 commonsourceibias.n478 commonsourceibias.n445 0.189894
R7947 commonsourceibias.n479 commonsourceibias.n478 0.189894
R7948 commonsourceibias.n479 commonsourceibias.n443 0.189894
R7949 commonsourceibias.n484 commonsourceibias.n443 0.189894
R7950 commonsourceibias.n485 commonsourceibias.n484 0.189894
R7951 commonsourceibias.n486 commonsourceibias.n485 0.189894
R7952 commonsourceibias.n486 commonsourceibias.n441 0.189894
R7953 commonsourceibias.n492 commonsourceibias.n441 0.189894
R7954 commonsourceibias.n493 commonsourceibias.n492 0.189894
R7955 commonsourceibias.n494 commonsourceibias.n493 0.189894
R7956 commonsourceibias.n494 commonsourceibias.n439 0.189894
R7957 commonsourceibias.n499 commonsourceibias.n439 0.189894
R7958 commonsourceibias.n500 commonsourceibias.n499 0.189894
R7959 commonsourceibias.n501 commonsourceibias.n500 0.189894
R7960 commonsourceibias.n501 commonsourceibias.n437 0.189894
R7961 commonsourceibias.n507 commonsourceibias.n437 0.189894
R7962 commonsourceibias.n508 commonsourceibias.n507 0.189894
R7963 commonsourceibias.n509 commonsourceibias.n508 0.189894
R7964 commonsourceibias.n509 commonsourceibias.n435 0.189894
R7965 commonsourceibias.n514 commonsourceibias.n435 0.189894
R7966 commonsourceibias.n515 commonsourceibias.n514 0.189894
R7967 commonsourceibias.n516 commonsourceibias.n515 0.189894
R7968 commonsourceibias.n516 commonsourceibias.n433 0.189894
R7969 commonsourceibias.n397 commonsourceibias.n396 0.189894
R7970 commonsourceibias.n397 commonsourceibias.n392 0.189894
R7971 commonsourceibias.n402 commonsourceibias.n392 0.189894
R7972 commonsourceibias.n403 commonsourceibias.n402 0.189894
R7973 commonsourceibias.n404 commonsourceibias.n403 0.189894
R7974 commonsourceibias.n404 commonsourceibias.n390 0.189894
R7975 commonsourceibias.n409 commonsourceibias.n390 0.189894
R7976 commonsourceibias.n410 commonsourceibias.n409 0.189894
R7977 commonsourceibias.n410 commonsourceibias.n388 0.189894
R7978 commonsourceibias.n414 commonsourceibias.n388 0.189894
R7979 commonsourceibias.n415 commonsourceibias.n414 0.189894
R7980 commonsourceibias.n415 commonsourceibias.n386 0.189894
R7981 commonsourceibias.n419 commonsourceibias.n386 0.189894
R7982 commonsourceibias.n420 commonsourceibias.n419 0.189894
R7983 commonsourceibias.n420 commonsourceibias.n384 0.189894
R7984 commonsourceibias.n425 commonsourceibias.n384 0.189894
R7985 commonsourceibias.n532 commonsourceibias.n382 0.189894
R7986 commonsourceibias.n538 commonsourceibias.n382 0.189894
R7987 commonsourceibias.n539 commonsourceibias.n538 0.189894
R7988 commonsourceibias.n540 commonsourceibias.n539 0.189894
R7989 commonsourceibias.n540 commonsourceibias.n380 0.189894
R7990 commonsourceibias.n545 commonsourceibias.n380 0.189894
R7991 commonsourceibias.n546 commonsourceibias.n545 0.189894
R7992 commonsourceibias.n547 commonsourceibias.n546 0.189894
R7993 commonsourceibias.n547 commonsourceibias.n378 0.189894
R7994 commonsourceibias.n553 commonsourceibias.n378 0.189894
R7995 commonsourceibias.n554 commonsourceibias.n553 0.189894
R7996 commonsourceibias.n555 commonsourceibias.n554 0.189894
R7997 commonsourceibias.n555 commonsourceibias.n376 0.189894
R7998 commonsourceibias.n560 commonsourceibias.n376 0.189894
R7999 commonsourceibias.n561 commonsourceibias.n560 0.189894
R8000 commonsourceibias.n562 commonsourceibias.n561 0.189894
R8001 commonsourceibias.n562 commonsourceibias.n374 0.189894
R8002 commonsourceibias.n681 commonsourceibias.n680 0.189894
R8003 commonsourceibias.n681 commonsourceibias.n676 0.189894
R8004 commonsourceibias.n686 commonsourceibias.n676 0.189894
R8005 commonsourceibias.n687 commonsourceibias.n686 0.189894
R8006 commonsourceibias.n688 commonsourceibias.n687 0.189894
R8007 commonsourceibias.n688 commonsourceibias.n674 0.189894
R8008 commonsourceibias.n693 commonsourceibias.n674 0.189894
R8009 commonsourceibias.n694 commonsourceibias.n693 0.189894
R8010 commonsourceibias.n694 commonsourceibias.n672 0.189894
R8011 commonsourceibias.n698 commonsourceibias.n672 0.189894
R8012 commonsourceibias.n699 commonsourceibias.n698 0.189894
R8013 commonsourceibias.n699 commonsourceibias.n670 0.189894
R8014 commonsourceibias.n703 commonsourceibias.n670 0.189894
R8015 commonsourceibias.n704 commonsourceibias.n703 0.189894
R8016 commonsourceibias.n704 commonsourceibias.n668 0.189894
R8017 commonsourceibias.n709 commonsourceibias.n668 0.189894
R8018 commonsourceibias.n710 commonsourceibias.n709 0.189894
R8019 commonsourceibias.n711 commonsourceibias.n710 0.189894
R8020 commonsourceibias.n711 commonsourceibias.n666 0.189894
R8021 commonsourceibias.n717 commonsourceibias.n666 0.189894
R8022 commonsourceibias.n718 commonsourceibias.n717 0.189894
R8023 commonsourceibias.n719 commonsourceibias.n718 0.189894
R8024 commonsourceibias.n719 commonsourceibias.n664 0.189894
R8025 commonsourceibias.n724 commonsourceibias.n664 0.189894
R8026 commonsourceibias.n725 commonsourceibias.n724 0.189894
R8027 commonsourceibias.n726 commonsourceibias.n725 0.189894
R8028 commonsourceibias.n726 commonsourceibias.n662 0.189894
R8029 commonsourceibias.n732 commonsourceibias.n662 0.189894
R8030 commonsourceibias.n733 commonsourceibias.n732 0.189894
R8031 commonsourceibias.n734 commonsourceibias.n733 0.189894
R8032 commonsourceibias.n734 commonsourceibias.n660 0.189894
R8033 commonsourceibias.n739 commonsourceibias.n660 0.189894
R8034 commonsourceibias.n740 commonsourceibias.n739 0.189894
R8035 commonsourceibias.n741 commonsourceibias.n740 0.189894
R8036 commonsourceibias.n741 commonsourceibias.n658 0.189894
R8037 commonsourceibias.n591 commonsourceibias.n590 0.189894
R8038 commonsourceibias.n591 commonsourceibias.n586 0.189894
R8039 commonsourceibias.n596 commonsourceibias.n586 0.189894
R8040 commonsourceibias.n597 commonsourceibias.n596 0.189894
R8041 commonsourceibias.n598 commonsourceibias.n597 0.189894
R8042 commonsourceibias.n598 commonsourceibias.n584 0.189894
R8043 commonsourceibias.n603 commonsourceibias.n584 0.189894
R8044 commonsourceibias.n604 commonsourceibias.n603 0.189894
R8045 commonsourceibias.n604 commonsourceibias.n582 0.189894
R8046 commonsourceibias.n608 commonsourceibias.n582 0.189894
R8047 commonsourceibias.n609 commonsourceibias.n608 0.189894
R8048 commonsourceibias.n609 commonsourceibias.n580 0.189894
R8049 commonsourceibias.n613 commonsourceibias.n580 0.189894
R8050 commonsourceibias.n614 commonsourceibias.n613 0.189894
R8051 commonsourceibias.n614 commonsourceibias.n578 0.189894
R8052 commonsourceibias.n619 commonsourceibias.n578 0.189894
R8053 commonsourceibias.n620 commonsourceibias.n619 0.189894
R8054 commonsourceibias.n621 commonsourceibias.n620 0.189894
R8055 commonsourceibias.n621 commonsourceibias.n576 0.189894
R8056 commonsourceibias.n627 commonsourceibias.n576 0.189894
R8057 commonsourceibias.n628 commonsourceibias.n627 0.189894
R8058 commonsourceibias.n629 commonsourceibias.n628 0.189894
R8059 commonsourceibias.n629 commonsourceibias.n574 0.189894
R8060 commonsourceibias.n634 commonsourceibias.n574 0.189894
R8061 commonsourceibias.n635 commonsourceibias.n634 0.189894
R8062 commonsourceibias.n636 commonsourceibias.n635 0.189894
R8063 commonsourceibias.n636 commonsourceibias.n572 0.189894
R8064 commonsourceibias.n642 commonsourceibias.n572 0.189894
R8065 commonsourceibias.n643 commonsourceibias.n642 0.189894
R8066 commonsourceibias.n644 commonsourceibias.n643 0.189894
R8067 commonsourceibias.n644 commonsourceibias.n570 0.189894
R8068 commonsourceibias.n649 commonsourceibias.n570 0.189894
R8069 commonsourceibias.n650 commonsourceibias.n649 0.189894
R8070 commonsourceibias.n651 commonsourceibias.n650 0.189894
R8071 commonsourceibias.n651 commonsourceibias.n568 0.189894
R8072 commonsourceibias.n159 commonsourceibias.n158 0.170955
R8073 commonsourceibias.n160 commonsourceibias.n159 0.170955
R8074 commonsourceibias.n531 commonsourceibias.n425 0.170955
R8075 commonsourceibias.n532 commonsourceibias.n531 0.170955
R8076 gnd.n7317 gnd.n7316 1810.87
R8077 gnd.n5236 gnd.n5235 927.927
R8078 gnd.n7808 gnd.n211 795.207
R8079 gnd.n352 gnd.n214 795.207
R8080 gnd.n3942 gnd.n1726 795.207
R8081 gnd.n4011 gnd.n1728 795.207
R8082 gnd.n4967 gnd.n1478 795.207
R8083 gnd.n3160 gnd.n1481 795.207
R8084 gnd.n1243 gnd.n1168 795.207
R8085 gnd.n5102 gnd.n1245 795.207
R8086 gnd.n3235 gnd.n2387 771.183
R8087 gnd.n4727 gnd.n1703 771.183
R8088 gnd.n3151 gnd.n2389 771.183
R8089 gnd.n4099 gnd.n1705 771.183
R8090 gnd.n6580 gnd.n1121 766.379
R8091 gnd.n6496 gnd.n1123 766.379
R8092 gnd.n5791 gnd.n5694 766.379
R8093 gnd.n5787 gnd.n5692 766.379
R8094 gnd.n6577 gnd.n5238 756.769
R8095 gnd.n6546 gnd.n1124 756.769
R8096 gnd.n5884 gnd.n5601 756.769
R8097 gnd.n5882 gnd.n5604 756.769
R8098 gnd.n7806 gnd.n216 739.952
R8099 gnd.n7697 gnd.n213 739.952
R8100 gnd.n4486 gnd.n1725 739.952
R8101 gnd.n4709 gnd.n1729 739.952
R8102 gnd.n4965 gnd.n1483 739.952
R8103 gnd.n2529 gnd.n1480 739.952
R8104 gnd.n5104 gnd.n1241 739.952
R8105 gnd.n5224 gnd.n1172 739.952
R8106 gnd.n6795 gnd.n871 737.549
R8107 gnd.n7315 gnd.n559 737.549
R8108 gnd.n7531 gnd.n432 737.549
R8109 gnd.n5234 gnd.n1126 737.549
R8110 gnd.n6795 gnd.n6794 585
R8111 gnd.n6796 gnd.n6795 585
R8112 gnd.n6793 gnd.n873 585
R8113 gnd.n873 gnd.n872 585
R8114 gnd.n6792 gnd.n6791 585
R8115 gnd.n6791 gnd.n6790 585
R8116 gnd.n878 gnd.n877 585
R8117 gnd.n6789 gnd.n878 585
R8118 gnd.n6787 gnd.n6786 585
R8119 gnd.n6788 gnd.n6787 585
R8120 gnd.n6785 gnd.n880 585
R8121 gnd.n880 gnd.n879 585
R8122 gnd.n6784 gnd.n6783 585
R8123 gnd.n6783 gnd.n6782 585
R8124 gnd.n886 gnd.n885 585
R8125 gnd.n6781 gnd.n886 585
R8126 gnd.n6779 gnd.n6778 585
R8127 gnd.n6780 gnd.n6779 585
R8128 gnd.n6777 gnd.n888 585
R8129 gnd.n888 gnd.n887 585
R8130 gnd.n6776 gnd.n6775 585
R8131 gnd.n6775 gnd.n6774 585
R8132 gnd.n894 gnd.n893 585
R8133 gnd.n6773 gnd.n894 585
R8134 gnd.n6771 gnd.n6770 585
R8135 gnd.n6772 gnd.n6771 585
R8136 gnd.n6769 gnd.n896 585
R8137 gnd.n896 gnd.n895 585
R8138 gnd.n6768 gnd.n6767 585
R8139 gnd.n6767 gnd.n6766 585
R8140 gnd.n902 gnd.n901 585
R8141 gnd.n6765 gnd.n902 585
R8142 gnd.n6763 gnd.n6762 585
R8143 gnd.n6764 gnd.n6763 585
R8144 gnd.n6761 gnd.n904 585
R8145 gnd.n904 gnd.n903 585
R8146 gnd.n6760 gnd.n6759 585
R8147 gnd.n6759 gnd.n6758 585
R8148 gnd.n910 gnd.n909 585
R8149 gnd.n6757 gnd.n910 585
R8150 gnd.n6755 gnd.n6754 585
R8151 gnd.n6756 gnd.n6755 585
R8152 gnd.n6753 gnd.n912 585
R8153 gnd.n912 gnd.n911 585
R8154 gnd.n6752 gnd.n6751 585
R8155 gnd.n6751 gnd.n6750 585
R8156 gnd.n918 gnd.n917 585
R8157 gnd.n6749 gnd.n918 585
R8158 gnd.n6747 gnd.n6746 585
R8159 gnd.n6748 gnd.n6747 585
R8160 gnd.n6745 gnd.n920 585
R8161 gnd.n920 gnd.n919 585
R8162 gnd.n6744 gnd.n6743 585
R8163 gnd.n6743 gnd.n6742 585
R8164 gnd.n926 gnd.n925 585
R8165 gnd.n6741 gnd.n926 585
R8166 gnd.n6739 gnd.n6738 585
R8167 gnd.n6740 gnd.n6739 585
R8168 gnd.n6737 gnd.n928 585
R8169 gnd.n928 gnd.n927 585
R8170 gnd.n6736 gnd.n6735 585
R8171 gnd.n6735 gnd.n6734 585
R8172 gnd.n934 gnd.n933 585
R8173 gnd.n6733 gnd.n934 585
R8174 gnd.n6731 gnd.n6730 585
R8175 gnd.n6732 gnd.n6731 585
R8176 gnd.n6729 gnd.n936 585
R8177 gnd.n936 gnd.n935 585
R8178 gnd.n6728 gnd.n6727 585
R8179 gnd.n6727 gnd.n6726 585
R8180 gnd.n942 gnd.n941 585
R8181 gnd.n6725 gnd.n942 585
R8182 gnd.n6723 gnd.n6722 585
R8183 gnd.n6724 gnd.n6723 585
R8184 gnd.n6721 gnd.n944 585
R8185 gnd.n944 gnd.n943 585
R8186 gnd.n6720 gnd.n6719 585
R8187 gnd.n6719 gnd.n6718 585
R8188 gnd.n950 gnd.n949 585
R8189 gnd.n6717 gnd.n950 585
R8190 gnd.n6715 gnd.n6714 585
R8191 gnd.n6716 gnd.n6715 585
R8192 gnd.n6713 gnd.n952 585
R8193 gnd.n952 gnd.n951 585
R8194 gnd.n6712 gnd.n6711 585
R8195 gnd.n6711 gnd.n6710 585
R8196 gnd.n958 gnd.n957 585
R8197 gnd.n6709 gnd.n958 585
R8198 gnd.n6707 gnd.n6706 585
R8199 gnd.n6708 gnd.n6707 585
R8200 gnd.n6705 gnd.n960 585
R8201 gnd.n960 gnd.n959 585
R8202 gnd.n6704 gnd.n6703 585
R8203 gnd.n6703 gnd.n6702 585
R8204 gnd.n966 gnd.n965 585
R8205 gnd.n6701 gnd.n966 585
R8206 gnd.n6699 gnd.n6698 585
R8207 gnd.n6700 gnd.n6699 585
R8208 gnd.n6697 gnd.n968 585
R8209 gnd.n968 gnd.n967 585
R8210 gnd.n6696 gnd.n6695 585
R8211 gnd.n6695 gnd.n6694 585
R8212 gnd.n974 gnd.n973 585
R8213 gnd.n6693 gnd.n974 585
R8214 gnd.n6691 gnd.n6690 585
R8215 gnd.n6692 gnd.n6691 585
R8216 gnd.n6689 gnd.n976 585
R8217 gnd.n976 gnd.n975 585
R8218 gnd.n6688 gnd.n6687 585
R8219 gnd.n6687 gnd.n6686 585
R8220 gnd.n982 gnd.n981 585
R8221 gnd.n6685 gnd.n982 585
R8222 gnd.n6683 gnd.n6682 585
R8223 gnd.n6684 gnd.n6683 585
R8224 gnd.n6681 gnd.n984 585
R8225 gnd.n984 gnd.n983 585
R8226 gnd.n6680 gnd.n6679 585
R8227 gnd.n6679 gnd.n6678 585
R8228 gnd.n990 gnd.n989 585
R8229 gnd.n6677 gnd.n990 585
R8230 gnd.n6675 gnd.n6674 585
R8231 gnd.n6676 gnd.n6675 585
R8232 gnd.n6673 gnd.n992 585
R8233 gnd.n992 gnd.n991 585
R8234 gnd.n6672 gnd.n6671 585
R8235 gnd.n6671 gnd.n6670 585
R8236 gnd.n998 gnd.n997 585
R8237 gnd.n6669 gnd.n998 585
R8238 gnd.n6667 gnd.n6666 585
R8239 gnd.n6668 gnd.n6667 585
R8240 gnd.n6665 gnd.n1000 585
R8241 gnd.n1000 gnd.n999 585
R8242 gnd.n6664 gnd.n6663 585
R8243 gnd.n6663 gnd.n6662 585
R8244 gnd.n1006 gnd.n1005 585
R8245 gnd.n6661 gnd.n1006 585
R8246 gnd.n6659 gnd.n6658 585
R8247 gnd.n6660 gnd.n6659 585
R8248 gnd.n6657 gnd.n1008 585
R8249 gnd.n1008 gnd.n1007 585
R8250 gnd.n6656 gnd.n6655 585
R8251 gnd.n6655 gnd.n6654 585
R8252 gnd.n1014 gnd.n1013 585
R8253 gnd.n6653 gnd.n1014 585
R8254 gnd.n6651 gnd.n6650 585
R8255 gnd.n6652 gnd.n6651 585
R8256 gnd.n6649 gnd.n1016 585
R8257 gnd.n1016 gnd.n1015 585
R8258 gnd.n6648 gnd.n6647 585
R8259 gnd.n6647 gnd.n6646 585
R8260 gnd.n1022 gnd.n1021 585
R8261 gnd.n6645 gnd.n1022 585
R8262 gnd.n6643 gnd.n6642 585
R8263 gnd.n6644 gnd.n6643 585
R8264 gnd.n6641 gnd.n1024 585
R8265 gnd.n1024 gnd.n1023 585
R8266 gnd.n6640 gnd.n6639 585
R8267 gnd.n6639 gnd.n6638 585
R8268 gnd.n1030 gnd.n1029 585
R8269 gnd.n6637 gnd.n1030 585
R8270 gnd.n6635 gnd.n6634 585
R8271 gnd.n6636 gnd.n6635 585
R8272 gnd.n6633 gnd.n1032 585
R8273 gnd.n1032 gnd.n1031 585
R8274 gnd.n6632 gnd.n6631 585
R8275 gnd.n6631 gnd.n6630 585
R8276 gnd.n1038 gnd.n1037 585
R8277 gnd.n6629 gnd.n1038 585
R8278 gnd.n871 gnd.n870 585
R8279 gnd.n6797 gnd.n871 585
R8280 gnd.n6800 gnd.n6799 585
R8281 gnd.n6799 gnd.n6798 585
R8282 gnd.n868 gnd.n867 585
R8283 gnd.n867 gnd.n866 585
R8284 gnd.n6805 gnd.n6804 585
R8285 gnd.n6806 gnd.n6805 585
R8286 gnd.n865 gnd.n864 585
R8287 gnd.n6807 gnd.n865 585
R8288 gnd.n6810 gnd.n6809 585
R8289 gnd.n6809 gnd.n6808 585
R8290 gnd.n862 gnd.n861 585
R8291 gnd.n861 gnd.n860 585
R8292 gnd.n6815 gnd.n6814 585
R8293 gnd.n6816 gnd.n6815 585
R8294 gnd.n859 gnd.n858 585
R8295 gnd.n6817 gnd.n859 585
R8296 gnd.n6820 gnd.n6819 585
R8297 gnd.n6819 gnd.n6818 585
R8298 gnd.n856 gnd.n855 585
R8299 gnd.n855 gnd.n854 585
R8300 gnd.n6825 gnd.n6824 585
R8301 gnd.n6826 gnd.n6825 585
R8302 gnd.n853 gnd.n852 585
R8303 gnd.n6827 gnd.n853 585
R8304 gnd.n6830 gnd.n6829 585
R8305 gnd.n6829 gnd.n6828 585
R8306 gnd.n850 gnd.n849 585
R8307 gnd.n849 gnd.n848 585
R8308 gnd.n6835 gnd.n6834 585
R8309 gnd.n6836 gnd.n6835 585
R8310 gnd.n847 gnd.n846 585
R8311 gnd.n6837 gnd.n847 585
R8312 gnd.n6840 gnd.n6839 585
R8313 gnd.n6839 gnd.n6838 585
R8314 gnd.n844 gnd.n843 585
R8315 gnd.n843 gnd.n842 585
R8316 gnd.n6845 gnd.n6844 585
R8317 gnd.n6846 gnd.n6845 585
R8318 gnd.n841 gnd.n840 585
R8319 gnd.n6847 gnd.n841 585
R8320 gnd.n6850 gnd.n6849 585
R8321 gnd.n6849 gnd.n6848 585
R8322 gnd.n838 gnd.n837 585
R8323 gnd.n837 gnd.n836 585
R8324 gnd.n6855 gnd.n6854 585
R8325 gnd.n6856 gnd.n6855 585
R8326 gnd.n835 gnd.n834 585
R8327 gnd.n6857 gnd.n835 585
R8328 gnd.n6860 gnd.n6859 585
R8329 gnd.n6859 gnd.n6858 585
R8330 gnd.n832 gnd.n831 585
R8331 gnd.n831 gnd.n830 585
R8332 gnd.n6865 gnd.n6864 585
R8333 gnd.n6866 gnd.n6865 585
R8334 gnd.n829 gnd.n828 585
R8335 gnd.n6867 gnd.n829 585
R8336 gnd.n6870 gnd.n6869 585
R8337 gnd.n6869 gnd.n6868 585
R8338 gnd.n826 gnd.n825 585
R8339 gnd.n825 gnd.n824 585
R8340 gnd.n6875 gnd.n6874 585
R8341 gnd.n6876 gnd.n6875 585
R8342 gnd.n823 gnd.n822 585
R8343 gnd.n6877 gnd.n823 585
R8344 gnd.n6880 gnd.n6879 585
R8345 gnd.n6879 gnd.n6878 585
R8346 gnd.n820 gnd.n819 585
R8347 gnd.n819 gnd.n818 585
R8348 gnd.n6885 gnd.n6884 585
R8349 gnd.n6886 gnd.n6885 585
R8350 gnd.n817 gnd.n816 585
R8351 gnd.n6887 gnd.n817 585
R8352 gnd.n6890 gnd.n6889 585
R8353 gnd.n6889 gnd.n6888 585
R8354 gnd.n814 gnd.n813 585
R8355 gnd.n813 gnd.n812 585
R8356 gnd.n6895 gnd.n6894 585
R8357 gnd.n6896 gnd.n6895 585
R8358 gnd.n811 gnd.n810 585
R8359 gnd.n6897 gnd.n811 585
R8360 gnd.n6900 gnd.n6899 585
R8361 gnd.n6899 gnd.n6898 585
R8362 gnd.n808 gnd.n807 585
R8363 gnd.n807 gnd.n806 585
R8364 gnd.n6905 gnd.n6904 585
R8365 gnd.n6906 gnd.n6905 585
R8366 gnd.n805 gnd.n804 585
R8367 gnd.n6907 gnd.n805 585
R8368 gnd.n6910 gnd.n6909 585
R8369 gnd.n6909 gnd.n6908 585
R8370 gnd.n802 gnd.n801 585
R8371 gnd.n801 gnd.n800 585
R8372 gnd.n6915 gnd.n6914 585
R8373 gnd.n6916 gnd.n6915 585
R8374 gnd.n799 gnd.n798 585
R8375 gnd.n6917 gnd.n799 585
R8376 gnd.n6920 gnd.n6919 585
R8377 gnd.n6919 gnd.n6918 585
R8378 gnd.n796 gnd.n795 585
R8379 gnd.n795 gnd.n794 585
R8380 gnd.n6925 gnd.n6924 585
R8381 gnd.n6926 gnd.n6925 585
R8382 gnd.n793 gnd.n792 585
R8383 gnd.n6927 gnd.n793 585
R8384 gnd.n6930 gnd.n6929 585
R8385 gnd.n6929 gnd.n6928 585
R8386 gnd.n790 gnd.n789 585
R8387 gnd.n789 gnd.n788 585
R8388 gnd.n6935 gnd.n6934 585
R8389 gnd.n6936 gnd.n6935 585
R8390 gnd.n787 gnd.n786 585
R8391 gnd.n6937 gnd.n787 585
R8392 gnd.n6940 gnd.n6939 585
R8393 gnd.n6939 gnd.n6938 585
R8394 gnd.n784 gnd.n783 585
R8395 gnd.n783 gnd.n782 585
R8396 gnd.n6945 gnd.n6944 585
R8397 gnd.n6946 gnd.n6945 585
R8398 gnd.n781 gnd.n780 585
R8399 gnd.n6947 gnd.n781 585
R8400 gnd.n6950 gnd.n6949 585
R8401 gnd.n6949 gnd.n6948 585
R8402 gnd.n778 gnd.n777 585
R8403 gnd.n777 gnd.n776 585
R8404 gnd.n6955 gnd.n6954 585
R8405 gnd.n6956 gnd.n6955 585
R8406 gnd.n775 gnd.n774 585
R8407 gnd.n6957 gnd.n775 585
R8408 gnd.n6960 gnd.n6959 585
R8409 gnd.n6959 gnd.n6958 585
R8410 gnd.n772 gnd.n771 585
R8411 gnd.n771 gnd.n770 585
R8412 gnd.n6965 gnd.n6964 585
R8413 gnd.n6966 gnd.n6965 585
R8414 gnd.n769 gnd.n768 585
R8415 gnd.n6967 gnd.n769 585
R8416 gnd.n6970 gnd.n6969 585
R8417 gnd.n6969 gnd.n6968 585
R8418 gnd.n766 gnd.n765 585
R8419 gnd.n765 gnd.n764 585
R8420 gnd.n6975 gnd.n6974 585
R8421 gnd.n6976 gnd.n6975 585
R8422 gnd.n763 gnd.n762 585
R8423 gnd.n6977 gnd.n763 585
R8424 gnd.n6980 gnd.n6979 585
R8425 gnd.n6979 gnd.n6978 585
R8426 gnd.n760 gnd.n759 585
R8427 gnd.n759 gnd.n758 585
R8428 gnd.n6985 gnd.n6984 585
R8429 gnd.n6986 gnd.n6985 585
R8430 gnd.n757 gnd.n756 585
R8431 gnd.n6987 gnd.n757 585
R8432 gnd.n6990 gnd.n6989 585
R8433 gnd.n6989 gnd.n6988 585
R8434 gnd.n754 gnd.n753 585
R8435 gnd.n753 gnd.n752 585
R8436 gnd.n6995 gnd.n6994 585
R8437 gnd.n6996 gnd.n6995 585
R8438 gnd.n751 gnd.n750 585
R8439 gnd.n6997 gnd.n751 585
R8440 gnd.n7000 gnd.n6999 585
R8441 gnd.n6999 gnd.n6998 585
R8442 gnd.n748 gnd.n747 585
R8443 gnd.n747 gnd.n746 585
R8444 gnd.n7005 gnd.n7004 585
R8445 gnd.n7006 gnd.n7005 585
R8446 gnd.n745 gnd.n744 585
R8447 gnd.n7007 gnd.n745 585
R8448 gnd.n7010 gnd.n7009 585
R8449 gnd.n7009 gnd.n7008 585
R8450 gnd.n742 gnd.n741 585
R8451 gnd.n741 gnd.n740 585
R8452 gnd.n7015 gnd.n7014 585
R8453 gnd.n7016 gnd.n7015 585
R8454 gnd.n739 gnd.n738 585
R8455 gnd.n7017 gnd.n739 585
R8456 gnd.n7020 gnd.n7019 585
R8457 gnd.n7019 gnd.n7018 585
R8458 gnd.n736 gnd.n735 585
R8459 gnd.n735 gnd.n734 585
R8460 gnd.n7025 gnd.n7024 585
R8461 gnd.n7026 gnd.n7025 585
R8462 gnd.n733 gnd.n732 585
R8463 gnd.n7027 gnd.n733 585
R8464 gnd.n7030 gnd.n7029 585
R8465 gnd.n7029 gnd.n7028 585
R8466 gnd.n730 gnd.n729 585
R8467 gnd.n729 gnd.n728 585
R8468 gnd.n7035 gnd.n7034 585
R8469 gnd.n7036 gnd.n7035 585
R8470 gnd.n727 gnd.n726 585
R8471 gnd.n7037 gnd.n727 585
R8472 gnd.n7040 gnd.n7039 585
R8473 gnd.n7039 gnd.n7038 585
R8474 gnd.n724 gnd.n723 585
R8475 gnd.n723 gnd.n722 585
R8476 gnd.n7045 gnd.n7044 585
R8477 gnd.n7046 gnd.n7045 585
R8478 gnd.n721 gnd.n720 585
R8479 gnd.n7047 gnd.n721 585
R8480 gnd.n7050 gnd.n7049 585
R8481 gnd.n7049 gnd.n7048 585
R8482 gnd.n718 gnd.n717 585
R8483 gnd.n717 gnd.n716 585
R8484 gnd.n7055 gnd.n7054 585
R8485 gnd.n7056 gnd.n7055 585
R8486 gnd.n715 gnd.n714 585
R8487 gnd.n7057 gnd.n715 585
R8488 gnd.n7060 gnd.n7059 585
R8489 gnd.n7059 gnd.n7058 585
R8490 gnd.n712 gnd.n711 585
R8491 gnd.n711 gnd.n710 585
R8492 gnd.n7065 gnd.n7064 585
R8493 gnd.n7066 gnd.n7065 585
R8494 gnd.n709 gnd.n708 585
R8495 gnd.n7067 gnd.n709 585
R8496 gnd.n7070 gnd.n7069 585
R8497 gnd.n7069 gnd.n7068 585
R8498 gnd.n706 gnd.n705 585
R8499 gnd.n705 gnd.n704 585
R8500 gnd.n7075 gnd.n7074 585
R8501 gnd.n7076 gnd.n7075 585
R8502 gnd.n703 gnd.n702 585
R8503 gnd.n7077 gnd.n703 585
R8504 gnd.n7080 gnd.n7079 585
R8505 gnd.n7079 gnd.n7078 585
R8506 gnd.n700 gnd.n699 585
R8507 gnd.n699 gnd.n698 585
R8508 gnd.n7085 gnd.n7084 585
R8509 gnd.n7086 gnd.n7085 585
R8510 gnd.n697 gnd.n696 585
R8511 gnd.n7087 gnd.n697 585
R8512 gnd.n7090 gnd.n7089 585
R8513 gnd.n7089 gnd.n7088 585
R8514 gnd.n694 gnd.n693 585
R8515 gnd.n693 gnd.n692 585
R8516 gnd.n7095 gnd.n7094 585
R8517 gnd.n7096 gnd.n7095 585
R8518 gnd.n691 gnd.n690 585
R8519 gnd.n7097 gnd.n691 585
R8520 gnd.n7100 gnd.n7099 585
R8521 gnd.n7099 gnd.n7098 585
R8522 gnd.n688 gnd.n687 585
R8523 gnd.n687 gnd.n686 585
R8524 gnd.n7105 gnd.n7104 585
R8525 gnd.n7106 gnd.n7105 585
R8526 gnd.n685 gnd.n684 585
R8527 gnd.n7107 gnd.n685 585
R8528 gnd.n7110 gnd.n7109 585
R8529 gnd.n7109 gnd.n7108 585
R8530 gnd.n682 gnd.n681 585
R8531 gnd.n681 gnd.n680 585
R8532 gnd.n7115 gnd.n7114 585
R8533 gnd.n7116 gnd.n7115 585
R8534 gnd.n679 gnd.n678 585
R8535 gnd.n7117 gnd.n679 585
R8536 gnd.n7120 gnd.n7119 585
R8537 gnd.n7119 gnd.n7118 585
R8538 gnd.n676 gnd.n675 585
R8539 gnd.n675 gnd.n674 585
R8540 gnd.n7125 gnd.n7124 585
R8541 gnd.n7126 gnd.n7125 585
R8542 gnd.n673 gnd.n672 585
R8543 gnd.n7127 gnd.n673 585
R8544 gnd.n7130 gnd.n7129 585
R8545 gnd.n7129 gnd.n7128 585
R8546 gnd.n670 gnd.n669 585
R8547 gnd.n669 gnd.n668 585
R8548 gnd.n7135 gnd.n7134 585
R8549 gnd.n7136 gnd.n7135 585
R8550 gnd.n667 gnd.n666 585
R8551 gnd.n7137 gnd.n667 585
R8552 gnd.n7140 gnd.n7139 585
R8553 gnd.n7139 gnd.n7138 585
R8554 gnd.n664 gnd.n663 585
R8555 gnd.n663 gnd.n662 585
R8556 gnd.n7145 gnd.n7144 585
R8557 gnd.n7146 gnd.n7145 585
R8558 gnd.n661 gnd.n660 585
R8559 gnd.n7147 gnd.n661 585
R8560 gnd.n7150 gnd.n7149 585
R8561 gnd.n7149 gnd.n7148 585
R8562 gnd.n658 gnd.n657 585
R8563 gnd.n657 gnd.n656 585
R8564 gnd.n7155 gnd.n7154 585
R8565 gnd.n7156 gnd.n7155 585
R8566 gnd.n655 gnd.n654 585
R8567 gnd.n7157 gnd.n655 585
R8568 gnd.n7160 gnd.n7159 585
R8569 gnd.n7159 gnd.n7158 585
R8570 gnd.n652 gnd.n651 585
R8571 gnd.n651 gnd.n650 585
R8572 gnd.n7165 gnd.n7164 585
R8573 gnd.n7166 gnd.n7165 585
R8574 gnd.n649 gnd.n648 585
R8575 gnd.n7167 gnd.n649 585
R8576 gnd.n7170 gnd.n7169 585
R8577 gnd.n7169 gnd.n7168 585
R8578 gnd.n646 gnd.n645 585
R8579 gnd.n645 gnd.n644 585
R8580 gnd.n7175 gnd.n7174 585
R8581 gnd.n7176 gnd.n7175 585
R8582 gnd.n643 gnd.n642 585
R8583 gnd.n7177 gnd.n643 585
R8584 gnd.n7180 gnd.n7179 585
R8585 gnd.n7179 gnd.n7178 585
R8586 gnd.n640 gnd.n639 585
R8587 gnd.n639 gnd.n638 585
R8588 gnd.n7185 gnd.n7184 585
R8589 gnd.n7186 gnd.n7185 585
R8590 gnd.n637 gnd.n636 585
R8591 gnd.n7187 gnd.n637 585
R8592 gnd.n7190 gnd.n7189 585
R8593 gnd.n7189 gnd.n7188 585
R8594 gnd.n634 gnd.n633 585
R8595 gnd.n633 gnd.n632 585
R8596 gnd.n7195 gnd.n7194 585
R8597 gnd.n7196 gnd.n7195 585
R8598 gnd.n631 gnd.n630 585
R8599 gnd.n7197 gnd.n631 585
R8600 gnd.n7200 gnd.n7199 585
R8601 gnd.n7199 gnd.n7198 585
R8602 gnd.n628 gnd.n627 585
R8603 gnd.n627 gnd.n626 585
R8604 gnd.n7205 gnd.n7204 585
R8605 gnd.n7206 gnd.n7205 585
R8606 gnd.n625 gnd.n624 585
R8607 gnd.n7207 gnd.n625 585
R8608 gnd.n7210 gnd.n7209 585
R8609 gnd.n7209 gnd.n7208 585
R8610 gnd.n622 gnd.n621 585
R8611 gnd.n621 gnd.n620 585
R8612 gnd.n7215 gnd.n7214 585
R8613 gnd.n7216 gnd.n7215 585
R8614 gnd.n619 gnd.n618 585
R8615 gnd.n7217 gnd.n619 585
R8616 gnd.n7220 gnd.n7219 585
R8617 gnd.n7219 gnd.n7218 585
R8618 gnd.n616 gnd.n615 585
R8619 gnd.n615 gnd.n614 585
R8620 gnd.n7225 gnd.n7224 585
R8621 gnd.n7226 gnd.n7225 585
R8622 gnd.n613 gnd.n612 585
R8623 gnd.n7227 gnd.n613 585
R8624 gnd.n7230 gnd.n7229 585
R8625 gnd.n7229 gnd.n7228 585
R8626 gnd.n610 gnd.n609 585
R8627 gnd.n609 gnd.n608 585
R8628 gnd.n7235 gnd.n7234 585
R8629 gnd.n7236 gnd.n7235 585
R8630 gnd.n607 gnd.n606 585
R8631 gnd.n7237 gnd.n607 585
R8632 gnd.n7240 gnd.n7239 585
R8633 gnd.n7239 gnd.n7238 585
R8634 gnd.n604 gnd.n603 585
R8635 gnd.n603 gnd.n602 585
R8636 gnd.n7245 gnd.n7244 585
R8637 gnd.n7246 gnd.n7245 585
R8638 gnd.n601 gnd.n600 585
R8639 gnd.n7247 gnd.n601 585
R8640 gnd.n7250 gnd.n7249 585
R8641 gnd.n7249 gnd.n7248 585
R8642 gnd.n598 gnd.n597 585
R8643 gnd.n597 gnd.n596 585
R8644 gnd.n7255 gnd.n7254 585
R8645 gnd.n7256 gnd.n7255 585
R8646 gnd.n595 gnd.n594 585
R8647 gnd.n7257 gnd.n595 585
R8648 gnd.n7260 gnd.n7259 585
R8649 gnd.n7259 gnd.n7258 585
R8650 gnd.n592 gnd.n591 585
R8651 gnd.n591 gnd.n590 585
R8652 gnd.n7265 gnd.n7264 585
R8653 gnd.n7266 gnd.n7265 585
R8654 gnd.n589 gnd.n588 585
R8655 gnd.n7267 gnd.n589 585
R8656 gnd.n7270 gnd.n7269 585
R8657 gnd.n7269 gnd.n7268 585
R8658 gnd.n586 gnd.n585 585
R8659 gnd.n585 gnd.n584 585
R8660 gnd.n7275 gnd.n7274 585
R8661 gnd.n7276 gnd.n7275 585
R8662 gnd.n583 gnd.n582 585
R8663 gnd.n7277 gnd.n583 585
R8664 gnd.n7280 gnd.n7279 585
R8665 gnd.n7279 gnd.n7278 585
R8666 gnd.n580 gnd.n579 585
R8667 gnd.n579 gnd.n578 585
R8668 gnd.n7285 gnd.n7284 585
R8669 gnd.n7286 gnd.n7285 585
R8670 gnd.n577 gnd.n576 585
R8671 gnd.n7287 gnd.n577 585
R8672 gnd.n7290 gnd.n7289 585
R8673 gnd.n7289 gnd.n7288 585
R8674 gnd.n574 gnd.n573 585
R8675 gnd.n573 gnd.n572 585
R8676 gnd.n7295 gnd.n7294 585
R8677 gnd.n7296 gnd.n7295 585
R8678 gnd.n571 gnd.n570 585
R8679 gnd.n7297 gnd.n571 585
R8680 gnd.n7300 gnd.n7299 585
R8681 gnd.n7299 gnd.n7298 585
R8682 gnd.n568 gnd.n567 585
R8683 gnd.n567 gnd.n566 585
R8684 gnd.n7305 gnd.n7304 585
R8685 gnd.n7306 gnd.n7305 585
R8686 gnd.n565 gnd.n564 585
R8687 gnd.n7307 gnd.n565 585
R8688 gnd.n7310 gnd.n7309 585
R8689 gnd.n7309 gnd.n7308 585
R8690 gnd.n562 gnd.n561 585
R8691 gnd.n561 gnd.n560 585
R8692 gnd.n7315 gnd.n7314 585
R8693 gnd.n7316 gnd.n7315 585
R8694 gnd.n7527 gnd.n7526 585
R8695 gnd.n7528 gnd.n7527 585
R8696 gnd.n436 gnd.n435 585
R8697 gnd.n435 gnd.n434 585
R8698 gnd.n7520 gnd.n7519 585
R8699 gnd.n7519 gnd.n7518 585
R8700 gnd.n439 gnd.n438 585
R8701 gnd.n7517 gnd.n439 585
R8702 gnd.n7515 gnd.n7514 585
R8703 gnd.n7516 gnd.n7515 585
R8704 gnd.n442 gnd.n441 585
R8705 gnd.n441 gnd.n440 585
R8706 gnd.n7510 gnd.n7509 585
R8707 gnd.n7509 gnd.n7508 585
R8708 gnd.n445 gnd.n444 585
R8709 gnd.n7507 gnd.n445 585
R8710 gnd.n7505 gnd.n7504 585
R8711 gnd.n7506 gnd.n7505 585
R8712 gnd.n448 gnd.n447 585
R8713 gnd.n447 gnd.n446 585
R8714 gnd.n7500 gnd.n7499 585
R8715 gnd.n7499 gnd.n7498 585
R8716 gnd.n451 gnd.n450 585
R8717 gnd.n7497 gnd.n451 585
R8718 gnd.n7495 gnd.n7494 585
R8719 gnd.n7496 gnd.n7495 585
R8720 gnd.n454 gnd.n453 585
R8721 gnd.n453 gnd.n452 585
R8722 gnd.n7490 gnd.n7489 585
R8723 gnd.n7489 gnd.n7488 585
R8724 gnd.n457 gnd.n456 585
R8725 gnd.n7487 gnd.n457 585
R8726 gnd.n7485 gnd.n7484 585
R8727 gnd.n7486 gnd.n7485 585
R8728 gnd.n460 gnd.n459 585
R8729 gnd.n459 gnd.n458 585
R8730 gnd.n7480 gnd.n7479 585
R8731 gnd.n7479 gnd.n7478 585
R8732 gnd.n463 gnd.n462 585
R8733 gnd.n7477 gnd.n463 585
R8734 gnd.n7475 gnd.n7474 585
R8735 gnd.n7476 gnd.n7475 585
R8736 gnd.n466 gnd.n465 585
R8737 gnd.n465 gnd.n464 585
R8738 gnd.n7470 gnd.n7469 585
R8739 gnd.n7469 gnd.n7468 585
R8740 gnd.n469 gnd.n468 585
R8741 gnd.n7467 gnd.n469 585
R8742 gnd.n7465 gnd.n7464 585
R8743 gnd.n7466 gnd.n7465 585
R8744 gnd.n472 gnd.n471 585
R8745 gnd.n471 gnd.n470 585
R8746 gnd.n7460 gnd.n7459 585
R8747 gnd.n7459 gnd.n7458 585
R8748 gnd.n475 gnd.n474 585
R8749 gnd.n7457 gnd.n475 585
R8750 gnd.n7455 gnd.n7454 585
R8751 gnd.n7456 gnd.n7455 585
R8752 gnd.n478 gnd.n477 585
R8753 gnd.n477 gnd.n476 585
R8754 gnd.n7450 gnd.n7449 585
R8755 gnd.n7449 gnd.n7448 585
R8756 gnd.n481 gnd.n480 585
R8757 gnd.n7447 gnd.n481 585
R8758 gnd.n7445 gnd.n7444 585
R8759 gnd.n7446 gnd.n7445 585
R8760 gnd.n484 gnd.n483 585
R8761 gnd.n483 gnd.n482 585
R8762 gnd.n7440 gnd.n7439 585
R8763 gnd.n7439 gnd.n7438 585
R8764 gnd.n487 gnd.n486 585
R8765 gnd.n7437 gnd.n487 585
R8766 gnd.n7435 gnd.n7434 585
R8767 gnd.n7436 gnd.n7435 585
R8768 gnd.n490 gnd.n489 585
R8769 gnd.n489 gnd.n488 585
R8770 gnd.n7430 gnd.n7429 585
R8771 gnd.n7429 gnd.n7428 585
R8772 gnd.n493 gnd.n492 585
R8773 gnd.n7427 gnd.n493 585
R8774 gnd.n7425 gnd.n7424 585
R8775 gnd.n7426 gnd.n7425 585
R8776 gnd.n496 gnd.n495 585
R8777 gnd.n495 gnd.n494 585
R8778 gnd.n7420 gnd.n7419 585
R8779 gnd.n7419 gnd.n7418 585
R8780 gnd.n499 gnd.n498 585
R8781 gnd.n7417 gnd.n499 585
R8782 gnd.n7415 gnd.n7414 585
R8783 gnd.n7416 gnd.n7415 585
R8784 gnd.n502 gnd.n501 585
R8785 gnd.n501 gnd.n500 585
R8786 gnd.n7410 gnd.n7409 585
R8787 gnd.n7409 gnd.n7408 585
R8788 gnd.n505 gnd.n504 585
R8789 gnd.n7407 gnd.n505 585
R8790 gnd.n7405 gnd.n7404 585
R8791 gnd.n7406 gnd.n7405 585
R8792 gnd.n508 gnd.n507 585
R8793 gnd.n507 gnd.n506 585
R8794 gnd.n7400 gnd.n7399 585
R8795 gnd.n7399 gnd.n7398 585
R8796 gnd.n511 gnd.n510 585
R8797 gnd.n7397 gnd.n511 585
R8798 gnd.n7395 gnd.n7394 585
R8799 gnd.n7396 gnd.n7395 585
R8800 gnd.n514 gnd.n513 585
R8801 gnd.n513 gnd.n512 585
R8802 gnd.n7390 gnd.n7389 585
R8803 gnd.n7389 gnd.n7388 585
R8804 gnd.n517 gnd.n516 585
R8805 gnd.n7387 gnd.n517 585
R8806 gnd.n7385 gnd.n7384 585
R8807 gnd.n7386 gnd.n7385 585
R8808 gnd.n520 gnd.n519 585
R8809 gnd.n519 gnd.n518 585
R8810 gnd.n7380 gnd.n7379 585
R8811 gnd.n7379 gnd.n7378 585
R8812 gnd.n523 gnd.n522 585
R8813 gnd.n7377 gnd.n523 585
R8814 gnd.n7375 gnd.n7374 585
R8815 gnd.n7376 gnd.n7375 585
R8816 gnd.n526 gnd.n525 585
R8817 gnd.n525 gnd.n524 585
R8818 gnd.n7370 gnd.n7369 585
R8819 gnd.n7369 gnd.n7368 585
R8820 gnd.n529 gnd.n528 585
R8821 gnd.n7367 gnd.n529 585
R8822 gnd.n7365 gnd.n7364 585
R8823 gnd.n7366 gnd.n7365 585
R8824 gnd.n532 gnd.n531 585
R8825 gnd.n531 gnd.n530 585
R8826 gnd.n7360 gnd.n7359 585
R8827 gnd.n7359 gnd.n7358 585
R8828 gnd.n535 gnd.n534 585
R8829 gnd.n7357 gnd.n535 585
R8830 gnd.n7355 gnd.n7354 585
R8831 gnd.n7356 gnd.n7355 585
R8832 gnd.n538 gnd.n537 585
R8833 gnd.n537 gnd.n536 585
R8834 gnd.n7350 gnd.n7349 585
R8835 gnd.n7349 gnd.n7348 585
R8836 gnd.n541 gnd.n540 585
R8837 gnd.n7347 gnd.n541 585
R8838 gnd.n7345 gnd.n7344 585
R8839 gnd.n7346 gnd.n7345 585
R8840 gnd.n544 gnd.n543 585
R8841 gnd.n543 gnd.n542 585
R8842 gnd.n7340 gnd.n7339 585
R8843 gnd.n7339 gnd.n7338 585
R8844 gnd.n547 gnd.n546 585
R8845 gnd.n7337 gnd.n547 585
R8846 gnd.n7335 gnd.n7334 585
R8847 gnd.n7336 gnd.n7335 585
R8848 gnd.n550 gnd.n549 585
R8849 gnd.n549 gnd.n548 585
R8850 gnd.n7330 gnd.n7329 585
R8851 gnd.n7329 gnd.n7328 585
R8852 gnd.n553 gnd.n552 585
R8853 gnd.n7327 gnd.n553 585
R8854 gnd.n7325 gnd.n7324 585
R8855 gnd.n7326 gnd.n7325 585
R8856 gnd.n556 gnd.n555 585
R8857 gnd.n555 gnd.n554 585
R8858 gnd.n7320 gnd.n7319 585
R8859 gnd.n7319 gnd.n7318 585
R8860 gnd.n559 gnd.n558 585
R8861 gnd.n7317 gnd.n559 585
R8862 gnd.n4968 gnd.n4967 585
R8863 gnd.n4967 gnd.n4966 585
R8864 gnd.n4969 gnd.n1474 585
R8865 gnd.n3140 gnd.n1474 585
R8866 gnd.n4971 gnd.n4970 585
R8867 gnd.n4972 gnd.n4971 585
R8868 gnd.n1458 gnd.n1457 585
R8869 gnd.n3133 gnd.n1458 585
R8870 gnd.n4980 gnd.n4979 585
R8871 gnd.n4979 gnd.n4978 585
R8872 gnd.n4981 gnd.n1453 585
R8873 gnd.n3124 gnd.n1453 585
R8874 gnd.n4983 gnd.n4982 585
R8875 gnd.n4984 gnd.n4983 585
R8876 gnd.n1438 gnd.n1437 585
R8877 gnd.n3118 gnd.n1438 585
R8878 gnd.n4992 gnd.n4991 585
R8879 gnd.n4991 gnd.n4990 585
R8880 gnd.n4993 gnd.n1433 585
R8881 gnd.n3049 gnd.n1433 585
R8882 gnd.n4995 gnd.n4994 585
R8883 gnd.n4996 gnd.n4995 585
R8884 gnd.n1418 gnd.n1417 585
R8885 gnd.n3043 gnd.n1418 585
R8886 gnd.n5004 gnd.n5003 585
R8887 gnd.n5003 gnd.n5002 585
R8888 gnd.n5005 gnd.n1413 585
R8889 gnd.n3037 gnd.n1413 585
R8890 gnd.n5007 gnd.n5006 585
R8891 gnd.n5008 gnd.n5007 585
R8892 gnd.n1398 gnd.n1397 585
R8893 gnd.n3066 gnd.n1398 585
R8894 gnd.n5016 gnd.n5015 585
R8895 gnd.n5015 gnd.n5014 585
R8896 gnd.n5017 gnd.n1393 585
R8897 gnd.n3030 gnd.n1393 585
R8898 gnd.n5019 gnd.n5018 585
R8899 gnd.n5020 gnd.n5019 585
R8900 gnd.n1379 gnd.n1378 585
R8901 gnd.n3022 gnd.n1379 585
R8902 gnd.n5028 gnd.n5027 585
R8903 gnd.n5027 gnd.n5026 585
R8904 gnd.n5029 gnd.n1373 585
R8905 gnd.n3015 gnd.n1373 585
R8906 gnd.n5031 gnd.n5030 585
R8907 gnd.n5032 gnd.n5031 585
R8908 gnd.n1374 gnd.n1372 585
R8909 gnd.n3007 gnd.n1372 585
R8910 gnd.n2968 gnd.n2656 585
R8911 gnd.n2978 gnd.n2656 585
R8912 gnd.n2969 gnd.n2665 585
R8913 gnd.n2665 gnd.n2654 585
R8914 gnd.n2971 gnd.n2970 585
R8915 gnd.n2972 gnd.n2971 585
R8916 gnd.n2666 gnd.n2664 585
R8917 gnd.n2959 gnd.n2664 585
R8918 gnd.n2941 gnd.n2940 585
R8919 gnd.n2942 gnd.n2941 585
R8920 gnd.n2685 gnd.n2681 585
R8921 gnd.n2945 gnd.n2681 585
R8922 gnd.n2933 gnd.n2932 585
R8923 gnd.n2934 gnd.n2933 585
R8924 gnd.n1350 gnd.n1349 585
R8925 gnd.n2690 gnd.n1350 585
R8926 gnd.n5042 gnd.n5041 585
R8927 gnd.n5041 gnd.n5040 585
R8928 gnd.n5043 gnd.n1345 585
R8929 gnd.n2883 gnd.n1345 585
R8930 gnd.n5045 gnd.n5044 585
R8931 gnd.n5046 gnd.n5045 585
R8932 gnd.n1329 gnd.n1328 585
R8933 gnd.n2889 gnd.n1329 585
R8934 gnd.n5054 gnd.n5053 585
R8935 gnd.n5053 gnd.n5052 585
R8936 gnd.n5055 gnd.n1324 585
R8937 gnd.n2895 gnd.n1324 585
R8938 gnd.n5057 gnd.n5056 585
R8939 gnd.n5058 gnd.n5057 585
R8940 gnd.n1309 gnd.n1308 585
R8941 gnd.n2901 gnd.n1309 585
R8942 gnd.n5066 gnd.n5065 585
R8943 gnd.n5065 gnd.n5064 585
R8944 gnd.n5067 gnd.n1304 585
R8945 gnd.n2862 gnd.n1304 585
R8946 gnd.n5069 gnd.n5068 585
R8947 gnd.n5070 gnd.n5069 585
R8948 gnd.n1288 gnd.n1287 585
R8949 gnd.n2853 gnd.n1288 585
R8950 gnd.n5078 gnd.n5077 585
R8951 gnd.n5077 gnd.n5076 585
R8952 gnd.n5079 gnd.n1283 585
R8953 gnd.n2846 gnd.n1283 585
R8954 gnd.n5081 gnd.n5080 585
R8955 gnd.n5082 gnd.n5081 585
R8956 gnd.n1268 gnd.n1267 585
R8957 gnd.n2838 gnd.n1268 585
R8958 gnd.n5090 gnd.n5089 585
R8959 gnd.n5089 gnd.n5088 585
R8960 gnd.n5091 gnd.n1262 585
R8961 gnd.n2788 gnd.n1262 585
R8962 gnd.n5093 gnd.n5092 585
R8963 gnd.n5094 gnd.n5093 585
R8964 gnd.n1263 gnd.n1246 585
R8965 gnd.n2780 gnd.n1246 585
R8966 gnd.n5101 gnd.n1247 585
R8967 gnd.n5101 gnd.n5100 585
R8968 gnd.n5102 gnd.n1238 585
R8969 gnd.n5103 gnd.n5102 585
R8970 gnd.n2732 gnd.n1245 585
R8971 gnd.n2734 gnd.n2733 585
R8972 gnd.n2736 gnd.n2735 585
R8973 gnd.n2740 gnd.n2730 585
R8974 gnd.n2742 gnd.n2741 585
R8975 gnd.n2744 gnd.n2743 585
R8976 gnd.n2746 gnd.n2745 585
R8977 gnd.n2750 gnd.n2728 585
R8978 gnd.n2752 gnd.n2751 585
R8979 gnd.n2754 gnd.n2753 585
R8980 gnd.n2756 gnd.n2755 585
R8981 gnd.n2760 gnd.n2726 585
R8982 gnd.n2762 gnd.n2761 585
R8983 gnd.n2764 gnd.n2763 585
R8984 gnd.n2766 gnd.n2765 585
R8985 gnd.n2723 gnd.n2722 585
R8986 gnd.n2770 gnd.n2724 585
R8987 gnd.n2771 gnd.n2719 585
R8988 gnd.n2772 gnd.n1168 585
R8989 gnd.n5226 gnd.n1168 585
R8990 gnd.n3161 gnd.n3160 585
R8991 gnd.n3162 gnd.n2606 585
R8992 gnd.n3163 gnd.n2602 585
R8993 gnd.n2600 gnd.n2591 585
R8994 gnd.n3170 gnd.n2590 585
R8995 gnd.n3171 gnd.n2588 585
R8996 gnd.n2587 gnd.n2580 585
R8997 gnd.n3178 gnd.n2579 585
R8998 gnd.n3179 gnd.n2578 585
R8999 gnd.n2576 gnd.n2568 585
R9000 gnd.n3186 gnd.n2567 585
R9001 gnd.n3187 gnd.n2565 585
R9002 gnd.n2564 gnd.n2557 585
R9003 gnd.n3194 gnd.n2556 585
R9004 gnd.n3195 gnd.n2555 585
R9005 gnd.n2553 gnd.n2545 585
R9006 gnd.n3202 gnd.n2544 585
R9007 gnd.n3203 gnd.n2542 585
R9008 gnd.n2541 gnd.n1478 585
R9009 gnd.n1487 gnd.n1478 585
R9010 gnd.n3143 gnd.n1481 585
R9011 gnd.n4966 gnd.n1481 585
R9012 gnd.n3142 gnd.n3141 585
R9013 gnd.n3141 gnd.n3140 585
R9014 gnd.n2609 gnd.n1472 585
R9015 gnd.n4972 gnd.n1472 585
R9016 gnd.n3132 gnd.n3131 585
R9017 gnd.n3133 gnd.n3132 585
R9018 gnd.n2612 gnd.n1461 585
R9019 gnd.n4978 gnd.n1461 585
R9020 gnd.n3126 gnd.n3125 585
R9021 gnd.n3125 gnd.n3124 585
R9022 gnd.n2614 gnd.n1451 585
R9023 gnd.n4984 gnd.n1451 585
R9024 gnd.n3052 gnd.n2617 585
R9025 gnd.n3118 gnd.n2617 585
R9026 gnd.n3053 gnd.n1441 585
R9027 gnd.n4990 gnd.n1441 585
R9028 gnd.n3054 gnd.n3050 585
R9029 gnd.n3050 gnd.n3049 585
R9030 gnd.n2636 gnd.n1431 585
R9031 gnd.n4996 gnd.n1431 585
R9032 gnd.n3058 gnd.n2635 585
R9033 gnd.n3043 gnd.n2635 585
R9034 gnd.n3059 gnd.n1421 585
R9035 gnd.n5002 gnd.n1421 585
R9036 gnd.n3060 gnd.n2634 585
R9037 gnd.n3037 gnd.n2634 585
R9038 gnd.n2631 gnd.n1411 585
R9039 gnd.n5008 gnd.n1411 585
R9040 gnd.n3065 gnd.n3064 585
R9041 gnd.n3066 gnd.n3065 585
R9042 gnd.n2630 gnd.n1401 585
R9043 gnd.n5014 gnd.n1401 585
R9044 gnd.n3029 gnd.n3028 585
R9045 gnd.n3030 gnd.n3029 585
R9046 gnd.n2639 gnd.n1391 585
R9047 gnd.n5020 gnd.n1391 585
R9048 gnd.n3024 gnd.n3023 585
R9049 gnd.n3023 gnd.n3022 585
R9050 gnd.n2641 gnd.n1382 585
R9051 gnd.n5026 gnd.n1382 585
R9052 gnd.n3014 gnd.n3013 585
R9053 gnd.n3015 gnd.n3014 585
R9054 gnd.n2644 gnd.n1370 585
R9055 gnd.n5032 gnd.n1370 585
R9056 gnd.n3009 gnd.n3008 585
R9057 gnd.n3008 gnd.n3007 585
R9058 gnd.n2647 gnd.n2646 585
R9059 gnd.n2978 gnd.n2647 585
R9060 gnd.n2952 gnd.n2951 585
R9061 gnd.n2951 gnd.n2654 585
R9062 gnd.n2956 gnd.n2662 585
R9063 gnd.n2972 gnd.n2662 585
R9064 gnd.n2958 gnd.n2957 585
R9065 gnd.n2959 gnd.n2958 585
R9066 gnd.n2674 gnd.n2673 585
R9067 gnd.n2942 gnd.n2673 585
R9068 gnd.n2947 gnd.n2946 585
R9069 gnd.n2946 gnd.n2945 585
R9070 gnd.n2677 gnd.n2676 585
R9071 gnd.n2934 gnd.n2677 585
R9072 gnd.n2878 gnd.n2877 585
R9073 gnd.n2877 gnd.n2690 585
R9074 gnd.n2879 gnd.n1353 585
R9075 gnd.n5040 gnd.n1353 585
R9076 gnd.n2885 gnd.n2884 585
R9077 gnd.n2884 gnd.n2883 585
R9078 gnd.n2886 gnd.n1343 585
R9079 gnd.n5046 gnd.n1343 585
R9080 gnd.n2888 gnd.n2887 585
R9081 gnd.n2889 gnd.n2888 585
R9082 gnd.n2706 gnd.n1332 585
R9083 gnd.n5052 gnd.n1332 585
R9084 gnd.n2897 gnd.n2896 585
R9085 gnd.n2896 gnd.n2895 585
R9086 gnd.n2898 gnd.n1322 585
R9087 gnd.n5058 gnd.n1322 585
R9088 gnd.n2900 gnd.n2899 585
R9089 gnd.n2901 gnd.n2900 585
R9090 gnd.n2702 gnd.n1312 585
R9091 gnd.n5064 gnd.n1312 585
R9092 gnd.n2861 gnd.n2860 585
R9093 gnd.n2862 gnd.n2861 585
R9094 gnd.n2708 gnd.n1302 585
R9095 gnd.n5070 gnd.n1302 585
R9096 gnd.n2855 gnd.n2854 585
R9097 gnd.n2854 gnd.n2853 585
R9098 gnd.n2710 gnd.n1291 585
R9099 gnd.n5076 gnd.n1291 585
R9100 gnd.n2845 gnd.n2844 585
R9101 gnd.n2846 gnd.n2845 585
R9102 gnd.n2712 gnd.n1281 585
R9103 gnd.n5082 gnd.n1281 585
R9104 gnd.n2840 gnd.n2839 585
R9105 gnd.n2839 gnd.n2838 585
R9106 gnd.n2714 gnd.n1271 585
R9107 gnd.n5088 gnd.n1271 585
R9108 gnd.n2787 gnd.n2786 585
R9109 gnd.n2788 gnd.n2787 585
R9110 gnd.n2716 gnd.n1260 585
R9111 gnd.n5094 gnd.n1260 585
R9112 gnd.n2782 gnd.n2781 585
R9113 gnd.n2781 gnd.n2780 585
R9114 gnd.n2776 gnd.n1248 585
R9115 gnd.n5100 gnd.n1248 585
R9116 gnd.n2775 gnd.n1243 585
R9117 gnd.n5103 gnd.n1243 585
R9118 gnd.n6581 gnd.n6580 585
R9119 gnd.n6580 gnd.n6579 585
R9120 gnd.n6582 gnd.n1116 585
R9121 gnd.n6489 gnd.n1116 585
R9122 gnd.n6584 gnd.n6583 585
R9123 gnd.n6585 gnd.n6584 585
R9124 gnd.n1117 gnd.n1115 585
R9125 gnd.n1115 gnd.n1111 585
R9126 gnd.n1096 gnd.n1095 585
R9127 gnd.n1100 gnd.n1096 585
R9128 gnd.n6595 gnd.n6594 585
R9129 gnd.n6594 gnd.n6593 585
R9130 gnd.n6596 gnd.n1090 585
R9131 gnd.n6478 gnd.n1090 585
R9132 gnd.n6598 gnd.n6597 585
R9133 gnd.n6599 gnd.n6598 585
R9134 gnd.n1091 gnd.n1089 585
R9135 gnd.n1089 gnd.n1085 585
R9136 gnd.n1071 gnd.n1070 585
R9137 gnd.n6471 gnd.n1071 585
R9138 gnd.n6609 gnd.n6608 585
R9139 gnd.n6608 gnd.n6607 585
R9140 gnd.n6610 gnd.n1065 585
R9141 gnd.n6138 gnd.n1065 585
R9142 gnd.n6612 gnd.n6611 585
R9143 gnd.n6613 gnd.n6612 585
R9144 gnd.n1066 gnd.n1064 585
R9145 gnd.n1064 gnd.n1060 585
R9146 gnd.n1048 gnd.n1047 585
R9147 gnd.n6146 gnd.n1048 585
R9148 gnd.n6623 gnd.n6622 585
R9149 gnd.n6622 gnd.n6621 585
R9150 gnd.n6624 gnd.n1042 585
R9151 gnd.n5330 gnd.n1042 585
R9152 gnd.n6626 gnd.n6625 585
R9153 gnd.n6627 gnd.n6626 585
R9154 gnd.n1043 gnd.n1041 585
R9155 gnd.n6155 gnd.n1041 585
R9156 gnd.n6120 gnd.n5346 585
R9157 gnd.n5346 gnd.n5336 585
R9158 gnd.n6122 gnd.n6121 585
R9159 gnd.n6123 gnd.n6122 585
R9160 gnd.n5347 gnd.n5345 585
R9161 gnd.n5355 gnd.n5345 585
R9162 gnd.n6096 gnd.n5367 585
R9163 gnd.n5367 gnd.n5354 585
R9164 gnd.n6098 gnd.n6097 585
R9165 gnd.n6099 gnd.n6098 585
R9166 gnd.n5368 gnd.n5366 585
R9167 gnd.n5366 gnd.n5362 585
R9168 gnd.n6084 gnd.n6083 585
R9169 gnd.n6083 gnd.n6082 585
R9170 gnd.n5373 gnd.n5372 585
R9171 gnd.n5382 gnd.n5373 585
R9172 gnd.n6073 gnd.n6072 585
R9173 gnd.n6072 gnd.n6071 585
R9174 gnd.n5380 gnd.n5379 585
R9175 gnd.n6059 gnd.n5380 585
R9176 gnd.n5497 gnd.n5496 585
R9177 gnd.n5497 gnd.n5389 585
R9178 gnd.n6016 gnd.n6015 585
R9179 gnd.n6015 gnd.n6014 585
R9180 gnd.n6017 gnd.n5491 585
R9181 gnd.n5502 gnd.n5491 585
R9182 gnd.n6019 gnd.n6018 585
R9183 gnd.n6020 gnd.n6019 585
R9184 gnd.n5492 gnd.n5490 585
R9185 gnd.n5515 gnd.n5490 585
R9186 gnd.n5475 gnd.n5474 585
R9187 gnd.n5478 gnd.n5475 585
R9188 gnd.n6030 gnd.n6029 585
R9189 gnd.n6029 gnd.n6028 585
R9190 gnd.n6031 gnd.n5469 585
R9191 gnd.n5990 gnd.n5469 585
R9192 gnd.n6033 gnd.n6032 585
R9193 gnd.n6034 gnd.n6033 585
R9194 gnd.n5470 gnd.n5468 585
R9195 gnd.n5529 gnd.n5468 585
R9196 gnd.n5982 gnd.n5981 585
R9197 gnd.n5981 gnd.n5980 585
R9198 gnd.n5526 gnd.n5525 585
R9199 gnd.n5964 gnd.n5526 585
R9200 gnd.n5951 gnd.n5545 585
R9201 gnd.n5545 gnd.n5544 585
R9202 gnd.n5953 gnd.n5952 585
R9203 gnd.n5954 gnd.n5953 585
R9204 gnd.n5546 gnd.n5543 585
R9205 gnd.n5552 gnd.n5543 585
R9206 gnd.n5932 gnd.n5931 585
R9207 gnd.n5933 gnd.n5932 585
R9208 gnd.n5563 gnd.n5562 585
R9209 gnd.n5562 gnd.n5558 585
R9210 gnd.n5922 gnd.n5921 585
R9211 gnd.n5923 gnd.n5922 585
R9212 gnd.n5573 gnd.n5572 585
R9213 gnd.n5578 gnd.n5572 585
R9214 gnd.n5900 gnd.n5591 585
R9215 gnd.n5591 gnd.n5577 585
R9216 gnd.n5902 gnd.n5901 585
R9217 gnd.n5903 gnd.n5902 585
R9218 gnd.n5592 gnd.n5590 585
R9219 gnd.n5590 gnd.n5586 585
R9220 gnd.n5891 gnd.n5890 585
R9221 gnd.n5892 gnd.n5891 585
R9222 gnd.n5599 gnd.n5598 585
R9223 gnd.n5603 gnd.n5598 585
R9224 gnd.n5868 gnd.n5620 585
R9225 gnd.n5620 gnd.n5602 585
R9226 gnd.n5870 gnd.n5869 585
R9227 gnd.n5871 gnd.n5870 585
R9228 gnd.n5621 gnd.n5619 585
R9229 gnd.n5619 gnd.n5610 585
R9230 gnd.n5863 gnd.n5862 585
R9231 gnd.n5862 gnd.n5861 585
R9232 gnd.n5668 gnd.n5667 585
R9233 gnd.n5669 gnd.n5668 585
R9234 gnd.n5822 gnd.n5821 585
R9235 gnd.n5823 gnd.n5822 585
R9236 gnd.n5678 gnd.n5677 585
R9237 gnd.n5677 gnd.n5676 585
R9238 gnd.n5817 gnd.n5816 585
R9239 gnd.n5816 gnd.n5815 585
R9240 gnd.n5681 gnd.n5680 585
R9241 gnd.n5682 gnd.n5681 585
R9242 gnd.n5806 gnd.n5805 585
R9243 gnd.n5807 gnd.n5806 585
R9244 gnd.n5689 gnd.n5688 585
R9245 gnd.n5798 gnd.n5688 585
R9246 gnd.n5801 gnd.n5800 585
R9247 gnd.n5800 gnd.n5799 585
R9248 gnd.n5692 gnd.n5691 585
R9249 gnd.n5693 gnd.n5692 585
R9250 gnd.n5787 gnd.n5786 585
R9251 gnd.n5785 gnd.n5711 585
R9252 gnd.n5784 gnd.n5710 585
R9253 gnd.n5789 gnd.n5710 585
R9254 gnd.n5783 gnd.n5782 585
R9255 gnd.n5781 gnd.n5780 585
R9256 gnd.n5779 gnd.n5778 585
R9257 gnd.n5777 gnd.n5776 585
R9258 gnd.n5775 gnd.n5774 585
R9259 gnd.n5773 gnd.n5772 585
R9260 gnd.n5771 gnd.n5770 585
R9261 gnd.n5769 gnd.n5768 585
R9262 gnd.n5767 gnd.n5766 585
R9263 gnd.n5765 gnd.n5764 585
R9264 gnd.n5763 gnd.n5762 585
R9265 gnd.n5761 gnd.n5760 585
R9266 gnd.n5759 gnd.n5758 585
R9267 gnd.n5757 gnd.n5756 585
R9268 gnd.n5755 gnd.n5754 585
R9269 gnd.n5753 gnd.n5752 585
R9270 gnd.n5751 gnd.n5750 585
R9271 gnd.n5749 gnd.n5748 585
R9272 gnd.n5747 gnd.n5746 585
R9273 gnd.n5745 gnd.n5744 585
R9274 gnd.n5743 gnd.n5742 585
R9275 gnd.n5741 gnd.n5740 585
R9276 gnd.n5698 gnd.n5697 585
R9277 gnd.n5792 gnd.n5791 585
R9278 gnd.n6497 gnd.n6496 585
R9279 gnd.n6498 gnd.n5315 585
R9280 gnd.n6500 gnd.n6499 585
R9281 gnd.n6502 gnd.n5314 585
R9282 gnd.n6504 gnd.n6503 585
R9283 gnd.n6505 gnd.n5305 585
R9284 gnd.n6507 gnd.n6506 585
R9285 gnd.n6509 gnd.n5303 585
R9286 gnd.n6511 gnd.n6510 585
R9287 gnd.n6512 gnd.n5298 585
R9288 gnd.n6514 gnd.n6513 585
R9289 gnd.n6516 gnd.n5296 585
R9290 gnd.n6518 gnd.n6517 585
R9291 gnd.n6519 gnd.n5291 585
R9292 gnd.n6521 gnd.n6520 585
R9293 gnd.n6523 gnd.n5289 585
R9294 gnd.n6525 gnd.n6524 585
R9295 gnd.n6526 gnd.n5284 585
R9296 gnd.n6528 gnd.n6527 585
R9297 gnd.n6530 gnd.n5282 585
R9298 gnd.n6532 gnd.n6531 585
R9299 gnd.n6533 gnd.n5277 585
R9300 gnd.n6535 gnd.n6534 585
R9301 gnd.n6537 gnd.n5275 585
R9302 gnd.n6539 gnd.n6538 585
R9303 gnd.n6540 gnd.n5273 585
R9304 gnd.n6541 gnd.n1121 585
R9305 gnd.n5236 gnd.n1121 585
R9306 gnd.n6492 gnd.n1123 585
R9307 gnd.n6579 gnd.n1123 585
R9308 gnd.n6491 gnd.n6490 585
R9309 gnd.n6490 gnd.n6489 585
R9310 gnd.n6488 gnd.n1113 585
R9311 gnd.n6585 gnd.n1113 585
R9312 gnd.n6482 gnd.n5320 585
R9313 gnd.n6482 gnd.n1111 585
R9314 gnd.n6484 gnd.n6483 585
R9315 gnd.n6483 gnd.n1100 585
R9316 gnd.n6481 gnd.n1098 585
R9317 gnd.n6593 gnd.n1098 585
R9318 gnd.n6480 gnd.n6479 585
R9319 gnd.n6479 gnd.n6478 585
R9320 gnd.n5322 gnd.n1087 585
R9321 gnd.n6599 gnd.n1087 585
R9322 gnd.n6474 gnd.n6473 585
R9323 gnd.n6473 gnd.n1085 585
R9324 gnd.n6472 gnd.n5324 585
R9325 gnd.n6472 gnd.n6471 585
R9326 gnd.n6137 gnd.n1073 585
R9327 gnd.n6607 gnd.n1073 585
R9328 gnd.n6140 gnd.n6139 585
R9329 gnd.n6139 gnd.n6138 585
R9330 gnd.n6141 gnd.n1062 585
R9331 gnd.n6613 gnd.n1062 585
R9332 gnd.n6143 gnd.n6142 585
R9333 gnd.n6143 gnd.n1060 585
R9334 gnd.n6148 gnd.n6147 585
R9335 gnd.n6147 gnd.n6146 585
R9336 gnd.n6149 gnd.n1050 585
R9337 gnd.n6621 gnd.n1050 585
R9338 gnd.n6151 gnd.n6150 585
R9339 gnd.n6150 gnd.n5330 585
R9340 gnd.n6152 gnd.n1040 585
R9341 gnd.n6627 gnd.n1040 585
R9342 gnd.n6154 gnd.n6153 585
R9343 gnd.n6155 gnd.n6154 585
R9344 gnd.n5339 gnd.n5338 585
R9345 gnd.n5338 gnd.n5336 585
R9346 gnd.n6125 gnd.n6124 585
R9347 gnd.n6124 gnd.n6123 585
R9348 gnd.n5342 gnd.n5341 585
R9349 gnd.n5355 gnd.n5342 585
R9350 gnd.n6047 gnd.n6046 585
R9351 gnd.n6046 gnd.n5354 585
R9352 gnd.n6048 gnd.n5364 585
R9353 gnd.n6099 gnd.n5364 585
R9354 gnd.n6050 gnd.n6049 585
R9355 gnd.n6049 gnd.n5362 585
R9356 gnd.n6051 gnd.n5375 585
R9357 gnd.n6082 gnd.n5375 585
R9358 gnd.n6053 gnd.n6052 585
R9359 gnd.n6052 gnd.n5382 585
R9360 gnd.n6054 gnd.n5381 585
R9361 gnd.n6071 gnd.n5381 585
R9362 gnd.n6056 gnd.n6055 585
R9363 gnd.n6059 gnd.n6056 585
R9364 gnd.n5392 gnd.n5391 585
R9365 gnd.n5391 gnd.n5389 585
R9366 gnd.n5499 gnd.n5498 585
R9367 gnd.n6014 gnd.n5498 585
R9368 gnd.n5501 gnd.n5500 585
R9369 gnd.n5502 gnd.n5501 585
R9370 gnd.n5512 gnd.n5488 585
R9371 gnd.n6020 gnd.n5488 585
R9372 gnd.n5514 gnd.n5513 585
R9373 gnd.n5515 gnd.n5514 585
R9374 gnd.n5511 gnd.n5510 585
R9375 gnd.n5511 gnd.n5478 585
R9376 gnd.n5509 gnd.n5476 585
R9377 gnd.n6028 gnd.n5476 585
R9378 gnd.n5465 gnd.n5463 585
R9379 gnd.n5990 gnd.n5465 585
R9380 gnd.n6036 gnd.n6035 585
R9381 gnd.n6035 gnd.n6034 585
R9382 gnd.n5464 gnd.n5462 585
R9383 gnd.n5529 gnd.n5464 585
R9384 gnd.n5961 gnd.n5528 585
R9385 gnd.n5980 gnd.n5528 585
R9386 gnd.n5963 gnd.n5962 585
R9387 gnd.n5964 gnd.n5963 585
R9388 gnd.n5538 gnd.n5537 585
R9389 gnd.n5544 gnd.n5537 585
R9390 gnd.n5956 gnd.n5955 585
R9391 gnd.n5955 gnd.n5954 585
R9392 gnd.n5541 gnd.n5540 585
R9393 gnd.n5552 gnd.n5541 585
R9394 gnd.n5841 gnd.n5560 585
R9395 gnd.n5933 gnd.n5560 585
R9396 gnd.n5843 gnd.n5842 585
R9397 gnd.n5842 gnd.n5558 585
R9398 gnd.n5844 gnd.n5571 585
R9399 gnd.n5923 gnd.n5571 585
R9400 gnd.n5846 gnd.n5845 585
R9401 gnd.n5846 gnd.n5578 585
R9402 gnd.n5848 gnd.n5847 585
R9403 gnd.n5847 gnd.n5577 585
R9404 gnd.n5849 gnd.n5588 585
R9405 gnd.n5903 gnd.n5588 585
R9406 gnd.n5851 gnd.n5850 585
R9407 gnd.n5850 gnd.n5586 585
R9408 gnd.n5852 gnd.n5597 585
R9409 gnd.n5892 gnd.n5597 585
R9410 gnd.n5854 gnd.n5853 585
R9411 gnd.n5854 gnd.n5603 585
R9412 gnd.n5856 gnd.n5855 585
R9413 gnd.n5855 gnd.n5602 585
R9414 gnd.n5857 gnd.n5618 585
R9415 gnd.n5871 gnd.n5618 585
R9416 gnd.n5858 gnd.n5671 585
R9417 gnd.n5671 gnd.n5610 585
R9418 gnd.n5860 gnd.n5859 585
R9419 gnd.n5861 gnd.n5860 585
R9420 gnd.n5672 gnd.n5670 585
R9421 gnd.n5670 gnd.n5669 585
R9422 gnd.n5825 gnd.n5824 585
R9423 gnd.n5824 gnd.n5823 585
R9424 gnd.n5675 gnd.n5674 585
R9425 gnd.n5676 gnd.n5675 585
R9426 gnd.n5814 gnd.n5813 585
R9427 gnd.n5815 gnd.n5814 585
R9428 gnd.n5684 gnd.n5683 585
R9429 gnd.n5683 gnd.n5682 585
R9430 gnd.n5809 gnd.n5808 585
R9431 gnd.n5808 gnd.n5807 585
R9432 gnd.n5687 gnd.n5686 585
R9433 gnd.n5798 gnd.n5687 585
R9434 gnd.n5797 gnd.n5796 585
R9435 gnd.n5799 gnd.n5797 585
R9436 gnd.n5695 gnd.n5694 585
R9437 gnd.n5694 gnd.n5693 585
R9438 gnd.n7809 gnd.n7808 585
R9439 gnd.n7808 gnd.n7807 585
R9440 gnd.n7810 gnd.n207 585
R9441 gnd.n7656 gnd.n207 585
R9442 gnd.n7812 gnd.n7811 585
R9443 gnd.n7813 gnd.n7812 585
R9444 gnd.n192 gnd.n191 585
R9445 gnd.n7649 gnd.n192 585
R9446 gnd.n7821 gnd.n7820 585
R9447 gnd.n7820 gnd.n7819 585
R9448 gnd.n7822 gnd.n187 585
R9449 gnd.n7640 gnd.n187 585
R9450 gnd.n7824 gnd.n7823 585
R9451 gnd.n7825 gnd.n7824 585
R9452 gnd.n171 gnd.n170 585
R9453 gnd.n7634 gnd.n171 585
R9454 gnd.n7833 gnd.n7832 585
R9455 gnd.n7832 gnd.n7831 585
R9456 gnd.n7834 gnd.n166 585
R9457 gnd.n7626 gnd.n166 585
R9458 gnd.n7836 gnd.n7835 585
R9459 gnd.n7837 gnd.n7836 585
R9460 gnd.n152 gnd.n151 585
R9461 gnd.n7620 gnd.n152 585
R9462 gnd.n7845 gnd.n7844 585
R9463 gnd.n7844 gnd.n7843 585
R9464 gnd.n7846 gnd.n147 585
R9465 gnd.n7612 gnd.n147 585
R9466 gnd.n7848 gnd.n7847 585
R9467 gnd.n7849 gnd.n7848 585
R9468 gnd.n131 gnd.n130 585
R9469 gnd.n7606 gnd.n131 585
R9470 gnd.n7857 gnd.n7856 585
R9471 gnd.n7856 gnd.n7855 585
R9472 gnd.n7858 gnd.n126 585
R9473 gnd.n7598 gnd.n126 585
R9474 gnd.n7860 gnd.n7859 585
R9475 gnd.n7861 gnd.n7860 585
R9476 gnd.n113 gnd.n112 585
R9477 gnd.n7592 gnd.n113 585
R9478 gnd.n7869 gnd.n7868 585
R9479 gnd.n7868 gnd.n7867 585
R9480 gnd.n7870 gnd.n107 585
R9481 gnd.n7584 gnd.n107 585
R9482 gnd.n7872 gnd.n7871 585
R9483 gnd.n7873 gnd.n7872 585
R9484 gnd.n108 gnd.n106 585
R9485 gnd.n7578 gnd.n106 585
R9486 gnd.n4595 gnd.n4594 585
R9487 gnd.n4594 gnd.n391 585
R9488 gnd.n4596 gnd.n88 585
R9489 gnd.n7881 gnd.n88 585
R9490 gnd.n4598 gnd.n4597 585
R9491 gnd.n4599 gnd.n4598 585
R9492 gnd.n4589 gnd.n4588 585
R9493 gnd.n4588 gnd.n1857 585
R9494 gnd.n1845 gnd.n1844 585
R9495 gnd.n4635 gnd.n1845 585
R9496 gnd.n4640 gnd.n4639 585
R9497 gnd.n4639 gnd.n4638 585
R9498 gnd.n4641 gnd.n1840 585
R9499 gnd.n4620 gnd.n1840 585
R9500 gnd.n4643 gnd.n4642 585
R9501 gnd.n4644 gnd.n4643 585
R9502 gnd.n1828 gnd.n1827 585
R9503 gnd.n4609 gnd.n1828 585
R9504 gnd.n4652 gnd.n4651 585
R9505 gnd.n4651 gnd.n4650 585
R9506 gnd.n4653 gnd.n1823 585
R9507 gnd.n4579 gnd.n1823 585
R9508 gnd.n4655 gnd.n4654 585
R9509 gnd.n4656 gnd.n4655 585
R9510 gnd.n1807 gnd.n1806 585
R9511 gnd.n4538 gnd.n1807 585
R9512 gnd.n4664 gnd.n4663 585
R9513 gnd.n4663 gnd.n4662 585
R9514 gnd.n4665 gnd.n1802 585
R9515 gnd.n4531 gnd.n1802 585
R9516 gnd.n4667 gnd.n4666 585
R9517 gnd.n4668 gnd.n4667 585
R9518 gnd.n1788 gnd.n1787 585
R9519 gnd.n4526 gnd.n1788 585
R9520 gnd.n4676 gnd.n4675 585
R9521 gnd.n4675 gnd.n4674 585
R9522 gnd.n4677 gnd.n1783 585
R9523 gnd.n4555 gnd.n1783 585
R9524 gnd.n4679 gnd.n4678 585
R9525 gnd.n4680 gnd.n4679 585
R9526 gnd.n1767 gnd.n1766 585
R9527 gnd.n4519 gnd.n1767 585
R9528 gnd.n4688 gnd.n4687 585
R9529 gnd.n4687 gnd.n4686 585
R9530 gnd.n4689 gnd.n1762 585
R9531 gnd.n4511 gnd.n1762 585
R9532 gnd.n4691 gnd.n4690 585
R9533 gnd.n4692 gnd.n4691 585
R9534 gnd.n1747 gnd.n1746 585
R9535 gnd.n4505 gnd.n1747 585
R9536 gnd.n4700 gnd.n4699 585
R9537 gnd.n4699 gnd.n4698 585
R9538 gnd.n4701 gnd.n1741 585
R9539 gnd.n4497 gnd.n1741 585
R9540 gnd.n4703 gnd.n4702 585
R9541 gnd.n4704 gnd.n4703 585
R9542 gnd.n1742 gnd.n1740 585
R9543 gnd.n3925 gnd.n1740 585
R9544 gnd.n4490 gnd.n1728 585
R9545 gnd.n4710 gnd.n1728 585
R9546 gnd.n4012 gnd.n4011 585
R9547 gnd.n3975 gnd.n3974 585
R9548 gnd.n4026 gnd.n4025 585
R9549 gnd.n4028 gnd.n3973 585
R9550 gnd.n4031 gnd.n4030 585
R9551 gnd.n3966 gnd.n3965 585
R9552 gnd.n4045 gnd.n4044 585
R9553 gnd.n4047 gnd.n3964 585
R9554 gnd.n4050 gnd.n4049 585
R9555 gnd.n3957 gnd.n3956 585
R9556 gnd.n4064 gnd.n4063 585
R9557 gnd.n4066 gnd.n3955 585
R9558 gnd.n4069 gnd.n4068 585
R9559 gnd.n3948 gnd.n3947 585
R9560 gnd.n4084 gnd.n4083 585
R9561 gnd.n4086 gnd.n3946 585
R9562 gnd.n4089 gnd.n4088 585
R9563 gnd.n4090 gnd.n3943 585
R9564 gnd.n3942 gnd.n3941 585
R9565 gnd.n3942 gnd.n1716 585
R9566 gnd.n353 gnd.n352 585
R9567 gnd.n7663 gnd.n348 585
R9568 gnd.n7665 gnd.n7664 585
R9569 gnd.n7667 gnd.n346 585
R9570 gnd.n7669 gnd.n7668 585
R9571 gnd.n7670 gnd.n341 585
R9572 gnd.n7672 gnd.n7671 585
R9573 gnd.n7674 gnd.n339 585
R9574 gnd.n7676 gnd.n7675 585
R9575 gnd.n7677 gnd.n334 585
R9576 gnd.n7679 gnd.n7678 585
R9577 gnd.n7681 gnd.n332 585
R9578 gnd.n7683 gnd.n7682 585
R9579 gnd.n7684 gnd.n327 585
R9580 gnd.n7686 gnd.n7685 585
R9581 gnd.n7688 gnd.n325 585
R9582 gnd.n7690 gnd.n7689 585
R9583 gnd.n7691 gnd.n323 585
R9584 gnd.n7692 gnd.n211 585
R9585 gnd.n223 gnd.n211 585
R9586 gnd.n7659 gnd.n214 585
R9587 gnd.n7807 gnd.n214 585
R9588 gnd.n7658 gnd.n7657 585
R9589 gnd.n7657 gnd.n7656 585
R9590 gnd.n357 gnd.n206 585
R9591 gnd.n7813 gnd.n206 585
R9592 gnd.n7648 gnd.n7647 585
R9593 gnd.n7649 gnd.n7648 585
R9594 gnd.n361 gnd.n195 585
R9595 gnd.n7819 gnd.n195 585
R9596 gnd.n7642 gnd.n7641 585
R9597 gnd.n7641 gnd.n7640 585
R9598 gnd.n363 gnd.n185 585
R9599 gnd.n7825 gnd.n185 585
R9600 gnd.n7633 gnd.n7632 585
R9601 gnd.n7634 gnd.n7633 585
R9602 gnd.n366 gnd.n174 585
R9603 gnd.n7831 gnd.n174 585
R9604 gnd.n7628 gnd.n7627 585
R9605 gnd.n7627 gnd.n7626 585
R9606 gnd.n368 gnd.n165 585
R9607 gnd.n7837 gnd.n165 585
R9608 gnd.n7619 gnd.n7618 585
R9609 gnd.n7620 gnd.n7619 585
R9610 gnd.n373 gnd.n155 585
R9611 gnd.n7843 gnd.n155 585
R9612 gnd.n7614 gnd.n7613 585
R9613 gnd.n7613 gnd.n7612 585
R9614 gnd.n375 gnd.n145 585
R9615 gnd.n7849 gnd.n145 585
R9616 gnd.n7605 gnd.n7604 585
R9617 gnd.n7606 gnd.n7605 585
R9618 gnd.n378 gnd.n134 585
R9619 gnd.n7855 gnd.n134 585
R9620 gnd.n7600 gnd.n7599 585
R9621 gnd.n7599 gnd.n7598 585
R9622 gnd.n380 gnd.n125 585
R9623 gnd.n7861 gnd.n125 585
R9624 gnd.n7591 gnd.n7590 585
R9625 gnd.n7592 gnd.n7591 585
R9626 gnd.n385 gnd.n116 585
R9627 gnd.n7867 gnd.n116 585
R9628 gnd.n7586 gnd.n7585 585
R9629 gnd.n7585 gnd.n7584 585
R9630 gnd.n387 gnd.n104 585
R9631 gnd.n7873 gnd.n104 585
R9632 gnd.n7577 gnd.n7576 585
R9633 gnd.n7578 gnd.n7577 585
R9634 gnd.n84 gnd.n83 585
R9635 gnd.n391 gnd.n84 585
R9636 gnd.n7883 gnd.n7882 585
R9637 gnd.n7882 gnd.n7881 585
R9638 gnd.n7884 gnd.n82 585
R9639 gnd.n4599 gnd.n82 585
R9640 gnd.n1856 gnd.n81 585
R9641 gnd.n1857 gnd.n1856 585
R9642 gnd.n4614 gnd.n1855 585
R9643 gnd.n4635 gnd.n1855 585
R9644 gnd.n1864 gnd.n1848 585
R9645 gnd.n4638 gnd.n1848 585
R9646 gnd.n4619 gnd.n4618 585
R9647 gnd.n4620 gnd.n4619 585
R9648 gnd.n1863 gnd.n1839 585
R9649 gnd.n4644 gnd.n1839 585
R9650 gnd.n4611 gnd.n4610 585
R9651 gnd.n4610 gnd.n4609 585
R9652 gnd.n1866 gnd.n1830 585
R9653 gnd.n4650 gnd.n1830 585
R9654 gnd.n4541 gnd.n1868 585
R9655 gnd.n4579 gnd.n1868 585
R9656 gnd.n4542 gnd.n1821 585
R9657 gnd.n4656 gnd.n1821 585
R9658 gnd.n4543 gnd.n4539 585
R9659 gnd.n4539 gnd.n4538 585
R9660 gnd.n1887 gnd.n1810 585
R9661 gnd.n4662 gnd.n1810 585
R9662 gnd.n4547 gnd.n1886 585
R9663 gnd.n4531 gnd.n1886 585
R9664 gnd.n4548 gnd.n1801 585
R9665 gnd.n4668 gnd.n1801 585
R9666 gnd.n4549 gnd.n1885 585
R9667 gnd.n4526 gnd.n1885 585
R9668 gnd.n1882 gnd.n1790 585
R9669 gnd.n4674 gnd.n1790 585
R9670 gnd.n4554 gnd.n4553 585
R9671 gnd.n4555 gnd.n4554 585
R9672 gnd.n1881 gnd.n1781 585
R9673 gnd.n4680 gnd.n1781 585
R9674 gnd.n4518 gnd.n4517 585
R9675 gnd.n4519 gnd.n4518 585
R9676 gnd.n1891 gnd.n1770 585
R9677 gnd.n4686 gnd.n1770 585
R9678 gnd.n4513 gnd.n4512 585
R9679 gnd.n4512 gnd.n4511 585
R9680 gnd.n1893 gnd.n1761 585
R9681 gnd.n4692 gnd.n1761 585
R9682 gnd.n4504 gnd.n4503 585
R9683 gnd.n4505 gnd.n4504 585
R9684 gnd.n1928 gnd.n1750 585
R9685 gnd.n4698 gnd.n1750 585
R9686 gnd.n4499 gnd.n4498 585
R9687 gnd.n4498 gnd.n4497 585
R9688 gnd.n1930 gnd.n1738 585
R9689 gnd.n4704 gnd.n1738 585
R9690 gnd.n3927 gnd.n3926 585
R9691 gnd.n3926 gnd.n3925 585
R9692 gnd.n3928 gnd.n1726 585
R9693 gnd.n4710 gnd.n1726 585
R9694 gnd.n6577 gnd.n6576 585
R9695 gnd.n6578 gnd.n6577 585
R9696 gnd.n5239 gnd.n5237 585
R9697 gnd.n5237 gnd.n1122 585
R9698 gnd.n1110 gnd.n1109 585
R9699 gnd.n1114 gnd.n1110 585
R9700 gnd.n6588 gnd.n6587 585
R9701 gnd.n6587 gnd.n6586 585
R9702 gnd.n6589 gnd.n1102 585
R9703 gnd.n6459 gnd.n1102 585
R9704 gnd.n6591 gnd.n6590 585
R9705 gnd.n6592 gnd.n6591 585
R9706 gnd.n1103 gnd.n1101 585
R9707 gnd.n1101 gnd.n1097 585
R9708 gnd.n1084 gnd.n1083 585
R9709 gnd.n1088 gnd.n1084 585
R9710 gnd.n6602 gnd.n6601 585
R9711 gnd.n6601 gnd.n6600 585
R9712 gnd.n6603 gnd.n1076 585
R9713 gnd.n6470 gnd.n1076 585
R9714 gnd.n6605 gnd.n6604 585
R9715 gnd.n6606 gnd.n6605 585
R9716 gnd.n1077 gnd.n1075 585
R9717 gnd.n1075 gnd.n1072 585
R9718 gnd.n1059 gnd.n1058 585
R9719 gnd.n1063 gnd.n1059 585
R9720 gnd.n6616 gnd.n6615 585
R9721 gnd.n6615 gnd.n6614 585
R9722 gnd.n6617 gnd.n1053 585
R9723 gnd.n6145 gnd.n1053 585
R9724 gnd.n6619 gnd.n6618 585
R9725 gnd.n6620 gnd.n6619 585
R9726 gnd.n1054 gnd.n1052 585
R9727 gnd.n1052 gnd.n1049 585
R9728 gnd.n6164 gnd.n6163 585
R9729 gnd.n6165 gnd.n6164 585
R9730 gnd.n5332 gnd.n5331 585
R9731 gnd.n5331 gnd.n1039 585
R9732 gnd.n6158 gnd.n6157 585
R9733 gnd.n6157 gnd.n6156 585
R9734 gnd.n5335 gnd.n5334 585
R9735 gnd.n5344 gnd.n5335 585
R9736 gnd.n6107 gnd.n5357 585
R9737 gnd.n5357 gnd.n5343 585
R9738 gnd.n6109 gnd.n6108 585
R9739 gnd.n6110 gnd.n6109 585
R9740 gnd.n5358 gnd.n5356 585
R9741 gnd.n5365 gnd.n5356 585
R9742 gnd.n6102 gnd.n6101 585
R9743 gnd.n6101 gnd.n6100 585
R9744 gnd.n5361 gnd.n5360 585
R9745 gnd.n6081 gnd.n5361 585
R9746 gnd.n6067 gnd.n5384 585
R9747 gnd.n5384 gnd.n5374 585
R9748 gnd.n6069 gnd.n6068 585
R9749 gnd.n6070 gnd.n6069 585
R9750 gnd.n5385 gnd.n5383 585
R9751 gnd.n6058 gnd.n5383 585
R9752 gnd.n6062 gnd.n6061 585
R9753 gnd.n6061 gnd.n6060 585
R9754 gnd.n5388 gnd.n5387 585
R9755 gnd.n6013 gnd.n5388 585
R9756 gnd.n5506 gnd.n5505 585
R9757 gnd.n5507 gnd.n5506 585
R9758 gnd.n5486 gnd.n5485 585
R9759 gnd.n5489 gnd.n5486 585
R9760 gnd.n6023 gnd.n6022 585
R9761 gnd.n6022 gnd.n6021 585
R9762 gnd.n6024 gnd.n5480 585
R9763 gnd.n5516 gnd.n5480 585
R9764 gnd.n6026 gnd.n6025 585
R9765 gnd.n6027 gnd.n6026 585
R9766 gnd.n5481 gnd.n5479 585
R9767 gnd.n5991 gnd.n5479 585
R9768 gnd.n5975 gnd.n5974 585
R9769 gnd.n5974 gnd.n5467 585
R9770 gnd.n5976 gnd.n5531 585
R9771 gnd.n5531 gnd.n5466 585
R9772 gnd.n5978 gnd.n5977 585
R9773 gnd.n5979 gnd.n5978 585
R9774 gnd.n5532 gnd.n5530 585
R9775 gnd.n5530 gnd.n5527 585
R9776 gnd.n5967 gnd.n5966 585
R9777 gnd.n5966 gnd.n5965 585
R9778 gnd.n5535 gnd.n5534 585
R9779 gnd.n5542 gnd.n5535 585
R9780 gnd.n5941 gnd.n5940 585
R9781 gnd.n5942 gnd.n5941 585
R9782 gnd.n5554 gnd.n5553 585
R9783 gnd.n5561 gnd.n5553 585
R9784 gnd.n5936 gnd.n5935 585
R9785 gnd.n5935 gnd.n5934 585
R9786 gnd.n5557 gnd.n5556 585
R9787 gnd.n5924 gnd.n5557 585
R9788 gnd.n5911 gnd.n5581 585
R9789 gnd.n5581 gnd.n5580 585
R9790 gnd.n5913 gnd.n5912 585
R9791 gnd.n5914 gnd.n5913 585
R9792 gnd.n5582 gnd.n5579 585
R9793 gnd.n5589 gnd.n5579 585
R9794 gnd.n5906 gnd.n5905 585
R9795 gnd.n5905 gnd.n5904 585
R9796 gnd.n5585 gnd.n5584 585
R9797 gnd.n5893 gnd.n5585 585
R9798 gnd.n5880 gnd.n5606 585
R9799 gnd.n5606 gnd.n5605 585
R9800 gnd.n5882 gnd.n5881 585
R9801 gnd.n5883 gnd.n5882 585
R9802 gnd.n5876 gnd.n5604 585
R9803 gnd.n5875 gnd.n5874 585
R9804 gnd.n5609 gnd.n5608 585
R9805 gnd.n5872 gnd.n5609 585
R9806 gnd.n5631 gnd.n5630 585
R9807 gnd.n5634 gnd.n5633 585
R9808 gnd.n5632 gnd.n5627 585
R9809 gnd.n5639 gnd.n5638 585
R9810 gnd.n5641 gnd.n5640 585
R9811 gnd.n5644 gnd.n5643 585
R9812 gnd.n5642 gnd.n5625 585
R9813 gnd.n5649 gnd.n5648 585
R9814 gnd.n5651 gnd.n5650 585
R9815 gnd.n5654 gnd.n5653 585
R9816 gnd.n5652 gnd.n5623 585
R9817 gnd.n5659 gnd.n5658 585
R9818 gnd.n5663 gnd.n5660 585
R9819 gnd.n5664 gnd.n5601 585
R9820 gnd.n6546 gnd.n6545 585
R9821 gnd.n6548 gnd.n5268 585
R9822 gnd.n6550 gnd.n6549 585
R9823 gnd.n6551 gnd.n5261 585
R9824 gnd.n6553 gnd.n6552 585
R9825 gnd.n6555 gnd.n5259 585
R9826 gnd.n6557 gnd.n6556 585
R9827 gnd.n6558 gnd.n5254 585
R9828 gnd.n6560 gnd.n6559 585
R9829 gnd.n6562 gnd.n5252 585
R9830 gnd.n6564 gnd.n6563 585
R9831 gnd.n6565 gnd.n5247 585
R9832 gnd.n6567 gnd.n6566 585
R9833 gnd.n6569 gnd.n5245 585
R9834 gnd.n6571 gnd.n6570 585
R9835 gnd.n6572 gnd.n5243 585
R9836 gnd.n6573 gnd.n5238 585
R9837 gnd.n5238 gnd.n5236 585
R9838 gnd.n6453 gnd.n1124 585
R9839 gnd.n6578 gnd.n1124 585
R9840 gnd.n6455 gnd.n6454 585
R9841 gnd.n6455 gnd.n1122 585
R9842 gnd.n6457 gnd.n6456 585
R9843 gnd.n6456 gnd.n1114 585
R9844 gnd.n6458 gnd.n1112 585
R9845 gnd.n6586 gnd.n1112 585
R9846 gnd.n6461 gnd.n6460 585
R9847 gnd.n6460 gnd.n6459 585
R9848 gnd.n6462 gnd.n1099 585
R9849 gnd.n6592 gnd.n1099 585
R9850 gnd.n6464 gnd.n6463 585
R9851 gnd.n6464 gnd.n1097 585
R9852 gnd.n6466 gnd.n6465 585
R9853 gnd.n6465 gnd.n1088 585
R9854 gnd.n6467 gnd.n1086 585
R9855 gnd.n6600 gnd.n1086 585
R9856 gnd.n6469 gnd.n6468 585
R9857 gnd.n6470 gnd.n6469 585
R9858 gnd.n6182 gnd.n1074 585
R9859 gnd.n6606 gnd.n1074 585
R9860 gnd.n6181 gnd.n6180 585
R9861 gnd.n6180 gnd.n1072 585
R9862 gnd.n6179 gnd.n6177 585
R9863 gnd.n6179 gnd.n1063 585
R9864 gnd.n6175 gnd.n1061 585
R9865 gnd.n6614 gnd.n1061 585
R9866 gnd.n6144 gnd.n5325 585
R9867 gnd.n6145 gnd.n6144 585
R9868 gnd.n6169 gnd.n1051 585
R9869 gnd.n6620 gnd.n1051 585
R9870 gnd.n6168 gnd.n6167 585
R9871 gnd.n6167 gnd.n1049 585
R9872 gnd.n6166 gnd.n5327 585
R9873 gnd.n6166 gnd.n6165 585
R9874 gnd.n6116 gnd.n5329 585
R9875 gnd.n5329 gnd.n1039 585
R9876 gnd.n6117 gnd.n5337 585
R9877 gnd.n6156 gnd.n5337 585
R9878 gnd.n6114 gnd.n6113 585
R9879 gnd.n6113 gnd.n5344 585
R9880 gnd.n6112 gnd.n5351 585
R9881 gnd.n6112 gnd.n5343 585
R9882 gnd.n6111 gnd.n5353 585
R9883 gnd.n6111 gnd.n6110 585
R9884 gnd.n6090 gnd.n5352 585
R9885 gnd.n5365 gnd.n5352 585
R9886 gnd.n6089 gnd.n5363 585
R9887 gnd.n6100 gnd.n5363 585
R9888 gnd.n6080 gnd.n5370 585
R9889 gnd.n6081 gnd.n6080 585
R9890 gnd.n6079 gnd.n6078 585
R9891 gnd.n6079 gnd.n5374 585
R9892 gnd.n6077 gnd.n5376 585
R9893 gnd.n6070 gnd.n5376 585
R9894 gnd.n6057 gnd.n5377 585
R9895 gnd.n6058 gnd.n6057 585
R9896 gnd.n6010 gnd.n5390 585
R9897 gnd.n6060 gnd.n5390 585
R9898 gnd.n6012 gnd.n6011 585
R9899 gnd.n6013 gnd.n6012 585
R9900 gnd.n6005 gnd.n5508 585
R9901 gnd.n5508 gnd.n5507 585
R9902 gnd.n6003 gnd.n6002 585
R9903 gnd.n6002 gnd.n5489 585
R9904 gnd.n6000 gnd.n5487 585
R9905 gnd.n6021 gnd.n5487 585
R9906 gnd.n5518 gnd.n5517 585
R9907 gnd.n5517 gnd.n5516 585
R9908 gnd.n5994 gnd.n5477 585
R9909 gnd.n6027 gnd.n5477 585
R9910 gnd.n5993 gnd.n5992 585
R9911 gnd.n5992 gnd.n5991 585
R9912 gnd.n5989 gnd.n5520 585
R9913 gnd.n5989 gnd.n5467 585
R9914 gnd.n5988 gnd.n5987 585
R9915 gnd.n5988 gnd.n5466 585
R9916 gnd.n5523 gnd.n5522 585
R9917 gnd.n5979 gnd.n5522 585
R9918 gnd.n5947 gnd.n5946 585
R9919 gnd.n5946 gnd.n5527 585
R9920 gnd.n5948 gnd.n5536 585
R9921 gnd.n5965 gnd.n5536 585
R9922 gnd.n5945 gnd.n5944 585
R9923 gnd.n5944 gnd.n5542 585
R9924 gnd.n5943 gnd.n5550 585
R9925 gnd.n5943 gnd.n5942 585
R9926 gnd.n5928 gnd.n5551 585
R9927 gnd.n5561 gnd.n5551 585
R9928 gnd.n5927 gnd.n5559 585
R9929 gnd.n5934 gnd.n5559 585
R9930 gnd.n5926 gnd.n5925 585
R9931 gnd.n5925 gnd.n5924 585
R9932 gnd.n5570 gnd.n5567 585
R9933 gnd.n5580 gnd.n5570 585
R9934 gnd.n5916 gnd.n5915 585
R9935 gnd.n5915 gnd.n5914 585
R9936 gnd.n5576 gnd.n5575 585
R9937 gnd.n5589 gnd.n5576 585
R9938 gnd.n5896 gnd.n5587 585
R9939 gnd.n5904 gnd.n5587 585
R9940 gnd.n5895 gnd.n5894 585
R9941 gnd.n5894 gnd.n5893 585
R9942 gnd.n5596 gnd.n5594 585
R9943 gnd.n5605 gnd.n5596 585
R9944 gnd.n5885 gnd.n5884 585
R9945 gnd.n5884 gnd.n5883 585
R9946 gnd.n4241 gnd.n4240 585
R9947 gnd.n4242 gnd.n4241 585
R9948 gnd.n4155 gnd.n2010 585
R9949 gnd.n2017 gnd.n2010 585
R9950 gnd.n4154 gnd.n4153 585
R9951 gnd.n4153 gnd.n4152 585
R9952 gnd.n2013 gnd.n2012 585
R9953 gnd.t60 gnd.n2013 585
R9954 gnd.n3889 gnd.n2078 585
R9955 gnd.n2078 gnd.n2077 585
R9956 gnd.n3891 gnd.n3890 585
R9957 gnd.n3892 gnd.n3891 585
R9958 gnd.n3888 gnd.n2076 585
R9959 gnd.n2084 gnd.n2076 585
R9960 gnd.n3887 gnd.n3886 585
R9961 gnd.n3886 gnd.n3885 585
R9962 gnd.n2080 gnd.n2079 585
R9963 gnd.n3752 gnd.n2080 585
R9964 gnd.n3867 gnd.n3866 585
R9965 gnd.n3868 gnd.n3867 585
R9966 gnd.n3865 gnd.n2096 585
R9967 gnd.n2096 gnd.n2092 585
R9968 gnd.n3864 gnd.n3863 585
R9969 gnd.n3863 gnd.n3862 585
R9970 gnd.n2098 gnd.n2097 585
R9971 gnd.n3760 gnd.n2098 585
R9972 gnd.n3842 gnd.n3841 585
R9973 gnd.n3843 gnd.n3842 585
R9974 gnd.n3840 gnd.n2110 585
R9975 gnd.n2110 gnd.n2107 585
R9976 gnd.n3839 gnd.n3838 585
R9977 gnd.n3838 gnd.n3837 585
R9978 gnd.n2112 gnd.n2111 585
R9979 gnd.n3768 gnd.n2112 585
R9980 gnd.n3824 gnd.n3823 585
R9981 gnd.n3825 gnd.n3824 585
R9982 gnd.n3822 gnd.n2122 585
R9983 gnd.n3817 gnd.n2122 585
R9984 gnd.n3821 gnd.n3820 585
R9985 gnd.n3820 gnd.n3819 585
R9986 gnd.n2124 gnd.n2123 585
R9987 gnd.n3775 gnd.n2124 585
R9988 gnd.n3793 gnd.n3792 585
R9989 gnd.n3792 gnd.n2136 585
R9990 gnd.n3794 gnd.n2145 585
R9991 gnd.n3780 gnd.n2145 585
R9992 gnd.n3796 gnd.n3795 585
R9993 gnd.n3797 gnd.n3796 585
R9994 gnd.n3791 gnd.n2144 585
R9995 gnd.n3786 gnd.n2144 585
R9996 gnd.n3790 gnd.n3789 585
R9997 gnd.n3789 gnd.n3788 585
R9998 gnd.n2147 gnd.n2146 585
R9999 gnd.n3746 gnd.n2147 585
R10000 gnd.n3732 gnd.n2165 585
R10001 gnd.n2165 gnd.n2164 585
R10002 gnd.n3734 gnd.n3733 585
R10003 gnd.n3735 gnd.n3734 585
R10004 gnd.n3731 gnd.n2163 585
R10005 gnd.n2163 gnd.n2159 585
R10006 gnd.n3730 gnd.n3729 585
R10007 gnd.n3729 gnd.n3728 585
R10008 gnd.n2167 gnd.n2166 585
R10009 gnd.n3666 gnd.n2167 585
R10010 gnd.n3707 gnd.n3706 585
R10011 gnd.n3708 gnd.n3707 585
R10012 gnd.n3705 gnd.n2179 585
R10013 gnd.n2179 gnd.n2176 585
R10014 gnd.n3704 gnd.n3703 585
R10015 gnd.n3703 gnd.n3702 585
R10016 gnd.n2181 gnd.n2180 585
R10017 gnd.n3674 gnd.n2181 585
R10018 gnd.n3689 gnd.n3688 585
R10019 gnd.n3690 gnd.n3689 585
R10020 gnd.n3687 gnd.n2192 585
R10021 gnd.n3680 gnd.n2192 585
R10022 gnd.n3686 gnd.n3685 585
R10023 gnd.n3685 gnd.n3684 585
R10024 gnd.n2194 gnd.n2193 585
R10025 gnd.n3656 gnd.n2194 585
R10026 gnd.n3642 gnd.n3641 585
R10027 gnd.n3641 gnd.n2200 585
R10028 gnd.n3643 gnd.n2209 585
R10029 gnd.n3575 gnd.n2209 585
R10030 gnd.n3645 gnd.n3644 585
R10031 gnd.n3646 gnd.n3645 585
R10032 gnd.n3640 gnd.n2208 585
R10033 gnd.n3635 gnd.n2208 585
R10034 gnd.n3639 gnd.n3638 585
R10035 gnd.n3638 gnd.n3637 585
R10036 gnd.n2211 gnd.n2210 585
R10037 gnd.n2223 gnd.n2211 585
R10038 gnd.n3599 gnd.n3598 585
R10039 gnd.n3598 gnd.n2222 585
R10040 gnd.n3600 gnd.n2233 585
R10041 gnd.n3586 gnd.n2233 585
R10042 gnd.n3602 gnd.n3601 585
R10043 gnd.n3603 gnd.n3602 585
R10044 gnd.n3597 gnd.n2232 585
R10045 gnd.n3592 gnd.n2232 585
R10046 gnd.n3596 gnd.n3595 585
R10047 gnd.n3595 gnd.n3594 585
R10048 gnd.n2235 gnd.n2234 585
R10049 gnd.n3569 gnd.n2235 585
R10050 gnd.n3555 gnd.n2250 585
R10051 gnd.n3533 gnd.n2250 585
R10052 gnd.n3557 gnd.n3556 585
R10053 gnd.n3558 gnd.n3557 585
R10054 gnd.n3554 gnd.n2249 585
R10055 gnd.n3548 gnd.n2249 585
R10056 gnd.n3553 gnd.n3552 585
R10057 gnd.n3552 gnd.n3551 585
R10058 gnd.n2252 gnd.n2251 585
R10059 gnd.n3541 gnd.n2252 585
R10060 gnd.n3517 gnd.n2269 585
R10061 gnd.n2269 gnd.n2268 585
R10062 gnd.n3519 gnd.n3518 585
R10063 gnd.n3520 gnd.n3519 585
R10064 gnd.n3516 gnd.n2266 585
R10065 gnd.n2266 gnd.n2263 585
R10066 gnd.n3515 gnd.n3514 585
R10067 gnd.n3514 gnd.n3513 585
R10068 gnd.n2271 gnd.n2270 585
R10069 gnd.n3429 gnd.n2271 585
R10070 gnd.n3497 gnd.n3496 585
R10071 gnd.n3498 gnd.n3497 585
R10072 gnd.n3495 gnd.n2284 585
R10073 gnd.n3490 gnd.n2284 585
R10074 gnd.n3494 gnd.n3493 585
R10075 gnd.n3493 gnd.n3492 585
R10076 gnd.n2286 gnd.n2285 585
R10077 gnd.n3478 gnd.n2286 585
R10078 gnd.n3465 gnd.n2308 585
R10079 gnd.n2308 gnd.n2296 585
R10080 gnd.n3467 gnd.n3466 585
R10081 gnd.n3468 gnd.n3467 585
R10082 gnd.n3464 gnd.n2307 585
R10083 gnd.n2307 gnd.n2303 585
R10084 gnd.n3463 gnd.n3462 585
R10085 gnd.n3462 gnd.n3461 585
R10086 gnd.n2310 gnd.n2309 585
R10087 gnd.n3444 gnd.n2310 585
R10088 gnd.n3450 gnd.n3449 585
R10089 gnd.n3451 gnd.n3450 585
R10090 gnd.n3448 gnd.n3447 585
R10091 gnd.n3447 gnd.n2319 585
R10092 gnd.n1614 gnd.n1613 585
R10093 gnd.n3420 gnd.n1614 585
R10094 gnd.n4829 gnd.n4828 585
R10095 gnd.n4828 gnd.n4827 585
R10096 gnd.n4830 gnd.n1611 585
R10097 gnd.n3409 gnd.n1611 585
R10098 gnd.n4832 gnd.n4831 585
R10099 gnd.n4833 gnd.n4832 585
R10100 gnd.n1612 gnd.n1610 585
R10101 gnd.n3402 gnd.n1610 585
R10102 gnd.n1596 gnd.n1595 585
R10103 gnd.n3400 gnd.n1596 585
R10104 gnd.n4843 gnd.n4842 585
R10105 gnd.n4842 gnd.n4841 585
R10106 gnd.n4844 gnd.n1574 585
R10107 gnd.n3394 gnd.n1574 585
R10108 gnd.n4909 gnd.n4908 585
R10109 gnd.n4907 gnd.n1573 585
R10110 gnd.n4906 gnd.n1572 585
R10111 gnd.n4911 gnd.n1572 585
R10112 gnd.n4905 gnd.n4904 585
R10113 gnd.n4903 gnd.n4902 585
R10114 gnd.n4901 gnd.n4900 585
R10115 gnd.n4899 gnd.n4898 585
R10116 gnd.n4897 gnd.n4896 585
R10117 gnd.n4895 gnd.n4894 585
R10118 gnd.n4893 gnd.n4892 585
R10119 gnd.n4891 gnd.n4890 585
R10120 gnd.n4889 gnd.n4888 585
R10121 gnd.n4887 gnd.n4886 585
R10122 gnd.n4885 gnd.n4884 585
R10123 gnd.n4883 gnd.n4882 585
R10124 gnd.n4881 gnd.n4880 585
R10125 gnd.n4879 gnd.n4878 585
R10126 gnd.n4877 gnd.n4876 585
R10127 gnd.n4875 gnd.n4874 585
R10128 gnd.n4873 gnd.n4872 585
R10129 gnd.n4871 gnd.n4870 585
R10130 gnd.n4869 gnd.n4868 585
R10131 gnd.n4867 gnd.n4866 585
R10132 gnd.n4865 gnd.n4864 585
R10133 gnd.n4863 gnd.n4862 585
R10134 gnd.n4861 gnd.n4860 585
R10135 gnd.n4859 gnd.n4858 585
R10136 gnd.n4857 gnd.n4856 585
R10137 gnd.n4855 gnd.n4854 585
R10138 gnd.n4853 gnd.n4852 585
R10139 gnd.n4851 gnd.n4850 585
R10140 gnd.n4849 gnd.n1536 585
R10141 gnd.n4914 gnd.n4913 585
R10142 gnd.n1538 gnd.n1535 585
R10143 gnd.n3331 gnd.n3330 585
R10144 gnd.n3333 gnd.n3332 585
R10145 gnd.n3336 gnd.n3335 585
R10146 gnd.n3338 gnd.n3337 585
R10147 gnd.n3340 gnd.n3339 585
R10148 gnd.n3342 gnd.n3341 585
R10149 gnd.n3344 gnd.n3343 585
R10150 gnd.n3346 gnd.n3345 585
R10151 gnd.n3348 gnd.n3347 585
R10152 gnd.n3350 gnd.n3349 585
R10153 gnd.n3352 gnd.n3351 585
R10154 gnd.n3354 gnd.n3353 585
R10155 gnd.n3356 gnd.n3355 585
R10156 gnd.n3358 gnd.n3357 585
R10157 gnd.n3360 gnd.n3359 585
R10158 gnd.n3362 gnd.n3361 585
R10159 gnd.n3364 gnd.n3363 585
R10160 gnd.n3366 gnd.n3365 585
R10161 gnd.n3368 gnd.n3367 585
R10162 gnd.n3370 gnd.n3369 585
R10163 gnd.n3372 gnd.n3371 585
R10164 gnd.n3374 gnd.n3373 585
R10165 gnd.n3376 gnd.n3375 585
R10166 gnd.n3378 gnd.n3377 585
R10167 gnd.n3380 gnd.n3379 585
R10168 gnd.n3382 gnd.n3381 585
R10169 gnd.n3384 gnd.n3383 585
R10170 gnd.n3386 gnd.n3385 585
R10171 gnd.n3388 gnd.n3387 585
R10172 gnd.n3390 gnd.n3389 585
R10173 gnd.n3392 gnd.n3391 585
R10174 gnd.n4245 gnd.n4244 585
R10175 gnd.n4247 gnd.n4246 585
R10176 gnd.n4249 gnd.n4248 585
R10177 gnd.n4251 gnd.n4250 585
R10178 gnd.n4253 gnd.n4252 585
R10179 gnd.n4255 gnd.n4254 585
R10180 gnd.n4257 gnd.n4256 585
R10181 gnd.n4259 gnd.n4258 585
R10182 gnd.n4261 gnd.n4260 585
R10183 gnd.n4263 gnd.n4262 585
R10184 gnd.n4265 gnd.n4264 585
R10185 gnd.n4267 gnd.n4266 585
R10186 gnd.n4269 gnd.n4268 585
R10187 gnd.n4271 gnd.n4270 585
R10188 gnd.n4273 gnd.n4272 585
R10189 gnd.n4275 gnd.n4274 585
R10190 gnd.n4277 gnd.n4276 585
R10191 gnd.n4279 gnd.n4278 585
R10192 gnd.n4281 gnd.n4280 585
R10193 gnd.n4283 gnd.n4282 585
R10194 gnd.n4285 gnd.n4284 585
R10195 gnd.n4287 gnd.n4286 585
R10196 gnd.n4289 gnd.n4288 585
R10197 gnd.n4291 gnd.n4290 585
R10198 gnd.n4293 gnd.n4292 585
R10199 gnd.n4295 gnd.n4294 585
R10200 gnd.n4297 gnd.n4296 585
R10201 gnd.n4299 gnd.n4298 585
R10202 gnd.n4301 gnd.n4300 585
R10203 gnd.n4303 gnd.n2003 585
R10204 gnd.n4305 gnd.n4304 585
R10205 gnd.n4307 gnd.n1967 585
R10206 gnd.n4309 gnd.n4308 585
R10207 gnd.n4312 gnd.n4311 585
R10208 gnd.n1970 gnd.n1968 585
R10209 gnd.n4178 gnd.n4177 585
R10210 gnd.n4180 gnd.n4179 585
R10211 gnd.n4183 gnd.n4182 585
R10212 gnd.n4185 gnd.n4184 585
R10213 gnd.n4187 gnd.n4186 585
R10214 gnd.n4189 gnd.n4188 585
R10215 gnd.n4191 gnd.n4190 585
R10216 gnd.n4193 gnd.n4192 585
R10217 gnd.n4195 gnd.n4194 585
R10218 gnd.n4197 gnd.n4196 585
R10219 gnd.n4199 gnd.n4198 585
R10220 gnd.n4201 gnd.n4200 585
R10221 gnd.n4203 gnd.n4202 585
R10222 gnd.n4205 gnd.n4204 585
R10223 gnd.n4207 gnd.n4206 585
R10224 gnd.n4209 gnd.n4208 585
R10225 gnd.n4211 gnd.n4210 585
R10226 gnd.n4213 gnd.n4212 585
R10227 gnd.n4215 gnd.n4214 585
R10228 gnd.n4217 gnd.n4216 585
R10229 gnd.n4219 gnd.n4218 585
R10230 gnd.n4221 gnd.n4220 585
R10231 gnd.n4223 gnd.n4222 585
R10232 gnd.n4225 gnd.n4224 585
R10233 gnd.n4227 gnd.n4226 585
R10234 gnd.n4229 gnd.n4228 585
R10235 gnd.n4231 gnd.n4230 585
R10236 gnd.n4233 gnd.n4232 585
R10237 gnd.n4235 gnd.n4234 585
R10238 gnd.n4237 gnd.n4236 585
R10239 gnd.n4238 gnd.n2011 585
R10240 gnd.n4243 gnd.n2006 585
R10241 gnd.n4243 gnd.n4242 585
R10242 gnd.n3896 gnd.n2007 585
R10243 gnd.n2017 gnd.n2007 585
R10244 gnd.n3897 gnd.n2015 585
R10245 gnd.n4152 gnd.n2015 585
R10246 gnd.n3899 gnd.n3898 585
R10247 gnd.t60 gnd.n3899 585
R10248 gnd.n3895 gnd.n2072 585
R10249 gnd.n2077 gnd.n2072 585
R10250 gnd.n3894 gnd.n3893 585
R10251 gnd.n3893 gnd.n3892 585
R10252 gnd.n2074 gnd.n2073 585
R10253 gnd.n2084 gnd.n2074 585
R10254 gnd.n3751 gnd.n2083 585
R10255 gnd.n3885 gnd.n2083 585
R10256 gnd.n3754 gnd.n3753 585
R10257 gnd.n3753 gnd.n3752 585
R10258 gnd.n3755 gnd.n2094 585
R10259 gnd.n3868 gnd.n2094 585
R10260 gnd.n3757 gnd.n3756 585
R10261 gnd.n3756 gnd.n2092 585
R10262 gnd.n3758 gnd.n2100 585
R10263 gnd.n3862 gnd.n2100 585
R10264 gnd.n3762 gnd.n3761 585
R10265 gnd.n3761 gnd.n3760 585
R10266 gnd.n3763 gnd.n2108 585
R10267 gnd.n3843 gnd.n2108 585
R10268 gnd.n3765 gnd.n3764 585
R10269 gnd.n3764 gnd.n2107 585
R10270 gnd.n3766 gnd.n2113 585
R10271 gnd.n3837 gnd.n2113 585
R10272 gnd.n3770 gnd.n3769 585
R10273 gnd.n3769 gnd.n3768 585
R10274 gnd.n3771 gnd.n2120 585
R10275 gnd.n3825 gnd.n2120 585
R10276 gnd.n3772 gnd.n2128 585
R10277 gnd.n3817 gnd.n2128 585
R10278 gnd.n3773 gnd.n2127 585
R10279 gnd.n3819 gnd.n2127 585
R10280 gnd.n3776 gnd.n3774 585
R10281 gnd.n3776 gnd.n3775 585
R10282 gnd.n3777 gnd.n3750 585
R10283 gnd.n3777 gnd.n2136 585
R10284 gnd.n3782 gnd.n3781 585
R10285 gnd.n3781 gnd.n3780 585
R10286 gnd.n3783 gnd.n2143 585
R10287 gnd.n3797 gnd.n2143 585
R10288 gnd.n3785 gnd.n3784 585
R10289 gnd.n3786 gnd.n3785 585
R10290 gnd.n3749 gnd.n2150 585
R10291 gnd.n3788 gnd.n2150 585
R10292 gnd.n3748 gnd.n3747 585
R10293 gnd.n3747 gnd.n3746 585
R10294 gnd.n2152 gnd.n2151 585
R10295 gnd.n2164 gnd.n2152 585
R10296 gnd.n3660 gnd.n2161 585
R10297 gnd.n3735 gnd.n2161 585
R10298 gnd.n3662 gnd.n3661 585
R10299 gnd.n3661 gnd.n2159 585
R10300 gnd.n3663 gnd.n2169 585
R10301 gnd.n3728 gnd.n2169 585
R10302 gnd.n3668 gnd.n3667 585
R10303 gnd.n3667 gnd.n3666 585
R10304 gnd.n3669 gnd.n2177 585
R10305 gnd.n3708 gnd.n2177 585
R10306 gnd.n3671 gnd.n3670 585
R10307 gnd.n3670 gnd.n2176 585
R10308 gnd.n3672 gnd.n2183 585
R10309 gnd.n3702 gnd.n2183 585
R10310 gnd.n3676 gnd.n3675 585
R10311 gnd.n3675 gnd.n3674 585
R10312 gnd.n3677 gnd.n2190 585
R10313 gnd.n3690 gnd.n2190 585
R10314 gnd.n3679 gnd.n3678 585
R10315 gnd.n3680 gnd.n3679 585
R10316 gnd.n3659 gnd.n2196 585
R10317 gnd.n3684 gnd.n2196 585
R10318 gnd.n3658 gnd.n3657 585
R10319 gnd.n3657 gnd.n3656 585
R10320 gnd.n2199 gnd.n2198 585
R10321 gnd.n2200 gnd.n2199 585
R10322 gnd.n3577 gnd.n3576 585
R10323 gnd.n3576 gnd.n3575 585
R10324 gnd.n3578 gnd.n2206 585
R10325 gnd.n3646 gnd.n2206 585
R10326 gnd.n3579 gnd.n2214 585
R10327 gnd.n3635 gnd.n2214 585
R10328 gnd.n3580 gnd.n2213 585
R10329 gnd.n3637 gnd.n2213 585
R10330 gnd.n3582 gnd.n3581 585
R10331 gnd.n3582 gnd.n2223 585
R10332 gnd.n3583 gnd.n3573 585
R10333 gnd.n3583 gnd.n2222 585
R10334 gnd.n3588 gnd.n3587 585
R10335 gnd.n3587 gnd.n3586 585
R10336 gnd.n3589 gnd.n2231 585
R10337 gnd.n3603 gnd.n2231 585
R10338 gnd.n3591 gnd.n3590 585
R10339 gnd.n3592 gnd.n3591 585
R10340 gnd.n3572 gnd.n2236 585
R10341 gnd.n3594 gnd.n2236 585
R10342 gnd.n3571 gnd.n3570 585
R10343 gnd.n3570 gnd.n3569 585
R10344 gnd.n2238 gnd.n2237 585
R10345 gnd.n3533 gnd.n2238 585
R10346 gnd.n3545 gnd.n2248 585
R10347 gnd.n3558 gnd.n2248 585
R10348 gnd.n3547 gnd.n3546 585
R10349 gnd.n3548 gnd.n3547 585
R10350 gnd.n3544 gnd.n2253 585
R10351 gnd.n3551 gnd.n2253 585
R10352 gnd.n3543 gnd.n3542 585
R10353 gnd.n3542 gnd.n3541 585
R10354 gnd.n2255 gnd.n2254 585
R10355 gnd.n2268 gnd.n2255 585
R10356 gnd.n3425 gnd.n2264 585
R10357 gnd.n3520 gnd.n2264 585
R10358 gnd.n3427 gnd.n3426 585
R10359 gnd.n3426 gnd.n2263 585
R10360 gnd.n3428 gnd.n2274 585
R10361 gnd.n3513 gnd.n2274 585
R10362 gnd.n3431 gnd.n3430 585
R10363 gnd.n3430 gnd.n3429 585
R10364 gnd.n3432 gnd.n2282 585
R10365 gnd.n3498 gnd.n2282 585
R10366 gnd.n3433 gnd.n2289 585
R10367 gnd.n3490 gnd.n2289 585
R10368 gnd.n3434 gnd.n2288 585
R10369 gnd.n3492 gnd.n2288 585
R10370 gnd.n3435 gnd.n2297 585
R10371 gnd.n3478 gnd.n2297 585
R10372 gnd.n3437 gnd.n3436 585
R10373 gnd.n3436 gnd.n2296 585
R10374 gnd.n3438 gnd.n2304 585
R10375 gnd.n3468 gnd.n2304 585
R10376 gnd.n3440 gnd.n3439 585
R10377 gnd.n3439 gnd.n2303 585
R10378 gnd.n3441 gnd.n2312 585
R10379 gnd.n3461 gnd.n2312 585
R10380 gnd.n3443 gnd.n3442 585
R10381 gnd.n3444 gnd.n3443 585
R10382 gnd.n3424 gnd.n2320 585
R10383 gnd.n3451 gnd.n2320 585
R10384 gnd.n3423 gnd.n3422 585
R10385 gnd.n3422 gnd.n2319 585
R10386 gnd.n3421 gnd.n2322 585
R10387 gnd.n3421 gnd.n3420 585
R10388 gnd.n3406 gnd.n1616 585
R10389 gnd.n4827 gnd.n1616 585
R10390 gnd.n3408 gnd.n3407 585
R10391 gnd.n3409 gnd.n3408 585
R10392 gnd.n3405 gnd.n1609 585
R10393 gnd.n4833 gnd.n1609 585
R10394 gnd.n3404 gnd.n3403 585
R10395 gnd.n3403 gnd.n3402 585
R10396 gnd.n3399 gnd.n3398 585
R10397 gnd.n3400 gnd.n3399 585
R10398 gnd.n3397 gnd.n1598 585
R10399 gnd.n4841 gnd.n1598 585
R10400 gnd.n3396 gnd.n3395 585
R10401 gnd.n3395 gnd.n3394 585
R10402 gnd.n4965 gnd.n4964 585
R10403 gnd.n4966 gnd.n4965 585
R10404 gnd.n1469 gnd.n1468 585
R10405 gnd.n3140 gnd.n1469 585
R10406 gnd.n4974 gnd.n4973 585
R10407 gnd.n4973 gnd.n4972 585
R10408 gnd.n4975 gnd.n1463 585
R10409 gnd.n3133 gnd.n1463 585
R10410 gnd.n4977 gnd.n4976 585
R10411 gnd.n4978 gnd.n4977 585
R10412 gnd.n1449 gnd.n1448 585
R10413 gnd.n3124 gnd.n1449 585
R10414 gnd.n4986 gnd.n4985 585
R10415 gnd.n4985 gnd.n4984 585
R10416 gnd.n4987 gnd.n1443 585
R10417 gnd.n3118 gnd.n1443 585
R10418 gnd.n4989 gnd.n4988 585
R10419 gnd.n4990 gnd.n4989 585
R10420 gnd.n1428 gnd.n1427 585
R10421 gnd.n3049 gnd.n1428 585
R10422 gnd.n4998 gnd.n4997 585
R10423 gnd.n4997 gnd.n4996 585
R10424 gnd.n4999 gnd.n1422 585
R10425 gnd.n3043 gnd.n1422 585
R10426 gnd.n5001 gnd.n5000 585
R10427 gnd.n5002 gnd.n5001 585
R10428 gnd.n1409 gnd.n1408 585
R10429 gnd.n3037 gnd.n1409 585
R10430 gnd.n5010 gnd.n5009 585
R10431 gnd.n5009 gnd.n5008 585
R10432 gnd.n5011 gnd.n1403 585
R10433 gnd.n3066 gnd.n1403 585
R10434 gnd.n5013 gnd.n5012 585
R10435 gnd.n5014 gnd.n5013 585
R10436 gnd.n1388 gnd.n1387 585
R10437 gnd.n3030 gnd.n1388 585
R10438 gnd.n5022 gnd.n5021 585
R10439 gnd.n5021 gnd.n5020 585
R10440 gnd.n5023 gnd.n1383 585
R10441 gnd.n3022 gnd.n1383 585
R10442 gnd.n5025 gnd.n5024 585
R10443 gnd.n5026 gnd.n5025 585
R10444 gnd.n1368 gnd.n1366 585
R10445 gnd.n3015 gnd.n1368 585
R10446 gnd.n5034 gnd.n5033 585
R10447 gnd.n5033 gnd.n5032 585
R10448 gnd.n1367 gnd.n1365 585
R10449 gnd.n3007 gnd.n1367 585
R10450 gnd.n2977 gnd.n2976 585
R10451 gnd.n2978 gnd.n2977 585
R10452 gnd.n2975 gnd.n2974 585
R10453 gnd.n2974 gnd.n2654 585
R10454 gnd.n2973 gnd.n2659 585
R10455 gnd.n2973 gnd.n2972 585
R10456 gnd.n2658 gnd.n2657 585
R10457 gnd.n2959 gnd.n2657 585
R10458 gnd.n2943 gnd.n2683 585
R10459 gnd.n2943 gnd.n2942 585
R10460 gnd.n2944 gnd.n1364 585
R10461 gnd.n2945 gnd.n2944 585
R10462 gnd.n2682 gnd.n1358 585
R10463 gnd.n2934 gnd.n2682 585
R10464 gnd.n5037 gnd.n1355 585
R10465 gnd.n2690 gnd.n1355 585
R10466 gnd.n5039 gnd.n5038 585
R10467 gnd.n5040 gnd.n5039 585
R10468 gnd.n1340 gnd.n1339 585
R10469 gnd.n2883 gnd.n1340 585
R10470 gnd.n5048 gnd.n5047 585
R10471 gnd.n5047 gnd.n5046 585
R10472 gnd.n5049 gnd.n1334 585
R10473 gnd.n2889 gnd.n1334 585
R10474 gnd.n5051 gnd.n5050 585
R10475 gnd.n5052 gnd.n5051 585
R10476 gnd.n1320 gnd.n1319 585
R10477 gnd.n2895 gnd.n1320 585
R10478 gnd.n5060 gnd.n5059 585
R10479 gnd.n5059 gnd.n5058 585
R10480 gnd.n5061 gnd.n1314 585
R10481 gnd.n2901 gnd.n1314 585
R10482 gnd.n5063 gnd.n5062 585
R10483 gnd.n5064 gnd.n5063 585
R10484 gnd.n1299 gnd.n1298 585
R10485 gnd.n2862 gnd.n1299 585
R10486 gnd.n5072 gnd.n5071 585
R10487 gnd.n5071 gnd.n5070 585
R10488 gnd.n5073 gnd.n1293 585
R10489 gnd.n2853 gnd.n1293 585
R10490 gnd.n5075 gnd.n5074 585
R10491 gnd.n5076 gnd.n5075 585
R10492 gnd.n1279 gnd.n1278 585
R10493 gnd.n2846 gnd.n1279 585
R10494 gnd.n5084 gnd.n5083 585
R10495 gnd.n5083 gnd.n5082 585
R10496 gnd.n5085 gnd.n1273 585
R10497 gnd.n2838 gnd.n1273 585
R10498 gnd.n5087 gnd.n5086 585
R10499 gnd.n5088 gnd.n5087 585
R10500 gnd.n1257 gnd.n1256 585
R10501 gnd.n2788 gnd.n1257 585
R10502 gnd.n5096 gnd.n5095 585
R10503 gnd.n5095 gnd.n5094 585
R10504 gnd.n5097 gnd.n1250 585
R10505 gnd.n2780 gnd.n1250 585
R10506 gnd.n5099 gnd.n5098 585
R10507 gnd.n5100 gnd.n5099 585
R10508 gnd.n1251 gnd.n1172 585
R10509 gnd.n5103 gnd.n1172 585
R10510 gnd.n5224 gnd.n5223 585
R10511 gnd.n5222 gnd.n1171 585
R10512 gnd.n5221 gnd.n1170 585
R10513 gnd.n5226 gnd.n1170 585
R10514 gnd.n5220 gnd.n5219 585
R10515 gnd.n5218 gnd.n5217 585
R10516 gnd.n5216 gnd.n5215 585
R10517 gnd.n5214 gnd.n5213 585
R10518 gnd.n5212 gnd.n5211 585
R10519 gnd.n5210 gnd.n5209 585
R10520 gnd.n5208 gnd.n5207 585
R10521 gnd.n5206 gnd.n5205 585
R10522 gnd.n5204 gnd.n5203 585
R10523 gnd.n5202 gnd.n5201 585
R10524 gnd.n5200 gnd.n5199 585
R10525 gnd.n5198 gnd.n5197 585
R10526 gnd.n5196 gnd.n5195 585
R10527 gnd.n5194 gnd.n5193 585
R10528 gnd.n5192 gnd.n5191 585
R10529 gnd.n5189 gnd.n5188 585
R10530 gnd.n5187 gnd.n5186 585
R10531 gnd.n5185 gnd.n5184 585
R10532 gnd.n5183 gnd.n5182 585
R10533 gnd.n5181 gnd.n5180 585
R10534 gnd.n5179 gnd.n5178 585
R10535 gnd.n5177 gnd.n5176 585
R10536 gnd.n5175 gnd.n5174 585
R10537 gnd.n5173 gnd.n5172 585
R10538 gnd.n5171 gnd.n5170 585
R10539 gnd.n5169 gnd.n5168 585
R10540 gnd.n5167 gnd.n5166 585
R10541 gnd.n5165 gnd.n5164 585
R10542 gnd.n5163 gnd.n5162 585
R10543 gnd.n5161 gnd.n5160 585
R10544 gnd.n5159 gnd.n5158 585
R10545 gnd.n5157 gnd.n5156 585
R10546 gnd.n5155 gnd.n5154 585
R10547 gnd.n5153 gnd.n5152 585
R10548 gnd.n5151 gnd.n5150 585
R10549 gnd.n5149 gnd.n5148 585
R10550 gnd.n5147 gnd.n5146 585
R10551 gnd.n5145 gnd.n5144 585
R10552 gnd.n5143 gnd.n5142 585
R10553 gnd.n5141 gnd.n5140 585
R10554 gnd.n5139 gnd.n5138 585
R10555 gnd.n5137 gnd.n5136 585
R10556 gnd.n5135 gnd.n5134 585
R10557 gnd.n5133 gnd.n5132 585
R10558 gnd.n5131 gnd.n5130 585
R10559 gnd.n5129 gnd.n5128 585
R10560 gnd.n5127 gnd.n5126 585
R10561 gnd.n5125 gnd.n5124 585
R10562 gnd.n5123 gnd.n5122 585
R10563 gnd.n5121 gnd.n5120 585
R10564 gnd.n5119 gnd.n5118 585
R10565 gnd.n5117 gnd.n5116 585
R10566 gnd.n5115 gnd.n5114 585
R10567 gnd.n5113 gnd.n5112 585
R10568 gnd.n5111 gnd.n5110 585
R10569 gnd.n1241 gnd.n1234 585
R10570 gnd.n2530 gnd.n2529 585
R10571 gnd.n2527 gnd.n2423 585
R10572 gnd.n2526 gnd.n2525 585
R10573 gnd.n2519 gnd.n2425 585
R10574 gnd.n2521 gnd.n2520 585
R10575 gnd.n2517 gnd.n2427 585
R10576 gnd.n2516 gnd.n2515 585
R10577 gnd.n2509 gnd.n2429 585
R10578 gnd.n2511 gnd.n2510 585
R10579 gnd.n2507 gnd.n2431 585
R10580 gnd.n2506 gnd.n2505 585
R10581 gnd.n2499 gnd.n2433 585
R10582 gnd.n2501 gnd.n2500 585
R10583 gnd.n2497 gnd.n2435 585
R10584 gnd.n2496 gnd.n2495 585
R10585 gnd.n2489 gnd.n2437 585
R10586 gnd.n2491 gnd.n2490 585
R10587 gnd.n2487 gnd.n2439 585
R10588 gnd.n2486 gnd.n2485 585
R10589 gnd.n2479 gnd.n2441 585
R10590 gnd.n2481 gnd.n2480 585
R10591 gnd.n2477 gnd.n2445 585
R10592 gnd.n2476 gnd.n2475 585
R10593 gnd.n2469 gnd.n2447 585
R10594 gnd.n2471 gnd.n2470 585
R10595 gnd.n2467 gnd.n2449 585
R10596 gnd.n2466 gnd.n2465 585
R10597 gnd.n2459 gnd.n2451 585
R10598 gnd.n2461 gnd.n2460 585
R10599 gnd.n2457 gnd.n2454 585
R10600 gnd.n2456 gnd.n1531 585
R10601 gnd.n4916 gnd.n1527 585
R10602 gnd.n4918 gnd.n4917 585
R10603 gnd.n4920 gnd.n1525 585
R10604 gnd.n4922 gnd.n4921 585
R10605 gnd.n4923 gnd.n1520 585
R10606 gnd.n4925 gnd.n4924 585
R10607 gnd.n4927 gnd.n1518 585
R10608 gnd.n4929 gnd.n4928 585
R10609 gnd.n4931 gnd.n1511 585
R10610 gnd.n4933 gnd.n4932 585
R10611 gnd.n4935 gnd.n1509 585
R10612 gnd.n4937 gnd.n4936 585
R10613 gnd.n4938 gnd.n1504 585
R10614 gnd.n4940 gnd.n4939 585
R10615 gnd.n4942 gnd.n1502 585
R10616 gnd.n4944 gnd.n4943 585
R10617 gnd.n4945 gnd.n1497 585
R10618 gnd.n4947 gnd.n4946 585
R10619 gnd.n4949 gnd.n1495 585
R10620 gnd.n4951 gnd.n4950 585
R10621 gnd.n4952 gnd.n1489 585
R10622 gnd.n4954 gnd.n4953 585
R10623 gnd.n4956 gnd.n1488 585
R10624 gnd.n4957 gnd.n1486 585
R10625 gnd.n4960 gnd.n4959 585
R10626 gnd.n4961 gnd.n1483 585
R10627 gnd.n1487 gnd.n1483 585
R10628 gnd.n3137 gnd.n1480 585
R10629 gnd.n4966 gnd.n1480 585
R10630 gnd.n3139 gnd.n3138 585
R10631 gnd.n3140 gnd.n3139 585
R10632 gnd.n3136 gnd.n1471 585
R10633 gnd.n4972 gnd.n1471 585
R10634 gnd.n3135 gnd.n3134 585
R10635 gnd.n3134 gnd.n3133 585
R10636 gnd.n2610 gnd.n1460 585
R10637 gnd.n4978 gnd.n1460 585
R10638 gnd.n3123 gnd.n3122 585
R10639 gnd.n3124 gnd.n3123 585
R10640 gnd.n3121 gnd.n1450 585
R10641 gnd.n4984 gnd.n1450 585
R10642 gnd.n3120 gnd.n3119 585
R10643 gnd.n3119 gnd.n3118 585
R10644 gnd.n2615 gnd.n1440 585
R10645 gnd.n4990 gnd.n1440 585
R10646 gnd.n3048 gnd.n3047 585
R10647 gnd.n3049 gnd.n3048 585
R10648 gnd.n3046 gnd.n1430 585
R10649 gnd.n4996 gnd.n1430 585
R10650 gnd.n3045 gnd.n3044 585
R10651 gnd.n3044 gnd.n3043 585
R10652 gnd.n3040 gnd.n1420 585
R10653 gnd.n5002 gnd.n1420 585
R10654 gnd.n3039 gnd.n3038 585
R10655 gnd.n3038 gnd.n3037 585
R10656 gnd.n3036 gnd.n1410 585
R10657 gnd.n5008 gnd.n1410 585
R10658 gnd.n3035 gnd.n2629 585
R10659 gnd.n3066 gnd.n2629 585
R10660 gnd.n3033 gnd.n1400 585
R10661 gnd.n5014 gnd.n1400 585
R10662 gnd.n3032 gnd.n3031 585
R10663 gnd.n3031 gnd.n3030 585
R10664 gnd.n2638 gnd.n1390 585
R10665 gnd.n5020 gnd.n1390 585
R10666 gnd.n3021 gnd.n3020 585
R10667 gnd.n3022 gnd.n3021 585
R10668 gnd.n3018 gnd.n1381 585
R10669 gnd.n5026 gnd.n1381 585
R10670 gnd.n3017 gnd.n3016 585
R10671 gnd.n3016 gnd.n3015 585
R10672 gnd.n2643 gnd.n1369 585
R10673 gnd.n5032 gnd.n1369 585
R10674 gnd.n2965 gnd.n2649 585
R10675 gnd.n3007 gnd.n2649 585
R10676 gnd.n2966 gnd.n2655 585
R10677 gnd.n2978 gnd.n2655 585
R10678 gnd.n2964 gnd.n2963 585
R10679 gnd.n2963 gnd.n2654 585
R10680 gnd.n2962 gnd.n2661 585
R10681 gnd.n2972 gnd.n2661 585
R10682 gnd.n2961 gnd.n2960 585
R10683 gnd.n2960 gnd.n2959 585
R10684 gnd.n2672 gnd.n2670 585
R10685 gnd.n2942 gnd.n2672 585
R10686 gnd.n2937 gnd.n2679 585
R10687 gnd.n2945 gnd.n2679 585
R10688 gnd.n2936 gnd.n2935 585
R10689 gnd.n2935 gnd.n2934 585
R10690 gnd.n2689 gnd.n2688 585
R10691 gnd.n2690 gnd.n2689 585
R10692 gnd.n2880 gnd.n1352 585
R10693 gnd.n5040 gnd.n1352 585
R10694 gnd.n2882 gnd.n2881 585
R10695 gnd.n2883 gnd.n2882 585
R10696 gnd.n2870 gnd.n1342 585
R10697 gnd.n5046 gnd.n1342 585
R10698 gnd.n2891 gnd.n2890 585
R10699 gnd.n2890 gnd.n2889 585
R10700 gnd.n2892 gnd.n1331 585
R10701 gnd.n5052 gnd.n1331 585
R10702 gnd.n2894 gnd.n2893 585
R10703 gnd.n2895 gnd.n2894 585
R10704 gnd.n2868 gnd.n1321 585
R10705 gnd.n5058 gnd.n1321 585
R10706 gnd.n2867 gnd.n2701 585
R10707 gnd.n2901 gnd.n2701 585
R10708 gnd.n2865 gnd.n1311 585
R10709 gnd.n5064 gnd.n1311 585
R10710 gnd.n2864 gnd.n2863 585
R10711 gnd.n2863 gnd.n2862 585
R10712 gnd.n2707 gnd.n1301 585
R10713 gnd.n5070 gnd.n1301 585
R10714 gnd.n2852 gnd.n2851 585
R10715 gnd.n2853 gnd.n2852 585
R10716 gnd.n2849 gnd.n1290 585
R10717 gnd.n5076 gnd.n1290 585
R10718 gnd.n2848 gnd.n2847 585
R10719 gnd.n2847 gnd.n2846 585
R10720 gnd.n2711 gnd.n1280 585
R10721 gnd.n5082 gnd.n1280 585
R10722 gnd.n2794 gnd.n2793 585
R10723 gnd.n2838 gnd.n2794 585
R10724 gnd.n2791 gnd.n1270 585
R10725 gnd.n5088 gnd.n1270 585
R10726 gnd.n2790 gnd.n2789 585
R10727 gnd.n2789 gnd.n2788 585
R10728 gnd.n2715 gnd.n1259 585
R10729 gnd.n5094 gnd.n1259 585
R10730 gnd.n2779 gnd.n2778 585
R10731 gnd.n2780 gnd.n2779 585
R10732 gnd.n1242 gnd.n1240 585
R10733 gnd.n5100 gnd.n1242 585
R10734 gnd.n5105 gnd.n5104 585
R10735 gnd.n5104 gnd.n5103 585
R10736 gnd.n7806 gnd.n7805 585
R10737 gnd.n7807 gnd.n7806 585
R10738 gnd.n203 gnd.n202 585
R10739 gnd.n7656 gnd.n203 585
R10740 gnd.n7815 gnd.n7814 585
R10741 gnd.n7814 gnd.n7813 585
R10742 gnd.n7816 gnd.n197 585
R10743 gnd.n7649 gnd.n197 585
R10744 gnd.n7818 gnd.n7817 585
R10745 gnd.n7819 gnd.n7818 585
R10746 gnd.n182 gnd.n181 585
R10747 gnd.n7640 gnd.n182 585
R10748 gnd.n7827 gnd.n7826 585
R10749 gnd.n7826 gnd.n7825 585
R10750 gnd.n7828 gnd.n176 585
R10751 gnd.n7634 gnd.n176 585
R10752 gnd.n7830 gnd.n7829 585
R10753 gnd.n7831 gnd.n7830 585
R10754 gnd.n162 gnd.n161 585
R10755 gnd.n7626 gnd.n162 585
R10756 gnd.n7839 gnd.n7838 585
R10757 gnd.n7838 gnd.n7837 585
R10758 gnd.n7840 gnd.n156 585
R10759 gnd.n7620 gnd.n156 585
R10760 gnd.n7842 gnd.n7841 585
R10761 gnd.n7843 gnd.n7842 585
R10762 gnd.n142 gnd.n141 585
R10763 gnd.n7612 gnd.n142 585
R10764 gnd.n7851 gnd.n7850 585
R10765 gnd.n7850 gnd.n7849 585
R10766 gnd.n7852 gnd.n136 585
R10767 gnd.n7606 gnd.n136 585
R10768 gnd.n7854 gnd.n7853 585
R10769 gnd.n7855 gnd.n7854 585
R10770 gnd.n122 gnd.n121 585
R10771 gnd.n7598 gnd.n122 585
R10772 gnd.n7863 gnd.n7862 585
R10773 gnd.n7862 gnd.n7861 585
R10774 gnd.n7864 gnd.n117 585
R10775 gnd.n7592 gnd.n117 585
R10776 gnd.n7866 gnd.n7865 585
R10777 gnd.n7867 gnd.n7866 585
R10778 gnd.n101 gnd.n99 585
R10779 gnd.n7584 gnd.n101 585
R10780 gnd.n7875 gnd.n7874 585
R10781 gnd.n7874 gnd.n7873 585
R10782 gnd.n100 gnd.n92 585
R10783 gnd.n7578 gnd.n100 585
R10784 gnd.n7878 gnd.n90 585
R10785 gnd.n391 gnd.n90 585
R10786 gnd.n7880 gnd.n7879 585
R10787 gnd.n7881 gnd.n7880 585
R10788 gnd.n1850 gnd.n89 585
R10789 gnd.n4599 gnd.n89 585
R10790 gnd.n1852 gnd.n1851 585
R10791 gnd.n1857 gnd.n1852 585
R10792 gnd.n4636 gnd.n1853 585
R10793 gnd.n4636 gnd.n4635 585
R10794 gnd.n4637 gnd.n97 585
R10795 gnd.n4638 gnd.n4637 585
R10796 gnd.n1836 gnd.n1835 585
R10797 gnd.n4620 gnd.n1836 585
R10798 gnd.n4646 gnd.n4645 585
R10799 gnd.n4645 gnd.n4644 585
R10800 gnd.n4647 gnd.n1832 585
R10801 gnd.n4609 gnd.n1832 585
R10802 gnd.n4649 gnd.n4648 585
R10803 gnd.n4650 gnd.n4649 585
R10804 gnd.n1818 gnd.n1817 585
R10805 gnd.n4579 gnd.n1818 585
R10806 gnd.n4658 gnd.n4657 585
R10807 gnd.n4657 gnd.n4656 585
R10808 gnd.n4659 gnd.n1812 585
R10809 gnd.n4538 gnd.n1812 585
R10810 gnd.n4661 gnd.n4660 585
R10811 gnd.n4662 gnd.n4661 585
R10812 gnd.n1798 gnd.n1797 585
R10813 gnd.n4531 gnd.n1798 585
R10814 gnd.n4670 gnd.n4669 585
R10815 gnd.n4669 gnd.n4668 585
R10816 gnd.n4671 gnd.n1792 585
R10817 gnd.n4526 gnd.n1792 585
R10818 gnd.n4673 gnd.n4672 585
R10819 gnd.n4674 gnd.n4673 585
R10820 gnd.n1778 gnd.n1777 585
R10821 gnd.n4555 gnd.n1778 585
R10822 gnd.n4682 gnd.n4681 585
R10823 gnd.n4681 gnd.n4680 585
R10824 gnd.n4683 gnd.n1772 585
R10825 gnd.n4519 gnd.n1772 585
R10826 gnd.n4685 gnd.n4684 585
R10827 gnd.n4686 gnd.n4685 585
R10828 gnd.n1758 gnd.n1757 585
R10829 gnd.n4511 gnd.n1758 585
R10830 gnd.n4694 gnd.n4693 585
R10831 gnd.n4693 gnd.n4692 585
R10832 gnd.n4695 gnd.n1752 585
R10833 gnd.n4505 gnd.n1752 585
R10834 gnd.n4697 gnd.n4696 585
R10835 gnd.n4698 gnd.n4697 585
R10836 gnd.n1735 gnd.n1734 585
R10837 gnd.n4497 gnd.n1735 585
R10838 gnd.n4706 gnd.n4705 585
R10839 gnd.n4705 gnd.n4704 585
R10840 gnd.n4707 gnd.n1730 585
R10841 gnd.n3925 gnd.n1730 585
R10842 gnd.n4709 gnd.n4708 585
R10843 gnd.n4710 gnd.n4709 585
R10844 gnd.n4338 gnd.n1729 585
R10845 gnd.n4343 gnd.n4341 585
R10846 gnd.n4344 gnd.n4337 585
R10847 gnd.n4344 gnd.n1716 585
R10848 gnd.n4347 gnd.n4346 585
R10849 gnd.n4335 gnd.n4334 585
R10850 gnd.n4352 gnd.n4351 585
R10851 gnd.n4354 gnd.n4333 585
R10852 gnd.n4357 gnd.n4356 585
R10853 gnd.n4331 gnd.n4330 585
R10854 gnd.n4362 gnd.n4361 585
R10855 gnd.n4364 gnd.n4329 585
R10856 gnd.n4367 gnd.n4366 585
R10857 gnd.n4327 gnd.n4326 585
R10858 gnd.n4372 gnd.n4371 585
R10859 gnd.n4374 gnd.n4325 585
R10860 gnd.n4377 gnd.n4376 585
R10861 gnd.n4323 gnd.n4322 585
R10862 gnd.n4385 gnd.n4384 585
R10863 gnd.n4387 gnd.n4321 585
R10864 gnd.n4390 gnd.n4389 585
R10865 gnd.n4319 gnd.n4318 585
R10866 gnd.n4395 gnd.n4394 585
R10867 gnd.n4397 gnd.n4317 585
R10868 gnd.n4400 gnd.n4399 585
R10869 gnd.n4315 gnd.n4314 585
R10870 gnd.n4406 gnd.n4405 585
R10871 gnd.n4410 gnd.n1966 585
R10872 gnd.n4413 gnd.n4412 585
R10873 gnd.n1964 gnd.n1963 585
R10874 gnd.n4418 gnd.n4417 585
R10875 gnd.n4420 gnd.n1962 585
R10876 gnd.n4423 gnd.n4422 585
R10877 gnd.n1960 gnd.n1959 585
R10878 gnd.n4428 gnd.n4427 585
R10879 gnd.n4430 gnd.n1958 585
R10880 gnd.n4435 gnd.n4432 585
R10881 gnd.n1956 gnd.n1955 585
R10882 gnd.n4440 gnd.n4439 585
R10883 gnd.n4442 gnd.n1954 585
R10884 gnd.n4445 gnd.n4444 585
R10885 gnd.n1952 gnd.n1951 585
R10886 gnd.n4450 gnd.n4449 585
R10887 gnd.n4452 gnd.n1950 585
R10888 gnd.n4455 gnd.n4454 585
R10889 gnd.n1948 gnd.n1947 585
R10890 gnd.n4460 gnd.n4459 585
R10891 gnd.n4462 gnd.n1946 585
R10892 gnd.n4465 gnd.n4464 585
R10893 gnd.n1944 gnd.n1943 585
R10894 gnd.n4470 gnd.n4469 585
R10895 gnd.n4472 gnd.n1942 585
R10896 gnd.n4475 gnd.n4474 585
R10897 gnd.n1940 gnd.n1939 585
R10898 gnd.n4481 gnd.n4480 585
R10899 gnd.n4483 gnd.n1938 585
R10900 gnd.n4484 gnd.n1937 585
R10901 gnd.n4487 gnd.n4486 585
R10902 gnd.n7697 gnd.n7696 585
R10903 gnd.n7699 gnd.n319 585
R10904 gnd.n7701 gnd.n7700 585
R10905 gnd.n7702 gnd.n312 585
R10906 gnd.n7704 gnd.n7703 585
R10907 gnd.n7706 gnd.n310 585
R10908 gnd.n7708 gnd.n7707 585
R10909 gnd.n7709 gnd.n305 585
R10910 gnd.n7711 gnd.n7710 585
R10911 gnd.n7713 gnd.n303 585
R10912 gnd.n7715 gnd.n7714 585
R10913 gnd.n7716 gnd.n298 585
R10914 gnd.n7718 gnd.n7717 585
R10915 gnd.n7720 gnd.n296 585
R10916 gnd.n7722 gnd.n7721 585
R10917 gnd.n7723 gnd.n291 585
R10918 gnd.n7725 gnd.n7724 585
R10919 gnd.n7727 gnd.n290 585
R10920 gnd.n7728 gnd.n287 585
R10921 gnd.n7731 gnd.n7730 585
R10922 gnd.n289 gnd.n283 585
R10923 gnd.n7735 gnd.n280 585
R10924 gnd.n7737 gnd.n7736 585
R10925 gnd.n7739 gnd.n278 585
R10926 gnd.n7741 gnd.n7740 585
R10927 gnd.n7742 gnd.n273 585
R10928 gnd.n7744 gnd.n7743 585
R10929 gnd.n7746 gnd.n271 585
R10930 gnd.n7748 gnd.n7747 585
R10931 gnd.n7749 gnd.n266 585
R10932 gnd.n7751 gnd.n7750 585
R10933 gnd.n7753 gnd.n264 585
R10934 gnd.n7755 gnd.n7754 585
R10935 gnd.n7756 gnd.n259 585
R10936 gnd.n7758 gnd.n7757 585
R10937 gnd.n7760 gnd.n257 585
R10938 gnd.n7762 gnd.n7761 585
R10939 gnd.n7763 gnd.n252 585
R10940 gnd.n7765 gnd.n7764 585
R10941 gnd.n7767 gnd.n250 585
R10942 gnd.n7769 gnd.n7768 585
R10943 gnd.n7773 gnd.n245 585
R10944 gnd.n7775 gnd.n7774 585
R10945 gnd.n7777 gnd.n243 585
R10946 gnd.n7779 gnd.n7778 585
R10947 gnd.n7780 gnd.n238 585
R10948 gnd.n7782 gnd.n7781 585
R10949 gnd.n7784 gnd.n236 585
R10950 gnd.n7786 gnd.n7785 585
R10951 gnd.n7787 gnd.n231 585
R10952 gnd.n7789 gnd.n7788 585
R10953 gnd.n7791 gnd.n229 585
R10954 gnd.n7793 gnd.n7792 585
R10955 gnd.n7794 gnd.n224 585
R10956 gnd.n7796 gnd.n7795 585
R10957 gnd.n7798 gnd.n221 585
R10958 gnd.n7800 gnd.n7799 585
R10959 gnd.n7801 gnd.n219 585
R10960 gnd.n7802 gnd.n216 585
R10961 gnd.n223 gnd.n216 585
R10962 gnd.n7653 gnd.n213 585
R10963 gnd.n7807 gnd.n213 585
R10964 gnd.n7655 gnd.n7654 585
R10965 gnd.n7656 gnd.n7655 585
R10966 gnd.n7652 gnd.n205 585
R10967 gnd.n7813 gnd.n205 585
R10968 gnd.n7651 gnd.n7650 585
R10969 gnd.n7650 gnd.n7649 585
R10970 gnd.n359 gnd.n194 585
R10971 gnd.n7819 gnd.n194 585
R10972 gnd.n7639 gnd.n7638 585
R10973 gnd.n7640 gnd.n7639 585
R10974 gnd.n7637 gnd.n184 585
R10975 gnd.n7825 gnd.n184 585
R10976 gnd.n7636 gnd.n7635 585
R10977 gnd.n7635 gnd.n7634 585
R10978 gnd.n364 gnd.n173 585
R10979 gnd.n7831 gnd.n173 585
R10980 gnd.n7625 gnd.n7624 585
R10981 gnd.n7626 gnd.n7625 585
R10982 gnd.n7623 gnd.n164 585
R10983 gnd.n7837 gnd.n164 585
R10984 gnd.n7622 gnd.n7621 585
R10985 gnd.n7621 gnd.n7620 585
R10986 gnd.n370 gnd.n154 585
R10987 gnd.n7843 gnd.n154 585
R10988 gnd.n7611 gnd.n7610 585
R10989 gnd.n7612 gnd.n7611 585
R10990 gnd.n7609 gnd.n144 585
R10991 gnd.n7849 gnd.n144 585
R10992 gnd.n7608 gnd.n7607 585
R10993 gnd.n7607 gnd.n7606 585
R10994 gnd.n376 gnd.n133 585
R10995 gnd.n7855 gnd.n133 585
R10996 gnd.n7597 gnd.n7596 585
R10997 gnd.n7598 gnd.n7597 585
R10998 gnd.n7595 gnd.n124 585
R10999 gnd.n7861 gnd.n124 585
R11000 gnd.n7594 gnd.n7593 585
R11001 gnd.n7593 gnd.n7592 585
R11002 gnd.n382 gnd.n115 585
R11003 gnd.n7867 gnd.n115 585
R11004 gnd.n7583 gnd.n7582 585
R11005 gnd.n7584 gnd.n7583 585
R11006 gnd.n7581 gnd.n103 585
R11007 gnd.n7873 gnd.n103 585
R11008 gnd.n7580 gnd.n7579 585
R11009 gnd.n7579 gnd.n7578 585
R11010 gnd.n390 gnd.n388 585
R11011 gnd.n391 gnd.n390 585
R11012 gnd.n4591 gnd.n86 585
R11013 gnd.n7881 gnd.n86 585
R11014 gnd.n4600 gnd.n4586 585
R11015 gnd.n4600 gnd.n4599 585
R11016 gnd.n4602 gnd.n4601 585
R11017 gnd.n4601 gnd.n1857 585
R11018 gnd.n4603 gnd.n1854 585
R11019 gnd.n4635 gnd.n1854 585
R11020 gnd.n4604 gnd.n1847 585
R11021 gnd.n4638 gnd.n1847 585
R11022 gnd.n4605 gnd.n1862 585
R11023 gnd.n4620 gnd.n1862 585
R11024 gnd.n4606 gnd.n1838 585
R11025 gnd.n4644 gnd.n1838 585
R11026 gnd.n4608 gnd.n4607 585
R11027 gnd.n4609 gnd.n4608 585
R11028 gnd.n4582 gnd.n1829 585
R11029 gnd.n4650 gnd.n1829 585
R11030 gnd.n4581 gnd.n4580 585
R11031 gnd.n4580 gnd.n4579 585
R11032 gnd.n1867 gnd.n1820 585
R11033 gnd.n4656 gnd.n1820 585
R11034 gnd.n4537 gnd.n4536 585
R11035 gnd.n4538 gnd.n4537 585
R11036 gnd.n4534 gnd.n1809 585
R11037 gnd.n4662 gnd.n1809 585
R11038 gnd.n4533 gnd.n4532 585
R11039 gnd.n4532 gnd.n4531 585
R11040 gnd.n4529 gnd.n1800 585
R11041 gnd.n4668 gnd.n1800 585
R11042 gnd.n4528 gnd.n4527 585
R11043 gnd.n4527 gnd.n4526 585
R11044 gnd.n4524 gnd.n1789 585
R11045 gnd.n4674 gnd.n1789 585
R11046 gnd.n4523 gnd.n1880 585
R11047 gnd.n4555 gnd.n1880 585
R11048 gnd.n4522 gnd.n1780 585
R11049 gnd.n4680 gnd.n1780 585
R11050 gnd.n4521 gnd.n4520 585
R11051 gnd.n4520 gnd.n4519 585
R11052 gnd.n1889 gnd.n1769 585
R11053 gnd.n4686 gnd.n1769 585
R11054 gnd.n4510 gnd.n4509 585
R11055 gnd.n4511 gnd.n4510 585
R11056 gnd.n4508 gnd.n1760 585
R11057 gnd.n4692 gnd.n1760 585
R11058 gnd.n4507 gnd.n4506 585
R11059 gnd.n4506 gnd.n4505 585
R11060 gnd.n1926 gnd.n1749 585
R11061 gnd.n4698 gnd.n1749 585
R11062 gnd.n4496 gnd.n4495 585
R11063 gnd.n4497 gnd.n4496 585
R11064 gnd.n4494 gnd.n1737 585
R11065 gnd.n4704 gnd.n1737 585
R11066 gnd.n4493 gnd.n1932 585
R11067 gnd.n3925 gnd.n1932 585
R11068 gnd.n1931 gnd.n1725 585
R11069 gnd.n4710 gnd.n1725 585
R11070 gnd.n5234 gnd.n5233 585
R11071 gnd.n5235 gnd.n5234 585
R11072 gnd.n7525 gnd.n432 585
R11073 gnd.n7529 gnd.n432 585
R11074 gnd.n7532 gnd.n7531 585
R11075 gnd.n7531 gnd.n7530 585
R11076 gnd.n7533 gnd.n427 585
R11077 gnd.n433 gnd.n427 585
R11078 gnd.n7535 gnd.n7534 585
R11079 gnd.n7535 gnd.n215 585
R11080 gnd.n7536 gnd.n426 585
R11081 gnd.n7536 gnd.n212 585
R11082 gnd.n7538 gnd.n7537 585
R11083 gnd.n7537 gnd.n358 585
R11084 gnd.n7539 gnd.n421 585
R11085 gnd.n421 gnd.n204 585
R11086 gnd.n7541 gnd.n7540 585
R11087 gnd.n7541 gnd.n196 585
R11088 gnd.n7542 gnd.n420 585
R11089 gnd.n7542 gnd.n193 585
R11090 gnd.n7544 gnd.n7543 585
R11091 gnd.n7543 gnd.n186 585
R11092 gnd.n7545 gnd.n415 585
R11093 gnd.n415 gnd.n183 585
R11094 gnd.n7547 gnd.n7546 585
R11095 gnd.n7547 gnd.n175 585
R11096 gnd.n7548 gnd.n414 585
R11097 gnd.n7548 gnd.n172 585
R11098 gnd.n7550 gnd.n7549 585
R11099 gnd.n7549 gnd.n369 585
R11100 gnd.n7551 gnd.n409 585
R11101 gnd.n409 gnd.n163 585
R11102 gnd.n7553 gnd.n7552 585
R11103 gnd.n7553 gnd.n372 585
R11104 gnd.n7554 gnd.n408 585
R11105 gnd.n7554 gnd.n153 585
R11106 gnd.n7556 gnd.n7555 585
R11107 gnd.n7555 gnd.n146 585
R11108 gnd.n7557 gnd.n403 585
R11109 gnd.n403 gnd.n143 585
R11110 gnd.n7559 gnd.n7558 585
R11111 gnd.n7559 gnd.n135 585
R11112 gnd.n7560 gnd.n402 585
R11113 gnd.n7560 gnd.n132 585
R11114 gnd.n7562 gnd.n7561 585
R11115 gnd.n7561 gnd.n381 585
R11116 gnd.n7563 gnd.n397 585
R11117 gnd.n397 gnd.n123 585
R11118 gnd.n7565 gnd.n7564 585
R11119 gnd.n7565 gnd.n384 585
R11120 gnd.n7566 gnd.n396 585
R11121 gnd.n7566 gnd.n114 585
R11122 gnd.n7568 gnd.n7567 585
R11123 gnd.n7567 gnd.n105 585
R11124 gnd.n7569 gnd.n393 585
R11125 gnd.n393 gnd.n102 585
R11126 gnd.n7572 gnd.n7571 585
R11127 gnd.n7573 gnd.n7572 585
R11128 gnd.n394 gnd.n392 585
R11129 gnd.n392 gnd.n87 585
R11130 gnd.n4629 gnd.n4628 585
R11131 gnd.n4628 gnd.n85 585
R11132 gnd.n4630 gnd.n1859 585
R11133 gnd.n4587 gnd.n1859 585
R11134 gnd.n4633 gnd.n4632 585
R11135 gnd.n4634 gnd.n4633 585
R11136 gnd.n4626 gnd.n1858 585
R11137 gnd.n1858 gnd.n1849 585
R11138 gnd.n4624 gnd.n4623 585
R11139 gnd.n4623 gnd.n1846 585
R11140 gnd.n4622 gnd.n1860 585
R11141 gnd.n4622 gnd.n4621 585
R11142 gnd.n4574 gnd.n1861 585
R11143 gnd.n1861 gnd.n1837 585
R11144 gnd.n4575 gnd.n1870 585
R11145 gnd.n1870 gnd.n1831 585
R11146 gnd.n4577 gnd.n4576 585
R11147 gnd.n4578 gnd.n4577 585
R11148 gnd.n1871 gnd.n1869 585
R11149 gnd.n1869 gnd.n1822 585
R11150 gnd.n4568 gnd.n4567 585
R11151 gnd.n4567 gnd.n1819 585
R11152 gnd.n4566 gnd.n1873 585
R11153 gnd.n4566 gnd.n1811 585
R11154 gnd.n4565 gnd.n4564 585
R11155 gnd.n4565 gnd.n1808 585
R11156 gnd.n1875 gnd.n1874 585
R11157 gnd.n4530 gnd.n1874 585
R11158 gnd.n4560 gnd.n4559 585
R11159 gnd.n4559 gnd.n1799 585
R11160 gnd.n4558 gnd.n1877 585
R11161 gnd.n4558 gnd.n1791 585
R11162 gnd.n4557 gnd.n1879 585
R11163 gnd.n4557 gnd.n4556 585
R11164 gnd.n1917 gnd.n1878 585
R11165 gnd.n1878 gnd.n1782 585
R11166 gnd.n1919 gnd.n1918 585
R11167 gnd.n1919 gnd.n1779 585
R11168 gnd.n1921 gnd.n1920 585
R11169 gnd.n1920 gnd.n1771 585
R11170 gnd.n1922 gnd.n1895 585
R11171 gnd.n1895 gnd.n1768 585
R11172 gnd.n1924 gnd.n1923 585
R11173 gnd.n1925 gnd.n1924 585
R11174 gnd.n1896 gnd.n1894 585
R11175 gnd.n1894 gnd.n1759 585
R11176 gnd.n1908 gnd.n1907 585
R11177 gnd.n1907 gnd.n1751 585
R11178 gnd.n1906 gnd.n1898 585
R11179 gnd.n1906 gnd.n1748 585
R11180 gnd.n1905 gnd.n1904 585
R11181 gnd.n1905 gnd.n1739 585
R11182 gnd.n1900 gnd.n1899 585
R11183 gnd.n1899 gnd.n1736 585
R11184 gnd.n1723 gnd.n1722 585
R11185 gnd.n1727 gnd.n1723 585
R11186 gnd.n4713 gnd.n4712 585
R11187 gnd.n4712 gnd.n4711 585
R11188 gnd.n4714 gnd.n1717 585
R11189 gnd.n1724 gnd.n1717 585
R11190 gnd.n4716 gnd.n4715 585
R11191 gnd.n4717 gnd.n4716 585
R11192 gnd.n1714 gnd.n1713 585
R11193 gnd.n4718 gnd.n1714 585
R11194 gnd.n4721 gnd.n4720 585
R11195 gnd.n4720 gnd.n4719 585
R11196 gnd.n4722 gnd.n1708 585
R11197 gnd.n1708 gnd.n1706 585
R11198 gnd.n4724 gnd.n4723 585
R11199 gnd.n4725 gnd.n4724 585
R11200 gnd.n1709 gnd.n1707 585
R11201 gnd.n1707 gnd.n1704 585
R11202 gnd.n4113 gnd.n4108 585
R11203 gnd.n4108 gnd.n4107 585
R11204 gnd.n4115 gnd.n4114 585
R11205 gnd.n4116 gnd.n4115 585
R11206 gnd.n2046 gnd.n2045 585
R11207 gnd.n4119 gnd.n2046 585
R11208 gnd.n4123 gnd.n4122 585
R11209 gnd.n4122 gnd.n4121 585
R11210 gnd.n4124 gnd.n2040 585
R11211 gnd.n2056 gnd.n2040 585
R11212 gnd.n4126 gnd.n4125 585
R11213 gnd.n4127 gnd.n4126 585
R11214 gnd.n2035 gnd.n2034 585
R11215 gnd.n4130 gnd.n2035 585
R11216 gnd.n4134 gnd.n4133 585
R11217 gnd.n4133 gnd.n4132 585
R11218 gnd.n4135 gnd.n2029 585
R11219 gnd.n2036 gnd.n2029 585
R11220 gnd.n4137 gnd.n4136 585
R11221 gnd.n4138 gnd.n4137 585
R11222 gnd.n2025 gnd.n2024 585
R11223 gnd.n4141 gnd.n2025 585
R11224 gnd.n4145 gnd.n4144 585
R11225 gnd.n4144 gnd.n4143 585
R11226 gnd.n4146 gnd.n2019 585
R11227 gnd.n2019 gnd.n2009 585
R11228 gnd.n4148 gnd.n4147 585
R11229 gnd.n4149 gnd.n4148 585
R11230 gnd.n2020 gnd.n2018 585
R11231 gnd.n2018 gnd.n2014 585
R11232 gnd.n3880 gnd.n3879 585
R11233 gnd.n3879 gnd.n2071 585
R11234 gnd.n3881 gnd.n2087 585
R11235 gnd.n2087 gnd.t114 585
R11236 gnd.n3883 gnd.n3882 585
R11237 gnd.n3884 gnd.n3883 585
R11238 gnd.n2088 gnd.n2086 585
R11239 gnd.n2095 gnd.n2086 585
R11240 gnd.n3872 gnd.n3871 585
R11241 gnd.n3871 gnd.n3870 585
R11242 gnd.n2091 gnd.n2090 585
R11243 gnd.n2099 gnd.n2091 585
R11244 gnd.n3833 gnd.n2115 585
R11245 gnd.n2115 gnd.n2109 585
R11246 gnd.n3835 gnd.n3834 585
R11247 gnd.n3836 gnd.n3835 585
R11248 gnd.n2116 gnd.n2114 585
R11249 gnd.n3767 gnd.n2114 585
R11250 gnd.n3828 gnd.n3827 585
R11251 gnd.n3827 gnd.n3826 585
R11252 gnd.n2119 gnd.n2118 585
R11253 gnd.n3818 gnd.n2119 585
R11254 gnd.n3805 gnd.n3804 585
R11255 gnd.n3806 gnd.n3805 585
R11256 gnd.n2138 gnd.n2137 585
R11257 gnd.n3779 gnd.n2137 585
R11258 gnd.n3800 gnd.n3799 585
R11259 gnd.n3799 gnd.n3798 585
R11260 gnd.n2141 gnd.n2140 585
R11261 gnd.n3787 gnd.n2141 585
R11262 gnd.n3744 gnd.n3743 585
R11263 gnd.n3745 gnd.n3744 585
R11264 gnd.n2155 gnd.n2154 585
R11265 gnd.n2162 gnd.n2154 585
R11266 gnd.n3739 gnd.n3738 585
R11267 gnd.n3738 gnd.n3737 585
R11268 gnd.n2158 gnd.n2157 585
R11269 gnd.n2168 gnd.n2158 585
R11270 gnd.n3698 gnd.n2185 585
R11271 gnd.n2185 gnd.n2178 585
R11272 gnd.n3700 gnd.n3699 585
R11273 gnd.n3701 gnd.n3700 585
R11274 gnd.n2186 gnd.n2184 585
R11275 gnd.n3673 gnd.n2184 585
R11276 gnd.n3693 gnd.n3692 585
R11277 gnd.n3692 gnd.n3691 585
R11278 gnd.n2189 gnd.n2188 585
R11279 gnd.n3683 gnd.n2189 585
R11280 gnd.n3654 gnd.n3653 585
R11281 gnd.n3655 gnd.n3654 585
R11282 gnd.n2202 gnd.n2201 585
R11283 gnd.n3574 gnd.n2201 585
R11284 gnd.n3649 gnd.n3648 585
R11285 gnd.n3648 gnd.n3647 585
R11286 gnd.n2205 gnd.n2204 585
R11287 gnd.n3636 gnd.n2205 585
R11288 gnd.n3611 gnd.n3610 585
R11289 gnd.n3612 gnd.n3611 585
R11290 gnd.n2225 gnd.n2224 585
R11291 gnd.n3585 gnd.n2224 585
R11292 gnd.n3606 gnd.n3605 585
R11293 gnd.n3605 gnd.n3604 585
R11294 gnd.n2228 gnd.n2227 585
R11295 gnd.n3593 gnd.n2228 585
R11296 gnd.n3531 gnd.n3530 585
R11297 gnd.n3531 gnd.n2239 585
R11298 gnd.n3536 gnd.n3535 585
R11299 gnd.n3535 gnd.n3534 585
R11300 gnd.n3537 gnd.n2258 585
R11301 gnd.n2258 gnd.n2247 585
R11302 gnd.n3539 gnd.n3538 585
R11303 gnd.n3540 gnd.n3539 585
R11304 gnd.n2259 gnd.n2257 585
R11305 gnd.n2267 gnd.n2257 585
R11306 gnd.n3523 gnd.n3522 585
R11307 gnd.n3522 gnd.n3521 585
R11308 gnd.n2262 gnd.n2261 585
R11309 gnd.n3512 gnd.n2262 585
R11310 gnd.n3486 gnd.n2291 585
R11311 gnd.n2291 gnd.n2283 585
R11312 gnd.n3488 gnd.n3487 585
R11313 gnd.n3489 gnd.n3488 585
R11314 gnd.n2292 gnd.n2290 585
R11315 gnd.n2290 gnd.n2287 585
R11316 gnd.n3481 gnd.n3480 585
R11317 gnd.n3480 gnd.n3479 585
R11318 gnd.n2295 gnd.n2294 585
R11319 gnd.n3469 gnd.n2295 585
R11320 gnd.n3459 gnd.n3458 585
R11321 gnd.n3460 gnd.n3459 585
R11322 gnd.n2314 gnd.n2313 585
R11323 gnd.n3445 gnd.n2313 585
R11324 gnd.n3454 gnd.n3453 585
R11325 gnd.n3453 gnd.n3452 585
R11326 gnd.n2318 gnd.n2317 585
R11327 gnd.n2318 gnd.n1618 585
R11328 gnd.n1607 gnd.n1606 585
R11329 gnd.n1615 gnd.n1607 585
R11330 gnd.n4836 gnd.n4835 585
R11331 gnd.n4835 gnd.n4834 585
R11332 gnd.n4837 gnd.n1601 585
R11333 gnd.n3401 gnd.n1601 585
R11334 gnd.n4839 gnd.n4838 585
R11335 gnd.n4840 gnd.n4839 585
R11336 gnd.n1602 gnd.n1600 585
R11337 gnd.n3393 gnd.n1600 585
R11338 gnd.n3295 gnd.n3294 585
R11339 gnd.n3294 gnd.n1539 585
R11340 gnd.n3296 gnd.n2344 585
R11341 gnd.n2344 gnd.n2332 585
R11342 gnd.n3298 gnd.n3297 585
R11343 gnd.n3299 gnd.n3298 585
R11344 gnd.n2345 gnd.n2343 585
R11345 gnd.n2343 gnd.n2340 585
R11346 gnd.n3287 gnd.n3286 585
R11347 gnd.n3286 gnd.n3285 585
R11348 gnd.n2348 gnd.n2347 585
R11349 gnd.n2357 gnd.n2348 585
R11350 gnd.n3260 gnd.n2369 585
R11351 gnd.n2369 gnd.n2356 585
R11352 gnd.n3262 gnd.n3261 585
R11353 gnd.n3263 gnd.n3262 585
R11354 gnd.n2370 gnd.n2368 585
R11355 gnd.n2368 gnd.n2365 585
R11356 gnd.n3255 gnd.n3254 585
R11357 gnd.n3254 gnd.n3253 585
R11358 gnd.n2373 gnd.n2372 585
R11359 gnd.n2381 gnd.n2373 585
R11360 gnd.n3230 gnd.n2393 585
R11361 gnd.n2393 gnd.n2392 585
R11362 gnd.n3232 gnd.n3231 585
R11363 gnd.n3233 gnd.n3232 585
R11364 gnd.n2394 gnd.n2391 585
R11365 gnd.n2391 gnd.n2388 585
R11366 gnd.n3225 gnd.n3224 585
R11367 gnd.n3224 gnd.n3223 585
R11368 gnd.n2397 gnd.n2396 585
R11369 gnd.n2398 gnd.n2397 585
R11370 gnd.n3100 gnd.n3099 585
R11371 gnd.n3099 gnd.n3098 585
R11372 gnd.n3101 gnd.n3092 585
R11373 gnd.n3097 gnd.n3092 585
R11374 gnd.n3104 gnd.n3102 585
R11375 gnd.n3104 gnd.n3103 585
R11376 gnd.n3105 gnd.n3091 585
R11377 gnd.n3105 gnd.n1482 585
R11378 gnd.n3107 gnd.n3106 585
R11379 gnd.n3106 gnd.n1479 585
R11380 gnd.n3108 gnd.n3086 585
R11381 gnd.n3086 gnd.n1473 585
R11382 gnd.n3110 gnd.n3109 585
R11383 gnd.n3110 gnd.n1470 585
R11384 gnd.n3111 gnd.n3085 585
R11385 gnd.n3111 gnd.n1462 585
R11386 gnd.n3113 gnd.n3112 585
R11387 gnd.n3112 gnd.n1459 585
R11388 gnd.n3114 gnd.n2619 585
R11389 gnd.n2619 gnd.n1452 585
R11390 gnd.n3116 gnd.n3115 585
R11391 gnd.n3117 gnd.n3116 585
R11392 gnd.n2620 gnd.n2618 585
R11393 gnd.n2618 gnd.n1442 585
R11394 gnd.n3079 gnd.n3078 585
R11395 gnd.n3078 gnd.n1439 585
R11396 gnd.n3077 gnd.n2622 585
R11397 gnd.n3077 gnd.n1432 585
R11398 gnd.n3076 gnd.n3075 585
R11399 gnd.n3076 gnd.n1429 585
R11400 gnd.n2624 gnd.n2623 585
R11401 gnd.n3042 gnd.n2623 585
R11402 gnd.n3071 gnd.n3070 585
R11403 gnd.n3070 gnd.n1419 585
R11404 gnd.n3069 gnd.n2626 585
R11405 gnd.n3069 gnd.n1412 585
R11406 gnd.n3068 gnd.n2628 585
R11407 gnd.n3068 gnd.n3067 585
R11408 gnd.n2993 gnd.n2627 585
R11409 gnd.n2627 gnd.n1402 585
R11410 gnd.n2995 gnd.n2994 585
R11411 gnd.n2994 gnd.n1399 585
R11412 gnd.n2996 gnd.n2986 585
R11413 gnd.n2986 gnd.n1392 585
R11414 gnd.n2998 gnd.n2997 585
R11415 gnd.n2998 gnd.n1389 585
R11416 gnd.n2999 gnd.n2985 585
R11417 gnd.n2999 gnd.n2642 585
R11418 gnd.n3001 gnd.n3000 585
R11419 gnd.n3000 gnd.n1380 585
R11420 gnd.n3002 gnd.n2651 585
R11421 gnd.n2651 gnd.n1371 585
R11422 gnd.n3005 gnd.n3004 585
R11423 gnd.n3006 gnd.n3005 585
R11424 gnd.n2983 gnd.n2650 585
R11425 gnd.n2650 gnd.n2648 585
R11426 gnd.n2981 gnd.n2980 585
R11427 gnd.n2980 gnd.n2979 585
R11428 gnd.n2653 gnd.n2652 585
R11429 gnd.n2663 gnd.n2653 585
R11430 gnd.n2922 gnd.n2920 585
R11431 gnd.n2920 gnd.n2660 585
R11432 gnd.n2924 gnd.n2923 585
R11433 gnd.n2924 gnd.n2684 585
R11434 gnd.n2926 gnd.n2925 585
R11435 gnd.n2925 gnd.n2680 585
R11436 gnd.n2927 gnd.n2692 585
R11437 gnd.n2692 gnd.n2678 585
R11438 gnd.n2930 gnd.n2929 585
R11439 gnd.n2931 gnd.n2930 585
R11440 gnd.n2918 gnd.n2691 585
R11441 gnd.n2691 gnd.n1354 585
R11442 gnd.n2912 gnd.n2693 585
R11443 gnd.n2912 gnd.n1351 585
R11444 gnd.n2914 gnd.n2913 585
R11445 gnd.n2913 gnd.n1344 585
R11446 gnd.n2911 gnd.n2695 585
R11447 gnd.n2911 gnd.n1341 585
R11448 gnd.n2910 gnd.n2909 585
R11449 gnd.n2910 gnd.n1333 585
R11450 gnd.n2697 gnd.n2696 585
R11451 gnd.n2696 gnd.n1330 585
R11452 gnd.n2905 gnd.n2904 585
R11453 gnd.n2904 gnd.n1323 585
R11454 gnd.n2903 gnd.n2699 585
R11455 gnd.n2903 gnd.n2902 585
R11456 gnd.n2825 gnd.n2700 585
R11457 gnd.n2700 gnd.n1313 585
R11458 gnd.n2827 gnd.n2826 585
R11459 gnd.n2826 gnd.n1310 585
R11460 gnd.n2828 gnd.n2819 585
R11461 gnd.n2819 gnd.n1303 585
R11462 gnd.n2830 gnd.n2829 585
R11463 gnd.n2830 gnd.n1300 585
R11464 gnd.n2831 gnd.n2818 585
R11465 gnd.n2831 gnd.n1292 585
R11466 gnd.n2833 gnd.n2832 585
R11467 gnd.n2832 gnd.n1289 585
R11468 gnd.n2834 gnd.n2796 585
R11469 gnd.n2796 gnd.n1282 585
R11470 gnd.n2836 gnd.n2835 585
R11471 gnd.n2837 gnd.n2836 585
R11472 gnd.n2797 gnd.n2795 585
R11473 gnd.n2795 gnd.n1272 585
R11474 gnd.n2812 gnd.n2811 585
R11475 gnd.n2811 gnd.n1269 585
R11476 gnd.n2810 gnd.n2799 585
R11477 gnd.n2810 gnd.n1261 585
R11478 gnd.n2809 gnd.n2808 585
R11479 gnd.n2809 gnd.n1258 585
R11480 gnd.n2801 gnd.n2800 585
R11481 gnd.n2800 gnd.n1249 585
R11482 gnd.n2804 gnd.n2803 585
R11483 gnd.n2803 gnd.n1244 585
R11484 gnd.n1130 gnd.n1129 585
R11485 gnd.n1169 gnd.n1130 585
R11486 gnd.n5229 gnd.n5228 585
R11487 gnd.n5228 gnd.n5227 585
R11488 gnd.n5230 gnd.n1126 585
R11489 gnd.n1126 gnd.n1125 585
R11490 gnd.n4728 gnd.n4727 585
R11491 gnd.n4727 gnd.n4726 585
R11492 gnd.n4729 gnd.n1701 585
R11493 gnd.n4106 gnd.n1701 585
R11494 gnd.n4730 gnd.n1700 585
R11495 gnd.n2050 gnd.n1700 585
R11496 gnd.n4117 gnd.n1698 585
R11497 gnd.n4118 gnd.n4117 585
R11498 gnd.n4734 gnd.n1697 585
R11499 gnd.n4120 gnd.n1697 585
R11500 gnd.n4735 gnd.n1696 585
R11501 gnd.n2047 gnd.n1696 585
R11502 gnd.n4736 gnd.n1695 585
R11503 gnd.n2057 gnd.n1695 585
R11504 gnd.n4128 gnd.n1693 585
R11505 gnd.n4129 gnd.n4128 585
R11506 gnd.n4740 gnd.n1692 585
R11507 gnd.n4131 gnd.n1692 585
R11508 gnd.n4741 gnd.n1691 585
R11509 gnd.n2037 gnd.n1691 585
R11510 gnd.n4742 gnd.n1690 585
R11511 gnd.n2028 gnd.n1690 585
R11512 gnd.n4139 gnd.n1688 585
R11513 gnd.n4140 gnd.n4139 585
R11514 gnd.n4746 gnd.n1687 585
R11515 gnd.n4142 gnd.n1687 585
R11516 gnd.n4747 gnd.n1686 585
R11517 gnd.n1971 gnd.n1686 585
R11518 gnd.n4748 gnd.n1685 585
R11519 gnd.n2008 gnd.n1685 585
R11520 gnd.n4150 gnd.n1683 585
R11521 gnd.n4151 gnd.n4150 585
R11522 gnd.n4752 gnd.n1682 585
R11523 gnd.n3900 gnd.n1682 585
R11524 gnd.n4753 gnd.n1681 585
R11525 gnd.n2075 gnd.n1681 585
R11526 gnd.n4754 gnd.n1680 585
R11527 gnd.n2085 gnd.n1680 585
R11528 gnd.n2081 gnd.n1678 585
R11529 gnd.n2082 gnd.n2081 585
R11530 gnd.n4758 gnd.n1677 585
R11531 gnd.n3869 gnd.n1677 585
R11532 gnd.n4759 gnd.n1676 585
R11533 gnd.n3861 gnd.n1676 585
R11534 gnd.n4760 gnd.n1675 585
R11535 gnd.n3759 gnd.n1675 585
R11536 gnd.n3844 gnd.n1673 585
R11537 gnd.n3845 gnd.n3844 585
R11538 gnd.n4764 gnd.n1672 585
R11539 gnd.n3837 gnd.n1672 585
R11540 gnd.n4765 gnd.n1671 585
R11541 gnd.n2121 gnd.n1671 585
R11542 gnd.n4766 gnd.n1670 585
R11543 gnd.n3816 gnd.n1670 585
R11544 gnd.n2125 gnd.n1668 585
R11545 gnd.n2126 gnd.n2125 585
R11546 gnd.n4770 gnd.n1667 585
R11547 gnd.n3807 gnd.n1667 585
R11548 gnd.n4771 gnd.n1666 585
R11549 gnd.n3778 gnd.n1666 585
R11550 gnd.n4772 gnd.n1665 585
R11551 gnd.n2142 gnd.n1665 585
R11552 gnd.n2148 gnd.n1663 585
R11553 gnd.n2149 gnd.n2148 585
R11554 gnd.n4776 gnd.n1662 585
R11555 gnd.n2153 gnd.n1662 585
R11556 gnd.n4777 gnd.n1661 585
R11557 gnd.n3736 gnd.n1661 585
R11558 gnd.n4778 gnd.n1660 585
R11559 gnd.n3727 gnd.n1660 585
R11560 gnd.n3664 gnd.n1658 585
R11561 gnd.n3665 gnd.n3664 585
R11562 gnd.n4782 gnd.n1657 585
R11563 gnd.n3709 gnd.n1657 585
R11564 gnd.n4783 gnd.n1656 585
R11565 gnd.n2182 gnd.n1656 585
R11566 gnd.n4784 gnd.n1655 585
R11567 gnd.n2191 gnd.n1655 585
R11568 gnd.n3681 gnd.n1653 585
R11569 gnd.n3682 gnd.n3681 585
R11570 gnd.n4788 gnd.n1652 585
R11571 gnd.n2195 gnd.n1652 585
R11572 gnd.n4789 gnd.n1651 585
R11573 gnd.n2200 gnd.n1651 585
R11574 gnd.n4790 gnd.n1650 585
R11575 gnd.n2207 gnd.n1650 585
R11576 gnd.n3633 gnd.n1648 585
R11577 gnd.n3634 gnd.n3633 585
R11578 gnd.n4794 gnd.n1647 585
R11579 gnd.n2212 gnd.n1647 585
R11580 gnd.n4795 gnd.n1646 585
R11581 gnd.n3613 gnd.n1646 585
R11582 gnd.n4796 gnd.n1645 585
R11583 gnd.n3584 gnd.n1645 585
R11584 gnd.n2229 gnd.n1643 585
R11585 gnd.n2230 gnd.n2229 585
R11586 gnd.n4800 gnd.n1642 585
R11587 gnd.n3568 gnd.n1642 585
R11588 gnd.n4801 gnd.n1641 585
R11589 gnd.n3532 gnd.n1641 585
R11590 gnd.n4802 gnd.n1640 585
R11591 gnd.n3559 gnd.n1640 585
R11592 gnd.n3549 gnd.n1638 585
R11593 gnd.n3550 gnd.n3549 585
R11594 gnd.n4806 gnd.n1637 585
R11595 gnd.n2256 gnd.n1637 585
R11596 gnd.n4807 gnd.n1636 585
R11597 gnd.n2265 gnd.n1636 585
R11598 gnd.n4808 gnd.n1635 585
R11599 gnd.n3511 gnd.n1635 585
R11600 gnd.n2272 gnd.n1633 585
R11601 gnd.n2273 gnd.n2272 585
R11602 gnd.n4812 gnd.n1632 585
R11603 gnd.n3499 gnd.n1632 585
R11604 gnd.n4813 gnd.n1631 585
R11605 gnd.n3491 gnd.n1631 585
R11606 gnd.n4814 gnd.n1630 585
R11607 gnd.n3478 gnd.n1630 585
R11608 gnd.n2305 gnd.n1628 585
R11609 gnd.n2306 gnd.n2305 585
R11610 gnd.n4818 gnd.n1627 585
R11611 gnd.n3470 gnd.n1627 585
R11612 gnd.n4819 gnd.n1626 585
R11613 gnd.n2311 gnd.n1626 585
R11614 gnd.n4820 gnd.n1625 585
R11615 gnd.n3446 gnd.n1625 585
R11616 gnd.n1622 gnd.n1620 585
R11617 gnd.n3419 gnd.n1620 585
R11618 gnd.n4825 gnd.n4824 585
R11619 gnd.n4826 gnd.n4825 585
R11620 gnd.n1621 gnd.n1619 585
R11621 gnd.n3410 gnd.n1619 585
R11622 gnd.n3310 gnd.n3308 585
R11623 gnd.n3308 gnd.n1608 585
R11624 gnd.n3311 gnd.n3307 585
R11625 gnd.n3307 gnd.n1599 585
R11626 gnd.n3312 gnd.n3306 585
R11627 gnd.n3306 gnd.n1597 585
R11628 gnd.n2336 gnd.n2334 585
R11629 gnd.n2334 gnd.n1571 585
R11630 gnd.n3317 gnd.n3316 585
R11631 gnd.n3318 gnd.n3317 585
R11632 gnd.n2335 gnd.n2333 585
R11633 gnd.n2342 gnd.n2333 585
R11634 gnd.n3302 gnd.n3301 585
R11635 gnd.n3301 gnd.n3300 585
R11636 gnd.n2339 gnd.n2338 585
R11637 gnd.n3284 gnd.n2339 585
R11638 gnd.n2361 gnd.n2359 585
R11639 gnd.n2359 gnd.n2349 585
R11640 gnd.n3272 gnd.n3271 585
R11641 gnd.n3273 gnd.n3272 585
R11642 gnd.n2360 gnd.n2358 585
R11643 gnd.n2367 gnd.n2358 585
R11644 gnd.n3266 gnd.n3265 585
R11645 gnd.n3265 gnd.n3264 585
R11646 gnd.n2364 gnd.n2363 585
R11647 gnd.n3252 gnd.n2364 585
R11648 gnd.n2385 gnd.n2383 585
R11649 gnd.n2383 gnd.n2374 585
R11650 gnd.n3242 gnd.n3241 585
R11651 gnd.n3243 gnd.n3242 585
R11652 gnd.n2384 gnd.n2382 585
R11653 gnd.n2390 gnd.n2382 585
R11654 gnd.n3236 gnd.n3235 585
R11655 gnd.n3235 gnd.n3234 585
R11656 gnd.n2413 gnd.n2387 585
R11657 gnd.n3220 gnd.n3219 585
R11658 gnd.n2414 gnd.n2412 585
R11659 gnd.n3222 gnd.n2412 585
R11660 gnd.n3215 gnd.n2416 585
R11661 gnd.n3214 gnd.n2417 585
R11662 gnd.n3213 gnd.n2418 585
R11663 gnd.n2534 gnd.n2419 585
R11664 gnd.n3208 gnd.n2535 585
R11665 gnd.n3207 gnd.n2536 585
R11666 gnd.n3206 gnd.n2537 585
R11667 gnd.n2547 gnd.n2538 585
R11668 gnd.n3199 gnd.n2548 585
R11669 gnd.n3198 gnd.n2549 585
R11670 gnd.n2551 gnd.n2550 585
R11671 gnd.n3191 gnd.n2559 585
R11672 gnd.n3190 gnd.n2560 585
R11673 gnd.n2570 gnd.n2561 585
R11674 gnd.n3183 gnd.n2571 585
R11675 gnd.n3182 gnd.n2572 585
R11676 gnd.n2574 gnd.n2573 585
R11677 gnd.n3175 gnd.n2582 585
R11678 gnd.n3174 gnd.n2583 585
R11679 gnd.n2593 gnd.n2584 585
R11680 gnd.n3167 gnd.n2594 585
R11681 gnd.n3166 gnd.n2595 585
R11682 gnd.n3147 gnd.n3146 585
R11683 gnd.n3149 gnd.n3148 585
R11684 gnd.n3156 gnd.n3150 585
R11685 gnd.n3155 gnd.n3151 585
R11686 gnd.n2053 gnd.n1705 585
R11687 gnd.n4726 gnd.n1705 585
R11688 gnd.n4105 gnd.n4104 585
R11689 gnd.n4106 gnd.n4105 585
R11690 gnd.n2052 gnd.n2051 585
R11691 gnd.n2051 gnd.n2050 585
R11692 gnd.n3921 gnd.n2049 585
R11693 gnd.n4118 gnd.n2049 585
R11694 gnd.n3920 gnd.n2048 585
R11695 gnd.n4120 gnd.n2048 585
R11696 gnd.n3919 gnd.n2059 585
R11697 gnd.n2059 gnd.n2047 585
R11698 gnd.n2058 gnd.n2055 585
R11699 gnd.n2058 gnd.n2057 585
R11700 gnd.n3915 gnd.n2039 585
R11701 gnd.n4129 gnd.n2039 585
R11702 gnd.n3914 gnd.n2038 585
R11703 gnd.n4131 gnd.n2038 585
R11704 gnd.n3913 gnd.n2063 585
R11705 gnd.n2063 gnd.n2037 585
R11706 gnd.n2062 gnd.n2061 585
R11707 gnd.n2062 gnd.n2028 585
R11708 gnd.n3909 gnd.n2027 585
R11709 gnd.n4140 gnd.n2027 585
R11710 gnd.n3908 gnd.n2026 585
R11711 gnd.n4142 gnd.n2026 585
R11712 gnd.n3907 gnd.n2067 585
R11713 gnd.n2067 gnd.n1971 585
R11714 gnd.n2066 gnd.n2065 585
R11715 gnd.n2066 gnd.n2008 585
R11716 gnd.n3903 gnd.n2016 585
R11717 gnd.n4151 gnd.n2016 585
R11718 gnd.n3902 gnd.n3901 585
R11719 gnd.n3901 gnd.n3900 585
R11720 gnd.n2070 gnd.n2069 585
R11721 gnd.n2075 gnd.n2070 585
R11722 gnd.n3854 gnd.n3853 585
R11723 gnd.n3853 gnd.n2085 585
R11724 gnd.n3855 gnd.n3852 585
R11725 gnd.n3852 gnd.n2082 585
R11726 gnd.n2103 gnd.n2093 585
R11727 gnd.n3869 gnd.n2093 585
R11728 gnd.n3860 gnd.n3859 585
R11729 gnd.n3861 gnd.n3860 585
R11730 gnd.n2102 gnd.n2101 585
R11731 gnd.n3759 gnd.n2101 585
R11732 gnd.n3847 gnd.n3846 585
R11733 gnd.n3846 gnd.n3845 585
R11734 gnd.n2106 gnd.n2105 585
R11735 gnd.n3837 gnd.n2106 585
R11736 gnd.n2132 gnd.n2130 585
R11737 gnd.n2130 gnd.n2121 585
R11738 gnd.n3815 gnd.n3814 585
R11739 gnd.n3816 gnd.n3815 585
R11740 gnd.n2131 gnd.n2129 585
R11741 gnd.n2129 gnd.n2126 585
R11742 gnd.n3809 gnd.n3808 585
R11743 gnd.n3808 gnd.n3807 585
R11744 gnd.n2135 gnd.n2134 585
R11745 gnd.n3778 gnd.n2135 585
R11746 gnd.n3719 gnd.n3717 585
R11747 gnd.n3717 gnd.n2142 585
R11748 gnd.n3720 gnd.n3716 585
R11749 gnd.n3716 gnd.n2149 585
R11750 gnd.n3721 gnd.n3715 585
R11751 gnd.n3715 gnd.n2153 585
R11752 gnd.n2172 gnd.n2160 585
R11753 gnd.n3736 gnd.n2160 585
R11754 gnd.n3726 gnd.n3725 585
R11755 gnd.n3727 gnd.n3726 585
R11756 gnd.n2171 gnd.n2170 585
R11757 gnd.n3665 gnd.n2170 585
R11758 gnd.n3711 gnd.n3710 585
R11759 gnd.n3710 gnd.n3709 585
R11760 gnd.n2175 gnd.n2174 585
R11761 gnd.n2182 gnd.n2175 585
R11762 gnd.n3622 gnd.n3621 585
R11763 gnd.n3621 gnd.n2191 585
R11764 gnd.n3625 gnd.n2197 585
R11765 gnd.n3682 gnd.n2197 585
R11766 gnd.n3626 gnd.n3620 585
R11767 gnd.n3620 gnd.n2195 585
R11768 gnd.n3627 gnd.n3619 585
R11769 gnd.n3619 gnd.n2200 585
R11770 gnd.n2218 gnd.n2216 585
R11771 gnd.n2216 gnd.n2207 585
R11772 gnd.n3632 gnd.n3631 585
R11773 gnd.n3634 gnd.n3632 585
R11774 gnd.n2217 gnd.n2215 585
R11775 gnd.n2215 gnd.n2212 585
R11776 gnd.n3615 gnd.n3614 585
R11777 gnd.n3614 gnd.n3613 585
R11778 gnd.n2221 gnd.n2220 585
R11779 gnd.n3584 gnd.n2221 585
R11780 gnd.n2243 gnd.n2241 585
R11781 gnd.n2241 gnd.n2230 585
R11782 gnd.n3567 gnd.n3566 585
R11783 gnd.n3568 gnd.n3567 585
R11784 gnd.n2242 gnd.n2240 585
R11785 gnd.n3532 gnd.n2240 585
R11786 gnd.n3561 gnd.n3560 585
R11787 gnd.n3560 gnd.n3559 585
R11788 gnd.n2246 gnd.n2245 585
R11789 gnd.n3550 gnd.n2246 585
R11790 gnd.n3505 gnd.n3504 585
R11791 gnd.n3504 gnd.n2256 585
R11792 gnd.n2278 gnd.n2276 585
R11793 gnd.n2276 gnd.n2265 585
R11794 gnd.n3510 gnd.n3509 585
R11795 gnd.n3511 gnd.n3510 585
R11796 gnd.n2277 gnd.n2275 585
R11797 gnd.n2275 gnd.n2273 585
R11798 gnd.n3501 gnd.n3500 585
R11799 gnd.n3500 gnd.n3499 585
R11800 gnd.n2281 gnd.n2280 585
R11801 gnd.n3491 gnd.n2281 585
R11802 gnd.n3477 gnd.n3476 585
R11803 gnd.n3478 gnd.n3477 585
R11804 gnd.n2299 gnd.n2298 585
R11805 gnd.n2306 gnd.n2298 585
R11806 gnd.n3472 gnd.n3471 585
R11807 gnd.n3471 gnd.n3470 585
R11808 gnd.n2302 gnd.n2301 585
R11809 gnd.n2311 gnd.n2302 585
R11810 gnd.n2324 gnd.n2321 585
R11811 gnd.n3446 gnd.n2321 585
R11812 gnd.n3418 gnd.n3417 585
R11813 gnd.n3419 gnd.n3418 585
R11814 gnd.n2323 gnd.n1617 585
R11815 gnd.n4826 gnd.n1617 585
R11816 gnd.n3412 gnd.n3411 585
R11817 gnd.n3411 gnd.n3410 585
R11818 gnd.n3327 gnd.n2326 585
R11819 gnd.n3327 gnd.n1608 585
R11820 gnd.n3326 gnd.n3325 585
R11821 gnd.n3326 gnd.n1599 585
R11822 gnd.n2328 gnd.n2327 585
R11823 gnd.n2327 gnd.n1597 585
R11824 gnd.n3321 gnd.n3320 585
R11825 gnd.n3320 gnd.n1571 585
R11826 gnd.n3319 gnd.n2330 585
R11827 gnd.n3319 gnd.n3318 585
R11828 gnd.n3278 gnd.n2331 585
R11829 gnd.n2342 gnd.n2331 585
R11830 gnd.n2352 gnd.n2341 585
R11831 gnd.n3300 gnd.n2341 585
R11832 gnd.n3283 gnd.n3282 585
R11833 gnd.n3284 gnd.n3283 585
R11834 gnd.n2351 gnd.n2350 585
R11835 gnd.n2350 gnd.n2349 585
R11836 gnd.n3275 gnd.n3274 585
R11837 gnd.n3274 gnd.n3273 585
R11838 gnd.n2355 gnd.n2354 585
R11839 gnd.n2367 gnd.n2355 585
R11840 gnd.n2377 gnd.n2366 585
R11841 gnd.n3264 gnd.n2366 585
R11842 gnd.n3251 gnd.n3250 585
R11843 gnd.n3252 gnd.n3251 585
R11844 gnd.n2376 gnd.n2375 585
R11845 gnd.n2375 gnd.n2374 585
R11846 gnd.n3245 gnd.n3244 585
R11847 gnd.n3244 gnd.n3243 585
R11848 gnd.n2380 gnd.n2379 585
R11849 gnd.n2390 gnd.n2380 585
R11850 gnd.n3152 gnd.n2389 585
R11851 gnd.n3234 gnd.n2389 585
R11852 gnd.n4079 gnd.n3933 585
R11853 gnd.n3933 gnd.n1715 585
R11854 gnd.n4080 gnd.n4077 585
R11855 gnd.n4075 gnd.n3951 585
R11856 gnd.n4074 gnd.n4073 585
R11857 gnd.n4058 gnd.n3953 585
R11858 gnd.n4060 gnd.n4059 585
R11859 gnd.n4056 gnd.n3960 585
R11860 gnd.n4055 gnd.n4054 585
R11861 gnd.n4039 gnd.n3962 585
R11862 gnd.n4041 gnd.n4040 585
R11863 gnd.n4037 gnd.n3969 585
R11864 gnd.n4036 gnd.n4035 585
R11865 gnd.n4020 gnd.n3971 585
R11866 gnd.n4022 gnd.n4021 585
R11867 gnd.n4018 gnd.n3978 585
R11868 gnd.n4017 gnd.n4016 585
R11869 gnd.n4005 gnd.n3980 585
R11870 gnd.n4007 gnd.n4006 585
R11871 gnd.n4003 gnd.n3981 585
R11872 gnd.n4002 gnd.n4001 585
R11873 gnd.n3994 gnd.n3983 585
R11874 gnd.n3996 gnd.n3995 585
R11875 gnd.n3992 gnd.n3985 585
R11876 gnd.n3991 gnd.n3990 585
R11877 gnd.n3987 gnd.n1703 585
R11878 gnd.n4100 gnd.n4099 585
R11879 gnd.n4097 gnd.n3931 585
R11880 gnd.n4096 gnd.n3932 585
R11881 gnd.n4094 gnd.n4093 585
R11882 gnd.n3328 gnd.t121 543.808
R11883 gnd.n2004 gnd.t118 543.808
R11884 gnd.n4846 gnd.t52 543.808
R11885 gnd.n4175 gnd.t45 543.808
R11886 gnd.n6797 gnd.n6796 540.215
R11887 gnd.n4241 gnd.n2011 458.866
R11888 gnd.n4244 gnd.n4243 458.866
R11889 gnd.n3395 gnd.n3392 458.866
R11890 gnd.n4909 gnd.n1574 458.866
R11891 gnd.n2596 gnd.t68 371.625
R11892 gnd.n3944 gnd.t88 371.625
R11893 gnd.n2603 gnd.t110 371.625
R11894 gnd.n4381 gnd.t85 371.625
R11895 gnd.n4433 gnd.t79 371.625
R11896 gnd.n1935 gnd.t19 371.625
R11897 gnd.n317 gnd.t107 371.625
R11898 gnd.n284 gnd.t27 371.625
R11899 gnd.n7770 gnd.t72 371.625
R11900 gnd.n354 gnd.t62 371.625
R11901 gnd.n1191 gnd.t38 371.625
R11902 gnd.n1213 gnd.t35 371.625
R11903 gnd.n1235 gnd.t23 371.625
R11904 gnd.n2720 gnd.t94 371.625
R11905 gnd.n1515 gnd.t100 371.625
R11906 gnd.n2421 gnd.t31 371.625
R11907 gnd.n2443 gnd.t65 371.625
R11908 gnd.n3934 gnd.t41 371.625
R11909 gnd.n7529 gnd.n7528 368.44
R11910 gnd.n5661 gnd.t75 323.425
R11911 gnd.n5266 gnd.t103 323.425
R11912 gnd.n7318 gnd.n7317 301.784
R11913 gnd.n7318 gnd.n554 301.784
R11914 gnd.n7326 gnd.n554 301.784
R11915 gnd.n7327 gnd.n7326 301.784
R11916 gnd.n7328 gnd.n7327 301.784
R11917 gnd.n7328 gnd.n548 301.784
R11918 gnd.n7336 gnd.n548 301.784
R11919 gnd.n7337 gnd.n7336 301.784
R11920 gnd.n7338 gnd.n7337 301.784
R11921 gnd.n7338 gnd.n542 301.784
R11922 gnd.n7346 gnd.n542 301.784
R11923 gnd.n7347 gnd.n7346 301.784
R11924 gnd.n7348 gnd.n7347 301.784
R11925 gnd.n7348 gnd.n536 301.784
R11926 gnd.n7356 gnd.n536 301.784
R11927 gnd.n7357 gnd.n7356 301.784
R11928 gnd.n7358 gnd.n7357 301.784
R11929 gnd.n7358 gnd.n530 301.784
R11930 gnd.n7366 gnd.n530 301.784
R11931 gnd.n7367 gnd.n7366 301.784
R11932 gnd.n7368 gnd.n7367 301.784
R11933 gnd.n7368 gnd.n524 301.784
R11934 gnd.n7376 gnd.n524 301.784
R11935 gnd.n7377 gnd.n7376 301.784
R11936 gnd.n7378 gnd.n7377 301.784
R11937 gnd.n7378 gnd.n518 301.784
R11938 gnd.n7386 gnd.n518 301.784
R11939 gnd.n7387 gnd.n7386 301.784
R11940 gnd.n7388 gnd.n7387 301.784
R11941 gnd.n7388 gnd.n512 301.784
R11942 gnd.n7396 gnd.n512 301.784
R11943 gnd.n7397 gnd.n7396 301.784
R11944 gnd.n7398 gnd.n7397 301.784
R11945 gnd.n7398 gnd.n506 301.784
R11946 gnd.n7406 gnd.n506 301.784
R11947 gnd.n7407 gnd.n7406 301.784
R11948 gnd.n7408 gnd.n7407 301.784
R11949 gnd.n7408 gnd.n500 301.784
R11950 gnd.n7416 gnd.n500 301.784
R11951 gnd.n7417 gnd.n7416 301.784
R11952 gnd.n7418 gnd.n7417 301.784
R11953 gnd.n7418 gnd.n494 301.784
R11954 gnd.n7426 gnd.n494 301.784
R11955 gnd.n7427 gnd.n7426 301.784
R11956 gnd.n7428 gnd.n7427 301.784
R11957 gnd.n7428 gnd.n488 301.784
R11958 gnd.n7436 gnd.n488 301.784
R11959 gnd.n7437 gnd.n7436 301.784
R11960 gnd.n7438 gnd.n7437 301.784
R11961 gnd.n7438 gnd.n482 301.784
R11962 gnd.n7446 gnd.n482 301.784
R11963 gnd.n7447 gnd.n7446 301.784
R11964 gnd.n7448 gnd.n7447 301.784
R11965 gnd.n7448 gnd.n476 301.784
R11966 gnd.n7456 gnd.n476 301.784
R11967 gnd.n7457 gnd.n7456 301.784
R11968 gnd.n7458 gnd.n7457 301.784
R11969 gnd.n7458 gnd.n470 301.784
R11970 gnd.n7466 gnd.n470 301.784
R11971 gnd.n7467 gnd.n7466 301.784
R11972 gnd.n7468 gnd.n7467 301.784
R11973 gnd.n7468 gnd.n464 301.784
R11974 gnd.n7476 gnd.n464 301.784
R11975 gnd.n7477 gnd.n7476 301.784
R11976 gnd.n7478 gnd.n7477 301.784
R11977 gnd.n7478 gnd.n458 301.784
R11978 gnd.n7486 gnd.n458 301.784
R11979 gnd.n7487 gnd.n7486 301.784
R11980 gnd.n7488 gnd.n7487 301.784
R11981 gnd.n7488 gnd.n452 301.784
R11982 gnd.n7496 gnd.n452 301.784
R11983 gnd.n7497 gnd.n7496 301.784
R11984 gnd.n7498 gnd.n7497 301.784
R11985 gnd.n7498 gnd.n446 301.784
R11986 gnd.n7506 gnd.n446 301.784
R11987 gnd.n7507 gnd.n7506 301.784
R11988 gnd.n7508 gnd.n7507 301.784
R11989 gnd.n7508 gnd.n440 301.784
R11990 gnd.n7516 gnd.n440 301.784
R11991 gnd.n7517 gnd.n7516 301.784
R11992 gnd.n7518 gnd.n7517 301.784
R11993 gnd.n7518 gnd.n434 301.784
R11994 gnd.n7528 gnd.n434 301.784
R11995 gnd.n6439 gnd.n6413 289.615
R11996 gnd.n6407 gnd.n6381 289.615
R11997 gnd.n6375 gnd.n6349 289.615
R11998 gnd.n6344 gnd.n6318 289.615
R11999 gnd.n6312 gnd.n6286 289.615
R12000 gnd.n6280 gnd.n6254 289.615
R12001 gnd.n6248 gnd.n6222 289.615
R12002 gnd.n6217 gnd.n6191 289.615
R12003 gnd.n5735 gnd.t12 279.217
R12004 gnd.n5310 gnd.t5 279.217
R12005 gnd.n1581 gnd.t18 260.649
R12006 gnd.n4167 gnd.t51 260.649
R12007 gnd.n4911 gnd.n4910 256.663
R12008 gnd.n4911 gnd.n1540 256.663
R12009 gnd.n4911 gnd.n1541 256.663
R12010 gnd.n4911 gnd.n1542 256.663
R12011 gnd.n4911 gnd.n1543 256.663
R12012 gnd.n4911 gnd.n1544 256.663
R12013 gnd.n4911 gnd.n1545 256.663
R12014 gnd.n4911 gnd.n1546 256.663
R12015 gnd.n4911 gnd.n1547 256.663
R12016 gnd.n4911 gnd.n1548 256.663
R12017 gnd.n4911 gnd.n1549 256.663
R12018 gnd.n4911 gnd.n1550 256.663
R12019 gnd.n4911 gnd.n1551 256.663
R12020 gnd.n4911 gnd.n1552 256.663
R12021 gnd.n4911 gnd.n1553 256.663
R12022 gnd.n4911 gnd.n1554 256.663
R12023 gnd.n4914 gnd.n1537 256.663
R12024 gnd.n4912 gnd.n4911 256.663
R12025 gnd.n4911 gnd.n1555 256.663
R12026 gnd.n4911 gnd.n1556 256.663
R12027 gnd.n4911 gnd.n1557 256.663
R12028 gnd.n4911 gnd.n1558 256.663
R12029 gnd.n4911 gnd.n1559 256.663
R12030 gnd.n4911 gnd.n1560 256.663
R12031 gnd.n4911 gnd.n1561 256.663
R12032 gnd.n4911 gnd.n1562 256.663
R12033 gnd.n4911 gnd.n1563 256.663
R12034 gnd.n4911 gnd.n1564 256.663
R12035 gnd.n4911 gnd.n1565 256.663
R12036 gnd.n4911 gnd.n1566 256.663
R12037 gnd.n4911 gnd.n1567 256.663
R12038 gnd.n4911 gnd.n1568 256.663
R12039 gnd.n4911 gnd.n1569 256.663
R12040 gnd.n4911 gnd.n1570 256.663
R12041 gnd.n4309 gnd.n1988 256.663
R12042 gnd.n4309 gnd.n1989 256.663
R12043 gnd.n4309 gnd.n1990 256.663
R12044 gnd.n4309 gnd.n1991 256.663
R12045 gnd.n4309 gnd.n1992 256.663
R12046 gnd.n4309 gnd.n1993 256.663
R12047 gnd.n4309 gnd.n1994 256.663
R12048 gnd.n4309 gnd.n1995 256.663
R12049 gnd.n4309 gnd.n1996 256.663
R12050 gnd.n4309 gnd.n1997 256.663
R12051 gnd.n4309 gnd.n1998 256.663
R12052 gnd.n4309 gnd.n1999 256.663
R12053 gnd.n4309 gnd.n2000 256.663
R12054 gnd.n4309 gnd.n2001 256.663
R12055 gnd.n4309 gnd.n2002 256.663
R12056 gnd.n4309 gnd.n4306 256.663
R12057 gnd.n4312 gnd.n1969 256.663
R12058 gnd.n4310 gnd.n4309 256.663
R12059 gnd.n4309 gnd.n1987 256.663
R12060 gnd.n4309 gnd.n1986 256.663
R12061 gnd.n4309 gnd.n1985 256.663
R12062 gnd.n4309 gnd.n1984 256.663
R12063 gnd.n4309 gnd.n1983 256.663
R12064 gnd.n4309 gnd.n1982 256.663
R12065 gnd.n4309 gnd.n1981 256.663
R12066 gnd.n4309 gnd.n1980 256.663
R12067 gnd.n4309 gnd.n1979 256.663
R12068 gnd.n4309 gnd.n1978 256.663
R12069 gnd.n4309 gnd.n1977 256.663
R12070 gnd.n4309 gnd.n1976 256.663
R12071 gnd.n4309 gnd.n1975 256.663
R12072 gnd.n4309 gnd.n1974 256.663
R12073 gnd.n4309 gnd.n1973 256.663
R12074 gnd.n4309 gnd.n1972 256.663
R12075 gnd.n5226 gnd.n1159 242.672
R12076 gnd.n5226 gnd.n1160 242.672
R12077 gnd.n5226 gnd.n1161 242.672
R12078 gnd.n5226 gnd.n1162 242.672
R12079 gnd.n5226 gnd.n1163 242.672
R12080 gnd.n5226 gnd.n1164 242.672
R12081 gnd.n5226 gnd.n1165 242.672
R12082 gnd.n5226 gnd.n1166 242.672
R12083 gnd.n5226 gnd.n1167 242.672
R12084 gnd.n3159 gnd.n1487 242.672
R12085 gnd.n2601 gnd.n1487 242.672
R12086 gnd.n2589 gnd.n1487 242.672
R12087 gnd.n2586 gnd.n1487 242.672
R12088 gnd.n2577 gnd.n1487 242.672
R12089 gnd.n2566 gnd.n1487 242.672
R12090 gnd.n2563 gnd.n1487 242.672
R12091 gnd.n2554 gnd.n1487 242.672
R12092 gnd.n2543 gnd.n1487 242.672
R12093 gnd.n5789 gnd.n5788 242.672
R12094 gnd.n5789 gnd.n5699 242.672
R12095 gnd.n5789 gnd.n5700 242.672
R12096 gnd.n5789 gnd.n5701 242.672
R12097 gnd.n5789 gnd.n5702 242.672
R12098 gnd.n5789 gnd.n5703 242.672
R12099 gnd.n5789 gnd.n5704 242.672
R12100 gnd.n5789 gnd.n5705 242.672
R12101 gnd.n5789 gnd.n5706 242.672
R12102 gnd.n5789 gnd.n5707 242.672
R12103 gnd.n5789 gnd.n5708 242.672
R12104 gnd.n5789 gnd.n5709 242.672
R12105 gnd.n5790 gnd.n5789 242.672
R12106 gnd.n6495 gnd.n5236 242.672
R12107 gnd.n6501 gnd.n5236 242.672
R12108 gnd.n5313 gnd.n5236 242.672
R12109 gnd.n6508 gnd.n5236 242.672
R12110 gnd.n5304 gnd.n5236 242.672
R12111 gnd.n6515 gnd.n5236 242.672
R12112 gnd.n5297 gnd.n5236 242.672
R12113 gnd.n6522 gnd.n5236 242.672
R12114 gnd.n5290 gnd.n5236 242.672
R12115 gnd.n6529 gnd.n5236 242.672
R12116 gnd.n5283 gnd.n5236 242.672
R12117 gnd.n6536 gnd.n5236 242.672
R12118 gnd.n5276 gnd.n5236 242.672
R12119 gnd.n4010 gnd.n1716 242.672
R12120 gnd.n4027 gnd.n1716 242.672
R12121 gnd.n4029 gnd.n1716 242.672
R12122 gnd.n4046 gnd.n1716 242.672
R12123 gnd.n4048 gnd.n1716 242.672
R12124 gnd.n4065 gnd.n1716 242.672
R12125 gnd.n4067 gnd.n1716 242.672
R12126 gnd.n4085 gnd.n1716 242.672
R12127 gnd.n4087 gnd.n1716 242.672
R12128 gnd.n351 gnd.n223 242.672
R12129 gnd.n7666 gnd.n223 242.672
R12130 gnd.n347 gnd.n223 242.672
R12131 gnd.n7673 gnd.n223 242.672
R12132 gnd.n340 gnd.n223 242.672
R12133 gnd.n7680 gnd.n223 242.672
R12134 gnd.n333 gnd.n223 242.672
R12135 gnd.n7687 gnd.n223 242.672
R12136 gnd.n326 gnd.n223 242.672
R12137 gnd.n5873 gnd.n5872 242.672
R12138 gnd.n5872 gnd.n5611 242.672
R12139 gnd.n5872 gnd.n5612 242.672
R12140 gnd.n5872 gnd.n5613 242.672
R12141 gnd.n5872 gnd.n5614 242.672
R12142 gnd.n5872 gnd.n5615 242.672
R12143 gnd.n5872 gnd.n5616 242.672
R12144 gnd.n5872 gnd.n5617 242.672
R12145 gnd.n6547 gnd.n5236 242.672
R12146 gnd.n5269 gnd.n5236 242.672
R12147 gnd.n6554 gnd.n5236 242.672
R12148 gnd.n5260 gnd.n5236 242.672
R12149 gnd.n6561 gnd.n5236 242.672
R12150 gnd.n5253 gnd.n5236 242.672
R12151 gnd.n6568 gnd.n5236 242.672
R12152 gnd.n5246 gnd.n5236 242.672
R12153 gnd.n5226 gnd.n5225 242.672
R12154 gnd.n5226 gnd.n1131 242.672
R12155 gnd.n5226 gnd.n1132 242.672
R12156 gnd.n5226 gnd.n1133 242.672
R12157 gnd.n5226 gnd.n1134 242.672
R12158 gnd.n5226 gnd.n1135 242.672
R12159 gnd.n5226 gnd.n1136 242.672
R12160 gnd.n5226 gnd.n1137 242.672
R12161 gnd.n5226 gnd.n1138 242.672
R12162 gnd.n5226 gnd.n1139 242.672
R12163 gnd.n5226 gnd.n1140 242.672
R12164 gnd.n5226 gnd.n1141 242.672
R12165 gnd.n5226 gnd.n1142 242.672
R12166 gnd.n5226 gnd.n1143 242.672
R12167 gnd.n5226 gnd.n1144 242.672
R12168 gnd.n5226 gnd.n1145 242.672
R12169 gnd.n5226 gnd.n1146 242.672
R12170 gnd.n5226 gnd.n1147 242.672
R12171 gnd.n5226 gnd.n1148 242.672
R12172 gnd.n5226 gnd.n1149 242.672
R12173 gnd.n5226 gnd.n1150 242.672
R12174 gnd.n5226 gnd.n1151 242.672
R12175 gnd.n5226 gnd.n1152 242.672
R12176 gnd.n5226 gnd.n1153 242.672
R12177 gnd.n5226 gnd.n1154 242.672
R12178 gnd.n5226 gnd.n1155 242.672
R12179 gnd.n5226 gnd.n1156 242.672
R12180 gnd.n5226 gnd.n1157 242.672
R12181 gnd.n5226 gnd.n1158 242.672
R12182 gnd.n2528 gnd.n1487 242.672
R12183 gnd.n2424 gnd.n1487 242.672
R12184 gnd.n2518 gnd.n1487 242.672
R12185 gnd.n2428 gnd.n1487 242.672
R12186 gnd.n2508 gnd.n1487 242.672
R12187 gnd.n2432 gnd.n1487 242.672
R12188 gnd.n2498 gnd.n1487 242.672
R12189 gnd.n2436 gnd.n1487 242.672
R12190 gnd.n2488 gnd.n1487 242.672
R12191 gnd.n2440 gnd.n1487 242.672
R12192 gnd.n2478 gnd.n1487 242.672
R12193 gnd.n2446 gnd.n1487 242.672
R12194 gnd.n2468 gnd.n1487 242.672
R12195 gnd.n2450 gnd.n1487 242.672
R12196 gnd.n2458 gnd.n1487 242.672
R12197 gnd.n2455 gnd.n1487 242.672
R12198 gnd.n4915 gnd.n1533 242.672
R12199 gnd.n1532 gnd.n1487 242.672
R12200 gnd.n4919 gnd.n1487 242.672
R12201 gnd.n1526 gnd.n1487 242.672
R12202 gnd.n4926 gnd.n1487 242.672
R12203 gnd.n1519 gnd.n1487 242.672
R12204 gnd.n4934 gnd.n1487 242.672
R12205 gnd.n1510 gnd.n1487 242.672
R12206 gnd.n4941 gnd.n1487 242.672
R12207 gnd.n1503 gnd.n1487 242.672
R12208 gnd.n4948 gnd.n1487 242.672
R12209 gnd.n1496 gnd.n1487 242.672
R12210 gnd.n4955 gnd.n1487 242.672
R12211 gnd.n4958 gnd.n1487 242.672
R12212 gnd.n4342 gnd.n1716 242.672
R12213 gnd.n4345 gnd.n1716 242.672
R12214 gnd.n4353 gnd.n1716 242.672
R12215 gnd.n4355 gnd.n1716 242.672
R12216 gnd.n4363 gnd.n1716 242.672
R12217 gnd.n4365 gnd.n1716 242.672
R12218 gnd.n4373 gnd.n1716 242.672
R12219 gnd.n4375 gnd.n1716 242.672
R12220 gnd.n4386 gnd.n1716 242.672
R12221 gnd.n4388 gnd.n1716 242.672
R12222 gnd.n4396 gnd.n1716 242.672
R12223 gnd.n4398 gnd.n1716 242.672
R12224 gnd.n4407 gnd.n1716 242.672
R12225 gnd.n4408 gnd.n4313 242.672
R12226 gnd.n4409 gnd.n1716 242.672
R12227 gnd.n4411 gnd.n1716 242.672
R12228 gnd.n4419 gnd.n1716 242.672
R12229 gnd.n4421 gnd.n1716 242.672
R12230 gnd.n4429 gnd.n1716 242.672
R12231 gnd.n4431 gnd.n1716 242.672
R12232 gnd.n4441 gnd.n1716 242.672
R12233 gnd.n4443 gnd.n1716 242.672
R12234 gnd.n4451 gnd.n1716 242.672
R12235 gnd.n4453 gnd.n1716 242.672
R12236 gnd.n4461 gnd.n1716 242.672
R12237 gnd.n4463 gnd.n1716 242.672
R12238 gnd.n4471 gnd.n1716 242.672
R12239 gnd.n4473 gnd.n1716 242.672
R12240 gnd.n4482 gnd.n1716 242.672
R12241 gnd.n4485 gnd.n1716 242.672
R12242 gnd.n7698 gnd.n223 242.672
R12243 gnd.n320 gnd.n223 242.672
R12244 gnd.n7705 gnd.n223 242.672
R12245 gnd.n311 gnd.n223 242.672
R12246 gnd.n7712 gnd.n223 242.672
R12247 gnd.n304 gnd.n223 242.672
R12248 gnd.n7719 gnd.n223 242.672
R12249 gnd.n297 gnd.n223 242.672
R12250 gnd.n7726 gnd.n223 242.672
R12251 gnd.n7729 gnd.n223 242.672
R12252 gnd.n288 gnd.n223 242.672
R12253 gnd.n7738 gnd.n223 242.672
R12254 gnd.n279 gnd.n223 242.672
R12255 gnd.n7745 gnd.n223 242.672
R12256 gnd.n272 gnd.n223 242.672
R12257 gnd.n7752 gnd.n223 242.672
R12258 gnd.n265 gnd.n223 242.672
R12259 gnd.n7759 gnd.n223 242.672
R12260 gnd.n258 gnd.n223 242.672
R12261 gnd.n7766 gnd.n223 242.672
R12262 gnd.n251 gnd.n223 242.672
R12263 gnd.n7776 gnd.n223 242.672
R12264 gnd.n244 gnd.n223 242.672
R12265 gnd.n7783 gnd.n223 242.672
R12266 gnd.n237 gnd.n223 242.672
R12267 gnd.n7790 gnd.n223 242.672
R12268 gnd.n230 gnd.n223 242.672
R12269 gnd.n7797 gnd.n223 242.672
R12270 gnd.n223 gnd.n222 242.672
R12271 gnd.n3222 gnd.n3221 242.672
R12272 gnd.n3222 gnd.n2399 242.672
R12273 gnd.n3222 gnd.n2400 242.672
R12274 gnd.n3222 gnd.n2401 242.672
R12275 gnd.n3222 gnd.n2402 242.672
R12276 gnd.n3222 gnd.n2403 242.672
R12277 gnd.n3222 gnd.n2404 242.672
R12278 gnd.n3222 gnd.n2405 242.672
R12279 gnd.n3222 gnd.n2406 242.672
R12280 gnd.n3222 gnd.n2407 242.672
R12281 gnd.n3222 gnd.n2408 242.672
R12282 gnd.n3222 gnd.n2409 242.672
R12283 gnd.n3222 gnd.n2410 242.672
R12284 gnd.n3222 gnd.n2411 242.672
R12285 gnd.n4076 gnd.n1715 242.672
R12286 gnd.n3952 gnd.n1715 242.672
R12287 gnd.n4057 gnd.n1715 242.672
R12288 gnd.n3961 gnd.n1715 242.672
R12289 gnd.n4038 gnd.n1715 242.672
R12290 gnd.n3970 gnd.n1715 242.672
R12291 gnd.n4019 gnd.n1715 242.672
R12292 gnd.n3979 gnd.n1715 242.672
R12293 gnd.n4004 gnd.n1715 242.672
R12294 gnd.n3982 gnd.n1715 242.672
R12295 gnd.n3993 gnd.n1715 242.672
R12296 gnd.n3986 gnd.n1715 242.672
R12297 gnd.n4098 gnd.n1715 242.672
R12298 gnd.n4095 gnd.n1715 242.672
R12299 gnd.n219 gnd.n216 240.244
R12300 gnd.n7799 gnd.n7798 240.244
R12301 gnd.n7796 gnd.n224 240.244
R12302 gnd.n7792 gnd.n7791 240.244
R12303 gnd.n7789 gnd.n231 240.244
R12304 gnd.n7785 gnd.n7784 240.244
R12305 gnd.n7782 gnd.n238 240.244
R12306 gnd.n7778 gnd.n7777 240.244
R12307 gnd.n7775 gnd.n245 240.244
R12308 gnd.n7768 gnd.n7767 240.244
R12309 gnd.n7765 gnd.n252 240.244
R12310 gnd.n7761 gnd.n7760 240.244
R12311 gnd.n7758 gnd.n259 240.244
R12312 gnd.n7754 gnd.n7753 240.244
R12313 gnd.n7751 gnd.n266 240.244
R12314 gnd.n7747 gnd.n7746 240.244
R12315 gnd.n7744 gnd.n273 240.244
R12316 gnd.n7740 gnd.n7739 240.244
R12317 gnd.n7737 gnd.n280 240.244
R12318 gnd.n7730 gnd.n289 240.244
R12319 gnd.n7728 gnd.n7727 240.244
R12320 gnd.n7725 gnd.n291 240.244
R12321 gnd.n7721 gnd.n7720 240.244
R12322 gnd.n7718 gnd.n298 240.244
R12323 gnd.n7714 gnd.n7713 240.244
R12324 gnd.n7711 gnd.n305 240.244
R12325 gnd.n7707 gnd.n7706 240.244
R12326 gnd.n7704 gnd.n312 240.244
R12327 gnd.n7700 gnd.n7699 240.244
R12328 gnd.n1932 gnd.n1725 240.244
R12329 gnd.n1932 gnd.n1737 240.244
R12330 gnd.n4496 gnd.n1737 240.244
R12331 gnd.n4496 gnd.n1749 240.244
R12332 gnd.n4506 gnd.n1749 240.244
R12333 gnd.n4506 gnd.n1760 240.244
R12334 gnd.n4510 gnd.n1760 240.244
R12335 gnd.n4510 gnd.n1769 240.244
R12336 gnd.n4520 gnd.n1769 240.244
R12337 gnd.n4520 gnd.n1780 240.244
R12338 gnd.n1880 gnd.n1780 240.244
R12339 gnd.n1880 gnd.n1789 240.244
R12340 gnd.n4527 gnd.n1789 240.244
R12341 gnd.n4527 gnd.n1800 240.244
R12342 gnd.n4532 gnd.n1800 240.244
R12343 gnd.n4532 gnd.n1809 240.244
R12344 gnd.n4537 gnd.n1809 240.244
R12345 gnd.n4537 gnd.n1820 240.244
R12346 gnd.n4580 gnd.n1820 240.244
R12347 gnd.n4580 gnd.n1829 240.244
R12348 gnd.n4608 gnd.n1829 240.244
R12349 gnd.n4608 gnd.n1838 240.244
R12350 gnd.n1862 gnd.n1838 240.244
R12351 gnd.n1862 gnd.n1847 240.244
R12352 gnd.n1854 gnd.n1847 240.244
R12353 gnd.n4601 gnd.n1854 240.244
R12354 gnd.n4601 gnd.n4600 240.244
R12355 gnd.n4600 gnd.n86 240.244
R12356 gnd.n390 gnd.n86 240.244
R12357 gnd.n7579 gnd.n390 240.244
R12358 gnd.n7579 gnd.n103 240.244
R12359 gnd.n7583 gnd.n103 240.244
R12360 gnd.n7583 gnd.n115 240.244
R12361 gnd.n7593 gnd.n115 240.244
R12362 gnd.n7593 gnd.n124 240.244
R12363 gnd.n7597 gnd.n124 240.244
R12364 gnd.n7597 gnd.n133 240.244
R12365 gnd.n7607 gnd.n133 240.244
R12366 gnd.n7607 gnd.n144 240.244
R12367 gnd.n7611 gnd.n144 240.244
R12368 gnd.n7611 gnd.n154 240.244
R12369 gnd.n7621 gnd.n154 240.244
R12370 gnd.n7621 gnd.n164 240.244
R12371 gnd.n7625 gnd.n164 240.244
R12372 gnd.n7625 gnd.n173 240.244
R12373 gnd.n7635 gnd.n173 240.244
R12374 gnd.n7635 gnd.n184 240.244
R12375 gnd.n7639 gnd.n184 240.244
R12376 gnd.n7639 gnd.n194 240.244
R12377 gnd.n7650 gnd.n194 240.244
R12378 gnd.n7650 gnd.n205 240.244
R12379 gnd.n7655 gnd.n205 240.244
R12380 gnd.n7655 gnd.n213 240.244
R12381 gnd.n4344 gnd.n4343 240.244
R12382 gnd.n4346 gnd.n4344 240.244
R12383 gnd.n4352 gnd.n4334 240.244
R12384 gnd.n4356 gnd.n4354 240.244
R12385 gnd.n4362 gnd.n4330 240.244
R12386 gnd.n4366 gnd.n4364 240.244
R12387 gnd.n4372 gnd.n4326 240.244
R12388 gnd.n4376 gnd.n4374 240.244
R12389 gnd.n4385 gnd.n4322 240.244
R12390 gnd.n4389 gnd.n4387 240.244
R12391 gnd.n4395 gnd.n4318 240.244
R12392 gnd.n4399 gnd.n4397 240.244
R12393 gnd.n4406 gnd.n4314 240.244
R12394 gnd.n4412 gnd.n4410 240.244
R12395 gnd.n4418 gnd.n1963 240.244
R12396 gnd.n4422 gnd.n4420 240.244
R12397 gnd.n4428 gnd.n1959 240.244
R12398 gnd.n4432 gnd.n4430 240.244
R12399 gnd.n4440 gnd.n1955 240.244
R12400 gnd.n4444 gnd.n4442 240.244
R12401 gnd.n4450 gnd.n1951 240.244
R12402 gnd.n4454 gnd.n4452 240.244
R12403 gnd.n4460 gnd.n1947 240.244
R12404 gnd.n4464 gnd.n4462 240.244
R12405 gnd.n4470 gnd.n1943 240.244
R12406 gnd.n4474 gnd.n4472 240.244
R12407 gnd.n4481 gnd.n1939 240.244
R12408 gnd.n4484 gnd.n4483 240.244
R12409 gnd.n4709 gnd.n1730 240.244
R12410 gnd.n4705 gnd.n1730 240.244
R12411 gnd.n4705 gnd.n1735 240.244
R12412 gnd.n4697 gnd.n1735 240.244
R12413 gnd.n4697 gnd.n1752 240.244
R12414 gnd.n4693 gnd.n1752 240.244
R12415 gnd.n4693 gnd.n1758 240.244
R12416 gnd.n4685 gnd.n1758 240.244
R12417 gnd.n4685 gnd.n1772 240.244
R12418 gnd.n4681 gnd.n1772 240.244
R12419 gnd.n4681 gnd.n1778 240.244
R12420 gnd.n4673 gnd.n1778 240.244
R12421 gnd.n4673 gnd.n1792 240.244
R12422 gnd.n4669 gnd.n1792 240.244
R12423 gnd.n4669 gnd.n1798 240.244
R12424 gnd.n4661 gnd.n1798 240.244
R12425 gnd.n4661 gnd.n1812 240.244
R12426 gnd.n4657 gnd.n1812 240.244
R12427 gnd.n4657 gnd.n1818 240.244
R12428 gnd.n4649 gnd.n1818 240.244
R12429 gnd.n4649 gnd.n1832 240.244
R12430 gnd.n4645 gnd.n1832 240.244
R12431 gnd.n4645 gnd.n1836 240.244
R12432 gnd.n4637 gnd.n1836 240.244
R12433 gnd.n4637 gnd.n4636 240.244
R12434 gnd.n4636 gnd.n1852 240.244
R12435 gnd.n1852 gnd.n89 240.244
R12436 gnd.n7880 gnd.n89 240.244
R12437 gnd.n7880 gnd.n90 240.244
R12438 gnd.n100 gnd.n90 240.244
R12439 gnd.n7874 gnd.n100 240.244
R12440 gnd.n7874 gnd.n101 240.244
R12441 gnd.n7866 gnd.n101 240.244
R12442 gnd.n7866 gnd.n117 240.244
R12443 gnd.n7862 gnd.n117 240.244
R12444 gnd.n7862 gnd.n122 240.244
R12445 gnd.n7854 gnd.n122 240.244
R12446 gnd.n7854 gnd.n136 240.244
R12447 gnd.n7850 gnd.n136 240.244
R12448 gnd.n7850 gnd.n142 240.244
R12449 gnd.n7842 gnd.n142 240.244
R12450 gnd.n7842 gnd.n156 240.244
R12451 gnd.n7838 gnd.n156 240.244
R12452 gnd.n7838 gnd.n162 240.244
R12453 gnd.n7830 gnd.n162 240.244
R12454 gnd.n7830 gnd.n176 240.244
R12455 gnd.n7826 gnd.n176 240.244
R12456 gnd.n7826 gnd.n182 240.244
R12457 gnd.n7818 gnd.n182 240.244
R12458 gnd.n7818 gnd.n197 240.244
R12459 gnd.n7814 gnd.n197 240.244
R12460 gnd.n7814 gnd.n203 240.244
R12461 gnd.n7806 gnd.n203 240.244
R12462 gnd.n4959 gnd.n1483 240.244
R12463 gnd.n4957 gnd.n4956 240.244
R12464 gnd.n4954 gnd.n1489 240.244
R12465 gnd.n4950 gnd.n4949 240.244
R12466 gnd.n4947 gnd.n1497 240.244
R12467 gnd.n4943 gnd.n4942 240.244
R12468 gnd.n4940 gnd.n1504 240.244
R12469 gnd.n4936 gnd.n4935 240.244
R12470 gnd.n4933 gnd.n1511 240.244
R12471 gnd.n4928 gnd.n4927 240.244
R12472 gnd.n4925 gnd.n1520 240.244
R12473 gnd.n4921 gnd.n4920 240.244
R12474 gnd.n4918 gnd.n1527 240.244
R12475 gnd.n2457 gnd.n2456 240.244
R12476 gnd.n2460 gnd.n2459 240.244
R12477 gnd.n2467 gnd.n2466 240.244
R12478 gnd.n2470 gnd.n2469 240.244
R12479 gnd.n2477 gnd.n2476 240.244
R12480 gnd.n2480 gnd.n2479 240.244
R12481 gnd.n2487 gnd.n2486 240.244
R12482 gnd.n2490 gnd.n2489 240.244
R12483 gnd.n2497 gnd.n2496 240.244
R12484 gnd.n2500 gnd.n2499 240.244
R12485 gnd.n2507 gnd.n2506 240.244
R12486 gnd.n2510 gnd.n2509 240.244
R12487 gnd.n2517 gnd.n2516 240.244
R12488 gnd.n2520 gnd.n2519 240.244
R12489 gnd.n2527 gnd.n2526 240.244
R12490 gnd.n5104 gnd.n1242 240.244
R12491 gnd.n2779 gnd.n1242 240.244
R12492 gnd.n2779 gnd.n1259 240.244
R12493 gnd.n2789 gnd.n1259 240.244
R12494 gnd.n2789 gnd.n1270 240.244
R12495 gnd.n2794 gnd.n1270 240.244
R12496 gnd.n2794 gnd.n1280 240.244
R12497 gnd.n2847 gnd.n1280 240.244
R12498 gnd.n2847 gnd.n1290 240.244
R12499 gnd.n2852 gnd.n1290 240.244
R12500 gnd.n2852 gnd.n1301 240.244
R12501 gnd.n2863 gnd.n1301 240.244
R12502 gnd.n2863 gnd.n1311 240.244
R12503 gnd.n2701 gnd.n1311 240.244
R12504 gnd.n2701 gnd.n1321 240.244
R12505 gnd.n2894 gnd.n1321 240.244
R12506 gnd.n2894 gnd.n1331 240.244
R12507 gnd.n2890 gnd.n1331 240.244
R12508 gnd.n2890 gnd.n1342 240.244
R12509 gnd.n2882 gnd.n1342 240.244
R12510 gnd.n2882 gnd.n1352 240.244
R12511 gnd.n2689 gnd.n1352 240.244
R12512 gnd.n2935 gnd.n2689 240.244
R12513 gnd.n2935 gnd.n2679 240.244
R12514 gnd.n2679 gnd.n2672 240.244
R12515 gnd.n2960 gnd.n2672 240.244
R12516 gnd.n2960 gnd.n2661 240.244
R12517 gnd.n2963 gnd.n2661 240.244
R12518 gnd.n2963 gnd.n2655 240.244
R12519 gnd.n2655 gnd.n2649 240.244
R12520 gnd.n2649 gnd.n1369 240.244
R12521 gnd.n3016 gnd.n1369 240.244
R12522 gnd.n3016 gnd.n1381 240.244
R12523 gnd.n3021 gnd.n1381 240.244
R12524 gnd.n3021 gnd.n1390 240.244
R12525 gnd.n3031 gnd.n1390 240.244
R12526 gnd.n3031 gnd.n1400 240.244
R12527 gnd.n2629 gnd.n1400 240.244
R12528 gnd.n2629 gnd.n1410 240.244
R12529 gnd.n3038 gnd.n1410 240.244
R12530 gnd.n3038 gnd.n1420 240.244
R12531 gnd.n3044 gnd.n1420 240.244
R12532 gnd.n3044 gnd.n1430 240.244
R12533 gnd.n3048 gnd.n1430 240.244
R12534 gnd.n3048 gnd.n1440 240.244
R12535 gnd.n3119 gnd.n1440 240.244
R12536 gnd.n3119 gnd.n1450 240.244
R12537 gnd.n3123 gnd.n1450 240.244
R12538 gnd.n3123 gnd.n1460 240.244
R12539 gnd.n3134 gnd.n1460 240.244
R12540 gnd.n3134 gnd.n1471 240.244
R12541 gnd.n3139 gnd.n1471 240.244
R12542 gnd.n3139 gnd.n1480 240.244
R12543 gnd.n1171 gnd.n1170 240.244
R12544 gnd.n5219 gnd.n1170 240.244
R12545 gnd.n5217 gnd.n5216 240.244
R12546 gnd.n5213 gnd.n5212 240.244
R12547 gnd.n5209 gnd.n5208 240.244
R12548 gnd.n5205 gnd.n5204 240.244
R12549 gnd.n5201 gnd.n5200 240.244
R12550 gnd.n5197 gnd.n5196 240.244
R12551 gnd.n5193 gnd.n5192 240.244
R12552 gnd.n5188 gnd.n5187 240.244
R12553 gnd.n5184 gnd.n5183 240.244
R12554 gnd.n5180 gnd.n5179 240.244
R12555 gnd.n5176 gnd.n5175 240.244
R12556 gnd.n5172 gnd.n5171 240.244
R12557 gnd.n5168 gnd.n5167 240.244
R12558 gnd.n5164 gnd.n5163 240.244
R12559 gnd.n5160 gnd.n5159 240.244
R12560 gnd.n5156 gnd.n5155 240.244
R12561 gnd.n5152 gnd.n5151 240.244
R12562 gnd.n5148 gnd.n5147 240.244
R12563 gnd.n5144 gnd.n5143 240.244
R12564 gnd.n5140 gnd.n5139 240.244
R12565 gnd.n5136 gnd.n5135 240.244
R12566 gnd.n5132 gnd.n5131 240.244
R12567 gnd.n5128 gnd.n5127 240.244
R12568 gnd.n5124 gnd.n5123 240.244
R12569 gnd.n5120 gnd.n5119 240.244
R12570 gnd.n5116 gnd.n5115 240.244
R12571 gnd.n5112 gnd.n5111 240.244
R12572 gnd.n5099 gnd.n1172 240.244
R12573 gnd.n5099 gnd.n1250 240.244
R12574 gnd.n5095 gnd.n1250 240.244
R12575 gnd.n5095 gnd.n1257 240.244
R12576 gnd.n5087 gnd.n1257 240.244
R12577 gnd.n5087 gnd.n1273 240.244
R12578 gnd.n5083 gnd.n1273 240.244
R12579 gnd.n5083 gnd.n1279 240.244
R12580 gnd.n5075 gnd.n1279 240.244
R12581 gnd.n5075 gnd.n1293 240.244
R12582 gnd.n5071 gnd.n1293 240.244
R12583 gnd.n5071 gnd.n1299 240.244
R12584 gnd.n5063 gnd.n1299 240.244
R12585 gnd.n5063 gnd.n1314 240.244
R12586 gnd.n5059 gnd.n1314 240.244
R12587 gnd.n5059 gnd.n1320 240.244
R12588 gnd.n5051 gnd.n1320 240.244
R12589 gnd.n5051 gnd.n1334 240.244
R12590 gnd.n5047 gnd.n1334 240.244
R12591 gnd.n5047 gnd.n1340 240.244
R12592 gnd.n5039 gnd.n1340 240.244
R12593 gnd.n5039 gnd.n1355 240.244
R12594 gnd.n2682 gnd.n1355 240.244
R12595 gnd.n2944 gnd.n2682 240.244
R12596 gnd.n2944 gnd.n2943 240.244
R12597 gnd.n2943 gnd.n2657 240.244
R12598 gnd.n2973 gnd.n2657 240.244
R12599 gnd.n2974 gnd.n2973 240.244
R12600 gnd.n2977 gnd.n2974 240.244
R12601 gnd.n2977 gnd.n1367 240.244
R12602 gnd.n5033 gnd.n1367 240.244
R12603 gnd.n5033 gnd.n1368 240.244
R12604 gnd.n5025 gnd.n1368 240.244
R12605 gnd.n5025 gnd.n1383 240.244
R12606 gnd.n5021 gnd.n1383 240.244
R12607 gnd.n5021 gnd.n1388 240.244
R12608 gnd.n5013 gnd.n1388 240.244
R12609 gnd.n5013 gnd.n1403 240.244
R12610 gnd.n5009 gnd.n1403 240.244
R12611 gnd.n5009 gnd.n1409 240.244
R12612 gnd.n5001 gnd.n1409 240.244
R12613 gnd.n5001 gnd.n1422 240.244
R12614 gnd.n4997 gnd.n1422 240.244
R12615 gnd.n4997 gnd.n1428 240.244
R12616 gnd.n4989 gnd.n1428 240.244
R12617 gnd.n4989 gnd.n1443 240.244
R12618 gnd.n4985 gnd.n1443 240.244
R12619 gnd.n4985 gnd.n1449 240.244
R12620 gnd.n4977 gnd.n1449 240.244
R12621 gnd.n4977 gnd.n1463 240.244
R12622 gnd.n4973 gnd.n1463 240.244
R12623 gnd.n4973 gnd.n1469 240.244
R12624 gnd.n4965 gnd.n1469 240.244
R12625 gnd.n5243 gnd.n5238 240.244
R12626 gnd.n6570 gnd.n6569 240.244
R12627 gnd.n6567 gnd.n5247 240.244
R12628 gnd.n6563 gnd.n6562 240.244
R12629 gnd.n6560 gnd.n5254 240.244
R12630 gnd.n6556 gnd.n6555 240.244
R12631 gnd.n6553 gnd.n5261 240.244
R12632 gnd.n6549 gnd.n6548 240.244
R12633 gnd.n5884 gnd.n5596 240.244
R12634 gnd.n5894 gnd.n5596 240.244
R12635 gnd.n5894 gnd.n5587 240.244
R12636 gnd.n5587 gnd.n5576 240.244
R12637 gnd.n5915 gnd.n5576 240.244
R12638 gnd.n5915 gnd.n5570 240.244
R12639 gnd.n5925 gnd.n5570 240.244
R12640 gnd.n5925 gnd.n5559 240.244
R12641 gnd.n5559 gnd.n5551 240.244
R12642 gnd.n5943 gnd.n5551 240.244
R12643 gnd.n5944 gnd.n5943 240.244
R12644 gnd.n5944 gnd.n5536 240.244
R12645 gnd.n5946 gnd.n5536 240.244
R12646 gnd.n5946 gnd.n5522 240.244
R12647 gnd.n5988 gnd.n5522 240.244
R12648 gnd.n5989 gnd.n5988 240.244
R12649 gnd.n5992 gnd.n5989 240.244
R12650 gnd.n5992 gnd.n5477 240.244
R12651 gnd.n5517 gnd.n5477 240.244
R12652 gnd.n5517 gnd.n5487 240.244
R12653 gnd.n6002 gnd.n5487 240.244
R12654 gnd.n6002 gnd.n5508 240.244
R12655 gnd.n6012 gnd.n5508 240.244
R12656 gnd.n6012 gnd.n5390 240.244
R12657 gnd.n6057 gnd.n5390 240.244
R12658 gnd.n6057 gnd.n5376 240.244
R12659 gnd.n6079 gnd.n5376 240.244
R12660 gnd.n6080 gnd.n6079 240.244
R12661 gnd.n6080 gnd.n5363 240.244
R12662 gnd.n5363 gnd.n5352 240.244
R12663 gnd.n6111 gnd.n5352 240.244
R12664 gnd.n6112 gnd.n6111 240.244
R12665 gnd.n6113 gnd.n6112 240.244
R12666 gnd.n6113 gnd.n5337 240.244
R12667 gnd.n5337 gnd.n5329 240.244
R12668 gnd.n6166 gnd.n5329 240.244
R12669 gnd.n6167 gnd.n6166 240.244
R12670 gnd.n6167 gnd.n1051 240.244
R12671 gnd.n6144 gnd.n1051 240.244
R12672 gnd.n6144 gnd.n1061 240.244
R12673 gnd.n6179 gnd.n1061 240.244
R12674 gnd.n6180 gnd.n6179 240.244
R12675 gnd.n6180 gnd.n1074 240.244
R12676 gnd.n6469 gnd.n1074 240.244
R12677 gnd.n6469 gnd.n1086 240.244
R12678 gnd.n6465 gnd.n1086 240.244
R12679 gnd.n6465 gnd.n6464 240.244
R12680 gnd.n6464 gnd.n1099 240.244
R12681 gnd.n6460 gnd.n1099 240.244
R12682 gnd.n6460 gnd.n1112 240.244
R12683 gnd.n6456 gnd.n1112 240.244
R12684 gnd.n6456 gnd.n6455 240.244
R12685 gnd.n6455 gnd.n1124 240.244
R12686 gnd.n5874 gnd.n5609 240.244
R12687 gnd.n5630 gnd.n5609 240.244
R12688 gnd.n5633 gnd.n5632 240.244
R12689 gnd.n5640 gnd.n5639 240.244
R12690 gnd.n5643 gnd.n5642 240.244
R12691 gnd.n5650 gnd.n5649 240.244
R12692 gnd.n5653 gnd.n5652 240.244
R12693 gnd.n5660 gnd.n5659 240.244
R12694 gnd.n5882 gnd.n5606 240.244
R12695 gnd.n5606 gnd.n5585 240.244
R12696 gnd.n5905 gnd.n5585 240.244
R12697 gnd.n5905 gnd.n5579 240.244
R12698 gnd.n5913 gnd.n5579 240.244
R12699 gnd.n5913 gnd.n5581 240.244
R12700 gnd.n5581 gnd.n5557 240.244
R12701 gnd.n5935 gnd.n5557 240.244
R12702 gnd.n5935 gnd.n5553 240.244
R12703 gnd.n5941 gnd.n5553 240.244
R12704 gnd.n5941 gnd.n5535 240.244
R12705 gnd.n5966 gnd.n5535 240.244
R12706 gnd.n5966 gnd.n5530 240.244
R12707 gnd.n5978 gnd.n5530 240.244
R12708 gnd.n5978 gnd.n5531 240.244
R12709 gnd.n5974 gnd.n5531 240.244
R12710 gnd.n5974 gnd.n5479 240.244
R12711 gnd.n6026 gnd.n5479 240.244
R12712 gnd.n6026 gnd.n5480 240.244
R12713 gnd.n6022 gnd.n5480 240.244
R12714 gnd.n6022 gnd.n5486 240.244
R12715 gnd.n5506 gnd.n5486 240.244
R12716 gnd.n5506 gnd.n5388 240.244
R12717 gnd.n6061 gnd.n5388 240.244
R12718 gnd.n6061 gnd.n5383 240.244
R12719 gnd.n6069 gnd.n5383 240.244
R12720 gnd.n6069 gnd.n5384 240.244
R12721 gnd.n5384 gnd.n5361 240.244
R12722 gnd.n6101 gnd.n5361 240.244
R12723 gnd.n6101 gnd.n5356 240.244
R12724 gnd.n6109 gnd.n5356 240.244
R12725 gnd.n6109 gnd.n5357 240.244
R12726 gnd.n5357 gnd.n5335 240.244
R12727 gnd.n6157 gnd.n5335 240.244
R12728 gnd.n6157 gnd.n5331 240.244
R12729 gnd.n6164 gnd.n5331 240.244
R12730 gnd.n6164 gnd.n1052 240.244
R12731 gnd.n6619 gnd.n1052 240.244
R12732 gnd.n6619 gnd.n1053 240.244
R12733 gnd.n6615 gnd.n1053 240.244
R12734 gnd.n6615 gnd.n1059 240.244
R12735 gnd.n1075 gnd.n1059 240.244
R12736 gnd.n6605 gnd.n1075 240.244
R12737 gnd.n6605 gnd.n1076 240.244
R12738 gnd.n6601 gnd.n1076 240.244
R12739 gnd.n6601 gnd.n1084 240.244
R12740 gnd.n1101 gnd.n1084 240.244
R12741 gnd.n6591 gnd.n1101 240.244
R12742 gnd.n6591 gnd.n1102 240.244
R12743 gnd.n6587 gnd.n1102 240.244
R12744 gnd.n6587 gnd.n1110 240.244
R12745 gnd.n5237 gnd.n1110 240.244
R12746 gnd.n6577 gnd.n5237 240.244
R12747 gnd.n323 gnd.n211 240.244
R12748 gnd.n7689 gnd.n7688 240.244
R12749 gnd.n7686 gnd.n327 240.244
R12750 gnd.n7682 gnd.n7681 240.244
R12751 gnd.n7679 gnd.n334 240.244
R12752 gnd.n7675 gnd.n7674 240.244
R12753 gnd.n7672 gnd.n341 240.244
R12754 gnd.n7668 gnd.n7667 240.244
R12755 gnd.n7665 gnd.n348 240.244
R12756 gnd.n3926 gnd.n1726 240.244
R12757 gnd.n3926 gnd.n1738 240.244
R12758 gnd.n4498 gnd.n1738 240.244
R12759 gnd.n4498 gnd.n1750 240.244
R12760 gnd.n4504 gnd.n1750 240.244
R12761 gnd.n4504 gnd.n1761 240.244
R12762 gnd.n4512 gnd.n1761 240.244
R12763 gnd.n4512 gnd.n1770 240.244
R12764 gnd.n4518 gnd.n1770 240.244
R12765 gnd.n4518 gnd.n1781 240.244
R12766 gnd.n4554 gnd.n1781 240.244
R12767 gnd.n4554 gnd.n1790 240.244
R12768 gnd.n1885 gnd.n1790 240.244
R12769 gnd.n1885 gnd.n1801 240.244
R12770 gnd.n1886 gnd.n1801 240.244
R12771 gnd.n1886 gnd.n1810 240.244
R12772 gnd.n4539 gnd.n1810 240.244
R12773 gnd.n4539 gnd.n1821 240.244
R12774 gnd.n1868 gnd.n1821 240.244
R12775 gnd.n1868 gnd.n1830 240.244
R12776 gnd.n4610 gnd.n1830 240.244
R12777 gnd.n4610 gnd.n1839 240.244
R12778 gnd.n4619 gnd.n1839 240.244
R12779 gnd.n4619 gnd.n1848 240.244
R12780 gnd.n1855 gnd.n1848 240.244
R12781 gnd.n1856 gnd.n1855 240.244
R12782 gnd.n1856 gnd.n82 240.244
R12783 gnd.n7882 gnd.n82 240.244
R12784 gnd.n7882 gnd.n84 240.244
R12785 gnd.n7577 gnd.n84 240.244
R12786 gnd.n7577 gnd.n104 240.244
R12787 gnd.n7585 gnd.n104 240.244
R12788 gnd.n7585 gnd.n116 240.244
R12789 gnd.n7591 gnd.n116 240.244
R12790 gnd.n7591 gnd.n125 240.244
R12791 gnd.n7599 gnd.n125 240.244
R12792 gnd.n7599 gnd.n134 240.244
R12793 gnd.n7605 gnd.n134 240.244
R12794 gnd.n7605 gnd.n145 240.244
R12795 gnd.n7613 gnd.n145 240.244
R12796 gnd.n7613 gnd.n155 240.244
R12797 gnd.n7619 gnd.n155 240.244
R12798 gnd.n7619 gnd.n165 240.244
R12799 gnd.n7627 gnd.n165 240.244
R12800 gnd.n7627 gnd.n174 240.244
R12801 gnd.n7633 gnd.n174 240.244
R12802 gnd.n7633 gnd.n185 240.244
R12803 gnd.n7641 gnd.n185 240.244
R12804 gnd.n7641 gnd.n195 240.244
R12805 gnd.n7648 gnd.n195 240.244
R12806 gnd.n7648 gnd.n206 240.244
R12807 gnd.n7657 gnd.n206 240.244
R12808 gnd.n7657 gnd.n214 240.244
R12809 gnd.n4026 gnd.n3974 240.244
R12810 gnd.n4030 gnd.n4028 240.244
R12811 gnd.n4045 gnd.n3965 240.244
R12812 gnd.n4049 gnd.n4047 240.244
R12813 gnd.n4064 gnd.n3956 240.244
R12814 gnd.n4068 gnd.n4066 240.244
R12815 gnd.n4084 gnd.n3947 240.244
R12816 gnd.n4088 gnd.n4086 240.244
R12817 gnd.n3943 gnd.n3942 240.244
R12818 gnd.n1740 gnd.n1728 240.244
R12819 gnd.n4703 gnd.n1740 240.244
R12820 gnd.n4703 gnd.n1741 240.244
R12821 gnd.n4699 gnd.n1741 240.244
R12822 gnd.n4699 gnd.n1747 240.244
R12823 gnd.n4691 gnd.n1747 240.244
R12824 gnd.n4691 gnd.n1762 240.244
R12825 gnd.n4687 gnd.n1762 240.244
R12826 gnd.n4687 gnd.n1767 240.244
R12827 gnd.n4679 gnd.n1767 240.244
R12828 gnd.n4679 gnd.n1783 240.244
R12829 gnd.n4675 gnd.n1783 240.244
R12830 gnd.n4675 gnd.n1788 240.244
R12831 gnd.n4667 gnd.n1788 240.244
R12832 gnd.n4667 gnd.n1802 240.244
R12833 gnd.n4663 gnd.n1802 240.244
R12834 gnd.n4663 gnd.n1807 240.244
R12835 gnd.n4655 gnd.n1807 240.244
R12836 gnd.n4655 gnd.n1823 240.244
R12837 gnd.n4651 gnd.n1823 240.244
R12838 gnd.n4651 gnd.n1828 240.244
R12839 gnd.n4643 gnd.n1828 240.244
R12840 gnd.n4643 gnd.n1840 240.244
R12841 gnd.n4639 gnd.n1840 240.244
R12842 gnd.n4639 gnd.n1845 240.244
R12843 gnd.n4588 gnd.n1845 240.244
R12844 gnd.n4598 gnd.n4588 240.244
R12845 gnd.n4598 gnd.n88 240.244
R12846 gnd.n4594 gnd.n88 240.244
R12847 gnd.n4594 gnd.n106 240.244
R12848 gnd.n7872 gnd.n106 240.244
R12849 gnd.n7872 gnd.n107 240.244
R12850 gnd.n7868 gnd.n107 240.244
R12851 gnd.n7868 gnd.n113 240.244
R12852 gnd.n7860 gnd.n113 240.244
R12853 gnd.n7860 gnd.n126 240.244
R12854 gnd.n7856 gnd.n126 240.244
R12855 gnd.n7856 gnd.n131 240.244
R12856 gnd.n7848 gnd.n131 240.244
R12857 gnd.n7848 gnd.n147 240.244
R12858 gnd.n7844 gnd.n147 240.244
R12859 gnd.n7844 gnd.n152 240.244
R12860 gnd.n7836 gnd.n152 240.244
R12861 gnd.n7836 gnd.n166 240.244
R12862 gnd.n7832 gnd.n166 240.244
R12863 gnd.n7832 gnd.n171 240.244
R12864 gnd.n7824 gnd.n171 240.244
R12865 gnd.n7824 gnd.n187 240.244
R12866 gnd.n7820 gnd.n187 240.244
R12867 gnd.n7820 gnd.n192 240.244
R12868 gnd.n7812 gnd.n192 240.244
R12869 gnd.n7812 gnd.n207 240.244
R12870 gnd.n7808 gnd.n207 240.244
R12871 gnd.n5273 gnd.n1121 240.244
R12872 gnd.n6538 gnd.n6537 240.244
R12873 gnd.n6535 gnd.n5277 240.244
R12874 gnd.n6531 gnd.n6530 240.244
R12875 gnd.n6528 gnd.n5284 240.244
R12876 gnd.n6524 gnd.n6523 240.244
R12877 gnd.n6521 gnd.n5291 240.244
R12878 gnd.n6517 gnd.n6516 240.244
R12879 gnd.n6514 gnd.n5298 240.244
R12880 gnd.n6510 gnd.n6509 240.244
R12881 gnd.n6507 gnd.n5305 240.244
R12882 gnd.n6503 gnd.n6502 240.244
R12883 gnd.n6500 gnd.n5315 240.244
R12884 gnd.n5797 gnd.n5694 240.244
R12885 gnd.n5797 gnd.n5687 240.244
R12886 gnd.n5808 gnd.n5687 240.244
R12887 gnd.n5808 gnd.n5683 240.244
R12888 gnd.n5814 gnd.n5683 240.244
R12889 gnd.n5814 gnd.n5675 240.244
R12890 gnd.n5824 gnd.n5675 240.244
R12891 gnd.n5824 gnd.n5670 240.244
R12892 gnd.n5860 gnd.n5670 240.244
R12893 gnd.n5860 gnd.n5671 240.244
R12894 gnd.n5671 gnd.n5618 240.244
R12895 gnd.n5855 gnd.n5618 240.244
R12896 gnd.n5855 gnd.n5854 240.244
R12897 gnd.n5854 gnd.n5597 240.244
R12898 gnd.n5850 gnd.n5597 240.244
R12899 gnd.n5850 gnd.n5588 240.244
R12900 gnd.n5847 gnd.n5588 240.244
R12901 gnd.n5847 gnd.n5846 240.244
R12902 gnd.n5846 gnd.n5571 240.244
R12903 gnd.n5842 gnd.n5571 240.244
R12904 gnd.n5842 gnd.n5560 240.244
R12905 gnd.n5560 gnd.n5541 240.244
R12906 gnd.n5955 gnd.n5541 240.244
R12907 gnd.n5955 gnd.n5537 240.244
R12908 gnd.n5963 gnd.n5537 240.244
R12909 gnd.n5963 gnd.n5528 240.244
R12910 gnd.n5528 gnd.n5464 240.244
R12911 gnd.n6035 gnd.n5464 240.244
R12912 gnd.n6035 gnd.n5465 240.244
R12913 gnd.n5476 gnd.n5465 240.244
R12914 gnd.n5511 gnd.n5476 240.244
R12915 gnd.n5514 gnd.n5511 240.244
R12916 gnd.n5514 gnd.n5488 240.244
R12917 gnd.n5501 gnd.n5488 240.244
R12918 gnd.n5501 gnd.n5498 240.244
R12919 gnd.n5498 gnd.n5391 240.244
R12920 gnd.n6056 gnd.n5391 240.244
R12921 gnd.n6056 gnd.n5381 240.244
R12922 gnd.n6052 gnd.n5381 240.244
R12923 gnd.n6052 gnd.n5375 240.244
R12924 gnd.n6049 gnd.n5375 240.244
R12925 gnd.n6049 gnd.n5364 240.244
R12926 gnd.n6046 gnd.n5364 240.244
R12927 gnd.n6046 gnd.n5342 240.244
R12928 gnd.n6124 gnd.n5342 240.244
R12929 gnd.n6124 gnd.n5338 240.244
R12930 gnd.n6154 gnd.n5338 240.244
R12931 gnd.n6154 gnd.n1040 240.244
R12932 gnd.n6150 gnd.n1040 240.244
R12933 gnd.n6150 gnd.n1050 240.244
R12934 gnd.n6147 gnd.n1050 240.244
R12935 gnd.n6147 gnd.n6143 240.244
R12936 gnd.n6143 gnd.n1062 240.244
R12937 gnd.n6139 gnd.n1062 240.244
R12938 gnd.n6139 gnd.n1073 240.244
R12939 gnd.n6472 gnd.n1073 240.244
R12940 gnd.n6473 gnd.n6472 240.244
R12941 gnd.n6473 gnd.n1087 240.244
R12942 gnd.n6479 gnd.n1087 240.244
R12943 gnd.n6479 gnd.n1098 240.244
R12944 gnd.n6483 gnd.n1098 240.244
R12945 gnd.n6483 gnd.n6482 240.244
R12946 gnd.n6482 gnd.n1113 240.244
R12947 gnd.n6490 gnd.n1113 240.244
R12948 gnd.n6490 gnd.n1123 240.244
R12949 gnd.n5711 gnd.n5710 240.244
R12950 gnd.n5782 gnd.n5710 240.244
R12951 gnd.n5780 gnd.n5779 240.244
R12952 gnd.n5776 gnd.n5775 240.244
R12953 gnd.n5772 gnd.n5771 240.244
R12954 gnd.n5768 gnd.n5767 240.244
R12955 gnd.n5764 gnd.n5763 240.244
R12956 gnd.n5760 gnd.n5759 240.244
R12957 gnd.n5756 gnd.n5755 240.244
R12958 gnd.n5752 gnd.n5751 240.244
R12959 gnd.n5748 gnd.n5747 240.244
R12960 gnd.n5744 gnd.n5743 240.244
R12961 gnd.n5740 gnd.n5698 240.244
R12962 gnd.n5800 gnd.n5692 240.244
R12963 gnd.n5800 gnd.n5688 240.244
R12964 gnd.n5806 gnd.n5688 240.244
R12965 gnd.n5806 gnd.n5681 240.244
R12966 gnd.n5816 gnd.n5681 240.244
R12967 gnd.n5816 gnd.n5677 240.244
R12968 gnd.n5822 gnd.n5677 240.244
R12969 gnd.n5822 gnd.n5668 240.244
R12970 gnd.n5862 gnd.n5668 240.244
R12971 gnd.n5862 gnd.n5619 240.244
R12972 gnd.n5870 gnd.n5619 240.244
R12973 gnd.n5870 gnd.n5620 240.244
R12974 gnd.n5620 gnd.n5598 240.244
R12975 gnd.n5891 gnd.n5598 240.244
R12976 gnd.n5891 gnd.n5590 240.244
R12977 gnd.n5902 gnd.n5590 240.244
R12978 gnd.n5902 gnd.n5591 240.244
R12979 gnd.n5591 gnd.n5572 240.244
R12980 gnd.n5922 gnd.n5572 240.244
R12981 gnd.n5922 gnd.n5562 240.244
R12982 gnd.n5932 gnd.n5562 240.244
R12983 gnd.n5932 gnd.n5543 240.244
R12984 gnd.n5953 gnd.n5543 240.244
R12985 gnd.n5953 gnd.n5545 240.244
R12986 gnd.n5545 gnd.n5526 240.244
R12987 gnd.n5981 gnd.n5526 240.244
R12988 gnd.n5981 gnd.n5468 240.244
R12989 gnd.n6033 gnd.n5468 240.244
R12990 gnd.n6033 gnd.n5469 240.244
R12991 gnd.n6029 gnd.n5469 240.244
R12992 gnd.n6029 gnd.n5475 240.244
R12993 gnd.n5490 gnd.n5475 240.244
R12994 gnd.n6019 gnd.n5490 240.244
R12995 gnd.n6019 gnd.n5491 240.244
R12996 gnd.n6015 gnd.n5491 240.244
R12997 gnd.n6015 gnd.n5497 240.244
R12998 gnd.n5497 gnd.n5380 240.244
R12999 gnd.n6072 gnd.n5380 240.244
R13000 gnd.n6072 gnd.n5373 240.244
R13001 gnd.n6083 gnd.n5373 240.244
R13002 gnd.n6083 gnd.n5366 240.244
R13003 gnd.n6098 gnd.n5366 240.244
R13004 gnd.n6098 gnd.n5367 240.244
R13005 gnd.n5367 gnd.n5345 240.244
R13006 gnd.n6122 gnd.n5345 240.244
R13007 gnd.n6122 gnd.n5346 240.244
R13008 gnd.n5346 gnd.n1041 240.244
R13009 gnd.n6626 gnd.n1041 240.244
R13010 gnd.n6626 gnd.n1042 240.244
R13011 gnd.n6622 gnd.n1042 240.244
R13012 gnd.n6622 gnd.n1048 240.244
R13013 gnd.n1064 gnd.n1048 240.244
R13014 gnd.n6612 gnd.n1064 240.244
R13015 gnd.n6612 gnd.n1065 240.244
R13016 gnd.n6608 gnd.n1065 240.244
R13017 gnd.n6608 gnd.n1071 240.244
R13018 gnd.n1089 gnd.n1071 240.244
R13019 gnd.n6598 gnd.n1089 240.244
R13020 gnd.n6598 gnd.n1090 240.244
R13021 gnd.n6594 gnd.n1090 240.244
R13022 gnd.n6594 gnd.n1096 240.244
R13023 gnd.n1115 gnd.n1096 240.244
R13024 gnd.n6584 gnd.n1115 240.244
R13025 gnd.n6584 gnd.n1116 240.244
R13026 gnd.n6580 gnd.n1116 240.244
R13027 gnd.n2542 gnd.n1478 240.244
R13028 gnd.n2553 gnd.n2544 240.244
R13029 gnd.n2556 gnd.n2555 240.244
R13030 gnd.n2565 gnd.n2564 240.244
R13031 gnd.n2576 gnd.n2567 240.244
R13032 gnd.n2579 gnd.n2578 240.244
R13033 gnd.n2588 gnd.n2587 240.244
R13034 gnd.n2600 gnd.n2590 240.244
R13035 gnd.n2606 gnd.n2602 240.244
R13036 gnd.n1248 gnd.n1243 240.244
R13037 gnd.n2781 gnd.n1248 240.244
R13038 gnd.n2781 gnd.n1260 240.244
R13039 gnd.n2787 gnd.n1260 240.244
R13040 gnd.n2787 gnd.n1271 240.244
R13041 gnd.n2839 gnd.n1271 240.244
R13042 gnd.n2839 gnd.n1281 240.244
R13043 gnd.n2845 gnd.n1281 240.244
R13044 gnd.n2845 gnd.n1291 240.244
R13045 gnd.n2854 gnd.n1291 240.244
R13046 gnd.n2854 gnd.n1302 240.244
R13047 gnd.n2861 gnd.n1302 240.244
R13048 gnd.n2861 gnd.n1312 240.244
R13049 gnd.n2900 gnd.n1312 240.244
R13050 gnd.n2900 gnd.n1322 240.244
R13051 gnd.n2896 gnd.n1322 240.244
R13052 gnd.n2896 gnd.n1332 240.244
R13053 gnd.n2888 gnd.n1332 240.244
R13054 gnd.n2888 gnd.n1343 240.244
R13055 gnd.n2884 gnd.n1343 240.244
R13056 gnd.n2884 gnd.n1353 240.244
R13057 gnd.n2877 gnd.n1353 240.244
R13058 gnd.n2877 gnd.n2677 240.244
R13059 gnd.n2946 gnd.n2677 240.244
R13060 gnd.n2946 gnd.n2673 240.244
R13061 gnd.n2958 gnd.n2673 240.244
R13062 gnd.n2958 gnd.n2662 240.244
R13063 gnd.n2951 gnd.n2662 240.244
R13064 gnd.n2951 gnd.n2647 240.244
R13065 gnd.n3008 gnd.n2647 240.244
R13066 gnd.n3008 gnd.n1370 240.244
R13067 gnd.n3014 gnd.n1370 240.244
R13068 gnd.n3014 gnd.n1382 240.244
R13069 gnd.n3023 gnd.n1382 240.244
R13070 gnd.n3023 gnd.n1391 240.244
R13071 gnd.n3029 gnd.n1391 240.244
R13072 gnd.n3029 gnd.n1401 240.244
R13073 gnd.n3065 gnd.n1401 240.244
R13074 gnd.n3065 gnd.n1411 240.244
R13075 gnd.n2634 gnd.n1411 240.244
R13076 gnd.n2634 gnd.n1421 240.244
R13077 gnd.n2635 gnd.n1421 240.244
R13078 gnd.n2635 gnd.n1431 240.244
R13079 gnd.n3050 gnd.n1431 240.244
R13080 gnd.n3050 gnd.n1441 240.244
R13081 gnd.n2617 gnd.n1441 240.244
R13082 gnd.n2617 gnd.n1451 240.244
R13083 gnd.n3125 gnd.n1451 240.244
R13084 gnd.n3125 gnd.n1461 240.244
R13085 gnd.n3132 gnd.n1461 240.244
R13086 gnd.n3132 gnd.n1472 240.244
R13087 gnd.n3141 gnd.n1472 240.244
R13088 gnd.n3141 gnd.n1481 240.244
R13089 gnd.n2735 gnd.n2734 240.244
R13090 gnd.n2741 gnd.n2740 240.244
R13091 gnd.n2745 gnd.n2744 240.244
R13092 gnd.n2751 gnd.n2750 240.244
R13093 gnd.n2755 gnd.n2754 240.244
R13094 gnd.n2761 gnd.n2760 240.244
R13095 gnd.n2765 gnd.n2764 240.244
R13096 gnd.n2724 gnd.n2723 240.244
R13097 gnd.n2719 gnd.n1168 240.244
R13098 gnd.n5102 gnd.n5101 240.244
R13099 gnd.n5101 gnd.n1246 240.244
R13100 gnd.n5093 gnd.n1246 240.244
R13101 gnd.n5093 gnd.n1262 240.244
R13102 gnd.n5089 gnd.n1262 240.244
R13103 gnd.n5089 gnd.n1268 240.244
R13104 gnd.n5081 gnd.n1268 240.244
R13105 gnd.n5081 gnd.n1283 240.244
R13106 gnd.n5077 gnd.n1283 240.244
R13107 gnd.n5077 gnd.n1288 240.244
R13108 gnd.n5069 gnd.n1288 240.244
R13109 gnd.n5069 gnd.n1304 240.244
R13110 gnd.n5065 gnd.n1304 240.244
R13111 gnd.n5065 gnd.n1309 240.244
R13112 gnd.n5057 gnd.n1309 240.244
R13113 gnd.n5057 gnd.n1324 240.244
R13114 gnd.n5053 gnd.n1324 240.244
R13115 gnd.n5053 gnd.n1329 240.244
R13116 gnd.n5045 gnd.n1329 240.244
R13117 gnd.n5045 gnd.n1345 240.244
R13118 gnd.n5041 gnd.n1345 240.244
R13119 gnd.n5041 gnd.n1350 240.244
R13120 gnd.n2933 gnd.n1350 240.244
R13121 gnd.n2933 gnd.n2681 240.244
R13122 gnd.n2941 gnd.n2681 240.244
R13123 gnd.n2941 gnd.n2664 240.244
R13124 gnd.n2971 gnd.n2664 240.244
R13125 gnd.n2971 gnd.n2665 240.244
R13126 gnd.n2665 gnd.n2656 240.244
R13127 gnd.n2656 gnd.n1372 240.244
R13128 gnd.n5031 gnd.n1372 240.244
R13129 gnd.n5031 gnd.n1373 240.244
R13130 gnd.n5027 gnd.n1373 240.244
R13131 gnd.n5027 gnd.n1379 240.244
R13132 gnd.n5019 gnd.n1379 240.244
R13133 gnd.n5019 gnd.n1393 240.244
R13134 gnd.n5015 gnd.n1393 240.244
R13135 gnd.n5015 gnd.n1398 240.244
R13136 gnd.n5007 gnd.n1398 240.244
R13137 gnd.n5007 gnd.n1413 240.244
R13138 gnd.n5003 gnd.n1413 240.244
R13139 gnd.n5003 gnd.n1418 240.244
R13140 gnd.n4995 gnd.n1418 240.244
R13141 gnd.n4995 gnd.n1433 240.244
R13142 gnd.n4991 gnd.n1433 240.244
R13143 gnd.n4991 gnd.n1438 240.244
R13144 gnd.n4983 gnd.n1438 240.244
R13145 gnd.n4983 gnd.n1453 240.244
R13146 gnd.n4979 gnd.n1453 240.244
R13147 gnd.n4979 gnd.n1458 240.244
R13148 gnd.n4971 gnd.n1458 240.244
R13149 gnd.n4971 gnd.n1474 240.244
R13150 gnd.n4967 gnd.n1474 240.244
R13151 gnd.n6799 gnd.n871 240.244
R13152 gnd.n6799 gnd.n867 240.244
R13153 gnd.n6805 gnd.n867 240.244
R13154 gnd.n6805 gnd.n865 240.244
R13155 gnd.n6809 gnd.n865 240.244
R13156 gnd.n6809 gnd.n861 240.244
R13157 gnd.n6815 gnd.n861 240.244
R13158 gnd.n6815 gnd.n859 240.244
R13159 gnd.n6819 gnd.n859 240.244
R13160 gnd.n6819 gnd.n855 240.244
R13161 gnd.n6825 gnd.n855 240.244
R13162 gnd.n6825 gnd.n853 240.244
R13163 gnd.n6829 gnd.n853 240.244
R13164 gnd.n6829 gnd.n849 240.244
R13165 gnd.n6835 gnd.n849 240.244
R13166 gnd.n6835 gnd.n847 240.244
R13167 gnd.n6839 gnd.n847 240.244
R13168 gnd.n6839 gnd.n843 240.244
R13169 gnd.n6845 gnd.n843 240.244
R13170 gnd.n6845 gnd.n841 240.244
R13171 gnd.n6849 gnd.n841 240.244
R13172 gnd.n6849 gnd.n837 240.244
R13173 gnd.n6855 gnd.n837 240.244
R13174 gnd.n6855 gnd.n835 240.244
R13175 gnd.n6859 gnd.n835 240.244
R13176 gnd.n6859 gnd.n831 240.244
R13177 gnd.n6865 gnd.n831 240.244
R13178 gnd.n6865 gnd.n829 240.244
R13179 gnd.n6869 gnd.n829 240.244
R13180 gnd.n6869 gnd.n825 240.244
R13181 gnd.n6875 gnd.n825 240.244
R13182 gnd.n6875 gnd.n823 240.244
R13183 gnd.n6879 gnd.n823 240.244
R13184 gnd.n6879 gnd.n819 240.244
R13185 gnd.n6885 gnd.n819 240.244
R13186 gnd.n6885 gnd.n817 240.244
R13187 gnd.n6889 gnd.n817 240.244
R13188 gnd.n6889 gnd.n813 240.244
R13189 gnd.n6895 gnd.n813 240.244
R13190 gnd.n6895 gnd.n811 240.244
R13191 gnd.n6899 gnd.n811 240.244
R13192 gnd.n6899 gnd.n807 240.244
R13193 gnd.n6905 gnd.n807 240.244
R13194 gnd.n6905 gnd.n805 240.244
R13195 gnd.n6909 gnd.n805 240.244
R13196 gnd.n6909 gnd.n801 240.244
R13197 gnd.n6915 gnd.n801 240.244
R13198 gnd.n6915 gnd.n799 240.244
R13199 gnd.n6919 gnd.n799 240.244
R13200 gnd.n6919 gnd.n795 240.244
R13201 gnd.n6925 gnd.n795 240.244
R13202 gnd.n6925 gnd.n793 240.244
R13203 gnd.n6929 gnd.n793 240.244
R13204 gnd.n6929 gnd.n789 240.244
R13205 gnd.n6935 gnd.n789 240.244
R13206 gnd.n6935 gnd.n787 240.244
R13207 gnd.n6939 gnd.n787 240.244
R13208 gnd.n6939 gnd.n783 240.244
R13209 gnd.n6945 gnd.n783 240.244
R13210 gnd.n6945 gnd.n781 240.244
R13211 gnd.n6949 gnd.n781 240.244
R13212 gnd.n6949 gnd.n777 240.244
R13213 gnd.n6955 gnd.n777 240.244
R13214 gnd.n6955 gnd.n775 240.244
R13215 gnd.n6959 gnd.n775 240.244
R13216 gnd.n6959 gnd.n771 240.244
R13217 gnd.n6965 gnd.n771 240.244
R13218 gnd.n6965 gnd.n769 240.244
R13219 gnd.n6969 gnd.n769 240.244
R13220 gnd.n6969 gnd.n765 240.244
R13221 gnd.n6975 gnd.n765 240.244
R13222 gnd.n6975 gnd.n763 240.244
R13223 gnd.n6979 gnd.n763 240.244
R13224 gnd.n6979 gnd.n759 240.244
R13225 gnd.n6985 gnd.n759 240.244
R13226 gnd.n6985 gnd.n757 240.244
R13227 gnd.n6989 gnd.n757 240.244
R13228 gnd.n6989 gnd.n753 240.244
R13229 gnd.n6995 gnd.n753 240.244
R13230 gnd.n6995 gnd.n751 240.244
R13231 gnd.n6999 gnd.n751 240.244
R13232 gnd.n6999 gnd.n747 240.244
R13233 gnd.n7005 gnd.n747 240.244
R13234 gnd.n7005 gnd.n745 240.244
R13235 gnd.n7009 gnd.n745 240.244
R13236 gnd.n7009 gnd.n741 240.244
R13237 gnd.n7015 gnd.n741 240.244
R13238 gnd.n7015 gnd.n739 240.244
R13239 gnd.n7019 gnd.n739 240.244
R13240 gnd.n7019 gnd.n735 240.244
R13241 gnd.n7025 gnd.n735 240.244
R13242 gnd.n7025 gnd.n733 240.244
R13243 gnd.n7029 gnd.n733 240.244
R13244 gnd.n7029 gnd.n729 240.244
R13245 gnd.n7035 gnd.n729 240.244
R13246 gnd.n7035 gnd.n727 240.244
R13247 gnd.n7039 gnd.n727 240.244
R13248 gnd.n7039 gnd.n723 240.244
R13249 gnd.n7045 gnd.n723 240.244
R13250 gnd.n7045 gnd.n721 240.244
R13251 gnd.n7049 gnd.n721 240.244
R13252 gnd.n7049 gnd.n717 240.244
R13253 gnd.n7055 gnd.n717 240.244
R13254 gnd.n7055 gnd.n715 240.244
R13255 gnd.n7059 gnd.n715 240.244
R13256 gnd.n7059 gnd.n711 240.244
R13257 gnd.n7065 gnd.n711 240.244
R13258 gnd.n7065 gnd.n709 240.244
R13259 gnd.n7069 gnd.n709 240.244
R13260 gnd.n7069 gnd.n705 240.244
R13261 gnd.n7075 gnd.n705 240.244
R13262 gnd.n7075 gnd.n703 240.244
R13263 gnd.n7079 gnd.n703 240.244
R13264 gnd.n7079 gnd.n699 240.244
R13265 gnd.n7085 gnd.n699 240.244
R13266 gnd.n7085 gnd.n697 240.244
R13267 gnd.n7089 gnd.n697 240.244
R13268 gnd.n7089 gnd.n693 240.244
R13269 gnd.n7095 gnd.n693 240.244
R13270 gnd.n7095 gnd.n691 240.244
R13271 gnd.n7099 gnd.n691 240.244
R13272 gnd.n7099 gnd.n687 240.244
R13273 gnd.n7105 gnd.n687 240.244
R13274 gnd.n7105 gnd.n685 240.244
R13275 gnd.n7109 gnd.n685 240.244
R13276 gnd.n7109 gnd.n681 240.244
R13277 gnd.n7115 gnd.n681 240.244
R13278 gnd.n7115 gnd.n679 240.244
R13279 gnd.n7119 gnd.n679 240.244
R13280 gnd.n7119 gnd.n675 240.244
R13281 gnd.n7125 gnd.n675 240.244
R13282 gnd.n7125 gnd.n673 240.244
R13283 gnd.n7129 gnd.n673 240.244
R13284 gnd.n7129 gnd.n669 240.244
R13285 gnd.n7135 gnd.n669 240.244
R13286 gnd.n7135 gnd.n667 240.244
R13287 gnd.n7139 gnd.n667 240.244
R13288 gnd.n7139 gnd.n663 240.244
R13289 gnd.n7145 gnd.n663 240.244
R13290 gnd.n7145 gnd.n661 240.244
R13291 gnd.n7149 gnd.n661 240.244
R13292 gnd.n7149 gnd.n657 240.244
R13293 gnd.n7155 gnd.n657 240.244
R13294 gnd.n7155 gnd.n655 240.244
R13295 gnd.n7159 gnd.n655 240.244
R13296 gnd.n7159 gnd.n651 240.244
R13297 gnd.n7165 gnd.n651 240.244
R13298 gnd.n7165 gnd.n649 240.244
R13299 gnd.n7169 gnd.n649 240.244
R13300 gnd.n7169 gnd.n645 240.244
R13301 gnd.n7175 gnd.n645 240.244
R13302 gnd.n7175 gnd.n643 240.244
R13303 gnd.n7179 gnd.n643 240.244
R13304 gnd.n7179 gnd.n639 240.244
R13305 gnd.n7185 gnd.n639 240.244
R13306 gnd.n7185 gnd.n637 240.244
R13307 gnd.n7189 gnd.n637 240.244
R13308 gnd.n7189 gnd.n633 240.244
R13309 gnd.n7195 gnd.n633 240.244
R13310 gnd.n7195 gnd.n631 240.244
R13311 gnd.n7199 gnd.n631 240.244
R13312 gnd.n7199 gnd.n627 240.244
R13313 gnd.n7205 gnd.n627 240.244
R13314 gnd.n7205 gnd.n625 240.244
R13315 gnd.n7209 gnd.n625 240.244
R13316 gnd.n7209 gnd.n621 240.244
R13317 gnd.n7215 gnd.n621 240.244
R13318 gnd.n7215 gnd.n619 240.244
R13319 gnd.n7219 gnd.n619 240.244
R13320 gnd.n7219 gnd.n615 240.244
R13321 gnd.n7225 gnd.n615 240.244
R13322 gnd.n7225 gnd.n613 240.244
R13323 gnd.n7229 gnd.n613 240.244
R13324 gnd.n7229 gnd.n609 240.244
R13325 gnd.n7235 gnd.n609 240.244
R13326 gnd.n7235 gnd.n607 240.244
R13327 gnd.n7239 gnd.n607 240.244
R13328 gnd.n7239 gnd.n603 240.244
R13329 gnd.n7245 gnd.n603 240.244
R13330 gnd.n7245 gnd.n601 240.244
R13331 gnd.n7249 gnd.n601 240.244
R13332 gnd.n7249 gnd.n597 240.244
R13333 gnd.n7255 gnd.n597 240.244
R13334 gnd.n7255 gnd.n595 240.244
R13335 gnd.n7259 gnd.n595 240.244
R13336 gnd.n7259 gnd.n591 240.244
R13337 gnd.n7265 gnd.n591 240.244
R13338 gnd.n7265 gnd.n589 240.244
R13339 gnd.n7269 gnd.n589 240.244
R13340 gnd.n7269 gnd.n585 240.244
R13341 gnd.n7275 gnd.n585 240.244
R13342 gnd.n7275 gnd.n583 240.244
R13343 gnd.n7279 gnd.n583 240.244
R13344 gnd.n7279 gnd.n579 240.244
R13345 gnd.n7285 gnd.n579 240.244
R13346 gnd.n7285 gnd.n577 240.244
R13347 gnd.n7289 gnd.n577 240.244
R13348 gnd.n7289 gnd.n573 240.244
R13349 gnd.n7295 gnd.n573 240.244
R13350 gnd.n7295 gnd.n571 240.244
R13351 gnd.n7299 gnd.n571 240.244
R13352 gnd.n7299 gnd.n567 240.244
R13353 gnd.n7305 gnd.n567 240.244
R13354 gnd.n7305 gnd.n565 240.244
R13355 gnd.n7309 gnd.n565 240.244
R13356 gnd.n7309 gnd.n561 240.244
R13357 gnd.n7315 gnd.n561 240.244
R13358 gnd.n7319 gnd.n559 240.244
R13359 gnd.n7319 gnd.n555 240.244
R13360 gnd.n7325 gnd.n555 240.244
R13361 gnd.n7325 gnd.n553 240.244
R13362 gnd.n7329 gnd.n553 240.244
R13363 gnd.n7329 gnd.n549 240.244
R13364 gnd.n7335 gnd.n549 240.244
R13365 gnd.n7335 gnd.n547 240.244
R13366 gnd.n7339 gnd.n547 240.244
R13367 gnd.n7339 gnd.n543 240.244
R13368 gnd.n7345 gnd.n543 240.244
R13369 gnd.n7345 gnd.n541 240.244
R13370 gnd.n7349 gnd.n541 240.244
R13371 gnd.n7349 gnd.n537 240.244
R13372 gnd.n7355 gnd.n537 240.244
R13373 gnd.n7355 gnd.n535 240.244
R13374 gnd.n7359 gnd.n535 240.244
R13375 gnd.n7359 gnd.n531 240.244
R13376 gnd.n7365 gnd.n531 240.244
R13377 gnd.n7365 gnd.n529 240.244
R13378 gnd.n7369 gnd.n529 240.244
R13379 gnd.n7369 gnd.n525 240.244
R13380 gnd.n7375 gnd.n525 240.244
R13381 gnd.n7375 gnd.n523 240.244
R13382 gnd.n7379 gnd.n523 240.244
R13383 gnd.n7379 gnd.n519 240.244
R13384 gnd.n7385 gnd.n519 240.244
R13385 gnd.n7385 gnd.n517 240.244
R13386 gnd.n7389 gnd.n517 240.244
R13387 gnd.n7389 gnd.n513 240.244
R13388 gnd.n7395 gnd.n513 240.244
R13389 gnd.n7395 gnd.n511 240.244
R13390 gnd.n7399 gnd.n511 240.244
R13391 gnd.n7399 gnd.n507 240.244
R13392 gnd.n7405 gnd.n507 240.244
R13393 gnd.n7405 gnd.n505 240.244
R13394 gnd.n7409 gnd.n505 240.244
R13395 gnd.n7409 gnd.n501 240.244
R13396 gnd.n7415 gnd.n501 240.244
R13397 gnd.n7415 gnd.n499 240.244
R13398 gnd.n7419 gnd.n499 240.244
R13399 gnd.n7419 gnd.n495 240.244
R13400 gnd.n7425 gnd.n495 240.244
R13401 gnd.n7425 gnd.n493 240.244
R13402 gnd.n7429 gnd.n493 240.244
R13403 gnd.n7429 gnd.n489 240.244
R13404 gnd.n7435 gnd.n489 240.244
R13405 gnd.n7435 gnd.n487 240.244
R13406 gnd.n7439 gnd.n487 240.244
R13407 gnd.n7439 gnd.n483 240.244
R13408 gnd.n7445 gnd.n483 240.244
R13409 gnd.n7445 gnd.n481 240.244
R13410 gnd.n7449 gnd.n481 240.244
R13411 gnd.n7449 gnd.n477 240.244
R13412 gnd.n7455 gnd.n477 240.244
R13413 gnd.n7455 gnd.n475 240.244
R13414 gnd.n7459 gnd.n475 240.244
R13415 gnd.n7459 gnd.n471 240.244
R13416 gnd.n7465 gnd.n471 240.244
R13417 gnd.n7465 gnd.n469 240.244
R13418 gnd.n7469 gnd.n469 240.244
R13419 gnd.n7469 gnd.n465 240.244
R13420 gnd.n7475 gnd.n465 240.244
R13421 gnd.n7475 gnd.n463 240.244
R13422 gnd.n7479 gnd.n463 240.244
R13423 gnd.n7479 gnd.n459 240.244
R13424 gnd.n7485 gnd.n459 240.244
R13425 gnd.n7485 gnd.n457 240.244
R13426 gnd.n7489 gnd.n457 240.244
R13427 gnd.n7489 gnd.n453 240.244
R13428 gnd.n7495 gnd.n453 240.244
R13429 gnd.n7495 gnd.n451 240.244
R13430 gnd.n7499 gnd.n451 240.244
R13431 gnd.n7499 gnd.n447 240.244
R13432 gnd.n7505 gnd.n447 240.244
R13433 gnd.n7505 gnd.n445 240.244
R13434 gnd.n7509 gnd.n445 240.244
R13435 gnd.n7509 gnd.n441 240.244
R13436 gnd.n7515 gnd.n441 240.244
R13437 gnd.n7515 gnd.n439 240.244
R13438 gnd.n7519 gnd.n439 240.244
R13439 gnd.n7519 gnd.n435 240.244
R13440 gnd.n7527 gnd.n435 240.244
R13441 gnd.n7527 gnd.n432 240.244
R13442 gnd.n5228 gnd.n1126 240.244
R13443 gnd.n5228 gnd.n1130 240.244
R13444 gnd.n2803 gnd.n1130 240.244
R13445 gnd.n2803 gnd.n2800 240.244
R13446 gnd.n2809 gnd.n2800 240.244
R13447 gnd.n2810 gnd.n2809 240.244
R13448 gnd.n2811 gnd.n2810 240.244
R13449 gnd.n2811 gnd.n2795 240.244
R13450 gnd.n2836 gnd.n2795 240.244
R13451 gnd.n2836 gnd.n2796 240.244
R13452 gnd.n2832 gnd.n2796 240.244
R13453 gnd.n2832 gnd.n2831 240.244
R13454 gnd.n2831 gnd.n2830 240.244
R13455 gnd.n2830 gnd.n2819 240.244
R13456 gnd.n2826 gnd.n2819 240.244
R13457 gnd.n2826 gnd.n2700 240.244
R13458 gnd.n2903 gnd.n2700 240.244
R13459 gnd.n2904 gnd.n2903 240.244
R13460 gnd.n2904 gnd.n2696 240.244
R13461 gnd.n2910 gnd.n2696 240.244
R13462 gnd.n2911 gnd.n2910 240.244
R13463 gnd.n2913 gnd.n2911 240.244
R13464 gnd.n2913 gnd.n2912 240.244
R13465 gnd.n2912 gnd.n2691 240.244
R13466 gnd.n2930 gnd.n2691 240.244
R13467 gnd.n2930 gnd.n2692 240.244
R13468 gnd.n2925 gnd.n2692 240.244
R13469 gnd.n2925 gnd.n2924 240.244
R13470 gnd.n2924 gnd.n2920 240.244
R13471 gnd.n2920 gnd.n2653 240.244
R13472 gnd.n2980 gnd.n2653 240.244
R13473 gnd.n2980 gnd.n2650 240.244
R13474 gnd.n3005 gnd.n2650 240.244
R13475 gnd.n3005 gnd.n2651 240.244
R13476 gnd.n3000 gnd.n2651 240.244
R13477 gnd.n3000 gnd.n2999 240.244
R13478 gnd.n2999 gnd.n2998 240.244
R13479 gnd.n2998 gnd.n2986 240.244
R13480 gnd.n2994 gnd.n2986 240.244
R13481 gnd.n2994 gnd.n2627 240.244
R13482 gnd.n3068 gnd.n2627 240.244
R13483 gnd.n3069 gnd.n3068 240.244
R13484 gnd.n3070 gnd.n3069 240.244
R13485 gnd.n3070 gnd.n2623 240.244
R13486 gnd.n3076 gnd.n2623 240.244
R13487 gnd.n3077 gnd.n3076 240.244
R13488 gnd.n3078 gnd.n3077 240.244
R13489 gnd.n3078 gnd.n2618 240.244
R13490 gnd.n3116 gnd.n2618 240.244
R13491 gnd.n3116 gnd.n2619 240.244
R13492 gnd.n3112 gnd.n2619 240.244
R13493 gnd.n3112 gnd.n3111 240.244
R13494 gnd.n3111 gnd.n3110 240.244
R13495 gnd.n3110 gnd.n3086 240.244
R13496 gnd.n3106 gnd.n3086 240.244
R13497 gnd.n3106 gnd.n3105 240.244
R13498 gnd.n3105 gnd.n3104 240.244
R13499 gnd.n3104 gnd.n3092 240.244
R13500 gnd.n3099 gnd.n3092 240.244
R13501 gnd.n3099 gnd.n2397 240.244
R13502 gnd.n3224 gnd.n2397 240.244
R13503 gnd.n3224 gnd.n2391 240.244
R13504 gnd.n3232 gnd.n2391 240.244
R13505 gnd.n3232 gnd.n2393 240.244
R13506 gnd.n2393 gnd.n2373 240.244
R13507 gnd.n3254 gnd.n2373 240.244
R13508 gnd.n3254 gnd.n2368 240.244
R13509 gnd.n3262 gnd.n2368 240.244
R13510 gnd.n3262 gnd.n2369 240.244
R13511 gnd.n2369 gnd.n2348 240.244
R13512 gnd.n3286 gnd.n2348 240.244
R13513 gnd.n3286 gnd.n2343 240.244
R13514 gnd.n3298 gnd.n2343 240.244
R13515 gnd.n3298 gnd.n2344 240.244
R13516 gnd.n3294 gnd.n2344 240.244
R13517 gnd.n3294 gnd.n1600 240.244
R13518 gnd.n4839 gnd.n1600 240.244
R13519 gnd.n4839 gnd.n1601 240.244
R13520 gnd.n4835 gnd.n1601 240.244
R13521 gnd.n4835 gnd.n1607 240.244
R13522 gnd.n2318 gnd.n1607 240.244
R13523 gnd.n3453 gnd.n2318 240.244
R13524 gnd.n3453 gnd.n2313 240.244
R13525 gnd.n3459 gnd.n2313 240.244
R13526 gnd.n3459 gnd.n2295 240.244
R13527 gnd.n3480 gnd.n2295 240.244
R13528 gnd.n3480 gnd.n2290 240.244
R13529 gnd.n3488 gnd.n2290 240.244
R13530 gnd.n3488 gnd.n2291 240.244
R13531 gnd.n2291 gnd.n2262 240.244
R13532 gnd.n3522 gnd.n2262 240.244
R13533 gnd.n3522 gnd.n2257 240.244
R13534 gnd.n3539 gnd.n2257 240.244
R13535 gnd.n3539 gnd.n2258 240.244
R13536 gnd.n3535 gnd.n2258 240.244
R13537 gnd.n3535 gnd.n3531 240.244
R13538 gnd.n3531 gnd.n2228 240.244
R13539 gnd.n3605 gnd.n2228 240.244
R13540 gnd.n3605 gnd.n2224 240.244
R13541 gnd.n3611 gnd.n2224 240.244
R13542 gnd.n3611 gnd.n2205 240.244
R13543 gnd.n3648 gnd.n2205 240.244
R13544 gnd.n3648 gnd.n2201 240.244
R13545 gnd.n3654 gnd.n2201 240.244
R13546 gnd.n3654 gnd.n2189 240.244
R13547 gnd.n3692 gnd.n2189 240.244
R13548 gnd.n3692 gnd.n2184 240.244
R13549 gnd.n3700 gnd.n2184 240.244
R13550 gnd.n3700 gnd.n2185 240.244
R13551 gnd.n2185 gnd.n2158 240.244
R13552 gnd.n3738 gnd.n2158 240.244
R13553 gnd.n3738 gnd.n2154 240.244
R13554 gnd.n3744 gnd.n2154 240.244
R13555 gnd.n3744 gnd.n2141 240.244
R13556 gnd.n3799 gnd.n2141 240.244
R13557 gnd.n3799 gnd.n2137 240.244
R13558 gnd.n3805 gnd.n2137 240.244
R13559 gnd.n3805 gnd.n2119 240.244
R13560 gnd.n3827 gnd.n2119 240.244
R13561 gnd.n3827 gnd.n2114 240.244
R13562 gnd.n3835 gnd.n2114 240.244
R13563 gnd.n3835 gnd.n2115 240.244
R13564 gnd.n2115 gnd.n2091 240.244
R13565 gnd.n3871 gnd.n2091 240.244
R13566 gnd.n3871 gnd.n2086 240.244
R13567 gnd.n3883 gnd.n2086 240.244
R13568 gnd.n3883 gnd.n2087 240.244
R13569 gnd.n3879 gnd.n2087 240.244
R13570 gnd.n3879 gnd.n2018 240.244
R13571 gnd.n4148 gnd.n2018 240.244
R13572 gnd.n4148 gnd.n2019 240.244
R13573 gnd.n4144 gnd.n2019 240.244
R13574 gnd.n4144 gnd.n2025 240.244
R13575 gnd.n4137 gnd.n2025 240.244
R13576 gnd.n4137 gnd.n2029 240.244
R13577 gnd.n4133 gnd.n2029 240.244
R13578 gnd.n4133 gnd.n2035 240.244
R13579 gnd.n4126 gnd.n2035 240.244
R13580 gnd.n4126 gnd.n2040 240.244
R13581 gnd.n4122 gnd.n2040 240.244
R13582 gnd.n4122 gnd.n2046 240.244
R13583 gnd.n4115 gnd.n2046 240.244
R13584 gnd.n4115 gnd.n4108 240.244
R13585 gnd.n4108 gnd.n1707 240.244
R13586 gnd.n4724 gnd.n1707 240.244
R13587 gnd.n4724 gnd.n1708 240.244
R13588 gnd.n4720 gnd.n1708 240.244
R13589 gnd.n4720 gnd.n1714 240.244
R13590 gnd.n4716 gnd.n1714 240.244
R13591 gnd.n4716 gnd.n1717 240.244
R13592 gnd.n4712 gnd.n1717 240.244
R13593 gnd.n4712 gnd.n1723 240.244
R13594 gnd.n1899 gnd.n1723 240.244
R13595 gnd.n1905 gnd.n1899 240.244
R13596 gnd.n1906 gnd.n1905 240.244
R13597 gnd.n1907 gnd.n1906 240.244
R13598 gnd.n1907 gnd.n1894 240.244
R13599 gnd.n1924 gnd.n1894 240.244
R13600 gnd.n1924 gnd.n1895 240.244
R13601 gnd.n1920 gnd.n1895 240.244
R13602 gnd.n1920 gnd.n1919 240.244
R13603 gnd.n1919 gnd.n1878 240.244
R13604 gnd.n4557 gnd.n1878 240.244
R13605 gnd.n4558 gnd.n4557 240.244
R13606 gnd.n4559 gnd.n4558 240.244
R13607 gnd.n4559 gnd.n1874 240.244
R13608 gnd.n4565 gnd.n1874 240.244
R13609 gnd.n4566 gnd.n4565 240.244
R13610 gnd.n4567 gnd.n4566 240.244
R13611 gnd.n4567 gnd.n1869 240.244
R13612 gnd.n4577 gnd.n1869 240.244
R13613 gnd.n4577 gnd.n1870 240.244
R13614 gnd.n1870 gnd.n1861 240.244
R13615 gnd.n4622 gnd.n1861 240.244
R13616 gnd.n4623 gnd.n4622 240.244
R13617 gnd.n4623 gnd.n1858 240.244
R13618 gnd.n4633 gnd.n1858 240.244
R13619 gnd.n4633 gnd.n1859 240.244
R13620 gnd.n4628 gnd.n1859 240.244
R13621 gnd.n4628 gnd.n392 240.244
R13622 gnd.n7572 gnd.n392 240.244
R13623 gnd.n7572 gnd.n393 240.244
R13624 gnd.n7567 gnd.n393 240.244
R13625 gnd.n7567 gnd.n7566 240.244
R13626 gnd.n7566 gnd.n7565 240.244
R13627 gnd.n7565 gnd.n397 240.244
R13628 gnd.n7561 gnd.n397 240.244
R13629 gnd.n7561 gnd.n7560 240.244
R13630 gnd.n7560 gnd.n7559 240.244
R13631 gnd.n7559 gnd.n403 240.244
R13632 gnd.n7555 gnd.n403 240.244
R13633 gnd.n7555 gnd.n7554 240.244
R13634 gnd.n7554 gnd.n7553 240.244
R13635 gnd.n7553 gnd.n409 240.244
R13636 gnd.n7549 gnd.n409 240.244
R13637 gnd.n7549 gnd.n7548 240.244
R13638 gnd.n7548 gnd.n7547 240.244
R13639 gnd.n7547 gnd.n415 240.244
R13640 gnd.n7543 gnd.n415 240.244
R13641 gnd.n7543 gnd.n7542 240.244
R13642 gnd.n7542 gnd.n7541 240.244
R13643 gnd.n7541 gnd.n421 240.244
R13644 gnd.n7537 gnd.n421 240.244
R13645 gnd.n7537 gnd.n7536 240.244
R13646 gnd.n7536 gnd.n7535 240.244
R13647 gnd.n7535 gnd.n427 240.244
R13648 gnd.n7531 gnd.n427 240.244
R13649 gnd.n6795 gnd.n873 240.244
R13650 gnd.n6791 gnd.n873 240.244
R13651 gnd.n6791 gnd.n878 240.244
R13652 gnd.n6787 gnd.n878 240.244
R13653 gnd.n6787 gnd.n880 240.244
R13654 gnd.n6783 gnd.n880 240.244
R13655 gnd.n6783 gnd.n886 240.244
R13656 gnd.n6779 gnd.n886 240.244
R13657 gnd.n6779 gnd.n888 240.244
R13658 gnd.n6775 gnd.n888 240.244
R13659 gnd.n6775 gnd.n894 240.244
R13660 gnd.n6771 gnd.n894 240.244
R13661 gnd.n6771 gnd.n896 240.244
R13662 gnd.n6767 gnd.n896 240.244
R13663 gnd.n6767 gnd.n902 240.244
R13664 gnd.n6763 gnd.n902 240.244
R13665 gnd.n6763 gnd.n904 240.244
R13666 gnd.n6759 gnd.n904 240.244
R13667 gnd.n6759 gnd.n910 240.244
R13668 gnd.n6755 gnd.n910 240.244
R13669 gnd.n6755 gnd.n912 240.244
R13670 gnd.n6751 gnd.n912 240.244
R13671 gnd.n6751 gnd.n918 240.244
R13672 gnd.n6747 gnd.n918 240.244
R13673 gnd.n6747 gnd.n920 240.244
R13674 gnd.n6743 gnd.n920 240.244
R13675 gnd.n6743 gnd.n926 240.244
R13676 gnd.n6739 gnd.n926 240.244
R13677 gnd.n6739 gnd.n928 240.244
R13678 gnd.n6735 gnd.n928 240.244
R13679 gnd.n6735 gnd.n934 240.244
R13680 gnd.n6731 gnd.n934 240.244
R13681 gnd.n6731 gnd.n936 240.244
R13682 gnd.n6727 gnd.n936 240.244
R13683 gnd.n6727 gnd.n942 240.244
R13684 gnd.n6723 gnd.n942 240.244
R13685 gnd.n6723 gnd.n944 240.244
R13686 gnd.n6719 gnd.n944 240.244
R13687 gnd.n6719 gnd.n950 240.244
R13688 gnd.n6715 gnd.n950 240.244
R13689 gnd.n6715 gnd.n952 240.244
R13690 gnd.n6711 gnd.n952 240.244
R13691 gnd.n6711 gnd.n958 240.244
R13692 gnd.n6707 gnd.n958 240.244
R13693 gnd.n6707 gnd.n960 240.244
R13694 gnd.n6703 gnd.n960 240.244
R13695 gnd.n6703 gnd.n966 240.244
R13696 gnd.n6699 gnd.n966 240.244
R13697 gnd.n6699 gnd.n968 240.244
R13698 gnd.n6695 gnd.n968 240.244
R13699 gnd.n6695 gnd.n974 240.244
R13700 gnd.n6691 gnd.n974 240.244
R13701 gnd.n6691 gnd.n976 240.244
R13702 gnd.n6687 gnd.n976 240.244
R13703 gnd.n6687 gnd.n982 240.244
R13704 gnd.n6683 gnd.n982 240.244
R13705 gnd.n6683 gnd.n984 240.244
R13706 gnd.n6679 gnd.n984 240.244
R13707 gnd.n6679 gnd.n990 240.244
R13708 gnd.n6675 gnd.n990 240.244
R13709 gnd.n6675 gnd.n992 240.244
R13710 gnd.n6671 gnd.n992 240.244
R13711 gnd.n6671 gnd.n998 240.244
R13712 gnd.n6667 gnd.n998 240.244
R13713 gnd.n6667 gnd.n1000 240.244
R13714 gnd.n6663 gnd.n1000 240.244
R13715 gnd.n6663 gnd.n1006 240.244
R13716 gnd.n6659 gnd.n1006 240.244
R13717 gnd.n6659 gnd.n1008 240.244
R13718 gnd.n6655 gnd.n1008 240.244
R13719 gnd.n6655 gnd.n1014 240.244
R13720 gnd.n6651 gnd.n1014 240.244
R13721 gnd.n6651 gnd.n1016 240.244
R13722 gnd.n6647 gnd.n1016 240.244
R13723 gnd.n6647 gnd.n1022 240.244
R13724 gnd.n6643 gnd.n1022 240.244
R13725 gnd.n6643 gnd.n1024 240.244
R13726 gnd.n6639 gnd.n1024 240.244
R13727 gnd.n6639 gnd.n1030 240.244
R13728 gnd.n6635 gnd.n1030 240.244
R13729 gnd.n6635 gnd.n1032 240.244
R13730 gnd.n6631 gnd.n1032 240.244
R13731 gnd.n6631 gnd.n1038 240.244
R13732 gnd.n5234 gnd.n1038 240.244
R13733 gnd.n3235 gnd.n2382 240.244
R13734 gnd.n3242 gnd.n2382 240.244
R13735 gnd.n3242 gnd.n2383 240.244
R13736 gnd.n2383 gnd.n2364 240.244
R13737 gnd.n3265 gnd.n2364 240.244
R13738 gnd.n3265 gnd.n2358 240.244
R13739 gnd.n3272 gnd.n2358 240.244
R13740 gnd.n3272 gnd.n2359 240.244
R13741 gnd.n2359 gnd.n2339 240.244
R13742 gnd.n3301 gnd.n2339 240.244
R13743 gnd.n3301 gnd.n2333 240.244
R13744 gnd.n3317 gnd.n2333 240.244
R13745 gnd.n3317 gnd.n2334 240.244
R13746 gnd.n3306 gnd.n2334 240.244
R13747 gnd.n3307 gnd.n3306 240.244
R13748 gnd.n3308 gnd.n3307 240.244
R13749 gnd.n3308 gnd.n1619 240.244
R13750 gnd.n4825 gnd.n1619 240.244
R13751 gnd.n4825 gnd.n1620 240.244
R13752 gnd.n1625 gnd.n1620 240.244
R13753 gnd.n1626 gnd.n1625 240.244
R13754 gnd.n1627 gnd.n1626 240.244
R13755 gnd.n2305 gnd.n1627 240.244
R13756 gnd.n2305 gnd.n1630 240.244
R13757 gnd.n1631 gnd.n1630 240.244
R13758 gnd.n1632 gnd.n1631 240.244
R13759 gnd.n2272 gnd.n1632 240.244
R13760 gnd.n2272 gnd.n1635 240.244
R13761 gnd.n1636 gnd.n1635 240.244
R13762 gnd.n1637 gnd.n1636 240.244
R13763 gnd.n3549 gnd.n1637 240.244
R13764 gnd.n3549 gnd.n1640 240.244
R13765 gnd.n1641 gnd.n1640 240.244
R13766 gnd.n1642 gnd.n1641 240.244
R13767 gnd.n2229 gnd.n1642 240.244
R13768 gnd.n2229 gnd.n1645 240.244
R13769 gnd.n1646 gnd.n1645 240.244
R13770 gnd.n1647 gnd.n1646 240.244
R13771 gnd.n3633 gnd.n1647 240.244
R13772 gnd.n3633 gnd.n1650 240.244
R13773 gnd.n1651 gnd.n1650 240.244
R13774 gnd.n1652 gnd.n1651 240.244
R13775 gnd.n3681 gnd.n1652 240.244
R13776 gnd.n3681 gnd.n1655 240.244
R13777 gnd.n1656 gnd.n1655 240.244
R13778 gnd.n1657 gnd.n1656 240.244
R13779 gnd.n3664 gnd.n1657 240.244
R13780 gnd.n3664 gnd.n1660 240.244
R13781 gnd.n1661 gnd.n1660 240.244
R13782 gnd.n1662 gnd.n1661 240.244
R13783 gnd.n2148 gnd.n1662 240.244
R13784 gnd.n2148 gnd.n1665 240.244
R13785 gnd.n1666 gnd.n1665 240.244
R13786 gnd.n1667 gnd.n1666 240.244
R13787 gnd.n2125 gnd.n1667 240.244
R13788 gnd.n2125 gnd.n1670 240.244
R13789 gnd.n1671 gnd.n1670 240.244
R13790 gnd.n1672 gnd.n1671 240.244
R13791 gnd.n3844 gnd.n1672 240.244
R13792 gnd.n3844 gnd.n1675 240.244
R13793 gnd.n1676 gnd.n1675 240.244
R13794 gnd.n1677 gnd.n1676 240.244
R13795 gnd.n2081 gnd.n1677 240.244
R13796 gnd.n2081 gnd.n1680 240.244
R13797 gnd.n1681 gnd.n1680 240.244
R13798 gnd.n1682 gnd.n1681 240.244
R13799 gnd.n4150 gnd.n1682 240.244
R13800 gnd.n4150 gnd.n1685 240.244
R13801 gnd.n1686 gnd.n1685 240.244
R13802 gnd.n1687 gnd.n1686 240.244
R13803 gnd.n4139 gnd.n1687 240.244
R13804 gnd.n4139 gnd.n1690 240.244
R13805 gnd.n1691 gnd.n1690 240.244
R13806 gnd.n1692 gnd.n1691 240.244
R13807 gnd.n4128 gnd.n1692 240.244
R13808 gnd.n4128 gnd.n1695 240.244
R13809 gnd.n1696 gnd.n1695 240.244
R13810 gnd.n1697 gnd.n1696 240.244
R13811 gnd.n4117 gnd.n1697 240.244
R13812 gnd.n4117 gnd.n1700 240.244
R13813 gnd.n1701 gnd.n1700 240.244
R13814 gnd.n4727 gnd.n1701 240.244
R13815 gnd.n3220 gnd.n2412 240.244
R13816 gnd.n2416 gnd.n2412 240.244
R13817 gnd.n2418 gnd.n2417 240.244
R13818 gnd.n2535 gnd.n2534 240.244
R13819 gnd.n2537 gnd.n2536 240.244
R13820 gnd.n2548 gnd.n2547 240.244
R13821 gnd.n2550 gnd.n2549 240.244
R13822 gnd.n2560 gnd.n2559 240.244
R13823 gnd.n2571 gnd.n2570 240.244
R13824 gnd.n2573 gnd.n2572 240.244
R13825 gnd.n2583 gnd.n2582 240.244
R13826 gnd.n2594 gnd.n2593 240.244
R13827 gnd.n3146 gnd.n2595 240.244
R13828 gnd.n3150 gnd.n3149 240.244
R13829 gnd.n2389 gnd.n2380 240.244
R13830 gnd.n3244 gnd.n2380 240.244
R13831 gnd.n3244 gnd.n2375 240.244
R13832 gnd.n3251 gnd.n2375 240.244
R13833 gnd.n3251 gnd.n2366 240.244
R13834 gnd.n2366 gnd.n2355 240.244
R13835 gnd.n3274 gnd.n2355 240.244
R13836 gnd.n3274 gnd.n2350 240.244
R13837 gnd.n3283 gnd.n2350 240.244
R13838 gnd.n3283 gnd.n2341 240.244
R13839 gnd.n2341 gnd.n2331 240.244
R13840 gnd.n3319 gnd.n2331 240.244
R13841 gnd.n3320 gnd.n3319 240.244
R13842 gnd.n3320 gnd.n2327 240.244
R13843 gnd.n3326 gnd.n2327 240.244
R13844 gnd.n3327 gnd.n3326 240.244
R13845 gnd.n3411 gnd.n3327 240.244
R13846 gnd.n3411 gnd.n1617 240.244
R13847 gnd.n3418 gnd.n1617 240.244
R13848 gnd.n3418 gnd.n2321 240.244
R13849 gnd.n2321 gnd.n2302 240.244
R13850 gnd.n3471 gnd.n2302 240.244
R13851 gnd.n3471 gnd.n2298 240.244
R13852 gnd.n3477 gnd.n2298 240.244
R13853 gnd.n3477 gnd.n2281 240.244
R13854 gnd.n3500 gnd.n2281 240.244
R13855 gnd.n3500 gnd.n2275 240.244
R13856 gnd.n3510 gnd.n2275 240.244
R13857 gnd.n3510 gnd.n2276 240.244
R13858 gnd.n3504 gnd.n2276 240.244
R13859 gnd.n3504 gnd.n2246 240.244
R13860 gnd.n3560 gnd.n2246 240.244
R13861 gnd.n3560 gnd.n2240 240.244
R13862 gnd.n3567 gnd.n2240 240.244
R13863 gnd.n3567 gnd.n2241 240.244
R13864 gnd.n2241 gnd.n2221 240.244
R13865 gnd.n3614 gnd.n2221 240.244
R13866 gnd.n3614 gnd.n2215 240.244
R13867 gnd.n3632 gnd.n2215 240.244
R13868 gnd.n3632 gnd.n2216 240.244
R13869 gnd.n3619 gnd.n2216 240.244
R13870 gnd.n3620 gnd.n3619 240.244
R13871 gnd.n3620 gnd.n2197 240.244
R13872 gnd.n3621 gnd.n2197 240.244
R13873 gnd.n3621 gnd.n2175 240.244
R13874 gnd.n3710 gnd.n2175 240.244
R13875 gnd.n3710 gnd.n2170 240.244
R13876 gnd.n3726 gnd.n2170 240.244
R13877 gnd.n3726 gnd.n2160 240.244
R13878 gnd.n3715 gnd.n2160 240.244
R13879 gnd.n3716 gnd.n3715 240.244
R13880 gnd.n3717 gnd.n3716 240.244
R13881 gnd.n3717 gnd.n2135 240.244
R13882 gnd.n3808 gnd.n2135 240.244
R13883 gnd.n3808 gnd.n2129 240.244
R13884 gnd.n3815 gnd.n2129 240.244
R13885 gnd.n3815 gnd.n2130 240.244
R13886 gnd.n2130 gnd.n2106 240.244
R13887 gnd.n3846 gnd.n2106 240.244
R13888 gnd.n3846 gnd.n2101 240.244
R13889 gnd.n3860 gnd.n2101 240.244
R13890 gnd.n3860 gnd.n2093 240.244
R13891 gnd.n3852 gnd.n2093 240.244
R13892 gnd.n3853 gnd.n3852 240.244
R13893 gnd.n3853 gnd.n2070 240.244
R13894 gnd.n3901 gnd.n2070 240.244
R13895 gnd.n3901 gnd.n2016 240.244
R13896 gnd.n2066 gnd.n2016 240.244
R13897 gnd.n2067 gnd.n2066 240.244
R13898 gnd.n2067 gnd.n2026 240.244
R13899 gnd.n2027 gnd.n2026 240.244
R13900 gnd.n2062 gnd.n2027 240.244
R13901 gnd.n2063 gnd.n2062 240.244
R13902 gnd.n2063 gnd.n2038 240.244
R13903 gnd.n2039 gnd.n2038 240.244
R13904 gnd.n2058 gnd.n2039 240.244
R13905 gnd.n2059 gnd.n2058 240.244
R13906 gnd.n2059 gnd.n2048 240.244
R13907 gnd.n2049 gnd.n2048 240.244
R13908 gnd.n2051 gnd.n2049 240.244
R13909 gnd.n4105 gnd.n2051 240.244
R13910 gnd.n4105 gnd.n1705 240.244
R13911 gnd.n3992 gnd.n3991 240.244
R13912 gnd.n3995 gnd.n3994 240.244
R13913 gnd.n4003 gnd.n4002 240.244
R13914 gnd.n4006 gnd.n4005 240.244
R13915 gnd.n4018 gnd.n4017 240.244
R13916 gnd.n4021 gnd.n4020 240.244
R13917 gnd.n4037 gnd.n4036 240.244
R13918 gnd.n4040 gnd.n4039 240.244
R13919 gnd.n4056 gnd.n4055 240.244
R13920 gnd.n4059 gnd.n4058 240.244
R13921 gnd.n4075 gnd.n4074 240.244
R13922 gnd.n4077 gnd.n3933 240.244
R13923 gnd.n4094 gnd.n3933 240.244
R13924 gnd.n4097 gnd.n4096 240.244
R13925 gnd.n1581 gnd.n1580 240.132
R13926 gnd.n4167 gnd.n4166 240.132
R13927 gnd.n6798 gnd.n6797 225.874
R13928 gnd.n6798 gnd.n866 225.874
R13929 gnd.n6806 gnd.n866 225.874
R13930 gnd.n6807 gnd.n6806 225.874
R13931 gnd.n6808 gnd.n6807 225.874
R13932 gnd.n6808 gnd.n860 225.874
R13933 gnd.n6816 gnd.n860 225.874
R13934 gnd.n6817 gnd.n6816 225.874
R13935 gnd.n6818 gnd.n6817 225.874
R13936 gnd.n6818 gnd.n854 225.874
R13937 gnd.n6826 gnd.n854 225.874
R13938 gnd.n6827 gnd.n6826 225.874
R13939 gnd.n6828 gnd.n6827 225.874
R13940 gnd.n6828 gnd.n848 225.874
R13941 gnd.n6836 gnd.n848 225.874
R13942 gnd.n6837 gnd.n6836 225.874
R13943 gnd.n6838 gnd.n6837 225.874
R13944 gnd.n6838 gnd.n842 225.874
R13945 gnd.n6846 gnd.n842 225.874
R13946 gnd.n6847 gnd.n6846 225.874
R13947 gnd.n6848 gnd.n6847 225.874
R13948 gnd.n6848 gnd.n836 225.874
R13949 gnd.n6856 gnd.n836 225.874
R13950 gnd.n6857 gnd.n6856 225.874
R13951 gnd.n6858 gnd.n6857 225.874
R13952 gnd.n6858 gnd.n830 225.874
R13953 gnd.n6866 gnd.n830 225.874
R13954 gnd.n6867 gnd.n6866 225.874
R13955 gnd.n6868 gnd.n6867 225.874
R13956 gnd.n6868 gnd.n824 225.874
R13957 gnd.n6876 gnd.n824 225.874
R13958 gnd.n6877 gnd.n6876 225.874
R13959 gnd.n6878 gnd.n6877 225.874
R13960 gnd.n6878 gnd.n818 225.874
R13961 gnd.n6886 gnd.n818 225.874
R13962 gnd.n6887 gnd.n6886 225.874
R13963 gnd.n6888 gnd.n6887 225.874
R13964 gnd.n6888 gnd.n812 225.874
R13965 gnd.n6896 gnd.n812 225.874
R13966 gnd.n6897 gnd.n6896 225.874
R13967 gnd.n6898 gnd.n6897 225.874
R13968 gnd.n6898 gnd.n806 225.874
R13969 gnd.n6906 gnd.n806 225.874
R13970 gnd.n6907 gnd.n6906 225.874
R13971 gnd.n6908 gnd.n6907 225.874
R13972 gnd.n6908 gnd.n800 225.874
R13973 gnd.n6916 gnd.n800 225.874
R13974 gnd.n6917 gnd.n6916 225.874
R13975 gnd.n6918 gnd.n6917 225.874
R13976 gnd.n6918 gnd.n794 225.874
R13977 gnd.n6926 gnd.n794 225.874
R13978 gnd.n6927 gnd.n6926 225.874
R13979 gnd.n6928 gnd.n6927 225.874
R13980 gnd.n6928 gnd.n788 225.874
R13981 gnd.n6936 gnd.n788 225.874
R13982 gnd.n6937 gnd.n6936 225.874
R13983 gnd.n6938 gnd.n6937 225.874
R13984 gnd.n6938 gnd.n782 225.874
R13985 gnd.n6946 gnd.n782 225.874
R13986 gnd.n6947 gnd.n6946 225.874
R13987 gnd.n6948 gnd.n6947 225.874
R13988 gnd.n6948 gnd.n776 225.874
R13989 gnd.n6956 gnd.n776 225.874
R13990 gnd.n6957 gnd.n6956 225.874
R13991 gnd.n6958 gnd.n6957 225.874
R13992 gnd.n6958 gnd.n770 225.874
R13993 gnd.n6966 gnd.n770 225.874
R13994 gnd.n6967 gnd.n6966 225.874
R13995 gnd.n6968 gnd.n6967 225.874
R13996 gnd.n6968 gnd.n764 225.874
R13997 gnd.n6976 gnd.n764 225.874
R13998 gnd.n6977 gnd.n6976 225.874
R13999 gnd.n6978 gnd.n6977 225.874
R14000 gnd.n6978 gnd.n758 225.874
R14001 gnd.n6986 gnd.n758 225.874
R14002 gnd.n6987 gnd.n6986 225.874
R14003 gnd.n6988 gnd.n6987 225.874
R14004 gnd.n6988 gnd.n752 225.874
R14005 gnd.n6996 gnd.n752 225.874
R14006 gnd.n6997 gnd.n6996 225.874
R14007 gnd.n6998 gnd.n6997 225.874
R14008 gnd.n6998 gnd.n746 225.874
R14009 gnd.n7006 gnd.n746 225.874
R14010 gnd.n7007 gnd.n7006 225.874
R14011 gnd.n7008 gnd.n7007 225.874
R14012 gnd.n7008 gnd.n740 225.874
R14013 gnd.n7016 gnd.n740 225.874
R14014 gnd.n7017 gnd.n7016 225.874
R14015 gnd.n7018 gnd.n7017 225.874
R14016 gnd.n7018 gnd.n734 225.874
R14017 gnd.n7026 gnd.n734 225.874
R14018 gnd.n7027 gnd.n7026 225.874
R14019 gnd.n7028 gnd.n7027 225.874
R14020 gnd.n7028 gnd.n728 225.874
R14021 gnd.n7036 gnd.n728 225.874
R14022 gnd.n7037 gnd.n7036 225.874
R14023 gnd.n7038 gnd.n7037 225.874
R14024 gnd.n7038 gnd.n722 225.874
R14025 gnd.n7046 gnd.n722 225.874
R14026 gnd.n7047 gnd.n7046 225.874
R14027 gnd.n7048 gnd.n7047 225.874
R14028 gnd.n7048 gnd.n716 225.874
R14029 gnd.n7056 gnd.n716 225.874
R14030 gnd.n7057 gnd.n7056 225.874
R14031 gnd.n7058 gnd.n7057 225.874
R14032 gnd.n7058 gnd.n710 225.874
R14033 gnd.n7066 gnd.n710 225.874
R14034 gnd.n7067 gnd.n7066 225.874
R14035 gnd.n7068 gnd.n7067 225.874
R14036 gnd.n7068 gnd.n704 225.874
R14037 gnd.n7076 gnd.n704 225.874
R14038 gnd.n7077 gnd.n7076 225.874
R14039 gnd.n7078 gnd.n7077 225.874
R14040 gnd.n7078 gnd.n698 225.874
R14041 gnd.n7086 gnd.n698 225.874
R14042 gnd.n7087 gnd.n7086 225.874
R14043 gnd.n7088 gnd.n7087 225.874
R14044 gnd.n7088 gnd.n692 225.874
R14045 gnd.n7096 gnd.n692 225.874
R14046 gnd.n7097 gnd.n7096 225.874
R14047 gnd.n7098 gnd.n7097 225.874
R14048 gnd.n7098 gnd.n686 225.874
R14049 gnd.n7106 gnd.n686 225.874
R14050 gnd.n7107 gnd.n7106 225.874
R14051 gnd.n7108 gnd.n7107 225.874
R14052 gnd.n7108 gnd.n680 225.874
R14053 gnd.n7116 gnd.n680 225.874
R14054 gnd.n7117 gnd.n7116 225.874
R14055 gnd.n7118 gnd.n7117 225.874
R14056 gnd.n7118 gnd.n674 225.874
R14057 gnd.n7126 gnd.n674 225.874
R14058 gnd.n7127 gnd.n7126 225.874
R14059 gnd.n7128 gnd.n7127 225.874
R14060 gnd.n7128 gnd.n668 225.874
R14061 gnd.n7136 gnd.n668 225.874
R14062 gnd.n7137 gnd.n7136 225.874
R14063 gnd.n7138 gnd.n7137 225.874
R14064 gnd.n7138 gnd.n662 225.874
R14065 gnd.n7146 gnd.n662 225.874
R14066 gnd.n7147 gnd.n7146 225.874
R14067 gnd.n7148 gnd.n7147 225.874
R14068 gnd.n7148 gnd.n656 225.874
R14069 gnd.n7156 gnd.n656 225.874
R14070 gnd.n7157 gnd.n7156 225.874
R14071 gnd.n7158 gnd.n7157 225.874
R14072 gnd.n7158 gnd.n650 225.874
R14073 gnd.n7166 gnd.n650 225.874
R14074 gnd.n7167 gnd.n7166 225.874
R14075 gnd.n7168 gnd.n7167 225.874
R14076 gnd.n7168 gnd.n644 225.874
R14077 gnd.n7176 gnd.n644 225.874
R14078 gnd.n7177 gnd.n7176 225.874
R14079 gnd.n7178 gnd.n7177 225.874
R14080 gnd.n7178 gnd.n638 225.874
R14081 gnd.n7186 gnd.n638 225.874
R14082 gnd.n7187 gnd.n7186 225.874
R14083 gnd.n7188 gnd.n7187 225.874
R14084 gnd.n7188 gnd.n632 225.874
R14085 gnd.n7196 gnd.n632 225.874
R14086 gnd.n7197 gnd.n7196 225.874
R14087 gnd.n7198 gnd.n7197 225.874
R14088 gnd.n7198 gnd.n626 225.874
R14089 gnd.n7206 gnd.n626 225.874
R14090 gnd.n7207 gnd.n7206 225.874
R14091 gnd.n7208 gnd.n7207 225.874
R14092 gnd.n7208 gnd.n620 225.874
R14093 gnd.n7216 gnd.n620 225.874
R14094 gnd.n7217 gnd.n7216 225.874
R14095 gnd.n7218 gnd.n7217 225.874
R14096 gnd.n7218 gnd.n614 225.874
R14097 gnd.n7226 gnd.n614 225.874
R14098 gnd.n7227 gnd.n7226 225.874
R14099 gnd.n7228 gnd.n7227 225.874
R14100 gnd.n7228 gnd.n608 225.874
R14101 gnd.n7236 gnd.n608 225.874
R14102 gnd.n7237 gnd.n7236 225.874
R14103 gnd.n7238 gnd.n7237 225.874
R14104 gnd.n7238 gnd.n602 225.874
R14105 gnd.n7246 gnd.n602 225.874
R14106 gnd.n7247 gnd.n7246 225.874
R14107 gnd.n7248 gnd.n7247 225.874
R14108 gnd.n7248 gnd.n596 225.874
R14109 gnd.n7256 gnd.n596 225.874
R14110 gnd.n7257 gnd.n7256 225.874
R14111 gnd.n7258 gnd.n7257 225.874
R14112 gnd.n7258 gnd.n590 225.874
R14113 gnd.n7266 gnd.n590 225.874
R14114 gnd.n7267 gnd.n7266 225.874
R14115 gnd.n7268 gnd.n7267 225.874
R14116 gnd.n7268 gnd.n584 225.874
R14117 gnd.n7276 gnd.n584 225.874
R14118 gnd.n7277 gnd.n7276 225.874
R14119 gnd.n7278 gnd.n7277 225.874
R14120 gnd.n7278 gnd.n578 225.874
R14121 gnd.n7286 gnd.n578 225.874
R14122 gnd.n7287 gnd.n7286 225.874
R14123 gnd.n7288 gnd.n7287 225.874
R14124 gnd.n7288 gnd.n572 225.874
R14125 gnd.n7296 gnd.n572 225.874
R14126 gnd.n7297 gnd.n7296 225.874
R14127 gnd.n7298 gnd.n7297 225.874
R14128 gnd.n7298 gnd.n566 225.874
R14129 gnd.n7306 gnd.n566 225.874
R14130 gnd.n7307 gnd.n7306 225.874
R14131 gnd.n7308 gnd.n7307 225.874
R14132 gnd.n7308 gnd.n560 225.874
R14133 gnd.n7316 gnd.n560 225.874
R14134 gnd.n5735 gnd.t15 224.174
R14135 gnd.n5310 gnd.t7 224.174
R14136 gnd.n4408 gnd.n4407 199.319
R14137 gnd.n4409 gnd.n4408 199.319
R14138 gnd.n1533 gnd.n1532 199.319
R14139 gnd.n2455 gnd.n1533 199.319
R14140 gnd.n1582 gnd.n1579 186.49
R14141 gnd.n4168 gnd.n4165 186.49
R14142 gnd.n6440 gnd.n6439 185
R14143 gnd.n6438 gnd.n6437 185
R14144 gnd.n6417 gnd.n6416 185
R14145 gnd.n6432 gnd.n6431 185
R14146 gnd.n6430 gnd.n6429 185
R14147 gnd.n6421 gnd.n6420 185
R14148 gnd.n6424 gnd.n6423 185
R14149 gnd.n6408 gnd.n6407 185
R14150 gnd.n6406 gnd.n6405 185
R14151 gnd.n6385 gnd.n6384 185
R14152 gnd.n6400 gnd.n6399 185
R14153 gnd.n6398 gnd.n6397 185
R14154 gnd.n6389 gnd.n6388 185
R14155 gnd.n6392 gnd.n6391 185
R14156 gnd.n6376 gnd.n6375 185
R14157 gnd.n6374 gnd.n6373 185
R14158 gnd.n6353 gnd.n6352 185
R14159 gnd.n6368 gnd.n6367 185
R14160 gnd.n6366 gnd.n6365 185
R14161 gnd.n6357 gnd.n6356 185
R14162 gnd.n6360 gnd.n6359 185
R14163 gnd.n6345 gnd.n6344 185
R14164 gnd.n6343 gnd.n6342 185
R14165 gnd.n6322 gnd.n6321 185
R14166 gnd.n6337 gnd.n6336 185
R14167 gnd.n6335 gnd.n6334 185
R14168 gnd.n6326 gnd.n6325 185
R14169 gnd.n6329 gnd.n6328 185
R14170 gnd.n6313 gnd.n6312 185
R14171 gnd.n6311 gnd.n6310 185
R14172 gnd.n6290 gnd.n6289 185
R14173 gnd.n6305 gnd.n6304 185
R14174 gnd.n6303 gnd.n6302 185
R14175 gnd.n6294 gnd.n6293 185
R14176 gnd.n6297 gnd.n6296 185
R14177 gnd.n6281 gnd.n6280 185
R14178 gnd.n6279 gnd.n6278 185
R14179 gnd.n6258 gnd.n6257 185
R14180 gnd.n6273 gnd.n6272 185
R14181 gnd.n6271 gnd.n6270 185
R14182 gnd.n6262 gnd.n6261 185
R14183 gnd.n6265 gnd.n6264 185
R14184 gnd.n6249 gnd.n6248 185
R14185 gnd.n6247 gnd.n6246 185
R14186 gnd.n6226 gnd.n6225 185
R14187 gnd.n6241 gnd.n6240 185
R14188 gnd.n6239 gnd.n6238 185
R14189 gnd.n6230 gnd.n6229 185
R14190 gnd.n6233 gnd.n6232 185
R14191 gnd.n6218 gnd.n6217 185
R14192 gnd.n6216 gnd.n6215 185
R14193 gnd.n6195 gnd.n6194 185
R14194 gnd.n6210 gnd.n6209 185
R14195 gnd.n6208 gnd.n6207 185
R14196 gnd.n6199 gnd.n6198 185
R14197 gnd.n6202 gnd.n6201 185
R14198 gnd.n5736 gnd.t14 178.987
R14199 gnd.n5311 gnd.t8 178.987
R14200 gnd.n1 gnd.t298 170.774
R14201 gnd.n7 gnd.t356 170.103
R14202 gnd.n6 gnd.t323 170.103
R14203 gnd.n5 gnd.t332 170.103
R14204 gnd.n4 gnd.t313 170.103
R14205 gnd.n3 gnd.t344 170.103
R14206 gnd.n2 gnd.t352 170.103
R14207 gnd.n1 gnd.t127 170.103
R14208 gnd.n4236 gnd.n4235 163.367
R14209 gnd.n4232 gnd.n4231 163.367
R14210 gnd.n4228 gnd.n4227 163.367
R14211 gnd.n4224 gnd.n4223 163.367
R14212 gnd.n4220 gnd.n4219 163.367
R14213 gnd.n4216 gnd.n4215 163.367
R14214 gnd.n4212 gnd.n4211 163.367
R14215 gnd.n4208 gnd.n4207 163.367
R14216 gnd.n4204 gnd.n4203 163.367
R14217 gnd.n4200 gnd.n4199 163.367
R14218 gnd.n4196 gnd.n4195 163.367
R14219 gnd.n4192 gnd.n4191 163.367
R14220 gnd.n4188 gnd.n4187 163.367
R14221 gnd.n4184 gnd.n4183 163.367
R14222 gnd.n4179 gnd.n4178 163.367
R14223 gnd.n4311 gnd.n1970 163.367
R14224 gnd.n4308 gnd.n4307 163.367
R14225 gnd.n4305 gnd.n2003 163.367
R14226 gnd.n4300 gnd.n4299 163.367
R14227 gnd.n4296 gnd.n4295 163.367
R14228 gnd.n4292 gnd.n4291 163.367
R14229 gnd.n4288 gnd.n4287 163.367
R14230 gnd.n4284 gnd.n4283 163.367
R14231 gnd.n4280 gnd.n4279 163.367
R14232 gnd.n4276 gnd.n4275 163.367
R14233 gnd.n4272 gnd.n4271 163.367
R14234 gnd.n4268 gnd.n4267 163.367
R14235 gnd.n4264 gnd.n4263 163.367
R14236 gnd.n4260 gnd.n4259 163.367
R14237 gnd.n4256 gnd.n4255 163.367
R14238 gnd.n4252 gnd.n4251 163.367
R14239 gnd.n4248 gnd.n4247 163.367
R14240 gnd.n3395 gnd.n1598 163.367
R14241 gnd.n3399 gnd.n1598 163.367
R14242 gnd.n3403 gnd.n3399 163.367
R14243 gnd.n3403 gnd.n1609 163.367
R14244 gnd.n3408 gnd.n1609 163.367
R14245 gnd.n3408 gnd.n1616 163.367
R14246 gnd.n3421 gnd.n1616 163.367
R14247 gnd.n3422 gnd.n3421 163.367
R14248 gnd.n3422 gnd.n2320 163.367
R14249 gnd.n3443 gnd.n2320 163.367
R14250 gnd.n3443 gnd.n2312 163.367
R14251 gnd.n3439 gnd.n2312 163.367
R14252 gnd.n3439 gnd.n2304 163.367
R14253 gnd.n3436 gnd.n2304 163.367
R14254 gnd.n3436 gnd.n2297 163.367
R14255 gnd.n2297 gnd.n2288 163.367
R14256 gnd.n2289 gnd.n2288 163.367
R14257 gnd.n2289 gnd.n2282 163.367
R14258 gnd.n3430 gnd.n2282 163.367
R14259 gnd.n3430 gnd.n2274 163.367
R14260 gnd.n3426 gnd.n2274 163.367
R14261 gnd.n3426 gnd.n2264 163.367
R14262 gnd.n2264 gnd.n2255 163.367
R14263 gnd.n3542 gnd.n2255 163.367
R14264 gnd.n3542 gnd.n2253 163.367
R14265 gnd.n3547 gnd.n2253 163.367
R14266 gnd.n3547 gnd.n2248 163.367
R14267 gnd.n2248 gnd.n2238 163.367
R14268 gnd.n3570 gnd.n2238 163.367
R14269 gnd.n3570 gnd.n2236 163.367
R14270 gnd.n3591 gnd.n2236 163.367
R14271 gnd.n3591 gnd.n2231 163.367
R14272 gnd.n3587 gnd.n2231 163.367
R14273 gnd.n3587 gnd.n3583 163.367
R14274 gnd.n3583 gnd.n3582 163.367
R14275 gnd.n3582 gnd.n2213 163.367
R14276 gnd.n2214 gnd.n2213 163.367
R14277 gnd.n2214 gnd.n2206 163.367
R14278 gnd.n3576 gnd.n2206 163.367
R14279 gnd.n3576 gnd.n2199 163.367
R14280 gnd.n3657 gnd.n2199 163.367
R14281 gnd.n3657 gnd.n2196 163.367
R14282 gnd.n3679 gnd.n2196 163.367
R14283 gnd.n3679 gnd.n2190 163.367
R14284 gnd.n3675 gnd.n2190 163.367
R14285 gnd.n3675 gnd.n2183 163.367
R14286 gnd.n3670 gnd.n2183 163.367
R14287 gnd.n3670 gnd.n2177 163.367
R14288 gnd.n3667 gnd.n2177 163.367
R14289 gnd.n3667 gnd.n2169 163.367
R14290 gnd.n3661 gnd.n2169 163.367
R14291 gnd.n3661 gnd.n2161 163.367
R14292 gnd.n2161 gnd.n2152 163.367
R14293 gnd.n3747 gnd.n2152 163.367
R14294 gnd.n3747 gnd.n2150 163.367
R14295 gnd.n3785 gnd.n2150 163.367
R14296 gnd.n3785 gnd.n2143 163.367
R14297 gnd.n3781 gnd.n2143 163.367
R14298 gnd.n3781 gnd.n3777 163.367
R14299 gnd.n3777 gnd.n3776 163.367
R14300 gnd.n3776 gnd.n2127 163.367
R14301 gnd.n2128 gnd.n2127 163.367
R14302 gnd.n2128 gnd.n2120 163.367
R14303 gnd.n3769 gnd.n2120 163.367
R14304 gnd.n3769 gnd.n2113 163.367
R14305 gnd.n3764 gnd.n2113 163.367
R14306 gnd.n3764 gnd.n2108 163.367
R14307 gnd.n3761 gnd.n2108 163.367
R14308 gnd.n3761 gnd.n2100 163.367
R14309 gnd.n3756 gnd.n2100 163.367
R14310 gnd.n3756 gnd.n2094 163.367
R14311 gnd.n3753 gnd.n2094 163.367
R14312 gnd.n3753 gnd.n2083 163.367
R14313 gnd.n2083 gnd.n2074 163.367
R14314 gnd.n3893 gnd.n2074 163.367
R14315 gnd.n3893 gnd.n2072 163.367
R14316 gnd.n3899 gnd.n2072 163.367
R14317 gnd.n3899 gnd.n2015 163.367
R14318 gnd.n2015 gnd.n2007 163.367
R14319 gnd.n4243 gnd.n2007 163.367
R14320 gnd.n1573 gnd.n1572 163.367
R14321 gnd.n4904 gnd.n1572 163.367
R14322 gnd.n4902 gnd.n4901 163.367
R14323 gnd.n4898 gnd.n4897 163.367
R14324 gnd.n4894 gnd.n4893 163.367
R14325 gnd.n4890 gnd.n4889 163.367
R14326 gnd.n4886 gnd.n4885 163.367
R14327 gnd.n4882 gnd.n4881 163.367
R14328 gnd.n4878 gnd.n4877 163.367
R14329 gnd.n4874 gnd.n4873 163.367
R14330 gnd.n4870 gnd.n4869 163.367
R14331 gnd.n4866 gnd.n4865 163.367
R14332 gnd.n4862 gnd.n4861 163.367
R14333 gnd.n4858 gnd.n4857 163.367
R14334 gnd.n4854 gnd.n4853 163.367
R14335 gnd.n4850 gnd.n4849 163.367
R14336 gnd.n4913 gnd.n1538 163.367
R14337 gnd.n3332 gnd.n3331 163.367
R14338 gnd.n3337 gnd.n3336 163.367
R14339 gnd.n3341 gnd.n3340 163.367
R14340 gnd.n3345 gnd.n3344 163.367
R14341 gnd.n3349 gnd.n3348 163.367
R14342 gnd.n3353 gnd.n3352 163.367
R14343 gnd.n3357 gnd.n3356 163.367
R14344 gnd.n3361 gnd.n3360 163.367
R14345 gnd.n3365 gnd.n3364 163.367
R14346 gnd.n3369 gnd.n3368 163.367
R14347 gnd.n3373 gnd.n3372 163.367
R14348 gnd.n3377 gnd.n3376 163.367
R14349 gnd.n3381 gnd.n3380 163.367
R14350 gnd.n3385 gnd.n3384 163.367
R14351 gnd.n3389 gnd.n3388 163.367
R14352 gnd.n4842 gnd.n1574 163.367
R14353 gnd.n4842 gnd.n1596 163.367
R14354 gnd.n1610 gnd.n1596 163.367
R14355 gnd.n4832 gnd.n1610 163.367
R14356 gnd.n4832 gnd.n1611 163.367
R14357 gnd.n4828 gnd.n1611 163.367
R14358 gnd.n4828 gnd.n1614 163.367
R14359 gnd.n3447 gnd.n1614 163.367
R14360 gnd.n3450 gnd.n3447 163.367
R14361 gnd.n3450 gnd.n2310 163.367
R14362 gnd.n3462 gnd.n2310 163.367
R14363 gnd.n3462 gnd.n2307 163.367
R14364 gnd.n3467 gnd.n2307 163.367
R14365 gnd.n3467 gnd.n2308 163.367
R14366 gnd.n2308 gnd.n2286 163.367
R14367 gnd.n3493 gnd.n2286 163.367
R14368 gnd.n3493 gnd.n2284 163.367
R14369 gnd.n3497 gnd.n2284 163.367
R14370 gnd.n3497 gnd.n2271 163.367
R14371 gnd.n3514 gnd.n2271 163.367
R14372 gnd.n3514 gnd.n2266 163.367
R14373 gnd.n3519 gnd.n2266 163.367
R14374 gnd.n3519 gnd.n2269 163.367
R14375 gnd.n2269 gnd.n2252 163.367
R14376 gnd.n3552 gnd.n2252 163.367
R14377 gnd.n3552 gnd.n2249 163.367
R14378 gnd.n3557 gnd.n2249 163.367
R14379 gnd.n3557 gnd.n2250 163.367
R14380 gnd.n2250 gnd.n2235 163.367
R14381 gnd.n3595 gnd.n2235 163.367
R14382 gnd.n3595 gnd.n2232 163.367
R14383 gnd.n3602 gnd.n2232 163.367
R14384 gnd.n3602 gnd.n2233 163.367
R14385 gnd.n3598 gnd.n2233 163.367
R14386 gnd.n3598 gnd.n2211 163.367
R14387 gnd.n3638 gnd.n2211 163.367
R14388 gnd.n3638 gnd.n2208 163.367
R14389 gnd.n3645 gnd.n2208 163.367
R14390 gnd.n3645 gnd.n2209 163.367
R14391 gnd.n3641 gnd.n2209 163.367
R14392 gnd.n3641 gnd.n2194 163.367
R14393 gnd.n3685 gnd.n2194 163.367
R14394 gnd.n3685 gnd.n2192 163.367
R14395 gnd.n3689 gnd.n2192 163.367
R14396 gnd.n3689 gnd.n2181 163.367
R14397 gnd.n3703 gnd.n2181 163.367
R14398 gnd.n3703 gnd.n2179 163.367
R14399 gnd.n3707 gnd.n2179 163.367
R14400 gnd.n3707 gnd.n2167 163.367
R14401 gnd.n3729 gnd.n2167 163.367
R14402 gnd.n3729 gnd.n2163 163.367
R14403 gnd.n3734 gnd.n2163 163.367
R14404 gnd.n3734 gnd.n2165 163.367
R14405 gnd.n2165 gnd.n2147 163.367
R14406 gnd.n3789 gnd.n2147 163.367
R14407 gnd.n3789 gnd.n2144 163.367
R14408 gnd.n3796 gnd.n2144 163.367
R14409 gnd.n3796 gnd.n2145 163.367
R14410 gnd.n3792 gnd.n2145 163.367
R14411 gnd.n3792 gnd.n2124 163.367
R14412 gnd.n3820 gnd.n2124 163.367
R14413 gnd.n3820 gnd.n2122 163.367
R14414 gnd.n3824 gnd.n2122 163.367
R14415 gnd.n3824 gnd.n2112 163.367
R14416 gnd.n3838 gnd.n2112 163.367
R14417 gnd.n3838 gnd.n2110 163.367
R14418 gnd.n3842 gnd.n2110 163.367
R14419 gnd.n3842 gnd.n2098 163.367
R14420 gnd.n3863 gnd.n2098 163.367
R14421 gnd.n3863 gnd.n2096 163.367
R14422 gnd.n3867 gnd.n2096 163.367
R14423 gnd.n3867 gnd.n2080 163.367
R14424 gnd.n3886 gnd.n2080 163.367
R14425 gnd.n3886 gnd.n2076 163.367
R14426 gnd.n3891 gnd.n2076 163.367
R14427 gnd.n3891 gnd.n2078 163.367
R14428 gnd.n2078 gnd.n2013 163.367
R14429 gnd.n4153 gnd.n2013 163.367
R14430 gnd.n4153 gnd.n2010 163.367
R14431 gnd.n4241 gnd.n2010 163.367
R14432 gnd.n4174 gnd.n4173 156.462
R14433 gnd.n6380 gnd.n6348 153.042
R14434 gnd.n6444 gnd.n6443 152.079
R14435 gnd.n6412 gnd.n6411 152.079
R14436 gnd.n6380 gnd.n6379 152.079
R14437 gnd.n1587 gnd.n1586 152
R14438 gnd.n1588 gnd.n1577 152
R14439 gnd.n1590 gnd.n1589 152
R14440 gnd.n1592 gnd.n1575 152
R14441 gnd.n1594 gnd.n1593 152
R14442 gnd.n4172 gnd.n4156 152
R14443 gnd.n4164 gnd.n4157 152
R14444 gnd.n4163 gnd.n4162 152
R14445 gnd.n4161 gnd.n4158 152
R14446 gnd.n4159 gnd.t49 150.546
R14447 gnd.t364 gnd.n6422 147.661
R14448 gnd.t360 gnd.n6390 147.661
R14449 gnd.t318 gnd.n6358 147.661
R14450 gnd.t338 gnd.n6327 147.661
R14451 gnd.t342 gnd.n6295 147.661
R14452 gnd.t349 gnd.n6263 147.661
R14453 gnd.t340 gnd.n6231 147.661
R14454 gnd.t347 gnd.n6200 147.661
R14455 gnd.n4310 gnd.n1969 143.351
R14456 gnd.n1554 gnd.n1537 143.351
R14457 gnd.n4912 gnd.n1537 143.351
R14458 gnd.n1584 gnd.t97 130.484
R14459 gnd.n1593 gnd.t16 126.766
R14460 gnd.n1591 gnd.t91 126.766
R14461 gnd.n1577 gnd.t116 126.766
R14462 gnd.n1585 gnd.t56 126.766
R14463 gnd.n4160 gnd.t113 126.766
R14464 gnd.n4162 gnd.t59 126.766
R14465 gnd.n4171 gnd.t9 126.766
R14466 gnd.n4173 gnd.t82 126.766
R14467 gnd.n4313 gnd.n4312 112.192
R14468 gnd.n4915 gnd.n4914 112.192
R14469 gnd.n6439 gnd.n6438 104.615
R14470 gnd.n6438 gnd.n6416 104.615
R14471 gnd.n6431 gnd.n6416 104.615
R14472 gnd.n6431 gnd.n6430 104.615
R14473 gnd.n6430 gnd.n6420 104.615
R14474 gnd.n6423 gnd.n6420 104.615
R14475 gnd.n6407 gnd.n6406 104.615
R14476 gnd.n6406 gnd.n6384 104.615
R14477 gnd.n6399 gnd.n6384 104.615
R14478 gnd.n6399 gnd.n6398 104.615
R14479 gnd.n6398 gnd.n6388 104.615
R14480 gnd.n6391 gnd.n6388 104.615
R14481 gnd.n6375 gnd.n6374 104.615
R14482 gnd.n6374 gnd.n6352 104.615
R14483 gnd.n6367 gnd.n6352 104.615
R14484 gnd.n6367 gnd.n6366 104.615
R14485 gnd.n6366 gnd.n6356 104.615
R14486 gnd.n6359 gnd.n6356 104.615
R14487 gnd.n6344 gnd.n6343 104.615
R14488 gnd.n6343 gnd.n6321 104.615
R14489 gnd.n6336 gnd.n6321 104.615
R14490 gnd.n6336 gnd.n6335 104.615
R14491 gnd.n6335 gnd.n6325 104.615
R14492 gnd.n6328 gnd.n6325 104.615
R14493 gnd.n6312 gnd.n6311 104.615
R14494 gnd.n6311 gnd.n6289 104.615
R14495 gnd.n6304 gnd.n6289 104.615
R14496 gnd.n6304 gnd.n6303 104.615
R14497 gnd.n6303 gnd.n6293 104.615
R14498 gnd.n6296 gnd.n6293 104.615
R14499 gnd.n6280 gnd.n6279 104.615
R14500 gnd.n6279 gnd.n6257 104.615
R14501 gnd.n6272 gnd.n6257 104.615
R14502 gnd.n6272 gnd.n6271 104.615
R14503 gnd.n6271 gnd.n6261 104.615
R14504 gnd.n6264 gnd.n6261 104.615
R14505 gnd.n6248 gnd.n6247 104.615
R14506 gnd.n6247 gnd.n6225 104.615
R14507 gnd.n6240 gnd.n6225 104.615
R14508 gnd.n6240 gnd.n6239 104.615
R14509 gnd.n6239 gnd.n6229 104.615
R14510 gnd.n6232 gnd.n6229 104.615
R14511 gnd.n6217 gnd.n6216 104.615
R14512 gnd.n6216 gnd.n6194 104.615
R14513 gnd.n6209 gnd.n6194 104.615
R14514 gnd.n6209 gnd.n6208 104.615
R14515 gnd.n6208 gnd.n6198 104.615
R14516 gnd.n6201 gnd.n6198 104.615
R14517 gnd.n5661 gnd.t78 100.632
R14518 gnd.n5266 gnd.t105 100.632
R14519 gnd.n7799 gnd.n222 99.6594
R14520 gnd.n7797 gnd.n7796 99.6594
R14521 gnd.n7792 gnd.n230 99.6594
R14522 gnd.n7790 gnd.n7789 99.6594
R14523 gnd.n7785 gnd.n237 99.6594
R14524 gnd.n7783 gnd.n7782 99.6594
R14525 gnd.n7778 gnd.n244 99.6594
R14526 gnd.n7776 gnd.n7775 99.6594
R14527 gnd.n7768 gnd.n251 99.6594
R14528 gnd.n7766 gnd.n7765 99.6594
R14529 gnd.n7761 gnd.n258 99.6594
R14530 gnd.n7759 gnd.n7758 99.6594
R14531 gnd.n7754 gnd.n265 99.6594
R14532 gnd.n7752 gnd.n7751 99.6594
R14533 gnd.n7747 gnd.n272 99.6594
R14534 gnd.n7745 gnd.n7744 99.6594
R14535 gnd.n7740 gnd.n279 99.6594
R14536 gnd.n7738 gnd.n7737 99.6594
R14537 gnd.n289 gnd.n288 99.6594
R14538 gnd.n7729 gnd.n7728 99.6594
R14539 gnd.n7726 gnd.n7725 99.6594
R14540 gnd.n7721 gnd.n297 99.6594
R14541 gnd.n7719 gnd.n7718 99.6594
R14542 gnd.n7714 gnd.n304 99.6594
R14543 gnd.n7712 gnd.n7711 99.6594
R14544 gnd.n7707 gnd.n311 99.6594
R14545 gnd.n7705 gnd.n7704 99.6594
R14546 gnd.n7700 gnd.n320 99.6594
R14547 gnd.n7698 gnd.n7697 99.6594
R14548 gnd.n4342 gnd.n1729 99.6594
R14549 gnd.n4346 gnd.n4345 99.6594
R14550 gnd.n4353 gnd.n4352 99.6594
R14551 gnd.n4356 gnd.n4355 99.6594
R14552 gnd.n4363 gnd.n4362 99.6594
R14553 gnd.n4366 gnd.n4365 99.6594
R14554 gnd.n4373 gnd.n4372 99.6594
R14555 gnd.n4376 gnd.n4375 99.6594
R14556 gnd.n4386 gnd.n4385 99.6594
R14557 gnd.n4389 gnd.n4388 99.6594
R14558 gnd.n4396 gnd.n4395 99.6594
R14559 gnd.n4399 gnd.n4398 99.6594
R14560 gnd.n4407 gnd.n4406 99.6594
R14561 gnd.n4412 gnd.n4411 99.6594
R14562 gnd.n4419 gnd.n4418 99.6594
R14563 gnd.n4422 gnd.n4421 99.6594
R14564 gnd.n4429 gnd.n4428 99.6594
R14565 gnd.n4432 gnd.n4431 99.6594
R14566 gnd.n4441 gnd.n4440 99.6594
R14567 gnd.n4444 gnd.n4443 99.6594
R14568 gnd.n4451 gnd.n4450 99.6594
R14569 gnd.n4454 gnd.n4453 99.6594
R14570 gnd.n4461 gnd.n4460 99.6594
R14571 gnd.n4464 gnd.n4463 99.6594
R14572 gnd.n4471 gnd.n4470 99.6594
R14573 gnd.n4474 gnd.n4473 99.6594
R14574 gnd.n4482 gnd.n4481 99.6594
R14575 gnd.n4485 gnd.n4484 99.6594
R14576 gnd.n4958 gnd.n4957 99.6594
R14577 gnd.n4955 gnd.n4954 99.6594
R14578 gnd.n4950 gnd.n1496 99.6594
R14579 gnd.n4948 gnd.n4947 99.6594
R14580 gnd.n4943 gnd.n1503 99.6594
R14581 gnd.n4941 gnd.n4940 99.6594
R14582 gnd.n4936 gnd.n1510 99.6594
R14583 gnd.n4934 gnd.n4933 99.6594
R14584 gnd.n4928 gnd.n1519 99.6594
R14585 gnd.n4926 gnd.n4925 99.6594
R14586 gnd.n4921 gnd.n1526 99.6594
R14587 gnd.n4919 gnd.n4918 99.6594
R14588 gnd.n2456 gnd.n2455 99.6594
R14589 gnd.n2460 gnd.n2458 99.6594
R14590 gnd.n2466 gnd.n2450 99.6594
R14591 gnd.n2470 gnd.n2468 99.6594
R14592 gnd.n2476 gnd.n2446 99.6594
R14593 gnd.n2480 gnd.n2478 99.6594
R14594 gnd.n2486 gnd.n2440 99.6594
R14595 gnd.n2490 gnd.n2488 99.6594
R14596 gnd.n2496 gnd.n2436 99.6594
R14597 gnd.n2500 gnd.n2498 99.6594
R14598 gnd.n2506 gnd.n2432 99.6594
R14599 gnd.n2510 gnd.n2508 99.6594
R14600 gnd.n2516 gnd.n2428 99.6594
R14601 gnd.n2520 gnd.n2518 99.6594
R14602 gnd.n2526 gnd.n2424 99.6594
R14603 gnd.n2529 gnd.n2528 99.6594
R14604 gnd.n5225 gnd.n5224 99.6594
R14605 gnd.n5219 gnd.n1131 99.6594
R14606 gnd.n5216 gnd.n1132 99.6594
R14607 gnd.n5212 gnd.n1133 99.6594
R14608 gnd.n5208 gnd.n1134 99.6594
R14609 gnd.n5204 gnd.n1135 99.6594
R14610 gnd.n5200 gnd.n1136 99.6594
R14611 gnd.n5196 gnd.n1137 99.6594
R14612 gnd.n5192 gnd.n1138 99.6594
R14613 gnd.n5187 gnd.n1139 99.6594
R14614 gnd.n5183 gnd.n1140 99.6594
R14615 gnd.n5179 gnd.n1141 99.6594
R14616 gnd.n5175 gnd.n1142 99.6594
R14617 gnd.n5171 gnd.n1143 99.6594
R14618 gnd.n5167 gnd.n1144 99.6594
R14619 gnd.n5163 gnd.n1145 99.6594
R14620 gnd.n5159 gnd.n1146 99.6594
R14621 gnd.n5155 gnd.n1147 99.6594
R14622 gnd.n5151 gnd.n1148 99.6594
R14623 gnd.n5147 gnd.n1149 99.6594
R14624 gnd.n5143 gnd.n1150 99.6594
R14625 gnd.n5139 gnd.n1151 99.6594
R14626 gnd.n5135 gnd.n1152 99.6594
R14627 gnd.n5131 gnd.n1153 99.6594
R14628 gnd.n5127 gnd.n1154 99.6594
R14629 gnd.n5123 gnd.n1155 99.6594
R14630 gnd.n5119 gnd.n1156 99.6594
R14631 gnd.n5115 gnd.n1157 99.6594
R14632 gnd.n5111 gnd.n1158 99.6594
R14633 gnd.n6570 gnd.n5246 99.6594
R14634 gnd.n6568 gnd.n6567 99.6594
R14635 gnd.n6563 gnd.n5253 99.6594
R14636 gnd.n6561 gnd.n6560 99.6594
R14637 gnd.n6556 gnd.n5260 99.6594
R14638 gnd.n6554 gnd.n6553 99.6594
R14639 gnd.n6549 gnd.n5269 99.6594
R14640 gnd.n6547 gnd.n6546 99.6594
R14641 gnd.n5873 gnd.n5604 99.6594
R14642 gnd.n5630 gnd.n5611 99.6594
R14643 gnd.n5632 gnd.n5612 99.6594
R14644 gnd.n5640 gnd.n5613 99.6594
R14645 gnd.n5642 gnd.n5614 99.6594
R14646 gnd.n5650 gnd.n5615 99.6594
R14647 gnd.n5652 gnd.n5616 99.6594
R14648 gnd.n5660 gnd.n5617 99.6594
R14649 gnd.n7689 gnd.n326 99.6594
R14650 gnd.n7687 gnd.n7686 99.6594
R14651 gnd.n7682 gnd.n333 99.6594
R14652 gnd.n7680 gnd.n7679 99.6594
R14653 gnd.n7675 gnd.n340 99.6594
R14654 gnd.n7673 gnd.n7672 99.6594
R14655 gnd.n7668 gnd.n347 99.6594
R14656 gnd.n7666 gnd.n7665 99.6594
R14657 gnd.n352 gnd.n351 99.6594
R14658 gnd.n4011 gnd.n4010 99.6594
R14659 gnd.n4027 gnd.n4026 99.6594
R14660 gnd.n4030 gnd.n4029 99.6594
R14661 gnd.n4046 gnd.n4045 99.6594
R14662 gnd.n4049 gnd.n4048 99.6594
R14663 gnd.n4065 gnd.n4064 99.6594
R14664 gnd.n4068 gnd.n4067 99.6594
R14665 gnd.n4085 gnd.n4084 99.6594
R14666 gnd.n4088 gnd.n4087 99.6594
R14667 gnd.n6538 gnd.n5276 99.6594
R14668 gnd.n6536 gnd.n6535 99.6594
R14669 gnd.n6531 gnd.n5283 99.6594
R14670 gnd.n6529 gnd.n6528 99.6594
R14671 gnd.n6524 gnd.n5290 99.6594
R14672 gnd.n6522 gnd.n6521 99.6594
R14673 gnd.n6517 gnd.n5297 99.6594
R14674 gnd.n6515 gnd.n6514 99.6594
R14675 gnd.n6510 gnd.n5304 99.6594
R14676 gnd.n6508 gnd.n6507 99.6594
R14677 gnd.n6503 gnd.n5313 99.6594
R14678 gnd.n6501 gnd.n6500 99.6594
R14679 gnd.n6496 gnd.n6495 99.6594
R14680 gnd.n5788 gnd.n5787 99.6594
R14681 gnd.n5782 gnd.n5699 99.6594
R14682 gnd.n5779 gnd.n5700 99.6594
R14683 gnd.n5775 gnd.n5701 99.6594
R14684 gnd.n5771 gnd.n5702 99.6594
R14685 gnd.n5767 gnd.n5703 99.6594
R14686 gnd.n5763 gnd.n5704 99.6594
R14687 gnd.n5759 gnd.n5705 99.6594
R14688 gnd.n5755 gnd.n5706 99.6594
R14689 gnd.n5751 gnd.n5707 99.6594
R14690 gnd.n5747 gnd.n5708 99.6594
R14691 gnd.n5743 gnd.n5709 99.6594
R14692 gnd.n5790 gnd.n5698 99.6594
R14693 gnd.n2544 gnd.n2543 99.6594
R14694 gnd.n2555 gnd.n2554 99.6594
R14695 gnd.n2564 gnd.n2563 99.6594
R14696 gnd.n2567 gnd.n2566 99.6594
R14697 gnd.n2578 gnd.n2577 99.6594
R14698 gnd.n2587 gnd.n2586 99.6594
R14699 gnd.n2590 gnd.n2589 99.6594
R14700 gnd.n2602 gnd.n2601 99.6594
R14701 gnd.n3160 gnd.n3159 99.6594
R14702 gnd.n1245 gnd.n1159 99.6594
R14703 gnd.n2735 gnd.n1160 99.6594
R14704 gnd.n2741 gnd.n1161 99.6594
R14705 gnd.n2745 gnd.n1162 99.6594
R14706 gnd.n2751 gnd.n1163 99.6594
R14707 gnd.n2755 gnd.n1164 99.6594
R14708 gnd.n2761 gnd.n1165 99.6594
R14709 gnd.n2765 gnd.n1166 99.6594
R14710 gnd.n2724 gnd.n1167 99.6594
R14711 gnd.n2734 gnd.n1159 99.6594
R14712 gnd.n2740 gnd.n1160 99.6594
R14713 gnd.n2744 gnd.n1161 99.6594
R14714 gnd.n2750 gnd.n1162 99.6594
R14715 gnd.n2754 gnd.n1163 99.6594
R14716 gnd.n2760 gnd.n1164 99.6594
R14717 gnd.n2764 gnd.n1165 99.6594
R14718 gnd.n2723 gnd.n1166 99.6594
R14719 gnd.n2719 gnd.n1167 99.6594
R14720 gnd.n3159 gnd.n2606 99.6594
R14721 gnd.n2601 gnd.n2600 99.6594
R14722 gnd.n2589 gnd.n2588 99.6594
R14723 gnd.n2586 gnd.n2579 99.6594
R14724 gnd.n2577 gnd.n2576 99.6594
R14725 gnd.n2566 gnd.n2565 99.6594
R14726 gnd.n2563 gnd.n2556 99.6594
R14727 gnd.n2554 gnd.n2553 99.6594
R14728 gnd.n2543 gnd.n2542 99.6594
R14729 gnd.n5788 gnd.n5711 99.6594
R14730 gnd.n5780 gnd.n5699 99.6594
R14731 gnd.n5776 gnd.n5700 99.6594
R14732 gnd.n5772 gnd.n5701 99.6594
R14733 gnd.n5768 gnd.n5702 99.6594
R14734 gnd.n5764 gnd.n5703 99.6594
R14735 gnd.n5760 gnd.n5704 99.6594
R14736 gnd.n5756 gnd.n5705 99.6594
R14737 gnd.n5752 gnd.n5706 99.6594
R14738 gnd.n5748 gnd.n5707 99.6594
R14739 gnd.n5744 gnd.n5708 99.6594
R14740 gnd.n5740 gnd.n5709 99.6594
R14741 gnd.n5791 gnd.n5790 99.6594
R14742 gnd.n6495 gnd.n5315 99.6594
R14743 gnd.n6502 gnd.n6501 99.6594
R14744 gnd.n5313 gnd.n5305 99.6594
R14745 gnd.n6509 gnd.n6508 99.6594
R14746 gnd.n5304 gnd.n5298 99.6594
R14747 gnd.n6516 gnd.n6515 99.6594
R14748 gnd.n5297 gnd.n5291 99.6594
R14749 gnd.n6523 gnd.n6522 99.6594
R14750 gnd.n5290 gnd.n5284 99.6594
R14751 gnd.n6530 gnd.n6529 99.6594
R14752 gnd.n5283 gnd.n5277 99.6594
R14753 gnd.n6537 gnd.n6536 99.6594
R14754 gnd.n5276 gnd.n5273 99.6594
R14755 gnd.n4010 gnd.n3974 99.6594
R14756 gnd.n4028 gnd.n4027 99.6594
R14757 gnd.n4029 gnd.n3965 99.6594
R14758 gnd.n4047 gnd.n4046 99.6594
R14759 gnd.n4048 gnd.n3956 99.6594
R14760 gnd.n4066 gnd.n4065 99.6594
R14761 gnd.n4067 gnd.n3947 99.6594
R14762 gnd.n4086 gnd.n4085 99.6594
R14763 gnd.n4087 gnd.n3943 99.6594
R14764 gnd.n351 gnd.n348 99.6594
R14765 gnd.n7667 gnd.n7666 99.6594
R14766 gnd.n347 gnd.n341 99.6594
R14767 gnd.n7674 gnd.n7673 99.6594
R14768 gnd.n340 gnd.n334 99.6594
R14769 gnd.n7681 gnd.n7680 99.6594
R14770 gnd.n333 gnd.n327 99.6594
R14771 gnd.n7688 gnd.n7687 99.6594
R14772 gnd.n326 gnd.n323 99.6594
R14773 gnd.n5874 gnd.n5873 99.6594
R14774 gnd.n5633 gnd.n5611 99.6594
R14775 gnd.n5639 gnd.n5612 99.6594
R14776 gnd.n5643 gnd.n5613 99.6594
R14777 gnd.n5649 gnd.n5614 99.6594
R14778 gnd.n5653 gnd.n5615 99.6594
R14779 gnd.n5659 gnd.n5616 99.6594
R14780 gnd.n5617 gnd.n5601 99.6594
R14781 gnd.n6548 gnd.n6547 99.6594
R14782 gnd.n5269 gnd.n5261 99.6594
R14783 gnd.n6555 gnd.n6554 99.6594
R14784 gnd.n5260 gnd.n5254 99.6594
R14785 gnd.n6562 gnd.n6561 99.6594
R14786 gnd.n5253 gnd.n5247 99.6594
R14787 gnd.n6569 gnd.n6568 99.6594
R14788 gnd.n5246 gnd.n5243 99.6594
R14789 gnd.n5225 gnd.n1171 99.6594
R14790 gnd.n5217 gnd.n1131 99.6594
R14791 gnd.n5213 gnd.n1132 99.6594
R14792 gnd.n5209 gnd.n1133 99.6594
R14793 gnd.n5205 gnd.n1134 99.6594
R14794 gnd.n5201 gnd.n1135 99.6594
R14795 gnd.n5197 gnd.n1136 99.6594
R14796 gnd.n5193 gnd.n1137 99.6594
R14797 gnd.n5188 gnd.n1138 99.6594
R14798 gnd.n5184 gnd.n1139 99.6594
R14799 gnd.n5180 gnd.n1140 99.6594
R14800 gnd.n5176 gnd.n1141 99.6594
R14801 gnd.n5172 gnd.n1142 99.6594
R14802 gnd.n5168 gnd.n1143 99.6594
R14803 gnd.n5164 gnd.n1144 99.6594
R14804 gnd.n5160 gnd.n1145 99.6594
R14805 gnd.n5156 gnd.n1146 99.6594
R14806 gnd.n5152 gnd.n1147 99.6594
R14807 gnd.n5148 gnd.n1148 99.6594
R14808 gnd.n5144 gnd.n1149 99.6594
R14809 gnd.n5140 gnd.n1150 99.6594
R14810 gnd.n5136 gnd.n1151 99.6594
R14811 gnd.n5132 gnd.n1152 99.6594
R14812 gnd.n5128 gnd.n1153 99.6594
R14813 gnd.n5124 gnd.n1154 99.6594
R14814 gnd.n5120 gnd.n1155 99.6594
R14815 gnd.n5116 gnd.n1156 99.6594
R14816 gnd.n5112 gnd.n1157 99.6594
R14817 gnd.n1241 gnd.n1158 99.6594
R14818 gnd.n2528 gnd.n2527 99.6594
R14819 gnd.n2519 gnd.n2424 99.6594
R14820 gnd.n2518 gnd.n2517 99.6594
R14821 gnd.n2509 gnd.n2428 99.6594
R14822 gnd.n2508 gnd.n2507 99.6594
R14823 gnd.n2499 gnd.n2432 99.6594
R14824 gnd.n2498 gnd.n2497 99.6594
R14825 gnd.n2489 gnd.n2436 99.6594
R14826 gnd.n2488 gnd.n2487 99.6594
R14827 gnd.n2479 gnd.n2440 99.6594
R14828 gnd.n2478 gnd.n2477 99.6594
R14829 gnd.n2469 gnd.n2446 99.6594
R14830 gnd.n2468 gnd.n2467 99.6594
R14831 gnd.n2459 gnd.n2450 99.6594
R14832 gnd.n2458 gnd.n2457 99.6594
R14833 gnd.n1532 gnd.n1527 99.6594
R14834 gnd.n4920 gnd.n4919 99.6594
R14835 gnd.n1526 gnd.n1520 99.6594
R14836 gnd.n4927 gnd.n4926 99.6594
R14837 gnd.n1519 gnd.n1511 99.6594
R14838 gnd.n4935 gnd.n4934 99.6594
R14839 gnd.n1510 gnd.n1504 99.6594
R14840 gnd.n4942 gnd.n4941 99.6594
R14841 gnd.n1503 gnd.n1497 99.6594
R14842 gnd.n4949 gnd.n4948 99.6594
R14843 gnd.n1496 gnd.n1489 99.6594
R14844 gnd.n4956 gnd.n4955 99.6594
R14845 gnd.n4959 gnd.n4958 99.6594
R14846 gnd.n4343 gnd.n4342 99.6594
R14847 gnd.n4345 gnd.n4334 99.6594
R14848 gnd.n4354 gnd.n4353 99.6594
R14849 gnd.n4355 gnd.n4330 99.6594
R14850 gnd.n4364 gnd.n4363 99.6594
R14851 gnd.n4365 gnd.n4326 99.6594
R14852 gnd.n4374 gnd.n4373 99.6594
R14853 gnd.n4375 gnd.n4322 99.6594
R14854 gnd.n4387 gnd.n4386 99.6594
R14855 gnd.n4388 gnd.n4318 99.6594
R14856 gnd.n4397 gnd.n4396 99.6594
R14857 gnd.n4398 gnd.n4314 99.6594
R14858 gnd.n4410 gnd.n4409 99.6594
R14859 gnd.n4411 gnd.n1963 99.6594
R14860 gnd.n4420 gnd.n4419 99.6594
R14861 gnd.n4421 gnd.n1959 99.6594
R14862 gnd.n4430 gnd.n4429 99.6594
R14863 gnd.n4431 gnd.n1955 99.6594
R14864 gnd.n4442 gnd.n4441 99.6594
R14865 gnd.n4443 gnd.n1951 99.6594
R14866 gnd.n4452 gnd.n4451 99.6594
R14867 gnd.n4453 gnd.n1947 99.6594
R14868 gnd.n4462 gnd.n4461 99.6594
R14869 gnd.n4463 gnd.n1943 99.6594
R14870 gnd.n4472 gnd.n4471 99.6594
R14871 gnd.n4473 gnd.n1939 99.6594
R14872 gnd.n4483 gnd.n4482 99.6594
R14873 gnd.n4486 gnd.n4485 99.6594
R14874 gnd.n7699 gnd.n7698 99.6594
R14875 gnd.n320 gnd.n312 99.6594
R14876 gnd.n7706 gnd.n7705 99.6594
R14877 gnd.n311 gnd.n305 99.6594
R14878 gnd.n7713 gnd.n7712 99.6594
R14879 gnd.n304 gnd.n298 99.6594
R14880 gnd.n7720 gnd.n7719 99.6594
R14881 gnd.n297 gnd.n291 99.6594
R14882 gnd.n7727 gnd.n7726 99.6594
R14883 gnd.n7730 gnd.n7729 99.6594
R14884 gnd.n288 gnd.n280 99.6594
R14885 gnd.n7739 gnd.n7738 99.6594
R14886 gnd.n279 gnd.n273 99.6594
R14887 gnd.n7746 gnd.n7745 99.6594
R14888 gnd.n272 gnd.n266 99.6594
R14889 gnd.n7753 gnd.n7752 99.6594
R14890 gnd.n265 gnd.n259 99.6594
R14891 gnd.n7760 gnd.n7759 99.6594
R14892 gnd.n258 gnd.n252 99.6594
R14893 gnd.n7767 gnd.n7766 99.6594
R14894 gnd.n251 gnd.n245 99.6594
R14895 gnd.n7777 gnd.n7776 99.6594
R14896 gnd.n244 gnd.n238 99.6594
R14897 gnd.n7784 gnd.n7783 99.6594
R14898 gnd.n237 gnd.n231 99.6594
R14899 gnd.n7791 gnd.n7790 99.6594
R14900 gnd.n230 gnd.n224 99.6594
R14901 gnd.n7798 gnd.n7797 99.6594
R14902 gnd.n222 gnd.n219 99.6594
R14903 gnd.n3221 gnd.n2387 99.6594
R14904 gnd.n2416 gnd.n2399 99.6594
R14905 gnd.n2418 gnd.n2400 99.6594
R14906 gnd.n2535 gnd.n2401 99.6594
R14907 gnd.n2537 gnd.n2402 99.6594
R14908 gnd.n2548 gnd.n2403 99.6594
R14909 gnd.n2550 gnd.n2404 99.6594
R14910 gnd.n2560 gnd.n2405 99.6594
R14911 gnd.n2571 gnd.n2406 99.6594
R14912 gnd.n2573 gnd.n2407 99.6594
R14913 gnd.n2583 gnd.n2408 99.6594
R14914 gnd.n2594 gnd.n2409 99.6594
R14915 gnd.n3146 gnd.n2410 99.6594
R14916 gnd.n3150 gnd.n2411 99.6594
R14917 gnd.n3221 gnd.n3220 99.6594
R14918 gnd.n2417 gnd.n2399 99.6594
R14919 gnd.n2534 gnd.n2400 99.6594
R14920 gnd.n2536 gnd.n2401 99.6594
R14921 gnd.n2547 gnd.n2402 99.6594
R14922 gnd.n2549 gnd.n2403 99.6594
R14923 gnd.n2559 gnd.n2404 99.6594
R14924 gnd.n2570 gnd.n2405 99.6594
R14925 gnd.n2572 gnd.n2406 99.6594
R14926 gnd.n2582 gnd.n2407 99.6594
R14927 gnd.n2593 gnd.n2408 99.6594
R14928 gnd.n2595 gnd.n2409 99.6594
R14929 gnd.n3149 gnd.n2410 99.6594
R14930 gnd.n3151 gnd.n2411 99.6594
R14931 gnd.n3991 gnd.n3986 99.6594
R14932 gnd.n3995 gnd.n3993 99.6594
R14933 gnd.n4002 gnd.n3982 99.6594
R14934 gnd.n4006 gnd.n4004 99.6594
R14935 gnd.n4017 gnd.n3979 99.6594
R14936 gnd.n4021 gnd.n4019 99.6594
R14937 gnd.n4036 gnd.n3970 99.6594
R14938 gnd.n4040 gnd.n4038 99.6594
R14939 gnd.n4055 gnd.n3961 99.6594
R14940 gnd.n4059 gnd.n4057 99.6594
R14941 gnd.n4074 gnd.n3952 99.6594
R14942 gnd.n4077 gnd.n4076 99.6594
R14943 gnd.n4095 gnd.n4094 99.6594
R14944 gnd.n4098 gnd.n4097 99.6594
R14945 gnd.n4076 gnd.n4075 99.6594
R14946 gnd.n4058 gnd.n3952 99.6594
R14947 gnd.n4057 gnd.n4056 99.6594
R14948 gnd.n4039 gnd.n3961 99.6594
R14949 gnd.n4038 gnd.n4037 99.6594
R14950 gnd.n4020 gnd.n3970 99.6594
R14951 gnd.n4019 gnd.n4018 99.6594
R14952 gnd.n4005 gnd.n3979 99.6594
R14953 gnd.n4004 gnd.n4003 99.6594
R14954 gnd.n3994 gnd.n3982 99.6594
R14955 gnd.n3993 gnd.n3992 99.6594
R14956 gnd.n3986 gnd.n1703 99.6594
R14957 gnd.n4099 gnd.n4098 99.6594
R14958 gnd.n4096 gnd.n4095 99.6594
R14959 gnd.n2596 gnd.t71 98.63
R14960 gnd.n3944 gnd.t90 98.63
R14961 gnd.n2603 gnd.t111 98.63
R14962 gnd.n4381 gnd.t87 98.63
R14963 gnd.n4433 gnd.t81 98.63
R14964 gnd.n1935 gnd.t22 98.63
R14965 gnd.n317 gnd.t108 98.63
R14966 gnd.n284 gnd.t29 98.63
R14967 gnd.n7770 gnd.t73 98.63
R14968 gnd.n354 gnd.t63 98.63
R14969 gnd.n1191 gnd.t40 98.63
R14970 gnd.n1213 gnd.t37 98.63
R14971 gnd.n1235 gnd.t26 98.63
R14972 gnd.n2720 gnd.t96 98.63
R14973 gnd.n1515 gnd.t101 98.63
R14974 gnd.n2421 gnd.t33 98.63
R14975 gnd.n2443 gnd.t66 98.63
R14976 gnd.n3934 gnd.t43 98.63
R14977 gnd.n3328 gnd.t123 88.9408
R14978 gnd.n2004 gnd.t119 88.9408
R14979 gnd.n4846 gnd.t55 88.933
R14980 gnd.n4175 gnd.t47 88.933
R14981 gnd.n1584 gnd.n1583 81.8399
R14982 gnd.n5662 gnd.t77 74.8376
R14983 gnd.n5267 gnd.t106 74.8376
R14984 gnd.n3329 gnd.t122 72.8438
R14985 gnd.n2005 gnd.t120 72.8438
R14986 gnd.n1585 gnd.n1578 72.8411
R14987 gnd.n1591 gnd.n1576 72.8411
R14988 gnd.n4171 gnd.n4170 72.8411
R14989 gnd.n2597 gnd.t70 72.836
R14990 gnd.n4847 gnd.t54 72.836
R14991 gnd.n4176 gnd.t48 72.836
R14992 gnd.n3945 gnd.t89 72.836
R14993 gnd.n2604 gnd.t112 72.836
R14994 gnd.n4382 gnd.t86 72.836
R14995 gnd.n4434 gnd.t80 72.836
R14996 gnd.n1936 gnd.t21 72.836
R14997 gnd.n318 gnd.t109 72.836
R14998 gnd.n285 gnd.t30 72.836
R14999 gnd.n7771 gnd.t74 72.836
R15000 gnd.n355 gnd.t64 72.836
R15001 gnd.n1192 gnd.t39 72.836
R15002 gnd.n1214 gnd.t36 72.836
R15003 gnd.n1236 gnd.t25 72.836
R15004 gnd.n2721 gnd.t95 72.836
R15005 gnd.n1516 gnd.t102 72.836
R15006 gnd.n2422 gnd.t34 72.836
R15007 gnd.n2444 gnd.t67 72.836
R15008 gnd.n3935 gnd.t44 72.836
R15009 gnd.n4236 gnd.n1972 71.676
R15010 gnd.n4232 gnd.n1973 71.676
R15011 gnd.n4228 gnd.n1974 71.676
R15012 gnd.n4224 gnd.n1975 71.676
R15013 gnd.n4220 gnd.n1976 71.676
R15014 gnd.n4216 gnd.n1977 71.676
R15015 gnd.n4212 gnd.n1978 71.676
R15016 gnd.n4208 gnd.n1979 71.676
R15017 gnd.n4204 gnd.n1980 71.676
R15018 gnd.n4200 gnd.n1981 71.676
R15019 gnd.n4196 gnd.n1982 71.676
R15020 gnd.n4192 gnd.n1983 71.676
R15021 gnd.n4188 gnd.n1984 71.676
R15022 gnd.n4184 gnd.n1985 71.676
R15023 gnd.n4179 gnd.n1986 71.676
R15024 gnd.n1987 gnd.n1970 71.676
R15025 gnd.n4308 gnd.n1969 71.676
R15026 gnd.n4306 gnd.n4305 71.676
R15027 gnd.n4300 gnd.n2002 71.676
R15028 gnd.n4296 gnd.n2001 71.676
R15029 gnd.n4292 gnd.n2000 71.676
R15030 gnd.n4288 gnd.n1999 71.676
R15031 gnd.n4284 gnd.n1998 71.676
R15032 gnd.n4280 gnd.n1997 71.676
R15033 gnd.n4276 gnd.n1996 71.676
R15034 gnd.n4272 gnd.n1995 71.676
R15035 gnd.n4268 gnd.n1994 71.676
R15036 gnd.n4264 gnd.n1993 71.676
R15037 gnd.n4260 gnd.n1992 71.676
R15038 gnd.n4256 gnd.n1991 71.676
R15039 gnd.n4252 gnd.n1990 71.676
R15040 gnd.n4248 gnd.n1989 71.676
R15041 gnd.n4244 gnd.n1988 71.676
R15042 gnd.n4910 gnd.n4909 71.676
R15043 gnd.n4904 gnd.n1540 71.676
R15044 gnd.n4901 gnd.n1541 71.676
R15045 gnd.n4897 gnd.n1542 71.676
R15046 gnd.n4893 gnd.n1543 71.676
R15047 gnd.n4889 gnd.n1544 71.676
R15048 gnd.n4885 gnd.n1545 71.676
R15049 gnd.n4881 gnd.n1546 71.676
R15050 gnd.n4877 gnd.n1547 71.676
R15051 gnd.n4873 gnd.n1548 71.676
R15052 gnd.n4869 gnd.n1549 71.676
R15053 gnd.n4865 gnd.n1550 71.676
R15054 gnd.n4861 gnd.n1551 71.676
R15055 gnd.n4857 gnd.n1552 71.676
R15056 gnd.n4853 gnd.n1553 71.676
R15057 gnd.n4849 gnd.n1554 71.676
R15058 gnd.n1555 gnd.n1538 71.676
R15059 gnd.n3332 gnd.n1556 71.676
R15060 gnd.n3337 gnd.n1557 71.676
R15061 gnd.n3341 gnd.n1558 71.676
R15062 gnd.n3345 gnd.n1559 71.676
R15063 gnd.n3349 gnd.n1560 71.676
R15064 gnd.n3353 gnd.n1561 71.676
R15065 gnd.n3357 gnd.n1562 71.676
R15066 gnd.n3361 gnd.n1563 71.676
R15067 gnd.n3365 gnd.n1564 71.676
R15068 gnd.n3369 gnd.n1565 71.676
R15069 gnd.n3373 gnd.n1566 71.676
R15070 gnd.n3377 gnd.n1567 71.676
R15071 gnd.n3381 gnd.n1568 71.676
R15072 gnd.n3385 gnd.n1569 71.676
R15073 gnd.n3389 gnd.n1570 71.676
R15074 gnd.n4910 gnd.n1573 71.676
R15075 gnd.n4902 gnd.n1540 71.676
R15076 gnd.n4898 gnd.n1541 71.676
R15077 gnd.n4894 gnd.n1542 71.676
R15078 gnd.n4890 gnd.n1543 71.676
R15079 gnd.n4886 gnd.n1544 71.676
R15080 gnd.n4882 gnd.n1545 71.676
R15081 gnd.n4878 gnd.n1546 71.676
R15082 gnd.n4874 gnd.n1547 71.676
R15083 gnd.n4870 gnd.n1548 71.676
R15084 gnd.n4866 gnd.n1549 71.676
R15085 gnd.n4862 gnd.n1550 71.676
R15086 gnd.n4858 gnd.n1551 71.676
R15087 gnd.n4854 gnd.n1552 71.676
R15088 gnd.n4850 gnd.n1553 71.676
R15089 gnd.n4913 gnd.n4912 71.676
R15090 gnd.n3331 gnd.n1555 71.676
R15091 gnd.n3336 gnd.n1556 71.676
R15092 gnd.n3340 gnd.n1557 71.676
R15093 gnd.n3344 gnd.n1558 71.676
R15094 gnd.n3348 gnd.n1559 71.676
R15095 gnd.n3352 gnd.n1560 71.676
R15096 gnd.n3356 gnd.n1561 71.676
R15097 gnd.n3360 gnd.n1562 71.676
R15098 gnd.n3364 gnd.n1563 71.676
R15099 gnd.n3368 gnd.n1564 71.676
R15100 gnd.n3372 gnd.n1565 71.676
R15101 gnd.n3376 gnd.n1566 71.676
R15102 gnd.n3380 gnd.n1567 71.676
R15103 gnd.n3384 gnd.n1568 71.676
R15104 gnd.n3388 gnd.n1569 71.676
R15105 gnd.n3392 gnd.n1570 71.676
R15106 gnd.n4247 gnd.n1988 71.676
R15107 gnd.n4251 gnd.n1989 71.676
R15108 gnd.n4255 gnd.n1990 71.676
R15109 gnd.n4259 gnd.n1991 71.676
R15110 gnd.n4263 gnd.n1992 71.676
R15111 gnd.n4267 gnd.n1993 71.676
R15112 gnd.n4271 gnd.n1994 71.676
R15113 gnd.n4275 gnd.n1995 71.676
R15114 gnd.n4279 gnd.n1996 71.676
R15115 gnd.n4283 gnd.n1997 71.676
R15116 gnd.n4287 gnd.n1998 71.676
R15117 gnd.n4291 gnd.n1999 71.676
R15118 gnd.n4295 gnd.n2000 71.676
R15119 gnd.n4299 gnd.n2001 71.676
R15120 gnd.n2003 gnd.n2002 71.676
R15121 gnd.n4307 gnd.n4306 71.676
R15122 gnd.n4311 gnd.n4310 71.676
R15123 gnd.n4178 gnd.n1987 71.676
R15124 gnd.n4183 gnd.n1986 71.676
R15125 gnd.n4187 gnd.n1985 71.676
R15126 gnd.n4191 gnd.n1984 71.676
R15127 gnd.n4195 gnd.n1983 71.676
R15128 gnd.n4199 gnd.n1982 71.676
R15129 gnd.n4203 gnd.n1981 71.676
R15130 gnd.n4207 gnd.n1980 71.676
R15131 gnd.n4211 gnd.n1979 71.676
R15132 gnd.n4215 gnd.n1978 71.676
R15133 gnd.n4219 gnd.n1977 71.676
R15134 gnd.n4223 gnd.n1976 71.676
R15135 gnd.n4227 gnd.n1975 71.676
R15136 gnd.n4231 gnd.n1974 71.676
R15137 gnd.n4235 gnd.n1973 71.676
R15138 gnd.n2011 gnd.n1972 71.676
R15139 gnd.n8 gnd.t358 69.1507
R15140 gnd.n14 gnd.t354 68.4792
R15141 gnd.n13 gnd.t334 68.4792
R15142 gnd.n12 gnd.t308 68.4792
R15143 gnd.n11 gnd.t362 68.4792
R15144 gnd.n10 gnd.t125 68.4792
R15145 gnd.n9 gnd.t366 68.4792
R15146 gnd.n8 gnd.t316 68.4792
R15147 gnd.n5789 gnd.n5693 64.369
R15148 gnd.n5235 gnd.n1125 59.5891
R15149 gnd.n7530 gnd.n7529 59.5891
R15150 gnd.n3334 gnd.n3329 59.5399
R15151 gnd.n4302 gnd.n2005 59.5399
R15152 gnd.n4848 gnd.n4847 59.5399
R15153 gnd.n4181 gnd.n4176 59.5399
R15154 gnd.n4845 gnd.n1594 59.1804
R15155 gnd.n6578 gnd.n5236 57.3586
R15156 gnd.n5444 gnd.t214 56.407
R15157 gnd.n5397 gnd.t277 56.407
R15158 gnd.n5412 gnd.t159 56.407
R15159 gnd.n5428 gnd.t266 56.407
R15160 gnd.n64 gnd.t180 56.407
R15161 gnd.n17 gnd.t168 56.407
R15162 gnd.n32 gnd.t289 56.407
R15163 gnd.n48 gnd.t230 56.407
R15164 gnd.n5457 gnd.t202 55.8337
R15165 gnd.n5410 gnd.t286 55.8337
R15166 gnd.n5425 gnd.t254 55.8337
R15167 gnd.n5441 gnd.t246 55.8337
R15168 gnd.n77 gnd.t140 55.8337
R15169 gnd.n30 gnd.t183 55.8337
R15170 gnd.n45 gnd.t241 55.8337
R15171 gnd.n61 gnd.t199 55.8337
R15172 gnd.n1582 gnd.n1581 54.358
R15173 gnd.n4168 gnd.n4167 54.358
R15174 gnd.n5444 gnd.n5443 53.0052
R15175 gnd.n5446 gnd.n5445 53.0052
R15176 gnd.n5448 gnd.n5447 53.0052
R15177 gnd.n5450 gnd.n5449 53.0052
R15178 gnd.n5452 gnd.n5451 53.0052
R15179 gnd.n5454 gnd.n5453 53.0052
R15180 gnd.n5456 gnd.n5455 53.0052
R15181 gnd.n5397 gnd.n5396 53.0052
R15182 gnd.n5399 gnd.n5398 53.0052
R15183 gnd.n5401 gnd.n5400 53.0052
R15184 gnd.n5403 gnd.n5402 53.0052
R15185 gnd.n5405 gnd.n5404 53.0052
R15186 gnd.n5407 gnd.n5406 53.0052
R15187 gnd.n5409 gnd.n5408 53.0052
R15188 gnd.n5412 gnd.n5411 53.0052
R15189 gnd.n5414 gnd.n5413 53.0052
R15190 gnd.n5416 gnd.n5415 53.0052
R15191 gnd.n5418 gnd.n5417 53.0052
R15192 gnd.n5420 gnd.n5419 53.0052
R15193 gnd.n5422 gnd.n5421 53.0052
R15194 gnd.n5424 gnd.n5423 53.0052
R15195 gnd.n5428 gnd.n5427 53.0052
R15196 gnd.n5430 gnd.n5429 53.0052
R15197 gnd.n5432 gnd.n5431 53.0052
R15198 gnd.n5434 gnd.n5433 53.0052
R15199 gnd.n5436 gnd.n5435 53.0052
R15200 gnd.n5438 gnd.n5437 53.0052
R15201 gnd.n5440 gnd.n5439 53.0052
R15202 gnd.n76 gnd.n75 53.0052
R15203 gnd.n74 gnd.n73 53.0052
R15204 gnd.n72 gnd.n71 53.0052
R15205 gnd.n70 gnd.n69 53.0052
R15206 gnd.n68 gnd.n67 53.0052
R15207 gnd.n66 gnd.n65 53.0052
R15208 gnd.n64 gnd.n63 53.0052
R15209 gnd.n29 gnd.n28 53.0052
R15210 gnd.n27 gnd.n26 53.0052
R15211 gnd.n25 gnd.n24 53.0052
R15212 gnd.n23 gnd.n22 53.0052
R15213 gnd.n21 gnd.n20 53.0052
R15214 gnd.n19 gnd.n18 53.0052
R15215 gnd.n17 gnd.n16 53.0052
R15216 gnd.n44 gnd.n43 53.0052
R15217 gnd.n42 gnd.n41 53.0052
R15218 gnd.n40 gnd.n39 53.0052
R15219 gnd.n38 gnd.n37 53.0052
R15220 gnd.n36 gnd.n35 53.0052
R15221 gnd.n34 gnd.n33 53.0052
R15222 gnd.n32 gnd.n31 53.0052
R15223 gnd.n60 gnd.n59 53.0052
R15224 gnd.n58 gnd.n57 53.0052
R15225 gnd.n56 gnd.n55 53.0052
R15226 gnd.n54 gnd.n53 53.0052
R15227 gnd.n52 gnd.n51 53.0052
R15228 gnd.n50 gnd.n49 53.0052
R15229 gnd.n48 gnd.n47 53.0052
R15230 gnd.n4159 gnd.n4158 52.4801
R15231 gnd.n6423 gnd.t364 52.3082
R15232 gnd.n6391 gnd.t360 52.3082
R15233 gnd.n6359 gnd.t318 52.3082
R15234 gnd.n6328 gnd.t338 52.3082
R15235 gnd.n6296 gnd.t342 52.3082
R15236 gnd.n6264 gnd.t349 52.3082
R15237 gnd.n6232 gnd.t340 52.3082
R15238 gnd.n6201 gnd.t347 52.3082
R15239 gnd.n6253 gnd.n6221 51.4173
R15240 gnd.n6317 gnd.n6316 50.455
R15241 gnd.n6285 gnd.n6284 50.455
R15242 gnd.n6253 gnd.n6252 50.455
R15243 gnd.n5736 gnd.n5735 45.1884
R15244 gnd.n5311 gnd.n5310 45.1884
R15245 gnd.n4239 gnd.n4174 44.3322
R15246 gnd.n1585 gnd.n1584 44.3189
R15247 gnd.n6796 gnd.n872 43.8952
R15248 gnd.n6790 gnd.n872 43.8952
R15249 gnd.n6790 gnd.n6789 43.8952
R15250 gnd.n6789 gnd.n6788 43.8952
R15251 gnd.n6788 gnd.n879 43.8952
R15252 gnd.n6782 gnd.n879 43.8952
R15253 gnd.n6782 gnd.n6781 43.8952
R15254 gnd.n6781 gnd.n6780 43.8952
R15255 gnd.n6780 gnd.n887 43.8952
R15256 gnd.n6774 gnd.n887 43.8952
R15257 gnd.n6774 gnd.n6773 43.8952
R15258 gnd.n6773 gnd.n6772 43.8952
R15259 gnd.n6772 gnd.n895 43.8952
R15260 gnd.n6766 gnd.n895 43.8952
R15261 gnd.n6766 gnd.n6765 43.8952
R15262 gnd.n6765 gnd.n6764 43.8952
R15263 gnd.n6764 gnd.n903 43.8952
R15264 gnd.n6758 gnd.n903 43.8952
R15265 gnd.n6758 gnd.n6757 43.8952
R15266 gnd.n6757 gnd.n6756 43.8952
R15267 gnd.n6756 gnd.n911 43.8952
R15268 gnd.n6750 gnd.n911 43.8952
R15269 gnd.n6750 gnd.n6749 43.8952
R15270 gnd.n6749 gnd.n6748 43.8952
R15271 gnd.n6748 gnd.n919 43.8952
R15272 gnd.n6742 gnd.n919 43.8952
R15273 gnd.n6742 gnd.n6741 43.8952
R15274 gnd.n6741 gnd.n6740 43.8952
R15275 gnd.n6740 gnd.n927 43.8952
R15276 gnd.n6734 gnd.n927 43.8952
R15277 gnd.n6734 gnd.n6733 43.8952
R15278 gnd.n6733 gnd.n6732 43.8952
R15279 gnd.n6732 gnd.n935 43.8952
R15280 gnd.n6726 gnd.n935 43.8952
R15281 gnd.n6726 gnd.n6725 43.8952
R15282 gnd.n6725 gnd.n6724 43.8952
R15283 gnd.n6724 gnd.n943 43.8952
R15284 gnd.n6718 gnd.n943 43.8952
R15285 gnd.n6718 gnd.n6717 43.8952
R15286 gnd.n6717 gnd.n6716 43.8952
R15287 gnd.n6716 gnd.n951 43.8952
R15288 gnd.n6710 gnd.n951 43.8952
R15289 gnd.n6710 gnd.n6709 43.8952
R15290 gnd.n6709 gnd.n6708 43.8952
R15291 gnd.n6708 gnd.n959 43.8952
R15292 gnd.n6702 gnd.n959 43.8952
R15293 gnd.n6702 gnd.n6701 43.8952
R15294 gnd.n6701 gnd.n6700 43.8952
R15295 gnd.n6700 gnd.n967 43.8952
R15296 gnd.n6694 gnd.n967 43.8952
R15297 gnd.n6694 gnd.n6693 43.8952
R15298 gnd.n6693 gnd.n6692 43.8952
R15299 gnd.n6692 gnd.n975 43.8952
R15300 gnd.n6686 gnd.n975 43.8952
R15301 gnd.n6686 gnd.n6685 43.8952
R15302 gnd.n6685 gnd.n6684 43.8952
R15303 gnd.n6684 gnd.n983 43.8952
R15304 gnd.n6678 gnd.n983 43.8952
R15305 gnd.n6678 gnd.n6677 43.8952
R15306 gnd.n6677 gnd.n6676 43.8952
R15307 gnd.n6676 gnd.n991 43.8952
R15308 gnd.n6670 gnd.n991 43.8952
R15309 gnd.n6670 gnd.n6669 43.8952
R15310 gnd.n6669 gnd.n6668 43.8952
R15311 gnd.n6668 gnd.n999 43.8952
R15312 gnd.n6662 gnd.n999 43.8952
R15313 gnd.n6662 gnd.n6661 43.8952
R15314 gnd.n6661 gnd.n6660 43.8952
R15315 gnd.n6660 gnd.n1007 43.8952
R15316 gnd.n6654 gnd.n1007 43.8952
R15317 gnd.n6654 gnd.n6653 43.8952
R15318 gnd.n6653 gnd.n6652 43.8952
R15319 gnd.n6652 gnd.n1015 43.8952
R15320 gnd.n6646 gnd.n1015 43.8952
R15321 gnd.n6646 gnd.n6645 43.8952
R15322 gnd.n6645 gnd.n6644 43.8952
R15323 gnd.n6644 gnd.n1023 43.8952
R15324 gnd.n6638 gnd.n1023 43.8952
R15325 gnd.n6638 gnd.n6637 43.8952
R15326 gnd.n6637 gnd.n6636 43.8952
R15327 gnd.n6636 gnd.n1031 43.8952
R15328 gnd.n6630 gnd.n1031 43.8952
R15329 gnd.n6630 gnd.n6629 43.8952
R15330 gnd.n2598 gnd.n2597 42.2793
R15331 gnd.n4090 gnd.n3945 42.2793
R15332 gnd.n5737 gnd.n5736 42.2793
R15333 gnd.n5312 gnd.n5311 42.2793
R15334 gnd.n5663 gnd.n5662 42.2793
R15335 gnd.n5268 gnd.n5267 42.2793
R15336 gnd.n3162 gnd.n2604 42.2793
R15337 gnd.n4383 gnd.n4382 42.2793
R15338 gnd.n4435 gnd.n4434 42.2793
R15339 gnd.n1937 gnd.n1936 42.2793
R15340 gnd.n319 gnd.n318 42.2793
R15341 gnd.n7735 gnd.n285 42.2793
R15342 gnd.n7772 gnd.n7771 42.2793
R15343 gnd.n7663 gnd.n355 42.2793
R15344 gnd.n5190 gnd.n1192 42.2793
R15345 gnd.n5150 gnd.n1214 42.2793
R15346 gnd.n5110 gnd.n1236 42.2793
R15347 gnd.n2771 gnd.n2721 42.2793
R15348 gnd.n4930 gnd.n1516 42.2793
R15349 gnd.n2423 gnd.n2422 42.2793
R15350 gnd.n2445 gnd.n2444 42.2793
R15351 gnd.n3936 gnd.n3935 42.2793
R15352 gnd.n1583 gnd.n1582 41.6274
R15353 gnd.n4169 gnd.n4168 41.6274
R15354 gnd.n1592 gnd.n1591 40.8975
R15355 gnd.n4172 gnd.n4171 40.8975
R15356 gnd.n1591 gnd.n1590 35.055
R15357 gnd.n1586 gnd.n1585 35.055
R15358 gnd.n4161 gnd.n4160 35.055
R15359 gnd.n4171 gnd.n4157 35.055
R15360 gnd.n5799 gnd.n5693 31.8661
R15361 gnd.n5799 gnd.n5798 31.8661
R15362 gnd.n5807 gnd.n5682 31.8661
R15363 gnd.n5815 gnd.n5682 31.8661
R15364 gnd.n5815 gnd.n5676 31.8661
R15365 gnd.n5823 gnd.n5676 31.8661
R15366 gnd.n5823 gnd.n5669 31.8661
R15367 gnd.n5861 gnd.n5669 31.8661
R15368 gnd.n5871 gnd.n5602 31.8661
R15369 gnd.n5227 gnd.n1125 31.8661
R15370 gnd.n3103 gnd.n1482 31.8661
R15371 gnd.n3098 gnd.n3097 31.8661
R15372 gnd.n3098 gnd.n2398 31.8661
R15373 gnd.n3223 gnd.n2388 31.8661
R15374 gnd.n4725 gnd.n1706 31.8661
R15375 gnd.n4719 gnd.n4718 31.8661
R15376 gnd.n4718 gnd.n4717 31.8661
R15377 gnd.n4711 gnd.n1724 31.8661
R15378 gnd.n7530 gnd.n433 31.8661
R15379 gnd.n5226 gnd.n1169 30.5915
R15380 gnd.n223 gnd.n215 30.5915
R15381 gnd.n4245 gnd.n2006 29.8151
R15382 gnd.n3396 gnd.n3391 29.8151
R15383 gnd.n5103 gnd.n1169 26.7676
R15384 gnd.n5100 gnd.n1244 26.7676
R15385 gnd.n5094 gnd.n1258 26.7676
R15386 gnd.n2788 gnd.n1261 26.7676
R15387 gnd.n5088 gnd.n1269 26.7676
R15388 gnd.n2838 gnd.n1272 26.7676
R15389 gnd.n2846 gnd.n1282 26.7676
R15390 gnd.n5076 gnd.n1289 26.7676
R15391 gnd.n5070 gnd.n1300 26.7676
R15392 gnd.n5064 gnd.n1310 26.7676
R15393 gnd.n2901 gnd.n1313 26.7676
R15394 gnd.n2895 gnd.n1323 26.7676
R15395 gnd.n5052 gnd.n1330 26.7676
R15396 gnd.n5046 gnd.n1341 26.7676
R15397 gnd.n5040 gnd.n1351 26.7676
R15398 gnd.n2690 gnd.n1354 26.7676
R15399 gnd.n2945 gnd.n2678 26.7676
R15400 gnd.n2942 gnd.n2680 26.7676
R15401 gnd.n2972 gnd.n2660 26.7676
R15402 gnd.n2979 gnd.n2978 26.7676
R15403 gnd.n3007 gnd.n2648 26.7676
R15404 gnd.n3015 gnd.n1371 26.7676
R15405 gnd.n5026 gnd.n1380 26.7676
R15406 gnd.n3022 gnd.n2642 26.7676
R15407 gnd.n5020 gnd.n1389 26.7676
R15408 gnd.n5014 gnd.n1399 26.7676
R15409 gnd.n3066 gnd.n1402 26.7676
R15410 gnd.n3037 gnd.n1412 26.7676
R15411 gnd.n5002 gnd.n1419 26.7676
R15412 gnd.n3043 gnd.n3042 26.7676
R15413 gnd.n4996 gnd.n1429 26.7676
R15414 gnd.n4990 gnd.n1439 26.7676
R15415 gnd.n3118 gnd.n1442 26.7676
R15416 gnd.n3124 gnd.n1452 26.7676
R15417 gnd.n4978 gnd.n1459 26.7676
R15418 gnd.n3133 gnd.n1462 26.7676
R15419 gnd.n4972 gnd.n1470 26.7676
R15420 gnd.n4966 gnd.n1479 26.7676
R15421 gnd.n4710 gnd.n1727 26.7676
R15422 gnd.n4704 gnd.n1739 26.7676
R15423 gnd.n4497 gnd.n1748 26.7676
R15424 gnd.n4698 gnd.n1751 26.7676
R15425 gnd.n4505 gnd.n1759 26.7676
R15426 gnd.n4511 gnd.n1768 26.7676
R15427 gnd.n4686 gnd.n1771 26.7676
R15428 gnd.n4680 gnd.n1782 26.7676
R15429 gnd.n4556 gnd.n4555 26.7676
R15430 gnd.n4674 gnd.n1791 26.7676
R15431 gnd.n4526 gnd.n1799 26.7676
R15432 gnd.n4531 gnd.n1808 26.7676
R15433 gnd.n4662 gnd.n1811 26.7676
R15434 gnd.n4656 gnd.n1822 26.7676
R15435 gnd.n4579 gnd.n4578 26.7676
R15436 gnd.n4650 gnd.n1831 26.7676
R15437 gnd.n4609 gnd.n1837 26.7676
R15438 gnd.n4620 gnd.n1846 26.7676
R15439 gnd.n4638 gnd.n1849 26.7676
R15440 gnd.n4587 gnd.n1857 26.7676
R15441 gnd.n7881 gnd.n87 26.7676
R15442 gnd.n7573 gnd.n391 26.7676
R15443 gnd.n7873 gnd.n105 26.7676
R15444 gnd.n7584 gnd.n114 26.7676
R15445 gnd.n7592 gnd.n123 26.7676
R15446 gnd.n7598 gnd.n132 26.7676
R15447 gnd.n7855 gnd.n135 26.7676
R15448 gnd.n7849 gnd.n146 26.7676
R15449 gnd.n7612 gnd.n153 26.7676
R15450 gnd.n7620 gnd.n163 26.7676
R15451 gnd.n7626 gnd.n172 26.7676
R15452 gnd.n7831 gnd.n175 26.7676
R15453 gnd.n7825 gnd.n186 26.7676
R15454 gnd.n7640 gnd.n193 26.7676
R15455 gnd.n7819 gnd.n196 26.7676
R15456 gnd.n7649 gnd.n204 26.7676
R15457 gnd.n7656 gnd.n212 26.7676
R15458 gnd.n7807 gnd.n215 26.7676
R15459 gnd.n2959 gnd.t216 26.4489
R15460 gnd.n4599 gnd.t181 26.4489
R15461 gnd.n6629 gnd.n6628 26.3373
R15462 gnd.n2889 gnd.t154 25.8116
R15463 gnd.n7861 gnd.t197 25.8116
R15464 gnd.n2597 gnd.n2596 25.7944
R15465 gnd.n3945 gnd.n3944 25.7944
R15466 gnd.n5662 gnd.n5661 25.7944
R15467 gnd.n5267 gnd.n5266 25.7944
R15468 gnd.n2604 gnd.n2603 25.7944
R15469 gnd.n4382 gnd.n4381 25.7944
R15470 gnd.n4434 gnd.n4433 25.7944
R15471 gnd.n1936 gnd.n1935 25.7944
R15472 gnd.n318 gnd.n317 25.7944
R15473 gnd.n285 gnd.n284 25.7944
R15474 gnd.n7771 gnd.n7770 25.7944
R15475 gnd.n355 gnd.n354 25.7944
R15476 gnd.n1192 gnd.n1191 25.7944
R15477 gnd.n1214 gnd.n1213 25.7944
R15478 gnd.n1236 gnd.n1235 25.7944
R15479 gnd.n2721 gnd.n2720 25.7944
R15480 gnd.n1516 gnd.n1515 25.7944
R15481 gnd.n2422 gnd.n2421 25.7944
R15482 gnd.n2444 gnd.n2443 25.7944
R15483 gnd.n3935 gnd.n3934 25.7944
R15484 gnd.n2853 gnd.t170 25.1743
R15485 gnd.n7837 gnd.t143 25.1743
R15486 gnd.n5883 gnd.n5603 24.8557
R15487 gnd.n5893 gnd.n5586 24.8557
R15488 gnd.n5589 gnd.n5577 24.8557
R15489 gnd.n5914 gnd.n5578 24.8557
R15490 gnd.n5924 gnd.n5558 24.8557
R15491 gnd.n5934 gnd.n5933 24.8557
R15492 gnd.n5544 gnd.n5542 24.8557
R15493 gnd.n5965 gnd.n5964 24.8557
R15494 gnd.n5980 gnd.n5527 24.8557
R15495 gnd.n6034 gnd.n5466 24.8557
R15496 gnd.n5990 gnd.n5467 24.8557
R15497 gnd.n6027 gnd.n5478 24.8557
R15498 gnd.n5516 gnd.n5515 24.8557
R15499 gnd.n6021 gnd.n6020 24.8557
R15500 gnd.n5502 gnd.n5489 24.8557
R15501 gnd.n6060 gnd.n6059 24.8557
R15502 gnd.n6070 gnd.n5382 24.8557
R15503 gnd.n6082 gnd.n5374 24.8557
R15504 gnd.n6081 gnd.n5362 24.8557
R15505 gnd.n6100 gnd.n6099 24.8557
R15506 gnd.n6110 gnd.n5355 24.8557
R15507 gnd.n6123 gnd.n5343 24.8557
R15508 gnd.n6156 gnd.n6155 24.8557
R15509 gnd.n6165 gnd.n5330 24.8557
R15510 gnd.n6621 gnd.n1049 24.8557
R15511 gnd.n6145 gnd.n1060 24.8557
R15512 gnd.n6614 gnd.n6613 24.8557
R15513 gnd.n6607 gnd.n1072 24.8557
R15514 gnd.n6470 gnd.n1085 24.8557
R15515 gnd.n6600 gnd.n6599 24.8557
R15516 gnd.n6593 gnd.n1097 24.8557
R15517 gnd.n6592 gnd.n1100 24.8557
R15518 gnd.n6459 gnd.n1111 24.8557
R15519 gnd.n6579 gnd.n1122 24.8557
R15520 gnd.n5904 gnd.t346 23.2624
R15521 gnd.n5605 gnd.t76 22.6251
R15522 gnd.t223 gnd.n1303 22.6251
R15523 gnd.n3140 gnd.t32 22.6251
R15524 gnd.n3925 gnd.t20 22.6251
R15525 gnd.n372 gnd.t189 22.6251
R15526 gnd.t203 gnd.n1344 21.9878
R15527 gnd.n384 gnd.t149 21.9878
R15528 gnd.t337 gnd.n5610 21.3504
R15529 gnd.n2663 gnd.t175 21.3504
R15530 gnd.t145 gnd.n4634 21.3504
R15531 gnd.n6138 gnd.t301 20.7131
R15532 gnd.t165 gnd.n1392 20.7131
R15533 gnd.t147 gnd.n1819 20.7131
R15534 gnd.n3103 gnd.n1487 20.3945
R15535 gnd.n1724 gnd.n1716 20.3945
R15536 gnd.t131 gnd.n5336 20.0758
R15537 gnd.t172 gnd.n1432 20.0758
R15538 gnd.t137 gnd.n1779 20.0758
R15539 gnd.n1580 gnd.t93 19.8005
R15540 gnd.n1580 gnd.t117 19.8005
R15541 gnd.n1579 gnd.t58 19.8005
R15542 gnd.n1579 gnd.t99 19.8005
R15543 gnd.n4166 gnd.t115 19.8005
R15544 gnd.n4166 gnd.t61 19.8005
R15545 gnd.n4165 gnd.t11 19.8005
R15546 gnd.n4165 gnd.t84 19.8005
R15547 gnd.n1576 gnd.n1575 19.5087
R15548 gnd.n1589 gnd.n1576 19.5087
R15549 gnd.n1587 gnd.n1578 19.5087
R15550 gnd.n4170 gnd.n4164 19.5087
R15551 gnd.n6071 gnd.t3 19.4385
R15552 gnd.n3152 gnd.n2379 19.3944
R15553 gnd.n3245 gnd.n2379 19.3944
R15554 gnd.n3245 gnd.n2376 19.3944
R15555 gnd.n3250 gnd.n2376 19.3944
R15556 gnd.n3250 gnd.n2377 19.3944
R15557 gnd.n2377 gnd.n2354 19.3944
R15558 gnd.n3275 gnd.n2354 19.3944
R15559 gnd.n3275 gnd.n2351 19.3944
R15560 gnd.n3282 gnd.n2351 19.3944
R15561 gnd.n3282 gnd.n2352 19.3944
R15562 gnd.n3278 gnd.n2352 19.3944
R15563 gnd.n3278 gnd.n2330 19.3944
R15564 gnd.n3321 gnd.n2330 19.3944
R15565 gnd.n3321 gnd.n2328 19.3944
R15566 gnd.n3325 gnd.n2328 19.3944
R15567 gnd.n3325 gnd.n2326 19.3944
R15568 gnd.n3412 gnd.n2326 19.3944
R15569 gnd.n3412 gnd.n2323 19.3944
R15570 gnd.n3417 gnd.n2323 19.3944
R15571 gnd.n3417 gnd.n2324 19.3944
R15572 gnd.n2324 gnd.n2301 19.3944
R15573 gnd.n3472 gnd.n2301 19.3944
R15574 gnd.n3472 gnd.n2299 19.3944
R15575 gnd.n3476 gnd.n2299 19.3944
R15576 gnd.n3476 gnd.n2280 19.3944
R15577 gnd.n3501 gnd.n2280 19.3944
R15578 gnd.n3501 gnd.n2277 19.3944
R15579 gnd.n3509 gnd.n2277 19.3944
R15580 gnd.n3509 gnd.n2278 19.3944
R15581 gnd.n3505 gnd.n2278 19.3944
R15582 gnd.n3505 gnd.n2245 19.3944
R15583 gnd.n3561 gnd.n2245 19.3944
R15584 gnd.n3561 gnd.n2242 19.3944
R15585 gnd.n3566 gnd.n2242 19.3944
R15586 gnd.n3566 gnd.n2243 19.3944
R15587 gnd.n2243 gnd.n2220 19.3944
R15588 gnd.n3615 gnd.n2220 19.3944
R15589 gnd.n3615 gnd.n2217 19.3944
R15590 gnd.n3631 gnd.n2217 19.3944
R15591 gnd.n3631 gnd.n2218 19.3944
R15592 gnd.n3627 gnd.n2218 19.3944
R15593 gnd.n3627 gnd.n3626 19.3944
R15594 gnd.n3626 gnd.n3625 19.3944
R15595 gnd.n3625 gnd.n3622 19.3944
R15596 gnd.n3622 gnd.n2174 19.3944
R15597 gnd.n3711 gnd.n2174 19.3944
R15598 gnd.n3711 gnd.n2171 19.3944
R15599 gnd.n3725 gnd.n2171 19.3944
R15600 gnd.n3725 gnd.n2172 19.3944
R15601 gnd.n3721 gnd.n2172 19.3944
R15602 gnd.n3721 gnd.n3720 19.3944
R15603 gnd.n3720 gnd.n3719 19.3944
R15604 gnd.n3719 gnd.n2134 19.3944
R15605 gnd.n3809 gnd.n2134 19.3944
R15606 gnd.n3809 gnd.n2131 19.3944
R15607 gnd.n3814 gnd.n2131 19.3944
R15608 gnd.n3814 gnd.n2132 19.3944
R15609 gnd.n2132 gnd.n2105 19.3944
R15610 gnd.n3847 gnd.n2105 19.3944
R15611 gnd.n3847 gnd.n2102 19.3944
R15612 gnd.n3859 gnd.n2102 19.3944
R15613 gnd.n3859 gnd.n2103 19.3944
R15614 gnd.n3855 gnd.n2103 19.3944
R15615 gnd.n3855 gnd.n3854 19.3944
R15616 gnd.n3854 gnd.n2069 19.3944
R15617 gnd.n3902 gnd.n2069 19.3944
R15618 gnd.n3903 gnd.n3902 19.3944
R15619 gnd.n3903 gnd.n2065 19.3944
R15620 gnd.n3907 gnd.n2065 19.3944
R15621 gnd.n3908 gnd.n3907 19.3944
R15622 gnd.n3909 gnd.n3908 19.3944
R15623 gnd.n3909 gnd.n2061 19.3944
R15624 gnd.n3913 gnd.n2061 19.3944
R15625 gnd.n3914 gnd.n3913 19.3944
R15626 gnd.n3915 gnd.n3914 19.3944
R15627 gnd.n3915 gnd.n2055 19.3944
R15628 gnd.n3919 gnd.n2055 19.3944
R15629 gnd.n3920 gnd.n3919 19.3944
R15630 gnd.n3921 gnd.n3920 19.3944
R15631 gnd.n3921 gnd.n2052 19.3944
R15632 gnd.n4104 gnd.n2052 19.3944
R15633 gnd.n4104 gnd.n2053 19.3944
R15634 gnd.n3148 gnd.n3147 19.3944
R15635 gnd.n3156 gnd.n3148 19.3944
R15636 gnd.n3156 gnd.n3155 19.3944
R15637 gnd.n3219 gnd.n2413 19.3944
R15638 gnd.n3219 gnd.n2414 19.3944
R15639 gnd.n3215 gnd.n2414 19.3944
R15640 gnd.n3215 gnd.n3214 19.3944
R15641 gnd.n3214 gnd.n3213 19.3944
R15642 gnd.n3213 gnd.n2419 19.3944
R15643 gnd.n3208 gnd.n2419 19.3944
R15644 gnd.n3208 gnd.n3207 19.3944
R15645 gnd.n3207 gnd.n3206 19.3944
R15646 gnd.n3206 gnd.n2538 19.3944
R15647 gnd.n3199 gnd.n2538 19.3944
R15648 gnd.n3199 gnd.n3198 19.3944
R15649 gnd.n3198 gnd.n2551 19.3944
R15650 gnd.n3191 gnd.n2551 19.3944
R15651 gnd.n3191 gnd.n3190 19.3944
R15652 gnd.n3190 gnd.n2561 19.3944
R15653 gnd.n3183 gnd.n2561 19.3944
R15654 gnd.n3183 gnd.n3182 19.3944
R15655 gnd.n3182 gnd.n2574 19.3944
R15656 gnd.n3175 gnd.n2574 19.3944
R15657 gnd.n3175 gnd.n3174 19.3944
R15658 gnd.n3174 gnd.n2584 19.3944
R15659 gnd.n3167 gnd.n2584 19.3944
R15660 gnd.n3167 gnd.n3166 19.3944
R15661 gnd.n4012 gnd.n3975 19.3944
R15662 gnd.n4025 gnd.n3975 19.3944
R15663 gnd.n4025 gnd.n3973 19.3944
R15664 gnd.n4031 gnd.n3973 19.3944
R15665 gnd.n4031 gnd.n3966 19.3944
R15666 gnd.n4044 gnd.n3966 19.3944
R15667 gnd.n4044 gnd.n3964 19.3944
R15668 gnd.n4050 gnd.n3964 19.3944
R15669 gnd.n4050 gnd.n3957 19.3944
R15670 gnd.n4063 gnd.n3957 19.3944
R15671 gnd.n4063 gnd.n3955 19.3944
R15672 gnd.n4069 gnd.n3955 19.3944
R15673 gnd.n4069 gnd.n3948 19.3944
R15674 gnd.n4083 gnd.n3948 19.3944
R15675 gnd.n4083 gnd.n3946 19.3944
R15676 gnd.n4089 gnd.n3946 19.3944
R15677 gnd.n5786 gnd.n5785 19.3944
R15678 gnd.n5785 gnd.n5784 19.3944
R15679 gnd.n5784 gnd.n5783 19.3944
R15680 gnd.n5783 gnd.n5781 19.3944
R15681 gnd.n5781 gnd.n5778 19.3944
R15682 gnd.n5778 gnd.n5777 19.3944
R15683 gnd.n5777 gnd.n5774 19.3944
R15684 gnd.n5774 gnd.n5773 19.3944
R15685 gnd.n5773 gnd.n5770 19.3944
R15686 gnd.n5770 gnd.n5769 19.3944
R15687 gnd.n5769 gnd.n5766 19.3944
R15688 gnd.n5766 gnd.n5765 19.3944
R15689 gnd.n5765 gnd.n5762 19.3944
R15690 gnd.n5762 gnd.n5761 19.3944
R15691 gnd.n5761 gnd.n5758 19.3944
R15692 gnd.n5758 gnd.n5757 19.3944
R15693 gnd.n5757 gnd.n5754 19.3944
R15694 gnd.n5754 gnd.n5753 19.3944
R15695 gnd.n5753 gnd.n5750 19.3944
R15696 gnd.n5750 gnd.n5749 19.3944
R15697 gnd.n5749 gnd.n5746 19.3944
R15698 gnd.n5746 gnd.n5745 19.3944
R15699 gnd.n5742 gnd.n5741 19.3944
R15700 gnd.n5741 gnd.n5697 19.3944
R15701 gnd.n5792 gnd.n5697 19.3944
R15702 gnd.n6499 gnd.n5314 19.3944
R15703 gnd.n6499 gnd.n6498 19.3944
R15704 gnd.n6498 gnd.n6497 19.3944
R15705 gnd.n6541 gnd.n6540 19.3944
R15706 gnd.n6540 gnd.n6539 19.3944
R15707 gnd.n6539 gnd.n5275 19.3944
R15708 gnd.n6534 gnd.n5275 19.3944
R15709 gnd.n6534 gnd.n6533 19.3944
R15710 gnd.n6533 gnd.n6532 19.3944
R15711 gnd.n6532 gnd.n5282 19.3944
R15712 gnd.n6527 gnd.n5282 19.3944
R15713 gnd.n6527 gnd.n6526 19.3944
R15714 gnd.n6526 gnd.n6525 19.3944
R15715 gnd.n6525 gnd.n5289 19.3944
R15716 gnd.n6520 gnd.n5289 19.3944
R15717 gnd.n6520 gnd.n6519 19.3944
R15718 gnd.n6519 gnd.n6518 19.3944
R15719 gnd.n6518 gnd.n5296 19.3944
R15720 gnd.n6513 gnd.n5296 19.3944
R15721 gnd.n6513 gnd.n6512 19.3944
R15722 gnd.n6512 gnd.n6511 19.3944
R15723 gnd.n6511 gnd.n5303 19.3944
R15724 gnd.n6506 gnd.n5303 19.3944
R15725 gnd.n6506 gnd.n6505 19.3944
R15726 gnd.n6505 gnd.n6504 19.3944
R15727 gnd.n5885 gnd.n5594 19.3944
R15728 gnd.n5895 gnd.n5594 19.3944
R15729 gnd.n5896 gnd.n5895 19.3944
R15730 gnd.n5896 gnd.n5575 19.3944
R15731 gnd.n5916 gnd.n5575 19.3944
R15732 gnd.n5916 gnd.n5567 19.3944
R15733 gnd.n5926 gnd.n5567 19.3944
R15734 gnd.n5927 gnd.n5926 19.3944
R15735 gnd.n5928 gnd.n5927 19.3944
R15736 gnd.n5928 gnd.n5550 19.3944
R15737 gnd.n5945 gnd.n5550 19.3944
R15738 gnd.n5948 gnd.n5945 19.3944
R15739 gnd.n5948 gnd.n5947 19.3944
R15740 gnd.n5947 gnd.n5523 19.3944
R15741 gnd.n5987 gnd.n5523 19.3944
R15742 gnd.n5987 gnd.n5520 19.3944
R15743 gnd.n5993 gnd.n5520 19.3944
R15744 gnd.n5994 gnd.n5993 19.3944
R15745 gnd.n5994 gnd.n5518 19.3944
R15746 gnd.n6000 gnd.n5518 19.3944
R15747 gnd.n6003 gnd.n6000 19.3944
R15748 gnd.n6005 gnd.n6003 19.3944
R15749 gnd.n6011 gnd.n6005 19.3944
R15750 gnd.n6011 gnd.n6010 19.3944
R15751 gnd.n6010 gnd.n5377 19.3944
R15752 gnd.n6077 gnd.n5377 19.3944
R15753 gnd.n6078 gnd.n6077 19.3944
R15754 gnd.n6078 gnd.n5370 19.3944
R15755 gnd.n6089 gnd.n5370 19.3944
R15756 gnd.n6090 gnd.n6089 19.3944
R15757 gnd.n6090 gnd.n5353 19.3944
R15758 gnd.n5353 gnd.n5351 19.3944
R15759 gnd.n6114 gnd.n5351 19.3944
R15760 gnd.n6117 gnd.n6114 19.3944
R15761 gnd.n6117 gnd.n6116 19.3944
R15762 gnd.n6116 gnd.n5327 19.3944
R15763 gnd.n6168 gnd.n5327 19.3944
R15764 gnd.n6169 gnd.n6168 19.3944
R15765 gnd.n6169 gnd.n5325 19.3944
R15766 gnd.n6175 gnd.n5325 19.3944
R15767 gnd.n6177 gnd.n6175 19.3944
R15768 gnd.n6181 gnd.n6177 19.3944
R15769 gnd.n6182 gnd.n6181 19.3944
R15770 gnd.n6468 gnd.n6182 19.3944
R15771 gnd.n6468 gnd.n6467 19.3944
R15772 gnd.n6467 gnd.n6466 19.3944
R15773 gnd.n6466 gnd.n6463 19.3944
R15774 gnd.n6463 gnd.n6462 19.3944
R15775 gnd.n6462 gnd.n6461 19.3944
R15776 gnd.n6461 gnd.n6458 19.3944
R15777 gnd.n6458 gnd.n6457 19.3944
R15778 gnd.n6457 gnd.n6454 19.3944
R15779 gnd.n6454 gnd.n6453 19.3944
R15780 gnd.n5876 gnd.n5875 19.3944
R15781 gnd.n5875 gnd.n5608 19.3944
R15782 gnd.n5631 gnd.n5608 19.3944
R15783 gnd.n5634 gnd.n5631 19.3944
R15784 gnd.n5634 gnd.n5627 19.3944
R15785 gnd.n5638 gnd.n5627 19.3944
R15786 gnd.n5641 gnd.n5638 19.3944
R15787 gnd.n5644 gnd.n5641 19.3944
R15788 gnd.n5644 gnd.n5625 19.3944
R15789 gnd.n5648 gnd.n5625 19.3944
R15790 gnd.n5651 gnd.n5648 19.3944
R15791 gnd.n5654 gnd.n5651 19.3944
R15792 gnd.n5654 gnd.n5623 19.3944
R15793 gnd.n5658 gnd.n5623 19.3944
R15794 gnd.n5881 gnd.n5880 19.3944
R15795 gnd.n5880 gnd.n5584 19.3944
R15796 gnd.n5906 gnd.n5584 19.3944
R15797 gnd.n5906 gnd.n5582 19.3944
R15798 gnd.n5912 gnd.n5582 19.3944
R15799 gnd.n5912 gnd.n5911 19.3944
R15800 gnd.n5911 gnd.n5556 19.3944
R15801 gnd.n5936 gnd.n5556 19.3944
R15802 gnd.n5936 gnd.n5554 19.3944
R15803 gnd.n5940 gnd.n5554 19.3944
R15804 gnd.n5940 gnd.n5534 19.3944
R15805 gnd.n5967 gnd.n5534 19.3944
R15806 gnd.n5967 gnd.n5532 19.3944
R15807 gnd.n5977 gnd.n5532 19.3944
R15808 gnd.n5977 gnd.n5976 19.3944
R15809 gnd.n5976 gnd.n5975 19.3944
R15810 gnd.n5975 gnd.n5481 19.3944
R15811 gnd.n6025 gnd.n5481 19.3944
R15812 gnd.n6025 gnd.n6024 19.3944
R15813 gnd.n6024 gnd.n6023 19.3944
R15814 gnd.n6023 gnd.n5485 19.3944
R15815 gnd.n5505 gnd.n5485 19.3944
R15816 gnd.n5505 gnd.n5387 19.3944
R15817 gnd.n6062 gnd.n5387 19.3944
R15818 gnd.n6062 gnd.n5385 19.3944
R15819 gnd.n6068 gnd.n5385 19.3944
R15820 gnd.n6068 gnd.n6067 19.3944
R15821 gnd.n6067 gnd.n5360 19.3944
R15822 gnd.n6102 gnd.n5360 19.3944
R15823 gnd.n6102 gnd.n5358 19.3944
R15824 gnd.n6108 gnd.n5358 19.3944
R15825 gnd.n6108 gnd.n6107 19.3944
R15826 gnd.n6107 gnd.n5334 19.3944
R15827 gnd.n6158 gnd.n5334 19.3944
R15828 gnd.n6158 gnd.n5332 19.3944
R15829 gnd.n6163 gnd.n5332 19.3944
R15830 gnd.n6163 gnd.n1054 19.3944
R15831 gnd.n6618 gnd.n1054 19.3944
R15832 gnd.n6618 gnd.n6617 19.3944
R15833 gnd.n6617 gnd.n6616 19.3944
R15834 gnd.n6616 gnd.n1058 19.3944
R15835 gnd.n1077 gnd.n1058 19.3944
R15836 gnd.n6604 gnd.n1077 19.3944
R15837 gnd.n6604 gnd.n6603 19.3944
R15838 gnd.n6603 gnd.n6602 19.3944
R15839 gnd.n6602 gnd.n1083 19.3944
R15840 gnd.n1103 gnd.n1083 19.3944
R15841 gnd.n6590 gnd.n1103 19.3944
R15842 gnd.n6590 gnd.n6589 19.3944
R15843 gnd.n6589 gnd.n6588 19.3944
R15844 gnd.n6588 gnd.n1109 19.3944
R15845 gnd.n5239 gnd.n1109 19.3944
R15846 gnd.n6576 gnd.n5239 19.3944
R15847 gnd.n6573 gnd.n6572 19.3944
R15848 gnd.n6572 gnd.n6571 19.3944
R15849 gnd.n6571 gnd.n5245 19.3944
R15850 gnd.n6566 gnd.n5245 19.3944
R15851 gnd.n6566 gnd.n6565 19.3944
R15852 gnd.n6565 gnd.n6564 19.3944
R15853 gnd.n6564 gnd.n5252 19.3944
R15854 gnd.n6559 gnd.n5252 19.3944
R15855 gnd.n6559 gnd.n6558 19.3944
R15856 gnd.n6558 gnd.n6557 19.3944
R15857 gnd.n6557 gnd.n5259 19.3944
R15858 gnd.n6552 gnd.n5259 19.3944
R15859 gnd.n6552 gnd.n6551 19.3944
R15860 gnd.n6551 gnd.n6550 19.3944
R15861 gnd.n5796 gnd.n5695 19.3944
R15862 gnd.n5796 gnd.n5686 19.3944
R15863 gnd.n5809 gnd.n5686 19.3944
R15864 gnd.n5809 gnd.n5684 19.3944
R15865 gnd.n5813 gnd.n5684 19.3944
R15866 gnd.n5813 gnd.n5674 19.3944
R15867 gnd.n5825 gnd.n5674 19.3944
R15868 gnd.n5825 gnd.n5672 19.3944
R15869 gnd.n5859 gnd.n5672 19.3944
R15870 gnd.n5859 gnd.n5858 19.3944
R15871 gnd.n5858 gnd.n5857 19.3944
R15872 gnd.n5857 gnd.n5856 19.3944
R15873 gnd.n5856 gnd.n5853 19.3944
R15874 gnd.n5853 gnd.n5852 19.3944
R15875 gnd.n5852 gnd.n5851 19.3944
R15876 gnd.n5851 gnd.n5849 19.3944
R15877 gnd.n5849 gnd.n5848 19.3944
R15878 gnd.n5848 gnd.n5845 19.3944
R15879 gnd.n5845 gnd.n5844 19.3944
R15880 gnd.n5844 gnd.n5843 19.3944
R15881 gnd.n5843 gnd.n5841 19.3944
R15882 gnd.n5841 gnd.n5540 19.3944
R15883 gnd.n5956 gnd.n5540 19.3944
R15884 gnd.n5956 gnd.n5538 19.3944
R15885 gnd.n5962 gnd.n5538 19.3944
R15886 gnd.n5962 gnd.n5961 19.3944
R15887 gnd.n5961 gnd.n5462 19.3944
R15888 gnd.n6036 gnd.n5462 19.3944
R15889 gnd.n6036 gnd.n5463 19.3944
R15890 gnd.n5510 gnd.n5509 19.3944
R15891 gnd.n5513 gnd.n5512 19.3944
R15892 gnd.n5500 gnd.n5499 19.3944
R15893 gnd.n6055 gnd.n5392 19.3944
R15894 gnd.n6055 gnd.n6054 19.3944
R15895 gnd.n6054 gnd.n6053 19.3944
R15896 gnd.n6053 gnd.n6051 19.3944
R15897 gnd.n6051 gnd.n6050 19.3944
R15898 gnd.n6050 gnd.n6048 19.3944
R15899 gnd.n6048 gnd.n6047 19.3944
R15900 gnd.n6047 gnd.n5341 19.3944
R15901 gnd.n6125 gnd.n5341 19.3944
R15902 gnd.n6125 gnd.n5339 19.3944
R15903 gnd.n6153 gnd.n5339 19.3944
R15904 gnd.n6153 gnd.n6152 19.3944
R15905 gnd.n6152 gnd.n6151 19.3944
R15906 gnd.n6151 gnd.n6149 19.3944
R15907 gnd.n6149 gnd.n6148 19.3944
R15908 gnd.n6148 gnd.n6142 19.3944
R15909 gnd.n6142 gnd.n6141 19.3944
R15910 gnd.n6141 gnd.n6140 19.3944
R15911 gnd.n6140 gnd.n6137 19.3944
R15912 gnd.n6137 gnd.n5324 19.3944
R15913 gnd.n6474 gnd.n5324 19.3944
R15914 gnd.n6474 gnd.n5322 19.3944
R15915 gnd.n6480 gnd.n5322 19.3944
R15916 gnd.n6481 gnd.n6480 19.3944
R15917 gnd.n6484 gnd.n6481 19.3944
R15918 gnd.n6484 gnd.n5320 19.3944
R15919 gnd.n6488 gnd.n5320 19.3944
R15920 gnd.n6491 gnd.n6488 19.3944
R15921 gnd.n6492 gnd.n6491 19.3944
R15922 gnd.n5801 gnd.n5691 19.3944
R15923 gnd.n5801 gnd.n5689 19.3944
R15924 gnd.n5805 gnd.n5689 19.3944
R15925 gnd.n5805 gnd.n5680 19.3944
R15926 gnd.n5817 gnd.n5680 19.3944
R15927 gnd.n5817 gnd.n5678 19.3944
R15928 gnd.n5821 gnd.n5678 19.3944
R15929 gnd.n5821 gnd.n5667 19.3944
R15930 gnd.n5863 gnd.n5667 19.3944
R15931 gnd.n5863 gnd.n5621 19.3944
R15932 gnd.n5869 gnd.n5621 19.3944
R15933 gnd.n5869 gnd.n5868 19.3944
R15934 gnd.n5868 gnd.n5599 19.3944
R15935 gnd.n5890 gnd.n5599 19.3944
R15936 gnd.n5890 gnd.n5592 19.3944
R15937 gnd.n5901 gnd.n5592 19.3944
R15938 gnd.n5901 gnd.n5900 19.3944
R15939 gnd.n5900 gnd.n5573 19.3944
R15940 gnd.n5921 gnd.n5573 19.3944
R15941 gnd.n5921 gnd.n5563 19.3944
R15942 gnd.n5931 gnd.n5563 19.3944
R15943 gnd.n5931 gnd.n5546 19.3944
R15944 gnd.n5952 gnd.n5546 19.3944
R15945 gnd.n5952 gnd.n5951 19.3944
R15946 gnd.n5951 gnd.n5525 19.3944
R15947 gnd.n5982 gnd.n5525 19.3944
R15948 gnd.n5982 gnd.n5470 19.3944
R15949 gnd.n6032 gnd.n5470 19.3944
R15950 gnd.n6032 gnd.n6031 19.3944
R15951 gnd.n6031 gnd.n6030 19.3944
R15952 gnd.n6030 gnd.n5474 19.3944
R15953 gnd.n5492 gnd.n5474 19.3944
R15954 gnd.n6018 gnd.n5492 19.3944
R15955 gnd.n6018 gnd.n6017 19.3944
R15956 gnd.n6017 gnd.n6016 19.3944
R15957 gnd.n6016 gnd.n5496 19.3944
R15958 gnd.n5496 gnd.n5379 19.3944
R15959 gnd.n6073 gnd.n5379 19.3944
R15960 gnd.n6073 gnd.n5372 19.3944
R15961 gnd.n6084 gnd.n5372 19.3944
R15962 gnd.n6084 gnd.n5368 19.3944
R15963 gnd.n6097 gnd.n5368 19.3944
R15964 gnd.n6097 gnd.n6096 19.3944
R15965 gnd.n6096 gnd.n5347 19.3944
R15966 gnd.n6121 gnd.n5347 19.3944
R15967 gnd.n6121 gnd.n6120 19.3944
R15968 gnd.n6120 gnd.n1043 19.3944
R15969 gnd.n6625 gnd.n1043 19.3944
R15970 gnd.n6625 gnd.n6624 19.3944
R15971 gnd.n6624 gnd.n6623 19.3944
R15972 gnd.n6623 gnd.n1047 19.3944
R15973 gnd.n1066 gnd.n1047 19.3944
R15974 gnd.n6611 gnd.n1066 19.3944
R15975 gnd.n6611 gnd.n6610 19.3944
R15976 gnd.n6610 gnd.n6609 19.3944
R15977 gnd.n6609 gnd.n1070 19.3944
R15978 gnd.n1091 gnd.n1070 19.3944
R15979 gnd.n6597 gnd.n1091 19.3944
R15980 gnd.n6597 gnd.n6596 19.3944
R15981 gnd.n6596 gnd.n6595 19.3944
R15982 gnd.n6595 gnd.n1095 19.3944
R15983 gnd.n1117 gnd.n1095 19.3944
R15984 gnd.n6583 gnd.n1117 19.3944
R15985 gnd.n6583 gnd.n6582 19.3944
R15986 gnd.n6582 gnd.n6581 19.3944
R15987 gnd.n3203 gnd.n2541 19.3944
R15988 gnd.n3203 gnd.n3202 19.3944
R15989 gnd.n3202 gnd.n2545 19.3944
R15990 gnd.n3195 gnd.n2545 19.3944
R15991 gnd.n3195 gnd.n3194 19.3944
R15992 gnd.n3194 gnd.n2557 19.3944
R15993 gnd.n3187 gnd.n2557 19.3944
R15994 gnd.n3187 gnd.n3186 19.3944
R15995 gnd.n3186 gnd.n2568 19.3944
R15996 gnd.n3179 gnd.n2568 19.3944
R15997 gnd.n3179 gnd.n3178 19.3944
R15998 gnd.n3178 gnd.n2580 19.3944
R15999 gnd.n3171 gnd.n2580 19.3944
R16000 gnd.n3171 gnd.n3170 19.3944
R16001 gnd.n3170 gnd.n2591 19.3944
R16002 gnd.n3163 gnd.n2591 19.3944
R16003 gnd.n7320 gnd.n558 19.3944
R16004 gnd.n7320 gnd.n556 19.3944
R16005 gnd.n7324 gnd.n556 19.3944
R16006 gnd.n7324 gnd.n552 19.3944
R16007 gnd.n7330 gnd.n552 19.3944
R16008 gnd.n7330 gnd.n550 19.3944
R16009 gnd.n7334 gnd.n550 19.3944
R16010 gnd.n7334 gnd.n546 19.3944
R16011 gnd.n7340 gnd.n546 19.3944
R16012 gnd.n7340 gnd.n544 19.3944
R16013 gnd.n7344 gnd.n544 19.3944
R16014 gnd.n7344 gnd.n540 19.3944
R16015 gnd.n7350 gnd.n540 19.3944
R16016 gnd.n7350 gnd.n538 19.3944
R16017 gnd.n7354 gnd.n538 19.3944
R16018 gnd.n7354 gnd.n534 19.3944
R16019 gnd.n7360 gnd.n534 19.3944
R16020 gnd.n7360 gnd.n532 19.3944
R16021 gnd.n7364 gnd.n532 19.3944
R16022 gnd.n7364 gnd.n528 19.3944
R16023 gnd.n7370 gnd.n528 19.3944
R16024 gnd.n7370 gnd.n526 19.3944
R16025 gnd.n7374 gnd.n526 19.3944
R16026 gnd.n7374 gnd.n522 19.3944
R16027 gnd.n7380 gnd.n522 19.3944
R16028 gnd.n7380 gnd.n520 19.3944
R16029 gnd.n7384 gnd.n520 19.3944
R16030 gnd.n7384 gnd.n516 19.3944
R16031 gnd.n7390 gnd.n516 19.3944
R16032 gnd.n7390 gnd.n514 19.3944
R16033 gnd.n7394 gnd.n514 19.3944
R16034 gnd.n7394 gnd.n510 19.3944
R16035 gnd.n7400 gnd.n510 19.3944
R16036 gnd.n7400 gnd.n508 19.3944
R16037 gnd.n7404 gnd.n508 19.3944
R16038 gnd.n7404 gnd.n504 19.3944
R16039 gnd.n7410 gnd.n504 19.3944
R16040 gnd.n7410 gnd.n502 19.3944
R16041 gnd.n7414 gnd.n502 19.3944
R16042 gnd.n7414 gnd.n498 19.3944
R16043 gnd.n7420 gnd.n498 19.3944
R16044 gnd.n7420 gnd.n496 19.3944
R16045 gnd.n7424 gnd.n496 19.3944
R16046 gnd.n7424 gnd.n492 19.3944
R16047 gnd.n7430 gnd.n492 19.3944
R16048 gnd.n7430 gnd.n490 19.3944
R16049 gnd.n7434 gnd.n490 19.3944
R16050 gnd.n7434 gnd.n486 19.3944
R16051 gnd.n7440 gnd.n486 19.3944
R16052 gnd.n7440 gnd.n484 19.3944
R16053 gnd.n7444 gnd.n484 19.3944
R16054 gnd.n7444 gnd.n480 19.3944
R16055 gnd.n7450 gnd.n480 19.3944
R16056 gnd.n7450 gnd.n478 19.3944
R16057 gnd.n7454 gnd.n478 19.3944
R16058 gnd.n7454 gnd.n474 19.3944
R16059 gnd.n7460 gnd.n474 19.3944
R16060 gnd.n7460 gnd.n472 19.3944
R16061 gnd.n7464 gnd.n472 19.3944
R16062 gnd.n7464 gnd.n468 19.3944
R16063 gnd.n7470 gnd.n468 19.3944
R16064 gnd.n7470 gnd.n466 19.3944
R16065 gnd.n7474 gnd.n466 19.3944
R16066 gnd.n7474 gnd.n462 19.3944
R16067 gnd.n7480 gnd.n462 19.3944
R16068 gnd.n7480 gnd.n460 19.3944
R16069 gnd.n7484 gnd.n460 19.3944
R16070 gnd.n7484 gnd.n456 19.3944
R16071 gnd.n7490 gnd.n456 19.3944
R16072 gnd.n7490 gnd.n454 19.3944
R16073 gnd.n7494 gnd.n454 19.3944
R16074 gnd.n7494 gnd.n450 19.3944
R16075 gnd.n7500 gnd.n450 19.3944
R16076 gnd.n7500 gnd.n448 19.3944
R16077 gnd.n7504 gnd.n448 19.3944
R16078 gnd.n7504 gnd.n444 19.3944
R16079 gnd.n7510 gnd.n444 19.3944
R16080 gnd.n7510 gnd.n442 19.3944
R16081 gnd.n7514 gnd.n442 19.3944
R16082 gnd.n7514 gnd.n438 19.3944
R16083 gnd.n7520 gnd.n438 19.3944
R16084 gnd.n7520 gnd.n436 19.3944
R16085 gnd.n7526 gnd.n436 19.3944
R16086 gnd.n7526 gnd.n7525 19.3944
R16087 gnd.n6800 gnd.n870 19.3944
R16088 gnd.n6800 gnd.n868 19.3944
R16089 gnd.n6804 gnd.n868 19.3944
R16090 gnd.n6804 gnd.n864 19.3944
R16091 gnd.n6810 gnd.n864 19.3944
R16092 gnd.n6810 gnd.n862 19.3944
R16093 gnd.n6814 gnd.n862 19.3944
R16094 gnd.n6814 gnd.n858 19.3944
R16095 gnd.n6820 gnd.n858 19.3944
R16096 gnd.n6820 gnd.n856 19.3944
R16097 gnd.n6824 gnd.n856 19.3944
R16098 gnd.n6824 gnd.n852 19.3944
R16099 gnd.n6830 gnd.n852 19.3944
R16100 gnd.n6830 gnd.n850 19.3944
R16101 gnd.n6834 gnd.n850 19.3944
R16102 gnd.n6834 gnd.n846 19.3944
R16103 gnd.n6840 gnd.n846 19.3944
R16104 gnd.n6840 gnd.n844 19.3944
R16105 gnd.n6844 gnd.n844 19.3944
R16106 gnd.n6844 gnd.n840 19.3944
R16107 gnd.n6850 gnd.n840 19.3944
R16108 gnd.n6850 gnd.n838 19.3944
R16109 gnd.n6854 gnd.n838 19.3944
R16110 gnd.n6854 gnd.n834 19.3944
R16111 gnd.n6860 gnd.n834 19.3944
R16112 gnd.n6860 gnd.n832 19.3944
R16113 gnd.n6864 gnd.n832 19.3944
R16114 gnd.n6864 gnd.n828 19.3944
R16115 gnd.n6870 gnd.n828 19.3944
R16116 gnd.n6870 gnd.n826 19.3944
R16117 gnd.n6874 gnd.n826 19.3944
R16118 gnd.n6874 gnd.n822 19.3944
R16119 gnd.n6880 gnd.n822 19.3944
R16120 gnd.n6880 gnd.n820 19.3944
R16121 gnd.n6884 gnd.n820 19.3944
R16122 gnd.n6884 gnd.n816 19.3944
R16123 gnd.n6890 gnd.n816 19.3944
R16124 gnd.n6890 gnd.n814 19.3944
R16125 gnd.n6894 gnd.n814 19.3944
R16126 gnd.n6894 gnd.n810 19.3944
R16127 gnd.n6900 gnd.n810 19.3944
R16128 gnd.n6900 gnd.n808 19.3944
R16129 gnd.n6904 gnd.n808 19.3944
R16130 gnd.n6904 gnd.n804 19.3944
R16131 gnd.n6910 gnd.n804 19.3944
R16132 gnd.n6910 gnd.n802 19.3944
R16133 gnd.n6914 gnd.n802 19.3944
R16134 gnd.n6914 gnd.n798 19.3944
R16135 gnd.n6920 gnd.n798 19.3944
R16136 gnd.n6920 gnd.n796 19.3944
R16137 gnd.n6924 gnd.n796 19.3944
R16138 gnd.n6924 gnd.n792 19.3944
R16139 gnd.n6930 gnd.n792 19.3944
R16140 gnd.n6930 gnd.n790 19.3944
R16141 gnd.n6934 gnd.n790 19.3944
R16142 gnd.n6934 gnd.n786 19.3944
R16143 gnd.n6940 gnd.n786 19.3944
R16144 gnd.n6940 gnd.n784 19.3944
R16145 gnd.n6944 gnd.n784 19.3944
R16146 gnd.n6944 gnd.n780 19.3944
R16147 gnd.n6950 gnd.n780 19.3944
R16148 gnd.n6950 gnd.n778 19.3944
R16149 gnd.n6954 gnd.n778 19.3944
R16150 gnd.n6954 gnd.n774 19.3944
R16151 gnd.n6960 gnd.n774 19.3944
R16152 gnd.n6960 gnd.n772 19.3944
R16153 gnd.n6964 gnd.n772 19.3944
R16154 gnd.n6964 gnd.n768 19.3944
R16155 gnd.n6970 gnd.n768 19.3944
R16156 gnd.n6970 gnd.n766 19.3944
R16157 gnd.n6974 gnd.n766 19.3944
R16158 gnd.n6974 gnd.n762 19.3944
R16159 gnd.n6980 gnd.n762 19.3944
R16160 gnd.n6980 gnd.n760 19.3944
R16161 gnd.n6984 gnd.n760 19.3944
R16162 gnd.n6984 gnd.n756 19.3944
R16163 gnd.n6990 gnd.n756 19.3944
R16164 gnd.n6990 gnd.n754 19.3944
R16165 gnd.n6994 gnd.n754 19.3944
R16166 gnd.n6994 gnd.n750 19.3944
R16167 gnd.n7000 gnd.n750 19.3944
R16168 gnd.n7000 gnd.n748 19.3944
R16169 gnd.n7004 gnd.n748 19.3944
R16170 gnd.n7004 gnd.n744 19.3944
R16171 gnd.n7010 gnd.n744 19.3944
R16172 gnd.n7010 gnd.n742 19.3944
R16173 gnd.n7014 gnd.n742 19.3944
R16174 gnd.n7014 gnd.n738 19.3944
R16175 gnd.n7020 gnd.n738 19.3944
R16176 gnd.n7020 gnd.n736 19.3944
R16177 gnd.n7024 gnd.n736 19.3944
R16178 gnd.n7024 gnd.n732 19.3944
R16179 gnd.n7030 gnd.n732 19.3944
R16180 gnd.n7030 gnd.n730 19.3944
R16181 gnd.n7034 gnd.n730 19.3944
R16182 gnd.n7034 gnd.n726 19.3944
R16183 gnd.n7040 gnd.n726 19.3944
R16184 gnd.n7040 gnd.n724 19.3944
R16185 gnd.n7044 gnd.n724 19.3944
R16186 gnd.n7044 gnd.n720 19.3944
R16187 gnd.n7050 gnd.n720 19.3944
R16188 gnd.n7050 gnd.n718 19.3944
R16189 gnd.n7054 gnd.n718 19.3944
R16190 gnd.n7054 gnd.n714 19.3944
R16191 gnd.n7060 gnd.n714 19.3944
R16192 gnd.n7060 gnd.n712 19.3944
R16193 gnd.n7064 gnd.n712 19.3944
R16194 gnd.n7064 gnd.n708 19.3944
R16195 gnd.n7070 gnd.n708 19.3944
R16196 gnd.n7070 gnd.n706 19.3944
R16197 gnd.n7074 gnd.n706 19.3944
R16198 gnd.n7074 gnd.n702 19.3944
R16199 gnd.n7080 gnd.n702 19.3944
R16200 gnd.n7080 gnd.n700 19.3944
R16201 gnd.n7084 gnd.n700 19.3944
R16202 gnd.n7084 gnd.n696 19.3944
R16203 gnd.n7090 gnd.n696 19.3944
R16204 gnd.n7090 gnd.n694 19.3944
R16205 gnd.n7094 gnd.n694 19.3944
R16206 gnd.n7094 gnd.n690 19.3944
R16207 gnd.n7100 gnd.n690 19.3944
R16208 gnd.n7100 gnd.n688 19.3944
R16209 gnd.n7104 gnd.n688 19.3944
R16210 gnd.n7104 gnd.n684 19.3944
R16211 gnd.n7110 gnd.n684 19.3944
R16212 gnd.n7110 gnd.n682 19.3944
R16213 gnd.n7114 gnd.n682 19.3944
R16214 gnd.n7114 gnd.n678 19.3944
R16215 gnd.n7120 gnd.n678 19.3944
R16216 gnd.n7120 gnd.n676 19.3944
R16217 gnd.n7124 gnd.n676 19.3944
R16218 gnd.n7124 gnd.n672 19.3944
R16219 gnd.n7130 gnd.n672 19.3944
R16220 gnd.n7130 gnd.n670 19.3944
R16221 gnd.n7134 gnd.n670 19.3944
R16222 gnd.n7134 gnd.n666 19.3944
R16223 gnd.n7140 gnd.n666 19.3944
R16224 gnd.n7140 gnd.n664 19.3944
R16225 gnd.n7144 gnd.n664 19.3944
R16226 gnd.n7144 gnd.n660 19.3944
R16227 gnd.n7150 gnd.n660 19.3944
R16228 gnd.n7150 gnd.n658 19.3944
R16229 gnd.n7154 gnd.n658 19.3944
R16230 gnd.n7154 gnd.n654 19.3944
R16231 gnd.n7160 gnd.n654 19.3944
R16232 gnd.n7160 gnd.n652 19.3944
R16233 gnd.n7164 gnd.n652 19.3944
R16234 gnd.n7164 gnd.n648 19.3944
R16235 gnd.n7170 gnd.n648 19.3944
R16236 gnd.n7170 gnd.n646 19.3944
R16237 gnd.n7174 gnd.n646 19.3944
R16238 gnd.n7174 gnd.n642 19.3944
R16239 gnd.n7180 gnd.n642 19.3944
R16240 gnd.n7180 gnd.n640 19.3944
R16241 gnd.n7184 gnd.n640 19.3944
R16242 gnd.n7184 gnd.n636 19.3944
R16243 gnd.n7190 gnd.n636 19.3944
R16244 gnd.n7190 gnd.n634 19.3944
R16245 gnd.n7194 gnd.n634 19.3944
R16246 gnd.n7194 gnd.n630 19.3944
R16247 gnd.n7200 gnd.n630 19.3944
R16248 gnd.n7200 gnd.n628 19.3944
R16249 gnd.n7204 gnd.n628 19.3944
R16250 gnd.n7204 gnd.n624 19.3944
R16251 gnd.n7210 gnd.n624 19.3944
R16252 gnd.n7210 gnd.n622 19.3944
R16253 gnd.n7214 gnd.n622 19.3944
R16254 gnd.n7214 gnd.n618 19.3944
R16255 gnd.n7220 gnd.n618 19.3944
R16256 gnd.n7220 gnd.n616 19.3944
R16257 gnd.n7224 gnd.n616 19.3944
R16258 gnd.n7224 gnd.n612 19.3944
R16259 gnd.n7230 gnd.n612 19.3944
R16260 gnd.n7230 gnd.n610 19.3944
R16261 gnd.n7234 gnd.n610 19.3944
R16262 gnd.n7234 gnd.n606 19.3944
R16263 gnd.n7240 gnd.n606 19.3944
R16264 gnd.n7240 gnd.n604 19.3944
R16265 gnd.n7244 gnd.n604 19.3944
R16266 gnd.n7244 gnd.n600 19.3944
R16267 gnd.n7250 gnd.n600 19.3944
R16268 gnd.n7250 gnd.n598 19.3944
R16269 gnd.n7254 gnd.n598 19.3944
R16270 gnd.n7254 gnd.n594 19.3944
R16271 gnd.n7260 gnd.n594 19.3944
R16272 gnd.n7260 gnd.n592 19.3944
R16273 gnd.n7264 gnd.n592 19.3944
R16274 gnd.n7264 gnd.n588 19.3944
R16275 gnd.n7270 gnd.n588 19.3944
R16276 gnd.n7270 gnd.n586 19.3944
R16277 gnd.n7274 gnd.n586 19.3944
R16278 gnd.n7274 gnd.n582 19.3944
R16279 gnd.n7280 gnd.n582 19.3944
R16280 gnd.n7280 gnd.n580 19.3944
R16281 gnd.n7284 gnd.n580 19.3944
R16282 gnd.n7284 gnd.n576 19.3944
R16283 gnd.n7290 gnd.n576 19.3944
R16284 gnd.n7290 gnd.n574 19.3944
R16285 gnd.n7294 gnd.n574 19.3944
R16286 gnd.n7294 gnd.n570 19.3944
R16287 gnd.n7300 gnd.n570 19.3944
R16288 gnd.n7300 gnd.n568 19.3944
R16289 gnd.n7304 gnd.n568 19.3944
R16290 gnd.n7304 gnd.n564 19.3944
R16291 gnd.n7310 gnd.n564 19.3944
R16292 gnd.n7310 gnd.n562 19.3944
R16293 gnd.n7314 gnd.n562 19.3944
R16294 gnd.n4341 gnd.n4338 19.3944
R16295 gnd.n4341 gnd.n4337 19.3944
R16296 gnd.n4347 gnd.n4337 19.3944
R16297 gnd.n4347 gnd.n4335 19.3944
R16298 gnd.n4351 gnd.n4335 19.3944
R16299 gnd.n4351 gnd.n4333 19.3944
R16300 gnd.n4357 gnd.n4333 19.3944
R16301 gnd.n4357 gnd.n4331 19.3944
R16302 gnd.n4361 gnd.n4331 19.3944
R16303 gnd.n4361 gnd.n4329 19.3944
R16304 gnd.n4367 gnd.n4329 19.3944
R16305 gnd.n4367 gnd.n4327 19.3944
R16306 gnd.n4371 gnd.n4327 19.3944
R16307 gnd.n4371 gnd.n4325 19.3944
R16308 gnd.n4377 gnd.n4325 19.3944
R16309 gnd.n4377 gnd.n4323 19.3944
R16310 gnd.n4384 gnd.n4323 19.3944
R16311 gnd.n4390 gnd.n4321 19.3944
R16312 gnd.n4390 gnd.n4319 19.3944
R16313 gnd.n4394 gnd.n4319 19.3944
R16314 gnd.n4394 gnd.n4317 19.3944
R16315 gnd.n4400 gnd.n4317 19.3944
R16316 gnd.n4400 gnd.n4315 19.3944
R16317 gnd.n4405 gnd.n4315 19.3944
R16318 gnd.n4413 gnd.n1966 19.3944
R16319 gnd.n4413 gnd.n1964 19.3944
R16320 gnd.n4417 gnd.n1964 19.3944
R16321 gnd.n4417 gnd.n1962 19.3944
R16322 gnd.n4423 gnd.n1962 19.3944
R16323 gnd.n4423 gnd.n1960 19.3944
R16324 gnd.n4427 gnd.n1960 19.3944
R16325 gnd.n4427 gnd.n1958 19.3944
R16326 gnd.n4439 gnd.n1956 19.3944
R16327 gnd.n4439 gnd.n1954 19.3944
R16328 gnd.n4445 gnd.n1954 19.3944
R16329 gnd.n4445 gnd.n1952 19.3944
R16330 gnd.n4449 gnd.n1952 19.3944
R16331 gnd.n4449 gnd.n1950 19.3944
R16332 gnd.n4455 gnd.n1950 19.3944
R16333 gnd.n4455 gnd.n1948 19.3944
R16334 gnd.n4459 gnd.n1948 19.3944
R16335 gnd.n4459 gnd.n1946 19.3944
R16336 gnd.n4465 gnd.n1946 19.3944
R16337 gnd.n4465 gnd.n1944 19.3944
R16338 gnd.n4469 gnd.n1944 19.3944
R16339 gnd.n4469 gnd.n1942 19.3944
R16340 gnd.n4475 gnd.n1942 19.3944
R16341 gnd.n4475 gnd.n1940 19.3944
R16342 gnd.n4480 gnd.n1940 19.3944
R16343 gnd.n4480 gnd.n1938 19.3944
R16344 gnd.n4493 gnd.n1931 19.3944
R16345 gnd.n4494 gnd.n4493 19.3944
R16346 gnd.n4495 gnd.n4494 19.3944
R16347 gnd.n4495 gnd.n1926 19.3944
R16348 gnd.n4507 gnd.n1926 19.3944
R16349 gnd.n4508 gnd.n4507 19.3944
R16350 gnd.n4509 gnd.n4508 19.3944
R16351 gnd.n4509 gnd.n1889 19.3944
R16352 gnd.n4521 gnd.n1889 19.3944
R16353 gnd.n4522 gnd.n4521 19.3944
R16354 gnd.n4523 gnd.n4522 19.3944
R16355 gnd.n4524 gnd.n4523 19.3944
R16356 gnd.n4528 gnd.n4524 19.3944
R16357 gnd.n4529 gnd.n4528 19.3944
R16358 gnd.n4533 gnd.n4529 19.3944
R16359 gnd.n4534 gnd.n4533 19.3944
R16360 gnd.n4536 gnd.n4534 19.3944
R16361 gnd.n4536 gnd.n1867 19.3944
R16362 gnd.n4581 gnd.n1867 19.3944
R16363 gnd.n4582 gnd.n4581 19.3944
R16364 gnd.n4607 gnd.n4582 19.3944
R16365 gnd.n4607 gnd.n4606 19.3944
R16366 gnd.n4606 gnd.n4605 19.3944
R16367 gnd.n4605 gnd.n4604 19.3944
R16368 gnd.n4604 gnd.n4603 19.3944
R16369 gnd.n4603 gnd.n4602 19.3944
R16370 gnd.n4602 gnd.n4586 19.3944
R16371 gnd.n4591 gnd.n4586 19.3944
R16372 gnd.n4591 gnd.n388 19.3944
R16373 gnd.n7580 gnd.n388 19.3944
R16374 gnd.n7581 gnd.n7580 19.3944
R16375 gnd.n7582 gnd.n7581 19.3944
R16376 gnd.n7582 gnd.n382 19.3944
R16377 gnd.n7594 gnd.n382 19.3944
R16378 gnd.n7595 gnd.n7594 19.3944
R16379 gnd.n7596 gnd.n7595 19.3944
R16380 gnd.n7596 gnd.n376 19.3944
R16381 gnd.n7608 gnd.n376 19.3944
R16382 gnd.n7609 gnd.n7608 19.3944
R16383 gnd.n7610 gnd.n7609 19.3944
R16384 gnd.n7610 gnd.n370 19.3944
R16385 gnd.n7622 gnd.n370 19.3944
R16386 gnd.n7623 gnd.n7622 19.3944
R16387 gnd.n7624 gnd.n7623 19.3944
R16388 gnd.n7624 gnd.n364 19.3944
R16389 gnd.n7636 gnd.n364 19.3944
R16390 gnd.n7637 gnd.n7636 19.3944
R16391 gnd.n7638 gnd.n7637 19.3944
R16392 gnd.n7638 gnd.n359 19.3944
R16393 gnd.n7651 gnd.n359 19.3944
R16394 gnd.n7652 gnd.n7651 19.3944
R16395 gnd.n7654 gnd.n7652 19.3944
R16396 gnd.n7654 gnd.n7653 19.3944
R16397 gnd.n4490 gnd.n1742 19.3944
R16398 gnd.n4702 gnd.n1742 19.3944
R16399 gnd.n4702 gnd.n4701 19.3944
R16400 gnd.n4701 gnd.n4700 19.3944
R16401 gnd.n4700 gnd.n1746 19.3944
R16402 gnd.n4690 gnd.n1746 19.3944
R16403 gnd.n4690 gnd.n4689 19.3944
R16404 gnd.n4689 gnd.n4688 19.3944
R16405 gnd.n4688 gnd.n1766 19.3944
R16406 gnd.n4678 gnd.n1766 19.3944
R16407 gnd.n4678 gnd.n4677 19.3944
R16408 gnd.n4677 gnd.n4676 19.3944
R16409 gnd.n4676 gnd.n1787 19.3944
R16410 gnd.n4666 gnd.n1787 19.3944
R16411 gnd.n4666 gnd.n4665 19.3944
R16412 gnd.n4665 gnd.n4664 19.3944
R16413 gnd.n4664 gnd.n1806 19.3944
R16414 gnd.n4654 gnd.n1806 19.3944
R16415 gnd.n4654 gnd.n4653 19.3944
R16416 gnd.n4653 gnd.n4652 19.3944
R16417 gnd.n4652 gnd.n1827 19.3944
R16418 gnd.n4642 gnd.n1827 19.3944
R16419 gnd.n4642 gnd.n4641 19.3944
R16420 gnd.n4641 gnd.n4640 19.3944
R16421 gnd.n4640 gnd.n1844 19.3944
R16422 gnd.n4589 gnd.n1844 19.3944
R16423 gnd.n4597 gnd.n4589 19.3944
R16424 gnd.n4597 gnd.n4596 19.3944
R16425 gnd.n4596 gnd.n4595 19.3944
R16426 gnd.n4595 gnd.n108 19.3944
R16427 gnd.n7871 gnd.n108 19.3944
R16428 gnd.n7871 gnd.n7870 19.3944
R16429 gnd.n7870 gnd.n7869 19.3944
R16430 gnd.n7869 gnd.n112 19.3944
R16431 gnd.n7859 gnd.n112 19.3944
R16432 gnd.n7859 gnd.n7858 19.3944
R16433 gnd.n7858 gnd.n7857 19.3944
R16434 gnd.n7857 gnd.n130 19.3944
R16435 gnd.n7847 gnd.n130 19.3944
R16436 gnd.n7847 gnd.n7846 19.3944
R16437 gnd.n7846 gnd.n7845 19.3944
R16438 gnd.n7845 gnd.n151 19.3944
R16439 gnd.n7835 gnd.n151 19.3944
R16440 gnd.n7835 gnd.n7834 19.3944
R16441 gnd.n7834 gnd.n7833 19.3944
R16442 gnd.n7833 gnd.n170 19.3944
R16443 gnd.n7823 gnd.n170 19.3944
R16444 gnd.n7823 gnd.n7822 19.3944
R16445 gnd.n7822 gnd.n7821 19.3944
R16446 gnd.n7821 gnd.n191 19.3944
R16447 gnd.n7811 gnd.n191 19.3944
R16448 gnd.n7811 gnd.n7810 19.3944
R16449 gnd.n7810 gnd.n7809 19.3944
R16450 gnd.n7731 gnd.n283 19.3944
R16451 gnd.n7731 gnd.n287 19.3944
R16452 gnd.n290 gnd.n287 19.3944
R16453 gnd.n7724 gnd.n290 19.3944
R16454 gnd.n7724 gnd.n7723 19.3944
R16455 gnd.n7723 gnd.n7722 19.3944
R16456 gnd.n7722 gnd.n296 19.3944
R16457 gnd.n7717 gnd.n296 19.3944
R16458 gnd.n7717 gnd.n7716 19.3944
R16459 gnd.n7716 gnd.n7715 19.3944
R16460 gnd.n7715 gnd.n303 19.3944
R16461 gnd.n7710 gnd.n303 19.3944
R16462 gnd.n7710 gnd.n7709 19.3944
R16463 gnd.n7709 gnd.n7708 19.3944
R16464 gnd.n7708 gnd.n310 19.3944
R16465 gnd.n7703 gnd.n310 19.3944
R16466 gnd.n7703 gnd.n7702 19.3944
R16467 gnd.n7702 gnd.n7701 19.3944
R16468 gnd.n7769 gnd.n250 19.3944
R16469 gnd.n7764 gnd.n250 19.3944
R16470 gnd.n7764 gnd.n7763 19.3944
R16471 gnd.n7763 gnd.n7762 19.3944
R16472 gnd.n7762 gnd.n257 19.3944
R16473 gnd.n7757 gnd.n257 19.3944
R16474 gnd.n7757 gnd.n7756 19.3944
R16475 gnd.n7756 gnd.n7755 19.3944
R16476 gnd.n7755 gnd.n264 19.3944
R16477 gnd.n7750 gnd.n264 19.3944
R16478 gnd.n7750 gnd.n7749 19.3944
R16479 gnd.n7749 gnd.n7748 19.3944
R16480 gnd.n7748 gnd.n271 19.3944
R16481 gnd.n7743 gnd.n271 19.3944
R16482 gnd.n7743 gnd.n7742 19.3944
R16483 gnd.n7742 gnd.n7741 19.3944
R16484 gnd.n7741 gnd.n278 19.3944
R16485 gnd.n7736 gnd.n278 19.3944
R16486 gnd.n7802 gnd.n7801 19.3944
R16487 gnd.n7801 gnd.n7800 19.3944
R16488 gnd.n7800 gnd.n221 19.3944
R16489 gnd.n7795 gnd.n221 19.3944
R16490 gnd.n7795 gnd.n7794 19.3944
R16491 gnd.n7794 gnd.n7793 19.3944
R16492 gnd.n7793 gnd.n229 19.3944
R16493 gnd.n7788 gnd.n229 19.3944
R16494 gnd.n7788 gnd.n7787 19.3944
R16495 gnd.n7787 gnd.n7786 19.3944
R16496 gnd.n7786 gnd.n236 19.3944
R16497 gnd.n7781 gnd.n236 19.3944
R16498 gnd.n7781 gnd.n7780 19.3944
R16499 gnd.n7780 gnd.n7779 19.3944
R16500 gnd.n7779 gnd.n243 19.3944
R16501 gnd.n7774 gnd.n243 19.3944
R16502 gnd.n7774 gnd.n7773 19.3944
R16503 gnd.n7692 gnd.n7691 19.3944
R16504 gnd.n7691 gnd.n7690 19.3944
R16505 gnd.n7690 gnd.n325 19.3944
R16506 gnd.n7685 gnd.n325 19.3944
R16507 gnd.n7685 gnd.n7684 19.3944
R16508 gnd.n7684 gnd.n7683 19.3944
R16509 gnd.n7683 gnd.n332 19.3944
R16510 gnd.n7678 gnd.n332 19.3944
R16511 gnd.n7678 gnd.n7677 19.3944
R16512 gnd.n7677 gnd.n7676 19.3944
R16513 gnd.n7676 gnd.n339 19.3944
R16514 gnd.n7671 gnd.n339 19.3944
R16515 gnd.n7671 gnd.n7670 19.3944
R16516 gnd.n7670 gnd.n7669 19.3944
R16517 gnd.n7669 gnd.n346 19.3944
R16518 gnd.n7664 gnd.n346 19.3944
R16519 gnd.n3928 gnd.n3927 19.3944
R16520 gnd.n3927 gnd.n1930 19.3944
R16521 gnd.n4499 gnd.n1930 19.3944
R16522 gnd.n4499 gnd.n1928 19.3944
R16523 gnd.n4503 gnd.n1928 19.3944
R16524 gnd.n4503 gnd.n1893 19.3944
R16525 gnd.n4513 gnd.n1893 19.3944
R16526 gnd.n4513 gnd.n1891 19.3944
R16527 gnd.n4517 gnd.n1891 19.3944
R16528 gnd.n4517 gnd.n1881 19.3944
R16529 gnd.n4553 gnd.n1881 19.3944
R16530 gnd.n4553 gnd.n1882 19.3944
R16531 gnd.n4549 gnd.n1882 19.3944
R16532 gnd.n4549 gnd.n4548 19.3944
R16533 gnd.n4548 gnd.n4547 19.3944
R16534 gnd.n4547 gnd.n1887 19.3944
R16535 gnd.n4543 gnd.n1887 19.3944
R16536 gnd.n4543 gnd.n4542 19.3944
R16537 gnd.n4542 gnd.n4541 19.3944
R16538 gnd.n4541 gnd.n1866 19.3944
R16539 gnd.n4611 gnd.n1866 19.3944
R16540 gnd.n4611 gnd.n1863 19.3944
R16541 gnd.n4618 gnd.n1863 19.3944
R16542 gnd.n4618 gnd.n1864 19.3944
R16543 gnd.n4614 gnd.n1864 19.3944
R16544 gnd.n4614 gnd.n81 19.3944
R16545 gnd.n7884 gnd.n81 19.3944
R16546 gnd.n7884 gnd.n7883 19.3944
R16547 gnd.n7883 gnd.n83 19.3944
R16548 gnd.n7576 gnd.n83 19.3944
R16549 gnd.n7576 gnd.n387 19.3944
R16550 gnd.n7586 gnd.n387 19.3944
R16551 gnd.n7586 gnd.n385 19.3944
R16552 gnd.n7590 gnd.n385 19.3944
R16553 gnd.n7590 gnd.n380 19.3944
R16554 gnd.n7600 gnd.n380 19.3944
R16555 gnd.n7600 gnd.n378 19.3944
R16556 gnd.n7604 gnd.n378 19.3944
R16557 gnd.n7604 gnd.n375 19.3944
R16558 gnd.n7614 gnd.n375 19.3944
R16559 gnd.n7614 gnd.n373 19.3944
R16560 gnd.n7618 gnd.n373 19.3944
R16561 gnd.n7618 gnd.n368 19.3944
R16562 gnd.n7628 gnd.n368 19.3944
R16563 gnd.n7628 gnd.n366 19.3944
R16564 gnd.n7632 gnd.n366 19.3944
R16565 gnd.n7632 gnd.n363 19.3944
R16566 gnd.n7642 gnd.n363 19.3944
R16567 gnd.n7642 gnd.n361 19.3944
R16568 gnd.n7647 gnd.n361 19.3944
R16569 gnd.n7647 gnd.n357 19.3944
R16570 gnd.n7658 gnd.n357 19.3944
R16571 gnd.n7659 gnd.n7658 19.3944
R16572 gnd.n4708 gnd.n4707 19.3944
R16573 gnd.n4707 gnd.n4706 19.3944
R16574 gnd.n4706 gnd.n1734 19.3944
R16575 gnd.n4696 gnd.n1734 19.3944
R16576 gnd.n4696 gnd.n4695 19.3944
R16577 gnd.n4695 gnd.n4694 19.3944
R16578 gnd.n4694 gnd.n1757 19.3944
R16579 gnd.n4684 gnd.n1757 19.3944
R16580 gnd.n4684 gnd.n4683 19.3944
R16581 gnd.n4683 gnd.n4682 19.3944
R16582 gnd.n4682 gnd.n1777 19.3944
R16583 gnd.n4672 gnd.n1777 19.3944
R16584 gnd.n4672 gnd.n4671 19.3944
R16585 gnd.n4671 gnd.n4670 19.3944
R16586 gnd.n4670 gnd.n1797 19.3944
R16587 gnd.n4660 gnd.n1797 19.3944
R16588 gnd.n4660 gnd.n4659 19.3944
R16589 gnd.n4659 gnd.n4658 19.3944
R16590 gnd.n4658 gnd.n1817 19.3944
R16591 gnd.n4648 gnd.n1817 19.3944
R16592 gnd.n4648 gnd.n4647 19.3944
R16593 gnd.n4647 gnd.n4646 19.3944
R16594 gnd.n1835 gnd.n97 19.3944
R16595 gnd.n1853 gnd.n97 19.3944
R16596 gnd.n1851 gnd.n1850 19.3944
R16597 gnd.n7879 gnd.n7878 19.3944
R16598 gnd.n7875 gnd.n92 19.3944
R16599 gnd.n7875 gnd.n99 19.3944
R16600 gnd.n7865 gnd.n99 19.3944
R16601 gnd.n7865 gnd.n7864 19.3944
R16602 gnd.n7864 gnd.n7863 19.3944
R16603 gnd.n7863 gnd.n121 19.3944
R16604 gnd.n7853 gnd.n121 19.3944
R16605 gnd.n7853 gnd.n7852 19.3944
R16606 gnd.n7852 gnd.n7851 19.3944
R16607 gnd.n7851 gnd.n141 19.3944
R16608 gnd.n7841 gnd.n141 19.3944
R16609 gnd.n7841 gnd.n7840 19.3944
R16610 gnd.n7840 gnd.n7839 19.3944
R16611 gnd.n7839 gnd.n161 19.3944
R16612 gnd.n7829 gnd.n161 19.3944
R16613 gnd.n7829 gnd.n7828 19.3944
R16614 gnd.n7828 gnd.n7827 19.3944
R16615 gnd.n7827 gnd.n181 19.3944
R16616 gnd.n7817 gnd.n181 19.3944
R16617 gnd.n7817 gnd.n7816 19.3944
R16618 gnd.n7816 gnd.n7815 19.3944
R16619 gnd.n7815 gnd.n202 19.3944
R16620 gnd.n7805 gnd.n202 19.3944
R16621 gnd.n5230 gnd.n5229 19.3944
R16622 gnd.n5229 gnd.n1129 19.3944
R16623 gnd.n2804 gnd.n1129 19.3944
R16624 gnd.n2804 gnd.n2801 19.3944
R16625 gnd.n2808 gnd.n2801 19.3944
R16626 gnd.n2808 gnd.n2799 19.3944
R16627 gnd.n2812 gnd.n2799 19.3944
R16628 gnd.n2812 gnd.n2797 19.3944
R16629 gnd.n2835 gnd.n2797 19.3944
R16630 gnd.n2835 gnd.n2834 19.3944
R16631 gnd.n2834 gnd.n2833 19.3944
R16632 gnd.n2833 gnd.n2818 19.3944
R16633 gnd.n2829 gnd.n2818 19.3944
R16634 gnd.n2829 gnd.n2828 19.3944
R16635 gnd.n2828 gnd.n2827 19.3944
R16636 gnd.n2827 gnd.n2825 19.3944
R16637 gnd.n2825 gnd.n2699 19.3944
R16638 gnd.n2905 gnd.n2699 19.3944
R16639 gnd.n2905 gnd.n2697 19.3944
R16640 gnd.n2909 gnd.n2697 19.3944
R16641 gnd.n2909 gnd.n2695 19.3944
R16642 gnd.n2914 gnd.n2695 19.3944
R16643 gnd.n2914 gnd.n2693 19.3944
R16644 gnd.n2918 gnd.n2693 19.3944
R16645 gnd.n2929 gnd.n2918 19.3944
R16646 gnd.n2927 gnd.n2926 19.3944
R16647 gnd.n2923 gnd.n2922 19.3944
R16648 gnd.n2981 gnd.n2652 19.3944
R16649 gnd.n3004 gnd.n2983 19.3944
R16650 gnd.n3002 gnd.n3001 19.3944
R16651 gnd.n3001 gnd.n2985 19.3944
R16652 gnd.n2997 gnd.n2985 19.3944
R16653 gnd.n2997 gnd.n2996 19.3944
R16654 gnd.n2996 gnd.n2995 19.3944
R16655 gnd.n2995 gnd.n2993 19.3944
R16656 gnd.n2993 gnd.n2628 19.3944
R16657 gnd.n2628 gnd.n2626 19.3944
R16658 gnd.n3071 gnd.n2626 19.3944
R16659 gnd.n3071 gnd.n2624 19.3944
R16660 gnd.n3075 gnd.n2624 19.3944
R16661 gnd.n3075 gnd.n2622 19.3944
R16662 gnd.n3079 gnd.n2622 19.3944
R16663 gnd.n3079 gnd.n2620 19.3944
R16664 gnd.n3115 gnd.n2620 19.3944
R16665 gnd.n3115 gnd.n3114 19.3944
R16666 gnd.n3114 gnd.n3113 19.3944
R16667 gnd.n3113 gnd.n3085 19.3944
R16668 gnd.n3109 gnd.n3085 19.3944
R16669 gnd.n3109 gnd.n3108 19.3944
R16670 gnd.n3108 gnd.n3107 19.3944
R16671 gnd.n3107 gnd.n3091 19.3944
R16672 gnd.n3102 gnd.n3091 19.3944
R16673 gnd.n3102 gnd.n3101 19.3944
R16674 gnd.n3101 gnd.n3100 19.3944
R16675 gnd.n3100 gnd.n2396 19.3944
R16676 gnd.n3225 gnd.n2396 19.3944
R16677 gnd.n3225 gnd.n2394 19.3944
R16678 gnd.n3231 gnd.n2394 19.3944
R16679 gnd.n3231 gnd.n3230 19.3944
R16680 gnd.n3230 gnd.n2372 19.3944
R16681 gnd.n3255 gnd.n2372 19.3944
R16682 gnd.n3255 gnd.n2370 19.3944
R16683 gnd.n3261 gnd.n2370 19.3944
R16684 gnd.n3261 gnd.n3260 19.3944
R16685 gnd.n3260 gnd.n2347 19.3944
R16686 gnd.n3287 gnd.n2347 19.3944
R16687 gnd.n3287 gnd.n2345 19.3944
R16688 gnd.n3297 gnd.n2345 19.3944
R16689 gnd.n3297 gnd.n3296 19.3944
R16690 gnd.n3296 gnd.n3295 19.3944
R16691 gnd.n3295 gnd.n1602 19.3944
R16692 gnd.n4838 gnd.n1602 19.3944
R16693 gnd.n4838 gnd.n4837 19.3944
R16694 gnd.n4837 gnd.n4836 19.3944
R16695 gnd.n4836 gnd.n1606 19.3944
R16696 gnd.n2317 gnd.n1606 19.3944
R16697 gnd.n3454 gnd.n2317 19.3944
R16698 gnd.n3454 gnd.n2314 19.3944
R16699 gnd.n3458 gnd.n2314 19.3944
R16700 gnd.n3458 gnd.n2294 19.3944
R16701 gnd.n3481 gnd.n2294 19.3944
R16702 gnd.n3481 gnd.n2292 19.3944
R16703 gnd.n3487 gnd.n2292 19.3944
R16704 gnd.n3487 gnd.n3486 19.3944
R16705 gnd.n3486 gnd.n2261 19.3944
R16706 gnd.n3523 gnd.n2261 19.3944
R16707 gnd.n3523 gnd.n2259 19.3944
R16708 gnd.n3538 gnd.n2259 19.3944
R16709 gnd.n3538 gnd.n3537 19.3944
R16710 gnd.n3537 gnd.n3536 19.3944
R16711 gnd.n3536 gnd.n3530 19.3944
R16712 gnd.n3530 gnd.n2227 19.3944
R16713 gnd.n3606 gnd.n2227 19.3944
R16714 gnd.n3606 gnd.n2225 19.3944
R16715 gnd.n3610 gnd.n2225 19.3944
R16716 gnd.n3610 gnd.n2204 19.3944
R16717 gnd.n3649 gnd.n2204 19.3944
R16718 gnd.n3649 gnd.n2202 19.3944
R16719 gnd.n3653 gnd.n2202 19.3944
R16720 gnd.n3653 gnd.n2188 19.3944
R16721 gnd.n3693 gnd.n2188 19.3944
R16722 gnd.n3693 gnd.n2186 19.3944
R16723 gnd.n3699 gnd.n2186 19.3944
R16724 gnd.n3699 gnd.n3698 19.3944
R16725 gnd.n3698 gnd.n2157 19.3944
R16726 gnd.n3739 gnd.n2157 19.3944
R16727 gnd.n3739 gnd.n2155 19.3944
R16728 gnd.n3743 gnd.n2155 19.3944
R16729 gnd.n3743 gnd.n2140 19.3944
R16730 gnd.n3800 gnd.n2140 19.3944
R16731 gnd.n3800 gnd.n2138 19.3944
R16732 gnd.n3804 gnd.n2138 19.3944
R16733 gnd.n3804 gnd.n2118 19.3944
R16734 gnd.n3828 gnd.n2118 19.3944
R16735 gnd.n3828 gnd.n2116 19.3944
R16736 gnd.n3834 gnd.n2116 19.3944
R16737 gnd.n3834 gnd.n3833 19.3944
R16738 gnd.n3833 gnd.n2090 19.3944
R16739 gnd.n3872 gnd.n2090 19.3944
R16740 gnd.n3872 gnd.n2088 19.3944
R16741 gnd.n3882 gnd.n2088 19.3944
R16742 gnd.n3882 gnd.n3881 19.3944
R16743 gnd.n3881 gnd.n3880 19.3944
R16744 gnd.n3880 gnd.n2020 19.3944
R16745 gnd.n4147 gnd.n2020 19.3944
R16746 gnd.n4147 gnd.n4146 19.3944
R16747 gnd.n4146 gnd.n4145 19.3944
R16748 gnd.n4145 gnd.n2024 19.3944
R16749 gnd.n4136 gnd.n2024 19.3944
R16750 gnd.n4136 gnd.n4135 19.3944
R16751 gnd.n4135 gnd.n4134 19.3944
R16752 gnd.n4134 gnd.n2034 19.3944
R16753 gnd.n4125 gnd.n2034 19.3944
R16754 gnd.n4125 gnd.n4124 19.3944
R16755 gnd.n4124 gnd.n4123 19.3944
R16756 gnd.n4123 gnd.n2045 19.3944
R16757 gnd.n4114 gnd.n2045 19.3944
R16758 gnd.n4114 gnd.n4113 19.3944
R16759 gnd.n4113 gnd.n1709 19.3944
R16760 gnd.n4723 gnd.n1709 19.3944
R16761 gnd.n4723 gnd.n4722 19.3944
R16762 gnd.n4722 gnd.n4721 19.3944
R16763 gnd.n4721 gnd.n1713 19.3944
R16764 gnd.n4715 gnd.n1713 19.3944
R16765 gnd.n4715 gnd.n4714 19.3944
R16766 gnd.n4714 gnd.n4713 19.3944
R16767 gnd.n4713 gnd.n1722 19.3944
R16768 gnd.n1900 gnd.n1722 19.3944
R16769 gnd.n1904 gnd.n1900 19.3944
R16770 gnd.n1904 gnd.n1898 19.3944
R16771 gnd.n1908 gnd.n1898 19.3944
R16772 gnd.n1908 gnd.n1896 19.3944
R16773 gnd.n1923 gnd.n1896 19.3944
R16774 gnd.n1923 gnd.n1922 19.3944
R16775 gnd.n1922 gnd.n1921 19.3944
R16776 gnd.n1921 gnd.n1918 19.3944
R16777 gnd.n1918 gnd.n1917 19.3944
R16778 gnd.n1917 gnd.n1879 19.3944
R16779 gnd.n1879 gnd.n1877 19.3944
R16780 gnd.n4560 gnd.n1877 19.3944
R16781 gnd.n4560 gnd.n1875 19.3944
R16782 gnd.n4564 gnd.n1875 19.3944
R16783 gnd.n4564 gnd.n1873 19.3944
R16784 gnd.n4568 gnd.n1873 19.3944
R16785 gnd.n4568 gnd.n1871 19.3944
R16786 gnd.n4576 gnd.n1871 19.3944
R16787 gnd.n4576 gnd.n4575 19.3944
R16788 gnd.n4575 gnd.n4574 19.3944
R16789 gnd.n4624 gnd.n1860 19.3944
R16790 gnd.n4632 gnd.n4626 19.3944
R16791 gnd.n4630 gnd.n4629 19.3944
R16792 gnd.n7571 gnd.n394 19.3944
R16793 gnd.n7569 gnd.n7568 19.3944
R16794 gnd.n7568 gnd.n396 19.3944
R16795 gnd.n7564 gnd.n396 19.3944
R16796 gnd.n7564 gnd.n7563 19.3944
R16797 gnd.n7563 gnd.n7562 19.3944
R16798 gnd.n7562 gnd.n402 19.3944
R16799 gnd.n7558 gnd.n402 19.3944
R16800 gnd.n7558 gnd.n7557 19.3944
R16801 gnd.n7557 gnd.n7556 19.3944
R16802 gnd.n7556 gnd.n408 19.3944
R16803 gnd.n7552 gnd.n408 19.3944
R16804 gnd.n7552 gnd.n7551 19.3944
R16805 gnd.n7551 gnd.n7550 19.3944
R16806 gnd.n7550 gnd.n414 19.3944
R16807 gnd.n7546 gnd.n414 19.3944
R16808 gnd.n7546 gnd.n7545 19.3944
R16809 gnd.n7545 gnd.n7544 19.3944
R16810 gnd.n7544 gnd.n420 19.3944
R16811 gnd.n7540 gnd.n420 19.3944
R16812 gnd.n7540 gnd.n7539 19.3944
R16813 gnd.n7539 gnd.n7538 19.3944
R16814 gnd.n7538 gnd.n426 19.3944
R16815 gnd.n7534 gnd.n426 19.3944
R16816 gnd.n7534 gnd.n7533 19.3944
R16817 gnd.n7533 gnd.n7532 19.3944
R16818 gnd.n5223 gnd.n5222 19.3944
R16819 gnd.n5222 gnd.n5221 19.3944
R16820 gnd.n5221 gnd.n5220 19.3944
R16821 gnd.n5220 gnd.n5218 19.3944
R16822 gnd.n5218 gnd.n5215 19.3944
R16823 gnd.n5215 gnd.n5214 19.3944
R16824 gnd.n5214 gnd.n5211 19.3944
R16825 gnd.n5211 gnd.n5210 19.3944
R16826 gnd.n5210 gnd.n5207 19.3944
R16827 gnd.n5207 gnd.n5206 19.3944
R16828 gnd.n5206 gnd.n5203 19.3944
R16829 gnd.n5203 gnd.n5202 19.3944
R16830 gnd.n5202 gnd.n5199 19.3944
R16831 gnd.n5199 gnd.n5198 19.3944
R16832 gnd.n5198 gnd.n5195 19.3944
R16833 gnd.n5195 gnd.n5194 19.3944
R16834 gnd.n5194 gnd.n5191 19.3944
R16835 gnd.n5189 gnd.n5186 19.3944
R16836 gnd.n5186 gnd.n5185 19.3944
R16837 gnd.n5185 gnd.n5182 19.3944
R16838 gnd.n5182 gnd.n5181 19.3944
R16839 gnd.n5181 gnd.n5178 19.3944
R16840 gnd.n5178 gnd.n5177 19.3944
R16841 gnd.n5177 gnd.n5174 19.3944
R16842 gnd.n5174 gnd.n5173 19.3944
R16843 gnd.n5173 gnd.n5170 19.3944
R16844 gnd.n5170 gnd.n5169 19.3944
R16845 gnd.n5169 gnd.n5166 19.3944
R16846 gnd.n5166 gnd.n5165 19.3944
R16847 gnd.n5165 gnd.n5162 19.3944
R16848 gnd.n5162 gnd.n5161 19.3944
R16849 gnd.n5161 gnd.n5158 19.3944
R16850 gnd.n5158 gnd.n5157 19.3944
R16851 gnd.n5157 gnd.n5154 19.3944
R16852 gnd.n5154 gnd.n5153 19.3944
R16853 gnd.n5149 gnd.n5146 19.3944
R16854 gnd.n5146 gnd.n5145 19.3944
R16855 gnd.n5145 gnd.n5142 19.3944
R16856 gnd.n5142 gnd.n5141 19.3944
R16857 gnd.n5141 gnd.n5138 19.3944
R16858 gnd.n5138 gnd.n5137 19.3944
R16859 gnd.n5137 gnd.n5134 19.3944
R16860 gnd.n5134 gnd.n5133 19.3944
R16861 gnd.n5133 gnd.n5130 19.3944
R16862 gnd.n5130 gnd.n5129 19.3944
R16863 gnd.n5129 gnd.n5126 19.3944
R16864 gnd.n5126 gnd.n5125 19.3944
R16865 gnd.n5125 gnd.n5122 19.3944
R16866 gnd.n5122 gnd.n5121 19.3944
R16867 gnd.n5121 gnd.n5118 19.3944
R16868 gnd.n5118 gnd.n5117 19.3944
R16869 gnd.n5117 gnd.n5114 19.3944
R16870 gnd.n5114 gnd.n5113 19.3944
R16871 gnd.n2733 gnd.n2732 19.3944
R16872 gnd.n2736 gnd.n2733 19.3944
R16873 gnd.n2736 gnd.n2730 19.3944
R16874 gnd.n2742 gnd.n2730 19.3944
R16875 gnd.n2743 gnd.n2742 19.3944
R16876 gnd.n2746 gnd.n2743 19.3944
R16877 gnd.n2746 gnd.n2728 19.3944
R16878 gnd.n2752 gnd.n2728 19.3944
R16879 gnd.n2753 gnd.n2752 19.3944
R16880 gnd.n2756 gnd.n2753 19.3944
R16881 gnd.n2756 gnd.n2726 19.3944
R16882 gnd.n2762 gnd.n2726 19.3944
R16883 gnd.n2763 gnd.n2762 19.3944
R16884 gnd.n2766 gnd.n2763 19.3944
R16885 gnd.n2766 gnd.n2722 19.3944
R16886 gnd.n2770 gnd.n2722 19.3944
R16887 gnd.n2776 gnd.n2775 19.3944
R16888 gnd.n2782 gnd.n2776 19.3944
R16889 gnd.n2782 gnd.n2716 19.3944
R16890 gnd.n2786 gnd.n2716 19.3944
R16891 gnd.n2786 gnd.n2714 19.3944
R16892 gnd.n2840 gnd.n2714 19.3944
R16893 gnd.n2840 gnd.n2712 19.3944
R16894 gnd.n2844 gnd.n2712 19.3944
R16895 gnd.n2844 gnd.n2710 19.3944
R16896 gnd.n2855 gnd.n2710 19.3944
R16897 gnd.n2855 gnd.n2708 19.3944
R16898 gnd.n2860 gnd.n2708 19.3944
R16899 gnd.n2860 gnd.n2702 19.3944
R16900 gnd.n2899 gnd.n2702 19.3944
R16901 gnd.n2899 gnd.n2898 19.3944
R16902 gnd.n2898 gnd.n2897 19.3944
R16903 gnd.n2897 gnd.n2706 19.3944
R16904 gnd.n2887 gnd.n2706 19.3944
R16905 gnd.n2887 gnd.n2886 19.3944
R16906 gnd.n2886 gnd.n2885 19.3944
R16907 gnd.n2885 gnd.n2879 19.3944
R16908 gnd.n2879 gnd.n2878 19.3944
R16909 gnd.n2878 gnd.n2676 19.3944
R16910 gnd.n2947 gnd.n2676 19.3944
R16911 gnd.n2947 gnd.n2674 19.3944
R16912 gnd.n2957 gnd.n2674 19.3944
R16913 gnd.n2957 gnd.n2956 19.3944
R16914 gnd.n2956 gnd.n2952 19.3944
R16915 gnd.n2952 gnd.n2646 19.3944
R16916 gnd.n3009 gnd.n2646 19.3944
R16917 gnd.n3009 gnd.n2644 19.3944
R16918 gnd.n3013 gnd.n2644 19.3944
R16919 gnd.n3013 gnd.n2641 19.3944
R16920 gnd.n3024 gnd.n2641 19.3944
R16921 gnd.n3024 gnd.n2639 19.3944
R16922 gnd.n3028 gnd.n2639 19.3944
R16923 gnd.n3028 gnd.n2630 19.3944
R16924 gnd.n3064 gnd.n2630 19.3944
R16925 gnd.n3064 gnd.n2631 19.3944
R16926 gnd.n3060 gnd.n2631 19.3944
R16927 gnd.n3060 gnd.n3059 19.3944
R16928 gnd.n3059 gnd.n3058 19.3944
R16929 gnd.n3058 gnd.n2636 19.3944
R16930 gnd.n3054 gnd.n2636 19.3944
R16931 gnd.n3054 gnd.n3053 19.3944
R16932 gnd.n3053 gnd.n3052 19.3944
R16933 gnd.n3052 gnd.n2614 19.3944
R16934 gnd.n3126 gnd.n2614 19.3944
R16935 gnd.n3126 gnd.n2612 19.3944
R16936 gnd.n3131 gnd.n2612 19.3944
R16937 gnd.n3131 gnd.n2609 19.3944
R16938 gnd.n3142 gnd.n2609 19.3944
R16939 gnd.n3143 gnd.n3142 19.3944
R16940 gnd.n5105 gnd.n1240 19.3944
R16941 gnd.n2778 gnd.n1240 19.3944
R16942 gnd.n2778 gnd.n2715 19.3944
R16943 gnd.n2790 gnd.n2715 19.3944
R16944 gnd.n2791 gnd.n2790 19.3944
R16945 gnd.n2793 gnd.n2791 19.3944
R16946 gnd.n2793 gnd.n2711 19.3944
R16947 gnd.n2848 gnd.n2711 19.3944
R16948 gnd.n2849 gnd.n2848 19.3944
R16949 gnd.n2851 gnd.n2849 19.3944
R16950 gnd.n2851 gnd.n2707 19.3944
R16951 gnd.n2864 gnd.n2707 19.3944
R16952 gnd.n2865 gnd.n2864 19.3944
R16953 gnd.n2867 gnd.n2865 19.3944
R16954 gnd.n2868 gnd.n2867 19.3944
R16955 gnd.n2893 gnd.n2868 19.3944
R16956 gnd.n2893 gnd.n2892 19.3944
R16957 gnd.n2892 gnd.n2891 19.3944
R16958 gnd.n2891 gnd.n2870 19.3944
R16959 gnd.n2881 gnd.n2870 19.3944
R16960 gnd.n2881 gnd.n2880 19.3944
R16961 gnd.n2880 gnd.n2688 19.3944
R16962 gnd.n2936 gnd.n2688 19.3944
R16963 gnd.n2937 gnd.n2936 19.3944
R16964 gnd.n2937 gnd.n2670 19.3944
R16965 gnd.n2961 gnd.n2670 19.3944
R16966 gnd.n2962 gnd.n2961 19.3944
R16967 gnd.n2964 gnd.n2962 19.3944
R16968 gnd.n2966 gnd.n2964 19.3944
R16969 gnd.n2966 gnd.n2965 19.3944
R16970 gnd.n2965 gnd.n2643 19.3944
R16971 gnd.n3017 gnd.n2643 19.3944
R16972 gnd.n3018 gnd.n3017 19.3944
R16973 gnd.n3020 gnd.n3018 19.3944
R16974 gnd.n3020 gnd.n2638 19.3944
R16975 gnd.n3032 gnd.n2638 19.3944
R16976 gnd.n3033 gnd.n3032 19.3944
R16977 gnd.n3035 gnd.n3033 19.3944
R16978 gnd.n3036 gnd.n3035 19.3944
R16979 gnd.n3039 gnd.n3036 19.3944
R16980 gnd.n3040 gnd.n3039 19.3944
R16981 gnd.n3045 gnd.n3040 19.3944
R16982 gnd.n3046 gnd.n3045 19.3944
R16983 gnd.n3047 gnd.n3046 19.3944
R16984 gnd.n3047 gnd.n2615 19.3944
R16985 gnd.n3120 gnd.n2615 19.3944
R16986 gnd.n3121 gnd.n3120 19.3944
R16987 gnd.n3122 gnd.n3121 19.3944
R16988 gnd.n3122 gnd.n2610 19.3944
R16989 gnd.n3135 gnd.n2610 19.3944
R16990 gnd.n3136 gnd.n3135 19.3944
R16991 gnd.n3138 gnd.n3136 19.3944
R16992 gnd.n3138 gnd.n3137 19.3944
R16993 gnd.n1247 gnd.n1238 19.3944
R16994 gnd.n1263 gnd.n1247 19.3944
R16995 gnd.n5092 gnd.n1263 19.3944
R16996 gnd.n5092 gnd.n5091 19.3944
R16997 gnd.n5091 gnd.n5090 19.3944
R16998 gnd.n5090 gnd.n1267 19.3944
R16999 gnd.n5080 gnd.n1267 19.3944
R17000 gnd.n5080 gnd.n5079 19.3944
R17001 gnd.n5079 gnd.n5078 19.3944
R17002 gnd.n5078 gnd.n1287 19.3944
R17003 gnd.n5068 gnd.n1287 19.3944
R17004 gnd.n5068 gnd.n5067 19.3944
R17005 gnd.n5067 gnd.n5066 19.3944
R17006 gnd.n5066 gnd.n1308 19.3944
R17007 gnd.n5056 gnd.n1308 19.3944
R17008 gnd.n5056 gnd.n5055 19.3944
R17009 gnd.n5055 gnd.n5054 19.3944
R17010 gnd.n5054 gnd.n1328 19.3944
R17011 gnd.n5044 gnd.n1328 19.3944
R17012 gnd.n5044 gnd.n5043 19.3944
R17013 gnd.n5043 gnd.n5042 19.3944
R17014 gnd.n5042 gnd.n1349 19.3944
R17015 gnd.n2932 gnd.n1349 19.3944
R17016 gnd.n2932 gnd.n2685 19.3944
R17017 gnd.n2940 gnd.n2685 19.3944
R17018 gnd.n2940 gnd.n2666 19.3944
R17019 gnd.n2970 gnd.n2666 19.3944
R17020 gnd.n2970 gnd.n2969 19.3944
R17021 gnd.n2969 gnd.n2968 19.3944
R17022 gnd.n2968 gnd.n1374 19.3944
R17023 gnd.n5030 gnd.n1374 19.3944
R17024 gnd.n5030 gnd.n5029 19.3944
R17025 gnd.n5029 gnd.n5028 19.3944
R17026 gnd.n5028 gnd.n1378 19.3944
R17027 gnd.n5018 gnd.n1378 19.3944
R17028 gnd.n5018 gnd.n5017 19.3944
R17029 gnd.n5017 gnd.n5016 19.3944
R17030 gnd.n5016 gnd.n1397 19.3944
R17031 gnd.n5006 gnd.n1397 19.3944
R17032 gnd.n5006 gnd.n5005 19.3944
R17033 gnd.n5005 gnd.n5004 19.3944
R17034 gnd.n5004 gnd.n1417 19.3944
R17035 gnd.n4994 gnd.n1417 19.3944
R17036 gnd.n4994 gnd.n4993 19.3944
R17037 gnd.n4993 gnd.n4992 19.3944
R17038 gnd.n4992 gnd.n1437 19.3944
R17039 gnd.n4982 gnd.n1437 19.3944
R17040 gnd.n4982 gnd.n4981 19.3944
R17041 gnd.n4981 gnd.n4980 19.3944
R17042 gnd.n4980 gnd.n1457 19.3944
R17043 gnd.n4970 gnd.n1457 19.3944
R17044 gnd.n4970 gnd.n4969 19.3944
R17045 gnd.n4969 gnd.n4968 19.3944
R17046 gnd.n4961 gnd.n4960 19.3944
R17047 gnd.n4960 gnd.n1486 19.3944
R17048 gnd.n1488 gnd.n1486 19.3944
R17049 gnd.n4953 gnd.n1488 19.3944
R17050 gnd.n4953 gnd.n4952 19.3944
R17051 gnd.n4952 gnd.n4951 19.3944
R17052 gnd.n4951 gnd.n1495 19.3944
R17053 gnd.n4946 gnd.n1495 19.3944
R17054 gnd.n4946 gnd.n4945 19.3944
R17055 gnd.n4945 gnd.n4944 19.3944
R17056 gnd.n4944 gnd.n1502 19.3944
R17057 gnd.n4939 gnd.n1502 19.3944
R17058 gnd.n4939 gnd.n4938 19.3944
R17059 gnd.n4938 gnd.n4937 19.3944
R17060 gnd.n4937 gnd.n1509 19.3944
R17061 gnd.n4932 gnd.n1509 19.3944
R17062 gnd.n4932 gnd.n4931 19.3944
R17063 gnd.n2481 gnd.n2441 19.3944
R17064 gnd.n2485 gnd.n2441 19.3944
R17065 gnd.n2485 gnd.n2439 19.3944
R17066 gnd.n2491 gnd.n2439 19.3944
R17067 gnd.n2491 gnd.n2437 19.3944
R17068 gnd.n2495 gnd.n2437 19.3944
R17069 gnd.n2495 gnd.n2435 19.3944
R17070 gnd.n2501 gnd.n2435 19.3944
R17071 gnd.n2501 gnd.n2433 19.3944
R17072 gnd.n2505 gnd.n2433 19.3944
R17073 gnd.n2505 gnd.n2431 19.3944
R17074 gnd.n2511 gnd.n2431 19.3944
R17075 gnd.n2511 gnd.n2429 19.3944
R17076 gnd.n2515 gnd.n2429 19.3944
R17077 gnd.n2515 gnd.n2427 19.3944
R17078 gnd.n2521 gnd.n2427 19.3944
R17079 gnd.n2521 gnd.n2425 19.3944
R17080 gnd.n2525 gnd.n2425 19.3944
R17081 gnd.n2454 gnd.n1531 19.3944
R17082 gnd.n2461 gnd.n2454 19.3944
R17083 gnd.n2461 gnd.n2451 19.3944
R17084 gnd.n2465 gnd.n2451 19.3944
R17085 gnd.n2465 gnd.n2449 19.3944
R17086 gnd.n2471 gnd.n2449 19.3944
R17087 gnd.n2471 gnd.n2447 19.3944
R17088 gnd.n2475 gnd.n2447 19.3944
R17089 gnd.n4929 gnd.n1518 19.3944
R17090 gnd.n4924 gnd.n1518 19.3944
R17091 gnd.n4924 gnd.n4923 19.3944
R17092 gnd.n4923 gnd.n4922 19.3944
R17093 gnd.n4922 gnd.n1525 19.3944
R17094 gnd.n4917 gnd.n1525 19.3944
R17095 gnd.n4917 gnd.n4916 19.3944
R17096 gnd.n5098 gnd.n1251 19.3944
R17097 gnd.n5098 gnd.n5097 19.3944
R17098 gnd.n5097 gnd.n5096 19.3944
R17099 gnd.n5096 gnd.n1256 19.3944
R17100 gnd.n5086 gnd.n1256 19.3944
R17101 gnd.n5086 gnd.n5085 19.3944
R17102 gnd.n5085 gnd.n5084 19.3944
R17103 gnd.n5084 gnd.n1278 19.3944
R17104 gnd.n5074 gnd.n1278 19.3944
R17105 gnd.n5074 gnd.n5073 19.3944
R17106 gnd.n5073 gnd.n5072 19.3944
R17107 gnd.n5072 gnd.n1298 19.3944
R17108 gnd.n5062 gnd.n1298 19.3944
R17109 gnd.n5062 gnd.n5061 19.3944
R17110 gnd.n5061 gnd.n5060 19.3944
R17111 gnd.n5060 gnd.n1319 19.3944
R17112 gnd.n5050 gnd.n1319 19.3944
R17113 gnd.n5050 gnd.n5049 19.3944
R17114 gnd.n5049 gnd.n5048 19.3944
R17115 gnd.n5048 gnd.n1339 19.3944
R17116 gnd.n5038 gnd.n1339 19.3944
R17117 gnd.n5038 gnd.n5037 19.3944
R17118 gnd.n1364 gnd.n1358 19.3944
R17119 gnd.n2683 gnd.n1364 19.3944
R17120 gnd.n2659 gnd.n2658 19.3944
R17121 gnd.n2976 gnd.n2975 19.3944
R17122 gnd.n5034 gnd.n1365 19.3944
R17123 gnd.n5034 gnd.n1366 19.3944
R17124 gnd.n5024 gnd.n1366 19.3944
R17125 gnd.n5024 gnd.n5023 19.3944
R17126 gnd.n5023 gnd.n5022 19.3944
R17127 gnd.n5022 gnd.n1387 19.3944
R17128 gnd.n5012 gnd.n1387 19.3944
R17129 gnd.n5012 gnd.n5011 19.3944
R17130 gnd.n5011 gnd.n5010 19.3944
R17131 gnd.n5010 gnd.n1408 19.3944
R17132 gnd.n5000 gnd.n1408 19.3944
R17133 gnd.n5000 gnd.n4999 19.3944
R17134 gnd.n4999 gnd.n4998 19.3944
R17135 gnd.n4998 gnd.n1427 19.3944
R17136 gnd.n4988 gnd.n1427 19.3944
R17137 gnd.n4988 gnd.n4987 19.3944
R17138 gnd.n4987 gnd.n4986 19.3944
R17139 gnd.n4986 gnd.n1448 19.3944
R17140 gnd.n4976 gnd.n1448 19.3944
R17141 gnd.n4976 gnd.n4975 19.3944
R17142 gnd.n4975 gnd.n4974 19.3944
R17143 gnd.n4974 gnd.n1468 19.3944
R17144 gnd.n4964 gnd.n1468 19.3944
R17145 gnd.n6794 gnd.n6793 19.3944
R17146 gnd.n6793 gnd.n6792 19.3944
R17147 gnd.n6792 gnd.n877 19.3944
R17148 gnd.n6786 gnd.n877 19.3944
R17149 gnd.n6786 gnd.n6785 19.3944
R17150 gnd.n6785 gnd.n6784 19.3944
R17151 gnd.n6784 gnd.n885 19.3944
R17152 gnd.n6778 gnd.n885 19.3944
R17153 gnd.n6778 gnd.n6777 19.3944
R17154 gnd.n6777 gnd.n6776 19.3944
R17155 gnd.n6776 gnd.n893 19.3944
R17156 gnd.n6770 gnd.n893 19.3944
R17157 gnd.n6770 gnd.n6769 19.3944
R17158 gnd.n6769 gnd.n6768 19.3944
R17159 gnd.n6768 gnd.n901 19.3944
R17160 gnd.n6762 gnd.n901 19.3944
R17161 gnd.n6762 gnd.n6761 19.3944
R17162 gnd.n6761 gnd.n6760 19.3944
R17163 gnd.n6760 gnd.n909 19.3944
R17164 gnd.n6754 gnd.n909 19.3944
R17165 gnd.n6754 gnd.n6753 19.3944
R17166 gnd.n6753 gnd.n6752 19.3944
R17167 gnd.n6752 gnd.n917 19.3944
R17168 gnd.n6746 gnd.n917 19.3944
R17169 gnd.n6746 gnd.n6745 19.3944
R17170 gnd.n6745 gnd.n6744 19.3944
R17171 gnd.n6744 gnd.n925 19.3944
R17172 gnd.n6738 gnd.n925 19.3944
R17173 gnd.n6738 gnd.n6737 19.3944
R17174 gnd.n6737 gnd.n6736 19.3944
R17175 gnd.n6736 gnd.n933 19.3944
R17176 gnd.n6730 gnd.n933 19.3944
R17177 gnd.n6730 gnd.n6729 19.3944
R17178 gnd.n6729 gnd.n6728 19.3944
R17179 gnd.n6728 gnd.n941 19.3944
R17180 gnd.n6722 gnd.n941 19.3944
R17181 gnd.n6722 gnd.n6721 19.3944
R17182 gnd.n6721 gnd.n6720 19.3944
R17183 gnd.n6720 gnd.n949 19.3944
R17184 gnd.n6714 gnd.n949 19.3944
R17185 gnd.n6714 gnd.n6713 19.3944
R17186 gnd.n6713 gnd.n6712 19.3944
R17187 gnd.n6712 gnd.n957 19.3944
R17188 gnd.n6706 gnd.n957 19.3944
R17189 gnd.n6706 gnd.n6705 19.3944
R17190 gnd.n6705 gnd.n6704 19.3944
R17191 gnd.n6704 gnd.n965 19.3944
R17192 gnd.n6698 gnd.n965 19.3944
R17193 gnd.n6698 gnd.n6697 19.3944
R17194 gnd.n6697 gnd.n6696 19.3944
R17195 gnd.n6696 gnd.n973 19.3944
R17196 gnd.n6690 gnd.n973 19.3944
R17197 gnd.n6690 gnd.n6689 19.3944
R17198 gnd.n6689 gnd.n6688 19.3944
R17199 gnd.n6688 gnd.n981 19.3944
R17200 gnd.n6682 gnd.n981 19.3944
R17201 gnd.n6682 gnd.n6681 19.3944
R17202 gnd.n6681 gnd.n6680 19.3944
R17203 gnd.n6680 gnd.n989 19.3944
R17204 gnd.n6674 gnd.n989 19.3944
R17205 gnd.n6674 gnd.n6673 19.3944
R17206 gnd.n6673 gnd.n6672 19.3944
R17207 gnd.n6672 gnd.n997 19.3944
R17208 gnd.n6666 gnd.n997 19.3944
R17209 gnd.n6666 gnd.n6665 19.3944
R17210 gnd.n6665 gnd.n6664 19.3944
R17211 gnd.n6664 gnd.n1005 19.3944
R17212 gnd.n6658 gnd.n1005 19.3944
R17213 gnd.n6658 gnd.n6657 19.3944
R17214 gnd.n6657 gnd.n6656 19.3944
R17215 gnd.n6656 gnd.n1013 19.3944
R17216 gnd.n6650 gnd.n1013 19.3944
R17217 gnd.n6650 gnd.n6649 19.3944
R17218 gnd.n6649 gnd.n6648 19.3944
R17219 gnd.n6648 gnd.n1021 19.3944
R17220 gnd.n6642 gnd.n1021 19.3944
R17221 gnd.n6642 gnd.n6641 19.3944
R17222 gnd.n6641 gnd.n6640 19.3944
R17223 gnd.n6640 gnd.n1029 19.3944
R17224 gnd.n6634 gnd.n1029 19.3944
R17225 gnd.n6634 gnd.n6633 19.3944
R17226 gnd.n6633 gnd.n6632 19.3944
R17227 gnd.n6632 gnd.n1037 19.3944
R17228 gnd.n5233 gnd.n1037 19.3944
R17229 gnd.n3236 gnd.n2384 19.3944
R17230 gnd.n3241 gnd.n2384 19.3944
R17231 gnd.n3241 gnd.n2385 19.3944
R17232 gnd.n2385 gnd.n2363 19.3944
R17233 gnd.n3266 gnd.n2363 19.3944
R17234 gnd.n3266 gnd.n2360 19.3944
R17235 gnd.n3271 gnd.n2360 19.3944
R17236 gnd.n3271 gnd.n2361 19.3944
R17237 gnd.n2361 gnd.n2338 19.3944
R17238 gnd.n3302 gnd.n2338 19.3944
R17239 gnd.n3302 gnd.n2335 19.3944
R17240 gnd.n3316 gnd.n2335 19.3944
R17241 gnd.n3316 gnd.n2336 19.3944
R17242 gnd.n3312 gnd.n2336 19.3944
R17243 gnd.n3312 gnd.n3311 19.3944
R17244 gnd.n3311 gnd.n3310 19.3944
R17245 gnd.n3310 gnd.n1621 19.3944
R17246 gnd.n4824 gnd.n1621 19.3944
R17247 gnd.n4824 gnd.n1622 19.3944
R17248 gnd.n4820 gnd.n1622 19.3944
R17249 gnd.n4820 gnd.n4819 19.3944
R17250 gnd.n4819 gnd.n4818 19.3944
R17251 gnd.n4818 gnd.n1628 19.3944
R17252 gnd.n4814 gnd.n1628 19.3944
R17253 gnd.n4814 gnd.n4813 19.3944
R17254 gnd.n4813 gnd.n4812 19.3944
R17255 gnd.n4812 gnd.n1633 19.3944
R17256 gnd.n4808 gnd.n1633 19.3944
R17257 gnd.n4808 gnd.n4807 19.3944
R17258 gnd.n4807 gnd.n4806 19.3944
R17259 gnd.n4806 gnd.n1638 19.3944
R17260 gnd.n4802 gnd.n1638 19.3944
R17261 gnd.n4802 gnd.n4801 19.3944
R17262 gnd.n4801 gnd.n4800 19.3944
R17263 gnd.n4800 gnd.n1643 19.3944
R17264 gnd.n4796 gnd.n1643 19.3944
R17265 gnd.n4796 gnd.n4795 19.3944
R17266 gnd.n4795 gnd.n4794 19.3944
R17267 gnd.n4794 gnd.n1648 19.3944
R17268 gnd.n4790 gnd.n1648 19.3944
R17269 gnd.n4790 gnd.n4789 19.3944
R17270 gnd.n4789 gnd.n4788 19.3944
R17271 gnd.n4788 gnd.n1653 19.3944
R17272 gnd.n4784 gnd.n1653 19.3944
R17273 gnd.n4784 gnd.n4783 19.3944
R17274 gnd.n4783 gnd.n4782 19.3944
R17275 gnd.n4782 gnd.n1658 19.3944
R17276 gnd.n4778 gnd.n1658 19.3944
R17277 gnd.n4778 gnd.n4777 19.3944
R17278 gnd.n4777 gnd.n4776 19.3944
R17279 gnd.n4776 gnd.n1663 19.3944
R17280 gnd.n4772 gnd.n1663 19.3944
R17281 gnd.n4772 gnd.n4771 19.3944
R17282 gnd.n4771 gnd.n4770 19.3944
R17283 gnd.n4770 gnd.n1668 19.3944
R17284 gnd.n4766 gnd.n1668 19.3944
R17285 gnd.n4766 gnd.n4765 19.3944
R17286 gnd.n4765 gnd.n4764 19.3944
R17287 gnd.n4764 gnd.n1673 19.3944
R17288 gnd.n4760 gnd.n1673 19.3944
R17289 gnd.n4760 gnd.n4759 19.3944
R17290 gnd.n4759 gnd.n4758 19.3944
R17291 gnd.n4758 gnd.n1678 19.3944
R17292 gnd.n4754 gnd.n1678 19.3944
R17293 gnd.n4754 gnd.n4753 19.3944
R17294 gnd.n4753 gnd.n4752 19.3944
R17295 gnd.n4752 gnd.n1683 19.3944
R17296 gnd.n4748 gnd.n1683 19.3944
R17297 gnd.n4748 gnd.n4747 19.3944
R17298 gnd.n4747 gnd.n4746 19.3944
R17299 gnd.n4746 gnd.n1688 19.3944
R17300 gnd.n4742 gnd.n1688 19.3944
R17301 gnd.n4742 gnd.n4741 19.3944
R17302 gnd.n4741 gnd.n4740 19.3944
R17303 gnd.n4740 gnd.n1693 19.3944
R17304 gnd.n4736 gnd.n1693 19.3944
R17305 gnd.n4736 gnd.n4735 19.3944
R17306 gnd.n4735 gnd.n4734 19.3944
R17307 gnd.n4734 gnd.n1698 19.3944
R17308 gnd.n4730 gnd.n1698 19.3944
R17309 gnd.n4730 gnd.n4729 19.3944
R17310 gnd.n4729 gnd.n4728 19.3944
R17311 gnd.n3990 gnd.n3987 19.3944
R17312 gnd.n3990 gnd.n3985 19.3944
R17313 gnd.n3996 gnd.n3985 19.3944
R17314 gnd.n3996 gnd.n3983 19.3944
R17315 gnd.n4001 gnd.n3983 19.3944
R17316 gnd.n4001 gnd.n3981 19.3944
R17317 gnd.n4007 gnd.n3981 19.3944
R17318 gnd.n4007 gnd.n3980 19.3944
R17319 gnd.n4016 gnd.n3980 19.3944
R17320 gnd.n4016 gnd.n3978 19.3944
R17321 gnd.n4022 gnd.n3978 19.3944
R17322 gnd.n4022 gnd.n3971 19.3944
R17323 gnd.n4035 gnd.n3971 19.3944
R17324 gnd.n4035 gnd.n3969 19.3944
R17325 gnd.n4041 gnd.n3969 19.3944
R17326 gnd.n4041 gnd.n3962 19.3944
R17327 gnd.n4054 gnd.n3962 19.3944
R17328 gnd.n4054 gnd.n3960 19.3944
R17329 gnd.n4060 gnd.n3960 19.3944
R17330 gnd.n4060 gnd.n3953 19.3944
R17331 gnd.n4073 gnd.n3953 19.3944
R17332 gnd.n4073 gnd.n3951 19.3944
R17333 gnd.n4080 gnd.n3951 19.3944
R17334 gnd.n4080 gnd.n4079 19.3944
R17335 gnd.n4093 gnd.n3932 19.3944
R17336 gnd.n3932 gnd.n3931 19.3944
R17337 gnd.n4100 gnd.n3931 19.3944
R17338 gnd.n6028 gnd.t1 18.8012
R17339 gnd.n6013 gnd.t359 18.8012
R17340 gnd.n5872 gnd.n5871 18.4825
R17341 gnd.n4405 gnd.n4313 18.4247
R17342 gnd.n4916 gnd.n4915 18.4247
R17343 gnd.n4090 gnd.n4089 18.2308
R17344 gnd.n3163 gnd.n3162 18.2308
R17345 gnd.n7664 gnd.n7663 18.2308
R17346 gnd.n2771 gnd.n2770 18.2308
R17347 gnd.t302 gnd.n5552 18.1639
R17348 gnd.n6628 gnd.n6627 18.1639
R17349 gnd.n4845 gnd.n4844 17.6395
R17350 gnd.n4240 gnd.n4239 17.6395
R17351 gnd.n5580 gnd.t2 17.5266
R17352 gnd.t24 gnd.n1249 17.5266
R17353 gnd.n4984 gnd.t158 17.5266
R17354 gnd.n4692 gnd.t167 17.5266
R17355 gnd.n358 gnd.t28 17.5266
R17356 gnd.n5979 gnd.t130 16.8893
R17357 gnd.n5008 gnd.t152 16.8893
R17358 gnd.n4668 gnd.t178 16.8893
R17359 gnd.n4435 gnd.n1958 16.6793
R17360 gnd.n7736 gnd.n7735 16.6793
R17361 gnd.n5153 gnd.n5150 16.6793
R17362 gnd.n2475 gnd.n2445 16.6793
R17363 gnd.n5807 gnd.t13 16.2519
R17364 gnd.n5507 gnd.t132 16.2519
R17365 gnd.n5032 gnd.t231 16.2519
R17366 gnd.n4644 gnd.t209 16.2519
R17367 gnd.n3329 gnd.n3328 16.0975
R17368 gnd.n2005 gnd.n2004 16.0975
R17369 gnd.n4847 gnd.n4846 16.0975
R17370 gnd.n4176 gnd.n4175 16.0975
R17371 gnd.n3222 gnd.n2398 15.9333
R17372 gnd.n3223 gnd.n3222 15.9333
R17373 gnd.n3234 gnd.n2388 15.9333
R17374 gnd.n3234 gnd.n3233 15.9333
R17375 gnd.n3233 gnd.n2390 15.9333
R17376 gnd.n2392 gnd.n2390 15.9333
R17377 gnd.n3243 gnd.n2381 15.9333
R17378 gnd.n2381 gnd.n2374 15.9333
R17379 gnd.n3253 gnd.n2374 15.9333
R17380 gnd.n3253 gnd.n3252 15.9333
R17381 gnd.n3252 gnd.n2365 15.9333
R17382 gnd.n3264 gnd.n2365 15.9333
R17383 gnd.n3264 gnd.n3263 15.9333
R17384 gnd.n3263 gnd.n2367 15.9333
R17385 gnd.n3273 gnd.n2356 15.9333
R17386 gnd.n3273 gnd.n2357 15.9333
R17387 gnd.n2357 gnd.n2349 15.9333
R17388 gnd.n3285 gnd.n2349 15.9333
R17389 gnd.n3285 gnd.n3284 15.9333
R17390 gnd.n3284 gnd.n2340 15.9333
R17391 gnd.n3300 gnd.n2340 15.9333
R17392 gnd.n3300 gnd.n3299 15.9333
R17393 gnd.n2342 gnd.n2332 15.9333
R17394 gnd.n3318 gnd.n2332 15.9333
R17395 gnd.n3318 gnd.n1539 15.9333
R17396 gnd.n3393 gnd.n1571 15.9333
R17397 gnd.n4840 gnd.n1599 15.9333
R17398 gnd.n4834 gnd.n1608 15.9333
R17399 gnd.n4826 gnd.n1618 15.9333
R17400 gnd.n3479 gnd.n3478 15.9333
R17401 gnd.n3512 gnd.n3511 15.9333
R17402 gnd.n2267 gnd.n2256 15.9333
R17403 gnd.n3559 gnd.n2247 15.9333
R17404 gnd.n3532 gnd.n2239 15.9333
R17405 gnd.n3604 gnd.n2230 15.9333
R17406 gnd.n3574 gnd.n2200 15.9333
R17407 gnd.n3655 gnd.n2200 15.9333
R17408 gnd.n3665 gnd.n2178 15.9333
R17409 gnd.n3737 gnd.n3736 15.9333
R17410 gnd.n3745 gnd.n2153 15.9333
R17411 gnd.n3798 gnd.n2142 15.9333
R17412 gnd.n3807 gnd.n3806 15.9333
R17413 gnd.n3837 gnd.n3836 15.9333
R17414 gnd.n3884 gnd.n2085 15.9333
R17415 gnd.n3900 gnd.n2071 15.9333
R17416 gnd.n4151 gnd.n4149 15.9333
R17417 gnd.n2009 gnd.n1971 15.9333
R17418 gnd.n4143 gnd.n4142 15.9333
R17419 gnd.n4142 gnd.n4141 15.9333
R17420 gnd.n4141 gnd.n4140 15.9333
R17421 gnd.n4138 gnd.n2028 15.9333
R17422 gnd.n2036 gnd.n2028 15.9333
R17423 gnd.n2037 gnd.n2036 15.9333
R17424 gnd.n4132 gnd.n2037 15.9333
R17425 gnd.n4132 gnd.n4131 15.9333
R17426 gnd.n4131 gnd.n4130 15.9333
R17427 gnd.n4130 gnd.n4129 15.9333
R17428 gnd.n4129 gnd.n4127 15.9333
R17429 gnd.n2057 gnd.n2056 15.9333
R17430 gnd.n2056 gnd.n2047 15.9333
R17431 gnd.n4121 gnd.n2047 15.9333
R17432 gnd.n4121 gnd.n4120 15.9333
R17433 gnd.n4120 gnd.n4119 15.9333
R17434 gnd.n4119 gnd.n4118 15.9333
R17435 gnd.n4118 gnd.n4116 15.9333
R17436 gnd.n4116 gnd.n2050 15.9333
R17437 gnd.n4107 gnd.n4106 15.9333
R17438 gnd.n4106 gnd.n1704 15.9333
R17439 gnd.n4726 gnd.n1704 15.9333
R17440 gnd.n4726 gnd.n4725 15.9333
R17441 gnd.n1715 gnd.n1706 15.9333
R17442 gnd.n4719 gnd.n1715 15.9333
R17443 gnd.n6424 gnd.n6422 15.6674
R17444 gnd.n6392 gnd.n6390 15.6674
R17445 gnd.n6360 gnd.n6358 15.6674
R17446 gnd.n6329 gnd.n6327 15.6674
R17447 gnd.n6297 gnd.n6295 15.6674
R17448 gnd.n6265 gnd.n6263 15.6674
R17449 gnd.n6233 gnd.n6231 15.6674
R17450 gnd.n6202 gnd.n6200 15.6674
R17451 gnd.n5798 gnd.t13 15.6146
R17452 gnd.t6 gnd.n6585 15.6146
R17453 gnd.n6489 gnd.t104 15.6146
R17454 gnd.n2934 gnd.t184 15.6146
R17455 gnd.n3243 gnd.t69 15.6146
R17456 gnd.t42 gnd.n2050 15.6146
R17457 gnd.n7578 gnd.t227 15.6146
R17458 gnd.n4487 gnd.n1937 15.3217
R17459 gnd.n7696 gnd.n319 15.3217
R17460 gnd.n5110 gnd.n1234 15.3217
R17461 gnd.n2530 gnd.n2423 15.3217
R17462 gnd.n4841 gnd.n1597 15.296
R17463 gnd.n3470 gnd.t319 15.296
R17464 gnd.n3550 gnd.n3548 15.296
R17465 gnd.n3569 gnd.n3568 15.296
R17466 gnd.n3727 gnd.n2159 15.296
R17467 gnd.n3746 gnd.n2149 15.296
R17468 gnd.n3759 gnd.t328 15.296
R17469 gnd.n4160 gnd.n4159 15.0827
R17470 gnd.n1583 gnd.n1578 15.0481
R17471 gnd.n4170 gnd.n4169 15.0481
R17472 gnd.n6620 gnd.t299 14.9773
R17473 gnd.n5058 gnd.t156 14.9773
R17474 gnd.n3299 gnd.t357 14.9773
R17475 gnd.t355 gnd.n4138 14.9773
R17476 gnd.n7606 gnd.t162 14.9773
R17477 gnd.n4833 gnd.t53 14.6587
R17478 gnd.n3460 gnd.n2303 14.6587
R17479 gnd.n3498 gnd.n2283 14.6587
R17480 gnd.n3818 gnd.n3817 14.6587
R17481 gnd.n3760 gnd.n2099 14.6587
R17482 gnd.n2077 gnd.t46 14.6587
R17483 gnd.n6606 gnd.t341 14.34
R17484 gnd.t4 gnd.n1088 14.34
R17485 gnd.n5082 gnd.t201 14.34
R17486 gnd.n7634 gnd.t139 14.34
R17487 gnd.n3885 gnd.n2082 14.0214
R17488 gnd.n5954 gnd.t317 13.7027
R17489 gnd.n5664 gnd.n5663 13.5763
R17490 gnd.n6545 gnd.n5268 13.5763
R17491 gnd.n5872 gnd.n5610 13.384
R17492 gnd.n3452 gnd.n3451 13.384
R17493 gnd.n3521 gnd.n2263 13.384
R17494 gnd.n3585 gnd.n2222 13.384
R17495 gnd.n3613 gnd.t321 13.384
R17496 gnd.n3647 gnd.t335 13.384
R17497 gnd.n3683 gnd.t350 13.384
R17498 gnd.t345 gnd.n2182 13.384
R17499 gnd.n3702 gnd.n3701 13.384
R17500 gnd.n3779 gnd.n2136 13.384
R17501 gnd.n3868 gnd.n2095 13.384
R17502 gnd.n1594 gnd.n1575 13.1884
R17503 gnd.n1589 gnd.n1588 13.1884
R17504 gnd.n1588 gnd.n1587 13.1884
R17505 gnd.n4163 gnd.n4158 13.1884
R17506 gnd.n4164 gnd.n4163 13.1884
R17507 gnd.n1590 gnd.n1577 13.146
R17508 gnd.n1586 gnd.n1577 13.146
R17509 gnd.n4162 gnd.n4161 13.146
R17510 gnd.n4162 gnd.n4157 13.146
R17511 gnd.n6425 gnd.n6421 12.8005
R17512 gnd.n6393 gnd.n6389 12.8005
R17513 gnd.n6361 gnd.n6357 12.8005
R17514 gnd.n6330 gnd.n6326 12.8005
R17515 gnd.n6298 gnd.n6294 12.8005
R17516 gnd.n6266 gnd.n6262 12.8005
R17517 gnd.n6234 gnd.n6230 12.8005
R17518 gnd.n6203 gnd.n6199 12.8005
R17519 gnd.n3513 gnd.n2273 12.7467
R17520 gnd.n2223 gnd.n2212 12.7467
R17521 gnd.n3674 gnd.n2191 12.7467
R17522 gnd.n3775 gnd.n2126 12.7467
R17523 gnd.n2837 gnd.t201 12.4281
R17524 gnd.t139 gnd.n183 12.4281
R17525 gnd.n5663 gnd.n5658 12.4126
R17526 gnd.n6550 gnd.n5268 12.4126
R17527 gnd.n4908 gnd.n4845 12.1761
R17528 gnd.n4239 gnd.n4238 12.1761
R17529 gnd.n4827 gnd.n1615 12.1094
R17530 gnd.n3541 gnd.n3540 12.1094
R17531 gnd.n3593 gnd.n3592 12.1094
R17532 gnd.n3666 gnd.n2168 12.1094
R17533 gnd.n3787 gnd.n3786 12.1094
R17534 gnd.n2084 gnd.t114 12.1094
R17535 gnd.n6429 gnd.n6428 12.0247
R17536 gnd.n6397 gnd.n6396 12.0247
R17537 gnd.n6365 gnd.n6364 12.0247
R17538 gnd.n6334 gnd.n6333 12.0247
R17539 gnd.n6302 gnd.n6301 12.0247
R17540 gnd.n6270 gnd.n6269 12.0247
R17541 gnd.n6238 gnd.n6237 12.0247
R17542 gnd.n6207 gnd.n6206 12.0247
R17543 gnd.n2902 gnd.t156 11.7908
R17544 gnd.t162 gnd.n143 11.7908
R17545 gnd.n3097 gnd.n1487 11.4721
R17546 gnd.t57 gnd.n3419 11.4721
R17547 gnd.n3468 gnd.n2306 11.4721
R17548 gnd.t134 gnd.n2287 11.4721
R17549 gnd.n3491 gnd.n3490 11.4721
R17550 gnd.n3646 gnd.n2207 11.4721
R17551 gnd.n3684 gnd.n2195 11.4721
R17552 gnd.n3825 gnd.n2121 11.4721
R17553 gnd.n3767 gnd.t330 11.4721
R17554 gnd.n3845 gnd.n3843 11.4721
R17555 gnd.n4717 gnd.n1716 11.4721
R17556 gnd.n6432 gnd.n6419 11.249
R17557 gnd.n6400 gnd.n6387 11.249
R17558 gnd.n6368 gnd.n6355 11.249
R17559 gnd.n6337 gnd.n6324 11.249
R17560 gnd.n6305 gnd.n6292 11.249
R17561 gnd.n6273 gnd.n6260 11.249
R17562 gnd.n6241 gnd.n6228 11.249
R17563 gnd.n6210 gnd.n6197 11.249
R17564 gnd.n5942 gnd.t317 11.1535
R17565 gnd.t184 gnd.n2931 11.1535
R17566 gnd.n2367 gnd.t297 11.1535
R17567 gnd.n2057 gnd.t353 11.1535
R17568 gnd.t227 gnd.n102 11.1535
R17569 gnd.n3534 gnd.n3533 10.8348
R17570 gnd.n3735 gnd.n2162 10.8348
R17571 gnd.n4152 gnd.n2014 10.8348
R17572 gnd.n1938 gnd.n1937 10.6672
R17573 gnd.n7701 gnd.n319 10.6672
R17574 gnd.n5113 gnd.n5110 10.6672
R17575 gnd.n2525 gnd.n2423 10.6672
R17576 gnd.n4304 gnd.n1967 10.6151
R17577 gnd.n4304 gnd.n4303 10.6151
R17578 gnd.n4301 gnd.n4298 10.6151
R17579 gnd.n4298 gnd.n4297 10.6151
R17580 gnd.n4297 gnd.n4294 10.6151
R17581 gnd.n4294 gnd.n4293 10.6151
R17582 gnd.n4293 gnd.n4290 10.6151
R17583 gnd.n4290 gnd.n4289 10.6151
R17584 gnd.n4289 gnd.n4286 10.6151
R17585 gnd.n4286 gnd.n4285 10.6151
R17586 gnd.n4285 gnd.n4282 10.6151
R17587 gnd.n4282 gnd.n4281 10.6151
R17588 gnd.n4281 gnd.n4278 10.6151
R17589 gnd.n4278 gnd.n4277 10.6151
R17590 gnd.n4277 gnd.n4274 10.6151
R17591 gnd.n4274 gnd.n4273 10.6151
R17592 gnd.n4273 gnd.n4270 10.6151
R17593 gnd.n4270 gnd.n4269 10.6151
R17594 gnd.n4269 gnd.n4266 10.6151
R17595 gnd.n4266 gnd.n4265 10.6151
R17596 gnd.n4265 gnd.n4262 10.6151
R17597 gnd.n4262 gnd.n4261 10.6151
R17598 gnd.n4261 gnd.n4258 10.6151
R17599 gnd.n4258 gnd.n4257 10.6151
R17600 gnd.n4257 gnd.n4254 10.6151
R17601 gnd.n4254 gnd.n4253 10.6151
R17602 gnd.n4253 gnd.n4250 10.6151
R17603 gnd.n4250 gnd.n4249 10.6151
R17604 gnd.n4249 gnd.n4246 10.6151
R17605 gnd.n4246 gnd.n4245 10.6151
R17606 gnd.n3397 gnd.n3396 10.6151
R17607 gnd.n3398 gnd.n3397 10.6151
R17608 gnd.n3404 gnd.n3398 10.6151
R17609 gnd.n3405 gnd.n3404 10.6151
R17610 gnd.n3407 gnd.n3405 10.6151
R17611 gnd.n3407 gnd.n3406 10.6151
R17612 gnd.n3406 gnd.n2322 10.6151
R17613 gnd.n3423 gnd.n2322 10.6151
R17614 gnd.n3424 gnd.n3423 10.6151
R17615 gnd.n3442 gnd.n3424 10.6151
R17616 gnd.n3442 gnd.n3441 10.6151
R17617 gnd.n3441 gnd.n3440 10.6151
R17618 gnd.n3440 gnd.n3438 10.6151
R17619 gnd.n3438 gnd.n3437 10.6151
R17620 gnd.n3437 gnd.n3435 10.6151
R17621 gnd.n3435 gnd.n3434 10.6151
R17622 gnd.n3434 gnd.n3433 10.6151
R17623 gnd.n3433 gnd.n3432 10.6151
R17624 gnd.n3432 gnd.n3431 10.6151
R17625 gnd.n3431 gnd.n3428 10.6151
R17626 gnd.n3428 gnd.n3427 10.6151
R17627 gnd.n3427 gnd.n3425 10.6151
R17628 gnd.n3425 gnd.n2254 10.6151
R17629 gnd.n3543 gnd.n2254 10.6151
R17630 gnd.n3544 gnd.n3543 10.6151
R17631 gnd.n3546 gnd.n3544 10.6151
R17632 gnd.n3546 gnd.n3545 10.6151
R17633 gnd.n3545 gnd.n2237 10.6151
R17634 gnd.n3571 gnd.n2237 10.6151
R17635 gnd.n3572 gnd.n3571 10.6151
R17636 gnd.n3590 gnd.n3572 10.6151
R17637 gnd.n3590 gnd.n3589 10.6151
R17638 gnd.n3589 gnd.n3588 10.6151
R17639 gnd.n3588 gnd.n3573 10.6151
R17640 gnd.n3581 gnd.n3573 10.6151
R17641 gnd.n3581 gnd.n3580 10.6151
R17642 gnd.n3580 gnd.n3579 10.6151
R17643 gnd.n3579 gnd.n3578 10.6151
R17644 gnd.n3578 gnd.n3577 10.6151
R17645 gnd.n3577 gnd.n2198 10.6151
R17646 gnd.n3658 gnd.n2198 10.6151
R17647 gnd.n3659 gnd.n3658 10.6151
R17648 gnd.n3678 gnd.n3659 10.6151
R17649 gnd.n3678 gnd.n3677 10.6151
R17650 gnd.n3677 gnd.n3676 10.6151
R17651 gnd.n3676 gnd.n3672 10.6151
R17652 gnd.n3672 gnd.n3671 10.6151
R17653 gnd.n3671 gnd.n3669 10.6151
R17654 gnd.n3669 gnd.n3668 10.6151
R17655 gnd.n3668 gnd.n3663 10.6151
R17656 gnd.n3663 gnd.n3662 10.6151
R17657 gnd.n3662 gnd.n3660 10.6151
R17658 gnd.n3660 gnd.n2151 10.6151
R17659 gnd.n3748 gnd.n2151 10.6151
R17660 gnd.n3749 gnd.n3748 10.6151
R17661 gnd.n3784 gnd.n3749 10.6151
R17662 gnd.n3784 gnd.n3783 10.6151
R17663 gnd.n3783 gnd.n3782 10.6151
R17664 gnd.n3782 gnd.n3750 10.6151
R17665 gnd.n3774 gnd.n3750 10.6151
R17666 gnd.n3774 gnd.n3773 10.6151
R17667 gnd.n3773 gnd.n3772 10.6151
R17668 gnd.n3772 gnd.n3771 10.6151
R17669 gnd.n3771 gnd.n3770 10.6151
R17670 gnd.n3770 gnd.n3766 10.6151
R17671 gnd.n3766 gnd.n3765 10.6151
R17672 gnd.n3765 gnd.n3763 10.6151
R17673 gnd.n3763 gnd.n3762 10.6151
R17674 gnd.n3762 gnd.n3758 10.6151
R17675 gnd.n3758 gnd.n3757 10.6151
R17676 gnd.n3757 gnd.n3755 10.6151
R17677 gnd.n3755 gnd.n3754 10.6151
R17678 gnd.n3754 gnd.n3751 10.6151
R17679 gnd.n3751 gnd.n2073 10.6151
R17680 gnd.n3894 gnd.n2073 10.6151
R17681 gnd.n3895 gnd.n3894 10.6151
R17682 gnd.n3898 gnd.n3895 10.6151
R17683 gnd.n3898 gnd.n3897 10.6151
R17684 gnd.n3897 gnd.n3896 10.6151
R17685 gnd.n3896 gnd.n2006 10.6151
R17686 gnd.n3330 gnd.n1535 10.6151
R17687 gnd.n3333 gnd.n3330 10.6151
R17688 gnd.n3338 gnd.n3335 10.6151
R17689 gnd.n3339 gnd.n3338 10.6151
R17690 gnd.n3342 gnd.n3339 10.6151
R17691 gnd.n3343 gnd.n3342 10.6151
R17692 gnd.n3346 gnd.n3343 10.6151
R17693 gnd.n3347 gnd.n3346 10.6151
R17694 gnd.n3350 gnd.n3347 10.6151
R17695 gnd.n3351 gnd.n3350 10.6151
R17696 gnd.n3354 gnd.n3351 10.6151
R17697 gnd.n3355 gnd.n3354 10.6151
R17698 gnd.n3358 gnd.n3355 10.6151
R17699 gnd.n3359 gnd.n3358 10.6151
R17700 gnd.n3362 gnd.n3359 10.6151
R17701 gnd.n3363 gnd.n3362 10.6151
R17702 gnd.n3366 gnd.n3363 10.6151
R17703 gnd.n3367 gnd.n3366 10.6151
R17704 gnd.n3370 gnd.n3367 10.6151
R17705 gnd.n3371 gnd.n3370 10.6151
R17706 gnd.n3374 gnd.n3371 10.6151
R17707 gnd.n3375 gnd.n3374 10.6151
R17708 gnd.n3378 gnd.n3375 10.6151
R17709 gnd.n3379 gnd.n3378 10.6151
R17710 gnd.n3382 gnd.n3379 10.6151
R17711 gnd.n3383 gnd.n3382 10.6151
R17712 gnd.n3386 gnd.n3383 10.6151
R17713 gnd.n3387 gnd.n3386 10.6151
R17714 gnd.n3390 gnd.n3387 10.6151
R17715 gnd.n3391 gnd.n3390 10.6151
R17716 gnd.n4908 gnd.n4907 10.6151
R17717 gnd.n4907 gnd.n4906 10.6151
R17718 gnd.n4906 gnd.n4905 10.6151
R17719 gnd.n4905 gnd.n4903 10.6151
R17720 gnd.n4903 gnd.n4900 10.6151
R17721 gnd.n4900 gnd.n4899 10.6151
R17722 gnd.n4899 gnd.n4896 10.6151
R17723 gnd.n4896 gnd.n4895 10.6151
R17724 gnd.n4895 gnd.n4892 10.6151
R17725 gnd.n4892 gnd.n4891 10.6151
R17726 gnd.n4891 gnd.n4888 10.6151
R17727 gnd.n4888 gnd.n4887 10.6151
R17728 gnd.n4887 gnd.n4884 10.6151
R17729 gnd.n4884 gnd.n4883 10.6151
R17730 gnd.n4883 gnd.n4880 10.6151
R17731 gnd.n4880 gnd.n4879 10.6151
R17732 gnd.n4879 gnd.n4876 10.6151
R17733 gnd.n4876 gnd.n4875 10.6151
R17734 gnd.n4875 gnd.n4872 10.6151
R17735 gnd.n4872 gnd.n4871 10.6151
R17736 gnd.n4871 gnd.n4868 10.6151
R17737 gnd.n4868 gnd.n4867 10.6151
R17738 gnd.n4867 gnd.n4864 10.6151
R17739 gnd.n4864 gnd.n4863 10.6151
R17740 gnd.n4863 gnd.n4860 10.6151
R17741 gnd.n4860 gnd.n4859 10.6151
R17742 gnd.n4859 gnd.n4856 10.6151
R17743 gnd.n4856 gnd.n4855 10.6151
R17744 gnd.n4852 gnd.n4851 10.6151
R17745 gnd.n4851 gnd.n1536 10.6151
R17746 gnd.n4238 gnd.n4237 10.6151
R17747 gnd.n4237 gnd.n4234 10.6151
R17748 gnd.n4234 gnd.n4233 10.6151
R17749 gnd.n4233 gnd.n4230 10.6151
R17750 gnd.n4230 gnd.n4229 10.6151
R17751 gnd.n4229 gnd.n4226 10.6151
R17752 gnd.n4226 gnd.n4225 10.6151
R17753 gnd.n4225 gnd.n4222 10.6151
R17754 gnd.n4222 gnd.n4221 10.6151
R17755 gnd.n4221 gnd.n4218 10.6151
R17756 gnd.n4218 gnd.n4217 10.6151
R17757 gnd.n4217 gnd.n4214 10.6151
R17758 gnd.n4214 gnd.n4213 10.6151
R17759 gnd.n4213 gnd.n4210 10.6151
R17760 gnd.n4210 gnd.n4209 10.6151
R17761 gnd.n4209 gnd.n4206 10.6151
R17762 gnd.n4206 gnd.n4205 10.6151
R17763 gnd.n4205 gnd.n4202 10.6151
R17764 gnd.n4202 gnd.n4201 10.6151
R17765 gnd.n4201 gnd.n4198 10.6151
R17766 gnd.n4198 gnd.n4197 10.6151
R17767 gnd.n4197 gnd.n4194 10.6151
R17768 gnd.n4194 gnd.n4193 10.6151
R17769 gnd.n4193 gnd.n4190 10.6151
R17770 gnd.n4190 gnd.n4189 10.6151
R17771 gnd.n4189 gnd.n4186 10.6151
R17772 gnd.n4186 gnd.n4185 10.6151
R17773 gnd.n4185 gnd.n4182 10.6151
R17774 gnd.n4180 gnd.n4177 10.6151
R17775 gnd.n4177 gnd.n1968 10.6151
R17776 gnd.n4844 gnd.n4843 10.6151
R17777 gnd.n4843 gnd.n1595 10.6151
R17778 gnd.n1612 gnd.n1595 10.6151
R17779 gnd.n4831 gnd.n1612 10.6151
R17780 gnd.n4831 gnd.n4830 10.6151
R17781 gnd.n4830 gnd.n4829 10.6151
R17782 gnd.n4829 gnd.n1613 10.6151
R17783 gnd.n3448 gnd.n1613 10.6151
R17784 gnd.n3449 gnd.n3448 10.6151
R17785 gnd.n3449 gnd.n2309 10.6151
R17786 gnd.n3463 gnd.n2309 10.6151
R17787 gnd.n3464 gnd.n3463 10.6151
R17788 gnd.n3466 gnd.n3464 10.6151
R17789 gnd.n3466 gnd.n3465 10.6151
R17790 gnd.n3465 gnd.n2285 10.6151
R17791 gnd.n3494 gnd.n2285 10.6151
R17792 gnd.n3495 gnd.n3494 10.6151
R17793 gnd.n3496 gnd.n3495 10.6151
R17794 gnd.n3496 gnd.n2270 10.6151
R17795 gnd.n3515 gnd.n2270 10.6151
R17796 gnd.n3516 gnd.n3515 10.6151
R17797 gnd.n3518 gnd.n3516 10.6151
R17798 gnd.n3518 gnd.n3517 10.6151
R17799 gnd.n3517 gnd.n2251 10.6151
R17800 gnd.n3553 gnd.n2251 10.6151
R17801 gnd.n3554 gnd.n3553 10.6151
R17802 gnd.n3556 gnd.n3554 10.6151
R17803 gnd.n3556 gnd.n3555 10.6151
R17804 gnd.n3555 gnd.n2234 10.6151
R17805 gnd.n3596 gnd.n2234 10.6151
R17806 gnd.n3597 gnd.n3596 10.6151
R17807 gnd.n3601 gnd.n3597 10.6151
R17808 gnd.n3601 gnd.n3600 10.6151
R17809 gnd.n3600 gnd.n3599 10.6151
R17810 gnd.n3599 gnd.n2210 10.6151
R17811 gnd.n3639 gnd.n2210 10.6151
R17812 gnd.n3640 gnd.n3639 10.6151
R17813 gnd.n3644 gnd.n3640 10.6151
R17814 gnd.n3644 gnd.n3643 10.6151
R17815 gnd.n3643 gnd.n3642 10.6151
R17816 gnd.n3642 gnd.n2193 10.6151
R17817 gnd.n3686 gnd.n2193 10.6151
R17818 gnd.n3687 gnd.n3686 10.6151
R17819 gnd.n3688 gnd.n3687 10.6151
R17820 gnd.n3688 gnd.n2180 10.6151
R17821 gnd.n3704 gnd.n2180 10.6151
R17822 gnd.n3705 gnd.n3704 10.6151
R17823 gnd.n3706 gnd.n3705 10.6151
R17824 gnd.n3706 gnd.n2166 10.6151
R17825 gnd.n3730 gnd.n2166 10.6151
R17826 gnd.n3731 gnd.n3730 10.6151
R17827 gnd.n3733 gnd.n3731 10.6151
R17828 gnd.n3733 gnd.n3732 10.6151
R17829 gnd.n3732 gnd.n2146 10.6151
R17830 gnd.n3790 gnd.n2146 10.6151
R17831 gnd.n3791 gnd.n3790 10.6151
R17832 gnd.n3795 gnd.n3791 10.6151
R17833 gnd.n3795 gnd.n3794 10.6151
R17834 gnd.n3794 gnd.n3793 10.6151
R17835 gnd.n3793 gnd.n2123 10.6151
R17836 gnd.n3821 gnd.n2123 10.6151
R17837 gnd.n3822 gnd.n3821 10.6151
R17838 gnd.n3823 gnd.n3822 10.6151
R17839 gnd.n3823 gnd.n2111 10.6151
R17840 gnd.n3839 gnd.n2111 10.6151
R17841 gnd.n3840 gnd.n3839 10.6151
R17842 gnd.n3841 gnd.n3840 10.6151
R17843 gnd.n3841 gnd.n2097 10.6151
R17844 gnd.n3864 gnd.n2097 10.6151
R17845 gnd.n3865 gnd.n3864 10.6151
R17846 gnd.n3866 gnd.n3865 10.6151
R17847 gnd.n3866 gnd.n2079 10.6151
R17848 gnd.n3887 gnd.n2079 10.6151
R17849 gnd.n3888 gnd.n3887 10.6151
R17850 gnd.n3890 gnd.n3888 10.6151
R17851 gnd.n3890 gnd.n3889 10.6151
R17852 gnd.n3889 gnd.n2012 10.6151
R17853 gnd.n4154 gnd.n2012 10.6151
R17854 gnd.n4155 gnd.n4154 10.6151
R17855 gnd.n4240 gnd.n4155 10.6151
R17856 gnd.n5861 gnd.t337 10.5161
R17857 gnd.n6471 gnd.t341 10.5161
R17858 gnd.n6478 gnd.t4 10.5161
R17859 gnd.n3006 gnd.t231 10.5161
R17860 gnd.n4911 gnd.n1571 10.5161
R17861 gnd.n4309 gnd.n1971 10.5161
R17862 gnd.n4621 gnd.t209 10.5161
R17863 gnd.n6433 gnd.n6417 10.4732
R17864 gnd.n6401 gnd.n6385 10.4732
R17865 gnd.n6369 gnd.n6353 10.4732
R17866 gnd.n6338 gnd.n6322 10.4732
R17867 gnd.n6306 gnd.n6290 10.4732
R17868 gnd.n6274 gnd.n6258 10.4732
R17869 gnd.n6242 gnd.n6226 10.4732
R17870 gnd.n6211 gnd.n6195 10.4732
R17871 gnd.n2306 gnd.n2296 10.1975
R17872 gnd.n2268 gnd.t133 10.1975
R17873 gnd.n3575 gnd.n2207 10.1975
R17874 gnd.n3656 gnd.n2195 10.1975
R17875 gnd.n3797 gnd.t310 10.1975
R17876 gnd.n3845 gnd.n2107 10.1975
R17877 gnd.n6146 gnd.t299 9.87883
R17878 gnd.n3067 gnd.t152 9.87883
R17879 gnd.n4530 gnd.t178 9.87883
R17880 gnd.n6437 gnd.n6436 9.69747
R17881 gnd.n6405 gnd.n6404 9.69747
R17882 gnd.n6373 gnd.n6372 9.69747
R17883 gnd.n6342 gnd.n6341 9.69747
R17884 gnd.n6310 gnd.n6309 9.69747
R17885 gnd.n6278 gnd.n6277 9.69747
R17886 gnd.n6246 gnd.n6245 9.69747
R17887 gnd.n6215 gnd.n6214 9.69747
R17888 gnd.n3409 gnd.n1615 9.56018
R17889 gnd.n3489 gnd.t327 9.56018
R17890 gnd.n3594 gnd.n3593 9.56018
R17891 gnd.n3728 gnd.n2168 9.56018
R17892 gnd.n3826 gnd.t329 9.56018
R17893 gnd.n3892 gnd.t114 9.56018
R17894 gnd.n2017 gnd.t10 9.56018
R17895 gnd.n4242 gnd.n2009 9.56018
R17896 gnd.n6443 gnd.n6442 9.45567
R17897 gnd.n6411 gnd.n6410 9.45567
R17898 gnd.n6379 gnd.n6378 9.45567
R17899 gnd.n6348 gnd.n6347 9.45567
R17900 gnd.n6316 gnd.n6315 9.45567
R17901 gnd.n6284 gnd.n6283 9.45567
R17902 gnd.n6252 gnd.n6251 9.45567
R17903 gnd.n6221 gnd.n6220 9.45567
R17904 gnd.n4435 gnd.n1956 9.30959
R17905 gnd.n7735 gnd.n283 9.30959
R17906 gnd.n5150 gnd.n5149 9.30959
R17907 gnd.n2481 gnd.n2445 9.30959
R17908 gnd.n6442 gnd.n6441 9.3005
R17909 gnd.n6415 gnd.n6414 9.3005
R17910 gnd.n6436 gnd.n6435 9.3005
R17911 gnd.n6434 gnd.n6433 9.3005
R17912 gnd.n6419 gnd.n6418 9.3005
R17913 gnd.n6428 gnd.n6427 9.3005
R17914 gnd.n6426 gnd.n6425 9.3005
R17915 gnd.n6410 gnd.n6409 9.3005
R17916 gnd.n6383 gnd.n6382 9.3005
R17917 gnd.n6404 gnd.n6403 9.3005
R17918 gnd.n6402 gnd.n6401 9.3005
R17919 gnd.n6387 gnd.n6386 9.3005
R17920 gnd.n6396 gnd.n6395 9.3005
R17921 gnd.n6394 gnd.n6393 9.3005
R17922 gnd.n6378 gnd.n6377 9.3005
R17923 gnd.n6351 gnd.n6350 9.3005
R17924 gnd.n6372 gnd.n6371 9.3005
R17925 gnd.n6370 gnd.n6369 9.3005
R17926 gnd.n6355 gnd.n6354 9.3005
R17927 gnd.n6364 gnd.n6363 9.3005
R17928 gnd.n6362 gnd.n6361 9.3005
R17929 gnd.n6347 gnd.n6346 9.3005
R17930 gnd.n6320 gnd.n6319 9.3005
R17931 gnd.n6341 gnd.n6340 9.3005
R17932 gnd.n6339 gnd.n6338 9.3005
R17933 gnd.n6324 gnd.n6323 9.3005
R17934 gnd.n6333 gnd.n6332 9.3005
R17935 gnd.n6331 gnd.n6330 9.3005
R17936 gnd.n6315 gnd.n6314 9.3005
R17937 gnd.n6288 gnd.n6287 9.3005
R17938 gnd.n6309 gnd.n6308 9.3005
R17939 gnd.n6307 gnd.n6306 9.3005
R17940 gnd.n6292 gnd.n6291 9.3005
R17941 gnd.n6301 gnd.n6300 9.3005
R17942 gnd.n6299 gnd.n6298 9.3005
R17943 gnd.n6283 gnd.n6282 9.3005
R17944 gnd.n6256 gnd.n6255 9.3005
R17945 gnd.n6277 gnd.n6276 9.3005
R17946 gnd.n6275 gnd.n6274 9.3005
R17947 gnd.n6260 gnd.n6259 9.3005
R17948 gnd.n6269 gnd.n6268 9.3005
R17949 gnd.n6267 gnd.n6266 9.3005
R17950 gnd.n6251 gnd.n6250 9.3005
R17951 gnd.n6224 gnd.n6223 9.3005
R17952 gnd.n6245 gnd.n6244 9.3005
R17953 gnd.n6243 gnd.n6242 9.3005
R17954 gnd.n6228 gnd.n6227 9.3005
R17955 gnd.n6237 gnd.n6236 9.3005
R17956 gnd.n6235 gnd.n6234 9.3005
R17957 gnd.n6220 gnd.n6219 9.3005
R17958 gnd.n6193 gnd.n6192 9.3005
R17959 gnd.n6214 gnd.n6213 9.3005
R17960 gnd.n6212 gnd.n6211 9.3005
R17961 gnd.n6197 gnd.n6196 9.3005
R17962 gnd.n6206 gnd.n6205 9.3005
R17963 gnd.n6204 gnd.n6203 9.3005
R17964 gnd.n6572 gnd.n5242 9.3005
R17965 gnd.n6571 gnd.n5244 9.3005
R17966 gnd.n5248 gnd.n5245 9.3005
R17967 gnd.n6566 gnd.n5249 9.3005
R17968 gnd.n6565 gnd.n5250 9.3005
R17969 gnd.n6564 gnd.n5251 9.3005
R17970 gnd.n5255 gnd.n5252 9.3005
R17971 gnd.n6559 gnd.n5256 9.3005
R17972 gnd.n6558 gnd.n5257 9.3005
R17973 gnd.n6557 gnd.n5258 9.3005
R17974 gnd.n5262 gnd.n5259 9.3005
R17975 gnd.n6552 gnd.n5263 9.3005
R17976 gnd.n6551 gnd.n5264 9.3005
R17977 gnd.n6550 gnd.n5265 9.3005
R17978 gnd.n5270 gnd.n5268 9.3005
R17979 gnd.n6545 gnd.n6544 9.3005
R17980 gnd.n6574 gnd.n6573 9.3005
R17981 gnd.n5880 gnd.n5879 9.3005
R17982 gnd.n5584 gnd.n5583 9.3005
R17983 gnd.n5907 gnd.n5906 9.3005
R17984 gnd.n5908 gnd.n5582 9.3005
R17985 gnd.n5912 gnd.n5909 9.3005
R17986 gnd.n5911 gnd.n5910 9.3005
R17987 gnd.n5556 gnd.n5555 9.3005
R17988 gnd.n5937 gnd.n5936 9.3005
R17989 gnd.n5938 gnd.n5554 9.3005
R17990 gnd.n5940 gnd.n5939 9.3005
R17991 gnd.n5534 gnd.n5533 9.3005
R17992 gnd.n5968 gnd.n5967 9.3005
R17993 gnd.n5969 gnd.n5532 9.3005
R17994 gnd.n5977 gnd.n5970 9.3005
R17995 gnd.n5976 gnd.n5971 9.3005
R17996 gnd.n5975 gnd.n5973 9.3005
R17997 gnd.n5972 gnd.n5481 9.3005
R17998 gnd.n6025 gnd.n5482 9.3005
R17999 gnd.n6024 gnd.n5483 9.3005
R18000 gnd.n6023 gnd.n5484 9.3005
R18001 gnd.n5503 gnd.n5485 9.3005
R18002 gnd.n5505 gnd.n5504 9.3005
R18003 gnd.n5387 gnd.n5386 9.3005
R18004 gnd.n6063 gnd.n6062 9.3005
R18005 gnd.n6064 gnd.n5385 9.3005
R18006 gnd.n6068 gnd.n6065 9.3005
R18007 gnd.n6067 gnd.n6066 9.3005
R18008 gnd.n5360 gnd.n5359 9.3005
R18009 gnd.n6103 gnd.n6102 9.3005
R18010 gnd.n6104 gnd.n5358 9.3005
R18011 gnd.n6108 gnd.n6105 9.3005
R18012 gnd.n6107 gnd.n6106 9.3005
R18013 gnd.n5334 gnd.n5333 9.3005
R18014 gnd.n6159 gnd.n6158 9.3005
R18015 gnd.n6160 gnd.n5332 9.3005
R18016 gnd.n6163 gnd.n6162 9.3005
R18017 gnd.n6161 gnd.n1054 9.3005
R18018 gnd.n6618 gnd.n1055 9.3005
R18019 gnd.n6617 gnd.n1056 9.3005
R18020 gnd.n6616 gnd.n1057 9.3005
R18021 gnd.n1078 gnd.n1058 9.3005
R18022 gnd.n1079 gnd.n1077 9.3005
R18023 gnd.n6604 gnd.n1080 9.3005
R18024 gnd.n6603 gnd.n1081 9.3005
R18025 gnd.n6602 gnd.n1082 9.3005
R18026 gnd.n1104 gnd.n1083 9.3005
R18027 gnd.n1105 gnd.n1103 9.3005
R18028 gnd.n6590 gnd.n1106 9.3005
R18029 gnd.n6589 gnd.n1107 9.3005
R18030 gnd.n6588 gnd.n1108 9.3005
R18031 gnd.n5240 gnd.n1109 9.3005
R18032 gnd.n5241 gnd.n5239 9.3005
R18033 gnd.n6576 gnd.n6575 9.3005
R18034 gnd.n5881 gnd.n5878 9.3005
R18035 gnd.n5663 gnd.n5622 9.3005
R18036 gnd.n5658 gnd.n5657 9.3005
R18037 gnd.n5656 gnd.n5623 9.3005
R18038 gnd.n5655 gnd.n5654 9.3005
R18039 gnd.n5651 gnd.n5624 9.3005
R18040 gnd.n5648 gnd.n5647 9.3005
R18041 gnd.n5646 gnd.n5625 9.3005
R18042 gnd.n5645 gnd.n5644 9.3005
R18043 gnd.n5641 gnd.n5626 9.3005
R18044 gnd.n5638 gnd.n5637 9.3005
R18045 gnd.n5636 gnd.n5627 9.3005
R18046 gnd.n5635 gnd.n5634 9.3005
R18047 gnd.n5631 gnd.n5629 9.3005
R18048 gnd.n5628 gnd.n5608 9.3005
R18049 gnd.n5875 gnd.n5607 9.3005
R18050 gnd.n5877 gnd.n5876 9.3005
R18051 gnd.n5665 gnd.n5664 9.3005
R18052 gnd.n5888 gnd.n5594 9.3005
R18053 gnd.n5895 gnd.n5595 9.3005
R18054 gnd.n5897 gnd.n5896 9.3005
R18055 gnd.n5898 gnd.n5575 9.3005
R18056 gnd.n5917 gnd.n5916 9.3005
R18057 gnd.n5919 gnd.n5567 9.3005
R18058 gnd.n5926 gnd.n5569 9.3005
R18059 gnd.n5927 gnd.n5564 9.3005
R18060 gnd.n5929 gnd.n5928 9.3005
R18061 gnd.n5565 gnd.n5550 9.3005
R18062 gnd.n5945 gnd.n5548 9.3005
R18063 gnd.n5949 gnd.n5948 9.3005
R18064 gnd.n5947 gnd.n5524 9.3005
R18065 gnd.n5984 gnd.n5523 9.3005
R18066 gnd.n5987 gnd.n5986 9.3005
R18067 gnd.n5520 gnd.n5519 9.3005
R18068 gnd.n5993 gnd.n5521 9.3005
R18069 gnd.n5995 gnd.n5994 9.3005
R18070 gnd.n5997 gnd.n5518 9.3005
R18071 gnd.n6000 gnd.n5999 9.3005
R18072 gnd.n6003 gnd.n6001 9.3005
R18073 gnd.n6005 gnd.n6004 9.3005
R18074 gnd.n6011 gnd.n6006 9.3005
R18075 gnd.n6010 gnd.n6009 9.3005
R18076 gnd.n5378 gnd.n5377 9.3005
R18077 gnd.n6077 gnd.n6076 9.3005
R18078 gnd.n6078 gnd.n5371 9.3005
R18079 gnd.n6086 gnd.n5370 9.3005
R18080 gnd.n6089 gnd.n6088 9.3005
R18081 gnd.n6091 gnd.n6090 9.3005
R18082 gnd.n6094 gnd.n5353 9.3005
R18083 gnd.n6092 gnd.n5351 9.3005
R18084 gnd.n6114 gnd.n5349 9.3005
R18085 gnd.n6118 gnd.n6117 9.3005
R18086 gnd.n6116 gnd.n6115 9.3005
R18087 gnd.n5327 gnd.n5326 9.3005
R18088 gnd.n6168 gnd.n5328 9.3005
R18089 gnd.n6170 gnd.n6169 9.3005
R18090 gnd.n6172 gnd.n5325 9.3005
R18091 gnd.n6175 gnd.n6174 9.3005
R18092 gnd.n6177 gnd.n6176 9.3005
R18093 gnd.n6181 gnd.n6178 9.3005
R18094 gnd.n6183 gnd.n6182 9.3005
R18095 gnd.n6468 gnd.n6185 9.3005
R18096 gnd.n6467 gnd.n6187 9.3005
R18097 gnd.n6466 gnd.n6188 9.3005
R18098 gnd.n6463 gnd.n6189 9.3005
R18099 gnd.n6462 gnd.n6190 9.3005
R18100 gnd.n6461 gnd.n6448 9.3005
R18101 gnd.n6458 gnd.n6450 9.3005
R18102 gnd.n6457 gnd.n6451 9.3005
R18103 gnd.n6454 gnd.n6452 9.3005
R18104 gnd.n6453 gnd.n5271 9.3005
R18105 gnd.n5886 gnd.n5885 9.3005
R18106 gnd.n6540 gnd.n5272 9.3005
R18107 gnd.n6539 gnd.n5274 9.3005
R18108 gnd.n5278 gnd.n5275 9.3005
R18109 gnd.n6534 gnd.n5279 9.3005
R18110 gnd.n6533 gnd.n5280 9.3005
R18111 gnd.n6532 gnd.n5281 9.3005
R18112 gnd.n5285 gnd.n5282 9.3005
R18113 gnd.n6527 gnd.n5286 9.3005
R18114 gnd.n6526 gnd.n5287 9.3005
R18115 gnd.n6525 gnd.n5288 9.3005
R18116 gnd.n5292 gnd.n5289 9.3005
R18117 gnd.n6520 gnd.n5293 9.3005
R18118 gnd.n6519 gnd.n5294 9.3005
R18119 gnd.n6518 gnd.n5295 9.3005
R18120 gnd.n5299 gnd.n5296 9.3005
R18121 gnd.n6513 gnd.n5300 9.3005
R18122 gnd.n6512 gnd.n5301 9.3005
R18123 gnd.n6511 gnd.n5302 9.3005
R18124 gnd.n5306 gnd.n5303 9.3005
R18125 gnd.n6506 gnd.n5307 9.3005
R18126 gnd.n6505 gnd.n5308 9.3005
R18127 gnd.n6504 gnd.n5309 9.3005
R18128 gnd.n5316 gnd.n5314 9.3005
R18129 gnd.n6499 gnd.n5317 9.3005
R18130 gnd.n6498 gnd.n5318 9.3005
R18131 gnd.n6497 gnd.n6494 9.3005
R18132 gnd.n6542 gnd.n6541 9.3005
R18133 gnd.n6055 gnd.n6039 9.3005
R18134 gnd.n6054 gnd.n6040 9.3005
R18135 gnd.n6053 gnd.n6041 9.3005
R18136 gnd.n6051 gnd.n6042 9.3005
R18137 gnd.n6050 gnd.n6043 9.3005
R18138 gnd.n6048 gnd.n6044 9.3005
R18139 gnd.n6047 gnd.n6045 9.3005
R18140 gnd.n5341 gnd.n5340 9.3005
R18141 gnd.n6126 gnd.n6125 9.3005
R18142 gnd.n6127 gnd.n5339 9.3005
R18143 gnd.n6153 gnd.n6128 9.3005
R18144 gnd.n6152 gnd.n6129 9.3005
R18145 gnd.n6151 gnd.n6130 9.3005
R18146 gnd.n6149 gnd.n6131 9.3005
R18147 gnd.n6148 gnd.n6132 9.3005
R18148 gnd.n6142 gnd.n6133 9.3005
R18149 gnd.n6141 gnd.n6134 9.3005
R18150 gnd.n6140 gnd.n6135 9.3005
R18151 gnd.n6137 gnd.n6136 9.3005
R18152 gnd.n5324 gnd.n5323 9.3005
R18153 gnd.n6475 gnd.n6474 9.3005
R18154 gnd.n6476 gnd.n5322 9.3005
R18155 gnd.n6480 gnd.n6477 9.3005
R18156 gnd.n6481 gnd.n5321 9.3005
R18157 gnd.n6485 gnd.n6484 9.3005
R18158 gnd.n6486 gnd.n5320 9.3005
R18159 gnd.n6488 gnd.n6487 9.3005
R18160 gnd.n6491 gnd.n5319 9.3005
R18161 gnd.n6493 gnd.n6492 9.3005
R18162 gnd.n5796 gnd.n5795 9.3005
R18163 gnd.n5686 gnd.n5685 9.3005
R18164 gnd.n5810 gnd.n5809 9.3005
R18165 gnd.n5811 gnd.n5684 9.3005
R18166 gnd.n5813 gnd.n5812 9.3005
R18167 gnd.n5674 gnd.n5673 9.3005
R18168 gnd.n5826 gnd.n5825 9.3005
R18169 gnd.n5827 gnd.n5672 9.3005
R18170 gnd.n5859 gnd.n5828 9.3005
R18171 gnd.n5858 gnd.n5829 9.3005
R18172 gnd.n5857 gnd.n5830 9.3005
R18173 gnd.n5856 gnd.n5831 9.3005
R18174 gnd.n5853 gnd.n5832 9.3005
R18175 gnd.n5852 gnd.n5833 9.3005
R18176 gnd.n5851 gnd.n5834 9.3005
R18177 gnd.n5849 gnd.n5835 9.3005
R18178 gnd.n5848 gnd.n5836 9.3005
R18179 gnd.n5845 gnd.n5837 9.3005
R18180 gnd.n5844 gnd.n5838 9.3005
R18181 gnd.n5843 gnd.n5839 9.3005
R18182 gnd.n5841 gnd.n5840 9.3005
R18183 gnd.n5540 gnd.n5539 9.3005
R18184 gnd.n5957 gnd.n5956 9.3005
R18185 gnd.n5958 gnd.n5538 9.3005
R18186 gnd.n5962 gnd.n5959 9.3005
R18187 gnd.n5961 gnd.n5960 9.3005
R18188 gnd.n5462 gnd.n5461 9.3005
R18189 gnd.n6037 gnd.n6036 9.3005
R18190 gnd.n5794 gnd.n5695 9.3005
R18191 gnd.n5697 gnd.n5696 9.3005
R18192 gnd.n5741 gnd.n5739 9.3005
R18193 gnd.n5742 gnd.n5738 9.3005
R18194 gnd.n5745 gnd.n5734 9.3005
R18195 gnd.n5746 gnd.n5733 9.3005
R18196 gnd.n5749 gnd.n5732 9.3005
R18197 gnd.n5750 gnd.n5731 9.3005
R18198 gnd.n5753 gnd.n5730 9.3005
R18199 gnd.n5754 gnd.n5729 9.3005
R18200 gnd.n5757 gnd.n5728 9.3005
R18201 gnd.n5758 gnd.n5727 9.3005
R18202 gnd.n5761 gnd.n5726 9.3005
R18203 gnd.n5762 gnd.n5725 9.3005
R18204 gnd.n5765 gnd.n5724 9.3005
R18205 gnd.n5766 gnd.n5723 9.3005
R18206 gnd.n5769 gnd.n5722 9.3005
R18207 gnd.n5770 gnd.n5721 9.3005
R18208 gnd.n5773 gnd.n5720 9.3005
R18209 gnd.n5774 gnd.n5719 9.3005
R18210 gnd.n5777 gnd.n5718 9.3005
R18211 gnd.n5778 gnd.n5717 9.3005
R18212 gnd.n5781 gnd.n5716 9.3005
R18213 gnd.n5783 gnd.n5715 9.3005
R18214 gnd.n5784 gnd.n5714 9.3005
R18215 gnd.n5785 gnd.n5713 9.3005
R18216 gnd.n5786 gnd.n5712 9.3005
R18217 gnd.n5793 gnd.n5792 9.3005
R18218 gnd.n5802 gnd.n5801 9.3005
R18219 gnd.n5803 gnd.n5689 9.3005
R18220 gnd.n5805 gnd.n5804 9.3005
R18221 gnd.n5680 gnd.n5679 9.3005
R18222 gnd.n5818 gnd.n5817 9.3005
R18223 gnd.n5819 gnd.n5678 9.3005
R18224 gnd.n5821 gnd.n5820 9.3005
R18225 gnd.n5667 gnd.n5666 9.3005
R18226 gnd.n5864 gnd.n5863 9.3005
R18227 gnd.n5865 gnd.n5621 9.3005
R18228 gnd.n5869 gnd.n5867 9.3005
R18229 gnd.n5868 gnd.n5600 9.3005
R18230 gnd.n5887 gnd.n5599 9.3005
R18231 gnd.n5890 gnd.n5889 9.3005
R18232 gnd.n5593 gnd.n5592 9.3005
R18233 gnd.n5901 gnd.n5899 9.3005
R18234 gnd.n5900 gnd.n5574 9.3005
R18235 gnd.n5918 gnd.n5573 9.3005
R18236 gnd.n5921 gnd.n5920 9.3005
R18237 gnd.n5568 gnd.n5563 9.3005
R18238 gnd.n5931 gnd.n5930 9.3005
R18239 gnd.n5566 gnd.n5546 9.3005
R18240 gnd.n5952 gnd.n5547 9.3005
R18241 gnd.n5951 gnd.n5950 9.3005
R18242 gnd.n5549 gnd.n5525 9.3005
R18243 gnd.n5983 gnd.n5982 9.3005
R18244 gnd.n5985 gnd.n5470 9.3005
R18245 gnd.n6032 gnd.n5471 9.3005
R18246 gnd.n6031 gnd.n5472 9.3005
R18247 gnd.n6030 gnd.n5473 9.3005
R18248 gnd.n5996 gnd.n5474 9.3005
R18249 gnd.n5998 gnd.n5492 9.3005
R18250 gnd.n6018 gnd.n5493 9.3005
R18251 gnd.n6017 gnd.n5494 9.3005
R18252 gnd.n6016 gnd.n5495 9.3005
R18253 gnd.n6007 gnd.n5496 9.3005
R18254 gnd.n6008 gnd.n5379 9.3005
R18255 gnd.n6074 gnd.n6073 9.3005
R18256 gnd.n6075 gnd.n5372 9.3005
R18257 gnd.n6085 gnd.n6084 9.3005
R18258 gnd.n6087 gnd.n5368 9.3005
R18259 gnd.n6097 gnd.n5369 9.3005
R18260 gnd.n6096 gnd.n6095 9.3005
R18261 gnd.n6093 gnd.n5347 9.3005
R18262 gnd.n6121 gnd.n5348 9.3005
R18263 gnd.n6120 gnd.n6119 9.3005
R18264 gnd.n5350 gnd.n1043 9.3005
R18265 gnd.n6625 gnd.n1044 9.3005
R18266 gnd.n6624 gnd.n1045 9.3005
R18267 gnd.n6623 gnd.n1046 9.3005
R18268 gnd.n6171 gnd.n1047 9.3005
R18269 gnd.n6173 gnd.n1066 9.3005
R18270 gnd.n6611 gnd.n1067 9.3005
R18271 gnd.n6610 gnd.n1068 9.3005
R18272 gnd.n6609 gnd.n1069 9.3005
R18273 gnd.n6184 gnd.n1070 9.3005
R18274 gnd.n6186 gnd.n1091 9.3005
R18275 gnd.n6597 gnd.n1092 9.3005
R18276 gnd.n6596 gnd.n1093 9.3005
R18277 gnd.n6595 gnd.n1094 9.3005
R18278 gnd.n6447 gnd.n1095 9.3005
R18279 gnd.n6449 gnd.n1117 9.3005
R18280 gnd.n6583 gnd.n1118 9.3005
R18281 gnd.n6582 gnd.n1119 9.3005
R18282 gnd.n6581 gnd.n1120 9.3005
R18283 gnd.n5691 gnd.n5690 9.3005
R18284 gnd.n870 gnd.n869 9.3005
R18285 gnd.n6801 gnd.n6800 9.3005
R18286 gnd.n6802 gnd.n868 9.3005
R18287 gnd.n6804 gnd.n6803 9.3005
R18288 gnd.n864 gnd.n863 9.3005
R18289 gnd.n6811 gnd.n6810 9.3005
R18290 gnd.n6812 gnd.n862 9.3005
R18291 gnd.n6814 gnd.n6813 9.3005
R18292 gnd.n858 gnd.n857 9.3005
R18293 gnd.n6821 gnd.n6820 9.3005
R18294 gnd.n6822 gnd.n856 9.3005
R18295 gnd.n6824 gnd.n6823 9.3005
R18296 gnd.n852 gnd.n851 9.3005
R18297 gnd.n6831 gnd.n6830 9.3005
R18298 gnd.n6832 gnd.n850 9.3005
R18299 gnd.n6834 gnd.n6833 9.3005
R18300 gnd.n846 gnd.n845 9.3005
R18301 gnd.n6841 gnd.n6840 9.3005
R18302 gnd.n6842 gnd.n844 9.3005
R18303 gnd.n6844 gnd.n6843 9.3005
R18304 gnd.n840 gnd.n839 9.3005
R18305 gnd.n6851 gnd.n6850 9.3005
R18306 gnd.n6852 gnd.n838 9.3005
R18307 gnd.n6854 gnd.n6853 9.3005
R18308 gnd.n834 gnd.n833 9.3005
R18309 gnd.n6861 gnd.n6860 9.3005
R18310 gnd.n6862 gnd.n832 9.3005
R18311 gnd.n6864 gnd.n6863 9.3005
R18312 gnd.n828 gnd.n827 9.3005
R18313 gnd.n6871 gnd.n6870 9.3005
R18314 gnd.n6872 gnd.n826 9.3005
R18315 gnd.n6874 gnd.n6873 9.3005
R18316 gnd.n822 gnd.n821 9.3005
R18317 gnd.n6881 gnd.n6880 9.3005
R18318 gnd.n6882 gnd.n820 9.3005
R18319 gnd.n6884 gnd.n6883 9.3005
R18320 gnd.n816 gnd.n815 9.3005
R18321 gnd.n6891 gnd.n6890 9.3005
R18322 gnd.n6892 gnd.n814 9.3005
R18323 gnd.n6894 gnd.n6893 9.3005
R18324 gnd.n810 gnd.n809 9.3005
R18325 gnd.n6901 gnd.n6900 9.3005
R18326 gnd.n6902 gnd.n808 9.3005
R18327 gnd.n6904 gnd.n6903 9.3005
R18328 gnd.n804 gnd.n803 9.3005
R18329 gnd.n6911 gnd.n6910 9.3005
R18330 gnd.n6912 gnd.n802 9.3005
R18331 gnd.n6914 gnd.n6913 9.3005
R18332 gnd.n798 gnd.n797 9.3005
R18333 gnd.n6921 gnd.n6920 9.3005
R18334 gnd.n6922 gnd.n796 9.3005
R18335 gnd.n6924 gnd.n6923 9.3005
R18336 gnd.n792 gnd.n791 9.3005
R18337 gnd.n6931 gnd.n6930 9.3005
R18338 gnd.n6932 gnd.n790 9.3005
R18339 gnd.n6934 gnd.n6933 9.3005
R18340 gnd.n786 gnd.n785 9.3005
R18341 gnd.n6941 gnd.n6940 9.3005
R18342 gnd.n6942 gnd.n784 9.3005
R18343 gnd.n6944 gnd.n6943 9.3005
R18344 gnd.n780 gnd.n779 9.3005
R18345 gnd.n6951 gnd.n6950 9.3005
R18346 gnd.n6952 gnd.n778 9.3005
R18347 gnd.n6954 gnd.n6953 9.3005
R18348 gnd.n774 gnd.n773 9.3005
R18349 gnd.n6961 gnd.n6960 9.3005
R18350 gnd.n6962 gnd.n772 9.3005
R18351 gnd.n6964 gnd.n6963 9.3005
R18352 gnd.n768 gnd.n767 9.3005
R18353 gnd.n6971 gnd.n6970 9.3005
R18354 gnd.n6972 gnd.n766 9.3005
R18355 gnd.n6974 gnd.n6973 9.3005
R18356 gnd.n762 gnd.n761 9.3005
R18357 gnd.n6981 gnd.n6980 9.3005
R18358 gnd.n6982 gnd.n760 9.3005
R18359 gnd.n6984 gnd.n6983 9.3005
R18360 gnd.n756 gnd.n755 9.3005
R18361 gnd.n6991 gnd.n6990 9.3005
R18362 gnd.n6992 gnd.n754 9.3005
R18363 gnd.n6994 gnd.n6993 9.3005
R18364 gnd.n750 gnd.n749 9.3005
R18365 gnd.n7001 gnd.n7000 9.3005
R18366 gnd.n7002 gnd.n748 9.3005
R18367 gnd.n7004 gnd.n7003 9.3005
R18368 gnd.n744 gnd.n743 9.3005
R18369 gnd.n7011 gnd.n7010 9.3005
R18370 gnd.n7012 gnd.n742 9.3005
R18371 gnd.n7014 gnd.n7013 9.3005
R18372 gnd.n738 gnd.n737 9.3005
R18373 gnd.n7021 gnd.n7020 9.3005
R18374 gnd.n7022 gnd.n736 9.3005
R18375 gnd.n7024 gnd.n7023 9.3005
R18376 gnd.n732 gnd.n731 9.3005
R18377 gnd.n7031 gnd.n7030 9.3005
R18378 gnd.n7032 gnd.n730 9.3005
R18379 gnd.n7034 gnd.n7033 9.3005
R18380 gnd.n726 gnd.n725 9.3005
R18381 gnd.n7041 gnd.n7040 9.3005
R18382 gnd.n7042 gnd.n724 9.3005
R18383 gnd.n7044 gnd.n7043 9.3005
R18384 gnd.n720 gnd.n719 9.3005
R18385 gnd.n7051 gnd.n7050 9.3005
R18386 gnd.n7052 gnd.n718 9.3005
R18387 gnd.n7054 gnd.n7053 9.3005
R18388 gnd.n714 gnd.n713 9.3005
R18389 gnd.n7061 gnd.n7060 9.3005
R18390 gnd.n7062 gnd.n712 9.3005
R18391 gnd.n7064 gnd.n7063 9.3005
R18392 gnd.n708 gnd.n707 9.3005
R18393 gnd.n7071 gnd.n7070 9.3005
R18394 gnd.n7072 gnd.n706 9.3005
R18395 gnd.n7074 gnd.n7073 9.3005
R18396 gnd.n702 gnd.n701 9.3005
R18397 gnd.n7081 gnd.n7080 9.3005
R18398 gnd.n7082 gnd.n700 9.3005
R18399 gnd.n7084 gnd.n7083 9.3005
R18400 gnd.n696 gnd.n695 9.3005
R18401 gnd.n7091 gnd.n7090 9.3005
R18402 gnd.n7092 gnd.n694 9.3005
R18403 gnd.n7094 gnd.n7093 9.3005
R18404 gnd.n690 gnd.n689 9.3005
R18405 gnd.n7101 gnd.n7100 9.3005
R18406 gnd.n7102 gnd.n688 9.3005
R18407 gnd.n7104 gnd.n7103 9.3005
R18408 gnd.n684 gnd.n683 9.3005
R18409 gnd.n7111 gnd.n7110 9.3005
R18410 gnd.n7112 gnd.n682 9.3005
R18411 gnd.n7114 gnd.n7113 9.3005
R18412 gnd.n678 gnd.n677 9.3005
R18413 gnd.n7121 gnd.n7120 9.3005
R18414 gnd.n7122 gnd.n676 9.3005
R18415 gnd.n7124 gnd.n7123 9.3005
R18416 gnd.n672 gnd.n671 9.3005
R18417 gnd.n7131 gnd.n7130 9.3005
R18418 gnd.n7132 gnd.n670 9.3005
R18419 gnd.n7134 gnd.n7133 9.3005
R18420 gnd.n666 gnd.n665 9.3005
R18421 gnd.n7141 gnd.n7140 9.3005
R18422 gnd.n7142 gnd.n664 9.3005
R18423 gnd.n7144 gnd.n7143 9.3005
R18424 gnd.n660 gnd.n659 9.3005
R18425 gnd.n7151 gnd.n7150 9.3005
R18426 gnd.n7152 gnd.n658 9.3005
R18427 gnd.n7154 gnd.n7153 9.3005
R18428 gnd.n654 gnd.n653 9.3005
R18429 gnd.n7161 gnd.n7160 9.3005
R18430 gnd.n7162 gnd.n652 9.3005
R18431 gnd.n7164 gnd.n7163 9.3005
R18432 gnd.n648 gnd.n647 9.3005
R18433 gnd.n7171 gnd.n7170 9.3005
R18434 gnd.n7172 gnd.n646 9.3005
R18435 gnd.n7174 gnd.n7173 9.3005
R18436 gnd.n642 gnd.n641 9.3005
R18437 gnd.n7181 gnd.n7180 9.3005
R18438 gnd.n7182 gnd.n640 9.3005
R18439 gnd.n7184 gnd.n7183 9.3005
R18440 gnd.n636 gnd.n635 9.3005
R18441 gnd.n7191 gnd.n7190 9.3005
R18442 gnd.n7192 gnd.n634 9.3005
R18443 gnd.n7194 gnd.n7193 9.3005
R18444 gnd.n630 gnd.n629 9.3005
R18445 gnd.n7201 gnd.n7200 9.3005
R18446 gnd.n7202 gnd.n628 9.3005
R18447 gnd.n7204 gnd.n7203 9.3005
R18448 gnd.n624 gnd.n623 9.3005
R18449 gnd.n7211 gnd.n7210 9.3005
R18450 gnd.n7212 gnd.n622 9.3005
R18451 gnd.n7214 gnd.n7213 9.3005
R18452 gnd.n618 gnd.n617 9.3005
R18453 gnd.n7221 gnd.n7220 9.3005
R18454 gnd.n7222 gnd.n616 9.3005
R18455 gnd.n7224 gnd.n7223 9.3005
R18456 gnd.n612 gnd.n611 9.3005
R18457 gnd.n7231 gnd.n7230 9.3005
R18458 gnd.n7232 gnd.n610 9.3005
R18459 gnd.n7234 gnd.n7233 9.3005
R18460 gnd.n606 gnd.n605 9.3005
R18461 gnd.n7241 gnd.n7240 9.3005
R18462 gnd.n7242 gnd.n604 9.3005
R18463 gnd.n7244 gnd.n7243 9.3005
R18464 gnd.n600 gnd.n599 9.3005
R18465 gnd.n7251 gnd.n7250 9.3005
R18466 gnd.n7252 gnd.n598 9.3005
R18467 gnd.n7254 gnd.n7253 9.3005
R18468 gnd.n594 gnd.n593 9.3005
R18469 gnd.n7261 gnd.n7260 9.3005
R18470 gnd.n7262 gnd.n592 9.3005
R18471 gnd.n7264 gnd.n7263 9.3005
R18472 gnd.n588 gnd.n587 9.3005
R18473 gnd.n7271 gnd.n7270 9.3005
R18474 gnd.n7272 gnd.n586 9.3005
R18475 gnd.n7274 gnd.n7273 9.3005
R18476 gnd.n582 gnd.n581 9.3005
R18477 gnd.n7281 gnd.n7280 9.3005
R18478 gnd.n7282 gnd.n580 9.3005
R18479 gnd.n7284 gnd.n7283 9.3005
R18480 gnd.n576 gnd.n575 9.3005
R18481 gnd.n7291 gnd.n7290 9.3005
R18482 gnd.n7292 gnd.n574 9.3005
R18483 gnd.n7294 gnd.n7293 9.3005
R18484 gnd.n570 gnd.n569 9.3005
R18485 gnd.n7301 gnd.n7300 9.3005
R18486 gnd.n7302 gnd.n568 9.3005
R18487 gnd.n7304 gnd.n7303 9.3005
R18488 gnd.n564 gnd.n563 9.3005
R18489 gnd.n7311 gnd.n7310 9.3005
R18490 gnd.n7312 gnd.n562 9.3005
R18491 gnd.n7314 gnd.n7313 9.3005
R18492 gnd.n7321 gnd.n7320 9.3005
R18493 gnd.n7322 gnd.n556 9.3005
R18494 gnd.n7324 gnd.n7323 9.3005
R18495 gnd.n552 gnd.n551 9.3005
R18496 gnd.n7331 gnd.n7330 9.3005
R18497 gnd.n7332 gnd.n550 9.3005
R18498 gnd.n7334 gnd.n7333 9.3005
R18499 gnd.n546 gnd.n545 9.3005
R18500 gnd.n7341 gnd.n7340 9.3005
R18501 gnd.n7342 gnd.n544 9.3005
R18502 gnd.n7344 gnd.n7343 9.3005
R18503 gnd.n540 gnd.n539 9.3005
R18504 gnd.n7351 gnd.n7350 9.3005
R18505 gnd.n7352 gnd.n538 9.3005
R18506 gnd.n7354 gnd.n7353 9.3005
R18507 gnd.n534 gnd.n533 9.3005
R18508 gnd.n7361 gnd.n7360 9.3005
R18509 gnd.n7362 gnd.n532 9.3005
R18510 gnd.n7364 gnd.n7363 9.3005
R18511 gnd.n528 gnd.n527 9.3005
R18512 gnd.n7371 gnd.n7370 9.3005
R18513 gnd.n7372 gnd.n526 9.3005
R18514 gnd.n7374 gnd.n7373 9.3005
R18515 gnd.n522 gnd.n521 9.3005
R18516 gnd.n7381 gnd.n7380 9.3005
R18517 gnd.n7382 gnd.n520 9.3005
R18518 gnd.n7384 gnd.n7383 9.3005
R18519 gnd.n516 gnd.n515 9.3005
R18520 gnd.n7391 gnd.n7390 9.3005
R18521 gnd.n7392 gnd.n514 9.3005
R18522 gnd.n7394 gnd.n7393 9.3005
R18523 gnd.n510 gnd.n509 9.3005
R18524 gnd.n7401 gnd.n7400 9.3005
R18525 gnd.n7402 gnd.n508 9.3005
R18526 gnd.n7404 gnd.n7403 9.3005
R18527 gnd.n504 gnd.n503 9.3005
R18528 gnd.n7411 gnd.n7410 9.3005
R18529 gnd.n7412 gnd.n502 9.3005
R18530 gnd.n7414 gnd.n7413 9.3005
R18531 gnd.n498 gnd.n497 9.3005
R18532 gnd.n7421 gnd.n7420 9.3005
R18533 gnd.n7422 gnd.n496 9.3005
R18534 gnd.n7424 gnd.n7423 9.3005
R18535 gnd.n492 gnd.n491 9.3005
R18536 gnd.n7431 gnd.n7430 9.3005
R18537 gnd.n7432 gnd.n490 9.3005
R18538 gnd.n7434 gnd.n7433 9.3005
R18539 gnd.n486 gnd.n485 9.3005
R18540 gnd.n7441 gnd.n7440 9.3005
R18541 gnd.n7442 gnd.n484 9.3005
R18542 gnd.n7444 gnd.n7443 9.3005
R18543 gnd.n480 gnd.n479 9.3005
R18544 gnd.n7451 gnd.n7450 9.3005
R18545 gnd.n7452 gnd.n478 9.3005
R18546 gnd.n7454 gnd.n7453 9.3005
R18547 gnd.n474 gnd.n473 9.3005
R18548 gnd.n7461 gnd.n7460 9.3005
R18549 gnd.n7462 gnd.n472 9.3005
R18550 gnd.n7464 gnd.n7463 9.3005
R18551 gnd.n468 gnd.n467 9.3005
R18552 gnd.n7471 gnd.n7470 9.3005
R18553 gnd.n7472 gnd.n466 9.3005
R18554 gnd.n7474 gnd.n7473 9.3005
R18555 gnd.n462 gnd.n461 9.3005
R18556 gnd.n7481 gnd.n7480 9.3005
R18557 gnd.n7482 gnd.n460 9.3005
R18558 gnd.n7484 gnd.n7483 9.3005
R18559 gnd.n456 gnd.n455 9.3005
R18560 gnd.n7491 gnd.n7490 9.3005
R18561 gnd.n7492 gnd.n454 9.3005
R18562 gnd.n7494 gnd.n7493 9.3005
R18563 gnd.n450 gnd.n449 9.3005
R18564 gnd.n7501 gnd.n7500 9.3005
R18565 gnd.n7502 gnd.n448 9.3005
R18566 gnd.n7504 gnd.n7503 9.3005
R18567 gnd.n444 gnd.n443 9.3005
R18568 gnd.n7511 gnd.n7510 9.3005
R18569 gnd.n7512 gnd.n442 9.3005
R18570 gnd.n7514 gnd.n7513 9.3005
R18571 gnd.n438 gnd.n437 9.3005
R18572 gnd.n7521 gnd.n7520 9.3005
R18573 gnd.n7522 gnd.n436 9.3005
R18574 gnd.n7526 gnd.n7523 9.3005
R18575 gnd.n7525 gnd.n7524 9.3005
R18576 gnd.n558 gnd.n557 9.3005
R18577 gnd.n7885 gnd.n7884 9.3005
R18578 gnd.n7883 gnd.n80 9.3005
R18579 gnd.n7574 gnd.n83 9.3005
R18580 gnd.n7576 gnd.n7575 9.3005
R18581 gnd.n387 gnd.n386 9.3005
R18582 gnd.n7587 gnd.n7586 9.3005
R18583 gnd.n7588 gnd.n385 9.3005
R18584 gnd.n7590 gnd.n7589 9.3005
R18585 gnd.n380 gnd.n379 9.3005
R18586 gnd.n7601 gnd.n7600 9.3005
R18587 gnd.n7602 gnd.n378 9.3005
R18588 gnd.n7604 gnd.n7603 9.3005
R18589 gnd.n375 gnd.n374 9.3005
R18590 gnd.n7615 gnd.n7614 9.3005
R18591 gnd.n7616 gnd.n373 9.3005
R18592 gnd.n7618 gnd.n7617 9.3005
R18593 gnd.n368 gnd.n367 9.3005
R18594 gnd.n7629 gnd.n7628 9.3005
R18595 gnd.n7630 gnd.n366 9.3005
R18596 gnd.n7632 gnd.n7631 9.3005
R18597 gnd.n363 gnd.n362 9.3005
R18598 gnd.n7643 gnd.n7642 9.3005
R18599 gnd.n7644 gnd.n361 9.3005
R18600 gnd.n7647 gnd.n7646 9.3005
R18601 gnd.n7645 gnd.n357 9.3005
R18602 gnd.n7658 gnd.n356 9.3005
R18603 gnd.n7660 gnd.n7659 9.3005
R18604 gnd.n7691 gnd.n322 9.3005
R18605 gnd.n7690 gnd.n324 9.3005
R18606 gnd.n328 gnd.n325 9.3005
R18607 gnd.n7685 gnd.n329 9.3005
R18608 gnd.n7684 gnd.n330 9.3005
R18609 gnd.n7683 gnd.n331 9.3005
R18610 gnd.n335 gnd.n332 9.3005
R18611 gnd.n7678 gnd.n336 9.3005
R18612 gnd.n7677 gnd.n337 9.3005
R18613 gnd.n7676 gnd.n338 9.3005
R18614 gnd.n342 gnd.n339 9.3005
R18615 gnd.n7671 gnd.n343 9.3005
R18616 gnd.n7670 gnd.n344 9.3005
R18617 gnd.n7669 gnd.n345 9.3005
R18618 gnd.n349 gnd.n346 9.3005
R18619 gnd.n7664 gnd.n350 9.3005
R18620 gnd.n7663 gnd.n7662 9.3005
R18621 gnd.n7661 gnd.n353 9.3005
R18622 gnd.n7693 gnd.n7692 9.3005
R18623 gnd.n7801 gnd.n218 9.3005
R18624 gnd.n7800 gnd.n220 9.3005
R18625 gnd.n225 gnd.n221 9.3005
R18626 gnd.n7795 gnd.n226 9.3005
R18627 gnd.n7794 gnd.n227 9.3005
R18628 gnd.n7793 gnd.n228 9.3005
R18629 gnd.n232 gnd.n229 9.3005
R18630 gnd.n7788 gnd.n233 9.3005
R18631 gnd.n7787 gnd.n234 9.3005
R18632 gnd.n7786 gnd.n235 9.3005
R18633 gnd.n239 gnd.n236 9.3005
R18634 gnd.n7781 gnd.n240 9.3005
R18635 gnd.n7780 gnd.n241 9.3005
R18636 gnd.n7779 gnd.n242 9.3005
R18637 gnd.n246 gnd.n243 9.3005
R18638 gnd.n7774 gnd.n247 9.3005
R18639 gnd.n7773 gnd.n248 9.3005
R18640 gnd.n7769 gnd.n249 9.3005
R18641 gnd.n253 gnd.n250 9.3005
R18642 gnd.n7764 gnd.n254 9.3005
R18643 gnd.n7763 gnd.n255 9.3005
R18644 gnd.n7762 gnd.n256 9.3005
R18645 gnd.n260 gnd.n257 9.3005
R18646 gnd.n7757 gnd.n261 9.3005
R18647 gnd.n7756 gnd.n262 9.3005
R18648 gnd.n7755 gnd.n263 9.3005
R18649 gnd.n267 gnd.n264 9.3005
R18650 gnd.n7750 gnd.n268 9.3005
R18651 gnd.n7749 gnd.n269 9.3005
R18652 gnd.n7748 gnd.n270 9.3005
R18653 gnd.n274 gnd.n271 9.3005
R18654 gnd.n7743 gnd.n275 9.3005
R18655 gnd.n7742 gnd.n276 9.3005
R18656 gnd.n7741 gnd.n277 9.3005
R18657 gnd.n281 gnd.n278 9.3005
R18658 gnd.n7736 gnd.n282 9.3005
R18659 gnd.n7735 gnd.n7734 9.3005
R18660 gnd.n7733 gnd.n283 9.3005
R18661 gnd.n7732 gnd.n7731 9.3005
R18662 gnd.n287 gnd.n286 9.3005
R18663 gnd.n292 gnd.n290 9.3005
R18664 gnd.n7724 gnd.n293 9.3005
R18665 gnd.n7723 gnd.n294 9.3005
R18666 gnd.n7722 gnd.n295 9.3005
R18667 gnd.n299 gnd.n296 9.3005
R18668 gnd.n7717 gnd.n300 9.3005
R18669 gnd.n7716 gnd.n301 9.3005
R18670 gnd.n7715 gnd.n302 9.3005
R18671 gnd.n306 gnd.n303 9.3005
R18672 gnd.n7710 gnd.n307 9.3005
R18673 gnd.n7709 gnd.n308 9.3005
R18674 gnd.n7708 gnd.n309 9.3005
R18675 gnd.n313 gnd.n310 9.3005
R18676 gnd.n7703 gnd.n314 9.3005
R18677 gnd.n7702 gnd.n315 9.3005
R18678 gnd.n7701 gnd.n316 9.3005
R18679 gnd.n321 gnd.n319 9.3005
R18680 gnd.n7696 gnd.n7695 9.3005
R18681 gnd.n7803 gnd.n7802 9.3005
R18682 gnd.n4492 gnd.n1742 9.3005
R18683 gnd.n4702 gnd.n1743 9.3005
R18684 gnd.n4701 gnd.n1744 9.3005
R18685 gnd.n4700 gnd.n1745 9.3005
R18686 gnd.n1927 gnd.n1746 9.3005
R18687 gnd.n4690 gnd.n1763 9.3005
R18688 gnd.n4689 gnd.n1764 9.3005
R18689 gnd.n4688 gnd.n1765 9.3005
R18690 gnd.n1890 gnd.n1766 9.3005
R18691 gnd.n4678 gnd.n1784 9.3005
R18692 gnd.n4677 gnd.n1785 9.3005
R18693 gnd.n4676 gnd.n1786 9.3005
R18694 gnd.n4525 gnd.n1787 9.3005
R18695 gnd.n4666 gnd.n1803 9.3005
R18696 gnd.n4665 gnd.n1804 9.3005
R18697 gnd.n4664 gnd.n1805 9.3005
R18698 gnd.n4535 gnd.n1806 9.3005
R18699 gnd.n4654 gnd.n1824 9.3005
R18700 gnd.n4653 gnd.n1825 9.3005
R18701 gnd.n4652 gnd.n1826 9.3005
R18702 gnd.n4583 gnd.n1827 9.3005
R18703 gnd.n4642 gnd.n1841 9.3005
R18704 gnd.n4641 gnd.n1842 9.3005
R18705 gnd.n4640 gnd.n1843 9.3005
R18706 gnd.n4584 gnd.n1844 9.3005
R18707 gnd.n4589 gnd.n4585 9.3005
R18708 gnd.n4597 gnd.n4590 9.3005
R18709 gnd.n4596 gnd.n4592 9.3005
R18710 gnd.n4595 gnd.n4593 9.3005
R18711 gnd.n389 gnd.n108 9.3005
R18712 gnd.n7871 gnd.n109 9.3005
R18713 gnd.n7870 gnd.n110 9.3005
R18714 gnd.n7869 gnd.n111 9.3005
R18715 gnd.n383 gnd.n112 9.3005
R18716 gnd.n7859 gnd.n127 9.3005
R18717 gnd.n7858 gnd.n128 9.3005
R18718 gnd.n7857 gnd.n129 9.3005
R18719 gnd.n377 gnd.n130 9.3005
R18720 gnd.n7847 gnd.n148 9.3005
R18721 gnd.n7846 gnd.n149 9.3005
R18722 gnd.n7845 gnd.n150 9.3005
R18723 gnd.n371 gnd.n151 9.3005
R18724 gnd.n7835 gnd.n167 9.3005
R18725 gnd.n7834 gnd.n168 9.3005
R18726 gnd.n7833 gnd.n169 9.3005
R18727 gnd.n365 gnd.n170 9.3005
R18728 gnd.n7823 gnd.n188 9.3005
R18729 gnd.n7822 gnd.n189 9.3005
R18730 gnd.n7821 gnd.n190 9.3005
R18731 gnd.n360 gnd.n191 9.3005
R18732 gnd.n7811 gnd.n208 9.3005
R18733 gnd.n7810 gnd.n209 9.3005
R18734 gnd.n7809 gnd.n210 9.3005
R18735 gnd.n4491 gnd.n4490 9.3005
R18736 gnd.n4493 gnd.n4492 9.3005
R18737 gnd.n4494 gnd.n1743 9.3005
R18738 gnd.n4495 gnd.n1744 9.3005
R18739 gnd.n1926 gnd.n1745 9.3005
R18740 gnd.n4507 gnd.n1927 9.3005
R18741 gnd.n4508 gnd.n1763 9.3005
R18742 gnd.n4509 gnd.n1764 9.3005
R18743 gnd.n1889 gnd.n1765 9.3005
R18744 gnd.n4521 gnd.n1890 9.3005
R18745 gnd.n4522 gnd.n1784 9.3005
R18746 gnd.n4523 gnd.n1785 9.3005
R18747 gnd.n4524 gnd.n1786 9.3005
R18748 gnd.n4528 gnd.n4525 9.3005
R18749 gnd.n4529 gnd.n1803 9.3005
R18750 gnd.n4533 gnd.n1804 9.3005
R18751 gnd.n4534 gnd.n1805 9.3005
R18752 gnd.n4536 gnd.n4535 9.3005
R18753 gnd.n1867 gnd.n1824 9.3005
R18754 gnd.n4581 gnd.n1825 9.3005
R18755 gnd.n4582 gnd.n1826 9.3005
R18756 gnd.n4607 gnd.n4583 9.3005
R18757 gnd.n4606 gnd.n1841 9.3005
R18758 gnd.n4605 gnd.n1842 9.3005
R18759 gnd.n4604 gnd.n1843 9.3005
R18760 gnd.n4603 gnd.n4584 9.3005
R18761 gnd.n4602 gnd.n4585 9.3005
R18762 gnd.n4590 gnd.n4586 9.3005
R18763 gnd.n4592 gnd.n4591 9.3005
R18764 gnd.n4593 gnd.n388 9.3005
R18765 gnd.n7580 gnd.n389 9.3005
R18766 gnd.n7581 gnd.n109 9.3005
R18767 gnd.n7582 gnd.n110 9.3005
R18768 gnd.n382 gnd.n111 9.3005
R18769 gnd.n7594 gnd.n383 9.3005
R18770 gnd.n7595 gnd.n127 9.3005
R18771 gnd.n7596 gnd.n128 9.3005
R18772 gnd.n376 gnd.n129 9.3005
R18773 gnd.n7608 gnd.n377 9.3005
R18774 gnd.n7609 gnd.n148 9.3005
R18775 gnd.n7610 gnd.n149 9.3005
R18776 gnd.n370 gnd.n150 9.3005
R18777 gnd.n7622 gnd.n371 9.3005
R18778 gnd.n7623 gnd.n167 9.3005
R18779 gnd.n7624 gnd.n168 9.3005
R18780 gnd.n364 gnd.n169 9.3005
R18781 gnd.n7636 gnd.n365 9.3005
R18782 gnd.n7637 gnd.n188 9.3005
R18783 gnd.n7638 gnd.n189 9.3005
R18784 gnd.n359 gnd.n190 9.3005
R18785 gnd.n7651 gnd.n360 9.3005
R18786 gnd.n7652 gnd.n208 9.3005
R18787 gnd.n7654 gnd.n209 9.3005
R18788 gnd.n7653 gnd.n210 9.3005
R18789 gnd.n4491 gnd.n1931 9.3005
R18790 gnd.n1937 gnd.n1934 9.3005
R18791 gnd.n4478 gnd.n1938 9.3005
R18792 gnd.n4480 gnd.n4479 9.3005
R18793 gnd.n4477 gnd.n1940 9.3005
R18794 gnd.n4476 gnd.n4475 9.3005
R18795 gnd.n1942 gnd.n1941 9.3005
R18796 gnd.n4469 gnd.n4468 9.3005
R18797 gnd.n4467 gnd.n1944 9.3005
R18798 gnd.n4466 gnd.n4465 9.3005
R18799 gnd.n1946 gnd.n1945 9.3005
R18800 gnd.n4459 gnd.n4458 9.3005
R18801 gnd.n4457 gnd.n1948 9.3005
R18802 gnd.n4456 gnd.n4455 9.3005
R18803 gnd.n1950 gnd.n1949 9.3005
R18804 gnd.n4449 gnd.n4448 9.3005
R18805 gnd.n4447 gnd.n1952 9.3005
R18806 gnd.n4446 gnd.n4445 9.3005
R18807 gnd.n1954 gnd.n1953 9.3005
R18808 gnd.n4439 gnd.n4438 9.3005
R18809 gnd.n4437 gnd.n1956 9.3005
R18810 gnd.n1958 gnd.n1957 9.3005
R18811 gnd.n4427 gnd.n4426 9.3005
R18812 gnd.n4425 gnd.n1960 9.3005
R18813 gnd.n4424 gnd.n4423 9.3005
R18814 gnd.n1962 gnd.n1961 9.3005
R18815 gnd.n4417 gnd.n4416 9.3005
R18816 gnd.n4415 gnd.n1964 9.3005
R18817 gnd.n4414 gnd.n4413 9.3005
R18818 gnd.n1966 gnd.n1965 9.3005
R18819 gnd.n4405 gnd.n4404 9.3005
R18820 gnd.n4402 gnd.n4315 9.3005
R18821 gnd.n4401 gnd.n4400 9.3005
R18822 gnd.n4317 gnd.n4316 9.3005
R18823 gnd.n4394 gnd.n4393 9.3005
R18824 gnd.n4392 gnd.n4319 9.3005
R18825 gnd.n4391 gnd.n4390 9.3005
R18826 gnd.n4321 gnd.n4320 9.3005
R18827 gnd.n4384 gnd.n4380 9.3005
R18828 gnd.n4379 gnd.n4323 9.3005
R18829 gnd.n4378 gnd.n4377 9.3005
R18830 gnd.n4325 gnd.n4324 9.3005
R18831 gnd.n4371 gnd.n4370 9.3005
R18832 gnd.n4369 gnd.n4327 9.3005
R18833 gnd.n4368 gnd.n4367 9.3005
R18834 gnd.n4329 gnd.n4328 9.3005
R18835 gnd.n4361 gnd.n4360 9.3005
R18836 gnd.n4359 gnd.n4331 9.3005
R18837 gnd.n4358 gnd.n4357 9.3005
R18838 gnd.n4333 gnd.n4332 9.3005
R18839 gnd.n4351 gnd.n4350 9.3005
R18840 gnd.n4349 gnd.n4335 9.3005
R18841 gnd.n4348 gnd.n4347 9.3005
R18842 gnd.n4337 gnd.n4336 9.3005
R18843 gnd.n4341 gnd.n4340 9.3005
R18844 gnd.n4339 gnd.n4338 9.3005
R18845 gnd.n4436 gnd.n4435 9.3005
R18846 gnd.n4488 gnd.n4487 9.3005
R18847 gnd.n4707 gnd.n1732 9.3005
R18848 gnd.n4706 gnd.n1733 9.3005
R18849 gnd.n1753 gnd.n1734 9.3005
R18850 gnd.n4696 gnd.n1754 9.3005
R18851 gnd.n4695 gnd.n1755 9.3005
R18852 gnd.n4694 gnd.n1756 9.3005
R18853 gnd.n1773 gnd.n1757 9.3005
R18854 gnd.n4684 gnd.n1774 9.3005
R18855 gnd.n4683 gnd.n1775 9.3005
R18856 gnd.n4682 gnd.n1776 9.3005
R18857 gnd.n1793 gnd.n1777 9.3005
R18858 gnd.n4672 gnd.n1794 9.3005
R18859 gnd.n4671 gnd.n1795 9.3005
R18860 gnd.n4670 gnd.n1796 9.3005
R18861 gnd.n1813 gnd.n1797 9.3005
R18862 gnd.n4660 gnd.n1814 9.3005
R18863 gnd.n4659 gnd.n1815 9.3005
R18864 gnd.n4658 gnd.n1816 9.3005
R18865 gnd.n1833 gnd.n1817 9.3005
R18866 gnd.n4648 gnd.n1834 9.3005
R18867 gnd.n4647 gnd.n94 9.3005
R18868 gnd.n99 gnd.n93 9.3005
R18869 gnd.n7865 gnd.n118 9.3005
R18870 gnd.n7864 gnd.n119 9.3005
R18871 gnd.n7863 gnd.n120 9.3005
R18872 gnd.n137 gnd.n121 9.3005
R18873 gnd.n7853 gnd.n138 9.3005
R18874 gnd.n7852 gnd.n139 9.3005
R18875 gnd.n7851 gnd.n140 9.3005
R18876 gnd.n157 gnd.n141 9.3005
R18877 gnd.n7841 gnd.n158 9.3005
R18878 gnd.n7840 gnd.n159 9.3005
R18879 gnd.n7839 gnd.n160 9.3005
R18880 gnd.n177 gnd.n161 9.3005
R18881 gnd.n7829 gnd.n178 9.3005
R18882 gnd.n7828 gnd.n179 9.3005
R18883 gnd.n7827 gnd.n180 9.3005
R18884 gnd.n198 gnd.n181 9.3005
R18885 gnd.n7817 gnd.n199 9.3005
R18886 gnd.n7816 gnd.n200 9.3005
R18887 gnd.n7815 gnd.n201 9.3005
R18888 gnd.n217 gnd.n202 9.3005
R18889 gnd.n7805 gnd.n7804 9.3005
R18890 gnd.n4708 gnd.n1731 9.3005
R18891 gnd.n7876 gnd.n97 9.3005
R18892 gnd.n7876 gnd.n7875 9.3005
R18893 gnd.n3001 gnd.n2984 9.3005
R18894 gnd.n2987 gnd.n2985 9.3005
R18895 gnd.n2997 gnd.n2988 9.3005
R18896 gnd.n2996 gnd.n2989 9.3005
R18897 gnd.n2995 gnd.n2990 9.3005
R18898 gnd.n2993 gnd.n2992 9.3005
R18899 gnd.n2991 gnd.n2628 9.3005
R18900 gnd.n2626 gnd.n2625 9.3005
R18901 gnd.n3072 gnd.n3071 9.3005
R18902 gnd.n3073 gnd.n2624 9.3005
R18903 gnd.n3075 gnd.n3074 9.3005
R18904 gnd.n2622 gnd.n2621 9.3005
R18905 gnd.n3080 gnd.n3079 9.3005
R18906 gnd.n3081 gnd.n2620 9.3005
R18907 gnd.n3115 gnd.n3082 9.3005
R18908 gnd.n3114 gnd.n3083 9.3005
R18909 gnd.n3113 gnd.n3084 9.3005
R18910 gnd.n3087 gnd.n3085 9.3005
R18911 gnd.n3109 gnd.n3088 9.3005
R18912 gnd.n3108 gnd.n3089 9.3005
R18913 gnd.n3107 gnd.n3090 9.3005
R18914 gnd.n3093 gnd.n3091 9.3005
R18915 gnd.n3102 gnd.n3094 9.3005
R18916 gnd.n3101 gnd.n3095 9.3005
R18917 gnd.n3100 gnd.n3096 9.3005
R18918 gnd.n2396 gnd.n2395 9.3005
R18919 gnd.n3226 gnd.n3225 9.3005
R18920 gnd.n3227 gnd.n2394 9.3005
R18921 gnd.n3231 gnd.n3228 9.3005
R18922 gnd.n3230 gnd.n3229 9.3005
R18923 gnd.n2372 gnd.n2371 9.3005
R18924 gnd.n3256 gnd.n3255 9.3005
R18925 gnd.n3257 gnd.n2370 9.3005
R18926 gnd.n3261 gnd.n3258 9.3005
R18927 gnd.n3260 gnd.n3259 9.3005
R18928 gnd.n2347 gnd.n2346 9.3005
R18929 gnd.n3288 gnd.n3287 9.3005
R18930 gnd.n3289 gnd.n2345 9.3005
R18931 gnd.n3297 gnd.n3290 9.3005
R18932 gnd.n3296 gnd.n3291 9.3005
R18933 gnd.n3295 gnd.n3293 9.3005
R18934 gnd.n3292 gnd.n1602 9.3005
R18935 gnd.n4838 gnd.n1603 9.3005
R18936 gnd.n4837 gnd.n1604 9.3005
R18937 gnd.n4836 gnd.n1605 9.3005
R18938 gnd.n2315 gnd.n1606 9.3005
R18939 gnd.n2317 gnd.n2316 9.3005
R18940 gnd.n3455 gnd.n3454 9.3005
R18941 gnd.n3456 gnd.n2314 9.3005
R18942 gnd.n3458 gnd.n3457 9.3005
R18943 gnd.n2294 gnd.n2293 9.3005
R18944 gnd.n3482 gnd.n3481 9.3005
R18945 gnd.n3483 gnd.n2292 9.3005
R18946 gnd.n3487 gnd.n3484 9.3005
R18947 gnd.n3486 gnd.n3485 9.3005
R18948 gnd.n2261 gnd.n2260 9.3005
R18949 gnd.n3524 gnd.n3523 9.3005
R18950 gnd.n3525 gnd.n2259 9.3005
R18951 gnd.n3538 gnd.n3526 9.3005
R18952 gnd.n3537 gnd.n3527 9.3005
R18953 gnd.n3536 gnd.n3528 9.3005
R18954 gnd.n3530 gnd.n3529 9.3005
R18955 gnd.n2227 gnd.n2226 9.3005
R18956 gnd.n3607 gnd.n3606 9.3005
R18957 gnd.n3608 gnd.n2225 9.3005
R18958 gnd.n3610 gnd.n3609 9.3005
R18959 gnd.n2204 gnd.n2203 9.3005
R18960 gnd.n3650 gnd.n3649 9.3005
R18961 gnd.n3651 gnd.n2202 9.3005
R18962 gnd.n3653 gnd.n3652 9.3005
R18963 gnd.n2188 gnd.n2187 9.3005
R18964 gnd.n3694 gnd.n3693 9.3005
R18965 gnd.n3695 gnd.n2186 9.3005
R18966 gnd.n3699 gnd.n3696 9.3005
R18967 gnd.n3698 gnd.n3697 9.3005
R18968 gnd.n2157 gnd.n2156 9.3005
R18969 gnd.n3740 gnd.n3739 9.3005
R18970 gnd.n3741 gnd.n2155 9.3005
R18971 gnd.n3743 gnd.n3742 9.3005
R18972 gnd.n2140 gnd.n2139 9.3005
R18973 gnd.n3801 gnd.n3800 9.3005
R18974 gnd.n3802 gnd.n2138 9.3005
R18975 gnd.n3804 gnd.n3803 9.3005
R18976 gnd.n2118 gnd.n2117 9.3005
R18977 gnd.n3829 gnd.n3828 9.3005
R18978 gnd.n3830 gnd.n2116 9.3005
R18979 gnd.n3834 gnd.n3831 9.3005
R18980 gnd.n3833 gnd.n3832 9.3005
R18981 gnd.n2090 gnd.n2089 9.3005
R18982 gnd.n3873 gnd.n3872 9.3005
R18983 gnd.n3874 gnd.n2088 9.3005
R18984 gnd.n3882 gnd.n3875 9.3005
R18985 gnd.n3881 gnd.n3876 9.3005
R18986 gnd.n3880 gnd.n3878 9.3005
R18987 gnd.n3877 gnd.n2020 9.3005
R18988 gnd.n4147 gnd.n2021 9.3005
R18989 gnd.n4146 gnd.n2022 9.3005
R18990 gnd.n4145 gnd.n2023 9.3005
R18991 gnd.n2030 gnd.n2024 9.3005
R18992 gnd.n4136 gnd.n2031 9.3005
R18993 gnd.n4135 gnd.n2032 9.3005
R18994 gnd.n4134 gnd.n2033 9.3005
R18995 gnd.n2041 gnd.n2034 9.3005
R18996 gnd.n4125 gnd.n2042 9.3005
R18997 gnd.n4124 gnd.n2043 9.3005
R18998 gnd.n4123 gnd.n2044 9.3005
R18999 gnd.n4109 gnd.n2045 9.3005
R19000 gnd.n4114 gnd.n4110 9.3005
R19001 gnd.n4113 gnd.n4112 9.3005
R19002 gnd.n4111 gnd.n1709 9.3005
R19003 gnd.n4723 gnd.n1710 9.3005
R19004 gnd.n4722 gnd.n1711 9.3005
R19005 gnd.n4721 gnd.n1712 9.3005
R19006 gnd.n1718 gnd.n1713 9.3005
R19007 gnd.n4715 gnd.n1719 9.3005
R19008 gnd.n4714 gnd.n1720 9.3005
R19009 gnd.n4713 gnd.n1721 9.3005
R19010 gnd.n1901 gnd.n1722 9.3005
R19011 gnd.n1902 gnd.n1900 9.3005
R19012 gnd.n1904 gnd.n1903 9.3005
R19013 gnd.n1898 gnd.n1897 9.3005
R19014 gnd.n1909 gnd.n1908 9.3005
R19015 gnd.n1910 gnd.n1896 9.3005
R19016 gnd.n1923 gnd.n1911 9.3005
R19017 gnd.n1922 gnd.n1912 9.3005
R19018 gnd.n1921 gnd.n1913 9.3005
R19019 gnd.n1918 gnd.n1914 9.3005
R19020 gnd.n1917 gnd.n1916 9.3005
R19021 gnd.n1915 gnd.n1879 9.3005
R19022 gnd.n1877 gnd.n1876 9.3005
R19023 gnd.n4561 gnd.n4560 9.3005
R19024 gnd.n4562 gnd.n1875 9.3005
R19025 gnd.n4564 gnd.n4563 9.3005
R19026 gnd.n1873 gnd.n1872 9.3005
R19027 gnd.n4569 gnd.n4568 9.3005
R19028 gnd.n4570 gnd.n1871 9.3005
R19029 gnd.n4576 gnd.n4571 9.3005
R19030 gnd.n4575 gnd.n4572 9.3005
R19031 gnd.n7568 gnd.n395 9.3005
R19032 gnd.n398 gnd.n396 9.3005
R19033 gnd.n7564 gnd.n399 9.3005
R19034 gnd.n7563 gnd.n400 9.3005
R19035 gnd.n7562 gnd.n401 9.3005
R19036 gnd.n404 gnd.n402 9.3005
R19037 gnd.n7558 gnd.n405 9.3005
R19038 gnd.n7557 gnd.n406 9.3005
R19039 gnd.n7556 gnd.n407 9.3005
R19040 gnd.n410 gnd.n408 9.3005
R19041 gnd.n7552 gnd.n411 9.3005
R19042 gnd.n7551 gnd.n412 9.3005
R19043 gnd.n7550 gnd.n413 9.3005
R19044 gnd.n416 gnd.n414 9.3005
R19045 gnd.n7546 gnd.n417 9.3005
R19046 gnd.n7545 gnd.n418 9.3005
R19047 gnd.n7544 gnd.n419 9.3005
R19048 gnd.n422 gnd.n420 9.3005
R19049 gnd.n7540 gnd.n423 9.3005
R19050 gnd.n7539 gnd.n424 9.3005
R19051 gnd.n7538 gnd.n425 9.3005
R19052 gnd.n428 gnd.n426 9.3005
R19053 gnd.n7534 gnd.n429 9.3005
R19054 gnd.n7533 gnd.n430 9.3005
R19055 gnd.n7532 gnd.n431 9.3005
R19056 gnd.n2776 gnd.n2717 9.3005
R19057 gnd.n2783 gnd.n2782 9.3005
R19058 gnd.n2784 gnd.n2716 9.3005
R19059 gnd.n2786 gnd.n2785 9.3005
R19060 gnd.n2714 gnd.n2713 9.3005
R19061 gnd.n2841 gnd.n2840 9.3005
R19062 gnd.n2842 gnd.n2712 9.3005
R19063 gnd.n2844 gnd.n2843 9.3005
R19064 gnd.n2710 gnd.n2709 9.3005
R19065 gnd.n2856 gnd.n2855 9.3005
R19066 gnd.n2857 gnd.n2708 9.3005
R19067 gnd.n2860 gnd.n2859 9.3005
R19068 gnd.n2858 gnd.n2702 9.3005
R19069 gnd.n2899 gnd.n2703 9.3005
R19070 gnd.n2898 gnd.n2704 9.3005
R19071 gnd.n2897 gnd.n2705 9.3005
R19072 gnd.n2871 gnd.n2706 9.3005
R19073 gnd.n2887 gnd.n2872 9.3005
R19074 gnd.n2886 gnd.n2873 9.3005
R19075 gnd.n2885 gnd.n2874 9.3005
R19076 gnd.n2879 gnd.n2875 9.3005
R19077 gnd.n2878 gnd.n2876 9.3005
R19078 gnd.n2676 gnd.n2675 9.3005
R19079 gnd.n2948 gnd.n2947 9.3005
R19080 gnd.n2949 gnd.n2674 9.3005
R19081 gnd.n2957 gnd.n2950 9.3005
R19082 gnd.n2775 gnd.n2774 9.3005
R19083 gnd.n2770 gnd.n2769 9.3005
R19084 gnd.n2768 gnd.n2722 9.3005
R19085 gnd.n2767 gnd.n2766 9.3005
R19086 gnd.n2763 gnd.n2725 9.3005
R19087 gnd.n2762 gnd.n2759 9.3005
R19088 gnd.n2758 gnd.n2726 9.3005
R19089 gnd.n2757 gnd.n2756 9.3005
R19090 gnd.n2753 gnd.n2727 9.3005
R19091 gnd.n2752 gnd.n2749 9.3005
R19092 gnd.n2748 gnd.n2728 9.3005
R19093 gnd.n2747 gnd.n2746 9.3005
R19094 gnd.n2743 gnd.n2729 9.3005
R19095 gnd.n2742 gnd.n2739 9.3005
R19096 gnd.n2738 gnd.n2730 9.3005
R19097 gnd.n2737 gnd.n2736 9.3005
R19098 gnd.n2733 gnd.n2731 9.3005
R19099 gnd.n2732 gnd.n1237 9.3005
R19100 gnd.n2771 gnd.n2718 9.3005
R19101 gnd.n2773 gnd.n2772 9.3005
R19102 gnd.n4916 gnd.n1530 9.3005
R19103 gnd.n4917 gnd.n1529 9.3005
R19104 gnd.n1528 gnd.n1525 9.3005
R19105 gnd.n4922 gnd.n1524 9.3005
R19106 gnd.n4923 gnd.n1523 9.3005
R19107 gnd.n4924 gnd.n1522 9.3005
R19108 gnd.n1521 gnd.n1518 9.3005
R19109 gnd.n4929 gnd.n1517 9.3005
R19110 gnd.n4931 gnd.n1514 9.3005
R19111 gnd.n4932 gnd.n1513 9.3005
R19112 gnd.n1512 gnd.n1509 9.3005
R19113 gnd.n4937 gnd.n1508 9.3005
R19114 gnd.n4938 gnd.n1507 9.3005
R19115 gnd.n4939 gnd.n1506 9.3005
R19116 gnd.n1505 gnd.n1502 9.3005
R19117 gnd.n4944 gnd.n1501 9.3005
R19118 gnd.n4945 gnd.n1500 9.3005
R19119 gnd.n4946 gnd.n1499 9.3005
R19120 gnd.n1498 gnd.n1495 9.3005
R19121 gnd.n4951 gnd.n1494 9.3005
R19122 gnd.n4952 gnd.n1493 9.3005
R19123 gnd.n4953 gnd.n1492 9.3005
R19124 gnd.n1491 gnd.n1488 9.3005
R19125 gnd.n1490 gnd.n1486 9.3005
R19126 gnd.n4960 gnd.n1485 9.3005
R19127 gnd.n4962 gnd.n4961 9.3005
R19128 gnd.n2454 gnd.n2453 9.3005
R19129 gnd.n2462 gnd.n2461 9.3005
R19130 gnd.n2463 gnd.n2451 9.3005
R19131 gnd.n2465 gnd.n2464 9.3005
R19132 gnd.n2449 gnd.n2448 9.3005
R19133 gnd.n2472 gnd.n2471 9.3005
R19134 gnd.n2473 gnd.n2447 9.3005
R19135 gnd.n2475 gnd.n2474 9.3005
R19136 gnd.n2445 gnd.n2442 9.3005
R19137 gnd.n2482 gnd.n2481 9.3005
R19138 gnd.n2483 gnd.n2441 9.3005
R19139 gnd.n2485 gnd.n2484 9.3005
R19140 gnd.n2439 gnd.n2438 9.3005
R19141 gnd.n2492 gnd.n2491 9.3005
R19142 gnd.n2493 gnd.n2437 9.3005
R19143 gnd.n2495 gnd.n2494 9.3005
R19144 gnd.n2435 gnd.n2434 9.3005
R19145 gnd.n2502 gnd.n2501 9.3005
R19146 gnd.n2503 gnd.n2433 9.3005
R19147 gnd.n2505 gnd.n2504 9.3005
R19148 gnd.n2431 gnd.n2430 9.3005
R19149 gnd.n2512 gnd.n2511 9.3005
R19150 gnd.n2513 gnd.n2429 9.3005
R19151 gnd.n2515 gnd.n2514 9.3005
R19152 gnd.n2427 gnd.n2426 9.3005
R19153 gnd.n2522 gnd.n2521 9.3005
R19154 gnd.n2523 gnd.n2425 9.3005
R19155 gnd.n2525 gnd.n2524 9.3005
R19156 gnd.n2423 gnd.n2420 9.3005
R19157 gnd.n2531 gnd.n2530 9.3005
R19158 gnd.n2452 gnd.n1531 9.3005
R19159 gnd.n1247 gnd.n1239 9.3005
R19160 gnd.n2777 gnd.n1263 9.3005
R19161 gnd.n5092 gnd.n1264 9.3005
R19162 gnd.n5091 gnd.n1265 9.3005
R19163 gnd.n5090 gnd.n1266 9.3005
R19164 gnd.n2792 gnd.n1267 9.3005
R19165 gnd.n5080 gnd.n1284 9.3005
R19166 gnd.n5079 gnd.n1285 9.3005
R19167 gnd.n5078 gnd.n1286 9.3005
R19168 gnd.n2850 gnd.n1287 9.3005
R19169 gnd.n5068 gnd.n1305 9.3005
R19170 gnd.n5067 gnd.n1306 9.3005
R19171 gnd.n5066 gnd.n1307 9.3005
R19172 gnd.n2866 gnd.n1308 9.3005
R19173 gnd.n5056 gnd.n1325 9.3005
R19174 gnd.n5055 gnd.n1326 9.3005
R19175 gnd.n5054 gnd.n1327 9.3005
R19176 gnd.n2869 gnd.n1328 9.3005
R19177 gnd.n5044 gnd.n1346 9.3005
R19178 gnd.n5043 gnd.n1347 9.3005
R19179 gnd.n5042 gnd.n1348 9.3005
R19180 gnd.n2687 gnd.n1349 9.3005
R19181 gnd.n2932 gnd.n2686 9.3005
R19182 gnd.n2938 gnd.n2685 9.3005
R19183 gnd.n2940 gnd.n2939 9.3005
R19184 gnd.n2671 gnd.n2666 9.3005
R19185 gnd.n2970 gnd.n2667 9.3005
R19186 gnd.n2969 gnd.n2668 9.3005
R19187 gnd.n2968 gnd.n2967 9.3005
R19188 gnd.n2669 gnd.n1374 9.3005
R19189 gnd.n5030 gnd.n1375 9.3005
R19190 gnd.n5029 gnd.n1376 9.3005
R19191 gnd.n5028 gnd.n1377 9.3005
R19192 gnd.n3019 gnd.n1378 9.3005
R19193 gnd.n5018 gnd.n1394 9.3005
R19194 gnd.n5017 gnd.n1395 9.3005
R19195 gnd.n5016 gnd.n1396 9.3005
R19196 gnd.n3034 gnd.n1397 9.3005
R19197 gnd.n5006 gnd.n1414 9.3005
R19198 gnd.n5005 gnd.n1415 9.3005
R19199 gnd.n5004 gnd.n1416 9.3005
R19200 gnd.n3041 gnd.n1417 9.3005
R19201 gnd.n4994 gnd.n1434 9.3005
R19202 gnd.n4993 gnd.n1435 9.3005
R19203 gnd.n4992 gnd.n1436 9.3005
R19204 gnd.n2616 gnd.n1437 9.3005
R19205 gnd.n4982 gnd.n1454 9.3005
R19206 gnd.n4981 gnd.n1455 9.3005
R19207 gnd.n4980 gnd.n1456 9.3005
R19208 gnd.n2611 gnd.n1457 9.3005
R19209 gnd.n4970 gnd.n1475 9.3005
R19210 gnd.n4969 gnd.n1476 9.3005
R19211 gnd.n4968 gnd.n1477 9.3005
R19212 gnd.n5106 gnd.n1238 9.3005
R19213 gnd.n1240 gnd.n1239 9.3005
R19214 gnd.n2778 gnd.n2777 9.3005
R19215 gnd.n2715 gnd.n1264 9.3005
R19216 gnd.n2790 gnd.n1265 9.3005
R19217 gnd.n2791 gnd.n1266 9.3005
R19218 gnd.n2793 gnd.n2792 9.3005
R19219 gnd.n2711 gnd.n1284 9.3005
R19220 gnd.n2848 gnd.n1285 9.3005
R19221 gnd.n2849 gnd.n1286 9.3005
R19222 gnd.n2851 gnd.n2850 9.3005
R19223 gnd.n2707 gnd.n1305 9.3005
R19224 gnd.n2864 gnd.n1306 9.3005
R19225 gnd.n2865 gnd.n1307 9.3005
R19226 gnd.n2867 gnd.n2866 9.3005
R19227 gnd.n2868 gnd.n1325 9.3005
R19228 gnd.n2893 gnd.n1326 9.3005
R19229 gnd.n2892 gnd.n1327 9.3005
R19230 gnd.n2891 gnd.n2869 9.3005
R19231 gnd.n2870 gnd.n1346 9.3005
R19232 gnd.n2881 gnd.n1347 9.3005
R19233 gnd.n2880 gnd.n1348 9.3005
R19234 gnd.n2688 gnd.n2687 9.3005
R19235 gnd.n2936 gnd.n2686 9.3005
R19236 gnd.n2938 gnd.n2937 9.3005
R19237 gnd.n2939 gnd.n2670 9.3005
R19238 gnd.n2961 gnd.n2671 9.3005
R19239 gnd.n2962 gnd.n2667 9.3005
R19240 gnd.n2964 gnd.n2668 9.3005
R19241 gnd.n2967 gnd.n2966 9.3005
R19242 gnd.n2965 gnd.n2669 9.3005
R19243 gnd.n2643 gnd.n1375 9.3005
R19244 gnd.n3017 gnd.n1376 9.3005
R19245 gnd.n3018 gnd.n1377 9.3005
R19246 gnd.n3020 gnd.n3019 9.3005
R19247 gnd.n2638 gnd.n1394 9.3005
R19248 gnd.n3032 gnd.n1395 9.3005
R19249 gnd.n3033 gnd.n1396 9.3005
R19250 gnd.n3035 gnd.n3034 9.3005
R19251 gnd.n3036 gnd.n1414 9.3005
R19252 gnd.n3039 gnd.n1415 9.3005
R19253 gnd.n3040 gnd.n1416 9.3005
R19254 gnd.n3045 gnd.n3041 9.3005
R19255 gnd.n3046 gnd.n1434 9.3005
R19256 gnd.n3047 gnd.n1435 9.3005
R19257 gnd.n2615 gnd.n1436 9.3005
R19258 gnd.n3120 gnd.n2616 9.3005
R19259 gnd.n3121 gnd.n1454 9.3005
R19260 gnd.n3122 gnd.n1455 9.3005
R19261 gnd.n2610 gnd.n1456 9.3005
R19262 gnd.n3135 gnd.n2611 9.3005
R19263 gnd.n3136 gnd.n1475 9.3005
R19264 gnd.n3138 gnd.n1476 9.3005
R19265 gnd.n3137 gnd.n1477 9.3005
R19266 gnd.n5106 gnd.n5105 9.3005
R19267 gnd.n5110 gnd.n5109 9.3005
R19268 gnd.n5113 gnd.n1233 9.3005
R19269 gnd.n5114 gnd.n1232 9.3005
R19270 gnd.n5117 gnd.n1231 9.3005
R19271 gnd.n5118 gnd.n1230 9.3005
R19272 gnd.n5121 gnd.n1229 9.3005
R19273 gnd.n5122 gnd.n1228 9.3005
R19274 gnd.n5125 gnd.n1227 9.3005
R19275 gnd.n5126 gnd.n1226 9.3005
R19276 gnd.n5129 gnd.n1225 9.3005
R19277 gnd.n5130 gnd.n1224 9.3005
R19278 gnd.n5133 gnd.n1223 9.3005
R19279 gnd.n5134 gnd.n1222 9.3005
R19280 gnd.n5137 gnd.n1221 9.3005
R19281 gnd.n5138 gnd.n1220 9.3005
R19282 gnd.n5141 gnd.n1219 9.3005
R19283 gnd.n5142 gnd.n1218 9.3005
R19284 gnd.n5145 gnd.n1217 9.3005
R19285 gnd.n5146 gnd.n1216 9.3005
R19286 gnd.n5149 gnd.n1215 9.3005
R19287 gnd.n5153 gnd.n1211 9.3005
R19288 gnd.n5154 gnd.n1210 9.3005
R19289 gnd.n5157 gnd.n1209 9.3005
R19290 gnd.n5158 gnd.n1208 9.3005
R19291 gnd.n5161 gnd.n1207 9.3005
R19292 gnd.n5162 gnd.n1206 9.3005
R19293 gnd.n5165 gnd.n1205 9.3005
R19294 gnd.n5166 gnd.n1204 9.3005
R19295 gnd.n5169 gnd.n1203 9.3005
R19296 gnd.n5170 gnd.n1202 9.3005
R19297 gnd.n5173 gnd.n1201 9.3005
R19298 gnd.n5174 gnd.n1200 9.3005
R19299 gnd.n5177 gnd.n1199 9.3005
R19300 gnd.n5178 gnd.n1198 9.3005
R19301 gnd.n5181 gnd.n1197 9.3005
R19302 gnd.n5182 gnd.n1196 9.3005
R19303 gnd.n5185 gnd.n1195 9.3005
R19304 gnd.n5186 gnd.n1194 9.3005
R19305 gnd.n5189 gnd.n1193 9.3005
R19306 gnd.n5191 gnd.n1190 9.3005
R19307 gnd.n5194 gnd.n1189 9.3005
R19308 gnd.n5195 gnd.n1188 9.3005
R19309 gnd.n5198 gnd.n1187 9.3005
R19310 gnd.n5199 gnd.n1186 9.3005
R19311 gnd.n5202 gnd.n1185 9.3005
R19312 gnd.n5203 gnd.n1184 9.3005
R19313 gnd.n5206 gnd.n1183 9.3005
R19314 gnd.n5207 gnd.n1182 9.3005
R19315 gnd.n5210 gnd.n1181 9.3005
R19316 gnd.n5211 gnd.n1180 9.3005
R19317 gnd.n5214 gnd.n1179 9.3005
R19318 gnd.n5215 gnd.n1178 9.3005
R19319 gnd.n5218 gnd.n1177 9.3005
R19320 gnd.n5220 gnd.n1176 9.3005
R19321 gnd.n5221 gnd.n1175 9.3005
R19322 gnd.n5222 gnd.n1174 9.3005
R19323 gnd.n5223 gnd.n1173 9.3005
R19324 gnd.n5150 gnd.n1212 9.3005
R19325 gnd.n5108 gnd.n1234 9.3005
R19326 gnd.n5098 gnd.n1253 9.3005
R19327 gnd.n5097 gnd.n1254 9.3005
R19328 gnd.n5096 gnd.n1255 9.3005
R19329 gnd.n1274 gnd.n1256 9.3005
R19330 gnd.n5086 gnd.n1275 9.3005
R19331 gnd.n5085 gnd.n1276 9.3005
R19332 gnd.n5084 gnd.n1277 9.3005
R19333 gnd.n1294 gnd.n1278 9.3005
R19334 gnd.n5074 gnd.n1295 9.3005
R19335 gnd.n5073 gnd.n1296 9.3005
R19336 gnd.n5072 gnd.n1297 9.3005
R19337 gnd.n1315 gnd.n1298 9.3005
R19338 gnd.n5062 gnd.n1316 9.3005
R19339 gnd.n5061 gnd.n1317 9.3005
R19340 gnd.n5060 gnd.n1318 9.3005
R19341 gnd.n1335 gnd.n1319 9.3005
R19342 gnd.n5050 gnd.n1336 9.3005
R19343 gnd.n5049 gnd.n1337 9.3005
R19344 gnd.n5048 gnd.n1338 9.3005
R19345 gnd.n1356 gnd.n1339 9.3005
R19346 gnd.n5038 gnd.n1357 9.3005
R19347 gnd.n1366 gnd.n1359 9.3005
R19348 gnd.n5024 gnd.n1384 9.3005
R19349 gnd.n5023 gnd.n1385 9.3005
R19350 gnd.n5022 gnd.n1386 9.3005
R19351 gnd.n1404 gnd.n1387 9.3005
R19352 gnd.n5012 gnd.n1405 9.3005
R19353 gnd.n5011 gnd.n1406 9.3005
R19354 gnd.n5010 gnd.n1407 9.3005
R19355 gnd.n1423 gnd.n1408 9.3005
R19356 gnd.n5000 gnd.n1424 9.3005
R19357 gnd.n4999 gnd.n1425 9.3005
R19358 gnd.n4998 gnd.n1426 9.3005
R19359 gnd.n1444 gnd.n1427 9.3005
R19360 gnd.n4988 gnd.n1445 9.3005
R19361 gnd.n4987 gnd.n1446 9.3005
R19362 gnd.n4986 gnd.n1447 9.3005
R19363 gnd.n1464 gnd.n1448 9.3005
R19364 gnd.n4976 gnd.n1465 9.3005
R19365 gnd.n4975 gnd.n1466 9.3005
R19366 gnd.n4974 gnd.n1467 9.3005
R19367 gnd.n1484 gnd.n1468 9.3005
R19368 gnd.n4964 gnd.n4963 9.3005
R19369 gnd.n1252 gnd.n1251 9.3005
R19370 gnd.n5035 gnd.n1364 9.3005
R19371 gnd.n5035 gnd.n5034 9.3005
R19372 gnd.n5229 gnd.n1128 9.3005
R19373 gnd.n2802 gnd.n1129 9.3005
R19374 gnd.n2805 gnd.n2804 9.3005
R19375 gnd.n2806 gnd.n2801 9.3005
R19376 gnd.n2808 gnd.n2807 9.3005
R19377 gnd.n2799 gnd.n2798 9.3005
R19378 gnd.n2813 gnd.n2812 9.3005
R19379 gnd.n2814 gnd.n2797 9.3005
R19380 gnd.n2835 gnd.n2815 9.3005
R19381 gnd.n2834 gnd.n2816 9.3005
R19382 gnd.n2833 gnd.n2817 9.3005
R19383 gnd.n2820 gnd.n2818 9.3005
R19384 gnd.n2829 gnd.n2821 9.3005
R19385 gnd.n2828 gnd.n2822 9.3005
R19386 gnd.n2827 gnd.n2823 9.3005
R19387 gnd.n2825 gnd.n2824 9.3005
R19388 gnd.n2699 gnd.n2698 9.3005
R19389 gnd.n2906 gnd.n2905 9.3005
R19390 gnd.n2907 gnd.n2697 9.3005
R19391 gnd.n2909 gnd.n2908 9.3005
R19392 gnd.n2695 gnd.n2694 9.3005
R19393 gnd.n2915 gnd.n2914 9.3005
R19394 gnd.n2916 gnd.n2693 9.3005
R19395 gnd.n2918 gnd.n2917 9.3005
R19396 gnd.n5231 gnd.n5230 9.3005
R19397 gnd.n1127 gnd.n1037 9.3005
R19398 gnd.n6632 gnd.n1036 9.3005
R19399 gnd.n6633 gnd.n1035 9.3005
R19400 gnd.n6634 gnd.n1034 9.3005
R19401 gnd.n1033 gnd.n1029 9.3005
R19402 gnd.n6640 gnd.n1028 9.3005
R19403 gnd.n6641 gnd.n1027 9.3005
R19404 gnd.n6642 gnd.n1026 9.3005
R19405 gnd.n1025 gnd.n1021 9.3005
R19406 gnd.n6648 gnd.n1020 9.3005
R19407 gnd.n6649 gnd.n1019 9.3005
R19408 gnd.n6650 gnd.n1018 9.3005
R19409 gnd.n1017 gnd.n1013 9.3005
R19410 gnd.n6656 gnd.n1012 9.3005
R19411 gnd.n6657 gnd.n1011 9.3005
R19412 gnd.n6658 gnd.n1010 9.3005
R19413 gnd.n1009 gnd.n1005 9.3005
R19414 gnd.n6664 gnd.n1004 9.3005
R19415 gnd.n6665 gnd.n1003 9.3005
R19416 gnd.n6666 gnd.n1002 9.3005
R19417 gnd.n1001 gnd.n997 9.3005
R19418 gnd.n6672 gnd.n996 9.3005
R19419 gnd.n6673 gnd.n995 9.3005
R19420 gnd.n6674 gnd.n994 9.3005
R19421 gnd.n993 gnd.n989 9.3005
R19422 gnd.n6680 gnd.n988 9.3005
R19423 gnd.n6681 gnd.n987 9.3005
R19424 gnd.n6682 gnd.n986 9.3005
R19425 gnd.n985 gnd.n981 9.3005
R19426 gnd.n6688 gnd.n980 9.3005
R19427 gnd.n6689 gnd.n979 9.3005
R19428 gnd.n6690 gnd.n978 9.3005
R19429 gnd.n977 gnd.n973 9.3005
R19430 gnd.n6696 gnd.n972 9.3005
R19431 gnd.n6697 gnd.n971 9.3005
R19432 gnd.n6698 gnd.n970 9.3005
R19433 gnd.n969 gnd.n965 9.3005
R19434 gnd.n6704 gnd.n964 9.3005
R19435 gnd.n6705 gnd.n963 9.3005
R19436 gnd.n6706 gnd.n962 9.3005
R19437 gnd.n961 gnd.n957 9.3005
R19438 gnd.n6712 gnd.n956 9.3005
R19439 gnd.n6713 gnd.n955 9.3005
R19440 gnd.n6714 gnd.n954 9.3005
R19441 gnd.n953 gnd.n949 9.3005
R19442 gnd.n6720 gnd.n948 9.3005
R19443 gnd.n6721 gnd.n947 9.3005
R19444 gnd.n6722 gnd.n946 9.3005
R19445 gnd.n945 gnd.n941 9.3005
R19446 gnd.n6728 gnd.n940 9.3005
R19447 gnd.n6729 gnd.n939 9.3005
R19448 gnd.n6730 gnd.n938 9.3005
R19449 gnd.n937 gnd.n933 9.3005
R19450 gnd.n6736 gnd.n932 9.3005
R19451 gnd.n6737 gnd.n931 9.3005
R19452 gnd.n6738 gnd.n930 9.3005
R19453 gnd.n929 gnd.n925 9.3005
R19454 gnd.n6744 gnd.n924 9.3005
R19455 gnd.n6745 gnd.n923 9.3005
R19456 gnd.n6746 gnd.n922 9.3005
R19457 gnd.n921 gnd.n917 9.3005
R19458 gnd.n6752 gnd.n916 9.3005
R19459 gnd.n6753 gnd.n915 9.3005
R19460 gnd.n6754 gnd.n914 9.3005
R19461 gnd.n913 gnd.n909 9.3005
R19462 gnd.n6760 gnd.n908 9.3005
R19463 gnd.n6761 gnd.n907 9.3005
R19464 gnd.n6762 gnd.n906 9.3005
R19465 gnd.n905 gnd.n901 9.3005
R19466 gnd.n6768 gnd.n900 9.3005
R19467 gnd.n6769 gnd.n899 9.3005
R19468 gnd.n6770 gnd.n898 9.3005
R19469 gnd.n897 gnd.n893 9.3005
R19470 gnd.n6776 gnd.n892 9.3005
R19471 gnd.n6777 gnd.n891 9.3005
R19472 gnd.n6778 gnd.n890 9.3005
R19473 gnd.n889 gnd.n885 9.3005
R19474 gnd.n6784 gnd.n884 9.3005
R19475 gnd.n6785 gnd.n883 9.3005
R19476 gnd.n6786 gnd.n882 9.3005
R19477 gnd.n881 gnd.n877 9.3005
R19478 gnd.n6792 gnd.n876 9.3005
R19479 gnd.n6793 gnd.n875 9.3005
R19480 gnd.n6794 gnd.n874 9.3005
R19481 gnd.n5233 gnd.n5232 9.3005
R19482 gnd.n4101 gnd.n4100 9.3005
R19483 gnd.n2379 gnd.n2378 9.3005
R19484 gnd.n3246 gnd.n3245 9.3005
R19485 gnd.n3247 gnd.n2376 9.3005
R19486 gnd.n3250 gnd.n3249 9.3005
R19487 gnd.n3248 gnd.n2377 9.3005
R19488 gnd.n2354 gnd.n2353 9.3005
R19489 gnd.n3276 gnd.n3275 9.3005
R19490 gnd.n3277 gnd.n2351 9.3005
R19491 gnd.n3282 gnd.n3281 9.3005
R19492 gnd.n3280 gnd.n2352 9.3005
R19493 gnd.n3279 gnd.n3278 9.3005
R19494 gnd.n2330 gnd.n2329 9.3005
R19495 gnd.n3322 gnd.n3321 9.3005
R19496 gnd.n3323 gnd.n2328 9.3005
R19497 gnd.n3325 gnd.n3324 9.3005
R19498 gnd.n2326 gnd.n2325 9.3005
R19499 gnd.n3413 gnd.n3412 9.3005
R19500 gnd.n3414 gnd.n2323 9.3005
R19501 gnd.n3417 gnd.n3416 9.3005
R19502 gnd.n3415 gnd.n2324 9.3005
R19503 gnd.n2301 gnd.n2300 9.3005
R19504 gnd.n3473 gnd.n3472 9.3005
R19505 gnd.n3474 gnd.n2299 9.3005
R19506 gnd.n3476 gnd.n3475 9.3005
R19507 gnd.n2280 gnd.n2279 9.3005
R19508 gnd.n3502 gnd.n3501 9.3005
R19509 gnd.n3503 gnd.n2277 9.3005
R19510 gnd.n3509 gnd.n3508 9.3005
R19511 gnd.n3507 gnd.n2278 9.3005
R19512 gnd.n3506 gnd.n3505 9.3005
R19513 gnd.n2245 gnd.n2244 9.3005
R19514 gnd.n3562 gnd.n3561 9.3005
R19515 gnd.n3563 gnd.n2242 9.3005
R19516 gnd.n3566 gnd.n3565 9.3005
R19517 gnd.n3564 gnd.n2243 9.3005
R19518 gnd.n2220 gnd.n2219 9.3005
R19519 gnd.n3616 gnd.n3615 9.3005
R19520 gnd.n3617 gnd.n2217 9.3005
R19521 gnd.n3631 gnd.n3630 9.3005
R19522 gnd.n3629 gnd.n2218 9.3005
R19523 gnd.n3628 gnd.n3627 9.3005
R19524 gnd.n3626 gnd.n3618 9.3005
R19525 gnd.n3625 gnd.n3624 9.3005
R19526 gnd.n3623 gnd.n3622 9.3005
R19527 gnd.n2174 gnd.n2173 9.3005
R19528 gnd.n3712 gnd.n3711 9.3005
R19529 gnd.n3713 gnd.n2171 9.3005
R19530 gnd.n3725 gnd.n3724 9.3005
R19531 gnd.n3723 gnd.n2172 9.3005
R19532 gnd.n3722 gnd.n3721 9.3005
R19533 gnd.n3720 gnd.n3714 9.3005
R19534 gnd.n3719 gnd.n3718 9.3005
R19535 gnd.n2134 gnd.n2133 9.3005
R19536 gnd.n3810 gnd.n3809 9.3005
R19537 gnd.n3811 gnd.n2131 9.3005
R19538 gnd.n3814 gnd.n3813 9.3005
R19539 gnd.n3812 gnd.n2132 9.3005
R19540 gnd.n2105 gnd.n2104 9.3005
R19541 gnd.n3848 gnd.n3847 9.3005
R19542 gnd.n3849 gnd.n2102 9.3005
R19543 gnd.n3859 gnd.n3858 9.3005
R19544 gnd.n3857 gnd.n2103 9.3005
R19545 gnd.n3856 gnd.n3855 9.3005
R19546 gnd.n3854 gnd.n3851 9.3005
R19547 gnd.n3850 gnd.n2069 9.3005
R19548 gnd.n3902 gnd.n2068 9.3005
R19549 gnd.n3904 gnd.n3903 9.3005
R19550 gnd.n3905 gnd.n2065 9.3005
R19551 gnd.n3907 gnd.n3906 9.3005
R19552 gnd.n3908 gnd.n2064 9.3005
R19553 gnd.n3910 gnd.n3909 9.3005
R19554 gnd.n3911 gnd.n2061 9.3005
R19555 gnd.n3913 gnd.n3912 9.3005
R19556 gnd.n3914 gnd.n2060 9.3005
R19557 gnd.n3916 gnd.n3915 9.3005
R19558 gnd.n3917 gnd.n2055 9.3005
R19559 gnd.n3919 gnd.n3918 9.3005
R19560 gnd.n3920 gnd.n2054 9.3005
R19561 gnd.n3922 gnd.n3921 9.3005
R19562 gnd.n3923 gnd.n2052 9.3005
R19563 gnd.n4104 gnd.n4103 9.3005
R19564 gnd.n4102 gnd.n2053 9.3005
R19565 gnd.n3153 gnd.n3152 9.3005
R19566 gnd.n3155 gnd.n3154 9.3005
R19567 gnd.n2956 gnd.n2955 9.3005
R19568 gnd.n2954 gnd.n2952 9.3005
R19569 gnd.n2646 gnd.n2645 9.3005
R19570 gnd.n3010 gnd.n3009 9.3005
R19571 gnd.n3011 gnd.n2644 9.3005
R19572 gnd.n3013 gnd.n3012 9.3005
R19573 gnd.n2641 gnd.n2640 9.3005
R19574 gnd.n3025 gnd.n3024 9.3005
R19575 gnd.n3026 gnd.n2639 9.3005
R19576 gnd.n3028 gnd.n3027 9.3005
R19577 gnd.n2632 gnd.n2630 9.3005
R19578 gnd.n3064 gnd.n3063 9.3005
R19579 gnd.n3062 gnd.n2631 9.3005
R19580 gnd.n3061 gnd.n3060 9.3005
R19581 gnd.n3059 gnd.n2633 9.3005
R19582 gnd.n3058 gnd.n3057 9.3005
R19583 gnd.n3056 gnd.n2636 9.3005
R19584 gnd.n3055 gnd.n3054 9.3005
R19585 gnd.n3053 gnd.n2637 9.3005
R19586 gnd.n3052 gnd.n3051 9.3005
R19587 gnd.n2614 gnd.n2613 9.3005
R19588 gnd.n3127 gnd.n3126 9.3005
R19589 gnd.n3128 gnd.n2612 9.3005
R19590 gnd.n3131 gnd.n3130 9.3005
R19591 gnd.n3129 gnd.n2609 9.3005
R19592 gnd.n3142 gnd.n2608 9.3005
R19593 gnd.n3144 gnd.n3143 9.3005
R19594 gnd.n3204 gnd.n3203 9.3005
R19595 gnd.n3202 gnd.n3201 9.3005
R19596 gnd.n2546 gnd.n2545 9.3005
R19597 gnd.n3196 gnd.n3195 9.3005
R19598 gnd.n3194 gnd.n3193 9.3005
R19599 gnd.n2558 gnd.n2557 9.3005
R19600 gnd.n3188 gnd.n3187 9.3005
R19601 gnd.n3186 gnd.n3185 9.3005
R19602 gnd.n2569 gnd.n2568 9.3005
R19603 gnd.n3180 gnd.n3179 9.3005
R19604 gnd.n3178 gnd.n3177 9.3005
R19605 gnd.n2581 gnd.n2580 9.3005
R19606 gnd.n3172 gnd.n3171 9.3005
R19607 gnd.n3170 gnd.n3169 9.3005
R19608 gnd.n2592 gnd.n2591 9.3005
R19609 gnd.n3164 gnd.n3163 9.3005
R19610 gnd.n3162 gnd.n2605 9.3005
R19611 gnd.n3161 gnd.n3158 9.3005
R19612 gnd.n2541 gnd.n2539 9.3005
R19613 gnd.n3157 gnd.n3156 9.3005
R19614 gnd.n3148 gnd.n2607 9.3005
R19615 gnd.n3147 gnd.n2599 9.3005
R19616 gnd.n3166 gnd.n3165 9.3005
R19617 gnd.n3168 gnd.n3167 9.3005
R19618 gnd.n2585 gnd.n2584 9.3005
R19619 gnd.n3174 gnd.n3173 9.3005
R19620 gnd.n3176 gnd.n3175 9.3005
R19621 gnd.n2575 gnd.n2574 9.3005
R19622 gnd.n3182 gnd.n3181 9.3005
R19623 gnd.n3184 gnd.n3183 9.3005
R19624 gnd.n2562 gnd.n2561 9.3005
R19625 gnd.n3190 gnd.n3189 9.3005
R19626 gnd.n3192 gnd.n3191 9.3005
R19627 gnd.n2552 gnd.n2551 9.3005
R19628 gnd.n3198 gnd.n3197 9.3005
R19629 gnd.n3200 gnd.n3199 9.3005
R19630 gnd.n2540 gnd.n2538 9.3005
R19631 gnd.n3206 gnd.n3205 9.3005
R19632 gnd.n3207 gnd.n2533 9.3005
R19633 gnd.n3209 gnd.n3208 9.3005
R19634 gnd.n3211 gnd.n2419 9.3005
R19635 gnd.n3213 gnd.n3212 9.3005
R19636 gnd.n3214 gnd.n2415 9.3005
R19637 gnd.n3216 gnd.n3215 9.3005
R19638 gnd.n3217 gnd.n2414 9.3005
R19639 gnd.n3219 gnd.n3218 9.3005
R19640 gnd.n2413 gnd.n2386 9.3005
R19641 gnd.n3238 gnd.n2384 9.3005
R19642 gnd.n3241 gnd.n3240 9.3005
R19643 gnd.n3239 gnd.n2385 9.3005
R19644 gnd.n2363 gnd.n2362 9.3005
R19645 gnd.n3267 gnd.n3266 9.3005
R19646 gnd.n3268 gnd.n2360 9.3005
R19647 gnd.n3271 gnd.n3270 9.3005
R19648 gnd.n3269 gnd.n2361 9.3005
R19649 gnd.n2338 gnd.n2337 9.3005
R19650 gnd.n3303 gnd.n3302 9.3005
R19651 gnd.n3304 gnd.n2335 9.3005
R19652 gnd.n3316 gnd.n3315 9.3005
R19653 gnd.n3314 gnd.n2336 9.3005
R19654 gnd.n3313 gnd.n3312 9.3005
R19655 gnd.n3311 gnd.n3305 9.3005
R19656 gnd.n3310 gnd.n3309 9.3005
R19657 gnd.n1623 gnd.n1621 9.3005
R19658 gnd.n4824 gnd.n4823 9.3005
R19659 gnd.n4822 gnd.n1622 9.3005
R19660 gnd.n4821 gnd.n4820 9.3005
R19661 gnd.n4819 gnd.n1624 9.3005
R19662 gnd.n4818 gnd.n4817 9.3005
R19663 gnd.n4816 gnd.n1628 9.3005
R19664 gnd.n4815 gnd.n4814 9.3005
R19665 gnd.n4813 gnd.n1629 9.3005
R19666 gnd.n4812 gnd.n4811 9.3005
R19667 gnd.n4810 gnd.n1633 9.3005
R19668 gnd.n4809 gnd.n4808 9.3005
R19669 gnd.n4807 gnd.n1634 9.3005
R19670 gnd.n4806 gnd.n4805 9.3005
R19671 gnd.n4804 gnd.n1638 9.3005
R19672 gnd.n4803 gnd.n4802 9.3005
R19673 gnd.n4801 gnd.n1639 9.3005
R19674 gnd.n4800 gnd.n4799 9.3005
R19675 gnd.n4798 gnd.n1643 9.3005
R19676 gnd.n4797 gnd.n4796 9.3005
R19677 gnd.n4795 gnd.n1644 9.3005
R19678 gnd.n4794 gnd.n4793 9.3005
R19679 gnd.n4792 gnd.n1648 9.3005
R19680 gnd.n4791 gnd.n4790 9.3005
R19681 gnd.n4789 gnd.n1649 9.3005
R19682 gnd.n4788 gnd.n4787 9.3005
R19683 gnd.n4786 gnd.n1653 9.3005
R19684 gnd.n4785 gnd.n4784 9.3005
R19685 gnd.n4783 gnd.n1654 9.3005
R19686 gnd.n4782 gnd.n4781 9.3005
R19687 gnd.n4780 gnd.n1658 9.3005
R19688 gnd.n4779 gnd.n4778 9.3005
R19689 gnd.n4777 gnd.n1659 9.3005
R19690 gnd.n4776 gnd.n4775 9.3005
R19691 gnd.n4774 gnd.n1663 9.3005
R19692 gnd.n4773 gnd.n4772 9.3005
R19693 gnd.n4771 gnd.n1664 9.3005
R19694 gnd.n4770 gnd.n4769 9.3005
R19695 gnd.n4768 gnd.n1668 9.3005
R19696 gnd.n4767 gnd.n4766 9.3005
R19697 gnd.n4765 gnd.n1669 9.3005
R19698 gnd.n4764 gnd.n4763 9.3005
R19699 gnd.n4762 gnd.n1673 9.3005
R19700 gnd.n4761 gnd.n4760 9.3005
R19701 gnd.n4759 gnd.n1674 9.3005
R19702 gnd.n4758 gnd.n4757 9.3005
R19703 gnd.n4756 gnd.n1678 9.3005
R19704 gnd.n4755 gnd.n4754 9.3005
R19705 gnd.n4753 gnd.n1679 9.3005
R19706 gnd.n4752 gnd.n4751 9.3005
R19707 gnd.n4750 gnd.n1683 9.3005
R19708 gnd.n4749 gnd.n4748 9.3005
R19709 gnd.n4747 gnd.n1684 9.3005
R19710 gnd.n4746 gnd.n4745 9.3005
R19711 gnd.n4744 gnd.n1688 9.3005
R19712 gnd.n4743 gnd.n4742 9.3005
R19713 gnd.n4741 gnd.n1689 9.3005
R19714 gnd.n4740 gnd.n4739 9.3005
R19715 gnd.n4738 gnd.n1693 9.3005
R19716 gnd.n4737 gnd.n4736 9.3005
R19717 gnd.n4735 gnd.n1694 9.3005
R19718 gnd.n4734 gnd.n4733 9.3005
R19719 gnd.n4732 gnd.n1698 9.3005
R19720 gnd.n4731 gnd.n4730 9.3005
R19721 gnd.n4729 gnd.n1699 9.3005
R19722 gnd.n4728 gnd.n1702 9.3005
R19723 gnd.n3237 gnd.n3236 9.3005
R19724 gnd.n3990 gnd.n3989 9.3005
R19725 gnd.n3985 gnd.n3984 9.3005
R19726 gnd.n3997 gnd.n3996 9.3005
R19727 gnd.n3998 gnd.n3983 9.3005
R19728 gnd.n4001 gnd.n4000 9.3005
R19729 gnd.n3999 gnd.n3981 9.3005
R19730 gnd.n3988 gnd.n3987 9.3005
R19731 gnd.n4089 gnd.n3937 9.3005
R19732 gnd.n3950 gnd.n3946 9.3005
R19733 gnd.n4083 gnd.n4082 9.3005
R19734 gnd.n4071 gnd.n3948 9.3005
R19735 gnd.n4070 gnd.n4069 9.3005
R19736 gnd.n3959 gnd.n3955 9.3005
R19737 gnd.n4063 gnd.n4062 9.3005
R19738 gnd.n4052 gnd.n3957 9.3005
R19739 gnd.n4051 gnd.n4050 9.3005
R19740 gnd.n3968 gnd.n3964 9.3005
R19741 gnd.n4044 gnd.n4043 9.3005
R19742 gnd.n4033 gnd.n3966 9.3005
R19743 gnd.n4032 gnd.n4031 9.3005
R19744 gnd.n3977 gnd.n3973 9.3005
R19745 gnd.n4025 gnd.n4024 9.3005
R19746 gnd.n4014 gnd.n3975 9.3005
R19747 gnd.n4013 gnd.n4012 9.3005
R19748 gnd.n4091 gnd.n4090 9.3005
R19749 gnd.n3941 gnd.n3940 9.3005
R19750 gnd.n4008 gnd.n4007 9.3005
R19751 gnd.n4009 gnd.n3980 9.3005
R19752 gnd.n4016 gnd.n4015 9.3005
R19753 gnd.n3978 gnd.n3976 9.3005
R19754 gnd.n4023 gnd.n4022 9.3005
R19755 gnd.n3972 gnd.n3971 9.3005
R19756 gnd.n4035 gnd.n4034 9.3005
R19757 gnd.n3969 gnd.n3967 9.3005
R19758 gnd.n4042 gnd.n4041 9.3005
R19759 gnd.n3963 gnd.n3962 9.3005
R19760 gnd.n4054 gnd.n4053 9.3005
R19761 gnd.n3960 gnd.n3958 9.3005
R19762 gnd.n4061 gnd.n4060 9.3005
R19763 gnd.n3954 gnd.n3953 9.3005
R19764 gnd.n4073 gnd.n4072 9.3005
R19765 gnd.n3951 gnd.n3949 9.3005
R19766 gnd.n4081 gnd.n4080 9.3005
R19767 gnd.n4079 gnd.n4078 9.3005
R19768 gnd.n4093 gnd.n4092 9.3005
R19769 gnd.n3938 gnd.n3932 9.3005
R19770 gnd.n3939 gnd.n3931 9.3005
R19771 gnd.n3927 gnd.n3924 9.3005
R19772 gnd.n1930 gnd.n1929 9.3005
R19773 gnd.n4500 gnd.n4499 9.3005
R19774 gnd.n4501 gnd.n1928 9.3005
R19775 gnd.n4503 gnd.n4502 9.3005
R19776 gnd.n1893 gnd.n1892 9.3005
R19777 gnd.n4514 gnd.n4513 9.3005
R19778 gnd.n4515 gnd.n1891 9.3005
R19779 gnd.n4517 gnd.n4516 9.3005
R19780 gnd.n1883 gnd.n1881 9.3005
R19781 gnd.n4553 gnd.n4552 9.3005
R19782 gnd.n4551 gnd.n1882 9.3005
R19783 gnd.n4550 gnd.n4549 9.3005
R19784 gnd.n4548 gnd.n1884 9.3005
R19785 gnd.n4547 gnd.n4546 9.3005
R19786 gnd.n4545 gnd.n1887 9.3005
R19787 gnd.n4544 gnd.n4543 9.3005
R19788 gnd.n4542 gnd.n1888 9.3005
R19789 gnd.n4541 gnd.n4540 9.3005
R19790 gnd.n1866 gnd.n1865 9.3005
R19791 gnd.n4612 gnd.n4611 9.3005
R19792 gnd.n4613 gnd.n1863 9.3005
R19793 gnd.n4618 gnd.n4617 9.3005
R19794 gnd.n4616 gnd.n1864 9.3005
R19795 gnd.n4615 gnd.n4614 9.3005
R19796 gnd.n81 gnd.n79 9.3005
R19797 gnd.n3929 gnd.n3928 9.3005
R19798 gnd.t326 gnd.n5354 9.24152
R19799 gnd.n6586 gnd.t6 9.24152
R19800 gnd.t104 gnd.n1114 9.24152
R19801 gnd.n2780 gnd.t24 9.24152
R19802 gnd.n3117 gnd.t158 9.24152
R19803 gnd.n3870 gnd.t322 9.24152
R19804 gnd.n1925 gnd.t167 9.24152
R19805 gnd.n7813 gnd.t28 9.24152
R19806 gnd.t348 gnd.t326 8.92286
R19807 gnd.n3461 gnd.n2311 8.92286
R19808 gnd.n3429 gnd.n2273 8.92286
R19809 gnd.n3540 gnd.t136 8.92286
R19810 gnd.n3558 gnd.t314 8.92286
R19811 gnd.n3637 gnd.n2212 8.92286
R19812 gnd.n3690 gnd.n2191 8.92286
R19813 gnd.n2164 gnd.t305 8.92286
R19814 gnd.t309 gnd.n3787 8.92286
R19815 gnd.n3819 gnd.n2126 8.92286
R19816 gnd.n3862 gnd.n3861 8.92286
R19817 gnd.n6440 gnd.n6415 8.92171
R19818 gnd.n6408 gnd.n6383 8.92171
R19819 gnd.n6376 gnd.n6351 8.92171
R19820 gnd.n6345 gnd.n6320 8.92171
R19821 gnd.n6313 gnd.n6288 8.92171
R19822 gnd.n6281 gnd.n6256 8.92171
R19823 gnd.n6249 gnd.n6224 8.92171
R19824 gnd.n6218 gnd.n6193 8.92171
R19825 gnd.n4174 gnd.n4156 8.72777
R19826 gnd.n6014 gnd.t132 8.60421
R19827 gnd.t124 gnd.n3635 8.60421
R19828 gnd.n3680 gnd.t312 8.60421
R19829 gnd.n5426 gnd.n5410 8.43656
R19830 gnd.n46 gnd.n30 8.43656
R19831 gnd.n3452 gnd.n2319 8.28555
R19832 gnd.n3521 gnd.n3520 8.28555
R19833 gnd.n3586 gnd.n3585 8.28555
R19834 gnd.n3701 gnd.n2176 8.28555
R19835 gnd.n3780 gnd.n3779 8.28555
R19836 gnd.n3752 gnd.n2095 8.28555
R19837 gnd.n6441 gnd.n6413 8.14595
R19838 gnd.n6409 gnd.n6381 8.14595
R19839 gnd.n6377 gnd.n6349 8.14595
R19840 gnd.n6346 gnd.n6318 8.14595
R19841 gnd.n6314 gnd.n6286 8.14595
R19842 gnd.n6282 gnd.n6254 8.14595
R19843 gnd.n6250 gnd.n6222 8.14595
R19844 gnd.n6219 gnd.n6191 8.14595
R19845 gnd.n2953 gnd.n0 8.10675
R19846 gnd.n7887 gnd.n7886 8.10675
R19847 gnd.n6446 gnd.n6445 7.97301
R19848 gnd.t130 gnd.n5529 7.9669
R19849 gnd.n3402 gnd.t126 7.9669
R19850 gnd.t60 gnd.t333 7.9669
R19851 gnd.n7887 gnd.n78 7.86902
R19852 gnd.n4090 gnd.n3941 7.75808
R19853 gnd.n3162 gnd.n3161 7.75808
R19854 gnd.n7663 gnd.n353 7.75808
R19855 gnd.n2772 gnd.n2771 7.75808
R19856 gnd.n3419 gnd.n2319 7.64824
R19857 gnd.n3520 gnd.n2265 7.64824
R19858 gnd.n3584 gnd.t128 7.64824
R19859 gnd.n3586 gnd.n3584 7.64824
R19860 gnd.n3709 gnd.n2176 7.64824
R19861 gnd.n3709 gnd.t306 7.64824
R19862 gnd.n3780 gnd.n3778 7.64824
R19863 gnd.n5459 gnd.n5458 7.53171
R19864 gnd.n5923 gnd.t2 7.32958
R19865 gnd.n1593 gnd.n1592 7.30353
R19866 gnd.n4173 gnd.n4172 7.30353
R19867 gnd.n5883 gnd.n5602 7.01093
R19868 gnd.n5605 gnd.n5603 7.01093
R19869 gnd.n5893 gnd.n5892 7.01093
R19870 gnd.n5904 gnd.n5586 7.01093
R19871 gnd.n5903 gnd.n5589 7.01093
R19872 gnd.n5914 gnd.n5577 7.01093
R19873 gnd.n5580 gnd.n5578 7.01093
R19874 gnd.n5924 gnd.n5923 7.01093
R19875 gnd.n5934 gnd.n5558 7.01093
R19876 gnd.n5933 gnd.n5561 7.01093
R19877 gnd.n5942 gnd.n5552 7.01093
R19878 gnd.n5954 gnd.n5542 7.01093
R19879 gnd.n5964 gnd.n5527 7.01093
R19880 gnd.n5980 gnd.n5979 7.01093
R19881 gnd.n5529 gnd.n5466 7.01093
R19882 gnd.n6034 gnd.n5467 7.01093
R19883 gnd.n6028 gnd.n6027 7.01093
R19884 gnd.n5516 gnd.n5478 7.01093
R19885 gnd.n6020 gnd.n5489 7.01093
R19886 gnd.n5507 gnd.n5502 7.01093
R19887 gnd.n6014 gnd.n6013 7.01093
R19888 gnd.n6060 gnd.n5389 7.01093
R19889 gnd.n6059 gnd.n6058 7.01093
R19890 gnd.n6071 gnd.n6070 7.01093
R19891 gnd.n5382 gnd.n5374 7.01093
R19892 gnd.n6100 gnd.n5362 7.01093
R19893 gnd.n6099 gnd.n5365 7.01093
R19894 gnd.n6110 gnd.n5354 7.01093
R19895 gnd.n5355 gnd.n5343 7.01093
R19896 gnd.n6123 gnd.n5344 7.01093
R19897 gnd.n6156 gnd.n5336 7.01093
R19898 gnd.n6155 gnd.n1039 7.01093
R19899 gnd.n6621 gnd.n6620 7.01093
R19900 gnd.n6146 gnd.n6145 7.01093
R19901 gnd.n6614 gnd.n1060 7.01093
R19902 gnd.n6613 gnd.n1063 7.01093
R19903 gnd.n6138 gnd.n1072 7.01093
R19904 gnd.n6607 gnd.n6606 7.01093
R19905 gnd.n6600 gnd.n1085 7.01093
R19906 gnd.n6599 gnd.n1088 7.01093
R19907 gnd.n6478 gnd.n1097 7.01093
R19908 gnd.n6593 gnd.n6592 7.01093
R19909 gnd.n6459 gnd.n1100 7.01093
R19910 gnd.n6586 gnd.n1111 7.01093
R19911 gnd.n6585 gnd.n1114 7.01093
R19912 gnd.n6489 gnd.n1122 7.01093
R19913 gnd.n6579 gnd.n6578 7.01093
R19914 gnd.n3444 gnd.t336 7.01093
R19915 gnd.n3461 gnd.n3460 7.01093
R19916 gnd.n3429 gnd.n2283 7.01093
R19917 gnd.n3637 gnd.n3636 7.01093
R19918 gnd.n3691 gnd.n3690 7.01093
R19919 gnd.n3819 gnd.n3818 7.01093
R19920 gnd.n3862 gnd.n2099 7.01093
R19921 gnd.t135 gnd.n2092 7.01093
R19922 gnd.n5561 gnd.t302 6.69227
R19923 gnd.n5365 gnd.t348 6.69227
R19924 gnd.n6628 gnd.n1039 6.69227
R19925 gnd.t303 gnd.n6470 6.69227
R19926 gnd.n3049 gnd.t172 6.69227
R19927 gnd.n3446 gnd.t315 6.69227
R19928 gnd.t322 gnd.n3869 6.69227
R19929 gnd.n4519 gnd.t137 6.69227
R19930 gnd.n4303 gnd.n4302 6.5566
R19931 gnd.n3334 gnd.n3333 6.5566
R19932 gnd.n4852 gnd.n4848 6.5566
R19933 gnd.n4181 gnd.n4180 6.5566
R19934 gnd.n3394 gnd.n1597 6.37362
R19935 gnd.n3410 gnd.n3409 6.37362
R19936 gnd.t98 gnd.n3445 6.37362
R19937 gnd.n3499 gnd.t327 6.37362
R19938 gnd.n3551 gnd.n3550 6.37362
R19939 gnd.n3603 gnd.t128 6.37362
R19940 gnd.t306 gnd.n3708 6.37362
R19941 gnd.n3788 gnd.n2149 6.37362
R19942 gnd.n3816 gnd.t329 6.37362
R19943 gnd.n3892 gnd.n2075 6.37362
R19944 gnd.n4242 gnd.n2008 6.37362
R19945 gnd.n3147 gnd.n2598 6.20656
R19946 gnd.n4093 gnd.n3936 6.20656
R19947 gnd.t339 gnd.n5990 6.05496
R19948 gnd.n5991 gnd.t1 6.05496
R19949 gnd.t359 gnd.n5389 6.05496
R19950 gnd.n6165 gnd.t0 6.05496
R19951 gnd.n3030 gnd.t165 6.05496
R19952 gnd.n3636 gnd.t124 6.05496
R19953 gnd.n3691 gnd.t312 6.05496
R19954 gnd.n4538 gnd.t147 6.05496
R19955 gnd.n6443 gnd.n6413 5.81868
R19956 gnd.n6411 gnd.n6381 5.81868
R19957 gnd.n6379 gnd.n6349 5.81868
R19958 gnd.n6348 gnd.n6318 5.81868
R19959 gnd.n6316 gnd.n6286 5.81868
R19960 gnd.n6284 gnd.n6254 5.81868
R19961 gnd.n6252 gnd.n6222 5.81868
R19962 gnd.n6221 gnd.n6191 5.81868
R19963 gnd.n3401 gnd.t92 5.73631
R19964 gnd.t336 gnd.n2311 5.73631
R19965 gnd.n3479 gnd.n2296 5.73631
R19966 gnd.n3492 gnd.n2287 5.73631
R19967 gnd.n3575 gnd.n3574 5.73631
R19968 gnd.n3656 gnd.n3655 5.73631
R19969 gnd.n3768 gnd.n3767 5.73631
R19970 gnd.n3836 gnd.n2107 5.73631
R19971 gnd.n3861 gnd.t135 5.73631
R19972 gnd.t10 gnd.n2008 5.73631
R19973 gnd.n4312 gnd.n1967 5.62001
R19974 gnd.n4914 gnd.n1535 5.62001
R19975 gnd.n4914 gnd.n1536 5.62001
R19976 gnd.n4312 gnd.n1968 5.62001
R19977 gnd.n5742 gnd.n5737 5.4308
R19978 gnd.n5314 gnd.n5312 5.4308
R19979 gnd.n6058 gnd.t3 5.41765
R19980 gnd.t300 gnd.n6081 5.41765
R19981 gnd.t363 gnd.n1049 5.41765
R19982 gnd.t175 gnd.n2654 5.41765
R19983 gnd.n4911 gnd.n1539 5.41765
R19984 gnd.t351 gnd.n3491 5.41765
R19985 gnd.t307 gnd.n2121 5.41765
R19986 gnd.n4635 gnd.t145 5.41765
R19987 gnd.n5103 gnd.n1244 5.09899
R19988 gnd.n5100 gnd.n1249 5.09899
R19989 gnd.n2780 gnd.n1258 5.09899
R19990 gnd.n5094 gnd.n1261 5.09899
R19991 gnd.n2788 gnd.n1269 5.09899
R19992 gnd.n5088 gnd.n1272 5.09899
R19993 gnd.n2838 gnd.n2837 5.09899
R19994 gnd.n5082 gnd.n1282 5.09899
R19995 gnd.n2846 gnd.n1289 5.09899
R19996 gnd.n5076 gnd.n1292 5.09899
R19997 gnd.n2853 gnd.n1300 5.09899
R19998 gnd.n5070 gnd.n1303 5.09899
R19999 gnd.n2862 gnd.n1310 5.09899
R20000 gnd.n5064 gnd.n1313 5.09899
R20001 gnd.n2902 gnd.n2901 5.09899
R20002 gnd.n5058 gnd.n1323 5.09899
R20003 gnd.n2895 gnd.n1330 5.09899
R20004 gnd.n5052 gnd.n1333 5.09899
R20005 gnd.n2889 gnd.n1341 5.09899
R20006 gnd.n5046 gnd.n1344 5.09899
R20007 gnd.n2883 gnd.n1351 5.09899
R20008 gnd.n5040 gnd.n1354 5.09899
R20009 gnd.n2931 gnd.n2690 5.09899
R20010 gnd.n2934 gnd.n2678 5.09899
R20011 gnd.n2945 gnd.n2680 5.09899
R20012 gnd.n2942 gnd.n2684 5.09899
R20013 gnd.n2959 gnd.n2660 5.09899
R20014 gnd.n2972 gnd.n2663 5.09899
R20015 gnd.n2979 gnd.n2654 5.09899
R20016 gnd.n2978 gnd.n2648 5.09899
R20017 gnd.n3007 gnd.n3006 5.09899
R20018 gnd.n5032 gnd.n1371 5.09899
R20019 gnd.n3015 gnd.n1380 5.09899
R20020 gnd.n3022 gnd.n1389 5.09899
R20021 gnd.n5020 gnd.n1392 5.09899
R20022 gnd.n3030 gnd.n1399 5.09899
R20023 gnd.n5014 gnd.n1402 5.09899
R20024 gnd.n3067 gnd.n3066 5.09899
R20025 gnd.n5008 gnd.n1412 5.09899
R20026 gnd.n3037 gnd.n1419 5.09899
R20027 gnd.n3043 gnd.n1429 5.09899
R20028 gnd.n4996 gnd.n1432 5.09899
R20029 gnd.n3049 gnd.n1439 5.09899
R20030 gnd.n4990 gnd.n1442 5.09899
R20031 gnd.n3118 gnd.n3117 5.09899
R20032 gnd.n4984 gnd.n1452 5.09899
R20033 gnd.n3124 gnd.n1459 5.09899
R20034 gnd.n4978 gnd.n1462 5.09899
R20035 gnd.n3133 gnd.n1470 5.09899
R20036 gnd.n4972 gnd.n1473 5.09899
R20037 gnd.n3140 gnd.n1479 5.09899
R20038 gnd.n4966 gnd.n1482 5.09899
R20039 gnd.t17 gnd.n3393 5.09899
R20040 gnd.n3400 gnd.n1599 5.09899
R20041 gnd.t92 gnd.n3400 5.09899
R20042 gnd.n3402 gnd.n1608 5.09899
R20043 gnd.n3559 gnd.n3558 5.09899
R20044 gnd.n3533 gnd.n3532 5.09899
R20045 gnd.n3736 gnd.n3735 5.09899
R20046 gnd.n2164 gnd.n2153 5.09899
R20047 gnd.t50 gnd.n2082 5.09899
R20048 gnd.n3900 gnd.t60 5.09899
R20049 gnd.n4152 gnd.n4151 5.09899
R20050 gnd.n4711 gnd.n4710 5.09899
R20051 gnd.n3925 gnd.n1727 5.09899
R20052 gnd.n4704 gnd.n1736 5.09899
R20053 gnd.n4497 gnd.n1739 5.09899
R20054 gnd.n4698 gnd.n1748 5.09899
R20055 gnd.n4505 gnd.n1751 5.09899
R20056 gnd.n4692 gnd.n1759 5.09899
R20057 gnd.n4511 gnd.n1925 5.09899
R20058 gnd.n4686 gnd.n1768 5.09899
R20059 gnd.n4519 gnd.n1771 5.09899
R20060 gnd.n4680 gnd.n1779 5.09899
R20061 gnd.n4555 gnd.n1782 5.09899
R20062 gnd.n4526 gnd.n1791 5.09899
R20063 gnd.n4668 gnd.n1799 5.09899
R20064 gnd.n4531 gnd.n4530 5.09899
R20065 gnd.n4662 gnd.n1808 5.09899
R20066 gnd.n4538 gnd.n1811 5.09899
R20067 gnd.n4656 gnd.n1819 5.09899
R20068 gnd.n4579 gnd.n1822 5.09899
R20069 gnd.n4609 gnd.n1831 5.09899
R20070 gnd.n4644 gnd.n1837 5.09899
R20071 gnd.n4621 gnd.n4620 5.09899
R20072 gnd.n4638 gnd.n1846 5.09899
R20073 gnd.n4635 gnd.n1849 5.09899
R20074 gnd.n4634 gnd.n1857 5.09899
R20075 gnd.n4599 gnd.n4587 5.09899
R20076 gnd.n7881 gnd.n85 5.09899
R20077 gnd.n391 gnd.n87 5.09899
R20078 gnd.n7578 gnd.n7573 5.09899
R20079 gnd.n7873 gnd.n102 5.09899
R20080 gnd.n7584 gnd.n105 5.09899
R20081 gnd.n7867 gnd.n114 5.09899
R20082 gnd.n7592 gnd.n384 5.09899
R20083 gnd.n7861 gnd.n123 5.09899
R20084 gnd.n7598 gnd.n381 5.09899
R20085 gnd.n7855 gnd.n132 5.09899
R20086 gnd.n7606 gnd.n135 5.09899
R20087 gnd.n7849 gnd.n143 5.09899
R20088 gnd.n7612 gnd.n146 5.09899
R20089 gnd.n7843 gnd.n153 5.09899
R20090 gnd.n7620 gnd.n372 5.09899
R20091 gnd.n7837 gnd.n163 5.09899
R20092 gnd.n7626 gnd.n369 5.09899
R20093 gnd.n7831 gnd.n172 5.09899
R20094 gnd.n7634 gnd.n175 5.09899
R20095 gnd.n7825 gnd.n183 5.09899
R20096 gnd.n7640 gnd.n186 5.09899
R20097 gnd.n7819 gnd.n193 5.09899
R20098 gnd.n7649 gnd.n196 5.09899
R20099 gnd.n7813 gnd.n204 5.09899
R20100 gnd.n7656 gnd.n358 5.09899
R20101 gnd.n7807 gnd.n212 5.09899
R20102 gnd.n6441 gnd.n6440 5.04292
R20103 gnd.n6409 gnd.n6408 5.04292
R20104 gnd.n6377 gnd.n6376 5.04292
R20105 gnd.n6346 gnd.n6345 5.04292
R20106 gnd.n6314 gnd.n6313 5.04292
R20107 gnd.n6282 gnd.n6281 5.04292
R20108 gnd.n6250 gnd.n6249 5.04292
R20109 gnd.n6219 gnd.n6218 5.04292
R20110 gnd.n6021 gnd.t325 4.78034
R20111 gnd.n5344 gnd.t131 4.78034
R20112 gnd.n2883 gnd.t203 4.78034
R20113 gnd.n5026 gnd.t218 4.78034
R20114 gnd.t297 gnd.n2356 4.78034
R20115 gnd.n3492 gnd.t351 4.78034
R20116 gnd.n3768 gnd.t307 4.78034
R20117 gnd.n4309 gnd.t83 4.78034
R20118 gnd.n4127 gnd.t353 4.78034
R20119 gnd.n4650 gnd.t186 4.78034
R20120 gnd.n7867 gnd.t149 4.78034
R20121 gnd.n5463 gnd.n5460 4.74817
R20122 gnd.n5513 gnd.n5395 4.74817
R20123 gnd.n5500 gnd.n5394 4.74817
R20124 gnd.n5393 gnd.n5392 4.74817
R20125 gnd.n5509 gnd.n5460 4.74817
R20126 gnd.n5510 gnd.n5395 4.74817
R20127 gnd.n5512 gnd.n5394 4.74817
R20128 gnd.n5499 gnd.n5393 4.74817
R20129 gnd.n4646 gnd.n98 4.74817
R20130 gnd.n1851 gnd.n96 4.74817
R20131 gnd.n7879 gnd.n91 4.74817
R20132 gnd.n7877 gnd.n92 4.74817
R20133 gnd.n1835 gnd.n98 4.74817
R20134 gnd.n1853 gnd.n96 4.74817
R20135 gnd.n1850 gnd.n91 4.74817
R20136 gnd.n7878 gnd.n7877 4.74817
R20137 gnd.n2929 gnd.n2928 4.74817
R20138 gnd.n2923 gnd.n2919 4.74817
R20139 gnd.n2921 gnd.n2652 4.74817
R20140 gnd.n2983 gnd.n2982 4.74817
R20141 gnd.n3003 gnd.n3002 4.74817
R20142 gnd.n4573 gnd.n1860 4.74817
R20143 gnd.n4626 gnd.n4625 4.74817
R20144 gnd.n4631 gnd.n4630 4.74817
R20145 gnd.n4627 gnd.n394 4.74817
R20146 gnd.n7570 gnd.n7569 4.74817
R20147 gnd.n4574 gnd.n4573 4.74817
R20148 gnd.n4625 gnd.n4624 4.74817
R20149 gnd.n4632 gnd.n4631 4.74817
R20150 gnd.n4629 gnd.n4627 4.74817
R20151 gnd.n7571 gnd.n7570 4.74817
R20152 gnd.n5037 gnd.n5036 4.74817
R20153 gnd.n2658 gnd.n1363 4.74817
R20154 gnd.n2975 gnd.n1362 4.74817
R20155 gnd.n1365 gnd.n1361 4.74817
R20156 gnd.n5036 gnd.n1358 4.74817
R20157 gnd.n2683 gnd.n1363 4.74817
R20158 gnd.n2659 gnd.n1362 4.74817
R20159 gnd.n2976 gnd.n1361 4.74817
R20160 gnd.n2928 gnd.n2927 4.74817
R20161 gnd.n2926 gnd.n2919 4.74817
R20162 gnd.n2922 gnd.n2921 4.74817
R20163 gnd.n2982 gnd.n2981 4.74817
R20164 gnd.n3004 gnd.n3003 4.74817
R20165 gnd.n5458 gnd.n5457 4.74296
R20166 gnd.n78 gnd.n77 4.74296
R20167 gnd.n5426 gnd.n5425 4.7074
R20168 gnd.n5442 gnd.n5441 4.7074
R20169 gnd.n46 gnd.n45 4.7074
R20170 gnd.n62 gnd.n61 4.7074
R20171 gnd.n5458 gnd.n5442 4.65959
R20172 gnd.n78 gnd.n62 4.65959
R20173 gnd.n4403 gnd.n4313 4.6132
R20174 gnd.n4915 gnd.n1534 4.6132
R20175 gnd.n3394 gnd.t17 4.46168
R20176 gnd.n3469 gnd.n3468 4.46168
R20177 gnd.n3478 gnd.t134 4.46168
R20178 gnd.n3490 gnd.n3489 4.46168
R20179 gnd.n3647 gnd.n3646 4.46168
R20180 gnd.n3684 gnd.n3683 4.46168
R20181 gnd.n3826 gnd.n3825 4.46168
R20182 gnd.n3837 gnd.t330 4.46168
R20183 gnd.n3843 gnd.n2109 4.46168
R20184 gnd.n4169 gnd.n4156 4.46111
R20185 gnd.n6426 gnd.n6422 4.38594
R20186 gnd.n6394 gnd.n6390 4.38594
R20187 gnd.n6362 gnd.n6358 4.38594
R20188 gnd.n6331 gnd.n6327 4.38594
R20189 gnd.n6299 gnd.n6295 4.38594
R20190 gnd.n6267 gnd.n6263 4.38594
R20191 gnd.n6235 gnd.n6231 4.38594
R20192 gnd.n6204 gnd.n6200 4.38594
R20193 gnd.n6437 gnd.n6415 4.26717
R20194 gnd.n6405 gnd.n6383 4.26717
R20195 gnd.n6373 gnd.n6351 4.26717
R20196 gnd.n6342 gnd.n6320 4.26717
R20197 gnd.n6310 gnd.n6288 4.26717
R20198 gnd.n6278 gnd.n6256 4.26717
R20199 gnd.n6246 gnd.n6224 4.26717
R20200 gnd.n6215 gnd.n6193 4.26717
R20201 gnd.n5965 gnd.t304 4.14303
R20202 gnd.t301 gnd.n1063 4.14303
R20203 gnd.n2862 gnd.t223 4.14303
R20204 gnd.n5002 gnd.t192 4.14303
R20205 gnd.t32 gnd.n1473 4.14303
R20206 gnd.t20 gnd.n1736 4.14303
R20207 gnd.n4674 gnd.t141 4.14303
R20208 gnd.n7843 gnd.t189 4.14303
R20209 gnd.n6445 gnd.n6444 4.08274
R20210 gnd.n4302 gnd.n4301 4.05904
R20211 gnd.n3335 gnd.n3334 4.05904
R20212 gnd.n4855 gnd.n4848 4.05904
R20213 gnd.n4182 gnd.n4181 4.05904
R20214 gnd.n15 gnd.n7 3.99943
R20215 gnd.n6038 gnd.n5459 3.83315
R20216 gnd.n4827 gnd.n4826 3.82437
R20217 gnd.t133 gnd.n2265 3.82437
R20218 gnd.n3541 gnd.n2256 3.82437
R20219 gnd.n3592 gnd.n2230 3.82437
R20220 gnd.n3666 gnd.n3665 3.82437
R20221 gnd.n3786 gnd.n2142 3.82437
R20222 gnd.n3778 gnd.t310 3.82437
R20223 gnd.n2085 gnd.n2084 3.82437
R20224 gnd.n5442 gnd.n5426 3.72967
R20225 gnd.n62 gnd.n46 3.72967
R20226 gnd.n6445 gnd.n6317 3.70378
R20227 gnd.n15 gnd.n14 3.60163
R20228 gnd.n6436 gnd.n6417 3.49141
R20229 gnd.n6404 gnd.n6385 3.49141
R20230 gnd.n6372 gnd.n6353 3.49141
R20231 gnd.n6341 gnd.n6322 3.49141
R20232 gnd.n6309 gnd.n6290 3.49141
R20233 gnd.n6277 gnd.n6258 3.49141
R20234 gnd.n6245 gnd.n6226 3.49141
R20235 gnd.n6214 gnd.n6195 3.49141
R20236 gnd.n4384 gnd.n4383 3.29747
R20237 gnd.n4383 gnd.n4321 3.29747
R20238 gnd.n7772 gnd.n7769 3.29747
R20239 gnd.n7773 gnd.n7772 3.29747
R20240 gnd.n5191 gnd.n5190 3.29747
R20241 gnd.n5190 gnd.n5189 3.29747
R20242 gnd.n4931 gnd.n4930 3.29747
R20243 gnd.n4930 gnd.n4929 3.29747
R20244 gnd.n3445 gnd.n3444 3.18706
R20245 gnd.n3594 gnd.t129 3.18706
R20246 gnd.n3612 gnd.n2223 3.18706
R20247 gnd.n3674 gnd.n3673 3.18706
R20248 gnd.n3728 gnd.t324 3.18706
R20249 gnd.n3870 gnd.n2092 3.18706
R20250 gnd.n5544 gnd.t304 2.8684
R20251 gnd.t126 gnd.n3401 2.8684
R20252 gnd.t315 gnd.t98 2.8684
R20253 gnd.t333 gnd.n2014 2.8684
R20254 gnd.n5443 gnd.t193 2.82907
R20255 gnd.n5443 gnd.t276 2.82907
R20256 gnd.n5445 gnd.t166 2.82907
R20257 gnd.n5445 gnd.t213 2.82907
R20258 gnd.n5447 gnd.t232 2.82907
R20259 gnd.n5447 gnd.t219 2.82907
R20260 gnd.n5449 gnd.t217 2.82907
R20261 gnd.n5449 gnd.t207 2.82907
R20262 gnd.n5451 gnd.t222 2.82907
R20263 gnd.n5451 gnd.t253 2.82907
R20264 gnd.n5453 gnd.t157 2.82907
R20265 gnd.n5453 gnd.t248 2.82907
R20266 gnd.n5455 gnd.t283 2.82907
R20267 gnd.n5455 gnd.t224 2.82907
R20268 gnd.n5396 gnd.t226 2.82907
R20269 gnd.n5396 gnd.t247 2.82907
R20270 gnd.n5398 gnd.t255 2.82907
R20271 gnd.n5398 gnd.t195 2.82907
R20272 gnd.n5400 gnd.t243 2.82907
R20273 gnd.n5400 gnd.t237 2.82907
R20274 gnd.n5402 gnd.t290 2.82907
R20275 gnd.n5402 gnd.t278 2.82907
R20276 gnd.n5404 gnd.t204 2.82907
R20277 gnd.n5404 gnd.t252 2.82907
R20278 gnd.n5406 gnd.t271 2.82907
R20279 gnd.n5406 gnd.t155 2.82907
R20280 gnd.n5408 gnd.t171 2.82907
R20281 gnd.n5408 gnd.t245 2.82907
R20282 gnd.n5411 gnd.t294 2.82907
R20283 gnd.n5411 gnd.t173 2.82907
R20284 gnd.n5413 gnd.t174 2.82907
R20285 gnd.n5413 gnd.t153 2.82907
R20286 gnd.n5415 gnd.t258 2.82907
R20287 gnd.n5415 gnd.t295 2.82907
R20288 gnd.n5417 gnd.t288 2.82907
R20289 gnd.n5417 gnd.t176 2.82907
R20290 gnd.n5419 gnd.t279 2.82907
R20291 gnd.n5419 gnd.t259 2.82907
R20292 gnd.n5421 gnd.t260 2.82907
R20293 gnd.n5421 gnd.t291 2.82907
R20294 gnd.n5423 gnd.t292 2.82907
R20295 gnd.n5423 gnd.t272 2.82907
R20296 gnd.n5427 gnd.t239 2.82907
R20297 gnd.n5427 gnd.t196 2.82907
R20298 gnd.n5429 gnd.t225 2.82907
R20299 gnd.n5429 gnd.t262 2.82907
R20300 gnd.n5431 gnd.t287 2.82907
R20301 gnd.n5431 gnd.t270 2.82907
R20302 gnd.n5433 gnd.t268 2.82907
R20303 gnd.n5433 gnd.t251 2.82907
R20304 gnd.n5435 gnd.t275 2.82907
R20305 gnd.n5435 gnd.t185 2.82907
R20306 gnd.n5437 gnd.t212 2.82907
R20307 gnd.n5437 gnd.t160 2.82907
R20308 gnd.n5439 gnd.t205 2.82907
R20309 gnd.n5439 gnd.t274 2.82907
R20310 gnd.n75 gnd.t190 2.82907
R20311 gnd.n75 gnd.t244 2.82907
R20312 gnd.n73 gnd.t198 2.82907
R20313 gnd.n73 gnd.t256 2.82907
R20314 gnd.n71 gnd.t228 2.82907
R20315 gnd.n71 gnd.t206 2.82907
R20316 gnd.n69 gnd.t161 2.82907
R20317 gnd.n69 gnd.t182 2.82907
R20318 gnd.n67 gnd.t187 2.82907
R20319 gnd.n67 gnd.t210 2.82907
R20320 gnd.n65 gnd.t179 2.82907
R20321 gnd.n65 gnd.t269 2.82907
R20322 gnd.n63 gnd.t238 2.82907
R20323 gnd.n63 gnd.t142 2.82907
R20324 gnd.n28 gnd.t280 2.82907
R20325 gnd.n28 gnd.t208 2.82907
R20326 gnd.n26 gnd.t200 2.82907
R20327 gnd.n26 gnd.t163 2.82907
R20328 gnd.n24 gnd.t296 2.82907
R20329 gnd.n24 gnd.t191 2.82907
R20330 gnd.n22 gnd.t169 2.82907
R20331 gnd.n22 gnd.t188 2.82907
R20332 gnd.n20 gnd.t267 2.82907
R20333 gnd.n20 gnd.t233 2.82907
R20334 gnd.n18 gnd.t221 2.82907
R20335 gnd.n18 gnd.t151 2.82907
R20336 gnd.n16 gnd.t285 2.82907
R20337 gnd.n16 gnd.t211 2.82907
R20338 gnd.n43 gnd.t250 2.82907
R20339 gnd.n43 gnd.t264 2.82907
R20340 gnd.n41 gnd.t265 2.82907
R20341 gnd.n41 gnd.t242 2.82907
R20342 gnd.n39 gnd.t240 2.82907
R20343 gnd.n39 gnd.t150 2.82907
R20344 gnd.n37 gnd.t146 2.82907
R20345 gnd.n37 gnd.t263 2.82907
R20346 gnd.n35 gnd.t273 2.82907
R20347 gnd.n35 gnd.t282 2.82907
R20348 gnd.n33 gnd.t281 2.82907
R20349 gnd.n33 gnd.t148 2.82907
R20350 gnd.n31 gnd.t138 2.82907
R20351 gnd.n31 gnd.t164 2.82907
R20352 gnd.n59 gnd.t236 2.82907
R20353 gnd.n59 gnd.t144 2.82907
R20354 gnd.n57 gnd.t261 2.82907
R20355 gnd.n57 gnd.t177 2.82907
R20356 gnd.n55 gnd.t284 2.82907
R20357 gnd.n55 gnd.t249 2.82907
R20358 gnd.n53 gnd.t220 2.82907
R20359 gnd.n53 gnd.t234 2.82907
R20360 gnd.n51 gnd.t235 2.82907
R20361 gnd.n51 gnd.t257 2.82907
R20362 gnd.n49 gnd.t229 2.82907
R20363 gnd.n49 gnd.t194 2.82907
R20364 gnd.n47 gnd.t293 2.82907
R20365 gnd.n47 gnd.t215 2.82907
R20366 gnd.n6433 gnd.n6432 2.71565
R20367 gnd.n6401 gnd.n6400 2.71565
R20368 gnd.n6369 gnd.n6368 2.71565
R20369 gnd.n6338 gnd.n6337 2.71565
R20370 gnd.n6306 gnd.n6305 2.71565
R20371 gnd.n6274 gnd.n6273 2.71565
R20372 gnd.n6242 gnd.n6241 2.71565
R20373 gnd.n6211 gnd.n6210 2.71565
R20374 gnd.n3420 gnd.t57 2.54975
R20375 gnd.n3451 gnd.n3446 2.54975
R20376 gnd.n3511 gnd.n2263 2.54975
R20377 gnd.n3613 gnd.n2222 2.54975
R20378 gnd.t321 gnd.n3612 2.54975
R20379 gnd.n3634 gnd.t335 2.54975
R20380 gnd.t350 gnd.n3682 2.54975
R20381 gnd.n3673 gnd.t345 2.54975
R20382 gnd.n3702 gnd.n2182 2.54975
R20383 gnd.n3807 gnd.n2136 2.54975
R20384 gnd.n3869 gnd.n3868 2.54975
R20385 gnd.n3752 gnd.t50 2.54975
R20386 gnd.n6038 gnd.n5460 2.27742
R20387 gnd.n6038 gnd.n5395 2.27742
R20388 gnd.n6038 gnd.n5394 2.27742
R20389 gnd.n6038 gnd.n5393 2.27742
R20390 gnd.n7876 gnd.n98 2.27742
R20391 gnd.n7876 gnd.n96 2.27742
R20392 gnd.n7876 gnd.n91 2.27742
R20393 gnd.n7877 gnd.n7876 2.27742
R20394 gnd.n4573 gnd.n95 2.27742
R20395 gnd.n4625 gnd.n95 2.27742
R20396 gnd.n4631 gnd.n95 2.27742
R20397 gnd.n4627 gnd.n95 2.27742
R20398 gnd.n7570 gnd.n95 2.27742
R20399 gnd.n5036 gnd.n5035 2.27742
R20400 gnd.n5035 gnd.n1363 2.27742
R20401 gnd.n5035 gnd.n1362 2.27742
R20402 gnd.n5035 gnd.n1361 2.27742
R20403 gnd.n2928 gnd.n1360 2.27742
R20404 gnd.n2919 gnd.n1360 2.27742
R20405 gnd.n2921 gnd.n1360 2.27742
R20406 gnd.n2982 gnd.n1360 2.27742
R20407 gnd.n3003 gnd.n1360 2.27742
R20408 gnd.n5892 gnd.t76 2.23109
R20409 gnd.n5515 gnd.t325 2.23109
R20410 gnd.n3568 gnd.t343 2.23109
R20411 gnd.t361 gnd.n3727 2.23109
R20412 gnd.n6429 gnd.n6419 1.93989
R20413 gnd.n6397 gnd.n6387 1.93989
R20414 gnd.n6365 gnd.n6355 1.93989
R20415 gnd.n6334 gnd.n6324 1.93989
R20416 gnd.n6302 gnd.n6292 1.93989
R20417 gnd.n6270 gnd.n6260 1.93989
R20418 gnd.n6238 gnd.n6228 1.93989
R20419 gnd.n6207 gnd.n6197 1.93989
R20420 gnd.n3420 gnd.n1618 1.91244
R20421 gnd.n3513 gnd.t320 1.91244
R20422 gnd.n3534 gnd.t314 1.91244
R20423 gnd.n3604 gnd.n3603 1.91244
R20424 gnd.n3708 gnd.n2178 1.91244
R20425 gnd.t305 gnd.n2162 1.91244
R20426 gnd.n3775 gnd.t311 1.91244
R20427 gnd.n3885 gnd.n3884 1.91244
R20428 gnd.t346 gnd.n5903 1.59378
R20429 gnd.n6082 gnd.t300 1.59378
R20430 gnd.n5330 gnd.t363 1.59378
R20431 gnd.t170 gnd.n1292 1.59378
R20432 gnd.t365 gnd.n2267 1.59378
R20433 gnd.n3798 gnd.t331 1.59378
R20434 gnd.n369 gnd.t143 1.59378
R20435 gnd.n5227 gnd.n5226 1.27512
R20436 gnd.n3470 gnd.n2303 1.27512
R20437 gnd.n3499 gnd.n3498 1.27512
R20438 gnd.t320 gnd.n3512 1.27512
R20439 gnd.n3635 gnd.n3634 1.27512
R20440 gnd.n3682 gnd.n3680 1.27512
R20441 gnd.n3806 gnd.t311 1.27512
R20442 gnd.n3817 gnd.n3816 1.27512
R20443 gnd.n3760 gnd.n3759 1.27512
R20444 gnd.n433 gnd.n223 1.27512
R20445 gnd.n5745 gnd.n5737 1.16414
R20446 gnd.n6504 gnd.n5312 1.16414
R20447 gnd.n6428 gnd.n6421 1.16414
R20448 gnd.n6396 gnd.n6389 1.16414
R20449 gnd.n6364 gnd.n6357 1.16414
R20450 gnd.n6333 gnd.n6326 1.16414
R20451 gnd.n6301 gnd.n6294 1.16414
R20452 gnd.n6269 gnd.n6262 1.16414
R20453 gnd.n6237 gnd.n6230 1.16414
R20454 gnd.n6206 gnd.n6199 1.16414
R20455 gnd.n4313 gnd.n1966 0.970197
R20456 gnd.n4915 gnd.n1531 0.970197
R20457 gnd.n6412 gnd.n6380 0.962709
R20458 gnd.n6444 gnd.n6412 0.962709
R20459 gnd.n6285 gnd.n6253 0.962709
R20460 gnd.n6317 gnd.n6285 0.962709
R20461 gnd.n5991 gnd.t339 0.956468
R20462 gnd.n6627 gnd.t0 0.956468
R20463 gnd.t154 gnd.n1333 0.956468
R20464 gnd.n3042 gnd.t192 0.956468
R20465 gnd.t357 gnd.n2342 0.956468
R20466 gnd.t343 gnd.t129 0.956468
R20467 gnd.t324 gnd.t361 0.956468
R20468 gnd.n4140 gnd.t355 0.956468
R20469 gnd.n4556 gnd.t141 0.956468
R20470 gnd.n381 gnd.t197 0.956468
R20471 gnd.n2 gnd.n1 0.672012
R20472 gnd.n3 gnd.n2 0.672012
R20473 gnd.n4 gnd.n3 0.672012
R20474 gnd.n5 gnd.n4 0.672012
R20475 gnd.n6 gnd.n5 0.672012
R20476 gnd.n7 gnd.n6 0.672012
R20477 gnd.n9 gnd.n8 0.672012
R20478 gnd.n10 gnd.n9 0.672012
R20479 gnd.n11 gnd.n10 0.672012
R20480 gnd.n12 gnd.n11 0.672012
R20481 gnd.n13 gnd.n12 0.672012
R20482 gnd.n14 gnd.n13 0.672012
R20483 gnd.n4841 gnd.n4840 0.637812
R20484 gnd.n4834 gnd.n4833 0.637812
R20485 gnd.n3410 gnd.t53 0.637812
R20486 gnd.t319 gnd.n3469 0.637812
R20487 gnd.n3551 gnd.t136 0.637812
R20488 gnd.n3548 gnd.n2247 0.637812
R20489 gnd.n3569 gnd.n2239 0.637812
R20490 gnd.n3737 gnd.n2159 0.637812
R20491 gnd.n3746 gnd.n3745 0.637812
R20492 gnd.n3788 gnd.t309 0.637812
R20493 gnd.t328 gnd.n2109 0.637812
R20494 gnd.t46 gnd.n2075 0.637812
R20495 gnd.n2077 gnd.n2071 0.637812
R20496 gnd.n4149 gnd.n2017 0.637812
R20497 gnd.n4143 gnd.t83 0.637812
R20498 gnd gnd.n0 0.59317
R20499 gnd.n5457 gnd.n5456 0.573776
R20500 gnd.n5456 gnd.n5454 0.573776
R20501 gnd.n5454 gnd.n5452 0.573776
R20502 gnd.n5452 gnd.n5450 0.573776
R20503 gnd.n5450 gnd.n5448 0.573776
R20504 gnd.n5448 gnd.n5446 0.573776
R20505 gnd.n5446 gnd.n5444 0.573776
R20506 gnd.n5410 gnd.n5409 0.573776
R20507 gnd.n5409 gnd.n5407 0.573776
R20508 gnd.n5407 gnd.n5405 0.573776
R20509 gnd.n5405 gnd.n5403 0.573776
R20510 gnd.n5403 gnd.n5401 0.573776
R20511 gnd.n5401 gnd.n5399 0.573776
R20512 gnd.n5399 gnd.n5397 0.573776
R20513 gnd.n5425 gnd.n5424 0.573776
R20514 gnd.n5424 gnd.n5422 0.573776
R20515 gnd.n5422 gnd.n5420 0.573776
R20516 gnd.n5420 gnd.n5418 0.573776
R20517 gnd.n5418 gnd.n5416 0.573776
R20518 gnd.n5416 gnd.n5414 0.573776
R20519 gnd.n5414 gnd.n5412 0.573776
R20520 gnd.n5441 gnd.n5440 0.573776
R20521 gnd.n5440 gnd.n5438 0.573776
R20522 gnd.n5438 gnd.n5436 0.573776
R20523 gnd.n5436 gnd.n5434 0.573776
R20524 gnd.n5434 gnd.n5432 0.573776
R20525 gnd.n5432 gnd.n5430 0.573776
R20526 gnd.n5430 gnd.n5428 0.573776
R20527 gnd.n66 gnd.n64 0.573776
R20528 gnd.n68 gnd.n66 0.573776
R20529 gnd.n70 gnd.n68 0.573776
R20530 gnd.n72 gnd.n70 0.573776
R20531 gnd.n74 gnd.n72 0.573776
R20532 gnd.n76 gnd.n74 0.573776
R20533 gnd.n77 gnd.n76 0.573776
R20534 gnd.n19 gnd.n17 0.573776
R20535 gnd.n21 gnd.n19 0.573776
R20536 gnd.n23 gnd.n21 0.573776
R20537 gnd.n25 gnd.n23 0.573776
R20538 gnd.n27 gnd.n25 0.573776
R20539 gnd.n29 gnd.n27 0.573776
R20540 gnd.n30 gnd.n29 0.573776
R20541 gnd.n34 gnd.n32 0.573776
R20542 gnd.n36 gnd.n34 0.573776
R20543 gnd.n38 gnd.n36 0.573776
R20544 gnd.n40 gnd.n38 0.573776
R20545 gnd.n42 gnd.n40 0.573776
R20546 gnd.n44 gnd.n42 0.573776
R20547 gnd.n45 gnd.n44 0.573776
R20548 gnd.n50 gnd.n48 0.573776
R20549 gnd.n52 gnd.n50 0.573776
R20550 gnd.n54 gnd.n52 0.573776
R20551 gnd.n56 gnd.n54 0.573776
R20552 gnd.n58 gnd.n56 0.573776
R20553 gnd.n60 gnd.n58 0.573776
R20554 gnd.n61 gnd.n60 0.573776
R20555 gnd.n7888 gnd.n7887 0.553533
R20556 gnd.n7661 gnd.n7660 0.505073
R20557 gnd.n2774 gnd.n2773 0.505073
R20558 gnd.n4102 gnd.n4101 0.489829
R20559 gnd.n3154 gnd.n3153 0.489829
R20560 gnd.n3237 gnd.n2386 0.489829
R20561 gnd.n3988 gnd.n1702 0.489829
R20562 gnd.n6494 gnd.n6493 0.486781
R20563 gnd.n5794 gnd.n5793 0.48678
R20564 gnd.n6575 gnd.n6574 0.480683
R20565 gnd.n5878 gnd.n5877 0.480683
R20566 gnd.n7804 gnd.n7803 0.470012
R20567 gnd.n4339 gnd.n1731 0.470012
R20568 gnd.n4963 gnd.n4962 0.470012
R20569 gnd.n1252 gnd.n1173 0.470012
R20570 gnd.n874 gnd.n869 0.468488
R20571 gnd.n7313 gnd.n557 0.468488
R20572 gnd.n7524 gnd.n431 0.468488
R20573 gnd.n5232 gnd.n5231 0.468488
R20574 gnd.n7876 gnd.n95 0.4255
R20575 gnd.n5035 gnd.n1360 0.4255
R20576 gnd.n3166 gnd.n2598 0.388379
R20577 gnd.n6425 gnd.n6424 0.388379
R20578 gnd.n6393 gnd.n6392 0.388379
R20579 gnd.n6361 gnd.n6360 0.388379
R20580 gnd.n6330 gnd.n6329 0.388379
R20581 gnd.n6298 gnd.n6297 0.388379
R20582 gnd.n6266 gnd.n6265 0.388379
R20583 gnd.n6234 gnd.n6233 0.388379
R20584 gnd.n6203 gnd.n6202 0.388379
R20585 gnd.n4079 gnd.n3936 0.388379
R20586 gnd.n7888 gnd.n15 0.374463
R20587 gnd.n6471 gnd.t303 0.319156
R20588 gnd.n2684 gnd.t216 0.319156
R20589 gnd.n2642 gnd.t218 0.319156
R20590 gnd.n2392 gnd.t69 0.319156
R20591 gnd.n2268 gnd.t365 0.319156
R20592 gnd.t331 gnd.n3797 0.319156
R20593 gnd.n4107 gnd.t42 0.319156
R20594 gnd.n4578 gnd.t186 0.319156
R20595 gnd.t181 gnd.n85 0.319156
R20596 gnd.n5712 gnd.n5690 0.311721
R20597 gnd gnd.n7888 0.295112
R20598 gnd.n7694 gnd.n7693 0.293183
R20599 gnd.n5107 gnd.n1237 0.293183
R20600 gnd.n3145 gnd.n3144 0.27489
R20601 gnd.n3930 gnd.n3929 0.27489
R20602 gnd.n6544 gnd.n6543 0.268793
R20603 gnd.n7695 gnd.n7694 0.258122
R20604 gnd.n4489 gnd.n4488 0.258122
R20605 gnd.n2532 gnd.n2531 0.258122
R20606 gnd.n5108 gnd.n5107 0.258122
R20607 gnd.n6543 gnd.n6542 0.241354
R20608 gnd.n4404 gnd.n4403 0.229039
R20609 gnd.n4403 gnd.n1965 0.229039
R20610 gnd.n1534 gnd.n1530 0.229039
R20611 gnd.n2452 gnd.n1534 0.229039
R20612 gnd.n5866 gnd.n5665 0.206293
R20613 gnd.n5459 gnd.n0 0.169152
R20614 gnd.n6442 gnd.n6414 0.155672
R20615 gnd.n6435 gnd.n6414 0.155672
R20616 gnd.n6435 gnd.n6434 0.155672
R20617 gnd.n6434 gnd.n6418 0.155672
R20618 gnd.n6427 gnd.n6418 0.155672
R20619 gnd.n6427 gnd.n6426 0.155672
R20620 gnd.n6410 gnd.n6382 0.155672
R20621 gnd.n6403 gnd.n6382 0.155672
R20622 gnd.n6403 gnd.n6402 0.155672
R20623 gnd.n6402 gnd.n6386 0.155672
R20624 gnd.n6395 gnd.n6386 0.155672
R20625 gnd.n6395 gnd.n6394 0.155672
R20626 gnd.n6378 gnd.n6350 0.155672
R20627 gnd.n6371 gnd.n6350 0.155672
R20628 gnd.n6371 gnd.n6370 0.155672
R20629 gnd.n6370 gnd.n6354 0.155672
R20630 gnd.n6363 gnd.n6354 0.155672
R20631 gnd.n6363 gnd.n6362 0.155672
R20632 gnd.n6347 gnd.n6319 0.155672
R20633 gnd.n6340 gnd.n6319 0.155672
R20634 gnd.n6340 gnd.n6339 0.155672
R20635 gnd.n6339 gnd.n6323 0.155672
R20636 gnd.n6332 gnd.n6323 0.155672
R20637 gnd.n6332 gnd.n6331 0.155672
R20638 gnd.n6315 gnd.n6287 0.155672
R20639 gnd.n6308 gnd.n6287 0.155672
R20640 gnd.n6308 gnd.n6307 0.155672
R20641 gnd.n6307 gnd.n6291 0.155672
R20642 gnd.n6300 gnd.n6291 0.155672
R20643 gnd.n6300 gnd.n6299 0.155672
R20644 gnd.n6283 gnd.n6255 0.155672
R20645 gnd.n6276 gnd.n6255 0.155672
R20646 gnd.n6276 gnd.n6275 0.155672
R20647 gnd.n6275 gnd.n6259 0.155672
R20648 gnd.n6268 gnd.n6259 0.155672
R20649 gnd.n6268 gnd.n6267 0.155672
R20650 gnd.n6251 gnd.n6223 0.155672
R20651 gnd.n6244 gnd.n6223 0.155672
R20652 gnd.n6244 gnd.n6243 0.155672
R20653 gnd.n6243 gnd.n6227 0.155672
R20654 gnd.n6236 gnd.n6227 0.155672
R20655 gnd.n6236 gnd.n6235 0.155672
R20656 gnd.n6220 gnd.n6192 0.155672
R20657 gnd.n6213 gnd.n6192 0.155672
R20658 gnd.n6213 gnd.n6212 0.155672
R20659 gnd.n6212 gnd.n6196 0.155672
R20660 gnd.n6205 gnd.n6196 0.155672
R20661 gnd.n6205 gnd.n6204 0.155672
R20662 gnd.n6574 gnd.n5242 0.152939
R20663 gnd.n5244 gnd.n5242 0.152939
R20664 gnd.n5248 gnd.n5244 0.152939
R20665 gnd.n5249 gnd.n5248 0.152939
R20666 gnd.n5250 gnd.n5249 0.152939
R20667 gnd.n5251 gnd.n5250 0.152939
R20668 gnd.n5255 gnd.n5251 0.152939
R20669 gnd.n5256 gnd.n5255 0.152939
R20670 gnd.n5257 gnd.n5256 0.152939
R20671 gnd.n5258 gnd.n5257 0.152939
R20672 gnd.n5262 gnd.n5258 0.152939
R20673 gnd.n5263 gnd.n5262 0.152939
R20674 gnd.n5264 gnd.n5263 0.152939
R20675 gnd.n5265 gnd.n5264 0.152939
R20676 gnd.n5270 gnd.n5265 0.152939
R20677 gnd.n6544 gnd.n5270 0.152939
R20678 gnd.n5879 gnd.n5878 0.152939
R20679 gnd.n5879 gnd.n5583 0.152939
R20680 gnd.n5907 gnd.n5583 0.152939
R20681 gnd.n5908 gnd.n5907 0.152939
R20682 gnd.n5909 gnd.n5908 0.152939
R20683 gnd.n5910 gnd.n5909 0.152939
R20684 gnd.n5910 gnd.n5555 0.152939
R20685 gnd.n5937 gnd.n5555 0.152939
R20686 gnd.n5938 gnd.n5937 0.152939
R20687 gnd.n5939 gnd.n5938 0.152939
R20688 gnd.n5939 gnd.n5533 0.152939
R20689 gnd.n5968 gnd.n5533 0.152939
R20690 gnd.n5969 gnd.n5968 0.152939
R20691 gnd.n5970 gnd.n5969 0.152939
R20692 gnd.n5971 gnd.n5970 0.152939
R20693 gnd.n5973 gnd.n5971 0.152939
R20694 gnd.n5973 gnd.n5972 0.152939
R20695 gnd.n5972 gnd.n5482 0.152939
R20696 gnd.n5483 gnd.n5482 0.152939
R20697 gnd.n5484 gnd.n5483 0.152939
R20698 gnd.n5503 gnd.n5484 0.152939
R20699 gnd.n5504 gnd.n5503 0.152939
R20700 gnd.n5504 gnd.n5386 0.152939
R20701 gnd.n6063 gnd.n5386 0.152939
R20702 gnd.n6064 gnd.n6063 0.152939
R20703 gnd.n6065 gnd.n6064 0.152939
R20704 gnd.n6066 gnd.n6065 0.152939
R20705 gnd.n6066 gnd.n5359 0.152939
R20706 gnd.n6103 gnd.n5359 0.152939
R20707 gnd.n6104 gnd.n6103 0.152939
R20708 gnd.n6105 gnd.n6104 0.152939
R20709 gnd.n6106 gnd.n6105 0.152939
R20710 gnd.n6106 gnd.n5333 0.152939
R20711 gnd.n6159 gnd.n5333 0.152939
R20712 gnd.n6160 gnd.n6159 0.152939
R20713 gnd.n6162 gnd.n6160 0.152939
R20714 gnd.n6162 gnd.n6161 0.152939
R20715 gnd.n6161 gnd.n1055 0.152939
R20716 gnd.n1056 gnd.n1055 0.152939
R20717 gnd.n1057 gnd.n1056 0.152939
R20718 gnd.n1078 gnd.n1057 0.152939
R20719 gnd.n1079 gnd.n1078 0.152939
R20720 gnd.n1080 gnd.n1079 0.152939
R20721 gnd.n1081 gnd.n1080 0.152939
R20722 gnd.n1082 gnd.n1081 0.152939
R20723 gnd.n1104 gnd.n1082 0.152939
R20724 gnd.n1105 gnd.n1104 0.152939
R20725 gnd.n1106 gnd.n1105 0.152939
R20726 gnd.n1107 gnd.n1106 0.152939
R20727 gnd.n1108 gnd.n1107 0.152939
R20728 gnd.n5240 gnd.n1108 0.152939
R20729 gnd.n5241 gnd.n5240 0.152939
R20730 gnd.n6575 gnd.n5241 0.152939
R20731 gnd.n5877 gnd.n5607 0.152939
R20732 gnd.n5628 gnd.n5607 0.152939
R20733 gnd.n5629 gnd.n5628 0.152939
R20734 gnd.n5635 gnd.n5629 0.152939
R20735 gnd.n5636 gnd.n5635 0.152939
R20736 gnd.n5637 gnd.n5636 0.152939
R20737 gnd.n5637 gnd.n5626 0.152939
R20738 gnd.n5645 gnd.n5626 0.152939
R20739 gnd.n5646 gnd.n5645 0.152939
R20740 gnd.n5647 gnd.n5646 0.152939
R20741 gnd.n5647 gnd.n5624 0.152939
R20742 gnd.n5655 gnd.n5624 0.152939
R20743 gnd.n5656 gnd.n5655 0.152939
R20744 gnd.n5657 gnd.n5656 0.152939
R20745 gnd.n5657 gnd.n5622 0.152939
R20746 gnd.n5665 gnd.n5622 0.152939
R20747 gnd.n6542 gnd.n5272 0.152939
R20748 gnd.n5274 gnd.n5272 0.152939
R20749 gnd.n5278 gnd.n5274 0.152939
R20750 gnd.n5279 gnd.n5278 0.152939
R20751 gnd.n5280 gnd.n5279 0.152939
R20752 gnd.n5281 gnd.n5280 0.152939
R20753 gnd.n5285 gnd.n5281 0.152939
R20754 gnd.n5286 gnd.n5285 0.152939
R20755 gnd.n5287 gnd.n5286 0.152939
R20756 gnd.n5288 gnd.n5287 0.152939
R20757 gnd.n5292 gnd.n5288 0.152939
R20758 gnd.n5293 gnd.n5292 0.152939
R20759 gnd.n5294 gnd.n5293 0.152939
R20760 gnd.n5295 gnd.n5294 0.152939
R20761 gnd.n5299 gnd.n5295 0.152939
R20762 gnd.n5300 gnd.n5299 0.152939
R20763 gnd.n5301 gnd.n5300 0.152939
R20764 gnd.n5302 gnd.n5301 0.152939
R20765 gnd.n5306 gnd.n5302 0.152939
R20766 gnd.n5307 gnd.n5306 0.152939
R20767 gnd.n5308 gnd.n5307 0.152939
R20768 gnd.n5309 gnd.n5308 0.152939
R20769 gnd.n5316 gnd.n5309 0.152939
R20770 gnd.n5317 gnd.n5316 0.152939
R20771 gnd.n5318 gnd.n5317 0.152939
R20772 gnd.n6494 gnd.n5318 0.152939
R20773 gnd.n6040 gnd.n6039 0.152939
R20774 gnd.n6041 gnd.n6040 0.152939
R20775 gnd.n6042 gnd.n6041 0.152939
R20776 gnd.n6043 gnd.n6042 0.152939
R20777 gnd.n6044 gnd.n6043 0.152939
R20778 gnd.n6045 gnd.n6044 0.152939
R20779 gnd.n6045 gnd.n5340 0.152939
R20780 gnd.n6126 gnd.n5340 0.152939
R20781 gnd.n6127 gnd.n6126 0.152939
R20782 gnd.n6128 gnd.n6127 0.152939
R20783 gnd.n6129 gnd.n6128 0.152939
R20784 gnd.n6130 gnd.n6129 0.152939
R20785 gnd.n6131 gnd.n6130 0.152939
R20786 gnd.n6132 gnd.n6131 0.152939
R20787 gnd.n6133 gnd.n6132 0.152939
R20788 gnd.n6134 gnd.n6133 0.152939
R20789 gnd.n6135 gnd.n6134 0.152939
R20790 gnd.n6136 gnd.n6135 0.152939
R20791 gnd.n6136 gnd.n5323 0.152939
R20792 gnd.n6475 gnd.n5323 0.152939
R20793 gnd.n6476 gnd.n6475 0.152939
R20794 gnd.n6477 gnd.n6476 0.152939
R20795 gnd.n6477 gnd.n5321 0.152939
R20796 gnd.n6485 gnd.n5321 0.152939
R20797 gnd.n6486 gnd.n6485 0.152939
R20798 gnd.n6487 gnd.n6486 0.152939
R20799 gnd.n6487 gnd.n5319 0.152939
R20800 gnd.n6493 gnd.n5319 0.152939
R20801 gnd.n5795 gnd.n5794 0.152939
R20802 gnd.n5795 gnd.n5685 0.152939
R20803 gnd.n5810 gnd.n5685 0.152939
R20804 gnd.n5811 gnd.n5810 0.152939
R20805 gnd.n5812 gnd.n5811 0.152939
R20806 gnd.n5812 gnd.n5673 0.152939
R20807 gnd.n5826 gnd.n5673 0.152939
R20808 gnd.n5827 gnd.n5826 0.152939
R20809 gnd.n5828 gnd.n5827 0.152939
R20810 gnd.n5829 gnd.n5828 0.152939
R20811 gnd.n5830 gnd.n5829 0.152939
R20812 gnd.n5831 gnd.n5830 0.152939
R20813 gnd.n5832 gnd.n5831 0.152939
R20814 gnd.n5833 gnd.n5832 0.152939
R20815 gnd.n5834 gnd.n5833 0.152939
R20816 gnd.n5835 gnd.n5834 0.152939
R20817 gnd.n5836 gnd.n5835 0.152939
R20818 gnd.n5837 gnd.n5836 0.152939
R20819 gnd.n5838 gnd.n5837 0.152939
R20820 gnd.n5839 gnd.n5838 0.152939
R20821 gnd.n5840 gnd.n5839 0.152939
R20822 gnd.n5840 gnd.n5539 0.152939
R20823 gnd.n5957 gnd.n5539 0.152939
R20824 gnd.n5958 gnd.n5957 0.152939
R20825 gnd.n5959 gnd.n5958 0.152939
R20826 gnd.n5960 gnd.n5959 0.152939
R20827 gnd.n5960 gnd.n5461 0.152939
R20828 gnd.n6037 gnd.n5461 0.152939
R20829 gnd.n5713 gnd.n5712 0.152939
R20830 gnd.n5714 gnd.n5713 0.152939
R20831 gnd.n5715 gnd.n5714 0.152939
R20832 gnd.n5716 gnd.n5715 0.152939
R20833 gnd.n5717 gnd.n5716 0.152939
R20834 gnd.n5718 gnd.n5717 0.152939
R20835 gnd.n5719 gnd.n5718 0.152939
R20836 gnd.n5720 gnd.n5719 0.152939
R20837 gnd.n5721 gnd.n5720 0.152939
R20838 gnd.n5722 gnd.n5721 0.152939
R20839 gnd.n5723 gnd.n5722 0.152939
R20840 gnd.n5724 gnd.n5723 0.152939
R20841 gnd.n5725 gnd.n5724 0.152939
R20842 gnd.n5726 gnd.n5725 0.152939
R20843 gnd.n5727 gnd.n5726 0.152939
R20844 gnd.n5728 gnd.n5727 0.152939
R20845 gnd.n5729 gnd.n5728 0.152939
R20846 gnd.n5730 gnd.n5729 0.152939
R20847 gnd.n5731 gnd.n5730 0.152939
R20848 gnd.n5732 gnd.n5731 0.152939
R20849 gnd.n5733 gnd.n5732 0.152939
R20850 gnd.n5734 gnd.n5733 0.152939
R20851 gnd.n5738 gnd.n5734 0.152939
R20852 gnd.n5739 gnd.n5738 0.152939
R20853 gnd.n5739 gnd.n5696 0.152939
R20854 gnd.n5793 gnd.n5696 0.152939
R20855 gnd.n6801 gnd.n869 0.152939
R20856 gnd.n6802 gnd.n6801 0.152939
R20857 gnd.n6803 gnd.n6802 0.152939
R20858 gnd.n6803 gnd.n863 0.152939
R20859 gnd.n6811 gnd.n863 0.152939
R20860 gnd.n6812 gnd.n6811 0.152939
R20861 gnd.n6813 gnd.n6812 0.152939
R20862 gnd.n6813 gnd.n857 0.152939
R20863 gnd.n6821 gnd.n857 0.152939
R20864 gnd.n6822 gnd.n6821 0.152939
R20865 gnd.n6823 gnd.n6822 0.152939
R20866 gnd.n6823 gnd.n851 0.152939
R20867 gnd.n6831 gnd.n851 0.152939
R20868 gnd.n6832 gnd.n6831 0.152939
R20869 gnd.n6833 gnd.n6832 0.152939
R20870 gnd.n6833 gnd.n845 0.152939
R20871 gnd.n6841 gnd.n845 0.152939
R20872 gnd.n6842 gnd.n6841 0.152939
R20873 gnd.n6843 gnd.n6842 0.152939
R20874 gnd.n6843 gnd.n839 0.152939
R20875 gnd.n6851 gnd.n839 0.152939
R20876 gnd.n6852 gnd.n6851 0.152939
R20877 gnd.n6853 gnd.n6852 0.152939
R20878 gnd.n6853 gnd.n833 0.152939
R20879 gnd.n6861 gnd.n833 0.152939
R20880 gnd.n6862 gnd.n6861 0.152939
R20881 gnd.n6863 gnd.n6862 0.152939
R20882 gnd.n6863 gnd.n827 0.152939
R20883 gnd.n6871 gnd.n827 0.152939
R20884 gnd.n6872 gnd.n6871 0.152939
R20885 gnd.n6873 gnd.n6872 0.152939
R20886 gnd.n6873 gnd.n821 0.152939
R20887 gnd.n6881 gnd.n821 0.152939
R20888 gnd.n6882 gnd.n6881 0.152939
R20889 gnd.n6883 gnd.n6882 0.152939
R20890 gnd.n6883 gnd.n815 0.152939
R20891 gnd.n6891 gnd.n815 0.152939
R20892 gnd.n6892 gnd.n6891 0.152939
R20893 gnd.n6893 gnd.n6892 0.152939
R20894 gnd.n6893 gnd.n809 0.152939
R20895 gnd.n6901 gnd.n809 0.152939
R20896 gnd.n6902 gnd.n6901 0.152939
R20897 gnd.n6903 gnd.n6902 0.152939
R20898 gnd.n6903 gnd.n803 0.152939
R20899 gnd.n6911 gnd.n803 0.152939
R20900 gnd.n6912 gnd.n6911 0.152939
R20901 gnd.n6913 gnd.n6912 0.152939
R20902 gnd.n6913 gnd.n797 0.152939
R20903 gnd.n6921 gnd.n797 0.152939
R20904 gnd.n6922 gnd.n6921 0.152939
R20905 gnd.n6923 gnd.n6922 0.152939
R20906 gnd.n6923 gnd.n791 0.152939
R20907 gnd.n6931 gnd.n791 0.152939
R20908 gnd.n6932 gnd.n6931 0.152939
R20909 gnd.n6933 gnd.n6932 0.152939
R20910 gnd.n6933 gnd.n785 0.152939
R20911 gnd.n6941 gnd.n785 0.152939
R20912 gnd.n6942 gnd.n6941 0.152939
R20913 gnd.n6943 gnd.n6942 0.152939
R20914 gnd.n6943 gnd.n779 0.152939
R20915 gnd.n6951 gnd.n779 0.152939
R20916 gnd.n6952 gnd.n6951 0.152939
R20917 gnd.n6953 gnd.n6952 0.152939
R20918 gnd.n6953 gnd.n773 0.152939
R20919 gnd.n6961 gnd.n773 0.152939
R20920 gnd.n6962 gnd.n6961 0.152939
R20921 gnd.n6963 gnd.n6962 0.152939
R20922 gnd.n6963 gnd.n767 0.152939
R20923 gnd.n6971 gnd.n767 0.152939
R20924 gnd.n6972 gnd.n6971 0.152939
R20925 gnd.n6973 gnd.n6972 0.152939
R20926 gnd.n6973 gnd.n761 0.152939
R20927 gnd.n6981 gnd.n761 0.152939
R20928 gnd.n6982 gnd.n6981 0.152939
R20929 gnd.n6983 gnd.n6982 0.152939
R20930 gnd.n6983 gnd.n755 0.152939
R20931 gnd.n6991 gnd.n755 0.152939
R20932 gnd.n6992 gnd.n6991 0.152939
R20933 gnd.n6993 gnd.n6992 0.152939
R20934 gnd.n6993 gnd.n749 0.152939
R20935 gnd.n7001 gnd.n749 0.152939
R20936 gnd.n7002 gnd.n7001 0.152939
R20937 gnd.n7003 gnd.n7002 0.152939
R20938 gnd.n7003 gnd.n743 0.152939
R20939 gnd.n7011 gnd.n743 0.152939
R20940 gnd.n7012 gnd.n7011 0.152939
R20941 gnd.n7013 gnd.n7012 0.152939
R20942 gnd.n7013 gnd.n737 0.152939
R20943 gnd.n7021 gnd.n737 0.152939
R20944 gnd.n7022 gnd.n7021 0.152939
R20945 gnd.n7023 gnd.n7022 0.152939
R20946 gnd.n7023 gnd.n731 0.152939
R20947 gnd.n7031 gnd.n731 0.152939
R20948 gnd.n7032 gnd.n7031 0.152939
R20949 gnd.n7033 gnd.n7032 0.152939
R20950 gnd.n7033 gnd.n725 0.152939
R20951 gnd.n7041 gnd.n725 0.152939
R20952 gnd.n7042 gnd.n7041 0.152939
R20953 gnd.n7043 gnd.n7042 0.152939
R20954 gnd.n7043 gnd.n719 0.152939
R20955 gnd.n7051 gnd.n719 0.152939
R20956 gnd.n7052 gnd.n7051 0.152939
R20957 gnd.n7053 gnd.n7052 0.152939
R20958 gnd.n7053 gnd.n713 0.152939
R20959 gnd.n7061 gnd.n713 0.152939
R20960 gnd.n7062 gnd.n7061 0.152939
R20961 gnd.n7063 gnd.n7062 0.152939
R20962 gnd.n7063 gnd.n707 0.152939
R20963 gnd.n7071 gnd.n707 0.152939
R20964 gnd.n7072 gnd.n7071 0.152939
R20965 gnd.n7073 gnd.n7072 0.152939
R20966 gnd.n7073 gnd.n701 0.152939
R20967 gnd.n7081 gnd.n701 0.152939
R20968 gnd.n7082 gnd.n7081 0.152939
R20969 gnd.n7083 gnd.n7082 0.152939
R20970 gnd.n7083 gnd.n695 0.152939
R20971 gnd.n7091 gnd.n695 0.152939
R20972 gnd.n7092 gnd.n7091 0.152939
R20973 gnd.n7093 gnd.n7092 0.152939
R20974 gnd.n7093 gnd.n689 0.152939
R20975 gnd.n7101 gnd.n689 0.152939
R20976 gnd.n7102 gnd.n7101 0.152939
R20977 gnd.n7103 gnd.n7102 0.152939
R20978 gnd.n7103 gnd.n683 0.152939
R20979 gnd.n7111 gnd.n683 0.152939
R20980 gnd.n7112 gnd.n7111 0.152939
R20981 gnd.n7113 gnd.n7112 0.152939
R20982 gnd.n7113 gnd.n677 0.152939
R20983 gnd.n7121 gnd.n677 0.152939
R20984 gnd.n7122 gnd.n7121 0.152939
R20985 gnd.n7123 gnd.n7122 0.152939
R20986 gnd.n7123 gnd.n671 0.152939
R20987 gnd.n7131 gnd.n671 0.152939
R20988 gnd.n7132 gnd.n7131 0.152939
R20989 gnd.n7133 gnd.n7132 0.152939
R20990 gnd.n7133 gnd.n665 0.152939
R20991 gnd.n7141 gnd.n665 0.152939
R20992 gnd.n7142 gnd.n7141 0.152939
R20993 gnd.n7143 gnd.n7142 0.152939
R20994 gnd.n7143 gnd.n659 0.152939
R20995 gnd.n7151 gnd.n659 0.152939
R20996 gnd.n7152 gnd.n7151 0.152939
R20997 gnd.n7153 gnd.n7152 0.152939
R20998 gnd.n7153 gnd.n653 0.152939
R20999 gnd.n7161 gnd.n653 0.152939
R21000 gnd.n7162 gnd.n7161 0.152939
R21001 gnd.n7163 gnd.n7162 0.152939
R21002 gnd.n7163 gnd.n647 0.152939
R21003 gnd.n7171 gnd.n647 0.152939
R21004 gnd.n7172 gnd.n7171 0.152939
R21005 gnd.n7173 gnd.n7172 0.152939
R21006 gnd.n7173 gnd.n641 0.152939
R21007 gnd.n7181 gnd.n641 0.152939
R21008 gnd.n7182 gnd.n7181 0.152939
R21009 gnd.n7183 gnd.n7182 0.152939
R21010 gnd.n7183 gnd.n635 0.152939
R21011 gnd.n7191 gnd.n635 0.152939
R21012 gnd.n7192 gnd.n7191 0.152939
R21013 gnd.n7193 gnd.n7192 0.152939
R21014 gnd.n7193 gnd.n629 0.152939
R21015 gnd.n7201 gnd.n629 0.152939
R21016 gnd.n7202 gnd.n7201 0.152939
R21017 gnd.n7203 gnd.n7202 0.152939
R21018 gnd.n7203 gnd.n623 0.152939
R21019 gnd.n7211 gnd.n623 0.152939
R21020 gnd.n7212 gnd.n7211 0.152939
R21021 gnd.n7213 gnd.n7212 0.152939
R21022 gnd.n7213 gnd.n617 0.152939
R21023 gnd.n7221 gnd.n617 0.152939
R21024 gnd.n7222 gnd.n7221 0.152939
R21025 gnd.n7223 gnd.n7222 0.152939
R21026 gnd.n7223 gnd.n611 0.152939
R21027 gnd.n7231 gnd.n611 0.152939
R21028 gnd.n7232 gnd.n7231 0.152939
R21029 gnd.n7233 gnd.n7232 0.152939
R21030 gnd.n7233 gnd.n605 0.152939
R21031 gnd.n7241 gnd.n605 0.152939
R21032 gnd.n7242 gnd.n7241 0.152939
R21033 gnd.n7243 gnd.n7242 0.152939
R21034 gnd.n7243 gnd.n599 0.152939
R21035 gnd.n7251 gnd.n599 0.152939
R21036 gnd.n7252 gnd.n7251 0.152939
R21037 gnd.n7253 gnd.n7252 0.152939
R21038 gnd.n7253 gnd.n593 0.152939
R21039 gnd.n7261 gnd.n593 0.152939
R21040 gnd.n7262 gnd.n7261 0.152939
R21041 gnd.n7263 gnd.n7262 0.152939
R21042 gnd.n7263 gnd.n587 0.152939
R21043 gnd.n7271 gnd.n587 0.152939
R21044 gnd.n7272 gnd.n7271 0.152939
R21045 gnd.n7273 gnd.n7272 0.152939
R21046 gnd.n7273 gnd.n581 0.152939
R21047 gnd.n7281 gnd.n581 0.152939
R21048 gnd.n7282 gnd.n7281 0.152939
R21049 gnd.n7283 gnd.n7282 0.152939
R21050 gnd.n7283 gnd.n575 0.152939
R21051 gnd.n7291 gnd.n575 0.152939
R21052 gnd.n7292 gnd.n7291 0.152939
R21053 gnd.n7293 gnd.n7292 0.152939
R21054 gnd.n7293 gnd.n569 0.152939
R21055 gnd.n7301 gnd.n569 0.152939
R21056 gnd.n7302 gnd.n7301 0.152939
R21057 gnd.n7303 gnd.n7302 0.152939
R21058 gnd.n7303 gnd.n563 0.152939
R21059 gnd.n7311 gnd.n563 0.152939
R21060 gnd.n7312 gnd.n7311 0.152939
R21061 gnd.n7313 gnd.n7312 0.152939
R21062 gnd.n7321 gnd.n557 0.152939
R21063 gnd.n7322 gnd.n7321 0.152939
R21064 gnd.n7323 gnd.n7322 0.152939
R21065 gnd.n7323 gnd.n551 0.152939
R21066 gnd.n7331 gnd.n551 0.152939
R21067 gnd.n7332 gnd.n7331 0.152939
R21068 gnd.n7333 gnd.n7332 0.152939
R21069 gnd.n7333 gnd.n545 0.152939
R21070 gnd.n7341 gnd.n545 0.152939
R21071 gnd.n7342 gnd.n7341 0.152939
R21072 gnd.n7343 gnd.n7342 0.152939
R21073 gnd.n7343 gnd.n539 0.152939
R21074 gnd.n7351 gnd.n539 0.152939
R21075 gnd.n7352 gnd.n7351 0.152939
R21076 gnd.n7353 gnd.n7352 0.152939
R21077 gnd.n7353 gnd.n533 0.152939
R21078 gnd.n7361 gnd.n533 0.152939
R21079 gnd.n7362 gnd.n7361 0.152939
R21080 gnd.n7363 gnd.n7362 0.152939
R21081 gnd.n7363 gnd.n527 0.152939
R21082 gnd.n7371 gnd.n527 0.152939
R21083 gnd.n7372 gnd.n7371 0.152939
R21084 gnd.n7373 gnd.n7372 0.152939
R21085 gnd.n7373 gnd.n521 0.152939
R21086 gnd.n7381 gnd.n521 0.152939
R21087 gnd.n7382 gnd.n7381 0.152939
R21088 gnd.n7383 gnd.n7382 0.152939
R21089 gnd.n7383 gnd.n515 0.152939
R21090 gnd.n7391 gnd.n515 0.152939
R21091 gnd.n7392 gnd.n7391 0.152939
R21092 gnd.n7393 gnd.n7392 0.152939
R21093 gnd.n7393 gnd.n509 0.152939
R21094 gnd.n7401 gnd.n509 0.152939
R21095 gnd.n7402 gnd.n7401 0.152939
R21096 gnd.n7403 gnd.n7402 0.152939
R21097 gnd.n7403 gnd.n503 0.152939
R21098 gnd.n7411 gnd.n503 0.152939
R21099 gnd.n7412 gnd.n7411 0.152939
R21100 gnd.n7413 gnd.n7412 0.152939
R21101 gnd.n7413 gnd.n497 0.152939
R21102 gnd.n7421 gnd.n497 0.152939
R21103 gnd.n7422 gnd.n7421 0.152939
R21104 gnd.n7423 gnd.n7422 0.152939
R21105 gnd.n7423 gnd.n491 0.152939
R21106 gnd.n7431 gnd.n491 0.152939
R21107 gnd.n7432 gnd.n7431 0.152939
R21108 gnd.n7433 gnd.n7432 0.152939
R21109 gnd.n7433 gnd.n485 0.152939
R21110 gnd.n7441 gnd.n485 0.152939
R21111 gnd.n7442 gnd.n7441 0.152939
R21112 gnd.n7443 gnd.n7442 0.152939
R21113 gnd.n7443 gnd.n479 0.152939
R21114 gnd.n7451 gnd.n479 0.152939
R21115 gnd.n7452 gnd.n7451 0.152939
R21116 gnd.n7453 gnd.n7452 0.152939
R21117 gnd.n7453 gnd.n473 0.152939
R21118 gnd.n7461 gnd.n473 0.152939
R21119 gnd.n7462 gnd.n7461 0.152939
R21120 gnd.n7463 gnd.n7462 0.152939
R21121 gnd.n7463 gnd.n467 0.152939
R21122 gnd.n7471 gnd.n467 0.152939
R21123 gnd.n7472 gnd.n7471 0.152939
R21124 gnd.n7473 gnd.n7472 0.152939
R21125 gnd.n7473 gnd.n461 0.152939
R21126 gnd.n7481 gnd.n461 0.152939
R21127 gnd.n7482 gnd.n7481 0.152939
R21128 gnd.n7483 gnd.n7482 0.152939
R21129 gnd.n7483 gnd.n455 0.152939
R21130 gnd.n7491 gnd.n455 0.152939
R21131 gnd.n7492 gnd.n7491 0.152939
R21132 gnd.n7493 gnd.n7492 0.152939
R21133 gnd.n7493 gnd.n449 0.152939
R21134 gnd.n7501 gnd.n449 0.152939
R21135 gnd.n7502 gnd.n7501 0.152939
R21136 gnd.n7503 gnd.n7502 0.152939
R21137 gnd.n7503 gnd.n443 0.152939
R21138 gnd.n7511 gnd.n443 0.152939
R21139 gnd.n7512 gnd.n7511 0.152939
R21140 gnd.n7513 gnd.n7512 0.152939
R21141 gnd.n7513 gnd.n437 0.152939
R21142 gnd.n7521 gnd.n437 0.152939
R21143 gnd.n7522 gnd.n7521 0.152939
R21144 gnd.n7523 gnd.n7522 0.152939
R21145 gnd.n7524 gnd.n7523 0.152939
R21146 gnd.n398 gnd.n395 0.152939
R21147 gnd.n399 gnd.n398 0.152939
R21148 gnd.n400 gnd.n399 0.152939
R21149 gnd.n401 gnd.n400 0.152939
R21150 gnd.n404 gnd.n401 0.152939
R21151 gnd.n405 gnd.n404 0.152939
R21152 gnd.n406 gnd.n405 0.152939
R21153 gnd.n407 gnd.n406 0.152939
R21154 gnd.n410 gnd.n407 0.152939
R21155 gnd.n411 gnd.n410 0.152939
R21156 gnd.n412 gnd.n411 0.152939
R21157 gnd.n413 gnd.n412 0.152939
R21158 gnd.n416 gnd.n413 0.152939
R21159 gnd.n417 gnd.n416 0.152939
R21160 gnd.n418 gnd.n417 0.152939
R21161 gnd.n419 gnd.n418 0.152939
R21162 gnd.n422 gnd.n419 0.152939
R21163 gnd.n423 gnd.n422 0.152939
R21164 gnd.n424 gnd.n423 0.152939
R21165 gnd.n425 gnd.n424 0.152939
R21166 gnd.n428 gnd.n425 0.152939
R21167 gnd.n429 gnd.n428 0.152939
R21168 gnd.n430 gnd.n429 0.152939
R21169 gnd.n431 gnd.n430 0.152939
R21170 gnd.n118 gnd.n93 0.152939
R21171 gnd.n119 gnd.n118 0.152939
R21172 gnd.n120 gnd.n119 0.152939
R21173 gnd.n137 gnd.n120 0.152939
R21174 gnd.n138 gnd.n137 0.152939
R21175 gnd.n139 gnd.n138 0.152939
R21176 gnd.n140 gnd.n139 0.152939
R21177 gnd.n157 gnd.n140 0.152939
R21178 gnd.n158 gnd.n157 0.152939
R21179 gnd.n159 gnd.n158 0.152939
R21180 gnd.n160 gnd.n159 0.152939
R21181 gnd.n177 gnd.n160 0.152939
R21182 gnd.n178 gnd.n177 0.152939
R21183 gnd.n179 gnd.n178 0.152939
R21184 gnd.n180 gnd.n179 0.152939
R21185 gnd.n198 gnd.n180 0.152939
R21186 gnd.n199 gnd.n198 0.152939
R21187 gnd.n200 gnd.n199 0.152939
R21188 gnd.n201 gnd.n200 0.152939
R21189 gnd.n217 gnd.n201 0.152939
R21190 gnd.n7804 gnd.n217 0.152939
R21191 gnd.n7885 gnd.n80 0.152939
R21192 gnd.n7574 gnd.n80 0.152939
R21193 gnd.n7575 gnd.n7574 0.152939
R21194 gnd.n7575 gnd.n386 0.152939
R21195 gnd.n7587 gnd.n386 0.152939
R21196 gnd.n7588 gnd.n7587 0.152939
R21197 gnd.n7589 gnd.n7588 0.152939
R21198 gnd.n7589 gnd.n379 0.152939
R21199 gnd.n7601 gnd.n379 0.152939
R21200 gnd.n7602 gnd.n7601 0.152939
R21201 gnd.n7603 gnd.n7602 0.152939
R21202 gnd.n7603 gnd.n374 0.152939
R21203 gnd.n7615 gnd.n374 0.152939
R21204 gnd.n7616 gnd.n7615 0.152939
R21205 gnd.n7617 gnd.n7616 0.152939
R21206 gnd.n7617 gnd.n367 0.152939
R21207 gnd.n7629 gnd.n367 0.152939
R21208 gnd.n7630 gnd.n7629 0.152939
R21209 gnd.n7631 gnd.n7630 0.152939
R21210 gnd.n7631 gnd.n362 0.152939
R21211 gnd.n7643 gnd.n362 0.152939
R21212 gnd.n7644 gnd.n7643 0.152939
R21213 gnd.n7646 gnd.n7644 0.152939
R21214 gnd.n7646 gnd.n7645 0.152939
R21215 gnd.n7645 gnd.n356 0.152939
R21216 gnd.n7660 gnd.n356 0.152939
R21217 gnd.n7693 gnd.n322 0.152939
R21218 gnd.n324 gnd.n322 0.152939
R21219 gnd.n328 gnd.n324 0.152939
R21220 gnd.n329 gnd.n328 0.152939
R21221 gnd.n330 gnd.n329 0.152939
R21222 gnd.n331 gnd.n330 0.152939
R21223 gnd.n335 gnd.n331 0.152939
R21224 gnd.n336 gnd.n335 0.152939
R21225 gnd.n337 gnd.n336 0.152939
R21226 gnd.n338 gnd.n337 0.152939
R21227 gnd.n342 gnd.n338 0.152939
R21228 gnd.n343 gnd.n342 0.152939
R21229 gnd.n344 gnd.n343 0.152939
R21230 gnd.n345 gnd.n344 0.152939
R21231 gnd.n349 gnd.n345 0.152939
R21232 gnd.n350 gnd.n349 0.152939
R21233 gnd.n7662 gnd.n350 0.152939
R21234 gnd.n7662 gnd.n7661 0.152939
R21235 gnd.n7803 gnd.n218 0.152939
R21236 gnd.n220 gnd.n218 0.152939
R21237 gnd.n225 gnd.n220 0.152939
R21238 gnd.n226 gnd.n225 0.152939
R21239 gnd.n227 gnd.n226 0.152939
R21240 gnd.n228 gnd.n227 0.152939
R21241 gnd.n232 gnd.n228 0.152939
R21242 gnd.n233 gnd.n232 0.152939
R21243 gnd.n234 gnd.n233 0.152939
R21244 gnd.n235 gnd.n234 0.152939
R21245 gnd.n239 gnd.n235 0.152939
R21246 gnd.n240 gnd.n239 0.152939
R21247 gnd.n241 gnd.n240 0.152939
R21248 gnd.n242 gnd.n241 0.152939
R21249 gnd.n246 gnd.n242 0.152939
R21250 gnd.n247 gnd.n246 0.152939
R21251 gnd.n248 gnd.n247 0.152939
R21252 gnd.n249 gnd.n248 0.152939
R21253 gnd.n253 gnd.n249 0.152939
R21254 gnd.n254 gnd.n253 0.152939
R21255 gnd.n255 gnd.n254 0.152939
R21256 gnd.n256 gnd.n255 0.152939
R21257 gnd.n260 gnd.n256 0.152939
R21258 gnd.n261 gnd.n260 0.152939
R21259 gnd.n262 gnd.n261 0.152939
R21260 gnd.n263 gnd.n262 0.152939
R21261 gnd.n267 gnd.n263 0.152939
R21262 gnd.n268 gnd.n267 0.152939
R21263 gnd.n269 gnd.n268 0.152939
R21264 gnd.n270 gnd.n269 0.152939
R21265 gnd.n274 gnd.n270 0.152939
R21266 gnd.n275 gnd.n274 0.152939
R21267 gnd.n276 gnd.n275 0.152939
R21268 gnd.n277 gnd.n276 0.152939
R21269 gnd.n281 gnd.n277 0.152939
R21270 gnd.n282 gnd.n281 0.152939
R21271 gnd.n7734 gnd.n282 0.152939
R21272 gnd.n7734 gnd.n7733 0.152939
R21273 gnd.n7733 gnd.n7732 0.152939
R21274 gnd.n7732 gnd.n286 0.152939
R21275 gnd.n292 gnd.n286 0.152939
R21276 gnd.n293 gnd.n292 0.152939
R21277 gnd.n294 gnd.n293 0.152939
R21278 gnd.n295 gnd.n294 0.152939
R21279 gnd.n299 gnd.n295 0.152939
R21280 gnd.n300 gnd.n299 0.152939
R21281 gnd.n301 gnd.n300 0.152939
R21282 gnd.n302 gnd.n301 0.152939
R21283 gnd.n306 gnd.n302 0.152939
R21284 gnd.n307 gnd.n306 0.152939
R21285 gnd.n308 gnd.n307 0.152939
R21286 gnd.n309 gnd.n308 0.152939
R21287 gnd.n313 gnd.n309 0.152939
R21288 gnd.n314 gnd.n313 0.152939
R21289 gnd.n315 gnd.n314 0.152939
R21290 gnd.n316 gnd.n315 0.152939
R21291 gnd.n321 gnd.n316 0.152939
R21292 gnd.n7695 gnd.n321 0.152939
R21293 gnd.n4340 gnd.n4339 0.152939
R21294 gnd.n4340 gnd.n4336 0.152939
R21295 gnd.n4348 gnd.n4336 0.152939
R21296 gnd.n4349 gnd.n4348 0.152939
R21297 gnd.n4350 gnd.n4349 0.152939
R21298 gnd.n4350 gnd.n4332 0.152939
R21299 gnd.n4358 gnd.n4332 0.152939
R21300 gnd.n4359 gnd.n4358 0.152939
R21301 gnd.n4360 gnd.n4359 0.152939
R21302 gnd.n4360 gnd.n4328 0.152939
R21303 gnd.n4368 gnd.n4328 0.152939
R21304 gnd.n4369 gnd.n4368 0.152939
R21305 gnd.n4370 gnd.n4369 0.152939
R21306 gnd.n4370 gnd.n4324 0.152939
R21307 gnd.n4378 gnd.n4324 0.152939
R21308 gnd.n4379 gnd.n4378 0.152939
R21309 gnd.n4380 gnd.n4379 0.152939
R21310 gnd.n4380 gnd.n4320 0.152939
R21311 gnd.n4391 gnd.n4320 0.152939
R21312 gnd.n4392 gnd.n4391 0.152939
R21313 gnd.n4393 gnd.n4392 0.152939
R21314 gnd.n4393 gnd.n4316 0.152939
R21315 gnd.n4401 gnd.n4316 0.152939
R21316 gnd.n4402 gnd.n4401 0.152939
R21317 gnd.n4404 gnd.n4402 0.152939
R21318 gnd.n4414 gnd.n1965 0.152939
R21319 gnd.n4415 gnd.n4414 0.152939
R21320 gnd.n4416 gnd.n4415 0.152939
R21321 gnd.n4416 gnd.n1961 0.152939
R21322 gnd.n4424 gnd.n1961 0.152939
R21323 gnd.n4425 gnd.n4424 0.152939
R21324 gnd.n4426 gnd.n4425 0.152939
R21325 gnd.n4426 gnd.n1957 0.152939
R21326 gnd.n4436 gnd.n1957 0.152939
R21327 gnd.n4437 gnd.n4436 0.152939
R21328 gnd.n4438 gnd.n4437 0.152939
R21329 gnd.n4438 gnd.n1953 0.152939
R21330 gnd.n4446 gnd.n1953 0.152939
R21331 gnd.n4447 gnd.n4446 0.152939
R21332 gnd.n4448 gnd.n4447 0.152939
R21333 gnd.n4448 gnd.n1949 0.152939
R21334 gnd.n4456 gnd.n1949 0.152939
R21335 gnd.n4457 gnd.n4456 0.152939
R21336 gnd.n4458 gnd.n4457 0.152939
R21337 gnd.n4458 gnd.n1945 0.152939
R21338 gnd.n4466 gnd.n1945 0.152939
R21339 gnd.n4467 gnd.n4466 0.152939
R21340 gnd.n4468 gnd.n4467 0.152939
R21341 gnd.n4468 gnd.n1941 0.152939
R21342 gnd.n4476 gnd.n1941 0.152939
R21343 gnd.n4477 gnd.n4476 0.152939
R21344 gnd.n4479 gnd.n4477 0.152939
R21345 gnd.n4479 gnd.n4478 0.152939
R21346 gnd.n4478 gnd.n1934 0.152939
R21347 gnd.n4488 gnd.n1934 0.152939
R21348 gnd.n1732 gnd.n1731 0.152939
R21349 gnd.n1733 gnd.n1732 0.152939
R21350 gnd.n1753 gnd.n1733 0.152939
R21351 gnd.n1754 gnd.n1753 0.152939
R21352 gnd.n1755 gnd.n1754 0.152939
R21353 gnd.n1756 gnd.n1755 0.152939
R21354 gnd.n1773 gnd.n1756 0.152939
R21355 gnd.n1774 gnd.n1773 0.152939
R21356 gnd.n1775 gnd.n1774 0.152939
R21357 gnd.n1776 gnd.n1775 0.152939
R21358 gnd.n1793 gnd.n1776 0.152939
R21359 gnd.n1794 gnd.n1793 0.152939
R21360 gnd.n1795 gnd.n1794 0.152939
R21361 gnd.n1796 gnd.n1795 0.152939
R21362 gnd.n1813 gnd.n1796 0.152939
R21363 gnd.n1814 gnd.n1813 0.152939
R21364 gnd.n1815 gnd.n1814 0.152939
R21365 gnd.n1816 gnd.n1815 0.152939
R21366 gnd.n1833 gnd.n1816 0.152939
R21367 gnd.n1834 gnd.n1833 0.152939
R21368 gnd.n1834 gnd.n94 0.152939
R21369 gnd.n2987 gnd.n2984 0.152939
R21370 gnd.n2988 gnd.n2987 0.152939
R21371 gnd.n2989 gnd.n2988 0.152939
R21372 gnd.n2990 gnd.n2989 0.152939
R21373 gnd.n2992 gnd.n2990 0.152939
R21374 gnd.n2992 gnd.n2991 0.152939
R21375 gnd.n2991 gnd.n2625 0.152939
R21376 gnd.n3072 gnd.n2625 0.152939
R21377 gnd.n3073 gnd.n3072 0.152939
R21378 gnd.n3074 gnd.n3073 0.152939
R21379 gnd.n3074 gnd.n2621 0.152939
R21380 gnd.n3080 gnd.n2621 0.152939
R21381 gnd.n3081 gnd.n3080 0.152939
R21382 gnd.n3082 gnd.n3081 0.152939
R21383 gnd.n3083 gnd.n3082 0.152939
R21384 gnd.n3084 gnd.n3083 0.152939
R21385 gnd.n3087 gnd.n3084 0.152939
R21386 gnd.n3088 gnd.n3087 0.152939
R21387 gnd.n3089 gnd.n3088 0.152939
R21388 gnd.n3090 gnd.n3089 0.152939
R21389 gnd.n3093 gnd.n3090 0.152939
R21390 gnd.n3094 gnd.n3093 0.152939
R21391 gnd.n3095 gnd.n3094 0.152939
R21392 gnd.n3096 gnd.n3095 0.152939
R21393 gnd.n3096 gnd.n2395 0.152939
R21394 gnd.n3226 gnd.n2395 0.152939
R21395 gnd.n3227 gnd.n3226 0.152939
R21396 gnd.n3228 gnd.n3227 0.152939
R21397 gnd.n3229 gnd.n3228 0.152939
R21398 gnd.n3229 gnd.n2371 0.152939
R21399 gnd.n3256 gnd.n2371 0.152939
R21400 gnd.n3257 gnd.n3256 0.152939
R21401 gnd.n3258 gnd.n3257 0.152939
R21402 gnd.n3259 gnd.n3258 0.152939
R21403 gnd.n3259 gnd.n2346 0.152939
R21404 gnd.n3288 gnd.n2346 0.152939
R21405 gnd.n3289 gnd.n3288 0.152939
R21406 gnd.n3290 gnd.n3289 0.152939
R21407 gnd.n3291 gnd.n3290 0.152939
R21408 gnd.n3293 gnd.n3291 0.152939
R21409 gnd.n3293 gnd.n3292 0.152939
R21410 gnd.n3292 gnd.n1603 0.152939
R21411 gnd.n1604 gnd.n1603 0.152939
R21412 gnd.n1605 gnd.n1604 0.152939
R21413 gnd.n2315 gnd.n1605 0.152939
R21414 gnd.n2316 gnd.n2315 0.152939
R21415 gnd.n3455 gnd.n2316 0.152939
R21416 gnd.n3456 gnd.n3455 0.152939
R21417 gnd.n3457 gnd.n3456 0.152939
R21418 gnd.n3457 gnd.n2293 0.152939
R21419 gnd.n3482 gnd.n2293 0.152939
R21420 gnd.n3483 gnd.n3482 0.152939
R21421 gnd.n3484 gnd.n3483 0.152939
R21422 gnd.n3485 gnd.n3484 0.152939
R21423 gnd.n3485 gnd.n2260 0.152939
R21424 gnd.n3524 gnd.n2260 0.152939
R21425 gnd.n3525 gnd.n3524 0.152939
R21426 gnd.n3526 gnd.n3525 0.152939
R21427 gnd.n3527 gnd.n3526 0.152939
R21428 gnd.n3528 gnd.n3527 0.152939
R21429 gnd.n3529 gnd.n3528 0.152939
R21430 gnd.n3529 gnd.n2226 0.152939
R21431 gnd.n3607 gnd.n2226 0.152939
R21432 gnd.n3608 gnd.n3607 0.152939
R21433 gnd.n3609 gnd.n3608 0.152939
R21434 gnd.n3609 gnd.n2203 0.152939
R21435 gnd.n3650 gnd.n2203 0.152939
R21436 gnd.n3651 gnd.n3650 0.152939
R21437 gnd.n3652 gnd.n3651 0.152939
R21438 gnd.n3652 gnd.n2187 0.152939
R21439 gnd.n3694 gnd.n2187 0.152939
R21440 gnd.n3695 gnd.n3694 0.152939
R21441 gnd.n3696 gnd.n3695 0.152939
R21442 gnd.n3697 gnd.n3696 0.152939
R21443 gnd.n3697 gnd.n2156 0.152939
R21444 gnd.n3740 gnd.n2156 0.152939
R21445 gnd.n3741 gnd.n3740 0.152939
R21446 gnd.n3742 gnd.n3741 0.152939
R21447 gnd.n3742 gnd.n2139 0.152939
R21448 gnd.n3801 gnd.n2139 0.152939
R21449 gnd.n3802 gnd.n3801 0.152939
R21450 gnd.n3803 gnd.n3802 0.152939
R21451 gnd.n3803 gnd.n2117 0.152939
R21452 gnd.n3829 gnd.n2117 0.152939
R21453 gnd.n3830 gnd.n3829 0.152939
R21454 gnd.n3831 gnd.n3830 0.152939
R21455 gnd.n3832 gnd.n3831 0.152939
R21456 gnd.n3832 gnd.n2089 0.152939
R21457 gnd.n3873 gnd.n2089 0.152939
R21458 gnd.n3874 gnd.n3873 0.152939
R21459 gnd.n3875 gnd.n3874 0.152939
R21460 gnd.n3876 gnd.n3875 0.152939
R21461 gnd.n3878 gnd.n3876 0.152939
R21462 gnd.n3878 gnd.n3877 0.152939
R21463 gnd.n3877 gnd.n2021 0.152939
R21464 gnd.n2022 gnd.n2021 0.152939
R21465 gnd.n2023 gnd.n2022 0.152939
R21466 gnd.n2030 gnd.n2023 0.152939
R21467 gnd.n2031 gnd.n2030 0.152939
R21468 gnd.n2032 gnd.n2031 0.152939
R21469 gnd.n2033 gnd.n2032 0.152939
R21470 gnd.n2041 gnd.n2033 0.152939
R21471 gnd.n2042 gnd.n2041 0.152939
R21472 gnd.n2043 gnd.n2042 0.152939
R21473 gnd.n2044 gnd.n2043 0.152939
R21474 gnd.n4109 gnd.n2044 0.152939
R21475 gnd.n4110 gnd.n4109 0.152939
R21476 gnd.n4112 gnd.n4110 0.152939
R21477 gnd.n4112 gnd.n4111 0.152939
R21478 gnd.n4111 gnd.n1710 0.152939
R21479 gnd.n1711 gnd.n1710 0.152939
R21480 gnd.n1712 gnd.n1711 0.152939
R21481 gnd.n1718 gnd.n1712 0.152939
R21482 gnd.n1719 gnd.n1718 0.152939
R21483 gnd.n1720 gnd.n1719 0.152939
R21484 gnd.n1721 gnd.n1720 0.152939
R21485 gnd.n1901 gnd.n1721 0.152939
R21486 gnd.n1902 gnd.n1901 0.152939
R21487 gnd.n1903 gnd.n1902 0.152939
R21488 gnd.n1903 gnd.n1897 0.152939
R21489 gnd.n1909 gnd.n1897 0.152939
R21490 gnd.n1910 gnd.n1909 0.152939
R21491 gnd.n1911 gnd.n1910 0.152939
R21492 gnd.n1912 gnd.n1911 0.152939
R21493 gnd.n1913 gnd.n1912 0.152939
R21494 gnd.n1914 gnd.n1913 0.152939
R21495 gnd.n1916 gnd.n1914 0.152939
R21496 gnd.n1916 gnd.n1915 0.152939
R21497 gnd.n1915 gnd.n1876 0.152939
R21498 gnd.n4561 gnd.n1876 0.152939
R21499 gnd.n4562 gnd.n4561 0.152939
R21500 gnd.n4563 gnd.n4562 0.152939
R21501 gnd.n4563 gnd.n1872 0.152939
R21502 gnd.n4569 gnd.n1872 0.152939
R21503 gnd.n4570 gnd.n4569 0.152939
R21504 gnd.n4571 gnd.n4570 0.152939
R21505 gnd.n4572 gnd.n4571 0.152939
R21506 gnd.n2774 gnd.n2717 0.152939
R21507 gnd.n2783 gnd.n2717 0.152939
R21508 gnd.n2784 gnd.n2783 0.152939
R21509 gnd.n2785 gnd.n2784 0.152939
R21510 gnd.n2785 gnd.n2713 0.152939
R21511 gnd.n2841 gnd.n2713 0.152939
R21512 gnd.n2842 gnd.n2841 0.152939
R21513 gnd.n2843 gnd.n2842 0.152939
R21514 gnd.n2843 gnd.n2709 0.152939
R21515 gnd.n2856 gnd.n2709 0.152939
R21516 gnd.n2857 gnd.n2856 0.152939
R21517 gnd.n2859 gnd.n2857 0.152939
R21518 gnd.n2859 gnd.n2858 0.152939
R21519 gnd.n2858 gnd.n2703 0.152939
R21520 gnd.n2704 gnd.n2703 0.152939
R21521 gnd.n2705 gnd.n2704 0.152939
R21522 gnd.n2871 gnd.n2705 0.152939
R21523 gnd.n2872 gnd.n2871 0.152939
R21524 gnd.n2873 gnd.n2872 0.152939
R21525 gnd.n2874 gnd.n2873 0.152939
R21526 gnd.n2875 gnd.n2874 0.152939
R21527 gnd.n2876 gnd.n2875 0.152939
R21528 gnd.n2876 gnd.n2675 0.152939
R21529 gnd.n2948 gnd.n2675 0.152939
R21530 gnd.n2949 gnd.n2948 0.152939
R21531 gnd.n2950 gnd.n2949 0.152939
R21532 gnd.n2731 gnd.n1237 0.152939
R21533 gnd.n2737 gnd.n2731 0.152939
R21534 gnd.n2738 gnd.n2737 0.152939
R21535 gnd.n2739 gnd.n2738 0.152939
R21536 gnd.n2739 gnd.n2729 0.152939
R21537 gnd.n2747 gnd.n2729 0.152939
R21538 gnd.n2748 gnd.n2747 0.152939
R21539 gnd.n2749 gnd.n2748 0.152939
R21540 gnd.n2749 gnd.n2727 0.152939
R21541 gnd.n2757 gnd.n2727 0.152939
R21542 gnd.n2758 gnd.n2757 0.152939
R21543 gnd.n2759 gnd.n2758 0.152939
R21544 gnd.n2759 gnd.n2725 0.152939
R21545 gnd.n2767 gnd.n2725 0.152939
R21546 gnd.n2768 gnd.n2767 0.152939
R21547 gnd.n2769 gnd.n2768 0.152939
R21548 gnd.n2769 gnd.n2718 0.152939
R21549 gnd.n2773 gnd.n2718 0.152939
R21550 gnd.n1384 gnd.n1359 0.152939
R21551 gnd.n1385 gnd.n1384 0.152939
R21552 gnd.n1386 gnd.n1385 0.152939
R21553 gnd.n1404 gnd.n1386 0.152939
R21554 gnd.n1405 gnd.n1404 0.152939
R21555 gnd.n1406 gnd.n1405 0.152939
R21556 gnd.n1407 gnd.n1406 0.152939
R21557 gnd.n1423 gnd.n1407 0.152939
R21558 gnd.n1424 gnd.n1423 0.152939
R21559 gnd.n1425 gnd.n1424 0.152939
R21560 gnd.n1426 gnd.n1425 0.152939
R21561 gnd.n1444 gnd.n1426 0.152939
R21562 gnd.n1445 gnd.n1444 0.152939
R21563 gnd.n1446 gnd.n1445 0.152939
R21564 gnd.n1447 gnd.n1446 0.152939
R21565 gnd.n1464 gnd.n1447 0.152939
R21566 gnd.n1465 gnd.n1464 0.152939
R21567 gnd.n1466 gnd.n1465 0.152939
R21568 gnd.n1467 gnd.n1466 0.152939
R21569 gnd.n1484 gnd.n1467 0.152939
R21570 gnd.n4963 gnd.n1484 0.152939
R21571 gnd.n4962 gnd.n1485 0.152939
R21572 gnd.n1490 gnd.n1485 0.152939
R21573 gnd.n1491 gnd.n1490 0.152939
R21574 gnd.n1492 gnd.n1491 0.152939
R21575 gnd.n1493 gnd.n1492 0.152939
R21576 gnd.n1494 gnd.n1493 0.152939
R21577 gnd.n1498 gnd.n1494 0.152939
R21578 gnd.n1499 gnd.n1498 0.152939
R21579 gnd.n1500 gnd.n1499 0.152939
R21580 gnd.n1501 gnd.n1500 0.152939
R21581 gnd.n1505 gnd.n1501 0.152939
R21582 gnd.n1506 gnd.n1505 0.152939
R21583 gnd.n1507 gnd.n1506 0.152939
R21584 gnd.n1508 gnd.n1507 0.152939
R21585 gnd.n1512 gnd.n1508 0.152939
R21586 gnd.n1513 gnd.n1512 0.152939
R21587 gnd.n1514 gnd.n1513 0.152939
R21588 gnd.n1517 gnd.n1514 0.152939
R21589 gnd.n1521 gnd.n1517 0.152939
R21590 gnd.n1522 gnd.n1521 0.152939
R21591 gnd.n1523 gnd.n1522 0.152939
R21592 gnd.n1524 gnd.n1523 0.152939
R21593 gnd.n1528 gnd.n1524 0.152939
R21594 gnd.n1529 gnd.n1528 0.152939
R21595 gnd.n1530 gnd.n1529 0.152939
R21596 gnd.n2453 gnd.n2452 0.152939
R21597 gnd.n2462 gnd.n2453 0.152939
R21598 gnd.n2463 gnd.n2462 0.152939
R21599 gnd.n2464 gnd.n2463 0.152939
R21600 gnd.n2464 gnd.n2448 0.152939
R21601 gnd.n2472 gnd.n2448 0.152939
R21602 gnd.n2473 gnd.n2472 0.152939
R21603 gnd.n2474 gnd.n2473 0.152939
R21604 gnd.n2474 gnd.n2442 0.152939
R21605 gnd.n2482 gnd.n2442 0.152939
R21606 gnd.n2483 gnd.n2482 0.152939
R21607 gnd.n2484 gnd.n2483 0.152939
R21608 gnd.n2484 gnd.n2438 0.152939
R21609 gnd.n2492 gnd.n2438 0.152939
R21610 gnd.n2493 gnd.n2492 0.152939
R21611 gnd.n2494 gnd.n2493 0.152939
R21612 gnd.n2494 gnd.n2434 0.152939
R21613 gnd.n2502 gnd.n2434 0.152939
R21614 gnd.n2503 gnd.n2502 0.152939
R21615 gnd.n2504 gnd.n2503 0.152939
R21616 gnd.n2504 gnd.n2430 0.152939
R21617 gnd.n2512 gnd.n2430 0.152939
R21618 gnd.n2513 gnd.n2512 0.152939
R21619 gnd.n2514 gnd.n2513 0.152939
R21620 gnd.n2514 gnd.n2426 0.152939
R21621 gnd.n2522 gnd.n2426 0.152939
R21622 gnd.n2523 gnd.n2522 0.152939
R21623 gnd.n2524 gnd.n2523 0.152939
R21624 gnd.n2524 gnd.n2420 0.152939
R21625 gnd.n2531 gnd.n2420 0.152939
R21626 gnd.n1174 gnd.n1173 0.152939
R21627 gnd.n1175 gnd.n1174 0.152939
R21628 gnd.n1176 gnd.n1175 0.152939
R21629 gnd.n1177 gnd.n1176 0.152939
R21630 gnd.n1178 gnd.n1177 0.152939
R21631 gnd.n1179 gnd.n1178 0.152939
R21632 gnd.n1180 gnd.n1179 0.152939
R21633 gnd.n1181 gnd.n1180 0.152939
R21634 gnd.n1182 gnd.n1181 0.152939
R21635 gnd.n1183 gnd.n1182 0.152939
R21636 gnd.n1184 gnd.n1183 0.152939
R21637 gnd.n1185 gnd.n1184 0.152939
R21638 gnd.n1186 gnd.n1185 0.152939
R21639 gnd.n1187 gnd.n1186 0.152939
R21640 gnd.n1188 gnd.n1187 0.152939
R21641 gnd.n1189 gnd.n1188 0.152939
R21642 gnd.n1190 gnd.n1189 0.152939
R21643 gnd.n1193 gnd.n1190 0.152939
R21644 gnd.n1194 gnd.n1193 0.152939
R21645 gnd.n1195 gnd.n1194 0.152939
R21646 gnd.n1196 gnd.n1195 0.152939
R21647 gnd.n1197 gnd.n1196 0.152939
R21648 gnd.n1198 gnd.n1197 0.152939
R21649 gnd.n1199 gnd.n1198 0.152939
R21650 gnd.n1200 gnd.n1199 0.152939
R21651 gnd.n1201 gnd.n1200 0.152939
R21652 gnd.n1202 gnd.n1201 0.152939
R21653 gnd.n1203 gnd.n1202 0.152939
R21654 gnd.n1204 gnd.n1203 0.152939
R21655 gnd.n1205 gnd.n1204 0.152939
R21656 gnd.n1206 gnd.n1205 0.152939
R21657 gnd.n1207 gnd.n1206 0.152939
R21658 gnd.n1208 gnd.n1207 0.152939
R21659 gnd.n1209 gnd.n1208 0.152939
R21660 gnd.n1210 gnd.n1209 0.152939
R21661 gnd.n1211 gnd.n1210 0.152939
R21662 gnd.n1212 gnd.n1211 0.152939
R21663 gnd.n1215 gnd.n1212 0.152939
R21664 gnd.n1216 gnd.n1215 0.152939
R21665 gnd.n1217 gnd.n1216 0.152939
R21666 gnd.n1218 gnd.n1217 0.152939
R21667 gnd.n1219 gnd.n1218 0.152939
R21668 gnd.n1220 gnd.n1219 0.152939
R21669 gnd.n1221 gnd.n1220 0.152939
R21670 gnd.n1222 gnd.n1221 0.152939
R21671 gnd.n1223 gnd.n1222 0.152939
R21672 gnd.n1224 gnd.n1223 0.152939
R21673 gnd.n1225 gnd.n1224 0.152939
R21674 gnd.n1226 gnd.n1225 0.152939
R21675 gnd.n1227 gnd.n1226 0.152939
R21676 gnd.n1228 gnd.n1227 0.152939
R21677 gnd.n1229 gnd.n1228 0.152939
R21678 gnd.n1230 gnd.n1229 0.152939
R21679 gnd.n1231 gnd.n1230 0.152939
R21680 gnd.n1232 gnd.n1231 0.152939
R21681 gnd.n1233 gnd.n1232 0.152939
R21682 gnd.n5109 gnd.n1233 0.152939
R21683 gnd.n5109 gnd.n5108 0.152939
R21684 gnd.n1253 gnd.n1252 0.152939
R21685 gnd.n1254 gnd.n1253 0.152939
R21686 gnd.n1255 gnd.n1254 0.152939
R21687 gnd.n1274 gnd.n1255 0.152939
R21688 gnd.n1275 gnd.n1274 0.152939
R21689 gnd.n1276 gnd.n1275 0.152939
R21690 gnd.n1277 gnd.n1276 0.152939
R21691 gnd.n1294 gnd.n1277 0.152939
R21692 gnd.n1295 gnd.n1294 0.152939
R21693 gnd.n1296 gnd.n1295 0.152939
R21694 gnd.n1297 gnd.n1296 0.152939
R21695 gnd.n1315 gnd.n1297 0.152939
R21696 gnd.n1316 gnd.n1315 0.152939
R21697 gnd.n1317 gnd.n1316 0.152939
R21698 gnd.n1318 gnd.n1317 0.152939
R21699 gnd.n1335 gnd.n1318 0.152939
R21700 gnd.n1336 gnd.n1335 0.152939
R21701 gnd.n1337 gnd.n1336 0.152939
R21702 gnd.n1338 gnd.n1337 0.152939
R21703 gnd.n1356 gnd.n1338 0.152939
R21704 gnd.n1357 gnd.n1356 0.152939
R21705 gnd.n5231 gnd.n1128 0.152939
R21706 gnd.n2802 gnd.n1128 0.152939
R21707 gnd.n2805 gnd.n2802 0.152939
R21708 gnd.n2806 gnd.n2805 0.152939
R21709 gnd.n2807 gnd.n2806 0.152939
R21710 gnd.n2807 gnd.n2798 0.152939
R21711 gnd.n2813 gnd.n2798 0.152939
R21712 gnd.n2814 gnd.n2813 0.152939
R21713 gnd.n2815 gnd.n2814 0.152939
R21714 gnd.n2816 gnd.n2815 0.152939
R21715 gnd.n2817 gnd.n2816 0.152939
R21716 gnd.n2820 gnd.n2817 0.152939
R21717 gnd.n2821 gnd.n2820 0.152939
R21718 gnd.n2822 gnd.n2821 0.152939
R21719 gnd.n2823 gnd.n2822 0.152939
R21720 gnd.n2824 gnd.n2823 0.152939
R21721 gnd.n2824 gnd.n2698 0.152939
R21722 gnd.n2906 gnd.n2698 0.152939
R21723 gnd.n2907 gnd.n2906 0.152939
R21724 gnd.n2908 gnd.n2907 0.152939
R21725 gnd.n2908 gnd.n2694 0.152939
R21726 gnd.n2915 gnd.n2694 0.152939
R21727 gnd.n2916 gnd.n2915 0.152939
R21728 gnd.n2917 gnd.n2916 0.152939
R21729 gnd.n875 gnd.n874 0.152939
R21730 gnd.n876 gnd.n875 0.152939
R21731 gnd.n881 gnd.n876 0.152939
R21732 gnd.n882 gnd.n881 0.152939
R21733 gnd.n883 gnd.n882 0.152939
R21734 gnd.n884 gnd.n883 0.152939
R21735 gnd.n889 gnd.n884 0.152939
R21736 gnd.n890 gnd.n889 0.152939
R21737 gnd.n891 gnd.n890 0.152939
R21738 gnd.n892 gnd.n891 0.152939
R21739 gnd.n897 gnd.n892 0.152939
R21740 gnd.n898 gnd.n897 0.152939
R21741 gnd.n899 gnd.n898 0.152939
R21742 gnd.n900 gnd.n899 0.152939
R21743 gnd.n905 gnd.n900 0.152939
R21744 gnd.n906 gnd.n905 0.152939
R21745 gnd.n907 gnd.n906 0.152939
R21746 gnd.n908 gnd.n907 0.152939
R21747 gnd.n913 gnd.n908 0.152939
R21748 gnd.n914 gnd.n913 0.152939
R21749 gnd.n915 gnd.n914 0.152939
R21750 gnd.n916 gnd.n915 0.152939
R21751 gnd.n921 gnd.n916 0.152939
R21752 gnd.n922 gnd.n921 0.152939
R21753 gnd.n923 gnd.n922 0.152939
R21754 gnd.n924 gnd.n923 0.152939
R21755 gnd.n929 gnd.n924 0.152939
R21756 gnd.n930 gnd.n929 0.152939
R21757 gnd.n931 gnd.n930 0.152939
R21758 gnd.n932 gnd.n931 0.152939
R21759 gnd.n937 gnd.n932 0.152939
R21760 gnd.n938 gnd.n937 0.152939
R21761 gnd.n939 gnd.n938 0.152939
R21762 gnd.n940 gnd.n939 0.152939
R21763 gnd.n945 gnd.n940 0.152939
R21764 gnd.n946 gnd.n945 0.152939
R21765 gnd.n947 gnd.n946 0.152939
R21766 gnd.n948 gnd.n947 0.152939
R21767 gnd.n953 gnd.n948 0.152939
R21768 gnd.n954 gnd.n953 0.152939
R21769 gnd.n955 gnd.n954 0.152939
R21770 gnd.n956 gnd.n955 0.152939
R21771 gnd.n961 gnd.n956 0.152939
R21772 gnd.n962 gnd.n961 0.152939
R21773 gnd.n963 gnd.n962 0.152939
R21774 gnd.n964 gnd.n963 0.152939
R21775 gnd.n969 gnd.n964 0.152939
R21776 gnd.n970 gnd.n969 0.152939
R21777 gnd.n971 gnd.n970 0.152939
R21778 gnd.n972 gnd.n971 0.152939
R21779 gnd.n977 gnd.n972 0.152939
R21780 gnd.n978 gnd.n977 0.152939
R21781 gnd.n979 gnd.n978 0.152939
R21782 gnd.n980 gnd.n979 0.152939
R21783 gnd.n985 gnd.n980 0.152939
R21784 gnd.n986 gnd.n985 0.152939
R21785 gnd.n987 gnd.n986 0.152939
R21786 gnd.n988 gnd.n987 0.152939
R21787 gnd.n993 gnd.n988 0.152939
R21788 gnd.n994 gnd.n993 0.152939
R21789 gnd.n995 gnd.n994 0.152939
R21790 gnd.n996 gnd.n995 0.152939
R21791 gnd.n1001 gnd.n996 0.152939
R21792 gnd.n1002 gnd.n1001 0.152939
R21793 gnd.n1003 gnd.n1002 0.152939
R21794 gnd.n1004 gnd.n1003 0.152939
R21795 gnd.n1009 gnd.n1004 0.152939
R21796 gnd.n1010 gnd.n1009 0.152939
R21797 gnd.n1011 gnd.n1010 0.152939
R21798 gnd.n1012 gnd.n1011 0.152939
R21799 gnd.n1017 gnd.n1012 0.152939
R21800 gnd.n1018 gnd.n1017 0.152939
R21801 gnd.n1019 gnd.n1018 0.152939
R21802 gnd.n1020 gnd.n1019 0.152939
R21803 gnd.n1025 gnd.n1020 0.152939
R21804 gnd.n1026 gnd.n1025 0.152939
R21805 gnd.n1027 gnd.n1026 0.152939
R21806 gnd.n1028 gnd.n1027 0.152939
R21807 gnd.n1033 gnd.n1028 0.152939
R21808 gnd.n1034 gnd.n1033 0.152939
R21809 gnd.n1035 gnd.n1034 0.152939
R21810 gnd.n1036 gnd.n1035 0.152939
R21811 gnd.n1127 gnd.n1036 0.152939
R21812 gnd.n5232 gnd.n1127 0.152939
R21813 gnd.n3153 gnd.n2378 0.152939
R21814 gnd.n3246 gnd.n2378 0.152939
R21815 gnd.n3247 gnd.n3246 0.152939
R21816 gnd.n3249 gnd.n3247 0.152939
R21817 gnd.n3249 gnd.n3248 0.152939
R21818 gnd.n3248 gnd.n2353 0.152939
R21819 gnd.n3276 gnd.n2353 0.152939
R21820 gnd.n3277 gnd.n3276 0.152939
R21821 gnd.n3281 gnd.n3277 0.152939
R21822 gnd.n3281 gnd.n3280 0.152939
R21823 gnd.n3280 gnd.n3279 0.152939
R21824 gnd.n3279 gnd.n2329 0.152939
R21825 gnd.n3322 gnd.n2329 0.152939
R21826 gnd.n3323 gnd.n3322 0.152939
R21827 gnd.n3324 gnd.n3323 0.152939
R21828 gnd.n3324 gnd.n2325 0.152939
R21829 gnd.n3413 gnd.n2325 0.152939
R21830 gnd.n3414 gnd.n3413 0.152939
R21831 gnd.n3416 gnd.n3414 0.152939
R21832 gnd.n3416 gnd.n3415 0.152939
R21833 gnd.n3415 gnd.n2300 0.152939
R21834 gnd.n3473 gnd.n2300 0.152939
R21835 gnd.n3474 gnd.n3473 0.152939
R21836 gnd.n3475 gnd.n3474 0.152939
R21837 gnd.n3475 gnd.n2279 0.152939
R21838 gnd.n3502 gnd.n2279 0.152939
R21839 gnd.n3503 gnd.n3502 0.152939
R21840 gnd.n3508 gnd.n3503 0.152939
R21841 gnd.n3508 gnd.n3507 0.152939
R21842 gnd.n3507 gnd.n3506 0.152939
R21843 gnd.n3506 gnd.n2244 0.152939
R21844 gnd.n3562 gnd.n2244 0.152939
R21845 gnd.n3563 gnd.n3562 0.152939
R21846 gnd.n3565 gnd.n3563 0.152939
R21847 gnd.n3565 gnd.n3564 0.152939
R21848 gnd.n3564 gnd.n2219 0.152939
R21849 gnd.n3616 gnd.n2219 0.152939
R21850 gnd.n3617 gnd.n3616 0.152939
R21851 gnd.n3630 gnd.n3617 0.152939
R21852 gnd.n3630 gnd.n3629 0.152939
R21853 gnd.n3629 gnd.n3628 0.152939
R21854 gnd.n3628 gnd.n3618 0.152939
R21855 gnd.n3624 gnd.n3618 0.152939
R21856 gnd.n3624 gnd.n3623 0.152939
R21857 gnd.n3623 gnd.n2173 0.152939
R21858 gnd.n3712 gnd.n2173 0.152939
R21859 gnd.n3713 gnd.n3712 0.152939
R21860 gnd.n3724 gnd.n3713 0.152939
R21861 gnd.n3724 gnd.n3723 0.152939
R21862 gnd.n3723 gnd.n3722 0.152939
R21863 gnd.n3722 gnd.n3714 0.152939
R21864 gnd.n3718 gnd.n3714 0.152939
R21865 gnd.n3718 gnd.n2133 0.152939
R21866 gnd.n3810 gnd.n2133 0.152939
R21867 gnd.n3811 gnd.n3810 0.152939
R21868 gnd.n3813 gnd.n3811 0.152939
R21869 gnd.n3813 gnd.n3812 0.152939
R21870 gnd.n3812 gnd.n2104 0.152939
R21871 gnd.n3848 gnd.n2104 0.152939
R21872 gnd.n3849 gnd.n3848 0.152939
R21873 gnd.n3858 gnd.n3849 0.152939
R21874 gnd.n3858 gnd.n3857 0.152939
R21875 gnd.n3857 gnd.n3856 0.152939
R21876 gnd.n3856 gnd.n3851 0.152939
R21877 gnd.n3851 gnd.n3850 0.152939
R21878 gnd.n3850 gnd.n2068 0.152939
R21879 gnd.n3904 gnd.n2068 0.152939
R21880 gnd.n3905 gnd.n3904 0.152939
R21881 gnd.n3906 gnd.n3905 0.152939
R21882 gnd.n3906 gnd.n2064 0.152939
R21883 gnd.n3910 gnd.n2064 0.152939
R21884 gnd.n3911 gnd.n3910 0.152939
R21885 gnd.n3912 gnd.n3911 0.152939
R21886 gnd.n3912 gnd.n2060 0.152939
R21887 gnd.n3916 gnd.n2060 0.152939
R21888 gnd.n3917 gnd.n3916 0.152939
R21889 gnd.n3918 gnd.n3917 0.152939
R21890 gnd.n3918 gnd.n2054 0.152939
R21891 gnd.n3922 gnd.n2054 0.152939
R21892 gnd.n3923 gnd.n3922 0.152939
R21893 gnd.n4103 gnd.n3923 0.152939
R21894 gnd.n4103 gnd.n4102 0.152939
R21895 gnd.n2955 gnd.n2954 0.152939
R21896 gnd.n2954 gnd.n2645 0.152939
R21897 gnd.n3010 gnd.n2645 0.152939
R21898 gnd.n3011 gnd.n3010 0.152939
R21899 gnd.n3012 gnd.n3011 0.152939
R21900 gnd.n3012 gnd.n2640 0.152939
R21901 gnd.n3025 gnd.n2640 0.152939
R21902 gnd.n3026 gnd.n3025 0.152939
R21903 gnd.n3027 gnd.n3026 0.152939
R21904 gnd.n3027 gnd.n2632 0.152939
R21905 gnd.n3063 gnd.n2632 0.152939
R21906 gnd.n3063 gnd.n3062 0.152939
R21907 gnd.n3062 gnd.n3061 0.152939
R21908 gnd.n3061 gnd.n2633 0.152939
R21909 gnd.n3057 gnd.n2633 0.152939
R21910 gnd.n3057 gnd.n3056 0.152939
R21911 gnd.n3056 gnd.n3055 0.152939
R21912 gnd.n3055 gnd.n2637 0.152939
R21913 gnd.n3051 gnd.n2637 0.152939
R21914 gnd.n3051 gnd.n2613 0.152939
R21915 gnd.n3127 gnd.n2613 0.152939
R21916 gnd.n3128 gnd.n3127 0.152939
R21917 gnd.n3130 gnd.n3128 0.152939
R21918 gnd.n3130 gnd.n3129 0.152939
R21919 gnd.n3129 gnd.n2608 0.152939
R21920 gnd.n3144 gnd.n2608 0.152939
R21921 gnd.n3218 gnd.n2386 0.152939
R21922 gnd.n3218 gnd.n3217 0.152939
R21923 gnd.n3217 gnd.n3216 0.152939
R21924 gnd.n3216 gnd.n2415 0.152939
R21925 gnd.n3212 gnd.n2415 0.152939
R21926 gnd.n3212 gnd.n3211 0.152939
R21927 gnd.n3238 gnd.n3237 0.152939
R21928 gnd.n3240 gnd.n3238 0.152939
R21929 gnd.n3240 gnd.n3239 0.152939
R21930 gnd.n3239 gnd.n2362 0.152939
R21931 gnd.n3267 gnd.n2362 0.152939
R21932 gnd.n3268 gnd.n3267 0.152939
R21933 gnd.n3270 gnd.n3268 0.152939
R21934 gnd.n3270 gnd.n3269 0.152939
R21935 gnd.n3269 gnd.n2337 0.152939
R21936 gnd.n3303 gnd.n2337 0.152939
R21937 gnd.n3304 gnd.n3303 0.152939
R21938 gnd.n3315 gnd.n3304 0.152939
R21939 gnd.n3315 gnd.n3314 0.152939
R21940 gnd.n3314 gnd.n3313 0.152939
R21941 gnd.n3313 gnd.n3305 0.152939
R21942 gnd.n3309 gnd.n3305 0.152939
R21943 gnd.n3309 gnd.n1623 0.152939
R21944 gnd.n4823 gnd.n1623 0.152939
R21945 gnd.n4823 gnd.n4822 0.152939
R21946 gnd.n4822 gnd.n4821 0.152939
R21947 gnd.n4821 gnd.n1624 0.152939
R21948 gnd.n4817 gnd.n1624 0.152939
R21949 gnd.n4817 gnd.n4816 0.152939
R21950 gnd.n4816 gnd.n4815 0.152939
R21951 gnd.n4815 gnd.n1629 0.152939
R21952 gnd.n4811 gnd.n1629 0.152939
R21953 gnd.n4811 gnd.n4810 0.152939
R21954 gnd.n4810 gnd.n4809 0.152939
R21955 gnd.n4809 gnd.n1634 0.152939
R21956 gnd.n4805 gnd.n1634 0.152939
R21957 gnd.n4805 gnd.n4804 0.152939
R21958 gnd.n4804 gnd.n4803 0.152939
R21959 gnd.n4803 gnd.n1639 0.152939
R21960 gnd.n4799 gnd.n1639 0.152939
R21961 gnd.n4799 gnd.n4798 0.152939
R21962 gnd.n4798 gnd.n4797 0.152939
R21963 gnd.n4797 gnd.n1644 0.152939
R21964 gnd.n4793 gnd.n1644 0.152939
R21965 gnd.n4793 gnd.n4792 0.152939
R21966 gnd.n4792 gnd.n4791 0.152939
R21967 gnd.n4791 gnd.n1649 0.152939
R21968 gnd.n4787 gnd.n1649 0.152939
R21969 gnd.n4787 gnd.n4786 0.152939
R21970 gnd.n4786 gnd.n4785 0.152939
R21971 gnd.n4785 gnd.n1654 0.152939
R21972 gnd.n4781 gnd.n1654 0.152939
R21973 gnd.n4781 gnd.n4780 0.152939
R21974 gnd.n4780 gnd.n4779 0.152939
R21975 gnd.n4779 gnd.n1659 0.152939
R21976 gnd.n4775 gnd.n1659 0.152939
R21977 gnd.n4775 gnd.n4774 0.152939
R21978 gnd.n4774 gnd.n4773 0.152939
R21979 gnd.n4773 gnd.n1664 0.152939
R21980 gnd.n4769 gnd.n1664 0.152939
R21981 gnd.n4769 gnd.n4768 0.152939
R21982 gnd.n4768 gnd.n4767 0.152939
R21983 gnd.n4767 gnd.n1669 0.152939
R21984 gnd.n4763 gnd.n1669 0.152939
R21985 gnd.n4763 gnd.n4762 0.152939
R21986 gnd.n4762 gnd.n4761 0.152939
R21987 gnd.n4761 gnd.n1674 0.152939
R21988 gnd.n4757 gnd.n1674 0.152939
R21989 gnd.n4757 gnd.n4756 0.152939
R21990 gnd.n4756 gnd.n4755 0.152939
R21991 gnd.n4755 gnd.n1679 0.152939
R21992 gnd.n4751 gnd.n1679 0.152939
R21993 gnd.n4751 gnd.n4750 0.152939
R21994 gnd.n4750 gnd.n4749 0.152939
R21995 gnd.n4749 gnd.n1684 0.152939
R21996 gnd.n4745 gnd.n1684 0.152939
R21997 gnd.n4745 gnd.n4744 0.152939
R21998 gnd.n4744 gnd.n4743 0.152939
R21999 gnd.n4743 gnd.n1689 0.152939
R22000 gnd.n4739 gnd.n1689 0.152939
R22001 gnd.n4739 gnd.n4738 0.152939
R22002 gnd.n4738 gnd.n4737 0.152939
R22003 gnd.n4737 gnd.n1694 0.152939
R22004 gnd.n4733 gnd.n1694 0.152939
R22005 gnd.n4733 gnd.n4732 0.152939
R22006 gnd.n4732 gnd.n4731 0.152939
R22007 gnd.n4731 gnd.n1699 0.152939
R22008 gnd.n1702 gnd.n1699 0.152939
R22009 gnd.n3989 gnd.n3988 0.152939
R22010 gnd.n3989 gnd.n3984 0.152939
R22011 gnd.n3997 gnd.n3984 0.152939
R22012 gnd.n3998 gnd.n3997 0.152939
R22013 gnd.n4000 gnd.n3998 0.152939
R22014 gnd.n4000 gnd.n3999 0.152939
R22015 gnd.n3929 gnd.n3924 0.152939
R22016 gnd.n3924 gnd.n1929 0.152939
R22017 gnd.n4500 gnd.n1929 0.152939
R22018 gnd.n4501 gnd.n4500 0.152939
R22019 gnd.n4502 gnd.n4501 0.152939
R22020 gnd.n4502 gnd.n1892 0.152939
R22021 gnd.n4514 gnd.n1892 0.152939
R22022 gnd.n4515 gnd.n4514 0.152939
R22023 gnd.n4516 gnd.n4515 0.152939
R22024 gnd.n4516 gnd.n1883 0.152939
R22025 gnd.n4552 gnd.n1883 0.152939
R22026 gnd.n4552 gnd.n4551 0.152939
R22027 gnd.n4551 gnd.n4550 0.152939
R22028 gnd.n4550 gnd.n1884 0.152939
R22029 gnd.n4546 gnd.n1884 0.152939
R22030 gnd.n4546 gnd.n4545 0.152939
R22031 gnd.n4545 gnd.n4544 0.152939
R22032 gnd.n4544 gnd.n1888 0.152939
R22033 gnd.n4540 gnd.n1888 0.152939
R22034 gnd.n4540 gnd.n1865 0.152939
R22035 gnd.n4612 gnd.n1865 0.152939
R22036 gnd.n4613 gnd.n4612 0.152939
R22037 gnd.n4617 gnd.n4613 0.152939
R22038 gnd.n4617 gnd.n4616 0.152939
R22039 gnd.n4616 gnd.n4615 0.152939
R22040 gnd.n4615 gnd.n79 0.152939
R22041 gnd.n3211 gnd.n3210 0.128549
R22042 gnd.n3999 gnd.n1933 0.128549
R22043 gnd.n2984 gnd.n1360 0.10111
R22044 gnd.n4572 gnd.n95 0.10111
R22045 gnd.n6039 gnd.n6038 0.0767195
R22046 gnd.n6038 gnd.n6037 0.0767195
R22047 gnd.n7876 gnd.n93 0.0767195
R22048 gnd.n7876 gnd.n94 0.0767195
R22049 gnd.n5035 gnd.n1359 0.0767195
R22050 gnd.n5035 gnd.n1357 0.0767195
R22051 gnd.n7886 gnd.n7885 0.0695946
R22052 gnd.n2953 gnd.n2950 0.0695946
R22053 gnd.n2955 gnd.n2953 0.0695946
R22054 gnd.n7886 gnd.n79 0.0695946
R22055 gnd.n3210 gnd.n2532 0.063
R22056 gnd.n4489 gnd.n1933 0.063
R22057 gnd.n395 gnd.n95 0.0523293
R22058 gnd.n2917 gnd.n1360 0.0523293
R22059 gnd.n6543 gnd.n5271 0.0477147
R22060 gnd.n4491 gnd.n4489 0.0477147
R22061 gnd.n7694 gnd.n210 0.0477147
R22062 gnd.n5107 gnd.n5106 0.0477147
R22063 gnd.n2532 gnd.n1477 0.0477147
R22064 gnd.n5802 gnd.n5690 0.0442063
R22065 gnd.n5803 gnd.n5802 0.0442063
R22066 gnd.n5804 gnd.n5803 0.0442063
R22067 gnd.n5804 gnd.n5679 0.0442063
R22068 gnd.n5818 gnd.n5679 0.0442063
R22069 gnd.n5819 gnd.n5818 0.0442063
R22070 gnd.n5820 gnd.n5819 0.0442063
R22071 gnd.n5820 gnd.n5666 0.0442063
R22072 gnd.n5864 gnd.n5666 0.0442063
R22073 gnd.n5865 gnd.n5864 0.0442063
R22074 gnd.n5867 gnd.n5600 0.0344674
R22075 gnd.n4492 gnd.n4491 0.0344674
R22076 gnd.n4492 gnd.n1743 0.0344674
R22077 gnd.n1744 gnd.n1743 0.0344674
R22078 gnd.n1745 gnd.n1744 0.0344674
R22079 gnd.n1927 gnd.n1745 0.0344674
R22080 gnd.n1927 gnd.n1763 0.0344674
R22081 gnd.n1764 gnd.n1763 0.0344674
R22082 gnd.n1765 gnd.n1764 0.0344674
R22083 gnd.n1890 gnd.n1765 0.0344674
R22084 gnd.n1890 gnd.n1784 0.0344674
R22085 gnd.n1785 gnd.n1784 0.0344674
R22086 gnd.n1786 gnd.n1785 0.0344674
R22087 gnd.n4525 gnd.n1786 0.0344674
R22088 gnd.n4525 gnd.n1803 0.0344674
R22089 gnd.n1804 gnd.n1803 0.0344674
R22090 gnd.n1805 gnd.n1804 0.0344674
R22091 gnd.n4535 gnd.n1805 0.0344674
R22092 gnd.n4535 gnd.n1824 0.0344674
R22093 gnd.n1825 gnd.n1824 0.0344674
R22094 gnd.n1826 gnd.n1825 0.0344674
R22095 gnd.n4583 gnd.n1826 0.0344674
R22096 gnd.n4583 gnd.n1841 0.0344674
R22097 gnd.n1842 gnd.n1841 0.0344674
R22098 gnd.n1843 gnd.n1842 0.0344674
R22099 gnd.n4584 gnd.n1843 0.0344674
R22100 gnd.n4585 gnd.n4584 0.0344674
R22101 gnd.n4590 gnd.n4585 0.0344674
R22102 gnd.n4592 gnd.n4590 0.0344674
R22103 gnd.n4593 gnd.n4592 0.0344674
R22104 gnd.n4593 gnd.n389 0.0344674
R22105 gnd.n389 gnd.n109 0.0344674
R22106 gnd.n110 gnd.n109 0.0344674
R22107 gnd.n111 gnd.n110 0.0344674
R22108 gnd.n383 gnd.n111 0.0344674
R22109 gnd.n383 gnd.n127 0.0344674
R22110 gnd.n128 gnd.n127 0.0344674
R22111 gnd.n129 gnd.n128 0.0344674
R22112 gnd.n377 gnd.n129 0.0344674
R22113 gnd.n377 gnd.n148 0.0344674
R22114 gnd.n149 gnd.n148 0.0344674
R22115 gnd.n150 gnd.n149 0.0344674
R22116 gnd.n371 gnd.n150 0.0344674
R22117 gnd.n371 gnd.n167 0.0344674
R22118 gnd.n168 gnd.n167 0.0344674
R22119 gnd.n169 gnd.n168 0.0344674
R22120 gnd.n365 gnd.n169 0.0344674
R22121 gnd.n365 gnd.n188 0.0344674
R22122 gnd.n189 gnd.n188 0.0344674
R22123 gnd.n190 gnd.n189 0.0344674
R22124 gnd.n360 gnd.n190 0.0344674
R22125 gnd.n360 gnd.n208 0.0344674
R22126 gnd.n209 gnd.n208 0.0344674
R22127 gnd.n210 gnd.n209 0.0344674
R22128 gnd.n5106 gnd.n1239 0.0344674
R22129 gnd.n2777 gnd.n1239 0.0344674
R22130 gnd.n2777 gnd.n1264 0.0344674
R22131 gnd.n1265 gnd.n1264 0.0344674
R22132 gnd.n1266 gnd.n1265 0.0344674
R22133 gnd.n2792 gnd.n1266 0.0344674
R22134 gnd.n2792 gnd.n1284 0.0344674
R22135 gnd.n1285 gnd.n1284 0.0344674
R22136 gnd.n1286 gnd.n1285 0.0344674
R22137 gnd.n2850 gnd.n1286 0.0344674
R22138 gnd.n2850 gnd.n1305 0.0344674
R22139 gnd.n1306 gnd.n1305 0.0344674
R22140 gnd.n1307 gnd.n1306 0.0344674
R22141 gnd.n2866 gnd.n1307 0.0344674
R22142 gnd.n2866 gnd.n1325 0.0344674
R22143 gnd.n1326 gnd.n1325 0.0344674
R22144 gnd.n1327 gnd.n1326 0.0344674
R22145 gnd.n2869 gnd.n1327 0.0344674
R22146 gnd.n2869 gnd.n1346 0.0344674
R22147 gnd.n1347 gnd.n1346 0.0344674
R22148 gnd.n1348 gnd.n1347 0.0344674
R22149 gnd.n2687 gnd.n1348 0.0344674
R22150 gnd.n2687 gnd.n2686 0.0344674
R22151 gnd.n2938 gnd.n2686 0.0344674
R22152 gnd.n2939 gnd.n2938 0.0344674
R22153 gnd.n2939 gnd.n2671 0.0344674
R22154 gnd.n2671 gnd.n2667 0.0344674
R22155 gnd.n2668 gnd.n2667 0.0344674
R22156 gnd.n2967 gnd.n2668 0.0344674
R22157 gnd.n2967 gnd.n2669 0.0344674
R22158 gnd.n2669 gnd.n1375 0.0344674
R22159 gnd.n1376 gnd.n1375 0.0344674
R22160 gnd.n1377 gnd.n1376 0.0344674
R22161 gnd.n3019 gnd.n1377 0.0344674
R22162 gnd.n3019 gnd.n1394 0.0344674
R22163 gnd.n1395 gnd.n1394 0.0344674
R22164 gnd.n1396 gnd.n1395 0.0344674
R22165 gnd.n3034 gnd.n1396 0.0344674
R22166 gnd.n3034 gnd.n1414 0.0344674
R22167 gnd.n1415 gnd.n1414 0.0344674
R22168 gnd.n1416 gnd.n1415 0.0344674
R22169 gnd.n3041 gnd.n1416 0.0344674
R22170 gnd.n3041 gnd.n1434 0.0344674
R22171 gnd.n1435 gnd.n1434 0.0344674
R22172 gnd.n1436 gnd.n1435 0.0344674
R22173 gnd.n2616 gnd.n1436 0.0344674
R22174 gnd.n2616 gnd.n1454 0.0344674
R22175 gnd.n1455 gnd.n1454 0.0344674
R22176 gnd.n1456 gnd.n1455 0.0344674
R22177 gnd.n2611 gnd.n1456 0.0344674
R22178 gnd.n2611 gnd.n1475 0.0344674
R22179 gnd.n1476 gnd.n1475 0.0344674
R22180 gnd.n1477 gnd.n1476 0.0344674
R22181 gnd.n3209 gnd.n2533 0.0344674
R22182 gnd.n4009 gnd.n4008 0.0344674
R22183 gnd.n3157 gnd.n3145 0.029712
R22184 gnd.n3939 gnd.n3930 0.029712
R22185 gnd.n5887 gnd.n5886 0.0269946
R22186 gnd.n5889 gnd.n5888 0.0269946
R22187 gnd.n5595 gnd.n5593 0.0269946
R22188 gnd.n5899 gnd.n5897 0.0269946
R22189 gnd.n5898 gnd.n5574 0.0269946
R22190 gnd.n5918 gnd.n5917 0.0269946
R22191 gnd.n5920 gnd.n5919 0.0269946
R22192 gnd.n5569 gnd.n5568 0.0269946
R22193 gnd.n5930 gnd.n5564 0.0269946
R22194 gnd.n5929 gnd.n5566 0.0269946
R22195 gnd.n5565 gnd.n5547 0.0269946
R22196 gnd.n5950 gnd.n5548 0.0269946
R22197 gnd.n5949 gnd.n5549 0.0269946
R22198 gnd.n5983 gnd.n5524 0.0269946
R22199 gnd.n5985 gnd.n5984 0.0269946
R22200 gnd.n5986 gnd.n5471 0.0269946
R22201 gnd.n5519 gnd.n5472 0.0269946
R22202 gnd.n5521 gnd.n5473 0.0269946
R22203 gnd.n5996 gnd.n5995 0.0269946
R22204 gnd.n5998 gnd.n5997 0.0269946
R22205 gnd.n5999 gnd.n5493 0.0269946
R22206 gnd.n6001 gnd.n5494 0.0269946
R22207 gnd.n6004 gnd.n5495 0.0269946
R22208 gnd.n6007 gnd.n6006 0.0269946
R22209 gnd.n6009 gnd.n6008 0.0269946
R22210 gnd.n6074 gnd.n5378 0.0269946
R22211 gnd.n6076 gnd.n6075 0.0269946
R22212 gnd.n6085 gnd.n5371 0.0269946
R22213 gnd.n6087 gnd.n6086 0.0269946
R22214 gnd.n6088 gnd.n5369 0.0269946
R22215 gnd.n6095 gnd.n6091 0.0269946
R22216 gnd.n6094 gnd.n6093 0.0269946
R22217 gnd.n6092 gnd.n5348 0.0269946
R22218 gnd.n6119 gnd.n5349 0.0269946
R22219 gnd.n6118 gnd.n5350 0.0269946
R22220 gnd.n6115 gnd.n1044 0.0269946
R22221 gnd.n5326 gnd.n1045 0.0269946
R22222 gnd.n5328 gnd.n1046 0.0269946
R22223 gnd.n6171 gnd.n6170 0.0269946
R22224 gnd.n6173 gnd.n6172 0.0269946
R22225 gnd.n6174 gnd.n1067 0.0269946
R22226 gnd.n6176 gnd.n1068 0.0269946
R22227 gnd.n6178 gnd.n1069 0.0269946
R22228 gnd.n6184 gnd.n6183 0.0269946
R22229 gnd.n6186 gnd.n6185 0.0269946
R22230 gnd.n6187 gnd.n1092 0.0269946
R22231 gnd.n6188 gnd.n1093 0.0269946
R22232 gnd.n6189 gnd.n1094 0.0269946
R22233 gnd.n6449 gnd.n6448 0.0269946
R22234 gnd.n6450 gnd.n1118 0.0269946
R22235 gnd.n6451 gnd.n1119 0.0269946
R22236 gnd.n6452 gnd.n1120 0.0269946
R22237 gnd.n3205 gnd.n2539 0.0225788
R22238 gnd.n3204 gnd.n2540 0.0225788
R22239 gnd.n3201 gnd.n3200 0.0225788
R22240 gnd.n3197 gnd.n2546 0.0225788
R22241 gnd.n3196 gnd.n2552 0.0225788
R22242 gnd.n3193 gnd.n3192 0.0225788
R22243 gnd.n3189 gnd.n2558 0.0225788
R22244 gnd.n3188 gnd.n2562 0.0225788
R22245 gnd.n3185 gnd.n3184 0.0225788
R22246 gnd.n3181 gnd.n2569 0.0225788
R22247 gnd.n3180 gnd.n2575 0.0225788
R22248 gnd.n3177 gnd.n3176 0.0225788
R22249 gnd.n3173 gnd.n2581 0.0225788
R22250 gnd.n3172 gnd.n2585 0.0225788
R22251 gnd.n3169 gnd.n3168 0.0225788
R22252 gnd.n3165 gnd.n2592 0.0225788
R22253 gnd.n3164 gnd.n2599 0.0225788
R22254 gnd.n2607 gnd.n2605 0.0225788
R22255 gnd.n3158 gnd.n3157 0.0225788
R22256 gnd.n4015 gnd.n4013 0.0225788
R22257 gnd.n4014 gnd.n3976 0.0225788
R22258 gnd.n4024 gnd.n4023 0.0225788
R22259 gnd.n3977 gnd.n3972 0.0225788
R22260 gnd.n4034 gnd.n4032 0.0225788
R22261 gnd.n4033 gnd.n3967 0.0225788
R22262 gnd.n4043 gnd.n4042 0.0225788
R22263 gnd.n3968 gnd.n3963 0.0225788
R22264 gnd.n4053 gnd.n4051 0.0225788
R22265 gnd.n4052 gnd.n3958 0.0225788
R22266 gnd.n4062 gnd.n4061 0.0225788
R22267 gnd.n3959 gnd.n3954 0.0225788
R22268 gnd.n4072 gnd.n4070 0.0225788
R22269 gnd.n4071 gnd.n3949 0.0225788
R22270 gnd.n4082 gnd.n4081 0.0225788
R22271 gnd.n4078 gnd.n3950 0.0225788
R22272 gnd.n4092 gnd.n3937 0.0225788
R22273 gnd.n4091 gnd.n3938 0.0225788
R22274 gnd.n3940 gnd.n3939 0.0225788
R22275 gnd.n4101 gnd.n3930 0.0218415
R22276 gnd.n3154 gnd.n3145 0.0218415
R22277 gnd.n5867 gnd.n5866 0.0202011
R22278 gnd.n5866 gnd.n5865 0.0148637
R22279 gnd.n6446 gnd.n6190 0.0144266
R22280 gnd.n6447 gnd.n6446 0.0130679
R22281 gnd.n2539 gnd.n2533 0.0123886
R22282 gnd.n3205 gnd.n3204 0.0123886
R22283 gnd.n3201 gnd.n2540 0.0123886
R22284 gnd.n3200 gnd.n2546 0.0123886
R22285 gnd.n3197 gnd.n3196 0.0123886
R22286 gnd.n3193 gnd.n2552 0.0123886
R22287 gnd.n3192 gnd.n2558 0.0123886
R22288 gnd.n3189 gnd.n3188 0.0123886
R22289 gnd.n3185 gnd.n2562 0.0123886
R22290 gnd.n3184 gnd.n2569 0.0123886
R22291 gnd.n3181 gnd.n3180 0.0123886
R22292 gnd.n3177 gnd.n2575 0.0123886
R22293 gnd.n3176 gnd.n2581 0.0123886
R22294 gnd.n3173 gnd.n3172 0.0123886
R22295 gnd.n3169 gnd.n2585 0.0123886
R22296 gnd.n3168 gnd.n2592 0.0123886
R22297 gnd.n3165 gnd.n3164 0.0123886
R22298 gnd.n2605 gnd.n2599 0.0123886
R22299 gnd.n3158 gnd.n2607 0.0123886
R22300 gnd.n4013 gnd.n4009 0.0123886
R22301 gnd.n4015 gnd.n4014 0.0123886
R22302 gnd.n4024 gnd.n3976 0.0123886
R22303 gnd.n4023 gnd.n3977 0.0123886
R22304 gnd.n4032 gnd.n3972 0.0123886
R22305 gnd.n4034 gnd.n4033 0.0123886
R22306 gnd.n4043 gnd.n3967 0.0123886
R22307 gnd.n4042 gnd.n3968 0.0123886
R22308 gnd.n4051 gnd.n3963 0.0123886
R22309 gnd.n4053 gnd.n4052 0.0123886
R22310 gnd.n4062 gnd.n3958 0.0123886
R22311 gnd.n4061 gnd.n3959 0.0123886
R22312 gnd.n4070 gnd.n3954 0.0123886
R22313 gnd.n4072 gnd.n4071 0.0123886
R22314 gnd.n4082 gnd.n3949 0.0123886
R22315 gnd.n4081 gnd.n3950 0.0123886
R22316 gnd.n4078 gnd.n3937 0.0123886
R22317 gnd.n4092 gnd.n4091 0.0123886
R22318 gnd.n3940 gnd.n3938 0.0123886
R22319 gnd.n5886 gnd.n5600 0.00797283
R22320 gnd.n5888 gnd.n5887 0.00797283
R22321 gnd.n5889 gnd.n5595 0.00797283
R22322 gnd.n5897 gnd.n5593 0.00797283
R22323 gnd.n5899 gnd.n5898 0.00797283
R22324 gnd.n5917 gnd.n5574 0.00797283
R22325 gnd.n5919 gnd.n5918 0.00797283
R22326 gnd.n5920 gnd.n5569 0.00797283
R22327 gnd.n5568 gnd.n5564 0.00797283
R22328 gnd.n5930 gnd.n5929 0.00797283
R22329 gnd.n5566 gnd.n5565 0.00797283
R22330 gnd.n5548 gnd.n5547 0.00797283
R22331 gnd.n5950 gnd.n5949 0.00797283
R22332 gnd.n5549 gnd.n5524 0.00797283
R22333 gnd.n5984 gnd.n5983 0.00797283
R22334 gnd.n5986 gnd.n5985 0.00797283
R22335 gnd.n5519 gnd.n5471 0.00797283
R22336 gnd.n5521 gnd.n5472 0.00797283
R22337 gnd.n5995 gnd.n5473 0.00797283
R22338 gnd.n5997 gnd.n5996 0.00797283
R22339 gnd.n5999 gnd.n5998 0.00797283
R22340 gnd.n6001 gnd.n5493 0.00797283
R22341 gnd.n6004 gnd.n5494 0.00797283
R22342 gnd.n6006 gnd.n5495 0.00797283
R22343 gnd.n6009 gnd.n6007 0.00797283
R22344 gnd.n6008 gnd.n5378 0.00797283
R22345 gnd.n6076 gnd.n6074 0.00797283
R22346 gnd.n6075 gnd.n5371 0.00797283
R22347 gnd.n6086 gnd.n6085 0.00797283
R22348 gnd.n6088 gnd.n6087 0.00797283
R22349 gnd.n6091 gnd.n5369 0.00797283
R22350 gnd.n6095 gnd.n6094 0.00797283
R22351 gnd.n6093 gnd.n6092 0.00797283
R22352 gnd.n5349 gnd.n5348 0.00797283
R22353 gnd.n6119 gnd.n6118 0.00797283
R22354 gnd.n6115 gnd.n5350 0.00797283
R22355 gnd.n5326 gnd.n1044 0.00797283
R22356 gnd.n5328 gnd.n1045 0.00797283
R22357 gnd.n6170 gnd.n1046 0.00797283
R22358 gnd.n6172 gnd.n6171 0.00797283
R22359 gnd.n6174 gnd.n6173 0.00797283
R22360 gnd.n6176 gnd.n1067 0.00797283
R22361 gnd.n6178 gnd.n1068 0.00797283
R22362 gnd.n6183 gnd.n1069 0.00797283
R22363 gnd.n6185 gnd.n6184 0.00797283
R22364 gnd.n6187 gnd.n6186 0.00797283
R22365 gnd.n6188 gnd.n1092 0.00797283
R22366 gnd.n6189 gnd.n1093 0.00797283
R22367 gnd.n6190 gnd.n1094 0.00797283
R22368 gnd.n6448 gnd.n6447 0.00797283
R22369 gnd.n6450 gnd.n6449 0.00797283
R22370 gnd.n6451 gnd.n1118 0.00797283
R22371 gnd.n6452 gnd.n1119 0.00797283
R22372 gnd.n5271 gnd.n1120 0.00797283
R22373 gnd.n3210 gnd.n3209 0.00593478
R22374 gnd.n4008 gnd.n1933 0.00593478
R22375 CSoutput.n19 CSoutput.t216 184.661
R22376 CSoutput.n78 CSoutput.n77 165.8
R22377 CSoutput.n76 CSoutput.n0 165.8
R22378 CSoutput.n75 CSoutput.n74 165.8
R22379 CSoutput.n73 CSoutput.n72 165.8
R22380 CSoutput.n71 CSoutput.n2 165.8
R22381 CSoutput.n69 CSoutput.n68 165.8
R22382 CSoutput.n67 CSoutput.n3 165.8
R22383 CSoutput.n66 CSoutput.n65 165.8
R22384 CSoutput.n63 CSoutput.n4 165.8
R22385 CSoutput.n61 CSoutput.n60 165.8
R22386 CSoutput.n59 CSoutput.n5 165.8
R22387 CSoutput.n58 CSoutput.n57 165.8
R22388 CSoutput.n55 CSoutput.n6 165.8
R22389 CSoutput.n54 CSoutput.n53 165.8
R22390 CSoutput.n52 CSoutput.n51 165.8
R22391 CSoutput.n50 CSoutput.n8 165.8
R22392 CSoutput.n48 CSoutput.n47 165.8
R22393 CSoutput.n46 CSoutput.n9 165.8
R22394 CSoutput.n45 CSoutput.n44 165.8
R22395 CSoutput.n42 CSoutput.n10 165.8
R22396 CSoutput.n41 CSoutput.n40 165.8
R22397 CSoutput.n39 CSoutput.n38 165.8
R22398 CSoutput.n37 CSoutput.n12 165.8
R22399 CSoutput.n35 CSoutput.n34 165.8
R22400 CSoutput.n33 CSoutput.n13 165.8
R22401 CSoutput.n32 CSoutput.n31 165.8
R22402 CSoutput.n29 CSoutput.n14 165.8
R22403 CSoutput.n28 CSoutput.n27 165.8
R22404 CSoutput.n26 CSoutput.n25 165.8
R22405 CSoutput.n24 CSoutput.n16 165.8
R22406 CSoutput.n22 CSoutput.n21 165.8
R22407 CSoutput.n20 CSoutput.n17 165.8
R22408 CSoutput.n77 CSoutput.t218 162.194
R22409 CSoutput.n18 CSoutput.t225 120.501
R22410 CSoutput.n23 CSoutput.t227 120.501
R22411 CSoutput.n15 CSoutput.t220 120.501
R22412 CSoutput.n30 CSoutput.t237 120.501
R22413 CSoutput.n36 CSoutput.t228 120.501
R22414 CSoutput.n11 CSoutput.t223 120.501
R22415 CSoutput.n43 CSoutput.t217 120.501
R22416 CSoutput.n49 CSoutput.t234 120.501
R22417 CSoutput.n7 CSoutput.t231 120.501
R22418 CSoutput.n56 CSoutput.t221 120.501
R22419 CSoutput.n62 CSoutput.t236 120.501
R22420 CSoutput.n64 CSoutput.t232 120.501
R22421 CSoutput.n70 CSoutput.t224 120.501
R22422 CSoutput.n1 CSoutput.t226 120.501
R22423 CSoutput.n330 CSoutput.n328 103.469
R22424 CSoutput.n310 CSoutput.n308 103.469
R22425 CSoutput.n291 CSoutput.n289 103.469
R22426 CSoutput.n120 CSoutput.n118 103.469
R22427 CSoutput.n100 CSoutput.n98 103.469
R22428 CSoutput.n81 CSoutput.n79 103.469
R22429 CSoutput.n344 CSoutput.n343 103.111
R22430 CSoutput.n342 CSoutput.n341 103.111
R22431 CSoutput.n340 CSoutput.n339 103.111
R22432 CSoutput.n338 CSoutput.n337 103.111
R22433 CSoutput.n336 CSoutput.n335 103.111
R22434 CSoutput.n334 CSoutput.n333 103.111
R22435 CSoutput.n332 CSoutput.n331 103.111
R22436 CSoutput.n330 CSoutput.n329 103.111
R22437 CSoutput.n326 CSoutput.n325 103.111
R22438 CSoutput.n324 CSoutput.n323 103.111
R22439 CSoutput.n322 CSoutput.n321 103.111
R22440 CSoutput.n320 CSoutput.n319 103.111
R22441 CSoutput.n318 CSoutput.n317 103.111
R22442 CSoutput.n316 CSoutput.n315 103.111
R22443 CSoutput.n314 CSoutput.n313 103.111
R22444 CSoutput.n312 CSoutput.n311 103.111
R22445 CSoutput.n310 CSoutput.n309 103.111
R22446 CSoutput.n307 CSoutput.n306 103.111
R22447 CSoutput.n305 CSoutput.n304 103.111
R22448 CSoutput.n303 CSoutput.n302 103.111
R22449 CSoutput.n301 CSoutput.n300 103.111
R22450 CSoutput.n299 CSoutput.n298 103.111
R22451 CSoutput.n297 CSoutput.n296 103.111
R22452 CSoutput.n295 CSoutput.n294 103.111
R22453 CSoutput.n293 CSoutput.n292 103.111
R22454 CSoutput.n291 CSoutput.n290 103.111
R22455 CSoutput.n120 CSoutput.n119 103.111
R22456 CSoutput.n122 CSoutput.n121 103.111
R22457 CSoutput.n124 CSoutput.n123 103.111
R22458 CSoutput.n126 CSoutput.n125 103.111
R22459 CSoutput.n128 CSoutput.n127 103.111
R22460 CSoutput.n130 CSoutput.n129 103.111
R22461 CSoutput.n132 CSoutput.n131 103.111
R22462 CSoutput.n134 CSoutput.n133 103.111
R22463 CSoutput.n136 CSoutput.n135 103.111
R22464 CSoutput.n100 CSoutput.n99 103.111
R22465 CSoutput.n102 CSoutput.n101 103.111
R22466 CSoutput.n104 CSoutput.n103 103.111
R22467 CSoutput.n106 CSoutput.n105 103.111
R22468 CSoutput.n108 CSoutput.n107 103.111
R22469 CSoutput.n110 CSoutput.n109 103.111
R22470 CSoutput.n112 CSoutput.n111 103.111
R22471 CSoutput.n114 CSoutput.n113 103.111
R22472 CSoutput.n116 CSoutput.n115 103.111
R22473 CSoutput.n81 CSoutput.n80 103.111
R22474 CSoutput.n83 CSoutput.n82 103.111
R22475 CSoutput.n85 CSoutput.n84 103.111
R22476 CSoutput.n87 CSoutput.n86 103.111
R22477 CSoutput.n89 CSoutput.n88 103.111
R22478 CSoutput.n91 CSoutput.n90 103.111
R22479 CSoutput.n93 CSoutput.n92 103.111
R22480 CSoutput.n95 CSoutput.n94 103.111
R22481 CSoutput.n97 CSoutput.n96 103.111
R22482 CSoutput.n346 CSoutput.n345 103.111
R22483 CSoutput.n382 CSoutput.n380 81.5057
R22484 CSoutput.n366 CSoutput.n364 81.5057
R22485 CSoutput.n351 CSoutput.n349 81.5057
R22486 CSoutput.n430 CSoutput.n428 81.5057
R22487 CSoutput.n414 CSoutput.n412 81.5057
R22488 CSoutput.n399 CSoutput.n397 81.5057
R22489 CSoutput.n394 CSoutput.n393 80.9324
R22490 CSoutput.n392 CSoutput.n391 80.9324
R22491 CSoutput.n390 CSoutput.n389 80.9324
R22492 CSoutput.n388 CSoutput.n387 80.9324
R22493 CSoutput.n386 CSoutput.n385 80.9324
R22494 CSoutput.n384 CSoutput.n383 80.9324
R22495 CSoutput.n382 CSoutput.n381 80.9324
R22496 CSoutput.n378 CSoutput.n377 80.9324
R22497 CSoutput.n376 CSoutput.n375 80.9324
R22498 CSoutput.n374 CSoutput.n373 80.9324
R22499 CSoutput.n372 CSoutput.n371 80.9324
R22500 CSoutput.n370 CSoutput.n369 80.9324
R22501 CSoutput.n368 CSoutput.n367 80.9324
R22502 CSoutput.n366 CSoutput.n365 80.9324
R22503 CSoutput.n363 CSoutput.n362 80.9324
R22504 CSoutput.n361 CSoutput.n360 80.9324
R22505 CSoutput.n359 CSoutput.n358 80.9324
R22506 CSoutput.n357 CSoutput.n356 80.9324
R22507 CSoutput.n355 CSoutput.n354 80.9324
R22508 CSoutput.n353 CSoutput.n352 80.9324
R22509 CSoutput.n351 CSoutput.n350 80.9324
R22510 CSoutput.n430 CSoutput.n429 80.9324
R22511 CSoutput.n432 CSoutput.n431 80.9324
R22512 CSoutput.n434 CSoutput.n433 80.9324
R22513 CSoutput.n436 CSoutput.n435 80.9324
R22514 CSoutput.n438 CSoutput.n437 80.9324
R22515 CSoutput.n440 CSoutput.n439 80.9324
R22516 CSoutput.n442 CSoutput.n441 80.9324
R22517 CSoutput.n414 CSoutput.n413 80.9324
R22518 CSoutput.n416 CSoutput.n415 80.9324
R22519 CSoutput.n418 CSoutput.n417 80.9324
R22520 CSoutput.n420 CSoutput.n419 80.9324
R22521 CSoutput.n422 CSoutput.n421 80.9324
R22522 CSoutput.n424 CSoutput.n423 80.9324
R22523 CSoutput.n426 CSoutput.n425 80.9324
R22524 CSoutput.n399 CSoutput.n398 80.9324
R22525 CSoutput.n401 CSoutput.n400 80.9324
R22526 CSoutput.n403 CSoutput.n402 80.9324
R22527 CSoutput.n405 CSoutput.n404 80.9324
R22528 CSoutput.n407 CSoutput.n406 80.9324
R22529 CSoutput.n409 CSoutput.n408 80.9324
R22530 CSoutput.n411 CSoutput.n410 80.9324
R22531 CSoutput.n25 CSoutput.n24 48.1486
R22532 CSoutput.n69 CSoutput.n3 48.1486
R22533 CSoutput.n38 CSoutput.n37 48.1486
R22534 CSoutput.n42 CSoutput.n41 48.1486
R22535 CSoutput.n51 CSoutput.n50 48.1486
R22536 CSoutput.n55 CSoutput.n54 48.1486
R22537 CSoutput.n22 CSoutput.n17 46.462
R22538 CSoutput.n72 CSoutput.n71 46.462
R22539 CSoutput.n20 CSoutput.n19 44.9055
R22540 CSoutput.n29 CSoutput.n28 43.7635
R22541 CSoutput.n65 CSoutput.n63 43.7635
R22542 CSoutput.n35 CSoutput.n13 41.7396
R22543 CSoutput.n57 CSoutput.n5 41.7396
R22544 CSoutput.n44 CSoutput.n9 37.0171
R22545 CSoutput.n48 CSoutput.n9 37.0171
R22546 CSoutput.n76 CSoutput.n75 34.9932
R22547 CSoutput.n31 CSoutput.n13 32.2947
R22548 CSoutput.n61 CSoutput.n5 32.2947
R22549 CSoutput.n30 CSoutput.n29 29.6014
R22550 CSoutput.n63 CSoutput.n62 29.6014
R22551 CSoutput.n19 CSoutput.n18 28.4085
R22552 CSoutput.n18 CSoutput.n17 25.1176
R22553 CSoutput.n72 CSoutput.n1 25.1176
R22554 CSoutput.n43 CSoutput.n42 22.0922
R22555 CSoutput.n50 CSoutput.n49 22.0922
R22556 CSoutput.n77 CSoutput.n76 21.8586
R22557 CSoutput.n37 CSoutput.n36 18.9681
R22558 CSoutput.n56 CSoutput.n55 18.9681
R22559 CSoutput.n25 CSoutput.n15 17.6292
R22560 CSoutput.n64 CSoutput.n3 17.6292
R22561 CSoutput.n24 CSoutput.n23 15.844
R22562 CSoutput.n70 CSoutput.n69 15.844
R22563 CSoutput.n38 CSoutput.n11 14.5051
R22564 CSoutput.n54 CSoutput.n7 14.5051
R22565 CSoutput.n445 CSoutput.n78 11.4967
R22566 CSoutput.n41 CSoutput.n11 11.3811
R22567 CSoutput.n51 CSoutput.n7 11.3811
R22568 CSoutput.n23 CSoutput.n22 10.0422
R22569 CSoutput.n71 CSoutput.n70 10.0422
R22570 CSoutput.n327 CSoutput.n307 9.25285
R22571 CSoutput.n117 CSoutput.n97 9.25285
R22572 CSoutput.n379 CSoutput.n363 8.98182
R22573 CSoutput.n427 CSoutput.n411 8.98182
R22574 CSoutput.n396 CSoutput.n348 8.55073
R22575 CSoutput.n28 CSoutput.n15 8.25698
R22576 CSoutput.n65 CSoutput.n64 8.25698
R22577 CSoutput.n348 CSoutput.n347 7.12641
R22578 CSoutput.n138 CSoutput.n137 7.12641
R22579 CSoutput.n36 CSoutput.n35 6.91809
R22580 CSoutput.n57 CSoutput.n56 6.91809
R22581 CSoutput.n396 CSoutput.n395 6.02792
R22582 CSoutput.n444 CSoutput.n443 6.02792
R22583 CSoutput.n395 CSoutput.n394 5.25266
R22584 CSoutput.n379 CSoutput.n378 5.25266
R22585 CSoutput.n443 CSoutput.n442 5.25266
R22586 CSoutput.n427 CSoutput.n426 5.25266
R22587 CSoutput.n347 CSoutput.n346 5.1449
R22588 CSoutput.n327 CSoutput.n326 5.1449
R22589 CSoutput.n137 CSoutput.n136 5.1449
R22590 CSoutput.n117 CSoutput.n116 5.1449
R22591 CSoutput.n445 CSoutput.n138 4.91834
R22592 CSoutput.n229 CSoutput.n182 4.5005
R22593 CSoutput.n198 CSoutput.n182 4.5005
R22594 CSoutput.n193 CSoutput.n177 4.5005
R22595 CSoutput.n193 CSoutput.n179 4.5005
R22596 CSoutput.n193 CSoutput.n176 4.5005
R22597 CSoutput.n193 CSoutput.n180 4.5005
R22598 CSoutput.n193 CSoutput.n175 4.5005
R22599 CSoutput.n193 CSoutput.t222 4.5005
R22600 CSoutput.n193 CSoutput.n174 4.5005
R22601 CSoutput.n193 CSoutput.n181 4.5005
R22602 CSoutput.n193 CSoutput.n182 4.5005
R22603 CSoutput.n191 CSoutput.n177 4.5005
R22604 CSoutput.n191 CSoutput.n179 4.5005
R22605 CSoutput.n191 CSoutput.n176 4.5005
R22606 CSoutput.n191 CSoutput.n180 4.5005
R22607 CSoutput.n191 CSoutput.n175 4.5005
R22608 CSoutput.n191 CSoutput.t222 4.5005
R22609 CSoutput.n191 CSoutput.n174 4.5005
R22610 CSoutput.n191 CSoutput.n181 4.5005
R22611 CSoutput.n191 CSoutput.n182 4.5005
R22612 CSoutput.n190 CSoutput.n177 4.5005
R22613 CSoutput.n190 CSoutput.n179 4.5005
R22614 CSoutput.n190 CSoutput.n176 4.5005
R22615 CSoutput.n190 CSoutput.n180 4.5005
R22616 CSoutput.n190 CSoutput.n175 4.5005
R22617 CSoutput.n190 CSoutput.t222 4.5005
R22618 CSoutput.n190 CSoutput.n174 4.5005
R22619 CSoutput.n190 CSoutput.n181 4.5005
R22620 CSoutput.n190 CSoutput.n182 4.5005
R22621 CSoutput.n275 CSoutput.n177 4.5005
R22622 CSoutput.n275 CSoutput.n179 4.5005
R22623 CSoutput.n275 CSoutput.n176 4.5005
R22624 CSoutput.n275 CSoutput.n180 4.5005
R22625 CSoutput.n275 CSoutput.n175 4.5005
R22626 CSoutput.n275 CSoutput.t222 4.5005
R22627 CSoutput.n275 CSoutput.n174 4.5005
R22628 CSoutput.n275 CSoutput.n181 4.5005
R22629 CSoutput.n275 CSoutput.n182 4.5005
R22630 CSoutput.n273 CSoutput.n177 4.5005
R22631 CSoutput.n273 CSoutput.n179 4.5005
R22632 CSoutput.n273 CSoutput.n176 4.5005
R22633 CSoutput.n273 CSoutput.n180 4.5005
R22634 CSoutput.n273 CSoutput.n175 4.5005
R22635 CSoutput.n273 CSoutput.t222 4.5005
R22636 CSoutput.n273 CSoutput.n174 4.5005
R22637 CSoutput.n273 CSoutput.n181 4.5005
R22638 CSoutput.n271 CSoutput.n177 4.5005
R22639 CSoutput.n271 CSoutput.n179 4.5005
R22640 CSoutput.n271 CSoutput.n176 4.5005
R22641 CSoutput.n271 CSoutput.n180 4.5005
R22642 CSoutput.n271 CSoutput.n175 4.5005
R22643 CSoutput.n271 CSoutput.t222 4.5005
R22644 CSoutput.n271 CSoutput.n174 4.5005
R22645 CSoutput.n271 CSoutput.n181 4.5005
R22646 CSoutput.n201 CSoutput.n177 4.5005
R22647 CSoutput.n201 CSoutput.n179 4.5005
R22648 CSoutput.n201 CSoutput.n176 4.5005
R22649 CSoutput.n201 CSoutput.n180 4.5005
R22650 CSoutput.n201 CSoutput.n175 4.5005
R22651 CSoutput.n201 CSoutput.t222 4.5005
R22652 CSoutput.n201 CSoutput.n174 4.5005
R22653 CSoutput.n201 CSoutput.n181 4.5005
R22654 CSoutput.n201 CSoutput.n182 4.5005
R22655 CSoutput.n200 CSoutput.n177 4.5005
R22656 CSoutput.n200 CSoutput.n179 4.5005
R22657 CSoutput.n200 CSoutput.n176 4.5005
R22658 CSoutput.n200 CSoutput.n180 4.5005
R22659 CSoutput.n200 CSoutput.n175 4.5005
R22660 CSoutput.n200 CSoutput.t222 4.5005
R22661 CSoutput.n200 CSoutput.n174 4.5005
R22662 CSoutput.n200 CSoutput.n181 4.5005
R22663 CSoutput.n200 CSoutput.n182 4.5005
R22664 CSoutput.n204 CSoutput.n177 4.5005
R22665 CSoutput.n204 CSoutput.n179 4.5005
R22666 CSoutput.n204 CSoutput.n176 4.5005
R22667 CSoutput.n204 CSoutput.n180 4.5005
R22668 CSoutput.n204 CSoutput.n175 4.5005
R22669 CSoutput.n204 CSoutput.t222 4.5005
R22670 CSoutput.n204 CSoutput.n174 4.5005
R22671 CSoutput.n204 CSoutput.n181 4.5005
R22672 CSoutput.n204 CSoutput.n182 4.5005
R22673 CSoutput.n203 CSoutput.n177 4.5005
R22674 CSoutput.n203 CSoutput.n179 4.5005
R22675 CSoutput.n203 CSoutput.n176 4.5005
R22676 CSoutput.n203 CSoutput.n180 4.5005
R22677 CSoutput.n203 CSoutput.n175 4.5005
R22678 CSoutput.n203 CSoutput.t222 4.5005
R22679 CSoutput.n203 CSoutput.n174 4.5005
R22680 CSoutput.n203 CSoutput.n181 4.5005
R22681 CSoutput.n203 CSoutput.n182 4.5005
R22682 CSoutput.n186 CSoutput.n177 4.5005
R22683 CSoutput.n186 CSoutput.n179 4.5005
R22684 CSoutput.n186 CSoutput.n176 4.5005
R22685 CSoutput.n186 CSoutput.n180 4.5005
R22686 CSoutput.n186 CSoutput.n175 4.5005
R22687 CSoutput.n186 CSoutput.t222 4.5005
R22688 CSoutput.n186 CSoutput.n174 4.5005
R22689 CSoutput.n186 CSoutput.n181 4.5005
R22690 CSoutput.n186 CSoutput.n182 4.5005
R22691 CSoutput.n278 CSoutput.n177 4.5005
R22692 CSoutput.n278 CSoutput.n179 4.5005
R22693 CSoutput.n278 CSoutput.n176 4.5005
R22694 CSoutput.n278 CSoutput.n180 4.5005
R22695 CSoutput.n278 CSoutput.n175 4.5005
R22696 CSoutput.n278 CSoutput.t222 4.5005
R22697 CSoutput.n278 CSoutput.n174 4.5005
R22698 CSoutput.n278 CSoutput.n181 4.5005
R22699 CSoutput.n278 CSoutput.n182 4.5005
R22700 CSoutput.n265 CSoutput.n236 4.5005
R22701 CSoutput.n265 CSoutput.n242 4.5005
R22702 CSoutput.n223 CSoutput.n212 4.5005
R22703 CSoutput.n223 CSoutput.n214 4.5005
R22704 CSoutput.n223 CSoutput.n211 4.5005
R22705 CSoutput.n223 CSoutput.n215 4.5005
R22706 CSoutput.n223 CSoutput.n210 4.5005
R22707 CSoutput.n223 CSoutput.t230 4.5005
R22708 CSoutput.n223 CSoutput.n209 4.5005
R22709 CSoutput.n223 CSoutput.n216 4.5005
R22710 CSoutput.n265 CSoutput.n223 4.5005
R22711 CSoutput.n244 CSoutput.n212 4.5005
R22712 CSoutput.n244 CSoutput.n214 4.5005
R22713 CSoutput.n244 CSoutput.n211 4.5005
R22714 CSoutput.n244 CSoutput.n215 4.5005
R22715 CSoutput.n244 CSoutput.n210 4.5005
R22716 CSoutput.n244 CSoutput.t230 4.5005
R22717 CSoutput.n244 CSoutput.n209 4.5005
R22718 CSoutput.n244 CSoutput.n216 4.5005
R22719 CSoutput.n265 CSoutput.n244 4.5005
R22720 CSoutput.n222 CSoutput.n212 4.5005
R22721 CSoutput.n222 CSoutput.n214 4.5005
R22722 CSoutput.n222 CSoutput.n211 4.5005
R22723 CSoutput.n222 CSoutput.n215 4.5005
R22724 CSoutput.n222 CSoutput.n210 4.5005
R22725 CSoutput.n222 CSoutput.t230 4.5005
R22726 CSoutput.n222 CSoutput.n209 4.5005
R22727 CSoutput.n222 CSoutput.n216 4.5005
R22728 CSoutput.n265 CSoutput.n222 4.5005
R22729 CSoutput.n246 CSoutput.n212 4.5005
R22730 CSoutput.n246 CSoutput.n214 4.5005
R22731 CSoutput.n246 CSoutput.n211 4.5005
R22732 CSoutput.n246 CSoutput.n215 4.5005
R22733 CSoutput.n246 CSoutput.n210 4.5005
R22734 CSoutput.n246 CSoutput.t230 4.5005
R22735 CSoutput.n246 CSoutput.n209 4.5005
R22736 CSoutput.n246 CSoutput.n216 4.5005
R22737 CSoutput.n265 CSoutput.n246 4.5005
R22738 CSoutput.n212 CSoutput.n207 4.5005
R22739 CSoutput.n214 CSoutput.n207 4.5005
R22740 CSoutput.n211 CSoutput.n207 4.5005
R22741 CSoutput.n215 CSoutput.n207 4.5005
R22742 CSoutput.n210 CSoutput.n207 4.5005
R22743 CSoutput.t230 CSoutput.n207 4.5005
R22744 CSoutput.n209 CSoutput.n207 4.5005
R22745 CSoutput.n216 CSoutput.n207 4.5005
R22746 CSoutput.n268 CSoutput.n212 4.5005
R22747 CSoutput.n268 CSoutput.n214 4.5005
R22748 CSoutput.n268 CSoutput.n211 4.5005
R22749 CSoutput.n268 CSoutput.n215 4.5005
R22750 CSoutput.n268 CSoutput.n210 4.5005
R22751 CSoutput.n268 CSoutput.t230 4.5005
R22752 CSoutput.n268 CSoutput.n209 4.5005
R22753 CSoutput.n268 CSoutput.n216 4.5005
R22754 CSoutput.n266 CSoutput.n212 4.5005
R22755 CSoutput.n266 CSoutput.n214 4.5005
R22756 CSoutput.n266 CSoutput.n211 4.5005
R22757 CSoutput.n266 CSoutput.n215 4.5005
R22758 CSoutput.n266 CSoutput.n210 4.5005
R22759 CSoutput.n266 CSoutput.t230 4.5005
R22760 CSoutput.n266 CSoutput.n209 4.5005
R22761 CSoutput.n266 CSoutput.n216 4.5005
R22762 CSoutput.n266 CSoutput.n265 4.5005
R22763 CSoutput.n248 CSoutput.n212 4.5005
R22764 CSoutput.n248 CSoutput.n214 4.5005
R22765 CSoutput.n248 CSoutput.n211 4.5005
R22766 CSoutput.n248 CSoutput.n215 4.5005
R22767 CSoutput.n248 CSoutput.n210 4.5005
R22768 CSoutput.n248 CSoutput.t230 4.5005
R22769 CSoutput.n248 CSoutput.n209 4.5005
R22770 CSoutput.n248 CSoutput.n216 4.5005
R22771 CSoutput.n265 CSoutput.n248 4.5005
R22772 CSoutput.n220 CSoutput.n212 4.5005
R22773 CSoutput.n220 CSoutput.n214 4.5005
R22774 CSoutput.n220 CSoutput.n211 4.5005
R22775 CSoutput.n220 CSoutput.n215 4.5005
R22776 CSoutput.n220 CSoutput.n210 4.5005
R22777 CSoutput.n220 CSoutput.t230 4.5005
R22778 CSoutput.n220 CSoutput.n209 4.5005
R22779 CSoutput.n220 CSoutput.n216 4.5005
R22780 CSoutput.n265 CSoutput.n220 4.5005
R22781 CSoutput.n250 CSoutput.n212 4.5005
R22782 CSoutput.n250 CSoutput.n214 4.5005
R22783 CSoutput.n250 CSoutput.n211 4.5005
R22784 CSoutput.n250 CSoutput.n215 4.5005
R22785 CSoutput.n250 CSoutput.n210 4.5005
R22786 CSoutput.n250 CSoutput.t230 4.5005
R22787 CSoutput.n250 CSoutput.n209 4.5005
R22788 CSoutput.n250 CSoutput.n216 4.5005
R22789 CSoutput.n265 CSoutput.n250 4.5005
R22790 CSoutput.n219 CSoutput.n212 4.5005
R22791 CSoutput.n219 CSoutput.n214 4.5005
R22792 CSoutput.n219 CSoutput.n211 4.5005
R22793 CSoutput.n219 CSoutput.n215 4.5005
R22794 CSoutput.n219 CSoutput.n210 4.5005
R22795 CSoutput.n219 CSoutput.t230 4.5005
R22796 CSoutput.n219 CSoutput.n209 4.5005
R22797 CSoutput.n219 CSoutput.n216 4.5005
R22798 CSoutput.n265 CSoutput.n219 4.5005
R22799 CSoutput.n264 CSoutput.n212 4.5005
R22800 CSoutput.n264 CSoutput.n214 4.5005
R22801 CSoutput.n264 CSoutput.n211 4.5005
R22802 CSoutput.n264 CSoutput.n215 4.5005
R22803 CSoutput.n264 CSoutput.n210 4.5005
R22804 CSoutput.n264 CSoutput.t230 4.5005
R22805 CSoutput.n264 CSoutput.n209 4.5005
R22806 CSoutput.n264 CSoutput.n216 4.5005
R22807 CSoutput.n265 CSoutput.n264 4.5005
R22808 CSoutput.n263 CSoutput.n148 4.5005
R22809 CSoutput.n164 CSoutput.n148 4.5005
R22810 CSoutput.n159 CSoutput.n143 4.5005
R22811 CSoutput.n159 CSoutput.n145 4.5005
R22812 CSoutput.n159 CSoutput.n142 4.5005
R22813 CSoutput.n159 CSoutput.n146 4.5005
R22814 CSoutput.n159 CSoutput.n141 4.5005
R22815 CSoutput.n159 CSoutput.t233 4.5005
R22816 CSoutput.n159 CSoutput.n140 4.5005
R22817 CSoutput.n159 CSoutput.n147 4.5005
R22818 CSoutput.n159 CSoutput.n148 4.5005
R22819 CSoutput.n157 CSoutput.n143 4.5005
R22820 CSoutput.n157 CSoutput.n145 4.5005
R22821 CSoutput.n157 CSoutput.n142 4.5005
R22822 CSoutput.n157 CSoutput.n146 4.5005
R22823 CSoutput.n157 CSoutput.n141 4.5005
R22824 CSoutput.n157 CSoutput.t233 4.5005
R22825 CSoutput.n157 CSoutput.n140 4.5005
R22826 CSoutput.n157 CSoutput.n147 4.5005
R22827 CSoutput.n157 CSoutput.n148 4.5005
R22828 CSoutput.n156 CSoutput.n143 4.5005
R22829 CSoutput.n156 CSoutput.n145 4.5005
R22830 CSoutput.n156 CSoutput.n142 4.5005
R22831 CSoutput.n156 CSoutput.n146 4.5005
R22832 CSoutput.n156 CSoutput.n141 4.5005
R22833 CSoutput.n156 CSoutput.t233 4.5005
R22834 CSoutput.n156 CSoutput.n140 4.5005
R22835 CSoutput.n156 CSoutput.n147 4.5005
R22836 CSoutput.n156 CSoutput.n148 4.5005
R22837 CSoutput.n285 CSoutput.n143 4.5005
R22838 CSoutput.n285 CSoutput.n145 4.5005
R22839 CSoutput.n285 CSoutput.n142 4.5005
R22840 CSoutput.n285 CSoutput.n146 4.5005
R22841 CSoutput.n285 CSoutput.n141 4.5005
R22842 CSoutput.n285 CSoutput.t233 4.5005
R22843 CSoutput.n285 CSoutput.n140 4.5005
R22844 CSoutput.n285 CSoutput.n147 4.5005
R22845 CSoutput.n285 CSoutput.n148 4.5005
R22846 CSoutput.n283 CSoutput.n143 4.5005
R22847 CSoutput.n283 CSoutput.n145 4.5005
R22848 CSoutput.n283 CSoutput.n142 4.5005
R22849 CSoutput.n283 CSoutput.n146 4.5005
R22850 CSoutput.n283 CSoutput.n141 4.5005
R22851 CSoutput.n283 CSoutput.t233 4.5005
R22852 CSoutput.n283 CSoutput.n140 4.5005
R22853 CSoutput.n283 CSoutput.n147 4.5005
R22854 CSoutput.n281 CSoutput.n143 4.5005
R22855 CSoutput.n281 CSoutput.n145 4.5005
R22856 CSoutput.n281 CSoutput.n142 4.5005
R22857 CSoutput.n281 CSoutput.n146 4.5005
R22858 CSoutput.n281 CSoutput.n141 4.5005
R22859 CSoutput.n281 CSoutput.t233 4.5005
R22860 CSoutput.n281 CSoutput.n140 4.5005
R22861 CSoutput.n281 CSoutput.n147 4.5005
R22862 CSoutput.n167 CSoutput.n143 4.5005
R22863 CSoutput.n167 CSoutput.n145 4.5005
R22864 CSoutput.n167 CSoutput.n142 4.5005
R22865 CSoutput.n167 CSoutput.n146 4.5005
R22866 CSoutput.n167 CSoutput.n141 4.5005
R22867 CSoutput.n167 CSoutput.t233 4.5005
R22868 CSoutput.n167 CSoutput.n140 4.5005
R22869 CSoutput.n167 CSoutput.n147 4.5005
R22870 CSoutput.n167 CSoutput.n148 4.5005
R22871 CSoutput.n166 CSoutput.n143 4.5005
R22872 CSoutput.n166 CSoutput.n145 4.5005
R22873 CSoutput.n166 CSoutput.n142 4.5005
R22874 CSoutput.n166 CSoutput.n146 4.5005
R22875 CSoutput.n166 CSoutput.n141 4.5005
R22876 CSoutput.n166 CSoutput.t233 4.5005
R22877 CSoutput.n166 CSoutput.n140 4.5005
R22878 CSoutput.n166 CSoutput.n147 4.5005
R22879 CSoutput.n166 CSoutput.n148 4.5005
R22880 CSoutput.n170 CSoutput.n143 4.5005
R22881 CSoutput.n170 CSoutput.n145 4.5005
R22882 CSoutput.n170 CSoutput.n142 4.5005
R22883 CSoutput.n170 CSoutput.n146 4.5005
R22884 CSoutput.n170 CSoutput.n141 4.5005
R22885 CSoutput.n170 CSoutput.t233 4.5005
R22886 CSoutput.n170 CSoutput.n140 4.5005
R22887 CSoutput.n170 CSoutput.n147 4.5005
R22888 CSoutput.n170 CSoutput.n148 4.5005
R22889 CSoutput.n169 CSoutput.n143 4.5005
R22890 CSoutput.n169 CSoutput.n145 4.5005
R22891 CSoutput.n169 CSoutput.n142 4.5005
R22892 CSoutput.n169 CSoutput.n146 4.5005
R22893 CSoutput.n169 CSoutput.n141 4.5005
R22894 CSoutput.n169 CSoutput.t233 4.5005
R22895 CSoutput.n169 CSoutput.n140 4.5005
R22896 CSoutput.n169 CSoutput.n147 4.5005
R22897 CSoutput.n169 CSoutput.n148 4.5005
R22898 CSoutput.n152 CSoutput.n143 4.5005
R22899 CSoutput.n152 CSoutput.n145 4.5005
R22900 CSoutput.n152 CSoutput.n142 4.5005
R22901 CSoutput.n152 CSoutput.n146 4.5005
R22902 CSoutput.n152 CSoutput.n141 4.5005
R22903 CSoutput.n152 CSoutput.t233 4.5005
R22904 CSoutput.n152 CSoutput.n140 4.5005
R22905 CSoutput.n152 CSoutput.n147 4.5005
R22906 CSoutput.n152 CSoutput.n148 4.5005
R22907 CSoutput.n288 CSoutput.n143 4.5005
R22908 CSoutput.n288 CSoutput.n145 4.5005
R22909 CSoutput.n288 CSoutput.n142 4.5005
R22910 CSoutput.n288 CSoutput.n146 4.5005
R22911 CSoutput.n288 CSoutput.n141 4.5005
R22912 CSoutput.n288 CSoutput.t233 4.5005
R22913 CSoutput.n288 CSoutput.n140 4.5005
R22914 CSoutput.n288 CSoutput.n147 4.5005
R22915 CSoutput.n288 CSoutput.n148 4.5005
R22916 CSoutput.n347 CSoutput.n327 4.10845
R22917 CSoutput.n137 CSoutput.n117 4.10845
R22918 CSoutput.n345 CSoutput.t185 4.06363
R22919 CSoutput.n345 CSoutput.t123 4.06363
R22920 CSoutput.n343 CSoutput.t139 4.06363
R22921 CSoutput.n343 CSoutput.t17 4.06363
R22922 CSoutput.n341 CSoutput.t128 4.06363
R22923 CSoutput.n341 CSoutput.t148 4.06363
R22924 CSoutput.n339 CSoutput.t125 4.06363
R22925 CSoutput.n339 CSoutput.t193 4.06363
R22926 CSoutput.n337 CSoutput.t135 4.06363
R22927 CSoutput.n337 CSoutput.t182 4.06363
R22928 CSoutput.n335 CSoutput.t120 4.06363
R22929 CSoutput.n335 CSoutput.t203 4.06363
R22930 CSoutput.n333 CSoutput.t209 4.06363
R22931 CSoutput.n333 CSoutput.t126 4.06363
R22932 CSoutput.n331 CSoutput.t16 4.06363
R22933 CSoutput.n331 CSoutput.t132 4.06363
R22934 CSoutput.n329 CSoutput.t187 4.06363
R22935 CSoutput.n329 CSoutput.t159 4.06363
R22936 CSoutput.n328 CSoutput.t129 4.06363
R22937 CSoutput.n328 CSoutput.t163 4.06363
R22938 CSoutput.n325 CSoutput.t205 4.06363
R22939 CSoutput.n325 CSoutput.t183 4.06363
R22940 CSoutput.n323 CSoutput.t186 4.06363
R22941 CSoutput.n323 CSoutput.t158 4.06363
R22942 CSoutput.n321 CSoutput.t178 4.06363
R22943 CSoutput.n321 CSoutput.t167 4.06363
R22944 CSoutput.n319 CSoutput.t181 4.06363
R22945 CSoutput.n319 CSoutput.t153 4.06363
R22946 CSoutput.n317 CSoutput.t12 4.06363
R22947 CSoutput.n317 CSoutput.t201 4.06363
R22948 CSoutput.n315 CSoutput.t137 4.06363
R22949 CSoutput.n315 CSoutput.t114 4.06363
R22950 CSoutput.n313 CSoutput.t5 4.06363
R22951 CSoutput.n313 CSoutput.t177 4.06363
R22952 CSoutput.n311 CSoutput.t213 4.06363
R22953 CSoutput.n311 CSoutput.t204 4.06363
R22954 CSoutput.n309 CSoutput.t166 4.06363
R22955 CSoutput.n309 CSoutput.t156 4.06363
R22956 CSoutput.n308 CSoutput.t179 4.06363
R22957 CSoutput.n308 CSoutput.t161 4.06363
R22958 CSoutput.n306 CSoutput.t10 4.06363
R22959 CSoutput.n306 CSoutput.t9 4.06363
R22960 CSoutput.n304 CSoutput.t130 4.06363
R22961 CSoutput.n304 CSoutput.t141 4.06363
R22962 CSoutput.n302 CSoutput.t162 4.06363
R22963 CSoutput.n302 CSoutput.t152 4.06363
R22964 CSoutput.n300 CSoutput.t196 4.06363
R22965 CSoutput.n300 CSoutput.t202 4.06363
R22966 CSoutput.n298 CSoutput.t176 4.06363
R22967 CSoutput.n298 CSoutput.t164 4.06363
R22968 CSoutput.n296 CSoutput.t11 4.06363
R22969 CSoutput.n296 CSoutput.t7 4.06363
R22970 CSoutput.n294 CSoutput.t134 4.06363
R22971 CSoutput.n294 CSoutput.t118 4.06363
R22972 CSoutput.n292 CSoutput.t1 4.06363
R22973 CSoutput.n292 CSoutput.t133 4.06363
R22974 CSoutput.n290 CSoutput.t212 4.06363
R22975 CSoutput.n290 CSoutput.t174 4.06363
R22976 CSoutput.n289 CSoutput.t4 4.06363
R22977 CSoutput.n289 CSoutput.t180 4.06363
R22978 CSoutput.n118 CSoutput.t211 4.06363
R22979 CSoutput.n118 CSoutput.t119 4.06363
R22980 CSoutput.n119 CSoutput.t2 4.06363
R22981 CSoutput.n119 CSoutput.t210 4.06363
R22982 CSoutput.n121 CSoutput.t155 4.06363
R22983 CSoutput.n121 CSoutput.t168 4.06363
R22984 CSoutput.n123 CSoutput.t3 4.06363
R22985 CSoutput.n123 CSoutput.t146 4.06363
R22986 CSoutput.n125 CSoutput.t194 4.06363
R22987 CSoutput.n125 CSoutput.t170 4.06363
R22988 CSoutput.n127 CSoutput.t124 4.06363
R22989 CSoutput.n127 CSoutput.t175 4.06363
R22990 CSoutput.n129 CSoutput.t214 4.06363
R22991 CSoutput.n129 CSoutput.t195 4.06363
R22992 CSoutput.n131 CSoutput.t154 4.06363
R22993 CSoutput.n131 CSoutput.t116 4.06363
R22994 CSoutput.n133 CSoutput.t169 4.06363
R22995 CSoutput.n133 CSoutput.t136 4.06363
R22996 CSoutput.n135 CSoutput.t190 4.06363
R22997 CSoutput.n135 CSoutput.t191 4.06363
R22998 CSoutput.n98 CSoutput.t189 4.06363
R22999 CSoutput.n98 CSoutput.t207 4.06363
R23000 CSoutput.n99 CSoutput.t144 4.06363
R23001 CSoutput.n99 CSoutput.t143 4.06363
R23002 CSoutput.n101 CSoutput.t151 4.06363
R23003 CSoutput.n101 CSoutput.t122 4.06363
R23004 CSoutput.n103 CSoutput.t145 4.06363
R23005 CSoutput.n103 CSoutput.t121 4.06363
R23006 CSoutput.n105 CSoutput.t13 4.06363
R23007 CSoutput.n105 CSoutput.t117 4.06363
R23008 CSoutput.n107 CSoutput.t115 4.06363
R23009 CSoutput.n107 CSoutput.t131 4.06363
R23010 CSoutput.n109 CSoutput.t160 4.06363
R23011 CSoutput.n109 CSoutput.t192 4.06363
R23012 CSoutput.n111 CSoutput.t188 4.06363
R23013 CSoutput.n111 CSoutput.t206 4.06363
R23014 CSoutput.n113 CSoutput.t184 4.06363
R23015 CSoutput.n113 CSoutput.t172 4.06363
R23016 CSoutput.n115 CSoutput.t150 4.06363
R23017 CSoutput.n115 CSoutput.t14 4.06363
R23018 CSoutput.n79 CSoutput.t200 4.06363
R23019 CSoutput.n79 CSoutput.t15 4.06363
R23020 CSoutput.n80 CSoutput.t147 4.06363
R23021 CSoutput.n80 CSoutput.t197 4.06363
R23022 CSoutput.n82 CSoutput.t149 4.06363
R23023 CSoutput.n82 CSoutput.t0 4.06363
R23024 CSoutput.n84 CSoutput.t140 4.06363
R23025 CSoutput.n84 CSoutput.t142 4.06363
R23026 CSoutput.n86 CSoutput.t6 4.06363
R23027 CSoutput.n86 CSoutput.t199 4.06363
R23028 CSoutput.n88 CSoutput.t165 4.06363
R23029 CSoutput.n88 CSoutput.t157 4.06363
R23030 CSoutput.n90 CSoutput.t171 4.06363
R23031 CSoutput.n90 CSoutput.t173 4.06363
R23032 CSoutput.n92 CSoutput.t208 4.06363
R23033 CSoutput.n92 CSoutput.t215 4.06363
R23034 CSoutput.n94 CSoutput.t138 4.06363
R23035 CSoutput.n94 CSoutput.t127 4.06363
R23036 CSoutput.n96 CSoutput.t8 4.06363
R23037 CSoutput.n96 CSoutput.t198 4.06363
R23038 CSoutput.n44 CSoutput.n43 3.79402
R23039 CSoutput.n49 CSoutput.n48 3.79402
R23040 CSoutput.n395 CSoutput.n379 3.72967
R23041 CSoutput.n443 CSoutput.n427 3.72967
R23042 CSoutput.n445 CSoutput.n444 3.61338
R23043 CSoutput.n348 CSoutput.n138 3.19963
R23044 CSoutput.n444 CSoutput.n396 3.08965
R23045 CSoutput.n393 CSoutput.t47 2.82907
R23046 CSoutput.n393 CSoutput.t37 2.82907
R23047 CSoutput.n391 CSoutput.t28 2.82907
R23048 CSoutput.n391 CSoutput.t98 2.82907
R23049 CSoutput.n389 CSoutput.t40 2.82907
R23050 CSoutput.n389 CSoutput.t44 2.82907
R23051 CSoutput.n387 CSoutput.t39 2.82907
R23052 CSoutput.n387 CSoutput.t113 2.82907
R23053 CSoutput.n385 CSoutput.t58 2.82907
R23054 CSoutput.n385 CSoutput.t31 2.82907
R23055 CSoutput.n383 CSoutput.t22 2.82907
R23056 CSoutput.n383 CSoutput.t87 2.82907
R23057 CSoutput.n381 CSoutput.t49 2.82907
R23058 CSoutput.n381 CSoutput.t53 2.82907
R23059 CSoutput.n380 CSoutput.t30 2.82907
R23060 CSoutput.n380 CSoutput.t102 2.82907
R23061 CSoutput.n377 CSoutput.t84 2.82907
R23062 CSoutput.n377 CSoutput.t65 2.82907
R23063 CSoutput.n375 CSoutput.t66 2.82907
R23064 CSoutput.n375 CSoutput.t72 2.82907
R23065 CSoutput.n373 CSoutput.t21 2.82907
R23066 CSoutput.n373 CSoutput.t85 2.82907
R23067 CSoutput.n371 CSoutput.t83 2.82907
R23068 CSoutput.n371 CSoutput.t64 2.82907
R23069 CSoutput.n369 CSoutput.t100 2.82907
R23070 CSoutput.n369 CSoutput.t19 2.82907
R23071 CSoutput.n367 CSoutput.t20 2.82907
R23072 CSoutput.n367 CSoutput.t92 2.82907
R23073 CSoutput.n365 CSoutput.t29 2.82907
R23074 CSoutput.n365 CSoutput.t99 2.82907
R23075 CSoutput.n364 CSoutput.t106 2.82907
R23076 CSoutput.n364 CSoutput.t18 2.82907
R23077 CSoutput.n362 CSoutput.t25 2.82907
R23078 CSoutput.n362 CSoutput.t48 2.82907
R23079 CSoutput.n360 CSoutput.t36 2.82907
R23080 CSoutput.n360 CSoutput.t61 2.82907
R23081 CSoutput.n358 CSoutput.t71 2.82907
R23082 CSoutput.n358 CSoutput.t81 2.82907
R23083 CSoutput.n356 CSoutput.t59 2.82907
R23084 CSoutput.n356 CSoutput.t101 2.82907
R23085 CSoutput.n354 CSoutput.t75 2.82907
R23086 CSoutput.n354 CSoutput.t52 2.82907
R23087 CSoutput.n352 CSoutput.t41 2.82907
R23088 CSoutput.n352 CSoutput.t60 2.82907
R23089 CSoutput.n350 CSoutput.t51 2.82907
R23090 CSoutput.n350 CSoutput.t56 2.82907
R23091 CSoutput.n349 CSoutput.t57 2.82907
R23092 CSoutput.n349 CSoutput.t110 2.82907
R23093 CSoutput.n428 CSoutput.t70 2.82907
R23094 CSoutput.n428 CSoutput.t95 2.82907
R23095 CSoutput.n429 CSoutput.t42 2.82907
R23096 CSoutput.n429 CSoutput.t55 2.82907
R23097 CSoutput.n431 CSoutput.t62 2.82907
R23098 CSoutput.n431 CSoutput.t76 2.82907
R23099 CSoutput.n433 CSoutput.t96 2.82907
R23100 CSoutput.n433 CSoutput.t67 2.82907
R23101 CSoutput.n435 CSoutput.t74 2.82907
R23102 CSoutput.n435 CSoutput.t107 2.82907
R23103 CSoutput.n437 CSoutput.t24 2.82907
R23104 CSoutput.n437 CSoutput.t45 2.82907
R23105 CSoutput.n439 CSoutput.t68 2.82907
R23106 CSoutput.n439 CSoutput.t90 2.82907
R23107 CSoutput.n441 CSoutput.t103 2.82907
R23108 CSoutput.n441 CSoutput.t32 2.82907
R23109 CSoutput.n412 CSoutput.t33 2.82907
R23110 CSoutput.n412 CSoutput.t26 2.82907
R23111 CSoutput.n413 CSoutput.t23 2.82907
R23112 CSoutput.n413 CSoutput.t111 2.82907
R23113 CSoutput.n415 CSoutput.t112 2.82907
R23114 CSoutput.n415 CSoutput.t34 2.82907
R23115 CSoutput.n417 CSoutput.t35 2.82907
R23116 CSoutput.n417 CSoutput.t77 2.82907
R23117 CSoutput.n419 CSoutput.t78 2.82907
R23118 CSoutput.n419 CSoutput.t105 2.82907
R23119 CSoutput.n421 CSoutput.t108 2.82907
R23120 CSoutput.n421 CSoutput.t97 2.82907
R23121 CSoutput.n423 CSoutput.t91 2.82907
R23122 CSoutput.n423 CSoutput.t79 2.82907
R23123 CSoutput.n425 CSoutput.t80 2.82907
R23124 CSoutput.n425 CSoutput.t109 2.82907
R23125 CSoutput.n397 CSoutput.t43 2.82907
R23126 CSoutput.n397 CSoutput.t86 2.82907
R23127 CSoutput.n398 CSoutput.t82 2.82907
R23128 CSoutput.n398 CSoutput.t63 2.82907
R23129 CSoutput.n400 CSoutput.t89 2.82907
R23130 CSoutput.n400 CSoutput.t54 2.82907
R23131 CSoutput.n402 CSoutput.t73 2.82907
R23132 CSoutput.n402 CSoutput.t104 2.82907
R23133 CSoutput.n404 CSoutput.t38 2.82907
R23134 CSoutput.n404 CSoutput.t88 2.82907
R23135 CSoutput.n406 CSoutput.t27 2.82907
R23136 CSoutput.n406 CSoutput.t94 2.82907
R23137 CSoutput.n408 CSoutput.t93 2.82907
R23138 CSoutput.n408 CSoutput.t50 2.82907
R23139 CSoutput.n410 CSoutput.t69 2.82907
R23140 CSoutput.n410 CSoutput.t46 2.82907
R23141 CSoutput.n75 CSoutput.n1 2.45513
R23142 CSoutput.n229 CSoutput.n227 2.251
R23143 CSoutput.n229 CSoutput.n226 2.251
R23144 CSoutput.n229 CSoutput.n225 2.251
R23145 CSoutput.n229 CSoutput.n224 2.251
R23146 CSoutput.n198 CSoutput.n197 2.251
R23147 CSoutput.n198 CSoutput.n196 2.251
R23148 CSoutput.n198 CSoutput.n195 2.251
R23149 CSoutput.n198 CSoutput.n194 2.251
R23150 CSoutput.n271 CSoutput.n270 2.251
R23151 CSoutput.n236 CSoutput.n234 2.251
R23152 CSoutput.n236 CSoutput.n233 2.251
R23153 CSoutput.n236 CSoutput.n232 2.251
R23154 CSoutput.n254 CSoutput.n236 2.251
R23155 CSoutput.n242 CSoutput.n241 2.251
R23156 CSoutput.n242 CSoutput.n240 2.251
R23157 CSoutput.n242 CSoutput.n239 2.251
R23158 CSoutput.n242 CSoutput.n238 2.251
R23159 CSoutput.n268 CSoutput.n208 2.251
R23160 CSoutput.n263 CSoutput.n261 2.251
R23161 CSoutput.n263 CSoutput.n260 2.251
R23162 CSoutput.n263 CSoutput.n259 2.251
R23163 CSoutput.n263 CSoutput.n258 2.251
R23164 CSoutput.n164 CSoutput.n163 2.251
R23165 CSoutput.n164 CSoutput.n162 2.251
R23166 CSoutput.n164 CSoutput.n161 2.251
R23167 CSoutput.n164 CSoutput.n160 2.251
R23168 CSoutput.n281 CSoutput.n280 2.251
R23169 CSoutput.n198 CSoutput.n178 2.2505
R23170 CSoutput.n193 CSoutput.n178 2.2505
R23171 CSoutput.n191 CSoutput.n178 2.2505
R23172 CSoutput.n190 CSoutput.n178 2.2505
R23173 CSoutput.n275 CSoutput.n178 2.2505
R23174 CSoutput.n273 CSoutput.n178 2.2505
R23175 CSoutput.n271 CSoutput.n178 2.2505
R23176 CSoutput.n201 CSoutput.n178 2.2505
R23177 CSoutput.n200 CSoutput.n178 2.2505
R23178 CSoutput.n204 CSoutput.n178 2.2505
R23179 CSoutput.n203 CSoutput.n178 2.2505
R23180 CSoutput.n186 CSoutput.n178 2.2505
R23181 CSoutput.n278 CSoutput.n178 2.2505
R23182 CSoutput.n278 CSoutput.n277 2.2505
R23183 CSoutput.n242 CSoutput.n213 2.2505
R23184 CSoutput.n223 CSoutput.n213 2.2505
R23185 CSoutput.n244 CSoutput.n213 2.2505
R23186 CSoutput.n222 CSoutput.n213 2.2505
R23187 CSoutput.n246 CSoutput.n213 2.2505
R23188 CSoutput.n213 CSoutput.n207 2.2505
R23189 CSoutput.n268 CSoutput.n213 2.2505
R23190 CSoutput.n266 CSoutput.n213 2.2505
R23191 CSoutput.n248 CSoutput.n213 2.2505
R23192 CSoutput.n220 CSoutput.n213 2.2505
R23193 CSoutput.n250 CSoutput.n213 2.2505
R23194 CSoutput.n219 CSoutput.n213 2.2505
R23195 CSoutput.n264 CSoutput.n213 2.2505
R23196 CSoutput.n264 CSoutput.n217 2.2505
R23197 CSoutput.n164 CSoutput.n144 2.2505
R23198 CSoutput.n159 CSoutput.n144 2.2505
R23199 CSoutput.n157 CSoutput.n144 2.2505
R23200 CSoutput.n156 CSoutput.n144 2.2505
R23201 CSoutput.n285 CSoutput.n144 2.2505
R23202 CSoutput.n283 CSoutput.n144 2.2505
R23203 CSoutput.n281 CSoutput.n144 2.2505
R23204 CSoutput.n167 CSoutput.n144 2.2505
R23205 CSoutput.n166 CSoutput.n144 2.2505
R23206 CSoutput.n170 CSoutput.n144 2.2505
R23207 CSoutput.n169 CSoutput.n144 2.2505
R23208 CSoutput.n152 CSoutput.n144 2.2505
R23209 CSoutput.n288 CSoutput.n144 2.2505
R23210 CSoutput.n288 CSoutput.n287 2.2505
R23211 CSoutput.n206 CSoutput.n199 2.25024
R23212 CSoutput.n206 CSoutput.n192 2.25024
R23213 CSoutput.n274 CSoutput.n206 2.25024
R23214 CSoutput.n206 CSoutput.n202 2.25024
R23215 CSoutput.n206 CSoutput.n205 2.25024
R23216 CSoutput.n206 CSoutput.n173 2.25024
R23217 CSoutput.n256 CSoutput.n253 2.25024
R23218 CSoutput.n256 CSoutput.n252 2.25024
R23219 CSoutput.n256 CSoutput.n251 2.25024
R23220 CSoutput.n256 CSoutput.n218 2.25024
R23221 CSoutput.n256 CSoutput.n255 2.25024
R23222 CSoutput.n257 CSoutput.n256 2.25024
R23223 CSoutput.n172 CSoutput.n165 2.25024
R23224 CSoutput.n172 CSoutput.n158 2.25024
R23225 CSoutput.n284 CSoutput.n172 2.25024
R23226 CSoutput.n172 CSoutput.n168 2.25024
R23227 CSoutput.n172 CSoutput.n171 2.25024
R23228 CSoutput.n172 CSoutput.n139 2.25024
R23229 CSoutput.n273 CSoutput.n183 1.50111
R23230 CSoutput.n221 CSoutput.n207 1.50111
R23231 CSoutput.n283 CSoutput.n149 1.50111
R23232 CSoutput.n229 CSoutput.n228 1.501
R23233 CSoutput.n236 CSoutput.n235 1.501
R23234 CSoutput.n263 CSoutput.n262 1.501
R23235 CSoutput.n277 CSoutput.n188 1.12536
R23236 CSoutput.n277 CSoutput.n189 1.12536
R23237 CSoutput.n277 CSoutput.n276 1.12536
R23238 CSoutput.n237 CSoutput.n217 1.12536
R23239 CSoutput.n243 CSoutput.n217 1.12536
R23240 CSoutput.n245 CSoutput.n217 1.12536
R23241 CSoutput.n287 CSoutput.n154 1.12536
R23242 CSoutput.n287 CSoutput.n155 1.12536
R23243 CSoutput.n287 CSoutput.n286 1.12536
R23244 CSoutput.n277 CSoutput.n184 1.12536
R23245 CSoutput.n277 CSoutput.n185 1.12536
R23246 CSoutput.n277 CSoutput.n187 1.12536
R23247 CSoutput.n267 CSoutput.n217 1.12536
R23248 CSoutput.n247 CSoutput.n217 1.12536
R23249 CSoutput.n249 CSoutput.n217 1.12536
R23250 CSoutput.n287 CSoutput.n150 1.12536
R23251 CSoutput.n287 CSoutput.n151 1.12536
R23252 CSoutput.n287 CSoutput.n153 1.12536
R23253 CSoutput.n31 CSoutput.n30 0.669944
R23254 CSoutput.n62 CSoutput.n61 0.669944
R23255 CSoutput.n384 CSoutput.n382 0.573776
R23256 CSoutput.n386 CSoutput.n384 0.573776
R23257 CSoutput.n388 CSoutput.n386 0.573776
R23258 CSoutput.n390 CSoutput.n388 0.573776
R23259 CSoutput.n392 CSoutput.n390 0.573776
R23260 CSoutput.n394 CSoutput.n392 0.573776
R23261 CSoutput.n368 CSoutput.n366 0.573776
R23262 CSoutput.n370 CSoutput.n368 0.573776
R23263 CSoutput.n372 CSoutput.n370 0.573776
R23264 CSoutput.n374 CSoutput.n372 0.573776
R23265 CSoutput.n376 CSoutput.n374 0.573776
R23266 CSoutput.n378 CSoutput.n376 0.573776
R23267 CSoutput.n353 CSoutput.n351 0.573776
R23268 CSoutput.n355 CSoutput.n353 0.573776
R23269 CSoutput.n357 CSoutput.n355 0.573776
R23270 CSoutput.n359 CSoutput.n357 0.573776
R23271 CSoutput.n361 CSoutput.n359 0.573776
R23272 CSoutput.n363 CSoutput.n361 0.573776
R23273 CSoutput.n442 CSoutput.n440 0.573776
R23274 CSoutput.n440 CSoutput.n438 0.573776
R23275 CSoutput.n438 CSoutput.n436 0.573776
R23276 CSoutput.n436 CSoutput.n434 0.573776
R23277 CSoutput.n434 CSoutput.n432 0.573776
R23278 CSoutput.n432 CSoutput.n430 0.573776
R23279 CSoutput.n426 CSoutput.n424 0.573776
R23280 CSoutput.n424 CSoutput.n422 0.573776
R23281 CSoutput.n422 CSoutput.n420 0.573776
R23282 CSoutput.n420 CSoutput.n418 0.573776
R23283 CSoutput.n418 CSoutput.n416 0.573776
R23284 CSoutput.n416 CSoutput.n414 0.573776
R23285 CSoutput.n411 CSoutput.n409 0.573776
R23286 CSoutput.n409 CSoutput.n407 0.573776
R23287 CSoutput.n407 CSoutput.n405 0.573776
R23288 CSoutput.n405 CSoutput.n403 0.573776
R23289 CSoutput.n403 CSoutput.n401 0.573776
R23290 CSoutput.n401 CSoutput.n399 0.573776
R23291 CSoutput.n445 CSoutput.n288 0.534303
R23292 CSoutput.n332 CSoutput.n330 0.358259
R23293 CSoutput.n334 CSoutput.n332 0.358259
R23294 CSoutput.n336 CSoutput.n334 0.358259
R23295 CSoutput.n338 CSoutput.n336 0.358259
R23296 CSoutput.n340 CSoutput.n338 0.358259
R23297 CSoutput.n342 CSoutput.n340 0.358259
R23298 CSoutput.n344 CSoutput.n342 0.358259
R23299 CSoutput.n346 CSoutput.n344 0.358259
R23300 CSoutput.n312 CSoutput.n310 0.358259
R23301 CSoutput.n314 CSoutput.n312 0.358259
R23302 CSoutput.n316 CSoutput.n314 0.358259
R23303 CSoutput.n318 CSoutput.n316 0.358259
R23304 CSoutput.n320 CSoutput.n318 0.358259
R23305 CSoutput.n322 CSoutput.n320 0.358259
R23306 CSoutput.n324 CSoutput.n322 0.358259
R23307 CSoutput.n326 CSoutput.n324 0.358259
R23308 CSoutput.n293 CSoutput.n291 0.358259
R23309 CSoutput.n295 CSoutput.n293 0.358259
R23310 CSoutput.n297 CSoutput.n295 0.358259
R23311 CSoutput.n299 CSoutput.n297 0.358259
R23312 CSoutput.n301 CSoutput.n299 0.358259
R23313 CSoutput.n303 CSoutput.n301 0.358259
R23314 CSoutput.n305 CSoutput.n303 0.358259
R23315 CSoutput.n307 CSoutput.n305 0.358259
R23316 CSoutput.n136 CSoutput.n134 0.358259
R23317 CSoutput.n134 CSoutput.n132 0.358259
R23318 CSoutput.n132 CSoutput.n130 0.358259
R23319 CSoutput.n130 CSoutput.n128 0.358259
R23320 CSoutput.n128 CSoutput.n126 0.358259
R23321 CSoutput.n126 CSoutput.n124 0.358259
R23322 CSoutput.n124 CSoutput.n122 0.358259
R23323 CSoutput.n122 CSoutput.n120 0.358259
R23324 CSoutput.n116 CSoutput.n114 0.358259
R23325 CSoutput.n114 CSoutput.n112 0.358259
R23326 CSoutput.n112 CSoutput.n110 0.358259
R23327 CSoutput.n110 CSoutput.n108 0.358259
R23328 CSoutput.n108 CSoutput.n106 0.358259
R23329 CSoutput.n106 CSoutput.n104 0.358259
R23330 CSoutput.n104 CSoutput.n102 0.358259
R23331 CSoutput.n102 CSoutput.n100 0.358259
R23332 CSoutput.n97 CSoutput.n95 0.358259
R23333 CSoutput.n95 CSoutput.n93 0.358259
R23334 CSoutput.n93 CSoutput.n91 0.358259
R23335 CSoutput.n91 CSoutput.n89 0.358259
R23336 CSoutput.n89 CSoutput.n87 0.358259
R23337 CSoutput.n87 CSoutput.n85 0.358259
R23338 CSoutput.n85 CSoutput.n83 0.358259
R23339 CSoutput.n83 CSoutput.n81 0.358259
R23340 CSoutput.n21 CSoutput.n20 0.169105
R23341 CSoutput.n21 CSoutput.n16 0.169105
R23342 CSoutput.n26 CSoutput.n16 0.169105
R23343 CSoutput.n27 CSoutput.n26 0.169105
R23344 CSoutput.n27 CSoutput.n14 0.169105
R23345 CSoutput.n32 CSoutput.n14 0.169105
R23346 CSoutput.n33 CSoutput.n32 0.169105
R23347 CSoutput.n34 CSoutput.n33 0.169105
R23348 CSoutput.n34 CSoutput.n12 0.169105
R23349 CSoutput.n39 CSoutput.n12 0.169105
R23350 CSoutput.n40 CSoutput.n39 0.169105
R23351 CSoutput.n40 CSoutput.n10 0.169105
R23352 CSoutput.n45 CSoutput.n10 0.169105
R23353 CSoutput.n46 CSoutput.n45 0.169105
R23354 CSoutput.n47 CSoutput.n46 0.169105
R23355 CSoutput.n47 CSoutput.n8 0.169105
R23356 CSoutput.n52 CSoutput.n8 0.169105
R23357 CSoutput.n53 CSoutput.n52 0.169105
R23358 CSoutput.n53 CSoutput.n6 0.169105
R23359 CSoutput.n58 CSoutput.n6 0.169105
R23360 CSoutput.n59 CSoutput.n58 0.169105
R23361 CSoutput.n60 CSoutput.n59 0.169105
R23362 CSoutput.n60 CSoutput.n4 0.169105
R23363 CSoutput.n66 CSoutput.n4 0.169105
R23364 CSoutput.n67 CSoutput.n66 0.169105
R23365 CSoutput.n68 CSoutput.n67 0.169105
R23366 CSoutput.n68 CSoutput.n2 0.169105
R23367 CSoutput.n73 CSoutput.n2 0.169105
R23368 CSoutput.n74 CSoutput.n73 0.169105
R23369 CSoutput.n74 CSoutput.n0 0.169105
R23370 CSoutput.n78 CSoutput.n0 0.169105
R23371 CSoutput.n231 CSoutput.n230 0.0910737
R23372 CSoutput.n282 CSoutput.n279 0.0723685
R23373 CSoutput.n236 CSoutput.n231 0.0522944
R23374 CSoutput.n279 CSoutput.n278 0.0499135
R23375 CSoutput.n230 CSoutput.n229 0.0499135
R23376 CSoutput.n264 CSoutput.n263 0.0464294
R23377 CSoutput.n272 CSoutput.n269 0.0391444
R23378 CSoutput.n231 CSoutput.t235 0.023435
R23379 CSoutput.n279 CSoutput.t219 0.02262
R23380 CSoutput.n230 CSoutput.t229 0.02262
R23381 CSoutput CSoutput.n445 0.0052
R23382 CSoutput.n201 CSoutput.n184 0.00365111
R23383 CSoutput.n204 CSoutput.n185 0.00365111
R23384 CSoutput.n187 CSoutput.n186 0.00365111
R23385 CSoutput.n229 CSoutput.n188 0.00365111
R23386 CSoutput.n193 CSoutput.n189 0.00365111
R23387 CSoutput.n276 CSoutput.n190 0.00365111
R23388 CSoutput.n267 CSoutput.n266 0.00365111
R23389 CSoutput.n247 CSoutput.n220 0.00365111
R23390 CSoutput.n249 CSoutput.n219 0.00365111
R23391 CSoutput.n237 CSoutput.n236 0.00365111
R23392 CSoutput.n243 CSoutput.n223 0.00365111
R23393 CSoutput.n245 CSoutput.n222 0.00365111
R23394 CSoutput.n167 CSoutput.n150 0.00365111
R23395 CSoutput.n170 CSoutput.n151 0.00365111
R23396 CSoutput.n153 CSoutput.n152 0.00365111
R23397 CSoutput.n263 CSoutput.n154 0.00365111
R23398 CSoutput.n159 CSoutput.n155 0.00365111
R23399 CSoutput.n286 CSoutput.n156 0.00365111
R23400 CSoutput.n198 CSoutput.n188 0.00340054
R23401 CSoutput.n191 CSoutput.n189 0.00340054
R23402 CSoutput.n276 CSoutput.n275 0.00340054
R23403 CSoutput.n271 CSoutput.n184 0.00340054
R23404 CSoutput.n200 CSoutput.n185 0.00340054
R23405 CSoutput.n203 CSoutput.n187 0.00340054
R23406 CSoutput.n242 CSoutput.n237 0.00340054
R23407 CSoutput.n244 CSoutput.n243 0.00340054
R23408 CSoutput.n246 CSoutput.n245 0.00340054
R23409 CSoutput.n268 CSoutput.n267 0.00340054
R23410 CSoutput.n248 CSoutput.n247 0.00340054
R23411 CSoutput.n250 CSoutput.n249 0.00340054
R23412 CSoutput.n164 CSoutput.n154 0.00340054
R23413 CSoutput.n157 CSoutput.n155 0.00340054
R23414 CSoutput.n286 CSoutput.n285 0.00340054
R23415 CSoutput.n281 CSoutput.n150 0.00340054
R23416 CSoutput.n166 CSoutput.n151 0.00340054
R23417 CSoutput.n169 CSoutput.n153 0.00340054
R23418 CSoutput.n199 CSoutput.n193 0.00252698
R23419 CSoutput.n192 CSoutput.n190 0.00252698
R23420 CSoutput.n274 CSoutput.n273 0.00252698
R23421 CSoutput.n202 CSoutput.n200 0.00252698
R23422 CSoutput.n205 CSoutput.n203 0.00252698
R23423 CSoutput.n278 CSoutput.n173 0.00252698
R23424 CSoutput.n199 CSoutput.n198 0.00252698
R23425 CSoutput.n192 CSoutput.n191 0.00252698
R23426 CSoutput.n275 CSoutput.n274 0.00252698
R23427 CSoutput.n202 CSoutput.n201 0.00252698
R23428 CSoutput.n205 CSoutput.n204 0.00252698
R23429 CSoutput.n186 CSoutput.n173 0.00252698
R23430 CSoutput.n253 CSoutput.n223 0.00252698
R23431 CSoutput.n252 CSoutput.n222 0.00252698
R23432 CSoutput.n251 CSoutput.n207 0.00252698
R23433 CSoutput.n248 CSoutput.n218 0.00252698
R23434 CSoutput.n255 CSoutput.n250 0.00252698
R23435 CSoutput.n264 CSoutput.n257 0.00252698
R23436 CSoutput.n253 CSoutput.n242 0.00252698
R23437 CSoutput.n252 CSoutput.n244 0.00252698
R23438 CSoutput.n251 CSoutput.n246 0.00252698
R23439 CSoutput.n266 CSoutput.n218 0.00252698
R23440 CSoutput.n255 CSoutput.n220 0.00252698
R23441 CSoutput.n257 CSoutput.n219 0.00252698
R23442 CSoutput.n165 CSoutput.n159 0.00252698
R23443 CSoutput.n158 CSoutput.n156 0.00252698
R23444 CSoutput.n284 CSoutput.n283 0.00252698
R23445 CSoutput.n168 CSoutput.n166 0.00252698
R23446 CSoutput.n171 CSoutput.n169 0.00252698
R23447 CSoutput.n288 CSoutput.n139 0.00252698
R23448 CSoutput.n165 CSoutput.n164 0.00252698
R23449 CSoutput.n158 CSoutput.n157 0.00252698
R23450 CSoutput.n285 CSoutput.n284 0.00252698
R23451 CSoutput.n168 CSoutput.n167 0.00252698
R23452 CSoutput.n171 CSoutput.n170 0.00252698
R23453 CSoutput.n152 CSoutput.n139 0.00252698
R23454 CSoutput.n273 CSoutput.n272 0.0020275
R23455 CSoutput.n272 CSoutput.n271 0.0020275
R23456 CSoutput.n269 CSoutput.n207 0.0020275
R23457 CSoutput.n269 CSoutput.n268 0.0020275
R23458 CSoutput.n283 CSoutput.n282 0.0020275
R23459 CSoutput.n282 CSoutput.n281 0.0020275
R23460 CSoutput.n183 CSoutput.n182 0.00166668
R23461 CSoutput.n265 CSoutput.n221 0.00166668
R23462 CSoutput.n149 CSoutput.n148 0.00166668
R23463 CSoutput.n287 CSoutput.n149 0.00133328
R23464 CSoutput.n221 CSoutput.n217 0.00133328
R23465 CSoutput.n277 CSoutput.n183 0.00133328
R23466 CSoutput.n280 CSoutput.n172 0.001
R23467 CSoutput.n258 CSoutput.n172 0.001
R23468 CSoutput.n160 CSoutput.n140 0.001
R23469 CSoutput.n259 CSoutput.n140 0.001
R23470 CSoutput.n161 CSoutput.n141 0.001
R23471 CSoutput.n260 CSoutput.n141 0.001
R23472 CSoutput.n162 CSoutput.n142 0.001
R23473 CSoutput.n261 CSoutput.n142 0.001
R23474 CSoutput.n163 CSoutput.n143 0.001
R23475 CSoutput.n262 CSoutput.n143 0.001
R23476 CSoutput.n256 CSoutput.n208 0.001
R23477 CSoutput.n256 CSoutput.n254 0.001
R23478 CSoutput.n238 CSoutput.n209 0.001
R23479 CSoutput.n232 CSoutput.n209 0.001
R23480 CSoutput.n239 CSoutput.n210 0.001
R23481 CSoutput.n233 CSoutput.n210 0.001
R23482 CSoutput.n240 CSoutput.n211 0.001
R23483 CSoutput.n234 CSoutput.n211 0.001
R23484 CSoutput.n241 CSoutput.n212 0.001
R23485 CSoutput.n235 CSoutput.n212 0.001
R23486 CSoutput.n270 CSoutput.n206 0.001
R23487 CSoutput.n224 CSoutput.n206 0.001
R23488 CSoutput.n194 CSoutput.n174 0.001
R23489 CSoutput.n225 CSoutput.n174 0.001
R23490 CSoutput.n195 CSoutput.n175 0.001
R23491 CSoutput.n226 CSoutput.n175 0.001
R23492 CSoutput.n196 CSoutput.n176 0.001
R23493 CSoutput.n227 CSoutput.n176 0.001
R23494 CSoutput.n197 CSoutput.n177 0.001
R23495 CSoutput.n228 CSoutput.n177 0.001
R23496 CSoutput.n228 CSoutput.n178 0.001
R23497 CSoutput.n227 CSoutput.n179 0.001
R23498 CSoutput.n226 CSoutput.n180 0.001
R23499 CSoutput.n225 CSoutput.t222 0.001
R23500 CSoutput.n224 CSoutput.n181 0.001
R23501 CSoutput.n197 CSoutput.n179 0.001
R23502 CSoutput.n196 CSoutput.n180 0.001
R23503 CSoutput.n195 CSoutput.t222 0.001
R23504 CSoutput.n194 CSoutput.n181 0.001
R23505 CSoutput.n270 CSoutput.n182 0.001
R23506 CSoutput.n235 CSoutput.n213 0.001
R23507 CSoutput.n234 CSoutput.n214 0.001
R23508 CSoutput.n233 CSoutput.n215 0.001
R23509 CSoutput.n232 CSoutput.t230 0.001
R23510 CSoutput.n254 CSoutput.n216 0.001
R23511 CSoutput.n241 CSoutput.n214 0.001
R23512 CSoutput.n240 CSoutput.n215 0.001
R23513 CSoutput.n239 CSoutput.t230 0.001
R23514 CSoutput.n238 CSoutput.n216 0.001
R23515 CSoutput.n265 CSoutput.n208 0.001
R23516 CSoutput.n262 CSoutput.n144 0.001
R23517 CSoutput.n261 CSoutput.n145 0.001
R23518 CSoutput.n260 CSoutput.n146 0.001
R23519 CSoutput.n259 CSoutput.t233 0.001
R23520 CSoutput.n258 CSoutput.n147 0.001
R23521 CSoutput.n163 CSoutput.n145 0.001
R23522 CSoutput.n162 CSoutput.n146 0.001
R23523 CSoutput.n161 CSoutput.t233 0.001
R23524 CSoutput.n160 CSoutput.n147 0.001
R23525 CSoutput.n280 CSoutput.n148 0.001
R23526 a_n9628_8799.n231 a_n9628_8799.t145 485.149
R23527 a_n9628_8799.n250 a_n9628_8799.t159 485.149
R23528 a_n9628_8799.n270 a_n9628_8799.t83 485.149
R23529 a_n9628_8799.n170 a_n9628_8799.t98 485.149
R23530 a_n9628_8799.n189 a_n9628_8799.t110 485.149
R23531 a_n9628_8799.n209 a_n9628_8799.t82 485.149
R23532 a_n9628_8799.n56 a_n9628_8799.t55 485.135
R23533 a_n9628_8799.n243 a_n9628_8799.t53 464.166
R23534 a_n9628_8799.n225 a_n9628_8799.t139 464.166
R23535 a_n9628_8799.n242 a_n9628_8799.t75 464.166
R23536 a_n9628_8799.n241 a_n9628_8799.t58 464.166
R23537 a_n9628_8799.n226 a_n9628_8799.t146 464.166
R23538 a_n9628_8799.n240 a_n9628_8799.t101 464.166
R23539 a_n9628_8799.n239 a_n9628_8799.t76 464.166
R23540 a_n9628_8799.n227 a_n9628_8799.t164 464.166
R23541 a_n9628_8799.n238 a_n9628_8799.t119 464.166
R23542 a_n9628_8799.n237 a_n9628_8799.t79 464.166
R23543 a_n9628_8799.n228 a_n9628_8799.t158 464.166
R23544 a_n9628_8799.n236 a_n9628_8799.t121 464.166
R23545 a_n9628_8799.n235 a_n9628_8799.t93 464.166
R23546 a_n9628_8799.n229 a_n9628_8799.t54 464.166
R23547 a_n9628_8799.n234 a_n9628_8799.t142 464.166
R23548 a_n9628_8799.n233 a_n9628_8799.t123 464.166
R23549 a_n9628_8799.n230 a_n9628_8799.t59 464.166
R23550 a_n9628_8799.n232 a_n9628_8799.t149 464.166
R23551 a_n9628_8799.n71 a_n9628_8799.t67 485.135
R23552 a_n9628_8799.n262 a_n9628_8799.t65 464.166
R23553 a_n9628_8799.n244 a_n9628_8799.t156 464.166
R23554 a_n9628_8799.n261 a_n9628_8799.t84 464.166
R23555 a_n9628_8799.n260 a_n9628_8799.t73 464.166
R23556 a_n9628_8799.n245 a_n9628_8799.t160 464.166
R23557 a_n9628_8799.n259 a_n9628_8799.t115 464.166
R23558 a_n9628_8799.n258 a_n9628_8799.t87 464.166
R23559 a_n9628_8799.n246 a_n9628_8799.t57 464.166
R23560 a_n9628_8799.n257 a_n9628_8799.t132 464.166
R23561 a_n9628_8799.n256 a_n9628_8799.t88 464.166
R23562 a_n9628_8799.n247 a_n9628_8799.t49 464.166
R23563 a_n9628_8799.n255 a_n9628_8799.t137 464.166
R23564 a_n9628_8799.n254 a_n9628_8799.t103 464.166
R23565 a_n9628_8799.n248 a_n9628_8799.t66 464.166
R23566 a_n9628_8799.n253 a_n9628_8799.t157 464.166
R23567 a_n9628_8799.n252 a_n9628_8799.t138 464.166
R23568 a_n9628_8799.n249 a_n9628_8799.t74 464.166
R23569 a_n9628_8799.n251 a_n9628_8799.t161 464.166
R23570 a_n9628_8799.n86 a_n9628_8799.t114 485.135
R23571 a_n9628_8799.n282 a_n9628_8799.t136 464.166
R23572 a_n9628_8799.n264 a_n9628_8799.t72 464.166
R23573 a_n9628_8799.n281 a_n9628_8799.t154 464.166
R23574 a_n9628_8799.n280 a_n9628_8799.t91 464.166
R23575 a_n9628_8799.n265 a_n9628_8799.t147 464.166
R23576 a_n9628_8799.n279 a_n9628_8799.t78 464.166
R23577 a_n9628_8799.n278 a_n9628_8799.t126 464.166
R23578 a_n9628_8799.n266 a_n9628_8799.t63 464.166
R23579 a_n9628_8799.n277 a_n9628_8799.t109 464.166
R23580 a_n9628_8799.n276 a_n9628_8799.t86 464.166
R23581 a_n9628_8799.n267 a_n9628_8799.t134 464.166
R23582 a_n9628_8799.n275 a_n9628_8799.t70 464.166
R23583 a_n9628_8799.n274 a_n9628_8799.t118 464.166
R23584 a_n9628_8799.n268 a_n9628_8799.t52 464.166
R23585 a_n9628_8799.n273 a_n9628_8799.t102 464.166
R23586 a_n9628_8799.n272 a_n9628_8799.t166 464.166
R23587 a_n9628_8799.n269 a_n9628_8799.t125 464.166
R23588 a_n9628_8799.n271 a_n9628_8799.t62 464.166
R23589 a_n9628_8799.n171 a_n9628_8799.t99 464.166
R23590 a_n9628_8799.n172 a_n9628_8799.t131 464.166
R23591 a_n9628_8799.n173 a_n9628_8799.t56 464.166
R23592 a_n9628_8799.n174 a_n9628_8799.t96 464.166
R23593 a_n9628_8799.n169 a_n9628_8799.t128 464.166
R23594 a_n9628_8799.n175 a_n9628_8799.t50 464.166
R23595 a_n9628_8799.n176 a_n9628_8799.t81 464.166
R23596 a_n9628_8799.n177 a_n9628_8799.t120 464.166
R23597 a_n9628_8799.n178 a_n9628_8799.t155 464.166
R23598 a_n9628_8799.n168 a_n9628_8799.t80 464.166
R23599 a_n9628_8799.n179 a_n9628_8799.t116 464.166
R23600 a_n9628_8799.n167 a_n9628_8799.t151 464.166
R23601 a_n9628_8799.n180 a_n9628_8799.t152 464.166
R23602 a_n9628_8799.n181 a_n9628_8799.t97 464.166
R23603 a_n9628_8799.n182 a_n9628_8799.t130 464.166
R23604 a_n9628_8799.n183 a_n9628_8799.t150 464.166
R23605 a_n9628_8799.n166 a_n9628_8799.t94 464.166
R23606 a_n9628_8799.n184 a_n9628_8799.t95 464.166
R23607 a_n9628_8799.n190 a_n9628_8799.t112 464.166
R23608 a_n9628_8799.n191 a_n9628_8799.t148 464.166
R23609 a_n9628_8799.n192 a_n9628_8799.t68 464.166
R23610 a_n9628_8799.n193 a_n9628_8799.t106 464.166
R23611 a_n9628_8799.n188 a_n9628_8799.t140 464.166
R23612 a_n9628_8799.n194 a_n9628_8799.t64 464.166
R23613 a_n9628_8799.n195 a_n9628_8799.t92 464.166
R23614 a_n9628_8799.n196 a_n9628_8799.t133 464.166
R23615 a_n9628_8799.n197 a_n9628_8799.t167 464.166
R23616 a_n9628_8799.n187 a_n9628_8799.t89 464.166
R23617 a_n9628_8799.n198 a_n9628_8799.t129 464.166
R23618 a_n9628_8799.n186 a_n9628_8799.t163 464.166
R23619 a_n9628_8799.n199 a_n9628_8799.t165 464.166
R23620 a_n9628_8799.n200 a_n9628_8799.t111 464.166
R23621 a_n9628_8799.n201 a_n9628_8799.t144 464.166
R23622 a_n9628_8799.n202 a_n9628_8799.t162 464.166
R23623 a_n9628_8799.n185 a_n9628_8799.t105 464.166
R23624 a_n9628_8799.n203 a_n9628_8799.t107 464.166
R23625 a_n9628_8799.n210 a_n9628_8799.t60 464.166
R23626 a_n9628_8799.n211 a_n9628_8799.t122 464.166
R23627 a_n9628_8799.n212 a_n9628_8799.t77 464.166
R23628 a_n9628_8799.n213 a_n9628_8799.t100 464.166
R23629 a_n9628_8799.n208 a_n9628_8799.t51 464.166
R23630 a_n9628_8799.n214 a_n9628_8799.t117 464.166
R23631 a_n9628_8799.n215 a_n9628_8799.t69 464.166
R23632 a_n9628_8799.n216 a_n9628_8799.t135 464.166
R23633 a_n9628_8799.n217 a_n9628_8799.t85 464.166
R23634 a_n9628_8799.n207 a_n9628_8799.t108 464.166
R23635 a_n9628_8799.n218 a_n9628_8799.t61 464.166
R23636 a_n9628_8799.n206 a_n9628_8799.t124 464.166
R23637 a_n9628_8799.n219 a_n9628_8799.t104 464.166
R23638 a_n9628_8799.n220 a_n9628_8799.t143 464.166
R23639 a_n9628_8799.n221 a_n9628_8799.t90 464.166
R23640 a_n9628_8799.n222 a_n9628_8799.t153 464.166
R23641 a_n9628_8799.n205 a_n9628_8799.t71 464.166
R23642 a_n9628_8799.n223 a_n9628_8799.t48 464.166
R23643 a_n9628_8799.n41 a_n9628_8799.n70 71.7212
R23644 a_n9628_8799.n70 a_n9628_8799.n230 17.8606
R23645 a_n9628_8799.n69 a_n9628_8799.n41 76.9909
R23646 a_n9628_8799.n233 a_n9628_8799.n69 7.32118
R23647 a_n9628_8799.n68 a_n9628_8799.n40 78.3454
R23648 a_n9628_8799.n40 a_n9628_8799.n67 72.8951
R23649 a_n9628_8799.n66 a_n9628_8799.n42 70.1674
R23650 a_n9628_8799.n236 a_n9628_8799.n66 20.9683
R23651 a_n9628_8799.n42 a_n9628_8799.n65 72.3034
R23652 a_n9628_8799.n65 a_n9628_8799.n228 16.6962
R23653 a_n9628_8799.n64 a_n9628_8799.n43 77.6622
R23654 a_n9628_8799.n237 a_n9628_8799.n64 5.97853
R23655 a_n9628_8799.n63 a_n9628_8799.n43 77.6622
R23656 a_n9628_8799.n44 a_n9628_8799.n62 72.3034
R23657 a_n9628_8799.n61 a_n9628_8799.n44 70.1674
R23658 a_n9628_8799.n240 a_n9628_8799.n61 20.9683
R23659 a_n9628_8799.n46 a_n9628_8799.n60 72.8951
R23660 a_n9628_8799.n60 a_n9628_8799.n226 15.5127
R23661 a_n9628_8799.n59 a_n9628_8799.n46 78.3454
R23662 a_n9628_8799.n241 a_n9628_8799.n59 4.61226
R23663 a_n9628_8799.n58 a_n9628_8799.n45 76.9909
R23664 a_n9628_8799.n45 a_n9628_8799.n57 71.7212
R23665 a_n9628_8799.n243 a_n9628_8799.n56 20.9683
R23666 a_n9628_8799.n47 a_n9628_8799.n56 70.1674
R23667 a_n9628_8799.n33 a_n9628_8799.n85 71.7212
R23668 a_n9628_8799.n85 a_n9628_8799.n249 17.8606
R23669 a_n9628_8799.n84 a_n9628_8799.n33 76.9909
R23670 a_n9628_8799.n252 a_n9628_8799.n84 7.32118
R23671 a_n9628_8799.n83 a_n9628_8799.n32 78.3454
R23672 a_n9628_8799.n32 a_n9628_8799.n82 72.8951
R23673 a_n9628_8799.n81 a_n9628_8799.n34 70.1674
R23674 a_n9628_8799.n255 a_n9628_8799.n81 20.9683
R23675 a_n9628_8799.n34 a_n9628_8799.n80 72.3034
R23676 a_n9628_8799.n80 a_n9628_8799.n247 16.6962
R23677 a_n9628_8799.n79 a_n9628_8799.n35 77.6622
R23678 a_n9628_8799.n256 a_n9628_8799.n79 5.97853
R23679 a_n9628_8799.n78 a_n9628_8799.n35 77.6622
R23680 a_n9628_8799.n36 a_n9628_8799.n77 72.3034
R23681 a_n9628_8799.n76 a_n9628_8799.n36 70.1674
R23682 a_n9628_8799.n259 a_n9628_8799.n76 20.9683
R23683 a_n9628_8799.n38 a_n9628_8799.n75 72.8951
R23684 a_n9628_8799.n75 a_n9628_8799.n245 15.5127
R23685 a_n9628_8799.n74 a_n9628_8799.n38 78.3454
R23686 a_n9628_8799.n260 a_n9628_8799.n74 4.61226
R23687 a_n9628_8799.n73 a_n9628_8799.n37 76.9909
R23688 a_n9628_8799.n37 a_n9628_8799.n72 71.7212
R23689 a_n9628_8799.n262 a_n9628_8799.n71 20.9683
R23690 a_n9628_8799.n39 a_n9628_8799.n71 70.1674
R23691 a_n9628_8799.n25 a_n9628_8799.n100 71.7212
R23692 a_n9628_8799.n100 a_n9628_8799.n269 17.8606
R23693 a_n9628_8799.n99 a_n9628_8799.n25 76.9909
R23694 a_n9628_8799.n272 a_n9628_8799.n99 7.32118
R23695 a_n9628_8799.n98 a_n9628_8799.n24 78.3454
R23696 a_n9628_8799.n24 a_n9628_8799.n97 72.8951
R23697 a_n9628_8799.n96 a_n9628_8799.n26 70.1674
R23698 a_n9628_8799.n275 a_n9628_8799.n96 20.9683
R23699 a_n9628_8799.n26 a_n9628_8799.n95 72.3034
R23700 a_n9628_8799.n95 a_n9628_8799.n267 16.6962
R23701 a_n9628_8799.n94 a_n9628_8799.n27 77.6622
R23702 a_n9628_8799.n276 a_n9628_8799.n94 5.97853
R23703 a_n9628_8799.n93 a_n9628_8799.n27 77.6622
R23704 a_n9628_8799.n28 a_n9628_8799.n92 72.3034
R23705 a_n9628_8799.n91 a_n9628_8799.n28 70.1674
R23706 a_n9628_8799.n279 a_n9628_8799.n91 20.9683
R23707 a_n9628_8799.n30 a_n9628_8799.n90 72.8951
R23708 a_n9628_8799.n90 a_n9628_8799.n265 15.5127
R23709 a_n9628_8799.n89 a_n9628_8799.n30 78.3454
R23710 a_n9628_8799.n280 a_n9628_8799.n89 4.61226
R23711 a_n9628_8799.n88 a_n9628_8799.n29 76.9909
R23712 a_n9628_8799.n29 a_n9628_8799.n87 71.7212
R23713 a_n9628_8799.n282 a_n9628_8799.n86 20.9683
R23714 a_n9628_8799.n31 a_n9628_8799.n86 70.1674
R23715 a_n9628_8799.n17 a_n9628_8799.n115 70.1674
R23716 a_n9628_8799.n184 a_n9628_8799.n115 20.9683
R23717 a_n9628_8799.n114 a_n9628_8799.n17 71.7212
R23718 a_n9628_8799.n114 a_n9628_8799.n166 17.8606
R23719 a_n9628_8799.n16 a_n9628_8799.n113 76.9909
R23720 a_n9628_8799.n183 a_n9628_8799.n113 7.32118
R23721 a_n9628_8799.n112 a_n9628_8799.n16 78.3454
R23722 a_n9628_8799.n18 a_n9628_8799.n111 72.8951
R23723 a_n9628_8799.n110 a_n9628_8799.n18 70.1674
R23724 a_n9628_8799.n110 a_n9628_8799.n167 20.9683
R23725 a_n9628_8799.n19 a_n9628_8799.n109 72.3034
R23726 a_n9628_8799.n179 a_n9628_8799.n109 16.6962
R23727 a_n9628_8799.n108 a_n9628_8799.n19 77.6622
R23728 a_n9628_8799.n108 a_n9628_8799.n168 5.97853
R23729 a_n9628_8799.n20 a_n9628_8799.n107 77.6622
R23730 a_n9628_8799.n106 a_n9628_8799.n20 72.3034
R23731 a_n9628_8799.n21 a_n9628_8799.n105 70.1674
R23732 a_n9628_8799.n175 a_n9628_8799.n105 20.9683
R23733 a_n9628_8799.n104 a_n9628_8799.n21 72.8951
R23734 a_n9628_8799.n104 a_n9628_8799.n169 15.5127
R23735 a_n9628_8799.n22 a_n9628_8799.n103 78.3454
R23736 a_n9628_8799.n174 a_n9628_8799.n103 4.61226
R23737 a_n9628_8799.n102 a_n9628_8799.n22 76.9909
R23738 a_n9628_8799.n101 a_n9628_8799.n172 17.8606
R23739 a_n9628_8799.n101 a_n9628_8799.n23 71.7212
R23740 a_n9628_8799.n9 a_n9628_8799.n130 70.1674
R23741 a_n9628_8799.n203 a_n9628_8799.n130 20.9683
R23742 a_n9628_8799.n129 a_n9628_8799.n9 71.7212
R23743 a_n9628_8799.n129 a_n9628_8799.n185 17.8606
R23744 a_n9628_8799.n8 a_n9628_8799.n128 76.9909
R23745 a_n9628_8799.n202 a_n9628_8799.n128 7.32118
R23746 a_n9628_8799.n127 a_n9628_8799.n8 78.3454
R23747 a_n9628_8799.n10 a_n9628_8799.n126 72.8951
R23748 a_n9628_8799.n125 a_n9628_8799.n10 70.1674
R23749 a_n9628_8799.n125 a_n9628_8799.n186 20.9683
R23750 a_n9628_8799.n11 a_n9628_8799.n124 72.3034
R23751 a_n9628_8799.n198 a_n9628_8799.n124 16.6962
R23752 a_n9628_8799.n123 a_n9628_8799.n11 77.6622
R23753 a_n9628_8799.n123 a_n9628_8799.n187 5.97853
R23754 a_n9628_8799.n12 a_n9628_8799.n122 77.6622
R23755 a_n9628_8799.n121 a_n9628_8799.n12 72.3034
R23756 a_n9628_8799.n13 a_n9628_8799.n120 70.1674
R23757 a_n9628_8799.n194 a_n9628_8799.n120 20.9683
R23758 a_n9628_8799.n119 a_n9628_8799.n13 72.8951
R23759 a_n9628_8799.n119 a_n9628_8799.n188 15.5127
R23760 a_n9628_8799.n14 a_n9628_8799.n118 78.3454
R23761 a_n9628_8799.n193 a_n9628_8799.n118 4.61226
R23762 a_n9628_8799.n117 a_n9628_8799.n14 76.9909
R23763 a_n9628_8799.n116 a_n9628_8799.n191 17.8606
R23764 a_n9628_8799.n116 a_n9628_8799.n15 71.7212
R23765 a_n9628_8799.n1 a_n9628_8799.n145 70.1674
R23766 a_n9628_8799.n223 a_n9628_8799.n145 20.9683
R23767 a_n9628_8799.n144 a_n9628_8799.n1 71.7212
R23768 a_n9628_8799.n144 a_n9628_8799.n205 17.8606
R23769 a_n9628_8799.n0 a_n9628_8799.n143 76.9909
R23770 a_n9628_8799.n222 a_n9628_8799.n143 7.32118
R23771 a_n9628_8799.n142 a_n9628_8799.n0 78.3454
R23772 a_n9628_8799.n2 a_n9628_8799.n141 72.8951
R23773 a_n9628_8799.n140 a_n9628_8799.n2 70.1674
R23774 a_n9628_8799.n140 a_n9628_8799.n206 20.9683
R23775 a_n9628_8799.n3 a_n9628_8799.n139 72.3034
R23776 a_n9628_8799.n218 a_n9628_8799.n139 16.6962
R23777 a_n9628_8799.n138 a_n9628_8799.n3 77.6622
R23778 a_n9628_8799.n138 a_n9628_8799.n207 5.97853
R23779 a_n9628_8799.n4 a_n9628_8799.n137 77.6622
R23780 a_n9628_8799.n136 a_n9628_8799.n4 72.3034
R23781 a_n9628_8799.n5 a_n9628_8799.n135 70.1674
R23782 a_n9628_8799.n214 a_n9628_8799.n135 20.9683
R23783 a_n9628_8799.n134 a_n9628_8799.n5 72.8951
R23784 a_n9628_8799.n134 a_n9628_8799.n208 15.5127
R23785 a_n9628_8799.n6 a_n9628_8799.n133 78.3454
R23786 a_n9628_8799.n213 a_n9628_8799.n133 4.61226
R23787 a_n9628_8799.n132 a_n9628_8799.n6 76.9909
R23788 a_n9628_8799.n131 a_n9628_8799.n211 17.8606
R23789 a_n9628_8799.n131 a_n9628_8799.n7 71.7212
R23790 a_n9628_8799.n291 a_n9628_8799.n146 98.9633
R23791 a_n9628_8799.n51 a_n9628_8799.n147 98.9631
R23792 a_n9628_8799.n53 a_n9628_8799.n287 98.6055
R23793 a_n9628_8799.n53 a_n9628_8799.n288 98.6055
R23794 a_n9628_8799.n54 a_n9628_8799.n289 98.6055
R23795 a_n9628_8799.n54 a_n9628_8799.n290 98.6055
R23796 a_n9628_8799.n51 a_n9628_8799.n148 98.6055
R23797 a_n9628_8799.n51 a_n9628_8799.n149 98.6055
R23798 a_n9628_8799.n52 a_n9628_8799.n150 98.6055
R23799 a_n9628_8799.n52 a_n9628_8799.n151 98.6055
R23800 a_n9628_8799.n153 a_n9628_8799.n152 98.6055
R23801 a_n9628_8799.n292 a_n9628_8799.n291 98.6054
R23802 a_n9628_8799.n49 a_n9628_8799.n154 81.2902
R23803 a_n9628_8799.n55 a_n9628_8799.n160 81.2902
R23804 a_n9628_8799.n48 a_n9628_8799.n157 81.2902
R23805 a_n9628_8799.n50 a_n9628_8799.n163 80.9324
R23806 a_n9628_8799.n50 a_n9628_8799.n164 80.9324
R23807 a_n9628_8799.n49 a_n9628_8799.n165 80.9324
R23808 a_n9628_8799.n49 a_n9628_8799.n156 80.9324
R23809 a_n9628_8799.n49 a_n9628_8799.n155 80.9324
R23810 a_n9628_8799.n55 a_n9628_8799.n161 80.9324
R23811 a_n9628_8799.n48 a_n9628_8799.n162 80.9324
R23812 a_n9628_8799.n48 a_n9628_8799.n159 80.9324
R23813 a_n9628_8799.n48 a_n9628_8799.n158 80.9324
R23814 a_n9628_8799.n41 a_n9628_8799.n231 70.4033
R23815 a_n9628_8799.n33 a_n9628_8799.n250 70.4033
R23816 a_n9628_8799.n25 a_n9628_8799.n270 70.4033
R23817 a_n9628_8799.n170 a_n9628_8799.n23 70.4033
R23818 a_n9628_8799.n189 a_n9628_8799.n15 70.4033
R23819 a_n9628_8799.n209 a_n9628_8799.n7 70.4033
R23820 a_n9628_8799.n242 a_n9628_8799.n241 48.2005
R23821 a_n9628_8799.n61 a_n9628_8799.n239 20.9683
R23822 a_n9628_8799.n238 a_n9628_8799.n237 48.2005
R23823 a_n9628_8799.n66 a_n9628_8799.n235 20.9683
R23824 a_n9628_8799.n234 a_n9628_8799.n233 48.2005
R23825 a_n9628_8799.n261 a_n9628_8799.n260 48.2005
R23826 a_n9628_8799.n76 a_n9628_8799.n258 20.9683
R23827 a_n9628_8799.n257 a_n9628_8799.n256 48.2005
R23828 a_n9628_8799.n81 a_n9628_8799.n254 20.9683
R23829 a_n9628_8799.n253 a_n9628_8799.n252 48.2005
R23830 a_n9628_8799.n281 a_n9628_8799.n280 48.2005
R23831 a_n9628_8799.n91 a_n9628_8799.n278 20.9683
R23832 a_n9628_8799.n277 a_n9628_8799.n276 48.2005
R23833 a_n9628_8799.n96 a_n9628_8799.n274 20.9683
R23834 a_n9628_8799.n273 a_n9628_8799.n272 48.2005
R23835 a_n9628_8799.n174 a_n9628_8799.n173 48.2005
R23836 a_n9628_8799.n176 a_n9628_8799.n105 20.9683
R23837 a_n9628_8799.n178 a_n9628_8799.n168 48.2005
R23838 a_n9628_8799.n180 a_n9628_8799.n110 20.9683
R23839 a_n9628_8799.n183 a_n9628_8799.n182 48.2005
R23840 a_n9628_8799.t127 a_n9628_8799.n115 485.135
R23841 a_n9628_8799.n193 a_n9628_8799.n192 48.2005
R23842 a_n9628_8799.n195 a_n9628_8799.n120 20.9683
R23843 a_n9628_8799.n197 a_n9628_8799.n187 48.2005
R23844 a_n9628_8799.n199 a_n9628_8799.n125 20.9683
R23845 a_n9628_8799.n202 a_n9628_8799.n201 48.2005
R23846 a_n9628_8799.t141 a_n9628_8799.n130 485.135
R23847 a_n9628_8799.n213 a_n9628_8799.n212 48.2005
R23848 a_n9628_8799.n215 a_n9628_8799.n135 20.9683
R23849 a_n9628_8799.n217 a_n9628_8799.n207 48.2005
R23850 a_n9628_8799.n219 a_n9628_8799.n140 20.9683
R23851 a_n9628_8799.n222 a_n9628_8799.n221 48.2005
R23852 a_n9628_8799.t113 a_n9628_8799.n145 485.135
R23853 a_n9628_8799.n57 a_n9628_8799.n225 17.8606
R23854 a_n9628_8799.n232 a_n9628_8799.n70 25.894
R23855 a_n9628_8799.n72 a_n9628_8799.n244 17.8606
R23856 a_n9628_8799.n251 a_n9628_8799.n85 25.894
R23857 a_n9628_8799.n87 a_n9628_8799.n264 17.8606
R23858 a_n9628_8799.n271 a_n9628_8799.n100 25.894
R23859 a_n9628_8799.n184 a_n9628_8799.n114 25.894
R23860 a_n9628_8799.n203 a_n9628_8799.n129 25.894
R23861 a_n9628_8799.n223 a_n9628_8799.n144 25.894
R23862 a_n9628_8799.n68 a_n9628_8799.n229 43.3183
R23863 a_n9628_8799.n83 a_n9628_8799.n248 43.3183
R23864 a_n9628_8799.n98 a_n9628_8799.n268 43.3183
R23865 a_n9628_8799.n181 a_n9628_8799.n112 43.3183
R23866 a_n9628_8799.n200 a_n9628_8799.n127 43.3183
R23867 a_n9628_8799.n220 a_n9628_8799.n142 43.3183
R23868 a_n9628_8799.n62 a_n9628_8799.n227 16.6962
R23869 a_n9628_8799.n236 a_n9628_8799.n65 27.6507
R23870 a_n9628_8799.n77 a_n9628_8799.n246 16.6962
R23871 a_n9628_8799.n255 a_n9628_8799.n80 27.6507
R23872 a_n9628_8799.n92 a_n9628_8799.n266 16.6962
R23873 a_n9628_8799.n275 a_n9628_8799.n95 27.6507
R23874 a_n9628_8799.n177 a_n9628_8799.n106 16.6962
R23875 a_n9628_8799.n167 a_n9628_8799.n109 27.6507
R23876 a_n9628_8799.n196 a_n9628_8799.n121 16.6962
R23877 a_n9628_8799.n186 a_n9628_8799.n124 27.6507
R23878 a_n9628_8799.n216 a_n9628_8799.n136 16.6962
R23879 a_n9628_8799.n206 a_n9628_8799.n139 27.6507
R23880 a_n9628_8799.n63 a_n9628_8799.n227 41.7634
R23881 a_n9628_8799.n78 a_n9628_8799.n246 41.7634
R23882 a_n9628_8799.n93 a_n9628_8799.n266 41.7634
R23883 a_n9628_8799.n107 a_n9628_8799.n177 41.7634
R23884 a_n9628_8799.n122 a_n9628_8799.n196 41.7634
R23885 a_n9628_8799.n137 a_n9628_8799.n216 41.7634
R23886 a_n9628_8799.n240 a_n9628_8799.n60 29.3885
R23887 a_n9628_8799.n67 a_n9628_8799.n229 15.5127
R23888 a_n9628_8799.n259 a_n9628_8799.n75 29.3885
R23889 a_n9628_8799.n82 a_n9628_8799.n248 15.5127
R23890 a_n9628_8799.n279 a_n9628_8799.n90 29.3885
R23891 a_n9628_8799.n97 a_n9628_8799.n268 15.5127
R23892 a_n9628_8799.n175 a_n9628_8799.n104 29.3885
R23893 a_n9628_8799.n181 a_n9628_8799.n111 15.5127
R23894 a_n9628_8799.n194 a_n9628_8799.n119 29.3885
R23895 a_n9628_8799.n200 a_n9628_8799.n126 15.5127
R23896 a_n9628_8799.n214 a_n9628_8799.n134 29.3885
R23897 a_n9628_8799.n220 a_n9628_8799.n141 15.5127
R23898 a_n9628_8799.n286 a_n9628_8799.n153 33.8967
R23899 a_n9628_8799.n58 a_n9628_8799.n225 40.1848
R23900 a_n9628_8799.n73 a_n9628_8799.n244 40.1848
R23901 a_n9628_8799.n88 a_n9628_8799.n264 40.1848
R23902 a_n9628_8799.n172 a_n9628_8799.n102 40.1848
R23903 a_n9628_8799.n191 a_n9628_8799.n117 40.1848
R23904 a_n9628_8799.n211 a_n9628_8799.n132 40.1848
R23905 a_n9628_8799.n50 a_n9628_8799.n48 32.5134
R23906 a_n9628_8799.n53 a_n9628_8799.n286 20.9925
R23907 a_n9628_8799.n232 a_n9628_8799.n231 20.9576
R23908 a_n9628_8799.n251 a_n9628_8799.n250 20.9576
R23909 a_n9628_8799.n271 a_n9628_8799.n270 20.9576
R23910 a_n9628_8799.n171 a_n9628_8799.n170 20.9576
R23911 a_n9628_8799.n190 a_n9628_8799.n189 20.9576
R23912 a_n9628_8799.n210 a_n9628_8799.n209 20.9576
R23913 a_n9628_8799.n58 a_n9628_8799.n242 7.32118
R23914 a_n9628_8799.n69 a_n9628_8799.n230 40.1848
R23915 a_n9628_8799.n73 a_n9628_8799.n261 7.32118
R23916 a_n9628_8799.n84 a_n9628_8799.n249 40.1848
R23917 a_n9628_8799.n88 a_n9628_8799.n281 7.32118
R23918 a_n9628_8799.n99 a_n9628_8799.n269 40.1848
R23919 a_n9628_8799.n173 a_n9628_8799.n102 7.32118
R23920 a_n9628_8799.n166 a_n9628_8799.n113 40.1848
R23921 a_n9628_8799.n192 a_n9628_8799.n117 7.32118
R23922 a_n9628_8799.n185 a_n9628_8799.n128 40.1848
R23923 a_n9628_8799.n212 a_n9628_8799.n132 7.32118
R23924 a_n9628_8799.n205 a_n9628_8799.n143 40.1848
R23925 a_n9628_8799.n235 a_n9628_8799.n67 29.3885
R23926 a_n9628_8799.n254 a_n9628_8799.n82 29.3885
R23927 a_n9628_8799.n274 a_n9628_8799.n97 29.3885
R23928 a_n9628_8799.n111 a_n9628_8799.n180 29.3885
R23929 a_n9628_8799.n126 a_n9628_8799.n199 29.3885
R23930 a_n9628_8799.n141 a_n9628_8799.n219 29.3885
R23931 a_n9628_8799.n63 a_n9628_8799.n238 5.97853
R23932 a_n9628_8799.n64 a_n9628_8799.n228 41.7634
R23933 a_n9628_8799.n78 a_n9628_8799.n257 5.97853
R23934 a_n9628_8799.n79 a_n9628_8799.n247 41.7634
R23935 a_n9628_8799.n93 a_n9628_8799.n277 5.97853
R23936 a_n9628_8799.n94 a_n9628_8799.n267 41.7634
R23937 a_n9628_8799.n178 a_n9628_8799.n107 5.97853
R23938 a_n9628_8799.n179 a_n9628_8799.n108 41.7634
R23939 a_n9628_8799.n197 a_n9628_8799.n122 5.97853
R23940 a_n9628_8799.n198 a_n9628_8799.n123 41.7634
R23941 a_n9628_8799.n217 a_n9628_8799.n137 5.97853
R23942 a_n9628_8799.n218 a_n9628_8799.n138 41.7634
R23943 a_n9628_8799.n285 a_n9628_8799.n49 12.3339
R23944 a_n9628_8799.n286 a_n9628_8799.n285 11.4887
R23945 a_n9628_8799.n239 a_n9628_8799.n62 27.6507
R23946 a_n9628_8799.n258 a_n9628_8799.n77 27.6507
R23947 a_n9628_8799.n278 a_n9628_8799.n92 27.6507
R23948 a_n9628_8799.n176 a_n9628_8799.n106 27.6507
R23949 a_n9628_8799.n195 a_n9628_8799.n121 27.6507
R23950 a_n9628_8799.n215 a_n9628_8799.n136 27.6507
R23951 a_n9628_8799.n59 a_n9628_8799.n226 43.3183
R23952 a_n9628_8799.n68 a_n9628_8799.n234 4.61226
R23953 a_n9628_8799.n74 a_n9628_8799.n245 43.3183
R23954 a_n9628_8799.n83 a_n9628_8799.n253 4.61226
R23955 a_n9628_8799.n89 a_n9628_8799.n265 43.3183
R23956 a_n9628_8799.n98 a_n9628_8799.n273 4.61226
R23957 a_n9628_8799.n169 a_n9628_8799.n103 43.3183
R23958 a_n9628_8799.n182 a_n9628_8799.n112 4.61226
R23959 a_n9628_8799.n188 a_n9628_8799.n118 43.3183
R23960 a_n9628_8799.n201 a_n9628_8799.n127 4.61226
R23961 a_n9628_8799.n208 a_n9628_8799.n133 43.3183
R23962 a_n9628_8799.n221 a_n9628_8799.n142 4.61226
R23963 a_n9628_8799.n263 a_n9628_8799.n47 9.04406
R23964 a_n9628_8799.n204 a_n9628_8799.n17 9.04406
R23965 a_n9628_8799.n243 a_n9628_8799.n57 25.894
R23966 a_n9628_8799.n262 a_n9628_8799.n72 25.894
R23967 a_n9628_8799.n282 a_n9628_8799.n87 25.894
R23968 a_n9628_8799.n101 a_n9628_8799.n171 25.894
R23969 a_n9628_8799.n116 a_n9628_8799.n190 25.894
R23970 a_n9628_8799.n131 a_n9628_8799.n210 25.894
R23971 a_n9628_8799.n284 a_n9628_8799.n224 7.1766
R23972 a_n9628_8799.n284 a_n9628_8799.n283 6.83037
R23973 a_n9628_8799.n263 a_n9628_8799.n39 4.93611
R23974 a_n9628_8799.n283 a_n9628_8799.n31 4.93611
R23975 a_n9628_8799.n204 a_n9628_8799.n9 4.93611
R23976 a_n9628_8799.n224 a_n9628_8799.n1 4.93611
R23977 a_n9628_8799.n283 a_n9628_8799.n263 4.10845
R23978 a_n9628_8799.n224 a_n9628_8799.n204 4.10845
R23979 a_n9628_8799.n287 a_n9628_8799.t32 3.61217
R23980 a_n9628_8799.n287 a_n9628_8799.t37 3.61217
R23981 a_n9628_8799.n288 a_n9628_8799.t33 3.61217
R23982 a_n9628_8799.n288 a_n9628_8799.t26 3.61217
R23983 a_n9628_8799.n289 a_n9628_8799.t43 3.61217
R23984 a_n9628_8799.n289 a_n9628_8799.t23 3.61217
R23985 a_n9628_8799.n290 a_n9628_8799.t36 3.61217
R23986 a_n9628_8799.n290 a_n9628_8799.t44 3.61217
R23987 a_n9628_8799.n146 a_n9628_8799.t41 3.61217
R23988 a_n9628_8799.n146 a_n9628_8799.t34 3.61217
R23989 a_n9628_8799.n147 a_n9628_8799.t27 3.61217
R23990 a_n9628_8799.n147 a_n9628_8799.t30 3.61217
R23991 a_n9628_8799.n148 a_n9628_8799.t24 3.61217
R23992 a_n9628_8799.n148 a_n9628_8799.t31 3.61217
R23993 a_n9628_8799.n149 a_n9628_8799.t35 3.61217
R23994 a_n9628_8799.n149 a_n9628_8799.t38 3.61217
R23995 a_n9628_8799.n150 a_n9628_8799.t39 3.61217
R23996 a_n9628_8799.n150 a_n9628_8799.t29 3.61217
R23997 a_n9628_8799.n151 a_n9628_8799.t22 3.61217
R23998 a_n9628_8799.n151 a_n9628_8799.t40 3.61217
R23999 a_n9628_8799.n152 a_n9628_8799.t42 3.61217
R24000 a_n9628_8799.n152 a_n9628_8799.t25 3.61217
R24001 a_n9628_8799.n292 a_n9628_8799.t28 3.61217
R24002 a_n9628_8799.t21 a_n9628_8799.n292 3.61217
R24003 a_n9628_8799.n285 a_n9628_8799.n284 3.4105
R24004 a_n9628_8799.n163 a_n9628_8799.t16 2.82907
R24005 a_n9628_8799.n163 a_n9628_8799.t18 2.82907
R24006 a_n9628_8799.n164 a_n9628_8799.t13 2.82907
R24007 a_n9628_8799.n164 a_n9628_8799.t14 2.82907
R24008 a_n9628_8799.n165 a_n9628_8799.t7 2.82907
R24009 a_n9628_8799.n165 a_n9628_8799.t8 2.82907
R24010 a_n9628_8799.n156 a_n9628_8799.t4 2.82907
R24011 a_n9628_8799.n156 a_n9628_8799.t6 2.82907
R24012 a_n9628_8799.n155 a_n9628_8799.t5 2.82907
R24013 a_n9628_8799.n155 a_n9628_8799.t15 2.82907
R24014 a_n9628_8799.n154 a_n9628_8799.t19 2.82907
R24015 a_n9628_8799.n154 a_n9628_8799.t47 2.82907
R24016 a_n9628_8799.n160 a_n9628_8799.t12 2.82907
R24017 a_n9628_8799.n160 a_n9628_8799.t17 2.82907
R24018 a_n9628_8799.n161 a_n9628_8799.t1 2.82907
R24019 a_n9628_8799.n161 a_n9628_8799.t0 2.82907
R24020 a_n9628_8799.n162 a_n9628_8799.t45 2.82907
R24021 a_n9628_8799.n162 a_n9628_8799.t9 2.82907
R24022 a_n9628_8799.n159 a_n9628_8799.t11 2.82907
R24023 a_n9628_8799.n159 a_n9628_8799.t2 2.82907
R24024 a_n9628_8799.n158 a_n9628_8799.t3 2.82907
R24025 a_n9628_8799.n158 a_n9628_8799.t46 2.82907
R24026 a_n9628_8799.n157 a_n9628_8799.t20 2.82907
R24027 a_n9628_8799.n157 a_n9628_8799.t10 2.82907
R24028 a_n9628_8799.n49 a_n9628_8799.n50 1.43153
R24029 a_n9628_8799.n41 a_n9628_8799.n40 1.13686
R24030 a_n9628_8799.n33 a_n9628_8799.n32 1.13686
R24031 a_n9628_8799.n25 a_n9628_8799.n24 1.13686
R24032 a_n9628_8799.n17 a_n9628_8799.n16 1.13686
R24033 a_n9628_8799.n9 a_n9628_8799.n8 1.13686
R24034 a_n9628_8799.n1 a_n9628_8799.n0 1.13686
R24035 a_n9628_8799.n48 a_n9628_8799.n55 1.07378
R24036 a_n9628_8799.n46 a_n9628_8799.n45 0.758076
R24037 a_n9628_8799.n46 a_n9628_8799.n44 0.758076
R24038 a_n9628_8799.n44 a_n9628_8799.n43 0.758076
R24039 a_n9628_8799.n43 a_n9628_8799.n42 0.758076
R24040 a_n9628_8799.n40 a_n9628_8799.n42 0.758076
R24041 a_n9628_8799.n38 a_n9628_8799.n37 0.758076
R24042 a_n9628_8799.n38 a_n9628_8799.n36 0.758076
R24043 a_n9628_8799.n36 a_n9628_8799.n35 0.758076
R24044 a_n9628_8799.n35 a_n9628_8799.n34 0.758076
R24045 a_n9628_8799.n32 a_n9628_8799.n34 0.758076
R24046 a_n9628_8799.n30 a_n9628_8799.n29 0.758076
R24047 a_n9628_8799.n30 a_n9628_8799.n28 0.758076
R24048 a_n9628_8799.n28 a_n9628_8799.n27 0.758076
R24049 a_n9628_8799.n27 a_n9628_8799.n26 0.758076
R24050 a_n9628_8799.n24 a_n9628_8799.n26 0.758076
R24051 a_n9628_8799.n21 a_n9628_8799.n22 0.758076
R24052 a_n9628_8799.n20 a_n9628_8799.n21 0.758076
R24053 a_n9628_8799.n19 a_n9628_8799.n20 0.758076
R24054 a_n9628_8799.n18 a_n9628_8799.n19 0.758076
R24055 a_n9628_8799.n16 a_n9628_8799.n18 0.758076
R24056 a_n9628_8799.n13 a_n9628_8799.n14 0.758076
R24057 a_n9628_8799.n12 a_n9628_8799.n13 0.758076
R24058 a_n9628_8799.n11 a_n9628_8799.n12 0.758076
R24059 a_n9628_8799.n10 a_n9628_8799.n11 0.758076
R24060 a_n9628_8799.n8 a_n9628_8799.n10 0.758076
R24061 a_n9628_8799.n5 a_n9628_8799.n6 0.758076
R24062 a_n9628_8799.n4 a_n9628_8799.n5 0.758076
R24063 a_n9628_8799.n3 a_n9628_8799.n4 0.758076
R24064 a_n9628_8799.n2 a_n9628_8799.n3 0.758076
R24065 a_n9628_8799.n0 a_n9628_8799.n2 0.758076
R24066 a_n9628_8799.n54 a_n9628_8799.n53 0.716017
R24067 a_n9628_8799.n291 a_n9628_8799.n54 0.716017
R24068 a_n9628_8799.n52 a_n9628_8799.n51 0.716017
R24069 a_n9628_8799.n153 a_n9628_8799.n52 0.716017
R24070 a_n9628_8799.n6 a_n9628_8799.n7 0.568682
R24071 a_n9628_8799.n14 a_n9628_8799.n15 0.568682
R24072 a_n9628_8799.n22 a_n9628_8799.n23 0.568682
R24073 a_n9628_8799.n29 a_n9628_8799.n31 0.568682
R24074 a_n9628_8799.n37 a_n9628_8799.n39 0.568682
R24075 a_n9628_8799.n45 a_n9628_8799.n47 0.568682
R24076 a_n2982_8322.n12 a_n2982_8322.t33 74.6477
R24077 a_n2982_8322.n1 a_n2982_8322.t12 74.6477
R24078 a_n2982_8322.n28 a_n2982_8322.t27 74.6474
R24079 a_n2982_8322.n20 a_n2982_8322.t7 74.2899
R24080 a_n2982_8322.n13 a_n2982_8322.t31 74.2899
R24081 a_n2982_8322.n14 a_n2982_8322.t34 74.2899
R24082 a_n2982_8322.n17 a_n2982_8322.t35 74.2899
R24083 a_n2982_8322.n10 a_n2982_8322.t6 74.2899
R24084 a_n2982_8322.n28 a_n2982_8322.n27 70.6783
R24085 a_n2982_8322.n26 a_n2982_8322.n25 70.6783
R24086 a_n2982_8322.n24 a_n2982_8322.n23 70.6783
R24087 a_n2982_8322.n22 a_n2982_8322.n21 70.6783
R24088 a_n2982_8322.n12 a_n2982_8322.n11 70.6783
R24089 a_n2982_8322.n16 a_n2982_8322.n15 70.6783
R24090 a_n2982_8322.n1 a_n2982_8322.n0 70.6783
R24091 a_n2982_8322.n3 a_n2982_8322.n2 70.6783
R24092 a_n2982_8322.n5 a_n2982_8322.n4 70.6783
R24093 a_n2982_8322.n7 a_n2982_8322.n6 70.6783
R24094 a_n2982_8322.n9 a_n2982_8322.n8 70.6783
R24095 a_n2982_8322.n30 a_n2982_8322.n29 70.6782
R24096 a_n2982_8322.n18 a_n2982_8322.n10 24.9022
R24097 a_n2982_8322.n19 a_n2982_8322.t0 9.69161
R24098 a_n2982_8322.n18 a_n2982_8322.n17 8.38735
R24099 a_n2982_8322.n20 a_n2982_8322.n19 6.90998
R24100 a_n2982_8322.n19 a_n2982_8322.n18 5.3452
R24101 a_n2982_8322.n27 a_n2982_8322.t20 3.61217
R24102 a_n2982_8322.n27 a_n2982_8322.t16 3.61217
R24103 a_n2982_8322.n25 a_n2982_8322.t26 3.61217
R24104 a_n2982_8322.n25 a_n2982_8322.t14 3.61217
R24105 a_n2982_8322.n23 a_n2982_8322.t11 3.61217
R24106 a_n2982_8322.n23 a_n2982_8322.t10 3.61217
R24107 a_n2982_8322.n21 a_n2982_8322.t24 3.61217
R24108 a_n2982_8322.n21 a_n2982_8322.t23 3.61217
R24109 a_n2982_8322.n11 a_n2982_8322.t37 3.61217
R24110 a_n2982_8322.n11 a_n2982_8322.t36 3.61217
R24111 a_n2982_8322.n15 a_n2982_8322.t32 3.61217
R24112 a_n2982_8322.n15 a_n2982_8322.t30 3.61217
R24113 a_n2982_8322.n0 a_n2982_8322.t25 3.61217
R24114 a_n2982_8322.n0 a_n2982_8322.t21 3.61217
R24115 a_n2982_8322.n2 a_n2982_8322.t28 3.61217
R24116 a_n2982_8322.n2 a_n2982_8322.t18 3.61217
R24117 a_n2982_8322.n4 a_n2982_8322.t9 3.61217
R24118 a_n2982_8322.n4 a_n2982_8322.t8 3.61217
R24119 a_n2982_8322.n6 a_n2982_8322.t22 3.61217
R24120 a_n2982_8322.n6 a_n2982_8322.t15 3.61217
R24121 a_n2982_8322.n8 a_n2982_8322.t19 3.61217
R24122 a_n2982_8322.n8 a_n2982_8322.t17 3.61217
R24123 a_n2982_8322.n30 a_n2982_8322.t13 3.61217
R24124 a_n2982_8322.t29 a_n2982_8322.n30 3.61217
R24125 a_n2982_8322.n17 a_n2982_8322.n16 0.358259
R24126 a_n2982_8322.n16 a_n2982_8322.n14 0.358259
R24127 a_n2982_8322.n13 a_n2982_8322.n12 0.358259
R24128 a_n2982_8322.n10 a_n2982_8322.n9 0.358259
R24129 a_n2982_8322.n9 a_n2982_8322.n7 0.358259
R24130 a_n2982_8322.n7 a_n2982_8322.n5 0.358259
R24131 a_n2982_8322.n5 a_n2982_8322.n3 0.358259
R24132 a_n2982_8322.n3 a_n2982_8322.n1 0.358259
R24133 a_n2982_8322.n22 a_n2982_8322.n20 0.358259
R24134 a_n2982_8322.n24 a_n2982_8322.n22 0.358259
R24135 a_n2982_8322.n26 a_n2982_8322.n24 0.358259
R24136 a_n2982_8322.n29 a_n2982_8322.n26 0.358259
R24137 a_n2982_8322.n29 a_n2982_8322.n28 0.358259
R24138 a_n2982_8322.n14 a_n2982_8322.n13 0.101793
R24139 a_n2982_8322.t5 a_n2982_8322.t1 0.0788333
R24140 a_n2982_8322.t4 a_n2982_8322.t2 0.0788333
R24141 a_n2982_8322.t0 a_n2982_8322.t3 0.0788333
R24142 a_n2982_8322.t4 a_n2982_8322.t5 0.0318333
R24143 a_n2982_8322.t0 a_n2982_8322.t2 0.0318333
R24144 a_n2982_8322.t1 a_n2982_8322.t2 0.0318333
R24145 a_n2982_8322.t3 a_n2982_8322.t4 0.0318333
R24146 output.n41 output.n15 289.615
R24147 output.n72 output.n46 289.615
R24148 output.n104 output.n78 289.615
R24149 output.n136 output.n110 289.615
R24150 output.n77 output.n45 197.26
R24151 output.n77 output.n76 196.298
R24152 output.n109 output.n108 196.298
R24153 output.n141 output.n140 196.298
R24154 output.n42 output.n41 185
R24155 output.n40 output.n39 185
R24156 output.n19 output.n18 185
R24157 output.n34 output.n33 185
R24158 output.n32 output.n31 185
R24159 output.n23 output.n22 185
R24160 output.n26 output.n25 185
R24161 output.n73 output.n72 185
R24162 output.n71 output.n70 185
R24163 output.n50 output.n49 185
R24164 output.n65 output.n64 185
R24165 output.n63 output.n62 185
R24166 output.n54 output.n53 185
R24167 output.n57 output.n56 185
R24168 output.n105 output.n104 185
R24169 output.n103 output.n102 185
R24170 output.n82 output.n81 185
R24171 output.n97 output.n96 185
R24172 output.n95 output.n94 185
R24173 output.n86 output.n85 185
R24174 output.n89 output.n88 185
R24175 output.n137 output.n136 185
R24176 output.n135 output.n134 185
R24177 output.n114 output.n113 185
R24178 output.n129 output.n128 185
R24179 output.n127 output.n126 185
R24180 output.n118 output.n117 185
R24181 output.n121 output.n120 185
R24182 output.t19 output.n24 147.661
R24183 output.t18 output.n55 147.661
R24184 output.t16 output.n87 147.661
R24185 output.t17 output.n119 147.661
R24186 output.n41 output.n40 104.615
R24187 output.n40 output.n18 104.615
R24188 output.n33 output.n18 104.615
R24189 output.n33 output.n32 104.615
R24190 output.n32 output.n22 104.615
R24191 output.n25 output.n22 104.615
R24192 output.n72 output.n71 104.615
R24193 output.n71 output.n49 104.615
R24194 output.n64 output.n49 104.615
R24195 output.n64 output.n63 104.615
R24196 output.n63 output.n53 104.615
R24197 output.n56 output.n53 104.615
R24198 output.n104 output.n103 104.615
R24199 output.n103 output.n81 104.615
R24200 output.n96 output.n81 104.615
R24201 output.n96 output.n95 104.615
R24202 output.n95 output.n85 104.615
R24203 output.n88 output.n85 104.615
R24204 output.n136 output.n135 104.615
R24205 output.n135 output.n113 104.615
R24206 output.n128 output.n113 104.615
R24207 output.n128 output.n127 104.615
R24208 output.n127 output.n117 104.615
R24209 output.n120 output.n117 104.615
R24210 output.n1 output.t13 77.056
R24211 output.n14 output.t15 76.6694
R24212 output.n1 output.n0 72.7095
R24213 output.n3 output.n2 72.7095
R24214 output.n5 output.n4 72.7095
R24215 output.n7 output.n6 72.7095
R24216 output.n9 output.n8 72.7095
R24217 output.n11 output.n10 72.7095
R24218 output.n13 output.n12 72.7095
R24219 output.n25 output.t19 52.3082
R24220 output.n56 output.t18 52.3082
R24221 output.n88 output.t16 52.3082
R24222 output.n120 output.t17 52.3082
R24223 output.n26 output.n24 15.6674
R24224 output.n57 output.n55 15.6674
R24225 output.n89 output.n87 15.6674
R24226 output.n121 output.n119 15.6674
R24227 output.n27 output.n23 12.8005
R24228 output.n58 output.n54 12.8005
R24229 output.n90 output.n86 12.8005
R24230 output.n122 output.n118 12.8005
R24231 output.n31 output.n30 12.0247
R24232 output.n62 output.n61 12.0247
R24233 output.n94 output.n93 12.0247
R24234 output.n126 output.n125 12.0247
R24235 output.n34 output.n21 11.249
R24236 output.n65 output.n52 11.249
R24237 output.n97 output.n84 11.249
R24238 output.n129 output.n116 11.249
R24239 output.n35 output.n19 10.4732
R24240 output.n66 output.n50 10.4732
R24241 output.n98 output.n82 10.4732
R24242 output.n130 output.n114 10.4732
R24243 output.n39 output.n38 9.69747
R24244 output.n70 output.n69 9.69747
R24245 output.n102 output.n101 9.69747
R24246 output.n134 output.n133 9.69747
R24247 output.n45 output.n44 9.45567
R24248 output.n76 output.n75 9.45567
R24249 output.n108 output.n107 9.45567
R24250 output.n140 output.n139 9.45567
R24251 output.n44 output.n43 9.3005
R24252 output.n17 output.n16 9.3005
R24253 output.n38 output.n37 9.3005
R24254 output.n36 output.n35 9.3005
R24255 output.n21 output.n20 9.3005
R24256 output.n30 output.n29 9.3005
R24257 output.n28 output.n27 9.3005
R24258 output.n75 output.n74 9.3005
R24259 output.n48 output.n47 9.3005
R24260 output.n69 output.n68 9.3005
R24261 output.n67 output.n66 9.3005
R24262 output.n52 output.n51 9.3005
R24263 output.n61 output.n60 9.3005
R24264 output.n59 output.n58 9.3005
R24265 output.n107 output.n106 9.3005
R24266 output.n80 output.n79 9.3005
R24267 output.n101 output.n100 9.3005
R24268 output.n99 output.n98 9.3005
R24269 output.n84 output.n83 9.3005
R24270 output.n93 output.n92 9.3005
R24271 output.n91 output.n90 9.3005
R24272 output.n139 output.n138 9.3005
R24273 output.n112 output.n111 9.3005
R24274 output.n133 output.n132 9.3005
R24275 output.n131 output.n130 9.3005
R24276 output.n116 output.n115 9.3005
R24277 output.n125 output.n124 9.3005
R24278 output.n123 output.n122 9.3005
R24279 output.n42 output.n17 8.92171
R24280 output.n73 output.n48 8.92171
R24281 output.n105 output.n80 8.92171
R24282 output.n137 output.n112 8.92171
R24283 output output.n141 8.15037
R24284 output.n43 output.n15 8.14595
R24285 output.n74 output.n46 8.14595
R24286 output.n106 output.n78 8.14595
R24287 output.n138 output.n110 8.14595
R24288 output.n45 output.n15 5.81868
R24289 output.n76 output.n46 5.81868
R24290 output.n108 output.n78 5.81868
R24291 output.n140 output.n110 5.81868
R24292 output.n43 output.n42 5.04292
R24293 output.n74 output.n73 5.04292
R24294 output.n106 output.n105 5.04292
R24295 output.n138 output.n137 5.04292
R24296 output.n28 output.n24 4.38594
R24297 output.n59 output.n55 4.38594
R24298 output.n91 output.n87 4.38594
R24299 output.n123 output.n119 4.38594
R24300 output.n39 output.n17 4.26717
R24301 output.n70 output.n48 4.26717
R24302 output.n102 output.n80 4.26717
R24303 output.n134 output.n112 4.26717
R24304 output.n0 output.t9 3.9605
R24305 output.n0 output.t7 3.9605
R24306 output.n2 output.t1 3.9605
R24307 output.n2 output.t3 3.9605
R24308 output.n4 output.t4 3.9605
R24309 output.n4 output.t11 3.9605
R24310 output.n6 output.t14 3.9605
R24311 output.n6 output.t2 3.9605
R24312 output.n8 output.t5 3.9605
R24313 output.n8 output.t10 3.9605
R24314 output.n10 output.t12 3.9605
R24315 output.n10 output.t0 3.9605
R24316 output.n12 output.t8 3.9605
R24317 output.n12 output.t6 3.9605
R24318 output.n38 output.n19 3.49141
R24319 output.n69 output.n50 3.49141
R24320 output.n101 output.n82 3.49141
R24321 output.n133 output.n114 3.49141
R24322 output.n35 output.n34 2.71565
R24323 output.n66 output.n65 2.71565
R24324 output.n98 output.n97 2.71565
R24325 output.n130 output.n129 2.71565
R24326 output.n31 output.n21 1.93989
R24327 output.n62 output.n52 1.93989
R24328 output.n94 output.n84 1.93989
R24329 output.n126 output.n116 1.93989
R24330 output.n30 output.n23 1.16414
R24331 output.n61 output.n54 1.16414
R24332 output.n93 output.n86 1.16414
R24333 output.n125 output.n118 1.16414
R24334 output.n141 output.n109 0.962709
R24335 output.n109 output.n77 0.962709
R24336 output.n27 output.n26 0.388379
R24337 output.n58 output.n57 0.388379
R24338 output.n90 output.n89 0.388379
R24339 output.n122 output.n121 0.388379
R24340 output.n14 output.n13 0.387128
R24341 output.n13 output.n11 0.387128
R24342 output.n11 output.n9 0.387128
R24343 output.n9 output.n7 0.387128
R24344 output.n7 output.n5 0.387128
R24345 output.n5 output.n3 0.387128
R24346 output.n3 output.n1 0.387128
R24347 output.n44 output.n16 0.155672
R24348 output.n37 output.n16 0.155672
R24349 output.n37 output.n36 0.155672
R24350 output.n36 output.n20 0.155672
R24351 output.n29 output.n20 0.155672
R24352 output.n29 output.n28 0.155672
R24353 output.n75 output.n47 0.155672
R24354 output.n68 output.n47 0.155672
R24355 output.n68 output.n67 0.155672
R24356 output.n67 output.n51 0.155672
R24357 output.n60 output.n51 0.155672
R24358 output.n60 output.n59 0.155672
R24359 output.n107 output.n79 0.155672
R24360 output.n100 output.n79 0.155672
R24361 output.n100 output.n99 0.155672
R24362 output.n99 output.n83 0.155672
R24363 output.n92 output.n83 0.155672
R24364 output.n92 output.n91 0.155672
R24365 output.n139 output.n111 0.155672
R24366 output.n132 output.n111 0.155672
R24367 output.n132 output.n131 0.155672
R24368 output.n131 output.n115 0.155672
R24369 output.n124 output.n115 0.155672
R24370 output.n124 output.n123 0.155672
R24371 output output.n14 0.126227
R24372 plus.n43 plus.t25 442.325
R24373 plus.n11 plus.t12 442.325
R24374 plus.n42 plus.t5 415.966
R24375 plus.n41 plus.t20 415.966
R24376 plus.n47 plus.t26 415.966
R24377 plus.n39 plus.t11 415.966
R24378 plus.n52 plus.t6 415.966
R24379 plus.n54 plus.t10 415.966
R24380 plus.n37 plus.t19 415.966
R24381 plus.n59 plus.t8 415.966
R24382 plus.n35 plus.t16 415.966
R24383 plus.n64 plus.t28 415.966
R24384 plus.n66 plus.t21 415.966
R24385 plus.n32 plus.t23 415.966
R24386 plus.n30 plus.t13 415.966
R24387 plus.n29 plus.t27 415.966
R24388 plus.n3 plus.t22 415.966
R24389 plus.n23 plus.t7 415.966
R24390 plus.n22 plus.t18 415.966
R24391 plus.n6 plus.t14 415.966
R24392 plus.n17 plus.t24 415.966
R24393 plus.n15 plus.t17 415.966
R24394 plus.n9 plus.t9 415.966
R24395 plus.n10 plus.t15 415.966
R24396 plus.n70 plus.t3 243.97
R24397 plus.n70 plus.n69 223.454
R24398 plus.n72 plus.n71 223.454
R24399 plus.n67 plus.n66 161.3
R24400 plus.n65 plus.n34 161.3
R24401 plus.n64 plus.n63 161.3
R24402 plus.n62 plus.n35 161.3
R24403 plus.n61 plus.n60 161.3
R24404 plus.n59 plus.n36 161.3
R24405 plus.n58 plus.n57 161.3
R24406 plus.n56 plus.n37 161.3
R24407 plus.n55 plus.n54 161.3
R24408 plus.n53 plus.n38 161.3
R24409 plus.n52 plus.n51 161.3
R24410 plus.n50 plus.n39 161.3
R24411 plus.n49 plus.n48 161.3
R24412 plus.n47 plus.n40 161.3
R24413 plus.n46 plus.n45 161.3
R24414 plus.n44 plus.n41 161.3
R24415 plus.n12 plus.n9 161.3
R24416 plus.n14 plus.n13 161.3
R24417 plus.n15 plus.n8 161.3
R24418 plus.n16 plus.n7 161.3
R24419 plus.n18 plus.n17 161.3
R24420 plus.n19 plus.n6 161.3
R24421 plus.n21 plus.n20 161.3
R24422 plus.n22 plus.n5 161.3
R24423 plus.n23 plus.n4 161.3
R24424 plus.n25 plus.n24 161.3
R24425 plus.n26 plus.n3 161.3
R24426 plus.n28 plus.n27 161.3
R24427 plus.n29 plus.n2 161.3
R24428 plus.n30 plus.n1 161.3
R24429 plus.n31 plus.n0 161.3
R24430 plus.n33 plus.n32 161.3
R24431 plus.n42 plus.n41 48.2005
R24432 plus.n52 plus.n39 48.2005
R24433 plus.n54 plus.n37 48.2005
R24434 plus.n64 plus.n35 48.2005
R24435 plus.n30 plus.n29 48.2005
R24436 plus.n23 plus.n22 48.2005
R24437 plus.n17 plus.n6 48.2005
R24438 plus.n10 plus.n9 48.2005
R24439 plus.n48 plus.n47 47.4702
R24440 plus.n59 plus.n58 47.4702
R24441 plus.n24 plus.n3 47.4702
R24442 plus.n16 plus.n15 47.4702
R24443 plus.n66 plus.n65 46.0096
R24444 plus.n32 plus.n31 46.0096
R24445 plus.n44 plus.n43 45.0871
R24446 plus.n12 plus.n11 45.0871
R24447 plus.n68 plus.n67 31.0554
R24448 plus.n47 plus.n46 25.5611
R24449 plus.n60 plus.n59 25.5611
R24450 plus.n28 plus.n3 25.5611
R24451 plus.n15 plus.n14 25.5611
R24452 plus.n53 plus.n52 24.1005
R24453 plus.n54 plus.n53 24.1005
R24454 plus.n22 plus.n21 24.1005
R24455 plus.n21 plus.n6 24.1005
R24456 plus.n46 plus.n41 22.6399
R24457 plus.n60 plus.n35 22.6399
R24458 plus.n29 plus.n28 22.6399
R24459 plus.n14 plus.n9 22.6399
R24460 plus.n69 plus.t4 19.8005
R24461 plus.n69 plus.t1 19.8005
R24462 plus.n71 plus.t0 19.8005
R24463 plus.n71 plus.t2 19.8005
R24464 plus plus.n73 14.4906
R24465 plus.n43 plus.n42 14.1472
R24466 plus.n11 plus.n10 14.1472
R24467 plus.n68 plus.n33 11.7259
R24468 plus.n73 plus.n72 5.40567
R24469 plus.n65 plus.n64 2.19141
R24470 plus.n31 plus.n30 2.19141
R24471 plus.n73 plus.n68 1.188
R24472 plus.n48 plus.n39 0.730803
R24473 plus.n58 plus.n37 0.730803
R24474 plus.n24 plus.n23 0.730803
R24475 plus.n17 plus.n16 0.730803
R24476 plus.n72 plus.n70 0.716017
R24477 plus.n45 plus.n44 0.189894
R24478 plus.n45 plus.n40 0.189894
R24479 plus.n49 plus.n40 0.189894
R24480 plus.n50 plus.n49 0.189894
R24481 plus.n51 plus.n50 0.189894
R24482 plus.n51 plus.n38 0.189894
R24483 plus.n55 plus.n38 0.189894
R24484 plus.n56 plus.n55 0.189894
R24485 plus.n57 plus.n56 0.189894
R24486 plus.n57 plus.n36 0.189894
R24487 plus.n61 plus.n36 0.189894
R24488 plus.n62 plus.n61 0.189894
R24489 plus.n63 plus.n62 0.189894
R24490 plus.n63 plus.n34 0.189894
R24491 plus.n67 plus.n34 0.189894
R24492 plus.n33 plus.n0 0.189894
R24493 plus.n1 plus.n0 0.189894
R24494 plus.n2 plus.n1 0.189894
R24495 plus.n27 plus.n2 0.189894
R24496 plus.n27 plus.n26 0.189894
R24497 plus.n26 plus.n25 0.189894
R24498 plus.n25 plus.n4 0.189894
R24499 plus.n5 plus.n4 0.189894
R24500 plus.n20 plus.n5 0.189894
R24501 plus.n20 plus.n19 0.189894
R24502 plus.n19 plus.n18 0.189894
R24503 plus.n18 plus.n7 0.189894
R24504 plus.n8 plus.n7 0.189894
R24505 plus.n13 plus.n8 0.189894
R24506 plus.n13 plus.n12 0.189894
R24507 a_n2903_n3924.n14 a_n2903_n3924.t3 214.994
R24508 a_n2903_n3924.n1 a_n2903_n3924.t51 214.493
R24509 a_n2903_n3924.n15 a_n2903_n3924.t7 214.321
R24510 a_n2903_n3924.n16 a_n2903_n3924.t36 214.321
R24511 a_n2903_n3924.n17 a_n2903_n3924.t5 214.321
R24512 a_n2903_n3924.n18 a_n2903_n3924.t43 214.321
R24513 a_n2903_n3924.n19 a_n2903_n3924.t50 214.321
R24514 a_n2903_n3924.n14 a_n2903_n3924.t0 214.321
R24515 a_n2903_n3924.n0 a_n2903_n3924.t13 55.8337
R24516 a_n2903_n3924.n2 a_n2903_n3924.t37 55.8337
R24517 a_n2903_n3924.n13 a_n2903_n3924.t38 55.8337
R24518 a_n2903_n3924.n47 a_n2903_n3924.t17 55.8335
R24519 a_n2903_n3924.n45 a_n2903_n3924.t1 55.8335
R24520 a_n2903_n3924.n34 a_n2903_n3924.t53 55.8335
R24521 a_n2903_n3924.n33 a_n2903_n3924.t26 55.8335
R24522 a_n2903_n3924.n22 a_n2903_n3924.t15 55.8335
R24523 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0052
R24524 a_n2903_n3924.n51 a_n2903_n3924.n50 53.0052
R24525 a_n2903_n3924.n53 a_n2903_n3924.n52 53.0052
R24526 a_n2903_n3924.n55 a_n2903_n3924.n54 53.0052
R24527 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R24528 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R24529 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R24530 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R24531 a_n2903_n3924.n12 a_n2903_n3924.n11 53.0052
R24532 a_n2903_n3924.n44 a_n2903_n3924.n43 53.0051
R24533 a_n2903_n3924.n42 a_n2903_n3924.n41 53.0051
R24534 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R24535 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R24536 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R24537 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R24538 a_n2903_n3924.n30 a_n2903_n3924.n29 53.0051
R24539 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R24540 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R24541 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R24542 a_n2903_n3924.n57 a_n2903_n3924.n56 53.0051
R24543 a_n2903_n3924.n21 a_n2903_n3924.n13 12.1555
R24544 a_n2903_n3924.n47 a_n2903_n3924.n46 12.1555
R24545 a_n2903_n3924.n22 a_n2903_n3924.n21 5.07593
R24546 a_n2903_n3924.n46 a_n2903_n3924.n45 5.07593
R24547 a_n2903_n3924.n48 a_n2903_n3924.t22 2.82907
R24548 a_n2903_n3924.n48 a_n2903_n3924.t10 2.82907
R24549 a_n2903_n3924.n50 a_n2903_n3924.t19 2.82907
R24550 a_n2903_n3924.n50 a_n2903_n3924.t30 2.82907
R24551 a_n2903_n3924.n52 a_n2903_n3924.t32 2.82907
R24552 a_n2903_n3924.n52 a_n2903_n3924.t28 2.82907
R24553 a_n2903_n3924.n54 a_n2903_n3924.t12 2.82907
R24554 a_n2903_n3924.n54 a_n2903_n3924.t27 2.82907
R24555 a_n2903_n3924.n3 a_n2903_n3924.t39 2.82907
R24556 a_n2903_n3924.n3 a_n2903_n3924.t49 2.82907
R24557 a_n2903_n3924.n5 a_n2903_n3924.t52 2.82907
R24558 a_n2903_n3924.n5 a_n2903_n3924.t48 2.82907
R24559 a_n2903_n3924.n7 a_n2903_n3924.t40 2.82907
R24560 a_n2903_n3924.n7 a_n2903_n3924.t2 2.82907
R24561 a_n2903_n3924.n9 a_n2903_n3924.t34 2.82907
R24562 a_n2903_n3924.n9 a_n2903_n3924.t46 2.82907
R24563 a_n2903_n3924.n11 a_n2903_n3924.t54 2.82907
R24564 a_n2903_n3924.n11 a_n2903_n3924.t4 2.82907
R24565 a_n2903_n3924.n43 a_n2903_n3924.t44 2.82907
R24566 a_n2903_n3924.n43 a_n2903_n3924.t35 2.82907
R24567 a_n2903_n3924.n41 a_n2903_n3924.t42 2.82907
R24568 a_n2903_n3924.n41 a_n2903_n3924.t55 2.82907
R24569 a_n2903_n3924.n39 a_n2903_n3924.t6 2.82907
R24570 a_n2903_n3924.n39 a_n2903_n3924.t47 2.82907
R24571 a_n2903_n3924.n37 a_n2903_n3924.t8 2.82907
R24572 a_n2903_n3924.n37 a_n2903_n3924.t41 2.82907
R24573 a_n2903_n3924.n35 a_n2903_n3924.t45 2.82907
R24574 a_n2903_n3924.n35 a_n2903_n3924.t9 2.82907
R24575 a_n2903_n3924.n31 a_n2903_n3924.t29 2.82907
R24576 a_n2903_n3924.n31 a_n2903_n3924.t23 2.82907
R24577 a_n2903_n3924.n29 a_n2903_n3924.t14 2.82907
R24578 a_n2903_n3924.n29 a_n2903_n3924.t21 2.82907
R24579 a_n2903_n3924.n27 a_n2903_n3924.t20 2.82907
R24580 a_n2903_n3924.n27 a_n2903_n3924.t24 2.82907
R24581 a_n2903_n3924.n25 a_n2903_n3924.t16 2.82907
R24582 a_n2903_n3924.n25 a_n2903_n3924.t31 2.82907
R24583 a_n2903_n3924.n23 a_n2903_n3924.t25 2.82907
R24584 a_n2903_n3924.n23 a_n2903_n3924.t11 2.82907
R24585 a_n2903_n3924.t33 a_n2903_n3924.n57 2.82907
R24586 a_n2903_n3924.n57 a_n2903_n3924.t18 2.82907
R24587 a_n2903_n3924.n46 a_n2903_n3924.n1 1.95694
R24588 a_n2903_n3924.n21 a_n2903_n3924.n20 1.95694
R24589 a_n2903_n3924.n19 a_n2903_n3924.n18 0.672012
R24590 a_n2903_n3924.n18 a_n2903_n3924.n17 0.672012
R24591 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R24592 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R24593 a_n2903_n3924.n20 a_n2903_n3924.n19 0.643669
R24594 a_n2903_n3924.n15 a_n2903_n3924.n1 0.501227
R24595 a_n2903_n3924.n24 a_n2903_n3924.n22 0.358259
R24596 a_n2903_n3924.n26 a_n2903_n3924.n24 0.358259
R24597 a_n2903_n3924.n28 a_n2903_n3924.n26 0.358259
R24598 a_n2903_n3924.n30 a_n2903_n3924.n28 0.358259
R24599 a_n2903_n3924.n32 a_n2903_n3924.n30 0.358259
R24600 a_n2903_n3924.n33 a_n2903_n3924.n32 0.358259
R24601 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R24602 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R24603 a_n2903_n3924.n40 a_n2903_n3924.n38 0.358259
R24604 a_n2903_n3924.n42 a_n2903_n3924.n40 0.358259
R24605 a_n2903_n3924.n44 a_n2903_n3924.n42 0.358259
R24606 a_n2903_n3924.n45 a_n2903_n3924.n44 0.358259
R24607 a_n2903_n3924.n13 a_n2903_n3924.n12 0.358259
R24608 a_n2903_n3924.n12 a_n2903_n3924.n10 0.358259
R24609 a_n2903_n3924.n10 a_n2903_n3924.n8 0.358259
R24610 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R24611 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R24612 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R24613 a_n2903_n3924.n56 a_n2903_n3924.n0 0.358259
R24614 a_n2903_n3924.n56 a_n2903_n3924.n55 0.358259
R24615 a_n2903_n3924.n55 a_n2903_n3924.n53 0.358259
R24616 a_n2903_n3924.n53 a_n2903_n3924.n51 0.358259
R24617 a_n2903_n3924.n51 a_n2903_n3924.n49 0.358259
R24618 a_n2903_n3924.n49 a_n2903_n3924.n47 0.358259
R24619 a_n2903_n3924.n34 a_n2903_n3924.n33 0.235414
R24620 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R24621 a_n2903_n3924.n20 a_n2903_n3924.n14 0.028843
R24622 minus.n45 minus.t26 442.325
R24623 minus.n9 minus.t12 442.325
R24624 minus.n66 minus.t16 415.966
R24625 minus.n64 minus.t28 415.966
R24626 minus.n63 minus.t21 415.966
R24627 minus.n37 minus.t14 415.966
R24628 minus.n57 minus.t23 415.966
R24629 minus.n56 minus.t11 415.966
R24630 minus.n40 minus.t5 415.966
R24631 minus.n51 minus.t17 415.966
R24632 minus.n49 minus.t10 415.966
R24633 minus.n43 minus.t25 415.966
R24634 minus.n44 minus.t7 415.966
R24635 minus.n8 minus.t18 415.966
R24636 minus.n7 minus.t8 415.966
R24637 minus.n13 minus.t13 415.966
R24638 minus.n5 minus.t24 415.966
R24639 minus.n18 minus.t19 415.966
R24640 minus.n20 minus.t22 415.966
R24641 minus.n3 minus.t6 415.966
R24642 minus.n25 minus.t20 415.966
R24643 minus.n1 minus.t27 415.966
R24644 minus.n30 minus.t15 415.966
R24645 minus.n32 minus.t9 415.966
R24646 minus.n72 minus.t3 243.255
R24647 minus.n71 minus.n69 224.169
R24648 minus.n71 minus.n70 223.454
R24649 minus.n46 minus.n43 161.3
R24650 minus.n48 minus.n47 161.3
R24651 minus.n49 minus.n42 161.3
R24652 minus.n50 minus.n41 161.3
R24653 minus.n52 minus.n51 161.3
R24654 minus.n53 minus.n40 161.3
R24655 minus.n55 minus.n54 161.3
R24656 minus.n56 minus.n39 161.3
R24657 minus.n57 minus.n38 161.3
R24658 minus.n59 minus.n58 161.3
R24659 minus.n60 minus.n37 161.3
R24660 minus.n62 minus.n61 161.3
R24661 minus.n63 minus.n36 161.3
R24662 minus.n64 minus.n35 161.3
R24663 minus.n65 minus.n34 161.3
R24664 minus.n67 minus.n66 161.3
R24665 minus.n33 minus.n32 161.3
R24666 minus.n31 minus.n0 161.3
R24667 minus.n30 minus.n29 161.3
R24668 minus.n28 minus.n1 161.3
R24669 minus.n27 minus.n26 161.3
R24670 minus.n25 minus.n2 161.3
R24671 minus.n24 minus.n23 161.3
R24672 minus.n22 minus.n3 161.3
R24673 minus.n21 minus.n20 161.3
R24674 minus.n19 minus.n4 161.3
R24675 minus.n18 minus.n17 161.3
R24676 minus.n16 minus.n5 161.3
R24677 minus.n15 minus.n14 161.3
R24678 minus.n13 minus.n6 161.3
R24679 minus.n12 minus.n11 161.3
R24680 minus.n10 minus.n7 161.3
R24681 minus.n64 minus.n63 48.2005
R24682 minus.n57 minus.n56 48.2005
R24683 minus.n51 minus.n40 48.2005
R24684 minus.n44 minus.n43 48.2005
R24685 minus.n8 minus.n7 48.2005
R24686 minus.n18 minus.n5 48.2005
R24687 minus.n20 minus.n3 48.2005
R24688 minus.n30 minus.n1 48.2005
R24689 minus.n58 minus.n37 47.4702
R24690 minus.n50 minus.n49 47.4702
R24691 minus.n14 minus.n13 47.4702
R24692 minus.n25 minus.n24 47.4702
R24693 minus.n66 minus.n65 46.0096
R24694 minus.n32 minus.n31 46.0096
R24695 minus.n10 minus.n9 45.0871
R24696 minus.n46 minus.n45 45.0871
R24697 minus.n68 minus.n67 31.2713
R24698 minus.n62 minus.n37 25.5611
R24699 minus.n49 minus.n48 25.5611
R24700 minus.n13 minus.n12 25.5611
R24701 minus.n26 minus.n25 25.5611
R24702 minus.n56 minus.n55 24.1005
R24703 minus.n55 minus.n40 24.1005
R24704 minus.n19 minus.n18 24.1005
R24705 minus.n20 minus.n19 24.1005
R24706 minus.n63 minus.n62 22.6399
R24707 minus.n48 minus.n43 22.6399
R24708 minus.n12 minus.n7 22.6399
R24709 minus.n26 minus.n1 22.6399
R24710 minus.n70 minus.t2 19.8005
R24711 minus.n70 minus.t0 19.8005
R24712 minus.n69 minus.t1 19.8005
R24713 minus.n69 minus.t4 19.8005
R24714 minus.n45 minus.n44 14.1472
R24715 minus.n9 minus.n8 14.1472
R24716 minus.n68 minus.n33 11.9418
R24717 minus minus.n73 11.6534
R24718 minus.n73 minus.n72 4.80222
R24719 minus.n65 minus.n64 2.19141
R24720 minus.n31 minus.n30 2.19141
R24721 minus.n73 minus.n68 0.972091
R24722 minus.n58 minus.n57 0.730803
R24723 minus.n51 minus.n50 0.730803
R24724 minus.n14 minus.n5 0.730803
R24725 minus.n24 minus.n3 0.730803
R24726 minus.n72 minus.n71 0.716017
R24727 minus.n67 minus.n34 0.189894
R24728 minus.n35 minus.n34 0.189894
R24729 minus.n36 minus.n35 0.189894
R24730 minus.n61 minus.n36 0.189894
R24731 minus.n61 minus.n60 0.189894
R24732 minus.n60 minus.n59 0.189894
R24733 minus.n59 minus.n38 0.189894
R24734 minus.n39 minus.n38 0.189894
R24735 minus.n54 minus.n39 0.189894
R24736 minus.n54 minus.n53 0.189894
R24737 minus.n53 minus.n52 0.189894
R24738 minus.n52 minus.n41 0.189894
R24739 minus.n42 minus.n41 0.189894
R24740 minus.n47 minus.n42 0.189894
R24741 minus.n47 minus.n46 0.189894
R24742 minus.n11 minus.n10 0.189894
R24743 minus.n11 minus.n6 0.189894
R24744 minus.n15 minus.n6 0.189894
R24745 minus.n16 minus.n15 0.189894
R24746 minus.n17 minus.n16 0.189894
R24747 minus.n17 minus.n4 0.189894
R24748 minus.n21 minus.n4 0.189894
R24749 minus.n22 minus.n21 0.189894
R24750 minus.n23 minus.n22 0.189894
R24751 minus.n23 minus.n2 0.189894
R24752 minus.n27 minus.n2 0.189894
R24753 minus.n28 minus.n27 0.189894
R24754 minus.n29 minus.n28 0.189894
R24755 minus.n29 minus.n0 0.189894
R24756 minus.n33 minus.n0 0.189894
R24757 diffpairibias.n0 diffpairibias.t18 436.822
R24758 diffpairibias.n21 diffpairibias.t19 435.479
R24759 diffpairibias.n20 diffpairibias.t16 435.479
R24760 diffpairibias.n19 diffpairibias.t17 435.479
R24761 diffpairibias.n18 diffpairibias.t21 435.479
R24762 diffpairibias.n0 diffpairibias.t22 435.479
R24763 diffpairibias.n1 diffpairibias.t20 435.479
R24764 diffpairibias.n2 diffpairibias.t23 435.479
R24765 diffpairibias.n10 diffpairibias.t0 377.536
R24766 diffpairibias.n10 diffpairibias.t8 376.193
R24767 diffpairibias.n11 diffpairibias.t10 376.193
R24768 diffpairibias.n12 diffpairibias.t6 376.193
R24769 diffpairibias.n13 diffpairibias.t2 376.193
R24770 diffpairibias.n14 diffpairibias.t12 376.193
R24771 diffpairibias.n15 diffpairibias.t4 376.193
R24772 diffpairibias.n16 diffpairibias.t14 376.193
R24773 diffpairibias.n3 diffpairibias.t1 113.368
R24774 diffpairibias.n3 diffpairibias.t9 112.698
R24775 diffpairibias.n4 diffpairibias.t11 112.698
R24776 diffpairibias.n5 diffpairibias.t7 112.698
R24777 diffpairibias.n6 diffpairibias.t3 112.698
R24778 diffpairibias.n7 diffpairibias.t13 112.698
R24779 diffpairibias.n8 diffpairibias.t5 112.698
R24780 diffpairibias.n9 diffpairibias.t15 112.698
R24781 diffpairibias.n17 diffpairibias.n16 4.77242
R24782 diffpairibias.n17 diffpairibias.n9 4.30807
R24783 diffpairibias.n18 diffpairibias.n17 4.13945
R24784 diffpairibias.n16 diffpairibias.n15 1.34352
R24785 diffpairibias.n15 diffpairibias.n14 1.34352
R24786 diffpairibias.n14 diffpairibias.n13 1.34352
R24787 diffpairibias.n13 diffpairibias.n12 1.34352
R24788 diffpairibias.n12 diffpairibias.n11 1.34352
R24789 diffpairibias.n11 diffpairibias.n10 1.34352
R24790 diffpairibias.n2 diffpairibias.n1 1.34352
R24791 diffpairibias.n1 diffpairibias.n0 1.34352
R24792 diffpairibias.n19 diffpairibias.n18 1.34352
R24793 diffpairibias.n20 diffpairibias.n19 1.34352
R24794 diffpairibias.n21 diffpairibias.n20 1.34352
R24795 diffpairibias.n22 diffpairibias.n21 0.862419
R24796 diffpairibias diffpairibias.n22 0.684875
R24797 diffpairibias.n9 diffpairibias.n8 0.672012
R24798 diffpairibias.n8 diffpairibias.n7 0.672012
R24799 diffpairibias.n7 diffpairibias.n6 0.672012
R24800 diffpairibias.n6 diffpairibias.n5 0.672012
R24801 diffpairibias.n5 diffpairibias.n4 0.672012
R24802 diffpairibias.n4 diffpairibias.n3 0.672012
R24803 diffpairibias.n22 diffpairibias.n2 0.190907
R24804 outputibias.n27 outputibias.n1 289.615
R24805 outputibias.n58 outputibias.n32 289.615
R24806 outputibias.n90 outputibias.n64 289.615
R24807 outputibias.n122 outputibias.n96 289.615
R24808 outputibias.n28 outputibias.n27 185
R24809 outputibias.n26 outputibias.n25 185
R24810 outputibias.n5 outputibias.n4 185
R24811 outputibias.n20 outputibias.n19 185
R24812 outputibias.n18 outputibias.n17 185
R24813 outputibias.n9 outputibias.n8 185
R24814 outputibias.n12 outputibias.n11 185
R24815 outputibias.n59 outputibias.n58 185
R24816 outputibias.n57 outputibias.n56 185
R24817 outputibias.n36 outputibias.n35 185
R24818 outputibias.n51 outputibias.n50 185
R24819 outputibias.n49 outputibias.n48 185
R24820 outputibias.n40 outputibias.n39 185
R24821 outputibias.n43 outputibias.n42 185
R24822 outputibias.n91 outputibias.n90 185
R24823 outputibias.n89 outputibias.n88 185
R24824 outputibias.n68 outputibias.n67 185
R24825 outputibias.n83 outputibias.n82 185
R24826 outputibias.n81 outputibias.n80 185
R24827 outputibias.n72 outputibias.n71 185
R24828 outputibias.n75 outputibias.n74 185
R24829 outputibias.n123 outputibias.n122 185
R24830 outputibias.n121 outputibias.n120 185
R24831 outputibias.n100 outputibias.n99 185
R24832 outputibias.n115 outputibias.n114 185
R24833 outputibias.n113 outputibias.n112 185
R24834 outputibias.n104 outputibias.n103 185
R24835 outputibias.n107 outputibias.n106 185
R24836 outputibias.n0 outputibias.t10 178.945
R24837 outputibias.n133 outputibias.t8 177.018
R24838 outputibias.n132 outputibias.t11 177.018
R24839 outputibias.n0 outputibias.t9 177.018
R24840 outputibias.t7 outputibias.n10 147.661
R24841 outputibias.t3 outputibias.n41 147.661
R24842 outputibias.t1 outputibias.n73 147.661
R24843 outputibias.t5 outputibias.n105 147.661
R24844 outputibias.n128 outputibias.t6 132.363
R24845 outputibias.n128 outputibias.t2 130.436
R24846 outputibias.n129 outputibias.t0 130.436
R24847 outputibias.n130 outputibias.t4 130.436
R24848 outputibias.n27 outputibias.n26 104.615
R24849 outputibias.n26 outputibias.n4 104.615
R24850 outputibias.n19 outputibias.n4 104.615
R24851 outputibias.n19 outputibias.n18 104.615
R24852 outputibias.n18 outputibias.n8 104.615
R24853 outputibias.n11 outputibias.n8 104.615
R24854 outputibias.n58 outputibias.n57 104.615
R24855 outputibias.n57 outputibias.n35 104.615
R24856 outputibias.n50 outputibias.n35 104.615
R24857 outputibias.n50 outputibias.n49 104.615
R24858 outputibias.n49 outputibias.n39 104.615
R24859 outputibias.n42 outputibias.n39 104.615
R24860 outputibias.n90 outputibias.n89 104.615
R24861 outputibias.n89 outputibias.n67 104.615
R24862 outputibias.n82 outputibias.n67 104.615
R24863 outputibias.n82 outputibias.n81 104.615
R24864 outputibias.n81 outputibias.n71 104.615
R24865 outputibias.n74 outputibias.n71 104.615
R24866 outputibias.n122 outputibias.n121 104.615
R24867 outputibias.n121 outputibias.n99 104.615
R24868 outputibias.n114 outputibias.n99 104.615
R24869 outputibias.n114 outputibias.n113 104.615
R24870 outputibias.n113 outputibias.n103 104.615
R24871 outputibias.n106 outputibias.n103 104.615
R24872 outputibias.n63 outputibias.n31 95.6354
R24873 outputibias.n63 outputibias.n62 94.6732
R24874 outputibias.n95 outputibias.n94 94.6732
R24875 outputibias.n127 outputibias.n126 94.6732
R24876 outputibias.n11 outputibias.t7 52.3082
R24877 outputibias.n42 outputibias.t3 52.3082
R24878 outputibias.n74 outputibias.t1 52.3082
R24879 outputibias.n106 outputibias.t5 52.3082
R24880 outputibias.n12 outputibias.n10 15.6674
R24881 outputibias.n43 outputibias.n41 15.6674
R24882 outputibias.n75 outputibias.n73 15.6674
R24883 outputibias.n107 outputibias.n105 15.6674
R24884 outputibias.n13 outputibias.n9 12.8005
R24885 outputibias.n44 outputibias.n40 12.8005
R24886 outputibias.n76 outputibias.n72 12.8005
R24887 outputibias.n108 outputibias.n104 12.8005
R24888 outputibias.n17 outputibias.n16 12.0247
R24889 outputibias.n48 outputibias.n47 12.0247
R24890 outputibias.n80 outputibias.n79 12.0247
R24891 outputibias.n112 outputibias.n111 12.0247
R24892 outputibias.n20 outputibias.n7 11.249
R24893 outputibias.n51 outputibias.n38 11.249
R24894 outputibias.n83 outputibias.n70 11.249
R24895 outputibias.n115 outputibias.n102 11.249
R24896 outputibias.n21 outputibias.n5 10.4732
R24897 outputibias.n52 outputibias.n36 10.4732
R24898 outputibias.n84 outputibias.n68 10.4732
R24899 outputibias.n116 outputibias.n100 10.4732
R24900 outputibias.n25 outputibias.n24 9.69747
R24901 outputibias.n56 outputibias.n55 9.69747
R24902 outputibias.n88 outputibias.n87 9.69747
R24903 outputibias.n120 outputibias.n119 9.69747
R24904 outputibias.n31 outputibias.n30 9.45567
R24905 outputibias.n62 outputibias.n61 9.45567
R24906 outputibias.n94 outputibias.n93 9.45567
R24907 outputibias.n126 outputibias.n125 9.45567
R24908 outputibias.n30 outputibias.n29 9.3005
R24909 outputibias.n3 outputibias.n2 9.3005
R24910 outputibias.n24 outputibias.n23 9.3005
R24911 outputibias.n22 outputibias.n21 9.3005
R24912 outputibias.n7 outputibias.n6 9.3005
R24913 outputibias.n16 outputibias.n15 9.3005
R24914 outputibias.n14 outputibias.n13 9.3005
R24915 outputibias.n61 outputibias.n60 9.3005
R24916 outputibias.n34 outputibias.n33 9.3005
R24917 outputibias.n55 outputibias.n54 9.3005
R24918 outputibias.n53 outputibias.n52 9.3005
R24919 outputibias.n38 outputibias.n37 9.3005
R24920 outputibias.n47 outputibias.n46 9.3005
R24921 outputibias.n45 outputibias.n44 9.3005
R24922 outputibias.n93 outputibias.n92 9.3005
R24923 outputibias.n66 outputibias.n65 9.3005
R24924 outputibias.n87 outputibias.n86 9.3005
R24925 outputibias.n85 outputibias.n84 9.3005
R24926 outputibias.n70 outputibias.n69 9.3005
R24927 outputibias.n79 outputibias.n78 9.3005
R24928 outputibias.n77 outputibias.n76 9.3005
R24929 outputibias.n125 outputibias.n124 9.3005
R24930 outputibias.n98 outputibias.n97 9.3005
R24931 outputibias.n119 outputibias.n118 9.3005
R24932 outputibias.n117 outputibias.n116 9.3005
R24933 outputibias.n102 outputibias.n101 9.3005
R24934 outputibias.n111 outputibias.n110 9.3005
R24935 outputibias.n109 outputibias.n108 9.3005
R24936 outputibias.n28 outputibias.n3 8.92171
R24937 outputibias.n59 outputibias.n34 8.92171
R24938 outputibias.n91 outputibias.n66 8.92171
R24939 outputibias.n123 outputibias.n98 8.92171
R24940 outputibias.n29 outputibias.n1 8.14595
R24941 outputibias.n60 outputibias.n32 8.14595
R24942 outputibias.n92 outputibias.n64 8.14595
R24943 outputibias.n124 outputibias.n96 8.14595
R24944 outputibias.n31 outputibias.n1 5.81868
R24945 outputibias.n62 outputibias.n32 5.81868
R24946 outputibias.n94 outputibias.n64 5.81868
R24947 outputibias.n126 outputibias.n96 5.81868
R24948 outputibias.n131 outputibias.n130 5.20947
R24949 outputibias.n29 outputibias.n28 5.04292
R24950 outputibias.n60 outputibias.n59 5.04292
R24951 outputibias.n92 outputibias.n91 5.04292
R24952 outputibias.n124 outputibias.n123 5.04292
R24953 outputibias.n131 outputibias.n127 4.42209
R24954 outputibias.n14 outputibias.n10 4.38594
R24955 outputibias.n45 outputibias.n41 4.38594
R24956 outputibias.n77 outputibias.n73 4.38594
R24957 outputibias.n109 outputibias.n105 4.38594
R24958 outputibias.n132 outputibias.n131 4.28454
R24959 outputibias.n25 outputibias.n3 4.26717
R24960 outputibias.n56 outputibias.n34 4.26717
R24961 outputibias.n88 outputibias.n66 4.26717
R24962 outputibias.n120 outputibias.n98 4.26717
R24963 outputibias.n24 outputibias.n5 3.49141
R24964 outputibias.n55 outputibias.n36 3.49141
R24965 outputibias.n87 outputibias.n68 3.49141
R24966 outputibias.n119 outputibias.n100 3.49141
R24967 outputibias.n21 outputibias.n20 2.71565
R24968 outputibias.n52 outputibias.n51 2.71565
R24969 outputibias.n84 outputibias.n83 2.71565
R24970 outputibias.n116 outputibias.n115 2.71565
R24971 outputibias.n17 outputibias.n7 1.93989
R24972 outputibias.n48 outputibias.n38 1.93989
R24973 outputibias.n80 outputibias.n70 1.93989
R24974 outputibias.n112 outputibias.n102 1.93989
R24975 outputibias.n130 outputibias.n129 1.9266
R24976 outputibias.n129 outputibias.n128 1.9266
R24977 outputibias.n133 outputibias.n132 1.92658
R24978 outputibias.n134 outputibias.n133 1.29913
R24979 outputibias.n16 outputibias.n9 1.16414
R24980 outputibias.n47 outputibias.n40 1.16414
R24981 outputibias.n79 outputibias.n72 1.16414
R24982 outputibias.n111 outputibias.n104 1.16414
R24983 outputibias.n127 outputibias.n95 0.962709
R24984 outputibias.n95 outputibias.n63 0.962709
R24985 outputibias.n13 outputibias.n12 0.388379
R24986 outputibias.n44 outputibias.n43 0.388379
R24987 outputibias.n76 outputibias.n75 0.388379
R24988 outputibias.n108 outputibias.n107 0.388379
R24989 outputibias.n134 outputibias.n0 0.337251
R24990 outputibias outputibias.n134 0.302375
R24991 outputibias.n30 outputibias.n2 0.155672
R24992 outputibias.n23 outputibias.n2 0.155672
R24993 outputibias.n23 outputibias.n22 0.155672
R24994 outputibias.n22 outputibias.n6 0.155672
R24995 outputibias.n15 outputibias.n6 0.155672
R24996 outputibias.n15 outputibias.n14 0.155672
R24997 outputibias.n61 outputibias.n33 0.155672
R24998 outputibias.n54 outputibias.n33 0.155672
R24999 outputibias.n54 outputibias.n53 0.155672
R25000 outputibias.n53 outputibias.n37 0.155672
R25001 outputibias.n46 outputibias.n37 0.155672
R25002 outputibias.n46 outputibias.n45 0.155672
R25003 outputibias.n93 outputibias.n65 0.155672
R25004 outputibias.n86 outputibias.n65 0.155672
R25005 outputibias.n86 outputibias.n85 0.155672
R25006 outputibias.n85 outputibias.n69 0.155672
R25007 outputibias.n78 outputibias.n69 0.155672
R25008 outputibias.n78 outputibias.n77 0.155672
R25009 outputibias.n125 outputibias.n97 0.155672
R25010 outputibias.n118 outputibias.n97 0.155672
R25011 outputibias.n118 outputibias.n117 0.155672
R25012 outputibias.n117 outputibias.n101 0.155672
R25013 outputibias.n110 outputibias.n101 0.155672
R25014 outputibias.n110 outputibias.n109 0.155672
C0 minus diffpairibias 2.98e-19
C1 commonsourceibias output 0.006829f
C2 CSoutput minus 2.85492f
C3 vdd plus 0.100442f
C4 commonsourceibias outputibias 0.003902f
C5 plus diffpairibias 2.75e-19
C6 vdd commonsourceibias 0.004262f
C7 CSoutput plus 0.859513f
C8 commonsourceibias diffpairibias 0.06482f
C9 CSoutput commonsourceibias 54.115f
C10 minus plus 9.23087f
C11 minus commonsourceibias 0.322616f
C12 plus commonsourceibias 0.276969f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13881f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 0.14236p
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.183644p
C22 plus gnd 33.4315f
C23 minus gnd 27.91584f
C24 CSoutput gnd 0.124285p
C25 vdd gnd 0.542244p
C26 outputibias.t9 gnd 0.11477f
C27 outputibias.t10 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t7 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t3 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t1 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t5 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t4 gnd 0.108319f
C161 outputibias.t0 gnd 0.108319f
C162 outputibias.t2 gnd 0.108319f
C163 outputibias.t6 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t11 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t8 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 minus.n0 gnd 0.032753f
C221 minus.t27 gnd 0.330896f
C222 minus.n1 gnd 0.152681f
C223 minus.n2 gnd 0.032753f
C224 minus.t6 gnd 0.330896f
C225 minus.n3 gnd 0.149652f
C226 minus.n4 gnd 0.032753f
C227 minus.t24 gnd 0.330896f
C228 minus.n5 gnd 0.149652f
C229 minus.n6 gnd 0.032753f
C230 minus.t8 gnd 0.330896f
C231 minus.n7 gnd 0.152681f
C232 minus.t12 gnd 0.339805f
C233 minus.t18 gnd 0.330896f
C234 minus.n8 gnd 0.156556f
C235 minus.n9 gnd 0.141715f
C236 minus.n10 gnd 0.132989f
C237 minus.n11 gnd 0.032753f
C238 minus.n12 gnd 0.007432f
C239 minus.t13 gnd 0.330896f
C240 minus.n13 gnd 0.152984f
C241 minus.n14 gnd 0.007432f
C242 minus.n15 gnd 0.032753f
C243 minus.n16 gnd 0.032753f
C244 minus.n17 gnd 0.032753f
C245 minus.t19 gnd 0.330896f
C246 minus.n18 gnd 0.152883f
C247 minus.n19 gnd 0.007432f
C248 minus.t22 gnd 0.330896f
C249 minus.n20 gnd 0.152883f
C250 minus.n21 gnd 0.032753f
C251 minus.n22 gnd 0.032753f
C252 minus.n23 gnd 0.032753f
C253 minus.n24 gnd 0.007432f
C254 minus.t20 gnd 0.330896f
C255 minus.n25 gnd 0.152984f
C256 minus.n26 gnd 0.007432f
C257 minus.n27 gnd 0.032753f
C258 minus.n28 gnd 0.032753f
C259 minus.n29 gnd 0.032753f
C260 minus.t15 gnd 0.330896f
C261 minus.n30 gnd 0.149854f
C262 minus.n31 gnd 0.007432f
C263 minus.t9 gnd 0.330896f
C264 minus.n32 gnd 0.149248f
C265 minus.n33 gnd 0.367575f
C266 minus.n34 gnd 0.032753f
C267 minus.t16 gnd 0.330896f
C268 minus.t28 gnd 0.330896f
C269 minus.n35 gnd 0.032753f
C270 minus.t21 gnd 0.330896f
C271 minus.n36 gnd 0.032753f
C272 minus.t14 gnd 0.330896f
C273 minus.n37 gnd 0.152984f
C274 minus.n38 gnd 0.032753f
C275 minus.t23 gnd 0.330896f
C276 minus.t11 gnd 0.330896f
C277 minus.n39 gnd 0.032753f
C278 minus.t5 gnd 0.330896f
C279 minus.n40 gnd 0.152883f
C280 minus.n41 gnd 0.032753f
C281 minus.t17 gnd 0.330896f
C282 minus.t10 gnd 0.330896f
C283 minus.n42 gnd 0.032753f
C284 minus.t25 gnd 0.330896f
C285 minus.n43 gnd 0.152681f
C286 minus.t26 gnd 0.339805f
C287 minus.t7 gnd 0.330896f
C288 minus.n44 gnd 0.156556f
C289 minus.n45 gnd 0.141715f
C290 minus.n46 gnd 0.132989f
C291 minus.n47 gnd 0.032753f
C292 minus.n48 gnd 0.007432f
C293 minus.n49 gnd 0.152984f
C294 minus.n50 gnd 0.007432f
C295 minus.n51 gnd 0.149652f
C296 minus.n52 gnd 0.032753f
C297 minus.n53 gnd 0.032753f
C298 minus.n54 gnd 0.032753f
C299 minus.n55 gnd 0.007432f
C300 minus.n56 gnd 0.152883f
C301 minus.n57 gnd 0.149652f
C302 minus.n58 gnd 0.007432f
C303 minus.n59 gnd 0.032753f
C304 minus.n60 gnd 0.032753f
C305 minus.n61 gnd 0.032753f
C306 minus.n62 gnd 0.007432f
C307 minus.n63 gnd 0.152681f
C308 minus.n64 gnd 0.149854f
C309 minus.n65 gnd 0.007432f
C310 minus.n66 gnd 0.149248f
C311 minus.n67 gnd 0.993889f
C312 minus.n68 gnd 1.50764f
C313 minus.t1 gnd 0.010097f
C314 minus.t4 gnd 0.010097f
C315 minus.n69 gnd 0.0332f
C316 minus.t2 gnd 0.010097f
C317 minus.t0 gnd 0.010097f
C318 minus.n70 gnd 0.032745f
C319 minus.n71 gnd 0.279466f
C320 minus.t3 gnd 0.056197f
C321 minus.n72 gnd 0.152502f
C322 minus.n73 gnd 2.13826f
C323 a_n2903_n3924.t18 gnd 0.108618f
C324 a_n2903_n3924.t13 gnd 1.12888f
C325 a_n2903_n3924.n0 gnd 0.383133f
C326 a_n2903_n3924.t51 gnd 1.40337f
C327 a_n2903_n3924.n1 gnd 1.48426f
C328 a_n2903_n3924.t37 gnd 1.12888f
C329 a_n2903_n3924.n2 gnd 0.383133f
C330 a_n2903_n3924.t39 gnd 0.108618f
C331 a_n2903_n3924.t49 gnd 0.108618f
C332 a_n2903_n3924.n3 gnd 0.887099f
C333 a_n2903_n3924.n4 gnd 0.359777f
C334 a_n2903_n3924.t52 gnd 0.108618f
C335 a_n2903_n3924.t48 gnd 0.108618f
C336 a_n2903_n3924.n5 gnd 0.887099f
C337 a_n2903_n3924.n6 gnd 0.359777f
C338 a_n2903_n3924.t40 gnd 0.108618f
C339 a_n2903_n3924.t2 gnd 0.108618f
C340 a_n2903_n3924.n7 gnd 0.887099f
C341 a_n2903_n3924.n8 gnd 0.359777f
C342 a_n2903_n3924.t34 gnd 0.108618f
C343 a_n2903_n3924.t46 gnd 0.108618f
C344 a_n2903_n3924.n9 gnd 0.887099f
C345 a_n2903_n3924.n10 gnd 0.359777f
C346 a_n2903_n3924.t54 gnd 0.108618f
C347 a_n2903_n3924.t4 gnd 0.108618f
C348 a_n2903_n3924.n11 gnd 0.887099f
C349 a_n2903_n3924.n12 gnd 0.359777f
C350 a_n2903_n3924.t38 gnd 1.12888f
C351 a_n2903_n3924.n13 gnd 0.974186f
C352 a_n2903_n3924.t3 gnd 1.40461f
C353 a_n2903_n3924.t0 gnd 1.40261f
C354 a_n2903_n3924.n14 gnd 1.26893f
C355 a_n2903_n3924.t7 gnd 1.40261f
C356 a_n2903_n3924.n15 gnd 0.892855f
C357 a_n2903_n3924.t36 gnd 1.40261f
C358 a_n2903_n3924.n16 gnd 0.987884f
C359 a_n2903_n3924.t5 gnd 1.40261f
C360 a_n2903_n3924.n17 gnd 0.987884f
C361 a_n2903_n3924.t43 gnd 1.40261f
C362 a_n2903_n3924.n18 gnd 0.987884f
C363 a_n2903_n3924.t50 gnd 1.40261f
C364 a_n2903_n3924.n19 gnd 0.972113f
C365 a_n2903_n3924.n20 gnd 0.533935f
C366 a_n2903_n3924.n21 gnd 1.01395f
C367 a_n2903_n3924.t15 gnd 1.12888f
C368 a_n2903_n3924.n22 gnd 0.619233f
C369 a_n2903_n3924.t25 gnd 0.108618f
C370 a_n2903_n3924.t11 gnd 0.108618f
C371 a_n2903_n3924.n23 gnd 0.887098f
C372 a_n2903_n3924.n24 gnd 0.359779f
C373 a_n2903_n3924.t16 gnd 0.108618f
C374 a_n2903_n3924.t31 gnd 0.108618f
C375 a_n2903_n3924.n25 gnd 0.887098f
C376 a_n2903_n3924.n26 gnd 0.359779f
C377 a_n2903_n3924.t20 gnd 0.108618f
C378 a_n2903_n3924.t24 gnd 0.108618f
C379 a_n2903_n3924.n27 gnd 0.887098f
C380 a_n2903_n3924.n28 gnd 0.359779f
C381 a_n2903_n3924.t14 gnd 0.108618f
C382 a_n2903_n3924.t21 gnd 0.108618f
C383 a_n2903_n3924.n29 gnd 0.887098f
C384 a_n2903_n3924.n30 gnd 0.359779f
C385 a_n2903_n3924.t29 gnd 0.108618f
C386 a_n2903_n3924.t23 gnd 0.108618f
C387 a_n2903_n3924.n31 gnd 0.887098f
C388 a_n2903_n3924.n32 gnd 0.359779f
C389 a_n2903_n3924.t26 gnd 1.12888f
C390 a_n2903_n3924.n33 gnd 0.383138f
C391 a_n2903_n3924.t53 gnd 1.12888f
C392 a_n2903_n3924.n34 gnd 0.383138f
C393 a_n2903_n3924.t45 gnd 0.108618f
C394 a_n2903_n3924.t9 gnd 0.108618f
C395 a_n2903_n3924.n35 gnd 0.887098f
C396 a_n2903_n3924.n36 gnd 0.359779f
C397 a_n2903_n3924.t8 gnd 0.108618f
C398 a_n2903_n3924.t41 gnd 0.108618f
C399 a_n2903_n3924.n37 gnd 0.887098f
C400 a_n2903_n3924.n38 gnd 0.359779f
C401 a_n2903_n3924.t6 gnd 0.108618f
C402 a_n2903_n3924.t47 gnd 0.108618f
C403 a_n2903_n3924.n39 gnd 0.887098f
C404 a_n2903_n3924.n40 gnd 0.359779f
C405 a_n2903_n3924.t42 gnd 0.108618f
C406 a_n2903_n3924.t55 gnd 0.108618f
C407 a_n2903_n3924.n41 gnd 0.887098f
C408 a_n2903_n3924.n42 gnd 0.359779f
C409 a_n2903_n3924.t44 gnd 0.108618f
C410 a_n2903_n3924.t35 gnd 0.108618f
C411 a_n2903_n3924.n43 gnd 0.887098f
C412 a_n2903_n3924.n44 gnd 0.359779f
C413 a_n2903_n3924.t1 gnd 1.12888f
C414 a_n2903_n3924.n45 gnd 0.619233f
C415 a_n2903_n3924.n46 gnd 1.01395f
C416 a_n2903_n3924.t17 gnd 1.12888f
C417 a_n2903_n3924.n47 gnd 0.97419f
C418 a_n2903_n3924.t22 gnd 0.108618f
C419 a_n2903_n3924.t10 gnd 0.108618f
C420 a_n2903_n3924.n48 gnd 0.887099f
C421 a_n2903_n3924.n49 gnd 0.359777f
C422 a_n2903_n3924.t19 gnd 0.108618f
C423 a_n2903_n3924.t30 gnd 0.108618f
C424 a_n2903_n3924.n50 gnd 0.887099f
C425 a_n2903_n3924.n51 gnd 0.359777f
C426 a_n2903_n3924.t32 gnd 0.108618f
C427 a_n2903_n3924.t28 gnd 0.108618f
C428 a_n2903_n3924.n52 gnd 0.887099f
C429 a_n2903_n3924.n53 gnd 0.359777f
C430 a_n2903_n3924.t12 gnd 0.108618f
C431 a_n2903_n3924.t27 gnd 0.108618f
C432 a_n2903_n3924.n54 gnd 0.887099f
C433 a_n2903_n3924.n55 gnd 0.359777f
C434 a_n2903_n3924.n56 gnd 0.359776f
C435 a_n2903_n3924.n57 gnd 0.887101f
C436 a_n2903_n3924.t33 gnd 0.108618f
C437 plus.n0 gnd 0.023738f
C438 plus.t23 gnd 0.239826f
C439 plus.n1 gnd 0.023738f
C440 plus.t13 gnd 0.239826f
C441 plus.n2 gnd 0.023738f
C442 plus.t27 gnd 0.239826f
C443 plus.t22 gnd 0.239826f
C444 plus.n3 gnd 0.110879f
C445 plus.n4 gnd 0.023738f
C446 plus.t7 gnd 0.239826f
C447 plus.n5 gnd 0.023738f
C448 plus.t18 gnd 0.239826f
C449 plus.t14 gnd 0.239826f
C450 plus.n6 gnd 0.110806f
C451 plus.n7 gnd 0.023738f
C452 plus.t24 gnd 0.239826f
C453 plus.n8 gnd 0.023738f
C454 plus.t17 gnd 0.239826f
C455 plus.t9 gnd 0.239826f
C456 plus.n9 gnd 0.11066f
C457 plus.t12 gnd 0.246283f
C458 plus.t15 gnd 0.239826f
C459 plus.n10 gnd 0.113468f
C460 plus.n11 gnd 0.102712f
C461 plus.n12 gnd 0.096387f
C462 plus.n13 gnd 0.023738f
C463 plus.n14 gnd 0.005387f
C464 plus.n15 gnd 0.110879f
C465 plus.n16 gnd 0.005387f
C466 plus.n17 gnd 0.108464f
C467 plus.n18 gnd 0.023738f
C468 plus.n19 gnd 0.023738f
C469 plus.n20 gnd 0.023738f
C470 plus.n21 gnd 0.005387f
C471 plus.n22 gnd 0.110806f
C472 plus.n23 gnd 0.108464f
C473 plus.n24 gnd 0.005387f
C474 plus.n25 gnd 0.023738f
C475 plus.n26 gnd 0.023738f
C476 plus.n27 gnd 0.023738f
C477 plus.n28 gnd 0.005387f
C478 plus.n29 gnd 0.11066f
C479 plus.n30 gnd 0.108611f
C480 plus.n31 gnd 0.005387f
C481 plus.n32 gnd 0.108172f
C482 plus.n33 gnd 0.260277f
C483 plus.n34 gnd 0.023738f
C484 plus.t16 gnd 0.239826f
C485 plus.n35 gnd 0.11066f
C486 plus.t28 gnd 0.239826f
C487 plus.n36 gnd 0.023738f
C488 plus.t19 gnd 0.239826f
C489 plus.n37 gnd 0.108464f
C490 plus.n38 gnd 0.023738f
C491 plus.t11 gnd 0.239826f
C492 plus.n39 gnd 0.108464f
C493 plus.t6 gnd 0.239826f
C494 plus.n40 gnd 0.023738f
C495 plus.t20 gnd 0.239826f
C496 plus.n41 gnd 0.11066f
C497 plus.t25 gnd 0.246283f
C498 plus.t5 gnd 0.239826f
C499 plus.n42 gnd 0.113468f
C500 plus.n43 gnd 0.102712f
C501 plus.n44 gnd 0.096387f
C502 plus.n45 gnd 0.023738f
C503 plus.n46 gnd 0.005387f
C504 plus.t26 gnd 0.239826f
C505 plus.n47 gnd 0.110879f
C506 plus.n48 gnd 0.005387f
C507 plus.n49 gnd 0.023738f
C508 plus.n50 gnd 0.023738f
C509 plus.n51 gnd 0.023738f
C510 plus.n52 gnd 0.110806f
C511 plus.n53 gnd 0.005387f
C512 plus.t10 gnd 0.239826f
C513 plus.n54 gnd 0.110806f
C514 plus.n55 gnd 0.023738f
C515 plus.n56 gnd 0.023738f
C516 plus.n57 gnd 0.023738f
C517 plus.n58 gnd 0.005387f
C518 plus.t8 gnd 0.239826f
C519 plus.n59 gnd 0.110879f
C520 plus.n60 gnd 0.005387f
C521 plus.n61 gnd 0.023738f
C522 plus.n62 gnd 0.023738f
C523 plus.n63 gnd 0.023738f
C524 plus.n64 gnd 0.108611f
C525 plus.n65 gnd 0.005387f
C526 plus.t21 gnd 0.239826f
C527 plus.n66 gnd 0.108172f
C528 plus.n67 gnd 0.710803f
C529 plus.n68 gnd 1.08335f
C530 plus.t3 gnd 0.040979f
C531 plus.t4 gnd 0.007318f
C532 plus.t1 gnd 0.007318f
C533 plus.n69 gnd 0.023733f
C534 plus.n70 gnd 0.184241f
C535 plus.t0 gnd 0.007318f
C536 plus.t2 gnd 0.007318f
C537 plus.n71 gnd 0.023733f
C538 plus.n72 gnd 0.138296f
C539 plus.n73 gnd 2.71566f
C540 output.t13 gnd 0.464308f
C541 output.t9 gnd 0.044422f
C542 output.t7 gnd 0.044422f
C543 output.n0 gnd 0.364624f
C544 output.n1 gnd 0.614102f
C545 output.t1 gnd 0.044422f
C546 output.t3 gnd 0.044422f
C547 output.n2 gnd 0.364624f
C548 output.n3 gnd 0.350265f
C549 output.t4 gnd 0.044422f
C550 output.t11 gnd 0.044422f
C551 output.n4 gnd 0.364624f
C552 output.n5 gnd 0.350265f
C553 output.t14 gnd 0.044422f
C554 output.t2 gnd 0.044422f
C555 output.n6 gnd 0.364624f
C556 output.n7 gnd 0.350265f
C557 output.t5 gnd 0.044422f
C558 output.t10 gnd 0.044422f
C559 output.n8 gnd 0.364624f
C560 output.n9 gnd 0.350265f
C561 output.t12 gnd 0.044422f
C562 output.t0 gnd 0.044422f
C563 output.n10 gnd 0.364624f
C564 output.n11 gnd 0.350265f
C565 output.t8 gnd 0.044422f
C566 output.t6 gnd 0.044422f
C567 output.n12 gnd 0.364624f
C568 output.n13 gnd 0.350265f
C569 output.t15 gnd 0.462979f
C570 output.n14 gnd 0.28994f
C571 output.n15 gnd 0.015803f
C572 output.n16 gnd 0.011243f
C573 output.n17 gnd 0.006041f
C574 output.n18 gnd 0.01428f
C575 output.n19 gnd 0.006397f
C576 output.n20 gnd 0.011243f
C577 output.n21 gnd 0.006041f
C578 output.n22 gnd 0.01428f
C579 output.n23 gnd 0.006397f
C580 output.n24 gnd 0.048111f
C581 output.t19 gnd 0.023274f
C582 output.n25 gnd 0.01071f
C583 output.n26 gnd 0.008435f
C584 output.n27 gnd 0.006041f
C585 output.n28 gnd 0.267512f
C586 output.n29 gnd 0.011243f
C587 output.n30 gnd 0.006041f
C588 output.n31 gnd 0.006397f
C589 output.n32 gnd 0.01428f
C590 output.n33 gnd 0.01428f
C591 output.n34 gnd 0.006397f
C592 output.n35 gnd 0.006041f
C593 output.n36 gnd 0.011243f
C594 output.n37 gnd 0.011243f
C595 output.n38 gnd 0.006041f
C596 output.n39 gnd 0.006397f
C597 output.n40 gnd 0.01428f
C598 output.n41 gnd 0.030913f
C599 output.n42 gnd 0.006397f
C600 output.n43 gnd 0.006041f
C601 output.n44 gnd 0.025987f
C602 output.n45 gnd 0.097665f
C603 output.n46 gnd 0.015803f
C604 output.n47 gnd 0.011243f
C605 output.n48 gnd 0.006041f
C606 output.n49 gnd 0.01428f
C607 output.n50 gnd 0.006397f
C608 output.n51 gnd 0.011243f
C609 output.n52 gnd 0.006041f
C610 output.n53 gnd 0.01428f
C611 output.n54 gnd 0.006397f
C612 output.n55 gnd 0.048111f
C613 output.t18 gnd 0.023274f
C614 output.n56 gnd 0.01071f
C615 output.n57 gnd 0.008435f
C616 output.n58 gnd 0.006041f
C617 output.n59 gnd 0.267512f
C618 output.n60 gnd 0.011243f
C619 output.n61 gnd 0.006041f
C620 output.n62 gnd 0.006397f
C621 output.n63 gnd 0.01428f
C622 output.n64 gnd 0.01428f
C623 output.n65 gnd 0.006397f
C624 output.n66 gnd 0.006041f
C625 output.n67 gnd 0.011243f
C626 output.n68 gnd 0.011243f
C627 output.n69 gnd 0.006041f
C628 output.n70 gnd 0.006397f
C629 output.n71 gnd 0.01428f
C630 output.n72 gnd 0.030913f
C631 output.n73 gnd 0.006397f
C632 output.n74 gnd 0.006041f
C633 output.n75 gnd 0.025987f
C634 output.n76 gnd 0.09306f
C635 output.n77 gnd 1.65264f
C636 output.n78 gnd 0.015803f
C637 output.n79 gnd 0.011243f
C638 output.n80 gnd 0.006041f
C639 output.n81 gnd 0.01428f
C640 output.n82 gnd 0.006397f
C641 output.n83 gnd 0.011243f
C642 output.n84 gnd 0.006041f
C643 output.n85 gnd 0.01428f
C644 output.n86 gnd 0.006397f
C645 output.n87 gnd 0.048111f
C646 output.t16 gnd 0.023274f
C647 output.n88 gnd 0.01071f
C648 output.n89 gnd 0.008435f
C649 output.n90 gnd 0.006041f
C650 output.n91 gnd 0.267512f
C651 output.n92 gnd 0.011243f
C652 output.n93 gnd 0.006041f
C653 output.n94 gnd 0.006397f
C654 output.n95 gnd 0.01428f
C655 output.n96 gnd 0.01428f
C656 output.n97 gnd 0.006397f
C657 output.n98 gnd 0.006041f
C658 output.n99 gnd 0.011243f
C659 output.n100 gnd 0.011243f
C660 output.n101 gnd 0.006041f
C661 output.n102 gnd 0.006397f
C662 output.n103 gnd 0.01428f
C663 output.n104 gnd 0.030913f
C664 output.n105 gnd 0.006397f
C665 output.n106 gnd 0.006041f
C666 output.n107 gnd 0.025987f
C667 output.n108 gnd 0.09306f
C668 output.n109 gnd 0.713089f
C669 output.n110 gnd 0.015803f
C670 output.n111 gnd 0.011243f
C671 output.n112 gnd 0.006041f
C672 output.n113 gnd 0.01428f
C673 output.n114 gnd 0.006397f
C674 output.n115 gnd 0.011243f
C675 output.n116 gnd 0.006041f
C676 output.n117 gnd 0.01428f
C677 output.n118 gnd 0.006397f
C678 output.n119 gnd 0.048111f
C679 output.t17 gnd 0.023274f
C680 output.n120 gnd 0.01071f
C681 output.n121 gnd 0.008435f
C682 output.n122 gnd 0.006041f
C683 output.n123 gnd 0.267512f
C684 output.n124 gnd 0.011243f
C685 output.n125 gnd 0.006041f
C686 output.n126 gnd 0.006397f
C687 output.n127 gnd 0.01428f
C688 output.n128 gnd 0.01428f
C689 output.n129 gnd 0.006397f
C690 output.n130 gnd 0.006041f
C691 output.n131 gnd 0.011243f
C692 output.n132 gnd 0.011243f
C693 output.n133 gnd 0.006041f
C694 output.n134 gnd 0.006397f
C695 output.n135 gnd 0.01428f
C696 output.n136 gnd 0.030913f
C697 output.n137 gnd 0.006397f
C698 output.n138 gnd 0.006041f
C699 output.n139 gnd 0.025987f
C700 output.n140 gnd 0.09306f
C701 output.n141 gnd 1.67353f
C702 a_n2982_8322.t13 gnd 0.100161f
C703 a_n2982_8322.t2 gnd 20.7793f
C704 a_n2982_8322.t1 gnd 20.633598f
C705 a_n2982_8322.t5 gnd 20.633598f
C706 a_n2982_8322.t4 gnd 20.7793f
C707 a_n2982_8322.t3 gnd 20.633598f
C708 a_n2982_8322.t0 gnd 28.9697f
C709 a_n2982_8322.t12 gnd 0.937857f
C710 a_n2982_8322.t25 gnd 0.100161f
C711 a_n2982_8322.t21 gnd 0.100161f
C712 a_n2982_8322.n0 gnd 0.705534f
C713 a_n2982_8322.n1 gnd 0.78833f
C714 a_n2982_8322.t28 gnd 0.100161f
C715 a_n2982_8322.t18 gnd 0.100161f
C716 a_n2982_8322.n2 gnd 0.705534f
C717 a_n2982_8322.n3 gnd 0.40054f
C718 a_n2982_8322.t9 gnd 0.100161f
C719 a_n2982_8322.t8 gnd 0.100161f
C720 a_n2982_8322.n4 gnd 0.705534f
C721 a_n2982_8322.n5 gnd 0.40054f
C722 a_n2982_8322.t22 gnd 0.100161f
C723 a_n2982_8322.t15 gnd 0.100161f
C724 a_n2982_8322.n6 gnd 0.705534f
C725 a_n2982_8322.n7 gnd 0.40054f
C726 a_n2982_8322.t19 gnd 0.100161f
C727 a_n2982_8322.t17 gnd 0.100161f
C728 a_n2982_8322.n8 gnd 0.705534f
C729 a_n2982_8322.n9 gnd 0.40054f
C730 a_n2982_8322.t6 gnd 0.935989f
C731 a_n2982_8322.n10 gnd 1.87142f
C732 a_n2982_8322.t33 gnd 0.937857f
C733 a_n2982_8322.t37 gnd 0.100161f
C734 a_n2982_8322.t36 gnd 0.100161f
C735 a_n2982_8322.n11 gnd 0.705534f
C736 a_n2982_8322.n12 gnd 0.78833f
C737 a_n2982_8322.t31 gnd 0.935989f
C738 a_n2982_8322.n13 gnd 0.396699f
C739 a_n2982_8322.t34 gnd 0.935989f
C740 a_n2982_8322.n14 gnd 0.396699f
C741 a_n2982_8322.t32 gnd 0.100161f
C742 a_n2982_8322.t30 gnd 0.100161f
C743 a_n2982_8322.n15 gnd 0.705534f
C744 a_n2982_8322.n16 gnd 0.40054f
C745 a_n2982_8322.t35 gnd 0.935989f
C746 a_n2982_8322.n17 gnd 1.47142f
C747 a_n2982_8322.n18 gnd 2.35138f
C748 a_n2982_8322.n19 gnd 3.33814f
C749 a_n2982_8322.t7 gnd 0.935989f
C750 a_n2982_8322.n20 gnd 1.11148f
C751 a_n2982_8322.t24 gnd 0.100161f
C752 a_n2982_8322.t23 gnd 0.100161f
C753 a_n2982_8322.n21 gnd 0.705534f
C754 a_n2982_8322.n22 gnd 0.40054f
C755 a_n2982_8322.t11 gnd 0.100161f
C756 a_n2982_8322.t10 gnd 0.100161f
C757 a_n2982_8322.n23 gnd 0.705534f
C758 a_n2982_8322.n24 gnd 0.40054f
C759 a_n2982_8322.t26 gnd 0.100161f
C760 a_n2982_8322.t14 gnd 0.100161f
C761 a_n2982_8322.n25 gnd 0.705534f
C762 a_n2982_8322.n26 gnd 0.40054f
C763 a_n2982_8322.t27 gnd 0.937854f
C764 a_n2982_8322.t20 gnd 0.100161f
C765 a_n2982_8322.t16 gnd 0.100161f
C766 a_n2982_8322.n27 gnd 0.705534f
C767 a_n2982_8322.n28 gnd 0.788332f
C768 a_n2982_8322.n29 gnd 0.400539f
C769 a_n2982_8322.n30 gnd 0.705536f
C770 a_n2982_8322.t29 gnd 0.100161f
C771 a_n9628_8799.n0 gnd 0.21338f
C772 a_n9628_8799.n1 gnd 0.292999f
C773 a_n9628_8799.n2 gnd 0.21338f
C774 a_n9628_8799.n3 gnd 0.21338f
C775 a_n9628_8799.n4 gnd 0.21338f
C776 a_n9628_8799.n5 gnd 0.21338f
C777 a_n9628_8799.n6 gnd 0.21338f
C778 a_n9628_8799.n7 gnd 0.221877f
C779 a_n9628_8799.n8 gnd 0.21338f
C780 a_n9628_8799.n9 gnd 0.292999f
C781 a_n9628_8799.n10 gnd 0.21338f
C782 a_n9628_8799.n11 gnd 0.21338f
C783 a_n9628_8799.n12 gnd 0.21338f
C784 a_n9628_8799.n13 gnd 0.21338f
C785 a_n9628_8799.n14 gnd 0.21338f
C786 a_n9628_8799.n15 gnd 0.221877f
C787 a_n9628_8799.n16 gnd 0.21338f
C788 a_n9628_8799.n17 gnd 0.462488f
C789 a_n9628_8799.n18 gnd 0.21338f
C790 a_n9628_8799.n19 gnd 0.21338f
C791 a_n9628_8799.n20 gnd 0.21338f
C792 a_n9628_8799.n21 gnd 0.21338f
C793 a_n9628_8799.n22 gnd 0.21338f
C794 a_n9628_8799.n23 gnd 0.221877f
C795 a_n9628_8799.n24 gnd 0.21338f
C796 a_n9628_8799.n25 gnd 0.328567f
C797 a_n9628_8799.n26 gnd 0.21338f
C798 a_n9628_8799.n27 gnd 0.21338f
C799 a_n9628_8799.n28 gnd 0.21338f
C800 a_n9628_8799.n29 gnd 0.21338f
C801 a_n9628_8799.n30 gnd 0.21338f
C802 a_n9628_8799.n31 gnd 0.186309f
C803 a_n9628_8799.n32 gnd 0.21338f
C804 a_n9628_8799.n33 gnd 0.328567f
C805 a_n9628_8799.n34 gnd 0.21338f
C806 a_n9628_8799.n35 gnd 0.21338f
C807 a_n9628_8799.n36 gnd 0.21338f
C808 a_n9628_8799.n37 gnd 0.21338f
C809 a_n9628_8799.n38 gnd 0.21338f
C810 a_n9628_8799.n39 gnd 0.186309f
C811 a_n9628_8799.n40 gnd 0.21338f
C812 a_n9628_8799.n41 gnd 0.328567f
C813 a_n9628_8799.n42 gnd 0.21338f
C814 a_n9628_8799.n43 gnd 0.21338f
C815 a_n9628_8799.n44 gnd 0.21338f
C816 a_n9628_8799.n45 gnd 0.21338f
C817 a_n9628_8799.n46 gnd 0.21338f
C818 a_n9628_8799.n47 gnd 0.355798f
C819 a_n9628_8799.n48 gnd 3.50187f
C820 a_n9628_8799.n49 gnd 1.78557f
C821 a_n9628_8799.n50 gnd 3.03803f
C822 a_n9628_8799.n51 gnd 1.56391f
C823 a_n9628_8799.n52 gnd 1.03271f
C824 a_n9628_8799.n53 gnd 3.09742f
C825 a_n9628_8799.n54 gnd 1.03271f
C826 a_n9628_8799.n55 gnd 0.718386f
C827 a_n9628_8799.n56 gnd 0.25689f
C828 a_n9628_8799.n57 gnd 0.003756f
C829 a_n9628_8799.n58 gnd 0.0099f
C830 a_n9628_8799.n59 gnd 0.010816f
C831 a_n9628_8799.n60 gnd 0.005716f
C832 a_n9628_8799.n62 gnd 0.004796f
C833 a_n9628_8799.n63 gnd 0.010372f
C834 a_n9628_8799.n64 gnd 0.010372f
C835 a_n9628_8799.n65 gnd 0.004796f
C836 a_n9628_8799.n67 gnd 0.005716f
C837 a_n9628_8799.n68 gnd 0.010816f
C838 a_n9628_8799.n69 gnd 0.0099f
C839 a_n9628_8799.n70 gnd 0.003756f
C840 a_n9628_8799.n71 gnd 0.25689f
C841 a_n9628_8799.n72 gnd 0.003756f
C842 a_n9628_8799.n73 gnd 0.0099f
C843 a_n9628_8799.n74 gnd 0.010816f
C844 a_n9628_8799.n75 gnd 0.005716f
C845 a_n9628_8799.n77 gnd 0.004796f
C846 a_n9628_8799.n78 gnd 0.010372f
C847 a_n9628_8799.n79 gnd 0.010372f
C848 a_n9628_8799.n80 gnd 0.004796f
C849 a_n9628_8799.n82 gnd 0.005716f
C850 a_n9628_8799.n83 gnd 0.010816f
C851 a_n9628_8799.n84 gnd 0.0099f
C852 a_n9628_8799.n85 gnd 0.003756f
C853 a_n9628_8799.n86 gnd 0.25689f
C854 a_n9628_8799.n87 gnd 0.003756f
C855 a_n9628_8799.n88 gnd 0.0099f
C856 a_n9628_8799.n89 gnd 0.010816f
C857 a_n9628_8799.n90 gnd 0.005716f
C858 a_n9628_8799.n92 gnd 0.004796f
C859 a_n9628_8799.n93 gnd 0.010372f
C860 a_n9628_8799.n94 gnd 0.010372f
C861 a_n9628_8799.n95 gnd 0.004796f
C862 a_n9628_8799.n97 gnd 0.005716f
C863 a_n9628_8799.n98 gnd 0.010816f
C864 a_n9628_8799.n99 gnd 0.0099f
C865 a_n9628_8799.n100 gnd 0.003756f
C866 a_n9628_8799.n101 gnd 0.003756f
C867 a_n9628_8799.n102 gnd 0.0099f
C868 a_n9628_8799.n103 gnd 0.010816f
C869 a_n9628_8799.n104 gnd 0.005716f
C870 a_n9628_8799.n106 gnd 0.004796f
C871 a_n9628_8799.n107 gnd 0.010372f
C872 a_n9628_8799.n108 gnd 0.010372f
C873 a_n9628_8799.n109 gnd 0.004796f
C874 a_n9628_8799.n111 gnd 0.005716f
C875 a_n9628_8799.n112 gnd 0.010816f
C876 a_n9628_8799.n113 gnd 0.0099f
C877 a_n9628_8799.n114 gnd 0.003756f
C878 a_n9628_8799.n115 gnd 0.25689f
C879 a_n9628_8799.n116 gnd 0.003756f
C880 a_n9628_8799.n117 gnd 0.0099f
C881 a_n9628_8799.n118 gnd 0.010816f
C882 a_n9628_8799.n119 gnd 0.005716f
C883 a_n9628_8799.n121 gnd 0.004796f
C884 a_n9628_8799.n122 gnd 0.010372f
C885 a_n9628_8799.n123 gnd 0.010372f
C886 a_n9628_8799.n124 gnd 0.004796f
C887 a_n9628_8799.n126 gnd 0.005716f
C888 a_n9628_8799.n127 gnd 0.010816f
C889 a_n9628_8799.n128 gnd 0.0099f
C890 a_n9628_8799.n129 gnd 0.003756f
C891 a_n9628_8799.n130 gnd 0.25689f
C892 a_n9628_8799.n131 gnd 0.003756f
C893 a_n9628_8799.n132 gnd 0.0099f
C894 a_n9628_8799.n133 gnd 0.010816f
C895 a_n9628_8799.n134 gnd 0.005716f
C896 a_n9628_8799.n136 gnd 0.004796f
C897 a_n9628_8799.n137 gnd 0.010372f
C898 a_n9628_8799.n138 gnd 0.010372f
C899 a_n9628_8799.n139 gnd 0.004796f
C900 a_n9628_8799.n141 gnd 0.005716f
C901 a_n9628_8799.n142 gnd 0.010816f
C902 a_n9628_8799.n143 gnd 0.0099f
C903 a_n9628_8799.n144 gnd 0.003756f
C904 a_n9628_8799.n145 gnd 0.25689f
C905 a_n9628_8799.t28 gnd 0.148003f
C906 a_n9628_8799.t41 gnd 0.148003f
C907 a_n9628_8799.t34 gnd 0.148003f
C908 a_n9628_8799.n146 gnd 1.16732f
C909 a_n9628_8799.t27 gnd 0.148003f
C910 a_n9628_8799.t30 gnd 0.148003f
C911 a_n9628_8799.n147 gnd 1.16732f
C912 a_n9628_8799.t24 gnd 0.148003f
C913 a_n9628_8799.t31 gnd 0.148003f
C914 a_n9628_8799.n148 gnd 1.1654f
C915 a_n9628_8799.t35 gnd 0.148003f
C916 a_n9628_8799.t38 gnd 0.148003f
C917 a_n9628_8799.n149 gnd 1.1654f
C918 a_n9628_8799.t39 gnd 0.148003f
C919 a_n9628_8799.t29 gnd 0.148003f
C920 a_n9628_8799.n150 gnd 1.1654f
C921 a_n9628_8799.t22 gnd 0.148003f
C922 a_n9628_8799.t40 gnd 0.148003f
C923 a_n9628_8799.n151 gnd 1.1654f
C924 a_n9628_8799.t42 gnd 0.148003f
C925 a_n9628_8799.t25 gnd 0.148003f
C926 a_n9628_8799.n152 gnd 1.1654f
C927 a_n9628_8799.n153 gnd 3.77696f
C928 a_n9628_8799.t19 gnd 0.115113f
C929 a_n9628_8799.t47 gnd 0.115113f
C930 a_n9628_8799.n154 gnd 1.0188f
C931 a_n9628_8799.t5 gnd 0.115113f
C932 a_n9628_8799.t15 gnd 0.115113f
C933 a_n9628_8799.n155 gnd 1.01718f
C934 a_n9628_8799.t4 gnd 0.115113f
C935 a_n9628_8799.t6 gnd 0.115113f
C936 a_n9628_8799.n156 gnd 1.01718f
C937 a_n9628_8799.t20 gnd 0.115113f
C938 a_n9628_8799.t10 gnd 0.115113f
C939 a_n9628_8799.n157 gnd 1.0188f
C940 a_n9628_8799.t3 gnd 0.115113f
C941 a_n9628_8799.t46 gnd 0.115113f
C942 a_n9628_8799.n158 gnd 1.01718f
C943 a_n9628_8799.t11 gnd 0.115113f
C944 a_n9628_8799.t2 gnd 0.115113f
C945 a_n9628_8799.n159 gnd 1.01718f
C946 a_n9628_8799.t12 gnd 0.115113f
C947 a_n9628_8799.t17 gnd 0.115113f
C948 a_n9628_8799.n160 gnd 1.0188f
C949 a_n9628_8799.t1 gnd 0.115113f
C950 a_n9628_8799.t0 gnd 0.115113f
C951 a_n9628_8799.n161 gnd 1.01718f
C952 a_n9628_8799.t45 gnd 0.115113f
C953 a_n9628_8799.t9 gnd 0.115113f
C954 a_n9628_8799.n162 gnd 1.01718f
C955 a_n9628_8799.t16 gnd 0.115113f
C956 a_n9628_8799.t18 gnd 0.115113f
C957 a_n9628_8799.n163 gnd 1.01718f
C958 a_n9628_8799.t13 gnd 0.115113f
C959 a_n9628_8799.t14 gnd 0.115113f
C960 a_n9628_8799.n164 gnd 1.01718f
C961 a_n9628_8799.t7 gnd 0.115113f
C962 a_n9628_8799.t8 gnd 0.115113f
C963 a_n9628_8799.n165 gnd 1.01718f
C964 a_n9628_8799.t94 gnd 0.613689f
C965 a_n9628_8799.n166 gnd 0.276291f
C966 a_n9628_8799.t130 gnd 0.613689f
C967 a_n9628_8799.t151 gnd 0.613689f
C968 a_n9628_8799.n167 gnd 0.27827f
C969 a_n9628_8799.t152 gnd 0.613689f
C970 a_n9628_8799.t80 gnd 0.613689f
C971 a_n9628_8799.n168 gnd 0.27129f
C972 a_n9628_8799.t120 gnd 0.613689f
C973 a_n9628_8799.t128 gnd 0.613689f
C974 a_n9628_8799.n169 gnd 0.275374f
C975 a_n9628_8799.t56 gnd 0.613689f
C976 a_n9628_8799.t99 gnd 0.613689f
C977 a_n9628_8799.t98 gnd 0.625304f
C978 a_n9628_8799.n170 gnd 0.257263f
C979 a_n9628_8799.n171 gnd 0.278653f
C980 a_n9628_8799.t131 gnd 0.613689f
C981 a_n9628_8799.n172 gnd 0.276291f
C982 a_n9628_8799.n173 gnd 0.271948f
C983 a_n9628_8799.t96 gnd 0.613689f
C984 a_n9628_8799.n174 gnd 0.270632f
C985 a_n9628_8799.t50 gnd 0.613689f
C986 a_n9628_8799.n175 gnd 0.278008f
C987 a_n9628_8799.t81 gnd 0.613689f
C988 a_n9628_8799.n176 gnd 0.27827f
C989 a_n9628_8799.n177 gnd 0.275818f
C990 a_n9628_8799.t155 gnd 0.613689f
C991 a_n9628_8799.n178 gnd 0.27129f
C992 a_n9628_8799.t116 gnd 0.613689f
C993 a_n9628_8799.n179 gnd 0.275818f
C994 a_n9628_8799.n180 gnd 0.278008f
C995 a_n9628_8799.t97 gnd 0.613689f
C996 a_n9628_8799.n181 gnd 0.275374f
C997 a_n9628_8799.n182 gnd 0.270632f
C998 a_n9628_8799.t150 gnd 0.613689f
C999 a_n9628_8799.n183 gnd 0.271948f
C1000 a_n9628_8799.t95 gnd 0.613689f
C1001 a_n9628_8799.n184 gnd 0.278653f
C1002 a_n9628_8799.t127 gnd 0.625294f
C1003 a_n9628_8799.t105 gnd 0.613689f
C1004 a_n9628_8799.n185 gnd 0.276291f
C1005 a_n9628_8799.t144 gnd 0.613689f
C1006 a_n9628_8799.t163 gnd 0.613689f
C1007 a_n9628_8799.n186 gnd 0.27827f
C1008 a_n9628_8799.t165 gnd 0.613689f
C1009 a_n9628_8799.t89 gnd 0.613689f
C1010 a_n9628_8799.n187 gnd 0.27129f
C1011 a_n9628_8799.t133 gnd 0.613689f
C1012 a_n9628_8799.t140 gnd 0.613689f
C1013 a_n9628_8799.n188 gnd 0.275374f
C1014 a_n9628_8799.t68 gnd 0.613689f
C1015 a_n9628_8799.t112 gnd 0.613689f
C1016 a_n9628_8799.t110 gnd 0.625304f
C1017 a_n9628_8799.n189 gnd 0.257263f
C1018 a_n9628_8799.n190 gnd 0.278653f
C1019 a_n9628_8799.t148 gnd 0.613689f
C1020 a_n9628_8799.n191 gnd 0.276291f
C1021 a_n9628_8799.n192 gnd 0.271948f
C1022 a_n9628_8799.t106 gnd 0.613689f
C1023 a_n9628_8799.n193 gnd 0.270632f
C1024 a_n9628_8799.t64 gnd 0.613689f
C1025 a_n9628_8799.n194 gnd 0.278008f
C1026 a_n9628_8799.t92 gnd 0.613689f
C1027 a_n9628_8799.n195 gnd 0.27827f
C1028 a_n9628_8799.n196 gnd 0.275818f
C1029 a_n9628_8799.t167 gnd 0.613689f
C1030 a_n9628_8799.n197 gnd 0.27129f
C1031 a_n9628_8799.t129 gnd 0.613689f
C1032 a_n9628_8799.n198 gnd 0.275818f
C1033 a_n9628_8799.n199 gnd 0.278008f
C1034 a_n9628_8799.t111 gnd 0.613689f
C1035 a_n9628_8799.n200 gnd 0.275374f
C1036 a_n9628_8799.n201 gnd 0.270632f
C1037 a_n9628_8799.t162 gnd 0.613689f
C1038 a_n9628_8799.n202 gnd 0.271948f
C1039 a_n9628_8799.t107 gnd 0.613689f
C1040 a_n9628_8799.n203 gnd 0.278653f
C1041 a_n9628_8799.t141 gnd 0.625294f
C1042 a_n9628_8799.n204 gnd 0.922596f
C1043 a_n9628_8799.t71 gnd 0.613689f
C1044 a_n9628_8799.n205 gnd 0.276291f
C1045 a_n9628_8799.t90 gnd 0.613689f
C1046 a_n9628_8799.t124 gnd 0.613689f
C1047 a_n9628_8799.n206 gnd 0.27827f
C1048 a_n9628_8799.t104 gnd 0.613689f
C1049 a_n9628_8799.t108 gnd 0.613689f
C1050 a_n9628_8799.n207 gnd 0.27129f
C1051 a_n9628_8799.t135 gnd 0.613689f
C1052 a_n9628_8799.t51 gnd 0.613689f
C1053 a_n9628_8799.n208 gnd 0.275374f
C1054 a_n9628_8799.t77 gnd 0.613689f
C1055 a_n9628_8799.t60 gnd 0.613689f
C1056 a_n9628_8799.t82 gnd 0.625304f
C1057 a_n9628_8799.n209 gnd 0.257263f
C1058 a_n9628_8799.n210 gnd 0.278653f
C1059 a_n9628_8799.t122 gnd 0.613689f
C1060 a_n9628_8799.n211 gnd 0.276291f
C1061 a_n9628_8799.n212 gnd 0.271948f
C1062 a_n9628_8799.t100 gnd 0.613689f
C1063 a_n9628_8799.n213 gnd 0.270632f
C1064 a_n9628_8799.t117 gnd 0.613689f
C1065 a_n9628_8799.n214 gnd 0.278008f
C1066 a_n9628_8799.t69 gnd 0.613689f
C1067 a_n9628_8799.n215 gnd 0.27827f
C1068 a_n9628_8799.n216 gnd 0.275818f
C1069 a_n9628_8799.t85 gnd 0.613689f
C1070 a_n9628_8799.n217 gnd 0.27129f
C1071 a_n9628_8799.t61 gnd 0.613689f
C1072 a_n9628_8799.n218 gnd 0.275818f
C1073 a_n9628_8799.n219 gnd 0.278008f
C1074 a_n9628_8799.t143 gnd 0.613689f
C1075 a_n9628_8799.n220 gnd 0.275374f
C1076 a_n9628_8799.n221 gnd 0.270632f
C1077 a_n9628_8799.t153 gnd 0.613689f
C1078 a_n9628_8799.n222 gnd 0.271948f
C1079 a_n9628_8799.t48 gnd 0.613689f
C1080 a_n9628_8799.n223 gnd 0.278653f
C1081 a_n9628_8799.t113 gnd 0.625294f
C1082 a_n9628_8799.n224 gnd 1.89486f
C1083 a_n9628_8799.t55 gnd 0.625294f
C1084 a_n9628_8799.t53 gnd 0.613689f
C1085 a_n9628_8799.t139 gnd 0.613689f
C1086 a_n9628_8799.n225 gnd 0.276291f
C1087 a_n9628_8799.t75 gnd 0.613689f
C1088 a_n9628_8799.t58 gnd 0.613689f
C1089 a_n9628_8799.t146 gnd 0.613689f
C1090 a_n9628_8799.n226 gnd 0.275374f
C1091 a_n9628_8799.t101 gnd 0.613689f
C1092 a_n9628_8799.t76 gnd 0.613689f
C1093 a_n9628_8799.t164 gnd 0.613689f
C1094 a_n9628_8799.n227 gnd 0.275818f
C1095 a_n9628_8799.t119 gnd 0.613689f
C1096 a_n9628_8799.t79 gnd 0.613689f
C1097 a_n9628_8799.t158 gnd 0.613689f
C1098 a_n9628_8799.n228 gnd 0.275818f
C1099 a_n9628_8799.t121 gnd 0.613689f
C1100 a_n9628_8799.t93 gnd 0.613689f
C1101 a_n9628_8799.t54 gnd 0.613689f
C1102 a_n9628_8799.n229 gnd 0.275374f
C1103 a_n9628_8799.t142 gnd 0.613689f
C1104 a_n9628_8799.t123 gnd 0.613689f
C1105 a_n9628_8799.t59 gnd 0.613689f
C1106 a_n9628_8799.n230 gnd 0.276291f
C1107 a_n9628_8799.t145 gnd 0.625304f
C1108 a_n9628_8799.n231 gnd 0.257263f
C1109 a_n9628_8799.t149 gnd 0.613689f
C1110 a_n9628_8799.n232 gnd 0.278653f
C1111 a_n9628_8799.n233 gnd 0.271948f
C1112 a_n9628_8799.n234 gnd 0.270632f
C1113 a_n9628_8799.n235 gnd 0.278008f
C1114 a_n9628_8799.n236 gnd 0.27827f
C1115 a_n9628_8799.n237 gnd 0.27129f
C1116 a_n9628_8799.n238 gnd 0.27129f
C1117 a_n9628_8799.n239 gnd 0.27827f
C1118 a_n9628_8799.n240 gnd 0.278008f
C1119 a_n9628_8799.n241 gnd 0.270632f
C1120 a_n9628_8799.n242 gnd 0.271948f
C1121 a_n9628_8799.n243 gnd 0.278653f
C1122 a_n9628_8799.t67 gnd 0.625294f
C1123 a_n9628_8799.t65 gnd 0.613689f
C1124 a_n9628_8799.t156 gnd 0.613689f
C1125 a_n9628_8799.n244 gnd 0.276291f
C1126 a_n9628_8799.t84 gnd 0.613689f
C1127 a_n9628_8799.t73 gnd 0.613689f
C1128 a_n9628_8799.t160 gnd 0.613689f
C1129 a_n9628_8799.n245 gnd 0.275374f
C1130 a_n9628_8799.t115 gnd 0.613689f
C1131 a_n9628_8799.t87 gnd 0.613689f
C1132 a_n9628_8799.t57 gnd 0.613689f
C1133 a_n9628_8799.n246 gnd 0.275818f
C1134 a_n9628_8799.t132 gnd 0.613689f
C1135 a_n9628_8799.t88 gnd 0.613689f
C1136 a_n9628_8799.t49 gnd 0.613689f
C1137 a_n9628_8799.n247 gnd 0.275818f
C1138 a_n9628_8799.t137 gnd 0.613689f
C1139 a_n9628_8799.t103 gnd 0.613689f
C1140 a_n9628_8799.t66 gnd 0.613689f
C1141 a_n9628_8799.n248 gnd 0.275374f
C1142 a_n9628_8799.t157 gnd 0.613689f
C1143 a_n9628_8799.t138 gnd 0.613689f
C1144 a_n9628_8799.t74 gnd 0.613689f
C1145 a_n9628_8799.n249 gnd 0.276291f
C1146 a_n9628_8799.t159 gnd 0.625304f
C1147 a_n9628_8799.n250 gnd 0.257263f
C1148 a_n9628_8799.t161 gnd 0.613689f
C1149 a_n9628_8799.n251 gnd 0.278653f
C1150 a_n9628_8799.n252 gnd 0.271948f
C1151 a_n9628_8799.n253 gnd 0.270632f
C1152 a_n9628_8799.n254 gnd 0.278008f
C1153 a_n9628_8799.n255 gnd 0.27827f
C1154 a_n9628_8799.n256 gnd 0.27129f
C1155 a_n9628_8799.n257 gnd 0.27129f
C1156 a_n9628_8799.n258 gnd 0.27827f
C1157 a_n9628_8799.n259 gnd 0.278008f
C1158 a_n9628_8799.n260 gnd 0.270632f
C1159 a_n9628_8799.n261 gnd 0.271948f
C1160 a_n9628_8799.n262 gnd 0.278653f
C1161 a_n9628_8799.n263 gnd 0.922596f
C1162 a_n9628_8799.t114 gnd 0.625294f
C1163 a_n9628_8799.t136 gnd 0.613689f
C1164 a_n9628_8799.t72 gnd 0.613689f
C1165 a_n9628_8799.n264 gnd 0.276291f
C1166 a_n9628_8799.t154 gnd 0.613689f
C1167 a_n9628_8799.t91 gnd 0.613689f
C1168 a_n9628_8799.t147 gnd 0.613689f
C1169 a_n9628_8799.n265 gnd 0.275374f
C1170 a_n9628_8799.t78 gnd 0.613689f
C1171 a_n9628_8799.t126 gnd 0.613689f
C1172 a_n9628_8799.t63 gnd 0.613689f
C1173 a_n9628_8799.n266 gnd 0.275818f
C1174 a_n9628_8799.t109 gnd 0.613689f
C1175 a_n9628_8799.t86 gnd 0.613689f
C1176 a_n9628_8799.t134 gnd 0.613689f
C1177 a_n9628_8799.n267 gnd 0.275818f
C1178 a_n9628_8799.t70 gnd 0.613689f
C1179 a_n9628_8799.t118 gnd 0.613689f
C1180 a_n9628_8799.t52 gnd 0.613689f
C1181 a_n9628_8799.n268 gnd 0.275374f
C1182 a_n9628_8799.t102 gnd 0.613689f
C1183 a_n9628_8799.t166 gnd 0.613689f
C1184 a_n9628_8799.t125 gnd 0.613689f
C1185 a_n9628_8799.n269 gnd 0.276291f
C1186 a_n9628_8799.t83 gnd 0.625304f
C1187 a_n9628_8799.n270 gnd 0.257263f
C1188 a_n9628_8799.t62 gnd 0.613689f
C1189 a_n9628_8799.n271 gnd 0.278653f
C1190 a_n9628_8799.n272 gnd 0.271948f
C1191 a_n9628_8799.n273 gnd 0.270632f
C1192 a_n9628_8799.n274 gnd 0.278008f
C1193 a_n9628_8799.n275 gnd 0.27827f
C1194 a_n9628_8799.n276 gnd 0.27129f
C1195 a_n9628_8799.n277 gnd 0.27129f
C1196 a_n9628_8799.n278 gnd 0.27827f
C1197 a_n9628_8799.n279 gnd 0.278008f
C1198 a_n9628_8799.n280 gnd 0.270632f
C1199 a_n9628_8799.n281 gnd 0.271948f
C1200 a_n9628_8799.n282 gnd 0.278653f
C1201 a_n9628_8799.n283 gnd 1.45394f
C1202 a_n9628_8799.n284 gnd 17.8366f
C1203 a_n9628_8799.n285 gnd 4.49131f
C1204 a_n9628_8799.n286 gnd 7.8322f
C1205 a_n9628_8799.t32 gnd 0.148003f
C1206 a_n9628_8799.t37 gnd 0.148003f
C1207 a_n9628_8799.n287 gnd 1.1654f
C1208 a_n9628_8799.t33 gnd 0.148003f
C1209 a_n9628_8799.t26 gnd 0.148003f
C1210 a_n9628_8799.n288 gnd 1.1654f
C1211 a_n9628_8799.t43 gnd 0.148003f
C1212 a_n9628_8799.t23 gnd 0.148003f
C1213 a_n9628_8799.n289 gnd 1.1654f
C1214 a_n9628_8799.t36 gnd 0.148003f
C1215 a_n9628_8799.t44 gnd 0.148003f
C1216 a_n9628_8799.n290 gnd 1.1654f
C1217 a_n9628_8799.n291 gnd 1.04755f
C1218 a_n9628_8799.n292 gnd 1.1654f
C1219 a_n9628_8799.t21 gnd 0.148003f
C1220 CSoutput.n0 gnd 0.049305f
C1221 CSoutput.t226 gnd 0.326143f
C1222 CSoutput.n1 gnd 0.14727f
C1223 CSoutput.n2 gnd 0.049305f
C1224 CSoutput.t224 gnd 0.326143f
C1225 CSoutput.n3 gnd 0.039078f
C1226 CSoutput.n4 gnd 0.049305f
C1227 CSoutput.t236 gnd 0.326143f
C1228 CSoutput.n5 gnd 0.033698f
C1229 CSoutput.n6 gnd 0.049305f
C1230 CSoutput.t221 gnd 0.326143f
C1231 CSoutput.t231 gnd 0.326143f
C1232 CSoutput.n7 gnd 0.145665f
C1233 CSoutput.n8 gnd 0.049305f
C1234 CSoutput.t234 gnd 0.326143f
C1235 CSoutput.n9 gnd 0.032129f
C1236 CSoutput.n10 gnd 0.049305f
C1237 CSoutput.t217 gnd 0.326143f
C1238 CSoutput.t223 gnd 0.326143f
C1239 CSoutput.n11 gnd 0.145665f
C1240 CSoutput.n12 gnd 0.049305f
C1241 CSoutput.t228 gnd 0.326143f
C1242 CSoutput.n13 gnd 0.033698f
C1243 CSoutput.n14 gnd 0.049305f
C1244 CSoutput.t237 gnd 0.326143f
C1245 CSoutput.t220 gnd 0.326143f
C1246 CSoutput.n15 gnd 0.145665f
C1247 CSoutput.n16 gnd 0.049305f
C1248 CSoutput.t227 gnd 0.326143f
C1249 CSoutput.n17 gnd 0.035991f
C1250 CSoutput.t216 gnd 0.38975f
C1251 CSoutput.t225 gnd 0.326143f
C1252 CSoutput.n18 gnd 0.185957f
C1253 CSoutput.n19 gnd 0.180443f
C1254 CSoutput.n20 gnd 0.209335f
C1255 CSoutput.n21 gnd 0.049305f
C1256 CSoutput.n22 gnd 0.041151f
C1257 CSoutput.n23 gnd 0.145665f
C1258 CSoutput.n24 gnd 0.039668f
C1259 CSoutput.n25 gnd 0.039078f
C1260 CSoutput.n26 gnd 0.049305f
C1261 CSoutput.n27 gnd 0.049305f
C1262 CSoutput.n28 gnd 0.040834f
C1263 CSoutput.n29 gnd 0.034669f
C1264 CSoutput.n30 gnd 0.148907f
C1265 CSoutput.n31 gnd 0.035147f
C1266 CSoutput.n32 gnd 0.049305f
C1267 CSoutput.n33 gnd 0.049305f
C1268 CSoutput.n34 gnd 0.049305f
C1269 CSoutput.n35 gnd 0.040399f
C1270 CSoutput.n36 gnd 0.145665f
C1271 CSoutput.n37 gnd 0.038636f
C1272 CSoutput.n38 gnd 0.04011f
C1273 CSoutput.n39 gnd 0.049305f
C1274 CSoutput.n40 gnd 0.049305f
C1275 CSoutput.n41 gnd 0.041142f
C1276 CSoutput.n42 gnd 0.037604f
C1277 CSoutput.n43 gnd 0.145665f
C1278 CSoutput.n44 gnd 0.038557f
C1279 CSoutput.n45 gnd 0.049305f
C1280 CSoutput.n46 gnd 0.049305f
C1281 CSoutput.n47 gnd 0.049305f
C1282 CSoutput.n48 gnd 0.038557f
C1283 CSoutput.n49 gnd 0.145665f
C1284 CSoutput.n50 gnd 0.037604f
C1285 CSoutput.n51 gnd 0.041142f
C1286 CSoutput.n52 gnd 0.049305f
C1287 CSoutput.n53 gnd 0.049305f
C1288 CSoutput.n54 gnd 0.04011f
C1289 CSoutput.n55 gnd 0.038636f
C1290 CSoutput.n56 gnd 0.145665f
C1291 CSoutput.n57 gnd 0.040399f
C1292 CSoutput.n58 gnd 0.049305f
C1293 CSoutput.n59 gnd 0.049305f
C1294 CSoutput.n60 gnd 0.049305f
C1295 CSoutput.n61 gnd 0.035147f
C1296 CSoutput.n62 gnd 0.148907f
C1297 CSoutput.n63 gnd 0.034669f
C1298 CSoutput.t232 gnd 0.326143f
C1299 CSoutput.n64 gnd 0.145665f
C1300 CSoutput.n65 gnd 0.040834f
C1301 CSoutput.n66 gnd 0.049305f
C1302 CSoutput.n67 gnd 0.049305f
C1303 CSoutput.n68 gnd 0.049305f
C1304 CSoutput.n69 gnd 0.039668f
C1305 CSoutput.n70 gnd 0.145665f
C1306 CSoutput.n71 gnd 0.041151f
C1307 CSoutput.n72 gnd 0.035991f
C1308 CSoutput.n73 gnd 0.049305f
C1309 CSoutput.n74 gnd 0.049305f
C1310 CSoutput.n75 gnd 0.037325f
C1311 CSoutput.n76 gnd 0.022167f
C1312 CSoutput.t218 gnd 0.366445f
C1313 CSoutput.n77 gnd 0.182035f
C1314 CSoutput.n78 gnd 0.744586f
C1315 CSoutput.t200 gnd 0.061501f
C1316 CSoutput.t15 gnd 0.061501f
C1317 CSoutput.n79 gnd 0.476163f
C1318 CSoutput.t147 gnd 0.061501f
C1319 CSoutput.t197 gnd 0.061501f
C1320 CSoutput.n80 gnd 0.475314f
C1321 CSoutput.n81 gnd 0.482443f
C1322 CSoutput.t149 gnd 0.061501f
C1323 CSoutput.t0 gnd 0.061501f
C1324 CSoutput.n82 gnd 0.475314f
C1325 CSoutput.n83 gnd 0.237728f
C1326 CSoutput.t140 gnd 0.061501f
C1327 CSoutput.t142 gnd 0.061501f
C1328 CSoutput.n84 gnd 0.475314f
C1329 CSoutput.n85 gnd 0.237728f
C1330 CSoutput.t6 gnd 0.061501f
C1331 CSoutput.t199 gnd 0.061501f
C1332 CSoutput.n86 gnd 0.475314f
C1333 CSoutput.n87 gnd 0.237728f
C1334 CSoutput.t165 gnd 0.061501f
C1335 CSoutput.t157 gnd 0.061501f
C1336 CSoutput.n88 gnd 0.475314f
C1337 CSoutput.n89 gnd 0.237728f
C1338 CSoutput.t171 gnd 0.061501f
C1339 CSoutput.t173 gnd 0.061501f
C1340 CSoutput.n90 gnd 0.475314f
C1341 CSoutput.n91 gnd 0.237728f
C1342 CSoutput.t208 gnd 0.061501f
C1343 CSoutput.t215 gnd 0.061501f
C1344 CSoutput.n92 gnd 0.475314f
C1345 CSoutput.n93 gnd 0.237728f
C1346 CSoutput.t138 gnd 0.061501f
C1347 CSoutput.t127 gnd 0.061501f
C1348 CSoutput.n94 gnd 0.475314f
C1349 CSoutput.n95 gnd 0.237728f
C1350 CSoutput.t8 gnd 0.061501f
C1351 CSoutput.t198 gnd 0.061501f
C1352 CSoutput.n96 gnd 0.475314f
C1353 CSoutput.n97 gnd 0.435938f
C1354 CSoutput.t189 gnd 0.061501f
C1355 CSoutput.t207 gnd 0.061501f
C1356 CSoutput.n98 gnd 0.476163f
C1357 CSoutput.t144 gnd 0.061501f
C1358 CSoutput.t143 gnd 0.061501f
C1359 CSoutput.n99 gnd 0.475314f
C1360 CSoutput.n100 gnd 0.482443f
C1361 CSoutput.t151 gnd 0.061501f
C1362 CSoutput.t122 gnd 0.061501f
C1363 CSoutput.n101 gnd 0.475314f
C1364 CSoutput.n102 gnd 0.237728f
C1365 CSoutput.t145 gnd 0.061501f
C1366 CSoutput.t121 gnd 0.061501f
C1367 CSoutput.n103 gnd 0.475314f
C1368 CSoutput.n104 gnd 0.237728f
C1369 CSoutput.t13 gnd 0.061501f
C1370 CSoutput.t117 gnd 0.061501f
C1371 CSoutput.n105 gnd 0.475314f
C1372 CSoutput.n106 gnd 0.237728f
C1373 CSoutput.t115 gnd 0.061501f
C1374 CSoutput.t131 gnd 0.061501f
C1375 CSoutput.n107 gnd 0.475314f
C1376 CSoutput.n108 gnd 0.237728f
C1377 CSoutput.t160 gnd 0.061501f
C1378 CSoutput.t192 gnd 0.061501f
C1379 CSoutput.n109 gnd 0.475314f
C1380 CSoutput.n110 gnd 0.237728f
C1381 CSoutput.t188 gnd 0.061501f
C1382 CSoutput.t206 gnd 0.061501f
C1383 CSoutput.n111 gnd 0.475314f
C1384 CSoutput.n112 gnd 0.237728f
C1385 CSoutput.t184 gnd 0.061501f
C1386 CSoutput.t172 gnd 0.061501f
C1387 CSoutput.n113 gnd 0.475314f
C1388 CSoutput.n114 gnd 0.237728f
C1389 CSoutput.t150 gnd 0.061501f
C1390 CSoutput.t14 gnd 0.061501f
C1391 CSoutput.n115 gnd 0.475314f
C1392 CSoutput.n116 gnd 0.354512f
C1393 CSoutput.n117 gnd 0.447037f
C1394 CSoutput.t211 gnd 0.061501f
C1395 CSoutput.t119 gnd 0.061501f
C1396 CSoutput.n118 gnd 0.476163f
C1397 CSoutput.t2 gnd 0.061501f
C1398 CSoutput.t210 gnd 0.061501f
C1399 CSoutput.n119 gnd 0.475314f
C1400 CSoutput.n120 gnd 0.482443f
C1401 CSoutput.t155 gnd 0.061501f
C1402 CSoutput.t168 gnd 0.061501f
C1403 CSoutput.n121 gnd 0.475314f
C1404 CSoutput.n122 gnd 0.237728f
C1405 CSoutput.t3 gnd 0.061501f
C1406 CSoutput.t146 gnd 0.061501f
C1407 CSoutput.n123 gnd 0.475314f
C1408 CSoutput.n124 gnd 0.237728f
C1409 CSoutput.t194 gnd 0.061501f
C1410 CSoutput.t170 gnd 0.061501f
C1411 CSoutput.n125 gnd 0.475314f
C1412 CSoutput.n126 gnd 0.237728f
C1413 CSoutput.t124 gnd 0.061501f
C1414 CSoutput.t175 gnd 0.061501f
C1415 CSoutput.n127 gnd 0.475314f
C1416 CSoutput.n128 gnd 0.237728f
C1417 CSoutput.t214 gnd 0.061501f
C1418 CSoutput.t195 gnd 0.061501f
C1419 CSoutput.n129 gnd 0.475314f
C1420 CSoutput.n130 gnd 0.237728f
C1421 CSoutput.t154 gnd 0.061501f
C1422 CSoutput.t116 gnd 0.061501f
C1423 CSoutput.n131 gnd 0.475314f
C1424 CSoutput.n132 gnd 0.237728f
C1425 CSoutput.t169 gnd 0.061501f
C1426 CSoutput.t136 gnd 0.061501f
C1427 CSoutput.n133 gnd 0.475314f
C1428 CSoutput.n134 gnd 0.237728f
C1429 CSoutput.t190 gnd 0.061501f
C1430 CSoutput.t191 gnd 0.061501f
C1431 CSoutput.n135 gnd 0.475314f
C1432 CSoutput.n136 gnd 0.354512f
C1433 CSoutput.n137 gnd 0.499673f
C1434 CSoutput.n138 gnd 9.571919f
C1435 CSoutput.n140 gnd 0.8722f
C1436 CSoutput.n141 gnd 0.65415f
C1437 CSoutput.n142 gnd 0.8722f
C1438 CSoutput.n143 gnd 0.8722f
C1439 CSoutput.n144 gnd 2.34823f
C1440 CSoutput.n145 gnd 0.8722f
C1441 CSoutput.n146 gnd 0.8722f
C1442 CSoutput.t233 gnd 1.09025f
C1443 CSoutput.n147 gnd 0.8722f
C1444 CSoutput.n148 gnd 0.8722f
C1445 CSoutput.n152 gnd 0.8722f
C1446 CSoutput.n156 gnd 0.8722f
C1447 CSoutput.n157 gnd 0.8722f
C1448 CSoutput.n159 gnd 0.8722f
C1449 CSoutput.n164 gnd 0.8722f
C1450 CSoutput.n166 gnd 0.8722f
C1451 CSoutput.n167 gnd 0.8722f
C1452 CSoutput.n169 gnd 0.8722f
C1453 CSoutput.n170 gnd 0.8722f
C1454 CSoutput.n172 gnd 0.8722f
C1455 CSoutput.t219 gnd 14.5744f
C1456 CSoutput.n174 gnd 0.8722f
C1457 CSoutput.n175 gnd 0.65415f
C1458 CSoutput.n176 gnd 0.8722f
C1459 CSoutput.n177 gnd 0.8722f
C1460 CSoutput.n178 gnd 2.34823f
C1461 CSoutput.n179 gnd 0.8722f
C1462 CSoutput.n180 gnd 0.8722f
C1463 CSoutput.t222 gnd 1.09025f
C1464 CSoutput.n181 gnd 0.8722f
C1465 CSoutput.n182 gnd 0.8722f
C1466 CSoutput.n186 gnd 0.8722f
C1467 CSoutput.n190 gnd 0.8722f
C1468 CSoutput.n191 gnd 0.8722f
C1469 CSoutput.n193 gnd 0.8722f
C1470 CSoutput.n198 gnd 0.8722f
C1471 CSoutput.n200 gnd 0.8722f
C1472 CSoutput.n201 gnd 0.8722f
C1473 CSoutput.n203 gnd 0.8722f
C1474 CSoutput.n204 gnd 0.8722f
C1475 CSoutput.n206 gnd 0.8722f
C1476 CSoutput.n207 gnd 0.65415f
C1477 CSoutput.n209 gnd 0.8722f
C1478 CSoutput.n210 gnd 0.65415f
C1479 CSoutput.n211 gnd 0.8722f
C1480 CSoutput.n212 gnd 0.8722f
C1481 CSoutput.n213 gnd 2.34823f
C1482 CSoutput.n214 gnd 0.8722f
C1483 CSoutput.n215 gnd 0.8722f
C1484 CSoutput.t230 gnd 1.09025f
C1485 CSoutput.n216 gnd 0.8722f
C1486 CSoutput.n217 gnd 2.34823f
C1487 CSoutput.n219 gnd 0.8722f
C1488 CSoutput.n220 gnd 0.8722f
C1489 CSoutput.n222 gnd 0.8722f
C1490 CSoutput.n223 gnd 0.8722f
C1491 CSoutput.t235 gnd 14.3368f
C1492 CSoutput.t229 gnd 14.5744f
C1493 CSoutput.n229 gnd 2.73622f
C1494 CSoutput.n230 gnd 11.1464f
C1495 CSoutput.n231 gnd 11.6128f
C1496 CSoutput.n236 gnd 2.96406f
C1497 CSoutput.n242 gnd 0.8722f
C1498 CSoutput.n244 gnd 0.8722f
C1499 CSoutput.n246 gnd 0.8722f
C1500 CSoutput.n248 gnd 0.8722f
C1501 CSoutput.n250 gnd 0.8722f
C1502 CSoutput.n256 gnd 0.8722f
C1503 CSoutput.n263 gnd 1.60015f
C1504 CSoutput.n264 gnd 1.60015f
C1505 CSoutput.n265 gnd 0.8722f
C1506 CSoutput.n266 gnd 0.8722f
C1507 CSoutput.n268 gnd 0.65415f
C1508 CSoutput.n269 gnd 0.560221f
C1509 CSoutput.n271 gnd 0.65415f
C1510 CSoutput.n272 gnd 0.560221f
C1511 CSoutput.n273 gnd 0.65415f
C1512 CSoutput.n275 gnd 0.8722f
C1513 CSoutput.n277 gnd 2.34823f
C1514 CSoutput.n278 gnd 2.73622f
C1515 CSoutput.n279 gnd 10.2518f
C1516 CSoutput.n281 gnd 0.65415f
C1517 CSoutput.n282 gnd 1.68317f
C1518 CSoutput.n283 gnd 0.65415f
C1519 CSoutput.n285 gnd 0.8722f
C1520 CSoutput.n287 gnd 2.34823f
C1521 CSoutput.n288 gnd 5.11428f
C1522 CSoutput.t4 gnd 0.061501f
C1523 CSoutput.t180 gnd 0.061501f
C1524 CSoutput.n289 gnd 0.476163f
C1525 CSoutput.t212 gnd 0.061501f
C1526 CSoutput.t174 gnd 0.061501f
C1527 CSoutput.n290 gnd 0.475314f
C1528 CSoutput.n291 gnd 0.482443f
C1529 CSoutput.t1 gnd 0.061501f
C1530 CSoutput.t133 gnd 0.061501f
C1531 CSoutput.n292 gnd 0.475314f
C1532 CSoutput.n293 gnd 0.237728f
C1533 CSoutput.t134 gnd 0.061501f
C1534 CSoutput.t118 gnd 0.061501f
C1535 CSoutput.n294 gnd 0.475314f
C1536 CSoutput.n295 gnd 0.237728f
C1537 CSoutput.t11 gnd 0.061501f
C1538 CSoutput.t7 gnd 0.061501f
C1539 CSoutput.n296 gnd 0.475314f
C1540 CSoutput.n297 gnd 0.237728f
C1541 CSoutput.t176 gnd 0.061501f
C1542 CSoutput.t164 gnd 0.061501f
C1543 CSoutput.n298 gnd 0.475314f
C1544 CSoutput.n299 gnd 0.237728f
C1545 CSoutput.t196 gnd 0.061501f
C1546 CSoutput.t202 gnd 0.061501f
C1547 CSoutput.n300 gnd 0.475314f
C1548 CSoutput.n301 gnd 0.237728f
C1549 CSoutput.t162 gnd 0.061501f
C1550 CSoutput.t152 gnd 0.061501f
C1551 CSoutput.n302 gnd 0.475314f
C1552 CSoutput.n303 gnd 0.237728f
C1553 CSoutput.t130 gnd 0.061501f
C1554 CSoutput.t141 gnd 0.061501f
C1555 CSoutput.n304 gnd 0.475314f
C1556 CSoutput.n305 gnd 0.237728f
C1557 CSoutput.t10 gnd 0.061501f
C1558 CSoutput.t9 gnd 0.061501f
C1559 CSoutput.n306 gnd 0.475314f
C1560 CSoutput.n307 gnd 0.435938f
C1561 CSoutput.t179 gnd 0.061501f
C1562 CSoutput.t161 gnd 0.061501f
C1563 CSoutput.n308 gnd 0.476163f
C1564 CSoutput.t166 gnd 0.061501f
C1565 CSoutput.t156 gnd 0.061501f
C1566 CSoutput.n309 gnd 0.475314f
C1567 CSoutput.n310 gnd 0.482443f
C1568 CSoutput.t213 gnd 0.061501f
C1569 CSoutput.t204 gnd 0.061501f
C1570 CSoutput.n311 gnd 0.475314f
C1571 CSoutput.n312 gnd 0.237728f
C1572 CSoutput.t5 gnd 0.061501f
C1573 CSoutput.t177 gnd 0.061501f
C1574 CSoutput.n313 gnd 0.475314f
C1575 CSoutput.n314 gnd 0.237728f
C1576 CSoutput.t137 gnd 0.061501f
C1577 CSoutput.t114 gnd 0.061501f
C1578 CSoutput.n315 gnd 0.475314f
C1579 CSoutput.n316 gnd 0.237728f
C1580 CSoutput.t12 gnd 0.061501f
C1581 CSoutput.t201 gnd 0.061501f
C1582 CSoutput.n317 gnd 0.475314f
C1583 CSoutput.n318 gnd 0.237728f
C1584 CSoutput.t181 gnd 0.061501f
C1585 CSoutput.t153 gnd 0.061501f
C1586 CSoutput.n319 gnd 0.475314f
C1587 CSoutput.n320 gnd 0.237728f
C1588 CSoutput.t178 gnd 0.061501f
C1589 CSoutput.t167 gnd 0.061501f
C1590 CSoutput.n321 gnd 0.475314f
C1591 CSoutput.n322 gnd 0.237728f
C1592 CSoutput.t186 gnd 0.061501f
C1593 CSoutput.t158 gnd 0.061501f
C1594 CSoutput.n323 gnd 0.475314f
C1595 CSoutput.n324 gnd 0.237728f
C1596 CSoutput.t205 gnd 0.061501f
C1597 CSoutput.t183 gnd 0.061501f
C1598 CSoutput.n325 gnd 0.475314f
C1599 CSoutput.n326 gnd 0.354512f
C1600 CSoutput.n327 gnd 0.447037f
C1601 CSoutput.t129 gnd 0.061501f
C1602 CSoutput.t163 gnd 0.061501f
C1603 CSoutput.n328 gnd 0.476163f
C1604 CSoutput.t187 gnd 0.061501f
C1605 CSoutput.t159 gnd 0.061501f
C1606 CSoutput.n329 gnd 0.475314f
C1607 CSoutput.n330 gnd 0.482443f
C1608 CSoutput.t16 gnd 0.061501f
C1609 CSoutput.t132 gnd 0.061501f
C1610 CSoutput.n331 gnd 0.475314f
C1611 CSoutput.n332 gnd 0.237728f
C1612 CSoutput.t209 gnd 0.061501f
C1613 CSoutput.t126 gnd 0.061501f
C1614 CSoutput.n333 gnd 0.475314f
C1615 CSoutput.n334 gnd 0.237728f
C1616 CSoutput.t120 gnd 0.061501f
C1617 CSoutput.t203 gnd 0.061501f
C1618 CSoutput.n335 gnd 0.475314f
C1619 CSoutput.n336 gnd 0.237728f
C1620 CSoutput.t135 gnd 0.061501f
C1621 CSoutput.t182 gnd 0.061501f
C1622 CSoutput.n337 gnd 0.475314f
C1623 CSoutput.n338 gnd 0.237728f
C1624 CSoutput.t125 gnd 0.061501f
C1625 CSoutput.t193 gnd 0.061501f
C1626 CSoutput.n339 gnd 0.475314f
C1627 CSoutput.n340 gnd 0.237728f
C1628 CSoutput.t128 gnd 0.061501f
C1629 CSoutput.t148 gnd 0.061501f
C1630 CSoutput.n341 gnd 0.475314f
C1631 CSoutput.n342 gnd 0.237728f
C1632 CSoutput.t139 gnd 0.061501f
C1633 CSoutput.t17 gnd 0.061501f
C1634 CSoutput.n343 gnd 0.475314f
C1635 CSoutput.n344 gnd 0.237728f
C1636 CSoutput.t185 gnd 0.061501f
C1637 CSoutput.t123 gnd 0.061501f
C1638 CSoutput.n345 gnd 0.475312f
C1639 CSoutput.n346 gnd 0.354513f
C1640 CSoutput.n347 gnd 0.499673f
C1641 CSoutput.n348 gnd 13.627701f
C1642 CSoutput.t57 gnd 0.053814f
C1643 CSoutput.t110 gnd 0.053814f
C1644 CSoutput.n349 gnd 0.477107f
C1645 CSoutput.t51 gnd 0.053814f
C1646 CSoutput.t56 gnd 0.053814f
C1647 CSoutput.n350 gnd 0.475516f
C1648 CSoutput.n351 gnd 0.443092f
C1649 CSoutput.t41 gnd 0.053814f
C1650 CSoutput.t60 gnd 0.053814f
C1651 CSoutput.n352 gnd 0.475516f
C1652 CSoutput.n353 gnd 0.218423f
C1653 CSoutput.t75 gnd 0.053814f
C1654 CSoutput.t52 gnd 0.053814f
C1655 CSoutput.n354 gnd 0.475516f
C1656 CSoutput.n355 gnd 0.218423f
C1657 CSoutput.t59 gnd 0.053814f
C1658 CSoutput.t101 gnd 0.053814f
C1659 CSoutput.n356 gnd 0.475516f
C1660 CSoutput.n357 gnd 0.218423f
C1661 CSoutput.t71 gnd 0.053814f
C1662 CSoutput.t81 gnd 0.053814f
C1663 CSoutput.n358 gnd 0.475516f
C1664 CSoutput.n359 gnd 0.218423f
C1665 CSoutput.t36 gnd 0.053814f
C1666 CSoutput.t61 gnd 0.053814f
C1667 CSoutput.n360 gnd 0.475516f
C1668 CSoutput.n361 gnd 0.218423f
C1669 CSoutput.t25 gnd 0.053814f
C1670 CSoutput.t48 gnd 0.053814f
C1671 CSoutput.n362 gnd 0.475516f
C1672 CSoutput.n363 gnd 0.40287f
C1673 CSoutput.t106 gnd 0.053814f
C1674 CSoutput.t18 gnd 0.053814f
C1675 CSoutput.n364 gnd 0.477107f
C1676 CSoutput.t29 gnd 0.053814f
C1677 CSoutput.t99 gnd 0.053814f
C1678 CSoutput.n365 gnd 0.475516f
C1679 CSoutput.n366 gnd 0.443092f
C1680 CSoutput.t20 gnd 0.053814f
C1681 CSoutput.t92 gnd 0.053814f
C1682 CSoutput.n367 gnd 0.475516f
C1683 CSoutput.n368 gnd 0.218423f
C1684 CSoutput.t100 gnd 0.053814f
C1685 CSoutput.t19 gnd 0.053814f
C1686 CSoutput.n369 gnd 0.475516f
C1687 CSoutput.n370 gnd 0.218423f
C1688 CSoutput.t83 gnd 0.053814f
C1689 CSoutput.t64 gnd 0.053814f
C1690 CSoutput.n371 gnd 0.475516f
C1691 CSoutput.n372 gnd 0.218423f
C1692 CSoutput.t21 gnd 0.053814f
C1693 CSoutput.t85 gnd 0.053814f
C1694 CSoutput.n373 gnd 0.475516f
C1695 CSoutput.n374 gnd 0.218423f
C1696 CSoutput.t66 gnd 0.053814f
C1697 CSoutput.t72 gnd 0.053814f
C1698 CSoutput.n375 gnd 0.475516f
C1699 CSoutput.n376 gnd 0.218423f
C1700 CSoutput.t84 gnd 0.053814f
C1701 CSoutput.t65 gnd 0.053814f
C1702 CSoutput.n377 gnd 0.475516f
C1703 CSoutput.n378 gnd 0.331614f
C1704 CSoutput.n379 gnd 0.418268f
C1705 CSoutput.t30 gnd 0.053814f
C1706 CSoutput.t102 gnd 0.053814f
C1707 CSoutput.n380 gnd 0.477107f
C1708 CSoutput.t49 gnd 0.053814f
C1709 CSoutput.t53 gnd 0.053814f
C1710 CSoutput.n381 gnd 0.475516f
C1711 CSoutput.n382 gnd 0.443092f
C1712 CSoutput.t22 gnd 0.053814f
C1713 CSoutput.t87 gnd 0.053814f
C1714 CSoutput.n383 gnd 0.475516f
C1715 CSoutput.n384 gnd 0.218423f
C1716 CSoutput.t58 gnd 0.053814f
C1717 CSoutput.t31 gnd 0.053814f
C1718 CSoutput.n385 gnd 0.475516f
C1719 CSoutput.n386 gnd 0.218423f
C1720 CSoutput.t39 gnd 0.053814f
C1721 CSoutput.t113 gnd 0.053814f
C1722 CSoutput.n387 gnd 0.475516f
C1723 CSoutput.n388 gnd 0.218423f
C1724 CSoutput.t40 gnd 0.053814f
C1725 CSoutput.t44 gnd 0.053814f
C1726 CSoutput.n389 gnd 0.475516f
C1727 CSoutput.n390 gnd 0.218423f
C1728 CSoutput.t28 gnd 0.053814f
C1729 CSoutput.t98 gnd 0.053814f
C1730 CSoutput.n391 gnd 0.475516f
C1731 CSoutput.n392 gnd 0.218423f
C1732 CSoutput.t47 gnd 0.053814f
C1733 CSoutput.t37 gnd 0.053814f
C1734 CSoutput.n393 gnd 0.475516f
C1735 CSoutput.n394 gnd 0.331614f
C1736 CSoutput.n395 gnd 0.449154f
C1737 CSoutput.n396 gnd 13.4951f
C1738 CSoutput.t43 gnd 0.053814f
C1739 CSoutput.t86 gnd 0.053814f
C1740 CSoutput.n397 gnd 0.477107f
C1741 CSoutput.t82 gnd 0.053814f
C1742 CSoutput.t63 gnd 0.053814f
C1743 CSoutput.n398 gnd 0.475516f
C1744 CSoutput.n399 gnd 0.443092f
C1745 CSoutput.t89 gnd 0.053814f
C1746 CSoutput.t54 gnd 0.053814f
C1747 CSoutput.n400 gnd 0.475516f
C1748 CSoutput.n401 gnd 0.218423f
C1749 CSoutput.t73 gnd 0.053814f
C1750 CSoutput.t104 gnd 0.053814f
C1751 CSoutput.n402 gnd 0.475516f
C1752 CSoutput.n403 gnd 0.218423f
C1753 CSoutput.t38 gnd 0.053814f
C1754 CSoutput.t88 gnd 0.053814f
C1755 CSoutput.n404 gnd 0.475516f
C1756 CSoutput.n405 gnd 0.218423f
C1757 CSoutput.t27 gnd 0.053814f
C1758 CSoutput.t94 gnd 0.053814f
C1759 CSoutput.n406 gnd 0.475516f
C1760 CSoutput.n407 gnd 0.218423f
C1761 CSoutput.t93 gnd 0.053814f
C1762 CSoutput.t50 gnd 0.053814f
C1763 CSoutput.n408 gnd 0.475516f
C1764 CSoutput.n409 gnd 0.218423f
C1765 CSoutput.t69 gnd 0.053814f
C1766 CSoutput.t46 gnd 0.053814f
C1767 CSoutput.n410 gnd 0.475516f
C1768 CSoutput.n411 gnd 0.40287f
C1769 CSoutput.t33 gnd 0.053814f
C1770 CSoutput.t26 gnd 0.053814f
C1771 CSoutput.n412 gnd 0.477107f
C1772 CSoutput.t23 gnd 0.053814f
C1773 CSoutput.t111 gnd 0.053814f
C1774 CSoutput.n413 gnd 0.475516f
C1775 CSoutput.n414 gnd 0.443092f
C1776 CSoutput.t112 gnd 0.053814f
C1777 CSoutput.t34 gnd 0.053814f
C1778 CSoutput.n415 gnd 0.475516f
C1779 CSoutput.n416 gnd 0.218423f
C1780 CSoutput.t35 gnd 0.053814f
C1781 CSoutput.t77 gnd 0.053814f
C1782 CSoutput.n417 gnd 0.475516f
C1783 CSoutput.n418 gnd 0.218423f
C1784 CSoutput.t78 gnd 0.053814f
C1785 CSoutput.t105 gnd 0.053814f
C1786 CSoutput.n419 gnd 0.475516f
C1787 CSoutput.n420 gnd 0.218423f
C1788 CSoutput.t108 gnd 0.053814f
C1789 CSoutput.t97 gnd 0.053814f
C1790 CSoutput.n421 gnd 0.475516f
C1791 CSoutput.n422 gnd 0.218423f
C1792 CSoutput.t91 gnd 0.053814f
C1793 CSoutput.t79 gnd 0.053814f
C1794 CSoutput.n423 gnd 0.475516f
C1795 CSoutput.n424 gnd 0.218423f
C1796 CSoutput.t80 gnd 0.053814f
C1797 CSoutput.t109 gnd 0.053814f
C1798 CSoutput.n425 gnd 0.475516f
C1799 CSoutput.n426 gnd 0.331614f
C1800 CSoutput.n427 gnd 0.418268f
C1801 CSoutput.t70 gnd 0.053814f
C1802 CSoutput.t95 gnd 0.053814f
C1803 CSoutput.n428 gnd 0.477107f
C1804 CSoutput.t42 gnd 0.053814f
C1805 CSoutput.t55 gnd 0.053814f
C1806 CSoutput.n429 gnd 0.475516f
C1807 CSoutput.n430 gnd 0.443092f
C1808 CSoutput.t62 gnd 0.053814f
C1809 CSoutput.t76 gnd 0.053814f
C1810 CSoutput.n431 gnd 0.475516f
C1811 CSoutput.n432 gnd 0.218423f
C1812 CSoutput.t96 gnd 0.053814f
C1813 CSoutput.t67 gnd 0.053814f
C1814 CSoutput.n433 gnd 0.475516f
C1815 CSoutput.n434 gnd 0.218423f
C1816 CSoutput.t74 gnd 0.053814f
C1817 CSoutput.t107 gnd 0.053814f
C1818 CSoutput.n435 gnd 0.475516f
C1819 CSoutput.n436 gnd 0.218423f
C1820 CSoutput.t24 gnd 0.053814f
C1821 CSoutput.t45 gnd 0.053814f
C1822 CSoutput.n437 gnd 0.475516f
C1823 CSoutput.n438 gnd 0.218423f
C1824 CSoutput.t68 gnd 0.053814f
C1825 CSoutput.t90 gnd 0.053814f
C1826 CSoutput.n439 gnd 0.475516f
C1827 CSoutput.n440 gnd 0.218423f
C1828 CSoutput.t103 gnd 0.053814f
C1829 CSoutput.t32 gnd 0.053814f
C1830 CSoutput.n441 gnd 0.475516f
C1831 CSoutput.n442 gnd 0.331614f
C1832 CSoutput.n443 gnd 0.449154f
C1833 CSoutput.n444 gnd 8.00328f
C1834 CSoutput.n445 gnd 14.821199f
C1835 commonsourceibias.n0 gnd 0.012609f
C1836 commonsourceibias.t120 gnd 0.190924f
C1837 commonsourceibias.t67 gnd 0.176537f
C1838 commonsourceibias.n1 gnd 0.00768f
C1839 commonsourceibias.n2 gnd 0.009449f
C1840 commonsourceibias.t126 gnd 0.176537f
C1841 commonsourceibias.n3 gnd 0.009585f
C1842 commonsourceibias.n4 gnd 0.009449f
C1843 commonsourceibias.t121 gnd 0.176537f
C1844 commonsourceibias.n5 gnd 0.070438f
C1845 commonsourceibias.t136 gnd 0.176537f
C1846 commonsourceibias.n6 gnd 0.007644f
C1847 commonsourceibias.n7 gnd 0.009449f
C1848 commonsourceibias.t117 gnd 0.176537f
C1849 commonsourceibias.n8 gnd 0.009122f
C1850 commonsourceibias.n9 gnd 0.009449f
C1851 commonsourceibias.t102 gnd 0.176537f
C1852 commonsourceibias.n10 gnd 0.070438f
C1853 commonsourceibias.t125 gnd 0.176537f
C1854 commonsourceibias.n11 gnd 0.007632f
C1855 commonsourceibias.n12 gnd 0.012609f
C1856 commonsourceibias.t20 gnd 0.190924f
C1857 commonsourceibias.t14 gnd 0.176537f
C1858 commonsourceibias.n13 gnd 0.00768f
C1859 commonsourceibias.n14 gnd 0.009449f
C1860 commonsourceibias.t58 gnd 0.176537f
C1861 commonsourceibias.n15 gnd 0.009585f
C1862 commonsourceibias.n16 gnd 0.009449f
C1863 commonsourceibias.t18 gnd 0.176537f
C1864 commonsourceibias.n17 gnd 0.070438f
C1865 commonsourceibias.t60 gnd 0.176537f
C1866 commonsourceibias.n18 gnd 0.007644f
C1867 commonsourceibias.n19 gnd 0.009449f
C1868 commonsourceibias.t24 gnd 0.176537f
C1869 commonsourceibias.n20 gnd 0.009122f
C1870 commonsourceibias.n21 gnd 0.009449f
C1871 commonsourceibias.t12 gnd 0.176537f
C1872 commonsourceibias.n22 gnd 0.070438f
C1873 commonsourceibias.t54 gnd 0.176537f
C1874 commonsourceibias.n23 gnd 0.007632f
C1875 commonsourceibias.n24 gnd 0.009449f
C1876 commonsourceibias.t22 gnd 0.176537f
C1877 commonsourceibias.t38 gnd 0.176537f
C1878 commonsourceibias.n25 gnd 0.070438f
C1879 commonsourceibias.n26 gnd 0.009449f
C1880 commonsourceibias.t8 gnd 0.176537f
C1881 commonsourceibias.n27 gnd 0.070438f
C1882 commonsourceibias.n28 gnd 0.009449f
C1883 commonsourceibias.t46 gnd 0.176537f
C1884 commonsourceibias.n29 gnd 0.070438f
C1885 commonsourceibias.n30 gnd 0.009449f
C1886 commonsourceibias.t62 gnd 0.176537f
C1887 commonsourceibias.n31 gnd 0.010741f
C1888 commonsourceibias.n32 gnd 0.009449f
C1889 commonsourceibias.t42 gnd 0.176537f
C1890 commonsourceibias.n33 gnd 0.012701f
C1891 commonsourceibias.t56 gnd 0.196658f
C1892 commonsourceibias.t16 gnd 0.176537f
C1893 commonsourceibias.n34 gnd 0.078486f
C1894 commonsourceibias.n35 gnd 0.084086f
C1895 commonsourceibias.n36 gnd 0.04022f
C1896 commonsourceibias.n37 gnd 0.009449f
C1897 commonsourceibias.n38 gnd 0.00768f
C1898 commonsourceibias.n39 gnd 0.013021f
C1899 commonsourceibias.n40 gnd 0.070438f
C1900 commonsourceibias.n41 gnd 0.013076f
C1901 commonsourceibias.n42 gnd 0.009449f
C1902 commonsourceibias.n43 gnd 0.009449f
C1903 commonsourceibias.n44 gnd 0.009449f
C1904 commonsourceibias.n45 gnd 0.009585f
C1905 commonsourceibias.n46 gnd 0.070438f
C1906 commonsourceibias.n47 gnd 0.011646f
C1907 commonsourceibias.n48 gnd 0.012884f
C1908 commonsourceibias.n49 gnd 0.009449f
C1909 commonsourceibias.n50 gnd 0.009449f
C1910 commonsourceibias.n51 gnd 0.0128f
C1911 commonsourceibias.n52 gnd 0.007644f
C1912 commonsourceibias.n53 gnd 0.012959f
C1913 commonsourceibias.n54 gnd 0.009449f
C1914 commonsourceibias.n55 gnd 0.009449f
C1915 commonsourceibias.n56 gnd 0.013038f
C1916 commonsourceibias.n57 gnd 0.011242f
C1917 commonsourceibias.n58 gnd 0.009122f
C1918 commonsourceibias.n59 gnd 0.009449f
C1919 commonsourceibias.n60 gnd 0.009449f
C1920 commonsourceibias.n61 gnd 0.011558f
C1921 commonsourceibias.n62 gnd 0.012972f
C1922 commonsourceibias.n63 gnd 0.070438f
C1923 commonsourceibias.n64 gnd 0.012885f
C1924 commonsourceibias.n65 gnd 0.009449f
C1925 commonsourceibias.n66 gnd 0.009449f
C1926 commonsourceibias.n67 gnd 0.009449f
C1927 commonsourceibias.n68 gnd 0.012885f
C1928 commonsourceibias.n69 gnd 0.070438f
C1929 commonsourceibias.n70 gnd 0.012972f
C1930 commonsourceibias.n71 gnd 0.011558f
C1931 commonsourceibias.n72 gnd 0.009449f
C1932 commonsourceibias.n73 gnd 0.009449f
C1933 commonsourceibias.n74 gnd 0.009449f
C1934 commonsourceibias.n75 gnd 0.011242f
C1935 commonsourceibias.n76 gnd 0.013038f
C1936 commonsourceibias.n77 gnd 0.070438f
C1937 commonsourceibias.n78 gnd 0.012959f
C1938 commonsourceibias.n79 gnd 0.009449f
C1939 commonsourceibias.n80 gnd 0.009449f
C1940 commonsourceibias.n81 gnd 0.009449f
C1941 commonsourceibias.n82 gnd 0.0128f
C1942 commonsourceibias.n83 gnd 0.070438f
C1943 commonsourceibias.n84 gnd 0.012884f
C1944 commonsourceibias.n85 gnd 0.011646f
C1945 commonsourceibias.n86 gnd 0.009449f
C1946 commonsourceibias.n87 gnd 0.009449f
C1947 commonsourceibias.n88 gnd 0.009449f
C1948 commonsourceibias.n89 gnd 0.010741f
C1949 commonsourceibias.n90 gnd 0.013076f
C1950 commonsourceibias.n91 gnd 0.070438f
C1951 commonsourceibias.n92 gnd 0.013021f
C1952 commonsourceibias.n93 gnd 0.009449f
C1953 commonsourceibias.n94 gnd 0.009449f
C1954 commonsourceibias.n95 gnd 0.009449f
C1955 commonsourceibias.n96 gnd 0.012701f
C1956 commonsourceibias.n97 gnd 0.070438f
C1957 commonsourceibias.n98 gnd 0.012732f
C1958 commonsourceibias.n99 gnd 0.084938f
C1959 commonsourceibias.n100 gnd 0.094974f
C1960 commonsourceibias.t21 gnd 0.02039f
C1961 commonsourceibias.t15 gnd 0.02039f
C1962 commonsourceibias.n101 gnd 0.180173f
C1963 commonsourceibias.n102 gnd 0.156069f
C1964 commonsourceibias.t59 gnd 0.02039f
C1965 commonsourceibias.t19 gnd 0.02039f
C1966 commonsourceibias.n103 gnd 0.180173f
C1967 commonsourceibias.n104 gnd 0.082761f
C1968 commonsourceibias.t61 gnd 0.02039f
C1969 commonsourceibias.t25 gnd 0.02039f
C1970 commonsourceibias.n105 gnd 0.180173f
C1971 commonsourceibias.n106 gnd 0.082761f
C1972 commonsourceibias.t13 gnd 0.02039f
C1973 commonsourceibias.t55 gnd 0.02039f
C1974 commonsourceibias.n107 gnd 0.180173f
C1975 commonsourceibias.n108 gnd 0.069143f
C1976 commonsourceibias.t17 gnd 0.02039f
C1977 commonsourceibias.t57 gnd 0.02039f
C1978 commonsourceibias.n109 gnd 0.180776f
C1979 commonsourceibias.t63 gnd 0.02039f
C1980 commonsourceibias.t43 gnd 0.02039f
C1981 commonsourceibias.n110 gnd 0.180173f
C1982 commonsourceibias.n111 gnd 0.167888f
C1983 commonsourceibias.t9 gnd 0.02039f
C1984 commonsourceibias.t47 gnd 0.02039f
C1985 commonsourceibias.n112 gnd 0.180173f
C1986 commonsourceibias.n113 gnd 0.082761f
C1987 commonsourceibias.t23 gnd 0.02039f
C1988 commonsourceibias.t39 gnd 0.02039f
C1989 commonsourceibias.n114 gnd 0.180173f
C1990 commonsourceibias.n115 gnd 0.069143f
C1991 commonsourceibias.n116 gnd 0.083724f
C1992 commonsourceibias.n117 gnd 0.009449f
C1993 commonsourceibias.t118 gnd 0.176537f
C1994 commonsourceibias.t76 gnd 0.176537f
C1995 commonsourceibias.n118 gnd 0.070438f
C1996 commonsourceibias.n119 gnd 0.009449f
C1997 commonsourceibias.t106 gnd 0.176537f
C1998 commonsourceibias.n120 gnd 0.070438f
C1999 commonsourceibias.n121 gnd 0.009449f
C2000 commonsourceibias.t96 gnd 0.176537f
C2001 commonsourceibias.n122 gnd 0.070438f
C2002 commonsourceibias.n123 gnd 0.009449f
C2003 commonsourceibias.t141 gnd 0.176537f
C2004 commonsourceibias.n124 gnd 0.010741f
C2005 commonsourceibias.n125 gnd 0.009449f
C2006 commonsourceibias.t116 gnd 0.176537f
C2007 commonsourceibias.n126 gnd 0.012701f
C2008 commonsourceibias.t129 gnd 0.196658f
C2009 commonsourceibias.t152 gnd 0.176537f
C2010 commonsourceibias.n127 gnd 0.078486f
C2011 commonsourceibias.n128 gnd 0.084086f
C2012 commonsourceibias.n129 gnd 0.04022f
C2013 commonsourceibias.n130 gnd 0.009449f
C2014 commonsourceibias.n131 gnd 0.00768f
C2015 commonsourceibias.n132 gnd 0.013021f
C2016 commonsourceibias.n133 gnd 0.070438f
C2017 commonsourceibias.n134 gnd 0.013076f
C2018 commonsourceibias.n135 gnd 0.009449f
C2019 commonsourceibias.n136 gnd 0.009449f
C2020 commonsourceibias.n137 gnd 0.009449f
C2021 commonsourceibias.n138 gnd 0.009585f
C2022 commonsourceibias.n139 gnd 0.070438f
C2023 commonsourceibias.n140 gnd 0.011646f
C2024 commonsourceibias.n141 gnd 0.012884f
C2025 commonsourceibias.n142 gnd 0.009449f
C2026 commonsourceibias.n143 gnd 0.009449f
C2027 commonsourceibias.n144 gnd 0.0128f
C2028 commonsourceibias.n145 gnd 0.007644f
C2029 commonsourceibias.n146 gnd 0.012959f
C2030 commonsourceibias.n147 gnd 0.009449f
C2031 commonsourceibias.n148 gnd 0.009449f
C2032 commonsourceibias.n149 gnd 0.013038f
C2033 commonsourceibias.n150 gnd 0.011242f
C2034 commonsourceibias.n151 gnd 0.009122f
C2035 commonsourceibias.n152 gnd 0.009449f
C2036 commonsourceibias.n153 gnd 0.009449f
C2037 commonsourceibias.n154 gnd 0.011558f
C2038 commonsourceibias.n155 gnd 0.012972f
C2039 commonsourceibias.n156 gnd 0.070438f
C2040 commonsourceibias.n157 gnd 0.012885f
C2041 commonsourceibias.n158 gnd 0.009404f
C2042 commonsourceibias.n159 gnd 0.068305f
C2043 commonsourceibias.n160 gnd 0.009404f
C2044 commonsourceibias.n161 gnd 0.012885f
C2045 commonsourceibias.n162 gnd 0.070438f
C2046 commonsourceibias.n163 gnd 0.012972f
C2047 commonsourceibias.n164 gnd 0.011558f
C2048 commonsourceibias.n165 gnd 0.009449f
C2049 commonsourceibias.n166 gnd 0.009449f
C2050 commonsourceibias.n167 gnd 0.009449f
C2051 commonsourceibias.n168 gnd 0.011242f
C2052 commonsourceibias.n169 gnd 0.013038f
C2053 commonsourceibias.n170 gnd 0.070438f
C2054 commonsourceibias.n171 gnd 0.012959f
C2055 commonsourceibias.n172 gnd 0.009449f
C2056 commonsourceibias.n173 gnd 0.009449f
C2057 commonsourceibias.n174 gnd 0.009449f
C2058 commonsourceibias.n175 gnd 0.0128f
C2059 commonsourceibias.n176 gnd 0.070438f
C2060 commonsourceibias.n177 gnd 0.012884f
C2061 commonsourceibias.n178 gnd 0.011646f
C2062 commonsourceibias.n179 gnd 0.009449f
C2063 commonsourceibias.n180 gnd 0.009449f
C2064 commonsourceibias.n181 gnd 0.009449f
C2065 commonsourceibias.n182 gnd 0.010741f
C2066 commonsourceibias.n183 gnd 0.013076f
C2067 commonsourceibias.n184 gnd 0.070438f
C2068 commonsourceibias.n185 gnd 0.013021f
C2069 commonsourceibias.n186 gnd 0.009449f
C2070 commonsourceibias.n187 gnd 0.009449f
C2071 commonsourceibias.n188 gnd 0.009449f
C2072 commonsourceibias.n189 gnd 0.012701f
C2073 commonsourceibias.n190 gnd 0.070438f
C2074 commonsourceibias.n191 gnd 0.012732f
C2075 commonsourceibias.n192 gnd 0.084938f
C2076 commonsourceibias.n193 gnd 0.056112f
C2077 commonsourceibias.n194 gnd 0.012609f
C2078 commonsourceibias.t71 gnd 0.190924f
C2079 commonsourceibias.t159 gnd 0.176537f
C2080 commonsourceibias.n195 gnd 0.00768f
C2081 commonsourceibias.n196 gnd 0.009449f
C2082 commonsourceibias.t148 gnd 0.176537f
C2083 commonsourceibias.n197 gnd 0.009585f
C2084 commonsourceibias.n198 gnd 0.009449f
C2085 commonsourceibias.t78 gnd 0.176537f
C2086 commonsourceibias.n199 gnd 0.070438f
C2087 commonsourceibias.t157 gnd 0.176537f
C2088 commonsourceibias.n200 gnd 0.007644f
C2089 commonsourceibias.n201 gnd 0.009449f
C2090 commonsourceibias.t85 gnd 0.176537f
C2091 commonsourceibias.n202 gnd 0.009122f
C2092 commonsourceibias.n203 gnd 0.009449f
C2093 commonsourceibias.t77 gnd 0.176537f
C2094 commonsourceibias.n204 gnd 0.070438f
C2095 commonsourceibias.t158 gnd 0.176537f
C2096 commonsourceibias.n205 gnd 0.007632f
C2097 commonsourceibias.n206 gnd 0.009449f
C2098 commonsourceibias.t94 gnd 0.176537f
C2099 commonsourceibias.t113 gnd 0.176537f
C2100 commonsourceibias.n207 gnd 0.070438f
C2101 commonsourceibias.n208 gnd 0.009449f
C2102 commonsourceibias.t156 gnd 0.176537f
C2103 commonsourceibias.n209 gnd 0.070438f
C2104 commonsourceibias.n210 gnd 0.009449f
C2105 commonsourceibias.t92 gnd 0.176537f
C2106 commonsourceibias.n211 gnd 0.070438f
C2107 commonsourceibias.n212 gnd 0.009449f
C2108 commonsourceibias.t111 gnd 0.176537f
C2109 commonsourceibias.n213 gnd 0.010741f
C2110 commonsourceibias.n214 gnd 0.009449f
C2111 commonsourceibias.t105 gnd 0.176537f
C2112 commonsourceibias.n215 gnd 0.012701f
C2113 commonsourceibias.t112 gnd 0.196658f
C2114 commonsourceibias.t93 gnd 0.176537f
C2115 commonsourceibias.n216 gnd 0.078486f
C2116 commonsourceibias.n217 gnd 0.084086f
C2117 commonsourceibias.n218 gnd 0.04022f
C2118 commonsourceibias.n219 gnd 0.009449f
C2119 commonsourceibias.n220 gnd 0.00768f
C2120 commonsourceibias.n221 gnd 0.013021f
C2121 commonsourceibias.n222 gnd 0.070438f
C2122 commonsourceibias.n223 gnd 0.013076f
C2123 commonsourceibias.n224 gnd 0.009449f
C2124 commonsourceibias.n225 gnd 0.009449f
C2125 commonsourceibias.n226 gnd 0.009449f
C2126 commonsourceibias.n227 gnd 0.009585f
C2127 commonsourceibias.n228 gnd 0.070438f
C2128 commonsourceibias.n229 gnd 0.011646f
C2129 commonsourceibias.n230 gnd 0.012884f
C2130 commonsourceibias.n231 gnd 0.009449f
C2131 commonsourceibias.n232 gnd 0.009449f
C2132 commonsourceibias.n233 gnd 0.0128f
C2133 commonsourceibias.n234 gnd 0.007644f
C2134 commonsourceibias.n235 gnd 0.012959f
C2135 commonsourceibias.n236 gnd 0.009449f
C2136 commonsourceibias.n237 gnd 0.009449f
C2137 commonsourceibias.n238 gnd 0.013038f
C2138 commonsourceibias.n239 gnd 0.011242f
C2139 commonsourceibias.n240 gnd 0.009122f
C2140 commonsourceibias.n241 gnd 0.009449f
C2141 commonsourceibias.n242 gnd 0.009449f
C2142 commonsourceibias.n243 gnd 0.011558f
C2143 commonsourceibias.n244 gnd 0.012972f
C2144 commonsourceibias.n245 gnd 0.070438f
C2145 commonsourceibias.n246 gnd 0.012885f
C2146 commonsourceibias.n247 gnd 0.009449f
C2147 commonsourceibias.n248 gnd 0.009449f
C2148 commonsourceibias.n249 gnd 0.009449f
C2149 commonsourceibias.n250 gnd 0.012885f
C2150 commonsourceibias.n251 gnd 0.070438f
C2151 commonsourceibias.n252 gnd 0.012972f
C2152 commonsourceibias.n253 gnd 0.011558f
C2153 commonsourceibias.n254 gnd 0.009449f
C2154 commonsourceibias.n255 gnd 0.009449f
C2155 commonsourceibias.n256 gnd 0.009449f
C2156 commonsourceibias.n257 gnd 0.011242f
C2157 commonsourceibias.n258 gnd 0.013038f
C2158 commonsourceibias.n259 gnd 0.070438f
C2159 commonsourceibias.n260 gnd 0.012959f
C2160 commonsourceibias.n261 gnd 0.009449f
C2161 commonsourceibias.n262 gnd 0.009449f
C2162 commonsourceibias.n263 gnd 0.009449f
C2163 commonsourceibias.n264 gnd 0.0128f
C2164 commonsourceibias.n265 gnd 0.070438f
C2165 commonsourceibias.n266 gnd 0.012884f
C2166 commonsourceibias.n267 gnd 0.011646f
C2167 commonsourceibias.n268 gnd 0.009449f
C2168 commonsourceibias.n269 gnd 0.009449f
C2169 commonsourceibias.n270 gnd 0.009449f
C2170 commonsourceibias.n271 gnd 0.010741f
C2171 commonsourceibias.n272 gnd 0.013076f
C2172 commonsourceibias.n273 gnd 0.070438f
C2173 commonsourceibias.n274 gnd 0.013021f
C2174 commonsourceibias.n275 gnd 0.009449f
C2175 commonsourceibias.n276 gnd 0.009449f
C2176 commonsourceibias.n277 gnd 0.009449f
C2177 commonsourceibias.n278 gnd 0.012701f
C2178 commonsourceibias.n279 gnd 0.070438f
C2179 commonsourceibias.n280 gnd 0.012732f
C2180 commonsourceibias.n281 gnd 0.084938f
C2181 commonsourceibias.n282 gnd 0.03031f
C2182 commonsourceibias.n283 gnd 0.151321f
C2183 commonsourceibias.n284 gnd 0.012609f
C2184 commonsourceibias.t75 gnd 0.176537f
C2185 commonsourceibias.n285 gnd 0.00768f
C2186 commonsourceibias.n286 gnd 0.009449f
C2187 commonsourceibias.t128 gnd 0.176537f
C2188 commonsourceibias.n287 gnd 0.009585f
C2189 commonsourceibias.n288 gnd 0.009449f
C2190 commonsourceibias.t124 gnd 0.176537f
C2191 commonsourceibias.n289 gnd 0.070438f
C2192 commonsourceibias.t155 gnd 0.176537f
C2193 commonsourceibias.n290 gnd 0.007644f
C2194 commonsourceibias.n291 gnd 0.009449f
C2195 commonsourceibias.t90 gnd 0.176537f
C2196 commonsourceibias.n292 gnd 0.009122f
C2197 commonsourceibias.n293 gnd 0.009449f
C2198 commonsourceibias.t119 gnd 0.176537f
C2199 commonsourceibias.n294 gnd 0.070438f
C2200 commonsourceibias.t146 gnd 0.176537f
C2201 commonsourceibias.n295 gnd 0.007632f
C2202 commonsourceibias.n296 gnd 0.009449f
C2203 commonsourceibias.t138 gnd 0.176537f
C2204 commonsourceibias.t64 gnd 0.176537f
C2205 commonsourceibias.n297 gnd 0.070438f
C2206 commonsourceibias.n298 gnd 0.009449f
C2207 commonsourceibias.t137 gnd 0.176537f
C2208 commonsourceibias.n299 gnd 0.070438f
C2209 commonsourceibias.n300 gnd 0.009449f
C2210 commonsourceibias.t133 gnd 0.176537f
C2211 commonsourceibias.n301 gnd 0.070438f
C2212 commonsourceibias.n302 gnd 0.009449f
C2213 commonsourceibias.t149 gnd 0.176537f
C2214 commonsourceibias.n303 gnd 0.010741f
C2215 commonsourceibias.n304 gnd 0.009449f
C2216 commonsourceibias.t79 gnd 0.176537f
C2217 commonsourceibias.n305 gnd 0.012701f
C2218 commonsourceibias.t140 gnd 0.196658f
C2219 commonsourceibias.t130 gnd 0.176537f
C2220 commonsourceibias.n306 gnd 0.078486f
C2221 commonsourceibias.n307 gnd 0.084086f
C2222 commonsourceibias.n308 gnd 0.04022f
C2223 commonsourceibias.n309 gnd 0.009449f
C2224 commonsourceibias.n310 gnd 0.00768f
C2225 commonsourceibias.n311 gnd 0.013021f
C2226 commonsourceibias.n312 gnd 0.070438f
C2227 commonsourceibias.n313 gnd 0.013076f
C2228 commonsourceibias.n314 gnd 0.009449f
C2229 commonsourceibias.n315 gnd 0.009449f
C2230 commonsourceibias.n316 gnd 0.009449f
C2231 commonsourceibias.n317 gnd 0.009585f
C2232 commonsourceibias.n318 gnd 0.070438f
C2233 commonsourceibias.n319 gnd 0.011646f
C2234 commonsourceibias.n320 gnd 0.012884f
C2235 commonsourceibias.n321 gnd 0.009449f
C2236 commonsourceibias.n322 gnd 0.009449f
C2237 commonsourceibias.n323 gnd 0.0128f
C2238 commonsourceibias.n324 gnd 0.007644f
C2239 commonsourceibias.n325 gnd 0.012959f
C2240 commonsourceibias.n326 gnd 0.009449f
C2241 commonsourceibias.n327 gnd 0.009449f
C2242 commonsourceibias.n328 gnd 0.013038f
C2243 commonsourceibias.n329 gnd 0.011242f
C2244 commonsourceibias.n330 gnd 0.009122f
C2245 commonsourceibias.n331 gnd 0.009449f
C2246 commonsourceibias.n332 gnd 0.009449f
C2247 commonsourceibias.n333 gnd 0.011558f
C2248 commonsourceibias.n334 gnd 0.012972f
C2249 commonsourceibias.n335 gnd 0.070438f
C2250 commonsourceibias.n336 gnd 0.012885f
C2251 commonsourceibias.n337 gnd 0.009449f
C2252 commonsourceibias.n338 gnd 0.009449f
C2253 commonsourceibias.n339 gnd 0.009449f
C2254 commonsourceibias.n340 gnd 0.012885f
C2255 commonsourceibias.n341 gnd 0.070438f
C2256 commonsourceibias.n342 gnd 0.012972f
C2257 commonsourceibias.n343 gnd 0.011558f
C2258 commonsourceibias.n344 gnd 0.009449f
C2259 commonsourceibias.n345 gnd 0.009449f
C2260 commonsourceibias.n346 gnd 0.009449f
C2261 commonsourceibias.n347 gnd 0.011242f
C2262 commonsourceibias.n348 gnd 0.013038f
C2263 commonsourceibias.n349 gnd 0.070438f
C2264 commonsourceibias.n350 gnd 0.012959f
C2265 commonsourceibias.n351 gnd 0.009449f
C2266 commonsourceibias.n352 gnd 0.009449f
C2267 commonsourceibias.n353 gnd 0.009449f
C2268 commonsourceibias.n354 gnd 0.0128f
C2269 commonsourceibias.n355 gnd 0.070438f
C2270 commonsourceibias.n356 gnd 0.012884f
C2271 commonsourceibias.n357 gnd 0.011646f
C2272 commonsourceibias.n358 gnd 0.009449f
C2273 commonsourceibias.n359 gnd 0.009449f
C2274 commonsourceibias.n360 gnd 0.009449f
C2275 commonsourceibias.n361 gnd 0.010741f
C2276 commonsourceibias.n362 gnd 0.013076f
C2277 commonsourceibias.n363 gnd 0.070438f
C2278 commonsourceibias.n364 gnd 0.013021f
C2279 commonsourceibias.n365 gnd 0.009449f
C2280 commonsourceibias.n366 gnd 0.009449f
C2281 commonsourceibias.n367 gnd 0.009449f
C2282 commonsourceibias.n368 gnd 0.012701f
C2283 commonsourceibias.n369 gnd 0.070438f
C2284 commonsourceibias.n370 gnd 0.012732f
C2285 commonsourceibias.t147 gnd 0.190924f
C2286 commonsourceibias.n371 gnd 0.084938f
C2287 commonsourceibias.n372 gnd 0.03031f
C2288 commonsourceibias.n373 gnd 0.449124f
C2289 commonsourceibias.n374 gnd 0.012609f
C2290 commonsourceibias.t91 gnd 0.190924f
C2291 commonsourceibias.t134 gnd 0.176537f
C2292 commonsourceibias.n375 gnd 0.00768f
C2293 commonsourceibias.n376 gnd 0.009449f
C2294 commonsourceibias.t114 gnd 0.176537f
C2295 commonsourceibias.n377 gnd 0.009585f
C2296 commonsourceibias.n378 gnd 0.009449f
C2297 commonsourceibias.t123 gnd 0.176537f
C2298 commonsourceibias.n379 gnd 0.007644f
C2299 commonsourceibias.n380 gnd 0.009449f
C2300 commonsourceibias.t88 gnd 0.176537f
C2301 commonsourceibias.n381 gnd 0.009122f
C2302 commonsourceibias.n382 gnd 0.009449f
C2303 commonsourceibias.t104 gnd 0.176537f
C2304 commonsourceibias.n383 gnd 0.007632f
C2305 commonsourceibias.n384 gnd 0.009449f
C2306 commonsourceibias.t89 gnd 0.176537f
C2307 commonsourceibias.t139 gnd 0.176537f
C2308 commonsourceibias.n385 gnd 0.070438f
C2309 commonsourceibias.n386 gnd 0.009449f
C2310 commonsourceibias.t83 gnd 0.176537f
C2311 commonsourceibias.n387 gnd 0.070438f
C2312 commonsourceibias.n388 gnd 0.009449f
C2313 commonsourceibias.t150 gnd 0.176537f
C2314 commonsourceibias.n389 gnd 0.070438f
C2315 commonsourceibias.n390 gnd 0.009449f
C2316 commonsourceibias.t127 gnd 0.176537f
C2317 commonsourceibias.n391 gnd 0.010741f
C2318 commonsourceibias.n392 gnd 0.009449f
C2319 commonsourceibias.t84 gnd 0.176537f
C2320 commonsourceibias.n393 gnd 0.012701f
C2321 commonsourceibias.t108 gnd 0.196658f
C2322 commonsourceibias.t131 gnd 0.176537f
C2323 commonsourceibias.n394 gnd 0.078486f
C2324 commonsourceibias.n395 gnd 0.084086f
C2325 commonsourceibias.n396 gnd 0.04022f
C2326 commonsourceibias.n397 gnd 0.009449f
C2327 commonsourceibias.n398 gnd 0.00768f
C2328 commonsourceibias.n399 gnd 0.013021f
C2329 commonsourceibias.n400 gnd 0.070438f
C2330 commonsourceibias.n401 gnd 0.013076f
C2331 commonsourceibias.n402 gnd 0.009449f
C2332 commonsourceibias.n403 gnd 0.009449f
C2333 commonsourceibias.n404 gnd 0.009449f
C2334 commonsourceibias.n405 gnd 0.009585f
C2335 commonsourceibias.n406 gnd 0.070438f
C2336 commonsourceibias.n407 gnd 0.011646f
C2337 commonsourceibias.n408 gnd 0.012884f
C2338 commonsourceibias.n409 gnd 0.009449f
C2339 commonsourceibias.n410 gnd 0.009449f
C2340 commonsourceibias.n411 gnd 0.0128f
C2341 commonsourceibias.n412 gnd 0.007644f
C2342 commonsourceibias.n413 gnd 0.012959f
C2343 commonsourceibias.n414 gnd 0.009449f
C2344 commonsourceibias.n415 gnd 0.009449f
C2345 commonsourceibias.n416 gnd 0.013038f
C2346 commonsourceibias.n417 gnd 0.011242f
C2347 commonsourceibias.n418 gnd 0.009122f
C2348 commonsourceibias.n419 gnd 0.009449f
C2349 commonsourceibias.n420 gnd 0.009449f
C2350 commonsourceibias.n421 gnd 0.011558f
C2351 commonsourceibias.n422 gnd 0.012972f
C2352 commonsourceibias.n423 gnd 0.070438f
C2353 commonsourceibias.n424 gnd 0.012885f
C2354 commonsourceibias.n425 gnd 0.009404f
C2355 commonsourceibias.t7 gnd 0.02039f
C2356 commonsourceibias.t51 gnd 0.02039f
C2357 commonsourceibias.n426 gnd 0.180776f
C2358 commonsourceibias.t37 gnd 0.02039f
C2359 commonsourceibias.t53 gnd 0.02039f
C2360 commonsourceibias.n427 gnd 0.180173f
C2361 commonsourceibias.n428 gnd 0.167888f
C2362 commonsourceibias.t1 gnd 0.02039f
C2363 commonsourceibias.t35 gnd 0.02039f
C2364 commonsourceibias.n429 gnd 0.180173f
C2365 commonsourceibias.n430 gnd 0.082761f
C2366 commonsourceibias.t3 gnd 0.02039f
C2367 commonsourceibias.t31 gnd 0.02039f
C2368 commonsourceibias.n431 gnd 0.180173f
C2369 commonsourceibias.n432 gnd 0.069143f
C2370 commonsourceibias.n433 gnd 0.012609f
C2371 commonsourceibias.t48 gnd 0.176537f
C2372 commonsourceibias.n434 gnd 0.00768f
C2373 commonsourceibias.n435 gnd 0.009449f
C2374 commonsourceibias.t44 gnd 0.176537f
C2375 commonsourceibias.n436 gnd 0.009585f
C2376 commonsourceibias.n437 gnd 0.009449f
C2377 commonsourceibias.t4 gnd 0.176537f
C2378 commonsourceibias.n438 gnd 0.007644f
C2379 commonsourceibias.n439 gnd 0.009449f
C2380 commonsourceibias.t32 gnd 0.176537f
C2381 commonsourceibias.n440 gnd 0.009122f
C2382 commonsourceibias.n441 gnd 0.009449f
C2383 commonsourceibias.t10 gnd 0.176537f
C2384 commonsourceibias.n442 gnd 0.007632f
C2385 commonsourceibias.n443 gnd 0.009449f
C2386 commonsourceibias.t30 gnd 0.176537f
C2387 commonsourceibias.t2 gnd 0.176537f
C2388 commonsourceibias.n444 gnd 0.070438f
C2389 commonsourceibias.n445 gnd 0.009449f
C2390 commonsourceibias.t34 gnd 0.176537f
C2391 commonsourceibias.n446 gnd 0.070438f
C2392 commonsourceibias.n447 gnd 0.009449f
C2393 commonsourceibias.t0 gnd 0.176537f
C2394 commonsourceibias.n448 gnd 0.070438f
C2395 commonsourceibias.n449 gnd 0.009449f
C2396 commonsourceibias.t52 gnd 0.176537f
C2397 commonsourceibias.n450 gnd 0.010741f
C2398 commonsourceibias.n451 gnd 0.009449f
C2399 commonsourceibias.t36 gnd 0.176537f
C2400 commonsourceibias.n452 gnd 0.012701f
C2401 commonsourceibias.t6 gnd 0.196658f
C2402 commonsourceibias.t50 gnd 0.176537f
C2403 commonsourceibias.n453 gnd 0.078486f
C2404 commonsourceibias.n454 gnd 0.084086f
C2405 commonsourceibias.n455 gnd 0.04022f
C2406 commonsourceibias.n456 gnd 0.009449f
C2407 commonsourceibias.n457 gnd 0.00768f
C2408 commonsourceibias.n458 gnd 0.013021f
C2409 commonsourceibias.n459 gnd 0.070438f
C2410 commonsourceibias.n460 gnd 0.013076f
C2411 commonsourceibias.n461 gnd 0.009449f
C2412 commonsourceibias.n462 gnd 0.009449f
C2413 commonsourceibias.n463 gnd 0.009449f
C2414 commonsourceibias.n464 gnd 0.009585f
C2415 commonsourceibias.n465 gnd 0.070438f
C2416 commonsourceibias.n466 gnd 0.011646f
C2417 commonsourceibias.n467 gnd 0.012884f
C2418 commonsourceibias.n468 gnd 0.009449f
C2419 commonsourceibias.n469 gnd 0.009449f
C2420 commonsourceibias.n470 gnd 0.0128f
C2421 commonsourceibias.n471 gnd 0.007644f
C2422 commonsourceibias.n472 gnd 0.012959f
C2423 commonsourceibias.n473 gnd 0.009449f
C2424 commonsourceibias.n474 gnd 0.009449f
C2425 commonsourceibias.n475 gnd 0.013038f
C2426 commonsourceibias.n476 gnd 0.011242f
C2427 commonsourceibias.n477 gnd 0.009122f
C2428 commonsourceibias.n478 gnd 0.009449f
C2429 commonsourceibias.n479 gnd 0.009449f
C2430 commonsourceibias.n480 gnd 0.011558f
C2431 commonsourceibias.n481 gnd 0.012972f
C2432 commonsourceibias.n482 gnd 0.070438f
C2433 commonsourceibias.n483 gnd 0.012885f
C2434 commonsourceibias.n484 gnd 0.009449f
C2435 commonsourceibias.n485 gnd 0.009449f
C2436 commonsourceibias.n486 gnd 0.009449f
C2437 commonsourceibias.n487 gnd 0.012885f
C2438 commonsourceibias.n488 gnd 0.070438f
C2439 commonsourceibias.n489 gnd 0.012972f
C2440 commonsourceibias.t40 gnd 0.176537f
C2441 commonsourceibias.n490 gnd 0.070438f
C2442 commonsourceibias.n491 gnd 0.011558f
C2443 commonsourceibias.n492 gnd 0.009449f
C2444 commonsourceibias.n493 gnd 0.009449f
C2445 commonsourceibias.n494 gnd 0.009449f
C2446 commonsourceibias.n495 gnd 0.011242f
C2447 commonsourceibias.n496 gnd 0.013038f
C2448 commonsourceibias.n497 gnd 0.070438f
C2449 commonsourceibias.n498 gnd 0.012959f
C2450 commonsourceibias.n499 gnd 0.009449f
C2451 commonsourceibias.n500 gnd 0.009449f
C2452 commonsourceibias.n501 gnd 0.009449f
C2453 commonsourceibias.n502 gnd 0.0128f
C2454 commonsourceibias.n503 gnd 0.070438f
C2455 commonsourceibias.n504 gnd 0.012884f
C2456 commonsourceibias.t26 gnd 0.176537f
C2457 commonsourceibias.n505 gnd 0.070438f
C2458 commonsourceibias.n506 gnd 0.011646f
C2459 commonsourceibias.n507 gnd 0.009449f
C2460 commonsourceibias.n508 gnd 0.009449f
C2461 commonsourceibias.n509 gnd 0.009449f
C2462 commonsourceibias.n510 gnd 0.010741f
C2463 commonsourceibias.n511 gnd 0.013076f
C2464 commonsourceibias.n512 gnd 0.070438f
C2465 commonsourceibias.n513 gnd 0.013021f
C2466 commonsourceibias.n514 gnd 0.009449f
C2467 commonsourceibias.n515 gnd 0.009449f
C2468 commonsourceibias.n516 gnd 0.009449f
C2469 commonsourceibias.n517 gnd 0.012701f
C2470 commonsourceibias.n518 gnd 0.070438f
C2471 commonsourceibias.n519 gnd 0.012732f
C2472 commonsourceibias.t28 gnd 0.190924f
C2473 commonsourceibias.n520 gnd 0.084938f
C2474 commonsourceibias.n521 gnd 0.094974f
C2475 commonsourceibias.t49 gnd 0.02039f
C2476 commonsourceibias.t29 gnd 0.02039f
C2477 commonsourceibias.n522 gnd 0.180173f
C2478 commonsourceibias.n523 gnd 0.156069f
C2479 commonsourceibias.t27 gnd 0.02039f
C2480 commonsourceibias.t45 gnd 0.02039f
C2481 commonsourceibias.n524 gnd 0.180173f
C2482 commonsourceibias.n525 gnd 0.082761f
C2483 commonsourceibias.t33 gnd 0.02039f
C2484 commonsourceibias.t5 gnd 0.02039f
C2485 commonsourceibias.n526 gnd 0.180173f
C2486 commonsourceibias.n527 gnd 0.082761f
C2487 commonsourceibias.t11 gnd 0.02039f
C2488 commonsourceibias.t41 gnd 0.02039f
C2489 commonsourceibias.n528 gnd 0.180173f
C2490 commonsourceibias.n529 gnd 0.069143f
C2491 commonsourceibias.n530 gnd 0.083724f
C2492 commonsourceibias.n531 gnd 0.068305f
C2493 commonsourceibias.n532 gnd 0.009404f
C2494 commonsourceibias.n533 gnd 0.012885f
C2495 commonsourceibias.n534 gnd 0.070438f
C2496 commonsourceibias.n535 gnd 0.012972f
C2497 commonsourceibias.t73 gnd 0.176537f
C2498 commonsourceibias.n536 gnd 0.070438f
C2499 commonsourceibias.n537 gnd 0.011558f
C2500 commonsourceibias.n538 gnd 0.009449f
C2501 commonsourceibias.n539 gnd 0.009449f
C2502 commonsourceibias.n540 gnd 0.009449f
C2503 commonsourceibias.n541 gnd 0.011242f
C2504 commonsourceibias.n542 gnd 0.013038f
C2505 commonsourceibias.n543 gnd 0.070438f
C2506 commonsourceibias.n544 gnd 0.012959f
C2507 commonsourceibias.n545 gnd 0.009449f
C2508 commonsourceibias.n546 gnd 0.009449f
C2509 commonsourceibias.n547 gnd 0.009449f
C2510 commonsourceibias.n548 gnd 0.0128f
C2511 commonsourceibias.n549 gnd 0.070438f
C2512 commonsourceibias.n550 gnd 0.012884f
C2513 commonsourceibias.t95 gnd 0.176537f
C2514 commonsourceibias.n551 gnd 0.070438f
C2515 commonsourceibias.n552 gnd 0.011646f
C2516 commonsourceibias.n553 gnd 0.009449f
C2517 commonsourceibias.n554 gnd 0.009449f
C2518 commonsourceibias.n555 gnd 0.009449f
C2519 commonsourceibias.n556 gnd 0.010741f
C2520 commonsourceibias.n557 gnd 0.013076f
C2521 commonsourceibias.n558 gnd 0.070438f
C2522 commonsourceibias.n559 gnd 0.013021f
C2523 commonsourceibias.n560 gnd 0.009449f
C2524 commonsourceibias.n561 gnd 0.009449f
C2525 commonsourceibias.n562 gnd 0.009449f
C2526 commonsourceibias.n563 gnd 0.012701f
C2527 commonsourceibias.n564 gnd 0.070438f
C2528 commonsourceibias.n565 gnd 0.012732f
C2529 commonsourceibias.n566 gnd 0.084938f
C2530 commonsourceibias.n567 gnd 0.056112f
C2531 commonsourceibias.n568 gnd 0.012609f
C2532 commonsourceibias.t144 gnd 0.176537f
C2533 commonsourceibias.n569 gnd 0.00768f
C2534 commonsourceibias.n570 gnd 0.009449f
C2535 commonsourceibias.t66 gnd 0.176537f
C2536 commonsourceibias.n571 gnd 0.009585f
C2537 commonsourceibias.n572 gnd 0.009449f
C2538 commonsourceibias.t143 gnd 0.176537f
C2539 commonsourceibias.n573 gnd 0.007644f
C2540 commonsourceibias.n574 gnd 0.009449f
C2541 commonsourceibias.t65 gnd 0.176537f
C2542 commonsourceibias.n575 gnd 0.009122f
C2543 commonsourceibias.n576 gnd 0.009449f
C2544 commonsourceibias.t142 gnd 0.176537f
C2545 commonsourceibias.n577 gnd 0.007632f
C2546 commonsourceibias.n578 gnd 0.009449f
C2547 commonsourceibias.t72 gnd 0.176537f
C2548 commonsourceibias.t99 gnd 0.176537f
C2549 commonsourceibias.n579 gnd 0.070438f
C2550 commonsourceibias.n580 gnd 0.009449f
C2551 commonsourceibias.t80 gnd 0.176537f
C2552 commonsourceibias.n581 gnd 0.070438f
C2553 commonsourceibias.n582 gnd 0.009449f
C2554 commonsourceibias.t69 gnd 0.176537f
C2555 commonsourceibias.n583 gnd 0.070438f
C2556 commonsourceibias.n584 gnd 0.009449f
C2557 commonsourceibias.t98 gnd 0.176537f
C2558 commonsourceibias.n585 gnd 0.010741f
C2559 commonsourceibias.n586 gnd 0.009449f
C2560 commonsourceibias.t86 gnd 0.176537f
C2561 commonsourceibias.n587 gnd 0.012701f
C2562 commonsourceibias.t97 gnd 0.196658f
C2563 commonsourceibias.t68 gnd 0.176537f
C2564 commonsourceibias.n588 gnd 0.078486f
C2565 commonsourceibias.n589 gnd 0.084086f
C2566 commonsourceibias.n590 gnd 0.04022f
C2567 commonsourceibias.n591 gnd 0.009449f
C2568 commonsourceibias.n592 gnd 0.00768f
C2569 commonsourceibias.n593 gnd 0.013021f
C2570 commonsourceibias.n594 gnd 0.070438f
C2571 commonsourceibias.n595 gnd 0.013076f
C2572 commonsourceibias.n596 gnd 0.009449f
C2573 commonsourceibias.n597 gnd 0.009449f
C2574 commonsourceibias.n598 gnd 0.009449f
C2575 commonsourceibias.n599 gnd 0.009585f
C2576 commonsourceibias.n600 gnd 0.070438f
C2577 commonsourceibias.n601 gnd 0.011646f
C2578 commonsourceibias.n602 gnd 0.012884f
C2579 commonsourceibias.n603 gnd 0.009449f
C2580 commonsourceibias.n604 gnd 0.009449f
C2581 commonsourceibias.n605 gnd 0.0128f
C2582 commonsourceibias.n606 gnd 0.007644f
C2583 commonsourceibias.n607 gnd 0.012959f
C2584 commonsourceibias.n608 gnd 0.009449f
C2585 commonsourceibias.n609 gnd 0.009449f
C2586 commonsourceibias.n610 gnd 0.013038f
C2587 commonsourceibias.n611 gnd 0.011242f
C2588 commonsourceibias.n612 gnd 0.009122f
C2589 commonsourceibias.n613 gnd 0.009449f
C2590 commonsourceibias.n614 gnd 0.009449f
C2591 commonsourceibias.n615 gnd 0.011558f
C2592 commonsourceibias.n616 gnd 0.012972f
C2593 commonsourceibias.n617 gnd 0.070438f
C2594 commonsourceibias.n618 gnd 0.012885f
C2595 commonsourceibias.n619 gnd 0.009449f
C2596 commonsourceibias.n620 gnd 0.009449f
C2597 commonsourceibias.n621 gnd 0.009449f
C2598 commonsourceibias.n622 gnd 0.012885f
C2599 commonsourceibias.n623 gnd 0.070438f
C2600 commonsourceibias.n624 gnd 0.012972f
C2601 commonsourceibias.t100 gnd 0.176537f
C2602 commonsourceibias.n625 gnd 0.070438f
C2603 commonsourceibias.n626 gnd 0.011558f
C2604 commonsourceibias.n627 gnd 0.009449f
C2605 commonsourceibias.n628 gnd 0.009449f
C2606 commonsourceibias.n629 gnd 0.009449f
C2607 commonsourceibias.n630 gnd 0.011242f
C2608 commonsourceibias.n631 gnd 0.013038f
C2609 commonsourceibias.n632 gnd 0.070438f
C2610 commonsourceibias.n633 gnd 0.012959f
C2611 commonsourceibias.n634 gnd 0.009449f
C2612 commonsourceibias.n635 gnd 0.009449f
C2613 commonsourceibias.n636 gnd 0.009449f
C2614 commonsourceibias.n637 gnd 0.0128f
C2615 commonsourceibias.n638 gnd 0.070438f
C2616 commonsourceibias.n639 gnd 0.012884f
C2617 commonsourceibias.t154 gnd 0.176537f
C2618 commonsourceibias.n640 gnd 0.070438f
C2619 commonsourceibias.n641 gnd 0.011646f
C2620 commonsourceibias.n642 gnd 0.009449f
C2621 commonsourceibias.n643 gnd 0.009449f
C2622 commonsourceibias.n644 gnd 0.009449f
C2623 commonsourceibias.n645 gnd 0.010741f
C2624 commonsourceibias.n646 gnd 0.013076f
C2625 commonsourceibias.n647 gnd 0.070438f
C2626 commonsourceibias.n648 gnd 0.013021f
C2627 commonsourceibias.n649 gnd 0.009449f
C2628 commonsourceibias.n650 gnd 0.009449f
C2629 commonsourceibias.n651 gnd 0.009449f
C2630 commonsourceibias.n652 gnd 0.012701f
C2631 commonsourceibias.n653 gnd 0.070438f
C2632 commonsourceibias.n654 gnd 0.012732f
C2633 commonsourceibias.t151 gnd 0.190924f
C2634 commonsourceibias.n655 gnd 0.084938f
C2635 commonsourceibias.n656 gnd 0.03031f
C2636 commonsourceibias.n657 gnd 0.151321f
C2637 commonsourceibias.n658 gnd 0.012609f
C2638 commonsourceibias.t107 gnd 0.176537f
C2639 commonsourceibias.n659 gnd 0.00768f
C2640 commonsourceibias.n660 gnd 0.009449f
C2641 commonsourceibias.t122 gnd 0.176537f
C2642 commonsourceibias.n661 gnd 0.009585f
C2643 commonsourceibias.n662 gnd 0.009449f
C2644 commonsourceibias.t101 gnd 0.176537f
C2645 commonsourceibias.n663 gnd 0.007644f
C2646 commonsourceibias.n664 gnd 0.009449f
C2647 commonsourceibias.t115 gnd 0.176537f
C2648 commonsourceibias.n665 gnd 0.009122f
C2649 commonsourceibias.n666 gnd 0.009449f
C2650 commonsourceibias.t81 gnd 0.176537f
C2651 commonsourceibias.n667 gnd 0.007632f
C2652 commonsourceibias.n668 gnd 0.009449f
C2653 commonsourceibias.t70 gnd 0.176537f
C2654 commonsourceibias.t103 gnd 0.176537f
C2655 commonsourceibias.n669 gnd 0.070438f
C2656 commonsourceibias.n670 gnd 0.009449f
C2657 commonsourceibias.t132 gnd 0.176537f
C2658 commonsourceibias.n671 gnd 0.070438f
C2659 commonsourceibias.n672 gnd 0.009449f
C2660 commonsourceibias.t153 gnd 0.176537f
C2661 commonsourceibias.n673 gnd 0.070438f
C2662 commonsourceibias.n674 gnd 0.009449f
C2663 commonsourceibias.t87 gnd 0.176537f
C2664 commonsourceibias.n675 gnd 0.010741f
C2665 commonsourceibias.n676 gnd 0.009449f
C2666 commonsourceibias.t109 gnd 0.176537f
C2667 commonsourceibias.n677 gnd 0.012701f
C2668 commonsourceibias.t74 gnd 0.196658f
C2669 commonsourceibias.t145 gnd 0.176537f
C2670 commonsourceibias.n678 gnd 0.078486f
C2671 commonsourceibias.n679 gnd 0.084086f
C2672 commonsourceibias.n680 gnd 0.04022f
C2673 commonsourceibias.n681 gnd 0.009449f
C2674 commonsourceibias.n682 gnd 0.00768f
C2675 commonsourceibias.n683 gnd 0.013021f
C2676 commonsourceibias.n684 gnd 0.070438f
C2677 commonsourceibias.n685 gnd 0.013076f
C2678 commonsourceibias.n686 gnd 0.009449f
C2679 commonsourceibias.n687 gnd 0.009449f
C2680 commonsourceibias.n688 gnd 0.009449f
C2681 commonsourceibias.n689 gnd 0.009585f
C2682 commonsourceibias.n690 gnd 0.070438f
C2683 commonsourceibias.n691 gnd 0.011646f
C2684 commonsourceibias.n692 gnd 0.012884f
C2685 commonsourceibias.n693 gnd 0.009449f
C2686 commonsourceibias.n694 gnd 0.009449f
C2687 commonsourceibias.n695 gnd 0.0128f
C2688 commonsourceibias.n696 gnd 0.007644f
C2689 commonsourceibias.n697 gnd 0.012959f
C2690 commonsourceibias.n698 gnd 0.009449f
C2691 commonsourceibias.n699 gnd 0.009449f
C2692 commonsourceibias.n700 gnd 0.013038f
C2693 commonsourceibias.n701 gnd 0.011242f
C2694 commonsourceibias.n702 gnd 0.009122f
C2695 commonsourceibias.n703 gnd 0.009449f
C2696 commonsourceibias.n704 gnd 0.009449f
C2697 commonsourceibias.n705 gnd 0.011558f
C2698 commonsourceibias.n706 gnd 0.012972f
C2699 commonsourceibias.n707 gnd 0.070438f
C2700 commonsourceibias.n708 gnd 0.012885f
C2701 commonsourceibias.n709 gnd 0.009449f
C2702 commonsourceibias.n710 gnd 0.009449f
C2703 commonsourceibias.n711 gnd 0.009449f
C2704 commonsourceibias.n712 gnd 0.012885f
C2705 commonsourceibias.n713 gnd 0.070438f
C2706 commonsourceibias.n714 gnd 0.012972f
C2707 commonsourceibias.t110 gnd 0.176537f
C2708 commonsourceibias.n715 gnd 0.070438f
C2709 commonsourceibias.n716 gnd 0.011558f
C2710 commonsourceibias.n717 gnd 0.009449f
C2711 commonsourceibias.n718 gnd 0.009449f
C2712 commonsourceibias.n719 gnd 0.009449f
C2713 commonsourceibias.n720 gnd 0.011242f
C2714 commonsourceibias.n721 gnd 0.013038f
C2715 commonsourceibias.n722 gnd 0.070438f
C2716 commonsourceibias.n723 gnd 0.012959f
C2717 commonsourceibias.n724 gnd 0.009449f
C2718 commonsourceibias.n725 gnd 0.009449f
C2719 commonsourceibias.n726 gnd 0.009449f
C2720 commonsourceibias.n727 gnd 0.0128f
C2721 commonsourceibias.n728 gnd 0.070438f
C2722 commonsourceibias.n729 gnd 0.012884f
C2723 commonsourceibias.t135 gnd 0.176537f
C2724 commonsourceibias.n730 gnd 0.070438f
C2725 commonsourceibias.n731 gnd 0.011646f
C2726 commonsourceibias.n732 gnd 0.009449f
C2727 commonsourceibias.n733 gnd 0.009449f
C2728 commonsourceibias.n734 gnd 0.009449f
C2729 commonsourceibias.n735 gnd 0.010741f
C2730 commonsourceibias.n736 gnd 0.013076f
C2731 commonsourceibias.n737 gnd 0.070438f
C2732 commonsourceibias.n738 gnd 0.013021f
C2733 commonsourceibias.n739 gnd 0.009449f
C2734 commonsourceibias.n740 gnd 0.009449f
C2735 commonsourceibias.n741 gnd 0.009449f
C2736 commonsourceibias.n742 gnd 0.012701f
C2737 commonsourceibias.n743 gnd 0.070438f
C2738 commonsourceibias.n744 gnd 0.012732f
C2739 commonsourceibias.t82 gnd 0.190924f
C2740 commonsourceibias.n745 gnd 0.084938f
C2741 commonsourceibias.n746 gnd 0.03031f
C2742 commonsourceibias.n747 gnd 0.199407f
C2743 commonsourceibias.n748 gnd 5.05322f
C2744 vdd.t185 gnd 0.037058f
C2745 vdd.t165 gnd 0.037058f
C2746 vdd.n0 gnd 0.29228f
C2747 vdd.t144 gnd 0.037058f
C2748 vdd.t181 gnd 0.037058f
C2749 vdd.n1 gnd 0.291797f
C2750 vdd.n2 gnd 0.269092f
C2751 vdd.t162 gnd 0.037058f
C2752 vdd.t192 gnd 0.037058f
C2753 vdd.n3 gnd 0.291797f
C2754 vdd.n4 gnd 0.13609f
C2755 vdd.t190 gnd 0.037058f
C2756 vdd.t170 gnd 0.037058f
C2757 vdd.n5 gnd 0.291797f
C2758 vdd.n6 gnd 0.127695f
C2759 vdd.t196 gnd 0.037058f
C2760 vdd.t160 gnd 0.037058f
C2761 vdd.n7 gnd 0.29228f
C2762 vdd.t168 gnd 0.037058f
C2763 vdd.t188 gnd 0.037058f
C2764 vdd.n8 gnd 0.291797f
C2765 vdd.n9 gnd 0.269093f
C2766 vdd.t177 gnd 0.037058f
C2767 vdd.t148 gnd 0.037058f
C2768 vdd.n10 gnd 0.291797f
C2769 vdd.n11 gnd 0.13609f
C2770 vdd.t157 gnd 0.037058f
C2771 vdd.t175 gnd 0.037058f
C2772 vdd.n12 gnd 0.291797f
C2773 vdd.n13 gnd 0.127695f
C2774 vdd.n14 gnd 0.090278f
C2775 vdd.t49 gnd 0.020588f
C2776 vdd.t8 gnd 0.020588f
C2777 vdd.n15 gnd 0.1895f
C2778 vdd.t45 gnd 0.020588f
C2779 vdd.t47 gnd 0.020588f
C2780 vdd.n16 gnd 0.188945f
C2781 vdd.n17 gnd 0.328824f
C2782 vdd.t40 gnd 0.020588f
C2783 vdd.t4 gnd 0.020588f
C2784 vdd.n18 gnd 0.188945f
C2785 vdd.n19 gnd 0.136039f
C2786 vdd.t6 gnd 0.020588f
C2787 vdd.t48 gnd 0.020588f
C2788 vdd.n20 gnd 0.1895f
C2789 vdd.t50 gnd 0.020588f
C2790 vdd.t39 gnd 0.020588f
C2791 vdd.n21 gnd 0.188945f
C2792 vdd.n22 gnd 0.328824f
C2793 vdd.t5 gnd 0.020588f
C2794 vdd.t83 gnd 0.020588f
C2795 vdd.n23 gnd 0.188945f
C2796 vdd.n24 gnd 0.136039f
C2797 vdd.t41 gnd 0.020588f
C2798 vdd.t7 gnd 0.020588f
C2799 vdd.n25 gnd 0.188945f
C2800 vdd.t46 gnd 0.020588f
C2801 vdd.t84 gnd 0.020588f
C2802 vdd.n26 gnd 0.188945f
C2803 vdd.n27 gnd 20.7697f
C2804 vdd.n28 gnd 8.3397f
C2805 vdd.n29 gnd 0.005615f
C2806 vdd.n30 gnd 0.005211f
C2807 vdd.n31 gnd 0.002882f
C2808 vdd.n32 gnd 0.006618f
C2809 vdd.n33 gnd 0.0028f
C2810 vdd.n34 gnd 0.002965f
C2811 vdd.n35 gnd 0.005211f
C2812 vdd.n36 gnd 0.0028f
C2813 vdd.n37 gnd 0.006618f
C2814 vdd.n38 gnd 0.002965f
C2815 vdd.n39 gnd 0.005211f
C2816 vdd.n40 gnd 0.0028f
C2817 vdd.n41 gnd 0.004963f
C2818 vdd.n42 gnd 0.004978f
C2819 vdd.t14 gnd 0.014218f
C2820 vdd.n43 gnd 0.031635f
C2821 vdd.n44 gnd 0.164637f
C2822 vdd.n45 gnd 0.0028f
C2823 vdd.n46 gnd 0.002965f
C2824 vdd.n47 gnd 0.006618f
C2825 vdd.n48 gnd 0.006618f
C2826 vdd.n49 gnd 0.002965f
C2827 vdd.n50 gnd 0.0028f
C2828 vdd.n51 gnd 0.005211f
C2829 vdd.n52 gnd 0.005211f
C2830 vdd.n53 gnd 0.0028f
C2831 vdd.n54 gnd 0.002965f
C2832 vdd.n55 gnd 0.006618f
C2833 vdd.n56 gnd 0.006618f
C2834 vdd.n57 gnd 0.002965f
C2835 vdd.n58 gnd 0.0028f
C2836 vdd.n59 gnd 0.005211f
C2837 vdd.n60 gnd 0.005211f
C2838 vdd.n61 gnd 0.0028f
C2839 vdd.n62 gnd 0.002965f
C2840 vdd.n63 gnd 0.006618f
C2841 vdd.n64 gnd 0.006618f
C2842 vdd.n65 gnd 0.015646f
C2843 vdd.n66 gnd 0.002882f
C2844 vdd.n67 gnd 0.0028f
C2845 vdd.n68 gnd 0.013467f
C2846 vdd.n69 gnd 0.009402f
C2847 vdd.t139 gnd 0.03294f
C2848 vdd.t228 gnd 0.03294f
C2849 vdd.n70 gnd 0.226387f
C2850 vdd.n71 gnd 0.178019f
C2851 vdd.t133 gnd 0.03294f
C2852 vdd.t3 gnd 0.03294f
C2853 vdd.n72 gnd 0.226387f
C2854 vdd.n73 gnd 0.14366f
C2855 vdd.t78 gnd 0.03294f
C2856 vdd.t79 gnd 0.03294f
C2857 vdd.n74 gnd 0.226387f
C2858 vdd.n75 gnd 0.14366f
C2859 vdd.t56 gnd 0.03294f
C2860 vdd.t28 gnd 0.03294f
C2861 vdd.n76 gnd 0.226387f
C2862 vdd.n77 gnd 0.14366f
C2863 vdd.t20 gnd 0.03294f
C2864 vdd.t135 gnd 0.03294f
C2865 vdd.n78 gnd 0.226387f
C2866 vdd.n79 gnd 0.14366f
C2867 vdd.t121 gnd 0.03294f
C2868 vdd.t212 gnd 0.03294f
C2869 vdd.n80 gnd 0.226387f
C2870 vdd.n81 gnd 0.14366f
C2871 vdd.t218 gnd 0.03294f
C2872 vdd.t118 gnd 0.03294f
C2873 vdd.n82 gnd 0.226387f
C2874 vdd.n83 gnd 0.14366f
C2875 vdd.t103 gnd 0.03294f
C2876 vdd.t73 gnd 0.03294f
C2877 vdd.n84 gnd 0.226387f
C2878 vdd.n85 gnd 0.14366f
C2879 vdd.t89 gnd 0.03294f
C2880 vdd.t26 gnd 0.03294f
C2881 vdd.n86 gnd 0.226387f
C2882 vdd.n87 gnd 0.14366f
C2883 vdd.n88 gnd 0.005615f
C2884 vdd.n89 gnd 0.005211f
C2885 vdd.n90 gnd 0.002882f
C2886 vdd.n91 gnd 0.006618f
C2887 vdd.n92 gnd 0.0028f
C2888 vdd.n93 gnd 0.002965f
C2889 vdd.n94 gnd 0.005211f
C2890 vdd.n95 gnd 0.0028f
C2891 vdd.n96 gnd 0.006618f
C2892 vdd.n97 gnd 0.002965f
C2893 vdd.n98 gnd 0.005211f
C2894 vdd.n99 gnd 0.0028f
C2895 vdd.n100 gnd 0.004963f
C2896 vdd.n101 gnd 0.004978f
C2897 vdd.t24 gnd 0.014218f
C2898 vdd.n102 gnd 0.031635f
C2899 vdd.n103 gnd 0.164637f
C2900 vdd.n104 gnd 0.0028f
C2901 vdd.n105 gnd 0.002965f
C2902 vdd.n106 gnd 0.006618f
C2903 vdd.n107 gnd 0.006618f
C2904 vdd.n108 gnd 0.002965f
C2905 vdd.n109 gnd 0.0028f
C2906 vdd.n110 gnd 0.005211f
C2907 vdd.n111 gnd 0.005211f
C2908 vdd.n112 gnd 0.0028f
C2909 vdd.n113 gnd 0.002965f
C2910 vdd.n114 gnd 0.006618f
C2911 vdd.n115 gnd 0.006618f
C2912 vdd.n116 gnd 0.002965f
C2913 vdd.n117 gnd 0.0028f
C2914 vdd.n118 gnd 0.005211f
C2915 vdd.n119 gnd 0.005211f
C2916 vdd.n120 gnd 0.0028f
C2917 vdd.n121 gnd 0.002965f
C2918 vdd.n122 gnd 0.006618f
C2919 vdd.n123 gnd 0.006618f
C2920 vdd.n124 gnd 0.015646f
C2921 vdd.n125 gnd 0.002882f
C2922 vdd.n126 gnd 0.0028f
C2923 vdd.n127 gnd 0.013467f
C2924 vdd.n128 gnd 0.009107f
C2925 vdd.n129 gnd 0.106884f
C2926 vdd.n130 gnd 0.005615f
C2927 vdd.n131 gnd 0.005211f
C2928 vdd.n132 gnd 0.002882f
C2929 vdd.n133 gnd 0.006618f
C2930 vdd.n134 gnd 0.0028f
C2931 vdd.n135 gnd 0.002965f
C2932 vdd.n136 gnd 0.005211f
C2933 vdd.n137 gnd 0.0028f
C2934 vdd.n138 gnd 0.006618f
C2935 vdd.n139 gnd 0.002965f
C2936 vdd.n140 gnd 0.005211f
C2937 vdd.n141 gnd 0.0028f
C2938 vdd.n142 gnd 0.004963f
C2939 vdd.n143 gnd 0.004978f
C2940 vdd.t138 gnd 0.014218f
C2941 vdd.n144 gnd 0.031635f
C2942 vdd.n145 gnd 0.164637f
C2943 vdd.n146 gnd 0.0028f
C2944 vdd.n147 gnd 0.002965f
C2945 vdd.n148 gnd 0.006618f
C2946 vdd.n149 gnd 0.006618f
C2947 vdd.n150 gnd 0.002965f
C2948 vdd.n151 gnd 0.0028f
C2949 vdd.n152 gnd 0.005211f
C2950 vdd.n153 gnd 0.005211f
C2951 vdd.n154 gnd 0.0028f
C2952 vdd.n155 gnd 0.002965f
C2953 vdd.n156 gnd 0.006618f
C2954 vdd.n157 gnd 0.006618f
C2955 vdd.n158 gnd 0.002965f
C2956 vdd.n159 gnd 0.0028f
C2957 vdd.n160 gnd 0.005211f
C2958 vdd.n161 gnd 0.005211f
C2959 vdd.n162 gnd 0.0028f
C2960 vdd.n163 gnd 0.002965f
C2961 vdd.n164 gnd 0.006618f
C2962 vdd.n165 gnd 0.006618f
C2963 vdd.n166 gnd 0.015646f
C2964 vdd.n167 gnd 0.002882f
C2965 vdd.n168 gnd 0.0028f
C2966 vdd.n169 gnd 0.013467f
C2967 vdd.n170 gnd 0.009402f
C2968 vdd.t117 gnd 0.03294f
C2969 vdd.t124 gnd 0.03294f
C2970 vdd.n171 gnd 0.226387f
C2971 vdd.n172 gnd 0.178019f
C2972 vdd.t110 gnd 0.03294f
C2973 vdd.t229 gnd 0.03294f
C2974 vdd.n173 gnd 0.226387f
C2975 vdd.n174 gnd 0.14366f
C2976 vdd.t220 gnd 0.03294f
C2977 vdd.t16 gnd 0.03294f
C2978 vdd.n175 gnd 0.226387f
C2979 vdd.n176 gnd 0.14366f
C2980 vdd.t136 gnd 0.03294f
C2981 vdd.t82 gnd 0.03294f
C2982 vdd.n177 gnd 0.226387f
C2983 vdd.n178 gnd 0.14366f
C2984 vdd.t42 gnd 0.03294f
C2985 vdd.t30 gnd 0.03294f
C2986 vdd.n179 gnd 0.226387f
C2987 vdd.n180 gnd 0.14366f
C2988 vdd.t217 gnd 0.03294f
C2989 vdd.t140 gnd 0.03294f
C2990 vdd.n181 gnd 0.226387f
C2991 vdd.n182 gnd 0.14366f
C2992 vdd.t105 gnd 0.03294f
C2993 vdd.t137 gnd 0.03294f
C2994 vdd.n183 gnd 0.226387f
C2995 vdd.n184 gnd 0.14366f
C2996 vdd.t125 gnd 0.03294f
C2997 vdd.t201 gnd 0.03294f
C2998 vdd.n185 gnd 0.226387f
C2999 vdd.n186 gnd 0.14366f
C3000 vdd.t112 gnd 0.03294f
C3001 vdd.t221 gnd 0.03294f
C3002 vdd.n187 gnd 0.226387f
C3003 vdd.n188 gnd 0.14366f
C3004 vdd.n189 gnd 0.005615f
C3005 vdd.n190 gnd 0.005211f
C3006 vdd.n191 gnd 0.002882f
C3007 vdd.n192 gnd 0.006618f
C3008 vdd.n193 gnd 0.0028f
C3009 vdd.n194 gnd 0.002965f
C3010 vdd.n195 gnd 0.005211f
C3011 vdd.n196 gnd 0.0028f
C3012 vdd.n197 gnd 0.006618f
C3013 vdd.n198 gnd 0.002965f
C3014 vdd.n199 gnd 0.005211f
C3015 vdd.n200 gnd 0.0028f
C3016 vdd.n201 gnd 0.004963f
C3017 vdd.n202 gnd 0.004978f
C3018 vdd.t198 gnd 0.014218f
C3019 vdd.n203 gnd 0.031635f
C3020 vdd.n204 gnd 0.164637f
C3021 vdd.n205 gnd 0.0028f
C3022 vdd.n206 gnd 0.002965f
C3023 vdd.n207 gnd 0.006618f
C3024 vdd.n208 gnd 0.006618f
C3025 vdd.n209 gnd 0.002965f
C3026 vdd.n210 gnd 0.0028f
C3027 vdd.n211 gnd 0.005211f
C3028 vdd.n212 gnd 0.005211f
C3029 vdd.n213 gnd 0.0028f
C3030 vdd.n214 gnd 0.002965f
C3031 vdd.n215 gnd 0.006618f
C3032 vdd.n216 gnd 0.006618f
C3033 vdd.n217 gnd 0.002965f
C3034 vdd.n218 gnd 0.0028f
C3035 vdd.n219 gnd 0.005211f
C3036 vdd.n220 gnd 0.005211f
C3037 vdd.n221 gnd 0.0028f
C3038 vdd.n222 gnd 0.002965f
C3039 vdd.n223 gnd 0.006618f
C3040 vdd.n224 gnd 0.006618f
C3041 vdd.n225 gnd 0.015646f
C3042 vdd.n226 gnd 0.002882f
C3043 vdd.n227 gnd 0.0028f
C3044 vdd.n228 gnd 0.013467f
C3045 vdd.n229 gnd 0.009107f
C3046 vdd.n230 gnd 0.063585f
C3047 vdd.n231 gnd 0.229114f
C3048 vdd.n232 gnd 0.005615f
C3049 vdd.n233 gnd 0.005211f
C3050 vdd.n234 gnd 0.002882f
C3051 vdd.n235 gnd 0.006618f
C3052 vdd.n236 gnd 0.0028f
C3053 vdd.n237 gnd 0.002965f
C3054 vdd.n238 gnd 0.005211f
C3055 vdd.n239 gnd 0.0028f
C3056 vdd.n240 gnd 0.006618f
C3057 vdd.n241 gnd 0.002965f
C3058 vdd.n242 gnd 0.005211f
C3059 vdd.n243 gnd 0.0028f
C3060 vdd.n244 gnd 0.004963f
C3061 vdd.n245 gnd 0.004978f
C3062 vdd.t71 gnd 0.014218f
C3063 vdd.n246 gnd 0.031635f
C3064 vdd.n247 gnd 0.164637f
C3065 vdd.n248 gnd 0.0028f
C3066 vdd.n249 gnd 0.002965f
C3067 vdd.n250 gnd 0.006618f
C3068 vdd.n251 gnd 0.006618f
C3069 vdd.n252 gnd 0.002965f
C3070 vdd.n253 gnd 0.0028f
C3071 vdd.n254 gnd 0.005211f
C3072 vdd.n255 gnd 0.005211f
C3073 vdd.n256 gnd 0.0028f
C3074 vdd.n257 gnd 0.002965f
C3075 vdd.n258 gnd 0.006618f
C3076 vdd.n259 gnd 0.006618f
C3077 vdd.n260 gnd 0.002965f
C3078 vdd.n261 gnd 0.0028f
C3079 vdd.n262 gnd 0.005211f
C3080 vdd.n263 gnd 0.005211f
C3081 vdd.n264 gnd 0.0028f
C3082 vdd.n265 gnd 0.002965f
C3083 vdd.n266 gnd 0.006618f
C3084 vdd.n267 gnd 0.006618f
C3085 vdd.n268 gnd 0.015646f
C3086 vdd.n269 gnd 0.002882f
C3087 vdd.n270 gnd 0.0028f
C3088 vdd.n271 gnd 0.013467f
C3089 vdd.n272 gnd 0.009402f
C3090 vdd.t119 gnd 0.03294f
C3091 vdd.t202 gnd 0.03294f
C3092 vdd.n273 gnd 0.226387f
C3093 vdd.n274 gnd 0.178019f
C3094 vdd.t113 gnd 0.03294f
C3095 vdd.t36 gnd 0.03294f
C3096 vdd.n275 gnd 0.226387f
C3097 vdd.n276 gnd 0.14366f
C3098 vdd.t77 gnd 0.03294f
C3099 vdd.t225 gnd 0.03294f
C3100 vdd.n277 gnd 0.226387f
C3101 vdd.n278 gnd 0.14366f
C3102 vdd.t66 gnd 0.03294f
C3103 vdd.t58 gnd 0.03294f
C3104 vdd.n279 gnd 0.226387f
C3105 vdd.n280 gnd 0.14366f
C3106 vdd.t219 gnd 0.03294f
C3107 vdd.t80 gnd 0.03294f
C3108 vdd.n281 gnd 0.226387f
C3109 vdd.n282 gnd 0.14366f
C3110 vdd.t197 gnd 0.03294f
C3111 vdd.t65 gnd 0.03294f
C3112 vdd.n283 gnd 0.226387f
C3113 vdd.n284 gnd 0.14366f
C3114 vdd.t209 gnd 0.03294f
C3115 vdd.t70 gnd 0.03294f
C3116 vdd.n285 gnd 0.226387f
C3117 vdd.n286 gnd 0.14366f
C3118 vdd.t98 gnd 0.03294f
C3119 vdd.t87 gnd 0.03294f
C3120 vdd.n287 gnd 0.226387f
C3121 vdd.n288 gnd 0.14366f
C3122 vdd.t38 gnd 0.03294f
C3123 vdd.t200 gnd 0.03294f
C3124 vdd.n289 gnd 0.226387f
C3125 vdd.n290 gnd 0.14366f
C3126 vdd.n291 gnd 0.005615f
C3127 vdd.n292 gnd 0.005211f
C3128 vdd.n293 gnd 0.002882f
C3129 vdd.n294 gnd 0.006618f
C3130 vdd.n295 gnd 0.0028f
C3131 vdd.n296 gnd 0.002965f
C3132 vdd.n297 gnd 0.005211f
C3133 vdd.n298 gnd 0.0028f
C3134 vdd.n299 gnd 0.006618f
C3135 vdd.n300 gnd 0.002965f
C3136 vdd.n301 gnd 0.005211f
C3137 vdd.n302 gnd 0.0028f
C3138 vdd.n303 gnd 0.004963f
C3139 vdd.n304 gnd 0.004978f
C3140 vdd.t62 gnd 0.014218f
C3141 vdd.n305 gnd 0.031635f
C3142 vdd.n306 gnd 0.164637f
C3143 vdd.n307 gnd 0.0028f
C3144 vdd.n308 gnd 0.002965f
C3145 vdd.n309 gnd 0.006618f
C3146 vdd.n310 gnd 0.006618f
C3147 vdd.n311 gnd 0.002965f
C3148 vdd.n312 gnd 0.0028f
C3149 vdd.n313 gnd 0.005211f
C3150 vdd.n314 gnd 0.005211f
C3151 vdd.n315 gnd 0.0028f
C3152 vdd.n316 gnd 0.002965f
C3153 vdd.n317 gnd 0.006618f
C3154 vdd.n318 gnd 0.006618f
C3155 vdd.n319 gnd 0.002965f
C3156 vdd.n320 gnd 0.0028f
C3157 vdd.n321 gnd 0.005211f
C3158 vdd.n322 gnd 0.005211f
C3159 vdd.n323 gnd 0.0028f
C3160 vdd.n324 gnd 0.002965f
C3161 vdd.n325 gnd 0.006618f
C3162 vdd.n326 gnd 0.006618f
C3163 vdd.n327 gnd 0.015646f
C3164 vdd.n328 gnd 0.002882f
C3165 vdd.n329 gnd 0.0028f
C3166 vdd.n330 gnd 0.013467f
C3167 vdd.n331 gnd 0.009107f
C3168 vdd.n332 gnd 0.063585f
C3169 vdd.n333 gnd 0.262286f
C3170 vdd.n334 gnd 0.007863f
C3171 vdd.n335 gnd 0.010231f
C3172 vdd.n336 gnd 0.008235f
C3173 vdd.n337 gnd 0.008235f
C3174 vdd.n338 gnd 0.010231f
C3175 vdd.n339 gnd 0.010231f
C3176 vdd.n340 gnd 0.747604f
C3177 vdd.n341 gnd 0.010231f
C3178 vdd.n342 gnd 0.010231f
C3179 vdd.n343 gnd 0.010231f
C3180 vdd.n344 gnd 0.810339f
C3181 vdd.n345 gnd 0.010231f
C3182 vdd.n346 gnd 0.010231f
C3183 vdd.n347 gnd 0.010231f
C3184 vdd.n348 gnd 0.010231f
C3185 vdd.n349 gnd 0.008235f
C3186 vdd.n350 gnd 0.010231f
C3187 vdd.t64 gnd 0.5228f
C3188 vdd.n351 gnd 0.010231f
C3189 vdd.n352 gnd 0.010231f
C3190 vdd.n353 gnd 0.010231f
C3191 vdd.t69 gnd 0.5228f
C3192 vdd.n354 gnd 0.010231f
C3193 vdd.n355 gnd 0.010231f
C3194 vdd.n356 gnd 0.010231f
C3195 vdd.n357 gnd 0.010231f
C3196 vdd.n358 gnd 0.010231f
C3197 vdd.n359 gnd 0.008235f
C3198 vdd.n360 gnd 0.010231f
C3199 vdd.n361 gnd 0.590764f
C3200 vdd.n362 gnd 0.010231f
C3201 vdd.n363 gnd 0.010231f
C3202 vdd.n364 gnd 0.010231f
C3203 vdd.t72 gnd 0.5228f
C3204 vdd.n365 gnd 0.010231f
C3205 vdd.n366 gnd 0.010231f
C3206 vdd.n367 gnd 0.010231f
C3207 vdd.n368 gnd 0.010231f
C3208 vdd.n369 gnd 0.010231f
C3209 vdd.n370 gnd 0.008235f
C3210 vdd.n371 gnd 0.010231f
C3211 vdd.t37 gnd 0.5228f
C3212 vdd.n372 gnd 0.010231f
C3213 vdd.n373 gnd 0.010231f
C3214 vdd.n374 gnd 0.010231f
C3215 vdd.n375 gnd 0.611676f
C3216 vdd.n376 gnd 0.010231f
C3217 vdd.n377 gnd 0.010231f
C3218 vdd.n378 gnd 0.010231f
C3219 vdd.n379 gnd 0.010231f
C3220 vdd.n380 gnd 0.010231f
C3221 vdd.n381 gnd 0.008235f
C3222 vdd.n382 gnd 0.010231f
C3223 vdd.t23 gnd 0.5228f
C3224 vdd.n383 gnd 0.010231f
C3225 vdd.n384 gnd 0.010231f
C3226 vdd.n385 gnd 0.010231f
C3227 vdd.n386 gnd 0.528028f
C3228 vdd.n387 gnd 0.010231f
C3229 vdd.n388 gnd 0.010231f
C3230 vdd.n389 gnd 0.010231f
C3231 vdd.n390 gnd 0.010231f
C3232 vdd.n391 gnd 0.024751f
C3233 vdd.n392 gnd 0.025281f
C3234 vdd.t245 gnd 0.5228f
C3235 vdd.n393 gnd 0.024751f
C3236 vdd.n425 gnd 0.010231f
C3237 vdd.t273 gnd 0.125873f
C3238 vdd.t272 gnd 0.134524f
C3239 vdd.t271 gnd 0.164388f
C3240 vdd.n426 gnd 0.210723f
C3241 vdd.n427 gnd 0.177869f
C3242 vdd.n428 gnd 0.013505f
C3243 vdd.n429 gnd 0.010231f
C3244 vdd.n430 gnd 0.008235f
C3245 vdd.n431 gnd 0.010231f
C3246 vdd.n432 gnd 0.008235f
C3247 vdd.n433 gnd 0.010231f
C3248 vdd.n434 gnd 0.008235f
C3249 vdd.n435 gnd 0.010231f
C3250 vdd.n436 gnd 0.008235f
C3251 vdd.n437 gnd 0.010231f
C3252 vdd.n438 gnd 0.008235f
C3253 vdd.n439 gnd 0.010231f
C3254 vdd.t247 gnd 0.125873f
C3255 vdd.t246 gnd 0.134524f
C3256 vdd.t244 gnd 0.164388f
C3257 vdd.n440 gnd 0.210723f
C3258 vdd.n441 gnd 0.177869f
C3259 vdd.n442 gnd 0.008235f
C3260 vdd.n443 gnd 0.010231f
C3261 vdd.n444 gnd 0.008235f
C3262 vdd.n445 gnd 0.010231f
C3263 vdd.n446 gnd 0.008235f
C3264 vdd.n447 gnd 0.010231f
C3265 vdd.n448 gnd 0.008235f
C3266 vdd.n449 gnd 0.010231f
C3267 vdd.n450 gnd 0.008235f
C3268 vdd.n451 gnd 0.010231f
C3269 vdd.t253 gnd 0.125873f
C3270 vdd.t252 gnd 0.134524f
C3271 vdd.t251 gnd 0.164388f
C3272 vdd.n452 gnd 0.210723f
C3273 vdd.n453 gnd 0.177869f
C3274 vdd.n454 gnd 0.017623f
C3275 vdd.n455 gnd 0.010231f
C3276 vdd.n456 gnd 0.008235f
C3277 vdd.n457 gnd 0.010231f
C3278 vdd.n458 gnd 0.008235f
C3279 vdd.n459 gnd 0.010231f
C3280 vdd.n460 gnd 0.008235f
C3281 vdd.n461 gnd 0.010231f
C3282 vdd.n462 gnd 0.008235f
C3283 vdd.n463 gnd 0.010231f
C3284 vdd.n464 gnd 0.025281f
C3285 vdd.n465 gnd 0.006835f
C3286 vdd.n466 gnd 0.008235f
C3287 vdd.n467 gnd 0.010231f
C3288 vdd.n468 gnd 0.010231f
C3289 vdd.n469 gnd 0.008235f
C3290 vdd.n470 gnd 0.010231f
C3291 vdd.n471 gnd 0.010231f
C3292 vdd.n472 gnd 0.010231f
C3293 vdd.n473 gnd 0.010231f
C3294 vdd.n474 gnd 0.010231f
C3295 vdd.n475 gnd 0.008235f
C3296 vdd.n476 gnd 0.008235f
C3297 vdd.n477 gnd 0.010231f
C3298 vdd.n478 gnd 0.010231f
C3299 vdd.n479 gnd 0.008235f
C3300 vdd.n480 gnd 0.010231f
C3301 vdd.n481 gnd 0.010231f
C3302 vdd.n482 gnd 0.010231f
C3303 vdd.n483 gnd 0.010231f
C3304 vdd.n484 gnd 0.010231f
C3305 vdd.n485 gnd 0.008235f
C3306 vdd.n486 gnd 0.008235f
C3307 vdd.n487 gnd 0.010231f
C3308 vdd.n488 gnd 0.010231f
C3309 vdd.n489 gnd 0.008235f
C3310 vdd.n490 gnd 0.010231f
C3311 vdd.n491 gnd 0.010231f
C3312 vdd.n492 gnd 0.010231f
C3313 vdd.n493 gnd 0.010231f
C3314 vdd.n494 gnd 0.010231f
C3315 vdd.n495 gnd 0.008235f
C3316 vdd.n496 gnd 0.008235f
C3317 vdd.n497 gnd 0.010231f
C3318 vdd.n498 gnd 0.010231f
C3319 vdd.n499 gnd 0.008235f
C3320 vdd.n500 gnd 0.010231f
C3321 vdd.n501 gnd 0.010231f
C3322 vdd.n502 gnd 0.010231f
C3323 vdd.n503 gnd 0.010231f
C3324 vdd.n504 gnd 0.010231f
C3325 vdd.n505 gnd 0.008235f
C3326 vdd.n506 gnd 0.008235f
C3327 vdd.n507 gnd 0.010231f
C3328 vdd.n508 gnd 0.010231f
C3329 vdd.n509 gnd 0.006876f
C3330 vdd.n510 gnd 0.010231f
C3331 vdd.n511 gnd 0.010231f
C3332 vdd.n512 gnd 0.010231f
C3333 vdd.n513 gnd 0.010231f
C3334 vdd.n514 gnd 0.010231f
C3335 vdd.n515 gnd 0.006876f
C3336 vdd.n516 gnd 0.008235f
C3337 vdd.n517 gnd 0.010231f
C3338 vdd.n518 gnd 0.010231f
C3339 vdd.n519 gnd 0.008235f
C3340 vdd.n520 gnd 0.010231f
C3341 vdd.n521 gnd 0.010231f
C3342 vdd.n522 gnd 0.010231f
C3343 vdd.n523 gnd 0.010231f
C3344 vdd.n524 gnd 0.010231f
C3345 vdd.n525 gnd 0.008235f
C3346 vdd.n526 gnd 0.008235f
C3347 vdd.n527 gnd 0.010231f
C3348 vdd.n528 gnd 0.010231f
C3349 vdd.n529 gnd 0.008235f
C3350 vdd.n530 gnd 0.010231f
C3351 vdd.n531 gnd 0.010231f
C3352 vdd.n532 gnd 0.010231f
C3353 vdd.n533 gnd 0.010231f
C3354 vdd.n534 gnd 0.010231f
C3355 vdd.n535 gnd 0.008235f
C3356 vdd.n536 gnd 0.008235f
C3357 vdd.n537 gnd 0.010231f
C3358 vdd.n538 gnd 0.010231f
C3359 vdd.n539 gnd 0.008235f
C3360 vdd.n540 gnd 0.010231f
C3361 vdd.n541 gnd 0.010231f
C3362 vdd.n542 gnd 0.010231f
C3363 vdd.n543 gnd 0.010231f
C3364 vdd.n544 gnd 0.010231f
C3365 vdd.n545 gnd 0.008235f
C3366 vdd.n546 gnd 0.008235f
C3367 vdd.n547 gnd 0.010231f
C3368 vdd.n548 gnd 0.010231f
C3369 vdd.n549 gnd 0.008235f
C3370 vdd.n550 gnd 0.010231f
C3371 vdd.n551 gnd 0.010231f
C3372 vdd.n552 gnd 0.010231f
C3373 vdd.n553 gnd 0.010231f
C3374 vdd.n554 gnd 0.010231f
C3375 vdd.n555 gnd 0.008235f
C3376 vdd.n556 gnd 0.008235f
C3377 vdd.n557 gnd 0.010231f
C3378 vdd.n558 gnd 0.010231f
C3379 vdd.n559 gnd 0.008235f
C3380 vdd.n560 gnd 0.010231f
C3381 vdd.n561 gnd 0.010231f
C3382 vdd.n562 gnd 0.010231f
C3383 vdd.n563 gnd 0.010231f
C3384 vdd.n564 gnd 0.010231f
C3385 vdd.n565 gnd 0.0056f
C3386 vdd.n566 gnd 0.017623f
C3387 vdd.n567 gnd 0.010231f
C3388 vdd.n568 gnd 0.010231f
C3389 vdd.n569 gnd 0.008153f
C3390 vdd.n570 gnd 0.010231f
C3391 vdd.n571 gnd 0.010231f
C3392 vdd.n572 gnd 0.010231f
C3393 vdd.n573 gnd 0.010231f
C3394 vdd.n574 gnd 0.010231f
C3395 vdd.n575 gnd 0.008235f
C3396 vdd.n576 gnd 0.008235f
C3397 vdd.n577 gnd 0.010231f
C3398 vdd.n578 gnd 0.010231f
C3399 vdd.n579 gnd 0.008235f
C3400 vdd.n580 gnd 0.010231f
C3401 vdd.n581 gnd 0.010231f
C3402 vdd.n582 gnd 0.010231f
C3403 vdd.n583 gnd 0.010231f
C3404 vdd.n584 gnd 0.010231f
C3405 vdd.n585 gnd 0.008235f
C3406 vdd.n586 gnd 0.008235f
C3407 vdd.n587 gnd 0.010231f
C3408 vdd.n588 gnd 0.010231f
C3409 vdd.n589 gnd 0.008235f
C3410 vdd.n590 gnd 0.010231f
C3411 vdd.n591 gnd 0.010231f
C3412 vdd.n592 gnd 0.010231f
C3413 vdd.n593 gnd 0.010231f
C3414 vdd.n594 gnd 0.010231f
C3415 vdd.n595 gnd 0.008235f
C3416 vdd.n596 gnd 0.008235f
C3417 vdd.n597 gnd 0.010231f
C3418 vdd.n598 gnd 0.010231f
C3419 vdd.n599 gnd 0.008235f
C3420 vdd.n600 gnd 0.010231f
C3421 vdd.n601 gnd 0.010231f
C3422 vdd.n602 gnd 0.010231f
C3423 vdd.n603 gnd 0.010231f
C3424 vdd.n604 gnd 0.010231f
C3425 vdd.n605 gnd 0.008235f
C3426 vdd.n606 gnd 0.008235f
C3427 vdd.n607 gnd 0.010231f
C3428 vdd.n608 gnd 0.010231f
C3429 vdd.n609 gnd 0.008235f
C3430 vdd.n610 gnd 0.010231f
C3431 vdd.n611 gnd 0.010231f
C3432 vdd.n612 gnd 0.010231f
C3433 vdd.n613 gnd 0.010231f
C3434 vdd.n614 gnd 0.010231f
C3435 vdd.n615 gnd 0.008235f
C3436 vdd.n616 gnd 0.010231f
C3437 vdd.n617 gnd 0.008235f
C3438 vdd.n618 gnd 0.004323f
C3439 vdd.n619 gnd 0.010231f
C3440 vdd.n620 gnd 0.010231f
C3441 vdd.n621 gnd 0.008235f
C3442 vdd.n622 gnd 0.010231f
C3443 vdd.n623 gnd 0.008235f
C3444 vdd.n624 gnd 0.010231f
C3445 vdd.n625 gnd 0.008235f
C3446 vdd.n626 gnd 0.010231f
C3447 vdd.n627 gnd 0.008235f
C3448 vdd.n628 gnd 0.010231f
C3449 vdd.n629 gnd 0.008235f
C3450 vdd.n630 gnd 0.010231f
C3451 vdd.n631 gnd 0.008235f
C3452 vdd.n632 gnd 0.010231f
C3453 vdd.n633 gnd 0.569852f
C3454 vdd.t19 gnd 0.5228f
C3455 vdd.n634 gnd 0.010231f
C3456 vdd.n635 gnd 0.008235f
C3457 vdd.n636 gnd 0.010231f
C3458 vdd.n637 gnd 0.008235f
C3459 vdd.n638 gnd 0.010231f
C3460 vdd.t55 gnd 0.5228f
C3461 vdd.n639 gnd 0.010231f
C3462 vdd.n640 gnd 0.008235f
C3463 vdd.n641 gnd 0.010231f
C3464 vdd.n642 gnd 0.008235f
C3465 vdd.n643 gnd 0.010231f
C3466 vdd.t15 gnd 0.5228f
C3467 vdd.n644 gnd 0.6535f
C3468 vdd.n645 gnd 0.010231f
C3469 vdd.n646 gnd 0.008235f
C3470 vdd.n647 gnd 0.010231f
C3471 vdd.n648 gnd 0.008235f
C3472 vdd.n649 gnd 0.010231f
C3473 vdd.t76 gnd 0.5228f
C3474 vdd.n650 gnd 0.010231f
C3475 vdd.n651 gnd 0.008235f
C3476 vdd.n652 gnd 0.010231f
C3477 vdd.n653 gnd 0.008235f
C3478 vdd.n654 gnd 0.010231f
C3479 vdd.n655 gnd 0.726692f
C3480 vdd.n656 gnd 0.867847f
C3481 vdd.t2 gnd 0.5228f
C3482 vdd.n657 gnd 0.010231f
C3483 vdd.n658 gnd 0.008235f
C3484 vdd.n659 gnd 0.010231f
C3485 vdd.n660 gnd 0.008235f
C3486 vdd.n661 gnd 0.010231f
C3487 vdd.n662 gnd 0.54894f
C3488 vdd.n663 gnd 0.010231f
C3489 vdd.n664 gnd 0.008235f
C3490 vdd.n665 gnd 0.010231f
C3491 vdd.n666 gnd 0.008235f
C3492 vdd.n667 gnd 0.010231f
C3493 vdd.t116 gnd 0.5228f
C3494 vdd.t123 gnd 0.5228f
C3495 vdd.n668 gnd 0.010231f
C3496 vdd.n669 gnd 0.008235f
C3497 vdd.n670 gnd 0.010231f
C3498 vdd.n671 gnd 0.008235f
C3499 vdd.n672 gnd 0.010231f
C3500 vdd.t13 gnd 0.5228f
C3501 vdd.n673 gnd 0.010231f
C3502 vdd.n674 gnd 0.008235f
C3503 vdd.n675 gnd 0.010231f
C3504 vdd.n676 gnd 0.008235f
C3505 vdd.n677 gnd 0.010231f
C3506 vdd.n678 gnd 1.0456f
C3507 vdd.n679 gnd 0.852163f
C3508 vdd.n680 gnd 0.010231f
C3509 vdd.n681 gnd 0.008235f
C3510 vdd.n682 gnd 0.024751f
C3511 vdd.n683 gnd 0.006835f
C3512 vdd.n684 gnd 0.024751f
C3513 vdd.t258 gnd 0.5228f
C3514 vdd.n685 gnd 0.024751f
C3515 vdd.n686 gnd 0.006835f
C3516 vdd.n687 gnd 0.008799f
C3517 vdd.t259 gnd 0.125873f
C3518 vdd.t260 gnd 0.134524f
C3519 vdd.t257 gnd 0.164388f
C3520 vdd.n688 gnd 0.210723f
C3521 vdd.n689 gnd 0.177045f
C3522 vdd.n690 gnd 0.012682f
C3523 vdd.n691 gnd 0.010231f
C3524 vdd.n692 gnd 12.3485f
C3525 vdd.n723 gnd 1.4377f
C3526 vdd.n724 gnd 0.010231f
C3527 vdd.n725 gnd 0.010231f
C3528 vdd.n726 gnd 0.025281f
C3529 vdd.n727 gnd 0.008799f
C3530 vdd.n728 gnd 0.010231f
C3531 vdd.n729 gnd 0.008235f
C3532 vdd.n730 gnd 0.006548f
C3533 vdd.n731 gnd 0.042961f
C3534 vdd.n732 gnd 0.008235f
C3535 vdd.n733 gnd 0.010231f
C3536 vdd.n734 gnd 0.010231f
C3537 vdd.n735 gnd 0.010231f
C3538 vdd.n736 gnd 0.010231f
C3539 vdd.n737 gnd 0.010231f
C3540 vdd.n738 gnd 0.010231f
C3541 vdd.n739 gnd 0.010231f
C3542 vdd.n740 gnd 0.010231f
C3543 vdd.n741 gnd 0.010231f
C3544 vdd.n742 gnd 0.010231f
C3545 vdd.n743 gnd 0.010231f
C3546 vdd.n744 gnd 0.010231f
C3547 vdd.n745 gnd 0.010231f
C3548 vdd.n746 gnd 0.010231f
C3549 vdd.n747 gnd 0.006876f
C3550 vdd.n748 gnd 0.010231f
C3551 vdd.n749 gnd 0.010231f
C3552 vdd.n750 gnd 0.010231f
C3553 vdd.n751 gnd 0.010231f
C3554 vdd.n752 gnd 0.010231f
C3555 vdd.n753 gnd 0.010231f
C3556 vdd.n754 gnd 0.010231f
C3557 vdd.n755 gnd 0.010231f
C3558 vdd.n756 gnd 0.010231f
C3559 vdd.n757 gnd 0.010231f
C3560 vdd.n758 gnd 0.010231f
C3561 vdd.n759 gnd 0.010231f
C3562 vdd.n760 gnd 0.010231f
C3563 vdd.n761 gnd 0.010231f
C3564 vdd.n762 gnd 0.010231f
C3565 vdd.n763 gnd 0.010231f
C3566 vdd.n764 gnd 0.010231f
C3567 vdd.n765 gnd 0.010231f
C3568 vdd.n766 gnd 0.010231f
C3569 vdd.n767 gnd 0.008153f
C3570 vdd.t269 gnd 0.125873f
C3571 vdd.t270 gnd 0.134524f
C3572 vdd.t268 gnd 0.164388f
C3573 vdd.n768 gnd 0.210723f
C3574 vdd.n769 gnd 0.177045f
C3575 vdd.n770 gnd 0.010231f
C3576 vdd.n771 gnd 0.010231f
C3577 vdd.n772 gnd 0.010231f
C3578 vdd.n773 gnd 0.010231f
C3579 vdd.n774 gnd 0.010231f
C3580 vdd.n775 gnd 0.010231f
C3581 vdd.n776 gnd 0.010231f
C3582 vdd.n777 gnd 0.010231f
C3583 vdd.n778 gnd 0.010231f
C3584 vdd.n779 gnd 0.010231f
C3585 vdd.n780 gnd 0.010231f
C3586 vdd.n781 gnd 0.010231f
C3587 vdd.n782 gnd 0.010231f
C3588 vdd.n783 gnd 0.006548f
C3589 vdd.n785 gnd 0.006957f
C3590 vdd.n786 gnd 0.006957f
C3591 vdd.n787 gnd 0.006957f
C3592 vdd.n788 gnd 0.006957f
C3593 vdd.n789 gnd 0.006957f
C3594 vdd.n790 gnd 0.006957f
C3595 vdd.n792 gnd 0.006957f
C3596 vdd.n793 gnd 0.006957f
C3597 vdd.n795 gnd 0.006957f
C3598 vdd.n796 gnd 0.005065f
C3599 vdd.n798 gnd 0.006957f
C3600 vdd.t235 gnd 0.281145f
C3601 vdd.t234 gnd 0.287787f
C3602 vdd.t232 gnd 0.183542f
C3603 vdd.n799 gnd 0.099195f
C3604 vdd.n800 gnd 0.056266f
C3605 vdd.n801 gnd 0.009943f
C3606 vdd.n802 gnd 0.015797f
C3607 vdd.n804 gnd 0.006957f
C3608 vdd.n805 gnd 0.711008f
C3609 vdd.n806 gnd 0.014897f
C3610 vdd.n807 gnd 0.014897f
C3611 vdd.n808 gnd 0.006957f
C3612 vdd.n809 gnd 0.015797f
C3613 vdd.n810 gnd 0.006957f
C3614 vdd.n811 gnd 0.006957f
C3615 vdd.n812 gnd 0.006957f
C3616 vdd.n813 gnd 0.006957f
C3617 vdd.n814 gnd 0.006957f
C3618 vdd.n816 gnd 0.006957f
C3619 vdd.n817 gnd 0.006957f
C3620 vdd.n819 gnd 0.006957f
C3621 vdd.n820 gnd 0.006957f
C3622 vdd.n822 gnd 0.006957f
C3623 vdd.n823 gnd 0.006957f
C3624 vdd.n825 gnd 0.006957f
C3625 vdd.n826 gnd 0.006957f
C3626 vdd.n828 gnd 0.006957f
C3627 vdd.n829 gnd 0.006957f
C3628 vdd.n831 gnd 0.006957f
C3629 vdd.t256 gnd 0.281145f
C3630 vdd.t255 gnd 0.287787f
C3631 vdd.t254 gnd 0.183542f
C3632 vdd.n832 gnd 0.099195f
C3633 vdd.n833 gnd 0.056266f
C3634 vdd.n834 gnd 0.006957f
C3635 vdd.n836 gnd 0.006957f
C3636 vdd.n837 gnd 0.006957f
C3637 vdd.t233 gnd 0.355504f
C3638 vdd.n838 gnd 0.006957f
C3639 vdd.n839 gnd 0.006957f
C3640 vdd.n840 gnd 0.006957f
C3641 vdd.n841 gnd 0.006957f
C3642 vdd.n842 gnd 0.006957f
C3643 vdd.n843 gnd 0.711008f
C3644 vdd.n844 gnd 0.006957f
C3645 vdd.n845 gnd 0.006957f
C3646 vdd.n846 gnd 0.559396f
C3647 vdd.n847 gnd 0.006957f
C3648 vdd.n848 gnd 0.006957f
C3649 vdd.n849 gnd 0.006957f
C3650 vdd.n850 gnd 0.006957f
C3651 vdd.n851 gnd 0.711008f
C3652 vdd.n852 gnd 0.006957f
C3653 vdd.n853 gnd 0.006957f
C3654 vdd.n854 gnd 0.006957f
C3655 vdd.n855 gnd 0.006957f
C3656 vdd.n856 gnd 0.006957f
C3657 vdd.t155 gnd 0.355504f
C3658 vdd.n857 gnd 0.006957f
C3659 vdd.n858 gnd 0.006957f
C3660 vdd.n859 gnd 0.006957f
C3661 vdd.n860 gnd 0.006957f
C3662 vdd.n861 gnd 0.006957f
C3663 vdd.t172 gnd 0.355504f
C3664 vdd.n862 gnd 0.006957f
C3665 vdd.n863 gnd 0.006957f
C3666 vdd.n864 gnd 0.684868f
C3667 vdd.n865 gnd 0.006957f
C3668 vdd.n866 gnd 0.006957f
C3669 vdd.n867 gnd 0.006957f
C3670 vdd.t171 gnd 0.355504f
C3671 vdd.n868 gnd 0.006957f
C3672 vdd.n869 gnd 0.006957f
C3673 vdd.n870 gnd 0.528028f
C3674 vdd.n871 gnd 0.006957f
C3675 vdd.n872 gnd 0.006957f
C3676 vdd.n873 gnd 0.006957f
C3677 vdd.n874 gnd 0.49666f
C3678 vdd.n875 gnd 0.006957f
C3679 vdd.n876 gnd 0.006957f
C3680 vdd.n877 gnd 0.371188f
C3681 vdd.n878 gnd 0.006957f
C3682 vdd.n879 gnd 0.006957f
C3683 vdd.n880 gnd 0.006957f
C3684 vdd.n881 gnd 0.6535f
C3685 vdd.n882 gnd 0.006957f
C3686 vdd.n883 gnd 0.006957f
C3687 vdd.t178 gnd 0.355504f
C3688 vdd.n884 gnd 0.006957f
C3689 vdd.n885 gnd 0.006957f
C3690 vdd.n886 gnd 0.006957f
C3691 vdd.n887 gnd 0.711008f
C3692 vdd.n888 gnd 0.006957f
C3693 vdd.n889 gnd 0.006957f
C3694 vdd.t179 gnd 0.355504f
C3695 vdd.n890 gnd 0.006957f
C3696 vdd.n891 gnd 0.006957f
C3697 vdd.n892 gnd 0.006957f
C3698 vdd.t149 gnd 0.355504f
C3699 vdd.n893 gnd 0.006957f
C3700 vdd.n894 gnd 0.006957f
C3701 vdd.n895 gnd 0.006957f
C3702 vdd.t263 gnd 0.287787f
C3703 vdd.t261 gnd 0.183542f
C3704 vdd.t264 gnd 0.287787f
C3705 vdd.n896 gnd 0.161748f
C3706 vdd.n897 gnd 0.020155f
C3707 vdd.n898 gnd 0.006957f
C3708 vdd.t262 gnd 0.256172f
C3709 vdd.n899 gnd 0.006957f
C3710 vdd.n900 gnd 0.006957f
C3711 vdd.n901 gnd 0.611676f
C3712 vdd.n902 gnd 0.006957f
C3713 vdd.n903 gnd 0.006957f
C3714 vdd.n904 gnd 0.006957f
C3715 vdd.n905 gnd 0.413012f
C3716 vdd.n906 gnd 0.006957f
C3717 vdd.n907 gnd 0.006957f
C3718 vdd.t150 gnd 0.146384f
C3719 vdd.n908 gnd 0.454836f
C3720 vdd.n909 gnd 0.006957f
C3721 vdd.n910 gnd 0.006957f
C3722 vdd.n911 gnd 0.006957f
C3723 vdd.n912 gnd 0.569852f
C3724 vdd.n913 gnd 0.006957f
C3725 vdd.n914 gnd 0.006957f
C3726 vdd.t163 gnd 0.355504f
C3727 vdd.n915 gnd 0.006957f
C3728 vdd.n916 gnd 0.006957f
C3729 vdd.n917 gnd 0.006957f
C3730 vdd.t159 gnd 0.355504f
C3731 vdd.n918 gnd 0.006957f
C3732 vdd.n919 gnd 0.006957f
C3733 vdd.t182 gnd 0.355504f
C3734 vdd.n920 gnd 0.006957f
C3735 vdd.n921 gnd 0.006957f
C3736 vdd.n922 gnd 0.006957f
C3737 vdd.t141 gnd 0.240488f
C3738 vdd.n923 gnd 0.006957f
C3739 vdd.n924 gnd 0.006957f
C3740 vdd.n925 gnd 0.62736f
C3741 vdd.n926 gnd 0.006957f
C3742 vdd.n927 gnd 0.006957f
C3743 vdd.n928 gnd 0.006957f
C3744 vdd.t183 gnd 0.355504f
C3745 vdd.n929 gnd 0.006957f
C3746 vdd.n930 gnd 0.006957f
C3747 vdd.t195 gnd 0.33982f
C3748 vdd.n931 gnd 0.47052f
C3749 vdd.n932 gnd 0.006957f
C3750 vdd.n933 gnd 0.006957f
C3751 vdd.n934 gnd 0.006957f
C3752 vdd.t145 gnd 0.355504f
C3753 vdd.n935 gnd 0.006957f
C3754 vdd.n936 gnd 0.006957f
C3755 vdd.t187 gnd 0.355504f
C3756 vdd.n937 gnd 0.006957f
C3757 vdd.n938 gnd 0.006957f
C3758 vdd.n939 gnd 0.006957f
C3759 vdd.n940 gnd 0.711008f
C3760 vdd.n941 gnd 0.006957f
C3761 vdd.n942 gnd 0.006957f
C3762 vdd.t167 gnd 0.355504f
C3763 vdd.n943 gnd 0.006957f
C3764 vdd.n944 gnd 0.006957f
C3765 vdd.n945 gnd 0.006957f
C3766 vdd.n946 gnd 0.491432f
C3767 vdd.n947 gnd 0.006957f
C3768 vdd.n948 gnd 0.006957f
C3769 vdd.n949 gnd 0.006957f
C3770 vdd.n950 gnd 0.006957f
C3771 vdd.n951 gnd 0.006957f
C3772 vdd.t285 gnd 0.355504f
C3773 vdd.n952 gnd 0.006957f
C3774 vdd.n953 gnd 0.006957f
C3775 vdd.t147 gnd 0.355504f
C3776 vdd.n954 gnd 0.006957f
C3777 vdd.n955 gnd 0.014897f
C3778 vdd.n956 gnd 0.014897f
C3779 vdd.n957 gnd 0.805111f
C3780 vdd.n958 gnd 0.006957f
C3781 vdd.n959 gnd 0.006957f
C3782 vdd.t176 gnd 0.355504f
C3783 vdd.n960 gnd 0.014897f
C3784 vdd.n961 gnd 0.006957f
C3785 vdd.n962 gnd 0.006957f
C3786 vdd.t189 gnd 0.606448f
C3787 vdd.n980 gnd 0.015797f
C3788 vdd.n998 gnd 0.014897f
C3789 vdd.n999 gnd 0.006957f
C3790 vdd.n1000 gnd 0.014897f
C3791 vdd.t301 gnd 0.281145f
C3792 vdd.t300 gnd 0.287787f
C3793 vdd.t299 gnd 0.183542f
C3794 vdd.n1001 gnd 0.099195f
C3795 vdd.n1002 gnd 0.056266f
C3796 vdd.n1003 gnd 0.015797f
C3797 vdd.n1004 gnd 0.006957f
C3798 vdd.n1005 gnd 0.41824f
C3799 vdd.n1006 gnd 0.014897f
C3800 vdd.n1007 gnd 0.006957f
C3801 vdd.n1008 gnd 0.015797f
C3802 vdd.n1009 gnd 0.006957f
C3803 vdd.t280 gnd 0.281145f
C3804 vdd.t279 gnd 0.287787f
C3805 vdd.t277 gnd 0.183542f
C3806 vdd.n1010 gnd 0.099195f
C3807 vdd.n1011 gnd 0.056266f
C3808 vdd.n1012 gnd 0.009943f
C3809 vdd.n1013 gnd 0.006957f
C3810 vdd.n1014 gnd 0.006957f
C3811 vdd.t278 gnd 0.355504f
C3812 vdd.n1015 gnd 0.006957f
C3813 vdd.t191 gnd 0.355504f
C3814 vdd.n1016 gnd 0.006957f
C3815 vdd.n1017 gnd 0.006957f
C3816 vdd.n1018 gnd 0.006957f
C3817 vdd.n1019 gnd 0.006957f
C3818 vdd.n1020 gnd 0.006957f
C3819 vdd.n1021 gnd 0.711008f
C3820 vdd.n1022 gnd 0.006957f
C3821 vdd.n1023 gnd 0.006957f
C3822 vdd.t161 gnd 0.355504f
C3823 vdd.n1024 gnd 0.006957f
C3824 vdd.n1025 gnd 0.006957f
C3825 vdd.n1026 gnd 0.006957f
C3826 vdd.n1027 gnd 0.006957f
C3827 vdd.n1028 gnd 0.512344f
C3828 vdd.n1029 gnd 0.006957f
C3829 vdd.n1030 gnd 0.006957f
C3830 vdd.n1031 gnd 0.006957f
C3831 vdd.n1032 gnd 0.006957f
C3832 vdd.n1033 gnd 0.006957f
C3833 vdd.t142 gnd 0.355504f
C3834 vdd.n1034 gnd 0.006957f
C3835 vdd.n1035 gnd 0.006957f
C3836 vdd.t180 gnd 0.355504f
C3837 vdd.n1036 gnd 0.006957f
C3838 vdd.n1037 gnd 0.006957f
C3839 vdd.n1038 gnd 0.006957f
C3840 vdd.t166 gnd 0.355504f
C3841 vdd.n1039 gnd 0.006957f
C3842 vdd.n1040 gnd 0.006957f
C3843 vdd.t143 gnd 0.355504f
C3844 vdd.n1041 gnd 0.006957f
C3845 vdd.n1042 gnd 0.006957f
C3846 vdd.n1043 gnd 0.006957f
C3847 vdd.t164 gnd 0.33982f
C3848 vdd.n1044 gnd 0.006957f
C3849 vdd.n1045 gnd 0.006957f
C3850 vdd.n1046 gnd 0.528028f
C3851 vdd.n1047 gnd 0.006957f
C3852 vdd.n1048 gnd 0.006957f
C3853 vdd.n1049 gnd 0.006957f
C3854 vdd.t184 gnd 0.355504f
C3855 vdd.n1050 gnd 0.006957f
C3856 vdd.n1051 gnd 0.006957f
C3857 vdd.t152 gnd 0.240488f
C3858 vdd.n1052 gnd 0.371188f
C3859 vdd.n1053 gnd 0.006957f
C3860 vdd.n1054 gnd 0.006957f
C3861 vdd.n1055 gnd 0.006957f
C3862 vdd.n1056 gnd 0.6535f
C3863 vdd.n1057 gnd 0.006957f
C3864 vdd.n1058 gnd 0.006957f
C3865 vdd.t193 gnd 0.355504f
C3866 vdd.n1059 gnd 0.006957f
C3867 vdd.n1060 gnd 0.006957f
C3868 vdd.n1061 gnd 0.006957f
C3869 vdd.n1062 gnd 0.711008f
C3870 vdd.n1063 gnd 0.006957f
C3871 vdd.n1064 gnd 0.006957f
C3872 vdd.t158 gnd 0.355504f
C3873 vdd.n1065 gnd 0.006957f
C3874 vdd.n1066 gnd 0.006957f
C3875 vdd.n1067 gnd 0.006957f
C3876 vdd.t151 gnd 0.146384f
C3877 vdd.n1068 gnd 0.006957f
C3878 vdd.n1069 gnd 0.006957f
C3879 vdd.n1070 gnd 0.006957f
C3880 vdd.t290 gnd 0.287787f
C3881 vdd.t288 gnd 0.183542f
C3882 vdd.t291 gnd 0.287787f
C3883 vdd.n1071 gnd 0.161748f
C3884 vdd.n1072 gnd 0.006957f
C3885 vdd.n1073 gnd 0.006957f
C3886 vdd.t173 gnd 0.355504f
C3887 vdd.n1074 gnd 0.006957f
C3888 vdd.n1075 gnd 0.006957f
C3889 vdd.t289 gnd 0.256172f
C3890 vdd.n1076 gnd 0.564624f
C3891 vdd.n1077 gnd 0.006957f
C3892 vdd.n1078 gnd 0.006957f
C3893 vdd.n1079 gnd 0.006957f
C3894 vdd.n1080 gnd 0.413012f
C3895 vdd.n1081 gnd 0.006957f
C3896 vdd.n1082 gnd 0.006957f
C3897 vdd.n1083 gnd 0.454836f
C3898 vdd.n1084 gnd 0.006957f
C3899 vdd.n1085 gnd 0.006957f
C3900 vdd.n1086 gnd 0.006957f
C3901 vdd.n1087 gnd 0.569852f
C3902 vdd.n1088 gnd 0.006957f
C3903 vdd.n1089 gnd 0.006957f
C3904 vdd.t153 gnd 0.355504f
C3905 vdd.n1090 gnd 0.006957f
C3906 vdd.n1091 gnd 0.006957f
C3907 vdd.n1092 gnd 0.006957f
C3908 vdd.n1093 gnd 0.711008f
C3909 vdd.n1094 gnd 0.006957f
C3910 vdd.n1095 gnd 0.006957f
C3911 vdd.t154 gnd 0.355504f
C3912 vdd.n1096 gnd 0.006957f
C3913 vdd.n1097 gnd 0.006957f
C3914 vdd.n1098 gnd 0.006957f
C3915 vdd.t194 gnd 0.355504f
C3916 vdd.n1099 gnd 0.006957f
C3917 vdd.n1100 gnd 0.006957f
C3918 vdd.n1101 gnd 0.006957f
C3919 vdd.n1102 gnd 0.006957f
C3920 vdd.n1103 gnd 0.006957f
C3921 vdd.t186 gnd 0.355504f
C3922 vdd.n1104 gnd 0.006957f
C3923 vdd.n1105 gnd 0.006957f
C3924 vdd.n1106 gnd 0.695324f
C3925 vdd.n1107 gnd 0.006957f
C3926 vdd.n1108 gnd 0.006957f
C3927 vdd.n1109 gnd 0.006957f
C3928 vdd.t146 gnd 0.355504f
C3929 vdd.n1110 gnd 0.006957f
C3930 vdd.n1111 gnd 0.006957f
C3931 vdd.n1112 gnd 0.538484f
C3932 vdd.n1113 gnd 0.006957f
C3933 vdd.n1114 gnd 0.006957f
C3934 vdd.n1115 gnd 0.006957f
C3935 vdd.n1116 gnd 0.711008f
C3936 vdd.n1117 gnd 0.006957f
C3937 vdd.n1118 gnd 0.006957f
C3938 vdd.n1119 gnd 0.381644f
C3939 vdd.n1120 gnd 0.006957f
C3940 vdd.n1121 gnd 0.006957f
C3941 vdd.n1122 gnd 0.006957f
C3942 vdd.n1123 gnd 0.711008f
C3943 vdd.n1124 gnd 0.006957f
C3944 vdd.n1125 gnd 0.006957f
C3945 vdd.n1126 gnd 0.006957f
C3946 vdd.n1127 gnd 0.006957f
C3947 vdd.n1128 gnd 0.006957f
C3948 vdd.t237 gnd 0.355504f
C3949 vdd.n1129 gnd 0.006957f
C3950 vdd.n1130 gnd 0.006957f
C3951 vdd.n1131 gnd 0.006957f
C3952 vdd.n1132 gnd 0.014897f
C3953 vdd.n1133 gnd 0.014897f
C3954 vdd.n1134 gnd 0.961951f
C3955 vdd.n1135 gnd 0.006957f
C3956 vdd.n1136 gnd 0.006957f
C3957 vdd.n1137 gnd 0.507116f
C3958 vdd.n1138 gnd 0.014897f
C3959 vdd.n1139 gnd 0.006957f
C3960 vdd.n1140 gnd 0.006957f
C3961 vdd.n1141 gnd 12.7668f
C3962 vdd.n1175 gnd 0.015797f
C3963 vdd.n1176 gnd 0.006957f
C3964 vdd.n1177 gnd 0.006957f
C3965 vdd.n1178 gnd 0.006548f
C3966 vdd.n1181 gnd 0.025281f
C3967 vdd.n1182 gnd 0.006835f
C3968 vdd.n1183 gnd 0.008235f
C3969 vdd.n1185 gnd 0.010231f
C3970 vdd.n1186 gnd 0.010231f
C3971 vdd.n1187 gnd 0.008235f
C3972 vdd.n1189 gnd 0.010231f
C3973 vdd.n1190 gnd 0.010231f
C3974 vdd.n1191 gnd 0.010231f
C3975 vdd.n1192 gnd 0.010231f
C3976 vdd.n1193 gnd 0.010231f
C3977 vdd.n1194 gnd 0.008235f
C3978 vdd.n1196 gnd 0.010231f
C3979 vdd.n1197 gnd 0.010231f
C3980 vdd.n1198 gnd 0.010231f
C3981 vdd.n1199 gnd 0.010231f
C3982 vdd.n1200 gnd 0.010231f
C3983 vdd.n1201 gnd 0.008235f
C3984 vdd.n1203 gnd 0.010231f
C3985 vdd.n1204 gnd 0.010231f
C3986 vdd.n1205 gnd 0.010231f
C3987 vdd.n1206 gnd 0.010231f
C3988 vdd.n1207 gnd 0.006876f
C3989 vdd.t250 gnd 0.125873f
C3990 vdd.t249 gnd 0.134524f
C3991 vdd.t248 gnd 0.164388f
C3992 vdd.n1208 gnd 0.210723f
C3993 vdd.n1209 gnd 0.177045f
C3994 vdd.n1211 gnd 0.010231f
C3995 vdd.n1212 gnd 0.010231f
C3996 vdd.n1213 gnd 0.008235f
C3997 vdd.n1214 gnd 0.010231f
C3998 vdd.n1216 gnd 0.010231f
C3999 vdd.n1217 gnd 0.010231f
C4000 vdd.n1218 gnd 0.010231f
C4001 vdd.n1219 gnd 0.010231f
C4002 vdd.n1220 gnd 0.008235f
C4003 vdd.n1222 gnd 0.010231f
C4004 vdd.n1223 gnd 0.010231f
C4005 vdd.n1224 gnd 0.010231f
C4006 vdd.n1225 gnd 0.010231f
C4007 vdd.n1226 gnd 0.010231f
C4008 vdd.n1227 gnd 0.008235f
C4009 vdd.n1229 gnd 0.010231f
C4010 vdd.n1230 gnd 0.010231f
C4011 vdd.n1231 gnd 0.010231f
C4012 vdd.n1232 gnd 0.010231f
C4013 vdd.n1233 gnd 0.010231f
C4014 vdd.n1234 gnd 0.008235f
C4015 vdd.n1236 gnd 0.010231f
C4016 vdd.n1237 gnd 0.010231f
C4017 vdd.n1238 gnd 0.010231f
C4018 vdd.n1239 gnd 0.010231f
C4019 vdd.n1240 gnd 0.010231f
C4020 vdd.n1241 gnd 0.008235f
C4021 vdd.n1243 gnd 0.010231f
C4022 vdd.n1244 gnd 0.010231f
C4023 vdd.n1245 gnd 0.010231f
C4024 vdd.n1246 gnd 0.010231f
C4025 vdd.n1247 gnd 0.008153f
C4026 vdd.t243 gnd 0.125873f
C4027 vdd.t242 gnd 0.134524f
C4028 vdd.t240 gnd 0.164388f
C4029 vdd.n1248 gnd 0.210723f
C4030 vdd.n1249 gnd 0.177045f
C4031 vdd.n1251 gnd 0.010231f
C4032 vdd.n1252 gnd 0.010231f
C4033 vdd.n1253 gnd 0.008235f
C4034 vdd.n1254 gnd 0.010231f
C4035 vdd.n1256 gnd 0.010231f
C4036 vdd.n1257 gnd 0.010231f
C4037 vdd.n1258 gnd 0.010231f
C4038 vdd.n1259 gnd 0.010231f
C4039 vdd.n1260 gnd 0.008235f
C4040 vdd.n1262 gnd 0.010231f
C4041 vdd.n1263 gnd 0.010231f
C4042 vdd.n1264 gnd 0.010231f
C4043 vdd.n1265 gnd 0.010231f
C4044 vdd.n1266 gnd 0.010231f
C4045 vdd.n1267 gnd 0.008235f
C4046 vdd.n1269 gnd 0.010231f
C4047 vdd.n1270 gnd 0.010231f
C4048 vdd.n1271 gnd 0.010231f
C4049 vdd.n1272 gnd 0.010231f
C4050 vdd.n1273 gnd 0.010231f
C4051 vdd.n1274 gnd 0.008235f
C4052 vdd.n1276 gnd 0.010231f
C4053 vdd.n1277 gnd 0.010231f
C4054 vdd.n1278 gnd 0.006548f
C4055 vdd.n1279 gnd 0.008235f
C4056 vdd.n1280 gnd 0.015797f
C4057 vdd.n1281 gnd 0.015797f
C4058 vdd.n1282 gnd 0.006957f
C4059 vdd.n1283 gnd 0.006957f
C4060 vdd.n1284 gnd 0.006957f
C4061 vdd.n1285 gnd 0.006957f
C4062 vdd.n1286 gnd 0.006957f
C4063 vdd.n1287 gnd 0.006957f
C4064 vdd.n1288 gnd 0.006957f
C4065 vdd.n1289 gnd 0.006957f
C4066 vdd.n1290 gnd 0.006957f
C4067 vdd.n1291 gnd 0.006957f
C4068 vdd.n1292 gnd 0.006957f
C4069 vdd.n1293 gnd 0.006957f
C4070 vdd.n1294 gnd 0.006957f
C4071 vdd.n1295 gnd 0.006957f
C4072 vdd.n1296 gnd 0.006957f
C4073 vdd.n1297 gnd 0.006957f
C4074 vdd.n1298 gnd 0.006957f
C4075 vdd.n1299 gnd 0.006957f
C4076 vdd.n1300 gnd 0.006957f
C4077 vdd.n1301 gnd 0.006957f
C4078 vdd.n1302 gnd 0.006957f
C4079 vdd.n1303 gnd 0.006957f
C4080 vdd.n1304 gnd 0.006957f
C4081 vdd.n1305 gnd 0.006957f
C4082 vdd.n1306 gnd 0.006957f
C4083 vdd.n1307 gnd 0.006957f
C4084 vdd.n1308 gnd 0.006957f
C4085 vdd.n1309 gnd 0.006957f
C4086 vdd.n1310 gnd 0.006957f
C4087 vdd.n1311 gnd 0.006957f
C4088 vdd.n1312 gnd 0.006957f
C4089 vdd.n1313 gnd 0.006957f
C4090 vdd.n1314 gnd 0.006957f
C4091 vdd.t238 gnd 0.281145f
C4092 vdd.t239 gnd 0.287787f
C4093 vdd.t236 gnd 0.183542f
C4094 vdd.n1315 gnd 0.099195f
C4095 vdd.n1316 gnd 0.056266f
C4096 vdd.n1317 gnd 0.009943f
C4097 vdd.n1318 gnd 0.006957f
C4098 vdd.t275 gnd 0.281145f
C4099 vdd.t276 gnd 0.287787f
C4100 vdd.t274 gnd 0.183542f
C4101 vdd.n1319 gnd 0.099195f
C4102 vdd.n1320 gnd 0.056266f
C4103 vdd.n1321 gnd 0.006957f
C4104 vdd.n1322 gnd 0.006957f
C4105 vdd.n1323 gnd 0.006957f
C4106 vdd.n1324 gnd 0.006957f
C4107 vdd.n1325 gnd 0.006957f
C4108 vdd.n1326 gnd 0.006957f
C4109 vdd.n1327 gnd 0.006957f
C4110 vdd.n1328 gnd 0.006957f
C4111 vdd.n1329 gnd 0.006957f
C4112 vdd.n1330 gnd 0.006957f
C4113 vdd.n1331 gnd 0.006957f
C4114 vdd.n1332 gnd 0.006957f
C4115 vdd.n1333 gnd 0.006957f
C4116 vdd.n1334 gnd 0.006957f
C4117 vdd.n1335 gnd 0.006957f
C4118 vdd.n1336 gnd 0.006957f
C4119 vdd.n1337 gnd 0.006957f
C4120 vdd.n1338 gnd 0.006957f
C4121 vdd.n1339 gnd 0.006957f
C4122 vdd.n1340 gnd 0.006957f
C4123 vdd.n1341 gnd 0.006957f
C4124 vdd.n1342 gnd 0.006957f
C4125 vdd.n1343 gnd 0.006957f
C4126 vdd.n1344 gnd 0.006957f
C4127 vdd.n1345 gnd 0.006957f
C4128 vdd.n1346 gnd 0.006957f
C4129 vdd.n1347 gnd 0.005065f
C4130 vdd.n1348 gnd 0.009943f
C4131 vdd.n1349 gnd 0.005371f
C4132 vdd.n1350 gnd 0.006957f
C4133 vdd.n1351 gnd 0.006957f
C4134 vdd.n1352 gnd 0.006957f
C4135 vdd.n1353 gnd 0.015797f
C4136 vdd.n1354 gnd 0.015797f
C4137 vdd.n1355 gnd 0.014897f
C4138 vdd.n1356 gnd 0.014897f
C4139 vdd.n1357 gnd 0.006957f
C4140 vdd.n1358 gnd 0.006957f
C4141 vdd.n1359 gnd 0.006957f
C4142 vdd.n1360 gnd 0.006957f
C4143 vdd.n1361 gnd 0.006957f
C4144 vdd.n1362 gnd 0.006957f
C4145 vdd.n1363 gnd 0.006957f
C4146 vdd.n1364 gnd 0.006957f
C4147 vdd.n1365 gnd 0.006957f
C4148 vdd.n1366 gnd 0.006957f
C4149 vdd.n1367 gnd 0.006957f
C4150 vdd.n1368 gnd 0.006957f
C4151 vdd.n1369 gnd 0.006957f
C4152 vdd.n1370 gnd 0.006957f
C4153 vdd.n1371 gnd 0.006957f
C4154 vdd.n1372 gnd 0.006957f
C4155 vdd.n1373 gnd 0.006957f
C4156 vdd.n1374 gnd 0.006957f
C4157 vdd.n1375 gnd 0.006957f
C4158 vdd.n1376 gnd 0.006957f
C4159 vdd.n1377 gnd 0.006957f
C4160 vdd.n1378 gnd 0.006957f
C4161 vdd.n1379 gnd 0.006957f
C4162 vdd.n1380 gnd 0.006957f
C4163 vdd.n1381 gnd 0.006957f
C4164 vdd.n1382 gnd 0.006957f
C4165 vdd.n1383 gnd 0.006957f
C4166 vdd.n1384 gnd 0.006957f
C4167 vdd.n1385 gnd 0.006957f
C4168 vdd.n1386 gnd 0.006957f
C4169 vdd.n1387 gnd 0.006957f
C4170 vdd.n1388 gnd 0.006957f
C4171 vdd.n1389 gnd 0.006957f
C4172 vdd.n1390 gnd 0.006957f
C4173 vdd.n1391 gnd 0.006957f
C4174 vdd.n1392 gnd 0.006957f
C4175 vdd.n1393 gnd 0.006957f
C4176 vdd.n1394 gnd 0.006957f
C4177 vdd.n1395 gnd 0.006957f
C4178 vdd.n1396 gnd 0.006957f
C4179 vdd.n1397 gnd 0.006957f
C4180 vdd.n1398 gnd 0.006957f
C4181 vdd.n1399 gnd 0.423468f
C4182 vdd.n1400 gnd 0.006957f
C4183 vdd.n1401 gnd 0.006957f
C4184 vdd.n1402 gnd 0.006957f
C4185 vdd.n1403 gnd 0.006957f
C4186 vdd.n1404 gnd 0.006957f
C4187 vdd.n1405 gnd 0.006957f
C4188 vdd.n1406 gnd 0.006957f
C4189 vdd.n1407 gnd 0.006957f
C4190 vdd.n1408 gnd 0.006957f
C4191 vdd.n1409 gnd 0.006957f
C4192 vdd.n1410 gnd 0.006957f
C4193 vdd.n1411 gnd 0.006957f
C4194 vdd.n1412 gnd 0.006957f
C4195 vdd.n1413 gnd 0.006957f
C4196 vdd.n1414 gnd 0.006957f
C4197 vdd.n1415 gnd 0.006957f
C4198 vdd.n1416 gnd 0.006957f
C4199 vdd.n1417 gnd 0.006957f
C4200 vdd.n1418 gnd 0.006957f
C4201 vdd.n1419 gnd 0.006957f
C4202 vdd.n1420 gnd 0.006957f
C4203 vdd.n1421 gnd 0.006957f
C4204 vdd.n1422 gnd 0.006957f
C4205 vdd.n1423 gnd 0.006957f
C4206 vdd.n1424 gnd 0.006957f
C4207 vdd.n1425 gnd 0.643044f
C4208 vdd.n1426 gnd 0.006957f
C4209 vdd.n1427 gnd 0.006957f
C4210 vdd.n1428 gnd 0.006957f
C4211 vdd.n1429 gnd 0.006957f
C4212 vdd.n1430 gnd 0.006957f
C4213 vdd.n1431 gnd 0.006957f
C4214 vdd.n1432 gnd 0.006957f
C4215 vdd.n1433 gnd 0.006957f
C4216 vdd.n1434 gnd 0.006957f
C4217 vdd.n1435 gnd 0.006957f
C4218 vdd.n1436 gnd 0.006957f
C4219 vdd.n1437 gnd 0.224804f
C4220 vdd.n1438 gnd 0.006957f
C4221 vdd.n1439 gnd 0.006957f
C4222 vdd.n1440 gnd 0.006957f
C4223 vdd.n1441 gnd 0.006957f
C4224 vdd.n1442 gnd 0.006957f
C4225 vdd.n1443 gnd 0.006957f
C4226 vdd.n1444 gnd 0.006957f
C4227 vdd.n1445 gnd 0.006957f
C4228 vdd.n1446 gnd 0.006957f
C4229 vdd.n1447 gnd 0.006957f
C4230 vdd.n1448 gnd 0.006957f
C4231 vdd.n1449 gnd 0.006957f
C4232 vdd.n1450 gnd 0.006957f
C4233 vdd.n1451 gnd 0.006957f
C4234 vdd.n1452 gnd 0.006957f
C4235 vdd.n1453 gnd 0.006957f
C4236 vdd.n1454 gnd 0.006957f
C4237 vdd.n1455 gnd 0.006957f
C4238 vdd.n1456 gnd 0.006957f
C4239 vdd.n1457 gnd 0.006957f
C4240 vdd.n1458 gnd 0.006957f
C4241 vdd.n1459 gnd 0.006957f
C4242 vdd.n1460 gnd 0.006957f
C4243 vdd.n1461 gnd 0.006957f
C4244 vdd.n1462 gnd 0.006957f
C4245 vdd.n1463 gnd 0.006957f
C4246 vdd.n1464 gnd 0.006957f
C4247 vdd.n1465 gnd 0.006957f
C4248 vdd.n1466 gnd 0.006957f
C4249 vdd.n1467 gnd 0.006957f
C4250 vdd.n1468 gnd 0.006957f
C4251 vdd.n1469 gnd 0.006957f
C4252 vdd.n1470 gnd 0.006957f
C4253 vdd.n1471 gnd 0.006957f
C4254 vdd.n1472 gnd 0.006957f
C4255 vdd.n1473 gnd 0.006957f
C4256 vdd.n1474 gnd 0.006957f
C4257 vdd.n1475 gnd 0.006957f
C4258 vdd.n1476 gnd 0.006957f
C4259 vdd.n1477 gnd 0.006957f
C4260 vdd.n1478 gnd 0.006957f
C4261 vdd.n1479 gnd 0.006957f
C4262 vdd.n1480 gnd 0.014897f
C4263 vdd.n1481 gnd 0.014897f
C4264 vdd.n1482 gnd 0.015797f
C4265 vdd.n1483 gnd 0.006957f
C4266 vdd.n1484 gnd 0.006957f
C4267 vdd.n1485 gnd 0.005371f
C4268 vdd.n1486 gnd 0.006957f
C4269 vdd.n1487 gnd 0.006957f
C4270 vdd.n1488 gnd 0.005065f
C4271 vdd.n1489 gnd 0.006957f
C4272 vdd.n1490 gnd 0.006957f
C4273 vdd.n1491 gnd 0.006957f
C4274 vdd.n1492 gnd 0.006957f
C4275 vdd.n1493 gnd 0.006957f
C4276 vdd.n1494 gnd 0.006957f
C4277 vdd.n1495 gnd 0.006957f
C4278 vdd.n1496 gnd 0.006957f
C4279 vdd.n1497 gnd 0.006957f
C4280 vdd.n1498 gnd 0.006957f
C4281 vdd.n1499 gnd 0.006957f
C4282 vdd.n1500 gnd 0.006957f
C4283 vdd.n1501 gnd 0.006957f
C4284 vdd.n1502 gnd 0.006957f
C4285 vdd.n1503 gnd 0.006957f
C4286 vdd.n1504 gnd 0.006957f
C4287 vdd.n1505 gnd 0.006957f
C4288 vdd.n1506 gnd 0.006957f
C4289 vdd.n1507 gnd 0.006957f
C4290 vdd.n1508 gnd 0.006957f
C4291 vdd.n1509 gnd 0.006957f
C4292 vdd.n1510 gnd 0.006957f
C4293 vdd.n1511 gnd 0.006957f
C4294 vdd.n1512 gnd 0.006957f
C4295 vdd.n1513 gnd 0.006957f
C4296 vdd.n1514 gnd 0.006957f
C4297 vdd.n1515 gnd 0.046868f
C4298 vdd.n1517 gnd 0.025281f
C4299 vdd.n1518 gnd 0.008235f
C4300 vdd.n1520 gnd 0.010231f
C4301 vdd.n1521 gnd 0.008235f
C4302 vdd.n1522 gnd 0.010231f
C4303 vdd.n1524 gnd 0.010231f
C4304 vdd.n1525 gnd 0.010231f
C4305 vdd.n1527 gnd 0.010231f
C4306 vdd.n1528 gnd 0.006835f
C4307 vdd.t241 gnd 0.5228f
C4308 vdd.n1529 gnd 0.010231f
C4309 vdd.n1530 gnd 0.025281f
C4310 vdd.n1531 gnd 0.008235f
C4311 vdd.n1532 gnd 0.010231f
C4312 vdd.n1533 gnd 0.008235f
C4313 vdd.n1534 gnd 0.010231f
C4314 vdd.n1535 gnd 1.0456f
C4315 vdd.n1536 gnd 0.010231f
C4316 vdd.n1537 gnd 0.008235f
C4317 vdd.n1538 gnd 0.008235f
C4318 vdd.n1539 gnd 0.010231f
C4319 vdd.n1540 gnd 0.008235f
C4320 vdd.n1541 gnd 0.010231f
C4321 vdd.t34 gnd 0.5228f
C4322 vdd.n1542 gnd 0.010231f
C4323 vdd.n1543 gnd 0.008235f
C4324 vdd.n1544 gnd 0.010231f
C4325 vdd.n1545 gnd 0.008235f
C4326 vdd.n1546 gnd 0.010231f
C4327 vdd.t204 gnd 0.5228f
C4328 vdd.n1547 gnd 0.010231f
C4329 vdd.n1548 gnd 0.008235f
C4330 vdd.n1549 gnd 0.010231f
C4331 vdd.n1550 gnd 0.008235f
C4332 vdd.n1551 gnd 0.010231f
C4333 vdd.n1552 gnd 0.841707f
C4334 vdd.n1553 gnd 0.867847f
C4335 vdd.t91 gnd 0.5228f
C4336 vdd.n1554 gnd 0.010231f
C4337 vdd.n1555 gnd 0.008235f
C4338 vdd.n1556 gnd 0.010231f
C4339 vdd.n1557 gnd 0.008235f
C4340 vdd.n1558 gnd 0.010231f
C4341 vdd.n1559 gnd 0.663956f
C4342 vdd.n1560 gnd 0.010231f
C4343 vdd.n1561 gnd 0.008235f
C4344 vdd.n1562 gnd 0.010231f
C4345 vdd.n1563 gnd 0.008235f
C4346 vdd.n1564 gnd 0.010231f
C4347 vdd.t99 gnd 0.5228f
C4348 vdd.t0 gnd 0.5228f
C4349 vdd.n1565 gnd 0.010231f
C4350 vdd.n1566 gnd 0.008235f
C4351 vdd.n1567 gnd 0.010231f
C4352 vdd.n1568 gnd 0.008235f
C4353 vdd.n1569 gnd 0.010231f
C4354 vdd.t59 gnd 0.5228f
C4355 vdd.n1570 gnd 0.010231f
C4356 vdd.n1571 gnd 0.008235f
C4357 vdd.n1572 gnd 0.010231f
C4358 vdd.n1573 gnd 0.008235f
C4359 vdd.n1574 gnd 0.010231f
C4360 vdd.t11 gnd 0.5228f
C4361 vdd.n1575 gnd 0.737148f
C4362 vdd.n1576 gnd 0.010231f
C4363 vdd.n1577 gnd 0.008235f
C4364 vdd.n1578 gnd 0.010231f
C4365 vdd.n1579 gnd 0.008235f
C4366 vdd.n1580 gnd 0.010231f
C4367 vdd.n1581 gnd 0.820795f
C4368 vdd.n1582 gnd 0.010231f
C4369 vdd.n1583 gnd 0.008235f
C4370 vdd.n1584 gnd 0.010231f
C4371 vdd.n1585 gnd 0.008235f
C4372 vdd.n1586 gnd 0.010231f
C4373 vdd.n1587 gnd 0.643044f
C4374 vdd.t17 gnd 0.5228f
C4375 vdd.n1588 gnd 0.010231f
C4376 vdd.n1589 gnd 0.008235f
C4377 vdd.n1590 gnd 0.010231f
C4378 vdd.n1591 gnd 0.008235f
C4379 vdd.n1592 gnd 0.010231f
C4380 vdd.t43 gnd 0.5228f
C4381 vdd.n1593 gnd 0.010231f
C4382 vdd.n1594 gnd 0.008235f
C4383 vdd.n1595 gnd 0.010231f
C4384 vdd.n1596 gnd 0.008235f
C4385 vdd.n1597 gnd 0.010231f
C4386 vdd.t131 gnd 0.5228f
C4387 vdd.n1598 gnd 0.580308f
C4388 vdd.n1599 gnd 0.010231f
C4389 vdd.n1600 gnd 0.008235f
C4390 vdd.n1601 gnd 0.010231f
C4391 vdd.n1602 gnd 0.008235f
C4392 vdd.n1603 gnd 0.010231f
C4393 vdd.t114 gnd 0.5228f
C4394 vdd.n1604 gnd 0.010231f
C4395 vdd.n1605 gnd 0.008235f
C4396 vdd.n1606 gnd 0.010231f
C4397 vdd.n1607 gnd 0.008235f
C4398 vdd.n1608 gnd 0.010231f
C4399 vdd.n1609 gnd 0.799883f
C4400 vdd.n1610 gnd 0.867847f
C4401 vdd.t51 gnd 0.5228f
C4402 vdd.n1611 gnd 0.010231f
C4403 vdd.n1612 gnd 0.008235f
C4404 vdd.n1613 gnd 0.010231f
C4405 vdd.n1614 gnd 0.008235f
C4406 vdd.n1615 gnd 0.010231f
C4407 vdd.n1616 gnd 0.622132f
C4408 vdd.n1617 gnd 0.010231f
C4409 vdd.n1618 gnd 0.008235f
C4410 vdd.n1619 gnd 0.010231f
C4411 vdd.n1620 gnd 0.008235f
C4412 vdd.n1621 gnd 0.010231f
C4413 vdd.t85 gnd 0.5228f
C4414 vdd.t67 gnd 0.5228f
C4415 vdd.n1622 gnd 0.010231f
C4416 vdd.n1623 gnd 0.008235f
C4417 vdd.n1624 gnd 0.010231f
C4418 vdd.n1625 gnd 0.008235f
C4419 vdd.n1626 gnd 0.010231f
C4420 vdd.t32 gnd 0.5228f
C4421 vdd.n1627 gnd 0.010231f
C4422 vdd.n1628 gnd 0.008235f
C4423 vdd.n1629 gnd 0.010231f
C4424 vdd.n1630 gnd 0.008235f
C4425 vdd.n1631 gnd 0.010231f
C4426 vdd.t21 gnd 0.5228f
C4427 vdd.n1632 gnd 0.778971f
C4428 vdd.n1633 gnd 0.010231f
C4429 vdd.n1634 gnd 0.008235f
C4430 vdd.n1635 gnd 0.010231f
C4431 vdd.n1636 gnd 0.008235f
C4432 vdd.n1637 gnd 0.010231f
C4433 vdd.n1638 gnd 1.0456f
C4434 vdd.n1639 gnd 0.010231f
C4435 vdd.n1640 gnd 0.008235f
C4436 vdd.n1641 gnd 0.024751f
C4437 vdd.n1642 gnd 0.006835f
C4438 vdd.n1643 gnd 0.024751f
C4439 vdd.t296 gnd 0.5228f
C4440 vdd.n1644 gnd 0.024751f
C4441 vdd.n1645 gnd 0.006835f
C4442 vdd.n1646 gnd 0.010231f
C4443 vdd.n1647 gnd 0.008235f
C4444 vdd.n1648 gnd 0.010231f
C4445 vdd.n1679 gnd 0.025281f
C4446 vdd.n1680 gnd 1.54226f
C4447 vdd.n1681 gnd 0.010231f
C4448 vdd.n1682 gnd 0.008235f
C4449 vdd.n1683 gnd 0.010231f
C4450 vdd.n1684 gnd 0.010231f
C4451 vdd.n1685 gnd 0.010231f
C4452 vdd.n1686 gnd 0.010231f
C4453 vdd.n1687 gnd 0.010231f
C4454 vdd.n1688 gnd 0.008235f
C4455 vdd.n1689 gnd 0.010231f
C4456 vdd.n1690 gnd 0.010231f
C4457 vdd.n1691 gnd 0.010231f
C4458 vdd.n1692 gnd 0.010231f
C4459 vdd.n1693 gnd 0.010231f
C4460 vdd.n1694 gnd 0.008235f
C4461 vdd.n1695 gnd 0.010231f
C4462 vdd.n1696 gnd 0.010231f
C4463 vdd.n1697 gnd 0.010231f
C4464 vdd.n1698 gnd 0.010231f
C4465 vdd.n1699 gnd 0.010231f
C4466 vdd.n1700 gnd 0.008235f
C4467 vdd.n1701 gnd 0.010231f
C4468 vdd.n1702 gnd 0.010231f
C4469 vdd.n1703 gnd 0.010231f
C4470 vdd.n1704 gnd 0.010231f
C4471 vdd.n1705 gnd 0.010231f
C4472 vdd.t306 gnd 0.125873f
C4473 vdd.t307 gnd 0.134524f
C4474 vdd.t305 gnd 0.164388f
C4475 vdd.n1706 gnd 0.210723f
C4476 vdd.n1707 gnd 0.177869f
C4477 vdd.n1708 gnd 0.017623f
C4478 vdd.n1709 gnd 0.010231f
C4479 vdd.n1710 gnd 0.010231f
C4480 vdd.n1711 gnd 0.010231f
C4481 vdd.n1712 gnd 0.010231f
C4482 vdd.n1713 gnd 0.010231f
C4483 vdd.n1714 gnd 0.008235f
C4484 vdd.n1715 gnd 0.010231f
C4485 vdd.n1716 gnd 0.010231f
C4486 vdd.n1717 gnd 0.010231f
C4487 vdd.n1718 gnd 0.010231f
C4488 vdd.n1719 gnd 0.010231f
C4489 vdd.n1720 gnd 0.008235f
C4490 vdd.n1721 gnd 0.010231f
C4491 vdd.n1722 gnd 0.010231f
C4492 vdd.n1723 gnd 0.010231f
C4493 vdd.n1724 gnd 0.010231f
C4494 vdd.n1725 gnd 0.010231f
C4495 vdd.n1726 gnd 0.008235f
C4496 vdd.n1727 gnd 0.010231f
C4497 vdd.n1728 gnd 0.010231f
C4498 vdd.n1729 gnd 0.010231f
C4499 vdd.n1730 gnd 0.010231f
C4500 vdd.n1731 gnd 0.010231f
C4501 vdd.n1732 gnd 0.008235f
C4502 vdd.n1733 gnd 0.010231f
C4503 vdd.n1734 gnd 0.010231f
C4504 vdd.n1735 gnd 0.010231f
C4505 vdd.n1736 gnd 0.010231f
C4506 vdd.n1737 gnd 0.010231f
C4507 vdd.n1738 gnd 0.008235f
C4508 vdd.n1739 gnd 0.010231f
C4509 vdd.n1740 gnd 0.010231f
C4510 vdd.n1741 gnd 0.010231f
C4511 vdd.n1742 gnd 0.010231f
C4512 vdd.n1743 gnd 0.008235f
C4513 vdd.n1744 gnd 0.010231f
C4514 vdd.n1745 gnd 0.010231f
C4515 vdd.n1746 gnd 0.010231f
C4516 vdd.n1747 gnd 0.010231f
C4517 vdd.n1748 gnd 0.010231f
C4518 vdd.n1749 gnd 0.008235f
C4519 vdd.n1750 gnd 0.010231f
C4520 vdd.n1751 gnd 0.010231f
C4521 vdd.n1752 gnd 0.010231f
C4522 vdd.n1753 gnd 0.010231f
C4523 vdd.n1754 gnd 0.010231f
C4524 vdd.n1755 gnd 0.008235f
C4525 vdd.n1756 gnd 0.010231f
C4526 vdd.n1757 gnd 0.010231f
C4527 vdd.n1758 gnd 0.010231f
C4528 vdd.n1759 gnd 0.010231f
C4529 vdd.n1760 gnd 0.010231f
C4530 vdd.n1761 gnd 0.008235f
C4531 vdd.n1762 gnd 0.010231f
C4532 vdd.n1763 gnd 0.010231f
C4533 vdd.n1764 gnd 0.010231f
C4534 vdd.n1765 gnd 0.010231f
C4535 vdd.n1766 gnd 0.010231f
C4536 vdd.n1767 gnd 0.008235f
C4537 vdd.n1768 gnd 0.010231f
C4538 vdd.n1769 gnd 0.010231f
C4539 vdd.n1770 gnd 0.010231f
C4540 vdd.n1771 gnd 0.010231f
C4541 vdd.t303 gnd 0.125873f
C4542 vdd.t304 gnd 0.134524f
C4543 vdd.t302 gnd 0.164388f
C4544 vdd.n1772 gnd 0.210723f
C4545 vdd.n1773 gnd 0.177869f
C4546 vdd.n1774 gnd 0.013505f
C4547 vdd.n1775 gnd 0.003912f
C4548 vdd.n1776 gnd 0.025281f
C4549 vdd.n1777 gnd 0.010231f
C4550 vdd.n1778 gnd 0.004323f
C4551 vdd.n1779 gnd 0.008235f
C4552 vdd.n1780 gnd 0.008235f
C4553 vdd.n1781 gnd 0.010231f
C4554 vdd.n1782 gnd 0.010231f
C4555 vdd.n1783 gnd 0.010231f
C4556 vdd.n1784 gnd 0.008235f
C4557 vdd.n1785 gnd 0.008235f
C4558 vdd.n1786 gnd 0.008235f
C4559 vdd.n1787 gnd 0.010231f
C4560 vdd.n1788 gnd 0.010231f
C4561 vdd.n1789 gnd 0.010231f
C4562 vdd.n1790 gnd 0.008235f
C4563 vdd.n1791 gnd 0.008235f
C4564 vdd.n1792 gnd 0.008235f
C4565 vdd.n1793 gnd 0.010231f
C4566 vdd.n1794 gnd 0.010231f
C4567 vdd.n1795 gnd 0.010231f
C4568 vdd.n1796 gnd 0.008235f
C4569 vdd.n1797 gnd 0.008235f
C4570 vdd.n1798 gnd 0.008235f
C4571 vdd.n1799 gnd 0.010231f
C4572 vdd.n1800 gnd 0.010231f
C4573 vdd.n1801 gnd 0.010231f
C4574 vdd.n1802 gnd 0.008235f
C4575 vdd.n1803 gnd 0.008235f
C4576 vdd.n1804 gnd 0.008235f
C4577 vdd.n1805 gnd 0.010231f
C4578 vdd.n1806 gnd 0.010231f
C4579 vdd.n1807 gnd 0.010231f
C4580 vdd.n1808 gnd 0.008153f
C4581 vdd.n1809 gnd 0.010231f
C4582 vdd.t297 gnd 0.125873f
C4583 vdd.t298 gnd 0.134524f
C4584 vdd.t295 gnd 0.164388f
C4585 vdd.n1810 gnd 0.210723f
C4586 vdd.n1811 gnd 0.177869f
C4587 vdd.n1812 gnd 0.017623f
C4588 vdd.n1813 gnd 0.0056f
C4589 vdd.n1814 gnd 0.010231f
C4590 vdd.n1815 gnd 0.010231f
C4591 vdd.n1816 gnd 0.010231f
C4592 vdd.n1817 gnd 0.008235f
C4593 vdd.n1818 gnd 0.008235f
C4594 vdd.n1819 gnd 0.008235f
C4595 vdd.n1820 gnd 0.010231f
C4596 vdd.n1821 gnd 0.010231f
C4597 vdd.n1822 gnd 0.010231f
C4598 vdd.n1823 gnd 0.008235f
C4599 vdd.n1824 gnd 0.008235f
C4600 vdd.n1825 gnd 0.008235f
C4601 vdd.n1826 gnd 0.010231f
C4602 vdd.n1827 gnd 0.010231f
C4603 vdd.n1828 gnd 0.010231f
C4604 vdd.n1829 gnd 0.008235f
C4605 vdd.n1830 gnd 0.008235f
C4606 vdd.n1831 gnd 0.008235f
C4607 vdd.n1832 gnd 0.010231f
C4608 vdd.n1833 gnd 0.010231f
C4609 vdd.n1834 gnd 0.010231f
C4610 vdd.n1835 gnd 0.008235f
C4611 vdd.n1836 gnd 0.008235f
C4612 vdd.n1837 gnd 0.008235f
C4613 vdd.n1838 gnd 0.010231f
C4614 vdd.n1839 gnd 0.010231f
C4615 vdd.n1840 gnd 0.010231f
C4616 vdd.n1841 gnd 0.008235f
C4617 vdd.n1842 gnd 0.008235f
C4618 vdd.n1843 gnd 0.006876f
C4619 vdd.n1844 gnd 0.010231f
C4620 vdd.n1845 gnd 0.010231f
C4621 vdd.n1846 gnd 0.010231f
C4622 vdd.n1847 gnd 0.006876f
C4623 vdd.n1848 gnd 0.008235f
C4624 vdd.n1849 gnd 0.008235f
C4625 vdd.n1850 gnd 0.010231f
C4626 vdd.n1851 gnd 0.010231f
C4627 vdd.n1852 gnd 0.010231f
C4628 vdd.n1853 gnd 0.008235f
C4629 vdd.n1854 gnd 0.008235f
C4630 vdd.n1855 gnd 0.008235f
C4631 vdd.n1856 gnd 0.010231f
C4632 vdd.n1857 gnd 0.010231f
C4633 vdd.n1858 gnd 0.010231f
C4634 vdd.n1859 gnd 0.008235f
C4635 vdd.n1860 gnd 0.008235f
C4636 vdd.n1861 gnd 0.008235f
C4637 vdd.n1862 gnd 0.010231f
C4638 vdd.n1863 gnd 0.010231f
C4639 vdd.n1864 gnd 0.010231f
C4640 vdd.n1865 gnd 0.008235f
C4641 vdd.n1866 gnd 0.008235f
C4642 vdd.n1867 gnd 0.008235f
C4643 vdd.n1868 gnd 0.010231f
C4644 vdd.n1869 gnd 0.010231f
C4645 vdd.n1870 gnd 0.010231f
C4646 vdd.n1871 gnd 0.008235f
C4647 vdd.n1872 gnd 0.010231f
C4648 vdd.n1873 gnd 2.47807f
C4649 vdd.n1875 gnd 0.025281f
C4650 vdd.n1876 gnd 0.006835f
C4651 vdd.n1877 gnd 0.025281f
C4652 vdd.n1878 gnd 0.024751f
C4653 vdd.n1879 gnd 0.010231f
C4654 vdd.n1880 gnd 0.008235f
C4655 vdd.n1881 gnd 0.010231f
C4656 vdd.n1882 gnd 0.528028f
C4657 vdd.n1883 gnd 0.010231f
C4658 vdd.n1884 gnd 0.008235f
C4659 vdd.n1885 gnd 0.010231f
C4660 vdd.n1886 gnd 0.010231f
C4661 vdd.n1887 gnd 0.010231f
C4662 vdd.n1888 gnd 0.008235f
C4663 vdd.n1889 gnd 0.010231f
C4664 vdd.n1890 gnd 0.956723f
C4665 vdd.n1891 gnd 1.0456f
C4666 vdd.n1892 gnd 0.010231f
C4667 vdd.n1893 gnd 0.008235f
C4668 vdd.n1894 gnd 0.010231f
C4669 vdd.n1895 gnd 0.010231f
C4670 vdd.n1896 gnd 0.010231f
C4671 vdd.n1897 gnd 0.008235f
C4672 vdd.n1898 gnd 0.010231f
C4673 vdd.n1899 gnd 0.611676f
C4674 vdd.n1900 gnd 0.010231f
C4675 vdd.n1901 gnd 0.008235f
C4676 vdd.n1902 gnd 0.010231f
C4677 vdd.n1903 gnd 0.010231f
C4678 vdd.n1904 gnd 0.010231f
C4679 vdd.n1905 gnd 0.008235f
C4680 vdd.n1906 gnd 0.010231f
C4681 vdd.n1907 gnd 0.60122f
C4682 vdd.n1908 gnd 0.789427f
C4683 vdd.n1909 gnd 0.010231f
C4684 vdd.n1910 gnd 0.008235f
C4685 vdd.n1911 gnd 0.010231f
C4686 vdd.n1912 gnd 0.010231f
C4687 vdd.n1913 gnd 0.010231f
C4688 vdd.n1914 gnd 0.008235f
C4689 vdd.n1915 gnd 0.010231f
C4690 vdd.n1916 gnd 0.867847f
C4691 vdd.n1917 gnd 0.010231f
C4692 vdd.n1918 gnd 0.008235f
C4693 vdd.n1919 gnd 0.010231f
C4694 vdd.n1920 gnd 0.010231f
C4695 vdd.n1921 gnd 0.010231f
C4696 vdd.n1922 gnd 0.008235f
C4697 vdd.n1923 gnd 0.010231f
C4698 vdd.t106 gnd 0.5228f
C4699 vdd.n1924 gnd 0.768516f
C4700 vdd.n1925 gnd 0.010231f
C4701 vdd.n1926 gnd 0.008235f
C4702 vdd.n1927 gnd 0.010231f
C4703 vdd.n1928 gnd 0.010231f
C4704 vdd.n1929 gnd 0.010231f
C4705 vdd.n1930 gnd 0.008235f
C4706 vdd.n1931 gnd 0.010231f
C4707 vdd.n1932 gnd 0.590764f
C4708 vdd.n1933 gnd 0.010231f
C4709 vdd.n1934 gnd 0.008235f
C4710 vdd.n1935 gnd 0.010231f
C4711 vdd.n1936 gnd 0.010231f
C4712 vdd.n1937 gnd 0.010231f
C4713 vdd.n1938 gnd 0.008235f
C4714 vdd.n1939 gnd 0.010231f
C4715 vdd.n1940 gnd 0.75806f
C4716 vdd.n1941 gnd 0.632588f
C4717 vdd.n1942 gnd 0.010231f
C4718 vdd.n1943 gnd 0.008235f
C4719 vdd.n1944 gnd 0.010231f
C4720 vdd.n1945 gnd 0.010231f
C4721 vdd.n1946 gnd 0.010231f
C4722 vdd.n1947 gnd 0.008235f
C4723 vdd.n1948 gnd 0.010231f
C4724 vdd.n1949 gnd 0.810339f
C4725 vdd.n1950 gnd 0.010231f
C4726 vdd.n1951 gnd 0.008235f
C4727 vdd.n1952 gnd 0.010231f
C4728 vdd.n1953 gnd 0.010231f
C4729 vdd.n1954 gnd 0.010231f
C4730 vdd.n1955 gnd 0.008235f
C4731 vdd.n1956 gnd 0.010231f
C4732 vdd.t74 gnd 0.5228f
C4733 vdd.n1957 gnd 0.867847f
C4734 vdd.n1958 gnd 0.010231f
C4735 vdd.n1959 gnd 0.008235f
C4736 vdd.n1960 gnd 0.010231f
C4737 vdd.n1961 gnd 0.007863f
C4738 vdd.n1962 gnd 0.005615f
C4739 vdd.n1963 gnd 0.005211f
C4740 vdd.n1964 gnd 0.002882f
C4741 vdd.n1965 gnd 0.006618f
C4742 vdd.n1966 gnd 0.0028f
C4743 vdd.n1967 gnd 0.002965f
C4744 vdd.n1968 gnd 0.005211f
C4745 vdd.n1969 gnd 0.0028f
C4746 vdd.n1970 gnd 0.006618f
C4747 vdd.n1971 gnd 0.002965f
C4748 vdd.n1972 gnd 0.005211f
C4749 vdd.n1973 gnd 0.0028f
C4750 vdd.n1974 gnd 0.004963f
C4751 vdd.n1975 gnd 0.004978f
C4752 vdd.t35 gnd 0.014218f
C4753 vdd.n1976 gnd 0.031635f
C4754 vdd.n1977 gnd 0.164637f
C4755 vdd.n1978 gnd 0.0028f
C4756 vdd.n1979 gnd 0.002965f
C4757 vdd.n1980 gnd 0.006618f
C4758 vdd.n1981 gnd 0.006618f
C4759 vdd.n1982 gnd 0.002965f
C4760 vdd.n1983 gnd 0.0028f
C4761 vdd.n1984 gnd 0.005211f
C4762 vdd.n1985 gnd 0.005211f
C4763 vdd.n1986 gnd 0.0028f
C4764 vdd.n1987 gnd 0.002965f
C4765 vdd.n1988 gnd 0.006618f
C4766 vdd.n1989 gnd 0.006618f
C4767 vdd.n1990 gnd 0.002965f
C4768 vdd.n1991 gnd 0.0028f
C4769 vdd.n1992 gnd 0.005211f
C4770 vdd.n1993 gnd 0.005211f
C4771 vdd.n1994 gnd 0.0028f
C4772 vdd.n1995 gnd 0.002965f
C4773 vdd.n1996 gnd 0.006618f
C4774 vdd.n1997 gnd 0.006618f
C4775 vdd.n1998 gnd 0.015646f
C4776 vdd.n1999 gnd 0.002882f
C4777 vdd.n2000 gnd 0.0028f
C4778 vdd.n2001 gnd 0.013467f
C4779 vdd.n2002 gnd 0.009402f
C4780 vdd.t213 gnd 0.03294f
C4781 vdd.t216 gnd 0.03294f
C4782 vdd.n2003 gnd 0.226387f
C4783 vdd.n2004 gnd 0.178019f
C4784 vdd.t1 gnd 0.03294f
C4785 vdd.t96 gnd 0.03294f
C4786 vdd.n2005 gnd 0.226387f
C4787 vdd.n2006 gnd 0.14366f
C4788 vdd.t90 gnd 0.03294f
C4789 vdd.t100 gnd 0.03294f
C4790 vdd.n2007 gnd 0.226387f
C4791 vdd.n2008 gnd 0.14366f
C4792 vdd.t215 gnd 0.03294f
C4793 vdd.t88 gnd 0.03294f
C4794 vdd.n2009 gnd 0.226387f
C4795 vdd.n2010 gnd 0.14366f
C4796 vdd.t111 gnd 0.03294f
C4797 vdd.t18 gnd 0.03294f
C4798 vdd.n2011 gnd 0.226387f
C4799 vdd.n2012 gnd 0.14366f
C4800 vdd.t132 gnd 0.03294f
C4801 vdd.t122 gnd 0.03294f
C4802 vdd.n2013 gnd 0.226387f
C4803 vdd.n2014 gnd 0.14366f
C4804 vdd.t231 gnd 0.03294f
C4805 vdd.t129 gnd 0.03294f
C4806 vdd.n2015 gnd 0.226387f
C4807 vdd.n2016 gnd 0.14366f
C4808 vdd.t68 gnd 0.03294f
C4809 vdd.t224 gnd 0.03294f
C4810 vdd.n2017 gnd 0.226387f
C4811 vdd.n2018 gnd 0.14366f
C4812 vdd.t214 gnd 0.03294f
C4813 vdd.t86 gnd 0.03294f
C4814 vdd.n2019 gnd 0.226387f
C4815 vdd.n2020 gnd 0.14366f
C4816 vdd.n2021 gnd 0.005615f
C4817 vdd.n2022 gnd 0.005211f
C4818 vdd.n2023 gnd 0.002882f
C4819 vdd.n2024 gnd 0.006618f
C4820 vdd.n2025 gnd 0.0028f
C4821 vdd.n2026 gnd 0.002965f
C4822 vdd.n2027 gnd 0.005211f
C4823 vdd.n2028 gnd 0.0028f
C4824 vdd.n2029 gnd 0.006618f
C4825 vdd.n2030 gnd 0.002965f
C4826 vdd.n2031 gnd 0.005211f
C4827 vdd.n2032 gnd 0.0028f
C4828 vdd.n2033 gnd 0.004963f
C4829 vdd.n2034 gnd 0.004978f
C4830 vdd.t22 gnd 0.014218f
C4831 vdd.n2035 gnd 0.031635f
C4832 vdd.n2036 gnd 0.164637f
C4833 vdd.n2037 gnd 0.0028f
C4834 vdd.n2038 gnd 0.002965f
C4835 vdd.n2039 gnd 0.006618f
C4836 vdd.n2040 gnd 0.006618f
C4837 vdd.n2041 gnd 0.002965f
C4838 vdd.n2042 gnd 0.0028f
C4839 vdd.n2043 gnd 0.005211f
C4840 vdd.n2044 gnd 0.005211f
C4841 vdd.n2045 gnd 0.0028f
C4842 vdd.n2046 gnd 0.002965f
C4843 vdd.n2047 gnd 0.006618f
C4844 vdd.n2048 gnd 0.006618f
C4845 vdd.n2049 gnd 0.002965f
C4846 vdd.n2050 gnd 0.0028f
C4847 vdd.n2051 gnd 0.005211f
C4848 vdd.n2052 gnd 0.005211f
C4849 vdd.n2053 gnd 0.0028f
C4850 vdd.n2054 gnd 0.002965f
C4851 vdd.n2055 gnd 0.006618f
C4852 vdd.n2056 gnd 0.006618f
C4853 vdd.n2057 gnd 0.015646f
C4854 vdd.n2058 gnd 0.002882f
C4855 vdd.n2059 gnd 0.0028f
C4856 vdd.n2060 gnd 0.013467f
C4857 vdd.n2061 gnd 0.009107f
C4858 vdd.n2062 gnd 0.106884f
C4859 vdd.n2063 gnd 0.005615f
C4860 vdd.n2064 gnd 0.005211f
C4861 vdd.n2065 gnd 0.002882f
C4862 vdd.n2066 gnd 0.006618f
C4863 vdd.n2067 gnd 0.0028f
C4864 vdd.n2068 gnd 0.002965f
C4865 vdd.n2069 gnd 0.005211f
C4866 vdd.n2070 gnd 0.0028f
C4867 vdd.n2071 gnd 0.006618f
C4868 vdd.n2072 gnd 0.002965f
C4869 vdd.n2073 gnd 0.005211f
C4870 vdd.n2074 gnd 0.0028f
C4871 vdd.n2075 gnd 0.004963f
C4872 vdd.n2076 gnd 0.004978f
C4873 vdd.t223 gnd 0.014218f
C4874 vdd.n2077 gnd 0.031635f
C4875 vdd.n2078 gnd 0.164637f
C4876 vdd.n2079 gnd 0.0028f
C4877 vdd.n2080 gnd 0.002965f
C4878 vdd.n2081 gnd 0.006618f
C4879 vdd.n2082 gnd 0.006618f
C4880 vdd.n2083 gnd 0.002965f
C4881 vdd.n2084 gnd 0.0028f
C4882 vdd.n2085 gnd 0.005211f
C4883 vdd.n2086 gnd 0.005211f
C4884 vdd.n2087 gnd 0.0028f
C4885 vdd.n2088 gnd 0.002965f
C4886 vdd.n2089 gnd 0.006618f
C4887 vdd.n2090 gnd 0.006618f
C4888 vdd.n2091 gnd 0.002965f
C4889 vdd.n2092 gnd 0.0028f
C4890 vdd.n2093 gnd 0.005211f
C4891 vdd.n2094 gnd 0.005211f
C4892 vdd.n2095 gnd 0.0028f
C4893 vdd.n2096 gnd 0.002965f
C4894 vdd.n2097 gnd 0.006618f
C4895 vdd.n2098 gnd 0.006618f
C4896 vdd.n2099 gnd 0.015646f
C4897 vdd.n2100 gnd 0.002882f
C4898 vdd.n2101 gnd 0.0028f
C4899 vdd.n2102 gnd 0.013467f
C4900 vdd.n2103 gnd 0.009402f
C4901 vdd.t92 gnd 0.03294f
C4902 vdd.t205 gnd 0.03294f
C4903 vdd.n2104 gnd 0.226387f
C4904 vdd.n2105 gnd 0.178019f
C4905 vdd.t61 gnd 0.03294f
C4906 vdd.t93 gnd 0.03294f
C4907 vdd.n2106 gnd 0.226387f
C4908 vdd.n2107 gnd 0.14366f
C4909 vdd.t60 gnd 0.03294f
C4910 vdd.t102 gnd 0.03294f
C4911 vdd.n2108 gnd 0.226387f
C4912 vdd.n2109 gnd 0.14366f
C4913 vdd.t54 gnd 0.03294f
C4914 vdd.t94 gnd 0.03294f
C4915 vdd.n2110 gnd 0.226387f
C4916 vdd.n2111 gnd 0.14366f
C4917 vdd.t75 gnd 0.03294f
C4918 vdd.t31 gnd 0.03294f
C4919 vdd.n2112 gnd 0.226387f
C4920 vdd.n2113 gnd 0.14366f
C4921 vdd.t208 gnd 0.03294f
C4922 vdd.t44 gnd 0.03294f
C4923 vdd.n2114 gnd 0.226387f
C4924 vdd.n2115 gnd 0.14366f
C4925 vdd.t222 gnd 0.03294f
C4926 vdd.t115 gnd 0.03294f
C4927 vdd.n2116 gnd 0.226387f
C4928 vdd.n2117 gnd 0.14366f
C4929 vdd.t130 gnd 0.03294f
C4930 vdd.t203 gnd 0.03294f
C4931 vdd.n2118 gnd 0.226387f
C4932 vdd.n2119 gnd 0.14366f
C4933 vdd.t33 gnd 0.03294f
C4934 vdd.t199 gnd 0.03294f
C4935 vdd.n2120 gnd 0.226387f
C4936 vdd.n2121 gnd 0.14366f
C4937 vdd.n2122 gnd 0.005615f
C4938 vdd.n2123 gnd 0.005211f
C4939 vdd.n2124 gnd 0.002882f
C4940 vdd.n2125 gnd 0.006618f
C4941 vdd.n2126 gnd 0.0028f
C4942 vdd.n2127 gnd 0.002965f
C4943 vdd.n2128 gnd 0.005211f
C4944 vdd.n2129 gnd 0.0028f
C4945 vdd.n2130 gnd 0.006618f
C4946 vdd.n2131 gnd 0.002965f
C4947 vdd.n2132 gnd 0.005211f
C4948 vdd.n2133 gnd 0.0028f
C4949 vdd.n2134 gnd 0.004963f
C4950 vdd.n2135 gnd 0.004978f
C4951 vdd.t101 gnd 0.014218f
C4952 vdd.n2136 gnd 0.031635f
C4953 vdd.n2137 gnd 0.164637f
C4954 vdd.n2138 gnd 0.0028f
C4955 vdd.n2139 gnd 0.002965f
C4956 vdd.n2140 gnd 0.006618f
C4957 vdd.n2141 gnd 0.006618f
C4958 vdd.n2142 gnd 0.002965f
C4959 vdd.n2143 gnd 0.0028f
C4960 vdd.n2144 gnd 0.005211f
C4961 vdd.n2145 gnd 0.005211f
C4962 vdd.n2146 gnd 0.0028f
C4963 vdd.n2147 gnd 0.002965f
C4964 vdd.n2148 gnd 0.006618f
C4965 vdd.n2149 gnd 0.006618f
C4966 vdd.n2150 gnd 0.002965f
C4967 vdd.n2151 gnd 0.0028f
C4968 vdd.n2152 gnd 0.005211f
C4969 vdd.n2153 gnd 0.005211f
C4970 vdd.n2154 gnd 0.0028f
C4971 vdd.n2155 gnd 0.002965f
C4972 vdd.n2156 gnd 0.006618f
C4973 vdd.n2157 gnd 0.006618f
C4974 vdd.n2158 gnd 0.015646f
C4975 vdd.n2159 gnd 0.002882f
C4976 vdd.n2160 gnd 0.0028f
C4977 vdd.n2161 gnd 0.013467f
C4978 vdd.n2162 gnd 0.009107f
C4979 vdd.n2163 gnd 0.063585f
C4980 vdd.n2164 gnd 0.229114f
C4981 vdd.n2165 gnd 0.005615f
C4982 vdd.n2166 gnd 0.005211f
C4983 vdd.n2167 gnd 0.002882f
C4984 vdd.n2168 gnd 0.006618f
C4985 vdd.n2169 gnd 0.0028f
C4986 vdd.n2170 gnd 0.002965f
C4987 vdd.n2171 gnd 0.005211f
C4988 vdd.n2172 gnd 0.0028f
C4989 vdd.n2173 gnd 0.006618f
C4990 vdd.n2174 gnd 0.002965f
C4991 vdd.n2175 gnd 0.005211f
C4992 vdd.n2176 gnd 0.0028f
C4993 vdd.n2177 gnd 0.004963f
C4994 vdd.n2178 gnd 0.004978f
C4995 vdd.t57 gnd 0.014218f
C4996 vdd.n2179 gnd 0.031635f
C4997 vdd.n2180 gnd 0.164637f
C4998 vdd.n2181 gnd 0.0028f
C4999 vdd.n2182 gnd 0.002965f
C5000 vdd.n2183 gnd 0.006618f
C5001 vdd.n2184 gnd 0.006618f
C5002 vdd.n2185 gnd 0.002965f
C5003 vdd.n2186 gnd 0.0028f
C5004 vdd.n2187 gnd 0.005211f
C5005 vdd.n2188 gnd 0.005211f
C5006 vdd.n2189 gnd 0.0028f
C5007 vdd.n2190 gnd 0.002965f
C5008 vdd.n2191 gnd 0.006618f
C5009 vdd.n2192 gnd 0.006618f
C5010 vdd.n2193 gnd 0.002965f
C5011 vdd.n2194 gnd 0.0028f
C5012 vdd.n2195 gnd 0.005211f
C5013 vdd.n2196 gnd 0.005211f
C5014 vdd.n2197 gnd 0.0028f
C5015 vdd.n2198 gnd 0.002965f
C5016 vdd.n2199 gnd 0.006618f
C5017 vdd.n2200 gnd 0.006618f
C5018 vdd.n2201 gnd 0.015646f
C5019 vdd.n2202 gnd 0.002882f
C5020 vdd.n2203 gnd 0.0028f
C5021 vdd.n2204 gnd 0.013467f
C5022 vdd.n2205 gnd 0.009402f
C5023 vdd.t226 gnd 0.03294f
C5024 vdd.t227 gnd 0.03294f
C5025 vdd.n2206 gnd 0.226387f
C5026 vdd.n2207 gnd 0.178019f
C5027 vdd.t126 gnd 0.03294f
C5028 vdd.t10 gnd 0.03294f
C5029 vdd.n2208 gnd 0.226387f
C5030 vdd.n2209 gnd 0.14366f
C5031 vdd.t95 gnd 0.03294f
C5032 vdd.t108 gnd 0.03294f
C5033 vdd.n2210 gnd 0.226387f
C5034 vdd.n2211 gnd 0.14366f
C5035 vdd.t128 gnd 0.03294f
C5036 vdd.t12 gnd 0.03294f
C5037 vdd.n2212 gnd 0.226387f
C5038 vdd.n2213 gnd 0.14366f
C5039 vdd.t134 gnd 0.03294f
C5040 vdd.t210 gnd 0.03294f
C5041 vdd.n2214 gnd 0.226387f
C5042 vdd.n2215 gnd 0.14366f
C5043 vdd.t211 gnd 0.03294f
C5044 vdd.t63 gnd 0.03294f
C5045 vdd.n2216 gnd 0.226387f
C5046 vdd.n2217 gnd 0.14366f
C5047 vdd.t52 gnd 0.03294f
C5048 vdd.t230 gnd 0.03294f
C5049 vdd.n2218 gnd 0.226387f
C5050 vdd.n2219 gnd 0.14366f
C5051 vdd.t81 gnd 0.03294f
C5052 vdd.t107 gnd 0.03294f
C5053 vdd.n2220 gnd 0.226387f
C5054 vdd.n2221 gnd 0.14366f
C5055 vdd.t207 gnd 0.03294f
C5056 vdd.t127 gnd 0.03294f
C5057 vdd.n2222 gnd 0.226387f
C5058 vdd.n2223 gnd 0.14366f
C5059 vdd.n2224 gnd 0.005615f
C5060 vdd.n2225 gnd 0.005211f
C5061 vdd.n2226 gnd 0.002882f
C5062 vdd.n2227 gnd 0.006618f
C5063 vdd.n2228 gnd 0.0028f
C5064 vdd.n2229 gnd 0.002965f
C5065 vdd.n2230 gnd 0.005211f
C5066 vdd.n2231 gnd 0.0028f
C5067 vdd.n2232 gnd 0.006618f
C5068 vdd.n2233 gnd 0.002965f
C5069 vdd.n2234 gnd 0.005211f
C5070 vdd.n2235 gnd 0.0028f
C5071 vdd.n2236 gnd 0.004963f
C5072 vdd.n2237 gnd 0.004978f
C5073 vdd.t206 gnd 0.014218f
C5074 vdd.n2238 gnd 0.031635f
C5075 vdd.n2239 gnd 0.164637f
C5076 vdd.n2240 gnd 0.0028f
C5077 vdd.n2241 gnd 0.002965f
C5078 vdd.n2242 gnd 0.006618f
C5079 vdd.n2243 gnd 0.006618f
C5080 vdd.n2244 gnd 0.002965f
C5081 vdd.n2245 gnd 0.0028f
C5082 vdd.n2246 gnd 0.005211f
C5083 vdd.n2247 gnd 0.005211f
C5084 vdd.n2248 gnd 0.0028f
C5085 vdd.n2249 gnd 0.002965f
C5086 vdd.n2250 gnd 0.006618f
C5087 vdd.n2251 gnd 0.006618f
C5088 vdd.n2252 gnd 0.002965f
C5089 vdd.n2253 gnd 0.0028f
C5090 vdd.n2254 gnd 0.005211f
C5091 vdd.n2255 gnd 0.005211f
C5092 vdd.n2256 gnd 0.0028f
C5093 vdd.n2257 gnd 0.002965f
C5094 vdd.n2258 gnd 0.006618f
C5095 vdd.n2259 gnd 0.006618f
C5096 vdd.n2260 gnd 0.015646f
C5097 vdd.n2261 gnd 0.002882f
C5098 vdd.n2262 gnd 0.0028f
C5099 vdd.n2263 gnd 0.013467f
C5100 vdd.n2264 gnd 0.009107f
C5101 vdd.n2265 gnd 0.063585f
C5102 vdd.n2266 gnd 0.262286f
C5103 vdd.n2267 gnd 2.99909f
C5104 vdd.n2268 gnd 0.603486f
C5105 vdd.n2269 gnd 0.007863f
C5106 vdd.n2270 gnd 0.008235f
C5107 vdd.n2271 gnd 0.010231f
C5108 vdd.n2272 gnd 0.747604f
C5109 vdd.n2273 gnd 0.010231f
C5110 vdd.n2274 gnd 0.008235f
C5111 vdd.n2275 gnd 0.010231f
C5112 vdd.n2276 gnd 0.010231f
C5113 vdd.n2277 gnd 0.010231f
C5114 vdd.n2278 gnd 0.008235f
C5115 vdd.n2279 gnd 0.010231f
C5116 vdd.n2280 gnd 0.867847f
C5117 vdd.t53 gnd 0.5228f
C5118 vdd.n2281 gnd 0.569852f
C5119 vdd.n2282 gnd 0.010231f
C5120 vdd.n2283 gnd 0.008235f
C5121 vdd.n2284 gnd 0.010231f
C5122 vdd.n2285 gnd 0.010231f
C5123 vdd.n2286 gnd 0.010231f
C5124 vdd.n2287 gnd 0.008235f
C5125 vdd.n2288 gnd 0.010231f
C5126 vdd.n2289 gnd 0.6535f
C5127 vdd.n2290 gnd 0.010231f
C5128 vdd.n2291 gnd 0.008235f
C5129 vdd.n2292 gnd 0.010231f
C5130 vdd.n2293 gnd 0.010231f
C5131 vdd.n2294 gnd 0.010231f
C5132 vdd.n2295 gnd 0.008235f
C5133 vdd.n2296 gnd 0.010231f
C5134 vdd.n2297 gnd 0.559396f
C5135 vdd.n2298 gnd 0.831251f
C5136 vdd.n2299 gnd 0.010231f
C5137 vdd.n2300 gnd 0.008235f
C5138 vdd.n2301 gnd 0.010231f
C5139 vdd.n2302 gnd 0.010231f
C5140 vdd.n2303 gnd 0.010231f
C5141 vdd.n2304 gnd 0.008235f
C5142 vdd.n2305 gnd 0.010231f
C5143 vdd.n2306 gnd 0.867847f
C5144 vdd.n2307 gnd 0.010231f
C5145 vdd.n2308 gnd 0.008235f
C5146 vdd.n2309 gnd 0.010231f
C5147 vdd.n2310 gnd 0.010231f
C5148 vdd.n2311 gnd 0.010231f
C5149 vdd.n2312 gnd 0.008235f
C5150 vdd.n2313 gnd 0.010231f
C5151 vdd.t9 gnd 0.5228f
C5152 vdd.n2314 gnd 0.726692f
C5153 vdd.n2315 gnd 0.010231f
C5154 vdd.n2316 gnd 0.008235f
C5155 vdd.n2317 gnd 0.010231f
C5156 vdd.n2318 gnd 0.010231f
C5157 vdd.n2319 gnd 0.010231f
C5158 vdd.n2320 gnd 0.008235f
C5159 vdd.n2321 gnd 0.010231f
C5160 vdd.n2322 gnd 0.54894f
C5161 vdd.n2323 gnd 0.010231f
C5162 vdd.n2324 gnd 0.008235f
C5163 vdd.n2325 gnd 0.010231f
C5164 vdd.n2326 gnd 0.010231f
C5165 vdd.n2327 gnd 0.010231f
C5166 vdd.n2328 gnd 0.008235f
C5167 vdd.n2329 gnd 0.010231f
C5168 vdd.n2330 gnd 0.716236f
C5169 vdd.n2331 gnd 0.674412f
C5170 vdd.n2332 gnd 0.010231f
C5171 vdd.n2333 gnd 0.008235f
C5172 vdd.n2334 gnd 0.010231f
C5173 vdd.n2335 gnd 0.010231f
C5174 vdd.n2336 gnd 0.010231f
C5175 vdd.n2337 gnd 0.008235f
C5176 vdd.n2338 gnd 0.010231f
C5177 vdd.n2339 gnd 0.852163f
C5178 vdd.n2340 gnd 0.010231f
C5179 vdd.n2341 gnd 0.008235f
C5180 vdd.n2342 gnd 0.010231f
C5181 vdd.n2343 gnd 0.010231f
C5182 vdd.n2344 gnd 0.024751f
C5183 vdd.n2345 gnd 0.010231f
C5184 vdd.n2346 gnd 0.010231f
C5185 vdd.n2347 gnd 0.008235f
C5186 vdd.n2348 gnd 0.010231f
C5187 vdd.n2349 gnd 0.632588f
C5188 vdd.n2350 gnd 1.0456f
C5189 vdd.n2351 gnd 0.010231f
C5190 vdd.n2352 gnd 0.008235f
C5191 vdd.n2353 gnd 0.010231f
C5192 vdd.n2354 gnd 0.010231f
C5193 vdd.n2355 gnd 0.024751f
C5194 vdd.n2356 gnd 0.006835f
C5195 vdd.n2357 gnd 0.024751f
C5196 vdd.n2358 gnd 1.4377f
C5197 vdd.n2359 gnd 0.024751f
C5198 vdd.n2360 gnd 0.025281f
C5199 vdd.n2361 gnd 0.003912f
C5200 vdd.t267 gnd 0.125873f
C5201 vdd.t266 gnd 0.134524f
C5202 vdd.t265 gnd 0.164388f
C5203 vdd.n2362 gnd 0.210723f
C5204 vdd.n2363 gnd 0.177045f
C5205 vdd.n2364 gnd 0.012682f
C5206 vdd.n2365 gnd 0.004323f
C5207 vdd.n2366 gnd 0.008799f
C5208 vdd.n2367 gnd 1.08617f
C5209 vdd.n2369 gnd 0.008235f
C5210 vdd.n2370 gnd 0.008235f
C5211 vdd.n2371 gnd 0.010231f
C5212 vdd.n2373 gnd 0.010231f
C5213 vdd.n2374 gnd 0.010231f
C5214 vdd.n2375 gnd 0.008235f
C5215 vdd.n2376 gnd 0.008235f
C5216 vdd.n2377 gnd 0.008235f
C5217 vdd.n2378 gnd 0.010231f
C5218 vdd.n2380 gnd 0.010231f
C5219 vdd.n2381 gnd 0.010231f
C5220 vdd.n2382 gnd 0.008235f
C5221 vdd.n2383 gnd 0.008235f
C5222 vdd.n2384 gnd 0.008235f
C5223 vdd.n2385 gnd 0.010231f
C5224 vdd.n2387 gnd 0.010231f
C5225 vdd.n2388 gnd 0.010231f
C5226 vdd.n2389 gnd 0.008235f
C5227 vdd.n2390 gnd 0.008235f
C5228 vdd.n2391 gnd 0.008235f
C5229 vdd.n2392 gnd 0.010231f
C5230 vdd.n2394 gnd 0.010231f
C5231 vdd.n2395 gnd 0.010231f
C5232 vdd.n2396 gnd 0.008235f
C5233 vdd.n2397 gnd 0.010231f
C5234 vdd.n2398 gnd 0.010231f
C5235 vdd.n2399 gnd 0.010231f
C5236 vdd.n2400 gnd 0.016799f
C5237 vdd.n2401 gnd 0.0056f
C5238 vdd.n2402 gnd 0.008235f
C5239 vdd.n2403 gnd 0.010231f
C5240 vdd.n2405 gnd 0.010231f
C5241 vdd.n2406 gnd 0.010231f
C5242 vdd.n2407 gnd 0.008235f
C5243 vdd.n2408 gnd 0.008235f
C5244 vdd.n2409 gnd 0.008235f
C5245 vdd.n2410 gnd 0.010231f
C5246 vdd.n2412 gnd 0.010231f
C5247 vdd.n2413 gnd 0.010231f
C5248 vdd.n2414 gnd 0.008235f
C5249 vdd.n2415 gnd 0.008235f
C5250 vdd.n2416 gnd 0.008235f
C5251 vdd.n2417 gnd 0.010231f
C5252 vdd.n2419 gnd 0.010231f
C5253 vdd.n2420 gnd 0.010231f
C5254 vdd.n2421 gnd 0.008235f
C5255 vdd.n2422 gnd 0.008235f
C5256 vdd.n2423 gnd 0.008235f
C5257 vdd.n2424 gnd 0.010231f
C5258 vdd.n2426 gnd 0.010231f
C5259 vdd.n2427 gnd 0.010231f
C5260 vdd.n2428 gnd 0.008235f
C5261 vdd.n2429 gnd 0.008235f
C5262 vdd.n2430 gnd 0.008235f
C5263 vdd.n2431 gnd 0.010231f
C5264 vdd.n2433 gnd 0.010231f
C5265 vdd.n2434 gnd 0.010231f
C5266 vdd.n2435 gnd 0.008235f
C5267 vdd.n2436 gnd 0.010231f
C5268 vdd.n2437 gnd 0.010231f
C5269 vdd.n2438 gnd 0.010231f
C5270 vdd.n2439 gnd 0.016799f
C5271 vdd.n2440 gnd 0.006876f
C5272 vdd.n2441 gnd 0.008235f
C5273 vdd.n2442 gnd 0.010231f
C5274 vdd.n2444 gnd 0.010231f
C5275 vdd.n2445 gnd 0.010231f
C5276 vdd.n2446 gnd 0.008235f
C5277 vdd.n2447 gnd 0.008235f
C5278 vdd.n2448 gnd 0.008235f
C5279 vdd.n2449 gnd 0.010231f
C5280 vdd.n2451 gnd 0.010231f
C5281 vdd.n2452 gnd 0.010231f
C5282 vdd.n2453 gnd 0.008235f
C5283 vdd.n2454 gnd 0.008235f
C5284 vdd.n2455 gnd 0.008235f
C5285 vdd.n2456 gnd 0.010231f
C5286 vdd.n2458 gnd 0.010231f
C5287 vdd.n2459 gnd 0.010231f
C5288 vdd.n2460 gnd 0.008235f
C5289 vdd.n2461 gnd 0.008235f
C5290 vdd.n2462 gnd 0.008235f
C5291 vdd.n2463 gnd 0.010231f
C5292 vdd.n2465 gnd 0.010231f
C5293 vdd.n2466 gnd 0.008235f
C5294 vdd.n2467 gnd 0.008235f
C5295 vdd.n2468 gnd 0.010231f
C5296 vdd.n2470 gnd 0.010231f
C5297 vdd.n2471 gnd 0.010231f
C5298 vdd.n2472 gnd 0.008235f
C5299 vdd.n2473 gnd 0.008799f
C5300 vdd.n2474 gnd 1.08617f
C5301 vdd.n2475 gnd 0.046868f
C5302 vdd.n2476 gnd 0.006957f
C5303 vdd.n2477 gnd 0.006957f
C5304 vdd.n2478 gnd 0.006957f
C5305 vdd.n2479 gnd 0.006957f
C5306 vdd.n2480 gnd 0.006957f
C5307 vdd.n2481 gnd 0.006957f
C5308 vdd.n2482 gnd 0.006957f
C5309 vdd.n2483 gnd 0.006957f
C5310 vdd.n2484 gnd 0.006957f
C5311 vdd.n2485 gnd 0.006957f
C5312 vdd.n2486 gnd 0.006957f
C5313 vdd.n2487 gnd 0.006957f
C5314 vdd.n2488 gnd 0.006957f
C5315 vdd.n2489 gnd 0.006957f
C5316 vdd.n2490 gnd 0.006957f
C5317 vdd.n2491 gnd 0.006957f
C5318 vdd.n2492 gnd 0.006957f
C5319 vdd.n2493 gnd 0.006957f
C5320 vdd.n2494 gnd 0.006957f
C5321 vdd.n2495 gnd 0.006957f
C5322 vdd.n2496 gnd 0.006957f
C5323 vdd.n2497 gnd 0.006957f
C5324 vdd.n2498 gnd 0.006957f
C5325 vdd.n2499 gnd 0.006957f
C5326 vdd.n2500 gnd 0.006957f
C5327 vdd.n2501 gnd 0.006957f
C5328 vdd.n2502 gnd 0.006957f
C5329 vdd.n2503 gnd 0.006957f
C5330 vdd.n2504 gnd 0.006957f
C5331 vdd.n2505 gnd 0.006957f
C5332 vdd.n2506 gnd 12.3485f
C5333 vdd.n2508 gnd 0.015797f
C5334 vdd.n2509 gnd 0.015797f
C5335 vdd.n2510 gnd 0.014897f
C5336 vdd.n2511 gnd 0.006957f
C5337 vdd.n2512 gnd 0.006957f
C5338 vdd.n2513 gnd 0.711008f
C5339 vdd.n2514 gnd 0.006957f
C5340 vdd.n2515 gnd 0.006957f
C5341 vdd.n2516 gnd 0.006957f
C5342 vdd.n2517 gnd 0.006957f
C5343 vdd.n2518 gnd 0.006957f
C5344 vdd.n2519 gnd 0.559396f
C5345 vdd.n2520 gnd 0.006957f
C5346 vdd.n2521 gnd 0.006957f
C5347 vdd.n2522 gnd 0.006957f
C5348 vdd.n2523 gnd 0.006957f
C5349 vdd.n2524 gnd 0.006957f
C5350 vdd.n2525 gnd 0.711008f
C5351 vdd.n2526 gnd 0.006957f
C5352 vdd.n2527 gnd 0.006957f
C5353 vdd.n2528 gnd 0.006957f
C5354 vdd.n2529 gnd 0.006957f
C5355 vdd.n2530 gnd 0.006957f
C5356 vdd.n2531 gnd 0.711008f
C5357 vdd.n2532 gnd 0.006957f
C5358 vdd.n2533 gnd 0.006957f
C5359 vdd.n2534 gnd 0.006957f
C5360 vdd.n2535 gnd 0.006957f
C5361 vdd.n2536 gnd 0.006957f
C5362 vdd.n2537 gnd 0.684868f
C5363 vdd.n2538 gnd 0.006957f
C5364 vdd.n2539 gnd 0.006957f
C5365 vdd.n2540 gnd 0.006957f
C5366 vdd.n2541 gnd 0.006957f
C5367 vdd.n2542 gnd 0.006957f
C5368 vdd.n2543 gnd 0.528028f
C5369 vdd.n2544 gnd 0.006957f
C5370 vdd.n2545 gnd 0.006957f
C5371 vdd.n2546 gnd 0.006957f
C5372 vdd.n2547 gnd 0.006957f
C5373 vdd.n2548 gnd 0.006957f
C5374 vdd.n2549 gnd 0.371188f
C5375 vdd.n2550 gnd 0.006957f
C5376 vdd.n2551 gnd 0.006957f
C5377 vdd.n2552 gnd 0.006957f
C5378 vdd.n2553 gnd 0.006957f
C5379 vdd.n2554 gnd 0.006957f
C5380 vdd.n2555 gnd 0.49666f
C5381 vdd.n2556 gnd 0.006957f
C5382 vdd.n2557 gnd 0.006957f
C5383 vdd.n2558 gnd 0.006957f
C5384 vdd.n2559 gnd 0.006957f
C5385 vdd.n2560 gnd 0.006957f
C5386 vdd.n2561 gnd 0.6535f
C5387 vdd.n2562 gnd 0.006957f
C5388 vdd.n2563 gnd 0.006957f
C5389 vdd.n2564 gnd 0.006957f
C5390 vdd.n2565 gnd 0.006957f
C5391 vdd.n2566 gnd 0.006957f
C5392 vdd.n2567 gnd 0.711008f
C5393 vdd.n2568 gnd 0.006957f
C5394 vdd.n2569 gnd 0.006957f
C5395 vdd.n2570 gnd 0.006957f
C5396 vdd.n2571 gnd 0.006957f
C5397 vdd.n2572 gnd 0.006957f
C5398 vdd.n2573 gnd 0.611676f
C5399 vdd.n2574 gnd 0.006957f
C5400 vdd.n2575 gnd 0.006957f
C5401 vdd.n2576 gnd 0.005525f
C5402 vdd.n2577 gnd 0.020155f
C5403 vdd.n2578 gnd 0.004911f
C5404 vdd.n2579 gnd 0.006957f
C5405 vdd.n2580 gnd 0.454836f
C5406 vdd.n2581 gnd 0.006957f
C5407 vdd.n2582 gnd 0.006957f
C5408 vdd.n2583 gnd 0.006957f
C5409 vdd.n2584 gnd 0.006957f
C5410 vdd.n2585 gnd 0.006957f
C5411 vdd.n2586 gnd 0.413012f
C5412 vdd.n2587 gnd 0.006957f
C5413 vdd.n2588 gnd 0.006957f
C5414 vdd.n2589 gnd 0.006957f
C5415 vdd.n2590 gnd 0.006957f
C5416 vdd.n2591 gnd 0.006957f
C5417 vdd.n2592 gnd 0.569852f
C5418 vdd.n2593 gnd 0.006957f
C5419 vdd.n2594 gnd 0.006957f
C5420 vdd.n2595 gnd 0.006957f
C5421 vdd.n2596 gnd 0.006957f
C5422 vdd.n2597 gnd 0.006957f
C5423 vdd.n2598 gnd 0.62736f
C5424 vdd.n2599 gnd 0.006957f
C5425 vdd.n2600 gnd 0.006957f
C5426 vdd.n2601 gnd 0.006957f
C5427 vdd.n2602 gnd 0.006957f
C5428 vdd.n2603 gnd 0.006957f
C5429 vdd.n2604 gnd 0.47052f
C5430 vdd.n2605 gnd 0.006957f
C5431 vdd.n2606 gnd 0.006957f
C5432 vdd.n2607 gnd 0.006957f
C5433 vdd.n2608 gnd 0.006957f
C5434 vdd.n2609 gnd 0.006957f
C5435 vdd.n2610 gnd 0.224804f
C5436 vdd.n2611 gnd 0.006957f
C5437 vdd.n2612 gnd 0.006957f
C5438 vdd.n2613 gnd 0.006957f
C5439 vdd.n2614 gnd 0.006957f
C5440 vdd.n2615 gnd 0.006957f
C5441 vdd.n2616 gnd 0.224804f
C5442 vdd.n2617 gnd 0.006957f
C5443 vdd.n2618 gnd 0.006957f
C5444 vdd.n2619 gnd 0.006957f
C5445 vdd.n2620 gnd 0.006957f
C5446 vdd.n2621 gnd 0.006957f
C5447 vdd.n2622 gnd 0.711008f
C5448 vdd.n2623 gnd 0.006957f
C5449 vdd.n2624 gnd 0.006957f
C5450 vdd.n2625 gnd 0.006957f
C5451 vdd.n2626 gnd 0.006957f
C5452 vdd.n2627 gnd 0.006957f
C5453 vdd.n2628 gnd 0.006957f
C5454 vdd.n2629 gnd 0.006957f
C5455 vdd.n2630 gnd 0.491432f
C5456 vdd.n2631 gnd 0.006957f
C5457 vdd.n2632 gnd 0.006957f
C5458 vdd.n2633 gnd 0.006957f
C5459 vdd.n2634 gnd 0.006957f
C5460 vdd.n2635 gnd 0.006957f
C5461 vdd.n2636 gnd 0.006957f
C5462 vdd.n2637 gnd 0.44438f
C5463 vdd.n2638 gnd 0.006957f
C5464 vdd.n2639 gnd 0.006957f
C5465 vdd.n2640 gnd 0.006957f
C5466 vdd.n2641 gnd 0.015797f
C5467 vdd.n2642 gnd 0.014897f
C5468 vdd.n2643 gnd 0.006957f
C5469 vdd.n2644 gnd 0.006957f
C5470 vdd.n2645 gnd 0.005371f
C5471 vdd.n2646 gnd 0.006957f
C5472 vdd.n2647 gnd 0.006957f
C5473 vdd.n2648 gnd 0.005065f
C5474 vdd.n2649 gnd 0.006957f
C5475 vdd.n2650 gnd 0.006957f
C5476 vdd.n2651 gnd 0.006957f
C5477 vdd.n2652 gnd 0.006957f
C5478 vdd.n2653 gnd 0.006957f
C5479 vdd.n2654 gnd 0.006957f
C5480 vdd.n2655 gnd 0.006957f
C5481 vdd.n2656 gnd 0.006957f
C5482 vdd.n2657 gnd 0.006957f
C5483 vdd.n2658 gnd 0.006957f
C5484 vdd.n2659 gnd 0.006957f
C5485 vdd.n2660 gnd 0.006957f
C5486 vdd.n2661 gnd 0.006957f
C5487 vdd.n2662 gnd 0.006957f
C5488 vdd.n2663 gnd 0.006957f
C5489 vdd.n2664 gnd 0.006957f
C5490 vdd.n2665 gnd 0.006957f
C5491 vdd.n2666 gnd 0.006957f
C5492 vdd.n2667 gnd 0.006957f
C5493 vdd.n2668 gnd 0.006957f
C5494 vdd.n2669 gnd 0.006957f
C5495 vdd.n2670 gnd 0.006957f
C5496 vdd.n2671 gnd 0.006957f
C5497 vdd.n2672 gnd 0.006957f
C5498 vdd.n2673 gnd 0.006957f
C5499 vdd.n2674 gnd 0.006957f
C5500 vdd.n2675 gnd 0.006957f
C5501 vdd.n2676 gnd 0.006957f
C5502 vdd.n2677 gnd 0.006957f
C5503 vdd.n2678 gnd 0.006957f
C5504 vdd.n2679 gnd 0.006957f
C5505 vdd.n2680 gnd 0.006957f
C5506 vdd.n2681 gnd 0.006957f
C5507 vdd.n2682 gnd 0.006957f
C5508 vdd.n2683 gnd 0.006957f
C5509 vdd.n2684 gnd 0.006957f
C5510 vdd.n2685 gnd 0.006957f
C5511 vdd.n2686 gnd 0.006957f
C5512 vdd.n2687 gnd 0.006957f
C5513 vdd.n2688 gnd 0.006957f
C5514 vdd.n2689 gnd 0.006957f
C5515 vdd.n2690 gnd 0.006957f
C5516 vdd.n2691 gnd 0.006957f
C5517 vdd.n2692 gnd 0.006957f
C5518 vdd.n2693 gnd 0.006957f
C5519 vdd.n2694 gnd 0.006957f
C5520 vdd.n2695 gnd 0.006957f
C5521 vdd.n2696 gnd 0.006957f
C5522 vdd.n2697 gnd 0.006957f
C5523 vdd.n2698 gnd 0.006957f
C5524 vdd.n2699 gnd 0.006957f
C5525 vdd.n2700 gnd 0.006957f
C5526 vdd.n2701 gnd 0.006957f
C5527 vdd.n2702 gnd 0.006957f
C5528 vdd.n2703 gnd 0.006957f
C5529 vdd.n2704 gnd 0.006957f
C5530 vdd.n2705 gnd 0.006957f
C5531 vdd.n2706 gnd 0.006957f
C5532 vdd.n2707 gnd 0.006957f
C5533 vdd.n2708 gnd 0.006957f
C5534 vdd.n2709 gnd 0.015797f
C5535 vdd.n2710 gnd 0.014897f
C5536 vdd.n2711 gnd 0.014897f
C5537 vdd.n2712 gnd 0.805111f
C5538 vdd.n2713 gnd 0.014897f
C5539 vdd.n2714 gnd 0.015797f
C5540 vdd.n2715 gnd 0.014897f
C5541 vdd.n2716 gnd 0.006957f
C5542 vdd.n2717 gnd 0.006957f
C5543 vdd.n2718 gnd 0.006957f
C5544 vdd.n2719 gnd 0.005371f
C5545 vdd.n2720 gnd 0.009943f
C5546 vdd.n2721 gnd 0.005065f
C5547 vdd.n2722 gnd 0.006957f
C5548 vdd.n2723 gnd 0.006957f
C5549 vdd.n2724 gnd 0.006957f
C5550 vdd.n2725 gnd 0.006957f
C5551 vdd.n2726 gnd 0.006957f
C5552 vdd.n2727 gnd 0.006957f
C5553 vdd.n2728 gnd 0.006957f
C5554 vdd.n2729 gnd 0.006957f
C5555 vdd.n2730 gnd 0.006957f
C5556 vdd.n2731 gnd 0.006957f
C5557 vdd.n2732 gnd 0.006957f
C5558 vdd.n2733 gnd 0.006957f
C5559 vdd.n2734 gnd 0.006957f
C5560 vdd.n2735 gnd 0.006957f
C5561 vdd.n2736 gnd 0.006957f
C5562 vdd.n2737 gnd 0.006957f
C5563 vdd.n2738 gnd 0.006957f
C5564 vdd.n2739 gnd 0.006957f
C5565 vdd.n2740 gnd 0.006957f
C5566 vdd.n2741 gnd 0.006957f
C5567 vdd.n2742 gnd 0.006957f
C5568 vdd.n2743 gnd 0.006957f
C5569 vdd.n2744 gnd 0.006957f
C5570 vdd.n2745 gnd 0.006957f
C5571 vdd.n2746 gnd 0.006957f
C5572 vdd.n2747 gnd 0.006957f
C5573 vdd.n2748 gnd 0.006957f
C5574 vdd.n2749 gnd 0.006957f
C5575 vdd.n2750 gnd 0.006957f
C5576 vdd.n2751 gnd 0.006957f
C5577 vdd.n2752 gnd 0.006957f
C5578 vdd.n2753 gnd 0.006957f
C5579 vdd.n2754 gnd 0.006957f
C5580 vdd.n2755 gnd 0.006957f
C5581 vdd.n2756 gnd 0.006957f
C5582 vdd.n2757 gnd 0.006957f
C5583 vdd.n2758 gnd 0.006957f
C5584 vdd.n2759 gnd 0.006957f
C5585 vdd.n2760 gnd 0.006957f
C5586 vdd.n2761 gnd 0.006957f
C5587 vdd.n2762 gnd 0.006957f
C5588 vdd.n2763 gnd 0.006957f
C5589 vdd.n2764 gnd 0.006957f
C5590 vdd.n2765 gnd 0.006957f
C5591 vdd.n2766 gnd 0.006957f
C5592 vdd.n2767 gnd 0.006957f
C5593 vdd.n2768 gnd 0.006957f
C5594 vdd.n2769 gnd 0.006957f
C5595 vdd.n2770 gnd 0.006957f
C5596 vdd.n2771 gnd 0.006957f
C5597 vdd.n2772 gnd 0.006957f
C5598 vdd.n2773 gnd 0.006957f
C5599 vdd.n2774 gnd 0.006957f
C5600 vdd.n2775 gnd 0.006957f
C5601 vdd.n2776 gnd 0.006957f
C5602 vdd.n2777 gnd 0.006957f
C5603 vdd.n2778 gnd 0.006957f
C5604 vdd.n2779 gnd 0.006957f
C5605 vdd.n2780 gnd 0.006957f
C5606 vdd.n2781 gnd 0.006957f
C5607 vdd.n2782 gnd 0.015797f
C5608 vdd.n2783 gnd 0.015797f
C5609 vdd.n2784 gnd 0.867847f
C5610 vdd.t169 gnd 3.08452f
C5611 vdd.t156 gnd 3.08452f
C5612 vdd.n2818 gnd 0.015797f
C5613 vdd.t174 gnd 0.606448f
C5614 vdd.n2819 gnd 0.006957f
C5615 vdd.t286 gnd 0.281145f
C5616 vdd.t287 gnd 0.287787f
C5617 vdd.t284 gnd 0.183542f
C5618 vdd.n2820 gnd 0.099195f
C5619 vdd.n2821 gnd 0.056266f
C5620 vdd.n2822 gnd 0.006957f
C5621 vdd.t293 gnd 0.281145f
C5622 vdd.t294 gnd 0.287787f
C5623 vdd.t292 gnd 0.183542f
C5624 vdd.n2823 gnd 0.099195f
C5625 vdd.n2824 gnd 0.056266f
C5626 vdd.n2825 gnd 0.009943f
C5627 vdd.n2826 gnd 0.015797f
C5628 vdd.n2827 gnd 0.015797f
C5629 vdd.n2828 gnd 0.006957f
C5630 vdd.n2829 gnd 0.006957f
C5631 vdd.n2830 gnd 0.006957f
C5632 vdd.n2831 gnd 0.006957f
C5633 vdd.n2832 gnd 0.006957f
C5634 vdd.n2833 gnd 0.006957f
C5635 vdd.n2834 gnd 0.006957f
C5636 vdd.n2835 gnd 0.006957f
C5637 vdd.n2836 gnd 0.006957f
C5638 vdd.n2837 gnd 0.006957f
C5639 vdd.n2838 gnd 0.006957f
C5640 vdd.n2839 gnd 0.006957f
C5641 vdd.n2840 gnd 0.006957f
C5642 vdd.n2841 gnd 0.006957f
C5643 vdd.n2842 gnd 0.006957f
C5644 vdd.n2843 gnd 0.006957f
C5645 vdd.n2844 gnd 0.006957f
C5646 vdd.n2845 gnd 0.006957f
C5647 vdd.n2846 gnd 0.006957f
C5648 vdd.n2847 gnd 0.006957f
C5649 vdd.n2848 gnd 0.006957f
C5650 vdd.n2849 gnd 0.006957f
C5651 vdd.n2850 gnd 0.006957f
C5652 vdd.n2851 gnd 0.006957f
C5653 vdd.n2852 gnd 0.006957f
C5654 vdd.n2853 gnd 0.006957f
C5655 vdd.n2854 gnd 0.006957f
C5656 vdd.n2855 gnd 0.006957f
C5657 vdd.n2856 gnd 0.006957f
C5658 vdd.n2857 gnd 0.006957f
C5659 vdd.n2858 gnd 0.006957f
C5660 vdd.n2859 gnd 0.006957f
C5661 vdd.n2860 gnd 0.006957f
C5662 vdd.n2861 gnd 0.006957f
C5663 vdd.n2862 gnd 0.006957f
C5664 vdd.n2863 gnd 0.006957f
C5665 vdd.n2864 gnd 0.006957f
C5666 vdd.n2865 gnd 0.006957f
C5667 vdd.n2866 gnd 0.006957f
C5668 vdd.n2867 gnd 0.006957f
C5669 vdd.n2868 gnd 0.006957f
C5670 vdd.n2869 gnd 0.006957f
C5671 vdd.n2870 gnd 0.006957f
C5672 vdd.n2871 gnd 0.006957f
C5673 vdd.n2872 gnd 0.006957f
C5674 vdd.n2873 gnd 0.006957f
C5675 vdd.n2874 gnd 0.006957f
C5676 vdd.n2875 gnd 0.006957f
C5677 vdd.n2876 gnd 0.006957f
C5678 vdd.n2877 gnd 0.006957f
C5679 vdd.n2878 gnd 0.006957f
C5680 vdd.n2879 gnd 0.006957f
C5681 vdd.n2880 gnd 0.006957f
C5682 vdd.n2881 gnd 0.006957f
C5683 vdd.n2882 gnd 0.006957f
C5684 vdd.n2883 gnd 0.006957f
C5685 vdd.n2884 gnd 0.006957f
C5686 vdd.n2885 gnd 0.006957f
C5687 vdd.n2886 gnd 0.006957f
C5688 vdd.n2887 gnd 0.006957f
C5689 vdd.n2888 gnd 0.005065f
C5690 vdd.n2889 gnd 0.006957f
C5691 vdd.n2890 gnd 0.006957f
C5692 vdd.n2891 gnd 0.005371f
C5693 vdd.n2892 gnd 0.006957f
C5694 vdd.n2893 gnd 0.006957f
C5695 vdd.n2894 gnd 0.015797f
C5696 vdd.n2895 gnd 0.014897f
C5697 vdd.n2896 gnd 0.014897f
C5698 vdd.n2897 gnd 0.006957f
C5699 vdd.n2898 gnd 0.006957f
C5700 vdd.n2899 gnd 0.006957f
C5701 vdd.n2900 gnd 0.006957f
C5702 vdd.n2901 gnd 0.006957f
C5703 vdd.n2902 gnd 0.006957f
C5704 vdd.n2903 gnd 0.006957f
C5705 vdd.n2904 gnd 0.006957f
C5706 vdd.n2905 gnd 0.006957f
C5707 vdd.n2906 gnd 0.006957f
C5708 vdd.n2907 gnd 0.006957f
C5709 vdd.n2908 gnd 0.006957f
C5710 vdd.n2909 gnd 0.006957f
C5711 vdd.n2910 gnd 0.006957f
C5712 vdd.n2911 gnd 0.006957f
C5713 vdd.n2912 gnd 0.006957f
C5714 vdd.n2913 gnd 0.006957f
C5715 vdd.n2914 gnd 0.006957f
C5716 vdd.n2915 gnd 0.006957f
C5717 vdd.n2916 gnd 0.006957f
C5718 vdd.n2917 gnd 0.006957f
C5719 vdd.n2918 gnd 0.006957f
C5720 vdd.n2919 gnd 0.006957f
C5721 vdd.n2920 gnd 0.006957f
C5722 vdd.n2921 gnd 0.006957f
C5723 vdd.n2922 gnd 0.006957f
C5724 vdd.n2923 gnd 0.006957f
C5725 vdd.n2924 gnd 0.006957f
C5726 vdd.n2925 gnd 0.006957f
C5727 vdd.n2926 gnd 0.006957f
C5728 vdd.n2927 gnd 0.006957f
C5729 vdd.n2928 gnd 0.006957f
C5730 vdd.n2929 gnd 0.006957f
C5731 vdd.n2930 gnd 0.006957f
C5732 vdd.n2931 gnd 0.006957f
C5733 vdd.n2932 gnd 0.006957f
C5734 vdd.n2933 gnd 0.006957f
C5735 vdd.n2934 gnd 0.006957f
C5736 vdd.n2935 gnd 0.006957f
C5737 vdd.n2936 gnd 0.006957f
C5738 vdd.n2937 gnd 0.006957f
C5739 vdd.n2938 gnd 0.006957f
C5740 vdd.n2939 gnd 0.006957f
C5741 vdd.n2940 gnd 0.006957f
C5742 vdd.n2941 gnd 0.006957f
C5743 vdd.n2942 gnd 0.006957f
C5744 vdd.n2943 gnd 0.006957f
C5745 vdd.n2944 gnd 0.006957f
C5746 vdd.n2945 gnd 0.006957f
C5747 vdd.n2946 gnd 0.006957f
C5748 vdd.n2947 gnd 0.006957f
C5749 vdd.n2948 gnd 0.006957f
C5750 vdd.n2949 gnd 0.006957f
C5751 vdd.n2950 gnd 0.006957f
C5752 vdd.n2951 gnd 0.006957f
C5753 vdd.n2952 gnd 0.006957f
C5754 vdd.n2953 gnd 0.006957f
C5755 vdd.n2954 gnd 0.006957f
C5756 vdd.n2955 gnd 0.006957f
C5757 vdd.n2956 gnd 0.006957f
C5758 vdd.n2957 gnd 0.006957f
C5759 vdd.n2958 gnd 0.006957f
C5760 vdd.n2959 gnd 0.006957f
C5761 vdd.n2960 gnd 0.006957f
C5762 vdd.n2961 gnd 0.006957f
C5763 vdd.n2962 gnd 0.006957f
C5764 vdd.n2963 gnd 0.006957f
C5765 vdd.n2964 gnd 0.006957f
C5766 vdd.n2965 gnd 0.006957f
C5767 vdd.n2966 gnd 0.006957f
C5768 vdd.n2967 gnd 0.006957f
C5769 vdd.n2968 gnd 0.006957f
C5770 vdd.n2969 gnd 0.006957f
C5771 vdd.n2970 gnd 0.006957f
C5772 vdd.n2971 gnd 0.006957f
C5773 vdd.n2972 gnd 0.006957f
C5774 vdd.n2973 gnd 0.006957f
C5775 vdd.n2974 gnd 0.006957f
C5776 vdd.n2975 gnd 0.006957f
C5777 vdd.n2976 gnd 0.006957f
C5778 vdd.n2977 gnd 0.006957f
C5779 vdd.n2978 gnd 0.006957f
C5780 vdd.n2979 gnd 0.006957f
C5781 vdd.n2980 gnd 0.006957f
C5782 vdd.n2981 gnd 0.006957f
C5783 vdd.n2982 gnd 0.006957f
C5784 vdd.n2983 gnd 0.006957f
C5785 vdd.n2984 gnd 0.006957f
C5786 vdd.n2985 gnd 0.006957f
C5787 vdd.n2986 gnd 0.006957f
C5788 vdd.n2987 gnd 0.006957f
C5789 vdd.n2988 gnd 0.006957f
C5790 vdd.n2989 gnd 0.006957f
C5791 vdd.n2990 gnd 0.006957f
C5792 vdd.n2991 gnd 0.006957f
C5793 vdd.n2992 gnd 0.006957f
C5794 vdd.n2993 gnd 0.006957f
C5795 vdd.n2994 gnd 0.006957f
C5796 vdd.n2995 gnd 0.006957f
C5797 vdd.n2996 gnd 0.006957f
C5798 vdd.n2997 gnd 0.006957f
C5799 vdd.n2998 gnd 0.224804f
C5800 vdd.n2999 gnd 0.006957f
C5801 vdd.n3000 gnd 0.006957f
C5802 vdd.n3001 gnd 0.006957f
C5803 vdd.n3002 gnd 0.006957f
C5804 vdd.n3003 gnd 0.006957f
C5805 vdd.n3004 gnd 0.224804f
C5806 vdd.n3005 gnd 0.006957f
C5807 vdd.n3006 gnd 0.006957f
C5808 vdd.n3007 gnd 0.006957f
C5809 vdd.n3008 gnd 0.006957f
C5810 vdd.n3009 gnd 0.006957f
C5811 vdd.n3010 gnd 0.006957f
C5812 vdd.n3011 gnd 0.006957f
C5813 vdd.n3012 gnd 0.006957f
C5814 vdd.n3013 gnd 0.006957f
C5815 vdd.n3014 gnd 0.006957f
C5816 vdd.n3015 gnd 0.006957f
C5817 vdd.n3016 gnd 0.44438f
C5818 vdd.n3017 gnd 0.006957f
C5819 vdd.n3018 gnd 0.006957f
C5820 vdd.n3019 gnd 0.006957f
C5821 vdd.n3020 gnd 0.014897f
C5822 vdd.n3021 gnd 0.014897f
C5823 vdd.n3022 gnd 0.015797f
C5824 vdd.n3023 gnd 0.015797f
C5825 vdd.n3024 gnd 0.006957f
C5826 vdd.n3025 gnd 0.006957f
C5827 vdd.n3026 gnd 0.006957f
C5828 vdd.n3027 gnd 0.005371f
C5829 vdd.n3028 gnd 0.009943f
C5830 vdd.n3029 gnd 0.005065f
C5831 vdd.n3030 gnd 0.006957f
C5832 vdd.n3031 gnd 0.006957f
C5833 vdd.n3032 gnd 0.006957f
C5834 vdd.n3033 gnd 0.006957f
C5835 vdd.n3034 gnd 0.006957f
C5836 vdd.n3035 gnd 0.006957f
C5837 vdd.n3036 gnd 0.006957f
C5838 vdd.n3037 gnd 0.006957f
C5839 vdd.n3038 gnd 0.006957f
C5840 vdd.n3039 gnd 0.006957f
C5841 vdd.n3040 gnd 0.006957f
C5842 vdd.n3041 gnd 0.006957f
C5843 vdd.n3042 gnd 0.006957f
C5844 vdd.n3043 gnd 0.006957f
C5845 vdd.n3044 gnd 0.006957f
C5846 vdd.n3045 gnd 0.006957f
C5847 vdd.n3046 gnd 0.006957f
C5848 vdd.n3047 gnd 0.006957f
C5849 vdd.n3048 gnd 0.006957f
C5850 vdd.n3049 gnd 0.006957f
C5851 vdd.n3050 gnd 0.006957f
C5852 vdd.n3051 gnd 0.006957f
C5853 vdd.n3052 gnd 0.006957f
C5854 vdd.n3053 gnd 0.006957f
C5855 vdd.n3054 gnd 0.006957f
C5856 vdd.n3055 gnd 0.006957f
C5857 vdd.n3056 gnd 0.006957f
C5858 vdd.n3057 gnd 0.006957f
C5859 vdd.n3058 gnd 0.006957f
C5860 vdd.n3059 gnd 0.006957f
C5861 vdd.n3060 gnd 0.006957f
C5862 vdd.n3061 gnd 0.006957f
C5863 vdd.n3062 gnd 0.006957f
C5864 vdd.n3063 gnd 0.006957f
C5865 vdd.n3064 gnd 0.006957f
C5866 vdd.n3065 gnd 0.006957f
C5867 vdd.n3066 gnd 0.006957f
C5868 vdd.n3067 gnd 0.006957f
C5869 vdd.n3068 gnd 0.006957f
C5870 vdd.n3069 gnd 0.006957f
C5871 vdd.n3070 gnd 0.006957f
C5872 vdd.n3071 gnd 0.006957f
C5873 vdd.n3072 gnd 0.006957f
C5874 vdd.n3073 gnd 0.006957f
C5875 vdd.n3074 gnd 0.006957f
C5876 vdd.n3075 gnd 0.006957f
C5877 vdd.n3076 gnd 0.006957f
C5878 vdd.n3077 gnd 0.006957f
C5879 vdd.n3078 gnd 0.006957f
C5880 vdd.n3079 gnd 0.006957f
C5881 vdd.n3080 gnd 0.006957f
C5882 vdd.n3081 gnd 0.006957f
C5883 vdd.n3082 gnd 0.006957f
C5884 vdd.n3083 gnd 0.006957f
C5885 vdd.n3084 gnd 0.006957f
C5886 vdd.n3085 gnd 0.006957f
C5887 vdd.n3086 gnd 0.006957f
C5888 vdd.n3087 gnd 0.006957f
C5889 vdd.n3088 gnd 0.867847f
C5890 vdd.n3090 gnd 0.015797f
C5891 vdd.n3091 gnd 0.015797f
C5892 vdd.n3092 gnd 0.014897f
C5893 vdd.n3093 gnd 0.006957f
C5894 vdd.n3094 gnd 0.006957f
C5895 vdd.n3095 gnd 0.41824f
C5896 vdd.n3096 gnd 0.006957f
C5897 vdd.n3097 gnd 0.006957f
C5898 vdd.n3098 gnd 0.006957f
C5899 vdd.n3099 gnd 0.006957f
C5900 vdd.n3100 gnd 0.006957f
C5901 vdd.n3101 gnd 0.423468f
C5902 vdd.n3102 gnd 0.006957f
C5903 vdd.n3103 gnd 0.006957f
C5904 vdd.n3104 gnd 0.006957f
C5905 vdd.n3105 gnd 0.006957f
C5906 vdd.n3106 gnd 0.006957f
C5907 vdd.n3107 gnd 0.711008f
C5908 vdd.n3108 gnd 0.006957f
C5909 vdd.n3109 gnd 0.006957f
C5910 vdd.n3110 gnd 0.006957f
C5911 vdd.n3111 gnd 0.006957f
C5912 vdd.n3112 gnd 0.006957f
C5913 vdd.n3113 gnd 0.512344f
C5914 vdd.n3114 gnd 0.006957f
C5915 vdd.n3115 gnd 0.006957f
C5916 vdd.n3116 gnd 0.006957f
C5917 vdd.n3117 gnd 0.006957f
C5918 vdd.n3118 gnd 0.006957f
C5919 vdd.n3119 gnd 0.643044f
C5920 vdd.n3120 gnd 0.006957f
C5921 vdd.n3121 gnd 0.006957f
C5922 vdd.n3122 gnd 0.006957f
C5923 vdd.n3123 gnd 0.006957f
C5924 vdd.n3124 gnd 0.006957f
C5925 vdd.n3125 gnd 0.528028f
C5926 vdd.n3126 gnd 0.006957f
C5927 vdd.n3127 gnd 0.006957f
C5928 vdd.n3128 gnd 0.006957f
C5929 vdd.n3129 gnd 0.006957f
C5930 vdd.n3130 gnd 0.006957f
C5931 vdd.n3131 gnd 0.371188f
C5932 vdd.n3132 gnd 0.006957f
C5933 vdd.n3133 gnd 0.006957f
C5934 vdd.n3134 gnd 0.006957f
C5935 vdd.n3135 gnd 0.006957f
C5936 vdd.n3136 gnd 0.006957f
C5937 vdd.n3137 gnd 0.224804f
C5938 vdd.n3138 gnd 0.006957f
C5939 vdd.n3139 gnd 0.006957f
C5940 vdd.n3140 gnd 0.006957f
C5941 vdd.n3141 gnd 0.006957f
C5942 vdd.n3142 gnd 0.006957f
C5943 vdd.n3143 gnd 0.6535f
C5944 vdd.n3144 gnd 0.006957f
C5945 vdd.n3145 gnd 0.006957f
C5946 vdd.n3146 gnd 0.006957f
C5947 vdd.n3147 gnd 0.004911f
C5948 vdd.n3148 gnd 0.006957f
C5949 vdd.n3149 gnd 0.006957f
C5950 vdd.n3150 gnd 0.711008f
C5951 vdd.n3151 gnd 0.006957f
C5952 vdd.n3152 gnd 0.006957f
C5953 vdd.n3153 gnd 0.006957f
C5954 vdd.n3154 gnd 0.006957f
C5955 vdd.n3155 gnd 0.006957f
C5956 vdd.n3156 gnd 0.564624f
C5957 vdd.n3157 gnd 0.006957f
C5958 vdd.n3158 gnd 0.005525f
C5959 vdd.n3159 gnd 0.006957f
C5960 vdd.n3160 gnd 0.006957f
C5961 vdd.n3161 gnd 0.006957f
C5962 vdd.n3162 gnd 0.454836f
C5963 vdd.n3163 gnd 0.006957f
C5964 vdd.n3164 gnd 0.006957f
C5965 vdd.n3165 gnd 0.006957f
C5966 vdd.n3166 gnd 0.006957f
C5967 vdd.n3167 gnd 0.006957f
C5968 vdd.n3168 gnd 0.413012f
C5969 vdd.n3169 gnd 0.006957f
C5970 vdd.n3170 gnd 0.006957f
C5971 vdd.n3171 gnd 0.006957f
C5972 vdd.n3172 gnd 0.006957f
C5973 vdd.n3173 gnd 0.006957f
C5974 vdd.n3174 gnd 0.569852f
C5975 vdd.n3175 gnd 0.006957f
C5976 vdd.n3176 gnd 0.006957f
C5977 vdd.n3177 gnd 0.006957f
C5978 vdd.n3178 gnd 0.006957f
C5979 vdd.n3179 gnd 0.006957f
C5980 vdd.n3180 gnd 0.711008f
C5981 vdd.n3181 gnd 0.006957f
C5982 vdd.n3182 gnd 0.006957f
C5983 vdd.n3183 gnd 0.006957f
C5984 vdd.n3184 gnd 0.006957f
C5985 vdd.n3185 gnd 0.006957f
C5986 vdd.n3186 gnd 0.695324f
C5987 vdd.n3187 gnd 0.006957f
C5988 vdd.n3188 gnd 0.006957f
C5989 vdd.n3189 gnd 0.006957f
C5990 vdd.n3190 gnd 0.006957f
C5991 vdd.n3191 gnd 0.006957f
C5992 vdd.n3192 gnd 0.538484f
C5993 vdd.n3193 gnd 0.006957f
C5994 vdd.n3194 gnd 0.006957f
C5995 vdd.n3195 gnd 0.006957f
C5996 vdd.n3196 gnd 0.006957f
C5997 vdd.n3197 gnd 0.006957f
C5998 vdd.n3198 gnd 0.381644f
C5999 vdd.n3199 gnd 0.006957f
C6000 vdd.n3200 gnd 0.006957f
C6001 vdd.n3201 gnd 0.006957f
C6002 vdd.n3202 gnd 0.006957f
C6003 vdd.n3203 gnd 0.006957f
C6004 vdd.n3204 gnd 0.711008f
C6005 vdd.n3205 gnd 0.006957f
C6006 vdd.n3206 gnd 0.006957f
C6007 vdd.n3207 gnd 0.006957f
C6008 vdd.n3208 gnd 0.006957f
C6009 vdd.n3209 gnd 0.006957f
C6010 vdd.n3210 gnd 0.006957f
C6011 vdd.n3212 gnd 0.006957f
C6012 vdd.n3213 gnd 0.006957f
C6013 vdd.n3215 gnd 0.006957f
C6014 vdd.n3216 gnd 0.006957f
C6015 vdd.n3219 gnd 0.006957f
C6016 vdd.n3220 gnd 0.006957f
C6017 vdd.n3221 gnd 0.006957f
C6018 vdd.n3222 gnd 0.006957f
C6019 vdd.n3224 gnd 0.006957f
C6020 vdd.n3225 gnd 0.006957f
C6021 vdd.n3226 gnd 0.006957f
C6022 vdd.n3227 gnd 0.006957f
C6023 vdd.n3228 gnd 0.006957f
C6024 vdd.n3229 gnd 0.006957f
C6025 vdd.n3231 gnd 0.006957f
C6026 vdd.n3232 gnd 0.006957f
C6027 vdd.n3233 gnd 0.006957f
C6028 vdd.n3234 gnd 0.006957f
C6029 vdd.n3235 gnd 0.006957f
C6030 vdd.n3236 gnd 0.006957f
C6031 vdd.n3238 gnd 0.006957f
C6032 vdd.n3239 gnd 0.006957f
C6033 vdd.n3240 gnd 0.006957f
C6034 vdd.n3241 gnd 0.006957f
C6035 vdd.n3242 gnd 0.006957f
C6036 vdd.n3243 gnd 0.006957f
C6037 vdd.n3245 gnd 0.006957f
C6038 vdd.n3246 gnd 0.015797f
C6039 vdd.n3247 gnd 0.015797f
C6040 vdd.n3248 gnd 0.014897f
C6041 vdd.n3249 gnd 0.006957f
C6042 vdd.n3250 gnd 0.006957f
C6043 vdd.n3251 gnd 0.006957f
C6044 vdd.n3252 gnd 0.006957f
C6045 vdd.n3253 gnd 0.006957f
C6046 vdd.n3254 gnd 0.006957f
C6047 vdd.n3255 gnd 0.711008f
C6048 vdd.n3256 gnd 0.006957f
C6049 vdd.n3257 gnd 0.006957f
C6050 vdd.n3258 gnd 0.006957f
C6051 vdd.n3259 gnd 0.006957f
C6052 vdd.n3260 gnd 0.006957f
C6053 vdd.n3261 gnd 0.507116f
C6054 vdd.n3262 gnd 0.006957f
C6055 vdd.n3263 gnd 0.006957f
C6056 vdd.n3264 gnd 0.006957f
C6057 vdd.n3265 gnd 0.015797f
C6058 vdd.n3266 gnd 0.014897f
C6059 vdd.n3267 gnd 0.015797f
C6060 vdd.n3269 gnd 0.006957f
C6061 vdd.n3270 gnd 0.006957f
C6062 vdd.n3271 gnd 0.005371f
C6063 vdd.n3272 gnd 0.009943f
C6064 vdd.n3273 gnd 0.005065f
C6065 vdd.n3274 gnd 0.006957f
C6066 vdd.n3275 gnd 0.006957f
C6067 vdd.n3277 gnd 0.006957f
C6068 vdd.n3278 gnd 0.006957f
C6069 vdd.n3279 gnd 0.006957f
C6070 vdd.n3280 gnd 0.006957f
C6071 vdd.n3281 gnd 0.006957f
C6072 vdd.n3282 gnd 0.006957f
C6073 vdd.n3284 gnd 0.006957f
C6074 vdd.n3285 gnd 0.006957f
C6075 vdd.n3286 gnd 0.006957f
C6076 vdd.n3287 gnd 0.006957f
C6077 vdd.n3288 gnd 0.006957f
C6078 vdd.n3289 gnd 0.006957f
C6079 vdd.n3291 gnd 0.006957f
C6080 vdd.n3292 gnd 0.006957f
C6081 vdd.n3293 gnd 0.006957f
C6082 vdd.n3294 gnd 0.006957f
C6083 vdd.n3295 gnd 0.006957f
C6084 vdd.n3296 gnd 0.006957f
C6085 vdd.n3298 gnd 0.006957f
C6086 vdd.n3299 gnd 0.006957f
C6087 vdd.n3300 gnd 0.006957f
C6088 vdd.n3302 gnd 0.006957f
C6089 vdd.n3303 gnd 0.006957f
C6090 vdd.n3304 gnd 0.006957f
C6091 vdd.n3305 gnd 0.006957f
C6092 vdd.n3306 gnd 0.006957f
C6093 vdd.n3307 gnd 0.006957f
C6094 vdd.n3309 gnd 0.006957f
C6095 vdd.n3310 gnd 0.006957f
C6096 vdd.n3311 gnd 0.006957f
C6097 vdd.n3312 gnd 0.006957f
C6098 vdd.n3313 gnd 0.006957f
C6099 vdd.n3314 gnd 0.006957f
C6100 vdd.n3316 gnd 0.006957f
C6101 vdd.n3317 gnd 0.006957f
C6102 vdd.n3318 gnd 0.006957f
C6103 vdd.n3319 gnd 0.006957f
C6104 vdd.n3320 gnd 0.006957f
C6105 vdd.n3321 gnd 0.006957f
C6106 vdd.n3323 gnd 0.006957f
C6107 vdd.n3324 gnd 0.006957f
C6108 vdd.n3326 gnd 0.006957f
C6109 vdd.n3327 gnd 0.006957f
C6110 vdd.n3328 gnd 0.015797f
C6111 vdd.n3329 gnd 0.014897f
C6112 vdd.n3330 gnd 0.014897f
C6113 vdd.n3331 gnd 0.961951f
C6114 vdd.n3332 gnd 0.014897f
C6115 vdd.n3333 gnd 0.015797f
C6116 vdd.n3334 gnd 0.014897f
C6117 vdd.n3335 gnd 0.006957f
C6118 vdd.n3336 gnd 0.005371f
C6119 vdd.n3337 gnd 0.006957f
C6120 vdd.n3339 gnd 0.006957f
C6121 vdd.n3340 gnd 0.006957f
C6122 vdd.n3341 gnd 0.006957f
C6123 vdd.n3342 gnd 0.006957f
C6124 vdd.n3343 gnd 0.006957f
C6125 vdd.n3344 gnd 0.006957f
C6126 vdd.n3346 gnd 0.006957f
C6127 vdd.n3347 gnd 0.006957f
C6128 vdd.n3348 gnd 0.006957f
C6129 vdd.n3349 gnd 0.006957f
C6130 vdd.n3350 gnd 0.006957f
C6131 vdd.n3351 gnd 0.006957f
C6132 vdd.n3353 gnd 0.006957f
C6133 vdd.n3354 gnd 0.006957f
C6134 vdd.n3355 gnd 0.006957f
C6135 vdd.n3356 gnd 0.006957f
C6136 vdd.n3357 gnd 0.006957f
C6137 vdd.n3358 gnd 0.006957f
C6138 vdd.n3360 gnd 0.006957f
C6139 vdd.n3361 gnd 0.006957f
C6140 vdd.n3363 gnd 0.006957f
C6141 vdd.n3364 gnd 0.042961f
C6142 vdd.n3365 gnd 1.09007f
C6143 vdd.n3367 gnd 0.004323f
C6144 vdd.n3368 gnd 0.008235f
C6145 vdd.n3369 gnd 0.010231f
C6146 vdd.n3370 gnd 0.010231f
C6147 vdd.n3371 gnd 0.008235f
C6148 vdd.n3372 gnd 0.008235f
C6149 vdd.n3373 gnd 0.010231f
C6150 vdd.n3374 gnd 0.010231f
C6151 vdd.n3375 gnd 0.008235f
C6152 vdd.n3376 gnd 0.008235f
C6153 vdd.n3377 gnd 0.010231f
C6154 vdd.n3378 gnd 0.010231f
C6155 vdd.n3379 gnd 0.008235f
C6156 vdd.n3380 gnd 0.008235f
C6157 vdd.n3381 gnd 0.010231f
C6158 vdd.n3382 gnd 0.010231f
C6159 vdd.n3383 gnd 0.008235f
C6160 vdd.n3384 gnd 0.008235f
C6161 vdd.n3385 gnd 0.010231f
C6162 vdd.n3386 gnd 0.010231f
C6163 vdd.n3387 gnd 0.008235f
C6164 vdd.n3388 gnd 0.008235f
C6165 vdd.n3389 gnd 0.010231f
C6166 vdd.n3390 gnd 0.010231f
C6167 vdd.n3391 gnd 0.008235f
C6168 vdd.n3392 gnd 0.008235f
C6169 vdd.n3393 gnd 0.010231f
C6170 vdd.n3394 gnd 0.010231f
C6171 vdd.n3395 gnd 0.008235f
C6172 vdd.n3396 gnd 0.008235f
C6173 vdd.n3397 gnd 0.010231f
C6174 vdd.n3398 gnd 0.010231f
C6175 vdd.n3399 gnd 0.008235f
C6176 vdd.n3400 gnd 0.008235f
C6177 vdd.n3401 gnd 0.010231f
C6178 vdd.n3402 gnd 0.010231f
C6179 vdd.n3403 gnd 0.008235f
C6180 vdd.n3404 gnd 0.010231f
C6181 vdd.n3405 gnd 0.010231f
C6182 vdd.n3406 gnd 0.008235f
C6183 vdd.n3407 gnd 0.010231f
C6184 vdd.n3408 gnd 0.010231f
C6185 vdd.n3409 gnd 0.010231f
C6186 vdd.n3410 gnd 0.016799f
C6187 vdd.n3411 gnd 0.010231f
C6188 vdd.n3412 gnd 0.010231f
C6189 vdd.n3413 gnd 0.0056f
C6190 vdd.n3414 gnd 0.008235f
C6191 vdd.n3415 gnd 0.010231f
C6192 vdd.n3416 gnd 0.010231f
C6193 vdd.n3417 gnd 0.008235f
C6194 vdd.n3418 gnd 0.008235f
C6195 vdd.n3419 gnd 0.010231f
C6196 vdd.n3420 gnd 0.010231f
C6197 vdd.n3421 gnd 0.008235f
C6198 vdd.n3422 gnd 0.008235f
C6199 vdd.n3423 gnd 0.010231f
C6200 vdd.n3424 gnd 0.010231f
C6201 vdd.n3425 gnd 0.008235f
C6202 vdd.n3426 gnd 0.008235f
C6203 vdd.n3427 gnd 0.010231f
C6204 vdd.n3428 gnd 0.010231f
C6205 vdd.n3429 gnd 0.008235f
C6206 vdd.n3430 gnd 0.008235f
C6207 vdd.n3431 gnd 0.010231f
C6208 vdd.n3432 gnd 0.010231f
C6209 vdd.n3433 gnd 0.008235f
C6210 vdd.n3434 gnd 0.008235f
C6211 vdd.n3435 gnd 0.010231f
C6212 vdd.n3436 gnd 0.010231f
C6213 vdd.n3437 gnd 0.008235f
C6214 vdd.n3438 gnd 0.008235f
C6215 vdd.n3439 gnd 0.010231f
C6216 vdd.n3440 gnd 0.010231f
C6217 vdd.n3441 gnd 0.008235f
C6218 vdd.n3442 gnd 0.008235f
C6219 vdd.n3443 gnd 0.010231f
C6220 vdd.n3444 gnd 0.010231f
C6221 vdd.n3445 gnd 0.008235f
C6222 vdd.n3446 gnd 0.008235f
C6223 vdd.n3447 gnd 0.010231f
C6224 vdd.n3448 gnd 0.010231f
C6225 vdd.n3449 gnd 0.008235f
C6226 vdd.n3450 gnd 0.010231f
C6227 vdd.n3451 gnd 0.010231f
C6228 vdd.n3452 gnd 0.008235f
C6229 vdd.n3453 gnd 0.010231f
C6230 vdd.n3454 gnd 0.010231f
C6231 vdd.n3455 gnd 0.010231f
C6232 vdd.t282 gnd 0.125873f
C6233 vdd.t283 gnd 0.134524f
C6234 vdd.t281 gnd 0.164388f
C6235 vdd.n3456 gnd 0.210723f
C6236 vdd.n3457 gnd 0.177045f
C6237 vdd.n3458 gnd 0.016799f
C6238 vdd.n3459 gnd 0.010231f
C6239 vdd.n3460 gnd 0.010231f
C6240 vdd.n3461 gnd 0.006876f
C6241 vdd.n3462 gnd 0.008235f
C6242 vdd.n3463 gnd 0.010231f
C6243 vdd.n3464 gnd 0.010231f
C6244 vdd.n3465 gnd 0.008235f
C6245 vdd.n3466 gnd 0.008235f
C6246 vdd.n3467 gnd 0.010231f
C6247 vdd.n3468 gnd 0.010231f
C6248 vdd.n3469 gnd 0.008235f
C6249 vdd.n3470 gnd 0.008235f
C6250 vdd.n3471 gnd 0.010231f
C6251 vdd.n3472 gnd 0.010231f
C6252 vdd.n3473 gnd 0.008235f
C6253 vdd.n3474 gnd 0.008235f
C6254 vdd.n3475 gnd 0.010231f
C6255 vdd.n3476 gnd 0.010231f
C6256 vdd.n3477 gnd 0.008235f
C6257 vdd.n3478 gnd 0.008235f
C6258 vdd.n3479 gnd 0.010231f
C6259 vdd.n3480 gnd 0.010231f
C6260 vdd.n3481 gnd 0.008235f
C6261 vdd.n3482 gnd 0.008235f
C6262 vdd.n3483 gnd 0.010231f
C6263 vdd.n3484 gnd 0.010231f
C6264 vdd.n3485 gnd 0.008235f
C6265 vdd.n3486 gnd 0.008235f
C6266 vdd.n3488 gnd 1.09007f
C6267 vdd.n3490 gnd 0.008235f
C6268 vdd.n3491 gnd 0.008235f
C6269 vdd.n3492 gnd 0.006835f
C6270 vdd.n3493 gnd 0.025281f
C6271 vdd.n3495 gnd 12.7668f
C6272 vdd.n3496 gnd 0.025281f
C6273 vdd.n3497 gnd 0.003912f
C6274 vdd.n3498 gnd 0.025281f
C6275 vdd.n3499 gnd 0.024751f
C6276 vdd.n3500 gnd 0.010231f
C6277 vdd.n3501 gnd 0.008235f
C6278 vdd.n3502 gnd 0.010231f
C6279 vdd.n3503 gnd 0.632588f
C6280 vdd.n3504 gnd 0.010231f
C6281 vdd.n3505 gnd 0.008235f
C6282 vdd.n3506 gnd 0.010231f
C6283 vdd.n3507 gnd 0.010231f
C6284 vdd.n3508 gnd 0.010231f
C6285 vdd.n3509 gnd 0.008235f
C6286 vdd.n3510 gnd 0.010231f
C6287 vdd.n3511 gnd 1.0456f
C6288 vdd.n3512 gnd 0.010231f
C6289 vdd.n3513 gnd 0.008235f
C6290 vdd.n3514 gnd 0.010231f
C6291 vdd.n3515 gnd 0.010231f
C6292 vdd.n3516 gnd 0.010231f
C6293 vdd.n3517 gnd 0.008235f
C6294 vdd.n3518 gnd 0.010231f
C6295 vdd.n3519 gnd 0.674412f
C6296 vdd.n3520 gnd 0.716236f
C6297 vdd.n3521 gnd 0.010231f
C6298 vdd.n3522 gnd 0.008235f
C6299 vdd.n3523 gnd 0.010231f
C6300 vdd.n3524 gnd 0.010231f
C6301 vdd.n3525 gnd 0.010231f
C6302 vdd.n3526 gnd 0.008235f
C6303 vdd.n3527 gnd 0.010231f
C6304 vdd.n3528 gnd 0.867847f
C6305 vdd.n3529 gnd 0.010231f
C6306 vdd.n3530 gnd 0.008235f
C6307 vdd.n3531 gnd 0.010231f
C6308 vdd.n3532 gnd 0.010231f
C6309 vdd.n3533 gnd 0.010231f
C6310 vdd.n3534 gnd 0.008235f
C6311 vdd.n3535 gnd 0.010231f
C6312 vdd.t109 gnd 0.5228f
C6313 vdd.n3536 gnd 0.841707f
C6314 vdd.n3537 gnd 0.010231f
C6315 vdd.n3538 gnd 0.008235f
C6316 vdd.n3539 gnd 0.010231f
C6317 vdd.n3540 gnd 0.010231f
C6318 vdd.n3541 gnd 0.010231f
C6319 vdd.n3542 gnd 0.008235f
C6320 vdd.n3543 gnd 0.010231f
C6321 vdd.n3544 gnd 0.663956f
C6322 vdd.n3545 gnd 0.010231f
C6323 vdd.n3546 gnd 0.008235f
C6324 vdd.n3547 gnd 0.010231f
C6325 vdd.n3548 gnd 0.010231f
C6326 vdd.n3549 gnd 0.010231f
C6327 vdd.n3550 gnd 0.008235f
C6328 vdd.n3551 gnd 0.010231f
C6329 vdd.n3552 gnd 0.831251f
C6330 vdd.n3553 gnd 0.559396f
C6331 vdd.n3554 gnd 0.010231f
C6332 vdd.n3555 gnd 0.008235f
C6333 vdd.n3556 gnd 0.010231f
C6334 vdd.n3557 gnd 0.010231f
C6335 vdd.n3558 gnd 0.010231f
C6336 vdd.n3559 gnd 0.008235f
C6337 vdd.n3560 gnd 0.010231f
C6338 vdd.n3561 gnd 0.737148f
C6339 vdd.n3562 gnd 0.010231f
C6340 vdd.n3563 gnd 0.008235f
C6341 vdd.n3564 gnd 0.010231f
C6342 vdd.n3565 gnd 0.010231f
C6343 vdd.n3566 gnd 0.010231f
C6344 vdd.n3567 gnd 0.010231f
C6345 vdd.n3568 gnd 0.010231f
C6346 vdd.n3569 gnd 0.008235f
C6347 vdd.n3570 gnd 0.008235f
C6348 vdd.n3571 gnd 0.010231f
C6349 vdd.t27 gnd 0.5228f
C6350 vdd.n3572 gnd 0.867847f
C6351 vdd.n3573 gnd 0.010231f
C6352 vdd.n3574 gnd 0.008235f
C6353 vdd.n3575 gnd 0.010231f
C6354 vdd.n3576 gnd 0.010231f
C6355 vdd.n3577 gnd 0.010231f
C6356 vdd.n3578 gnd 0.008235f
C6357 vdd.n3579 gnd 0.010231f
C6358 vdd.n3580 gnd 0.820795f
C6359 vdd.n3581 gnd 0.010231f
C6360 vdd.n3582 gnd 0.010231f
C6361 vdd.n3583 gnd 0.008235f
C6362 vdd.n3584 gnd 0.008235f
C6363 vdd.n3585 gnd 0.010231f
C6364 vdd.n3586 gnd 0.010231f
C6365 vdd.n3587 gnd 0.010231f
C6366 vdd.n3588 gnd 0.008235f
C6367 vdd.n3589 gnd 0.010231f
C6368 vdd.n3590 gnd 0.008235f
C6369 vdd.n3591 gnd 0.008235f
C6370 vdd.n3592 gnd 0.010231f
C6371 vdd.n3593 gnd 0.010231f
C6372 vdd.n3594 gnd 0.010231f
C6373 vdd.n3595 gnd 0.008235f
C6374 vdd.n3596 gnd 0.010231f
C6375 vdd.n3597 gnd 0.008235f
C6376 vdd.n3598 gnd 0.008235f
C6377 vdd.n3599 gnd 0.010231f
C6378 vdd.n3600 gnd 0.010231f
C6379 vdd.n3601 gnd 0.010231f
C6380 vdd.n3602 gnd 0.008235f
C6381 vdd.n3603 gnd 0.867847f
C6382 vdd.n3604 gnd 0.010231f
C6383 vdd.n3605 gnd 0.008235f
C6384 vdd.n3606 gnd 0.008235f
C6385 vdd.n3607 gnd 0.010231f
C6386 vdd.n3608 gnd 0.010231f
C6387 vdd.n3609 gnd 0.010231f
C6388 vdd.n3610 gnd 0.008235f
C6389 vdd.n3611 gnd 0.010231f
C6390 vdd.n3612 gnd 0.008235f
C6391 vdd.n3613 gnd 0.008235f
C6392 vdd.n3614 gnd 0.010231f
C6393 vdd.n3615 gnd 0.010231f
C6394 vdd.n3616 gnd 0.010231f
C6395 vdd.n3617 gnd 0.008235f
C6396 vdd.n3618 gnd 0.010231f
C6397 vdd.n3619 gnd 0.008235f
C6398 vdd.n3620 gnd 0.006835f
C6399 vdd.n3621 gnd 0.024751f
C6400 vdd.n3622 gnd 0.025281f
C6401 vdd.n3623 gnd 0.003912f
C6402 vdd.n3624 gnd 0.025281f
C6403 vdd.n3626 gnd 2.47807f
C6404 vdd.n3627 gnd 1.54226f
C6405 vdd.n3628 gnd 0.024751f
C6406 vdd.n3629 gnd 0.006835f
C6407 vdd.n3630 gnd 0.008235f
C6408 vdd.n3631 gnd 0.008235f
C6409 vdd.n3632 gnd 0.010231f
C6410 vdd.n3633 gnd 1.0456f
C6411 vdd.n3634 gnd 1.0456f
C6412 vdd.n3635 gnd 0.956723f
C6413 vdd.n3636 gnd 0.010231f
C6414 vdd.n3637 gnd 0.008235f
C6415 vdd.n3638 gnd 0.008235f
C6416 vdd.n3639 gnd 0.008235f
C6417 vdd.n3640 gnd 0.010231f
C6418 vdd.n3641 gnd 0.778971f
C6419 vdd.t25 gnd 0.5228f
C6420 vdd.n3642 gnd 0.789427f
C6421 vdd.n3643 gnd 0.60122f
C6422 vdd.n3644 gnd 0.010231f
C6423 vdd.n3645 gnd 0.008235f
C6424 vdd.n3646 gnd 0.008235f
C6425 vdd.n3647 gnd 0.008235f
C6426 vdd.n3648 gnd 0.010231f
C6427 vdd.n3649 gnd 0.622132f
C6428 vdd.n3650 gnd 0.768516f
C6429 vdd.t97 gnd 0.5228f
C6430 vdd.n3651 gnd 0.799883f
C6431 vdd.n3652 gnd 0.010231f
C6432 vdd.n3653 gnd 0.008235f
C6433 vdd.n3654 gnd 0.008235f
C6434 vdd.n3655 gnd 0.008235f
C6435 vdd.n3656 gnd 0.010231f
C6436 vdd.n3657 gnd 0.867847f
C6437 vdd.t104 gnd 0.5228f
C6438 vdd.n3658 gnd 0.632588f
C6439 vdd.n3659 gnd 0.75806f
C6440 vdd.n3660 gnd 0.010231f
C6441 vdd.n3661 gnd 0.008235f
C6442 vdd.n3662 gnd 0.008235f
C6443 vdd.n3663 gnd 0.008235f
C6444 vdd.n3664 gnd 0.010231f
C6445 vdd.n3665 gnd 0.580308f
C6446 vdd.t120 gnd 0.5228f
C6447 vdd.n3666 gnd 0.867847f
C6448 vdd.t29 gnd 0.5228f
C6449 vdd.n3667 gnd 0.643044f
C6450 vdd.n3668 gnd 0.010231f
C6451 vdd.n3669 gnd 0.008235f
C6452 vdd.n3670 gnd 0.007863f
C6453 vdd.n3671 gnd 0.603486f
C6454 vdd.n3672 gnd 2.98812f
C6455 a_n2804_13878.t23 gnd 0.194878f
C6456 a_n2804_13878.t10 gnd 0.194878f
C6457 a_n2804_13878.t20 gnd 0.194878f
C6458 a_n2804_13878.n0 gnd 1.53612f
C6459 a_n2804_13878.t25 gnd 0.194878f
C6460 a_n2804_13878.t15 gnd 0.194878f
C6461 a_n2804_13878.n1 gnd 1.5345f
C6462 a_n2804_13878.n2 gnd 2.14416f
C6463 a_n2804_13878.t21 gnd 0.194878f
C6464 a_n2804_13878.t14 gnd 0.194878f
C6465 a_n2804_13878.n3 gnd 1.5345f
C6466 a_n2804_13878.n4 gnd 1.04587f
C6467 a_n2804_13878.t8 gnd 0.194878f
C6468 a_n2804_13878.t11 gnd 0.194878f
C6469 a_n2804_13878.n5 gnd 1.5345f
C6470 a_n2804_13878.n6 gnd 1.04587f
C6471 a_n2804_13878.t24 gnd 0.194878f
C6472 a_n2804_13878.t9 gnd 0.194878f
C6473 a_n2804_13878.n7 gnd 1.5345f
C6474 a_n2804_13878.n8 gnd 1.04587f
C6475 a_n2804_13878.t19 gnd 0.194878f
C6476 a_n2804_13878.t7 gnd 0.194878f
C6477 a_n2804_13878.n9 gnd 1.5345f
C6478 a_n2804_13878.n10 gnd 4.90989f
C6479 a_n2804_13878.t30 gnd 1.82474f
C6480 a_n2804_13878.t3 gnd 0.194878f
C6481 a_n2804_13878.t4 gnd 0.194878f
C6482 a_n2804_13878.n11 gnd 1.37272f
C6483 a_n2804_13878.n12 gnd 1.53381f
C6484 a_n2804_13878.t5 gnd 1.8211f
C6485 a_n2804_13878.n13 gnd 0.771835f
C6486 a_n2804_13878.t1 gnd 1.8211f
C6487 a_n2804_13878.n14 gnd 0.771835f
C6488 a_n2804_13878.t2 gnd 0.194878f
C6489 a_n2804_13878.t0 gnd 0.194878f
C6490 a_n2804_13878.n15 gnd 1.37272f
C6491 a_n2804_13878.n16 gnd 0.77931f
C6492 a_n2804_13878.t31 gnd 1.8211f
C6493 a_n2804_13878.n17 gnd 2.86287f
C6494 a_n2804_13878.n18 gnd 3.75497f
C6495 a_n2804_13878.t13 gnd 0.194878f
C6496 a_n2804_13878.t22 gnd 0.194878f
C6497 a_n2804_13878.n19 gnd 1.53449f
C6498 a_n2804_13878.n20 gnd 2.50654f
C6499 a_n2804_13878.t26 gnd 0.194878f
C6500 a_n2804_13878.t12 gnd 0.194878f
C6501 a_n2804_13878.n21 gnd 1.5345f
C6502 a_n2804_13878.n22 gnd 0.679894f
C6503 a_n2804_13878.t16 gnd 0.194878f
C6504 a_n2804_13878.t17 gnd 0.194878f
C6505 a_n2804_13878.n23 gnd 1.5345f
C6506 a_n2804_13878.n24 gnd 0.679894f
C6507 a_n2804_13878.t27 gnd 0.194878f
C6508 a_n2804_13878.t28 gnd 0.194878f
C6509 a_n2804_13878.n25 gnd 1.5345f
C6510 a_n2804_13878.n26 gnd 0.679894f
C6511 a_n2804_13878.t6 gnd 0.194878f
C6512 a_n2804_13878.t18 gnd 0.194878f
C6513 a_n2804_13878.n27 gnd 1.5345f
C6514 a_n2804_13878.n28 gnd 1.37932f
C6515 a_n2804_13878.n29 gnd 1.53704f
C6516 a_n2804_13878.t29 gnd 0.194878f
C6517 a_n2982_13878.n0 gnd 0.930299f
C6518 a_n2982_13878.n1 gnd 0.204505f
C6519 a_n2982_13878.n2 gnd 0.150622f
C6520 a_n2982_13878.n3 gnd 0.23673f
C6521 a_n2982_13878.n4 gnd 0.182847f
C6522 a_n2982_13878.n5 gnd 0.204505f
C6523 a_n2982_13878.n6 gnd 0.150622f
C6524 a_n2982_13878.n7 gnd 0.984182f
C6525 a_n2982_13878.n8 gnd 0.215533f
C6526 a_n2982_13878.n9 gnd 0.758602f
C6527 a_n2982_13878.n10 gnd 0.215533f
C6528 a_n2982_13878.n11 gnd 0.215533f
C6529 a_n2982_13878.n12 gnd 0.490874f
C6530 a_n2982_13878.n13 gnd 0.282596f
C6531 a_n2982_13878.n14 gnd 0.215533f
C6532 a_n2982_13878.n15 gnd 0.544757f
C6533 a_n2982_13878.n16 gnd 0.215533f
C6534 a_n2982_13878.n17 gnd 0.215533f
C6535 a_n2982_13878.n18 gnd 0.958966f
C6536 a_n2982_13878.n19 gnd 0.282596f
C6537 a_n2982_13878.n20 gnd 3.20753f
C6538 a_n2982_13878.n21 gnd 0.215533f
C6539 a_n2982_13878.n22 gnd 0.215533f
C6540 a_n2982_13878.n23 gnd 0.868451f
C6541 a_n2982_13878.n24 gnd 0.215533f
C6542 a_n2982_13878.n25 gnd 0.282596f
C6543 a_n2982_13878.n26 gnd 1.00004f
C6544 a_n2982_13878.n27 gnd 0.215533f
C6545 a_n2982_13878.n28 gnd 0.215533f
C6546 a_n2982_13878.n29 gnd 0.490874f
C6547 a_n2982_13878.n30 gnd 0.215533f
C6548 a_n2982_13878.n31 gnd 0.282596f
C6549 a_n2982_13878.n32 gnd 3.4865f
C6550 a_n2982_13878.n33 gnd 2.65557f
C6551 a_n2982_13878.n34 gnd 3.74061f
C6552 a_n2982_13878.n35 gnd 1.19566f
C6553 a_n2982_13878.n36 gnd 2.1833f
C6554 a_n2982_13878.n37 gnd 1.77446f
C6555 a_n2982_13878.n38 gnd 1.77446f
C6556 a_n2982_13878.n39 gnd 2.38801f
C6557 a_n2982_13878.n40 gnd 1.19566f
C6558 a_n2982_13878.n41 gnd 0.725631f
C6559 a_n2982_13878.n42 gnd 0.725634f
C6560 a_n2982_13878.n43 gnd 0.008648f
C6561 a_n2982_13878.n44 gnd 4.17e-19
C6562 a_n2982_13878.n46 gnd 0.008345f
C6563 a_n2982_13878.n47 gnd 0.012134f
C6564 a_n2982_13878.n48 gnd 0.008028f
C6565 a_n2982_13878.n50 gnd 1.69354f
C6566 a_n2982_13878.n51 gnd 0.285885f
C6567 a_n2982_13878.n52 gnd 0.008648f
C6568 a_n2982_13878.n53 gnd 4.17e-19
C6569 a_n2982_13878.n55 gnd 0.008345f
C6570 a_n2982_13878.n56 gnd 0.012134f
C6571 a_n2982_13878.n57 gnd 0.008028f
C6572 a_n2982_13878.n59 gnd 0.008648f
C6573 a_n2982_13878.n60 gnd 4.17e-19
C6574 a_n2982_13878.n62 gnd 0.008345f
C6575 a_n2982_13878.n63 gnd 0.012134f
C6576 a_n2982_13878.n64 gnd 0.008028f
C6577 a_n2982_13878.n66 gnd 0.285885f
C6578 a_n2982_13878.n67 gnd 0.008648f
C6579 a_n2982_13878.n68 gnd 4.17e-19
C6580 a_n2982_13878.n70 gnd 0.008345f
C6581 a_n2982_13878.n71 gnd 0.012134f
C6582 a_n2982_13878.n72 gnd 0.008028f
C6583 a_n2982_13878.n74 gnd 0.285885f
C6584 a_n2982_13878.n75 gnd 0.008345f
C6585 a_n2982_13878.n76 gnd 0.284719f
C6586 a_n2982_13878.n77 gnd 0.008345f
C6587 a_n2982_13878.n78 gnd 0.284719f
C6588 a_n2982_13878.n79 gnd 0.008345f
C6589 a_n2982_13878.n80 gnd 0.284719f
C6590 a_n2982_13878.n81 gnd 0.008345f
C6591 a_n2982_13878.n82 gnd 0.284719f
C6592 a_n2982_13878.n83 gnd 0.285885f
C6593 a_n2982_13878.t55 gnd 0.149496f
C6594 a_n2982_13878.t51 gnd 1.39981f
C6595 a_n2982_13878.t53 gnd 0.149496f
C6596 a_n2982_13878.t29 gnd 0.149496f
C6597 a_n2982_13878.n84 gnd 1.05305f
C6598 a_n2982_13878.t25 gnd 0.149496f
C6599 a_n2982_13878.t57 gnd 0.149496f
C6600 a_n2982_13878.n85 gnd 1.05305f
C6601 a_n2982_13878.t36 gnd 0.695384f
C6602 a_n2982_13878.n86 gnd 0.305719f
C6603 a_n2982_13878.t64 gnd 0.695384f
C6604 a_n2982_13878.t48 gnd 0.695384f
C6605 a_n2982_13878.n87 gnd 0.296537f
C6606 a_n2982_13878.t56 gnd 0.695384f
C6607 a_n2982_13878.n88 gnd 0.308347f
C6608 a_n2982_13878.t54 gnd 0.695384f
C6609 a_n2982_13878.t28 gnd 0.695384f
C6610 a_n2982_13878.n89 gnd 0.30152f
C6611 a_n2982_13878.t50 gnd 0.70986f
C6612 a_n2982_13878.t86 gnd 0.695384f
C6613 a_n2982_13878.n90 gnd 0.305719f
C6614 a_n2982_13878.t95 gnd 0.695384f
C6615 a_n2982_13878.t101 gnd 0.695384f
C6616 a_n2982_13878.n91 gnd 0.296537f
C6617 a_n2982_13878.t105 gnd 0.695384f
C6618 a_n2982_13878.n92 gnd 0.308347f
C6619 a_n2982_13878.t76 gnd 0.695384f
C6620 a_n2982_13878.t79 gnd 0.695384f
C6621 a_n2982_13878.n93 gnd 0.30152f
C6622 a_n2982_13878.t109 gnd 0.70986f
C6623 a_n2982_13878.t44 gnd 0.70986f
C6624 a_n2982_13878.t32 gnd 0.695384f
C6625 a_n2982_13878.t60 gnd 0.695384f
C6626 a_n2982_13878.t40 gnd 0.695384f
C6627 a_n2982_13878.n94 gnd 0.305597f
C6628 a_n2982_13878.t22 gnd 0.695384f
C6629 a_n2982_13878.t30 gnd 0.695384f
C6630 a_n2982_13878.t66 gnd 0.695384f
C6631 a_n2982_13878.n95 gnd 0.301852f
C6632 a_n2982_13878.t42 gnd 0.695384f
C6633 a_n2982_13878.t62 gnd 0.695384f
C6634 a_n2982_13878.t34 gnd 0.695384f
C6635 a_n2982_13878.n96 gnd 0.305719f
C6636 a_n2982_13878.t26 gnd 0.695384f
C6637 a_n2982_13878.t38 gnd 0.70657f
C6638 a_n2982_13878.t69 gnd 0.116275f
C6639 a_n2982_13878.t15 gnd 0.116275f
C6640 a_n2982_13878.n97 gnd 1.02908f
C6641 a_n2982_13878.t5 gnd 0.116275f
C6642 a_n2982_13878.t4 gnd 0.116275f
C6643 a_n2982_13878.n98 gnd 1.02744f
C6644 a_n2982_13878.t12 gnd 0.116275f
C6645 a_n2982_13878.t3 gnd 0.116275f
C6646 a_n2982_13878.n99 gnd 1.02744f
C6647 a_n2982_13878.t7 gnd 0.116275f
C6648 a_n2982_13878.t0 gnd 0.116275f
C6649 a_n2982_13878.n100 gnd 1.02908f
C6650 a_n2982_13878.t71 gnd 0.116275f
C6651 a_n2982_13878.t14 gnd 0.116275f
C6652 a_n2982_13878.n101 gnd 1.02744f
C6653 a_n2982_13878.t17 gnd 0.116275f
C6654 a_n2982_13878.t13 gnd 0.116275f
C6655 a_n2982_13878.n102 gnd 1.02744f
C6656 a_n2982_13878.t9 gnd 0.116275f
C6657 a_n2982_13878.t70 gnd 0.116275f
C6658 a_n2982_13878.n103 gnd 1.02744f
C6659 a_n2982_13878.t2 gnd 0.116275f
C6660 a_n2982_13878.t6 gnd 0.116275f
C6661 a_n2982_13878.n104 gnd 1.02744f
C6662 a_n2982_13878.t16 gnd 0.116275f
C6663 a_n2982_13878.t11 gnd 0.116275f
C6664 a_n2982_13878.n105 gnd 1.02744f
C6665 a_n2982_13878.t19 gnd 0.116275f
C6666 a_n2982_13878.t8 gnd 0.116275f
C6667 a_n2982_13878.n106 gnd 1.02908f
C6668 a_n2982_13878.t18 gnd 0.116275f
C6669 a_n2982_13878.t10 gnd 0.116275f
C6670 a_n2982_13878.n107 gnd 1.02744f
C6671 a_n2982_13878.t1 gnd 0.116275f
C6672 a_n2982_13878.t68 gnd 0.116275f
C6673 a_n2982_13878.n108 gnd 1.02744f
C6674 a_n2982_13878.t110 gnd 0.70986f
C6675 a_n2982_13878.t87 gnd 0.695384f
C6676 a_n2982_13878.t92 gnd 0.695384f
C6677 a_n2982_13878.t80 gnd 0.695384f
C6678 a_n2982_13878.n109 gnd 0.305597f
C6679 a_n2982_13878.t97 gnd 0.695384f
C6680 a_n2982_13878.t106 gnd 0.695384f
C6681 a_n2982_13878.t107 gnd 0.695384f
C6682 a_n2982_13878.n110 gnd 0.301852f
C6683 a_n2982_13878.t74 gnd 0.695384f
C6684 a_n2982_13878.t89 gnd 0.695384f
C6685 a_n2982_13878.t77 gnd 0.695384f
C6686 a_n2982_13878.n111 gnd 0.305719f
C6687 a_n2982_13878.t84 gnd 0.695384f
C6688 a_n2982_13878.t103 gnd 0.70657f
C6689 a_n2982_13878.n112 gnd 0.307896f
C6690 a_n2982_13878.n113 gnd 0.302112f
C6691 a_n2982_13878.n114 gnd 0.296537f
C6692 a_n2982_13878.n115 gnd 0.305735f
C6693 a_n2982_13878.n116 gnd 0.308347f
C6694 a_n2982_13878.n117 gnd 0.30152f
C6695 a_n2982_13878.n118 gnd 0.307896f
C6696 a_n2982_13878.n119 gnd 0.307896f
C6697 a_n2982_13878.n120 gnd 0.302112f
C6698 a_n2982_13878.n121 gnd 0.296537f
C6699 a_n2982_13878.n122 gnd 0.305735f
C6700 a_n2982_13878.n123 gnd 0.308347f
C6701 a_n2982_13878.n124 gnd 0.30152f
C6702 a_n2982_13878.n125 gnd 0.307896f
C6703 a_n2982_13878.t39 gnd 1.39981f
C6704 a_n2982_13878.t35 gnd 0.149496f
C6705 a_n2982_13878.t27 gnd 0.149496f
C6706 a_n2982_13878.n126 gnd 1.05305f
C6707 a_n2982_13878.t43 gnd 0.149496f
C6708 a_n2982_13878.t63 gnd 0.149496f
C6709 a_n2982_13878.n127 gnd 1.05305f
C6710 a_n2982_13878.t31 gnd 0.149496f
C6711 a_n2982_13878.t67 gnd 0.149496f
C6712 a_n2982_13878.n128 gnd 1.05305f
C6713 a_n2982_13878.t41 gnd 0.149496f
C6714 a_n2982_13878.t23 gnd 0.149496f
C6715 a_n2982_13878.n129 gnd 1.05305f
C6716 a_n2982_13878.t33 gnd 0.149496f
C6717 a_n2982_13878.t61 gnd 0.149496f
C6718 a_n2982_13878.n130 gnd 1.05305f
C6719 a_n2982_13878.t45 gnd 1.39702f
C6720 a_n2982_13878.n131 gnd 1.0237f
C6721 a_n2982_13878.t85 gnd 0.695384f
C6722 a_n2982_13878.t96 gnd 0.695384f
C6723 a_n2982_13878.t111 gnd 0.695384f
C6724 a_n2982_13878.n132 gnd 0.305735f
C6725 a_n2982_13878.t98 gnd 0.695384f
C6726 a_n2982_13878.t81 gnd 0.695384f
C6727 a_n2982_13878.t82 gnd 0.695384f
C6728 a_n2982_13878.n133 gnd 0.305735f
C6729 a_n2982_13878.t102 gnd 0.695384f
C6730 a_n2982_13878.t91 gnd 0.695384f
C6731 a_n2982_13878.t90 gnd 0.695384f
C6732 a_n2982_13878.n134 gnd 0.305735f
C6733 a_n2982_13878.t94 gnd 0.695384f
C6734 a_n2982_13878.t83 gnd 0.695384f
C6735 a_n2982_13878.t72 gnd 0.695384f
C6736 a_n2982_13878.n135 gnd 0.305735f
C6737 a_n2982_13878.t99 gnd 0.707035f
C6738 a_n2982_13878.n136 gnd 0.301852f
C6739 a_n2982_13878.n137 gnd 0.296371f
C6740 a_n2982_13878.t108 gnd 0.707035f
C6741 a_n2982_13878.n138 gnd 0.301852f
C6742 a_n2982_13878.n139 gnd 0.296371f
C6743 a_n2982_13878.t93 gnd 0.707035f
C6744 a_n2982_13878.n140 gnd 0.301852f
C6745 a_n2982_13878.n141 gnd 0.296371f
C6746 a_n2982_13878.t88 gnd 0.707035f
C6747 a_n2982_13878.n142 gnd 0.301852f
C6748 a_n2982_13878.n143 gnd 0.296371f
C6749 a_n2982_13878.n144 gnd 1.36231f
C6750 a_n2982_13878.t78 gnd 0.695384f
C6751 a_n2982_13878.n145 gnd 0.307896f
C6752 a_n2982_13878.t104 gnd 0.695384f
C6753 a_n2982_13878.n146 gnd 0.305597f
C6754 a_n2982_13878.n147 gnd 0.305735f
C6755 a_n2982_13878.t100 gnd 0.695384f
C6756 a_n2982_13878.n148 gnd 0.301852f
C6757 a_n2982_13878.t73 gnd 0.695384f
C6758 a_n2982_13878.n149 gnd 0.302112f
C6759 a_n2982_13878.n150 gnd 0.307896f
C6760 a_n2982_13878.t75 gnd 0.70657f
C6761 a_n2982_13878.t52 gnd 0.695384f
C6762 a_n2982_13878.n151 gnd 0.307896f
C6763 a_n2982_13878.t24 gnd 0.695384f
C6764 a_n2982_13878.n152 gnd 0.305597f
C6765 a_n2982_13878.n153 gnd 0.305735f
C6766 a_n2982_13878.t20 gnd 0.695384f
C6767 a_n2982_13878.n154 gnd 0.301852f
C6768 a_n2982_13878.t58 gnd 0.695384f
C6769 a_n2982_13878.n155 gnd 0.302112f
C6770 a_n2982_13878.n156 gnd 0.307896f
C6771 a_n2982_13878.t46 gnd 0.70657f
C6772 a_n2982_13878.n157 gnd 1.34634f
C6773 a_n2982_13878.t47 gnd 1.39701f
C6774 a_n2982_13878.t37 gnd 0.149496f
C6775 a_n2982_13878.t65 gnd 0.149496f
C6776 a_n2982_13878.n158 gnd 1.05305f
C6777 a_n2982_13878.t49 gnd 0.149496f
C6778 a_n2982_13878.t59 gnd 0.149496f
C6779 a_n2982_13878.n159 gnd 1.05305f
C6780 a_n2982_13878.n160 gnd 1.05305f
C6781 a_n2982_13878.t21 gnd 0.149496f
.ends

