* NGSPICE file created from opamp48.ext - technology: sky130A

.subckt opamp48 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 CSoutput.t169 a_n6308_8799.t36 vdd.t227 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X1 gnd.t413 commonsourceibias.t28 commonsourceibias.t29 gnd.t316 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n6308_8799.t21 plus.t5 a_n3827_n3924.t51 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X3 a_n1808_13878.t19 a_n2408_n452.t21 a_n2408_n452.t22 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t78 vdd.t76 vdd.t77 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X5 a_n1808_13878.t7 a_n2408_n452.t48 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 gnd.t146 gnd.t144 gnd.t145 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X7 gnd.t412 commonsourceibias.t80 CSoutput.t56 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t411 commonsourceibias.t81 CSoutput.t191 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 CSoutput.t64 commonsourceibias.t82 gnd.t410 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 CSoutput.t168 a_n6308_8799.t37 vdd.t222 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 commonsourceibias.t27 commonsourceibias.t26 gnd.t409 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 gnd.t408 commonsourceibias.t83 CSoutput.t62 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t143 gnd.t141 minus.t4 gnd.t142 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X14 gnd.t407 commonsourceibias.t36 commonsourceibias.t37 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 a_n3827_n3924.t55 diffpairibias.t20 gnd.t205 gnd.t204 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X16 CSoutput.t82 commonsourceibias.t84 gnd.t406 gnd.t354 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 CSoutput.t167 a_n6308_8799.t38 vdd.t226 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 a_n3827_n3924.t50 plus.t6 a_n6308_8799.t24 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X19 gnd.t405 commonsourceibias.t34 commonsourceibias.t35 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 a_n3827_n3924.t10 minus.t5 a_n2408_n452.t10 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X21 a_n1986_8322.t19 a_n2408_n452.t49 a_n6308_8799.t4 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X22 commonsourceibias.t33 commonsourceibias.t32 gnd.t404 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 gnd.t403 commonsourceibias.t85 CSoutput.t11 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 a_n2408_n452.t12 minus.t6 a_n3827_n3924.t13 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X25 gnd.t140 gnd.t138 gnd.t139 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X26 CSoutput.t67 commonsourceibias.t86 gnd.t402 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 vdd.t221 a_n6308_8799.t39 CSoutput.t166 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 gnd.t137 gnd.t134 gnd.t136 gnd.t135 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X29 CSoutput.t3 commonsourceibias.t87 gnd.t401 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 a_n2408_n452.t7 minus.t7 a_n3827_n3924.t7 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X31 CSoutput.t165 a_n6308_8799.t40 vdd.t220 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 vdd.t225 a_n6308_8799.t41 CSoutput.t164 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 commonsourceibias.t31 commonsourceibias.t30 gnd.t400 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 a_n6308_8799.t27 a_n2408_n452.t50 a_n1986_8322.t18 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X35 CSoutput.t163 a_n6308_8799.t42 vdd.t224 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X36 gnd.t399 commonsourceibias.t88 CSoutput.t96 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 gnd.t133 gnd.t131 gnd.t132 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X38 CSoutput.t44 commonsourceibias.t89 gnd.t398 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X39 vdd.t75 vdd.t73 vdd.t74 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X40 a_n3827_n3924.t2 minus.t8 a_n2408_n452.t2 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X41 CSoutput.t182 commonsourceibias.t90 gnd.t397 gnd.t354 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 gnd.t396 commonsourceibias.t18 commonsourceibias.t19 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X43 outputibias.t7 outputibias.t6 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X44 gnd.t395 commonsourceibias.t16 commonsourceibias.t17 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X45 CSoutput.t190 commonsourceibias.t91 gnd.t386 gnd.t318 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 CSoutput.t162 a_n6308_8799.t43 vdd.t223 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 vdd.t72 vdd.t70 vdd.t71 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X48 CSoutput.t161 a_n6308_8799.t44 vdd.t219 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 a_n3827_n3924.t11 diffpairibias.t21 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X50 commonsourceibias.t15 commonsourceibias.t14 gnd.t394 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t187 commonsourceibias.t92 gnd.t393 gnd.t318 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t160 a_n6308_8799.t45 vdd.t218 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 a_n3827_n3924.t49 plus.t7 a_n6308_8799.t16 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X54 gnd.t392 commonsourceibias.t12 commonsourceibias.t13 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X55 CSoutput.t177 commonsourceibias.t93 gnd.t391 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X56 a_n1808_13878.t18 a_n2408_n452.t31 a_n2408_n452.t32 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X57 vdd.t217 a_n6308_8799.t46 CSoutput.t159 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 a_n6308_8799.t31 plus.t8 a_n3827_n3924.t48 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X59 CSoutput.t158 a_n6308_8799.t47 vdd.t216 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X60 a_n2408_n452.t30 a_n2408_n452.t29 a_n1808_13878.t17 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X61 a_n6308_8799.t11 plus.t9 a_n3827_n3924.t47 gnd.t153 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X62 vdd.t69 vdd.t67 vdd.t68 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X63 CSoutput.t30 commonsourceibias.t94 gnd.t390 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X64 vdd.t123 CSoutput.t192 output.t19 gnd.t197 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X65 gnd.t389 commonsourceibias.t95 CSoutput.t73 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X66 diffpairibias.t19 diffpairibias.t18 gnd.t179 gnd.t178 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X67 CSoutput.t94 commonsourceibias.t96 gnd.t385 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 a_n3827_n3924.t46 plus.t10 a_n6308_8799.t20 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X69 a_n2408_n452.t11 minus.t9 a_n3827_n3924.t12 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X70 CSoutput.t91 commonsourceibias.t97 gnd.t388 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X71 CSoutput.t95 commonsourceibias.t98 gnd.t387 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 commonsourceibias.t39 commonsourceibias.t38 gnd.t384 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 gnd.t130 gnd.t128 plus.t4 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X74 gnd.t127 gnd.t125 gnd.t126 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X75 CSoutput.t7 commonsourceibias.t99 gnd.t383 gnd.t354 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 vdd.t215 a_n6308_8799.t48 CSoutput.t157 vdd.t214 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 vdd.t213 a_n6308_8799.t49 CSoutput.t156 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 diffpairibias.t17 diffpairibias.t16 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 CSoutput.t155 a_n6308_8799.t50 vdd.t212 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X80 gnd.t124 gnd.t122 gnd.t123 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X81 CSoutput.t85 commonsourceibias.t100 gnd.t382 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X82 vdd.t211 a_n6308_8799.t51 CSoutput.t154 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 CSoutput.t31 commonsourceibias.t101 gnd.t381 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 CSoutput.t153 a_n6308_8799.t52 vdd.t204 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 gnd.t121 gnd.t119 gnd.t120 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X86 CSoutput.t152 a_n6308_8799.t53 vdd.t210 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 CSoutput.t151 a_n6308_8799.t54 vdd.t209 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X88 vdd.t208 a_n6308_8799.t55 CSoutput.t150 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 gnd.t380 commonsourceibias.t102 CSoutput.t53 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 gnd.t118 gnd.t116 gnd.t117 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X91 gnd.t115 gnd.t113 plus.t3 gnd.t114 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X92 CSoutput.t37 commonsourceibias.t103 gnd.t379 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 gnd.t378 commonsourceibias.t104 CSoutput.t46 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X94 a_n3827_n3924.t45 plus.t11 a_n6308_8799.t15 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X95 gnd.t112 gnd.t110 gnd.t111 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X96 output.t3 outputibias.t8 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X97 a_n3827_n3924.t54 diffpairibias.t22 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X98 CSoutput.t183 commonsourceibias.t105 gnd.t377 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 a_n2408_n452.t42 a_n2408_n452.t41 a_n1808_13878.t16 vdd.t81 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 vdd.t207 a_n6308_8799.t56 CSoutput.t149 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 vdd.t206 a_n6308_8799.t57 CSoutput.t148 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n6308_8799.t28 a_n2408_n452.t51 a_n1986_8322.t17 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X103 a_n2408_n452.t26 a_n2408_n452.t25 a_n1808_13878.t15 vdd.t97 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X104 gnd.t376 commonsourceibias.t106 CSoutput.t75 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X105 vdd.t89 CSoutput.t193 output.t18 gnd.t196 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X106 vdd.t205 a_n6308_8799.t58 CSoutput.t147 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 commonsourceibias.t41 commonsourceibias.t40 gnd.t375 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t374 commonsourceibias.t107 CSoutput.t22 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 gnd.t109 gnd.t106 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X110 CSoutput.t43 commonsourceibias.t108 gnd.t373 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X111 vdd.t203 a_n6308_8799.t59 CSoutput.t146 vdd.t155 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X112 CSoutput.t194 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X113 gnd.t372 commonsourceibias.t46 commonsourceibias.t47 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 CSoutput.t145 a_n6308_8799.t60 vdd.t202 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 CSoutput.t58 commonsourceibias.t109 gnd.t371 gnd.t318 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X116 diffpairibias.t15 diffpairibias.t14 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X117 a_n2408_n452.t45 minus.t10 a_n3827_n3924.t26 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X118 vdd.t66 vdd.t64 vdd.t65 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X119 vdd.t201 a_n6308_8799.t61 CSoutput.t144 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 vdd.t63 vdd.t60 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 gnd.t370 commonsourceibias.t110 CSoutput.t40 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 a_n3827_n3924.t25 minus.t11 a_n2408_n452.t44 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X123 vdd.t59 vdd.t57 vdd.t58 vdd.t8 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X124 vdd.t56 vdd.t54 vdd.t55 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X125 vdd.t120 a_n2408_n452.t52 a_n1986_8322.t7 vdd.t119 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 gnd.t369 commonsourceibias.t44 commonsourceibias.t45 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 CSoutput.t26 commonsourceibias.t111 gnd.t368 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 CSoutput.t14 commonsourceibias.t112 gnd.t367 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X129 a_n1986_8322.t6 a_n2408_n452.t53 vdd.t122 vdd.t121 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 a_n3827_n3924.t23 diffpairibias.t23 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X131 CSoutput.t143 a_n6308_8799.t62 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X132 gnd.t366 commonsourceibias.t113 CSoutput.t29 gnd.t316 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 vdd.t198 a_n6308_8799.t63 CSoutput.t142 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 a_n3827_n3924.t4 minus.t12 a_n2408_n452.t4 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X135 a_n3827_n3924.t8 minus.t13 a_n2408_n452.t8 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X136 commonsourceibias.t43 commonsourceibias.t42 gnd.t365 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X137 vdd.t104 a_n2408_n452.t54 a_n1808_13878.t6 vdd.t103 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X138 gnd.t364 commonsourceibias.t114 CSoutput.t23 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X139 commonsourceibias.t79 commonsourceibias.t78 gnd.t363 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 a_n2408_n452.t3 minus.t14 a_n3827_n3924.t3 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X141 a_n3827_n3924.t44 plus.t12 a_n6308_8799.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X142 a_n3827_n3924.t43 plus.t13 a_n6308_8799.t32 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X143 vdd.t53 vdd.t50 vdd.t52 vdd.t51 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 gnd.t362 commonsourceibias.t76 commonsourceibias.t77 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X145 output.t17 CSoutput.t195 vdd.t90 gnd.t195 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X146 CSoutput.t60 commonsourceibias.t115 gnd.t361 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 gnd.t360 commonsourceibias.t116 CSoutput.t172 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X148 a_n2408_n452.t43 minus.t15 a_n3827_n3924.t24 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X149 vdd.t49 vdd.t46 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X150 vdd.t196 a_n6308_8799.t64 CSoutput.t141 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 gnd.t105 gnd.t103 plus.t2 gnd.t104 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X152 CSoutput.t49 commonsourceibias.t117 gnd.t359 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n6308_8799.t26 plus.t14 a_n3827_n3924.t42 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X154 a_n6308_8799.t19 plus.t15 a_n3827_n3924.t41 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X155 commonsourceibias.t75 commonsourceibias.t74 gnd.t358 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X156 vdd.t45 vdd.t42 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X157 a_n1986_8322.t5 a_n2408_n452.t55 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X158 a_n6308_8799.t22 a_n2408_n452.t56 a_n1986_8322.t16 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X159 gnd.t357 commonsourceibias.t118 CSoutput.t83 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X160 diffpairibias.t13 diffpairibias.t12 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X161 CSoutput.t196 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X162 a_n2408_n452.t1 minus.t16 a_n3827_n3924.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X163 a_n2408_n452.t40 a_n2408_n452.t39 a_n1808_13878.t14 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X164 vdd.t194 a_n6308_8799.t65 CSoutput.t140 vdd.t155 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X165 a_n6308_8799.t23 a_n2408_n452.t57 a_n1986_8322.t15 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X166 CSoutput.t139 a_n6308_8799.t66 vdd.t193 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 gnd.t356 commonsourceibias.t72 commonsourceibias.t73 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 a_n1808_13878.t13 a_n2408_n452.t37 a_n2408_n452.t38 vdd.t113 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X169 commonsourceibias.t71 commonsourceibias.t70 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 a_n3827_n3924.t27 minus.t17 a_n2408_n452.t46 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X171 gnd.t353 commonsourceibias.t119 CSoutput.t65 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 gnd.t102 gnd.t100 gnd.t101 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X173 output.t16 CSoutput.t197 vdd.t91 gnd.t194 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X174 gnd.t352 commonsourceibias.t120 CSoutput.t78 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 gnd.t99 gnd.t96 gnd.t98 gnd.t97 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X176 vdd.t86 a_n2408_n452.t58 a_n1986_8322.t4 vdd.t85 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X177 output.t2 outputibias.t9 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X178 gnd.t95 gnd.t93 gnd.t94 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X179 output.t15 CSoutput.t198 vdd.t92 gnd.t193 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X180 minus.t3 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X181 CSoutput.t138 a_n6308_8799.t67 vdd.t192 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X182 vdd.t93 CSoutput.t199 output.t14 gnd.t192 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X183 vdd.t191 a_n6308_8799.t68 CSoutput.t137 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X184 CSoutput.t54 commonsourceibias.t121 gnd.t351 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 gnd.t350 commonsourceibias.t122 CSoutput.t174 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 commonsourceibias.t49 commonsourceibias.t48 gnd.t349 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 gnd.t348 commonsourceibias.t123 CSoutput.t45 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 a_n3827_n3924.t40 plus.t16 a_n6308_8799.t10 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X189 gnd.t347 commonsourceibias.t124 CSoutput.t93 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X190 a_n3827_n3924.t52 diffpairibias.t24 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X191 a_n3827_n3924.t17 diffpairibias.t25 gnd.t148 gnd.t147 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X192 vdd.t190 a_n6308_8799.t69 CSoutput.t136 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X193 a_n6308_8799.t9 plus.t17 a_n3827_n3924.t39 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X194 CSoutput.t200 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X195 CSoutput.t135 a_n6308_8799.t70 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X196 CSoutput.t134 a_n6308_8799.t71 vdd.t187 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t201 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X198 CSoutput.t79 commonsourceibias.t125 gnd.t346 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 output.t13 CSoutput.t202 vdd.t0 gnd.t191 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X200 gnd.t89 gnd.t87 gnd.t88 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X201 gnd.t345 commonsourceibias.t126 CSoutput.t17 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 diffpairibias.t11 diffpairibias.t10 gnd.t166 gnd.t165 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X203 gnd.t86 gnd.t84 gnd.t85 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X204 a_n1808_13878.t5 a_n2408_n452.t59 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X205 vdd.t41 vdd.t39 vdd.t40 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X206 vdd.t95 a_n2408_n452.t60 a_n1808_13878.t4 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X207 gnd.t344 commonsourceibias.t127 CSoutput.t72 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 gnd.t343 commonsourceibias.t128 CSoutput.t48 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 CSoutput.t10 commonsourceibias.t129 gnd.t342 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X210 output.t12 CSoutput.t203 vdd.t1 gnd.t190 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X211 outputibias.t5 outputibias.t4 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X212 plus.t1 gnd.t81 gnd.t83 gnd.t82 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X213 diffpairibias.t9 diffpairibias.t8 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X214 gnd.t231 commonsourceibias.t130 CSoutput.t61 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 a_n3827_n3924.t56 minus.t18 a_n2408_n452.t47 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X216 CSoutput.t133 a_n6308_8799.t72 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 gnd.t341 commonsourceibias.t131 CSoutput.t66 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 vdd.t186 a_n6308_8799.t73 CSoutput.t132 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X219 commonsourceibias.t11 commonsourceibias.t10 gnd.t340 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 a_n2408_n452.t18 minus.t19 a_n3827_n3924.t21 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X221 a_n1986_8322.t14 a_n2408_n452.t61 a_n6308_8799.t6 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X222 diffpairibias.t7 diffpairibias.t6 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X223 a_n2408_n452.t17 minus.t20 a_n3827_n3924.t20 gnd.t153 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X224 CSoutput.t131 a_n6308_8799.t74 vdd.t185 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 a_n2408_n452.t14 minus.t21 a_n3827_n3924.t16 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X226 vdd.t184 a_n6308_8799.t75 CSoutput.t130 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 vdd.t229 a_n2408_n452.t62 a_n1986_8322.t3 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X228 vdd.t180 a_n6308_8799.t76 CSoutput.t129 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 a_n3827_n3924.t6 minus.t22 a_n2408_n452.t6 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X230 CSoutput.t89 commonsourceibias.t132 gnd.t339 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X231 a_n6308_8799.t33 plus.t18 a_n3827_n3924.t38 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X232 gnd.t80 gnd.t78 gnd.t79 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X233 commonsourceibias.t9 commonsourceibias.t8 gnd.t338 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X234 commonsourceibias.t7 commonsourceibias.t6 gnd.t337 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 a_n3827_n3924.t5 minus.t23 a_n2408_n452.t5 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X236 gnd.t77 gnd.t74 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X237 gnd.t73 gnd.t70 gnd.t72 gnd.t71 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X238 a_n1808_13878.t3 a_n2408_n452.t63 vdd.t231 vdd.t230 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X239 vdd.t2 CSoutput.t204 output.t11 gnd.t189 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X240 CSoutput.t5 commonsourceibias.t133 gnd.t336 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 vdd.t179 a_n6308_8799.t77 CSoutput.t128 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 vdd.t38 vdd.t36 vdd.t37 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X243 gnd.t328 commonsourceibias.t134 CSoutput.t4 gnd.t316 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 CSoutput.t127 a_n6308_8799.t78 vdd.t178 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 CSoutput.t126 a_n6308_8799.t79 vdd.t177 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 gnd.t335 commonsourceibias.t50 commonsourceibias.t51 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X247 gnd.t69 gnd.t67 minus.t2 gnd.t68 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X248 gnd.t334 commonsourceibias.t135 CSoutput.t175 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t51 commonsourceibias.t136 gnd.t333 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 gnd.t66 gnd.t63 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X251 CSoutput.t16 commonsourceibias.t137 gnd.t332 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 gnd.t331 commonsourceibias.t138 CSoutput.t8 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 CSoutput.t80 commonsourceibias.t139 gnd.t330 gnd.t329 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t62 gnd.t60 gnd.t61 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X255 vdd.t35 vdd.t33 vdd.t34 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X256 a_n3827_n3924.t14 diffpairibias.t26 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X257 gnd.t327 commonsourceibias.t140 CSoutput.t19 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X258 a_n1986_8322.t13 a_n2408_n452.t64 a_n6308_8799.t12 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X259 commonsourceibias.t55 commonsourceibias.t54 gnd.t326 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 vdd.t126 CSoutput.t205 output.t10 gnd.t188 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X261 vdd.t102 a_n2408_n452.t65 a_n1986_8322.t2 vdd.t101 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X262 CSoutput.t125 a_n6308_8799.t80 vdd.t176 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 vdd.t174 a_n6308_8799.t81 CSoutput.t124 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X264 CSoutput.t21 commonsourceibias.t141 gnd.t325 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 CSoutput.t123 a_n6308_8799.t82 vdd.t173 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X266 gnd.t324 commonsourceibias.t142 CSoutput.t74 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 vdd.t172 a_n6308_8799.t83 CSoutput.t122 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 vdd.t171 a_n6308_8799.t84 CSoutput.t121 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 a_n6308_8799.t2 plus.t19 a_n3827_n3924.t37 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X270 CSoutput.t92 commonsourceibias.t143 gnd.t323 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 outputibias.t3 outputibias.t2 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X272 gnd.t322 commonsourceibias.t144 CSoutput.t38 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X273 gnd.t321 commonsourceibias.t145 CSoutput.t50 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X274 CSoutput.t170 commonsourceibias.t146 gnd.t320 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 gnd.t59 gnd.t56 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X276 commonsourceibias.t53 commonsourceibias.t52 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X277 vdd.t32 vdd.t29 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X278 a_n3827_n3924.t36 plus.t20 a_n6308_8799.t25 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X279 a_n1808_13878.t12 a_n2408_n452.t35 a_n2408_n452.t36 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X280 CSoutput.t32 commonsourceibias.t147 gnd.t297 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n1986_8322.t12 a_n2408_n452.t66 a_n6308_8799.t5 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 output.t1 outputibias.t10 gnd.t174 gnd.t173 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X283 diffpairibias.t5 diffpairibias.t4 gnd.t415 gnd.t414 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X284 gnd.t317 commonsourceibias.t148 CSoutput.t179 gnd.t316 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 CSoutput.t188 commonsourceibias.t149 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X286 gnd.t313 commonsourceibias.t58 commonsourceibias.t59 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 gnd.t55 gnd.t52 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X288 outputibias.t1 outputibias.t0 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X289 commonsourceibias.t57 commonsourceibias.t56 gnd.t312 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 CSoutput.t120 a_n6308_8799.t85 vdd.t170 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 gnd.t311 commonsourceibias.t150 CSoutput.t81 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 a_n3827_n3924.t22 diffpairibias.t27 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X293 vdd.t143 a_n6308_8799.t86 CSoutput.t119 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X294 gnd.t310 commonsourceibias.t151 CSoutput.t9 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 gnd.t309 commonsourceibias.t152 CSoutput.t34 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 gnd.t307 commonsourceibias.t153 CSoutput.t57 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X297 CSoutput.t206 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X298 vdd.t28 vdd.t26 vdd.t27 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X299 vdd.t168 a_n6308_8799.t87 CSoutput.t118 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 a_n1986_8322.t1 a_n2408_n452.t67 vdd.t84 vdd.t83 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X301 gnd.t306 commonsourceibias.t154 CSoutput.t39 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 CSoutput.t181 commonsourceibias.t155 gnd.t305 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 CSoutput.t117 a_n6308_8799.t88 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 output.t9 CSoutput.t207 vdd.t127 gnd.t187 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X305 gnd.t304 commonsourceibias.t62 commonsourceibias.t63 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 commonsourceibias.t61 commonsourceibias.t60 gnd.t303 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 vdd.t108 a_n2408_n452.t68 a_n1808_13878.t2 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X308 plus.t0 gnd.t49 gnd.t51 gnd.t50 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X309 gnd.t302 commonsourceibias.t156 CSoutput.t86 gnd.t301 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 CSoutput.t84 commonsourceibias.t157 gnd.t300 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 CSoutput.t116 a_n6308_8799.t89 vdd.t166 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X312 CSoutput.t59 commonsourceibias.t158 gnd.t299 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 gnd.t296 commonsourceibias.t159 CSoutput.t71 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 commonsourceibias.t23 commonsourceibias.t22 gnd.t295 gnd.t294 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 gnd.t293 commonsourceibias.t160 CSoutput.t0 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X316 a_n3827_n3924.t35 plus.t21 a_n6308_8799.t18 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.7
X317 vdd.t165 a_n6308_8799.t90 CSoutput.t115 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 vdd.t145 a_n6308_8799.t91 CSoutput.t114 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 vdd.t25 vdd.t22 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X320 gnd.t292 commonsourceibias.t20 commonsourceibias.t21 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 a_n3827_n3924.t0 minus.t24 a_n2408_n452.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X322 a_n1986_8322.t11 a_n2408_n452.t69 a_n6308_8799.t13 vdd.t109 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X323 vdd.t21 vdd.t19 vdd.t20 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X324 CSoutput.t113 a_n6308_8799.t92 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 a_n6308_8799.t14 a_n2408_n452.t70 a_n1986_8322.t10 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X326 output.t0 outputibias.t11 gnd.t213 gnd.t212 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X327 gnd.t291 commonsourceibias.t161 CSoutput.t63 gnd.t290 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X328 a_n6308_8799.t1 plus.t22 a_n3827_n3924.t34 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X329 vdd.t162 a_n6308_8799.t93 CSoutput.t112 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 a_n1808_13878.t1 a_n2408_n452.t71 vdd.t112 vdd.t111 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X331 CSoutput.t6 commonsourceibias.t162 gnd.t289 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 CSoutput.t12 commonsourceibias.t163 gnd.t288 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 gnd.t287 commonsourceibias.t164 CSoutput.t18 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 CSoutput.t42 commonsourceibias.t165 gnd.t286 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 a_n2408_n452.t16 minus.t25 a_n3827_n3924.t19 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X336 vdd.t128 CSoutput.t208 output.t8 gnd.t186 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X337 gnd.t284 commonsourceibias.t64 commonsourceibias.t65 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 CSoutput.t87 commonsourceibias.t166 gnd.t283 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X339 CSoutput.t2 commonsourceibias.t167 gnd.t282 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 CSoutput.t25 commonsourceibias.t168 gnd.t281 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 gnd.t280 commonsourceibias.t169 CSoutput.t35 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X342 a_n6308_8799.t35 plus.t23 a_n3827_n3924.t33 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X343 gnd.t48 gnd.t45 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.7
X344 CSoutput.t97 commonsourceibias.t170 gnd.t279 gnd.t278 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 gnd.t44 gnd.t42 minus.t1 gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X346 a_n3827_n3924.t9 minus.t26 a_n2408_n452.t9 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X347 CSoutput.t47 commonsourceibias.t171 gnd.t277 gnd.t276 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 CSoutput.t36 commonsourceibias.t172 gnd.t275 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 gnd.t274 commonsourceibias.t173 CSoutput.t184 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X350 CSoutput.t111 a_n6308_8799.t94 vdd.t160 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 a_n1808_13878.t11 a_n2408_n452.t23 a_n2408_n452.t24 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X352 output.t7 CSoutput.t209 vdd.t129 gnd.t185 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X353 a_n3827_n3924.t32 plus.t24 a_n6308_8799.t3 gnd.t12 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X354 gnd.t273 commonsourceibias.t4 commonsourceibias.t5 gnd.t272 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 CSoutput.t210 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X356 gnd.t271 commonsourceibias.t2 commonsourceibias.t3 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 gnd.t269 commonsourceibias.t0 commonsourceibias.t1 gnd.t268 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 CSoutput.t110 a_n6308_8799.t95 vdd.t159 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X359 a_n3827_n3924.t53 diffpairibias.t28 gnd.t201 gnd.t200 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X360 vdd.t158 a_n6308_8799.t96 CSoutput.t109 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X361 CSoutput.t15 commonsourceibias.t174 gnd.t267 gnd.t266 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 gnd.t265 commonsourceibias.t175 CSoutput.t90 gnd.t230 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 a_n2408_n452.t34 a_n2408_n452.t33 a_n1808_13878.t10 vdd.t109 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X364 a_n6308_8799.t29 a_n2408_n452.t72 a_n1986_8322.t9 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X365 CSoutput.t28 commonsourceibias.t176 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 a_n6308_8799.t34 plus.t25 a_n3827_n3924.t31 gnd.t177 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X367 vdd.t157 a_n6308_8799.t97 CSoutput.t108 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd.t41 gnd.t38 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X369 gnd.t262 commonsourceibias.t177 CSoutput.t55 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X370 gnd.t261 commonsourceibias.t178 CSoutput.t13 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 gnd.t259 commonsourceibias.t179 CSoutput.t180 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 diffpairibias.t3 diffpairibias.t2 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X373 gnd.t257 commonsourceibias.t180 CSoutput.t173 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X374 vdd.t156 a_n6308_8799.t98 CSoutput.t107 vdd.t155 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X375 vdd.t18 vdd.t15 vdd.t17 vdd.t16 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X376 CSoutput.t88 commonsourceibias.t181 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 CSoutput.t106 a_n6308_8799.t99 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X378 output.t6 CSoutput.t211 vdd.t130 gnd.t184 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X379 vdd.t131 CSoutput.t212 output.t5 gnd.t183 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X380 a_n3827_n3924.t30 plus.t26 a_n6308_8799.t17 gnd.t170 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X381 gnd.t254 commonsourceibias.t182 CSoutput.t176 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 gnd.t252 commonsourceibias.t183 CSoutput.t171 gnd.t251 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X383 gnd.t37 gnd.t34 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X384 gnd.t33 gnd.t30 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X385 diffpairibias.t1 diffpairibias.t0 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X386 CSoutput.t52 commonsourceibias.t184 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X387 CSoutput.t20 commonsourceibias.t185 gnd.t248 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X388 gnd.t246 commonsourceibias.t24 commonsourceibias.t25 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X389 a_n3827_n3924.t29 plus.t27 a_n6308_8799.t30 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X390 gnd.t244 commonsourceibias.t186 CSoutput.t33 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X391 vdd.t125 a_n2408_n452.t73 a_n1808_13878.t0 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X392 a_n6308_8799.t7 plus.t28 a_n3827_n3924.t28 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X393 a_n3827_n3924.t15 minus.t27 a_n2408_n452.t13 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.7
X394 CSoutput.t105 a_n6308_8799.t100 vdd.t151 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 vdd.t152 a_n6308_8799.t101 CSoutput.t104 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 gnd.t243 commonsourceibias.t187 CSoutput.t27 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 CSoutput.t103 a_n6308_8799.t102 vdd.t149 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X398 gnd.t241 commonsourceibias.t66 commonsourceibias.t67 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 gnd.t239 commonsourceibias.t188 CSoutput.t77 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X400 CSoutput.t178 commonsourceibias.t189 gnd.t238 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X401 gnd.t237 commonsourceibias.t190 CSoutput.t189 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 a_n2408_n452.t15 minus.t28 a_n3827_n3924.t18 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.7
X403 CSoutput.t102 a_n6308_8799.t103 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X404 a_n1986_8322.t8 a_n2408_n452.t74 a_n6308_8799.t8 vdd.t97 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X405 CSoutput.t68 commonsourceibias.t191 gnd.t235 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X406 CSoutput.t70 commonsourceibias.t192 gnd.t233 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X407 vdd.t139 a_n6308_8799.t104 CSoutput.t101 vdd.t138 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X408 CSoutput.t100 a_n6308_8799.t105 vdd.t137 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X409 vdd.t135 a_n6308_8799.t106 CSoutput.t99 vdd.t134 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X410 gnd.t229 commonsourceibias.t193 CSoutput.t41 gnd.t228 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 commonsourceibias.t69 commonsourceibias.t68 gnd.t227 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X412 gnd.t225 commonsourceibias.t194 CSoutput.t76 gnd.t224 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 CSoutput.t24 commonsourceibias.t195 gnd.t223 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X414 a_n1986_8322.t0 a_n2408_n452.t75 vdd.t99 vdd.t98 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X415 vdd.t14 vdd.t11 vdd.t13 vdd.t12 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X416 gnd.t221 commonsourceibias.t196 CSoutput.t185 gnd.t220 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X417 a_n1808_13878.t9 a_n2408_n452.t27 a_n2408_n452.t28 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X418 vdd.t116 CSoutput.t213 output.t4 gnd.t182 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X419 vdd.t133 a_n6308_8799.t107 CSoutput.t98 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X420 minus.t0 gnd.t27 gnd.t29 gnd.t28 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X421 a_n3827_n3924.t57 diffpairibias.t29 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X422 CSoutput.t186 commonsourceibias.t197 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X423 CSoutput.t69 commonsourceibias.t198 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 a_n2408_n452.t20 a_n2408_n452.t19 a_n1808_13878.t8 vdd.t96 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X425 gnd.t215 commonsourceibias.t199 CSoutput.t1 gnd.t214 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X426 vdd.t10 vdd.t7 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X427 vdd.t6 vdd.t3 vdd.t5 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
R0 a_n6308_8799.n138 a_n6308_8799.t82 490.524
R1 a_n6308_8799.n149 a_n6308_8799.t89 490.524
R2 a_n6308_8799.n161 a_n6308_8799.t99 490.524
R3 a_n6308_8799.n104 a_n6308_8799.t59 490.524
R4 a_n6308_8799.n115 a_n6308_8799.t65 490.524
R5 a_n6308_8799.n127 a_n6308_8799.t98 490.524
R6 a_n6308_8799.n30 a_n6308_8799.t68 484.3
R7 a_n6308_8799.n144 a_n6308_8799.t67 464.166
R8 a_n6308_8799.n143 a_n6308_8799.t49 464.166
R9 a_n6308_8799.n134 a_n6308_8799.t95 464.166
R10 a_n6308_8799.n142 a_n6308_8799.t69 464.166
R11 a_n6308_8799.n141 a_n6308_8799.t54 464.166
R12 a_n6308_8799.n135 a_n6308_8799.t97 464.166
R13 a_n6308_8799.n140 a_n6308_8799.t79 464.166
R14 a_n6308_8799.n139 a_n6308_8799.t77 464.166
R15 a_n6308_8799.n136 a_n6308_8799.t38 464.166
R16 a_n6308_8799.n137 a_n6308_8799.t83 464.166
R17 a_n6308_8799.n39 a_n6308_8799.t73 484.3
R18 a_n6308_8799.n155 a_n6308_8799.t72 464.166
R19 a_n6308_8799.n154 a_n6308_8799.t61 464.166
R20 a_n6308_8799.n145 a_n6308_8799.t103 464.166
R21 a_n6308_8799.n153 a_n6308_8799.t76 464.166
R22 a_n6308_8799.n152 a_n6308_8799.t62 464.166
R23 a_n6308_8799.n146 a_n6308_8799.t107 464.166
R24 a_n6308_8799.n151 a_n6308_8799.t88 464.166
R25 a_n6308_8799.n150 a_n6308_8799.t87 464.166
R26 a_n6308_8799.n147 a_n6308_8799.t45 464.166
R27 a_n6308_8799.n148 a_n6308_8799.t90 464.166
R28 a_n6308_8799.n48 a_n6308_8799.t106 484.3
R29 a_n6308_8799.n167 a_n6308_8799.t47 464.166
R30 a_n6308_8799.n166 a_n6308_8799.t75 464.166
R31 a_n6308_8799.n157 a_n6308_8799.t37 464.166
R32 a_n6308_8799.n165 a_n6308_8799.t93 464.166
R33 a_n6308_8799.n164 a_n6308_8799.t52 464.166
R34 a_n6308_8799.n158 a_n6308_8799.t81 464.166
R35 a_n6308_8799.n163 a_n6308_8799.t40 464.166
R36 a_n6308_8799.n162 a_n6308_8799.t56 464.166
R37 a_n6308_8799.n159 a_n6308_8799.t102 464.166
R38 a_n6308_8799.n160 a_n6308_8799.t86 464.166
R39 a_n6308_8799.n103 a_n6308_8799.t60 464.166
R40 a_n6308_8799.n102 a_n6308_8799.t84 464.166
R41 a_n6308_8799.n105 a_n6308_8799.t36 464.166
R42 a_n6308_8799.n101 a_n6308_8799.t57 464.166
R43 a_n6308_8799.n106 a_n6308_8799.t71 464.166
R44 a_n6308_8799.n107 a_n6308_8799.t96 464.166
R45 a_n6308_8799.n100 a_n6308_8799.t44 464.166
R46 a_n6308_8799.n108 a_n6308_8799.t55 464.166
R47 a_n6308_8799.n99 a_n6308_8799.t94 464.166
R48 a_n6308_8799.n109 a_n6308_8799.t41 464.166
R49 a_n6308_8799.n114 a_n6308_8799.t66 464.166
R50 a_n6308_8799.n113 a_n6308_8799.t91 464.166
R51 a_n6308_8799.n116 a_n6308_8799.t43 464.166
R52 a_n6308_8799.n112 a_n6308_8799.t64 464.166
R53 a_n6308_8799.n117 a_n6308_8799.t78 464.166
R54 a_n6308_8799.n118 a_n6308_8799.t104 464.166
R55 a_n6308_8799.n111 a_n6308_8799.t53 464.166
R56 a_n6308_8799.n119 a_n6308_8799.t63 464.166
R57 a_n6308_8799.n110 a_n6308_8799.t100 464.166
R58 a_n6308_8799.n120 a_n6308_8799.t48 464.166
R59 a_n6308_8799.n126 a_n6308_8799.t85 464.166
R60 a_n6308_8799.n125 a_n6308_8799.t101 464.166
R61 a_n6308_8799.n128 a_n6308_8799.t70 464.166
R62 a_n6308_8799.n124 a_n6308_8799.t39 464.166
R63 a_n6308_8799.n129 a_n6308_8799.t80 464.166
R64 a_n6308_8799.n130 a_n6308_8799.t51 464.166
R65 a_n6308_8799.n123 a_n6308_8799.t92 464.166
R66 a_n6308_8799.n131 a_n6308_8799.t58 464.166
R67 a_n6308_8799.n122 a_n6308_8799.t74 464.166
R68 a_n6308_8799.n132 a_n6308_8799.t46 464.166
R69 a_n6308_8799.n38 a_n6308_8799.n37 75.3623
R70 a_n6308_8799.n36 a_n6308_8799.n24 70.3058
R71 a_n6308_8799.n24 a_n6308_8799.n35 70.1674
R72 a_n6308_8799.n35 a_n6308_8799.n135 20.9683
R73 a_n6308_8799.n34 a_n6308_8799.n25 75.0448
R74 a_n6308_8799.n141 a_n6308_8799.n34 11.2134
R75 a_n6308_8799.n33 a_n6308_8799.n25 80.4688
R76 a_n6308_8799.n27 a_n6308_8799.n32 74.73
R77 a_n6308_8799.n31 a_n6308_8799.n27 70.1674
R78 a_n6308_8799.n144 a_n6308_8799.n31 20.9683
R79 a_n6308_8799.n26 a_n6308_8799.n30 70.5844
R80 a_n6308_8799.n47 a_n6308_8799.n46 75.3623
R81 a_n6308_8799.n45 a_n6308_8799.n20 70.3058
R82 a_n6308_8799.n20 a_n6308_8799.n44 70.1674
R83 a_n6308_8799.n44 a_n6308_8799.n146 20.9683
R84 a_n6308_8799.n43 a_n6308_8799.n21 75.0448
R85 a_n6308_8799.n152 a_n6308_8799.n43 11.2134
R86 a_n6308_8799.n42 a_n6308_8799.n21 80.4688
R87 a_n6308_8799.n23 a_n6308_8799.n41 74.73
R88 a_n6308_8799.n40 a_n6308_8799.n23 70.1674
R89 a_n6308_8799.n155 a_n6308_8799.n40 20.9683
R90 a_n6308_8799.n22 a_n6308_8799.n39 70.5844
R91 a_n6308_8799.n56 a_n6308_8799.n55 75.3623
R92 a_n6308_8799.n54 a_n6308_8799.n16 70.3058
R93 a_n6308_8799.n16 a_n6308_8799.n53 70.1674
R94 a_n6308_8799.n53 a_n6308_8799.n158 20.9683
R95 a_n6308_8799.n52 a_n6308_8799.n17 75.0448
R96 a_n6308_8799.n164 a_n6308_8799.n52 11.2134
R97 a_n6308_8799.n51 a_n6308_8799.n17 80.4688
R98 a_n6308_8799.n19 a_n6308_8799.n50 74.73
R99 a_n6308_8799.n49 a_n6308_8799.n19 70.1674
R100 a_n6308_8799.n167 a_n6308_8799.n49 20.9683
R101 a_n6308_8799.n18 a_n6308_8799.n48 70.5844
R102 a_n6308_8799.n12 a_n6308_8799.n65 70.5844
R103 a_n6308_8799.n64 a_n6308_8799.n13 70.1674
R104 a_n6308_8799.n64 a_n6308_8799.n99 20.9683
R105 a_n6308_8799.n13 a_n6308_8799.n63 74.73
R106 a_n6308_8799.n108 a_n6308_8799.n63 11.843
R107 a_n6308_8799.n62 a_n6308_8799.n14 80.4688
R108 a_n6308_8799.n62 a_n6308_8799.n100 0.365327
R109 a_n6308_8799.n14 a_n6308_8799.n61 75.0448
R110 a_n6308_8799.n60 a_n6308_8799.n15 70.1674
R111 a_n6308_8799.n60 a_n6308_8799.n101 20.9683
R112 a_n6308_8799.n15 a_n6308_8799.n59 70.3058
R113 a_n6308_8799.n105 a_n6308_8799.n59 20.6913
R114 a_n6308_8799.n58 a_n6308_8799.n57 75.3623
R115 a_n6308_8799.n8 a_n6308_8799.n74 70.5844
R116 a_n6308_8799.n73 a_n6308_8799.n9 70.1674
R117 a_n6308_8799.n73 a_n6308_8799.n110 20.9683
R118 a_n6308_8799.n9 a_n6308_8799.n72 74.73
R119 a_n6308_8799.n119 a_n6308_8799.n72 11.843
R120 a_n6308_8799.n71 a_n6308_8799.n10 80.4688
R121 a_n6308_8799.n71 a_n6308_8799.n111 0.365327
R122 a_n6308_8799.n10 a_n6308_8799.n70 75.0448
R123 a_n6308_8799.n69 a_n6308_8799.n11 70.1674
R124 a_n6308_8799.n69 a_n6308_8799.n112 20.9683
R125 a_n6308_8799.n11 a_n6308_8799.n68 70.3058
R126 a_n6308_8799.n116 a_n6308_8799.n68 20.6913
R127 a_n6308_8799.n67 a_n6308_8799.n66 75.3623
R128 a_n6308_8799.n4 a_n6308_8799.n83 70.5844
R129 a_n6308_8799.n82 a_n6308_8799.n5 70.1674
R130 a_n6308_8799.n82 a_n6308_8799.n122 20.9683
R131 a_n6308_8799.n5 a_n6308_8799.n81 74.73
R132 a_n6308_8799.n131 a_n6308_8799.n81 11.843
R133 a_n6308_8799.n80 a_n6308_8799.n6 80.4688
R134 a_n6308_8799.n80 a_n6308_8799.n123 0.365327
R135 a_n6308_8799.n6 a_n6308_8799.n79 75.0448
R136 a_n6308_8799.n78 a_n6308_8799.n7 70.1674
R137 a_n6308_8799.n78 a_n6308_8799.n124 20.9683
R138 a_n6308_8799.n7 a_n6308_8799.n77 70.3058
R139 a_n6308_8799.n128 a_n6308_8799.n77 20.6913
R140 a_n6308_8799.n76 a_n6308_8799.n75 75.3623
R141 a_n6308_8799.n28 a_n6308_8799.n84 98.9633
R142 a_n6308_8799.n29 a_n6308_8799.n173 98.9631
R143 a_n6308_8799.n29 a_n6308_8799.n172 98.6055
R144 a_n6308_8799.n28 a_n6308_8799.n86 98.6055
R145 a_n6308_8799.n28 a_n6308_8799.n85 98.6055
R146 a_n6308_8799.n174 a_n6308_8799.n29 98.6054
R147 a_n6308_8799.n1 a_n6308_8799.n87 81.3764
R148 a_n6308_8799.n3 a_n6308_8799.n93 81.3764
R149 a_n6308_8799.n0 a_n6308_8799.n90 81.3764
R150 a_n6308_8799.n2 a_n6308_8799.n96 80.9324
R151 a_n6308_8799.n2 a_n6308_8799.n97 80.9324
R152 a_n6308_8799.n1 a_n6308_8799.n98 80.9324
R153 a_n6308_8799.n1 a_n6308_8799.n89 80.9324
R154 a_n6308_8799.n1 a_n6308_8799.n88 80.9324
R155 a_n6308_8799.n3 a_n6308_8799.n94 80.9324
R156 a_n6308_8799.n0 a_n6308_8799.n95 80.9324
R157 a_n6308_8799.n0 a_n6308_8799.n92 80.9324
R158 a_n6308_8799.n0 a_n6308_8799.n91 80.9324
R159 a_n6308_8799.n31 a_n6308_8799.n143 20.9683
R160 a_n6308_8799.n142 a_n6308_8799.n141 48.2005
R161 a_n6308_8799.n140 a_n6308_8799.n35 20.9683
R162 a_n6308_8799.n137 a_n6308_8799.n136 48.2005
R163 a_n6308_8799.n40 a_n6308_8799.n154 20.9683
R164 a_n6308_8799.n153 a_n6308_8799.n152 48.2005
R165 a_n6308_8799.n151 a_n6308_8799.n44 20.9683
R166 a_n6308_8799.n148 a_n6308_8799.n147 48.2005
R167 a_n6308_8799.n49 a_n6308_8799.n166 20.9683
R168 a_n6308_8799.n165 a_n6308_8799.n164 48.2005
R169 a_n6308_8799.n163 a_n6308_8799.n53 20.9683
R170 a_n6308_8799.n160 a_n6308_8799.n159 48.2005
R171 a_n6308_8799.n103 a_n6308_8799.n102 48.2005
R172 a_n6308_8799.n106 a_n6308_8799.n60 20.9683
R173 a_n6308_8799.n107 a_n6308_8799.n100 48.2005
R174 a_n6308_8799.n109 a_n6308_8799.n64 20.9683
R175 a_n6308_8799.n114 a_n6308_8799.n113 48.2005
R176 a_n6308_8799.n117 a_n6308_8799.n69 20.9683
R177 a_n6308_8799.n118 a_n6308_8799.n111 48.2005
R178 a_n6308_8799.n120 a_n6308_8799.n73 20.9683
R179 a_n6308_8799.n126 a_n6308_8799.n125 48.2005
R180 a_n6308_8799.n129 a_n6308_8799.n78 20.9683
R181 a_n6308_8799.n130 a_n6308_8799.n123 48.2005
R182 a_n6308_8799.n132 a_n6308_8799.n82 20.9683
R183 a_n6308_8799.n33 a_n6308_8799.n134 47.835
R184 a_n6308_8799.n36 a_n6308_8799.n139 20.6913
R185 a_n6308_8799.n42 a_n6308_8799.n145 47.835
R186 a_n6308_8799.n45 a_n6308_8799.n150 20.6913
R187 a_n6308_8799.n51 a_n6308_8799.n157 47.835
R188 a_n6308_8799.n54 a_n6308_8799.n162 20.6913
R189 a_n6308_8799.n101 a_n6308_8799.n59 21.4216
R190 a_n6308_8799.n112 a_n6308_8799.n68 21.4216
R191 a_n6308_8799.n124 a_n6308_8799.n77 21.4216
R192 a_n6308_8799.t42 a_n6308_8799.n65 484.3
R193 a_n6308_8799.t50 a_n6308_8799.n74 484.3
R194 a_n6308_8799.t105 a_n6308_8799.n83 484.3
R195 a_n6308_8799.n58 a_n6308_8799.n104 45.0871
R196 a_n6308_8799.n67 a_n6308_8799.n115 45.0871
R197 a_n6308_8799.n76 a_n6308_8799.n127 45.0871
R198 a_n6308_8799.n38 a_n6308_8799.n138 45.0871
R199 a_n6308_8799.n47 a_n6308_8799.n149 45.0871
R200 a_n6308_8799.n56 a_n6308_8799.n161 45.0871
R201 a_n6308_8799.n2 a_n6308_8799.n0 33.4185
R202 a_n6308_8799.n32 a_n6308_8799.n134 11.843
R203 a_n6308_8799.n139 a_n6308_8799.n37 36.139
R204 a_n6308_8799.n41 a_n6308_8799.n145 11.843
R205 a_n6308_8799.n150 a_n6308_8799.n46 36.139
R206 a_n6308_8799.n50 a_n6308_8799.n157 11.843
R207 a_n6308_8799.n162 a_n6308_8799.n55 36.139
R208 a_n6308_8799.n105 a_n6308_8799.n57 36.139
R209 a_n6308_8799.n99 a_n6308_8799.n63 34.4824
R210 a_n6308_8799.n116 a_n6308_8799.n66 36.139
R211 a_n6308_8799.n110 a_n6308_8799.n72 34.4824
R212 a_n6308_8799.n128 a_n6308_8799.n75 36.139
R213 a_n6308_8799.n122 a_n6308_8799.n81 34.4824
R214 a_n6308_8799.n34 a_n6308_8799.n135 35.3134
R215 a_n6308_8799.n43 a_n6308_8799.n146 35.3134
R216 a_n6308_8799.n52 a_n6308_8799.n158 35.3134
R217 a_n6308_8799.n61 a_n6308_8799.n106 35.3134
R218 a_n6308_8799.n107 a_n6308_8799.n61 11.2134
R219 a_n6308_8799.n70 a_n6308_8799.n117 35.3134
R220 a_n6308_8799.n118 a_n6308_8799.n70 11.2134
R221 a_n6308_8799.n79 a_n6308_8799.n129 35.3134
R222 a_n6308_8799.n130 a_n6308_8799.n79 11.2134
R223 a_n6308_8799.n143 a_n6308_8799.n32 34.4824
R224 a_n6308_8799.n37 a_n6308_8799.n136 10.5784
R225 a_n6308_8799.n154 a_n6308_8799.n41 34.4824
R226 a_n6308_8799.n46 a_n6308_8799.n147 10.5784
R227 a_n6308_8799.n166 a_n6308_8799.n50 34.4824
R228 a_n6308_8799.n55 a_n6308_8799.n159 10.5784
R229 a_n6308_8799.n57 a_n6308_8799.n102 10.5784
R230 a_n6308_8799.n66 a_n6308_8799.n113 10.5784
R231 a_n6308_8799.n75 a_n6308_8799.n125 10.5784
R232 a_n6308_8799.n138 a_n6308_8799.n137 14.1472
R233 a_n6308_8799.n149 a_n6308_8799.n148 14.1472
R234 a_n6308_8799.n161 a_n6308_8799.n160 14.1472
R235 a_n6308_8799.n104 a_n6308_8799.n103 14.1472
R236 a_n6308_8799.n115 a_n6308_8799.n114 14.1472
R237 a_n6308_8799.n127 a_n6308_8799.n126 14.1472
R238 a_n6308_8799.n170 a_n6308_8799.n1 12.3339
R239 a_n6308_8799.n171 a_n6308_8799.n170 11.4887
R240 a_n6308_8799.n156 a_n6308_8799.n26 9.01755
R241 a_n6308_8799.n121 a_n6308_8799.n12 9.01755
R242 a_n6308_8799.n169 a_n6308_8799.n133 6.90212
R243 a_n6308_8799.n169 a_n6308_8799.n168 6.48069
R244 a_n6308_8799.n156 a_n6308_8799.n22 4.90959
R245 a_n6308_8799.n168 a_n6308_8799.n18 4.90959
R246 a_n6308_8799.n121 a_n6308_8799.n8 4.90959
R247 a_n6308_8799.n133 a_n6308_8799.n4 4.90959
R248 a_n6308_8799.n168 a_n6308_8799.n156 4.10845
R249 a_n6308_8799.n133 a_n6308_8799.n121 4.10845
R250 a_n6308_8799.n173 a_n6308_8799.t12 3.61217
R251 a_n6308_8799.n173 a_n6308_8799.t27 3.61217
R252 a_n6308_8799.n172 a_n6308_8799.t13 3.61217
R253 a_n6308_8799.n172 a_n6308_8799.t14 3.61217
R254 a_n6308_8799.n86 a_n6308_8799.t5 3.61217
R255 a_n6308_8799.n86 a_n6308_8799.t29 3.61217
R256 a_n6308_8799.n85 a_n6308_8799.t6 3.61217
R257 a_n6308_8799.n85 a_n6308_8799.t28 3.61217
R258 a_n6308_8799.n84 a_n6308_8799.t8 3.61217
R259 a_n6308_8799.n84 a_n6308_8799.t23 3.61217
R260 a_n6308_8799.t4 a_n6308_8799.n174 3.61217
R261 a_n6308_8799.n174 a_n6308_8799.t22 3.61217
R262 a_n6308_8799.n170 a_n6308_8799.n169 3.4105
R263 a_n6308_8799.n96 a_n6308_8799.t20 2.82907
R264 a_n6308_8799.n96 a_n6308_8799.t31 2.82907
R265 a_n6308_8799.n97 a_n6308_8799.t0 2.82907
R266 a_n6308_8799.n97 a_n6308_8799.t7 2.82907
R267 a_n6308_8799.n98 a_n6308_8799.t16 2.82907
R268 a_n6308_8799.n98 a_n6308_8799.t26 2.82907
R269 a_n6308_8799.n89 a_n6308_8799.t30 2.82907
R270 a_n6308_8799.n89 a_n6308_8799.t11 2.82907
R271 a_n6308_8799.n88 a_n6308_8799.t17 2.82907
R272 a_n6308_8799.n88 a_n6308_8799.t34 2.82907
R273 a_n6308_8799.n87 a_n6308_8799.t25 2.82907
R274 a_n6308_8799.n87 a_n6308_8799.t2 2.82907
R275 a_n6308_8799.n93 a_n6308_8799.t32 2.82907
R276 a_n6308_8799.n93 a_n6308_8799.t19 2.82907
R277 a_n6308_8799.n94 a_n6308_8799.t3 2.82907
R278 a_n6308_8799.n94 a_n6308_8799.t33 2.82907
R279 a_n6308_8799.n95 a_n6308_8799.t24 2.82907
R280 a_n6308_8799.n95 a_n6308_8799.t35 2.82907
R281 a_n6308_8799.n92 a_n6308_8799.t15 2.82907
R282 a_n6308_8799.n92 a_n6308_8799.t21 2.82907
R283 a_n6308_8799.n91 a_n6308_8799.t10 2.82907
R284 a_n6308_8799.n91 a_n6308_8799.t9 2.82907
R285 a_n6308_8799.n90 a_n6308_8799.t18 2.82907
R286 a_n6308_8799.n90 a_n6308_8799.t1 2.82907
R287 a_n6308_8799.n30 a_n6308_8799.n144 22.3251
R288 a_n6308_8799.n39 a_n6308_8799.n155 22.3251
R289 a_n6308_8799.n48 a_n6308_8799.n167 22.3251
R290 a_n6308_8799.n65 a_n6308_8799.n109 22.3251
R291 a_n6308_8799.n74 a_n6308_8799.n120 22.3251
R292 a_n6308_8799.n83 a_n6308_8799.n132 22.3251
R293 a_n6308_8799.n33 a_n6308_8799.n142 0.365327
R294 a_n6308_8799.n140 a_n6308_8799.n36 21.4216
R295 a_n6308_8799.n42 a_n6308_8799.n153 0.365327
R296 a_n6308_8799.n151 a_n6308_8799.n45 21.4216
R297 a_n6308_8799.n51 a_n6308_8799.n165 0.365327
R298 a_n6308_8799.n163 a_n6308_8799.n54 21.4216
R299 a_n6308_8799.n108 a_n6308_8799.n62 47.835
R300 a_n6308_8799.n119 a_n6308_8799.n71 47.835
R301 a_n6308_8799.n131 a_n6308_8799.n80 47.835
R302 a_n6308_8799.n29 a_n6308_8799.n171 31.2933
R303 a_n6308_8799.n171 a_n6308_8799.n28 17.8718
R304 a_n6308_8799.n1 a_n6308_8799.n2 1.77636
R305 a_n6308_8799.n0 a_n6308_8799.n3 1.3324
R306 a_n6308_8799.n27 a_n6308_8799.n25 0.758076
R307 a_n6308_8799.n25 a_n6308_8799.n24 0.758076
R308 a_n6308_8799.n38 a_n6308_8799.n24 0.758076
R309 a_n6308_8799.n23 a_n6308_8799.n21 0.758076
R310 a_n6308_8799.n21 a_n6308_8799.n20 0.758076
R311 a_n6308_8799.n47 a_n6308_8799.n20 0.758076
R312 a_n6308_8799.n19 a_n6308_8799.n17 0.758076
R313 a_n6308_8799.n17 a_n6308_8799.n16 0.758076
R314 a_n6308_8799.n56 a_n6308_8799.n16 0.758076
R315 a_n6308_8799.n15 a_n6308_8799.n14 0.758076
R316 a_n6308_8799.n14 a_n6308_8799.n13 0.758076
R317 a_n6308_8799.n13 a_n6308_8799.n12 0.758076
R318 a_n6308_8799.n11 a_n6308_8799.n10 0.758076
R319 a_n6308_8799.n10 a_n6308_8799.n9 0.758076
R320 a_n6308_8799.n9 a_n6308_8799.n8 0.758076
R321 a_n6308_8799.n7 a_n6308_8799.n6 0.758076
R322 a_n6308_8799.n6 a_n6308_8799.n5 0.758076
R323 a_n6308_8799.n5 a_n6308_8799.n4 0.758076
R324 a_n6308_8799.n76 a_n6308_8799.n7 0.568682
R325 a_n6308_8799.n67 a_n6308_8799.n11 0.568682
R326 a_n6308_8799.n58 a_n6308_8799.n15 0.568682
R327 a_n6308_8799.n19 a_n6308_8799.n18 0.568682
R328 a_n6308_8799.n23 a_n6308_8799.n22 0.568682
R329 a_n6308_8799.n27 a_n6308_8799.n26 0.568682
R330 vdd.n303 vdd.n267 756.745
R331 vdd.n252 vdd.n216 756.745
R332 vdd.n209 vdd.n173 756.745
R333 vdd.n158 vdd.n122 756.745
R334 vdd.n116 vdd.n80 756.745
R335 vdd.n65 vdd.n29 756.745
R336 vdd.n1498 vdd.n1462 756.745
R337 vdd.n1549 vdd.n1513 756.745
R338 vdd.n1404 vdd.n1368 756.745
R339 vdd.n1455 vdd.n1419 756.745
R340 vdd.n1311 vdd.n1275 756.745
R341 vdd.n1362 vdd.n1326 756.745
R342 vdd.n1889 vdd.t57 640.208
R343 vdd.n793 vdd.t42 640.208
R344 vdd.n1863 vdd.t7 640.208
R345 vdd.n785 vdd.t67 640.208
R346 vdd.n2634 vdd.t29 640.208
R347 vdd.n2354 vdd.t64 640.208
R348 vdd.n661 vdd.t46 640.208
R349 vdd.n2351 vdd.t50 640.208
R350 vdd.n625 vdd.t54 640.208
R351 vdd.n855 vdd.t60 640.208
R352 vdd.n1110 vdd.t3 592.009
R353 vdd.n1147 vdd.t26 592.009
R354 vdd.n1021 vdd.t36 592.009
R355 vdd.n2045 vdd.t22 592.009
R356 vdd.n1682 vdd.t33 592.009
R357 vdd.n1642 vdd.t39 592.009
R358 vdd.n3021 vdd.t76 592.009
R359 vdd.n427 vdd.t73 592.009
R360 vdd.n387 vdd.t11 592.009
R361 vdd.n580 vdd.t15 592.009
R362 vdd.n543 vdd.t19 592.009
R363 vdd.n2808 vdd.t70 592.009
R364 vdd.n304 vdd.n303 585
R365 vdd.n302 vdd.n269 585
R366 vdd.n301 vdd.n300 585
R367 vdd.n272 vdd.n270 585
R368 vdd.n295 vdd.n294 585
R369 vdd.n293 vdd.n292 585
R370 vdd.n276 vdd.n275 585
R371 vdd.n287 vdd.n286 585
R372 vdd.n285 vdd.n284 585
R373 vdd.n280 vdd.n279 585
R374 vdd.n253 vdd.n252 585
R375 vdd.n251 vdd.n218 585
R376 vdd.n250 vdd.n249 585
R377 vdd.n221 vdd.n219 585
R378 vdd.n244 vdd.n243 585
R379 vdd.n242 vdd.n241 585
R380 vdd.n225 vdd.n224 585
R381 vdd.n236 vdd.n235 585
R382 vdd.n234 vdd.n233 585
R383 vdd.n229 vdd.n228 585
R384 vdd.n210 vdd.n209 585
R385 vdd.n208 vdd.n175 585
R386 vdd.n207 vdd.n206 585
R387 vdd.n178 vdd.n176 585
R388 vdd.n201 vdd.n200 585
R389 vdd.n199 vdd.n198 585
R390 vdd.n182 vdd.n181 585
R391 vdd.n193 vdd.n192 585
R392 vdd.n191 vdd.n190 585
R393 vdd.n186 vdd.n185 585
R394 vdd.n159 vdd.n158 585
R395 vdd.n157 vdd.n124 585
R396 vdd.n156 vdd.n155 585
R397 vdd.n127 vdd.n125 585
R398 vdd.n150 vdd.n149 585
R399 vdd.n148 vdd.n147 585
R400 vdd.n131 vdd.n130 585
R401 vdd.n142 vdd.n141 585
R402 vdd.n140 vdd.n139 585
R403 vdd.n135 vdd.n134 585
R404 vdd.n117 vdd.n116 585
R405 vdd.n115 vdd.n82 585
R406 vdd.n114 vdd.n113 585
R407 vdd.n85 vdd.n83 585
R408 vdd.n108 vdd.n107 585
R409 vdd.n106 vdd.n105 585
R410 vdd.n89 vdd.n88 585
R411 vdd.n100 vdd.n99 585
R412 vdd.n98 vdd.n97 585
R413 vdd.n93 vdd.n92 585
R414 vdd.n66 vdd.n65 585
R415 vdd.n64 vdd.n31 585
R416 vdd.n63 vdd.n62 585
R417 vdd.n34 vdd.n32 585
R418 vdd.n57 vdd.n56 585
R419 vdd.n55 vdd.n54 585
R420 vdd.n38 vdd.n37 585
R421 vdd.n49 vdd.n48 585
R422 vdd.n47 vdd.n46 585
R423 vdd.n42 vdd.n41 585
R424 vdd.n1499 vdd.n1498 585
R425 vdd.n1497 vdd.n1464 585
R426 vdd.n1496 vdd.n1495 585
R427 vdd.n1467 vdd.n1465 585
R428 vdd.n1490 vdd.n1489 585
R429 vdd.n1488 vdd.n1487 585
R430 vdd.n1471 vdd.n1470 585
R431 vdd.n1482 vdd.n1481 585
R432 vdd.n1480 vdd.n1479 585
R433 vdd.n1475 vdd.n1474 585
R434 vdd.n1550 vdd.n1549 585
R435 vdd.n1548 vdd.n1515 585
R436 vdd.n1547 vdd.n1546 585
R437 vdd.n1518 vdd.n1516 585
R438 vdd.n1541 vdd.n1540 585
R439 vdd.n1539 vdd.n1538 585
R440 vdd.n1522 vdd.n1521 585
R441 vdd.n1533 vdd.n1532 585
R442 vdd.n1531 vdd.n1530 585
R443 vdd.n1526 vdd.n1525 585
R444 vdd.n1405 vdd.n1404 585
R445 vdd.n1403 vdd.n1370 585
R446 vdd.n1402 vdd.n1401 585
R447 vdd.n1373 vdd.n1371 585
R448 vdd.n1396 vdd.n1395 585
R449 vdd.n1394 vdd.n1393 585
R450 vdd.n1377 vdd.n1376 585
R451 vdd.n1388 vdd.n1387 585
R452 vdd.n1386 vdd.n1385 585
R453 vdd.n1381 vdd.n1380 585
R454 vdd.n1456 vdd.n1455 585
R455 vdd.n1454 vdd.n1421 585
R456 vdd.n1453 vdd.n1452 585
R457 vdd.n1424 vdd.n1422 585
R458 vdd.n1447 vdd.n1446 585
R459 vdd.n1445 vdd.n1444 585
R460 vdd.n1428 vdd.n1427 585
R461 vdd.n1439 vdd.n1438 585
R462 vdd.n1437 vdd.n1436 585
R463 vdd.n1432 vdd.n1431 585
R464 vdd.n1312 vdd.n1311 585
R465 vdd.n1310 vdd.n1277 585
R466 vdd.n1309 vdd.n1308 585
R467 vdd.n1280 vdd.n1278 585
R468 vdd.n1303 vdd.n1302 585
R469 vdd.n1301 vdd.n1300 585
R470 vdd.n1284 vdd.n1283 585
R471 vdd.n1295 vdd.n1294 585
R472 vdd.n1293 vdd.n1292 585
R473 vdd.n1288 vdd.n1287 585
R474 vdd.n1363 vdd.n1362 585
R475 vdd.n1361 vdd.n1328 585
R476 vdd.n1360 vdd.n1359 585
R477 vdd.n1331 vdd.n1329 585
R478 vdd.n1354 vdd.n1353 585
R479 vdd.n1352 vdd.n1351 585
R480 vdd.n1335 vdd.n1334 585
R481 vdd.n1346 vdd.n1345 585
R482 vdd.n1344 vdd.n1343 585
R483 vdd.n1339 vdd.n1338 585
R484 vdd.n3137 vdd.n352 488.781
R485 vdd.n3019 vdd.n350 488.781
R486 vdd.n2941 vdd.n515 488.781
R487 vdd.n2939 vdd.n517 488.781
R488 vdd.n2040 vdd.n903 488.781
R489 vdd.n2043 vdd.n2042 488.781
R490 vdd.n1216 vdd.n981 488.781
R491 vdd.n1214 vdd.n984 488.781
R492 vdd.n281 vdd.t173 329.043
R493 vdd.n230 vdd.t191 329.043
R494 vdd.n187 vdd.t166 329.043
R495 vdd.n136 vdd.t186 329.043
R496 vdd.n94 vdd.t154 329.043
R497 vdd.n43 vdd.t135 329.043
R498 vdd.n1476 vdd.t224 329.043
R499 vdd.n1527 vdd.t203 329.043
R500 vdd.n1382 vdd.t212 329.043
R501 vdd.n1433 vdd.t194 329.043
R502 vdd.n1289 vdd.t137 329.043
R503 vdd.n1340 vdd.t156 329.043
R504 vdd.n1110 vdd.t6 319.788
R505 vdd.n1147 vdd.t28 319.788
R506 vdd.n1021 vdd.t38 319.788
R507 vdd.n2045 vdd.t24 319.788
R508 vdd.n1682 vdd.t34 319.788
R509 vdd.n1642 vdd.t40 319.788
R510 vdd.n3021 vdd.t77 319.788
R511 vdd.n427 vdd.t74 319.788
R512 vdd.n387 vdd.t13 319.788
R513 vdd.n580 vdd.t18 319.788
R514 vdd.n543 vdd.t21 319.788
R515 vdd.n2808 vdd.t72 319.788
R516 vdd.n1111 vdd.t5 303.69
R517 vdd.n1148 vdd.t27 303.69
R518 vdd.n1022 vdd.t37 303.69
R519 vdd.n2046 vdd.t25 303.69
R520 vdd.n1683 vdd.t35 303.69
R521 vdd.n1643 vdd.t41 303.69
R522 vdd.n3022 vdd.t78 303.69
R523 vdd.n428 vdd.t75 303.69
R524 vdd.n388 vdd.t14 303.69
R525 vdd.n581 vdd.t17 303.69
R526 vdd.n544 vdd.t20 303.69
R527 vdd.n2809 vdd.t71 303.69
R528 vdd.n2577 vdd.n741 297.074
R529 vdd.n2770 vdd.n635 297.074
R530 vdd.n2707 vdd.n632 297.074
R531 vdd.n2500 vdd.n742 297.074
R532 vdd.n2315 vdd.n782 297.074
R533 vdd.n2246 vdd.n2245 297.074
R534 vdd.n1992 vdd.n878 297.074
R535 vdd.n2088 vdd.n876 297.074
R536 vdd.n2686 vdd.n633 297.074
R537 vdd.n2773 vdd.n2772 297.074
R538 vdd.n2349 vdd.n743 297.074
R539 vdd.n2575 vdd.n744 297.074
R540 vdd.n2243 vdd.n791 297.074
R541 vdd.n789 vdd.n764 297.074
R542 vdd.n1929 vdd.n879 297.074
R543 vdd.n2086 vdd.n880 297.074
R544 vdd.n2688 vdd.n633 185
R545 vdd.n2771 vdd.n633 185
R546 vdd.n2690 vdd.n2689 185
R547 vdd.n2689 vdd.n631 185
R548 vdd.n2691 vdd.n667 185
R549 vdd.n2701 vdd.n667 185
R550 vdd.n2692 vdd.n676 185
R551 vdd.n676 vdd.n674 185
R552 vdd.n2694 vdd.n2693 185
R553 vdd.n2695 vdd.n2694 185
R554 vdd.n2647 vdd.n675 185
R555 vdd.n675 vdd.n671 185
R556 vdd.n2646 vdd.n2645 185
R557 vdd.n2645 vdd.n2644 185
R558 vdd.n678 vdd.n677 185
R559 vdd.n679 vdd.n678 185
R560 vdd.n2637 vdd.n2636 185
R561 vdd.n2638 vdd.n2637 185
R562 vdd.n2633 vdd.n688 185
R563 vdd.n688 vdd.n685 185
R564 vdd.n2632 vdd.n2631 185
R565 vdd.n2631 vdd.n2630 185
R566 vdd.n690 vdd.n689 185
R567 vdd.n698 vdd.n690 185
R568 vdd.n2623 vdd.n2622 185
R569 vdd.n2624 vdd.n2623 185
R570 vdd.n2621 vdd.n699 185
R571 vdd.n2472 vdd.n699 185
R572 vdd.n2620 vdd.n2619 185
R573 vdd.n2619 vdd.n2618 185
R574 vdd.n701 vdd.n700 185
R575 vdd.n702 vdd.n701 185
R576 vdd.n2611 vdd.n2610 185
R577 vdd.n2612 vdd.n2611 185
R578 vdd.n2609 vdd.n711 185
R579 vdd.n711 vdd.n708 185
R580 vdd.n2608 vdd.n2607 185
R581 vdd.n2607 vdd.n2606 185
R582 vdd.n713 vdd.n712 185
R583 vdd.n721 vdd.n713 185
R584 vdd.n2599 vdd.n2598 185
R585 vdd.n2600 vdd.n2599 185
R586 vdd.n2597 vdd.n722 185
R587 vdd.n728 vdd.n722 185
R588 vdd.n2596 vdd.n2595 185
R589 vdd.n2595 vdd.n2594 185
R590 vdd.n724 vdd.n723 185
R591 vdd.n725 vdd.n724 185
R592 vdd.n2587 vdd.n2586 185
R593 vdd.n2588 vdd.n2587 185
R594 vdd.n2585 vdd.n734 185
R595 vdd.n2493 vdd.n734 185
R596 vdd.n2584 vdd.n2583 185
R597 vdd.n2583 vdd.n2582 185
R598 vdd.n736 vdd.n735 185
R599 vdd.t87 vdd.n736 185
R600 vdd.n2575 vdd.n2574 185
R601 vdd.n2576 vdd.n2575 185
R602 vdd.n2573 vdd.n744 185
R603 vdd.n2572 vdd.n2571 185
R604 vdd.n746 vdd.n745 185
R605 vdd.n2358 vdd.n2357 185
R606 vdd.n2360 vdd.n2359 185
R607 vdd.n2362 vdd.n2361 185
R608 vdd.n2364 vdd.n2363 185
R609 vdd.n2366 vdd.n2365 185
R610 vdd.n2368 vdd.n2367 185
R611 vdd.n2370 vdd.n2369 185
R612 vdd.n2372 vdd.n2371 185
R613 vdd.n2374 vdd.n2373 185
R614 vdd.n2376 vdd.n2375 185
R615 vdd.n2378 vdd.n2377 185
R616 vdd.n2380 vdd.n2379 185
R617 vdd.n2382 vdd.n2381 185
R618 vdd.n2384 vdd.n2383 185
R619 vdd.n2386 vdd.n2385 185
R620 vdd.n2388 vdd.n2387 185
R621 vdd.n2390 vdd.n2389 185
R622 vdd.n2392 vdd.n2391 185
R623 vdd.n2394 vdd.n2393 185
R624 vdd.n2396 vdd.n2395 185
R625 vdd.n2398 vdd.n2397 185
R626 vdd.n2400 vdd.n2399 185
R627 vdd.n2402 vdd.n2401 185
R628 vdd.n2404 vdd.n2403 185
R629 vdd.n2406 vdd.n2405 185
R630 vdd.n2408 vdd.n2407 185
R631 vdd.n2410 vdd.n2409 185
R632 vdd.n2412 vdd.n2411 185
R633 vdd.n2414 vdd.n2413 185
R634 vdd.n2416 vdd.n2415 185
R635 vdd.n2418 vdd.n2417 185
R636 vdd.n2419 vdd.n2349 185
R637 vdd.n2569 vdd.n2349 185
R638 vdd.n2774 vdd.n2773 185
R639 vdd.n2775 vdd.n624 185
R640 vdd.n2777 vdd.n2776 185
R641 vdd.n2779 vdd.n622 185
R642 vdd.n2781 vdd.n2780 185
R643 vdd.n2782 vdd.n621 185
R644 vdd.n2784 vdd.n2783 185
R645 vdd.n2786 vdd.n619 185
R646 vdd.n2788 vdd.n2787 185
R647 vdd.n2789 vdd.n618 185
R648 vdd.n2791 vdd.n2790 185
R649 vdd.n2793 vdd.n616 185
R650 vdd.n2795 vdd.n2794 185
R651 vdd.n2796 vdd.n615 185
R652 vdd.n2798 vdd.n2797 185
R653 vdd.n2800 vdd.n614 185
R654 vdd.n2801 vdd.n611 185
R655 vdd.n2804 vdd.n2803 185
R656 vdd.n612 vdd.n610 185
R657 vdd.n2660 vdd.n2659 185
R658 vdd.n2662 vdd.n2661 185
R659 vdd.n2664 vdd.n2656 185
R660 vdd.n2666 vdd.n2665 185
R661 vdd.n2667 vdd.n2655 185
R662 vdd.n2669 vdd.n2668 185
R663 vdd.n2671 vdd.n2653 185
R664 vdd.n2673 vdd.n2672 185
R665 vdd.n2674 vdd.n2652 185
R666 vdd.n2676 vdd.n2675 185
R667 vdd.n2678 vdd.n2650 185
R668 vdd.n2680 vdd.n2679 185
R669 vdd.n2681 vdd.n2649 185
R670 vdd.n2683 vdd.n2682 185
R671 vdd.n2685 vdd.n2648 185
R672 vdd.n2687 vdd.n2686 185
R673 vdd.n2686 vdd.n613 185
R674 vdd.n2772 vdd.n628 185
R675 vdd.n2772 vdd.n2771 185
R676 vdd.n2424 vdd.n630 185
R677 vdd.n631 vdd.n630 185
R678 vdd.n2425 vdd.n666 185
R679 vdd.n2701 vdd.n666 185
R680 vdd.n2427 vdd.n2426 185
R681 vdd.n2426 vdd.n674 185
R682 vdd.n2428 vdd.n673 185
R683 vdd.n2695 vdd.n673 185
R684 vdd.n2430 vdd.n2429 185
R685 vdd.n2429 vdd.n671 185
R686 vdd.n2431 vdd.n681 185
R687 vdd.n2644 vdd.n681 185
R688 vdd.n2433 vdd.n2432 185
R689 vdd.n2432 vdd.n679 185
R690 vdd.n2434 vdd.n687 185
R691 vdd.n2638 vdd.n687 185
R692 vdd.n2436 vdd.n2435 185
R693 vdd.n2435 vdd.n685 185
R694 vdd.n2437 vdd.n692 185
R695 vdd.n2630 vdd.n692 185
R696 vdd.n2439 vdd.n2438 185
R697 vdd.n2438 vdd.n698 185
R698 vdd.n2440 vdd.n697 185
R699 vdd.n2624 vdd.n697 185
R700 vdd.n2474 vdd.n2473 185
R701 vdd.n2473 vdd.n2472 185
R702 vdd.n2475 vdd.n704 185
R703 vdd.n2618 vdd.n704 185
R704 vdd.n2477 vdd.n2476 185
R705 vdd.n2476 vdd.n702 185
R706 vdd.n2478 vdd.n710 185
R707 vdd.n2612 vdd.n710 185
R708 vdd.n2480 vdd.n2479 185
R709 vdd.n2479 vdd.n708 185
R710 vdd.n2481 vdd.n715 185
R711 vdd.n2606 vdd.n715 185
R712 vdd.n2483 vdd.n2482 185
R713 vdd.n2482 vdd.n721 185
R714 vdd.n2484 vdd.n720 185
R715 vdd.n2600 vdd.n720 185
R716 vdd.n2486 vdd.n2485 185
R717 vdd.n2485 vdd.n728 185
R718 vdd.n2487 vdd.n727 185
R719 vdd.n2594 vdd.n727 185
R720 vdd.n2489 vdd.n2488 185
R721 vdd.n2488 vdd.n725 185
R722 vdd.n2490 vdd.n733 185
R723 vdd.n2588 vdd.n733 185
R724 vdd.n2492 vdd.n2491 185
R725 vdd.n2493 vdd.n2492 185
R726 vdd.n2423 vdd.n738 185
R727 vdd.n2582 vdd.n738 185
R728 vdd.n2422 vdd.n2421 185
R729 vdd.n2421 vdd.t87 185
R730 vdd.n2420 vdd.n743 185
R731 vdd.n2576 vdd.n743 185
R732 vdd.n2040 vdd.n2039 185
R733 vdd.n2041 vdd.n2040 185
R734 vdd.n904 vdd.n902 185
R735 vdd.n1606 vdd.n902 185
R736 vdd.n1609 vdd.n1608 185
R737 vdd.n1608 vdd.n1607 185
R738 vdd.n907 vdd.n906 185
R739 vdd.n908 vdd.n907 185
R740 vdd.n1595 vdd.n1594 185
R741 vdd.n1596 vdd.n1595 185
R742 vdd.n916 vdd.n915 185
R743 vdd.n1587 vdd.n915 185
R744 vdd.n1590 vdd.n1589 185
R745 vdd.n1589 vdd.n1588 185
R746 vdd.n919 vdd.n918 185
R747 vdd.n925 vdd.n919 185
R748 vdd.n1578 vdd.n1577 185
R749 vdd.n1579 vdd.n1578 185
R750 vdd.n927 vdd.n926 185
R751 vdd.n1570 vdd.n926 185
R752 vdd.n1573 vdd.n1572 185
R753 vdd.n1572 vdd.n1571 185
R754 vdd.n930 vdd.n929 185
R755 vdd.n931 vdd.n930 185
R756 vdd.n1561 vdd.n1560 185
R757 vdd.n1562 vdd.n1561 185
R758 vdd.n939 vdd.n938 185
R759 vdd.n938 vdd.n937 185
R760 vdd.n1274 vdd.n1273 185
R761 vdd.n1273 vdd.n1272 185
R762 vdd.n942 vdd.n941 185
R763 vdd.n948 vdd.n942 185
R764 vdd.n1263 vdd.n1262 185
R765 vdd.n1264 vdd.n1263 185
R766 vdd.n950 vdd.n949 185
R767 vdd.n1255 vdd.n949 185
R768 vdd.n1258 vdd.n1257 185
R769 vdd.n1257 vdd.n1256 185
R770 vdd.n953 vdd.n952 185
R771 vdd.n960 vdd.n953 185
R772 vdd.n1246 vdd.n1245 185
R773 vdd.n1247 vdd.n1246 185
R774 vdd.n962 vdd.n961 185
R775 vdd.n961 vdd.n959 185
R776 vdd.n1241 vdd.n1240 185
R777 vdd.n1240 vdd.n1239 185
R778 vdd.n965 vdd.n964 185
R779 vdd.n966 vdd.n965 185
R780 vdd.n1230 vdd.n1229 185
R781 vdd.n1231 vdd.n1230 185
R782 vdd.n974 vdd.n973 185
R783 vdd.n973 vdd.n972 185
R784 vdd.n1225 vdd.n1224 185
R785 vdd.n1224 vdd.n1223 185
R786 vdd.n977 vdd.n976 185
R787 vdd.n983 vdd.n977 185
R788 vdd.n1214 vdd.n1213 185
R789 vdd.n1215 vdd.n1214 185
R790 vdd.n1210 vdd.n984 185
R791 vdd.n1209 vdd.n987 185
R792 vdd.n1208 vdd.n988 185
R793 vdd.n988 vdd.n982 185
R794 vdd.n991 vdd.n989 185
R795 vdd.n1204 vdd.n993 185
R796 vdd.n1203 vdd.n994 185
R797 vdd.n1202 vdd.n996 185
R798 vdd.n999 vdd.n997 185
R799 vdd.n1198 vdd.n1001 185
R800 vdd.n1197 vdd.n1002 185
R801 vdd.n1196 vdd.n1004 185
R802 vdd.n1007 vdd.n1005 185
R803 vdd.n1192 vdd.n1009 185
R804 vdd.n1191 vdd.n1010 185
R805 vdd.n1190 vdd.n1012 185
R806 vdd.n1015 vdd.n1013 185
R807 vdd.n1186 vdd.n1017 185
R808 vdd.n1185 vdd.n1018 185
R809 vdd.n1184 vdd.n1020 185
R810 vdd.n1025 vdd.n1023 185
R811 vdd.n1180 vdd.n1027 185
R812 vdd.n1179 vdd.n1028 185
R813 vdd.n1178 vdd.n1030 185
R814 vdd.n1033 vdd.n1031 185
R815 vdd.n1174 vdd.n1035 185
R816 vdd.n1173 vdd.n1036 185
R817 vdd.n1172 vdd.n1038 185
R818 vdd.n1041 vdd.n1039 185
R819 vdd.n1168 vdd.n1043 185
R820 vdd.n1167 vdd.n1044 185
R821 vdd.n1166 vdd.n1046 185
R822 vdd.n1049 vdd.n1047 185
R823 vdd.n1162 vdd.n1051 185
R824 vdd.n1161 vdd.n1052 185
R825 vdd.n1160 vdd.n1054 185
R826 vdd.n1057 vdd.n1055 185
R827 vdd.n1156 vdd.n1059 185
R828 vdd.n1155 vdd.n1060 185
R829 vdd.n1154 vdd.n1062 185
R830 vdd.n1065 vdd.n1063 185
R831 vdd.n1150 vdd.n1067 185
R832 vdd.n1149 vdd.n1146 185
R833 vdd.n1144 vdd.n1068 185
R834 vdd.n1143 vdd.n1142 185
R835 vdd.n1073 vdd.n1070 185
R836 vdd.n1138 vdd.n1074 185
R837 vdd.n1137 vdd.n1076 185
R838 vdd.n1136 vdd.n1077 185
R839 vdd.n1081 vdd.n1078 185
R840 vdd.n1132 vdd.n1082 185
R841 vdd.n1131 vdd.n1084 185
R842 vdd.n1130 vdd.n1085 185
R843 vdd.n1089 vdd.n1086 185
R844 vdd.n1126 vdd.n1090 185
R845 vdd.n1125 vdd.n1092 185
R846 vdd.n1124 vdd.n1093 185
R847 vdd.n1097 vdd.n1094 185
R848 vdd.n1120 vdd.n1098 185
R849 vdd.n1119 vdd.n1100 185
R850 vdd.n1118 vdd.n1101 185
R851 vdd.n1105 vdd.n1102 185
R852 vdd.n1114 vdd.n1106 185
R853 vdd.n1113 vdd.n1108 185
R854 vdd.n1109 vdd.n981 185
R855 vdd.n982 vdd.n981 185
R856 vdd.n2044 vdd.n2043 185
R857 vdd.n2048 vdd.n897 185
R858 vdd.n1711 vdd.n896 185
R859 vdd.n1714 vdd.n1713 185
R860 vdd.n1716 vdd.n1715 185
R861 vdd.n1719 vdd.n1718 185
R862 vdd.n1721 vdd.n1720 185
R863 vdd.n1723 vdd.n1709 185
R864 vdd.n1725 vdd.n1724 185
R865 vdd.n1726 vdd.n1703 185
R866 vdd.n1728 vdd.n1727 185
R867 vdd.n1730 vdd.n1701 185
R868 vdd.n1732 vdd.n1731 185
R869 vdd.n1733 vdd.n1696 185
R870 vdd.n1735 vdd.n1734 185
R871 vdd.n1737 vdd.n1694 185
R872 vdd.n1739 vdd.n1738 185
R873 vdd.n1740 vdd.n1690 185
R874 vdd.n1742 vdd.n1741 185
R875 vdd.n1744 vdd.n1687 185
R876 vdd.n1746 vdd.n1745 185
R877 vdd.n1688 vdd.n1681 185
R878 vdd.n1750 vdd.n1685 185
R879 vdd.n1751 vdd.n1677 185
R880 vdd.n1753 vdd.n1752 185
R881 vdd.n1755 vdd.n1675 185
R882 vdd.n1757 vdd.n1756 185
R883 vdd.n1758 vdd.n1670 185
R884 vdd.n1760 vdd.n1759 185
R885 vdd.n1762 vdd.n1668 185
R886 vdd.n1764 vdd.n1763 185
R887 vdd.n1765 vdd.n1663 185
R888 vdd.n1767 vdd.n1766 185
R889 vdd.n1769 vdd.n1661 185
R890 vdd.n1771 vdd.n1770 185
R891 vdd.n1772 vdd.n1656 185
R892 vdd.n1774 vdd.n1773 185
R893 vdd.n1776 vdd.n1654 185
R894 vdd.n1778 vdd.n1777 185
R895 vdd.n1779 vdd.n1650 185
R896 vdd.n1781 vdd.n1780 185
R897 vdd.n1783 vdd.n1647 185
R898 vdd.n1785 vdd.n1784 185
R899 vdd.n1648 vdd.n1641 185
R900 vdd.n1789 vdd.n1645 185
R901 vdd.n1790 vdd.n1637 185
R902 vdd.n1792 vdd.n1791 185
R903 vdd.n1794 vdd.n1635 185
R904 vdd.n1796 vdd.n1795 185
R905 vdd.n1797 vdd.n1630 185
R906 vdd.n1799 vdd.n1798 185
R907 vdd.n1801 vdd.n1628 185
R908 vdd.n1803 vdd.n1802 185
R909 vdd.n1804 vdd.n1623 185
R910 vdd.n1806 vdd.n1805 185
R911 vdd.n1808 vdd.n1622 185
R912 vdd.n1809 vdd.n1619 185
R913 vdd.n1812 vdd.n1811 185
R914 vdd.n1621 vdd.n1617 185
R915 vdd.n2029 vdd.n1615 185
R916 vdd.n2031 vdd.n2030 185
R917 vdd.n2033 vdd.n1613 185
R918 vdd.n2035 vdd.n2034 185
R919 vdd.n2036 vdd.n903 185
R920 vdd.n2042 vdd.n900 185
R921 vdd.n2042 vdd.n2041 185
R922 vdd.n911 vdd.n899 185
R923 vdd.n1606 vdd.n899 185
R924 vdd.n1605 vdd.n1604 185
R925 vdd.n1607 vdd.n1605 185
R926 vdd.n910 vdd.n909 185
R927 vdd.n909 vdd.n908 185
R928 vdd.n1598 vdd.n1597 185
R929 vdd.n1597 vdd.n1596 185
R930 vdd.n914 vdd.n913 185
R931 vdd.n1587 vdd.n914 185
R932 vdd.n1586 vdd.n1585 185
R933 vdd.n1588 vdd.n1586 185
R934 vdd.n921 vdd.n920 185
R935 vdd.n925 vdd.n920 185
R936 vdd.n1581 vdd.n1580 185
R937 vdd.n1580 vdd.n1579 185
R938 vdd.n924 vdd.n923 185
R939 vdd.n1570 vdd.n924 185
R940 vdd.n1569 vdd.n1568 185
R941 vdd.n1571 vdd.n1569 185
R942 vdd.n933 vdd.n932 185
R943 vdd.n932 vdd.n931 185
R944 vdd.n1564 vdd.n1563 185
R945 vdd.n1563 vdd.n1562 185
R946 vdd.n936 vdd.n935 185
R947 vdd.n937 vdd.n936 185
R948 vdd.n1271 vdd.n1270 185
R949 vdd.n1272 vdd.n1271 185
R950 vdd.n944 vdd.n943 185
R951 vdd.n948 vdd.n943 185
R952 vdd.n1266 vdd.n1265 185
R953 vdd.n1265 vdd.n1264 185
R954 vdd.n947 vdd.n946 185
R955 vdd.n1255 vdd.n947 185
R956 vdd.n1254 vdd.n1253 185
R957 vdd.n1256 vdd.n1254 185
R958 vdd.n955 vdd.n954 185
R959 vdd.n960 vdd.n954 185
R960 vdd.n1249 vdd.n1248 185
R961 vdd.n1248 vdd.n1247 185
R962 vdd.n958 vdd.n957 185
R963 vdd.n959 vdd.n958 185
R964 vdd.n1238 vdd.n1237 185
R965 vdd.n1239 vdd.n1238 185
R966 vdd.n968 vdd.n967 185
R967 vdd.n967 vdd.n966 185
R968 vdd.n1233 vdd.n1232 185
R969 vdd.n1232 vdd.n1231 185
R970 vdd.n971 vdd.n970 185
R971 vdd.n972 vdd.n971 185
R972 vdd.n1222 vdd.n1221 185
R973 vdd.n1223 vdd.n1222 185
R974 vdd.n979 vdd.n978 185
R975 vdd.n983 vdd.n978 185
R976 vdd.n1217 vdd.n1216 185
R977 vdd.n1216 vdd.n1215 185
R978 vdd.n784 vdd.n782 185
R979 vdd.n2244 vdd.n782 185
R980 vdd.n2166 vdd.n801 185
R981 vdd.n801 vdd.t119 185
R982 vdd.n2168 vdd.n2167 185
R983 vdd.n2169 vdd.n2168 185
R984 vdd.n2165 vdd.n800 185
R985 vdd.n1868 vdd.n800 185
R986 vdd.n2164 vdd.n2163 185
R987 vdd.n2163 vdd.n2162 185
R988 vdd.n803 vdd.n802 185
R989 vdd.n804 vdd.n803 185
R990 vdd.n2153 vdd.n2152 185
R991 vdd.n2154 vdd.n2153 185
R992 vdd.n2151 vdd.n814 185
R993 vdd.n814 vdd.n811 185
R994 vdd.n2150 vdd.n2149 185
R995 vdd.n2149 vdd.n2148 185
R996 vdd.n816 vdd.n815 185
R997 vdd.n817 vdd.n816 185
R998 vdd.n2141 vdd.n2140 185
R999 vdd.n2142 vdd.n2141 185
R1000 vdd.n2139 vdd.n825 185
R1001 vdd.n830 vdd.n825 185
R1002 vdd.n2138 vdd.n2137 185
R1003 vdd.n2137 vdd.n2136 185
R1004 vdd.n827 vdd.n826 185
R1005 vdd.n836 vdd.n827 185
R1006 vdd.n2129 vdd.n2128 185
R1007 vdd.n2130 vdd.n2129 185
R1008 vdd.n2127 vdd.n837 185
R1009 vdd.n1969 vdd.n837 185
R1010 vdd.n2126 vdd.n2125 185
R1011 vdd.n2125 vdd.n2124 185
R1012 vdd.n839 vdd.n838 185
R1013 vdd.n840 vdd.n839 185
R1014 vdd.n2117 vdd.n2116 185
R1015 vdd.n2118 vdd.n2117 185
R1016 vdd.n2115 vdd.n849 185
R1017 vdd.n849 vdd.n846 185
R1018 vdd.n2114 vdd.n2113 185
R1019 vdd.n2113 vdd.n2112 185
R1020 vdd.n851 vdd.n850 185
R1021 vdd.n861 vdd.n851 185
R1022 vdd.n2104 vdd.n2103 185
R1023 vdd.n2105 vdd.n2104 185
R1024 vdd.n2102 vdd.n862 185
R1025 vdd.n862 vdd.n858 185
R1026 vdd.n2101 vdd.n2100 185
R1027 vdd.n2100 vdd.n2099 185
R1028 vdd.n864 vdd.n863 185
R1029 vdd.n865 vdd.n864 185
R1030 vdd.n2092 vdd.n2091 185
R1031 vdd.n2093 vdd.n2092 185
R1032 vdd.n2090 vdd.n874 185
R1033 vdd.n874 vdd.n871 185
R1034 vdd.n2089 vdd.n2088 185
R1035 vdd.n2088 vdd.n2087 185
R1036 vdd.n876 vdd.n875 185
R1037 vdd.n1824 vdd.n1823 185
R1038 vdd.n1825 vdd.n1821 185
R1039 vdd.n1821 vdd.n877 185
R1040 vdd.n1827 vdd.n1826 185
R1041 vdd.n1829 vdd.n1820 185
R1042 vdd.n1832 vdd.n1831 185
R1043 vdd.n1833 vdd.n1819 185
R1044 vdd.n1835 vdd.n1834 185
R1045 vdd.n1837 vdd.n1818 185
R1046 vdd.n1840 vdd.n1839 185
R1047 vdd.n1841 vdd.n1817 185
R1048 vdd.n1843 vdd.n1842 185
R1049 vdd.n1845 vdd.n1816 185
R1050 vdd.n1848 vdd.n1847 185
R1051 vdd.n1849 vdd.n1815 185
R1052 vdd.n1851 vdd.n1850 185
R1053 vdd.n1853 vdd.n1814 185
R1054 vdd.n2026 vdd.n1854 185
R1055 vdd.n2025 vdd.n2024 185
R1056 vdd.n2022 vdd.n1855 185
R1057 vdd.n2020 vdd.n2019 185
R1058 vdd.n2018 vdd.n1856 185
R1059 vdd.n2017 vdd.n2016 185
R1060 vdd.n2014 vdd.n1857 185
R1061 vdd.n2012 vdd.n2011 185
R1062 vdd.n2010 vdd.n1858 185
R1063 vdd.n2009 vdd.n2008 185
R1064 vdd.n2006 vdd.n1859 185
R1065 vdd.n2004 vdd.n2003 185
R1066 vdd.n2002 vdd.n1860 185
R1067 vdd.n2001 vdd.n2000 185
R1068 vdd.n1998 vdd.n1861 185
R1069 vdd.n1996 vdd.n1995 185
R1070 vdd.n1994 vdd.n1862 185
R1071 vdd.n1993 vdd.n1992 185
R1072 vdd.n2247 vdd.n2246 185
R1073 vdd.n2249 vdd.n2248 185
R1074 vdd.n2251 vdd.n2250 185
R1075 vdd.n2254 vdd.n2253 185
R1076 vdd.n2256 vdd.n2255 185
R1077 vdd.n2258 vdd.n2257 185
R1078 vdd.n2260 vdd.n2259 185
R1079 vdd.n2262 vdd.n2261 185
R1080 vdd.n2264 vdd.n2263 185
R1081 vdd.n2266 vdd.n2265 185
R1082 vdd.n2268 vdd.n2267 185
R1083 vdd.n2270 vdd.n2269 185
R1084 vdd.n2272 vdd.n2271 185
R1085 vdd.n2274 vdd.n2273 185
R1086 vdd.n2276 vdd.n2275 185
R1087 vdd.n2278 vdd.n2277 185
R1088 vdd.n2280 vdd.n2279 185
R1089 vdd.n2282 vdd.n2281 185
R1090 vdd.n2284 vdd.n2283 185
R1091 vdd.n2286 vdd.n2285 185
R1092 vdd.n2288 vdd.n2287 185
R1093 vdd.n2290 vdd.n2289 185
R1094 vdd.n2292 vdd.n2291 185
R1095 vdd.n2294 vdd.n2293 185
R1096 vdd.n2296 vdd.n2295 185
R1097 vdd.n2298 vdd.n2297 185
R1098 vdd.n2300 vdd.n2299 185
R1099 vdd.n2302 vdd.n2301 185
R1100 vdd.n2304 vdd.n2303 185
R1101 vdd.n2306 vdd.n2305 185
R1102 vdd.n2308 vdd.n2307 185
R1103 vdd.n2310 vdd.n2309 185
R1104 vdd.n2312 vdd.n2311 185
R1105 vdd.n2313 vdd.n783 185
R1106 vdd.n2315 vdd.n2314 185
R1107 vdd.n2316 vdd.n2315 185
R1108 vdd.n2245 vdd.n787 185
R1109 vdd.n2245 vdd.n2244 185
R1110 vdd.n1866 vdd.n788 185
R1111 vdd.t119 vdd.n788 185
R1112 vdd.n1867 vdd.n798 185
R1113 vdd.n2169 vdd.n798 185
R1114 vdd.n1870 vdd.n1869 185
R1115 vdd.n1869 vdd.n1868 185
R1116 vdd.n1871 vdd.n805 185
R1117 vdd.n2162 vdd.n805 185
R1118 vdd.n1873 vdd.n1872 185
R1119 vdd.n1872 vdd.n804 185
R1120 vdd.n1874 vdd.n812 185
R1121 vdd.n2154 vdd.n812 185
R1122 vdd.n1876 vdd.n1875 185
R1123 vdd.n1875 vdd.n811 185
R1124 vdd.n1877 vdd.n818 185
R1125 vdd.n2148 vdd.n818 185
R1126 vdd.n1879 vdd.n1878 185
R1127 vdd.n1878 vdd.n817 185
R1128 vdd.n1880 vdd.n823 185
R1129 vdd.n2142 vdd.n823 185
R1130 vdd.n1882 vdd.n1881 185
R1131 vdd.n1881 vdd.n830 185
R1132 vdd.n1883 vdd.n828 185
R1133 vdd.n2136 vdd.n828 185
R1134 vdd.n1885 vdd.n1884 185
R1135 vdd.n1884 vdd.n836 185
R1136 vdd.n1886 vdd.n834 185
R1137 vdd.n2130 vdd.n834 185
R1138 vdd.n1971 vdd.n1970 185
R1139 vdd.n1970 vdd.n1969 185
R1140 vdd.n1972 vdd.n841 185
R1141 vdd.n2124 vdd.n841 185
R1142 vdd.n1974 vdd.n1973 185
R1143 vdd.n1973 vdd.n840 185
R1144 vdd.n1975 vdd.n847 185
R1145 vdd.n2118 vdd.n847 185
R1146 vdd.n1977 vdd.n1976 185
R1147 vdd.n1976 vdd.n846 185
R1148 vdd.n1978 vdd.n852 185
R1149 vdd.n2112 vdd.n852 185
R1150 vdd.n1980 vdd.n1979 185
R1151 vdd.n1979 vdd.n861 185
R1152 vdd.n1981 vdd.n859 185
R1153 vdd.n2105 vdd.n859 185
R1154 vdd.n1983 vdd.n1982 185
R1155 vdd.n1982 vdd.n858 185
R1156 vdd.n1984 vdd.n866 185
R1157 vdd.n2099 vdd.n866 185
R1158 vdd.n1986 vdd.n1985 185
R1159 vdd.n1985 vdd.n865 185
R1160 vdd.n1987 vdd.n872 185
R1161 vdd.n2093 vdd.n872 185
R1162 vdd.n1989 vdd.n1988 185
R1163 vdd.n1988 vdd.n871 185
R1164 vdd.n1990 vdd.n878 185
R1165 vdd.n2087 vdd.n878 185
R1166 vdd.n3137 vdd.n3136 185
R1167 vdd.n3138 vdd.n3137 185
R1168 vdd.n347 vdd.n346 185
R1169 vdd.n3139 vdd.n347 185
R1170 vdd.n3142 vdd.n3141 185
R1171 vdd.n3141 vdd.n3140 185
R1172 vdd.n3143 vdd.n341 185
R1173 vdd.n341 vdd.n340 185
R1174 vdd.n3145 vdd.n3144 185
R1175 vdd.n3146 vdd.n3145 185
R1176 vdd.n336 vdd.n335 185
R1177 vdd.n3147 vdd.n336 185
R1178 vdd.n3150 vdd.n3149 185
R1179 vdd.n3149 vdd.n3148 185
R1180 vdd.n3151 vdd.n330 185
R1181 vdd.n330 vdd.n329 185
R1182 vdd.n3153 vdd.n3152 185
R1183 vdd.n3154 vdd.n3153 185
R1184 vdd.n324 vdd.n323 185
R1185 vdd.n3155 vdd.n324 185
R1186 vdd.n3158 vdd.n3157 185
R1187 vdd.n3157 vdd.n3156 185
R1188 vdd.n3159 vdd.n319 185
R1189 vdd.n325 vdd.n319 185
R1190 vdd.n3161 vdd.n3160 185
R1191 vdd.n3162 vdd.n3161 185
R1192 vdd.n315 vdd.n313 185
R1193 vdd.n3163 vdd.n315 185
R1194 vdd.n3166 vdd.n3165 185
R1195 vdd.n3165 vdd.n3164 185
R1196 vdd.n314 vdd.n312 185
R1197 vdd.n481 vdd.n314 185
R1198 vdd.n2988 vdd.n2987 185
R1199 vdd.n2989 vdd.n2988 185
R1200 vdd.n483 vdd.n482 185
R1201 vdd.n2980 vdd.n482 185
R1202 vdd.n2983 vdd.n2982 185
R1203 vdd.n2982 vdd.n2981 185
R1204 vdd.n486 vdd.n485 185
R1205 vdd.n493 vdd.n486 185
R1206 vdd.n2971 vdd.n2970 185
R1207 vdd.n2972 vdd.n2971 185
R1208 vdd.n495 vdd.n494 185
R1209 vdd.n494 vdd.n492 185
R1210 vdd.n2966 vdd.n2965 185
R1211 vdd.n2965 vdd.n2964 185
R1212 vdd.n498 vdd.n497 185
R1213 vdd.n499 vdd.n498 185
R1214 vdd.n2955 vdd.n2954 185
R1215 vdd.n2956 vdd.n2955 185
R1216 vdd.n507 vdd.n506 185
R1217 vdd.n506 vdd.n505 185
R1218 vdd.n2950 vdd.n2949 185
R1219 vdd.n2949 vdd.n2948 185
R1220 vdd.n510 vdd.n509 185
R1221 vdd.n511 vdd.n510 185
R1222 vdd.n2939 vdd.n2938 185
R1223 vdd.n2940 vdd.n2939 185
R1224 vdd.n2935 vdd.n517 185
R1225 vdd.n2934 vdd.n2933 185
R1226 vdd.n2931 vdd.n519 185
R1227 vdd.n2931 vdd.n516 185
R1228 vdd.n2930 vdd.n2929 185
R1229 vdd.n2928 vdd.n2927 185
R1230 vdd.n2926 vdd.n2925 185
R1231 vdd.n2924 vdd.n2923 185
R1232 vdd.n2922 vdd.n525 185
R1233 vdd.n2920 vdd.n2919 185
R1234 vdd.n2918 vdd.n526 185
R1235 vdd.n2917 vdd.n2916 185
R1236 vdd.n2914 vdd.n531 185
R1237 vdd.n2912 vdd.n2911 185
R1238 vdd.n2910 vdd.n532 185
R1239 vdd.n2909 vdd.n2908 185
R1240 vdd.n2906 vdd.n537 185
R1241 vdd.n2904 vdd.n2903 185
R1242 vdd.n2902 vdd.n538 185
R1243 vdd.n2901 vdd.n2900 185
R1244 vdd.n2898 vdd.n545 185
R1245 vdd.n2896 vdd.n2895 185
R1246 vdd.n2894 vdd.n546 185
R1247 vdd.n2893 vdd.n2892 185
R1248 vdd.n2890 vdd.n551 185
R1249 vdd.n2888 vdd.n2887 185
R1250 vdd.n2886 vdd.n552 185
R1251 vdd.n2885 vdd.n2884 185
R1252 vdd.n2882 vdd.n557 185
R1253 vdd.n2880 vdd.n2879 185
R1254 vdd.n2878 vdd.n558 185
R1255 vdd.n2877 vdd.n2876 185
R1256 vdd.n2874 vdd.n563 185
R1257 vdd.n2872 vdd.n2871 185
R1258 vdd.n2870 vdd.n564 185
R1259 vdd.n2869 vdd.n2868 185
R1260 vdd.n2866 vdd.n569 185
R1261 vdd.n2864 vdd.n2863 185
R1262 vdd.n2862 vdd.n570 185
R1263 vdd.n2861 vdd.n2860 185
R1264 vdd.n2858 vdd.n575 185
R1265 vdd.n2856 vdd.n2855 185
R1266 vdd.n2854 vdd.n576 185
R1267 vdd.n585 vdd.n579 185
R1268 vdd.n2850 vdd.n2849 185
R1269 vdd.n2847 vdd.n583 185
R1270 vdd.n2846 vdd.n2845 185
R1271 vdd.n2844 vdd.n2843 185
R1272 vdd.n2842 vdd.n589 185
R1273 vdd.n2840 vdd.n2839 185
R1274 vdd.n2838 vdd.n590 185
R1275 vdd.n2837 vdd.n2836 185
R1276 vdd.n2834 vdd.n595 185
R1277 vdd.n2832 vdd.n2831 185
R1278 vdd.n2830 vdd.n596 185
R1279 vdd.n2829 vdd.n2828 185
R1280 vdd.n2826 vdd.n601 185
R1281 vdd.n2824 vdd.n2823 185
R1282 vdd.n2822 vdd.n602 185
R1283 vdd.n2821 vdd.n2820 185
R1284 vdd.n2818 vdd.n2817 185
R1285 vdd.n2816 vdd.n2815 185
R1286 vdd.n2814 vdd.n2813 185
R1287 vdd.n2812 vdd.n2811 185
R1288 vdd.n2807 vdd.n515 185
R1289 vdd.n516 vdd.n515 185
R1290 vdd.n3020 vdd.n3019 185
R1291 vdd.n3024 vdd.n462 185
R1292 vdd.n3026 vdd.n3025 185
R1293 vdd.n3028 vdd.n460 185
R1294 vdd.n3030 vdd.n3029 185
R1295 vdd.n3031 vdd.n455 185
R1296 vdd.n3033 vdd.n3032 185
R1297 vdd.n3035 vdd.n453 185
R1298 vdd.n3037 vdd.n3036 185
R1299 vdd.n3038 vdd.n448 185
R1300 vdd.n3040 vdd.n3039 185
R1301 vdd.n3042 vdd.n446 185
R1302 vdd.n3044 vdd.n3043 185
R1303 vdd.n3045 vdd.n441 185
R1304 vdd.n3047 vdd.n3046 185
R1305 vdd.n3049 vdd.n439 185
R1306 vdd.n3051 vdd.n3050 185
R1307 vdd.n3052 vdd.n435 185
R1308 vdd.n3054 vdd.n3053 185
R1309 vdd.n3056 vdd.n432 185
R1310 vdd.n3058 vdd.n3057 185
R1311 vdd.n433 vdd.n426 185
R1312 vdd.n3062 vdd.n430 185
R1313 vdd.n3063 vdd.n422 185
R1314 vdd.n3065 vdd.n3064 185
R1315 vdd.n3067 vdd.n420 185
R1316 vdd.n3069 vdd.n3068 185
R1317 vdd.n3070 vdd.n415 185
R1318 vdd.n3072 vdd.n3071 185
R1319 vdd.n3074 vdd.n413 185
R1320 vdd.n3076 vdd.n3075 185
R1321 vdd.n3077 vdd.n408 185
R1322 vdd.n3079 vdd.n3078 185
R1323 vdd.n3081 vdd.n406 185
R1324 vdd.n3083 vdd.n3082 185
R1325 vdd.n3084 vdd.n401 185
R1326 vdd.n3086 vdd.n3085 185
R1327 vdd.n3088 vdd.n399 185
R1328 vdd.n3090 vdd.n3089 185
R1329 vdd.n3091 vdd.n395 185
R1330 vdd.n3093 vdd.n3092 185
R1331 vdd.n3095 vdd.n392 185
R1332 vdd.n3097 vdd.n3096 185
R1333 vdd.n393 vdd.n386 185
R1334 vdd.n3101 vdd.n390 185
R1335 vdd.n3102 vdd.n382 185
R1336 vdd.n3104 vdd.n3103 185
R1337 vdd.n3106 vdd.n380 185
R1338 vdd.n3108 vdd.n3107 185
R1339 vdd.n3109 vdd.n375 185
R1340 vdd.n3111 vdd.n3110 185
R1341 vdd.n3113 vdd.n373 185
R1342 vdd.n3115 vdd.n3114 185
R1343 vdd.n3116 vdd.n368 185
R1344 vdd.n3118 vdd.n3117 185
R1345 vdd.n3120 vdd.n366 185
R1346 vdd.n3122 vdd.n3121 185
R1347 vdd.n3123 vdd.n360 185
R1348 vdd.n3125 vdd.n3124 185
R1349 vdd.n3127 vdd.n359 185
R1350 vdd.n3128 vdd.n358 185
R1351 vdd.n3131 vdd.n3130 185
R1352 vdd.n3132 vdd.n356 185
R1353 vdd.n3133 vdd.n352 185
R1354 vdd.n3015 vdd.n350 185
R1355 vdd.n3138 vdd.n350 185
R1356 vdd.n3014 vdd.n349 185
R1357 vdd.n3139 vdd.n349 185
R1358 vdd.n3013 vdd.n348 185
R1359 vdd.n3140 vdd.n348 185
R1360 vdd.n468 vdd.n467 185
R1361 vdd.n467 vdd.n340 185
R1362 vdd.n3009 vdd.n339 185
R1363 vdd.n3146 vdd.n339 185
R1364 vdd.n3008 vdd.n338 185
R1365 vdd.n3147 vdd.n338 185
R1366 vdd.n3007 vdd.n337 185
R1367 vdd.n3148 vdd.n337 185
R1368 vdd.n471 vdd.n470 185
R1369 vdd.n470 vdd.n329 185
R1370 vdd.n3003 vdd.n328 185
R1371 vdd.n3154 vdd.n328 185
R1372 vdd.n3002 vdd.n327 185
R1373 vdd.n3155 vdd.n327 185
R1374 vdd.n3001 vdd.n326 185
R1375 vdd.n3156 vdd.n326 185
R1376 vdd.n474 vdd.n473 185
R1377 vdd.n473 vdd.n325 185
R1378 vdd.n2997 vdd.n318 185
R1379 vdd.n3162 vdd.n318 185
R1380 vdd.n2996 vdd.n317 185
R1381 vdd.n3163 vdd.n317 185
R1382 vdd.n2995 vdd.n316 185
R1383 vdd.n3164 vdd.n316 185
R1384 vdd.n480 vdd.n476 185
R1385 vdd.n481 vdd.n480 185
R1386 vdd.n2991 vdd.n2990 185
R1387 vdd.n2990 vdd.n2989 185
R1388 vdd.n479 vdd.n478 185
R1389 vdd.n2980 vdd.n479 185
R1390 vdd.n2979 vdd.n2978 185
R1391 vdd.n2981 vdd.n2979 185
R1392 vdd.n488 vdd.n487 185
R1393 vdd.n493 vdd.n487 185
R1394 vdd.n2974 vdd.n2973 185
R1395 vdd.n2973 vdd.n2972 185
R1396 vdd.n491 vdd.n490 185
R1397 vdd.n492 vdd.n491 185
R1398 vdd.n2963 vdd.n2962 185
R1399 vdd.n2964 vdd.n2963 185
R1400 vdd.n501 vdd.n500 185
R1401 vdd.n500 vdd.n499 185
R1402 vdd.n2958 vdd.n2957 185
R1403 vdd.n2957 vdd.n2956 185
R1404 vdd.n504 vdd.n503 185
R1405 vdd.n505 vdd.n504 185
R1406 vdd.n2947 vdd.n2946 185
R1407 vdd.n2948 vdd.n2947 185
R1408 vdd.n513 vdd.n512 185
R1409 vdd.n512 vdd.n511 185
R1410 vdd.n2942 vdd.n2941 185
R1411 vdd.n2941 vdd.n2940 185
R1412 vdd.n741 vdd.n740 185
R1413 vdd.n2567 vdd.n2566 185
R1414 vdd.n2565 vdd.n2350 185
R1415 vdd.n2569 vdd.n2350 185
R1416 vdd.n2564 vdd.n2563 185
R1417 vdd.n2562 vdd.n2561 185
R1418 vdd.n2560 vdd.n2559 185
R1419 vdd.n2558 vdd.n2557 185
R1420 vdd.n2556 vdd.n2555 185
R1421 vdd.n2554 vdd.n2553 185
R1422 vdd.n2552 vdd.n2551 185
R1423 vdd.n2550 vdd.n2549 185
R1424 vdd.n2548 vdd.n2547 185
R1425 vdd.n2546 vdd.n2545 185
R1426 vdd.n2544 vdd.n2543 185
R1427 vdd.n2542 vdd.n2541 185
R1428 vdd.n2540 vdd.n2539 185
R1429 vdd.n2538 vdd.n2537 185
R1430 vdd.n2536 vdd.n2535 185
R1431 vdd.n2534 vdd.n2533 185
R1432 vdd.n2532 vdd.n2531 185
R1433 vdd.n2530 vdd.n2529 185
R1434 vdd.n2528 vdd.n2527 185
R1435 vdd.n2526 vdd.n2525 185
R1436 vdd.n2524 vdd.n2523 185
R1437 vdd.n2522 vdd.n2521 185
R1438 vdd.n2520 vdd.n2519 185
R1439 vdd.n2518 vdd.n2517 185
R1440 vdd.n2516 vdd.n2515 185
R1441 vdd.n2514 vdd.n2513 185
R1442 vdd.n2512 vdd.n2511 185
R1443 vdd.n2510 vdd.n2509 185
R1444 vdd.n2508 vdd.n2507 185
R1445 vdd.n2505 vdd.n2504 185
R1446 vdd.n2503 vdd.n2502 185
R1447 vdd.n2501 vdd.n2500 185
R1448 vdd.n2708 vdd.n2707 185
R1449 vdd.n2709 vdd.n660 185
R1450 vdd.n2711 vdd.n2710 185
R1451 vdd.n2713 vdd.n658 185
R1452 vdd.n2715 vdd.n2714 185
R1453 vdd.n2716 vdd.n657 185
R1454 vdd.n2718 vdd.n2717 185
R1455 vdd.n2720 vdd.n655 185
R1456 vdd.n2722 vdd.n2721 185
R1457 vdd.n2723 vdd.n654 185
R1458 vdd.n2725 vdd.n2724 185
R1459 vdd.n2727 vdd.n652 185
R1460 vdd.n2729 vdd.n2728 185
R1461 vdd.n2730 vdd.n651 185
R1462 vdd.n2732 vdd.n2731 185
R1463 vdd.n2734 vdd.n649 185
R1464 vdd.n2736 vdd.n2735 185
R1465 vdd.n2738 vdd.n648 185
R1466 vdd.n2740 vdd.n2739 185
R1467 vdd.n2742 vdd.n646 185
R1468 vdd.n2744 vdd.n2743 185
R1469 vdd.n2745 vdd.n645 185
R1470 vdd.n2747 vdd.n2746 185
R1471 vdd.n2749 vdd.n643 185
R1472 vdd.n2751 vdd.n2750 185
R1473 vdd.n2752 vdd.n642 185
R1474 vdd.n2754 vdd.n2753 185
R1475 vdd.n2756 vdd.n640 185
R1476 vdd.n2758 vdd.n2757 185
R1477 vdd.n2759 vdd.n639 185
R1478 vdd.n2761 vdd.n2760 185
R1479 vdd.n2763 vdd.n638 185
R1480 vdd.n2764 vdd.n637 185
R1481 vdd.n2767 vdd.n2766 185
R1482 vdd.n2768 vdd.n635 185
R1483 vdd.n635 vdd.n613 185
R1484 vdd.n2705 vdd.n632 185
R1485 vdd.n2771 vdd.n632 185
R1486 vdd.n2704 vdd.n2703 185
R1487 vdd.n2703 vdd.n631 185
R1488 vdd.n2702 vdd.n664 185
R1489 vdd.n2702 vdd.n2701 185
R1490 vdd.n2456 vdd.n665 185
R1491 vdd.n674 vdd.n665 185
R1492 vdd.n2457 vdd.n672 185
R1493 vdd.n2695 vdd.n672 185
R1494 vdd.n2459 vdd.n2458 185
R1495 vdd.n2458 vdd.n671 185
R1496 vdd.n2460 vdd.n680 185
R1497 vdd.n2644 vdd.n680 185
R1498 vdd.n2462 vdd.n2461 185
R1499 vdd.n2461 vdd.n679 185
R1500 vdd.n2463 vdd.n686 185
R1501 vdd.n2638 vdd.n686 185
R1502 vdd.n2465 vdd.n2464 185
R1503 vdd.n2464 vdd.n685 185
R1504 vdd.n2466 vdd.n691 185
R1505 vdd.n2630 vdd.n691 185
R1506 vdd.n2468 vdd.n2467 185
R1507 vdd.n2467 vdd.n698 185
R1508 vdd.n2469 vdd.n696 185
R1509 vdd.n2624 vdd.n696 185
R1510 vdd.n2471 vdd.n2470 185
R1511 vdd.n2472 vdd.n2471 185
R1512 vdd.n2455 vdd.n703 185
R1513 vdd.n2618 vdd.n703 185
R1514 vdd.n2454 vdd.n2453 185
R1515 vdd.n2453 vdd.n702 185
R1516 vdd.n2452 vdd.n709 185
R1517 vdd.n2612 vdd.n709 185
R1518 vdd.n2451 vdd.n2450 185
R1519 vdd.n2450 vdd.n708 185
R1520 vdd.n2449 vdd.n714 185
R1521 vdd.n2606 vdd.n714 185
R1522 vdd.n2448 vdd.n2447 185
R1523 vdd.n2447 vdd.n721 185
R1524 vdd.n2446 vdd.n719 185
R1525 vdd.n2600 vdd.n719 185
R1526 vdd.n2445 vdd.n2444 185
R1527 vdd.n2444 vdd.n728 185
R1528 vdd.n2443 vdd.n726 185
R1529 vdd.n2594 vdd.n726 185
R1530 vdd.n2442 vdd.n2441 185
R1531 vdd.n2441 vdd.n725 185
R1532 vdd.n2353 vdd.n732 185
R1533 vdd.n2588 vdd.n732 185
R1534 vdd.n2495 vdd.n2494 185
R1535 vdd.n2494 vdd.n2493 185
R1536 vdd.n2496 vdd.n737 185
R1537 vdd.n2582 vdd.n737 185
R1538 vdd.n2498 vdd.n2497 185
R1539 vdd.n2497 vdd.t87 185
R1540 vdd.n2499 vdd.n742 185
R1541 vdd.n2576 vdd.n742 185
R1542 vdd.n2578 vdd.n2577 185
R1543 vdd.n2577 vdd.n2576 185
R1544 vdd.n2579 vdd.n739 185
R1545 vdd.n739 vdd.t87 185
R1546 vdd.n2581 vdd.n2580 185
R1547 vdd.n2582 vdd.n2581 185
R1548 vdd.n731 vdd.n730 185
R1549 vdd.n2493 vdd.n731 185
R1550 vdd.n2590 vdd.n2589 185
R1551 vdd.n2589 vdd.n2588 185
R1552 vdd.n2591 vdd.n729 185
R1553 vdd.n729 vdd.n725 185
R1554 vdd.n2593 vdd.n2592 185
R1555 vdd.n2594 vdd.n2593 185
R1556 vdd.n718 vdd.n717 185
R1557 vdd.n728 vdd.n718 185
R1558 vdd.n2602 vdd.n2601 185
R1559 vdd.n2601 vdd.n2600 185
R1560 vdd.n2603 vdd.n716 185
R1561 vdd.n721 vdd.n716 185
R1562 vdd.n2605 vdd.n2604 185
R1563 vdd.n2606 vdd.n2605 185
R1564 vdd.n707 vdd.n706 185
R1565 vdd.n708 vdd.n707 185
R1566 vdd.n2614 vdd.n2613 185
R1567 vdd.n2613 vdd.n2612 185
R1568 vdd.n2615 vdd.n705 185
R1569 vdd.n705 vdd.n702 185
R1570 vdd.n2617 vdd.n2616 185
R1571 vdd.n2618 vdd.n2617 185
R1572 vdd.n695 vdd.n694 185
R1573 vdd.n2472 vdd.n695 185
R1574 vdd.n2626 vdd.n2625 185
R1575 vdd.n2625 vdd.n2624 185
R1576 vdd.n2627 vdd.n693 185
R1577 vdd.n698 vdd.n693 185
R1578 vdd.n2629 vdd.n2628 185
R1579 vdd.n2630 vdd.n2629 185
R1580 vdd.n684 vdd.n683 185
R1581 vdd.n685 vdd.n684 185
R1582 vdd.n2640 vdd.n2639 185
R1583 vdd.n2639 vdd.n2638 185
R1584 vdd.n2641 vdd.n682 185
R1585 vdd.n682 vdd.n679 185
R1586 vdd.n2643 vdd.n2642 185
R1587 vdd.n2644 vdd.n2643 185
R1588 vdd.n670 vdd.n669 185
R1589 vdd.n671 vdd.n670 185
R1590 vdd.n2697 vdd.n2696 185
R1591 vdd.n2696 vdd.n2695 185
R1592 vdd.n2698 vdd.n668 185
R1593 vdd.n674 vdd.n668 185
R1594 vdd.n2700 vdd.n2699 185
R1595 vdd.n2701 vdd.n2700 185
R1596 vdd.n636 vdd.n634 185
R1597 vdd.n634 vdd.n631 185
R1598 vdd.n2770 vdd.n2769 185
R1599 vdd.n2771 vdd.n2770 185
R1600 vdd.n2243 vdd.n2242 185
R1601 vdd.n2244 vdd.n2243 185
R1602 vdd.n792 vdd.n790 185
R1603 vdd.n790 vdd.t119 185
R1604 vdd.n2158 vdd.n799 185
R1605 vdd.n2169 vdd.n799 185
R1606 vdd.n2159 vdd.n808 185
R1607 vdd.n1868 vdd.n808 185
R1608 vdd.n2161 vdd.n2160 185
R1609 vdd.n2162 vdd.n2161 185
R1610 vdd.n2157 vdd.n807 185
R1611 vdd.n807 vdd.n804 185
R1612 vdd.n2156 vdd.n2155 185
R1613 vdd.n2155 vdd.n2154 185
R1614 vdd.n810 vdd.n809 185
R1615 vdd.n811 vdd.n810 185
R1616 vdd.n2147 vdd.n2146 185
R1617 vdd.n2148 vdd.n2147 185
R1618 vdd.n2145 vdd.n820 185
R1619 vdd.n820 vdd.n817 185
R1620 vdd.n2144 vdd.n2143 185
R1621 vdd.n2143 vdd.n2142 185
R1622 vdd.n822 vdd.n821 185
R1623 vdd.n830 vdd.n822 185
R1624 vdd.n2135 vdd.n2134 185
R1625 vdd.n2136 vdd.n2135 185
R1626 vdd.n2133 vdd.n831 185
R1627 vdd.n836 vdd.n831 185
R1628 vdd.n2132 vdd.n2131 185
R1629 vdd.n2131 vdd.n2130 185
R1630 vdd.n833 vdd.n832 185
R1631 vdd.n1969 vdd.n833 185
R1632 vdd.n2123 vdd.n2122 185
R1633 vdd.n2124 vdd.n2123 185
R1634 vdd.n2121 vdd.n843 185
R1635 vdd.n843 vdd.n840 185
R1636 vdd.n2120 vdd.n2119 185
R1637 vdd.n2119 vdd.n2118 185
R1638 vdd.n845 vdd.n844 185
R1639 vdd.n846 vdd.n845 185
R1640 vdd.n2111 vdd.n2110 185
R1641 vdd.n2112 vdd.n2111 185
R1642 vdd.n2108 vdd.n854 185
R1643 vdd.n861 vdd.n854 185
R1644 vdd.n2107 vdd.n2106 185
R1645 vdd.n2106 vdd.n2105 185
R1646 vdd.n857 vdd.n856 185
R1647 vdd.n858 vdd.n857 185
R1648 vdd.n2098 vdd.n2097 185
R1649 vdd.n2099 vdd.n2098 185
R1650 vdd.n2096 vdd.n868 185
R1651 vdd.n868 vdd.n865 185
R1652 vdd.n2095 vdd.n2094 185
R1653 vdd.n2094 vdd.n2093 185
R1654 vdd.n870 vdd.n869 185
R1655 vdd.n871 vdd.n870 185
R1656 vdd.n2086 vdd.n2085 185
R1657 vdd.n2087 vdd.n2086 185
R1658 vdd.n2174 vdd.n764 185
R1659 vdd.n2316 vdd.n764 185
R1660 vdd.n2176 vdd.n2175 185
R1661 vdd.n2178 vdd.n2177 185
R1662 vdd.n2180 vdd.n2179 185
R1663 vdd.n2182 vdd.n2181 185
R1664 vdd.n2184 vdd.n2183 185
R1665 vdd.n2186 vdd.n2185 185
R1666 vdd.n2188 vdd.n2187 185
R1667 vdd.n2190 vdd.n2189 185
R1668 vdd.n2192 vdd.n2191 185
R1669 vdd.n2194 vdd.n2193 185
R1670 vdd.n2196 vdd.n2195 185
R1671 vdd.n2198 vdd.n2197 185
R1672 vdd.n2200 vdd.n2199 185
R1673 vdd.n2202 vdd.n2201 185
R1674 vdd.n2204 vdd.n2203 185
R1675 vdd.n2206 vdd.n2205 185
R1676 vdd.n2208 vdd.n2207 185
R1677 vdd.n2210 vdd.n2209 185
R1678 vdd.n2212 vdd.n2211 185
R1679 vdd.n2214 vdd.n2213 185
R1680 vdd.n2216 vdd.n2215 185
R1681 vdd.n2218 vdd.n2217 185
R1682 vdd.n2220 vdd.n2219 185
R1683 vdd.n2222 vdd.n2221 185
R1684 vdd.n2224 vdd.n2223 185
R1685 vdd.n2226 vdd.n2225 185
R1686 vdd.n2228 vdd.n2227 185
R1687 vdd.n2230 vdd.n2229 185
R1688 vdd.n2232 vdd.n2231 185
R1689 vdd.n2234 vdd.n2233 185
R1690 vdd.n2236 vdd.n2235 185
R1691 vdd.n2238 vdd.n2237 185
R1692 vdd.n2240 vdd.n2239 185
R1693 vdd.n2241 vdd.n791 185
R1694 vdd.n2173 vdd.n789 185
R1695 vdd.n2244 vdd.n789 185
R1696 vdd.n2172 vdd.n2171 185
R1697 vdd.n2171 vdd.t119 185
R1698 vdd.n2170 vdd.n796 185
R1699 vdd.n2170 vdd.n2169 185
R1700 vdd.n1950 vdd.n797 185
R1701 vdd.n1868 vdd.n797 185
R1702 vdd.n1951 vdd.n806 185
R1703 vdd.n2162 vdd.n806 185
R1704 vdd.n1953 vdd.n1952 185
R1705 vdd.n1952 vdd.n804 185
R1706 vdd.n1954 vdd.n813 185
R1707 vdd.n2154 vdd.n813 185
R1708 vdd.n1956 vdd.n1955 185
R1709 vdd.n1955 vdd.n811 185
R1710 vdd.n1957 vdd.n819 185
R1711 vdd.n2148 vdd.n819 185
R1712 vdd.n1959 vdd.n1958 185
R1713 vdd.n1958 vdd.n817 185
R1714 vdd.n1960 vdd.n824 185
R1715 vdd.n2142 vdd.n824 185
R1716 vdd.n1962 vdd.n1961 185
R1717 vdd.n1961 vdd.n830 185
R1718 vdd.n1963 vdd.n829 185
R1719 vdd.n2136 vdd.n829 185
R1720 vdd.n1965 vdd.n1964 185
R1721 vdd.n1964 vdd.n836 185
R1722 vdd.n1966 vdd.n835 185
R1723 vdd.n2130 vdd.n835 185
R1724 vdd.n1968 vdd.n1967 185
R1725 vdd.n1969 vdd.n1968 185
R1726 vdd.n1949 vdd.n842 185
R1727 vdd.n2124 vdd.n842 185
R1728 vdd.n1948 vdd.n1947 185
R1729 vdd.n1947 vdd.n840 185
R1730 vdd.n1946 vdd.n848 185
R1731 vdd.n2118 vdd.n848 185
R1732 vdd.n1945 vdd.n1944 185
R1733 vdd.n1944 vdd.n846 185
R1734 vdd.n1943 vdd.n853 185
R1735 vdd.n2112 vdd.n853 185
R1736 vdd.n1942 vdd.n1941 185
R1737 vdd.n1941 vdd.n861 185
R1738 vdd.n1940 vdd.n860 185
R1739 vdd.n2105 vdd.n860 185
R1740 vdd.n1939 vdd.n1938 185
R1741 vdd.n1938 vdd.n858 185
R1742 vdd.n1937 vdd.n867 185
R1743 vdd.n2099 vdd.n867 185
R1744 vdd.n1936 vdd.n1935 185
R1745 vdd.n1935 vdd.n865 185
R1746 vdd.n1934 vdd.n873 185
R1747 vdd.n2093 vdd.n873 185
R1748 vdd.n1933 vdd.n1932 185
R1749 vdd.n1932 vdd.n871 185
R1750 vdd.n1931 vdd.n879 185
R1751 vdd.n2087 vdd.n879 185
R1752 vdd.n2084 vdd.n880 185
R1753 vdd.n2083 vdd.n2082 185
R1754 vdd.n2080 vdd.n881 185
R1755 vdd.n2078 vdd.n2077 185
R1756 vdd.n2076 vdd.n882 185
R1757 vdd.n2075 vdd.n2074 185
R1758 vdd.n2072 vdd.n883 185
R1759 vdd.n2070 vdd.n2069 185
R1760 vdd.n2068 vdd.n884 185
R1761 vdd.n2067 vdd.n2066 185
R1762 vdd.n2064 vdd.n885 185
R1763 vdd.n2062 vdd.n2061 185
R1764 vdd.n2060 vdd.n886 185
R1765 vdd.n2059 vdd.n2058 185
R1766 vdd.n2056 vdd.n887 185
R1767 vdd.n2054 vdd.n2053 185
R1768 vdd.n2052 vdd.n888 185
R1769 vdd.n2051 vdd.n890 185
R1770 vdd.n1896 vdd.n891 185
R1771 vdd.n1899 vdd.n1898 185
R1772 vdd.n1901 vdd.n1900 185
R1773 vdd.n1903 vdd.n1895 185
R1774 vdd.n1906 vdd.n1905 185
R1775 vdd.n1907 vdd.n1894 185
R1776 vdd.n1909 vdd.n1908 185
R1777 vdd.n1911 vdd.n1893 185
R1778 vdd.n1914 vdd.n1913 185
R1779 vdd.n1915 vdd.n1892 185
R1780 vdd.n1917 vdd.n1916 185
R1781 vdd.n1919 vdd.n1891 185
R1782 vdd.n1922 vdd.n1921 185
R1783 vdd.n1923 vdd.n1888 185
R1784 vdd.n1926 vdd.n1925 185
R1785 vdd.n1928 vdd.n1887 185
R1786 vdd.n1930 vdd.n1929 185
R1787 vdd.n1929 vdd.n877 185
R1788 vdd.n303 vdd.n302 171.744
R1789 vdd.n302 vdd.n301 171.744
R1790 vdd.n301 vdd.n270 171.744
R1791 vdd.n294 vdd.n270 171.744
R1792 vdd.n294 vdd.n293 171.744
R1793 vdd.n293 vdd.n275 171.744
R1794 vdd.n286 vdd.n275 171.744
R1795 vdd.n286 vdd.n285 171.744
R1796 vdd.n285 vdd.n279 171.744
R1797 vdd.n252 vdd.n251 171.744
R1798 vdd.n251 vdd.n250 171.744
R1799 vdd.n250 vdd.n219 171.744
R1800 vdd.n243 vdd.n219 171.744
R1801 vdd.n243 vdd.n242 171.744
R1802 vdd.n242 vdd.n224 171.744
R1803 vdd.n235 vdd.n224 171.744
R1804 vdd.n235 vdd.n234 171.744
R1805 vdd.n234 vdd.n228 171.744
R1806 vdd.n209 vdd.n208 171.744
R1807 vdd.n208 vdd.n207 171.744
R1808 vdd.n207 vdd.n176 171.744
R1809 vdd.n200 vdd.n176 171.744
R1810 vdd.n200 vdd.n199 171.744
R1811 vdd.n199 vdd.n181 171.744
R1812 vdd.n192 vdd.n181 171.744
R1813 vdd.n192 vdd.n191 171.744
R1814 vdd.n191 vdd.n185 171.744
R1815 vdd.n158 vdd.n157 171.744
R1816 vdd.n157 vdd.n156 171.744
R1817 vdd.n156 vdd.n125 171.744
R1818 vdd.n149 vdd.n125 171.744
R1819 vdd.n149 vdd.n148 171.744
R1820 vdd.n148 vdd.n130 171.744
R1821 vdd.n141 vdd.n130 171.744
R1822 vdd.n141 vdd.n140 171.744
R1823 vdd.n140 vdd.n134 171.744
R1824 vdd.n116 vdd.n115 171.744
R1825 vdd.n115 vdd.n114 171.744
R1826 vdd.n114 vdd.n83 171.744
R1827 vdd.n107 vdd.n83 171.744
R1828 vdd.n107 vdd.n106 171.744
R1829 vdd.n106 vdd.n88 171.744
R1830 vdd.n99 vdd.n88 171.744
R1831 vdd.n99 vdd.n98 171.744
R1832 vdd.n98 vdd.n92 171.744
R1833 vdd.n65 vdd.n64 171.744
R1834 vdd.n64 vdd.n63 171.744
R1835 vdd.n63 vdd.n32 171.744
R1836 vdd.n56 vdd.n32 171.744
R1837 vdd.n56 vdd.n55 171.744
R1838 vdd.n55 vdd.n37 171.744
R1839 vdd.n48 vdd.n37 171.744
R1840 vdd.n48 vdd.n47 171.744
R1841 vdd.n47 vdd.n41 171.744
R1842 vdd.n1498 vdd.n1497 171.744
R1843 vdd.n1497 vdd.n1496 171.744
R1844 vdd.n1496 vdd.n1465 171.744
R1845 vdd.n1489 vdd.n1465 171.744
R1846 vdd.n1489 vdd.n1488 171.744
R1847 vdd.n1488 vdd.n1470 171.744
R1848 vdd.n1481 vdd.n1470 171.744
R1849 vdd.n1481 vdd.n1480 171.744
R1850 vdd.n1480 vdd.n1474 171.744
R1851 vdd.n1549 vdd.n1548 171.744
R1852 vdd.n1548 vdd.n1547 171.744
R1853 vdd.n1547 vdd.n1516 171.744
R1854 vdd.n1540 vdd.n1516 171.744
R1855 vdd.n1540 vdd.n1539 171.744
R1856 vdd.n1539 vdd.n1521 171.744
R1857 vdd.n1532 vdd.n1521 171.744
R1858 vdd.n1532 vdd.n1531 171.744
R1859 vdd.n1531 vdd.n1525 171.744
R1860 vdd.n1404 vdd.n1403 171.744
R1861 vdd.n1403 vdd.n1402 171.744
R1862 vdd.n1402 vdd.n1371 171.744
R1863 vdd.n1395 vdd.n1371 171.744
R1864 vdd.n1395 vdd.n1394 171.744
R1865 vdd.n1394 vdd.n1376 171.744
R1866 vdd.n1387 vdd.n1376 171.744
R1867 vdd.n1387 vdd.n1386 171.744
R1868 vdd.n1386 vdd.n1380 171.744
R1869 vdd.n1455 vdd.n1454 171.744
R1870 vdd.n1454 vdd.n1453 171.744
R1871 vdd.n1453 vdd.n1422 171.744
R1872 vdd.n1446 vdd.n1422 171.744
R1873 vdd.n1446 vdd.n1445 171.744
R1874 vdd.n1445 vdd.n1427 171.744
R1875 vdd.n1438 vdd.n1427 171.744
R1876 vdd.n1438 vdd.n1437 171.744
R1877 vdd.n1437 vdd.n1431 171.744
R1878 vdd.n1311 vdd.n1310 171.744
R1879 vdd.n1310 vdd.n1309 171.744
R1880 vdd.n1309 vdd.n1278 171.744
R1881 vdd.n1302 vdd.n1278 171.744
R1882 vdd.n1302 vdd.n1301 171.744
R1883 vdd.n1301 vdd.n1283 171.744
R1884 vdd.n1294 vdd.n1283 171.744
R1885 vdd.n1294 vdd.n1293 171.744
R1886 vdd.n1293 vdd.n1287 171.744
R1887 vdd.n1362 vdd.n1361 171.744
R1888 vdd.n1361 vdd.n1360 171.744
R1889 vdd.n1360 vdd.n1329 171.744
R1890 vdd.n1353 vdd.n1329 171.744
R1891 vdd.n1353 vdd.n1352 171.744
R1892 vdd.n1352 vdd.n1334 171.744
R1893 vdd.n1345 vdd.n1334 171.744
R1894 vdd.n1345 vdd.n1344 171.744
R1895 vdd.n1344 vdd.n1338 171.744
R1896 vdd.n3130 vdd.n356 146.341
R1897 vdd.n3128 vdd.n3127 146.341
R1898 vdd.n3125 vdd.n360 146.341
R1899 vdd.n3121 vdd.n3120 146.341
R1900 vdd.n3118 vdd.n368 146.341
R1901 vdd.n3114 vdd.n3113 146.341
R1902 vdd.n3111 vdd.n375 146.341
R1903 vdd.n3107 vdd.n3106 146.341
R1904 vdd.n3104 vdd.n382 146.341
R1905 vdd.n393 vdd.n390 146.341
R1906 vdd.n3096 vdd.n3095 146.341
R1907 vdd.n3093 vdd.n395 146.341
R1908 vdd.n3089 vdd.n3088 146.341
R1909 vdd.n3086 vdd.n401 146.341
R1910 vdd.n3082 vdd.n3081 146.341
R1911 vdd.n3079 vdd.n408 146.341
R1912 vdd.n3075 vdd.n3074 146.341
R1913 vdd.n3072 vdd.n415 146.341
R1914 vdd.n3068 vdd.n3067 146.341
R1915 vdd.n3065 vdd.n422 146.341
R1916 vdd.n433 vdd.n430 146.341
R1917 vdd.n3057 vdd.n3056 146.341
R1918 vdd.n3054 vdd.n435 146.341
R1919 vdd.n3050 vdd.n3049 146.341
R1920 vdd.n3047 vdd.n441 146.341
R1921 vdd.n3043 vdd.n3042 146.341
R1922 vdd.n3040 vdd.n448 146.341
R1923 vdd.n3036 vdd.n3035 146.341
R1924 vdd.n3033 vdd.n455 146.341
R1925 vdd.n3029 vdd.n3028 146.341
R1926 vdd.n3026 vdd.n462 146.341
R1927 vdd.n2941 vdd.n512 146.341
R1928 vdd.n2947 vdd.n512 146.341
R1929 vdd.n2947 vdd.n504 146.341
R1930 vdd.n2957 vdd.n504 146.341
R1931 vdd.n2957 vdd.n500 146.341
R1932 vdd.n2963 vdd.n500 146.341
R1933 vdd.n2963 vdd.n491 146.341
R1934 vdd.n2973 vdd.n491 146.341
R1935 vdd.n2973 vdd.n487 146.341
R1936 vdd.n2979 vdd.n487 146.341
R1937 vdd.n2979 vdd.n479 146.341
R1938 vdd.n2990 vdd.n479 146.341
R1939 vdd.n2990 vdd.n480 146.341
R1940 vdd.n480 vdd.n316 146.341
R1941 vdd.n317 vdd.n316 146.341
R1942 vdd.n318 vdd.n317 146.341
R1943 vdd.n473 vdd.n318 146.341
R1944 vdd.n473 vdd.n326 146.341
R1945 vdd.n327 vdd.n326 146.341
R1946 vdd.n328 vdd.n327 146.341
R1947 vdd.n470 vdd.n328 146.341
R1948 vdd.n470 vdd.n337 146.341
R1949 vdd.n338 vdd.n337 146.341
R1950 vdd.n339 vdd.n338 146.341
R1951 vdd.n467 vdd.n339 146.341
R1952 vdd.n467 vdd.n348 146.341
R1953 vdd.n349 vdd.n348 146.341
R1954 vdd.n350 vdd.n349 146.341
R1955 vdd.n2933 vdd.n2931 146.341
R1956 vdd.n2931 vdd.n2930 146.341
R1957 vdd.n2927 vdd.n2926 146.341
R1958 vdd.n2923 vdd.n2922 146.341
R1959 vdd.n2920 vdd.n526 146.341
R1960 vdd.n2916 vdd.n2914 146.341
R1961 vdd.n2912 vdd.n532 146.341
R1962 vdd.n2908 vdd.n2906 146.341
R1963 vdd.n2904 vdd.n538 146.341
R1964 vdd.n2900 vdd.n2898 146.341
R1965 vdd.n2896 vdd.n546 146.341
R1966 vdd.n2892 vdd.n2890 146.341
R1967 vdd.n2888 vdd.n552 146.341
R1968 vdd.n2884 vdd.n2882 146.341
R1969 vdd.n2880 vdd.n558 146.341
R1970 vdd.n2876 vdd.n2874 146.341
R1971 vdd.n2872 vdd.n564 146.341
R1972 vdd.n2868 vdd.n2866 146.341
R1973 vdd.n2864 vdd.n570 146.341
R1974 vdd.n2860 vdd.n2858 146.341
R1975 vdd.n2856 vdd.n576 146.341
R1976 vdd.n2849 vdd.n585 146.341
R1977 vdd.n2847 vdd.n2846 146.341
R1978 vdd.n2843 vdd.n2842 146.341
R1979 vdd.n2840 vdd.n590 146.341
R1980 vdd.n2836 vdd.n2834 146.341
R1981 vdd.n2832 vdd.n596 146.341
R1982 vdd.n2828 vdd.n2826 146.341
R1983 vdd.n2824 vdd.n602 146.341
R1984 vdd.n2820 vdd.n2818 146.341
R1985 vdd.n2815 vdd.n2814 146.341
R1986 vdd.n2811 vdd.n515 146.341
R1987 vdd.n2939 vdd.n510 146.341
R1988 vdd.n2949 vdd.n510 146.341
R1989 vdd.n2949 vdd.n506 146.341
R1990 vdd.n2955 vdd.n506 146.341
R1991 vdd.n2955 vdd.n498 146.341
R1992 vdd.n2965 vdd.n498 146.341
R1993 vdd.n2965 vdd.n494 146.341
R1994 vdd.n2971 vdd.n494 146.341
R1995 vdd.n2971 vdd.n486 146.341
R1996 vdd.n2982 vdd.n486 146.341
R1997 vdd.n2982 vdd.n482 146.341
R1998 vdd.n2988 vdd.n482 146.341
R1999 vdd.n2988 vdd.n314 146.341
R2000 vdd.n3165 vdd.n314 146.341
R2001 vdd.n3165 vdd.n315 146.341
R2002 vdd.n3161 vdd.n315 146.341
R2003 vdd.n3161 vdd.n319 146.341
R2004 vdd.n3157 vdd.n319 146.341
R2005 vdd.n3157 vdd.n324 146.341
R2006 vdd.n3153 vdd.n324 146.341
R2007 vdd.n3153 vdd.n330 146.341
R2008 vdd.n3149 vdd.n330 146.341
R2009 vdd.n3149 vdd.n336 146.341
R2010 vdd.n3145 vdd.n336 146.341
R2011 vdd.n3145 vdd.n341 146.341
R2012 vdd.n3141 vdd.n341 146.341
R2013 vdd.n3141 vdd.n347 146.341
R2014 vdd.n3137 vdd.n347 146.341
R2015 vdd.n2034 vdd.n2033 146.341
R2016 vdd.n2031 vdd.n1615 146.341
R2017 vdd.n1811 vdd.n1621 146.341
R2018 vdd.n1809 vdd.n1808 146.341
R2019 vdd.n1806 vdd.n1623 146.341
R2020 vdd.n1802 vdd.n1801 146.341
R2021 vdd.n1799 vdd.n1630 146.341
R2022 vdd.n1795 vdd.n1794 146.341
R2023 vdd.n1792 vdd.n1637 146.341
R2024 vdd.n1648 vdd.n1645 146.341
R2025 vdd.n1784 vdd.n1783 146.341
R2026 vdd.n1781 vdd.n1650 146.341
R2027 vdd.n1777 vdd.n1776 146.341
R2028 vdd.n1774 vdd.n1656 146.341
R2029 vdd.n1770 vdd.n1769 146.341
R2030 vdd.n1767 vdd.n1663 146.341
R2031 vdd.n1763 vdd.n1762 146.341
R2032 vdd.n1760 vdd.n1670 146.341
R2033 vdd.n1756 vdd.n1755 146.341
R2034 vdd.n1753 vdd.n1677 146.341
R2035 vdd.n1688 vdd.n1685 146.341
R2036 vdd.n1745 vdd.n1744 146.341
R2037 vdd.n1742 vdd.n1690 146.341
R2038 vdd.n1738 vdd.n1737 146.341
R2039 vdd.n1735 vdd.n1696 146.341
R2040 vdd.n1731 vdd.n1730 146.341
R2041 vdd.n1728 vdd.n1703 146.341
R2042 vdd.n1724 vdd.n1723 146.341
R2043 vdd.n1721 vdd.n1718 146.341
R2044 vdd.n1716 vdd.n1713 146.341
R2045 vdd.n1711 vdd.n897 146.341
R2046 vdd.n1216 vdd.n978 146.341
R2047 vdd.n1222 vdd.n978 146.341
R2048 vdd.n1222 vdd.n971 146.341
R2049 vdd.n1232 vdd.n971 146.341
R2050 vdd.n1232 vdd.n967 146.341
R2051 vdd.n1238 vdd.n967 146.341
R2052 vdd.n1238 vdd.n958 146.341
R2053 vdd.n1248 vdd.n958 146.341
R2054 vdd.n1248 vdd.n954 146.341
R2055 vdd.n1254 vdd.n954 146.341
R2056 vdd.n1254 vdd.n947 146.341
R2057 vdd.n1265 vdd.n947 146.341
R2058 vdd.n1265 vdd.n943 146.341
R2059 vdd.n1271 vdd.n943 146.341
R2060 vdd.n1271 vdd.n936 146.341
R2061 vdd.n1563 vdd.n936 146.341
R2062 vdd.n1563 vdd.n932 146.341
R2063 vdd.n1569 vdd.n932 146.341
R2064 vdd.n1569 vdd.n924 146.341
R2065 vdd.n1580 vdd.n924 146.341
R2066 vdd.n1580 vdd.n920 146.341
R2067 vdd.n1586 vdd.n920 146.341
R2068 vdd.n1586 vdd.n914 146.341
R2069 vdd.n1597 vdd.n914 146.341
R2070 vdd.n1597 vdd.n909 146.341
R2071 vdd.n1605 vdd.n909 146.341
R2072 vdd.n1605 vdd.n899 146.341
R2073 vdd.n2042 vdd.n899 146.341
R2074 vdd.n988 vdd.n987 146.341
R2075 vdd.n991 vdd.n988 146.341
R2076 vdd.n994 vdd.n993 146.341
R2077 vdd.n999 vdd.n996 146.341
R2078 vdd.n1002 vdd.n1001 146.341
R2079 vdd.n1007 vdd.n1004 146.341
R2080 vdd.n1010 vdd.n1009 146.341
R2081 vdd.n1015 vdd.n1012 146.341
R2082 vdd.n1018 vdd.n1017 146.341
R2083 vdd.n1025 vdd.n1020 146.341
R2084 vdd.n1028 vdd.n1027 146.341
R2085 vdd.n1033 vdd.n1030 146.341
R2086 vdd.n1036 vdd.n1035 146.341
R2087 vdd.n1041 vdd.n1038 146.341
R2088 vdd.n1044 vdd.n1043 146.341
R2089 vdd.n1049 vdd.n1046 146.341
R2090 vdd.n1052 vdd.n1051 146.341
R2091 vdd.n1057 vdd.n1054 146.341
R2092 vdd.n1060 vdd.n1059 146.341
R2093 vdd.n1065 vdd.n1062 146.341
R2094 vdd.n1146 vdd.n1067 146.341
R2095 vdd.n1144 vdd.n1143 146.341
R2096 vdd.n1074 vdd.n1073 146.341
R2097 vdd.n1077 vdd.n1076 146.341
R2098 vdd.n1082 vdd.n1081 146.341
R2099 vdd.n1085 vdd.n1084 146.341
R2100 vdd.n1090 vdd.n1089 146.341
R2101 vdd.n1093 vdd.n1092 146.341
R2102 vdd.n1098 vdd.n1097 146.341
R2103 vdd.n1101 vdd.n1100 146.341
R2104 vdd.n1106 vdd.n1105 146.341
R2105 vdd.n1108 vdd.n981 146.341
R2106 vdd.n1214 vdd.n977 146.341
R2107 vdd.n1224 vdd.n977 146.341
R2108 vdd.n1224 vdd.n973 146.341
R2109 vdd.n1230 vdd.n973 146.341
R2110 vdd.n1230 vdd.n965 146.341
R2111 vdd.n1240 vdd.n965 146.341
R2112 vdd.n1240 vdd.n961 146.341
R2113 vdd.n1246 vdd.n961 146.341
R2114 vdd.n1246 vdd.n953 146.341
R2115 vdd.n1257 vdd.n953 146.341
R2116 vdd.n1257 vdd.n949 146.341
R2117 vdd.n1263 vdd.n949 146.341
R2118 vdd.n1263 vdd.n942 146.341
R2119 vdd.n1273 vdd.n942 146.341
R2120 vdd.n1273 vdd.n938 146.341
R2121 vdd.n1561 vdd.n938 146.341
R2122 vdd.n1561 vdd.n930 146.341
R2123 vdd.n1572 vdd.n930 146.341
R2124 vdd.n1572 vdd.n926 146.341
R2125 vdd.n1578 vdd.n926 146.341
R2126 vdd.n1578 vdd.n919 146.341
R2127 vdd.n1589 vdd.n919 146.341
R2128 vdd.n1589 vdd.n915 146.341
R2129 vdd.n1595 vdd.n915 146.341
R2130 vdd.n1595 vdd.n907 146.341
R2131 vdd.n1608 vdd.n907 146.341
R2132 vdd.n1608 vdd.n902 146.341
R2133 vdd.n2040 vdd.n902 146.341
R2134 vdd.n901 vdd.n877 141.707
R2135 vdd.n613 vdd.n516 141.707
R2136 vdd.n1889 vdd.t59 127.284
R2137 vdd.n793 vdd.t44 127.284
R2138 vdd.n1863 vdd.t10 127.284
R2139 vdd.n785 vdd.t68 127.284
R2140 vdd.n2634 vdd.t31 127.284
R2141 vdd.n2634 vdd.t32 127.284
R2142 vdd.n2354 vdd.t66 127.284
R2143 vdd.n661 vdd.t48 127.284
R2144 vdd.n2351 vdd.t53 127.284
R2145 vdd.n625 vdd.t55 127.284
R2146 vdd.n855 vdd.t62 127.284
R2147 vdd.n855 vdd.t63 127.284
R2148 vdd.n22 vdd.n20 117.314
R2149 vdd.n17 vdd.n15 117.314
R2150 vdd.n27 vdd.n26 116.927
R2151 vdd.n24 vdd.n23 116.927
R2152 vdd.n22 vdd.n21 116.927
R2153 vdd.n17 vdd.n16 116.927
R2154 vdd.n19 vdd.n18 116.927
R2155 vdd.n27 vdd.n25 116.927
R2156 vdd.n1890 vdd.t58 111.188
R2157 vdd.n794 vdd.t45 111.188
R2158 vdd.n1864 vdd.t9 111.188
R2159 vdd.n786 vdd.t69 111.188
R2160 vdd.n2355 vdd.t65 111.188
R2161 vdd.n662 vdd.t49 111.188
R2162 vdd.n2352 vdd.t52 111.188
R2163 vdd.n626 vdd.t56 111.188
R2164 vdd.n2577 vdd.n739 99.5127
R2165 vdd.n2581 vdd.n739 99.5127
R2166 vdd.n2581 vdd.n731 99.5127
R2167 vdd.n2589 vdd.n731 99.5127
R2168 vdd.n2589 vdd.n729 99.5127
R2169 vdd.n2593 vdd.n729 99.5127
R2170 vdd.n2593 vdd.n718 99.5127
R2171 vdd.n2601 vdd.n718 99.5127
R2172 vdd.n2601 vdd.n716 99.5127
R2173 vdd.n2605 vdd.n716 99.5127
R2174 vdd.n2605 vdd.n707 99.5127
R2175 vdd.n2613 vdd.n707 99.5127
R2176 vdd.n2613 vdd.n705 99.5127
R2177 vdd.n2617 vdd.n705 99.5127
R2178 vdd.n2617 vdd.n695 99.5127
R2179 vdd.n2625 vdd.n695 99.5127
R2180 vdd.n2625 vdd.n693 99.5127
R2181 vdd.n2629 vdd.n693 99.5127
R2182 vdd.n2629 vdd.n684 99.5127
R2183 vdd.n2639 vdd.n684 99.5127
R2184 vdd.n2639 vdd.n682 99.5127
R2185 vdd.n2643 vdd.n682 99.5127
R2186 vdd.n2643 vdd.n670 99.5127
R2187 vdd.n2696 vdd.n670 99.5127
R2188 vdd.n2696 vdd.n668 99.5127
R2189 vdd.n2700 vdd.n668 99.5127
R2190 vdd.n2700 vdd.n634 99.5127
R2191 vdd.n2770 vdd.n634 99.5127
R2192 vdd.n2766 vdd.n635 99.5127
R2193 vdd.n2764 vdd.n2763 99.5127
R2194 vdd.n2761 vdd.n639 99.5127
R2195 vdd.n2757 vdd.n2756 99.5127
R2196 vdd.n2754 vdd.n642 99.5127
R2197 vdd.n2750 vdd.n2749 99.5127
R2198 vdd.n2747 vdd.n645 99.5127
R2199 vdd.n2743 vdd.n2742 99.5127
R2200 vdd.n2740 vdd.n648 99.5127
R2201 vdd.n2735 vdd.n2734 99.5127
R2202 vdd.n2732 vdd.n651 99.5127
R2203 vdd.n2728 vdd.n2727 99.5127
R2204 vdd.n2725 vdd.n654 99.5127
R2205 vdd.n2721 vdd.n2720 99.5127
R2206 vdd.n2718 vdd.n657 99.5127
R2207 vdd.n2714 vdd.n2713 99.5127
R2208 vdd.n2711 vdd.n660 99.5127
R2209 vdd.n2497 vdd.n742 99.5127
R2210 vdd.n2497 vdd.n737 99.5127
R2211 vdd.n2494 vdd.n737 99.5127
R2212 vdd.n2494 vdd.n732 99.5127
R2213 vdd.n2441 vdd.n732 99.5127
R2214 vdd.n2441 vdd.n726 99.5127
R2215 vdd.n2444 vdd.n726 99.5127
R2216 vdd.n2444 vdd.n719 99.5127
R2217 vdd.n2447 vdd.n719 99.5127
R2218 vdd.n2447 vdd.n714 99.5127
R2219 vdd.n2450 vdd.n714 99.5127
R2220 vdd.n2450 vdd.n709 99.5127
R2221 vdd.n2453 vdd.n709 99.5127
R2222 vdd.n2453 vdd.n703 99.5127
R2223 vdd.n2471 vdd.n703 99.5127
R2224 vdd.n2471 vdd.n696 99.5127
R2225 vdd.n2467 vdd.n696 99.5127
R2226 vdd.n2467 vdd.n691 99.5127
R2227 vdd.n2464 vdd.n691 99.5127
R2228 vdd.n2464 vdd.n686 99.5127
R2229 vdd.n2461 vdd.n686 99.5127
R2230 vdd.n2461 vdd.n680 99.5127
R2231 vdd.n2458 vdd.n680 99.5127
R2232 vdd.n2458 vdd.n672 99.5127
R2233 vdd.n672 vdd.n665 99.5127
R2234 vdd.n2702 vdd.n665 99.5127
R2235 vdd.n2703 vdd.n2702 99.5127
R2236 vdd.n2703 vdd.n632 99.5127
R2237 vdd.n2567 vdd.n2350 99.5127
R2238 vdd.n2563 vdd.n2350 99.5127
R2239 vdd.n2561 vdd.n2560 99.5127
R2240 vdd.n2557 vdd.n2556 99.5127
R2241 vdd.n2553 vdd.n2552 99.5127
R2242 vdd.n2549 vdd.n2548 99.5127
R2243 vdd.n2545 vdd.n2544 99.5127
R2244 vdd.n2541 vdd.n2540 99.5127
R2245 vdd.n2537 vdd.n2536 99.5127
R2246 vdd.n2533 vdd.n2532 99.5127
R2247 vdd.n2529 vdd.n2528 99.5127
R2248 vdd.n2525 vdd.n2524 99.5127
R2249 vdd.n2521 vdd.n2520 99.5127
R2250 vdd.n2517 vdd.n2516 99.5127
R2251 vdd.n2513 vdd.n2512 99.5127
R2252 vdd.n2509 vdd.n2508 99.5127
R2253 vdd.n2504 vdd.n2503 99.5127
R2254 vdd.n2315 vdd.n783 99.5127
R2255 vdd.n2311 vdd.n2310 99.5127
R2256 vdd.n2307 vdd.n2306 99.5127
R2257 vdd.n2303 vdd.n2302 99.5127
R2258 vdd.n2299 vdd.n2298 99.5127
R2259 vdd.n2295 vdd.n2294 99.5127
R2260 vdd.n2291 vdd.n2290 99.5127
R2261 vdd.n2287 vdd.n2286 99.5127
R2262 vdd.n2283 vdd.n2282 99.5127
R2263 vdd.n2279 vdd.n2278 99.5127
R2264 vdd.n2275 vdd.n2274 99.5127
R2265 vdd.n2271 vdd.n2270 99.5127
R2266 vdd.n2267 vdd.n2266 99.5127
R2267 vdd.n2263 vdd.n2262 99.5127
R2268 vdd.n2259 vdd.n2258 99.5127
R2269 vdd.n2255 vdd.n2254 99.5127
R2270 vdd.n2250 vdd.n2249 99.5127
R2271 vdd.n1988 vdd.n878 99.5127
R2272 vdd.n1988 vdd.n872 99.5127
R2273 vdd.n1985 vdd.n872 99.5127
R2274 vdd.n1985 vdd.n866 99.5127
R2275 vdd.n1982 vdd.n866 99.5127
R2276 vdd.n1982 vdd.n859 99.5127
R2277 vdd.n1979 vdd.n859 99.5127
R2278 vdd.n1979 vdd.n852 99.5127
R2279 vdd.n1976 vdd.n852 99.5127
R2280 vdd.n1976 vdd.n847 99.5127
R2281 vdd.n1973 vdd.n847 99.5127
R2282 vdd.n1973 vdd.n841 99.5127
R2283 vdd.n1970 vdd.n841 99.5127
R2284 vdd.n1970 vdd.n834 99.5127
R2285 vdd.n1884 vdd.n834 99.5127
R2286 vdd.n1884 vdd.n828 99.5127
R2287 vdd.n1881 vdd.n828 99.5127
R2288 vdd.n1881 vdd.n823 99.5127
R2289 vdd.n1878 vdd.n823 99.5127
R2290 vdd.n1878 vdd.n818 99.5127
R2291 vdd.n1875 vdd.n818 99.5127
R2292 vdd.n1875 vdd.n812 99.5127
R2293 vdd.n1872 vdd.n812 99.5127
R2294 vdd.n1872 vdd.n805 99.5127
R2295 vdd.n1869 vdd.n805 99.5127
R2296 vdd.n1869 vdd.n798 99.5127
R2297 vdd.n798 vdd.n788 99.5127
R2298 vdd.n2245 vdd.n788 99.5127
R2299 vdd.n1823 vdd.n1821 99.5127
R2300 vdd.n1827 vdd.n1821 99.5127
R2301 vdd.n1831 vdd.n1829 99.5127
R2302 vdd.n1835 vdd.n1819 99.5127
R2303 vdd.n1839 vdd.n1837 99.5127
R2304 vdd.n1843 vdd.n1817 99.5127
R2305 vdd.n1847 vdd.n1845 99.5127
R2306 vdd.n1851 vdd.n1815 99.5127
R2307 vdd.n1854 vdd.n1853 99.5127
R2308 vdd.n2024 vdd.n2022 99.5127
R2309 vdd.n2020 vdd.n1856 99.5127
R2310 vdd.n2016 vdd.n2014 99.5127
R2311 vdd.n2012 vdd.n1858 99.5127
R2312 vdd.n2008 vdd.n2006 99.5127
R2313 vdd.n2004 vdd.n1860 99.5127
R2314 vdd.n2000 vdd.n1998 99.5127
R2315 vdd.n1996 vdd.n1862 99.5127
R2316 vdd.n2088 vdd.n874 99.5127
R2317 vdd.n2092 vdd.n874 99.5127
R2318 vdd.n2092 vdd.n864 99.5127
R2319 vdd.n2100 vdd.n864 99.5127
R2320 vdd.n2100 vdd.n862 99.5127
R2321 vdd.n2104 vdd.n862 99.5127
R2322 vdd.n2104 vdd.n851 99.5127
R2323 vdd.n2113 vdd.n851 99.5127
R2324 vdd.n2113 vdd.n849 99.5127
R2325 vdd.n2117 vdd.n849 99.5127
R2326 vdd.n2117 vdd.n839 99.5127
R2327 vdd.n2125 vdd.n839 99.5127
R2328 vdd.n2125 vdd.n837 99.5127
R2329 vdd.n2129 vdd.n837 99.5127
R2330 vdd.n2129 vdd.n827 99.5127
R2331 vdd.n2137 vdd.n827 99.5127
R2332 vdd.n2137 vdd.n825 99.5127
R2333 vdd.n2141 vdd.n825 99.5127
R2334 vdd.n2141 vdd.n816 99.5127
R2335 vdd.n2149 vdd.n816 99.5127
R2336 vdd.n2149 vdd.n814 99.5127
R2337 vdd.n2153 vdd.n814 99.5127
R2338 vdd.n2153 vdd.n803 99.5127
R2339 vdd.n2163 vdd.n803 99.5127
R2340 vdd.n2163 vdd.n800 99.5127
R2341 vdd.n2168 vdd.n800 99.5127
R2342 vdd.n2168 vdd.n801 99.5127
R2343 vdd.n801 vdd.n782 99.5127
R2344 vdd.n2686 vdd.n2685 99.5127
R2345 vdd.n2683 vdd.n2649 99.5127
R2346 vdd.n2679 vdd.n2678 99.5127
R2347 vdd.n2676 vdd.n2652 99.5127
R2348 vdd.n2672 vdd.n2671 99.5127
R2349 vdd.n2669 vdd.n2655 99.5127
R2350 vdd.n2665 vdd.n2664 99.5127
R2351 vdd.n2662 vdd.n2659 99.5127
R2352 vdd.n2803 vdd.n612 99.5127
R2353 vdd.n2801 vdd.n2800 99.5127
R2354 vdd.n2798 vdd.n615 99.5127
R2355 vdd.n2794 vdd.n2793 99.5127
R2356 vdd.n2791 vdd.n618 99.5127
R2357 vdd.n2787 vdd.n2786 99.5127
R2358 vdd.n2784 vdd.n621 99.5127
R2359 vdd.n2780 vdd.n2779 99.5127
R2360 vdd.n2777 vdd.n624 99.5127
R2361 vdd.n2421 vdd.n743 99.5127
R2362 vdd.n2421 vdd.n738 99.5127
R2363 vdd.n2492 vdd.n738 99.5127
R2364 vdd.n2492 vdd.n733 99.5127
R2365 vdd.n2488 vdd.n733 99.5127
R2366 vdd.n2488 vdd.n727 99.5127
R2367 vdd.n2485 vdd.n727 99.5127
R2368 vdd.n2485 vdd.n720 99.5127
R2369 vdd.n2482 vdd.n720 99.5127
R2370 vdd.n2482 vdd.n715 99.5127
R2371 vdd.n2479 vdd.n715 99.5127
R2372 vdd.n2479 vdd.n710 99.5127
R2373 vdd.n2476 vdd.n710 99.5127
R2374 vdd.n2476 vdd.n704 99.5127
R2375 vdd.n2473 vdd.n704 99.5127
R2376 vdd.n2473 vdd.n697 99.5127
R2377 vdd.n2438 vdd.n697 99.5127
R2378 vdd.n2438 vdd.n692 99.5127
R2379 vdd.n2435 vdd.n692 99.5127
R2380 vdd.n2435 vdd.n687 99.5127
R2381 vdd.n2432 vdd.n687 99.5127
R2382 vdd.n2432 vdd.n681 99.5127
R2383 vdd.n2429 vdd.n681 99.5127
R2384 vdd.n2429 vdd.n673 99.5127
R2385 vdd.n2426 vdd.n673 99.5127
R2386 vdd.n2426 vdd.n666 99.5127
R2387 vdd.n666 vdd.n630 99.5127
R2388 vdd.n2772 vdd.n630 99.5127
R2389 vdd.n2571 vdd.n746 99.5127
R2390 vdd.n2359 vdd.n2358 99.5127
R2391 vdd.n2363 vdd.n2362 99.5127
R2392 vdd.n2367 vdd.n2366 99.5127
R2393 vdd.n2371 vdd.n2370 99.5127
R2394 vdd.n2375 vdd.n2374 99.5127
R2395 vdd.n2379 vdd.n2378 99.5127
R2396 vdd.n2383 vdd.n2382 99.5127
R2397 vdd.n2387 vdd.n2386 99.5127
R2398 vdd.n2391 vdd.n2390 99.5127
R2399 vdd.n2395 vdd.n2394 99.5127
R2400 vdd.n2399 vdd.n2398 99.5127
R2401 vdd.n2403 vdd.n2402 99.5127
R2402 vdd.n2407 vdd.n2406 99.5127
R2403 vdd.n2411 vdd.n2410 99.5127
R2404 vdd.n2415 vdd.n2414 99.5127
R2405 vdd.n2417 vdd.n2349 99.5127
R2406 vdd.n2575 vdd.n736 99.5127
R2407 vdd.n2583 vdd.n736 99.5127
R2408 vdd.n2583 vdd.n734 99.5127
R2409 vdd.n2587 vdd.n734 99.5127
R2410 vdd.n2587 vdd.n724 99.5127
R2411 vdd.n2595 vdd.n724 99.5127
R2412 vdd.n2595 vdd.n722 99.5127
R2413 vdd.n2599 vdd.n722 99.5127
R2414 vdd.n2599 vdd.n713 99.5127
R2415 vdd.n2607 vdd.n713 99.5127
R2416 vdd.n2607 vdd.n711 99.5127
R2417 vdd.n2611 vdd.n711 99.5127
R2418 vdd.n2611 vdd.n701 99.5127
R2419 vdd.n2619 vdd.n701 99.5127
R2420 vdd.n2619 vdd.n699 99.5127
R2421 vdd.n2623 vdd.n699 99.5127
R2422 vdd.n2623 vdd.n690 99.5127
R2423 vdd.n2631 vdd.n690 99.5127
R2424 vdd.n2631 vdd.n688 99.5127
R2425 vdd.n2637 vdd.n688 99.5127
R2426 vdd.n2637 vdd.n678 99.5127
R2427 vdd.n2645 vdd.n678 99.5127
R2428 vdd.n2645 vdd.n675 99.5127
R2429 vdd.n2694 vdd.n675 99.5127
R2430 vdd.n2694 vdd.n676 99.5127
R2431 vdd.n676 vdd.n667 99.5127
R2432 vdd.n2689 vdd.n667 99.5127
R2433 vdd.n2689 vdd.n633 99.5127
R2434 vdd.n2239 vdd.n2238 99.5127
R2435 vdd.n2235 vdd.n2234 99.5127
R2436 vdd.n2231 vdd.n2230 99.5127
R2437 vdd.n2227 vdd.n2226 99.5127
R2438 vdd.n2223 vdd.n2222 99.5127
R2439 vdd.n2219 vdd.n2218 99.5127
R2440 vdd.n2215 vdd.n2214 99.5127
R2441 vdd.n2211 vdd.n2210 99.5127
R2442 vdd.n2207 vdd.n2206 99.5127
R2443 vdd.n2203 vdd.n2202 99.5127
R2444 vdd.n2199 vdd.n2198 99.5127
R2445 vdd.n2195 vdd.n2194 99.5127
R2446 vdd.n2191 vdd.n2190 99.5127
R2447 vdd.n2187 vdd.n2186 99.5127
R2448 vdd.n2183 vdd.n2182 99.5127
R2449 vdd.n2179 vdd.n2178 99.5127
R2450 vdd.n2175 vdd.n764 99.5127
R2451 vdd.n1932 vdd.n879 99.5127
R2452 vdd.n1932 vdd.n873 99.5127
R2453 vdd.n1935 vdd.n873 99.5127
R2454 vdd.n1935 vdd.n867 99.5127
R2455 vdd.n1938 vdd.n867 99.5127
R2456 vdd.n1938 vdd.n860 99.5127
R2457 vdd.n1941 vdd.n860 99.5127
R2458 vdd.n1941 vdd.n853 99.5127
R2459 vdd.n1944 vdd.n853 99.5127
R2460 vdd.n1944 vdd.n848 99.5127
R2461 vdd.n1947 vdd.n848 99.5127
R2462 vdd.n1947 vdd.n842 99.5127
R2463 vdd.n1968 vdd.n842 99.5127
R2464 vdd.n1968 vdd.n835 99.5127
R2465 vdd.n1964 vdd.n835 99.5127
R2466 vdd.n1964 vdd.n829 99.5127
R2467 vdd.n1961 vdd.n829 99.5127
R2468 vdd.n1961 vdd.n824 99.5127
R2469 vdd.n1958 vdd.n824 99.5127
R2470 vdd.n1958 vdd.n819 99.5127
R2471 vdd.n1955 vdd.n819 99.5127
R2472 vdd.n1955 vdd.n813 99.5127
R2473 vdd.n1952 vdd.n813 99.5127
R2474 vdd.n1952 vdd.n806 99.5127
R2475 vdd.n806 vdd.n797 99.5127
R2476 vdd.n2170 vdd.n797 99.5127
R2477 vdd.n2171 vdd.n2170 99.5127
R2478 vdd.n2171 vdd.n789 99.5127
R2479 vdd.n2082 vdd.n2080 99.5127
R2480 vdd.n2078 vdd.n882 99.5127
R2481 vdd.n2074 vdd.n2072 99.5127
R2482 vdd.n2070 vdd.n884 99.5127
R2483 vdd.n2066 vdd.n2064 99.5127
R2484 vdd.n2062 vdd.n886 99.5127
R2485 vdd.n2058 vdd.n2056 99.5127
R2486 vdd.n2054 vdd.n888 99.5127
R2487 vdd.n1896 vdd.n890 99.5127
R2488 vdd.n1901 vdd.n1898 99.5127
R2489 vdd.n1905 vdd.n1903 99.5127
R2490 vdd.n1909 vdd.n1894 99.5127
R2491 vdd.n1913 vdd.n1911 99.5127
R2492 vdd.n1917 vdd.n1892 99.5127
R2493 vdd.n1921 vdd.n1919 99.5127
R2494 vdd.n1926 vdd.n1888 99.5127
R2495 vdd.n1929 vdd.n1928 99.5127
R2496 vdd.n2086 vdd.n870 99.5127
R2497 vdd.n2094 vdd.n870 99.5127
R2498 vdd.n2094 vdd.n868 99.5127
R2499 vdd.n2098 vdd.n868 99.5127
R2500 vdd.n2098 vdd.n857 99.5127
R2501 vdd.n2106 vdd.n857 99.5127
R2502 vdd.n2106 vdd.n854 99.5127
R2503 vdd.n2111 vdd.n854 99.5127
R2504 vdd.n2111 vdd.n845 99.5127
R2505 vdd.n2119 vdd.n845 99.5127
R2506 vdd.n2119 vdd.n843 99.5127
R2507 vdd.n2123 vdd.n843 99.5127
R2508 vdd.n2123 vdd.n833 99.5127
R2509 vdd.n2131 vdd.n833 99.5127
R2510 vdd.n2131 vdd.n831 99.5127
R2511 vdd.n2135 vdd.n831 99.5127
R2512 vdd.n2135 vdd.n822 99.5127
R2513 vdd.n2143 vdd.n822 99.5127
R2514 vdd.n2143 vdd.n820 99.5127
R2515 vdd.n2147 vdd.n820 99.5127
R2516 vdd.n2147 vdd.n810 99.5127
R2517 vdd.n2155 vdd.n810 99.5127
R2518 vdd.n2155 vdd.n807 99.5127
R2519 vdd.n2161 vdd.n807 99.5127
R2520 vdd.n2161 vdd.n808 99.5127
R2521 vdd.n808 vdd.n799 99.5127
R2522 vdd.n799 vdd.n790 99.5127
R2523 vdd.n2243 vdd.n790 99.5127
R2524 vdd.n9 vdd.n7 98.9633
R2525 vdd.n2 vdd.n0 98.9633
R2526 vdd.n9 vdd.n8 98.6055
R2527 vdd.n11 vdd.n10 98.6055
R2528 vdd.n13 vdd.n12 98.6055
R2529 vdd.n6 vdd.n5 98.6055
R2530 vdd.n4 vdd.n3 98.6055
R2531 vdd.n2 vdd.n1 98.6055
R2532 vdd.t173 vdd.n279 85.8723
R2533 vdd.t191 vdd.n228 85.8723
R2534 vdd.t166 vdd.n185 85.8723
R2535 vdd.t186 vdd.n134 85.8723
R2536 vdd.t154 vdd.n92 85.8723
R2537 vdd.t135 vdd.n41 85.8723
R2538 vdd.t224 vdd.n1474 85.8723
R2539 vdd.t203 vdd.n1525 85.8723
R2540 vdd.t212 vdd.n1380 85.8723
R2541 vdd.t194 vdd.n1431 85.8723
R2542 vdd.t137 vdd.n1287 85.8723
R2543 vdd.t156 vdd.n1338 85.8723
R2544 vdd.n2635 vdd.n2634 78.546
R2545 vdd.n2109 vdd.n855 78.546
R2546 vdd.n266 vdd.n265 75.1835
R2547 vdd.n264 vdd.n263 75.1835
R2548 vdd.n262 vdd.n261 75.1835
R2549 vdd.n260 vdd.n259 75.1835
R2550 vdd.n258 vdd.n257 75.1835
R2551 vdd.n172 vdd.n171 75.1835
R2552 vdd.n170 vdd.n169 75.1835
R2553 vdd.n168 vdd.n167 75.1835
R2554 vdd.n166 vdd.n165 75.1835
R2555 vdd.n164 vdd.n163 75.1835
R2556 vdd.n79 vdd.n78 75.1835
R2557 vdd.n77 vdd.n76 75.1835
R2558 vdd.n75 vdd.n74 75.1835
R2559 vdd.n73 vdd.n72 75.1835
R2560 vdd.n71 vdd.n70 75.1835
R2561 vdd.n1504 vdd.n1503 75.1835
R2562 vdd.n1506 vdd.n1505 75.1835
R2563 vdd.n1508 vdd.n1507 75.1835
R2564 vdd.n1510 vdd.n1509 75.1835
R2565 vdd.n1512 vdd.n1511 75.1835
R2566 vdd.n1410 vdd.n1409 75.1835
R2567 vdd.n1412 vdd.n1411 75.1835
R2568 vdd.n1414 vdd.n1413 75.1835
R2569 vdd.n1416 vdd.n1415 75.1835
R2570 vdd.n1418 vdd.n1417 75.1835
R2571 vdd.n1317 vdd.n1316 75.1835
R2572 vdd.n1319 vdd.n1318 75.1835
R2573 vdd.n1321 vdd.n1320 75.1835
R2574 vdd.n1323 vdd.n1322 75.1835
R2575 vdd.n1325 vdd.n1324 75.1835
R2576 vdd.n2570 vdd.n2569 72.8958
R2577 vdd.n2569 vdd.n2333 72.8958
R2578 vdd.n2569 vdd.n2334 72.8958
R2579 vdd.n2569 vdd.n2335 72.8958
R2580 vdd.n2569 vdd.n2336 72.8958
R2581 vdd.n2569 vdd.n2337 72.8958
R2582 vdd.n2569 vdd.n2338 72.8958
R2583 vdd.n2569 vdd.n2339 72.8958
R2584 vdd.n2569 vdd.n2340 72.8958
R2585 vdd.n2569 vdd.n2341 72.8958
R2586 vdd.n2569 vdd.n2342 72.8958
R2587 vdd.n2569 vdd.n2343 72.8958
R2588 vdd.n2569 vdd.n2344 72.8958
R2589 vdd.n2569 vdd.n2345 72.8958
R2590 vdd.n2569 vdd.n2346 72.8958
R2591 vdd.n2569 vdd.n2347 72.8958
R2592 vdd.n2569 vdd.n2348 72.8958
R2593 vdd.n629 vdd.n613 72.8958
R2594 vdd.n2778 vdd.n613 72.8958
R2595 vdd.n623 vdd.n613 72.8958
R2596 vdd.n2785 vdd.n613 72.8958
R2597 vdd.n620 vdd.n613 72.8958
R2598 vdd.n2792 vdd.n613 72.8958
R2599 vdd.n617 vdd.n613 72.8958
R2600 vdd.n2799 vdd.n613 72.8958
R2601 vdd.n2802 vdd.n613 72.8958
R2602 vdd.n2658 vdd.n613 72.8958
R2603 vdd.n2663 vdd.n613 72.8958
R2604 vdd.n2657 vdd.n613 72.8958
R2605 vdd.n2670 vdd.n613 72.8958
R2606 vdd.n2654 vdd.n613 72.8958
R2607 vdd.n2677 vdd.n613 72.8958
R2608 vdd.n2651 vdd.n613 72.8958
R2609 vdd.n2684 vdd.n613 72.8958
R2610 vdd.n1822 vdd.n877 72.8958
R2611 vdd.n1828 vdd.n877 72.8958
R2612 vdd.n1830 vdd.n877 72.8958
R2613 vdd.n1836 vdd.n877 72.8958
R2614 vdd.n1838 vdd.n877 72.8958
R2615 vdd.n1844 vdd.n877 72.8958
R2616 vdd.n1846 vdd.n877 72.8958
R2617 vdd.n1852 vdd.n877 72.8958
R2618 vdd.n2023 vdd.n877 72.8958
R2619 vdd.n2021 vdd.n877 72.8958
R2620 vdd.n2015 vdd.n877 72.8958
R2621 vdd.n2013 vdd.n877 72.8958
R2622 vdd.n2007 vdd.n877 72.8958
R2623 vdd.n2005 vdd.n877 72.8958
R2624 vdd.n1999 vdd.n877 72.8958
R2625 vdd.n1997 vdd.n877 72.8958
R2626 vdd.n1991 vdd.n877 72.8958
R2627 vdd.n2316 vdd.n765 72.8958
R2628 vdd.n2316 vdd.n766 72.8958
R2629 vdd.n2316 vdd.n767 72.8958
R2630 vdd.n2316 vdd.n768 72.8958
R2631 vdd.n2316 vdd.n769 72.8958
R2632 vdd.n2316 vdd.n770 72.8958
R2633 vdd.n2316 vdd.n771 72.8958
R2634 vdd.n2316 vdd.n772 72.8958
R2635 vdd.n2316 vdd.n773 72.8958
R2636 vdd.n2316 vdd.n774 72.8958
R2637 vdd.n2316 vdd.n775 72.8958
R2638 vdd.n2316 vdd.n776 72.8958
R2639 vdd.n2316 vdd.n777 72.8958
R2640 vdd.n2316 vdd.n778 72.8958
R2641 vdd.n2316 vdd.n779 72.8958
R2642 vdd.n2316 vdd.n780 72.8958
R2643 vdd.n2316 vdd.n781 72.8958
R2644 vdd.n2569 vdd.n2568 72.8958
R2645 vdd.n2569 vdd.n2317 72.8958
R2646 vdd.n2569 vdd.n2318 72.8958
R2647 vdd.n2569 vdd.n2319 72.8958
R2648 vdd.n2569 vdd.n2320 72.8958
R2649 vdd.n2569 vdd.n2321 72.8958
R2650 vdd.n2569 vdd.n2322 72.8958
R2651 vdd.n2569 vdd.n2323 72.8958
R2652 vdd.n2569 vdd.n2324 72.8958
R2653 vdd.n2569 vdd.n2325 72.8958
R2654 vdd.n2569 vdd.n2326 72.8958
R2655 vdd.n2569 vdd.n2327 72.8958
R2656 vdd.n2569 vdd.n2328 72.8958
R2657 vdd.n2569 vdd.n2329 72.8958
R2658 vdd.n2569 vdd.n2330 72.8958
R2659 vdd.n2569 vdd.n2331 72.8958
R2660 vdd.n2569 vdd.n2332 72.8958
R2661 vdd.n2706 vdd.n613 72.8958
R2662 vdd.n2712 vdd.n613 72.8958
R2663 vdd.n659 vdd.n613 72.8958
R2664 vdd.n2719 vdd.n613 72.8958
R2665 vdd.n656 vdd.n613 72.8958
R2666 vdd.n2726 vdd.n613 72.8958
R2667 vdd.n653 vdd.n613 72.8958
R2668 vdd.n2733 vdd.n613 72.8958
R2669 vdd.n650 vdd.n613 72.8958
R2670 vdd.n2741 vdd.n613 72.8958
R2671 vdd.n647 vdd.n613 72.8958
R2672 vdd.n2748 vdd.n613 72.8958
R2673 vdd.n644 vdd.n613 72.8958
R2674 vdd.n2755 vdd.n613 72.8958
R2675 vdd.n641 vdd.n613 72.8958
R2676 vdd.n2762 vdd.n613 72.8958
R2677 vdd.n2765 vdd.n613 72.8958
R2678 vdd.n2316 vdd.n763 72.8958
R2679 vdd.n2316 vdd.n762 72.8958
R2680 vdd.n2316 vdd.n761 72.8958
R2681 vdd.n2316 vdd.n760 72.8958
R2682 vdd.n2316 vdd.n759 72.8958
R2683 vdd.n2316 vdd.n758 72.8958
R2684 vdd.n2316 vdd.n757 72.8958
R2685 vdd.n2316 vdd.n756 72.8958
R2686 vdd.n2316 vdd.n755 72.8958
R2687 vdd.n2316 vdd.n754 72.8958
R2688 vdd.n2316 vdd.n753 72.8958
R2689 vdd.n2316 vdd.n752 72.8958
R2690 vdd.n2316 vdd.n751 72.8958
R2691 vdd.n2316 vdd.n750 72.8958
R2692 vdd.n2316 vdd.n749 72.8958
R2693 vdd.n2316 vdd.n748 72.8958
R2694 vdd.n2316 vdd.n747 72.8958
R2695 vdd.n2081 vdd.n877 72.8958
R2696 vdd.n2079 vdd.n877 72.8958
R2697 vdd.n2073 vdd.n877 72.8958
R2698 vdd.n2071 vdd.n877 72.8958
R2699 vdd.n2065 vdd.n877 72.8958
R2700 vdd.n2063 vdd.n877 72.8958
R2701 vdd.n2057 vdd.n877 72.8958
R2702 vdd.n2055 vdd.n877 72.8958
R2703 vdd.n889 vdd.n877 72.8958
R2704 vdd.n1897 vdd.n877 72.8958
R2705 vdd.n1902 vdd.n877 72.8958
R2706 vdd.n1904 vdd.n877 72.8958
R2707 vdd.n1910 vdd.n877 72.8958
R2708 vdd.n1912 vdd.n877 72.8958
R2709 vdd.n1918 vdd.n877 72.8958
R2710 vdd.n1920 vdd.n877 72.8958
R2711 vdd.n1927 vdd.n877 72.8958
R2712 vdd.n986 vdd.n982 66.2847
R2713 vdd.n992 vdd.n982 66.2847
R2714 vdd.n995 vdd.n982 66.2847
R2715 vdd.n1000 vdd.n982 66.2847
R2716 vdd.n1003 vdd.n982 66.2847
R2717 vdd.n1008 vdd.n982 66.2847
R2718 vdd.n1011 vdd.n982 66.2847
R2719 vdd.n1016 vdd.n982 66.2847
R2720 vdd.n1019 vdd.n982 66.2847
R2721 vdd.n1026 vdd.n982 66.2847
R2722 vdd.n1029 vdd.n982 66.2847
R2723 vdd.n1034 vdd.n982 66.2847
R2724 vdd.n1037 vdd.n982 66.2847
R2725 vdd.n1042 vdd.n982 66.2847
R2726 vdd.n1045 vdd.n982 66.2847
R2727 vdd.n1050 vdd.n982 66.2847
R2728 vdd.n1053 vdd.n982 66.2847
R2729 vdd.n1058 vdd.n982 66.2847
R2730 vdd.n1061 vdd.n982 66.2847
R2731 vdd.n1066 vdd.n982 66.2847
R2732 vdd.n1145 vdd.n982 66.2847
R2733 vdd.n1069 vdd.n982 66.2847
R2734 vdd.n1075 vdd.n982 66.2847
R2735 vdd.n1080 vdd.n982 66.2847
R2736 vdd.n1083 vdd.n982 66.2847
R2737 vdd.n1088 vdd.n982 66.2847
R2738 vdd.n1091 vdd.n982 66.2847
R2739 vdd.n1096 vdd.n982 66.2847
R2740 vdd.n1099 vdd.n982 66.2847
R2741 vdd.n1104 vdd.n982 66.2847
R2742 vdd.n1107 vdd.n982 66.2847
R2743 vdd.n901 vdd.n898 66.2847
R2744 vdd.n1712 vdd.n901 66.2847
R2745 vdd.n1717 vdd.n901 66.2847
R2746 vdd.n1722 vdd.n901 66.2847
R2747 vdd.n1710 vdd.n901 66.2847
R2748 vdd.n1729 vdd.n901 66.2847
R2749 vdd.n1702 vdd.n901 66.2847
R2750 vdd.n1736 vdd.n901 66.2847
R2751 vdd.n1695 vdd.n901 66.2847
R2752 vdd.n1743 vdd.n901 66.2847
R2753 vdd.n1689 vdd.n901 66.2847
R2754 vdd.n1684 vdd.n901 66.2847
R2755 vdd.n1754 vdd.n901 66.2847
R2756 vdd.n1676 vdd.n901 66.2847
R2757 vdd.n1761 vdd.n901 66.2847
R2758 vdd.n1669 vdd.n901 66.2847
R2759 vdd.n1768 vdd.n901 66.2847
R2760 vdd.n1662 vdd.n901 66.2847
R2761 vdd.n1775 vdd.n901 66.2847
R2762 vdd.n1655 vdd.n901 66.2847
R2763 vdd.n1782 vdd.n901 66.2847
R2764 vdd.n1649 vdd.n901 66.2847
R2765 vdd.n1644 vdd.n901 66.2847
R2766 vdd.n1793 vdd.n901 66.2847
R2767 vdd.n1636 vdd.n901 66.2847
R2768 vdd.n1800 vdd.n901 66.2847
R2769 vdd.n1629 vdd.n901 66.2847
R2770 vdd.n1807 vdd.n901 66.2847
R2771 vdd.n1810 vdd.n901 66.2847
R2772 vdd.n1620 vdd.n901 66.2847
R2773 vdd.n2032 vdd.n901 66.2847
R2774 vdd.n1614 vdd.n901 66.2847
R2775 vdd.n2932 vdd.n516 66.2847
R2776 vdd.n520 vdd.n516 66.2847
R2777 vdd.n523 vdd.n516 66.2847
R2778 vdd.n2921 vdd.n516 66.2847
R2779 vdd.n2915 vdd.n516 66.2847
R2780 vdd.n2913 vdd.n516 66.2847
R2781 vdd.n2907 vdd.n516 66.2847
R2782 vdd.n2905 vdd.n516 66.2847
R2783 vdd.n2899 vdd.n516 66.2847
R2784 vdd.n2897 vdd.n516 66.2847
R2785 vdd.n2891 vdd.n516 66.2847
R2786 vdd.n2889 vdd.n516 66.2847
R2787 vdd.n2883 vdd.n516 66.2847
R2788 vdd.n2881 vdd.n516 66.2847
R2789 vdd.n2875 vdd.n516 66.2847
R2790 vdd.n2873 vdd.n516 66.2847
R2791 vdd.n2867 vdd.n516 66.2847
R2792 vdd.n2865 vdd.n516 66.2847
R2793 vdd.n2859 vdd.n516 66.2847
R2794 vdd.n2857 vdd.n516 66.2847
R2795 vdd.n584 vdd.n516 66.2847
R2796 vdd.n2848 vdd.n516 66.2847
R2797 vdd.n586 vdd.n516 66.2847
R2798 vdd.n2841 vdd.n516 66.2847
R2799 vdd.n2835 vdd.n516 66.2847
R2800 vdd.n2833 vdd.n516 66.2847
R2801 vdd.n2827 vdd.n516 66.2847
R2802 vdd.n2825 vdd.n516 66.2847
R2803 vdd.n2819 vdd.n516 66.2847
R2804 vdd.n607 vdd.n516 66.2847
R2805 vdd.n609 vdd.n516 66.2847
R2806 vdd.n3018 vdd.n351 66.2847
R2807 vdd.n3027 vdd.n351 66.2847
R2808 vdd.n461 vdd.n351 66.2847
R2809 vdd.n3034 vdd.n351 66.2847
R2810 vdd.n454 vdd.n351 66.2847
R2811 vdd.n3041 vdd.n351 66.2847
R2812 vdd.n447 vdd.n351 66.2847
R2813 vdd.n3048 vdd.n351 66.2847
R2814 vdd.n440 vdd.n351 66.2847
R2815 vdd.n3055 vdd.n351 66.2847
R2816 vdd.n434 vdd.n351 66.2847
R2817 vdd.n429 vdd.n351 66.2847
R2818 vdd.n3066 vdd.n351 66.2847
R2819 vdd.n421 vdd.n351 66.2847
R2820 vdd.n3073 vdd.n351 66.2847
R2821 vdd.n414 vdd.n351 66.2847
R2822 vdd.n3080 vdd.n351 66.2847
R2823 vdd.n407 vdd.n351 66.2847
R2824 vdd.n3087 vdd.n351 66.2847
R2825 vdd.n400 vdd.n351 66.2847
R2826 vdd.n3094 vdd.n351 66.2847
R2827 vdd.n394 vdd.n351 66.2847
R2828 vdd.n389 vdd.n351 66.2847
R2829 vdd.n3105 vdd.n351 66.2847
R2830 vdd.n381 vdd.n351 66.2847
R2831 vdd.n3112 vdd.n351 66.2847
R2832 vdd.n374 vdd.n351 66.2847
R2833 vdd.n3119 vdd.n351 66.2847
R2834 vdd.n367 vdd.n351 66.2847
R2835 vdd.n3126 vdd.n351 66.2847
R2836 vdd.n3129 vdd.n351 66.2847
R2837 vdd.n355 vdd.n351 66.2847
R2838 vdd.n356 vdd.n355 52.4337
R2839 vdd.n3129 vdd.n3128 52.4337
R2840 vdd.n3126 vdd.n3125 52.4337
R2841 vdd.n3121 vdd.n367 52.4337
R2842 vdd.n3119 vdd.n3118 52.4337
R2843 vdd.n3114 vdd.n374 52.4337
R2844 vdd.n3112 vdd.n3111 52.4337
R2845 vdd.n3107 vdd.n381 52.4337
R2846 vdd.n3105 vdd.n3104 52.4337
R2847 vdd.n390 vdd.n389 52.4337
R2848 vdd.n3096 vdd.n394 52.4337
R2849 vdd.n3094 vdd.n3093 52.4337
R2850 vdd.n3089 vdd.n400 52.4337
R2851 vdd.n3087 vdd.n3086 52.4337
R2852 vdd.n3082 vdd.n407 52.4337
R2853 vdd.n3080 vdd.n3079 52.4337
R2854 vdd.n3075 vdd.n414 52.4337
R2855 vdd.n3073 vdd.n3072 52.4337
R2856 vdd.n3068 vdd.n421 52.4337
R2857 vdd.n3066 vdd.n3065 52.4337
R2858 vdd.n430 vdd.n429 52.4337
R2859 vdd.n3057 vdd.n434 52.4337
R2860 vdd.n3055 vdd.n3054 52.4337
R2861 vdd.n3050 vdd.n440 52.4337
R2862 vdd.n3048 vdd.n3047 52.4337
R2863 vdd.n3043 vdd.n447 52.4337
R2864 vdd.n3041 vdd.n3040 52.4337
R2865 vdd.n3036 vdd.n454 52.4337
R2866 vdd.n3034 vdd.n3033 52.4337
R2867 vdd.n3029 vdd.n461 52.4337
R2868 vdd.n3027 vdd.n3026 52.4337
R2869 vdd.n3019 vdd.n3018 52.4337
R2870 vdd.n2932 vdd.n517 52.4337
R2871 vdd.n2930 vdd.n520 52.4337
R2872 vdd.n2926 vdd.n523 52.4337
R2873 vdd.n2922 vdd.n2921 52.4337
R2874 vdd.n2915 vdd.n526 52.4337
R2875 vdd.n2914 vdd.n2913 52.4337
R2876 vdd.n2907 vdd.n532 52.4337
R2877 vdd.n2906 vdd.n2905 52.4337
R2878 vdd.n2899 vdd.n538 52.4337
R2879 vdd.n2898 vdd.n2897 52.4337
R2880 vdd.n2891 vdd.n546 52.4337
R2881 vdd.n2890 vdd.n2889 52.4337
R2882 vdd.n2883 vdd.n552 52.4337
R2883 vdd.n2882 vdd.n2881 52.4337
R2884 vdd.n2875 vdd.n558 52.4337
R2885 vdd.n2874 vdd.n2873 52.4337
R2886 vdd.n2867 vdd.n564 52.4337
R2887 vdd.n2866 vdd.n2865 52.4337
R2888 vdd.n2859 vdd.n570 52.4337
R2889 vdd.n2858 vdd.n2857 52.4337
R2890 vdd.n584 vdd.n576 52.4337
R2891 vdd.n2849 vdd.n2848 52.4337
R2892 vdd.n2846 vdd.n586 52.4337
R2893 vdd.n2842 vdd.n2841 52.4337
R2894 vdd.n2835 vdd.n590 52.4337
R2895 vdd.n2834 vdd.n2833 52.4337
R2896 vdd.n2827 vdd.n596 52.4337
R2897 vdd.n2826 vdd.n2825 52.4337
R2898 vdd.n2819 vdd.n602 52.4337
R2899 vdd.n2818 vdd.n607 52.4337
R2900 vdd.n2814 vdd.n609 52.4337
R2901 vdd.n2034 vdd.n1614 52.4337
R2902 vdd.n2032 vdd.n2031 52.4337
R2903 vdd.n1621 vdd.n1620 52.4337
R2904 vdd.n1810 vdd.n1809 52.4337
R2905 vdd.n1807 vdd.n1806 52.4337
R2906 vdd.n1802 vdd.n1629 52.4337
R2907 vdd.n1800 vdd.n1799 52.4337
R2908 vdd.n1795 vdd.n1636 52.4337
R2909 vdd.n1793 vdd.n1792 52.4337
R2910 vdd.n1645 vdd.n1644 52.4337
R2911 vdd.n1784 vdd.n1649 52.4337
R2912 vdd.n1782 vdd.n1781 52.4337
R2913 vdd.n1777 vdd.n1655 52.4337
R2914 vdd.n1775 vdd.n1774 52.4337
R2915 vdd.n1770 vdd.n1662 52.4337
R2916 vdd.n1768 vdd.n1767 52.4337
R2917 vdd.n1763 vdd.n1669 52.4337
R2918 vdd.n1761 vdd.n1760 52.4337
R2919 vdd.n1756 vdd.n1676 52.4337
R2920 vdd.n1754 vdd.n1753 52.4337
R2921 vdd.n1685 vdd.n1684 52.4337
R2922 vdd.n1745 vdd.n1689 52.4337
R2923 vdd.n1743 vdd.n1742 52.4337
R2924 vdd.n1738 vdd.n1695 52.4337
R2925 vdd.n1736 vdd.n1735 52.4337
R2926 vdd.n1731 vdd.n1702 52.4337
R2927 vdd.n1729 vdd.n1728 52.4337
R2928 vdd.n1724 vdd.n1710 52.4337
R2929 vdd.n1722 vdd.n1721 52.4337
R2930 vdd.n1717 vdd.n1716 52.4337
R2931 vdd.n1712 vdd.n1711 52.4337
R2932 vdd.n2043 vdd.n898 52.4337
R2933 vdd.n986 vdd.n984 52.4337
R2934 vdd.n992 vdd.n991 52.4337
R2935 vdd.n995 vdd.n994 52.4337
R2936 vdd.n1000 vdd.n999 52.4337
R2937 vdd.n1003 vdd.n1002 52.4337
R2938 vdd.n1008 vdd.n1007 52.4337
R2939 vdd.n1011 vdd.n1010 52.4337
R2940 vdd.n1016 vdd.n1015 52.4337
R2941 vdd.n1019 vdd.n1018 52.4337
R2942 vdd.n1026 vdd.n1025 52.4337
R2943 vdd.n1029 vdd.n1028 52.4337
R2944 vdd.n1034 vdd.n1033 52.4337
R2945 vdd.n1037 vdd.n1036 52.4337
R2946 vdd.n1042 vdd.n1041 52.4337
R2947 vdd.n1045 vdd.n1044 52.4337
R2948 vdd.n1050 vdd.n1049 52.4337
R2949 vdd.n1053 vdd.n1052 52.4337
R2950 vdd.n1058 vdd.n1057 52.4337
R2951 vdd.n1061 vdd.n1060 52.4337
R2952 vdd.n1066 vdd.n1065 52.4337
R2953 vdd.n1146 vdd.n1145 52.4337
R2954 vdd.n1143 vdd.n1069 52.4337
R2955 vdd.n1075 vdd.n1074 52.4337
R2956 vdd.n1080 vdd.n1077 52.4337
R2957 vdd.n1083 vdd.n1082 52.4337
R2958 vdd.n1088 vdd.n1085 52.4337
R2959 vdd.n1091 vdd.n1090 52.4337
R2960 vdd.n1096 vdd.n1093 52.4337
R2961 vdd.n1099 vdd.n1098 52.4337
R2962 vdd.n1104 vdd.n1101 52.4337
R2963 vdd.n1107 vdd.n1106 52.4337
R2964 vdd.n987 vdd.n986 52.4337
R2965 vdd.n993 vdd.n992 52.4337
R2966 vdd.n996 vdd.n995 52.4337
R2967 vdd.n1001 vdd.n1000 52.4337
R2968 vdd.n1004 vdd.n1003 52.4337
R2969 vdd.n1009 vdd.n1008 52.4337
R2970 vdd.n1012 vdd.n1011 52.4337
R2971 vdd.n1017 vdd.n1016 52.4337
R2972 vdd.n1020 vdd.n1019 52.4337
R2973 vdd.n1027 vdd.n1026 52.4337
R2974 vdd.n1030 vdd.n1029 52.4337
R2975 vdd.n1035 vdd.n1034 52.4337
R2976 vdd.n1038 vdd.n1037 52.4337
R2977 vdd.n1043 vdd.n1042 52.4337
R2978 vdd.n1046 vdd.n1045 52.4337
R2979 vdd.n1051 vdd.n1050 52.4337
R2980 vdd.n1054 vdd.n1053 52.4337
R2981 vdd.n1059 vdd.n1058 52.4337
R2982 vdd.n1062 vdd.n1061 52.4337
R2983 vdd.n1067 vdd.n1066 52.4337
R2984 vdd.n1145 vdd.n1144 52.4337
R2985 vdd.n1073 vdd.n1069 52.4337
R2986 vdd.n1076 vdd.n1075 52.4337
R2987 vdd.n1081 vdd.n1080 52.4337
R2988 vdd.n1084 vdd.n1083 52.4337
R2989 vdd.n1089 vdd.n1088 52.4337
R2990 vdd.n1092 vdd.n1091 52.4337
R2991 vdd.n1097 vdd.n1096 52.4337
R2992 vdd.n1100 vdd.n1099 52.4337
R2993 vdd.n1105 vdd.n1104 52.4337
R2994 vdd.n1108 vdd.n1107 52.4337
R2995 vdd.n898 vdd.n897 52.4337
R2996 vdd.n1713 vdd.n1712 52.4337
R2997 vdd.n1718 vdd.n1717 52.4337
R2998 vdd.n1723 vdd.n1722 52.4337
R2999 vdd.n1710 vdd.n1703 52.4337
R3000 vdd.n1730 vdd.n1729 52.4337
R3001 vdd.n1702 vdd.n1696 52.4337
R3002 vdd.n1737 vdd.n1736 52.4337
R3003 vdd.n1695 vdd.n1690 52.4337
R3004 vdd.n1744 vdd.n1743 52.4337
R3005 vdd.n1689 vdd.n1688 52.4337
R3006 vdd.n1684 vdd.n1677 52.4337
R3007 vdd.n1755 vdd.n1754 52.4337
R3008 vdd.n1676 vdd.n1670 52.4337
R3009 vdd.n1762 vdd.n1761 52.4337
R3010 vdd.n1669 vdd.n1663 52.4337
R3011 vdd.n1769 vdd.n1768 52.4337
R3012 vdd.n1662 vdd.n1656 52.4337
R3013 vdd.n1776 vdd.n1775 52.4337
R3014 vdd.n1655 vdd.n1650 52.4337
R3015 vdd.n1783 vdd.n1782 52.4337
R3016 vdd.n1649 vdd.n1648 52.4337
R3017 vdd.n1644 vdd.n1637 52.4337
R3018 vdd.n1794 vdd.n1793 52.4337
R3019 vdd.n1636 vdd.n1630 52.4337
R3020 vdd.n1801 vdd.n1800 52.4337
R3021 vdd.n1629 vdd.n1623 52.4337
R3022 vdd.n1808 vdd.n1807 52.4337
R3023 vdd.n1811 vdd.n1810 52.4337
R3024 vdd.n1620 vdd.n1615 52.4337
R3025 vdd.n2033 vdd.n2032 52.4337
R3026 vdd.n1614 vdd.n903 52.4337
R3027 vdd.n2933 vdd.n2932 52.4337
R3028 vdd.n2927 vdd.n520 52.4337
R3029 vdd.n2923 vdd.n523 52.4337
R3030 vdd.n2921 vdd.n2920 52.4337
R3031 vdd.n2916 vdd.n2915 52.4337
R3032 vdd.n2913 vdd.n2912 52.4337
R3033 vdd.n2908 vdd.n2907 52.4337
R3034 vdd.n2905 vdd.n2904 52.4337
R3035 vdd.n2900 vdd.n2899 52.4337
R3036 vdd.n2897 vdd.n2896 52.4337
R3037 vdd.n2892 vdd.n2891 52.4337
R3038 vdd.n2889 vdd.n2888 52.4337
R3039 vdd.n2884 vdd.n2883 52.4337
R3040 vdd.n2881 vdd.n2880 52.4337
R3041 vdd.n2876 vdd.n2875 52.4337
R3042 vdd.n2873 vdd.n2872 52.4337
R3043 vdd.n2868 vdd.n2867 52.4337
R3044 vdd.n2865 vdd.n2864 52.4337
R3045 vdd.n2860 vdd.n2859 52.4337
R3046 vdd.n2857 vdd.n2856 52.4337
R3047 vdd.n585 vdd.n584 52.4337
R3048 vdd.n2848 vdd.n2847 52.4337
R3049 vdd.n2843 vdd.n586 52.4337
R3050 vdd.n2841 vdd.n2840 52.4337
R3051 vdd.n2836 vdd.n2835 52.4337
R3052 vdd.n2833 vdd.n2832 52.4337
R3053 vdd.n2828 vdd.n2827 52.4337
R3054 vdd.n2825 vdd.n2824 52.4337
R3055 vdd.n2820 vdd.n2819 52.4337
R3056 vdd.n2815 vdd.n607 52.4337
R3057 vdd.n2811 vdd.n609 52.4337
R3058 vdd.n3018 vdd.n462 52.4337
R3059 vdd.n3028 vdd.n3027 52.4337
R3060 vdd.n461 vdd.n455 52.4337
R3061 vdd.n3035 vdd.n3034 52.4337
R3062 vdd.n454 vdd.n448 52.4337
R3063 vdd.n3042 vdd.n3041 52.4337
R3064 vdd.n447 vdd.n441 52.4337
R3065 vdd.n3049 vdd.n3048 52.4337
R3066 vdd.n440 vdd.n435 52.4337
R3067 vdd.n3056 vdd.n3055 52.4337
R3068 vdd.n434 vdd.n433 52.4337
R3069 vdd.n429 vdd.n422 52.4337
R3070 vdd.n3067 vdd.n3066 52.4337
R3071 vdd.n421 vdd.n415 52.4337
R3072 vdd.n3074 vdd.n3073 52.4337
R3073 vdd.n414 vdd.n408 52.4337
R3074 vdd.n3081 vdd.n3080 52.4337
R3075 vdd.n407 vdd.n401 52.4337
R3076 vdd.n3088 vdd.n3087 52.4337
R3077 vdd.n400 vdd.n395 52.4337
R3078 vdd.n3095 vdd.n3094 52.4337
R3079 vdd.n394 vdd.n393 52.4337
R3080 vdd.n389 vdd.n382 52.4337
R3081 vdd.n3106 vdd.n3105 52.4337
R3082 vdd.n381 vdd.n375 52.4337
R3083 vdd.n3113 vdd.n3112 52.4337
R3084 vdd.n374 vdd.n368 52.4337
R3085 vdd.n3120 vdd.n3119 52.4337
R3086 vdd.n367 vdd.n360 52.4337
R3087 vdd.n3127 vdd.n3126 52.4337
R3088 vdd.n3130 vdd.n3129 52.4337
R3089 vdd.n355 vdd.n352 52.4337
R3090 vdd.t111 vdd.t228 51.4683
R3091 vdd.n258 vdd.n256 42.0461
R3092 vdd.n164 vdd.n162 42.0461
R3093 vdd.n71 vdd.n69 42.0461
R3094 vdd.n1504 vdd.n1502 42.0461
R3095 vdd.n1410 vdd.n1408 42.0461
R3096 vdd.n1317 vdd.n1315 42.0461
R3097 vdd.n308 vdd.n307 41.6884
R3098 vdd.n214 vdd.n213 41.6884
R3099 vdd.n121 vdd.n120 41.6884
R3100 vdd.n1554 vdd.n1553 41.6884
R3101 vdd.n1460 vdd.n1459 41.6884
R3102 vdd.n1367 vdd.n1366 41.6884
R3103 vdd.n1112 vdd.n1111 41.1157
R3104 vdd.n1149 vdd.n1148 41.1157
R3105 vdd.n1023 vdd.n1022 41.1157
R3106 vdd.n3023 vdd.n3022 41.1157
R3107 vdd.n3062 vdd.n428 41.1157
R3108 vdd.n3101 vdd.n388 41.1157
R3109 vdd.n2765 vdd.n2764 39.2114
R3110 vdd.n2762 vdd.n2761 39.2114
R3111 vdd.n2757 vdd.n641 39.2114
R3112 vdd.n2755 vdd.n2754 39.2114
R3113 vdd.n2750 vdd.n644 39.2114
R3114 vdd.n2748 vdd.n2747 39.2114
R3115 vdd.n2743 vdd.n647 39.2114
R3116 vdd.n2741 vdd.n2740 39.2114
R3117 vdd.n2735 vdd.n650 39.2114
R3118 vdd.n2733 vdd.n2732 39.2114
R3119 vdd.n2728 vdd.n653 39.2114
R3120 vdd.n2726 vdd.n2725 39.2114
R3121 vdd.n2721 vdd.n656 39.2114
R3122 vdd.n2719 vdd.n2718 39.2114
R3123 vdd.n2714 vdd.n659 39.2114
R3124 vdd.n2712 vdd.n2711 39.2114
R3125 vdd.n2707 vdd.n2706 39.2114
R3126 vdd.n2568 vdd.n741 39.2114
R3127 vdd.n2563 vdd.n2317 39.2114
R3128 vdd.n2560 vdd.n2318 39.2114
R3129 vdd.n2556 vdd.n2319 39.2114
R3130 vdd.n2552 vdd.n2320 39.2114
R3131 vdd.n2548 vdd.n2321 39.2114
R3132 vdd.n2544 vdd.n2322 39.2114
R3133 vdd.n2540 vdd.n2323 39.2114
R3134 vdd.n2536 vdd.n2324 39.2114
R3135 vdd.n2532 vdd.n2325 39.2114
R3136 vdd.n2528 vdd.n2326 39.2114
R3137 vdd.n2524 vdd.n2327 39.2114
R3138 vdd.n2520 vdd.n2328 39.2114
R3139 vdd.n2516 vdd.n2329 39.2114
R3140 vdd.n2512 vdd.n2330 39.2114
R3141 vdd.n2508 vdd.n2331 39.2114
R3142 vdd.n2503 vdd.n2332 39.2114
R3143 vdd.n2311 vdd.n781 39.2114
R3144 vdd.n2307 vdd.n780 39.2114
R3145 vdd.n2303 vdd.n779 39.2114
R3146 vdd.n2299 vdd.n778 39.2114
R3147 vdd.n2295 vdd.n777 39.2114
R3148 vdd.n2291 vdd.n776 39.2114
R3149 vdd.n2287 vdd.n775 39.2114
R3150 vdd.n2283 vdd.n774 39.2114
R3151 vdd.n2279 vdd.n773 39.2114
R3152 vdd.n2275 vdd.n772 39.2114
R3153 vdd.n2271 vdd.n771 39.2114
R3154 vdd.n2267 vdd.n770 39.2114
R3155 vdd.n2263 vdd.n769 39.2114
R3156 vdd.n2259 vdd.n768 39.2114
R3157 vdd.n2255 vdd.n767 39.2114
R3158 vdd.n2250 vdd.n766 39.2114
R3159 vdd.n2246 vdd.n765 39.2114
R3160 vdd.n1822 vdd.n876 39.2114
R3161 vdd.n1828 vdd.n1827 39.2114
R3162 vdd.n1831 vdd.n1830 39.2114
R3163 vdd.n1836 vdd.n1835 39.2114
R3164 vdd.n1839 vdd.n1838 39.2114
R3165 vdd.n1844 vdd.n1843 39.2114
R3166 vdd.n1847 vdd.n1846 39.2114
R3167 vdd.n1852 vdd.n1851 39.2114
R3168 vdd.n2023 vdd.n1854 39.2114
R3169 vdd.n2022 vdd.n2021 39.2114
R3170 vdd.n2015 vdd.n1856 39.2114
R3171 vdd.n2014 vdd.n2013 39.2114
R3172 vdd.n2007 vdd.n1858 39.2114
R3173 vdd.n2006 vdd.n2005 39.2114
R3174 vdd.n1999 vdd.n1860 39.2114
R3175 vdd.n1998 vdd.n1997 39.2114
R3176 vdd.n1991 vdd.n1862 39.2114
R3177 vdd.n2684 vdd.n2683 39.2114
R3178 vdd.n2679 vdd.n2651 39.2114
R3179 vdd.n2677 vdd.n2676 39.2114
R3180 vdd.n2672 vdd.n2654 39.2114
R3181 vdd.n2670 vdd.n2669 39.2114
R3182 vdd.n2665 vdd.n2657 39.2114
R3183 vdd.n2663 vdd.n2662 39.2114
R3184 vdd.n2658 vdd.n612 39.2114
R3185 vdd.n2802 vdd.n2801 39.2114
R3186 vdd.n2799 vdd.n2798 39.2114
R3187 vdd.n2794 vdd.n617 39.2114
R3188 vdd.n2792 vdd.n2791 39.2114
R3189 vdd.n2787 vdd.n620 39.2114
R3190 vdd.n2785 vdd.n2784 39.2114
R3191 vdd.n2780 vdd.n623 39.2114
R3192 vdd.n2778 vdd.n2777 39.2114
R3193 vdd.n2773 vdd.n629 39.2114
R3194 vdd.n2570 vdd.n744 39.2114
R3195 vdd.n2333 vdd.n746 39.2114
R3196 vdd.n2359 vdd.n2334 39.2114
R3197 vdd.n2363 vdd.n2335 39.2114
R3198 vdd.n2367 vdd.n2336 39.2114
R3199 vdd.n2371 vdd.n2337 39.2114
R3200 vdd.n2375 vdd.n2338 39.2114
R3201 vdd.n2379 vdd.n2339 39.2114
R3202 vdd.n2383 vdd.n2340 39.2114
R3203 vdd.n2387 vdd.n2341 39.2114
R3204 vdd.n2391 vdd.n2342 39.2114
R3205 vdd.n2395 vdd.n2343 39.2114
R3206 vdd.n2399 vdd.n2344 39.2114
R3207 vdd.n2403 vdd.n2345 39.2114
R3208 vdd.n2407 vdd.n2346 39.2114
R3209 vdd.n2411 vdd.n2347 39.2114
R3210 vdd.n2415 vdd.n2348 39.2114
R3211 vdd.n2571 vdd.n2570 39.2114
R3212 vdd.n2358 vdd.n2333 39.2114
R3213 vdd.n2362 vdd.n2334 39.2114
R3214 vdd.n2366 vdd.n2335 39.2114
R3215 vdd.n2370 vdd.n2336 39.2114
R3216 vdd.n2374 vdd.n2337 39.2114
R3217 vdd.n2378 vdd.n2338 39.2114
R3218 vdd.n2382 vdd.n2339 39.2114
R3219 vdd.n2386 vdd.n2340 39.2114
R3220 vdd.n2390 vdd.n2341 39.2114
R3221 vdd.n2394 vdd.n2342 39.2114
R3222 vdd.n2398 vdd.n2343 39.2114
R3223 vdd.n2402 vdd.n2344 39.2114
R3224 vdd.n2406 vdd.n2345 39.2114
R3225 vdd.n2410 vdd.n2346 39.2114
R3226 vdd.n2414 vdd.n2347 39.2114
R3227 vdd.n2417 vdd.n2348 39.2114
R3228 vdd.n629 vdd.n624 39.2114
R3229 vdd.n2779 vdd.n2778 39.2114
R3230 vdd.n623 vdd.n621 39.2114
R3231 vdd.n2786 vdd.n2785 39.2114
R3232 vdd.n620 vdd.n618 39.2114
R3233 vdd.n2793 vdd.n2792 39.2114
R3234 vdd.n617 vdd.n615 39.2114
R3235 vdd.n2800 vdd.n2799 39.2114
R3236 vdd.n2803 vdd.n2802 39.2114
R3237 vdd.n2659 vdd.n2658 39.2114
R3238 vdd.n2664 vdd.n2663 39.2114
R3239 vdd.n2657 vdd.n2655 39.2114
R3240 vdd.n2671 vdd.n2670 39.2114
R3241 vdd.n2654 vdd.n2652 39.2114
R3242 vdd.n2678 vdd.n2677 39.2114
R3243 vdd.n2651 vdd.n2649 39.2114
R3244 vdd.n2685 vdd.n2684 39.2114
R3245 vdd.n1823 vdd.n1822 39.2114
R3246 vdd.n1829 vdd.n1828 39.2114
R3247 vdd.n1830 vdd.n1819 39.2114
R3248 vdd.n1837 vdd.n1836 39.2114
R3249 vdd.n1838 vdd.n1817 39.2114
R3250 vdd.n1845 vdd.n1844 39.2114
R3251 vdd.n1846 vdd.n1815 39.2114
R3252 vdd.n1853 vdd.n1852 39.2114
R3253 vdd.n2024 vdd.n2023 39.2114
R3254 vdd.n2021 vdd.n2020 39.2114
R3255 vdd.n2016 vdd.n2015 39.2114
R3256 vdd.n2013 vdd.n2012 39.2114
R3257 vdd.n2008 vdd.n2007 39.2114
R3258 vdd.n2005 vdd.n2004 39.2114
R3259 vdd.n2000 vdd.n1999 39.2114
R3260 vdd.n1997 vdd.n1996 39.2114
R3261 vdd.n1992 vdd.n1991 39.2114
R3262 vdd.n2249 vdd.n765 39.2114
R3263 vdd.n2254 vdd.n766 39.2114
R3264 vdd.n2258 vdd.n767 39.2114
R3265 vdd.n2262 vdd.n768 39.2114
R3266 vdd.n2266 vdd.n769 39.2114
R3267 vdd.n2270 vdd.n770 39.2114
R3268 vdd.n2274 vdd.n771 39.2114
R3269 vdd.n2278 vdd.n772 39.2114
R3270 vdd.n2282 vdd.n773 39.2114
R3271 vdd.n2286 vdd.n774 39.2114
R3272 vdd.n2290 vdd.n775 39.2114
R3273 vdd.n2294 vdd.n776 39.2114
R3274 vdd.n2298 vdd.n777 39.2114
R3275 vdd.n2302 vdd.n778 39.2114
R3276 vdd.n2306 vdd.n779 39.2114
R3277 vdd.n2310 vdd.n780 39.2114
R3278 vdd.n783 vdd.n781 39.2114
R3279 vdd.n2568 vdd.n2567 39.2114
R3280 vdd.n2561 vdd.n2317 39.2114
R3281 vdd.n2557 vdd.n2318 39.2114
R3282 vdd.n2553 vdd.n2319 39.2114
R3283 vdd.n2549 vdd.n2320 39.2114
R3284 vdd.n2545 vdd.n2321 39.2114
R3285 vdd.n2541 vdd.n2322 39.2114
R3286 vdd.n2537 vdd.n2323 39.2114
R3287 vdd.n2533 vdd.n2324 39.2114
R3288 vdd.n2529 vdd.n2325 39.2114
R3289 vdd.n2525 vdd.n2326 39.2114
R3290 vdd.n2521 vdd.n2327 39.2114
R3291 vdd.n2517 vdd.n2328 39.2114
R3292 vdd.n2513 vdd.n2329 39.2114
R3293 vdd.n2509 vdd.n2330 39.2114
R3294 vdd.n2504 vdd.n2331 39.2114
R3295 vdd.n2500 vdd.n2332 39.2114
R3296 vdd.n2706 vdd.n660 39.2114
R3297 vdd.n2713 vdd.n2712 39.2114
R3298 vdd.n659 vdd.n657 39.2114
R3299 vdd.n2720 vdd.n2719 39.2114
R3300 vdd.n656 vdd.n654 39.2114
R3301 vdd.n2727 vdd.n2726 39.2114
R3302 vdd.n653 vdd.n651 39.2114
R3303 vdd.n2734 vdd.n2733 39.2114
R3304 vdd.n650 vdd.n648 39.2114
R3305 vdd.n2742 vdd.n2741 39.2114
R3306 vdd.n647 vdd.n645 39.2114
R3307 vdd.n2749 vdd.n2748 39.2114
R3308 vdd.n644 vdd.n642 39.2114
R3309 vdd.n2756 vdd.n2755 39.2114
R3310 vdd.n641 vdd.n639 39.2114
R3311 vdd.n2763 vdd.n2762 39.2114
R3312 vdd.n2766 vdd.n2765 39.2114
R3313 vdd.n791 vdd.n747 39.2114
R3314 vdd.n2238 vdd.n748 39.2114
R3315 vdd.n2234 vdd.n749 39.2114
R3316 vdd.n2230 vdd.n750 39.2114
R3317 vdd.n2226 vdd.n751 39.2114
R3318 vdd.n2222 vdd.n752 39.2114
R3319 vdd.n2218 vdd.n753 39.2114
R3320 vdd.n2214 vdd.n754 39.2114
R3321 vdd.n2210 vdd.n755 39.2114
R3322 vdd.n2206 vdd.n756 39.2114
R3323 vdd.n2202 vdd.n757 39.2114
R3324 vdd.n2198 vdd.n758 39.2114
R3325 vdd.n2194 vdd.n759 39.2114
R3326 vdd.n2190 vdd.n760 39.2114
R3327 vdd.n2186 vdd.n761 39.2114
R3328 vdd.n2182 vdd.n762 39.2114
R3329 vdd.n2178 vdd.n763 39.2114
R3330 vdd.n2081 vdd.n880 39.2114
R3331 vdd.n2080 vdd.n2079 39.2114
R3332 vdd.n2073 vdd.n882 39.2114
R3333 vdd.n2072 vdd.n2071 39.2114
R3334 vdd.n2065 vdd.n884 39.2114
R3335 vdd.n2064 vdd.n2063 39.2114
R3336 vdd.n2057 vdd.n886 39.2114
R3337 vdd.n2056 vdd.n2055 39.2114
R3338 vdd.n889 vdd.n888 39.2114
R3339 vdd.n1897 vdd.n1896 39.2114
R3340 vdd.n1902 vdd.n1901 39.2114
R3341 vdd.n1905 vdd.n1904 39.2114
R3342 vdd.n1910 vdd.n1909 39.2114
R3343 vdd.n1913 vdd.n1912 39.2114
R3344 vdd.n1918 vdd.n1917 39.2114
R3345 vdd.n1921 vdd.n1920 39.2114
R3346 vdd.n1927 vdd.n1926 39.2114
R3347 vdd.n2175 vdd.n763 39.2114
R3348 vdd.n2179 vdd.n762 39.2114
R3349 vdd.n2183 vdd.n761 39.2114
R3350 vdd.n2187 vdd.n760 39.2114
R3351 vdd.n2191 vdd.n759 39.2114
R3352 vdd.n2195 vdd.n758 39.2114
R3353 vdd.n2199 vdd.n757 39.2114
R3354 vdd.n2203 vdd.n756 39.2114
R3355 vdd.n2207 vdd.n755 39.2114
R3356 vdd.n2211 vdd.n754 39.2114
R3357 vdd.n2215 vdd.n753 39.2114
R3358 vdd.n2219 vdd.n752 39.2114
R3359 vdd.n2223 vdd.n751 39.2114
R3360 vdd.n2227 vdd.n750 39.2114
R3361 vdd.n2231 vdd.n749 39.2114
R3362 vdd.n2235 vdd.n748 39.2114
R3363 vdd.n2239 vdd.n747 39.2114
R3364 vdd.n2082 vdd.n2081 39.2114
R3365 vdd.n2079 vdd.n2078 39.2114
R3366 vdd.n2074 vdd.n2073 39.2114
R3367 vdd.n2071 vdd.n2070 39.2114
R3368 vdd.n2066 vdd.n2065 39.2114
R3369 vdd.n2063 vdd.n2062 39.2114
R3370 vdd.n2058 vdd.n2057 39.2114
R3371 vdd.n2055 vdd.n2054 39.2114
R3372 vdd.n890 vdd.n889 39.2114
R3373 vdd.n1898 vdd.n1897 39.2114
R3374 vdd.n1903 vdd.n1902 39.2114
R3375 vdd.n1904 vdd.n1894 39.2114
R3376 vdd.n1911 vdd.n1910 39.2114
R3377 vdd.n1912 vdd.n1892 39.2114
R3378 vdd.n1919 vdd.n1918 39.2114
R3379 vdd.n1920 vdd.n1888 39.2114
R3380 vdd.n1928 vdd.n1927 39.2114
R3381 vdd.n2047 vdd.n2046 37.2369
R3382 vdd.n1750 vdd.n1683 37.2369
R3383 vdd.n1789 vdd.n1643 37.2369
R3384 vdd.n2854 vdd.n581 37.2369
R3385 vdd.n545 vdd.n544 37.2369
R3386 vdd.n2810 vdd.n2809 37.2369
R3387 vdd.n2089 vdd.n875 31.6883
R3388 vdd.n2314 vdd.n784 31.6883
R3389 vdd.n2247 vdd.n787 31.6883
R3390 vdd.n1993 vdd.n1990 31.6883
R3391 vdd.n2501 vdd.n2499 31.6883
R3392 vdd.n2708 vdd.n2705 31.6883
R3393 vdd.n2578 vdd.n740 31.6883
R3394 vdd.n2769 vdd.n2768 31.6883
R3395 vdd.n2688 vdd.n2687 31.6883
R3396 vdd.n2774 vdd.n628 31.6883
R3397 vdd.n2420 vdd.n2419 31.6883
R3398 vdd.n2574 vdd.n2573 31.6883
R3399 vdd.n2085 vdd.n2084 31.6883
R3400 vdd.n2242 vdd.n2241 31.6883
R3401 vdd.n2174 vdd.n2173 31.6883
R3402 vdd.n1931 vdd.n1930 31.6883
R3403 vdd.n1924 vdd.n1890 30.449
R3404 vdd.n795 vdd.n794 30.449
R3405 vdd.n1865 vdd.n1864 30.449
R3406 vdd.n2252 vdd.n786 30.449
R3407 vdd.n2356 vdd.n2355 30.449
R3408 vdd.n663 vdd.n662 30.449
R3409 vdd.n2506 vdd.n2352 30.449
R3410 vdd.n627 vdd.n626 30.449
R3411 vdd.n1215 vdd.n982 20.633
R3412 vdd.n2041 vdd.n901 20.633
R3413 vdd.n2940 vdd.n516 20.633
R3414 vdd.n3138 vdd.n351 20.633
R3415 vdd.n1217 vdd.n979 19.3944
R3416 vdd.n1221 vdd.n979 19.3944
R3417 vdd.n1221 vdd.n970 19.3944
R3418 vdd.n1233 vdd.n970 19.3944
R3419 vdd.n1233 vdd.n968 19.3944
R3420 vdd.n1237 vdd.n968 19.3944
R3421 vdd.n1237 vdd.n957 19.3944
R3422 vdd.n1249 vdd.n957 19.3944
R3423 vdd.n1249 vdd.n955 19.3944
R3424 vdd.n1253 vdd.n955 19.3944
R3425 vdd.n1253 vdd.n946 19.3944
R3426 vdd.n1266 vdd.n946 19.3944
R3427 vdd.n1266 vdd.n944 19.3944
R3428 vdd.n1270 vdd.n944 19.3944
R3429 vdd.n1270 vdd.n935 19.3944
R3430 vdd.n1564 vdd.n935 19.3944
R3431 vdd.n1564 vdd.n933 19.3944
R3432 vdd.n1568 vdd.n933 19.3944
R3433 vdd.n1568 vdd.n923 19.3944
R3434 vdd.n1581 vdd.n923 19.3944
R3435 vdd.n1581 vdd.n921 19.3944
R3436 vdd.n1585 vdd.n921 19.3944
R3437 vdd.n1585 vdd.n913 19.3944
R3438 vdd.n1598 vdd.n913 19.3944
R3439 vdd.n1598 vdd.n910 19.3944
R3440 vdd.n1604 vdd.n910 19.3944
R3441 vdd.n1604 vdd.n911 19.3944
R3442 vdd.n911 vdd.n900 19.3944
R3443 vdd.n1142 vdd.n1068 19.3944
R3444 vdd.n1142 vdd.n1070 19.3944
R3445 vdd.n1138 vdd.n1070 19.3944
R3446 vdd.n1138 vdd.n1137 19.3944
R3447 vdd.n1137 vdd.n1136 19.3944
R3448 vdd.n1136 vdd.n1078 19.3944
R3449 vdd.n1132 vdd.n1078 19.3944
R3450 vdd.n1132 vdd.n1131 19.3944
R3451 vdd.n1131 vdd.n1130 19.3944
R3452 vdd.n1130 vdd.n1086 19.3944
R3453 vdd.n1126 vdd.n1086 19.3944
R3454 vdd.n1126 vdd.n1125 19.3944
R3455 vdd.n1125 vdd.n1124 19.3944
R3456 vdd.n1124 vdd.n1094 19.3944
R3457 vdd.n1120 vdd.n1094 19.3944
R3458 vdd.n1120 vdd.n1119 19.3944
R3459 vdd.n1119 vdd.n1118 19.3944
R3460 vdd.n1118 vdd.n1102 19.3944
R3461 vdd.n1114 vdd.n1102 19.3944
R3462 vdd.n1114 vdd.n1113 19.3944
R3463 vdd.n1180 vdd.n1179 19.3944
R3464 vdd.n1179 vdd.n1178 19.3944
R3465 vdd.n1178 vdd.n1031 19.3944
R3466 vdd.n1174 vdd.n1031 19.3944
R3467 vdd.n1174 vdd.n1173 19.3944
R3468 vdd.n1173 vdd.n1172 19.3944
R3469 vdd.n1172 vdd.n1039 19.3944
R3470 vdd.n1168 vdd.n1039 19.3944
R3471 vdd.n1168 vdd.n1167 19.3944
R3472 vdd.n1167 vdd.n1166 19.3944
R3473 vdd.n1166 vdd.n1047 19.3944
R3474 vdd.n1162 vdd.n1047 19.3944
R3475 vdd.n1162 vdd.n1161 19.3944
R3476 vdd.n1161 vdd.n1160 19.3944
R3477 vdd.n1160 vdd.n1055 19.3944
R3478 vdd.n1156 vdd.n1055 19.3944
R3479 vdd.n1156 vdd.n1155 19.3944
R3480 vdd.n1155 vdd.n1154 19.3944
R3481 vdd.n1154 vdd.n1063 19.3944
R3482 vdd.n1150 vdd.n1063 19.3944
R3483 vdd.n1210 vdd.n1209 19.3944
R3484 vdd.n1209 vdd.n1208 19.3944
R3485 vdd.n1208 vdd.n989 19.3944
R3486 vdd.n1204 vdd.n989 19.3944
R3487 vdd.n1204 vdd.n1203 19.3944
R3488 vdd.n1203 vdd.n1202 19.3944
R3489 vdd.n1202 vdd.n997 19.3944
R3490 vdd.n1198 vdd.n997 19.3944
R3491 vdd.n1198 vdd.n1197 19.3944
R3492 vdd.n1197 vdd.n1196 19.3944
R3493 vdd.n1196 vdd.n1005 19.3944
R3494 vdd.n1192 vdd.n1005 19.3944
R3495 vdd.n1192 vdd.n1191 19.3944
R3496 vdd.n1191 vdd.n1190 19.3944
R3497 vdd.n1190 vdd.n1013 19.3944
R3498 vdd.n1186 vdd.n1013 19.3944
R3499 vdd.n1186 vdd.n1185 19.3944
R3500 vdd.n1185 vdd.n1184 19.3944
R3501 vdd.n1746 vdd.n1681 19.3944
R3502 vdd.n1746 vdd.n1687 19.3944
R3503 vdd.n1741 vdd.n1687 19.3944
R3504 vdd.n1741 vdd.n1740 19.3944
R3505 vdd.n1740 vdd.n1739 19.3944
R3506 vdd.n1739 vdd.n1694 19.3944
R3507 vdd.n1734 vdd.n1694 19.3944
R3508 vdd.n1734 vdd.n1733 19.3944
R3509 vdd.n1733 vdd.n1732 19.3944
R3510 vdd.n1732 vdd.n1701 19.3944
R3511 vdd.n1727 vdd.n1701 19.3944
R3512 vdd.n1727 vdd.n1726 19.3944
R3513 vdd.n1726 vdd.n1725 19.3944
R3514 vdd.n1725 vdd.n1709 19.3944
R3515 vdd.n1720 vdd.n1709 19.3944
R3516 vdd.n1720 vdd.n1719 19.3944
R3517 vdd.n1715 vdd.n1714 19.3944
R3518 vdd.n2048 vdd.n896 19.3944
R3519 vdd.n1785 vdd.n1641 19.3944
R3520 vdd.n1785 vdd.n1647 19.3944
R3521 vdd.n1780 vdd.n1647 19.3944
R3522 vdd.n1780 vdd.n1779 19.3944
R3523 vdd.n1779 vdd.n1778 19.3944
R3524 vdd.n1778 vdd.n1654 19.3944
R3525 vdd.n1773 vdd.n1654 19.3944
R3526 vdd.n1773 vdd.n1772 19.3944
R3527 vdd.n1772 vdd.n1771 19.3944
R3528 vdd.n1771 vdd.n1661 19.3944
R3529 vdd.n1766 vdd.n1661 19.3944
R3530 vdd.n1766 vdd.n1765 19.3944
R3531 vdd.n1765 vdd.n1764 19.3944
R3532 vdd.n1764 vdd.n1668 19.3944
R3533 vdd.n1759 vdd.n1668 19.3944
R3534 vdd.n1759 vdd.n1758 19.3944
R3535 vdd.n1758 vdd.n1757 19.3944
R3536 vdd.n1757 vdd.n1675 19.3944
R3537 vdd.n1752 vdd.n1675 19.3944
R3538 vdd.n1752 vdd.n1751 19.3944
R3539 vdd.n2036 vdd.n2035 19.3944
R3540 vdd.n2035 vdd.n1613 19.3944
R3541 vdd.n2030 vdd.n2029 19.3944
R3542 vdd.n1812 vdd.n1617 19.3944
R3543 vdd.n1812 vdd.n1619 19.3944
R3544 vdd.n1622 vdd.n1619 19.3944
R3545 vdd.n1805 vdd.n1622 19.3944
R3546 vdd.n1805 vdd.n1804 19.3944
R3547 vdd.n1804 vdd.n1803 19.3944
R3548 vdd.n1803 vdd.n1628 19.3944
R3549 vdd.n1798 vdd.n1628 19.3944
R3550 vdd.n1798 vdd.n1797 19.3944
R3551 vdd.n1797 vdd.n1796 19.3944
R3552 vdd.n1796 vdd.n1635 19.3944
R3553 vdd.n1791 vdd.n1635 19.3944
R3554 vdd.n1791 vdd.n1790 19.3944
R3555 vdd.n1213 vdd.n976 19.3944
R3556 vdd.n1225 vdd.n976 19.3944
R3557 vdd.n1225 vdd.n974 19.3944
R3558 vdd.n1229 vdd.n974 19.3944
R3559 vdd.n1229 vdd.n964 19.3944
R3560 vdd.n1241 vdd.n964 19.3944
R3561 vdd.n1241 vdd.n962 19.3944
R3562 vdd.n1245 vdd.n962 19.3944
R3563 vdd.n1245 vdd.n952 19.3944
R3564 vdd.n1258 vdd.n952 19.3944
R3565 vdd.n1258 vdd.n950 19.3944
R3566 vdd.n1262 vdd.n950 19.3944
R3567 vdd.n1262 vdd.n941 19.3944
R3568 vdd.n1274 vdd.n941 19.3944
R3569 vdd.n1274 vdd.n939 19.3944
R3570 vdd.n1560 vdd.n939 19.3944
R3571 vdd.n1560 vdd.n929 19.3944
R3572 vdd.n1573 vdd.n929 19.3944
R3573 vdd.n1573 vdd.n927 19.3944
R3574 vdd.n1577 vdd.n927 19.3944
R3575 vdd.n1577 vdd.n918 19.3944
R3576 vdd.n1590 vdd.n918 19.3944
R3577 vdd.n1590 vdd.n916 19.3944
R3578 vdd.n1594 vdd.n916 19.3944
R3579 vdd.n1594 vdd.n906 19.3944
R3580 vdd.n1609 vdd.n906 19.3944
R3581 vdd.n1609 vdd.n904 19.3944
R3582 vdd.n2039 vdd.n904 19.3944
R3583 vdd.n2942 vdd.n513 19.3944
R3584 vdd.n2946 vdd.n513 19.3944
R3585 vdd.n2946 vdd.n503 19.3944
R3586 vdd.n2958 vdd.n503 19.3944
R3587 vdd.n2958 vdd.n501 19.3944
R3588 vdd.n2962 vdd.n501 19.3944
R3589 vdd.n2962 vdd.n490 19.3944
R3590 vdd.n2974 vdd.n490 19.3944
R3591 vdd.n2974 vdd.n488 19.3944
R3592 vdd.n2978 vdd.n488 19.3944
R3593 vdd.n2978 vdd.n478 19.3944
R3594 vdd.n2991 vdd.n478 19.3944
R3595 vdd.n2991 vdd.n476 19.3944
R3596 vdd.n2995 vdd.n476 19.3944
R3597 vdd.n2996 vdd.n2995 19.3944
R3598 vdd.n2997 vdd.n2996 19.3944
R3599 vdd.n2997 vdd.n474 19.3944
R3600 vdd.n3001 vdd.n474 19.3944
R3601 vdd.n3002 vdd.n3001 19.3944
R3602 vdd.n3003 vdd.n3002 19.3944
R3603 vdd.n3003 vdd.n471 19.3944
R3604 vdd.n3007 vdd.n471 19.3944
R3605 vdd.n3008 vdd.n3007 19.3944
R3606 vdd.n3009 vdd.n3008 19.3944
R3607 vdd.n3009 vdd.n468 19.3944
R3608 vdd.n3013 vdd.n468 19.3944
R3609 vdd.n3014 vdd.n3013 19.3944
R3610 vdd.n3015 vdd.n3014 19.3944
R3611 vdd.n3058 vdd.n426 19.3944
R3612 vdd.n3058 vdd.n432 19.3944
R3613 vdd.n3053 vdd.n432 19.3944
R3614 vdd.n3053 vdd.n3052 19.3944
R3615 vdd.n3052 vdd.n3051 19.3944
R3616 vdd.n3051 vdd.n439 19.3944
R3617 vdd.n3046 vdd.n439 19.3944
R3618 vdd.n3046 vdd.n3045 19.3944
R3619 vdd.n3045 vdd.n3044 19.3944
R3620 vdd.n3044 vdd.n446 19.3944
R3621 vdd.n3039 vdd.n446 19.3944
R3622 vdd.n3039 vdd.n3038 19.3944
R3623 vdd.n3038 vdd.n3037 19.3944
R3624 vdd.n3037 vdd.n453 19.3944
R3625 vdd.n3032 vdd.n453 19.3944
R3626 vdd.n3032 vdd.n3031 19.3944
R3627 vdd.n3031 vdd.n3030 19.3944
R3628 vdd.n3030 vdd.n460 19.3944
R3629 vdd.n3025 vdd.n460 19.3944
R3630 vdd.n3025 vdd.n3024 19.3944
R3631 vdd.n3097 vdd.n386 19.3944
R3632 vdd.n3097 vdd.n392 19.3944
R3633 vdd.n3092 vdd.n392 19.3944
R3634 vdd.n3092 vdd.n3091 19.3944
R3635 vdd.n3091 vdd.n3090 19.3944
R3636 vdd.n3090 vdd.n399 19.3944
R3637 vdd.n3085 vdd.n399 19.3944
R3638 vdd.n3085 vdd.n3084 19.3944
R3639 vdd.n3084 vdd.n3083 19.3944
R3640 vdd.n3083 vdd.n406 19.3944
R3641 vdd.n3078 vdd.n406 19.3944
R3642 vdd.n3078 vdd.n3077 19.3944
R3643 vdd.n3077 vdd.n3076 19.3944
R3644 vdd.n3076 vdd.n413 19.3944
R3645 vdd.n3071 vdd.n413 19.3944
R3646 vdd.n3071 vdd.n3070 19.3944
R3647 vdd.n3070 vdd.n3069 19.3944
R3648 vdd.n3069 vdd.n420 19.3944
R3649 vdd.n3064 vdd.n420 19.3944
R3650 vdd.n3064 vdd.n3063 19.3944
R3651 vdd.n3133 vdd.n3132 19.3944
R3652 vdd.n3132 vdd.n3131 19.3944
R3653 vdd.n3131 vdd.n358 19.3944
R3654 vdd.n359 vdd.n358 19.3944
R3655 vdd.n3124 vdd.n359 19.3944
R3656 vdd.n3124 vdd.n3123 19.3944
R3657 vdd.n3123 vdd.n3122 19.3944
R3658 vdd.n3122 vdd.n366 19.3944
R3659 vdd.n3117 vdd.n366 19.3944
R3660 vdd.n3117 vdd.n3116 19.3944
R3661 vdd.n3116 vdd.n3115 19.3944
R3662 vdd.n3115 vdd.n373 19.3944
R3663 vdd.n3110 vdd.n373 19.3944
R3664 vdd.n3110 vdd.n3109 19.3944
R3665 vdd.n3109 vdd.n3108 19.3944
R3666 vdd.n3108 vdd.n380 19.3944
R3667 vdd.n3103 vdd.n380 19.3944
R3668 vdd.n3103 vdd.n3102 19.3944
R3669 vdd.n2938 vdd.n509 19.3944
R3670 vdd.n2950 vdd.n509 19.3944
R3671 vdd.n2950 vdd.n507 19.3944
R3672 vdd.n2954 vdd.n507 19.3944
R3673 vdd.n2954 vdd.n497 19.3944
R3674 vdd.n2966 vdd.n497 19.3944
R3675 vdd.n2966 vdd.n495 19.3944
R3676 vdd.n2970 vdd.n495 19.3944
R3677 vdd.n2970 vdd.n485 19.3944
R3678 vdd.n2983 vdd.n485 19.3944
R3679 vdd.n2983 vdd.n483 19.3944
R3680 vdd.n2987 vdd.n483 19.3944
R3681 vdd.n2987 vdd.n312 19.3944
R3682 vdd.n3166 vdd.n312 19.3944
R3683 vdd.n3166 vdd.n313 19.3944
R3684 vdd.n3160 vdd.n313 19.3944
R3685 vdd.n3160 vdd.n3159 19.3944
R3686 vdd.n3159 vdd.n3158 19.3944
R3687 vdd.n3158 vdd.n323 19.3944
R3688 vdd.n3152 vdd.n323 19.3944
R3689 vdd.n3152 vdd.n3151 19.3944
R3690 vdd.n3151 vdd.n3150 19.3944
R3691 vdd.n3150 vdd.n335 19.3944
R3692 vdd.n3144 vdd.n335 19.3944
R3693 vdd.n3144 vdd.n3143 19.3944
R3694 vdd.n3143 vdd.n3142 19.3944
R3695 vdd.n3142 vdd.n346 19.3944
R3696 vdd.n3136 vdd.n346 19.3944
R3697 vdd.n2895 vdd.n2894 19.3944
R3698 vdd.n2894 vdd.n2893 19.3944
R3699 vdd.n2893 vdd.n551 19.3944
R3700 vdd.n2887 vdd.n551 19.3944
R3701 vdd.n2887 vdd.n2886 19.3944
R3702 vdd.n2886 vdd.n2885 19.3944
R3703 vdd.n2885 vdd.n557 19.3944
R3704 vdd.n2879 vdd.n557 19.3944
R3705 vdd.n2879 vdd.n2878 19.3944
R3706 vdd.n2878 vdd.n2877 19.3944
R3707 vdd.n2877 vdd.n563 19.3944
R3708 vdd.n2871 vdd.n563 19.3944
R3709 vdd.n2871 vdd.n2870 19.3944
R3710 vdd.n2870 vdd.n2869 19.3944
R3711 vdd.n2869 vdd.n569 19.3944
R3712 vdd.n2863 vdd.n569 19.3944
R3713 vdd.n2863 vdd.n2862 19.3944
R3714 vdd.n2862 vdd.n2861 19.3944
R3715 vdd.n2861 vdd.n575 19.3944
R3716 vdd.n2855 vdd.n575 19.3944
R3717 vdd.n2935 vdd.n2934 19.3944
R3718 vdd.n2934 vdd.n519 19.3944
R3719 vdd.n2929 vdd.n2928 19.3944
R3720 vdd.n2925 vdd.n2924 19.3944
R3721 vdd.n2924 vdd.n525 19.3944
R3722 vdd.n2919 vdd.n525 19.3944
R3723 vdd.n2919 vdd.n2918 19.3944
R3724 vdd.n2918 vdd.n2917 19.3944
R3725 vdd.n2917 vdd.n531 19.3944
R3726 vdd.n2911 vdd.n531 19.3944
R3727 vdd.n2911 vdd.n2910 19.3944
R3728 vdd.n2910 vdd.n2909 19.3944
R3729 vdd.n2909 vdd.n537 19.3944
R3730 vdd.n2903 vdd.n537 19.3944
R3731 vdd.n2903 vdd.n2902 19.3944
R3732 vdd.n2902 vdd.n2901 19.3944
R3733 vdd.n2850 vdd.n579 19.3944
R3734 vdd.n2850 vdd.n583 19.3944
R3735 vdd.n2845 vdd.n583 19.3944
R3736 vdd.n2845 vdd.n2844 19.3944
R3737 vdd.n2844 vdd.n589 19.3944
R3738 vdd.n2839 vdd.n589 19.3944
R3739 vdd.n2839 vdd.n2838 19.3944
R3740 vdd.n2838 vdd.n2837 19.3944
R3741 vdd.n2837 vdd.n595 19.3944
R3742 vdd.n2831 vdd.n595 19.3944
R3743 vdd.n2831 vdd.n2830 19.3944
R3744 vdd.n2830 vdd.n2829 19.3944
R3745 vdd.n2829 vdd.n601 19.3944
R3746 vdd.n2823 vdd.n601 19.3944
R3747 vdd.n2823 vdd.n2822 19.3944
R3748 vdd.n2822 vdd.n2821 19.3944
R3749 vdd.n2817 vdd.n2816 19.3944
R3750 vdd.n2813 vdd.n2812 19.3944
R3751 vdd.n1149 vdd.n1068 19.0066
R3752 vdd.n1750 vdd.n1681 19.0066
R3753 vdd.n3062 vdd.n426 19.0066
R3754 vdd.n2854 vdd.n579 19.0066
R3755 vdd.n1890 vdd.n1889 16.0975
R3756 vdd.n794 vdd.n793 16.0975
R3757 vdd.n1111 vdd.n1110 16.0975
R3758 vdd.n1148 vdd.n1147 16.0975
R3759 vdd.n1022 vdd.n1021 16.0975
R3760 vdd.n2046 vdd.n2045 16.0975
R3761 vdd.n1683 vdd.n1682 16.0975
R3762 vdd.n1643 vdd.n1642 16.0975
R3763 vdd.n1864 vdd.n1863 16.0975
R3764 vdd.n786 vdd.n785 16.0975
R3765 vdd.n2355 vdd.n2354 16.0975
R3766 vdd.n3022 vdd.n3021 16.0975
R3767 vdd.n428 vdd.n427 16.0975
R3768 vdd.n388 vdd.n387 16.0975
R3769 vdd.n581 vdd.n580 16.0975
R3770 vdd.n544 vdd.n543 16.0975
R3771 vdd.n662 vdd.n661 16.0975
R3772 vdd.n2352 vdd.n2351 16.0975
R3773 vdd.n2809 vdd.n2808 16.0975
R3774 vdd.n626 vdd.n625 16.0975
R3775 vdd.t228 vdd.n2316 15.4182
R3776 vdd.n2569 vdd.t111 15.4182
R3777 vdd.n28 vdd.n27 14.8792
R3778 vdd.n2087 vdd.n877 14.5112
R3779 vdd.n2771 vdd.n613 14.5112
R3780 vdd.n304 vdd.n269 13.1884
R3781 vdd.n253 vdd.n218 13.1884
R3782 vdd.n210 vdd.n175 13.1884
R3783 vdd.n159 vdd.n124 13.1884
R3784 vdd.n117 vdd.n82 13.1884
R3785 vdd.n66 vdd.n31 13.1884
R3786 vdd.n1499 vdd.n1464 13.1884
R3787 vdd.n1550 vdd.n1515 13.1884
R3788 vdd.n1405 vdd.n1370 13.1884
R3789 vdd.n1456 vdd.n1421 13.1884
R3790 vdd.n1312 vdd.n1277 13.1884
R3791 vdd.n1363 vdd.n1328 13.1884
R3792 vdd.n1180 vdd.n1023 12.9944
R3793 vdd.n1184 vdd.n1023 12.9944
R3794 vdd.n1789 vdd.n1641 12.9944
R3795 vdd.n1790 vdd.n1789 12.9944
R3796 vdd.n3101 vdd.n386 12.9944
R3797 vdd.n3102 vdd.n3101 12.9944
R3798 vdd.n2895 vdd.n545 12.9944
R3799 vdd.n2901 vdd.n545 12.9944
R3800 vdd.n305 vdd.n267 12.8005
R3801 vdd.n300 vdd.n271 12.8005
R3802 vdd.n254 vdd.n216 12.8005
R3803 vdd.n249 vdd.n220 12.8005
R3804 vdd.n211 vdd.n173 12.8005
R3805 vdd.n206 vdd.n177 12.8005
R3806 vdd.n160 vdd.n122 12.8005
R3807 vdd.n155 vdd.n126 12.8005
R3808 vdd.n118 vdd.n80 12.8005
R3809 vdd.n113 vdd.n84 12.8005
R3810 vdd.n67 vdd.n29 12.8005
R3811 vdd.n62 vdd.n33 12.8005
R3812 vdd.n1500 vdd.n1462 12.8005
R3813 vdd.n1495 vdd.n1466 12.8005
R3814 vdd.n1551 vdd.n1513 12.8005
R3815 vdd.n1546 vdd.n1517 12.8005
R3816 vdd.n1406 vdd.n1368 12.8005
R3817 vdd.n1401 vdd.n1372 12.8005
R3818 vdd.n1457 vdd.n1419 12.8005
R3819 vdd.n1452 vdd.n1423 12.8005
R3820 vdd.n1313 vdd.n1275 12.8005
R3821 vdd.n1308 vdd.n1279 12.8005
R3822 vdd.n1364 vdd.n1326 12.8005
R3823 vdd.n1359 vdd.n1330 12.8005
R3824 vdd.n299 vdd.n272 12.0247
R3825 vdd.n248 vdd.n221 12.0247
R3826 vdd.n205 vdd.n178 12.0247
R3827 vdd.n154 vdd.n127 12.0247
R3828 vdd.n112 vdd.n85 12.0247
R3829 vdd.n61 vdd.n34 12.0247
R3830 vdd.n1494 vdd.n1467 12.0247
R3831 vdd.n1545 vdd.n1518 12.0247
R3832 vdd.n1400 vdd.n1373 12.0247
R3833 vdd.n1451 vdd.n1424 12.0247
R3834 vdd.n1307 vdd.n1280 12.0247
R3835 vdd.n1358 vdd.n1331 12.0247
R3836 vdd.n1215 vdd.n983 11.337
R3837 vdd.n1223 vdd.n972 11.337
R3838 vdd.n1231 vdd.n972 11.337
R3839 vdd.n1239 vdd.n966 11.337
R3840 vdd.n1247 vdd.n959 11.337
R3841 vdd.n1256 vdd.n1255 11.337
R3842 vdd.n1264 vdd.n948 11.337
R3843 vdd.n1562 vdd.n937 11.337
R3844 vdd.n1571 vdd.n931 11.337
R3845 vdd.n1579 vdd.n925 11.337
R3846 vdd.n1588 vdd.n1587 11.337
R3847 vdd.n1596 vdd.n908 11.337
R3848 vdd.n1607 vdd.n908 11.337
R3849 vdd.n1607 vdd.n1606 11.337
R3850 vdd.n2948 vdd.n511 11.337
R3851 vdd.n2948 vdd.n505 11.337
R3852 vdd.n2956 vdd.n505 11.337
R3853 vdd.n2964 vdd.n499 11.337
R3854 vdd.n2972 vdd.n492 11.337
R3855 vdd.n2981 vdd.n2980 11.337
R3856 vdd.n2989 vdd.n481 11.337
R3857 vdd.n3163 vdd.n3162 11.337
R3858 vdd.n3156 vdd.n325 11.337
R3859 vdd.n3154 vdd.n329 11.337
R3860 vdd.n3148 vdd.n3147 11.337
R3861 vdd.n3146 vdd.n340 11.337
R3862 vdd.n3140 vdd.n340 11.337
R3863 vdd.n3139 vdd.n3138 11.337
R3864 vdd.n296 vdd.n295 11.249
R3865 vdd.n245 vdd.n244 11.249
R3866 vdd.n202 vdd.n201 11.249
R3867 vdd.n151 vdd.n150 11.249
R3868 vdd.n109 vdd.n108 11.249
R3869 vdd.n58 vdd.n57 11.249
R3870 vdd.n1491 vdd.n1490 11.249
R3871 vdd.n1542 vdd.n1541 11.249
R3872 vdd.n1397 vdd.n1396 11.249
R3873 vdd.n1448 vdd.n1447 11.249
R3874 vdd.n1304 vdd.n1303 11.249
R3875 vdd.n1355 vdd.n1354 11.249
R3876 vdd.n2244 vdd.t121 11.1103
R3877 vdd.n2576 vdd.t94 11.1103
R3878 vdd.n1231 vdd.t155 10.9969
R3879 vdd.t153 vdd.n3146 10.9969
R3880 vdd.n960 vdd.t188 10.7702
R3881 vdd.t167 vdd.n3155 10.7702
R3882 vdd.n281 vdd.n280 10.7238
R3883 vdd.n230 vdd.n229 10.7238
R3884 vdd.n187 vdd.n186 10.7238
R3885 vdd.n136 vdd.n135 10.7238
R3886 vdd.n94 vdd.n93 10.7238
R3887 vdd.n43 vdd.n42 10.7238
R3888 vdd.n1476 vdd.n1475 10.7238
R3889 vdd.n1527 vdd.n1526 10.7238
R3890 vdd.n1382 vdd.n1381 10.7238
R3891 vdd.n1433 vdd.n1432 10.7238
R3892 vdd.n1289 vdd.n1288 10.7238
R3893 vdd.n1340 vdd.n1339 10.7238
R3894 vdd.n2090 vdd.n2089 10.6151
R3895 vdd.n2091 vdd.n2090 10.6151
R3896 vdd.n2091 vdd.n863 10.6151
R3897 vdd.n2101 vdd.n863 10.6151
R3898 vdd.n2102 vdd.n2101 10.6151
R3899 vdd.n2103 vdd.n2102 10.6151
R3900 vdd.n2103 vdd.n850 10.6151
R3901 vdd.n2114 vdd.n850 10.6151
R3902 vdd.n2115 vdd.n2114 10.6151
R3903 vdd.n2116 vdd.n2115 10.6151
R3904 vdd.n2116 vdd.n838 10.6151
R3905 vdd.n2126 vdd.n838 10.6151
R3906 vdd.n2127 vdd.n2126 10.6151
R3907 vdd.n2128 vdd.n2127 10.6151
R3908 vdd.n2128 vdd.n826 10.6151
R3909 vdd.n2138 vdd.n826 10.6151
R3910 vdd.n2139 vdd.n2138 10.6151
R3911 vdd.n2140 vdd.n2139 10.6151
R3912 vdd.n2140 vdd.n815 10.6151
R3913 vdd.n2150 vdd.n815 10.6151
R3914 vdd.n2151 vdd.n2150 10.6151
R3915 vdd.n2152 vdd.n2151 10.6151
R3916 vdd.n2152 vdd.n802 10.6151
R3917 vdd.n2164 vdd.n802 10.6151
R3918 vdd.n2165 vdd.n2164 10.6151
R3919 vdd.n2167 vdd.n2165 10.6151
R3920 vdd.n2167 vdd.n2166 10.6151
R3921 vdd.n2166 vdd.n784 10.6151
R3922 vdd.n2314 vdd.n2313 10.6151
R3923 vdd.n2313 vdd.n2312 10.6151
R3924 vdd.n2312 vdd.n2309 10.6151
R3925 vdd.n2309 vdd.n2308 10.6151
R3926 vdd.n2308 vdd.n2305 10.6151
R3927 vdd.n2305 vdd.n2304 10.6151
R3928 vdd.n2304 vdd.n2301 10.6151
R3929 vdd.n2301 vdd.n2300 10.6151
R3930 vdd.n2300 vdd.n2297 10.6151
R3931 vdd.n2297 vdd.n2296 10.6151
R3932 vdd.n2296 vdd.n2293 10.6151
R3933 vdd.n2293 vdd.n2292 10.6151
R3934 vdd.n2292 vdd.n2289 10.6151
R3935 vdd.n2289 vdd.n2288 10.6151
R3936 vdd.n2288 vdd.n2285 10.6151
R3937 vdd.n2285 vdd.n2284 10.6151
R3938 vdd.n2284 vdd.n2281 10.6151
R3939 vdd.n2281 vdd.n2280 10.6151
R3940 vdd.n2280 vdd.n2277 10.6151
R3941 vdd.n2277 vdd.n2276 10.6151
R3942 vdd.n2276 vdd.n2273 10.6151
R3943 vdd.n2273 vdd.n2272 10.6151
R3944 vdd.n2272 vdd.n2269 10.6151
R3945 vdd.n2269 vdd.n2268 10.6151
R3946 vdd.n2268 vdd.n2265 10.6151
R3947 vdd.n2265 vdd.n2264 10.6151
R3948 vdd.n2264 vdd.n2261 10.6151
R3949 vdd.n2261 vdd.n2260 10.6151
R3950 vdd.n2260 vdd.n2257 10.6151
R3951 vdd.n2257 vdd.n2256 10.6151
R3952 vdd.n2256 vdd.n2253 10.6151
R3953 vdd.n2251 vdd.n2248 10.6151
R3954 vdd.n2248 vdd.n2247 10.6151
R3955 vdd.n1990 vdd.n1989 10.6151
R3956 vdd.n1989 vdd.n1987 10.6151
R3957 vdd.n1987 vdd.n1986 10.6151
R3958 vdd.n1986 vdd.n1984 10.6151
R3959 vdd.n1984 vdd.n1983 10.6151
R3960 vdd.n1983 vdd.n1981 10.6151
R3961 vdd.n1981 vdd.n1980 10.6151
R3962 vdd.n1980 vdd.n1978 10.6151
R3963 vdd.n1978 vdd.n1977 10.6151
R3964 vdd.n1977 vdd.n1975 10.6151
R3965 vdd.n1975 vdd.n1974 10.6151
R3966 vdd.n1974 vdd.n1972 10.6151
R3967 vdd.n1972 vdd.n1971 10.6151
R3968 vdd.n1971 vdd.n1886 10.6151
R3969 vdd.n1886 vdd.n1885 10.6151
R3970 vdd.n1885 vdd.n1883 10.6151
R3971 vdd.n1883 vdd.n1882 10.6151
R3972 vdd.n1882 vdd.n1880 10.6151
R3973 vdd.n1880 vdd.n1879 10.6151
R3974 vdd.n1879 vdd.n1877 10.6151
R3975 vdd.n1877 vdd.n1876 10.6151
R3976 vdd.n1876 vdd.n1874 10.6151
R3977 vdd.n1874 vdd.n1873 10.6151
R3978 vdd.n1873 vdd.n1871 10.6151
R3979 vdd.n1871 vdd.n1870 10.6151
R3980 vdd.n1870 vdd.n1867 10.6151
R3981 vdd.n1867 vdd.n1866 10.6151
R3982 vdd.n1866 vdd.n787 10.6151
R3983 vdd.n1824 vdd.n875 10.6151
R3984 vdd.n1825 vdd.n1824 10.6151
R3985 vdd.n1826 vdd.n1825 10.6151
R3986 vdd.n1826 vdd.n1820 10.6151
R3987 vdd.n1832 vdd.n1820 10.6151
R3988 vdd.n1833 vdd.n1832 10.6151
R3989 vdd.n1834 vdd.n1833 10.6151
R3990 vdd.n1834 vdd.n1818 10.6151
R3991 vdd.n1840 vdd.n1818 10.6151
R3992 vdd.n1841 vdd.n1840 10.6151
R3993 vdd.n1842 vdd.n1841 10.6151
R3994 vdd.n1842 vdd.n1816 10.6151
R3995 vdd.n1848 vdd.n1816 10.6151
R3996 vdd.n1849 vdd.n1848 10.6151
R3997 vdd.n1850 vdd.n1849 10.6151
R3998 vdd.n1850 vdd.n1814 10.6151
R3999 vdd.n2026 vdd.n1814 10.6151
R4000 vdd.n2026 vdd.n2025 10.6151
R4001 vdd.n2025 vdd.n1855 10.6151
R4002 vdd.n2019 vdd.n1855 10.6151
R4003 vdd.n2019 vdd.n2018 10.6151
R4004 vdd.n2018 vdd.n2017 10.6151
R4005 vdd.n2017 vdd.n1857 10.6151
R4006 vdd.n2011 vdd.n1857 10.6151
R4007 vdd.n2011 vdd.n2010 10.6151
R4008 vdd.n2010 vdd.n2009 10.6151
R4009 vdd.n2009 vdd.n1859 10.6151
R4010 vdd.n2003 vdd.n1859 10.6151
R4011 vdd.n2003 vdd.n2002 10.6151
R4012 vdd.n2002 vdd.n2001 10.6151
R4013 vdd.n2001 vdd.n1861 10.6151
R4014 vdd.n1995 vdd.n1994 10.6151
R4015 vdd.n1994 vdd.n1993 10.6151
R4016 vdd.n2499 vdd.n2498 10.6151
R4017 vdd.n2498 vdd.n2496 10.6151
R4018 vdd.n2496 vdd.n2495 10.6151
R4019 vdd.n2495 vdd.n2353 10.6151
R4020 vdd.n2442 vdd.n2353 10.6151
R4021 vdd.n2443 vdd.n2442 10.6151
R4022 vdd.n2445 vdd.n2443 10.6151
R4023 vdd.n2446 vdd.n2445 10.6151
R4024 vdd.n2448 vdd.n2446 10.6151
R4025 vdd.n2449 vdd.n2448 10.6151
R4026 vdd.n2451 vdd.n2449 10.6151
R4027 vdd.n2452 vdd.n2451 10.6151
R4028 vdd.n2454 vdd.n2452 10.6151
R4029 vdd.n2455 vdd.n2454 10.6151
R4030 vdd.n2470 vdd.n2455 10.6151
R4031 vdd.n2470 vdd.n2469 10.6151
R4032 vdd.n2469 vdd.n2468 10.6151
R4033 vdd.n2468 vdd.n2466 10.6151
R4034 vdd.n2466 vdd.n2465 10.6151
R4035 vdd.n2465 vdd.n2463 10.6151
R4036 vdd.n2463 vdd.n2462 10.6151
R4037 vdd.n2462 vdd.n2460 10.6151
R4038 vdd.n2460 vdd.n2459 10.6151
R4039 vdd.n2459 vdd.n2457 10.6151
R4040 vdd.n2457 vdd.n2456 10.6151
R4041 vdd.n2456 vdd.n664 10.6151
R4042 vdd.n2704 vdd.n664 10.6151
R4043 vdd.n2705 vdd.n2704 10.6151
R4044 vdd.n2566 vdd.n740 10.6151
R4045 vdd.n2566 vdd.n2565 10.6151
R4046 vdd.n2565 vdd.n2564 10.6151
R4047 vdd.n2564 vdd.n2562 10.6151
R4048 vdd.n2562 vdd.n2559 10.6151
R4049 vdd.n2559 vdd.n2558 10.6151
R4050 vdd.n2558 vdd.n2555 10.6151
R4051 vdd.n2555 vdd.n2554 10.6151
R4052 vdd.n2554 vdd.n2551 10.6151
R4053 vdd.n2551 vdd.n2550 10.6151
R4054 vdd.n2550 vdd.n2547 10.6151
R4055 vdd.n2547 vdd.n2546 10.6151
R4056 vdd.n2546 vdd.n2543 10.6151
R4057 vdd.n2543 vdd.n2542 10.6151
R4058 vdd.n2542 vdd.n2539 10.6151
R4059 vdd.n2539 vdd.n2538 10.6151
R4060 vdd.n2538 vdd.n2535 10.6151
R4061 vdd.n2535 vdd.n2534 10.6151
R4062 vdd.n2534 vdd.n2531 10.6151
R4063 vdd.n2531 vdd.n2530 10.6151
R4064 vdd.n2530 vdd.n2527 10.6151
R4065 vdd.n2527 vdd.n2526 10.6151
R4066 vdd.n2526 vdd.n2523 10.6151
R4067 vdd.n2523 vdd.n2522 10.6151
R4068 vdd.n2522 vdd.n2519 10.6151
R4069 vdd.n2519 vdd.n2518 10.6151
R4070 vdd.n2518 vdd.n2515 10.6151
R4071 vdd.n2515 vdd.n2514 10.6151
R4072 vdd.n2514 vdd.n2511 10.6151
R4073 vdd.n2511 vdd.n2510 10.6151
R4074 vdd.n2510 vdd.n2507 10.6151
R4075 vdd.n2505 vdd.n2502 10.6151
R4076 vdd.n2502 vdd.n2501 10.6151
R4077 vdd.n2579 vdd.n2578 10.6151
R4078 vdd.n2580 vdd.n2579 10.6151
R4079 vdd.n2580 vdd.n730 10.6151
R4080 vdd.n2590 vdd.n730 10.6151
R4081 vdd.n2591 vdd.n2590 10.6151
R4082 vdd.n2592 vdd.n2591 10.6151
R4083 vdd.n2592 vdd.n717 10.6151
R4084 vdd.n2602 vdd.n717 10.6151
R4085 vdd.n2603 vdd.n2602 10.6151
R4086 vdd.n2604 vdd.n2603 10.6151
R4087 vdd.n2604 vdd.n706 10.6151
R4088 vdd.n2614 vdd.n706 10.6151
R4089 vdd.n2615 vdd.n2614 10.6151
R4090 vdd.n2616 vdd.n2615 10.6151
R4091 vdd.n2616 vdd.n694 10.6151
R4092 vdd.n2626 vdd.n694 10.6151
R4093 vdd.n2627 vdd.n2626 10.6151
R4094 vdd.n2628 vdd.n2627 10.6151
R4095 vdd.n2628 vdd.n683 10.6151
R4096 vdd.n2640 vdd.n683 10.6151
R4097 vdd.n2641 vdd.n2640 10.6151
R4098 vdd.n2642 vdd.n2641 10.6151
R4099 vdd.n2642 vdd.n669 10.6151
R4100 vdd.n2697 vdd.n669 10.6151
R4101 vdd.n2698 vdd.n2697 10.6151
R4102 vdd.n2699 vdd.n2698 10.6151
R4103 vdd.n2699 vdd.n636 10.6151
R4104 vdd.n2769 vdd.n636 10.6151
R4105 vdd.n2768 vdd.n2767 10.6151
R4106 vdd.n2767 vdd.n637 10.6151
R4107 vdd.n638 vdd.n637 10.6151
R4108 vdd.n2760 vdd.n638 10.6151
R4109 vdd.n2760 vdd.n2759 10.6151
R4110 vdd.n2759 vdd.n2758 10.6151
R4111 vdd.n2758 vdd.n640 10.6151
R4112 vdd.n2753 vdd.n640 10.6151
R4113 vdd.n2753 vdd.n2752 10.6151
R4114 vdd.n2752 vdd.n2751 10.6151
R4115 vdd.n2751 vdd.n643 10.6151
R4116 vdd.n2746 vdd.n643 10.6151
R4117 vdd.n2746 vdd.n2745 10.6151
R4118 vdd.n2745 vdd.n2744 10.6151
R4119 vdd.n2744 vdd.n646 10.6151
R4120 vdd.n2739 vdd.n646 10.6151
R4121 vdd.n2739 vdd.n2738 10.6151
R4122 vdd.n2738 vdd.n2736 10.6151
R4123 vdd.n2736 vdd.n649 10.6151
R4124 vdd.n2731 vdd.n649 10.6151
R4125 vdd.n2731 vdd.n2730 10.6151
R4126 vdd.n2730 vdd.n2729 10.6151
R4127 vdd.n2729 vdd.n652 10.6151
R4128 vdd.n2724 vdd.n652 10.6151
R4129 vdd.n2724 vdd.n2723 10.6151
R4130 vdd.n2723 vdd.n2722 10.6151
R4131 vdd.n2722 vdd.n655 10.6151
R4132 vdd.n2717 vdd.n655 10.6151
R4133 vdd.n2717 vdd.n2716 10.6151
R4134 vdd.n2716 vdd.n2715 10.6151
R4135 vdd.n2715 vdd.n658 10.6151
R4136 vdd.n2710 vdd.n2709 10.6151
R4137 vdd.n2709 vdd.n2708 10.6151
R4138 vdd.n2687 vdd.n2648 10.6151
R4139 vdd.n2682 vdd.n2648 10.6151
R4140 vdd.n2682 vdd.n2681 10.6151
R4141 vdd.n2681 vdd.n2680 10.6151
R4142 vdd.n2680 vdd.n2650 10.6151
R4143 vdd.n2675 vdd.n2650 10.6151
R4144 vdd.n2675 vdd.n2674 10.6151
R4145 vdd.n2674 vdd.n2673 10.6151
R4146 vdd.n2673 vdd.n2653 10.6151
R4147 vdd.n2668 vdd.n2653 10.6151
R4148 vdd.n2668 vdd.n2667 10.6151
R4149 vdd.n2667 vdd.n2666 10.6151
R4150 vdd.n2666 vdd.n2656 10.6151
R4151 vdd.n2661 vdd.n2656 10.6151
R4152 vdd.n2661 vdd.n2660 10.6151
R4153 vdd.n2660 vdd.n610 10.6151
R4154 vdd.n2804 vdd.n610 10.6151
R4155 vdd.n2804 vdd.n611 10.6151
R4156 vdd.n614 vdd.n611 10.6151
R4157 vdd.n2797 vdd.n614 10.6151
R4158 vdd.n2797 vdd.n2796 10.6151
R4159 vdd.n2796 vdd.n2795 10.6151
R4160 vdd.n2795 vdd.n616 10.6151
R4161 vdd.n2790 vdd.n616 10.6151
R4162 vdd.n2790 vdd.n2789 10.6151
R4163 vdd.n2789 vdd.n2788 10.6151
R4164 vdd.n2788 vdd.n619 10.6151
R4165 vdd.n2783 vdd.n619 10.6151
R4166 vdd.n2783 vdd.n2782 10.6151
R4167 vdd.n2782 vdd.n2781 10.6151
R4168 vdd.n2781 vdd.n622 10.6151
R4169 vdd.n2776 vdd.n2775 10.6151
R4170 vdd.n2775 vdd.n2774 10.6151
R4171 vdd.n2422 vdd.n2420 10.6151
R4172 vdd.n2423 vdd.n2422 10.6151
R4173 vdd.n2491 vdd.n2423 10.6151
R4174 vdd.n2491 vdd.n2490 10.6151
R4175 vdd.n2490 vdd.n2489 10.6151
R4176 vdd.n2489 vdd.n2487 10.6151
R4177 vdd.n2487 vdd.n2486 10.6151
R4178 vdd.n2486 vdd.n2484 10.6151
R4179 vdd.n2484 vdd.n2483 10.6151
R4180 vdd.n2483 vdd.n2481 10.6151
R4181 vdd.n2481 vdd.n2480 10.6151
R4182 vdd.n2480 vdd.n2478 10.6151
R4183 vdd.n2478 vdd.n2477 10.6151
R4184 vdd.n2477 vdd.n2475 10.6151
R4185 vdd.n2475 vdd.n2474 10.6151
R4186 vdd.n2474 vdd.n2440 10.6151
R4187 vdd.n2440 vdd.n2439 10.6151
R4188 vdd.n2439 vdd.n2437 10.6151
R4189 vdd.n2437 vdd.n2436 10.6151
R4190 vdd.n2436 vdd.n2434 10.6151
R4191 vdd.n2434 vdd.n2433 10.6151
R4192 vdd.n2433 vdd.n2431 10.6151
R4193 vdd.n2431 vdd.n2430 10.6151
R4194 vdd.n2430 vdd.n2428 10.6151
R4195 vdd.n2428 vdd.n2427 10.6151
R4196 vdd.n2427 vdd.n2425 10.6151
R4197 vdd.n2425 vdd.n2424 10.6151
R4198 vdd.n2424 vdd.n628 10.6151
R4199 vdd.n2573 vdd.n2572 10.6151
R4200 vdd.n2572 vdd.n745 10.6151
R4201 vdd.n2357 vdd.n745 10.6151
R4202 vdd.n2360 vdd.n2357 10.6151
R4203 vdd.n2361 vdd.n2360 10.6151
R4204 vdd.n2364 vdd.n2361 10.6151
R4205 vdd.n2365 vdd.n2364 10.6151
R4206 vdd.n2368 vdd.n2365 10.6151
R4207 vdd.n2369 vdd.n2368 10.6151
R4208 vdd.n2372 vdd.n2369 10.6151
R4209 vdd.n2373 vdd.n2372 10.6151
R4210 vdd.n2376 vdd.n2373 10.6151
R4211 vdd.n2377 vdd.n2376 10.6151
R4212 vdd.n2380 vdd.n2377 10.6151
R4213 vdd.n2381 vdd.n2380 10.6151
R4214 vdd.n2384 vdd.n2381 10.6151
R4215 vdd.n2385 vdd.n2384 10.6151
R4216 vdd.n2388 vdd.n2385 10.6151
R4217 vdd.n2389 vdd.n2388 10.6151
R4218 vdd.n2392 vdd.n2389 10.6151
R4219 vdd.n2393 vdd.n2392 10.6151
R4220 vdd.n2396 vdd.n2393 10.6151
R4221 vdd.n2397 vdd.n2396 10.6151
R4222 vdd.n2400 vdd.n2397 10.6151
R4223 vdd.n2401 vdd.n2400 10.6151
R4224 vdd.n2404 vdd.n2401 10.6151
R4225 vdd.n2405 vdd.n2404 10.6151
R4226 vdd.n2408 vdd.n2405 10.6151
R4227 vdd.n2409 vdd.n2408 10.6151
R4228 vdd.n2412 vdd.n2409 10.6151
R4229 vdd.n2413 vdd.n2412 10.6151
R4230 vdd.n2418 vdd.n2416 10.6151
R4231 vdd.n2419 vdd.n2418 10.6151
R4232 vdd.n2574 vdd.n735 10.6151
R4233 vdd.n2584 vdd.n735 10.6151
R4234 vdd.n2585 vdd.n2584 10.6151
R4235 vdd.n2586 vdd.n2585 10.6151
R4236 vdd.n2586 vdd.n723 10.6151
R4237 vdd.n2596 vdd.n723 10.6151
R4238 vdd.n2597 vdd.n2596 10.6151
R4239 vdd.n2598 vdd.n2597 10.6151
R4240 vdd.n2598 vdd.n712 10.6151
R4241 vdd.n2608 vdd.n712 10.6151
R4242 vdd.n2609 vdd.n2608 10.6151
R4243 vdd.n2610 vdd.n2609 10.6151
R4244 vdd.n2610 vdd.n700 10.6151
R4245 vdd.n2620 vdd.n700 10.6151
R4246 vdd.n2621 vdd.n2620 10.6151
R4247 vdd.n2622 vdd.n2621 10.6151
R4248 vdd.n2622 vdd.n689 10.6151
R4249 vdd.n2632 vdd.n689 10.6151
R4250 vdd.n2633 vdd.n2632 10.6151
R4251 vdd.n2636 vdd.n2633 10.6151
R4252 vdd.n2646 vdd.n677 10.6151
R4253 vdd.n2647 vdd.n2646 10.6151
R4254 vdd.n2693 vdd.n2647 10.6151
R4255 vdd.n2693 vdd.n2692 10.6151
R4256 vdd.n2692 vdd.n2691 10.6151
R4257 vdd.n2691 vdd.n2690 10.6151
R4258 vdd.n2690 vdd.n2688 10.6151
R4259 vdd.n2085 vdd.n869 10.6151
R4260 vdd.n2095 vdd.n869 10.6151
R4261 vdd.n2096 vdd.n2095 10.6151
R4262 vdd.n2097 vdd.n2096 10.6151
R4263 vdd.n2097 vdd.n856 10.6151
R4264 vdd.n2107 vdd.n856 10.6151
R4265 vdd.n2108 vdd.n2107 10.6151
R4266 vdd.n2110 vdd.n844 10.6151
R4267 vdd.n2120 vdd.n844 10.6151
R4268 vdd.n2121 vdd.n2120 10.6151
R4269 vdd.n2122 vdd.n2121 10.6151
R4270 vdd.n2122 vdd.n832 10.6151
R4271 vdd.n2132 vdd.n832 10.6151
R4272 vdd.n2133 vdd.n2132 10.6151
R4273 vdd.n2134 vdd.n2133 10.6151
R4274 vdd.n2134 vdd.n821 10.6151
R4275 vdd.n2144 vdd.n821 10.6151
R4276 vdd.n2145 vdd.n2144 10.6151
R4277 vdd.n2146 vdd.n2145 10.6151
R4278 vdd.n2146 vdd.n809 10.6151
R4279 vdd.n2156 vdd.n809 10.6151
R4280 vdd.n2157 vdd.n2156 10.6151
R4281 vdd.n2160 vdd.n2157 10.6151
R4282 vdd.n2160 vdd.n2159 10.6151
R4283 vdd.n2159 vdd.n2158 10.6151
R4284 vdd.n2158 vdd.n792 10.6151
R4285 vdd.n2242 vdd.n792 10.6151
R4286 vdd.n2241 vdd.n2240 10.6151
R4287 vdd.n2240 vdd.n2237 10.6151
R4288 vdd.n2237 vdd.n2236 10.6151
R4289 vdd.n2236 vdd.n2233 10.6151
R4290 vdd.n2233 vdd.n2232 10.6151
R4291 vdd.n2232 vdd.n2229 10.6151
R4292 vdd.n2229 vdd.n2228 10.6151
R4293 vdd.n2228 vdd.n2225 10.6151
R4294 vdd.n2225 vdd.n2224 10.6151
R4295 vdd.n2224 vdd.n2221 10.6151
R4296 vdd.n2221 vdd.n2220 10.6151
R4297 vdd.n2220 vdd.n2217 10.6151
R4298 vdd.n2217 vdd.n2216 10.6151
R4299 vdd.n2216 vdd.n2213 10.6151
R4300 vdd.n2213 vdd.n2212 10.6151
R4301 vdd.n2212 vdd.n2209 10.6151
R4302 vdd.n2209 vdd.n2208 10.6151
R4303 vdd.n2208 vdd.n2205 10.6151
R4304 vdd.n2205 vdd.n2204 10.6151
R4305 vdd.n2204 vdd.n2201 10.6151
R4306 vdd.n2201 vdd.n2200 10.6151
R4307 vdd.n2200 vdd.n2197 10.6151
R4308 vdd.n2197 vdd.n2196 10.6151
R4309 vdd.n2196 vdd.n2193 10.6151
R4310 vdd.n2193 vdd.n2192 10.6151
R4311 vdd.n2192 vdd.n2189 10.6151
R4312 vdd.n2189 vdd.n2188 10.6151
R4313 vdd.n2188 vdd.n2185 10.6151
R4314 vdd.n2185 vdd.n2184 10.6151
R4315 vdd.n2184 vdd.n2181 10.6151
R4316 vdd.n2181 vdd.n2180 10.6151
R4317 vdd.n2177 vdd.n2176 10.6151
R4318 vdd.n2176 vdd.n2174 10.6151
R4319 vdd.n1933 vdd.n1931 10.6151
R4320 vdd.n1934 vdd.n1933 10.6151
R4321 vdd.n1936 vdd.n1934 10.6151
R4322 vdd.n1937 vdd.n1936 10.6151
R4323 vdd.n1939 vdd.n1937 10.6151
R4324 vdd.n1940 vdd.n1939 10.6151
R4325 vdd.n1942 vdd.n1940 10.6151
R4326 vdd.n1943 vdd.n1942 10.6151
R4327 vdd.n1945 vdd.n1943 10.6151
R4328 vdd.n1946 vdd.n1945 10.6151
R4329 vdd.n1948 vdd.n1946 10.6151
R4330 vdd.n1949 vdd.n1948 10.6151
R4331 vdd.n1967 vdd.n1949 10.6151
R4332 vdd.n1967 vdd.n1966 10.6151
R4333 vdd.n1966 vdd.n1965 10.6151
R4334 vdd.n1965 vdd.n1963 10.6151
R4335 vdd.n1963 vdd.n1962 10.6151
R4336 vdd.n1962 vdd.n1960 10.6151
R4337 vdd.n1960 vdd.n1959 10.6151
R4338 vdd.n1959 vdd.n1957 10.6151
R4339 vdd.n1957 vdd.n1956 10.6151
R4340 vdd.n1956 vdd.n1954 10.6151
R4341 vdd.n1954 vdd.n1953 10.6151
R4342 vdd.n1953 vdd.n1951 10.6151
R4343 vdd.n1951 vdd.n1950 10.6151
R4344 vdd.n1950 vdd.n796 10.6151
R4345 vdd.n2172 vdd.n796 10.6151
R4346 vdd.n2173 vdd.n2172 10.6151
R4347 vdd.n2084 vdd.n2083 10.6151
R4348 vdd.n2083 vdd.n881 10.6151
R4349 vdd.n2077 vdd.n881 10.6151
R4350 vdd.n2077 vdd.n2076 10.6151
R4351 vdd.n2076 vdd.n2075 10.6151
R4352 vdd.n2075 vdd.n883 10.6151
R4353 vdd.n2069 vdd.n883 10.6151
R4354 vdd.n2069 vdd.n2068 10.6151
R4355 vdd.n2068 vdd.n2067 10.6151
R4356 vdd.n2067 vdd.n885 10.6151
R4357 vdd.n2061 vdd.n885 10.6151
R4358 vdd.n2061 vdd.n2060 10.6151
R4359 vdd.n2060 vdd.n2059 10.6151
R4360 vdd.n2059 vdd.n887 10.6151
R4361 vdd.n2053 vdd.n887 10.6151
R4362 vdd.n2053 vdd.n2052 10.6151
R4363 vdd.n2052 vdd.n2051 10.6151
R4364 vdd.n2051 vdd.n891 10.6151
R4365 vdd.n1899 vdd.n891 10.6151
R4366 vdd.n1900 vdd.n1899 10.6151
R4367 vdd.n1900 vdd.n1895 10.6151
R4368 vdd.n1906 vdd.n1895 10.6151
R4369 vdd.n1907 vdd.n1906 10.6151
R4370 vdd.n1908 vdd.n1907 10.6151
R4371 vdd.n1908 vdd.n1893 10.6151
R4372 vdd.n1914 vdd.n1893 10.6151
R4373 vdd.n1915 vdd.n1914 10.6151
R4374 vdd.n1916 vdd.n1915 10.6151
R4375 vdd.n1916 vdd.n1891 10.6151
R4376 vdd.n1922 vdd.n1891 10.6151
R4377 vdd.n1923 vdd.n1922 10.6151
R4378 vdd.n1925 vdd.n1887 10.6151
R4379 vdd.n1930 vdd.n1887 10.6151
R4380 vdd.n1272 vdd.t138 10.5435
R4381 vdd.n2041 vdd.t23 10.5435
R4382 vdd.n2940 vdd.t16 10.5435
R4383 vdd.n3164 vdd.t199 10.5435
R4384 vdd.n292 vdd.n274 10.4732
R4385 vdd.n241 vdd.n223 10.4732
R4386 vdd.n198 vdd.n180 10.4732
R4387 vdd.n147 vdd.n129 10.4732
R4388 vdd.n105 vdd.n87 10.4732
R4389 vdd.n54 vdd.n36 10.4732
R4390 vdd.n1487 vdd.n1469 10.4732
R4391 vdd.n1538 vdd.n1520 10.4732
R4392 vdd.n1393 vdd.n1375 10.4732
R4393 vdd.n1444 vdd.n1426 10.4732
R4394 vdd.n1300 vdd.n1282 10.4732
R4395 vdd.n1351 vdd.n1333 10.4732
R4396 vdd.n1570 vdd.t150 10.3167
R4397 vdd.t183 vdd.n493 10.3167
R4398 vdd.n1223 vdd.t4 9.86327
R4399 vdd.n3140 vdd.t12 9.86327
R4400 vdd.n291 vdd.n276 9.69747
R4401 vdd.n240 vdd.n225 9.69747
R4402 vdd.n197 vdd.n182 9.69747
R4403 vdd.n146 vdd.n131 9.69747
R4404 vdd.n104 vdd.n89 9.69747
R4405 vdd.n53 vdd.n38 9.69747
R4406 vdd.n1486 vdd.n1471 9.69747
R4407 vdd.n1537 vdd.n1522 9.69747
R4408 vdd.n1392 vdd.n1377 9.69747
R4409 vdd.n1443 vdd.n1428 9.69747
R4410 vdd.n1299 vdd.n1284 9.69747
R4411 vdd.n1350 vdd.n1335 9.69747
R4412 vdd.n2027 vdd.n2026 9.67831
R4413 vdd.n2738 vdd.n2737 9.67831
R4414 vdd.n2805 vdd.n2804 9.67831
R4415 vdd.n2051 vdd.n2050 9.67831
R4416 vdd.n307 vdd.n306 9.45567
R4417 vdd.n256 vdd.n255 9.45567
R4418 vdd.n213 vdd.n212 9.45567
R4419 vdd.n162 vdd.n161 9.45567
R4420 vdd.n120 vdd.n119 9.45567
R4421 vdd.n69 vdd.n68 9.45567
R4422 vdd.n1502 vdd.n1501 9.45567
R4423 vdd.n1553 vdd.n1552 9.45567
R4424 vdd.n1408 vdd.n1407 9.45567
R4425 vdd.n1459 vdd.n1458 9.45567
R4426 vdd.n1315 vdd.n1314 9.45567
R4427 vdd.n1366 vdd.n1365 9.45567
R4428 vdd.n1787 vdd.n1641 9.3005
R4429 vdd.n1786 vdd.n1785 9.3005
R4430 vdd.n1647 vdd.n1646 9.3005
R4431 vdd.n1780 vdd.n1651 9.3005
R4432 vdd.n1779 vdd.n1652 9.3005
R4433 vdd.n1778 vdd.n1653 9.3005
R4434 vdd.n1657 vdd.n1654 9.3005
R4435 vdd.n1773 vdd.n1658 9.3005
R4436 vdd.n1772 vdd.n1659 9.3005
R4437 vdd.n1771 vdd.n1660 9.3005
R4438 vdd.n1664 vdd.n1661 9.3005
R4439 vdd.n1766 vdd.n1665 9.3005
R4440 vdd.n1765 vdd.n1666 9.3005
R4441 vdd.n1764 vdd.n1667 9.3005
R4442 vdd.n1671 vdd.n1668 9.3005
R4443 vdd.n1759 vdd.n1672 9.3005
R4444 vdd.n1758 vdd.n1673 9.3005
R4445 vdd.n1757 vdd.n1674 9.3005
R4446 vdd.n1678 vdd.n1675 9.3005
R4447 vdd.n1752 vdd.n1679 9.3005
R4448 vdd.n1751 vdd.n1680 9.3005
R4449 vdd.n1750 vdd.n1749 9.3005
R4450 vdd.n1748 vdd.n1681 9.3005
R4451 vdd.n1747 vdd.n1746 9.3005
R4452 vdd.n1687 vdd.n1686 9.3005
R4453 vdd.n1741 vdd.n1691 9.3005
R4454 vdd.n1740 vdd.n1692 9.3005
R4455 vdd.n1739 vdd.n1693 9.3005
R4456 vdd.n1697 vdd.n1694 9.3005
R4457 vdd.n1734 vdd.n1698 9.3005
R4458 vdd.n1733 vdd.n1699 9.3005
R4459 vdd.n1732 vdd.n1700 9.3005
R4460 vdd.n1704 vdd.n1701 9.3005
R4461 vdd.n1727 vdd.n1705 9.3005
R4462 vdd.n1726 vdd.n1706 9.3005
R4463 vdd.n1725 vdd.n1707 9.3005
R4464 vdd.n1709 vdd.n1708 9.3005
R4465 vdd.n1720 vdd.n892 9.3005
R4466 vdd.n1789 vdd.n1788 9.3005
R4467 vdd.n1813 vdd.n1812 9.3005
R4468 vdd.n1619 vdd.n1618 9.3005
R4469 vdd.n1624 vdd.n1622 9.3005
R4470 vdd.n1805 vdd.n1625 9.3005
R4471 vdd.n1804 vdd.n1626 9.3005
R4472 vdd.n1803 vdd.n1627 9.3005
R4473 vdd.n1631 vdd.n1628 9.3005
R4474 vdd.n1798 vdd.n1632 9.3005
R4475 vdd.n1797 vdd.n1633 9.3005
R4476 vdd.n1796 vdd.n1634 9.3005
R4477 vdd.n1638 vdd.n1635 9.3005
R4478 vdd.n1791 vdd.n1639 9.3005
R4479 vdd.n1790 vdd.n1640 9.3005
R4480 vdd.n2035 vdd.n1612 9.3005
R4481 vdd.n2037 vdd.n2036 9.3005
R4482 vdd.n1558 vdd.n939 9.3005
R4483 vdd.n1560 vdd.n1559 9.3005
R4484 vdd.n929 vdd.n928 9.3005
R4485 vdd.n1574 vdd.n1573 9.3005
R4486 vdd.n1575 vdd.n927 9.3005
R4487 vdd.n1577 vdd.n1576 9.3005
R4488 vdd.n918 vdd.n917 9.3005
R4489 vdd.n1591 vdd.n1590 9.3005
R4490 vdd.n1592 vdd.n916 9.3005
R4491 vdd.n1594 vdd.n1593 9.3005
R4492 vdd.n906 vdd.n905 9.3005
R4493 vdd.n1610 vdd.n1609 9.3005
R4494 vdd.n1611 vdd.n904 9.3005
R4495 vdd.n2039 vdd.n2038 9.3005
R4496 vdd.n283 vdd.n282 9.3005
R4497 vdd.n278 vdd.n277 9.3005
R4498 vdd.n289 vdd.n288 9.3005
R4499 vdd.n291 vdd.n290 9.3005
R4500 vdd.n274 vdd.n273 9.3005
R4501 vdd.n297 vdd.n296 9.3005
R4502 vdd.n299 vdd.n298 9.3005
R4503 vdd.n271 vdd.n268 9.3005
R4504 vdd.n306 vdd.n305 9.3005
R4505 vdd.n232 vdd.n231 9.3005
R4506 vdd.n227 vdd.n226 9.3005
R4507 vdd.n238 vdd.n237 9.3005
R4508 vdd.n240 vdd.n239 9.3005
R4509 vdd.n223 vdd.n222 9.3005
R4510 vdd.n246 vdd.n245 9.3005
R4511 vdd.n248 vdd.n247 9.3005
R4512 vdd.n220 vdd.n217 9.3005
R4513 vdd.n255 vdd.n254 9.3005
R4514 vdd.n189 vdd.n188 9.3005
R4515 vdd.n184 vdd.n183 9.3005
R4516 vdd.n195 vdd.n194 9.3005
R4517 vdd.n197 vdd.n196 9.3005
R4518 vdd.n180 vdd.n179 9.3005
R4519 vdd.n203 vdd.n202 9.3005
R4520 vdd.n205 vdd.n204 9.3005
R4521 vdd.n177 vdd.n174 9.3005
R4522 vdd.n212 vdd.n211 9.3005
R4523 vdd.n138 vdd.n137 9.3005
R4524 vdd.n133 vdd.n132 9.3005
R4525 vdd.n144 vdd.n143 9.3005
R4526 vdd.n146 vdd.n145 9.3005
R4527 vdd.n129 vdd.n128 9.3005
R4528 vdd.n152 vdd.n151 9.3005
R4529 vdd.n154 vdd.n153 9.3005
R4530 vdd.n126 vdd.n123 9.3005
R4531 vdd.n161 vdd.n160 9.3005
R4532 vdd.n96 vdd.n95 9.3005
R4533 vdd.n91 vdd.n90 9.3005
R4534 vdd.n102 vdd.n101 9.3005
R4535 vdd.n104 vdd.n103 9.3005
R4536 vdd.n87 vdd.n86 9.3005
R4537 vdd.n110 vdd.n109 9.3005
R4538 vdd.n112 vdd.n111 9.3005
R4539 vdd.n84 vdd.n81 9.3005
R4540 vdd.n119 vdd.n118 9.3005
R4541 vdd.n45 vdd.n44 9.3005
R4542 vdd.n40 vdd.n39 9.3005
R4543 vdd.n51 vdd.n50 9.3005
R4544 vdd.n53 vdd.n52 9.3005
R4545 vdd.n36 vdd.n35 9.3005
R4546 vdd.n59 vdd.n58 9.3005
R4547 vdd.n61 vdd.n60 9.3005
R4548 vdd.n33 vdd.n30 9.3005
R4549 vdd.n68 vdd.n67 9.3005
R4550 vdd.n2854 vdd.n2853 9.3005
R4551 vdd.n2855 vdd.n578 9.3005
R4552 vdd.n577 vdd.n575 9.3005
R4553 vdd.n2861 vdd.n574 9.3005
R4554 vdd.n2862 vdd.n573 9.3005
R4555 vdd.n2863 vdd.n572 9.3005
R4556 vdd.n571 vdd.n569 9.3005
R4557 vdd.n2869 vdd.n568 9.3005
R4558 vdd.n2870 vdd.n567 9.3005
R4559 vdd.n2871 vdd.n566 9.3005
R4560 vdd.n565 vdd.n563 9.3005
R4561 vdd.n2877 vdd.n562 9.3005
R4562 vdd.n2878 vdd.n561 9.3005
R4563 vdd.n2879 vdd.n560 9.3005
R4564 vdd.n559 vdd.n557 9.3005
R4565 vdd.n2885 vdd.n556 9.3005
R4566 vdd.n2886 vdd.n555 9.3005
R4567 vdd.n2887 vdd.n554 9.3005
R4568 vdd.n553 vdd.n551 9.3005
R4569 vdd.n2893 vdd.n550 9.3005
R4570 vdd.n2894 vdd.n549 9.3005
R4571 vdd.n2895 vdd.n548 9.3005
R4572 vdd.n547 vdd.n545 9.3005
R4573 vdd.n2901 vdd.n542 9.3005
R4574 vdd.n2902 vdd.n541 9.3005
R4575 vdd.n2903 vdd.n540 9.3005
R4576 vdd.n539 vdd.n537 9.3005
R4577 vdd.n2909 vdd.n536 9.3005
R4578 vdd.n2910 vdd.n535 9.3005
R4579 vdd.n2911 vdd.n534 9.3005
R4580 vdd.n533 vdd.n531 9.3005
R4581 vdd.n2917 vdd.n530 9.3005
R4582 vdd.n2918 vdd.n529 9.3005
R4583 vdd.n2919 vdd.n528 9.3005
R4584 vdd.n527 vdd.n525 9.3005
R4585 vdd.n2924 vdd.n524 9.3005
R4586 vdd.n2934 vdd.n518 9.3005
R4587 vdd.n2936 vdd.n2935 9.3005
R4588 vdd.n509 vdd.n508 9.3005
R4589 vdd.n2951 vdd.n2950 9.3005
R4590 vdd.n2952 vdd.n507 9.3005
R4591 vdd.n2954 vdd.n2953 9.3005
R4592 vdd.n497 vdd.n496 9.3005
R4593 vdd.n2967 vdd.n2966 9.3005
R4594 vdd.n2968 vdd.n495 9.3005
R4595 vdd.n2970 vdd.n2969 9.3005
R4596 vdd.n485 vdd.n484 9.3005
R4597 vdd.n2984 vdd.n2983 9.3005
R4598 vdd.n2985 vdd.n483 9.3005
R4599 vdd.n2987 vdd.n2986 9.3005
R4600 vdd.n312 vdd.n310 9.3005
R4601 vdd.n2938 vdd.n2937 9.3005
R4602 vdd.n3167 vdd.n3166 9.3005
R4603 vdd.n313 vdd.n311 9.3005
R4604 vdd.n3160 vdd.n320 9.3005
R4605 vdd.n3159 vdd.n321 9.3005
R4606 vdd.n3158 vdd.n322 9.3005
R4607 vdd.n331 vdd.n323 9.3005
R4608 vdd.n3152 vdd.n332 9.3005
R4609 vdd.n3151 vdd.n333 9.3005
R4610 vdd.n3150 vdd.n334 9.3005
R4611 vdd.n342 vdd.n335 9.3005
R4612 vdd.n3144 vdd.n343 9.3005
R4613 vdd.n3143 vdd.n344 9.3005
R4614 vdd.n3142 vdd.n345 9.3005
R4615 vdd.n353 vdd.n346 9.3005
R4616 vdd.n3136 vdd.n3135 9.3005
R4617 vdd.n3132 vdd.n354 9.3005
R4618 vdd.n3131 vdd.n357 9.3005
R4619 vdd.n361 vdd.n358 9.3005
R4620 vdd.n362 vdd.n359 9.3005
R4621 vdd.n3124 vdd.n363 9.3005
R4622 vdd.n3123 vdd.n364 9.3005
R4623 vdd.n3122 vdd.n365 9.3005
R4624 vdd.n369 vdd.n366 9.3005
R4625 vdd.n3117 vdd.n370 9.3005
R4626 vdd.n3116 vdd.n371 9.3005
R4627 vdd.n3115 vdd.n372 9.3005
R4628 vdd.n376 vdd.n373 9.3005
R4629 vdd.n3110 vdd.n377 9.3005
R4630 vdd.n3109 vdd.n378 9.3005
R4631 vdd.n3108 vdd.n379 9.3005
R4632 vdd.n383 vdd.n380 9.3005
R4633 vdd.n3103 vdd.n384 9.3005
R4634 vdd.n3102 vdd.n385 9.3005
R4635 vdd.n3101 vdd.n3100 9.3005
R4636 vdd.n3099 vdd.n386 9.3005
R4637 vdd.n3098 vdd.n3097 9.3005
R4638 vdd.n392 vdd.n391 9.3005
R4639 vdd.n3092 vdd.n396 9.3005
R4640 vdd.n3091 vdd.n397 9.3005
R4641 vdd.n3090 vdd.n398 9.3005
R4642 vdd.n402 vdd.n399 9.3005
R4643 vdd.n3085 vdd.n403 9.3005
R4644 vdd.n3084 vdd.n404 9.3005
R4645 vdd.n3083 vdd.n405 9.3005
R4646 vdd.n409 vdd.n406 9.3005
R4647 vdd.n3078 vdd.n410 9.3005
R4648 vdd.n3077 vdd.n411 9.3005
R4649 vdd.n3076 vdd.n412 9.3005
R4650 vdd.n416 vdd.n413 9.3005
R4651 vdd.n3071 vdd.n417 9.3005
R4652 vdd.n3070 vdd.n418 9.3005
R4653 vdd.n3069 vdd.n419 9.3005
R4654 vdd.n423 vdd.n420 9.3005
R4655 vdd.n3064 vdd.n424 9.3005
R4656 vdd.n3063 vdd.n425 9.3005
R4657 vdd.n3062 vdd.n3061 9.3005
R4658 vdd.n3060 vdd.n426 9.3005
R4659 vdd.n3059 vdd.n3058 9.3005
R4660 vdd.n432 vdd.n431 9.3005
R4661 vdd.n3053 vdd.n436 9.3005
R4662 vdd.n3052 vdd.n437 9.3005
R4663 vdd.n3051 vdd.n438 9.3005
R4664 vdd.n442 vdd.n439 9.3005
R4665 vdd.n3046 vdd.n443 9.3005
R4666 vdd.n3045 vdd.n444 9.3005
R4667 vdd.n3044 vdd.n445 9.3005
R4668 vdd.n449 vdd.n446 9.3005
R4669 vdd.n3039 vdd.n450 9.3005
R4670 vdd.n3038 vdd.n451 9.3005
R4671 vdd.n3037 vdd.n452 9.3005
R4672 vdd.n456 vdd.n453 9.3005
R4673 vdd.n3032 vdd.n457 9.3005
R4674 vdd.n3031 vdd.n458 9.3005
R4675 vdd.n3030 vdd.n459 9.3005
R4676 vdd.n463 vdd.n460 9.3005
R4677 vdd.n3025 vdd.n464 9.3005
R4678 vdd.n3024 vdd.n465 9.3005
R4679 vdd.n3020 vdd.n3017 9.3005
R4680 vdd.n3134 vdd.n3133 9.3005
R4681 vdd.n2944 vdd.n513 9.3005
R4682 vdd.n2946 vdd.n2945 9.3005
R4683 vdd.n503 vdd.n502 9.3005
R4684 vdd.n2959 vdd.n2958 9.3005
R4685 vdd.n2960 vdd.n501 9.3005
R4686 vdd.n2962 vdd.n2961 9.3005
R4687 vdd.n490 vdd.n489 9.3005
R4688 vdd.n2975 vdd.n2974 9.3005
R4689 vdd.n2976 vdd.n488 9.3005
R4690 vdd.n2978 vdd.n2977 9.3005
R4691 vdd.n478 vdd.n477 9.3005
R4692 vdd.n2992 vdd.n2991 9.3005
R4693 vdd.n2993 vdd.n476 9.3005
R4694 vdd.n2995 vdd.n2994 9.3005
R4695 vdd.n2996 vdd.n475 9.3005
R4696 vdd.n2998 vdd.n2997 9.3005
R4697 vdd.n2999 vdd.n474 9.3005
R4698 vdd.n3001 vdd.n3000 9.3005
R4699 vdd.n3002 vdd.n472 9.3005
R4700 vdd.n3004 vdd.n3003 9.3005
R4701 vdd.n3005 vdd.n471 9.3005
R4702 vdd.n3007 vdd.n3006 9.3005
R4703 vdd.n3008 vdd.n469 9.3005
R4704 vdd.n3010 vdd.n3009 9.3005
R4705 vdd.n3011 vdd.n468 9.3005
R4706 vdd.n3013 vdd.n3012 9.3005
R4707 vdd.n3014 vdd.n466 9.3005
R4708 vdd.n3016 vdd.n3015 9.3005
R4709 vdd.n2943 vdd.n2942 9.3005
R4710 vdd.n2807 vdd.n514 9.3005
R4711 vdd.n2812 vdd.n2806 9.3005
R4712 vdd.n2822 vdd.n605 9.3005
R4713 vdd.n2823 vdd.n604 9.3005
R4714 vdd.n603 vdd.n601 9.3005
R4715 vdd.n2829 vdd.n600 9.3005
R4716 vdd.n2830 vdd.n599 9.3005
R4717 vdd.n2831 vdd.n598 9.3005
R4718 vdd.n597 vdd.n595 9.3005
R4719 vdd.n2837 vdd.n594 9.3005
R4720 vdd.n2838 vdd.n593 9.3005
R4721 vdd.n2839 vdd.n592 9.3005
R4722 vdd.n591 vdd.n589 9.3005
R4723 vdd.n2844 vdd.n588 9.3005
R4724 vdd.n2845 vdd.n587 9.3005
R4725 vdd.n583 vdd.n582 9.3005
R4726 vdd.n2851 vdd.n2850 9.3005
R4727 vdd.n2852 vdd.n579 9.3005
R4728 vdd.n2049 vdd.n2048 9.3005
R4729 vdd.n2044 vdd.n895 9.3005
R4730 vdd.n1219 vdd.n979 9.3005
R4731 vdd.n1221 vdd.n1220 9.3005
R4732 vdd.n970 vdd.n969 9.3005
R4733 vdd.n1234 vdd.n1233 9.3005
R4734 vdd.n1235 vdd.n968 9.3005
R4735 vdd.n1237 vdd.n1236 9.3005
R4736 vdd.n957 vdd.n956 9.3005
R4737 vdd.n1250 vdd.n1249 9.3005
R4738 vdd.n1251 vdd.n955 9.3005
R4739 vdd.n1253 vdd.n1252 9.3005
R4740 vdd.n946 vdd.n945 9.3005
R4741 vdd.n1267 vdd.n1266 9.3005
R4742 vdd.n1268 vdd.n944 9.3005
R4743 vdd.n1270 vdd.n1269 9.3005
R4744 vdd.n935 vdd.n934 9.3005
R4745 vdd.n1565 vdd.n1564 9.3005
R4746 vdd.n1566 vdd.n933 9.3005
R4747 vdd.n1568 vdd.n1567 9.3005
R4748 vdd.n923 vdd.n922 9.3005
R4749 vdd.n1582 vdd.n1581 9.3005
R4750 vdd.n1583 vdd.n921 9.3005
R4751 vdd.n1585 vdd.n1584 9.3005
R4752 vdd.n913 vdd.n912 9.3005
R4753 vdd.n1599 vdd.n1598 9.3005
R4754 vdd.n1600 vdd.n910 9.3005
R4755 vdd.n1604 vdd.n1603 9.3005
R4756 vdd.n1602 vdd.n911 9.3005
R4757 vdd.n1601 vdd.n900 9.3005
R4758 vdd.n1218 vdd.n1217 9.3005
R4759 vdd.n1113 vdd.n1103 9.3005
R4760 vdd.n1115 vdd.n1114 9.3005
R4761 vdd.n1116 vdd.n1102 9.3005
R4762 vdd.n1118 vdd.n1117 9.3005
R4763 vdd.n1119 vdd.n1095 9.3005
R4764 vdd.n1121 vdd.n1120 9.3005
R4765 vdd.n1122 vdd.n1094 9.3005
R4766 vdd.n1124 vdd.n1123 9.3005
R4767 vdd.n1125 vdd.n1087 9.3005
R4768 vdd.n1127 vdd.n1126 9.3005
R4769 vdd.n1128 vdd.n1086 9.3005
R4770 vdd.n1130 vdd.n1129 9.3005
R4771 vdd.n1131 vdd.n1079 9.3005
R4772 vdd.n1133 vdd.n1132 9.3005
R4773 vdd.n1134 vdd.n1078 9.3005
R4774 vdd.n1136 vdd.n1135 9.3005
R4775 vdd.n1137 vdd.n1072 9.3005
R4776 vdd.n1139 vdd.n1138 9.3005
R4777 vdd.n1140 vdd.n1070 9.3005
R4778 vdd.n1142 vdd.n1141 9.3005
R4779 vdd.n1071 vdd.n1068 9.3005
R4780 vdd.n1149 vdd.n1064 9.3005
R4781 vdd.n1151 vdd.n1150 9.3005
R4782 vdd.n1152 vdd.n1063 9.3005
R4783 vdd.n1154 vdd.n1153 9.3005
R4784 vdd.n1155 vdd.n1056 9.3005
R4785 vdd.n1157 vdd.n1156 9.3005
R4786 vdd.n1158 vdd.n1055 9.3005
R4787 vdd.n1160 vdd.n1159 9.3005
R4788 vdd.n1161 vdd.n1048 9.3005
R4789 vdd.n1163 vdd.n1162 9.3005
R4790 vdd.n1164 vdd.n1047 9.3005
R4791 vdd.n1166 vdd.n1165 9.3005
R4792 vdd.n1167 vdd.n1040 9.3005
R4793 vdd.n1169 vdd.n1168 9.3005
R4794 vdd.n1170 vdd.n1039 9.3005
R4795 vdd.n1172 vdd.n1171 9.3005
R4796 vdd.n1173 vdd.n1032 9.3005
R4797 vdd.n1175 vdd.n1174 9.3005
R4798 vdd.n1176 vdd.n1031 9.3005
R4799 vdd.n1178 vdd.n1177 9.3005
R4800 vdd.n1179 vdd.n1024 9.3005
R4801 vdd.n1181 vdd.n1180 9.3005
R4802 vdd.n1182 vdd.n1023 9.3005
R4803 vdd.n1184 vdd.n1183 9.3005
R4804 vdd.n1185 vdd.n1014 9.3005
R4805 vdd.n1187 vdd.n1186 9.3005
R4806 vdd.n1188 vdd.n1013 9.3005
R4807 vdd.n1190 vdd.n1189 9.3005
R4808 vdd.n1191 vdd.n1006 9.3005
R4809 vdd.n1193 vdd.n1192 9.3005
R4810 vdd.n1194 vdd.n1005 9.3005
R4811 vdd.n1196 vdd.n1195 9.3005
R4812 vdd.n1197 vdd.n998 9.3005
R4813 vdd.n1199 vdd.n1198 9.3005
R4814 vdd.n1200 vdd.n997 9.3005
R4815 vdd.n1202 vdd.n1201 9.3005
R4816 vdd.n1203 vdd.n990 9.3005
R4817 vdd.n1205 vdd.n1204 9.3005
R4818 vdd.n1206 vdd.n989 9.3005
R4819 vdd.n1208 vdd.n1207 9.3005
R4820 vdd.n1209 vdd.n985 9.3005
R4821 vdd.n1211 vdd.n1210 9.3005
R4822 vdd.n1109 vdd.n980 9.3005
R4823 vdd.n976 vdd.n975 9.3005
R4824 vdd.n1226 vdd.n1225 9.3005
R4825 vdd.n1227 vdd.n974 9.3005
R4826 vdd.n1229 vdd.n1228 9.3005
R4827 vdd.n964 vdd.n963 9.3005
R4828 vdd.n1242 vdd.n1241 9.3005
R4829 vdd.n1243 vdd.n962 9.3005
R4830 vdd.n1245 vdd.n1244 9.3005
R4831 vdd.n952 vdd.n951 9.3005
R4832 vdd.n1259 vdd.n1258 9.3005
R4833 vdd.n1260 vdd.n950 9.3005
R4834 vdd.n1262 vdd.n1261 9.3005
R4835 vdd.n941 vdd.n940 9.3005
R4836 vdd.n1213 vdd.n1212 9.3005
R4837 vdd.n1557 vdd.n1274 9.3005
R4838 vdd.n1478 vdd.n1477 9.3005
R4839 vdd.n1473 vdd.n1472 9.3005
R4840 vdd.n1484 vdd.n1483 9.3005
R4841 vdd.n1486 vdd.n1485 9.3005
R4842 vdd.n1469 vdd.n1468 9.3005
R4843 vdd.n1492 vdd.n1491 9.3005
R4844 vdd.n1494 vdd.n1493 9.3005
R4845 vdd.n1466 vdd.n1463 9.3005
R4846 vdd.n1501 vdd.n1500 9.3005
R4847 vdd.n1529 vdd.n1528 9.3005
R4848 vdd.n1524 vdd.n1523 9.3005
R4849 vdd.n1535 vdd.n1534 9.3005
R4850 vdd.n1537 vdd.n1536 9.3005
R4851 vdd.n1520 vdd.n1519 9.3005
R4852 vdd.n1543 vdd.n1542 9.3005
R4853 vdd.n1545 vdd.n1544 9.3005
R4854 vdd.n1517 vdd.n1514 9.3005
R4855 vdd.n1552 vdd.n1551 9.3005
R4856 vdd.n1384 vdd.n1383 9.3005
R4857 vdd.n1379 vdd.n1378 9.3005
R4858 vdd.n1390 vdd.n1389 9.3005
R4859 vdd.n1392 vdd.n1391 9.3005
R4860 vdd.n1375 vdd.n1374 9.3005
R4861 vdd.n1398 vdd.n1397 9.3005
R4862 vdd.n1400 vdd.n1399 9.3005
R4863 vdd.n1372 vdd.n1369 9.3005
R4864 vdd.n1407 vdd.n1406 9.3005
R4865 vdd.n1435 vdd.n1434 9.3005
R4866 vdd.n1430 vdd.n1429 9.3005
R4867 vdd.n1441 vdd.n1440 9.3005
R4868 vdd.n1443 vdd.n1442 9.3005
R4869 vdd.n1426 vdd.n1425 9.3005
R4870 vdd.n1449 vdd.n1448 9.3005
R4871 vdd.n1451 vdd.n1450 9.3005
R4872 vdd.n1423 vdd.n1420 9.3005
R4873 vdd.n1458 vdd.n1457 9.3005
R4874 vdd.n1291 vdd.n1290 9.3005
R4875 vdd.n1286 vdd.n1285 9.3005
R4876 vdd.n1297 vdd.n1296 9.3005
R4877 vdd.n1299 vdd.n1298 9.3005
R4878 vdd.n1282 vdd.n1281 9.3005
R4879 vdd.n1305 vdd.n1304 9.3005
R4880 vdd.n1307 vdd.n1306 9.3005
R4881 vdd.n1279 vdd.n1276 9.3005
R4882 vdd.n1314 vdd.n1313 9.3005
R4883 vdd.n1342 vdd.n1341 9.3005
R4884 vdd.n1337 vdd.n1336 9.3005
R4885 vdd.n1348 vdd.n1347 9.3005
R4886 vdd.n1350 vdd.n1349 9.3005
R4887 vdd.n1333 vdd.n1332 9.3005
R4888 vdd.n1356 vdd.n1355 9.3005
R4889 vdd.n1358 vdd.n1357 9.3005
R4890 vdd.n1330 vdd.n1327 9.3005
R4891 vdd.n1365 vdd.n1364 9.3005
R4892 vdd.n288 vdd.n287 8.92171
R4893 vdd.n237 vdd.n236 8.92171
R4894 vdd.n194 vdd.n193 8.92171
R4895 vdd.n143 vdd.n142 8.92171
R4896 vdd.n101 vdd.n100 8.92171
R4897 vdd.n50 vdd.n49 8.92171
R4898 vdd.n1483 vdd.n1482 8.92171
R4899 vdd.n1534 vdd.n1533 8.92171
R4900 vdd.n1389 vdd.n1388 8.92171
R4901 vdd.n1440 vdd.n1439 8.92171
R4902 vdd.n1296 vdd.n1295 8.92171
R4903 vdd.n1347 vdd.n1346 8.92171
R4904 vdd.n215 vdd.n121 8.81535
R4905 vdd.n1461 vdd.n1367 8.81535
R4906 vdd.n1596 vdd.t136 8.72962
R4907 vdd.n2956 vdd.t134 8.72962
R4908 vdd.t197 vdd.n1570 8.50289
R4909 vdd.n493 vdd.t146 8.50289
R4910 vdd.n28 vdd.n14 8.42249
R4911 vdd.n1272 vdd.t175 8.27616
R4912 vdd.n3164 vdd.t132 8.27616
R4913 vdd.n3168 vdd.n3167 8.16225
R4914 vdd.n1557 vdd.n1556 8.16225
R4915 vdd.n284 vdd.n278 8.14595
R4916 vdd.n233 vdd.n227 8.14595
R4917 vdd.n190 vdd.n184 8.14595
R4918 vdd.n139 vdd.n133 8.14595
R4919 vdd.n97 vdd.n91 8.14595
R4920 vdd.n46 vdd.n40 8.14595
R4921 vdd.n1479 vdd.n1473 8.14595
R4922 vdd.n1530 vdd.n1524 8.14595
R4923 vdd.n1385 vdd.n1379 8.14595
R4924 vdd.n1436 vdd.n1430 8.14595
R4925 vdd.n1292 vdd.n1286 8.14595
R4926 vdd.n1343 vdd.n1337 8.14595
R4927 vdd.n2635 vdd.n677 8.11757
R4928 vdd.n2109 vdd.n2108 8.11757
R4929 vdd.t144 vdd.n960 8.04943
R4930 vdd.n3155 vdd.t148 8.04943
R4931 vdd.n2087 vdd.n871 7.70933
R4932 vdd.n2093 vdd.n871 7.70933
R4933 vdd.n2099 vdd.n865 7.70933
R4934 vdd.n2099 vdd.n858 7.70933
R4935 vdd.n2105 vdd.n858 7.70933
R4936 vdd.n2105 vdd.n861 7.70933
R4937 vdd.n2112 vdd.n846 7.70933
R4938 vdd.n2118 vdd.n846 7.70933
R4939 vdd.n2124 vdd.n840 7.70933
R4940 vdd.n2130 vdd.n836 7.70933
R4941 vdd.n2136 vdd.n830 7.70933
R4942 vdd.n2148 vdd.n817 7.70933
R4943 vdd.n2154 vdd.n811 7.70933
R4944 vdd.n2154 vdd.n804 7.70933
R4945 vdd.n2162 vdd.n804 7.70933
R4946 vdd.n2169 vdd.t119 7.70933
R4947 vdd.n2244 vdd.t119 7.70933
R4948 vdd.n2576 vdd.t87 7.70933
R4949 vdd.n2582 vdd.t87 7.70933
R4950 vdd.n2588 vdd.n725 7.70933
R4951 vdd.n2594 vdd.n725 7.70933
R4952 vdd.n2594 vdd.n728 7.70933
R4953 vdd.n2600 vdd.n721 7.70933
R4954 vdd.n2612 vdd.n708 7.70933
R4955 vdd.n2618 vdd.n702 7.70933
R4956 vdd.n2624 vdd.n698 7.70933
R4957 vdd.n2630 vdd.n685 7.70933
R4958 vdd.n2638 vdd.n685 7.70933
R4959 vdd.n2644 vdd.n679 7.70933
R4960 vdd.n2644 vdd.n671 7.70933
R4961 vdd.n2695 vdd.n671 7.70933
R4962 vdd.n2695 vdd.n674 7.70933
R4963 vdd.n2701 vdd.n631 7.70933
R4964 vdd.n2771 vdd.n631 7.70933
R4965 vdd.n283 vdd.n280 7.3702
R4966 vdd.n232 vdd.n229 7.3702
R4967 vdd.n189 vdd.n186 7.3702
R4968 vdd.n138 vdd.n135 7.3702
R4969 vdd.n96 vdd.n93 7.3702
R4970 vdd.n45 vdd.n42 7.3702
R4971 vdd.n1478 vdd.n1475 7.3702
R4972 vdd.n1529 vdd.n1526 7.3702
R4973 vdd.n1384 vdd.n1381 7.3702
R4974 vdd.n1435 vdd.n1432 7.3702
R4975 vdd.n1291 vdd.n1288 7.3702
R4976 vdd.n1342 vdd.n1339 7.3702
R4977 vdd.n1239 vdd.t169 7.1425
R4978 vdd.n3148 vdd.t142 7.1425
R4979 vdd.n1150 vdd.n1149 6.98232
R4980 vdd.n1751 vdd.n1750 6.98232
R4981 vdd.n3063 vdd.n3062 6.98232
R4982 vdd.n2855 vdd.n2854 6.98232
R4983 vdd.n1255 vdd.t195 6.91577
R4984 vdd.n325 vdd.t140 6.91577
R4985 vdd.n1562 vdd.t163 6.68904
R4986 vdd.n2989 vdd.t161 6.68904
R4987 vdd.n925 vdd.t214 6.46231
R4988 vdd.t181 vdd.n492 6.46231
R4989 vdd.n3168 vdd.n309 6.27748
R4990 vdd.n1556 vdd.n1555 6.27748
R4991 vdd.n2124 vdd.t81 6.00885
R4992 vdd.n2624 vdd.t113 6.00885
R4993 vdd.n861 vdd.t61 5.89549
R4994 vdd.t30 vdd.n679 5.89549
R4995 vdd.n284 vdd.n283 5.81868
R4996 vdd.n233 vdd.n232 5.81868
R4997 vdd.n190 vdd.n189 5.81868
R4998 vdd.n139 vdd.n138 5.81868
R4999 vdd.n97 vdd.n96 5.81868
R5000 vdd.n46 vdd.n45 5.81868
R5001 vdd.n1479 vdd.n1478 5.81868
R5002 vdd.n1530 vdd.n1529 5.81868
R5003 vdd.n1385 vdd.n1384 5.81868
R5004 vdd.n1436 vdd.n1435 5.81868
R5005 vdd.n1292 vdd.n1291 5.81868
R5006 vdd.n1343 vdd.n1342 5.81868
R5007 vdd.t8 vdd.n865 5.78212
R5008 vdd.n1868 vdd.t43 5.78212
R5009 vdd.n2493 vdd.t51 5.78212
R5010 vdd.n674 vdd.t47 5.78212
R5011 vdd.n2252 vdd.n2251 5.77611
R5012 vdd.n1995 vdd.n1865 5.77611
R5013 vdd.n2506 vdd.n2505 5.77611
R5014 vdd.n2710 vdd.n663 5.77611
R5015 vdd.n2776 vdd.n627 5.77611
R5016 vdd.n2416 vdd.n2356 5.77611
R5017 vdd.n2177 vdd.n795 5.77611
R5018 vdd.n1925 vdd.n1924 5.77611
R5019 vdd.n1112 vdd.n1109 5.62474
R5020 vdd.n2047 vdd.n2044 5.62474
R5021 vdd.n3023 vdd.n3020 5.62474
R5022 vdd.n2810 vdd.n2807 5.62474
R5023 vdd.t98 vdd.n817 5.44203
R5024 vdd.n721 vdd.t103 5.44203
R5025 vdd.t110 vdd.n840 5.10193
R5026 vdd.n830 vdd.t100 5.10193
R5027 vdd.t118 vdd.n708 5.10193
R5028 vdd.n698 vdd.t82 5.10193
R5029 vdd.n287 vdd.n278 5.04292
R5030 vdd.n236 vdd.n227 5.04292
R5031 vdd.n193 vdd.n184 5.04292
R5032 vdd.n142 vdd.n133 5.04292
R5033 vdd.n100 vdd.n91 5.04292
R5034 vdd.n49 vdd.n40 5.04292
R5035 vdd.n1482 vdd.n1473 5.04292
R5036 vdd.n1533 vdd.n1524 5.04292
R5037 vdd.n1388 vdd.n1379 5.04292
R5038 vdd.n1439 vdd.n1430 5.04292
R5039 vdd.n1295 vdd.n1286 5.04292
R5040 vdd.n1346 vdd.n1337 5.04292
R5041 vdd.n1588 vdd.t214 4.8752
R5042 vdd.t117 vdd.t101 4.8752
R5043 vdd.t115 vdd.t85 4.8752
R5044 vdd.t230 vdd.t97 4.8752
R5045 vdd.t79 vdd.t96 4.8752
R5046 vdd.n2964 vdd.t181 4.8752
R5047 vdd.n2253 vdd.n2252 4.83952
R5048 vdd.n1865 vdd.n1861 4.83952
R5049 vdd.n2507 vdd.n2506 4.83952
R5050 vdd.n663 vdd.n658 4.83952
R5051 vdd.n627 vdd.n622 4.83952
R5052 vdd.n2413 vdd.n2356 4.83952
R5053 vdd.n2180 vdd.n795 4.83952
R5054 vdd.n1924 vdd.n1923 4.83952
R5055 vdd.n1719 vdd.n893 4.74817
R5056 vdd.n1714 vdd.n894 4.74817
R5057 vdd.n1616 vdd.n1613 4.74817
R5058 vdd.n2028 vdd.n1617 4.74817
R5059 vdd.n2030 vdd.n1616 4.74817
R5060 vdd.n2029 vdd.n2028 4.74817
R5061 vdd.n521 vdd.n519 4.74817
R5062 vdd.n2925 vdd.n522 4.74817
R5063 vdd.n2928 vdd.n522 4.74817
R5064 vdd.n2929 vdd.n521 4.74817
R5065 vdd.n2817 vdd.n606 4.74817
R5066 vdd.n2813 vdd.n608 4.74817
R5067 vdd.n2816 vdd.n608 4.74817
R5068 vdd.n2821 vdd.n606 4.74817
R5069 vdd.n1715 vdd.n893 4.74817
R5070 vdd.n896 vdd.n894 4.74817
R5071 vdd.n309 vdd.n308 4.7074
R5072 vdd.n215 vdd.n214 4.7074
R5073 vdd.n1555 vdd.n1554 4.7074
R5074 vdd.n1461 vdd.n1460 4.7074
R5075 vdd.t163 vdd.n931 4.64847
R5076 vdd.n2980 vdd.t161 4.64847
R5077 vdd.n2130 vdd.t105 4.53511
R5078 vdd.n2618 vdd.t107 4.53511
R5079 vdd.n1264 vdd.t195 4.42174
R5080 vdd.n3162 vdd.t140 4.42174
R5081 vdd.n2162 vdd.t83 4.30838
R5082 vdd.n2588 vdd.t124 4.30838
R5083 vdd.n288 vdd.n276 4.26717
R5084 vdd.n237 vdd.n225 4.26717
R5085 vdd.n194 vdd.n182 4.26717
R5086 vdd.n143 vdd.n131 4.26717
R5087 vdd.n101 vdd.n89 4.26717
R5088 vdd.n50 vdd.n38 4.26717
R5089 vdd.n1483 vdd.n1471 4.26717
R5090 vdd.n1534 vdd.n1522 4.26717
R5091 vdd.n1389 vdd.n1377 4.26717
R5092 vdd.n1440 vdd.n1428 4.26717
R5093 vdd.n1296 vdd.n1284 4.26717
R5094 vdd.n1347 vdd.n1335 4.26717
R5095 vdd.t169 vdd.n959 4.19501
R5096 vdd.t142 vdd.n329 4.19501
R5097 vdd.n309 vdd.n215 4.10845
R5098 vdd.n1555 vdd.n1461 4.10845
R5099 vdd.n265 vdd.t226 4.06363
R5100 vdd.n265 vdd.t172 4.06363
R5101 vdd.n263 vdd.t177 4.06363
R5102 vdd.n263 vdd.t179 4.06363
R5103 vdd.n261 vdd.t209 4.06363
R5104 vdd.n261 vdd.t157 4.06363
R5105 vdd.n259 vdd.t159 4.06363
R5106 vdd.n259 vdd.t190 4.06363
R5107 vdd.n257 vdd.t192 4.06363
R5108 vdd.n257 vdd.t213 4.06363
R5109 vdd.n171 vdd.t218 4.06363
R5110 vdd.n171 vdd.t165 4.06363
R5111 vdd.n169 vdd.t141 4.06363
R5112 vdd.n169 vdd.t168 4.06363
R5113 vdd.n167 vdd.t200 4.06363
R5114 vdd.n167 vdd.t133 4.06363
R5115 vdd.n165 vdd.t147 4.06363
R5116 vdd.n165 vdd.t180 4.06363
R5117 vdd.n163 vdd.t182 4.06363
R5118 vdd.n163 vdd.t201 4.06363
R5119 vdd.n78 vdd.t149 4.06363
R5120 vdd.n78 vdd.t143 4.06363
R5121 vdd.n76 vdd.t220 4.06363
R5122 vdd.n76 vdd.t207 4.06363
R5123 vdd.n74 vdd.t204 4.06363
R5124 vdd.n74 vdd.t174 4.06363
R5125 vdd.n72 vdd.t222 4.06363
R5126 vdd.n72 vdd.t162 4.06363
R5127 vdd.n70 vdd.t216 4.06363
R5128 vdd.n70 vdd.t184 4.06363
R5129 vdd.n1503 vdd.t160 4.06363
R5130 vdd.n1503 vdd.t225 4.06363
R5131 vdd.n1505 vdd.t219 4.06363
R5132 vdd.n1505 vdd.t208 4.06363
R5133 vdd.n1507 vdd.t187 4.06363
R5134 vdd.n1507 vdd.t158 4.06363
R5135 vdd.n1509 vdd.t227 4.06363
R5136 vdd.n1509 vdd.t206 4.06363
R5137 vdd.n1511 vdd.t202 4.06363
R5138 vdd.n1511 vdd.t171 4.06363
R5139 vdd.n1409 vdd.t151 4.06363
R5140 vdd.n1409 vdd.t215 4.06363
R5141 vdd.n1411 vdd.t210 4.06363
R5142 vdd.n1411 vdd.t198 4.06363
R5143 vdd.n1413 vdd.t178 4.06363
R5144 vdd.n1413 vdd.t139 4.06363
R5145 vdd.n1415 vdd.t223 4.06363
R5146 vdd.n1415 vdd.t196 4.06363
R5147 vdd.n1417 vdd.t193 4.06363
R5148 vdd.n1417 vdd.t145 4.06363
R5149 vdd.n1316 vdd.t185 4.06363
R5150 vdd.n1316 vdd.t217 4.06363
R5151 vdd.n1318 vdd.t164 4.06363
R5152 vdd.n1318 vdd.t205 4.06363
R5153 vdd.n1320 vdd.t176 4.06363
R5154 vdd.n1320 vdd.t211 4.06363
R5155 vdd.n1322 vdd.t189 4.06363
R5156 vdd.n1322 vdd.t221 4.06363
R5157 vdd.n1324 vdd.t170 4.06363
R5158 vdd.n1324 vdd.t152 4.06363
R5159 vdd.n26 vdd.t130 3.9605
R5160 vdd.n26 vdd.t93 3.9605
R5161 vdd.n23 vdd.t127 3.9605
R5162 vdd.n23 vdd.t128 3.9605
R5163 vdd.n21 vdd.t92 3.9605
R5164 vdd.n21 vdd.t89 3.9605
R5165 vdd.n20 vdd.t129 3.9605
R5166 vdd.n20 vdd.t126 3.9605
R5167 vdd.n15 vdd.t91 3.9605
R5168 vdd.n15 vdd.t131 3.9605
R5169 vdd.n16 vdd.t1 3.9605
R5170 vdd.n16 vdd.t2 3.9605
R5171 vdd.n18 vdd.t0 3.9605
R5172 vdd.n18 vdd.t116 3.9605
R5173 vdd.n25 vdd.t90 3.9605
R5174 vdd.n25 vdd.t123 3.9605
R5175 vdd.n7 vdd.t80 3.61217
R5176 vdd.n7 vdd.t108 3.61217
R5177 vdd.n8 vdd.t231 3.61217
R5178 vdd.n8 vdd.t104 3.61217
R5179 vdd.n10 vdd.t88 3.61217
R5180 vdd.n10 vdd.t125 3.61217
R5181 vdd.n12 vdd.t112 3.61217
R5182 vdd.n12 vdd.t95 3.61217
R5183 vdd.n5 vdd.t122 3.61217
R5184 vdd.n5 vdd.t229 3.61217
R5185 vdd.n3 vdd.t84 3.61217
R5186 vdd.n3 vdd.t120 3.61217
R5187 vdd.n1 vdd.t99 3.61217
R5188 vdd.n1 vdd.t86 3.61217
R5189 vdd.n0 vdd.t106 3.61217
R5190 vdd.n0 vdd.t102 3.61217
R5191 vdd.n292 vdd.n291 3.49141
R5192 vdd.n241 vdd.n240 3.49141
R5193 vdd.n198 vdd.n197 3.49141
R5194 vdd.n147 vdd.n146 3.49141
R5195 vdd.n105 vdd.n104 3.49141
R5196 vdd.n54 vdd.n53 3.49141
R5197 vdd.n1487 vdd.n1486 3.49141
R5198 vdd.n1538 vdd.n1537 3.49141
R5199 vdd.n1393 vdd.n1392 3.49141
R5200 vdd.n1444 vdd.n1443 3.49141
R5201 vdd.n1300 vdd.n1299 3.49141
R5202 vdd.n1351 vdd.n1350 3.49141
R5203 vdd.n1868 vdd.t83 3.40145
R5204 vdd.n2316 vdd.t121 3.40145
R5205 vdd.n2569 vdd.t94 3.40145
R5206 vdd.n2493 vdd.t124 3.40145
R5207 vdd.n1247 vdd.t144 3.28809
R5208 vdd.t148 vdd.n3154 3.28809
R5209 vdd.n1969 vdd.t105 3.17472
R5210 vdd.n2472 vdd.t107 3.17472
R5211 vdd.n948 vdd.t175 3.06136
R5212 vdd.t132 vdd.n3163 3.06136
R5213 vdd.n1571 vdd.t197 2.83463
R5214 vdd.n2981 vdd.t146 2.83463
R5215 vdd.n295 vdd.n274 2.71565
R5216 vdd.n244 vdd.n223 2.71565
R5217 vdd.n201 vdd.n180 2.71565
R5218 vdd.n150 vdd.n129 2.71565
R5219 vdd.n108 vdd.n87 2.71565
R5220 vdd.n57 vdd.n36 2.71565
R5221 vdd.n1490 vdd.n1469 2.71565
R5222 vdd.n1541 vdd.n1520 2.71565
R5223 vdd.n1396 vdd.n1375 2.71565
R5224 vdd.n1447 vdd.n1426 2.71565
R5225 vdd.n1303 vdd.n1282 2.71565
R5226 vdd.n1354 vdd.n1333 2.71565
R5227 vdd.n1587 vdd.t136 2.6079
R5228 vdd.n2118 vdd.t110 2.6079
R5229 vdd.n2142 vdd.t100 2.6079
R5230 vdd.n2606 vdd.t118 2.6079
R5231 vdd.n2630 vdd.t82 2.6079
R5232 vdd.t134 vdd.n499 2.6079
R5233 vdd.n2636 vdd.n2635 2.49806
R5234 vdd.n2110 vdd.n2109 2.49806
R5235 vdd.n282 vdd.n281 2.4129
R5236 vdd.n231 vdd.n230 2.4129
R5237 vdd.n188 vdd.n187 2.4129
R5238 vdd.n137 vdd.n136 2.4129
R5239 vdd.n95 vdd.n94 2.4129
R5240 vdd.n44 vdd.n43 2.4129
R5241 vdd.n1477 vdd.n1476 2.4129
R5242 vdd.n1528 vdd.n1527 2.4129
R5243 vdd.n1383 vdd.n1382 2.4129
R5244 vdd.n1434 vdd.n1433 2.4129
R5245 vdd.n1290 vdd.n1289 2.4129
R5246 vdd.n1341 vdd.n1340 2.4129
R5247 vdd.n2027 vdd.n1616 2.27742
R5248 vdd.n2028 vdd.n2027 2.27742
R5249 vdd.n2737 vdd.n522 2.27742
R5250 vdd.n2737 vdd.n521 2.27742
R5251 vdd.n2805 vdd.n608 2.27742
R5252 vdd.n2805 vdd.n606 2.27742
R5253 vdd.n2050 vdd.n893 2.27742
R5254 vdd.n2050 vdd.n894 2.27742
R5255 vdd.n2142 vdd.t98 2.2678
R5256 vdd.n2606 vdd.t103 2.2678
R5257 vdd.t85 vdd.n811 2.04107
R5258 vdd.n728 vdd.t230 2.04107
R5259 vdd.n296 vdd.n272 1.93989
R5260 vdd.n245 vdd.n221 1.93989
R5261 vdd.n202 vdd.n178 1.93989
R5262 vdd.n151 vdd.n127 1.93989
R5263 vdd.n109 vdd.n85 1.93989
R5264 vdd.n58 vdd.n34 1.93989
R5265 vdd.n1491 vdd.n1467 1.93989
R5266 vdd.n1542 vdd.n1518 1.93989
R5267 vdd.n1397 vdd.n1373 1.93989
R5268 vdd.n1448 vdd.n1424 1.93989
R5269 vdd.n1304 vdd.n1280 1.93989
R5270 vdd.n1355 vdd.n1331 1.93989
R5271 vdd.n2093 vdd.t8 1.92771
R5272 vdd.n2169 vdd.t43 1.92771
R5273 vdd.n2582 vdd.t51 1.92771
R5274 vdd.n2701 vdd.t47 1.92771
R5275 vdd.n1969 vdd.t81 1.70098
R5276 vdd.n836 vdd.t117 1.70098
R5277 vdd.t96 vdd.n702 1.70098
R5278 vdd.n2472 vdd.t113 1.70098
R5279 vdd.n983 vdd.t4 1.47425
R5280 vdd.t12 vdd.n3139 1.47425
R5281 vdd.n307 vdd.n267 1.16414
R5282 vdd.n300 vdd.n299 1.16414
R5283 vdd.n256 vdd.n216 1.16414
R5284 vdd.n249 vdd.n248 1.16414
R5285 vdd.n213 vdd.n173 1.16414
R5286 vdd.n206 vdd.n205 1.16414
R5287 vdd.n162 vdd.n122 1.16414
R5288 vdd.n155 vdd.n154 1.16414
R5289 vdd.n120 vdd.n80 1.16414
R5290 vdd.n113 vdd.n112 1.16414
R5291 vdd.n69 vdd.n29 1.16414
R5292 vdd.n62 vdd.n61 1.16414
R5293 vdd.n1502 vdd.n1462 1.16414
R5294 vdd.n1495 vdd.n1494 1.16414
R5295 vdd.n1553 vdd.n1513 1.16414
R5296 vdd.n1546 vdd.n1545 1.16414
R5297 vdd.n1408 vdd.n1368 1.16414
R5298 vdd.n1401 vdd.n1400 1.16414
R5299 vdd.n1459 vdd.n1419 1.16414
R5300 vdd.n1452 vdd.n1451 1.16414
R5301 vdd.n1315 vdd.n1275 1.16414
R5302 vdd.n1308 vdd.n1307 1.16414
R5303 vdd.n1366 vdd.n1326 1.16414
R5304 vdd.n1359 vdd.n1358 1.16414
R5305 vdd.n2136 vdd.t101 1.13415
R5306 vdd.n2612 vdd.t79 1.13415
R5307 vdd.n1579 vdd.t150 1.02079
R5308 vdd.t61 vdd.t109 1.02079
R5309 vdd.t114 vdd.t30 1.02079
R5310 vdd.n2972 vdd.t183 1.02079
R5311 vdd.n1113 vdd.n1112 0.970197
R5312 vdd.n2048 vdd.n2047 0.970197
R5313 vdd.n3024 vdd.n3023 0.970197
R5314 vdd.n2812 vdd.n2810 0.970197
R5315 vdd.n1556 vdd.n28 0.800283
R5316 vdd.t138 vdd.n937 0.794056
R5317 vdd.n1606 vdd.t23 0.794056
R5318 vdd.n2112 vdd.t109 0.794056
R5319 vdd.n2148 vdd.t115 0.794056
R5320 vdd.n2600 vdd.t97 0.794056
R5321 vdd.n2638 vdd.t114 0.794056
R5322 vdd.t16 vdd.n511 0.794056
R5323 vdd.n481 vdd.t199 0.794056
R5324 vdd vdd.n3168 0.79245
R5325 vdd.n1256 vdd.t188 0.567326
R5326 vdd.n3156 vdd.t167 0.567326
R5327 vdd.n2038 vdd.n2037 0.509646
R5328 vdd.n2937 vdd.n2936 0.509646
R5329 vdd.n3135 vdd.n3134 0.509646
R5330 vdd.n3017 vdd.n3016 0.509646
R5331 vdd.n2943 vdd.n514 0.509646
R5332 vdd.n1601 vdd.n895 0.509646
R5333 vdd.n1218 vdd.n980 0.509646
R5334 vdd.n1212 vdd.n1211 0.509646
R5335 vdd.n4 vdd.n2 0.459552
R5336 vdd.n11 vdd.n9 0.459552
R5337 vdd.n305 vdd.n304 0.388379
R5338 vdd.n271 vdd.n269 0.388379
R5339 vdd.n254 vdd.n253 0.388379
R5340 vdd.n220 vdd.n218 0.388379
R5341 vdd.n211 vdd.n210 0.388379
R5342 vdd.n177 vdd.n175 0.388379
R5343 vdd.n160 vdd.n159 0.388379
R5344 vdd.n126 vdd.n124 0.388379
R5345 vdd.n118 vdd.n117 0.388379
R5346 vdd.n84 vdd.n82 0.388379
R5347 vdd.n67 vdd.n66 0.388379
R5348 vdd.n33 vdd.n31 0.388379
R5349 vdd.n1500 vdd.n1499 0.388379
R5350 vdd.n1466 vdd.n1464 0.388379
R5351 vdd.n1551 vdd.n1550 0.388379
R5352 vdd.n1517 vdd.n1515 0.388379
R5353 vdd.n1406 vdd.n1405 0.388379
R5354 vdd.n1372 vdd.n1370 0.388379
R5355 vdd.n1457 vdd.n1456 0.388379
R5356 vdd.n1423 vdd.n1421 0.388379
R5357 vdd.n1313 vdd.n1312 0.388379
R5358 vdd.n1279 vdd.n1277 0.388379
R5359 vdd.n1364 vdd.n1363 0.388379
R5360 vdd.n1330 vdd.n1328 0.388379
R5361 vdd.n19 vdd.n17 0.387128
R5362 vdd.n24 vdd.n22 0.387128
R5363 vdd.n6 vdd.n4 0.358259
R5364 vdd.n13 vdd.n11 0.358259
R5365 vdd.n260 vdd.n258 0.358259
R5366 vdd.n262 vdd.n260 0.358259
R5367 vdd.n264 vdd.n262 0.358259
R5368 vdd.n266 vdd.n264 0.358259
R5369 vdd.n308 vdd.n266 0.358259
R5370 vdd.n166 vdd.n164 0.358259
R5371 vdd.n168 vdd.n166 0.358259
R5372 vdd.n170 vdd.n168 0.358259
R5373 vdd.n172 vdd.n170 0.358259
R5374 vdd.n214 vdd.n172 0.358259
R5375 vdd.n73 vdd.n71 0.358259
R5376 vdd.n75 vdd.n73 0.358259
R5377 vdd.n77 vdd.n75 0.358259
R5378 vdd.n79 vdd.n77 0.358259
R5379 vdd.n121 vdd.n79 0.358259
R5380 vdd.n1554 vdd.n1512 0.358259
R5381 vdd.n1512 vdd.n1510 0.358259
R5382 vdd.n1510 vdd.n1508 0.358259
R5383 vdd.n1508 vdd.n1506 0.358259
R5384 vdd.n1506 vdd.n1504 0.358259
R5385 vdd.n1460 vdd.n1418 0.358259
R5386 vdd.n1418 vdd.n1416 0.358259
R5387 vdd.n1416 vdd.n1414 0.358259
R5388 vdd.n1414 vdd.n1412 0.358259
R5389 vdd.n1412 vdd.n1410 0.358259
R5390 vdd.n1367 vdd.n1325 0.358259
R5391 vdd.n1325 vdd.n1323 0.358259
R5392 vdd.n1323 vdd.n1321 0.358259
R5393 vdd.n1321 vdd.n1319 0.358259
R5394 vdd.n1319 vdd.n1317 0.358259
R5395 vdd.t155 vdd.n966 0.340595
R5396 vdd.n3147 vdd.t153 0.340595
R5397 vdd.n14 vdd.n6 0.334552
R5398 vdd.n14 vdd.n13 0.334552
R5399 vdd.n27 vdd.n19 0.21707
R5400 vdd.n27 vdd.n24 0.21707
R5401 vdd.n306 vdd.n268 0.155672
R5402 vdd.n298 vdd.n268 0.155672
R5403 vdd.n298 vdd.n297 0.155672
R5404 vdd.n297 vdd.n273 0.155672
R5405 vdd.n290 vdd.n273 0.155672
R5406 vdd.n290 vdd.n289 0.155672
R5407 vdd.n289 vdd.n277 0.155672
R5408 vdd.n282 vdd.n277 0.155672
R5409 vdd.n255 vdd.n217 0.155672
R5410 vdd.n247 vdd.n217 0.155672
R5411 vdd.n247 vdd.n246 0.155672
R5412 vdd.n246 vdd.n222 0.155672
R5413 vdd.n239 vdd.n222 0.155672
R5414 vdd.n239 vdd.n238 0.155672
R5415 vdd.n238 vdd.n226 0.155672
R5416 vdd.n231 vdd.n226 0.155672
R5417 vdd.n212 vdd.n174 0.155672
R5418 vdd.n204 vdd.n174 0.155672
R5419 vdd.n204 vdd.n203 0.155672
R5420 vdd.n203 vdd.n179 0.155672
R5421 vdd.n196 vdd.n179 0.155672
R5422 vdd.n196 vdd.n195 0.155672
R5423 vdd.n195 vdd.n183 0.155672
R5424 vdd.n188 vdd.n183 0.155672
R5425 vdd.n161 vdd.n123 0.155672
R5426 vdd.n153 vdd.n123 0.155672
R5427 vdd.n153 vdd.n152 0.155672
R5428 vdd.n152 vdd.n128 0.155672
R5429 vdd.n145 vdd.n128 0.155672
R5430 vdd.n145 vdd.n144 0.155672
R5431 vdd.n144 vdd.n132 0.155672
R5432 vdd.n137 vdd.n132 0.155672
R5433 vdd.n119 vdd.n81 0.155672
R5434 vdd.n111 vdd.n81 0.155672
R5435 vdd.n111 vdd.n110 0.155672
R5436 vdd.n110 vdd.n86 0.155672
R5437 vdd.n103 vdd.n86 0.155672
R5438 vdd.n103 vdd.n102 0.155672
R5439 vdd.n102 vdd.n90 0.155672
R5440 vdd.n95 vdd.n90 0.155672
R5441 vdd.n68 vdd.n30 0.155672
R5442 vdd.n60 vdd.n30 0.155672
R5443 vdd.n60 vdd.n59 0.155672
R5444 vdd.n59 vdd.n35 0.155672
R5445 vdd.n52 vdd.n35 0.155672
R5446 vdd.n52 vdd.n51 0.155672
R5447 vdd.n51 vdd.n39 0.155672
R5448 vdd.n44 vdd.n39 0.155672
R5449 vdd.n1501 vdd.n1463 0.155672
R5450 vdd.n1493 vdd.n1463 0.155672
R5451 vdd.n1493 vdd.n1492 0.155672
R5452 vdd.n1492 vdd.n1468 0.155672
R5453 vdd.n1485 vdd.n1468 0.155672
R5454 vdd.n1485 vdd.n1484 0.155672
R5455 vdd.n1484 vdd.n1472 0.155672
R5456 vdd.n1477 vdd.n1472 0.155672
R5457 vdd.n1552 vdd.n1514 0.155672
R5458 vdd.n1544 vdd.n1514 0.155672
R5459 vdd.n1544 vdd.n1543 0.155672
R5460 vdd.n1543 vdd.n1519 0.155672
R5461 vdd.n1536 vdd.n1519 0.155672
R5462 vdd.n1536 vdd.n1535 0.155672
R5463 vdd.n1535 vdd.n1523 0.155672
R5464 vdd.n1528 vdd.n1523 0.155672
R5465 vdd.n1407 vdd.n1369 0.155672
R5466 vdd.n1399 vdd.n1369 0.155672
R5467 vdd.n1399 vdd.n1398 0.155672
R5468 vdd.n1398 vdd.n1374 0.155672
R5469 vdd.n1391 vdd.n1374 0.155672
R5470 vdd.n1391 vdd.n1390 0.155672
R5471 vdd.n1390 vdd.n1378 0.155672
R5472 vdd.n1383 vdd.n1378 0.155672
R5473 vdd.n1458 vdd.n1420 0.155672
R5474 vdd.n1450 vdd.n1420 0.155672
R5475 vdd.n1450 vdd.n1449 0.155672
R5476 vdd.n1449 vdd.n1425 0.155672
R5477 vdd.n1442 vdd.n1425 0.155672
R5478 vdd.n1442 vdd.n1441 0.155672
R5479 vdd.n1441 vdd.n1429 0.155672
R5480 vdd.n1434 vdd.n1429 0.155672
R5481 vdd.n1314 vdd.n1276 0.155672
R5482 vdd.n1306 vdd.n1276 0.155672
R5483 vdd.n1306 vdd.n1305 0.155672
R5484 vdd.n1305 vdd.n1281 0.155672
R5485 vdd.n1298 vdd.n1281 0.155672
R5486 vdd.n1298 vdd.n1297 0.155672
R5487 vdd.n1297 vdd.n1285 0.155672
R5488 vdd.n1290 vdd.n1285 0.155672
R5489 vdd.n1365 vdd.n1327 0.155672
R5490 vdd.n1357 vdd.n1327 0.155672
R5491 vdd.n1357 vdd.n1356 0.155672
R5492 vdd.n1356 vdd.n1332 0.155672
R5493 vdd.n1349 vdd.n1332 0.155672
R5494 vdd.n1349 vdd.n1348 0.155672
R5495 vdd.n1348 vdd.n1336 0.155672
R5496 vdd.n1341 vdd.n1336 0.155672
R5497 vdd.n1813 vdd.n1618 0.152939
R5498 vdd.n1624 vdd.n1618 0.152939
R5499 vdd.n1625 vdd.n1624 0.152939
R5500 vdd.n1626 vdd.n1625 0.152939
R5501 vdd.n1627 vdd.n1626 0.152939
R5502 vdd.n1631 vdd.n1627 0.152939
R5503 vdd.n1632 vdd.n1631 0.152939
R5504 vdd.n1633 vdd.n1632 0.152939
R5505 vdd.n1634 vdd.n1633 0.152939
R5506 vdd.n1638 vdd.n1634 0.152939
R5507 vdd.n1639 vdd.n1638 0.152939
R5508 vdd.n1640 vdd.n1639 0.152939
R5509 vdd.n1788 vdd.n1640 0.152939
R5510 vdd.n1788 vdd.n1787 0.152939
R5511 vdd.n1787 vdd.n1786 0.152939
R5512 vdd.n1786 vdd.n1646 0.152939
R5513 vdd.n1651 vdd.n1646 0.152939
R5514 vdd.n1652 vdd.n1651 0.152939
R5515 vdd.n1653 vdd.n1652 0.152939
R5516 vdd.n1657 vdd.n1653 0.152939
R5517 vdd.n1658 vdd.n1657 0.152939
R5518 vdd.n1659 vdd.n1658 0.152939
R5519 vdd.n1660 vdd.n1659 0.152939
R5520 vdd.n1664 vdd.n1660 0.152939
R5521 vdd.n1665 vdd.n1664 0.152939
R5522 vdd.n1666 vdd.n1665 0.152939
R5523 vdd.n1667 vdd.n1666 0.152939
R5524 vdd.n1671 vdd.n1667 0.152939
R5525 vdd.n1672 vdd.n1671 0.152939
R5526 vdd.n1673 vdd.n1672 0.152939
R5527 vdd.n1674 vdd.n1673 0.152939
R5528 vdd.n1678 vdd.n1674 0.152939
R5529 vdd.n1679 vdd.n1678 0.152939
R5530 vdd.n1680 vdd.n1679 0.152939
R5531 vdd.n1749 vdd.n1680 0.152939
R5532 vdd.n1749 vdd.n1748 0.152939
R5533 vdd.n1748 vdd.n1747 0.152939
R5534 vdd.n1747 vdd.n1686 0.152939
R5535 vdd.n1691 vdd.n1686 0.152939
R5536 vdd.n1692 vdd.n1691 0.152939
R5537 vdd.n1693 vdd.n1692 0.152939
R5538 vdd.n1697 vdd.n1693 0.152939
R5539 vdd.n1698 vdd.n1697 0.152939
R5540 vdd.n1699 vdd.n1698 0.152939
R5541 vdd.n1700 vdd.n1699 0.152939
R5542 vdd.n1704 vdd.n1700 0.152939
R5543 vdd.n1705 vdd.n1704 0.152939
R5544 vdd.n1706 vdd.n1705 0.152939
R5545 vdd.n1707 vdd.n1706 0.152939
R5546 vdd.n1708 vdd.n1707 0.152939
R5547 vdd.n1708 vdd.n892 0.152939
R5548 vdd.n2037 vdd.n1612 0.152939
R5549 vdd.n1559 vdd.n1558 0.152939
R5550 vdd.n1559 vdd.n928 0.152939
R5551 vdd.n1574 vdd.n928 0.152939
R5552 vdd.n1575 vdd.n1574 0.152939
R5553 vdd.n1576 vdd.n1575 0.152939
R5554 vdd.n1576 vdd.n917 0.152939
R5555 vdd.n1591 vdd.n917 0.152939
R5556 vdd.n1592 vdd.n1591 0.152939
R5557 vdd.n1593 vdd.n1592 0.152939
R5558 vdd.n1593 vdd.n905 0.152939
R5559 vdd.n1610 vdd.n905 0.152939
R5560 vdd.n1611 vdd.n1610 0.152939
R5561 vdd.n2038 vdd.n1611 0.152939
R5562 vdd.n527 vdd.n524 0.152939
R5563 vdd.n528 vdd.n527 0.152939
R5564 vdd.n529 vdd.n528 0.152939
R5565 vdd.n530 vdd.n529 0.152939
R5566 vdd.n533 vdd.n530 0.152939
R5567 vdd.n534 vdd.n533 0.152939
R5568 vdd.n535 vdd.n534 0.152939
R5569 vdd.n536 vdd.n535 0.152939
R5570 vdd.n539 vdd.n536 0.152939
R5571 vdd.n540 vdd.n539 0.152939
R5572 vdd.n541 vdd.n540 0.152939
R5573 vdd.n542 vdd.n541 0.152939
R5574 vdd.n547 vdd.n542 0.152939
R5575 vdd.n548 vdd.n547 0.152939
R5576 vdd.n549 vdd.n548 0.152939
R5577 vdd.n550 vdd.n549 0.152939
R5578 vdd.n553 vdd.n550 0.152939
R5579 vdd.n554 vdd.n553 0.152939
R5580 vdd.n555 vdd.n554 0.152939
R5581 vdd.n556 vdd.n555 0.152939
R5582 vdd.n559 vdd.n556 0.152939
R5583 vdd.n560 vdd.n559 0.152939
R5584 vdd.n561 vdd.n560 0.152939
R5585 vdd.n562 vdd.n561 0.152939
R5586 vdd.n565 vdd.n562 0.152939
R5587 vdd.n566 vdd.n565 0.152939
R5588 vdd.n567 vdd.n566 0.152939
R5589 vdd.n568 vdd.n567 0.152939
R5590 vdd.n571 vdd.n568 0.152939
R5591 vdd.n572 vdd.n571 0.152939
R5592 vdd.n573 vdd.n572 0.152939
R5593 vdd.n574 vdd.n573 0.152939
R5594 vdd.n577 vdd.n574 0.152939
R5595 vdd.n578 vdd.n577 0.152939
R5596 vdd.n2853 vdd.n578 0.152939
R5597 vdd.n2853 vdd.n2852 0.152939
R5598 vdd.n2852 vdd.n2851 0.152939
R5599 vdd.n2851 vdd.n582 0.152939
R5600 vdd.n587 vdd.n582 0.152939
R5601 vdd.n588 vdd.n587 0.152939
R5602 vdd.n591 vdd.n588 0.152939
R5603 vdd.n592 vdd.n591 0.152939
R5604 vdd.n593 vdd.n592 0.152939
R5605 vdd.n594 vdd.n593 0.152939
R5606 vdd.n597 vdd.n594 0.152939
R5607 vdd.n598 vdd.n597 0.152939
R5608 vdd.n599 vdd.n598 0.152939
R5609 vdd.n600 vdd.n599 0.152939
R5610 vdd.n603 vdd.n600 0.152939
R5611 vdd.n604 vdd.n603 0.152939
R5612 vdd.n605 vdd.n604 0.152939
R5613 vdd.n2936 vdd.n518 0.152939
R5614 vdd.n2937 vdd.n508 0.152939
R5615 vdd.n2951 vdd.n508 0.152939
R5616 vdd.n2952 vdd.n2951 0.152939
R5617 vdd.n2953 vdd.n2952 0.152939
R5618 vdd.n2953 vdd.n496 0.152939
R5619 vdd.n2967 vdd.n496 0.152939
R5620 vdd.n2968 vdd.n2967 0.152939
R5621 vdd.n2969 vdd.n2968 0.152939
R5622 vdd.n2969 vdd.n484 0.152939
R5623 vdd.n2984 vdd.n484 0.152939
R5624 vdd.n2985 vdd.n2984 0.152939
R5625 vdd.n2986 vdd.n2985 0.152939
R5626 vdd.n2986 vdd.n310 0.152939
R5627 vdd.n320 vdd.n311 0.152939
R5628 vdd.n321 vdd.n320 0.152939
R5629 vdd.n322 vdd.n321 0.152939
R5630 vdd.n331 vdd.n322 0.152939
R5631 vdd.n332 vdd.n331 0.152939
R5632 vdd.n333 vdd.n332 0.152939
R5633 vdd.n334 vdd.n333 0.152939
R5634 vdd.n342 vdd.n334 0.152939
R5635 vdd.n343 vdd.n342 0.152939
R5636 vdd.n344 vdd.n343 0.152939
R5637 vdd.n345 vdd.n344 0.152939
R5638 vdd.n353 vdd.n345 0.152939
R5639 vdd.n3135 vdd.n353 0.152939
R5640 vdd.n3134 vdd.n354 0.152939
R5641 vdd.n357 vdd.n354 0.152939
R5642 vdd.n361 vdd.n357 0.152939
R5643 vdd.n362 vdd.n361 0.152939
R5644 vdd.n363 vdd.n362 0.152939
R5645 vdd.n364 vdd.n363 0.152939
R5646 vdd.n365 vdd.n364 0.152939
R5647 vdd.n369 vdd.n365 0.152939
R5648 vdd.n370 vdd.n369 0.152939
R5649 vdd.n371 vdd.n370 0.152939
R5650 vdd.n372 vdd.n371 0.152939
R5651 vdd.n376 vdd.n372 0.152939
R5652 vdd.n377 vdd.n376 0.152939
R5653 vdd.n378 vdd.n377 0.152939
R5654 vdd.n379 vdd.n378 0.152939
R5655 vdd.n383 vdd.n379 0.152939
R5656 vdd.n384 vdd.n383 0.152939
R5657 vdd.n385 vdd.n384 0.152939
R5658 vdd.n3100 vdd.n385 0.152939
R5659 vdd.n3100 vdd.n3099 0.152939
R5660 vdd.n3099 vdd.n3098 0.152939
R5661 vdd.n3098 vdd.n391 0.152939
R5662 vdd.n396 vdd.n391 0.152939
R5663 vdd.n397 vdd.n396 0.152939
R5664 vdd.n398 vdd.n397 0.152939
R5665 vdd.n402 vdd.n398 0.152939
R5666 vdd.n403 vdd.n402 0.152939
R5667 vdd.n404 vdd.n403 0.152939
R5668 vdd.n405 vdd.n404 0.152939
R5669 vdd.n409 vdd.n405 0.152939
R5670 vdd.n410 vdd.n409 0.152939
R5671 vdd.n411 vdd.n410 0.152939
R5672 vdd.n412 vdd.n411 0.152939
R5673 vdd.n416 vdd.n412 0.152939
R5674 vdd.n417 vdd.n416 0.152939
R5675 vdd.n418 vdd.n417 0.152939
R5676 vdd.n419 vdd.n418 0.152939
R5677 vdd.n423 vdd.n419 0.152939
R5678 vdd.n424 vdd.n423 0.152939
R5679 vdd.n425 vdd.n424 0.152939
R5680 vdd.n3061 vdd.n425 0.152939
R5681 vdd.n3061 vdd.n3060 0.152939
R5682 vdd.n3060 vdd.n3059 0.152939
R5683 vdd.n3059 vdd.n431 0.152939
R5684 vdd.n436 vdd.n431 0.152939
R5685 vdd.n437 vdd.n436 0.152939
R5686 vdd.n438 vdd.n437 0.152939
R5687 vdd.n442 vdd.n438 0.152939
R5688 vdd.n443 vdd.n442 0.152939
R5689 vdd.n444 vdd.n443 0.152939
R5690 vdd.n445 vdd.n444 0.152939
R5691 vdd.n449 vdd.n445 0.152939
R5692 vdd.n450 vdd.n449 0.152939
R5693 vdd.n451 vdd.n450 0.152939
R5694 vdd.n452 vdd.n451 0.152939
R5695 vdd.n456 vdd.n452 0.152939
R5696 vdd.n457 vdd.n456 0.152939
R5697 vdd.n458 vdd.n457 0.152939
R5698 vdd.n459 vdd.n458 0.152939
R5699 vdd.n463 vdd.n459 0.152939
R5700 vdd.n464 vdd.n463 0.152939
R5701 vdd.n465 vdd.n464 0.152939
R5702 vdd.n3017 vdd.n465 0.152939
R5703 vdd.n2944 vdd.n2943 0.152939
R5704 vdd.n2945 vdd.n2944 0.152939
R5705 vdd.n2945 vdd.n502 0.152939
R5706 vdd.n2959 vdd.n502 0.152939
R5707 vdd.n2960 vdd.n2959 0.152939
R5708 vdd.n2961 vdd.n2960 0.152939
R5709 vdd.n2961 vdd.n489 0.152939
R5710 vdd.n2975 vdd.n489 0.152939
R5711 vdd.n2976 vdd.n2975 0.152939
R5712 vdd.n2977 vdd.n2976 0.152939
R5713 vdd.n2977 vdd.n477 0.152939
R5714 vdd.n2992 vdd.n477 0.152939
R5715 vdd.n2993 vdd.n2992 0.152939
R5716 vdd.n2994 vdd.n2993 0.152939
R5717 vdd.n2994 vdd.n475 0.152939
R5718 vdd.n2998 vdd.n475 0.152939
R5719 vdd.n2999 vdd.n2998 0.152939
R5720 vdd.n3000 vdd.n2999 0.152939
R5721 vdd.n3000 vdd.n472 0.152939
R5722 vdd.n3004 vdd.n472 0.152939
R5723 vdd.n3005 vdd.n3004 0.152939
R5724 vdd.n3006 vdd.n3005 0.152939
R5725 vdd.n3006 vdd.n469 0.152939
R5726 vdd.n3010 vdd.n469 0.152939
R5727 vdd.n3011 vdd.n3010 0.152939
R5728 vdd.n3012 vdd.n3011 0.152939
R5729 vdd.n3012 vdd.n466 0.152939
R5730 vdd.n3016 vdd.n466 0.152939
R5731 vdd.n2806 vdd.n514 0.152939
R5732 vdd.n2049 vdd.n895 0.152939
R5733 vdd.n1219 vdd.n1218 0.152939
R5734 vdd.n1220 vdd.n1219 0.152939
R5735 vdd.n1220 vdd.n969 0.152939
R5736 vdd.n1234 vdd.n969 0.152939
R5737 vdd.n1235 vdd.n1234 0.152939
R5738 vdd.n1236 vdd.n1235 0.152939
R5739 vdd.n1236 vdd.n956 0.152939
R5740 vdd.n1250 vdd.n956 0.152939
R5741 vdd.n1251 vdd.n1250 0.152939
R5742 vdd.n1252 vdd.n1251 0.152939
R5743 vdd.n1252 vdd.n945 0.152939
R5744 vdd.n1267 vdd.n945 0.152939
R5745 vdd.n1268 vdd.n1267 0.152939
R5746 vdd.n1269 vdd.n1268 0.152939
R5747 vdd.n1269 vdd.n934 0.152939
R5748 vdd.n1565 vdd.n934 0.152939
R5749 vdd.n1566 vdd.n1565 0.152939
R5750 vdd.n1567 vdd.n1566 0.152939
R5751 vdd.n1567 vdd.n922 0.152939
R5752 vdd.n1582 vdd.n922 0.152939
R5753 vdd.n1583 vdd.n1582 0.152939
R5754 vdd.n1584 vdd.n1583 0.152939
R5755 vdd.n1584 vdd.n912 0.152939
R5756 vdd.n1599 vdd.n912 0.152939
R5757 vdd.n1600 vdd.n1599 0.152939
R5758 vdd.n1603 vdd.n1600 0.152939
R5759 vdd.n1603 vdd.n1602 0.152939
R5760 vdd.n1602 vdd.n1601 0.152939
R5761 vdd.n1211 vdd.n985 0.152939
R5762 vdd.n1207 vdd.n985 0.152939
R5763 vdd.n1207 vdd.n1206 0.152939
R5764 vdd.n1206 vdd.n1205 0.152939
R5765 vdd.n1205 vdd.n990 0.152939
R5766 vdd.n1201 vdd.n990 0.152939
R5767 vdd.n1201 vdd.n1200 0.152939
R5768 vdd.n1200 vdd.n1199 0.152939
R5769 vdd.n1199 vdd.n998 0.152939
R5770 vdd.n1195 vdd.n998 0.152939
R5771 vdd.n1195 vdd.n1194 0.152939
R5772 vdd.n1194 vdd.n1193 0.152939
R5773 vdd.n1193 vdd.n1006 0.152939
R5774 vdd.n1189 vdd.n1006 0.152939
R5775 vdd.n1189 vdd.n1188 0.152939
R5776 vdd.n1188 vdd.n1187 0.152939
R5777 vdd.n1187 vdd.n1014 0.152939
R5778 vdd.n1183 vdd.n1014 0.152939
R5779 vdd.n1183 vdd.n1182 0.152939
R5780 vdd.n1182 vdd.n1181 0.152939
R5781 vdd.n1181 vdd.n1024 0.152939
R5782 vdd.n1177 vdd.n1024 0.152939
R5783 vdd.n1177 vdd.n1176 0.152939
R5784 vdd.n1176 vdd.n1175 0.152939
R5785 vdd.n1175 vdd.n1032 0.152939
R5786 vdd.n1171 vdd.n1032 0.152939
R5787 vdd.n1171 vdd.n1170 0.152939
R5788 vdd.n1170 vdd.n1169 0.152939
R5789 vdd.n1169 vdd.n1040 0.152939
R5790 vdd.n1165 vdd.n1040 0.152939
R5791 vdd.n1165 vdd.n1164 0.152939
R5792 vdd.n1164 vdd.n1163 0.152939
R5793 vdd.n1163 vdd.n1048 0.152939
R5794 vdd.n1159 vdd.n1048 0.152939
R5795 vdd.n1159 vdd.n1158 0.152939
R5796 vdd.n1158 vdd.n1157 0.152939
R5797 vdd.n1157 vdd.n1056 0.152939
R5798 vdd.n1153 vdd.n1056 0.152939
R5799 vdd.n1153 vdd.n1152 0.152939
R5800 vdd.n1152 vdd.n1151 0.152939
R5801 vdd.n1151 vdd.n1064 0.152939
R5802 vdd.n1071 vdd.n1064 0.152939
R5803 vdd.n1141 vdd.n1071 0.152939
R5804 vdd.n1141 vdd.n1140 0.152939
R5805 vdd.n1140 vdd.n1139 0.152939
R5806 vdd.n1139 vdd.n1072 0.152939
R5807 vdd.n1135 vdd.n1072 0.152939
R5808 vdd.n1135 vdd.n1134 0.152939
R5809 vdd.n1134 vdd.n1133 0.152939
R5810 vdd.n1133 vdd.n1079 0.152939
R5811 vdd.n1129 vdd.n1079 0.152939
R5812 vdd.n1129 vdd.n1128 0.152939
R5813 vdd.n1128 vdd.n1127 0.152939
R5814 vdd.n1127 vdd.n1087 0.152939
R5815 vdd.n1123 vdd.n1087 0.152939
R5816 vdd.n1123 vdd.n1122 0.152939
R5817 vdd.n1122 vdd.n1121 0.152939
R5818 vdd.n1121 vdd.n1095 0.152939
R5819 vdd.n1117 vdd.n1095 0.152939
R5820 vdd.n1117 vdd.n1116 0.152939
R5821 vdd.n1116 vdd.n1115 0.152939
R5822 vdd.n1115 vdd.n1103 0.152939
R5823 vdd.n1103 vdd.n980 0.152939
R5824 vdd.n1212 vdd.n975 0.152939
R5825 vdd.n1226 vdd.n975 0.152939
R5826 vdd.n1227 vdd.n1226 0.152939
R5827 vdd.n1228 vdd.n1227 0.152939
R5828 vdd.n1228 vdd.n963 0.152939
R5829 vdd.n1242 vdd.n963 0.152939
R5830 vdd.n1243 vdd.n1242 0.152939
R5831 vdd.n1244 vdd.n1243 0.152939
R5832 vdd.n1244 vdd.n951 0.152939
R5833 vdd.n1259 vdd.n951 0.152939
R5834 vdd.n1260 vdd.n1259 0.152939
R5835 vdd.n1261 vdd.n1260 0.152939
R5836 vdd.n1261 vdd.n940 0.152939
R5837 vdd.n1558 vdd.n1557 0.145814
R5838 vdd.n3167 vdd.n310 0.145814
R5839 vdd.n3167 vdd.n311 0.145814
R5840 vdd.n1557 vdd.n940 0.145814
R5841 vdd.n2027 vdd.n1612 0.110256
R5842 vdd.n2737 vdd.n518 0.110256
R5843 vdd.n2806 vdd.n2805 0.110256
R5844 vdd.n2050 vdd.n2049 0.110256
R5845 vdd.n2027 vdd.n1813 0.0431829
R5846 vdd.n2050 vdd.n892 0.0431829
R5847 vdd.n2737 vdd.n524 0.0431829
R5848 vdd.n2805 vdd.n605 0.0431829
R5849 vdd vdd.n28 0.00833333
R5850 CSoutput.n19 CSoutput.t209 184.661
R5851 CSoutput.n78 CSoutput.n77 165.8
R5852 CSoutput.n76 CSoutput.n0 165.8
R5853 CSoutput.n75 CSoutput.n74 165.8
R5854 CSoutput.n73 CSoutput.n72 165.8
R5855 CSoutput.n71 CSoutput.n2 165.8
R5856 CSoutput.n69 CSoutput.n68 165.8
R5857 CSoutput.n67 CSoutput.n3 165.8
R5858 CSoutput.n66 CSoutput.n65 165.8
R5859 CSoutput.n63 CSoutput.n4 165.8
R5860 CSoutput.n61 CSoutput.n60 165.8
R5861 CSoutput.n59 CSoutput.n5 165.8
R5862 CSoutput.n58 CSoutput.n57 165.8
R5863 CSoutput.n55 CSoutput.n6 165.8
R5864 CSoutput.n54 CSoutput.n53 165.8
R5865 CSoutput.n52 CSoutput.n51 165.8
R5866 CSoutput.n50 CSoutput.n8 165.8
R5867 CSoutput.n48 CSoutput.n47 165.8
R5868 CSoutput.n46 CSoutput.n9 165.8
R5869 CSoutput.n45 CSoutput.n44 165.8
R5870 CSoutput.n42 CSoutput.n10 165.8
R5871 CSoutput.n41 CSoutput.n40 165.8
R5872 CSoutput.n39 CSoutput.n38 165.8
R5873 CSoutput.n37 CSoutput.n12 165.8
R5874 CSoutput.n35 CSoutput.n34 165.8
R5875 CSoutput.n33 CSoutput.n13 165.8
R5876 CSoutput.n32 CSoutput.n31 165.8
R5877 CSoutput.n29 CSoutput.n14 165.8
R5878 CSoutput.n28 CSoutput.n27 165.8
R5879 CSoutput.n26 CSoutput.n25 165.8
R5880 CSoutput.n24 CSoutput.n16 165.8
R5881 CSoutput.n22 CSoutput.n21 165.8
R5882 CSoutput.n20 CSoutput.n17 165.8
R5883 CSoutput.n77 CSoutput.t212 162.194
R5884 CSoutput.n18 CSoutput.t205 120.501
R5885 CSoutput.n23 CSoutput.t198 120.501
R5886 CSoutput.n15 CSoutput.t193 120.501
R5887 CSoutput.n30 CSoutput.t207 120.501
R5888 CSoutput.n36 CSoutput.t208 120.501
R5889 CSoutput.n11 CSoutput.t195 120.501
R5890 CSoutput.n43 CSoutput.t192 120.501
R5891 CSoutput.n49 CSoutput.t211 120.501
R5892 CSoutput.n7 CSoutput.t199 120.501
R5893 CSoutput.n56 CSoutput.t202 120.501
R5894 CSoutput.n62 CSoutput.t213 120.501
R5895 CSoutput.n64 CSoutput.t203 120.501
R5896 CSoutput.n70 CSoutput.t204 120.501
R5897 CSoutput.n1 CSoutput.t197 120.501
R5898 CSoutput.n290 CSoutput.n288 103.469
R5899 CSoutput.n278 CSoutput.n276 103.469
R5900 CSoutput.n267 CSoutput.n265 103.469
R5901 CSoutput.n104 CSoutput.n102 103.469
R5902 CSoutput.n92 CSoutput.n90 103.469
R5903 CSoutput.n81 CSoutput.n79 103.469
R5904 CSoutput.n296 CSoutput.n295 103.111
R5905 CSoutput.n294 CSoutput.n293 103.111
R5906 CSoutput.n292 CSoutput.n291 103.111
R5907 CSoutput.n290 CSoutput.n289 103.111
R5908 CSoutput.n286 CSoutput.n285 103.111
R5909 CSoutput.n284 CSoutput.n283 103.111
R5910 CSoutput.n282 CSoutput.n281 103.111
R5911 CSoutput.n280 CSoutput.n279 103.111
R5912 CSoutput.n278 CSoutput.n277 103.111
R5913 CSoutput.n275 CSoutput.n274 103.111
R5914 CSoutput.n273 CSoutput.n272 103.111
R5915 CSoutput.n271 CSoutput.n270 103.111
R5916 CSoutput.n269 CSoutput.n268 103.111
R5917 CSoutput.n267 CSoutput.n266 103.111
R5918 CSoutput.n104 CSoutput.n103 103.111
R5919 CSoutput.n106 CSoutput.n105 103.111
R5920 CSoutput.n108 CSoutput.n107 103.111
R5921 CSoutput.n110 CSoutput.n109 103.111
R5922 CSoutput.n112 CSoutput.n111 103.111
R5923 CSoutput.n92 CSoutput.n91 103.111
R5924 CSoutput.n94 CSoutput.n93 103.111
R5925 CSoutput.n96 CSoutput.n95 103.111
R5926 CSoutput.n98 CSoutput.n97 103.111
R5927 CSoutput.n100 CSoutput.n99 103.111
R5928 CSoutput.n81 CSoutput.n80 103.111
R5929 CSoutput.n83 CSoutput.n82 103.111
R5930 CSoutput.n85 CSoutput.n84 103.111
R5931 CSoutput.n87 CSoutput.n86 103.111
R5932 CSoutput.n89 CSoutput.n88 103.111
R5933 CSoutput.n298 CSoutput.n297 103.111
R5934 CSoutput.n342 CSoutput.n340 81.5057
R5935 CSoutput.n322 CSoutput.n320 81.5057
R5936 CSoutput.n303 CSoutput.n301 81.5057
R5937 CSoutput.n402 CSoutput.n400 81.5057
R5938 CSoutput.n382 CSoutput.n380 81.5057
R5939 CSoutput.n363 CSoutput.n361 81.5057
R5940 CSoutput.n358 CSoutput.n357 80.9324
R5941 CSoutput.n356 CSoutput.n355 80.9324
R5942 CSoutput.n354 CSoutput.n353 80.9324
R5943 CSoutput.n352 CSoutput.n351 80.9324
R5944 CSoutput.n350 CSoutput.n349 80.9324
R5945 CSoutput.n348 CSoutput.n347 80.9324
R5946 CSoutput.n346 CSoutput.n345 80.9324
R5947 CSoutput.n344 CSoutput.n343 80.9324
R5948 CSoutput.n342 CSoutput.n341 80.9324
R5949 CSoutput.n338 CSoutput.n337 80.9324
R5950 CSoutput.n336 CSoutput.n335 80.9324
R5951 CSoutput.n334 CSoutput.n333 80.9324
R5952 CSoutput.n332 CSoutput.n331 80.9324
R5953 CSoutput.n330 CSoutput.n329 80.9324
R5954 CSoutput.n328 CSoutput.n327 80.9324
R5955 CSoutput.n326 CSoutput.n325 80.9324
R5956 CSoutput.n324 CSoutput.n323 80.9324
R5957 CSoutput.n322 CSoutput.n321 80.9324
R5958 CSoutput.n319 CSoutput.n318 80.9324
R5959 CSoutput.n317 CSoutput.n316 80.9324
R5960 CSoutput.n315 CSoutput.n314 80.9324
R5961 CSoutput.n313 CSoutput.n312 80.9324
R5962 CSoutput.n311 CSoutput.n310 80.9324
R5963 CSoutput.n309 CSoutput.n308 80.9324
R5964 CSoutput.n307 CSoutput.n306 80.9324
R5965 CSoutput.n305 CSoutput.n304 80.9324
R5966 CSoutput.n303 CSoutput.n302 80.9324
R5967 CSoutput.n402 CSoutput.n401 80.9324
R5968 CSoutput.n404 CSoutput.n403 80.9324
R5969 CSoutput.n406 CSoutput.n405 80.9324
R5970 CSoutput.n408 CSoutput.n407 80.9324
R5971 CSoutput.n410 CSoutput.n409 80.9324
R5972 CSoutput.n412 CSoutput.n411 80.9324
R5973 CSoutput.n414 CSoutput.n413 80.9324
R5974 CSoutput.n416 CSoutput.n415 80.9324
R5975 CSoutput.n418 CSoutput.n417 80.9324
R5976 CSoutput.n382 CSoutput.n381 80.9324
R5977 CSoutput.n384 CSoutput.n383 80.9324
R5978 CSoutput.n386 CSoutput.n385 80.9324
R5979 CSoutput.n388 CSoutput.n387 80.9324
R5980 CSoutput.n390 CSoutput.n389 80.9324
R5981 CSoutput.n392 CSoutput.n391 80.9324
R5982 CSoutput.n394 CSoutput.n393 80.9324
R5983 CSoutput.n396 CSoutput.n395 80.9324
R5984 CSoutput.n398 CSoutput.n397 80.9324
R5985 CSoutput.n363 CSoutput.n362 80.9324
R5986 CSoutput.n365 CSoutput.n364 80.9324
R5987 CSoutput.n367 CSoutput.n366 80.9324
R5988 CSoutput.n369 CSoutput.n368 80.9324
R5989 CSoutput.n371 CSoutput.n370 80.9324
R5990 CSoutput.n373 CSoutput.n372 80.9324
R5991 CSoutput.n375 CSoutput.n374 80.9324
R5992 CSoutput.n377 CSoutput.n376 80.9324
R5993 CSoutput.n379 CSoutput.n378 80.9324
R5994 CSoutput.n25 CSoutput.n24 48.1486
R5995 CSoutput.n69 CSoutput.n3 48.1486
R5996 CSoutput.n38 CSoutput.n37 48.1486
R5997 CSoutput.n42 CSoutput.n41 48.1486
R5998 CSoutput.n51 CSoutput.n50 48.1486
R5999 CSoutput.n55 CSoutput.n54 48.1486
R6000 CSoutput.n22 CSoutput.n17 46.462
R6001 CSoutput.n72 CSoutput.n71 46.462
R6002 CSoutput.n20 CSoutput.n19 44.9055
R6003 CSoutput.n29 CSoutput.n28 43.7635
R6004 CSoutput.n65 CSoutput.n63 43.7635
R6005 CSoutput.n35 CSoutput.n13 41.7396
R6006 CSoutput.n57 CSoutput.n5 41.7396
R6007 CSoutput.n44 CSoutput.n9 37.0171
R6008 CSoutput.n48 CSoutput.n9 37.0171
R6009 CSoutput.n76 CSoutput.n75 34.9932
R6010 CSoutput.n31 CSoutput.n13 32.2947
R6011 CSoutput.n61 CSoutput.n5 32.2947
R6012 CSoutput.n30 CSoutput.n29 29.6014
R6013 CSoutput.n63 CSoutput.n62 29.6014
R6014 CSoutput.n19 CSoutput.n18 28.4085
R6015 CSoutput.n18 CSoutput.n17 25.1176
R6016 CSoutput.n72 CSoutput.n1 25.1176
R6017 CSoutput.n43 CSoutput.n42 22.0922
R6018 CSoutput.n50 CSoutput.n49 22.0922
R6019 CSoutput.n77 CSoutput.n76 21.8586
R6020 CSoutput.n37 CSoutput.n36 18.9681
R6021 CSoutput.n56 CSoutput.n55 18.9681
R6022 CSoutput.n25 CSoutput.n15 17.6292
R6023 CSoutput.n64 CSoutput.n3 17.6292
R6024 CSoutput.n24 CSoutput.n23 15.844
R6025 CSoutput.n70 CSoutput.n69 15.844
R6026 CSoutput.n38 CSoutput.n11 14.5051
R6027 CSoutput.n54 CSoutput.n7 14.5051
R6028 CSoutput.n421 CSoutput.n78 11.4982
R6029 CSoutput.n41 CSoutput.n11 11.3811
R6030 CSoutput.n51 CSoutput.n7 11.3811
R6031 CSoutput.n23 CSoutput.n22 10.0422
R6032 CSoutput.n71 CSoutput.n70 10.0422
R6033 CSoutput.n360 CSoutput.n300 9.30273
R6034 CSoutput.n287 CSoutput.n275 9.25285
R6035 CSoutput.n101 CSoutput.n89 9.25285
R6036 CSoutput.n339 CSoutput.n319 8.98182
R6037 CSoutput.n399 CSoutput.n379 8.98182
R6038 CSoutput.n28 CSoutput.n15 8.25698
R6039 CSoutput.n65 CSoutput.n64 8.25698
R6040 CSoutput.n300 CSoutput.n299 7.12641
R6041 CSoutput.n114 CSoutput.n113 7.12641
R6042 CSoutput.n36 CSoutput.n35 6.91809
R6043 CSoutput.n57 CSoutput.n56 6.91809
R6044 CSoutput.n360 CSoutput.n359 6.02792
R6045 CSoutput.n420 CSoutput.n419 6.02792
R6046 CSoutput.n421 CSoutput.n114 5.71029
R6047 CSoutput.n359 CSoutput.n358 5.25266
R6048 CSoutput.n339 CSoutput.n338 5.25266
R6049 CSoutput.n419 CSoutput.n418 5.25266
R6050 CSoutput.n399 CSoutput.n398 5.25266
R6051 CSoutput.n299 CSoutput.n298 5.1449
R6052 CSoutput.n287 CSoutput.n286 5.1449
R6053 CSoutput.n113 CSoutput.n112 5.1449
R6054 CSoutput.n101 CSoutput.n100 5.1449
R6055 CSoutput.n205 CSoutput.n158 4.5005
R6056 CSoutput.n174 CSoutput.n158 4.5005
R6057 CSoutput.n169 CSoutput.n153 4.5005
R6058 CSoutput.n169 CSoutput.n155 4.5005
R6059 CSoutput.n169 CSoutput.n152 4.5005
R6060 CSoutput.n169 CSoutput.n156 4.5005
R6061 CSoutput.n169 CSoutput.n151 4.5005
R6062 CSoutput.n169 CSoutput.t196 4.5005
R6063 CSoutput.n169 CSoutput.n150 4.5005
R6064 CSoutput.n169 CSoutput.n157 4.5005
R6065 CSoutput.n169 CSoutput.n158 4.5005
R6066 CSoutput.n167 CSoutput.n153 4.5005
R6067 CSoutput.n167 CSoutput.n155 4.5005
R6068 CSoutput.n167 CSoutput.n152 4.5005
R6069 CSoutput.n167 CSoutput.n156 4.5005
R6070 CSoutput.n167 CSoutput.n151 4.5005
R6071 CSoutput.n167 CSoutput.t196 4.5005
R6072 CSoutput.n167 CSoutput.n150 4.5005
R6073 CSoutput.n167 CSoutput.n157 4.5005
R6074 CSoutput.n167 CSoutput.n158 4.5005
R6075 CSoutput.n166 CSoutput.n153 4.5005
R6076 CSoutput.n166 CSoutput.n155 4.5005
R6077 CSoutput.n166 CSoutput.n152 4.5005
R6078 CSoutput.n166 CSoutput.n156 4.5005
R6079 CSoutput.n166 CSoutput.n151 4.5005
R6080 CSoutput.n166 CSoutput.t196 4.5005
R6081 CSoutput.n166 CSoutput.n150 4.5005
R6082 CSoutput.n166 CSoutput.n157 4.5005
R6083 CSoutput.n166 CSoutput.n158 4.5005
R6084 CSoutput.n251 CSoutput.n153 4.5005
R6085 CSoutput.n251 CSoutput.n155 4.5005
R6086 CSoutput.n251 CSoutput.n152 4.5005
R6087 CSoutput.n251 CSoutput.n156 4.5005
R6088 CSoutput.n251 CSoutput.n151 4.5005
R6089 CSoutput.n251 CSoutput.t196 4.5005
R6090 CSoutput.n251 CSoutput.n150 4.5005
R6091 CSoutput.n251 CSoutput.n157 4.5005
R6092 CSoutput.n251 CSoutput.n158 4.5005
R6093 CSoutput.n249 CSoutput.n153 4.5005
R6094 CSoutput.n249 CSoutput.n155 4.5005
R6095 CSoutput.n249 CSoutput.n152 4.5005
R6096 CSoutput.n249 CSoutput.n156 4.5005
R6097 CSoutput.n249 CSoutput.n151 4.5005
R6098 CSoutput.n249 CSoutput.t196 4.5005
R6099 CSoutput.n249 CSoutput.n150 4.5005
R6100 CSoutput.n249 CSoutput.n157 4.5005
R6101 CSoutput.n247 CSoutput.n153 4.5005
R6102 CSoutput.n247 CSoutput.n155 4.5005
R6103 CSoutput.n247 CSoutput.n152 4.5005
R6104 CSoutput.n247 CSoutput.n156 4.5005
R6105 CSoutput.n247 CSoutput.n151 4.5005
R6106 CSoutput.n247 CSoutput.t196 4.5005
R6107 CSoutput.n247 CSoutput.n150 4.5005
R6108 CSoutput.n247 CSoutput.n157 4.5005
R6109 CSoutput.n177 CSoutput.n153 4.5005
R6110 CSoutput.n177 CSoutput.n155 4.5005
R6111 CSoutput.n177 CSoutput.n152 4.5005
R6112 CSoutput.n177 CSoutput.n156 4.5005
R6113 CSoutput.n177 CSoutput.n151 4.5005
R6114 CSoutput.n177 CSoutput.t196 4.5005
R6115 CSoutput.n177 CSoutput.n150 4.5005
R6116 CSoutput.n177 CSoutput.n157 4.5005
R6117 CSoutput.n177 CSoutput.n158 4.5005
R6118 CSoutput.n176 CSoutput.n153 4.5005
R6119 CSoutput.n176 CSoutput.n155 4.5005
R6120 CSoutput.n176 CSoutput.n152 4.5005
R6121 CSoutput.n176 CSoutput.n156 4.5005
R6122 CSoutput.n176 CSoutput.n151 4.5005
R6123 CSoutput.n176 CSoutput.t196 4.5005
R6124 CSoutput.n176 CSoutput.n150 4.5005
R6125 CSoutput.n176 CSoutput.n157 4.5005
R6126 CSoutput.n176 CSoutput.n158 4.5005
R6127 CSoutput.n180 CSoutput.n153 4.5005
R6128 CSoutput.n180 CSoutput.n155 4.5005
R6129 CSoutput.n180 CSoutput.n152 4.5005
R6130 CSoutput.n180 CSoutput.n156 4.5005
R6131 CSoutput.n180 CSoutput.n151 4.5005
R6132 CSoutput.n180 CSoutput.t196 4.5005
R6133 CSoutput.n180 CSoutput.n150 4.5005
R6134 CSoutput.n180 CSoutput.n157 4.5005
R6135 CSoutput.n180 CSoutput.n158 4.5005
R6136 CSoutput.n179 CSoutput.n153 4.5005
R6137 CSoutput.n179 CSoutput.n155 4.5005
R6138 CSoutput.n179 CSoutput.n152 4.5005
R6139 CSoutput.n179 CSoutput.n156 4.5005
R6140 CSoutput.n179 CSoutput.n151 4.5005
R6141 CSoutput.n179 CSoutput.t196 4.5005
R6142 CSoutput.n179 CSoutput.n150 4.5005
R6143 CSoutput.n179 CSoutput.n157 4.5005
R6144 CSoutput.n179 CSoutput.n158 4.5005
R6145 CSoutput.n162 CSoutput.n153 4.5005
R6146 CSoutput.n162 CSoutput.n155 4.5005
R6147 CSoutput.n162 CSoutput.n152 4.5005
R6148 CSoutput.n162 CSoutput.n156 4.5005
R6149 CSoutput.n162 CSoutput.n151 4.5005
R6150 CSoutput.n162 CSoutput.t196 4.5005
R6151 CSoutput.n162 CSoutput.n150 4.5005
R6152 CSoutput.n162 CSoutput.n157 4.5005
R6153 CSoutput.n162 CSoutput.n158 4.5005
R6154 CSoutput.n254 CSoutput.n153 4.5005
R6155 CSoutput.n254 CSoutput.n155 4.5005
R6156 CSoutput.n254 CSoutput.n152 4.5005
R6157 CSoutput.n254 CSoutput.n156 4.5005
R6158 CSoutput.n254 CSoutput.n151 4.5005
R6159 CSoutput.n254 CSoutput.t196 4.5005
R6160 CSoutput.n254 CSoutput.n150 4.5005
R6161 CSoutput.n254 CSoutput.n157 4.5005
R6162 CSoutput.n254 CSoutput.n158 4.5005
R6163 CSoutput.n241 CSoutput.n212 4.5005
R6164 CSoutput.n241 CSoutput.n218 4.5005
R6165 CSoutput.n199 CSoutput.n188 4.5005
R6166 CSoutput.n199 CSoutput.n190 4.5005
R6167 CSoutput.n199 CSoutput.n187 4.5005
R6168 CSoutput.n199 CSoutput.n191 4.5005
R6169 CSoutput.n199 CSoutput.n186 4.5005
R6170 CSoutput.n199 CSoutput.t200 4.5005
R6171 CSoutput.n199 CSoutput.n185 4.5005
R6172 CSoutput.n199 CSoutput.n192 4.5005
R6173 CSoutput.n241 CSoutput.n199 4.5005
R6174 CSoutput.n220 CSoutput.n188 4.5005
R6175 CSoutput.n220 CSoutput.n190 4.5005
R6176 CSoutput.n220 CSoutput.n187 4.5005
R6177 CSoutput.n220 CSoutput.n191 4.5005
R6178 CSoutput.n220 CSoutput.n186 4.5005
R6179 CSoutput.n220 CSoutput.t200 4.5005
R6180 CSoutput.n220 CSoutput.n185 4.5005
R6181 CSoutput.n220 CSoutput.n192 4.5005
R6182 CSoutput.n241 CSoutput.n220 4.5005
R6183 CSoutput.n198 CSoutput.n188 4.5005
R6184 CSoutput.n198 CSoutput.n190 4.5005
R6185 CSoutput.n198 CSoutput.n187 4.5005
R6186 CSoutput.n198 CSoutput.n191 4.5005
R6187 CSoutput.n198 CSoutput.n186 4.5005
R6188 CSoutput.n198 CSoutput.t200 4.5005
R6189 CSoutput.n198 CSoutput.n185 4.5005
R6190 CSoutput.n198 CSoutput.n192 4.5005
R6191 CSoutput.n241 CSoutput.n198 4.5005
R6192 CSoutput.n222 CSoutput.n188 4.5005
R6193 CSoutput.n222 CSoutput.n190 4.5005
R6194 CSoutput.n222 CSoutput.n187 4.5005
R6195 CSoutput.n222 CSoutput.n191 4.5005
R6196 CSoutput.n222 CSoutput.n186 4.5005
R6197 CSoutput.n222 CSoutput.t200 4.5005
R6198 CSoutput.n222 CSoutput.n185 4.5005
R6199 CSoutput.n222 CSoutput.n192 4.5005
R6200 CSoutput.n241 CSoutput.n222 4.5005
R6201 CSoutput.n188 CSoutput.n183 4.5005
R6202 CSoutput.n190 CSoutput.n183 4.5005
R6203 CSoutput.n187 CSoutput.n183 4.5005
R6204 CSoutput.n191 CSoutput.n183 4.5005
R6205 CSoutput.n186 CSoutput.n183 4.5005
R6206 CSoutput.t200 CSoutput.n183 4.5005
R6207 CSoutput.n185 CSoutput.n183 4.5005
R6208 CSoutput.n192 CSoutput.n183 4.5005
R6209 CSoutput.n244 CSoutput.n188 4.5005
R6210 CSoutput.n244 CSoutput.n190 4.5005
R6211 CSoutput.n244 CSoutput.n187 4.5005
R6212 CSoutput.n244 CSoutput.n191 4.5005
R6213 CSoutput.n244 CSoutput.n186 4.5005
R6214 CSoutput.n244 CSoutput.t200 4.5005
R6215 CSoutput.n244 CSoutput.n185 4.5005
R6216 CSoutput.n244 CSoutput.n192 4.5005
R6217 CSoutput.n242 CSoutput.n188 4.5005
R6218 CSoutput.n242 CSoutput.n190 4.5005
R6219 CSoutput.n242 CSoutput.n187 4.5005
R6220 CSoutput.n242 CSoutput.n191 4.5005
R6221 CSoutput.n242 CSoutput.n186 4.5005
R6222 CSoutput.n242 CSoutput.t200 4.5005
R6223 CSoutput.n242 CSoutput.n185 4.5005
R6224 CSoutput.n242 CSoutput.n192 4.5005
R6225 CSoutput.n242 CSoutput.n241 4.5005
R6226 CSoutput.n224 CSoutput.n188 4.5005
R6227 CSoutput.n224 CSoutput.n190 4.5005
R6228 CSoutput.n224 CSoutput.n187 4.5005
R6229 CSoutput.n224 CSoutput.n191 4.5005
R6230 CSoutput.n224 CSoutput.n186 4.5005
R6231 CSoutput.n224 CSoutput.t200 4.5005
R6232 CSoutput.n224 CSoutput.n185 4.5005
R6233 CSoutput.n224 CSoutput.n192 4.5005
R6234 CSoutput.n241 CSoutput.n224 4.5005
R6235 CSoutput.n196 CSoutput.n188 4.5005
R6236 CSoutput.n196 CSoutput.n190 4.5005
R6237 CSoutput.n196 CSoutput.n187 4.5005
R6238 CSoutput.n196 CSoutput.n191 4.5005
R6239 CSoutput.n196 CSoutput.n186 4.5005
R6240 CSoutput.n196 CSoutput.t200 4.5005
R6241 CSoutput.n196 CSoutput.n185 4.5005
R6242 CSoutput.n196 CSoutput.n192 4.5005
R6243 CSoutput.n241 CSoutput.n196 4.5005
R6244 CSoutput.n226 CSoutput.n188 4.5005
R6245 CSoutput.n226 CSoutput.n190 4.5005
R6246 CSoutput.n226 CSoutput.n187 4.5005
R6247 CSoutput.n226 CSoutput.n191 4.5005
R6248 CSoutput.n226 CSoutput.n186 4.5005
R6249 CSoutput.n226 CSoutput.t200 4.5005
R6250 CSoutput.n226 CSoutput.n185 4.5005
R6251 CSoutput.n226 CSoutput.n192 4.5005
R6252 CSoutput.n241 CSoutput.n226 4.5005
R6253 CSoutput.n195 CSoutput.n188 4.5005
R6254 CSoutput.n195 CSoutput.n190 4.5005
R6255 CSoutput.n195 CSoutput.n187 4.5005
R6256 CSoutput.n195 CSoutput.n191 4.5005
R6257 CSoutput.n195 CSoutput.n186 4.5005
R6258 CSoutput.n195 CSoutput.t200 4.5005
R6259 CSoutput.n195 CSoutput.n185 4.5005
R6260 CSoutput.n195 CSoutput.n192 4.5005
R6261 CSoutput.n241 CSoutput.n195 4.5005
R6262 CSoutput.n240 CSoutput.n188 4.5005
R6263 CSoutput.n240 CSoutput.n190 4.5005
R6264 CSoutput.n240 CSoutput.n187 4.5005
R6265 CSoutput.n240 CSoutput.n191 4.5005
R6266 CSoutput.n240 CSoutput.n186 4.5005
R6267 CSoutput.n240 CSoutput.t200 4.5005
R6268 CSoutput.n240 CSoutput.n185 4.5005
R6269 CSoutput.n240 CSoutput.n192 4.5005
R6270 CSoutput.n241 CSoutput.n240 4.5005
R6271 CSoutput.n239 CSoutput.n124 4.5005
R6272 CSoutput.n140 CSoutput.n124 4.5005
R6273 CSoutput.n135 CSoutput.n119 4.5005
R6274 CSoutput.n135 CSoutput.n121 4.5005
R6275 CSoutput.n135 CSoutput.n118 4.5005
R6276 CSoutput.n135 CSoutput.n122 4.5005
R6277 CSoutput.n135 CSoutput.n117 4.5005
R6278 CSoutput.n135 CSoutput.t201 4.5005
R6279 CSoutput.n135 CSoutput.n116 4.5005
R6280 CSoutput.n135 CSoutput.n123 4.5005
R6281 CSoutput.n135 CSoutput.n124 4.5005
R6282 CSoutput.n133 CSoutput.n119 4.5005
R6283 CSoutput.n133 CSoutput.n121 4.5005
R6284 CSoutput.n133 CSoutput.n118 4.5005
R6285 CSoutput.n133 CSoutput.n122 4.5005
R6286 CSoutput.n133 CSoutput.n117 4.5005
R6287 CSoutput.n133 CSoutput.t201 4.5005
R6288 CSoutput.n133 CSoutput.n116 4.5005
R6289 CSoutput.n133 CSoutput.n123 4.5005
R6290 CSoutput.n133 CSoutput.n124 4.5005
R6291 CSoutput.n132 CSoutput.n119 4.5005
R6292 CSoutput.n132 CSoutput.n121 4.5005
R6293 CSoutput.n132 CSoutput.n118 4.5005
R6294 CSoutput.n132 CSoutput.n122 4.5005
R6295 CSoutput.n132 CSoutput.n117 4.5005
R6296 CSoutput.n132 CSoutput.t201 4.5005
R6297 CSoutput.n132 CSoutput.n116 4.5005
R6298 CSoutput.n132 CSoutput.n123 4.5005
R6299 CSoutput.n132 CSoutput.n124 4.5005
R6300 CSoutput.n261 CSoutput.n119 4.5005
R6301 CSoutput.n261 CSoutput.n121 4.5005
R6302 CSoutput.n261 CSoutput.n118 4.5005
R6303 CSoutput.n261 CSoutput.n122 4.5005
R6304 CSoutput.n261 CSoutput.n117 4.5005
R6305 CSoutput.n261 CSoutput.t201 4.5005
R6306 CSoutput.n261 CSoutput.n116 4.5005
R6307 CSoutput.n261 CSoutput.n123 4.5005
R6308 CSoutput.n261 CSoutput.n124 4.5005
R6309 CSoutput.n259 CSoutput.n119 4.5005
R6310 CSoutput.n259 CSoutput.n121 4.5005
R6311 CSoutput.n259 CSoutput.n118 4.5005
R6312 CSoutput.n259 CSoutput.n122 4.5005
R6313 CSoutput.n259 CSoutput.n117 4.5005
R6314 CSoutput.n259 CSoutput.t201 4.5005
R6315 CSoutput.n259 CSoutput.n116 4.5005
R6316 CSoutput.n259 CSoutput.n123 4.5005
R6317 CSoutput.n257 CSoutput.n119 4.5005
R6318 CSoutput.n257 CSoutput.n121 4.5005
R6319 CSoutput.n257 CSoutput.n118 4.5005
R6320 CSoutput.n257 CSoutput.n122 4.5005
R6321 CSoutput.n257 CSoutput.n117 4.5005
R6322 CSoutput.n257 CSoutput.t201 4.5005
R6323 CSoutput.n257 CSoutput.n116 4.5005
R6324 CSoutput.n257 CSoutput.n123 4.5005
R6325 CSoutput.n143 CSoutput.n119 4.5005
R6326 CSoutput.n143 CSoutput.n121 4.5005
R6327 CSoutput.n143 CSoutput.n118 4.5005
R6328 CSoutput.n143 CSoutput.n122 4.5005
R6329 CSoutput.n143 CSoutput.n117 4.5005
R6330 CSoutput.n143 CSoutput.t201 4.5005
R6331 CSoutput.n143 CSoutput.n116 4.5005
R6332 CSoutput.n143 CSoutput.n123 4.5005
R6333 CSoutput.n143 CSoutput.n124 4.5005
R6334 CSoutput.n142 CSoutput.n119 4.5005
R6335 CSoutput.n142 CSoutput.n121 4.5005
R6336 CSoutput.n142 CSoutput.n118 4.5005
R6337 CSoutput.n142 CSoutput.n122 4.5005
R6338 CSoutput.n142 CSoutput.n117 4.5005
R6339 CSoutput.n142 CSoutput.t201 4.5005
R6340 CSoutput.n142 CSoutput.n116 4.5005
R6341 CSoutput.n142 CSoutput.n123 4.5005
R6342 CSoutput.n142 CSoutput.n124 4.5005
R6343 CSoutput.n146 CSoutput.n119 4.5005
R6344 CSoutput.n146 CSoutput.n121 4.5005
R6345 CSoutput.n146 CSoutput.n118 4.5005
R6346 CSoutput.n146 CSoutput.n122 4.5005
R6347 CSoutput.n146 CSoutput.n117 4.5005
R6348 CSoutput.n146 CSoutput.t201 4.5005
R6349 CSoutput.n146 CSoutput.n116 4.5005
R6350 CSoutput.n146 CSoutput.n123 4.5005
R6351 CSoutput.n146 CSoutput.n124 4.5005
R6352 CSoutput.n145 CSoutput.n119 4.5005
R6353 CSoutput.n145 CSoutput.n121 4.5005
R6354 CSoutput.n145 CSoutput.n118 4.5005
R6355 CSoutput.n145 CSoutput.n122 4.5005
R6356 CSoutput.n145 CSoutput.n117 4.5005
R6357 CSoutput.n145 CSoutput.t201 4.5005
R6358 CSoutput.n145 CSoutput.n116 4.5005
R6359 CSoutput.n145 CSoutput.n123 4.5005
R6360 CSoutput.n145 CSoutput.n124 4.5005
R6361 CSoutput.n128 CSoutput.n119 4.5005
R6362 CSoutput.n128 CSoutput.n121 4.5005
R6363 CSoutput.n128 CSoutput.n118 4.5005
R6364 CSoutput.n128 CSoutput.n122 4.5005
R6365 CSoutput.n128 CSoutput.n117 4.5005
R6366 CSoutput.n128 CSoutput.t201 4.5005
R6367 CSoutput.n128 CSoutput.n116 4.5005
R6368 CSoutput.n128 CSoutput.n123 4.5005
R6369 CSoutput.n128 CSoutput.n124 4.5005
R6370 CSoutput.n264 CSoutput.n119 4.5005
R6371 CSoutput.n264 CSoutput.n121 4.5005
R6372 CSoutput.n264 CSoutput.n118 4.5005
R6373 CSoutput.n264 CSoutput.n122 4.5005
R6374 CSoutput.n264 CSoutput.n117 4.5005
R6375 CSoutput.n264 CSoutput.t201 4.5005
R6376 CSoutput.n264 CSoutput.n116 4.5005
R6377 CSoutput.n264 CSoutput.n123 4.5005
R6378 CSoutput.n264 CSoutput.n124 4.5005
R6379 CSoutput.n299 CSoutput.n287 4.10845
R6380 CSoutput.n113 CSoutput.n101 4.10845
R6381 CSoutput.n297 CSoutput.t122 4.06363
R6382 CSoutput.n297 CSoutput.t123 4.06363
R6383 CSoutput.n295 CSoutput.t128 4.06363
R6384 CSoutput.n295 CSoutput.t167 4.06363
R6385 CSoutput.n293 CSoutput.t108 4.06363
R6386 CSoutput.n293 CSoutput.t126 4.06363
R6387 CSoutput.n291 CSoutput.t136 4.06363
R6388 CSoutput.n291 CSoutput.t151 4.06363
R6389 CSoutput.n289 CSoutput.t156 4.06363
R6390 CSoutput.n289 CSoutput.t110 4.06363
R6391 CSoutput.n288 CSoutput.t137 4.06363
R6392 CSoutput.n288 CSoutput.t138 4.06363
R6393 CSoutput.n285 CSoutput.t115 4.06363
R6394 CSoutput.n285 CSoutput.t116 4.06363
R6395 CSoutput.n283 CSoutput.t118 4.06363
R6396 CSoutput.n283 CSoutput.t160 4.06363
R6397 CSoutput.n281 CSoutput.t98 4.06363
R6398 CSoutput.n281 CSoutput.t117 4.06363
R6399 CSoutput.n279 CSoutput.t129 4.06363
R6400 CSoutput.n279 CSoutput.t143 4.06363
R6401 CSoutput.n277 CSoutput.t144 4.06363
R6402 CSoutput.n277 CSoutput.t102 4.06363
R6403 CSoutput.n276 CSoutput.t132 4.06363
R6404 CSoutput.n276 CSoutput.t133 4.06363
R6405 CSoutput.n274 CSoutput.t119 4.06363
R6406 CSoutput.n274 CSoutput.t106 4.06363
R6407 CSoutput.n272 CSoutput.t149 4.06363
R6408 CSoutput.n272 CSoutput.t103 4.06363
R6409 CSoutput.n270 CSoutput.t124 4.06363
R6410 CSoutput.n270 CSoutput.t165 4.06363
R6411 CSoutput.n268 CSoutput.t112 4.06363
R6412 CSoutput.n268 CSoutput.t153 4.06363
R6413 CSoutput.n266 CSoutput.t130 4.06363
R6414 CSoutput.n266 CSoutput.t168 4.06363
R6415 CSoutput.n265 CSoutput.t99 4.06363
R6416 CSoutput.n265 CSoutput.t158 4.06363
R6417 CSoutput.n102 CSoutput.t164 4.06363
R6418 CSoutput.n102 CSoutput.t163 4.06363
R6419 CSoutput.n103 CSoutput.t150 4.06363
R6420 CSoutput.n103 CSoutput.t111 4.06363
R6421 CSoutput.n105 CSoutput.t109 4.06363
R6422 CSoutput.n105 CSoutput.t161 4.06363
R6423 CSoutput.n107 CSoutput.t148 4.06363
R6424 CSoutput.n107 CSoutput.t134 4.06363
R6425 CSoutput.n109 CSoutput.t121 4.06363
R6426 CSoutput.n109 CSoutput.t169 4.06363
R6427 CSoutput.n111 CSoutput.t146 4.06363
R6428 CSoutput.n111 CSoutput.t145 4.06363
R6429 CSoutput.n90 CSoutput.t157 4.06363
R6430 CSoutput.n90 CSoutput.t155 4.06363
R6431 CSoutput.n91 CSoutput.t142 4.06363
R6432 CSoutput.n91 CSoutput.t105 4.06363
R6433 CSoutput.n93 CSoutput.t101 4.06363
R6434 CSoutput.n93 CSoutput.t152 4.06363
R6435 CSoutput.n95 CSoutput.t141 4.06363
R6436 CSoutput.n95 CSoutput.t127 4.06363
R6437 CSoutput.n97 CSoutput.t114 4.06363
R6438 CSoutput.n97 CSoutput.t162 4.06363
R6439 CSoutput.n99 CSoutput.t140 4.06363
R6440 CSoutput.n99 CSoutput.t139 4.06363
R6441 CSoutput.n79 CSoutput.t159 4.06363
R6442 CSoutput.n79 CSoutput.t100 4.06363
R6443 CSoutput.n80 CSoutput.t147 4.06363
R6444 CSoutput.n80 CSoutput.t131 4.06363
R6445 CSoutput.n82 CSoutput.t154 4.06363
R6446 CSoutput.n82 CSoutput.t113 4.06363
R6447 CSoutput.n84 CSoutput.t166 4.06363
R6448 CSoutput.n84 CSoutput.t125 4.06363
R6449 CSoutput.n86 CSoutput.t104 4.06363
R6450 CSoutput.n86 CSoutput.t135 4.06363
R6451 CSoutput.n88 CSoutput.t107 4.06363
R6452 CSoutput.n88 CSoutput.t120 4.06363
R6453 CSoutput.n44 CSoutput.n43 3.79402
R6454 CSoutput.n49 CSoutput.n48 3.79402
R6455 CSoutput.n359 CSoutput.n339 3.72967
R6456 CSoutput.n419 CSoutput.n399 3.72967
R6457 CSoutput.n420 CSoutput.n360 3.71319
R6458 CSoutput.n421 CSoutput.n420 3.57343
R6459 CSoutput.n357 CSoutput.t9 2.82907
R6460 CSoutput.n357 CSoutput.t52 2.82907
R6461 CSoutput.n355 CSoutput.t191 2.82907
R6462 CSoutput.n355 CSoutput.t7 2.82907
R6463 CSoutput.n353 CSoutput.t55 2.82907
R6464 CSoutput.n353 CSoutput.t97 2.82907
R6465 CSoutput.n351 CSoutput.t33 2.82907
R6466 CSoutput.n351 CSoutput.t187 2.82907
R6467 CSoutput.n349 CSoutput.t61 2.82907
R6468 CSoutput.n349 CSoutput.t69 2.82907
R6469 CSoutput.n347 CSoutput.t96 2.82907
R6470 CSoutput.n347 CSoutput.t43 2.82907
R6471 CSoutput.n345 CSoutput.t81 2.82907
R6472 CSoutput.n345 CSoutput.t21 2.82907
R6473 CSoutput.n343 CSoutput.t1 2.82907
R6474 CSoutput.n343 CSoutput.t95 2.82907
R6475 CSoutput.n341 CSoutput.t22 2.82907
R6476 CSoutput.n341 CSoutput.t25 2.82907
R6477 CSoutput.n340 CSoutput.t171 2.82907
R6478 CSoutput.n340 CSoutput.t44 2.82907
R6479 CSoutput.n337 CSoutput.t56 2.82907
R6480 CSoutput.n337 CSoutput.t30 2.82907
R6481 CSoutput.n335 CSoutput.t73 2.82907
R6482 CSoutput.n335 CSoutput.t182 2.82907
R6483 CSoutput.n333 CSoutput.t35 2.82907
R6484 CSoutput.n333 CSoutput.t64 2.82907
R6485 CSoutput.n331 CSoutput.t189 2.82907
R6486 CSoutput.n331 CSoutput.t190 2.82907
R6487 CSoutput.n329 CSoutput.t90 2.82907
R6488 CSoutput.n329 CSoutput.t84 2.82907
R6489 CSoutput.n327 CSoutput.t71 2.82907
R6490 CSoutput.n327 CSoutput.t20 2.82907
R6491 CSoutput.n325 CSoutput.t38 2.82907
R6492 CSoutput.n325 CSoutput.t15 2.82907
R6493 CSoutput.n323 CSoutput.t184 2.82907
R6494 CSoutput.n323 CSoutput.t59 2.82907
R6495 CSoutput.n321 CSoutput.t0 2.82907
R6496 CSoutput.n321 CSoutput.t170 2.82907
R6497 CSoutput.n320 CSoutput.t50 2.82907
R6498 CSoutput.n320 CSoutput.t36 2.82907
R6499 CSoutput.n318 CSoutput.t66 2.82907
R6500 CSoutput.n318 CSoutput.t85 2.82907
R6501 CSoutput.n316 CSoutput.t45 2.82907
R6502 CSoutput.n316 CSoutput.t82 2.82907
R6503 CSoutput.n314 CSoutput.t176 2.82907
R6504 CSoutput.n314 CSoutput.t87 2.82907
R6505 CSoutput.n312 CSoutput.t19 2.82907
R6506 CSoutput.n312 CSoutput.t58 2.82907
R6507 CSoutput.n310 CSoutput.t65 2.82907
R6508 CSoutput.n310 CSoutput.t181 2.82907
R6509 CSoutput.n308 CSoutput.t41 2.82907
R6510 CSoutput.n308 CSoutput.t51 2.82907
R6511 CSoutput.n306 CSoutput.t86 2.82907
R6512 CSoutput.n306 CSoutput.t92 2.82907
R6513 CSoutput.n304 CSoutput.t74 2.82907
R6514 CSoutput.n304 CSoutput.t31 2.82907
R6515 CSoutput.n302 CSoutput.t93 2.82907
R6516 CSoutput.n302 CSoutput.t186 2.82907
R6517 CSoutput.n301 CSoutput.t46 2.82907
R6518 CSoutput.n301 CSoutput.t88 2.82907
R6519 CSoutput.n400 CSoutput.t29 2.82907
R6520 CSoutput.n400 CSoutput.t177 2.82907
R6521 CSoutput.n401 CSoutput.t11 2.82907
R6522 CSoutput.n401 CSoutput.t79 2.82907
R6523 CSoutput.n403 CSoutput.t78 2.82907
R6524 CSoutput.n403 CSoutput.t37 2.82907
R6525 CSoutput.n405 CSoutput.t180 2.82907
R6526 CSoutput.n405 CSoutput.t5 2.82907
R6527 CSoutput.n407 CSoutput.t17 2.82907
R6528 CSoutput.n407 CSoutput.t14 2.82907
R6529 CSoutput.n409 CSoutput.t53 2.82907
R6530 CSoutput.n409 CSoutput.t54 2.82907
R6531 CSoutput.n411 CSoutput.t172 2.82907
R6532 CSoutput.n411 CSoutput.t94 2.82907
R6533 CSoutput.n413 CSoutput.t13 2.82907
R6534 CSoutput.n413 CSoutput.t2 2.82907
R6535 CSoutput.n415 CSoutput.t75 2.82907
R6536 CSoutput.n415 CSoutput.t3 2.82907
R6537 CSoutput.n417 CSoutput.t185 2.82907
R6538 CSoutput.n417 CSoutput.t42 2.82907
R6539 CSoutput.n380 CSoutput.t179 2.82907
R6540 CSoutput.n380 CSoutput.t10 2.82907
R6541 CSoutput.n381 CSoutput.t48 2.82907
R6542 CSoutput.n381 CSoutput.t80 2.82907
R6543 CSoutput.n383 CSoutput.t8 2.82907
R6544 CSoutput.n383 CSoutput.t32 2.82907
R6545 CSoutput.n385 CSoutput.t39 2.82907
R6546 CSoutput.n385 CSoutput.t6 2.82907
R6547 CSoutput.n387 CSoutput.t63 2.82907
R6548 CSoutput.n387 CSoutput.t16 2.82907
R6549 CSoutput.n389 CSoutput.t175 2.82907
R6550 CSoutput.n389 CSoutput.t24 2.82907
R6551 CSoutput.n391 CSoutput.t76 2.82907
R6552 CSoutput.n391 CSoutput.t47 2.82907
R6553 CSoutput.n393 CSoutput.t18 2.82907
R6554 CSoutput.n393 CSoutput.t28 2.82907
R6555 CSoutput.n395 CSoutput.t173 2.82907
R6556 CSoutput.n395 CSoutput.t178 2.82907
R6557 CSoutput.n397 CSoutput.t77 2.82907
R6558 CSoutput.n397 CSoutput.t12 2.82907
R6559 CSoutput.n361 CSoutput.t4 2.82907
R6560 CSoutput.n361 CSoutput.t68 2.82907
R6561 CSoutput.n362 CSoutput.t34 2.82907
R6562 CSoutput.n362 CSoutput.t91 2.82907
R6563 CSoutput.n364 CSoutput.t27 2.82907
R6564 CSoutput.n364 CSoutput.t49 2.82907
R6565 CSoutput.n366 CSoutput.t83 2.82907
R6566 CSoutput.n366 CSoutput.t89 2.82907
R6567 CSoutput.n368 CSoutput.t23 2.82907
R6568 CSoutput.n368 CSoutput.t188 2.82907
R6569 CSoutput.n370 CSoutput.t174 2.82907
R6570 CSoutput.n370 CSoutput.t183 2.82907
R6571 CSoutput.n372 CSoutput.t62 2.82907
R6572 CSoutput.n372 CSoutput.t60 2.82907
R6573 CSoutput.n374 CSoutput.t40 2.82907
R6574 CSoutput.n374 CSoutput.t26 2.82907
R6575 CSoutput.n376 CSoutput.t72 2.82907
R6576 CSoutput.n376 CSoutput.t70 2.82907
R6577 CSoutput.n378 CSoutput.t57 2.82907
R6578 CSoutput.n378 CSoutput.t67 2.82907
R6579 CSoutput.n75 CSoutput.n1 2.45513
R6580 CSoutput.n205 CSoutput.n203 2.251
R6581 CSoutput.n205 CSoutput.n202 2.251
R6582 CSoutput.n205 CSoutput.n201 2.251
R6583 CSoutput.n205 CSoutput.n200 2.251
R6584 CSoutput.n174 CSoutput.n173 2.251
R6585 CSoutput.n174 CSoutput.n172 2.251
R6586 CSoutput.n174 CSoutput.n171 2.251
R6587 CSoutput.n174 CSoutput.n170 2.251
R6588 CSoutput.n247 CSoutput.n246 2.251
R6589 CSoutput.n212 CSoutput.n210 2.251
R6590 CSoutput.n212 CSoutput.n209 2.251
R6591 CSoutput.n212 CSoutput.n208 2.251
R6592 CSoutput.n230 CSoutput.n212 2.251
R6593 CSoutput.n218 CSoutput.n217 2.251
R6594 CSoutput.n218 CSoutput.n216 2.251
R6595 CSoutput.n218 CSoutput.n215 2.251
R6596 CSoutput.n218 CSoutput.n214 2.251
R6597 CSoutput.n244 CSoutput.n184 2.251
R6598 CSoutput.n239 CSoutput.n237 2.251
R6599 CSoutput.n239 CSoutput.n236 2.251
R6600 CSoutput.n239 CSoutput.n235 2.251
R6601 CSoutput.n239 CSoutput.n234 2.251
R6602 CSoutput.n140 CSoutput.n139 2.251
R6603 CSoutput.n140 CSoutput.n138 2.251
R6604 CSoutput.n140 CSoutput.n137 2.251
R6605 CSoutput.n140 CSoutput.n136 2.251
R6606 CSoutput.n257 CSoutput.n256 2.251
R6607 CSoutput.n174 CSoutput.n154 2.2505
R6608 CSoutput.n169 CSoutput.n154 2.2505
R6609 CSoutput.n167 CSoutput.n154 2.2505
R6610 CSoutput.n166 CSoutput.n154 2.2505
R6611 CSoutput.n251 CSoutput.n154 2.2505
R6612 CSoutput.n249 CSoutput.n154 2.2505
R6613 CSoutput.n247 CSoutput.n154 2.2505
R6614 CSoutput.n177 CSoutput.n154 2.2505
R6615 CSoutput.n176 CSoutput.n154 2.2505
R6616 CSoutput.n180 CSoutput.n154 2.2505
R6617 CSoutput.n179 CSoutput.n154 2.2505
R6618 CSoutput.n162 CSoutput.n154 2.2505
R6619 CSoutput.n254 CSoutput.n154 2.2505
R6620 CSoutput.n254 CSoutput.n253 2.2505
R6621 CSoutput.n218 CSoutput.n189 2.2505
R6622 CSoutput.n199 CSoutput.n189 2.2505
R6623 CSoutput.n220 CSoutput.n189 2.2505
R6624 CSoutput.n198 CSoutput.n189 2.2505
R6625 CSoutput.n222 CSoutput.n189 2.2505
R6626 CSoutput.n189 CSoutput.n183 2.2505
R6627 CSoutput.n244 CSoutput.n189 2.2505
R6628 CSoutput.n242 CSoutput.n189 2.2505
R6629 CSoutput.n224 CSoutput.n189 2.2505
R6630 CSoutput.n196 CSoutput.n189 2.2505
R6631 CSoutput.n226 CSoutput.n189 2.2505
R6632 CSoutput.n195 CSoutput.n189 2.2505
R6633 CSoutput.n240 CSoutput.n189 2.2505
R6634 CSoutput.n240 CSoutput.n193 2.2505
R6635 CSoutput.n140 CSoutput.n120 2.2505
R6636 CSoutput.n135 CSoutput.n120 2.2505
R6637 CSoutput.n133 CSoutput.n120 2.2505
R6638 CSoutput.n132 CSoutput.n120 2.2505
R6639 CSoutput.n261 CSoutput.n120 2.2505
R6640 CSoutput.n259 CSoutput.n120 2.2505
R6641 CSoutput.n257 CSoutput.n120 2.2505
R6642 CSoutput.n143 CSoutput.n120 2.2505
R6643 CSoutput.n142 CSoutput.n120 2.2505
R6644 CSoutput.n146 CSoutput.n120 2.2505
R6645 CSoutput.n145 CSoutput.n120 2.2505
R6646 CSoutput.n128 CSoutput.n120 2.2505
R6647 CSoutput.n264 CSoutput.n120 2.2505
R6648 CSoutput.n264 CSoutput.n263 2.2505
R6649 CSoutput.n182 CSoutput.n175 2.25024
R6650 CSoutput.n182 CSoutput.n168 2.25024
R6651 CSoutput.n250 CSoutput.n182 2.25024
R6652 CSoutput.n182 CSoutput.n178 2.25024
R6653 CSoutput.n182 CSoutput.n181 2.25024
R6654 CSoutput.n182 CSoutput.n149 2.25024
R6655 CSoutput.n232 CSoutput.n229 2.25024
R6656 CSoutput.n232 CSoutput.n228 2.25024
R6657 CSoutput.n232 CSoutput.n227 2.25024
R6658 CSoutput.n232 CSoutput.n194 2.25024
R6659 CSoutput.n232 CSoutput.n231 2.25024
R6660 CSoutput.n233 CSoutput.n232 2.25024
R6661 CSoutput.n148 CSoutput.n141 2.25024
R6662 CSoutput.n148 CSoutput.n134 2.25024
R6663 CSoutput.n260 CSoutput.n148 2.25024
R6664 CSoutput.n148 CSoutput.n144 2.25024
R6665 CSoutput.n148 CSoutput.n147 2.25024
R6666 CSoutput.n148 CSoutput.n115 2.25024
R6667 CSoutput.n300 CSoutput.n114 2.15937
R6668 CSoutput.n249 CSoutput.n159 1.50111
R6669 CSoutput.n197 CSoutput.n183 1.50111
R6670 CSoutput.n259 CSoutput.n125 1.50111
R6671 CSoutput.n205 CSoutput.n204 1.501
R6672 CSoutput.n212 CSoutput.n211 1.501
R6673 CSoutput.n239 CSoutput.n238 1.501
R6674 CSoutput.n253 CSoutput.n164 1.12536
R6675 CSoutput.n253 CSoutput.n165 1.12536
R6676 CSoutput.n253 CSoutput.n252 1.12536
R6677 CSoutput.n213 CSoutput.n193 1.12536
R6678 CSoutput.n219 CSoutput.n193 1.12536
R6679 CSoutput.n221 CSoutput.n193 1.12536
R6680 CSoutput.n263 CSoutput.n130 1.12536
R6681 CSoutput.n263 CSoutput.n131 1.12536
R6682 CSoutput.n263 CSoutput.n262 1.12536
R6683 CSoutput.n253 CSoutput.n160 1.12536
R6684 CSoutput.n253 CSoutput.n161 1.12536
R6685 CSoutput.n253 CSoutput.n163 1.12536
R6686 CSoutput.n243 CSoutput.n193 1.12536
R6687 CSoutput.n223 CSoutput.n193 1.12536
R6688 CSoutput.n225 CSoutput.n193 1.12536
R6689 CSoutput.n263 CSoutput.n126 1.12536
R6690 CSoutput.n263 CSoutput.n127 1.12536
R6691 CSoutput.n263 CSoutput.n129 1.12536
R6692 CSoutput.n31 CSoutput.n30 0.669944
R6693 CSoutput.n62 CSoutput.n61 0.669944
R6694 CSoutput.n344 CSoutput.n342 0.573776
R6695 CSoutput.n346 CSoutput.n344 0.573776
R6696 CSoutput.n348 CSoutput.n346 0.573776
R6697 CSoutput.n350 CSoutput.n348 0.573776
R6698 CSoutput.n352 CSoutput.n350 0.573776
R6699 CSoutput.n354 CSoutput.n352 0.573776
R6700 CSoutput.n356 CSoutput.n354 0.573776
R6701 CSoutput.n358 CSoutput.n356 0.573776
R6702 CSoutput.n324 CSoutput.n322 0.573776
R6703 CSoutput.n326 CSoutput.n324 0.573776
R6704 CSoutput.n328 CSoutput.n326 0.573776
R6705 CSoutput.n330 CSoutput.n328 0.573776
R6706 CSoutput.n332 CSoutput.n330 0.573776
R6707 CSoutput.n334 CSoutput.n332 0.573776
R6708 CSoutput.n336 CSoutput.n334 0.573776
R6709 CSoutput.n338 CSoutput.n336 0.573776
R6710 CSoutput.n305 CSoutput.n303 0.573776
R6711 CSoutput.n307 CSoutput.n305 0.573776
R6712 CSoutput.n309 CSoutput.n307 0.573776
R6713 CSoutput.n311 CSoutput.n309 0.573776
R6714 CSoutput.n313 CSoutput.n311 0.573776
R6715 CSoutput.n315 CSoutput.n313 0.573776
R6716 CSoutput.n317 CSoutput.n315 0.573776
R6717 CSoutput.n319 CSoutput.n317 0.573776
R6718 CSoutput.n418 CSoutput.n416 0.573776
R6719 CSoutput.n416 CSoutput.n414 0.573776
R6720 CSoutput.n414 CSoutput.n412 0.573776
R6721 CSoutput.n412 CSoutput.n410 0.573776
R6722 CSoutput.n410 CSoutput.n408 0.573776
R6723 CSoutput.n408 CSoutput.n406 0.573776
R6724 CSoutput.n406 CSoutput.n404 0.573776
R6725 CSoutput.n404 CSoutput.n402 0.573776
R6726 CSoutput.n398 CSoutput.n396 0.573776
R6727 CSoutput.n396 CSoutput.n394 0.573776
R6728 CSoutput.n394 CSoutput.n392 0.573776
R6729 CSoutput.n392 CSoutput.n390 0.573776
R6730 CSoutput.n390 CSoutput.n388 0.573776
R6731 CSoutput.n388 CSoutput.n386 0.573776
R6732 CSoutput.n386 CSoutput.n384 0.573776
R6733 CSoutput.n384 CSoutput.n382 0.573776
R6734 CSoutput.n379 CSoutput.n377 0.573776
R6735 CSoutput.n377 CSoutput.n375 0.573776
R6736 CSoutput.n375 CSoutput.n373 0.573776
R6737 CSoutput.n373 CSoutput.n371 0.573776
R6738 CSoutput.n371 CSoutput.n369 0.573776
R6739 CSoutput.n369 CSoutput.n367 0.573776
R6740 CSoutput.n367 CSoutput.n365 0.573776
R6741 CSoutput.n365 CSoutput.n363 0.573776
R6742 CSoutput.n421 CSoutput.n264 0.53442
R6743 CSoutput.n292 CSoutput.n290 0.358259
R6744 CSoutput.n294 CSoutput.n292 0.358259
R6745 CSoutput.n296 CSoutput.n294 0.358259
R6746 CSoutput.n298 CSoutput.n296 0.358259
R6747 CSoutput.n280 CSoutput.n278 0.358259
R6748 CSoutput.n282 CSoutput.n280 0.358259
R6749 CSoutput.n284 CSoutput.n282 0.358259
R6750 CSoutput.n286 CSoutput.n284 0.358259
R6751 CSoutput.n269 CSoutput.n267 0.358259
R6752 CSoutput.n271 CSoutput.n269 0.358259
R6753 CSoutput.n273 CSoutput.n271 0.358259
R6754 CSoutput.n275 CSoutput.n273 0.358259
R6755 CSoutput.n112 CSoutput.n110 0.358259
R6756 CSoutput.n110 CSoutput.n108 0.358259
R6757 CSoutput.n108 CSoutput.n106 0.358259
R6758 CSoutput.n106 CSoutput.n104 0.358259
R6759 CSoutput.n100 CSoutput.n98 0.358259
R6760 CSoutput.n98 CSoutput.n96 0.358259
R6761 CSoutput.n96 CSoutput.n94 0.358259
R6762 CSoutput.n94 CSoutput.n92 0.358259
R6763 CSoutput.n89 CSoutput.n87 0.358259
R6764 CSoutput.n87 CSoutput.n85 0.358259
R6765 CSoutput.n85 CSoutput.n83 0.358259
R6766 CSoutput.n83 CSoutput.n81 0.358259
R6767 CSoutput.n21 CSoutput.n20 0.169105
R6768 CSoutput.n21 CSoutput.n16 0.169105
R6769 CSoutput.n26 CSoutput.n16 0.169105
R6770 CSoutput.n27 CSoutput.n26 0.169105
R6771 CSoutput.n27 CSoutput.n14 0.169105
R6772 CSoutput.n32 CSoutput.n14 0.169105
R6773 CSoutput.n33 CSoutput.n32 0.169105
R6774 CSoutput.n34 CSoutput.n33 0.169105
R6775 CSoutput.n34 CSoutput.n12 0.169105
R6776 CSoutput.n39 CSoutput.n12 0.169105
R6777 CSoutput.n40 CSoutput.n39 0.169105
R6778 CSoutput.n40 CSoutput.n10 0.169105
R6779 CSoutput.n45 CSoutput.n10 0.169105
R6780 CSoutput.n46 CSoutput.n45 0.169105
R6781 CSoutput.n47 CSoutput.n46 0.169105
R6782 CSoutput.n47 CSoutput.n8 0.169105
R6783 CSoutput.n52 CSoutput.n8 0.169105
R6784 CSoutput.n53 CSoutput.n52 0.169105
R6785 CSoutput.n53 CSoutput.n6 0.169105
R6786 CSoutput.n58 CSoutput.n6 0.169105
R6787 CSoutput.n59 CSoutput.n58 0.169105
R6788 CSoutput.n60 CSoutput.n59 0.169105
R6789 CSoutput.n60 CSoutput.n4 0.169105
R6790 CSoutput.n66 CSoutput.n4 0.169105
R6791 CSoutput.n67 CSoutput.n66 0.169105
R6792 CSoutput.n68 CSoutput.n67 0.169105
R6793 CSoutput.n68 CSoutput.n2 0.169105
R6794 CSoutput.n73 CSoutput.n2 0.169105
R6795 CSoutput.n74 CSoutput.n73 0.169105
R6796 CSoutput.n74 CSoutput.n0 0.169105
R6797 CSoutput.n78 CSoutput.n0 0.169105
R6798 CSoutput.n207 CSoutput.n206 0.0910737
R6799 CSoutput.n258 CSoutput.n255 0.0723685
R6800 CSoutput.n212 CSoutput.n207 0.0522944
R6801 CSoutput.n255 CSoutput.n254 0.0499135
R6802 CSoutput.n206 CSoutput.n205 0.0499135
R6803 CSoutput.n240 CSoutput.n239 0.0464294
R6804 CSoutput.n248 CSoutput.n245 0.0391444
R6805 CSoutput.n207 CSoutput.t210 0.023435
R6806 CSoutput.n255 CSoutput.t194 0.02262
R6807 CSoutput.n206 CSoutput.t206 0.02262
R6808 CSoutput CSoutput.n421 0.0052
R6809 CSoutput.n177 CSoutput.n160 0.00365111
R6810 CSoutput.n180 CSoutput.n161 0.00365111
R6811 CSoutput.n163 CSoutput.n162 0.00365111
R6812 CSoutput.n205 CSoutput.n164 0.00365111
R6813 CSoutput.n169 CSoutput.n165 0.00365111
R6814 CSoutput.n252 CSoutput.n166 0.00365111
R6815 CSoutput.n243 CSoutput.n242 0.00365111
R6816 CSoutput.n223 CSoutput.n196 0.00365111
R6817 CSoutput.n225 CSoutput.n195 0.00365111
R6818 CSoutput.n213 CSoutput.n212 0.00365111
R6819 CSoutput.n219 CSoutput.n199 0.00365111
R6820 CSoutput.n221 CSoutput.n198 0.00365111
R6821 CSoutput.n143 CSoutput.n126 0.00365111
R6822 CSoutput.n146 CSoutput.n127 0.00365111
R6823 CSoutput.n129 CSoutput.n128 0.00365111
R6824 CSoutput.n239 CSoutput.n130 0.00365111
R6825 CSoutput.n135 CSoutput.n131 0.00365111
R6826 CSoutput.n262 CSoutput.n132 0.00365111
R6827 CSoutput.n174 CSoutput.n164 0.00340054
R6828 CSoutput.n167 CSoutput.n165 0.00340054
R6829 CSoutput.n252 CSoutput.n251 0.00340054
R6830 CSoutput.n247 CSoutput.n160 0.00340054
R6831 CSoutput.n176 CSoutput.n161 0.00340054
R6832 CSoutput.n179 CSoutput.n163 0.00340054
R6833 CSoutput.n218 CSoutput.n213 0.00340054
R6834 CSoutput.n220 CSoutput.n219 0.00340054
R6835 CSoutput.n222 CSoutput.n221 0.00340054
R6836 CSoutput.n244 CSoutput.n243 0.00340054
R6837 CSoutput.n224 CSoutput.n223 0.00340054
R6838 CSoutput.n226 CSoutput.n225 0.00340054
R6839 CSoutput.n140 CSoutput.n130 0.00340054
R6840 CSoutput.n133 CSoutput.n131 0.00340054
R6841 CSoutput.n262 CSoutput.n261 0.00340054
R6842 CSoutput.n257 CSoutput.n126 0.00340054
R6843 CSoutput.n142 CSoutput.n127 0.00340054
R6844 CSoutput.n145 CSoutput.n129 0.00340054
R6845 CSoutput.n175 CSoutput.n169 0.00252698
R6846 CSoutput.n168 CSoutput.n166 0.00252698
R6847 CSoutput.n250 CSoutput.n249 0.00252698
R6848 CSoutput.n178 CSoutput.n176 0.00252698
R6849 CSoutput.n181 CSoutput.n179 0.00252698
R6850 CSoutput.n254 CSoutput.n149 0.00252698
R6851 CSoutput.n175 CSoutput.n174 0.00252698
R6852 CSoutput.n168 CSoutput.n167 0.00252698
R6853 CSoutput.n251 CSoutput.n250 0.00252698
R6854 CSoutput.n178 CSoutput.n177 0.00252698
R6855 CSoutput.n181 CSoutput.n180 0.00252698
R6856 CSoutput.n162 CSoutput.n149 0.00252698
R6857 CSoutput.n229 CSoutput.n199 0.00252698
R6858 CSoutput.n228 CSoutput.n198 0.00252698
R6859 CSoutput.n227 CSoutput.n183 0.00252698
R6860 CSoutput.n224 CSoutput.n194 0.00252698
R6861 CSoutput.n231 CSoutput.n226 0.00252698
R6862 CSoutput.n240 CSoutput.n233 0.00252698
R6863 CSoutput.n229 CSoutput.n218 0.00252698
R6864 CSoutput.n228 CSoutput.n220 0.00252698
R6865 CSoutput.n227 CSoutput.n222 0.00252698
R6866 CSoutput.n242 CSoutput.n194 0.00252698
R6867 CSoutput.n231 CSoutput.n196 0.00252698
R6868 CSoutput.n233 CSoutput.n195 0.00252698
R6869 CSoutput.n141 CSoutput.n135 0.00252698
R6870 CSoutput.n134 CSoutput.n132 0.00252698
R6871 CSoutput.n260 CSoutput.n259 0.00252698
R6872 CSoutput.n144 CSoutput.n142 0.00252698
R6873 CSoutput.n147 CSoutput.n145 0.00252698
R6874 CSoutput.n264 CSoutput.n115 0.00252698
R6875 CSoutput.n141 CSoutput.n140 0.00252698
R6876 CSoutput.n134 CSoutput.n133 0.00252698
R6877 CSoutput.n261 CSoutput.n260 0.00252698
R6878 CSoutput.n144 CSoutput.n143 0.00252698
R6879 CSoutput.n147 CSoutput.n146 0.00252698
R6880 CSoutput.n128 CSoutput.n115 0.00252698
R6881 CSoutput.n249 CSoutput.n248 0.0020275
R6882 CSoutput.n248 CSoutput.n247 0.0020275
R6883 CSoutput.n245 CSoutput.n183 0.0020275
R6884 CSoutput.n245 CSoutput.n244 0.0020275
R6885 CSoutput.n259 CSoutput.n258 0.0020275
R6886 CSoutput.n258 CSoutput.n257 0.0020275
R6887 CSoutput.n159 CSoutput.n158 0.00166668
R6888 CSoutput.n241 CSoutput.n197 0.00166668
R6889 CSoutput.n125 CSoutput.n124 0.00166668
R6890 CSoutput.n263 CSoutput.n125 0.00133328
R6891 CSoutput.n197 CSoutput.n193 0.00133328
R6892 CSoutput.n253 CSoutput.n159 0.00133328
R6893 CSoutput.n256 CSoutput.n148 0.001
R6894 CSoutput.n234 CSoutput.n148 0.001
R6895 CSoutput.n136 CSoutput.n116 0.001
R6896 CSoutput.n235 CSoutput.n116 0.001
R6897 CSoutput.n137 CSoutput.n117 0.001
R6898 CSoutput.n236 CSoutput.n117 0.001
R6899 CSoutput.n138 CSoutput.n118 0.001
R6900 CSoutput.n237 CSoutput.n118 0.001
R6901 CSoutput.n139 CSoutput.n119 0.001
R6902 CSoutput.n238 CSoutput.n119 0.001
R6903 CSoutput.n232 CSoutput.n184 0.001
R6904 CSoutput.n232 CSoutput.n230 0.001
R6905 CSoutput.n214 CSoutput.n185 0.001
R6906 CSoutput.n208 CSoutput.n185 0.001
R6907 CSoutput.n215 CSoutput.n186 0.001
R6908 CSoutput.n209 CSoutput.n186 0.001
R6909 CSoutput.n216 CSoutput.n187 0.001
R6910 CSoutput.n210 CSoutput.n187 0.001
R6911 CSoutput.n217 CSoutput.n188 0.001
R6912 CSoutput.n211 CSoutput.n188 0.001
R6913 CSoutput.n246 CSoutput.n182 0.001
R6914 CSoutput.n200 CSoutput.n182 0.001
R6915 CSoutput.n170 CSoutput.n150 0.001
R6916 CSoutput.n201 CSoutput.n150 0.001
R6917 CSoutput.n171 CSoutput.n151 0.001
R6918 CSoutput.n202 CSoutput.n151 0.001
R6919 CSoutput.n172 CSoutput.n152 0.001
R6920 CSoutput.n203 CSoutput.n152 0.001
R6921 CSoutput.n173 CSoutput.n153 0.001
R6922 CSoutput.n204 CSoutput.n153 0.001
R6923 CSoutput.n204 CSoutput.n154 0.001
R6924 CSoutput.n203 CSoutput.n155 0.001
R6925 CSoutput.n202 CSoutput.n156 0.001
R6926 CSoutput.n201 CSoutput.t196 0.001
R6927 CSoutput.n200 CSoutput.n157 0.001
R6928 CSoutput.n173 CSoutput.n155 0.001
R6929 CSoutput.n172 CSoutput.n156 0.001
R6930 CSoutput.n171 CSoutput.t196 0.001
R6931 CSoutput.n170 CSoutput.n157 0.001
R6932 CSoutput.n246 CSoutput.n158 0.001
R6933 CSoutput.n211 CSoutput.n189 0.001
R6934 CSoutput.n210 CSoutput.n190 0.001
R6935 CSoutput.n209 CSoutput.n191 0.001
R6936 CSoutput.n208 CSoutput.t200 0.001
R6937 CSoutput.n230 CSoutput.n192 0.001
R6938 CSoutput.n217 CSoutput.n190 0.001
R6939 CSoutput.n216 CSoutput.n191 0.001
R6940 CSoutput.n215 CSoutput.t200 0.001
R6941 CSoutput.n214 CSoutput.n192 0.001
R6942 CSoutput.n241 CSoutput.n184 0.001
R6943 CSoutput.n238 CSoutput.n120 0.001
R6944 CSoutput.n237 CSoutput.n121 0.001
R6945 CSoutput.n236 CSoutput.n122 0.001
R6946 CSoutput.n235 CSoutput.t201 0.001
R6947 CSoutput.n234 CSoutput.n123 0.001
R6948 CSoutput.n139 CSoutput.n121 0.001
R6949 CSoutput.n138 CSoutput.n122 0.001
R6950 CSoutput.n137 CSoutput.t201 0.001
R6951 CSoutput.n136 CSoutput.n123 0.001
R6952 CSoutput.n256 CSoutput.n124 0.001
R6953 commonsourceibias.n397 commonsourceibias.t184 222.032
R6954 commonsourceibias.n281 commonsourceibias.t94 222.032
R6955 commonsourceibias.n44 commonsourceibias.t8 222.032
R6956 commonsourceibias.n166 commonsourceibias.t100 222.032
R6957 commonsourceibias.n875 commonsourceibias.t196 222.032
R6958 commonsourceibias.n759 commonsourceibias.t188 222.032
R6959 commonsourceibias.n529 commonsourceibias.t16 222.032
R6960 commonsourceibias.n645 commonsourceibias.t153 222.032
R6961 commonsourceibias.n480 commonsourceibias.t183 207.983
R6962 commonsourceibias.n364 commonsourceibias.t145 207.983
R6963 commonsourceibias.n127 commonsourceibias.t50 207.983
R6964 commonsourceibias.n249 commonsourceibias.t104 207.983
R6965 commonsourceibias.n963 commonsourceibias.t93 207.983
R6966 commonsourceibias.n847 commonsourceibias.t129 207.983
R6967 commonsourceibias.n617 commonsourceibias.t42 207.983
R6968 commonsourceibias.n732 commonsourceibias.t191 207.983
R6969 commonsourceibias.n396 commonsourceibias.t151 168.701
R6970 commonsourceibias.n402 commonsourceibias.t99 168.701
R6971 commonsourceibias.n408 commonsourceibias.t81 168.701
R6972 commonsourceibias.n392 commonsourceibias.t170 168.701
R6973 commonsourceibias.n416 commonsourceibias.t177 168.701
R6974 commonsourceibias.n422 commonsourceibias.t92 168.701
R6975 commonsourceibias.n387 commonsourceibias.t186 168.701
R6976 commonsourceibias.n430 commonsourceibias.t198 168.701
R6977 commonsourceibias.n436 commonsourceibias.t130 168.701
R6978 commonsourceibias.n382 commonsourceibias.t108 168.701
R6979 commonsourceibias.n444 commonsourceibias.t88 168.701
R6980 commonsourceibias.n450 commonsourceibias.t141 168.701
R6981 commonsourceibias.n377 commonsourceibias.t150 168.701
R6982 commonsourceibias.n458 commonsourceibias.t98 168.701
R6983 commonsourceibias.n464 commonsourceibias.t199 168.701
R6984 commonsourceibias.n372 commonsourceibias.t168 168.701
R6985 commonsourceibias.n472 commonsourceibias.t107 168.701
R6986 commonsourceibias.n478 commonsourceibias.t89 168.701
R6987 commonsourceibias.n362 commonsourceibias.t172 168.701
R6988 commonsourceibias.n356 commonsourceibias.t160 168.701
R6989 commonsourceibias.n256 commonsourceibias.t146 168.701
R6990 commonsourceibias.n348 commonsourceibias.t173 168.701
R6991 commonsourceibias.n342 commonsourceibias.t158 168.701
R6992 commonsourceibias.n261 commonsourceibias.t144 168.701
R6993 commonsourceibias.n334 commonsourceibias.t174 168.701
R6994 commonsourceibias.n328 commonsourceibias.t159 168.701
R6995 commonsourceibias.n266 commonsourceibias.t185 168.701
R6996 commonsourceibias.n320 commonsourceibias.t175 168.701
R6997 commonsourceibias.n314 commonsourceibias.t157 168.701
R6998 commonsourceibias.n271 commonsourceibias.t190 168.701
R6999 commonsourceibias.n306 commonsourceibias.t91 168.701
R7000 commonsourceibias.n300 commonsourceibias.t169 168.701
R7001 commonsourceibias.n276 commonsourceibias.t82 168.701
R7002 commonsourceibias.n292 commonsourceibias.t95 168.701
R7003 commonsourceibias.n286 commonsourceibias.t90 168.701
R7004 commonsourceibias.n280 commonsourceibias.t80 168.701
R7005 commonsourceibias.n125 commonsourceibias.t40 168.701
R7006 commonsourceibias.n119 commonsourceibias.t0 168.701
R7007 commonsourceibias.n19 commonsourceibias.t74 168.701
R7008 commonsourceibias.n111 commonsourceibias.t34 168.701
R7009 commonsourceibias.n105 commonsourceibias.t6 168.701
R7010 commonsourceibias.n24 commonsourceibias.t12 168.701
R7011 commonsourceibias.n97 commonsourceibias.t32 168.701
R7012 commonsourceibias.n91 commonsourceibias.t76 168.701
R7013 commonsourceibias.n29 commonsourceibias.t26 168.701
R7014 commonsourceibias.n83 commonsourceibias.t64 168.701
R7015 commonsourceibias.n77 commonsourceibias.t14 168.701
R7016 commonsourceibias.n34 commonsourceibias.t36 168.701
R7017 commonsourceibias.n69 commonsourceibias.t52 168.701
R7018 commonsourceibias.n63 commonsourceibias.t46 168.701
R7019 commonsourceibias.n39 commonsourceibias.t38 168.701
R7020 commonsourceibias.n55 commonsourceibias.t2 168.701
R7021 commonsourceibias.n49 commonsourceibias.t70 168.701
R7022 commonsourceibias.n43 commonsourceibias.t66 168.701
R7023 commonsourceibias.n247 commonsourceibias.t181 168.701
R7024 commonsourceibias.n241 commonsourceibias.t124 168.701
R7025 commonsourceibias.n5 commonsourceibias.t197 168.701
R7026 commonsourceibias.n233 commonsourceibias.t142 168.701
R7027 commonsourceibias.n227 commonsourceibias.t101 168.701
R7028 commonsourceibias.n10 commonsourceibias.t156 168.701
R7029 commonsourceibias.n219 commonsourceibias.t143 168.701
R7030 commonsourceibias.n213 commonsourceibias.t193 168.701
R7031 commonsourceibias.n150 commonsourceibias.t136 168.701
R7032 commonsourceibias.n151 commonsourceibias.t119 168.701
R7033 commonsourceibias.n153 commonsourceibias.t155 168.701
R7034 commonsourceibias.n155 commonsourceibias.t140 168.701
R7035 commonsourceibias.n191 commonsourceibias.t109 168.701
R7036 commonsourceibias.n185 commonsourceibias.t182 168.701
R7037 commonsourceibias.n161 commonsourceibias.t166 168.701
R7038 commonsourceibias.n177 commonsourceibias.t123 168.701
R7039 commonsourceibias.n171 commonsourceibias.t84 168.701
R7040 commonsourceibias.n165 commonsourceibias.t131 168.701
R7041 commonsourceibias.n874 commonsourceibias.t165 168.701
R7042 commonsourceibias.n880 commonsourceibias.t106 168.701
R7043 commonsourceibias.n886 commonsourceibias.t87 168.701
R7044 commonsourceibias.n888 commonsourceibias.t178 168.701
R7045 commonsourceibias.n895 commonsourceibias.t167 168.701
R7046 commonsourceibias.n901 commonsourceibias.t116 168.701
R7047 commonsourceibias.n903 commonsourceibias.t96 168.701
R7048 commonsourceibias.n910 commonsourceibias.t102 168.701
R7049 commonsourceibias.n916 commonsourceibias.t121 168.701
R7050 commonsourceibias.n918 commonsourceibias.t126 168.701
R7051 commonsourceibias.n925 commonsourceibias.t112 168.701
R7052 commonsourceibias.n931 commonsourceibias.t179 168.701
R7053 commonsourceibias.n933 commonsourceibias.t133 168.701
R7054 commonsourceibias.n940 commonsourceibias.t120 168.701
R7055 commonsourceibias.n946 commonsourceibias.t103 168.701
R7056 commonsourceibias.n948 commonsourceibias.t85 168.701
R7057 commonsourceibias.n955 commonsourceibias.t125 168.701
R7058 commonsourceibias.n961 commonsourceibias.t113 168.701
R7059 commonsourceibias.n758 commonsourceibias.t163 168.701
R7060 commonsourceibias.n764 commonsourceibias.t180 168.701
R7061 commonsourceibias.n770 commonsourceibias.t189 168.701
R7062 commonsourceibias.n772 commonsourceibias.t164 168.701
R7063 commonsourceibias.n779 commonsourceibias.t176 168.701
R7064 commonsourceibias.n785 commonsourceibias.t194 168.701
R7065 commonsourceibias.n787 commonsourceibias.t171 168.701
R7066 commonsourceibias.n794 commonsourceibias.t135 168.701
R7067 commonsourceibias.n800 commonsourceibias.t195 168.701
R7068 commonsourceibias.n802 commonsourceibias.t161 168.701
R7069 commonsourceibias.n809 commonsourceibias.t137 168.701
R7070 commonsourceibias.n815 commonsourceibias.t154 168.701
R7071 commonsourceibias.n817 commonsourceibias.t162 168.701
R7072 commonsourceibias.n824 commonsourceibias.t138 168.701
R7073 commonsourceibias.n830 commonsourceibias.t147 168.701
R7074 commonsourceibias.n832 commonsourceibias.t128 168.701
R7075 commonsourceibias.n839 commonsourceibias.t139 168.701
R7076 commonsourceibias.n845 commonsourceibias.t148 168.701
R7077 commonsourceibias.n528 commonsourceibias.t48 168.701
R7078 commonsourceibias.n534 commonsourceibias.t24 168.701
R7079 commonsourceibias.n540 commonsourceibias.t78 168.701
R7080 commonsourceibias.n542 commonsourceibias.t58 168.701
R7081 commonsourceibias.n549 commonsourceibias.t56 168.701
R7082 commonsourceibias.n555 commonsourceibias.t72 168.701
R7083 commonsourceibias.n557 commonsourceibias.t60 168.701
R7084 commonsourceibias.n564 commonsourceibias.t4 168.701
R7085 commonsourceibias.n570 commonsourceibias.t54 168.701
R7086 commonsourceibias.n572 commonsourceibias.t62 168.701
R7087 commonsourceibias.n579 commonsourceibias.t30 168.701
R7088 commonsourceibias.n585 commonsourceibias.t20 168.701
R7089 commonsourceibias.n587 commonsourceibias.t68 168.701
R7090 commonsourceibias.n594 commonsourceibias.t44 168.701
R7091 commonsourceibias.n600 commonsourceibias.t22 168.701
R7092 commonsourceibias.n602 commonsourceibias.t18 168.701
R7093 commonsourceibias.n609 commonsourceibias.t10 168.701
R7094 commonsourceibias.n615 commonsourceibias.t28 168.701
R7095 commonsourceibias.n730 commonsourceibias.t134 168.701
R7096 commonsourceibias.n724 commonsourceibias.t97 168.701
R7097 commonsourceibias.n717 commonsourceibias.t152 168.701
R7098 commonsourceibias.n715 commonsourceibias.t117 168.701
R7099 commonsourceibias.n709 commonsourceibias.t187 168.701
R7100 commonsourceibias.n702 commonsourceibias.t132 168.701
R7101 commonsourceibias.n700 commonsourceibias.t118 168.701
R7102 commonsourceibias.n694 commonsourceibias.t149 168.701
R7103 commonsourceibias.n687 commonsourceibias.t114 168.701
R7104 commonsourceibias.n644 commonsourceibias.t86 168.701
R7105 commonsourceibias.n650 commonsourceibias.t127 168.701
R7106 commonsourceibias.n656 commonsourceibias.t192 168.701
R7107 commonsourceibias.n658 commonsourceibias.t110 168.701
R7108 commonsourceibias.n665 commonsourceibias.t111 168.701
R7109 commonsourceibias.n671 commonsourceibias.t83 168.701
R7110 commonsourceibias.n635 commonsourceibias.t115 168.701
R7111 commonsourceibias.n633 commonsourceibias.t122 168.701
R7112 commonsourceibias.n631 commonsourceibias.t105 168.701
R7113 commonsourceibias.n479 commonsourceibias.n367 161.3
R7114 commonsourceibias.n477 commonsourceibias.n476 161.3
R7115 commonsourceibias.n475 commonsourceibias.n368 161.3
R7116 commonsourceibias.n474 commonsourceibias.n473 161.3
R7117 commonsourceibias.n471 commonsourceibias.n369 161.3
R7118 commonsourceibias.n470 commonsourceibias.n469 161.3
R7119 commonsourceibias.n468 commonsourceibias.n370 161.3
R7120 commonsourceibias.n467 commonsourceibias.n466 161.3
R7121 commonsourceibias.n465 commonsourceibias.n371 161.3
R7122 commonsourceibias.n463 commonsourceibias.n462 161.3
R7123 commonsourceibias.n461 commonsourceibias.n373 161.3
R7124 commonsourceibias.n460 commonsourceibias.n459 161.3
R7125 commonsourceibias.n457 commonsourceibias.n374 161.3
R7126 commonsourceibias.n456 commonsourceibias.n455 161.3
R7127 commonsourceibias.n454 commonsourceibias.n375 161.3
R7128 commonsourceibias.n453 commonsourceibias.n452 161.3
R7129 commonsourceibias.n451 commonsourceibias.n376 161.3
R7130 commonsourceibias.n449 commonsourceibias.n448 161.3
R7131 commonsourceibias.n447 commonsourceibias.n378 161.3
R7132 commonsourceibias.n446 commonsourceibias.n445 161.3
R7133 commonsourceibias.n443 commonsourceibias.n379 161.3
R7134 commonsourceibias.n442 commonsourceibias.n441 161.3
R7135 commonsourceibias.n440 commonsourceibias.n380 161.3
R7136 commonsourceibias.n439 commonsourceibias.n438 161.3
R7137 commonsourceibias.n437 commonsourceibias.n381 161.3
R7138 commonsourceibias.n435 commonsourceibias.n434 161.3
R7139 commonsourceibias.n433 commonsourceibias.n383 161.3
R7140 commonsourceibias.n432 commonsourceibias.n431 161.3
R7141 commonsourceibias.n429 commonsourceibias.n384 161.3
R7142 commonsourceibias.n428 commonsourceibias.n427 161.3
R7143 commonsourceibias.n426 commonsourceibias.n385 161.3
R7144 commonsourceibias.n425 commonsourceibias.n424 161.3
R7145 commonsourceibias.n423 commonsourceibias.n386 161.3
R7146 commonsourceibias.n421 commonsourceibias.n420 161.3
R7147 commonsourceibias.n419 commonsourceibias.n388 161.3
R7148 commonsourceibias.n418 commonsourceibias.n417 161.3
R7149 commonsourceibias.n415 commonsourceibias.n389 161.3
R7150 commonsourceibias.n414 commonsourceibias.n413 161.3
R7151 commonsourceibias.n412 commonsourceibias.n390 161.3
R7152 commonsourceibias.n411 commonsourceibias.n410 161.3
R7153 commonsourceibias.n409 commonsourceibias.n391 161.3
R7154 commonsourceibias.n407 commonsourceibias.n406 161.3
R7155 commonsourceibias.n405 commonsourceibias.n393 161.3
R7156 commonsourceibias.n404 commonsourceibias.n403 161.3
R7157 commonsourceibias.n401 commonsourceibias.n394 161.3
R7158 commonsourceibias.n400 commonsourceibias.n399 161.3
R7159 commonsourceibias.n398 commonsourceibias.n395 161.3
R7160 commonsourceibias.n282 commonsourceibias.n279 161.3
R7161 commonsourceibias.n284 commonsourceibias.n283 161.3
R7162 commonsourceibias.n285 commonsourceibias.n278 161.3
R7163 commonsourceibias.n288 commonsourceibias.n287 161.3
R7164 commonsourceibias.n289 commonsourceibias.n277 161.3
R7165 commonsourceibias.n291 commonsourceibias.n290 161.3
R7166 commonsourceibias.n293 commonsourceibias.n275 161.3
R7167 commonsourceibias.n295 commonsourceibias.n294 161.3
R7168 commonsourceibias.n296 commonsourceibias.n274 161.3
R7169 commonsourceibias.n298 commonsourceibias.n297 161.3
R7170 commonsourceibias.n299 commonsourceibias.n273 161.3
R7171 commonsourceibias.n302 commonsourceibias.n301 161.3
R7172 commonsourceibias.n303 commonsourceibias.n272 161.3
R7173 commonsourceibias.n305 commonsourceibias.n304 161.3
R7174 commonsourceibias.n307 commonsourceibias.n270 161.3
R7175 commonsourceibias.n309 commonsourceibias.n308 161.3
R7176 commonsourceibias.n310 commonsourceibias.n269 161.3
R7177 commonsourceibias.n312 commonsourceibias.n311 161.3
R7178 commonsourceibias.n313 commonsourceibias.n268 161.3
R7179 commonsourceibias.n316 commonsourceibias.n315 161.3
R7180 commonsourceibias.n317 commonsourceibias.n267 161.3
R7181 commonsourceibias.n319 commonsourceibias.n318 161.3
R7182 commonsourceibias.n321 commonsourceibias.n265 161.3
R7183 commonsourceibias.n323 commonsourceibias.n322 161.3
R7184 commonsourceibias.n324 commonsourceibias.n264 161.3
R7185 commonsourceibias.n326 commonsourceibias.n325 161.3
R7186 commonsourceibias.n327 commonsourceibias.n263 161.3
R7187 commonsourceibias.n330 commonsourceibias.n329 161.3
R7188 commonsourceibias.n331 commonsourceibias.n262 161.3
R7189 commonsourceibias.n333 commonsourceibias.n332 161.3
R7190 commonsourceibias.n335 commonsourceibias.n260 161.3
R7191 commonsourceibias.n337 commonsourceibias.n336 161.3
R7192 commonsourceibias.n338 commonsourceibias.n259 161.3
R7193 commonsourceibias.n340 commonsourceibias.n339 161.3
R7194 commonsourceibias.n341 commonsourceibias.n258 161.3
R7195 commonsourceibias.n344 commonsourceibias.n343 161.3
R7196 commonsourceibias.n345 commonsourceibias.n257 161.3
R7197 commonsourceibias.n347 commonsourceibias.n346 161.3
R7198 commonsourceibias.n349 commonsourceibias.n255 161.3
R7199 commonsourceibias.n351 commonsourceibias.n350 161.3
R7200 commonsourceibias.n352 commonsourceibias.n254 161.3
R7201 commonsourceibias.n354 commonsourceibias.n353 161.3
R7202 commonsourceibias.n355 commonsourceibias.n253 161.3
R7203 commonsourceibias.n358 commonsourceibias.n357 161.3
R7204 commonsourceibias.n359 commonsourceibias.n252 161.3
R7205 commonsourceibias.n361 commonsourceibias.n360 161.3
R7206 commonsourceibias.n363 commonsourceibias.n251 161.3
R7207 commonsourceibias.n45 commonsourceibias.n42 161.3
R7208 commonsourceibias.n47 commonsourceibias.n46 161.3
R7209 commonsourceibias.n48 commonsourceibias.n41 161.3
R7210 commonsourceibias.n51 commonsourceibias.n50 161.3
R7211 commonsourceibias.n52 commonsourceibias.n40 161.3
R7212 commonsourceibias.n54 commonsourceibias.n53 161.3
R7213 commonsourceibias.n56 commonsourceibias.n38 161.3
R7214 commonsourceibias.n58 commonsourceibias.n57 161.3
R7215 commonsourceibias.n59 commonsourceibias.n37 161.3
R7216 commonsourceibias.n61 commonsourceibias.n60 161.3
R7217 commonsourceibias.n62 commonsourceibias.n36 161.3
R7218 commonsourceibias.n65 commonsourceibias.n64 161.3
R7219 commonsourceibias.n66 commonsourceibias.n35 161.3
R7220 commonsourceibias.n68 commonsourceibias.n67 161.3
R7221 commonsourceibias.n70 commonsourceibias.n33 161.3
R7222 commonsourceibias.n72 commonsourceibias.n71 161.3
R7223 commonsourceibias.n73 commonsourceibias.n32 161.3
R7224 commonsourceibias.n75 commonsourceibias.n74 161.3
R7225 commonsourceibias.n76 commonsourceibias.n31 161.3
R7226 commonsourceibias.n79 commonsourceibias.n78 161.3
R7227 commonsourceibias.n80 commonsourceibias.n30 161.3
R7228 commonsourceibias.n82 commonsourceibias.n81 161.3
R7229 commonsourceibias.n84 commonsourceibias.n28 161.3
R7230 commonsourceibias.n86 commonsourceibias.n85 161.3
R7231 commonsourceibias.n87 commonsourceibias.n27 161.3
R7232 commonsourceibias.n89 commonsourceibias.n88 161.3
R7233 commonsourceibias.n90 commonsourceibias.n26 161.3
R7234 commonsourceibias.n93 commonsourceibias.n92 161.3
R7235 commonsourceibias.n94 commonsourceibias.n25 161.3
R7236 commonsourceibias.n96 commonsourceibias.n95 161.3
R7237 commonsourceibias.n98 commonsourceibias.n23 161.3
R7238 commonsourceibias.n100 commonsourceibias.n99 161.3
R7239 commonsourceibias.n101 commonsourceibias.n22 161.3
R7240 commonsourceibias.n103 commonsourceibias.n102 161.3
R7241 commonsourceibias.n104 commonsourceibias.n21 161.3
R7242 commonsourceibias.n107 commonsourceibias.n106 161.3
R7243 commonsourceibias.n108 commonsourceibias.n20 161.3
R7244 commonsourceibias.n110 commonsourceibias.n109 161.3
R7245 commonsourceibias.n112 commonsourceibias.n18 161.3
R7246 commonsourceibias.n114 commonsourceibias.n113 161.3
R7247 commonsourceibias.n115 commonsourceibias.n17 161.3
R7248 commonsourceibias.n117 commonsourceibias.n116 161.3
R7249 commonsourceibias.n118 commonsourceibias.n16 161.3
R7250 commonsourceibias.n121 commonsourceibias.n120 161.3
R7251 commonsourceibias.n122 commonsourceibias.n15 161.3
R7252 commonsourceibias.n124 commonsourceibias.n123 161.3
R7253 commonsourceibias.n126 commonsourceibias.n14 161.3
R7254 commonsourceibias.n167 commonsourceibias.n164 161.3
R7255 commonsourceibias.n169 commonsourceibias.n168 161.3
R7256 commonsourceibias.n170 commonsourceibias.n163 161.3
R7257 commonsourceibias.n173 commonsourceibias.n172 161.3
R7258 commonsourceibias.n174 commonsourceibias.n162 161.3
R7259 commonsourceibias.n176 commonsourceibias.n175 161.3
R7260 commonsourceibias.n178 commonsourceibias.n160 161.3
R7261 commonsourceibias.n180 commonsourceibias.n179 161.3
R7262 commonsourceibias.n181 commonsourceibias.n159 161.3
R7263 commonsourceibias.n183 commonsourceibias.n182 161.3
R7264 commonsourceibias.n184 commonsourceibias.n158 161.3
R7265 commonsourceibias.n187 commonsourceibias.n186 161.3
R7266 commonsourceibias.n188 commonsourceibias.n157 161.3
R7267 commonsourceibias.n190 commonsourceibias.n189 161.3
R7268 commonsourceibias.n192 commonsourceibias.n156 161.3
R7269 commonsourceibias.n194 commonsourceibias.n193 161.3
R7270 commonsourceibias.n196 commonsourceibias.n195 161.3
R7271 commonsourceibias.n197 commonsourceibias.n154 161.3
R7272 commonsourceibias.n199 commonsourceibias.n198 161.3
R7273 commonsourceibias.n201 commonsourceibias.n200 161.3
R7274 commonsourceibias.n202 commonsourceibias.n152 161.3
R7275 commonsourceibias.n204 commonsourceibias.n203 161.3
R7276 commonsourceibias.n206 commonsourceibias.n205 161.3
R7277 commonsourceibias.n208 commonsourceibias.n207 161.3
R7278 commonsourceibias.n209 commonsourceibias.n13 161.3
R7279 commonsourceibias.n211 commonsourceibias.n210 161.3
R7280 commonsourceibias.n212 commonsourceibias.n12 161.3
R7281 commonsourceibias.n215 commonsourceibias.n214 161.3
R7282 commonsourceibias.n216 commonsourceibias.n11 161.3
R7283 commonsourceibias.n218 commonsourceibias.n217 161.3
R7284 commonsourceibias.n220 commonsourceibias.n9 161.3
R7285 commonsourceibias.n222 commonsourceibias.n221 161.3
R7286 commonsourceibias.n223 commonsourceibias.n8 161.3
R7287 commonsourceibias.n225 commonsourceibias.n224 161.3
R7288 commonsourceibias.n226 commonsourceibias.n7 161.3
R7289 commonsourceibias.n229 commonsourceibias.n228 161.3
R7290 commonsourceibias.n230 commonsourceibias.n6 161.3
R7291 commonsourceibias.n232 commonsourceibias.n231 161.3
R7292 commonsourceibias.n234 commonsourceibias.n4 161.3
R7293 commonsourceibias.n236 commonsourceibias.n235 161.3
R7294 commonsourceibias.n237 commonsourceibias.n3 161.3
R7295 commonsourceibias.n239 commonsourceibias.n238 161.3
R7296 commonsourceibias.n240 commonsourceibias.n2 161.3
R7297 commonsourceibias.n243 commonsourceibias.n242 161.3
R7298 commonsourceibias.n244 commonsourceibias.n1 161.3
R7299 commonsourceibias.n246 commonsourceibias.n245 161.3
R7300 commonsourceibias.n248 commonsourceibias.n0 161.3
R7301 commonsourceibias.n962 commonsourceibias.n850 161.3
R7302 commonsourceibias.n960 commonsourceibias.n959 161.3
R7303 commonsourceibias.n958 commonsourceibias.n851 161.3
R7304 commonsourceibias.n957 commonsourceibias.n956 161.3
R7305 commonsourceibias.n954 commonsourceibias.n852 161.3
R7306 commonsourceibias.n953 commonsourceibias.n952 161.3
R7307 commonsourceibias.n951 commonsourceibias.n853 161.3
R7308 commonsourceibias.n950 commonsourceibias.n949 161.3
R7309 commonsourceibias.n947 commonsourceibias.n854 161.3
R7310 commonsourceibias.n945 commonsourceibias.n944 161.3
R7311 commonsourceibias.n943 commonsourceibias.n855 161.3
R7312 commonsourceibias.n942 commonsourceibias.n941 161.3
R7313 commonsourceibias.n939 commonsourceibias.n856 161.3
R7314 commonsourceibias.n938 commonsourceibias.n937 161.3
R7315 commonsourceibias.n936 commonsourceibias.n857 161.3
R7316 commonsourceibias.n935 commonsourceibias.n934 161.3
R7317 commonsourceibias.n932 commonsourceibias.n858 161.3
R7318 commonsourceibias.n930 commonsourceibias.n929 161.3
R7319 commonsourceibias.n928 commonsourceibias.n859 161.3
R7320 commonsourceibias.n927 commonsourceibias.n926 161.3
R7321 commonsourceibias.n924 commonsourceibias.n860 161.3
R7322 commonsourceibias.n923 commonsourceibias.n922 161.3
R7323 commonsourceibias.n921 commonsourceibias.n861 161.3
R7324 commonsourceibias.n920 commonsourceibias.n919 161.3
R7325 commonsourceibias.n917 commonsourceibias.n862 161.3
R7326 commonsourceibias.n915 commonsourceibias.n914 161.3
R7327 commonsourceibias.n913 commonsourceibias.n863 161.3
R7328 commonsourceibias.n912 commonsourceibias.n911 161.3
R7329 commonsourceibias.n909 commonsourceibias.n864 161.3
R7330 commonsourceibias.n908 commonsourceibias.n907 161.3
R7331 commonsourceibias.n906 commonsourceibias.n865 161.3
R7332 commonsourceibias.n905 commonsourceibias.n904 161.3
R7333 commonsourceibias.n902 commonsourceibias.n866 161.3
R7334 commonsourceibias.n900 commonsourceibias.n899 161.3
R7335 commonsourceibias.n898 commonsourceibias.n867 161.3
R7336 commonsourceibias.n897 commonsourceibias.n896 161.3
R7337 commonsourceibias.n894 commonsourceibias.n868 161.3
R7338 commonsourceibias.n893 commonsourceibias.n892 161.3
R7339 commonsourceibias.n891 commonsourceibias.n869 161.3
R7340 commonsourceibias.n890 commonsourceibias.n889 161.3
R7341 commonsourceibias.n887 commonsourceibias.n870 161.3
R7342 commonsourceibias.n885 commonsourceibias.n884 161.3
R7343 commonsourceibias.n883 commonsourceibias.n871 161.3
R7344 commonsourceibias.n882 commonsourceibias.n881 161.3
R7345 commonsourceibias.n879 commonsourceibias.n872 161.3
R7346 commonsourceibias.n878 commonsourceibias.n877 161.3
R7347 commonsourceibias.n876 commonsourceibias.n873 161.3
R7348 commonsourceibias.n846 commonsourceibias.n734 161.3
R7349 commonsourceibias.n844 commonsourceibias.n843 161.3
R7350 commonsourceibias.n842 commonsourceibias.n735 161.3
R7351 commonsourceibias.n841 commonsourceibias.n840 161.3
R7352 commonsourceibias.n838 commonsourceibias.n736 161.3
R7353 commonsourceibias.n837 commonsourceibias.n836 161.3
R7354 commonsourceibias.n835 commonsourceibias.n737 161.3
R7355 commonsourceibias.n834 commonsourceibias.n833 161.3
R7356 commonsourceibias.n831 commonsourceibias.n738 161.3
R7357 commonsourceibias.n829 commonsourceibias.n828 161.3
R7358 commonsourceibias.n827 commonsourceibias.n739 161.3
R7359 commonsourceibias.n826 commonsourceibias.n825 161.3
R7360 commonsourceibias.n823 commonsourceibias.n740 161.3
R7361 commonsourceibias.n822 commonsourceibias.n821 161.3
R7362 commonsourceibias.n820 commonsourceibias.n741 161.3
R7363 commonsourceibias.n819 commonsourceibias.n818 161.3
R7364 commonsourceibias.n816 commonsourceibias.n742 161.3
R7365 commonsourceibias.n814 commonsourceibias.n813 161.3
R7366 commonsourceibias.n812 commonsourceibias.n743 161.3
R7367 commonsourceibias.n811 commonsourceibias.n810 161.3
R7368 commonsourceibias.n808 commonsourceibias.n744 161.3
R7369 commonsourceibias.n807 commonsourceibias.n806 161.3
R7370 commonsourceibias.n805 commonsourceibias.n745 161.3
R7371 commonsourceibias.n804 commonsourceibias.n803 161.3
R7372 commonsourceibias.n801 commonsourceibias.n746 161.3
R7373 commonsourceibias.n799 commonsourceibias.n798 161.3
R7374 commonsourceibias.n797 commonsourceibias.n747 161.3
R7375 commonsourceibias.n796 commonsourceibias.n795 161.3
R7376 commonsourceibias.n793 commonsourceibias.n748 161.3
R7377 commonsourceibias.n792 commonsourceibias.n791 161.3
R7378 commonsourceibias.n790 commonsourceibias.n749 161.3
R7379 commonsourceibias.n789 commonsourceibias.n788 161.3
R7380 commonsourceibias.n786 commonsourceibias.n750 161.3
R7381 commonsourceibias.n784 commonsourceibias.n783 161.3
R7382 commonsourceibias.n782 commonsourceibias.n751 161.3
R7383 commonsourceibias.n781 commonsourceibias.n780 161.3
R7384 commonsourceibias.n778 commonsourceibias.n752 161.3
R7385 commonsourceibias.n777 commonsourceibias.n776 161.3
R7386 commonsourceibias.n775 commonsourceibias.n753 161.3
R7387 commonsourceibias.n774 commonsourceibias.n773 161.3
R7388 commonsourceibias.n771 commonsourceibias.n754 161.3
R7389 commonsourceibias.n769 commonsourceibias.n768 161.3
R7390 commonsourceibias.n767 commonsourceibias.n755 161.3
R7391 commonsourceibias.n766 commonsourceibias.n765 161.3
R7392 commonsourceibias.n763 commonsourceibias.n756 161.3
R7393 commonsourceibias.n762 commonsourceibias.n761 161.3
R7394 commonsourceibias.n760 commonsourceibias.n757 161.3
R7395 commonsourceibias.n616 commonsourceibias.n504 161.3
R7396 commonsourceibias.n614 commonsourceibias.n613 161.3
R7397 commonsourceibias.n612 commonsourceibias.n505 161.3
R7398 commonsourceibias.n611 commonsourceibias.n610 161.3
R7399 commonsourceibias.n608 commonsourceibias.n506 161.3
R7400 commonsourceibias.n607 commonsourceibias.n606 161.3
R7401 commonsourceibias.n605 commonsourceibias.n507 161.3
R7402 commonsourceibias.n604 commonsourceibias.n603 161.3
R7403 commonsourceibias.n601 commonsourceibias.n508 161.3
R7404 commonsourceibias.n599 commonsourceibias.n598 161.3
R7405 commonsourceibias.n597 commonsourceibias.n509 161.3
R7406 commonsourceibias.n596 commonsourceibias.n595 161.3
R7407 commonsourceibias.n593 commonsourceibias.n510 161.3
R7408 commonsourceibias.n592 commonsourceibias.n591 161.3
R7409 commonsourceibias.n590 commonsourceibias.n511 161.3
R7410 commonsourceibias.n589 commonsourceibias.n588 161.3
R7411 commonsourceibias.n586 commonsourceibias.n512 161.3
R7412 commonsourceibias.n584 commonsourceibias.n583 161.3
R7413 commonsourceibias.n582 commonsourceibias.n513 161.3
R7414 commonsourceibias.n581 commonsourceibias.n580 161.3
R7415 commonsourceibias.n578 commonsourceibias.n514 161.3
R7416 commonsourceibias.n577 commonsourceibias.n576 161.3
R7417 commonsourceibias.n575 commonsourceibias.n515 161.3
R7418 commonsourceibias.n574 commonsourceibias.n573 161.3
R7419 commonsourceibias.n571 commonsourceibias.n516 161.3
R7420 commonsourceibias.n569 commonsourceibias.n568 161.3
R7421 commonsourceibias.n567 commonsourceibias.n517 161.3
R7422 commonsourceibias.n566 commonsourceibias.n565 161.3
R7423 commonsourceibias.n563 commonsourceibias.n518 161.3
R7424 commonsourceibias.n562 commonsourceibias.n561 161.3
R7425 commonsourceibias.n560 commonsourceibias.n519 161.3
R7426 commonsourceibias.n559 commonsourceibias.n558 161.3
R7427 commonsourceibias.n556 commonsourceibias.n520 161.3
R7428 commonsourceibias.n554 commonsourceibias.n553 161.3
R7429 commonsourceibias.n552 commonsourceibias.n521 161.3
R7430 commonsourceibias.n551 commonsourceibias.n550 161.3
R7431 commonsourceibias.n548 commonsourceibias.n522 161.3
R7432 commonsourceibias.n547 commonsourceibias.n546 161.3
R7433 commonsourceibias.n545 commonsourceibias.n523 161.3
R7434 commonsourceibias.n544 commonsourceibias.n543 161.3
R7435 commonsourceibias.n541 commonsourceibias.n524 161.3
R7436 commonsourceibias.n539 commonsourceibias.n538 161.3
R7437 commonsourceibias.n537 commonsourceibias.n525 161.3
R7438 commonsourceibias.n536 commonsourceibias.n535 161.3
R7439 commonsourceibias.n533 commonsourceibias.n526 161.3
R7440 commonsourceibias.n532 commonsourceibias.n531 161.3
R7441 commonsourceibias.n530 commonsourceibias.n527 161.3
R7442 commonsourceibias.n686 commonsourceibias.n685 161.3
R7443 commonsourceibias.n684 commonsourceibias.n683 161.3
R7444 commonsourceibias.n682 commonsourceibias.n632 161.3
R7445 commonsourceibias.n681 commonsourceibias.n680 161.3
R7446 commonsourceibias.n679 commonsourceibias.n678 161.3
R7447 commonsourceibias.n677 commonsourceibias.n634 161.3
R7448 commonsourceibias.n676 commonsourceibias.n675 161.3
R7449 commonsourceibias.n674 commonsourceibias.n673 161.3
R7450 commonsourceibias.n672 commonsourceibias.n636 161.3
R7451 commonsourceibias.n670 commonsourceibias.n669 161.3
R7452 commonsourceibias.n668 commonsourceibias.n637 161.3
R7453 commonsourceibias.n667 commonsourceibias.n666 161.3
R7454 commonsourceibias.n664 commonsourceibias.n638 161.3
R7455 commonsourceibias.n663 commonsourceibias.n662 161.3
R7456 commonsourceibias.n661 commonsourceibias.n639 161.3
R7457 commonsourceibias.n660 commonsourceibias.n659 161.3
R7458 commonsourceibias.n657 commonsourceibias.n640 161.3
R7459 commonsourceibias.n655 commonsourceibias.n654 161.3
R7460 commonsourceibias.n653 commonsourceibias.n641 161.3
R7461 commonsourceibias.n652 commonsourceibias.n651 161.3
R7462 commonsourceibias.n649 commonsourceibias.n642 161.3
R7463 commonsourceibias.n648 commonsourceibias.n647 161.3
R7464 commonsourceibias.n646 commonsourceibias.n643 161.3
R7465 commonsourceibias.n731 commonsourceibias.n483 161.3
R7466 commonsourceibias.n729 commonsourceibias.n728 161.3
R7467 commonsourceibias.n727 commonsourceibias.n484 161.3
R7468 commonsourceibias.n726 commonsourceibias.n725 161.3
R7469 commonsourceibias.n723 commonsourceibias.n485 161.3
R7470 commonsourceibias.n722 commonsourceibias.n721 161.3
R7471 commonsourceibias.n720 commonsourceibias.n486 161.3
R7472 commonsourceibias.n719 commonsourceibias.n718 161.3
R7473 commonsourceibias.n716 commonsourceibias.n487 161.3
R7474 commonsourceibias.n714 commonsourceibias.n713 161.3
R7475 commonsourceibias.n712 commonsourceibias.n488 161.3
R7476 commonsourceibias.n711 commonsourceibias.n710 161.3
R7477 commonsourceibias.n708 commonsourceibias.n489 161.3
R7478 commonsourceibias.n707 commonsourceibias.n706 161.3
R7479 commonsourceibias.n705 commonsourceibias.n490 161.3
R7480 commonsourceibias.n704 commonsourceibias.n703 161.3
R7481 commonsourceibias.n701 commonsourceibias.n491 161.3
R7482 commonsourceibias.n699 commonsourceibias.n698 161.3
R7483 commonsourceibias.n697 commonsourceibias.n492 161.3
R7484 commonsourceibias.n696 commonsourceibias.n695 161.3
R7485 commonsourceibias.n693 commonsourceibias.n493 161.3
R7486 commonsourceibias.n692 commonsourceibias.n691 161.3
R7487 commonsourceibias.n690 commonsourceibias.n494 161.3
R7488 commonsourceibias.n689 commonsourceibias.n688 161.3
R7489 commonsourceibias.n141 commonsourceibias.n139 81.5057
R7490 commonsourceibias.n497 commonsourceibias.n495 81.5057
R7491 commonsourceibias.n141 commonsourceibias.n140 80.9324
R7492 commonsourceibias.n143 commonsourceibias.n142 80.9324
R7493 commonsourceibias.n145 commonsourceibias.n144 80.9324
R7494 commonsourceibias.n147 commonsourceibias.n146 80.9324
R7495 commonsourceibias.n138 commonsourceibias.n137 80.9324
R7496 commonsourceibias.n136 commonsourceibias.n135 80.9324
R7497 commonsourceibias.n134 commonsourceibias.n133 80.9324
R7498 commonsourceibias.n132 commonsourceibias.n131 80.9324
R7499 commonsourceibias.n130 commonsourceibias.n129 80.9324
R7500 commonsourceibias.n620 commonsourceibias.n619 80.9324
R7501 commonsourceibias.n622 commonsourceibias.n621 80.9324
R7502 commonsourceibias.n624 commonsourceibias.n623 80.9324
R7503 commonsourceibias.n626 commonsourceibias.n625 80.9324
R7504 commonsourceibias.n628 commonsourceibias.n627 80.9324
R7505 commonsourceibias.n503 commonsourceibias.n502 80.9324
R7506 commonsourceibias.n501 commonsourceibias.n500 80.9324
R7507 commonsourceibias.n499 commonsourceibias.n498 80.9324
R7508 commonsourceibias.n497 commonsourceibias.n496 80.9324
R7509 commonsourceibias.n481 commonsourceibias.n480 80.6037
R7510 commonsourceibias.n365 commonsourceibias.n364 80.6037
R7511 commonsourceibias.n128 commonsourceibias.n127 80.6037
R7512 commonsourceibias.n250 commonsourceibias.n249 80.6037
R7513 commonsourceibias.n964 commonsourceibias.n963 80.6037
R7514 commonsourceibias.n848 commonsourceibias.n847 80.6037
R7515 commonsourceibias.n618 commonsourceibias.n617 80.6037
R7516 commonsourceibias.n733 commonsourceibias.n732 80.6037
R7517 commonsourceibias.n438 commonsourceibias.n437 56.5617
R7518 commonsourceibias.n452 commonsourceibias.n451 56.5617
R7519 commonsourceibias.n322 commonsourceibias.n321 56.5617
R7520 commonsourceibias.n308 commonsourceibias.n307 56.5617
R7521 commonsourceibias.n85 commonsourceibias.n84 56.5617
R7522 commonsourceibias.n71 commonsourceibias.n70 56.5617
R7523 commonsourceibias.n207 commonsourceibias.n206 56.5617
R7524 commonsourceibias.n193 commonsourceibias.n192 56.5617
R7525 commonsourceibias.n919 commonsourceibias.n917 56.5617
R7526 commonsourceibias.n934 commonsourceibias.n932 56.5617
R7527 commonsourceibias.n803 commonsourceibias.n801 56.5617
R7528 commonsourceibias.n818 commonsourceibias.n816 56.5617
R7529 commonsourceibias.n573 commonsourceibias.n571 56.5617
R7530 commonsourceibias.n588 commonsourceibias.n586 56.5617
R7531 commonsourceibias.n688 commonsourceibias.n686 56.5617
R7532 commonsourceibias.n410 commonsourceibias.n409 56.5617
R7533 commonsourceibias.n424 commonsourceibias.n423 56.5617
R7534 commonsourceibias.n466 commonsourceibias.n465 56.5617
R7535 commonsourceibias.n350 commonsourceibias.n349 56.5617
R7536 commonsourceibias.n336 commonsourceibias.n335 56.5617
R7537 commonsourceibias.n294 commonsourceibias.n293 56.5617
R7538 commonsourceibias.n113 commonsourceibias.n112 56.5617
R7539 commonsourceibias.n99 commonsourceibias.n98 56.5617
R7540 commonsourceibias.n57 commonsourceibias.n56 56.5617
R7541 commonsourceibias.n235 commonsourceibias.n234 56.5617
R7542 commonsourceibias.n221 commonsourceibias.n220 56.5617
R7543 commonsourceibias.n179 commonsourceibias.n178 56.5617
R7544 commonsourceibias.n889 commonsourceibias.n887 56.5617
R7545 commonsourceibias.n904 commonsourceibias.n902 56.5617
R7546 commonsourceibias.n949 commonsourceibias.n947 56.5617
R7547 commonsourceibias.n773 commonsourceibias.n771 56.5617
R7548 commonsourceibias.n788 commonsourceibias.n786 56.5617
R7549 commonsourceibias.n833 commonsourceibias.n831 56.5617
R7550 commonsourceibias.n543 commonsourceibias.n541 56.5617
R7551 commonsourceibias.n558 commonsourceibias.n556 56.5617
R7552 commonsourceibias.n603 commonsourceibias.n601 56.5617
R7553 commonsourceibias.n718 commonsourceibias.n716 56.5617
R7554 commonsourceibias.n703 commonsourceibias.n701 56.5617
R7555 commonsourceibias.n659 commonsourceibias.n657 56.5617
R7556 commonsourceibias.n673 commonsourceibias.n672 56.5617
R7557 commonsourceibias.n401 commonsourceibias.n400 51.2335
R7558 commonsourceibias.n473 commonsourceibias.n368 51.2335
R7559 commonsourceibias.n357 commonsourceibias.n252 51.2335
R7560 commonsourceibias.n285 commonsourceibias.n284 51.2335
R7561 commonsourceibias.n120 commonsourceibias.n15 51.2335
R7562 commonsourceibias.n48 commonsourceibias.n47 51.2335
R7563 commonsourceibias.n242 commonsourceibias.n1 51.2335
R7564 commonsourceibias.n170 commonsourceibias.n169 51.2335
R7565 commonsourceibias.n879 commonsourceibias.n878 51.2335
R7566 commonsourceibias.n956 commonsourceibias.n851 51.2335
R7567 commonsourceibias.n763 commonsourceibias.n762 51.2335
R7568 commonsourceibias.n840 commonsourceibias.n735 51.2335
R7569 commonsourceibias.n533 commonsourceibias.n532 51.2335
R7570 commonsourceibias.n610 commonsourceibias.n505 51.2335
R7571 commonsourceibias.n725 commonsourceibias.n484 51.2335
R7572 commonsourceibias.n649 commonsourceibias.n648 51.2335
R7573 commonsourceibias.n480 commonsourceibias.n479 50.9056
R7574 commonsourceibias.n364 commonsourceibias.n363 50.9056
R7575 commonsourceibias.n127 commonsourceibias.n126 50.9056
R7576 commonsourceibias.n249 commonsourceibias.n248 50.9056
R7577 commonsourceibias.n963 commonsourceibias.n962 50.9056
R7578 commonsourceibias.n847 commonsourceibias.n846 50.9056
R7579 commonsourceibias.n617 commonsourceibias.n616 50.9056
R7580 commonsourceibias.n732 commonsourceibias.n731 50.9056
R7581 commonsourceibias.n415 commonsourceibias.n414 50.2647
R7582 commonsourceibias.n459 commonsourceibias.n373 50.2647
R7583 commonsourceibias.n343 commonsourceibias.n257 50.2647
R7584 commonsourceibias.n299 commonsourceibias.n298 50.2647
R7585 commonsourceibias.n106 commonsourceibias.n20 50.2647
R7586 commonsourceibias.n62 commonsourceibias.n61 50.2647
R7587 commonsourceibias.n228 commonsourceibias.n6 50.2647
R7588 commonsourceibias.n184 commonsourceibias.n183 50.2647
R7589 commonsourceibias.n894 commonsourceibias.n893 50.2647
R7590 commonsourceibias.n941 commonsourceibias.n855 50.2647
R7591 commonsourceibias.n778 commonsourceibias.n777 50.2647
R7592 commonsourceibias.n825 commonsourceibias.n739 50.2647
R7593 commonsourceibias.n548 commonsourceibias.n547 50.2647
R7594 commonsourceibias.n595 commonsourceibias.n509 50.2647
R7595 commonsourceibias.n710 commonsourceibias.n488 50.2647
R7596 commonsourceibias.n664 commonsourceibias.n663 50.2647
R7597 commonsourceibias.n397 commonsourceibias.n396 49.9027
R7598 commonsourceibias.n281 commonsourceibias.n280 49.9027
R7599 commonsourceibias.n44 commonsourceibias.n43 49.9027
R7600 commonsourceibias.n166 commonsourceibias.n165 49.9027
R7601 commonsourceibias.n875 commonsourceibias.n874 49.9027
R7602 commonsourceibias.n759 commonsourceibias.n758 49.9027
R7603 commonsourceibias.n529 commonsourceibias.n528 49.9027
R7604 commonsourceibias.n645 commonsourceibias.n644 49.9027
R7605 commonsourceibias.n429 commonsourceibias.n428 49.296
R7606 commonsourceibias.n445 commonsourceibias.n378 49.296
R7607 commonsourceibias.n329 commonsourceibias.n262 49.296
R7608 commonsourceibias.n313 commonsourceibias.n312 49.296
R7609 commonsourceibias.n92 commonsourceibias.n25 49.296
R7610 commonsourceibias.n76 commonsourceibias.n75 49.296
R7611 commonsourceibias.n214 commonsourceibias.n11 49.296
R7612 commonsourceibias.n198 commonsourceibias.n197 49.296
R7613 commonsourceibias.n909 commonsourceibias.n908 49.296
R7614 commonsourceibias.n926 commonsourceibias.n859 49.296
R7615 commonsourceibias.n793 commonsourceibias.n792 49.296
R7616 commonsourceibias.n810 commonsourceibias.n743 49.296
R7617 commonsourceibias.n563 commonsourceibias.n562 49.296
R7618 commonsourceibias.n580 commonsourceibias.n513 49.296
R7619 commonsourceibias.n695 commonsourceibias.n492 49.296
R7620 commonsourceibias.n678 commonsourceibias.n677 49.296
R7621 commonsourceibias.n431 commonsourceibias.n383 48.3272
R7622 commonsourceibias.n443 commonsourceibias.n442 48.3272
R7623 commonsourceibias.n327 commonsourceibias.n326 48.3272
R7624 commonsourceibias.n315 commonsourceibias.n267 48.3272
R7625 commonsourceibias.n90 commonsourceibias.n89 48.3272
R7626 commonsourceibias.n78 commonsourceibias.n30 48.3272
R7627 commonsourceibias.n212 commonsourceibias.n211 48.3272
R7628 commonsourceibias.n202 commonsourceibias.n201 48.3272
R7629 commonsourceibias.n911 commonsourceibias.n863 48.3272
R7630 commonsourceibias.n924 commonsourceibias.n923 48.3272
R7631 commonsourceibias.n795 commonsourceibias.n747 48.3272
R7632 commonsourceibias.n808 commonsourceibias.n807 48.3272
R7633 commonsourceibias.n565 commonsourceibias.n517 48.3272
R7634 commonsourceibias.n578 commonsourceibias.n577 48.3272
R7635 commonsourceibias.n693 commonsourceibias.n692 48.3272
R7636 commonsourceibias.n682 commonsourceibias.n681 48.3272
R7637 commonsourceibias.n417 commonsourceibias.n388 47.3584
R7638 commonsourceibias.n457 commonsourceibias.n456 47.3584
R7639 commonsourceibias.n341 commonsourceibias.n340 47.3584
R7640 commonsourceibias.n301 commonsourceibias.n272 47.3584
R7641 commonsourceibias.n104 commonsourceibias.n103 47.3584
R7642 commonsourceibias.n64 commonsourceibias.n35 47.3584
R7643 commonsourceibias.n226 commonsourceibias.n225 47.3584
R7644 commonsourceibias.n186 commonsourceibias.n157 47.3584
R7645 commonsourceibias.n896 commonsourceibias.n867 47.3584
R7646 commonsourceibias.n939 commonsourceibias.n938 47.3584
R7647 commonsourceibias.n780 commonsourceibias.n751 47.3584
R7648 commonsourceibias.n823 commonsourceibias.n822 47.3584
R7649 commonsourceibias.n550 commonsourceibias.n521 47.3584
R7650 commonsourceibias.n593 commonsourceibias.n592 47.3584
R7651 commonsourceibias.n708 commonsourceibias.n707 47.3584
R7652 commonsourceibias.n666 commonsourceibias.n637 47.3584
R7653 commonsourceibias.n403 commonsourceibias.n393 46.3896
R7654 commonsourceibias.n471 commonsourceibias.n470 46.3896
R7655 commonsourceibias.n355 commonsourceibias.n354 46.3896
R7656 commonsourceibias.n287 commonsourceibias.n277 46.3896
R7657 commonsourceibias.n118 commonsourceibias.n117 46.3896
R7658 commonsourceibias.n50 commonsourceibias.n40 46.3896
R7659 commonsourceibias.n240 commonsourceibias.n239 46.3896
R7660 commonsourceibias.n172 commonsourceibias.n162 46.3896
R7661 commonsourceibias.n881 commonsourceibias.n871 46.3896
R7662 commonsourceibias.n954 commonsourceibias.n953 46.3896
R7663 commonsourceibias.n765 commonsourceibias.n755 46.3896
R7664 commonsourceibias.n838 commonsourceibias.n837 46.3896
R7665 commonsourceibias.n535 commonsourceibias.n525 46.3896
R7666 commonsourceibias.n608 commonsourceibias.n607 46.3896
R7667 commonsourceibias.n723 commonsourceibias.n722 46.3896
R7668 commonsourceibias.n651 commonsourceibias.n641 46.3896
R7669 commonsourceibias.n398 commonsourceibias.n397 44.7059
R7670 commonsourceibias.n876 commonsourceibias.n875 44.7059
R7671 commonsourceibias.n760 commonsourceibias.n759 44.7059
R7672 commonsourceibias.n530 commonsourceibias.n529 44.7059
R7673 commonsourceibias.n646 commonsourceibias.n645 44.7059
R7674 commonsourceibias.n282 commonsourceibias.n281 44.7059
R7675 commonsourceibias.n45 commonsourceibias.n44 44.7059
R7676 commonsourceibias.n167 commonsourceibias.n166 44.7059
R7677 commonsourceibias.n407 commonsourceibias.n393 34.7644
R7678 commonsourceibias.n470 commonsourceibias.n370 34.7644
R7679 commonsourceibias.n354 commonsourceibias.n254 34.7644
R7680 commonsourceibias.n291 commonsourceibias.n277 34.7644
R7681 commonsourceibias.n117 commonsourceibias.n17 34.7644
R7682 commonsourceibias.n54 commonsourceibias.n40 34.7644
R7683 commonsourceibias.n239 commonsourceibias.n3 34.7644
R7684 commonsourceibias.n176 commonsourceibias.n162 34.7644
R7685 commonsourceibias.n885 commonsourceibias.n871 34.7644
R7686 commonsourceibias.n953 commonsourceibias.n853 34.7644
R7687 commonsourceibias.n769 commonsourceibias.n755 34.7644
R7688 commonsourceibias.n837 commonsourceibias.n737 34.7644
R7689 commonsourceibias.n539 commonsourceibias.n525 34.7644
R7690 commonsourceibias.n607 commonsourceibias.n507 34.7644
R7691 commonsourceibias.n722 commonsourceibias.n486 34.7644
R7692 commonsourceibias.n655 commonsourceibias.n641 34.7644
R7693 commonsourceibias.n421 commonsourceibias.n388 33.7956
R7694 commonsourceibias.n456 commonsourceibias.n375 33.7956
R7695 commonsourceibias.n340 commonsourceibias.n259 33.7956
R7696 commonsourceibias.n305 commonsourceibias.n272 33.7956
R7697 commonsourceibias.n103 commonsourceibias.n22 33.7956
R7698 commonsourceibias.n68 commonsourceibias.n35 33.7956
R7699 commonsourceibias.n225 commonsourceibias.n8 33.7956
R7700 commonsourceibias.n190 commonsourceibias.n157 33.7956
R7701 commonsourceibias.n900 commonsourceibias.n867 33.7956
R7702 commonsourceibias.n938 commonsourceibias.n857 33.7956
R7703 commonsourceibias.n784 commonsourceibias.n751 33.7956
R7704 commonsourceibias.n822 commonsourceibias.n741 33.7956
R7705 commonsourceibias.n554 commonsourceibias.n521 33.7956
R7706 commonsourceibias.n592 commonsourceibias.n511 33.7956
R7707 commonsourceibias.n707 commonsourceibias.n490 33.7956
R7708 commonsourceibias.n670 commonsourceibias.n637 33.7956
R7709 commonsourceibias.n435 commonsourceibias.n383 32.8269
R7710 commonsourceibias.n442 commonsourceibias.n380 32.8269
R7711 commonsourceibias.n326 commonsourceibias.n264 32.8269
R7712 commonsourceibias.n319 commonsourceibias.n267 32.8269
R7713 commonsourceibias.n89 commonsourceibias.n27 32.8269
R7714 commonsourceibias.n82 commonsourceibias.n30 32.8269
R7715 commonsourceibias.n211 commonsourceibias.n13 32.8269
R7716 commonsourceibias.n203 commonsourceibias.n202 32.8269
R7717 commonsourceibias.n915 commonsourceibias.n863 32.8269
R7718 commonsourceibias.n923 commonsourceibias.n861 32.8269
R7719 commonsourceibias.n799 commonsourceibias.n747 32.8269
R7720 commonsourceibias.n807 commonsourceibias.n745 32.8269
R7721 commonsourceibias.n569 commonsourceibias.n517 32.8269
R7722 commonsourceibias.n577 commonsourceibias.n515 32.8269
R7723 commonsourceibias.n692 commonsourceibias.n494 32.8269
R7724 commonsourceibias.n683 commonsourceibias.n682 32.8269
R7725 commonsourceibias.n428 commonsourceibias.n385 31.8581
R7726 commonsourceibias.n449 commonsourceibias.n378 31.8581
R7727 commonsourceibias.n333 commonsourceibias.n262 31.8581
R7728 commonsourceibias.n312 commonsourceibias.n269 31.8581
R7729 commonsourceibias.n96 commonsourceibias.n25 31.8581
R7730 commonsourceibias.n75 commonsourceibias.n32 31.8581
R7731 commonsourceibias.n218 commonsourceibias.n11 31.8581
R7732 commonsourceibias.n197 commonsourceibias.n196 31.8581
R7733 commonsourceibias.n908 commonsourceibias.n865 31.8581
R7734 commonsourceibias.n930 commonsourceibias.n859 31.8581
R7735 commonsourceibias.n792 commonsourceibias.n749 31.8581
R7736 commonsourceibias.n814 commonsourceibias.n743 31.8581
R7737 commonsourceibias.n562 commonsourceibias.n519 31.8581
R7738 commonsourceibias.n584 commonsourceibias.n513 31.8581
R7739 commonsourceibias.n699 commonsourceibias.n492 31.8581
R7740 commonsourceibias.n677 commonsourceibias.n676 31.8581
R7741 commonsourceibias.n414 commonsourceibias.n390 30.8893
R7742 commonsourceibias.n463 commonsourceibias.n373 30.8893
R7743 commonsourceibias.n347 commonsourceibias.n257 30.8893
R7744 commonsourceibias.n298 commonsourceibias.n274 30.8893
R7745 commonsourceibias.n110 commonsourceibias.n20 30.8893
R7746 commonsourceibias.n61 commonsourceibias.n37 30.8893
R7747 commonsourceibias.n232 commonsourceibias.n6 30.8893
R7748 commonsourceibias.n183 commonsourceibias.n159 30.8893
R7749 commonsourceibias.n893 commonsourceibias.n869 30.8893
R7750 commonsourceibias.n945 commonsourceibias.n855 30.8893
R7751 commonsourceibias.n777 commonsourceibias.n753 30.8893
R7752 commonsourceibias.n829 commonsourceibias.n739 30.8893
R7753 commonsourceibias.n547 commonsourceibias.n523 30.8893
R7754 commonsourceibias.n599 commonsourceibias.n509 30.8893
R7755 commonsourceibias.n714 commonsourceibias.n488 30.8893
R7756 commonsourceibias.n663 commonsourceibias.n639 30.8893
R7757 commonsourceibias.n400 commonsourceibias.n395 29.9206
R7758 commonsourceibias.n477 commonsourceibias.n368 29.9206
R7759 commonsourceibias.n361 commonsourceibias.n252 29.9206
R7760 commonsourceibias.n284 commonsourceibias.n279 29.9206
R7761 commonsourceibias.n124 commonsourceibias.n15 29.9206
R7762 commonsourceibias.n47 commonsourceibias.n42 29.9206
R7763 commonsourceibias.n246 commonsourceibias.n1 29.9206
R7764 commonsourceibias.n169 commonsourceibias.n164 29.9206
R7765 commonsourceibias.n878 commonsourceibias.n873 29.9206
R7766 commonsourceibias.n960 commonsourceibias.n851 29.9206
R7767 commonsourceibias.n762 commonsourceibias.n757 29.9206
R7768 commonsourceibias.n844 commonsourceibias.n735 29.9206
R7769 commonsourceibias.n532 commonsourceibias.n527 29.9206
R7770 commonsourceibias.n614 commonsourceibias.n505 29.9206
R7771 commonsourceibias.n729 commonsourceibias.n484 29.9206
R7772 commonsourceibias.n648 commonsourceibias.n643 29.9206
R7773 commonsourceibias.n479 commonsourceibias.n478 21.8872
R7774 commonsourceibias.n363 commonsourceibias.n362 21.8872
R7775 commonsourceibias.n126 commonsourceibias.n125 21.8872
R7776 commonsourceibias.n248 commonsourceibias.n247 21.8872
R7777 commonsourceibias.n962 commonsourceibias.n961 21.8872
R7778 commonsourceibias.n846 commonsourceibias.n845 21.8872
R7779 commonsourceibias.n616 commonsourceibias.n615 21.8872
R7780 commonsourceibias.n731 commonsourceibias.n730 21.8872
R7781 commonsourceibias.n410 commonsourceibias.n392 21.3954
R7782 commonsourceibias.n465 commonsourceibias.n464 21.3954
R7783 commonsourceibias.n349 commonsourceibias.n348 21.3954
R7784 commonsourceibias.n294 commonsourceibias.n276 21.3954
R7785 commonsourceibias.n112 commonsourceibias.n111 21.3954
R7786 commonsourceibias.n57 commonsourceibias.n39 21.3954
R7787 commonsourceibias.n234 commonsourceibias.n233 21.3954
R7788 commonsourceibias.n179 commonsourceibias.n161 21.3954
R7789 commonsourceibias.n889 commonsourceibias.n888 21.3954
R7790 commonsourceibias.n947 commonsourceibias.n946 21.3954
R7791 commonsourceibias.n773 commonsourceibias.n772 21.3954
R7792 commonsourceibias.n831 commonsourceibias.n830 21.3954
R7793 commonsourceibias.n543 commonsourceibias.n542 21.3954
R7794 commonsourceibias.n601 commonsourceibias.n600 21.3954
R7795 commonsourceibias.n716 commonsourceibias.n715 21.3954
R7796 commonsourceibias.n659 commonsourceibias.n658 21.3954
R7797 commonsourceibias.n424 commonsourceibias.n387 20.9036
R7798 commonsourceibias.n451 commonsourceibias.n450 20.9036
R7799 commonsourceibias.n335 commonsourceibias.n334 20.9036
R7800 commonsourceibias.n308 commonsourceibias.n271 20.9036
R7801 commonsourceibias.n98 commonsourceibias.n97 20.9036
R7802 commonsourceibias.n71 commonsourceibias.n34 20.9036
R7803 commonsourceibias.n220 commonsourceibias.n219 20.9036
R7804 commonsourceibias.n193 commonsourceibias.n155 20.9036
R7805 commonsourceibias.n904 commonsourceibias.n903 20.9036
R7806 commonsourceibias.n932 commonsourceibias.n931 20.9036
R7807 commonsourceibias.n788 commonsourceibias.n787 20.9036
R7808 commonsourceibias.n816 commonsourceibias.n815 20.9036
R7809 commonsourceibias.n558 commonsourceibias.n557 20.9036
R7810 commonsourceibias.n586 commonsourceibias.n585 20.9036
R7811 commonsourceibias.n701 commonsourceibias.n700 20.9036
R7812 commonsourceibias.n673 commonsourceibias.n635 20.9036
R7813 commonsourceibias.n437 commonsourceibias.n436 20.4117
R7814 commonsourceibias.n438 commonsourceibias.n382 20.4117
R7815 commonsourceibias.n322 commonsourceibias.n266 20.4117
R7816 commonsourceibias.n321 commonsourceibias.n320 20.4117
R7817 commonsourceibias.n85 commonsourceibias.n29 20.4117
R7818 commonsourceibias.n84 commonsourceibias.n83 20.4117
R7819 commonsourceibias.n207 commonsourceibias.n150 20.4117
R7820 commonsourceibias.n206 commonsourceibias.n151 20.4117
R7821 commonsourceibias.n917 commonsourceibias.n916 20.4117
R7822 commonsourceibias.n919 commonsourceibias.n918 20.4117
R7823 commonsourceibias.n801 commonsourceibias.n800 20.4117
R7824 commonsourceibias.n803 commonsourceibias.n802 20.4117
R7825 commonsourceibias.n571 commonsourceibias.n570 20.4117
R7826 commonsourceibias.n573 commonsourceibias.n572 20.4117
R7827 commonsourceibias.n688 commonsourceibias.n687 20.4117
R7828 commonsourceibias.n686 commonsourceibias.n631 20.4117
R7829 commonsourceibias.n423 commonsourceibias.n422 19.9199
R7830 commonsourceibias.n452 commonsourceibias.n377 19.9199
R7831 commonsourceibias.n336 commonsourceibias.n261 19.9199
R7832 commonsourceibias.n307 commonsourceibias.n306 19.9199
R7833 commonsourceibias.n99 commonsourceibias.n24 19.9199
R7834 commonsourceibias.n70 commonsourceibias.n69 19.9199
R7835 commonsourceibias.n221 commonsourceibias.n10 19.9199
R7836 commonsourceibias.n192 commonsourceibias.n191 19.9199
R7837 commonsourceibias.n902 commonsourceibias.n901 19.9199
R7838 commonsourceibias.n934 commonsourceibias.n933 19.9199
R7839 commonsourceibias.n786 commonsourceibias.n785 19.9199
R7840 commonsourceibias.n818 commonsourceibias.n817 19.9199
R7841 commonsourceibias.n556 commonsourceibias.n555 19.9199
R7842 commonsourceibias.n588 commonsourceibias.n587 19.9199
R7843 commonsourceibias.n703 commonsourceibias.n702 19.9199
R7844 commonsourceibias.n672 commonsourceibias.n671 19.9199
R7845 commonsourceibias.n409 commonsourceibias.n408 19.4281
R7846 commonsourceibias.n466 commonsourceibias.n372 19.4281
R7847 commonsourceibias.n350 commonsourceibias.n256 19.4281
R7848 commonsourceibias.n293 commonsourceibias.n292 19.4281
R7849 commonsourceibias.n113 commonsourceibias.n19 19.4281
R7850 commonsourceibias.n56 commonsourceibias.n55 19.4281
R7851 commonsourceibias.n235 commonsourceibias.n5 19.4281
R7852 commonsourceibias.n178 commonsourceibias.n177 19.4281
R7853 commonsourceibias.n887 commonsourceibias.n886 19.4281
R7854 commonsourceibias.n949 commonsourceibias.n948 19.4281
R7855 commonsourceibias.n771 commonsourceibias.n770 19.4281
R7856 commonsourceibias.n833 commonsourceibias.n832 19.4281
R7857 commonsourceibias.n541 commonsourceibias.n540 19.4281
R7858 commonsourceibias.n603 commonsourceibias.n602 19.4281
R7859 commonsourceibias.n718 commonsourceibias.n717 19.4281
R7860 commonsourceibias.n657 commonsourceibias.n656 19.4281
R7861 commonsourceibias.n402 commonsourceibias.n401 13.526
R7862 commonsourceibias.n473 commonsourceibias.n472 13.526
R7863 commonsourceibias.n357 commonsourceibias.n356 13.526
R7864 commonsourceibias.n286 commonsourceibias.n285 13.526
R7865 commonsourceibias.n120 commonsourceibias.n119 13.526
R7866 commonsourceibias.n49 commonsourceibias.n48 13.526
R7867 commonsourceibias.n242 commonsourceibias.n241 13.526
R7868 commonsourceibias.n171 commonsourceibias.n170 13.526
R7869 commonsourceibias.n880 commonsourceibias.n879 13.526
R7870 commonsourceibias.n956 commonsourceibias.n955 13.526
R7871 commonsourceibias.n764 commonsourceibias.n763 13.526
R7872 commonsourceibias.n840 commonsourceibias.n839 13.526
R7873 commonsourceibias.n534 commonsourceibias.n533 13.526
R7874 commonsourceibias.n610 commonsourceibias.n609 13.526
R7875 commonsourceibias.n725 commonsourceibias.n724 13.526
R7876 commonsourceibias.n650 commonsourceibias.n649 13.526
R7877 commonsourceibias.n130 commonsourceibias.n128 13.2322
R7878 commonsourceibias.n620 commonsourceibias.n618 13.2322
R7879 commonsourceibias.n416 commonsourceibias.n415 13.0342
R7880 commonsourceibias.n459 commonsourceibias.n458 13.0342
R7881 commonsourceibias.n343 commonsourceibias.n342 13.0342
R7882 commonsourceibias.n300 commonsourceibias.n299 13.0342
R7883 commonsourceibias.n106 commonsourceibias.n105 13.0342
R7884 commonsourceibias.n63 commonsourceibias.n62 13.0342
R7885 commonsourceibias.n228 commonsourceibias.n227 13.0342
R7886 commonsourceibias.n185 commonsourceibias.n184 13.0342
R7887 commonsourceibias.n895 commonsourceibias.n894 13.0342
R7888 commonsourceibias.n941 commonsourceibias.n940 13.0342
R7889 commonsourceibias.n779 commonsourceibias.n778 13.0342
R7890 commonsourceibias.n825 commonsourceibias.n824 13.0342
R7891 commonsourceibias.n549 commonsourceibias.n548 13.0342
R7892 commonsourceibias.n595 commonsourceibias.n594 13.0342
R7893 commonsourceibias.n710 commonsourceibias.n709 13.0342
R7894 commonsourceibias.n665 commonsourceibias.n664 13.0342
R7895 commonsourceibias.n430 commonsourceibias.n429 12.5423
R7896 commonsourceibias.n445 commonsourceibias.n444 12.5423
R7897 commonsourceibias.n329 commonsourceibias.n328 12.5423
R7898 commonsourceibias.n314 commonsourceibias.n313 12.5423
R7899 commonsourceibias.n92 commonsourceibias.n91 12.5423
R7900 commonsourceibias.n77 commonsourceibias.n76 12.5423
R7901 commonsourceibias.n214 commonsourceibias.n213 12.5423
R7902 commonsourceibias.n198 commonsourceibias.n153 12.5423
R7903 commonsourceibias.n910 commonsourceibias.n909 12.5423
R7904 commonsourceibias.n926 commonsourceibias.n925 12.5423
R7905 commonsourceibias.n794 commonsourceibias.n793 12.5423
R7906 commonsourceibias.n810 commonsourceibias.n809 12.5423
R7907 commonsourceibias.n564 commonsourceibias.n563 12.5423
R7908 commonsourceibias.n580 commonsourceibias.n579 12.5423
R7909 commonsourceibias.n695 commonsourceibias.n694 12.5423
R7910 commonsourceibias.n678 commonsourceibias.n633 12.5423
R7911 commonsourceibias.n431 commonsourceibias.n430 12.0505
R7912 commonsourceibias.n444 commonsourceibias.n443 12.0505
R7913 commonsourceibias.n328 commonsourceibias.n327 12.0505
R7914 commonsourceibias.n315 commonsourceibias.n314 12.0505
R7915 commonsourceibias.n91 commonsourceibias.n90 12.0505
R7916 commonsourceibias.n78 commonsourceibias.n77 12.0505
R7917 commonsourceibias.n213 commonsourceibias.n212 12.0505
R7918 commonsourceibias.n201 commonsourceibias.n153 12.0505
R7919 commonsourceibias.n911 commonsourceibias.n910 12.0505
R7920 commonsourceibias.n925 commonsourceibias.n924 12.0505
R7921 commonsourceibias.n795 commonsourceibias.n794 12.0505
R7922 commonsourceibias.n809 commonsourceibias.n808 12.0505
R7923 commonsourceibias.n565 commonsourceibias.n564 12.0505
R7924 commonsourceibias.n579 commonsourceibias.n578 12.0505
R7925 commonsourceibias.n694 commonsourceibias.n693 12.0505
R7926 commonsourceibias.n681 commonsourceibias.n633 12.0505
R7927 commonsourceibias.n417 commonsourceibias.n416 11.5587
R7928 commonsourceibias.n458 commonsourceibias.n457 11.5587
R7929 commonsourceibias.n342 commonsourceibias.n341 11.5587
R7930 commonsourceibias.n301 commonsourceibias.n300 11.5587
R7931 commonsourceibias.n105 commonsourceibias.n104 11.5587
R7932 commonsourceibias.n64 commonsourceibias.n63 11.5587
R7933 commonsourceibias.n227 commonsourceibias.n226 11.5587
R7934 commonsourceibias.n186 commonsourceibias.n185 11.5587
R7935 commonsourceibias.n896 commonsourceibias.n895 11.5587
R7936 commonsourceibias.n940 commonsourceibias.n939 11.5587
R7937 commonsourceibias.n780 commonsourceibias.n779 11.5587
R7938 commonsourceibias.n824 commonsourceibias.n823 11.5587
R7939 commonsourceibias.n550 commonsourceibias.n549 11.5587
R7940 commonsourceibias.n594 commonsourceibias.n593 11.5587
R7941 commonsourceibias.n709 commonsourceibias.n708 11.5587
R7942 commonsourceibias.n666 commonsourceibias.n665 11.5587
R7943 commonsourceibias.n403 commonsourceibias.n402 11.0668
R7944 commonsourceibias.n472 commonsourceibias.n471 11.0668
R7945 commonsourceibias.n356 commonsourceibias.n355 11.0668
R7946 commonsourceibias.n287 commonsourceibias.n286 11.0668
R7947 commonsourceibias.n119 commonsourceibias.n118 11.0668
R7948 commonsourceibias.n50 commonsourceibias.n49 11.0668
R7949 commonsourceibias.n241 commonsourceibias.n240 11.0668
R7950 commonsourceibias.n172 commonsourceibias.n171 11.0668
R7951 commonsourceibias.n881 commonsourceibias.n880 11.0668
R7952 commonsourceibias.n955 commonsourceibias.n954 11.0668
R7953 commonsourceibias.n765 commonsourceibias.n764 11.0668
R7954 commonsourceibias.n839 commonsourceibias.n838 11.0668
R7955 commonsourceibias.n535 commonsourceibias.n534 11.0668
R7956 commonsourceibias.n609 commonsourceibias.n608 11.0668
R7957 commonsourceibias.n724 commonsourceibias.n723 11.0668
R7958 commonsourceibias.n651 commonsourceibias.n650 11.0668
R7959 commonsourceibias.n966 commonsourceibias.n482 10.4122
R7960 commonsourceibias.n149 commonsourceibias.n148 9.50363
R7961 commonsourceibias.n630 commonsourceibias.n629 9.50363
R7962 commonsourceibias.n366 commonsourceibias.n250 8.76042
R7963 commonsourceibias.n849 commonsourceibias.n733 8.76042
R7964 commonsourceibias.n966 commonsourceibias.n965 8.46921
R7965 commonsourceibias.n408 commonsourceibias.n407 5.16479
R7966 commonsourceibias.n372 commonsourceibias.n370 5.16479
R7967 commonsourceibias.n256 commonsourceibias.n254 5.16479
R7968 commonsourceibias.n292 commonsourceibias.n291 5.16479
R7969 commonsourceibias.n19 commonsourceibias.n17 5.16479
R7970 commonsourceibias.n55 commonsourceibias.n54 5.16479
R7971 commonsourceibias.n5 commonsourceibias.n3 5.16479
R7972 commonsourceibias.n177 commonsourceibias.n176 5.16479
R7973 commonsourceibias.n886 commonsourceibias.n885 5.16479
R7974 commonsourceibias.n948 commonsourceibias.n853 5.16479
R7975 commonsourceibias.n770 commonsourceibias.n769 5.16479
R7976 commonsourceibias.n832 commonsourceibias.n737 5.16479
R7977 commonsourceibias.n540 commonsourceibias.n539 5.16479
R7978 commonsourceibias.n602 commonsourceibias.n507 5.16479
R7979 commonsourceibias.n717 commonsourceibias.n486 5.16479
R7980 commonsourceibias.n656 commonsourceibias.n655 5.16479
R7981 commonsourceibias.n482 commonsourceibias.n481 5.03125
R7982 commonsourceibias.n366 commonsourceibias.n365 5.03125
R7983 commonsourceibias.n965 commonsourceibias.n964 5.03125
R7984 commonsourceibias.n849 commonsourceibias.n848 5.03125
R7985 commonsourceibias.n422 commonsourceibias.n421 4.67295
R7986 commonsourceibias.n377 commonsourceibias.n375 4.67295
R7987 commonsourceibias.n261 commonsourceibias.n259 4.67295
R7988 commonsourceibias.n306 commonsourceibias.n305 4.67295
R7989 commonsourceibias.n24 commonsourceibias.n22 4.67295
R7990 commonsourceibias.n69 commonsourceibias.n68 4.67295
R7991 commonsourceibias.n10 commonsourceibias.n8 4.67295
R7992 commonsourceibias.n191 commonsourceibias.n190 4.67295
R7993 commonsourceibias.n901 commonsourceibias.n900 4.67295
R7994 commonsourceibias.n933 commonsourceibias.n857 4.67295
R7995 commonsourceibias.n785 commonsourceibias.n784 4.67295
R7996 commonsourceibias.n817 commonsourceibias.n741 4.67295
R7997 commonsourceibias.n555 commonsourceibias.n554 4.67295
R7998 commonsourceibias.n587 commonsourceibias.n511 4.67295
R7999 commonsourceibias.n702 commonsourceibias.n490 4.67295
R8000 commonsourceibias.n671 commonsourceibias.n670 4.67295
R8001 commonsourceibias commonsourceibias.n966 4.20978
R8002 commonsourceibias.n436 commonsourceibias.n435 4.18111
R8003 commonsourceibias.n382 commonsourceibias.n380 4.18111
R8004 commonsourceibias.n266 commonsourceibias.n264 4.18111
R8005 commonsourceibias.n320 commonsourceibias.n319 4.18111
R8006 commonsourceibias.n29 commonsourceibias.n27 4.18111
R8007 commonsourceibias.n83 commonsourceibias.n82 4.18111
R8008 commonsourceibias.n150 commonsourceibias.n13 4.18111
R8009 commonsourceibias.n203 commonsourceibias.n151 4.18111
R8010 commonsourceibias.n916 commonsourceibias.n915 4.18111
R8011 commonsourceibias.n918 commonsourceibias.n861 4.18111
R8012 commonsourceibias.n800 commonsourceibias.n799 4.18111
R8013 commonsourceibias.n802 commonsourceibias.n745 4.18111
R8014 commonsourceibias.n570 commonsourceibias.n569 4.18111
R8015 commonsourceibias.n572 commonsourceibias.n515 4.18111
R8016 commonsourceibias.n687 commonsourceibias.n494 4.18111
R8017 commonsourceibias.n683 commonsourceibias.n631 4.18111
R8018 commonsourceibias.n482 commonsourceibias.n366 3.72967
R8019 commonsourceibias.n965 commonsourceibias.n849 3.72967
R8020 commonsourceibias.n387 commonsourceibias.n385 3.68928
R8021 commonsourceibias.n450 commonsourceibias.n449 3.68928
R8022 commonsourceibias.n334 commonsourceibias.n333 3.68928
R8023 commonsourceibias.n271 commonsourceibias.n269 3.68928
R8024 commonsourceibias.n97 commonsourceibias.n96 3.68928
R8025 commonsourceibias.n34 commonsourceibias.n32 3.68928
R8026 commonsourceibias.n219 commonsourceibias.n218 3.68928
R8027 commonsourceibias.n196 commonsourceibias.n155 3.68928
R8028 commonsourceibias.n903 commonsourceibias.n865 3.68928
R8029 commonsourceibias.n931 commonsourceibias.n930 3.68928
R8030 commonsourceibias.n787 commonsourceibias.n749 3.68928
R8031 commonsourceibias.n815 commonsourceibias.n814 3.68928
R8032 commonsourceibias.n557 commonsourceibias.n519 3.68928
R8033 commonsourceibias.n585 commonsourceibias.n584 3.68928
R8034 commonsourceibias.n700 commonsourceibias.n699 3.68928
R8035 commonsourceibias.n676 commonsourceibias.n635 3.68928
R8036 commonsourceibias.n392 commonsourceibias.n390 3.19744
R8037 commonsourceibias.n464 commonsourceibias.n463 3.19744
R8038 commonsourceibias.n348 commonsourceibias.n347 3.19744
R8039 commonsourceibias.n276 commonsourceibias.n274 3.19744
R8040 commonsourceibias.n111 commonsourceibias.n110 3.19744
R8041 commonsourceibias.n39 commonsourceibias.n37 3.19744
R8042 commonsourceibias.n233 commonsourceibias.n232 3.19744
R8043 commonsourceibias.n161 commonsourceibias.n159 3.19744
R8044 commonsourceibias.n888 commonsourceibias.n869 3.19744
R8045 commonsourceibias.n946 commonsourceibias.n945 3.19744
R8046 commonsourceibias.n772 commonsourceibias.n753 3.19744
R8047 commonsourceibias.n830 commonsourceibias.n829 3.19744
R8048 commonsourceibias.n542 commonsourceibias.n523 3.19744
R8049 commonsourceibias.n600 commonsourceibias.n599 3.19744
R8050 commonsourceibias.n715 commonsourceibias.n714 3.19744
R8051 commonsourceibias.n658 commonsourceibias.n639 3.19744
R8052 commonsourceibias.n139 commonsourceibias.t67 2.82907
R8053 commonsourceibias.n139 commonsourceibias.t9 2.82907
R8054 commonsourceibias.n140 commonsourceibias.t3 2.82907
R8055 commonsourceibias.n140 commonsourceibias.t71 2.82907
R8056 commonsourceibias.n142 commonsourceibias.t47 2.82907
R8057 commonsourceibias.n142 commonsourceibias.t39 2.82907
R8058 commonsourceibias.n144 commonsourceibias.t37 2.82907
R8059 commonsourceibias.n144 commonsourceibias.t53 2.82907
R8060 commonsourceibias.n146 commonsourceibias.t65 2.82907
R8061 commonsourceibias.n146 commonsourceibias.t15 2.82907
R8062 commonsourceibias.n137 commonsourceibias.t77 2.82907
R8063 commonsourceibias.n137 commonsourceibias.t27 2.82907
R8064 commonsourceibias.n135 commonsourceibias.t13 2.82907
R8065 commonsourceibias.n135 commonsourceibias.t33 2.82907
R8066 commonsourceibias.n133 commonsourceibias.t35 2.82907
R8067 commonsourceibias.n133 commonsourceibias.t7 2.82907
R8068 commonsourceibias.n131 commonsourceibias.t1 2.82907
R8069 commonsourceibias.n131 commonsourceibias.t75 2.82907
R8070 commonsourceibias.n129 commonsourceibias.t51 2.82907
R8071 commonsourceibias.n129 commonsourceibias.t41 2.82907
R8072 commonsourceibias.n619 commonsourceibias.t29 2.82907
R8073 commonsourceibias.n619 commonsourceibias.t43 2.82907
R8074 commonsourceibias.n621 commonsourceibias.t19 2.82907
R8075 commonsourceibias.n621 commonsourceibias.t11 2.82907
R8076 commonsourceibias.n623 commonsourceibias.t45 2.82907
R8077 commonsourceibias.n623 commonsourceibias.t23 2.82907
R8078 commonsourceibias.n625 commonsourceibias.t21 2.82907
R8079 commonsourceibias.n625 commonsourceibias.t69 2.82907
R8080 commonsourceibias.n627 commonsourceibias.t63 2.82907
R8081 commonsourceibias.n627 commonsourceibias.t31 2.82907
R8082 commonsourceibias.n502 commonsourceibias.t5 2.82907
R8083 commonsourceibias.n502 commonsourceibias.t55 2.82907
R8084 commonsourceibias.n500 commonsourceibias.t73 2.82907
R8085 commonsourceibias.n500 commonsourceibias.t61 2.82907
R8086 commonsourceibias.n498 commonsourceibias.t59 2.82907
R8087 commonsourceibias.n498 commonsourceibias.t57 2.82907
R8088 commonsourceibias.n496 commonsourceibias.t25 2.82907
R8089 commonsourceibias.n496 commonsourceibias.t79 2.82907
R8090 commonsourceibias.n495 commonsourceibias.t17 2.82907
R8091 commonsourceibias.n495 commonsourceibias.t49 2.82907
R8092 commonsourceibias.n396 commonsourceibias.n395 2.7056
R8093 commonsourceibias.n478 commonsourceibias.n477 2.7056
R8094 commonsourceibias.n362 commonsourceibias.n361 2.7056
R8095 commonsourceibias.n280 commonsourceibias.n279 2.7056
R8096 commonsourceibias.n125 commonsourceibias.n124 2.7056
R8097 commonsourceibias.n43 commonsourceibias.n42 2.7056
R8098 commonsourceibias.n247 commonsourceibias.n246 2.7056
R8099 commonsourceibias.n165 commonsourceibias.n164 2.7056
R8100 commonsourceibias.n874 commonsourceibias.n873 2.7056
R8101 commonsourceibias.n961 commonsourceibias.n960 2.7056
R8102 commonsourceibias.n758 commonsourceibias.n757 2.7056
R8103 commonsourceibias.n845 commonsourceibias.n844 2.7056
R8104 commonsourceibias.n528 commonsourceibias.n527 2.7056
R8105 commonsourceibias.n615 commonsourceibias.n614 2.7056
R8106 commonsourceibias.n730 commonsourceibias.n729 2.7056
R8107 commonsourceibias.n644 commonsourceibias.n643 2.7056
R8108 commonsourceibias.n132 commonsourceibias.n130 0.573776
R8109 commonsourceibias.n134 commonsourceibias.n132 0.573776
R8110 commonsourceibias.n136 commonsourceibias.n134 0.573776
R8111 commonsourceibias.n138 commonsourceibias.n136 0.573776
R8112 commonsourceibias.n147 commonsourceibias.n145 0.573776
R8113 commonsourceibias.n145 commonsourceibias.n143 0.573776
R8114 commonsourceibias.n143 commonsourceibias.n141 0.573776
R8115 commonsourceibias.n499 commonsourceibias.n497 0.573776
R8116 commonsourceibias.n501 commonsourceibias.n499 0.573776
R8117 commonsourceibias.n503 commonsourceibias.n501 0.573776
R8118 commonsourceibias.n628 commonsourceibias.n626 0.573776
R8119 commonsourceibias.n626 commonsourceibias.n624 0.573776
R8120 commonsourceibias.n624 commonsourceibias.n622 0.573776
R8121 commonsourceibias.n622 commonsourceibias.n620 0.573776
R8122 commonsourceibias.n148 commonsourceibias.n138 0.287138
R8123 commonsourceibias.n148 commonsourceibias.n147 0.287138
R8124 commonsourceibias.n629 commonsourceibias.n503 0.287138
R8125 commonsourceibias.n629 commonsourceibias.n628 0.287138
R8126 commonsourceibias.n481 commonsourceibias.n367 0.285035
R8127 commonsourceibias.n365 commonsourceibias.n251 0.285035
R8128 commonsourceibias.n128 commonsourceibias.n14 0.285035
R8129 commonsourceibias.n250 commonsourceibias.n0 0.285035
R8130 commonsourceibias.n964 commonsourceibias.n850 0.285035
R8131 commonsourceibias.n848 commonsourceibias.n734 0.285035
R8132 commonsourceibias.n618 commonsourceibias.n504 0.285035
R8133 commonsourceibias.n733 commonsourceibias.n483 0.285035
R8134 commonsourceibias.n476 commonsourceibias.n367 0.189894
R8135 commonsourceibias.n476 commonsourceibias.n475 0.189894
R8136 commonsourceibias.n475 commonsourceibias.n474 0.189894
R8137 commonsourceibias.n474 commonsourceibias.n369 0.189894
R8138 commonsourceibias.n469 commonsourceibias.n369 0.189894
R8139 commonsourceibias.n469 commonsourceibias.n468 0.189894
R8140 commonsourceibias.n468 commonsourceibias.n467 0.189894
R8141 commonsourceibias.n467 commonsourceibias.n371 0.189894
R8142 commonsourceibias.n462 commonsourceibias.n371 0.189894
R8143 commonsourceibias.n462 commonsourceibias.n461 0.189894
R8144 commonsourceibias.n461 commonsourceibias.n460 0.189894
R8145 commonsourceibias.n460 commonsourceibias.n374 0.189894
R8146 commonsourceibias.n455 commonsourceibias.n374 0.189894
R8147 commonsourceibias.n455 commonsourceibias.n454 0.189894
R8148 commonsourceibias.n454 commonsourceibias.n453 0.189894
R8149 commonsourceibias.n453 commonsourceibias.n376 0.189894
R8150 commonsourceibias.n448 commonsourceibias.n376 0.189894
R8151 commonsourceibias.n448 commonsourceibias.n447 0.189894
R8152 commonsourceibias.n447 commonsourceibias.n446 0.189894
R8153 commonsourceibias.n446 commonsourceibias.n379 0.189894
R8154 commonsourceibias.n441 commonsourceibias.n379 0.189894
R8155 commonsourceibias.n441 commonsourceibias.n440 0.189894
R8156 commonsourceibias.n440 commonsourceibias.n439 0.189894
R8157 commonsourceibias.n439 commonsourceibias.n381 0.189894
R8158 commonsourceibias.n434 commonsourceibias.n381 0.189894
R8159 commonsourceibias.n434 commonsourceibias.n433 0.189894
R8160 commonsourceibias.n433 commonsourceibias.n432 0.189894
R8161 commonsourceibias.n432 commonsourceibias.n384 0.189894
R8162 commonsourceibias.n427 commonsourceibias.n384 0.189894
R8163 commonsourceibias.n427 commonsourceibias.n426 0.189894
R8164 commonsourceibias.n426 commonsourceibias.n425 0.189894
R8165 commonsourceibias.n425 commonsourceibias.n386 0.189894
R8166 commonsourceibias.n420 commonsourceibias.n386 0.189894
R8167 commonsourceibias.n420 commonsourceibias.n419 0.189894
R8168 commonsourceibias.n419 commonsourceibias.n418 0.189894
R8169 commonsourceibias.n418 commonsourceibias.n389 0.189894
R8170 commonsourceibias.n413 commonsourceibias.n389 0.189894
R8171 commonsourceibias.n413 commonsourceibias.n412 0.189894
R8172 commonsourceibias.n412 commonsourceibias.n411 0.189894
R8173 commonsourceibias.n411 commonsourceibias.n391 0.189894
R8174 commonsourceibias.n406 commonsourceibias.n391 0.189894
R8175 commonsourceibias.n406 commonsourceibias.n405 0.189894
R8176 commonsourceibias.n405 commonsourceibias.n404 0.189894
R8177 commonsourceibias.n404 commonsourceibias.n394 0.189894
R8178 commonsourceibias.n399 commonsourceibias.n394 0.189894
R8179 commonsourceibias.n399 commonsourceibias.n398 0.189894
R8180 commonsourceibias.n360 commonsourceibias.n251 0.189894
R8181 commonsourceibias.n360 commonsourceibias.n359 0.189894
R8182 commonsourceibias.n359 commonsourceibias.n358 0.189894
R8183 commonsourceibias.n358 commonsourceibias.n253 0.189894
R8184 commonsourceibias.n353 commonsourceibias.n253 0.189894
R8185 commonsourceibias.n353 commonsourceibias.n352 0.189894
R8186 commonsourceibias.n352 commonsourceibias.n351 0.189894
R8187 commonsourceibias.n351 commonsourceibias.n255 0.189894
R8188 commonsourceibias.n346 commonsourceibias.n255 0.189894
R8189 commonsourceibias.n346 commonsourceibias.n345 0.189894
R8190 commonsourceibias.n345 commonsourceibias.n344 0.189894
R8191 commonsourceibias.n344 commonsourceibias.n258 0.189894
R8192 commonsourceibias.n339 commonsourceibias.n258 0.189894
R8193 commonsourceibias.n339 commonsourceibias.n338 0.189894
R8194 commonsourceibias.n338 commonsourceibias.n337 0.189894
R8195 commonsourceibias.n337 commonsourceibias.n260 0.189894
R8196 commonsourceibias.n332 commonsourceibias.n260 0.189894
R8197 commonsourceibias.n332 commonsourceibias.n331 0.189894
R8198 commonsourceibias.n331 commonsourceibias.n330 0.189894
R8199 commonsourceibias.n330 commonsourceibias.n263 0.189894
R8200 commonsourceibias.n325 commonsourceibias.n263 0.189894
R8201 commonsourceibias.n325 commonsourceibias.n324 0.189894
R8202 commonsourceibias.n324 commonsourceibias.n323 0.189894
R8203 commonsourceibias.n323 commonsourceibias.n265 0.189894
R8204 commonsourceibias.n318 commonsourceibias.n265 0.189894
R8205 commonsourceibias.n318 commonsourceibias.n317 0.189894
R8206 commonsourceibias.n317 commonsourceibias.n316 0.189894
R8207 commonsourceibias.n316 commonsourceibias.n268 0.189894
R8208 commonsourceibias.n311 commonsourceibias.n268 0.189894
R8209 commonsourceibias.n311 commonsourceibias.n310 0.189894
R8210 commonsourceibias.n310 commonsourceibias.n309 0.189894
R8211 commonsourceibias.n309 commonsourceibias.n270 0.189894
R8212 commonsourceibias.n304 commonsourceibias.n270 0.189894
R8213 commonsourceibias.n304 commonsourceibias.n303 0.189894
R8214 commonsourceibias.n303 commonsourceibias.n302 0.189894
R8215 commonsourceibias.n302 commonsourceibias.n273 0.189894
R8216 commonsourceibias.n297 commonsourceibias.n273 0.189894
R8217 commonsourceibias.n297 commonsourceibias.n296 0.189894
R8218 commonsourceibias.n296 commonsourceibias.n295 0.189894
R8219 commonsourceibias.n295 commonsourceibias.n275 0.189894
R8220 commonsourceibias.n290 commonsourceibias.n275 0.189894
R8221 commonsourceibias.n290 commonsourceibias.n289 0.189894
R8222 commonsourceibias.n289 commonsourceibias.n288 0.189894
R8223 commonsourceibias.n288 commonsourceibias.n278 0.189894
R8224 commonsourceibias.n283 commonsourceibias.n278 0.189894
R8225 commonsourceibias.n283 commonsourceibias.n282 0.189894
R8226 commonsourceibias.n123 commonsourceibias.n14 0.189894
R8227 commonsourceibias.n123 commonsourceibias.n122 0.189894
R8228 commonsourceibias.n122 commonsourceibias.n121 0.189894
R8229 commonsourceibias.n121 commonsourceibias.n16 0.189894
R8230 commonsourceibias.n116 commonsourceibias.n16 0.189894
R8231 commonsourceibias.n116 commonsourceibias.n115 0.189894
R8232 commonsourceibias.n115 commonsourceibias.n114 0.189894
R8233 commonsourceibias.n114 commonsourceibias.n18 0.189894
R8234 commonsourceibias.n109 commonsourceibias.n18 0.189894
R8235 commonsourceibias.n109 commonsourceibias.n108 0.189894
R8236 commonsourceibias.n108 commonsourceibias.n107 0.189894
R8237 commonsourceibias.n107 commonsourceibias.n21 0.189894
R8238 commonsourceibias.n102 commonsourceibias.n21 0.189894
R8239 commonsourceibias.n102 commonsourceibias.n101 0.189894
R8240 commonsourceibias.n101 commonsourceibias.n100 0.189894
R8241 commonsourceibias.n100 commonsourceibias.n23 0.189894
R8242 commonsourceibias.n95 commonsourceibias.n23 0.189894
R8243 commonsourceibias.n95 commonsourceibias.n94 0.189894
R8244 commonsourceibias.n94 commonsourceibias.n93 0.189894
R8245 commonsourceibias.n93 commonsourceibias.n26 0.189894
R8246 commonsourceibias.n88 commonsourceibias.n26 0.189894
R8247 commonsourceibias.n88 commonsourceibias.n87 0.189894
R8248 commonsourceibias.n87 commonsourceibias.n86 0.189894
R8249 commonsourceibias.n86 commonsourceibias.n28 0.189894
R8250 commonsourceibias.n81 commonsourceibias.n28 0.189894
R8251 commonsourceibias.n81 commonsourceibias.n80 0.189894
R8252 commonsourceibias.n80 commonsourceibias.n79 0.189894
R8253 commonsourceibias.n79 commonsourceibias.n31 0.189894
R8254 commonsourceibias.n74 commonsourceibias.n31 0.189894
R8255 commonsourceibias.n74 commonsourceibias.n73 0.189894
R8256 commonsourceibias.n73 commonsourceibias.n72 0.189894
R8257 commonsourceibias.n72 commonsourceibias.n33 0.189894
R8258 commonsourceibias.n67 commonsourceibias.n33 0.189894
R8259 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8260 commonsourceibias.n66 commonsourceibias.n65 0.189894
R8261 commonsourceibias.n65 commonsourceibias.n36 0.189894
R8262 commonsourceibias.n60 commonsourceibias.n36 0.189894
R8263 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8264 commonsourceibias.n59 commonsourceibias.n58 0.189894
R8265 commonsourceibias.n58 commonsourceibias.n38 0.189894
R8266 commonsourceibias.n53 commonsourceibias.n38 0.189894
R8267 commonsourceibias.n53 commonsourceibias.n52 0.189894
R8268 commonsourceibias.n52 commonsourceibias.n51 0.189894
R8269 commonsourceibias.n51 commonsourceibias.n41 0.189894
R8270 commonsourceibias.n46 commonsourceibias.n41 0.189894
R8271 commonsourceibias.n46 commonsourceibias.n45 0.189894
R8272 commonsourceibias.n205 commonsourceibias.n204 0.189894
R8273 commonsourceibias.n204 commonsourceibias.n152 0.189894
R8274 commonsourceibias.n200 commonsourceibias.n152 0.189894
R8275 commonsourceibias.n200 commonsourceibias.n199 0.189894
R8276 commonsourceibias.n199 commonsourceibias.n154 0.189894
R8277 commonsourceibias.n195 commonsourceibias.n154 0.189894
R8278 commonsourceibias.n195 commonsourceibias.n194 0.189894
R8279 commonsourceibias.n194 commonsourceibias.n156 0.189894
R8280 commonsourceibias.n189 commonsourceibias.n156 0.189894
R8281 commonsourceibias.n189 commonsourceibias.n188 0.189894
R8282 commonsourceibias.n188 commonsourceibias.n187 0.189894
R8283 commonsourceibias.n187 commonsourceibias.n158 0.189894
R8284 commonsourceibias.n182 commonsourceibias.n158 0.189894
R8285 commonsourceibias.n182 commonsourceibias.n181 0.189894
R8286 commonsourceibias.n181 commonsourceibias.n180 0.189894
R8287 commonsourceibias.n180 commonsourceibias.n160 0.189894
R8288 commonsourceibias.n175 commonsourceibias.n160 0.189894
R8289 commonsourceibias.n175 commonsourceibias.n174 0.189894
R8290 commonsourceibias.n174 commonsourceibias.n173 0.189894
R8291 commonsourceibias.n173 commonsourceibias.n163 0.189894
R8292 commonsourceibias.n168 commonsourceibias.n163 0.189894
R8293 commonsourceibias.n168 commonsourceibias.n167 0.189894
R8294 commonsourceibias.n245 commonsourceibias.n0 0.189894
R8295 commonsourceibias.n245 commonsourceibias.n244 0.189894
R8296 commonsourceibias.n244 commonsourceibias.n243 0.189894
R8297 commonsourceibias.n243 commonsourceibias.n2 0.189894
R8298 commonsourceibias.n238 commonsourceibias.n2 0.189894
R8299 commonsourceibias.n238 commonsourceibias.n237 0.189894
R8300 commonsourceibias.n237 commonsourceibias.n236 0.189894
R8301 commonsourceibias.n236 commonsourceibias.n4 0.189894
R8302 commonsourceibias.n231 commonsourceibias.n4 0.189894
R8303 commonsourceibias.n231 commonsourceibias.n230 0.189894
R8304 commonsourceibias.n230 commonsourceibias.n229 0.189894
R8305 commonsourceibias.n229 commonsourceibias.n7 0.189894
R8306 commonsourceibias.n224 commonsourceibias.n7 0.189894
R8307 commonsourceibias.n224 commonsourceibias.n223 0.189894
R8308 commonsourceibias.n223 commonsourceibias.n222 0.189894
R8309 commonsourceibias.n222 commonsourceibias.n9 0.189894
R8310 commonsourceibias.n217 commonsourceibias.n9 0.189894
R8311 commonsourceibias.n217 commonsourceibias.n216 0.189894
R8312 commonsourceibias.n216 commonsourceibias.n215 0.189894
R8313 commonsourceibias.n215 commonsourceibias.n12 0.189894
R8314 commonsourceibias.n210 commonsourceibias.n12 0.189894
R8315 commonsourceibias.n210 commonsourceibias.n209 0.189894
R8316 commonsourceibias.n209 commonsourceibias.n208 0.189894
R8317 commonsourceibias.n877 commonsourceibias.n876 0.189894
R8318 commonsourceibias.n877 commonsourceibias.n872 0.189894
R8319 commonsourceibias.n882 commonsourceibias.n872 0.189894
R8320 commonsourceibias.n883 commonsourceibias.n882 0.189894
R8321 commonsourceibias.n884 commonsourceibias.n883 0.189894
R8322 commonsourceibias.n884 commonsourceibias.n870 0.189894
R8323 commonsourceibias.n890 commonsourceibias.n870 0.189894
R8324 commonsourceibias.n891 commonsourceibias.n890 0.189894
R8325 commonsourceibias.n892 commonsourceibias.n891 0.189894
R8326 commonsourceibias.n892 commonsourceibias.n868 0.189894
R8327 commonsourceibias.n897 commonsourceibias.n868 0.189894
R8328 commonsourceibias.n898 commonsourceibias.n897 0.189894
R8329 commonsourceibias.n899 commonsourceibias.n898 0.189894
R8330 commonsourceibias.n899 commonsourceibias.n866 0.189894
R8331 commonsourceibias.n905 commonsourceibias.n866 0.189894
R8332 commonsourceibias.n906 commonsourceibias.n905 0.189894
R8333 commonsourceibias.n907 commonsourceibias.n906 0.189894
R8334 commonsourceibias.n907 commonsourceibias.n864 0.189894
R8335 commonsourceibias.n912 commonsourceibias.n864 0.189894
R8336 commonsourceibias.n913 commonsourceibias.n912 0.189894
R8337 commonsourceibias.n914 commonsourceibias.n913 0.189894
R8338 commonsourceibias.n914 commonsourceibias.n862 0.189894
R8339 commonsourceibias.n920 commonsourceibias.n862 0.189894
R8340 commonsourceibias.n921 commonsourceibias.n920 0.189894
R8341 commonsourceibias.n922 commonsourceibias.n921 0.189894
R8342 commonsourceibias.n922 commonsourceibias.n860 0.189894
R8343 commonsourceibias.n927 commonsourceibias.n860 0.189894
R8344 commonsourceibias.n928 commonsourceibias.n927 0.189894
R8345 commonsourceibias.n929 commonsourceibias.n928 0.189894
R8346 commonsourceibias.n929 commonsourceibias.n858 0.189894
R8347 commonsourceibias.n935 commonsourceibias.n858 0.189894
R8348 commonsourceibias.n936 commonsourceibias.n935 0.189894
R8349 commonsourceibias.n937 commonsourceibias.n936 0.189894
R8350 commonsourceibias.n937 commonsourceibias.n856 0.189894
R8351 commonsourceibias.n942 commonsourceibias.n856 0.189894
R8352 commonsourceibias.n943 commonsourceibias.n942 0.189894
R8353 commonsourceibias.n944 commonsourceibias.n943 0.189894
R8354 commonsourceibias.n944 commonsourceibias.n854 0.189894
R8355 commonsourceibias.n950 commonsourceibias.n854 0.189894
R8356 commonsourceibias.n951 commonsourceibias.n950 0.189894
R8357 commonsourceibias.n952 commonsourceibias.n951 0.189894
R8358 commonsourceibias.n952 commonsourceibias.n852 0.189894
R8359 commonsourceibias.n957 commonsourceibias.n852 0.189894
R8360 commonsourceibias.n958 commonsourceibias.n957 0.189894
R8361 commonsourceibias.n959 commonsourceibias.n958 0.189894
R8362 commonsourceibias.n959 commonsourceibias.n850 0.189894
R8363 commonsourceibias.n761 commonsourceibias.n760 0.189894
R8364 commonsourceibias.n761 commonsourceibias.n756 0.189894
R8365 commonsourceibias.n766 commonsourceibias.n756 0.189894
R8366 commonsourceibias.n767 commonsourceibias.n766 0.189894
R8367 commonsourceibias.n768 commonsourceibias.n767 0.189894
R8368 commonsourceibias.n768 commonsourceibias.n754 0.189894
R8369 commonsourceibias.n774 commonsourceibias.n754 0.189894
R8370 commonsourceibias.n775 commonsourceibias.n774 0.189894
R8371 commonsourceibias.n776 commonsourceibias.n775 0.189894
R8372 commonsourceibias.n776 commonsourceibias.n752 0.189894
R8373 commonsourceibias.n781 commonsourceibias.n752 0.189894
R8374 commonsourceibias.n782 commonsourceibias.n781 0.189894
R8375 commonsourceibias.n783 commonsourceibias.n782 0.189894
R8376 commonsourceibias.n783 commonsourceibias.n750 0.189894
R8377 commonsourceibias.n789 commonsourceibias.n750 0.189894
R8378 commonsourceibias.n790 commonsourceibias.n789 0.189894
R8379 commonsourceibias.n791 commonsourceibias.n790 0.189894
R8380 commonsourceibias.n791 commonsourceibias.n748 0.189894
R8381 commonsourceibias.n796 commonsourceibias.n748 0.189894
R8382 commonsourceibias.n797 commonsourceibias.n796 0.189894
R8383 commonsourceibias.n798 commonsourceibias.n797 0.189894
R8384 commonsourceibias.n798 commonsourceibias.n746 0.189894
R8385 commonsourceibias.n804 commonsourceibias.n746 0.189894
R8386 commonsourceibias.n805 commonsourceibias.n804 0.189894
R8387 commonsourceibias.n806 commonsourceibias.n805 0.189894
R8388 commonsourceibias.n806 commonsourceibias.n744 0.189894
R8389 commonsourceibias.n811 commonsourceibias.n744 0.189894
R8390 commonsourceibias.n812 commonsourceibias.n811 0.189894
R8391 commonsourceibias.n813 commonsourceibias.n812 0.189894
R8392 commonsourceibias.n813 commonsourceibias.n742 0.189894
R8393 commonsourceibias.n819 commonsourceibias.n742 0.189894
R8394 commonsourceibias.n820 commonsourceibias.n819 0.189894
R8395 commonsourceibias.n821 commonsourceibias.n820 0.189894
R8396 commonsourceibias.n821 commonsourceibias.n740 0.189894
R8397 commonsourceibias.n826 commonsourceibias.n740 0.189894
R8398 commonsourceibias.n827 commonsourceibias.n826 0.189894
R8399 commonsourceibias.n828 commonsourceibias.n827 0.189894
R8400 commonsourceibias.n828 commonsourceibias.n738 0.189894
R8401 commonsourceibias.n834 commonsourceibias.n738 0.189894
R8402 commonsourceibias.n835 commonsourceibias.n834 0.189894
R8403 commonsourceibias.n836 commonsourceibias.n835 0.189894
R8404 commonsourceibias.n836 commonsourceibias.n736 0.189894
R8405 commonsourceibias.n841 commonsourceibias.n736 0.189894
R8406 commonsourceibias.n842 commonsourceibias.n841 0.189894
R8407 commonsourceibias.n843 commonsourceibias.n842 0.189894
R8408 commonsourceibias.n843 commonsourceibias.n734 0.189894
R8409 commonsourceibias.n531 commonsourceibias.n530 0.189894
R8410 commonsourceibias.n531 commonsourceibias.n526 0.189894
R8411 commonsourceibias.n536 commonsourceibias.n526 0.189894
R8412 commonsourceibias.n537 commonsourceibias.n536 0.189894
R8413 commonsourceibias.n538 commonsourceibias.n537 0.189894
R8414 commonsourceibias.n538 commonsourceibias.n524 0.189894
R8415 commonsourceibias.n544 commonsourceibias.n524 0.189894
R8416 commonsourceibias.n545 commonsourceibias.n544 0.189894
R8417 commonsourceibias.n546 commonsourceibias.n545 0.189894
R8418 commonsourceibias.n546 commonsourceibias.n522 0.189894
R8419 commonsourceibias.n551 commonsourceibias.n522 0.189894
R8420 commonsourceibias.n552 commonsourceibias.n551 0.189894
R8421 commonsourceibias.n553 commonsourceibias.n552 0.189894
R8422 commonsourceibias.n553 commonsourceibias.n520 0.189894
R8423 commonsourceibias.n559 commonsourceibias.n520 0.189894
R8424 commonsourceibias.n560 commonsourceibias.n559 0.189894
R8425 commonsourceibias.n561 commonsourceibias.n560 0.189894
R8426 commonsourceibias.n561 commonsourceibias.n518 0.189894
R8427 commonsourceibias.n566 commonsourceibias.n518 0.189894
R8428 commonsourceibias.n567 commonsourceibias.n566 0.189894
R8429 commonsourceibias.n568 commonsourceibias.n567 0.189894
R8430 commonsourceibias.n568 commonsourceibias.n516 0.189894
R8431 commonsourceibias.n574 commonsourceibias.n516 0.189894
R8432 commonsourceibias.n575 commonsourceibias.n574 0.189894
R8433 commonsourceibias.n576 commonsourceibias.n575 0.189894
R8434 commonsourceibias.n576 commonsourceibias.n514 0.189894
R8435 commonsourceibias.n581 commonsourceibias.n514 0.189894
R8436 commonsourceibias.n582 commonsourceibias.n581 0.189894
R8437 commonsourceibias.n583 commonsourceibias.n582 0.189894
R8438 commonsourceibias.n583 commonsourceibias.n512 0.189894
R8439 commonsourceibias.n589 commonsourceibias.n512 0.189894
R8440 commonsourceibias.n590 commonsourceibias.n589 0.189894
R8441 commonsourceibias.n591 commonsourceibias.n590 0.189894
R8442 commonsourceibias.n591 commonsourceibias.n510 0.189894
R8443 commonsourceibias.n596 commonsourceibias.n510 0.189894
R8444 commonsourceibias.n597 commonsourceibias.n596 0.189894
R8445 commonsourceibias.n598 commonsourceibias.n597 0.189894
R8446 commonsourceibias.n598 commonsourceibias.n508 0.189894
R8447 commonsourceibias.n604 commonsourceibias.n508 0.189894
R8448 commonsourceibias.n605 commonsourceibias.n604 0.189894
R8449 commonsourceibias.n606 commonsourceibias.n605 0.189894
R8450 commonsourceibias.n606 commonsourceibias.n506 0.189894
R8451 commonsourceibias.n611 commonsourceibias.n506 0.189894
R8452 commonsourceibias.n612 commonsourceibias.n611 0.189894
R8453 commonsourceibias.n613 commonsourceibias.n612 0.189894
R8454 commonsourceibias.n613 commonsourceibias.n504 0.189894
R8455 commonsourceibias.n647 commonsourceibias.n646 0.189894
R8456 commonsourceibias.n647 commonsourceibias.n642 0.189894
R8457 commonsourceibias.n652 commonsourceibias.n642 0.189894
R8458 commonsourceibias.n653 commonsourceibias.n652 0.189894
R8459 commonsourceibias.n654 commonsourceibias.n653 0.189894
R8460 commonsourceibias.n654 commonsourceibias.n640 0.189894
R8461 commonsourceibias.n660 commonsourceibias.n640 0.189894
R8462 commonsourceibias.n661 commonsourceibias.n660 0.189894
R8463 commonsourceibias.n662 commonsourceibias.n661 0.189894
R8464 commonsourceibias.n662 commonsourceibias.n638 0.189894
R8465 commonsourceibias.n667 commonsourceibias.n638 0.189894
R8466 commonsourceibias.n668 commonsourceibias.n667 0.189894
R8467 commonsourceibias.n669 commonsourceibias.n668 0.189894
R8468 commonsourceibias.n669 commonsourceibias.n636 0.189894
R8469 commonsourceibias.n674 commonsourceibias.n636 0.189894
R8470 commonsourceibias.n675 commonsourceibias.n674 0.189894
R8471 commonsourceibias.n675 commonsourceibias.n634 0.189894
R8472 commonsourceibias.n679 commonsourceibias.n634 0.189894
R8473 commonsourceibias.n680 commonsourceibias.n679 0.189894
R8474 commonsourceibias.n680 commonsourceibias.n632 0.189894
R8475 commonsourceibias.n684 commonsourceibias.n632 0.189894
R8476 commonsourceibias.n685 commonsourceibias.n684 0.189894
R8477 commonsourceibias.n690 commonsourceibias.n689 0.189894
R8478 commonsourceibias.n691 commonsourceibias.n690 0.189894
R8479 commonsourceibias.n691 commonsourceibias.n493 0.189894
R8480 commonsourceibias.n696 commonsourceibias.n493 0.189894
R8481 commonsourceibias.n697 commonsourceibias.n696 0.189894
R8482 commonsourceibias.n698 commonsourceibias.n697 0.189894
R8483 commonsourceibias.n698 commonsourceibias.n491 0.189894
R8484 commonsourceibias.n704 commonsourceibias.n491 0.189894
R8485 commonsourceibias.n705 commonsourceibias.n704 0.189894
R8486 commonsourceibias.n706 commonsourceibias.n705 0.189894
R8487 commonsourceibias.n706 commonsourceibias.n489 0.189894
R8488 commonsourceibias.n711 commonsourceibias.n489 0.189894
R8489 commonsourceibias.n712 commonsourceibias.n711 0.189894
R8490 commonsourceibias.n713 commonsourceibias.n712 0.189894
R8491 commonsourceibias.n713 commonsourceibias.n487 0.189894
R8492 commonsourceibias.n719 commonsourceibias.n487 0.189894
R8493 commonsourceibias.n720 commonsourceibias.n719 0.189894
R8494 commonsourceibias.n721 commonsourceibias.n720 0.189894
R8495 commonsourceibias.n721 commonsourceibias.n485 0.189894
R8496 commonsourceibias.n726 commonsourceibias.n485 0.189894
R8497 commonsourceibias.n727 commonsourceibias.n726 0.189894
R8498 commonsourceibias.n728 commonsourceibias.n727 0.189894
R8499 commonsourceibias.n728 commonsourceibias.n483 0.189894
R8500 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R8501 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R8502 commonsourceibias.n685 commonsourceibias.n630 0.0762576
R8503 commonsourceibias.n689 commonsourceibias.n630 0.0762576
R8504 gnd.n3813 gnd.n2413 766.379
R8505 gnd.n3816 gnd.n3815 766.379
R8506 gnd.n3055 gnd.n2958 766.379
R8507 gnd.n3051 gnd.n2956 766.379
R8508 gnd.n3904 gnd.n2435 756.769
R8509 gnd.n3807 gnd.n3806 756.769
R8510 gnd.n3148 gnd.n2865 756.769
R8511 gnd.n3146 gnd.n2868 756.769
R8512 gnd.n7644 gnd.n254 751.963
R8513 gnd.n7319 gnd.n252 751.963
R8514 gnd.n1154 gnd.n1030 751.963
R8515 gnd.n6012 gnd.n6011 751.963
R8516 gnd.n2080 gnd.n833 751.963
R8517 gnd.n4942 gnd.n842 751.963
R8518 gnd.n4213 gnd.n3908 751.963
R8519 gnd.n4261 gnd.n3910 751.963
R8520 gnd.n6813 gnd.n538 730.245
R8521 gnd.n5007 gnd.n862 711.122
R8522 gnd.n5914 gnd.n1168 711.122
R8523 gnd.n6384 gnd.n864 711.122
R8524 gnd.n6228 gnd.n995 711.122
R8525 gnd.n7646 gnd.n249 696.707
R8526 gnd.n7638 gnd.n251 696.707
R8527 gnd.n1153 gnd.n1152 696.707
R8528 gnd.n6213 gnd.n1072 696.707
R8529 gnd.n1782 gnd.n828 696.707
R8530 gnd.n6402 gnd.n6401 696.707
R8531 gnd.n4120 gnd.n3907 696.707
R8532 gnd.n4263 gnd.n2411 696.707
R8533 gnd.n6455 gnd.n751 689.5
R8534 gnd.n6812 gnd.n539 689.5
R8535 gnd.n7025 gnd.n7024 689.5
R8536 gnd.n4868 gnd.n4571 689.5
R8537 gnd.n4550 gnd.n756 585
R8538 gnd.n6452 gnd.n756 585
R8539 gnd.n4549 gnd.n4548 585
R8540 gnd.n4548 gnd.n4547 585
R8541 gnd.n2184 gnd.n2183 585
R8542 gnd.n2185 gnd.n2184 585
R8543 gnd.n4520 gnd.n2195 585
R8544 gnd.n4535 gnd.n2195 585
R8545 gnd.n4521 gnd.n2205 585
R8546 gnd.n2205 gnd.n2193 585
R8547 gnd.n4523 gnd.n4522 585
R8548 gnd.n4524 gnd.n4523 585
R8549 gnd.n2206 gnd.n2204 585
R8550 gnd.n4508 gnd.n2204 585
R8551 gnd.n4484 gnd.n4483 585
R8552 gnd.n4483 gnd.n2212 585
R8553 gnd.n4485 gnd.n2221 585
R8554 gnd.n4499 gnd.n2221 585
R8555 gnd.n4486 gnd.n2231 585
R8556 gnd.n2231 gnd.n2219 585
R8557 gnd.n4488 gnd.n4487 585
R8558 gnd.n4489 gnd.n4488 585
R8559 gnd.n2232 gnd.n2230 585
R8560 gnd.n4474 gnd.n2230 585
R8561 gnd.n4450 gnd.n4449 585
R8562 gnd.n4449 gnd.n2238 585
R8563 gnd.n4451 gnd.n2246 585
R8564 gnd.n4465 gnd.n2246 585
R8565 gnd.n4452 gnd.n2257 585
R8566 gnd.n2257 gnd.n2255 585
R8567 gnd.n4454 gnd.n4453 585
R8568 gnd.n4455 gnd.n4454 585
R8569 gnd.n2258 gnd.n2256 585
R8570 gnd.n4440 gnd.n2256 585
R8571 gnd.n4416 gnd.n4415 585
R8572 gnd.n4415 gnd.n2264 585
R8573 gnd.n4417 gnd.n2272 585
R8574 gnd.n4431 gnd.n2272 585
R8575 gnd.n4418 gnd.n2283 585
R8576 gnd.n2283 gnd.n2281 585
R8577 gnd.n4420 gnd.n4419 585
R8578 gnd.n4421 gnd.n4420 585
R8579 gnd.n2284 gnd.n2282 585
R8580 gnd.n4406 gnd.n2282 585
R8581 gnd.n4381 gnd.n4380 585
R8582 gnd.n4380 gnd.n2290 585
R8583 gnd.n4382 gnd.n2297 585
R8584 gnd.n4396 gnd.n2297 585
R8585 gnd.n4383 gnd.n2309 585
R8586 gnd.n2309 gnd.n2307 585
R8587 gnd.n4385 gnd.n4384 585
R8588 gnd.n4386 gnd.n4385 585
R8589 gnd.n2310 gnd.n2308 585
R8590 gnd.n2308 gnd.n2304 585
R8591 gnd.n4358 gnd.n2318 585
R8592 gnd.n4370 gnd.n2318 585
R8593 gnd.n4359 gnd.n2328 585
R8594 gnd.n2328 gnd.n2316 585
R8595 gnd.n4361 gnd.n4360 585
R8596 gnd.n4362 gnd.n4361 585
R8597 gnd.n2329 gnd.n2327 585
R8598 gnd.n2327 gnd.n2324 585
R8599 gnd.n4338 gnd.n2335 585
R8600 gnd.n4350 gnd.n2335 585
R8601 gnd.n4339 gnd.n2346 585
R8602 gnd.n2346 gnd.n2344 585
R8603 gnd.n4341 gnd.n4340 585
R8604 gnd.n4342 gnd.n4341 585
R8605 gnd.n2347 gnd.n2345 585
R8606 gnd.n2345 gnd.n2341 585
R8607 gnd.n4318 gnd.n2354 585
R8608 gnd.n4330 gnd.n2354 585
R8609 gnd.n4319 gnd.n2364 585
R8610 gnd.n2364 gnd.n2352 585
R8611 gnd.n4321 gnd.n4320 585
R8612 gnd.n4322 gnd.n4321 585
R8613 gnd.n2365 gnd.n2363 585
R8614 gnd.n2363 gnd.n2360 585
R8615 gnd.n4298 gnd.n2371 585
R8616 gnd.n4310 gnd.n2371 585
R8617 gnd.n4299 gnd.n2382 585
R8618 gnd.n2382 gnd.n2380 585
R8619 gnd.n4301 gnd.n4300 585
R8620 gnd.n4302 gnd.n4301 585
R8621 gnd.n2383 gnd.n2381 585
R8622 gnd.n2381 gnd.n2377 585
R8623 gnd.n4278 gnd.n2390 585
R8624 gnd.n4290 gnd.n2390 585
R8625 gnd.n4279 gnd.n2400 585
R8626 gnd.n2400 gnd.n2388 585
R8627 gnd.n4281 gnd.n4280 585
R8628 gnd.n4282 gnd.n4281 585
R8629 gnd.n2401 gnd.n2399 585
R8630 gnd.n2399 gnd.n2396 585
R8631 gnd.n4258 gnd.n2407 585
R8632 gnd.n4270 gnd.n2407 585
R8633 gnd.n4259 gnd.n3911 585
R8634 gnd.n3911 gnd.n3909 585
R8635 gnd.n4261 gnd.n4260 585
R8636 gnd.n4262 gnd.n4261 585
R8637 gnd.n4250 gnd.n3910 585
R8638 gnd.n4249 gnd.n4248 585
R8639 gnd.n4246 gnd.n4124 585
R8640 gnd.n4244 gnd.n4243 585
R8641 gnd.n4242 gnd.n4125 585
R8642 gnd.n4241 gnd.n4240 585
R8643 gnd.n4238 gnd.n4130 585
R8644 gnd.n4236 gnd.n4235 585
R8645 gnd.n4234 gnd.n4131 585
R8646 gnd.n4233 gnd.n4232 585
R8647 gnd.n4230 gnd.n4136 585
R8648 gnd.n4228 gnd.n4227 585
R8649 gnd.n4226 gnd.n4137 585
R8650 gnd.n4225 gnd.n4224 585
R8651 gnd.n4222 gnd.n4142 585
R8652 gnd.n4220 gnd.n4219 585
R8653 gnd.n4218 gnd.n4143 585
R8654 gnd.n4212 gnd.n4148 585
R8655 gnd.n4214 gnd.n4213 585
R8656 gnd.n4213 gnd.n3906 585
R8657 gnd.n2189 gnd.n755 585
R8658 gnd.n6452 gnd.n755 585
R8659 gnd.n4546 gnd.n4545 585
R8660 gnd.n4547 gnd.n4546 585
R8661 gnd.n2188 gnd.n2187 585
R8662 gnd.n2187 gnd.n2185 585
R8663 gnd.n4537 gnd.n4536 585
R8664 gnd.n4536 gnd.n4535 585
R8665 gnd.n2192 gnd.n2191 585
R8666 gnd.n2193 gnd.n2192 585
R8667 gnd.n2215 gnd.n2203 585
R8668 gnd.n4524 gnd.n2203 585
R8669 gnd.n4507 gnd.n4506 585
R8670 gnd.n4508 gnd.n4507 585
R8671 gnd.n2214 gnd.n2213 585
R8672 gnd.n2213 gnd.n2212 585
R8673 gnd.n4501 gnd.n4500 585
R8674 gnd.n4500 gnd.n4499 585
R8675 gnd.n2218 gnd.n2217 585
R8676 gnd.n2219 gnd.n2218 585
R8677 gnd.n2241 gnd.n2229 585
R8678 gnd.n4489 gnd.n2229 585
R8679 gnd.n4473 gnd.n4472 585
R8680 gnd.n4474 gnd.n4473 585
R8681 gnd.n2240 gnd.n2239 585
R8682 gnd.n2239 gnd.n2238 585
R8683 gnd.n4467 gnd.n4466 585
R8684 gnd.n4466 gnd.n4465 585
R8685 gnd.n2244 gnd.n2243 585
R8686 gnd.n2255 gnd.n2244 585
R8687 gnd.n2267 gnd.n2254 585
R8688 gnd.n4455 gnd.n2254 585
R8689 gnd.n4439 gnd.n4438 585
R8690 gnd.n4440 gnd.n4439 585
R8691 gnd.n2266 gnd.n2265 585
R8692 gnd.n2265 gnd.n2264 585
R8693 gnd.n4433 gnd.n4432 585
R8694 gnd.n4432 gnd.n4431 585
R8695 gnd.n2270 gnd.n2269 585
R8696 gnd.n2281 gnd.n2270 585
R8697 gnd.n4403 gnd.n2280 585
R8698 gnd.n4421 gnd.n2280 585
R8699 gnd.n4405 gnd.n4404 585
R8700 gnd.n4406 gnd.n4405 585
R8701 gnd.n2292 gnd.n2291 585
R8702 gnd.n2291 gnd.n2290 585
R8703 gnd.n4398 gnd.n4397 585
R8704 gnd.n4397 gnd.n4396 585
R8705 gnd.n2295 gnd.n2294 585
R8706 gnd.n2307 gnd.n2295 585
R8707 gnd.n4173 gnd.n2306 585
R8708 gnd.n4386 gnd.n2306 585
R8709 gnd.n4175 gnd.n4174 585
R8710 gnd.n4174 gnd.n2304 585
R8711 gnd.n4176 gnd.n2317 585
R8712 gnd.n4370 gnd.n2317 585
R8713 gnd.n4178 gnd.n4177 585
R8714 gnd.n4177 gnd.n2316 585
R8715 gnd.n4179 gnd.n2326 585
R8716 gnd.n4362 gnd.n2326 585
R8717 gnd.n4181 gnd.n4180 585
R8718 gnd.n4180 gnd.n2324 585
R8719 gnd.n4182 gnd.n2334 585
R8720 gnd.n4350 gnd.n2334 585
R8721 gnd.n4184 gnd.n4183 585
R8722 gnd.n4183 gnd.n2344 585
R8723 gnd.n4185 gnd.n2343 585
R8724 gnd.n4342 gnd.n2343 585
R8725 gnd.n4187 gnd.n4186 585
R8726 gnd.n4186 gnd.n2341 585
R8727 gnd.n4188 gnd.n2353 585
R8728 gnd.n4330 gnd.n2353 585
R8729 gnd.n4190 gnd.n4189 585
R8730 gnd.n4189 gnd.n2352 585
R8731 gnd.n4191 gnd.n2362 585
R8732 gnd.n4322 gnd.n2362 585
R8733 gnd.n4193 gnd.n4192 585
R8734 gnd.n4192 gnd.n2360 585
R8735 gnd.n4194 gnd.n2370 585
R8736 gnd.n4310 gnd.n2370 585
R8737 gnd.n4196 gnd.n4195 585
R8738 gnd.n4195 gnd.n2380 585
R8739 gnd.n4197 gnd.n2379 585
R8740 gnd.n4302 gnd.n2379 585
R8741 gnd.n4199 gnd.n4198 585
R8742 gnd.n4198 gnd.n2377 585
R8743 gnd.n4200 gnd.n2389 585
R8744 gnd.n4290 gnd.n2389 585
R8745 gnd.n4202 gnd.n4201 585
R8746 gnd.n4201 gnd.n2388 585
R8747 gnd.n4203 gnd.n2398 585
R8748 gnd.n4282 gnd.n2398 585
R8749 gnd.n4205 gnd.n4204 585
R8750 gnd.n4204 gnd.n2396 585
R8751 gnd.n4206 gnd.n2406 585
R8752 gnd.n4270 gnd.n2406 585
R8753 gnd.n4208 gnd.n4207 585
R8754 gnd.n4207 gnd.n3909 585
R8755 gnd.n4209 gnd.n3908 585
R8756 gnd.n4262 gnd.n3908 585
R8757 gnd.n3813 gnd.n3812 585
R8758 gnd.n3814 gnd.n3813 585
R8759 gnd.n2488 gnd.n2487 585
R8760 gnd.n2494 gnd.n2487 585
R8761 gnd.n3788 gnd.n2506 585
R8762 gnd.n2506 gnd.n2493 585
R8763 gnd.n3790 gnd.n3789 585
R8764 gnd.n3791 gnd.n3790 585
R8765 gnd.n2507 gnd.n2505 585
R8766 gnd.n2505 gnd.n2501 585
R8767 gnd.n3522 gnd.n3521 585
R8768 gnd.n3521 gnd.n3520 585
R8769 gnd.n2512 gnd.n2511 585
R8770 gnd.n3491 gnd.n2512 585
R8771 gnd.n3511 gnd.n3510 585
R8772 gnd.n3510 gnd.n3509 585
R8773 gnd.n2519 gnd.n2518 585
R8774 gnd.n3497 gnd.n2519 585
R8775 gnd.n3467 gnd.n2539 585
R8776 gnd.n2539 gnd.n2538 585
R8777 gnd.n3469 gnd.n3468 585
R8778 gnd.n3470 gnd.n3469 585
R8779 gnd.n2540 gnd.n2537 585
R8780 gnd.n2548 gnd.n2537 585
R8781 gnd.n3445 gnd.n2560 585
R8782 gnd.n2560 gnd.n2547 585
R8783 gnd.n3447 gnd.n3446 585
R8784 gnd.n3448 gnd.n3447 585
R8785 gnd.n2561 gnd.n2559 585
R8786 gnd.n2559 gnd.n2555 585
R8787 gnd.n3433 gnd.n3432 585
R8788 gnd.n3432 gnd.n3431 585
R8789 gnd.n2566 gnd.n2565 585
R8790 gnd.n2576 gnd.n2566 585
R8791 gnd.n3422 gnd.n3421 585
R8792 gnd.n3421 gnd.n3420 585
R8793 gnd.n2573 gnd.n2572 585
R8794 gnd.n3408 gnd.n2573 585
R8795 gnd.n3382 gnd.n2594 585
R8796 gnd.n2594 gnd.n2583 585
R8797 gnd.n3384 gnd.n3383 585
R8798 gnd.n3385 gnd.n3384 585
R8799 gnd.n2595 gnd.n2593 585
R8800 gnd.n2603 gnd.n2593 585
R8801 gnd.n3360 gnd.n2615 585
R8802 gnd.n2615 gnd.n2602 585
R8803 gnd.n3362 gnd.n3361 585
R8804 gnd.n3363 gnd.n3362 585
R8805 gnd.n2616 gnd.n2614 585
R8806 gnd.n2614 gnd.n2610 585
R8807 gnd.n3348 gnd.n3347 585
R8808 gnd.n3347 gnd.n3346 585
R8809 gnd.n2621 gnd.n2620 585
R8810 gnd.n2630 gnd.n2621 585
R8811 gnd.n3337 gnd.n3336 585
R8812 gnd.n3336 gnd.n3335 585
R8813 gnd.n2628 gnd.n2627 585
R8814 gnd.n3323 gnd.n2628 585
R8815 gnd.n2761 gnd.n2760 585
R8816 gnd.n2761 gnd.n2637 585
R8817 gnd.n3280 gnd.n3279 585
R8818 gnd.n3279 gnd.n3278 585
R8819 gnd.n3281 gnd.n2755 585
R8820 gnd.n2766 gnd.n2755 585
R8821 gnd.n3283 gnd.n3282 585
R8822 gnd.n3284 gnd.n3283 585
R8823 gnd.n2756 gnd.n2754 585
R8824 gnd.n2779 gnd.n2754 585
R8825 gnd.n2739 gnd.n2738 585
R8826 gnd.n2742 gnd.n2739 585
R8827 gnd.n3294 gnd.n3293 585
R8828 gnd.n3293 gnd.n3292 585
R8829 gnd.n3295 gnd.n2733 585
R8830 gnd.n3254 gnd.n2733 585
R8831 gnd.n3297 gnd.n3296 585
R8832 gnd.n3298 gnd.n3297 585
R8833 gnd.n2734 gnd.n2732 585
R8834 gnd.n2793 gnd.n2732 585
R8835 gnd.n3246 gnd.n3245 585
R8836 gnd.n3245 gnd.n3244 585
R8837 gnd.n2790 gnd.n2789 585
R8838 gnd.n3228 gnd.n2790 585
R8839 gnd.n3215 gnd.n2809 585
R8840 gnd.n2809 gnd.n2808 585
R8841 gnd.n3217 gnd.n3216 585
R8842 gnd.n3218 gnd.n3217 585
R8843 gnd.n2810 gnd.n2807 585
R8844 gnd.n2816 gnd.n2807 585
R8845 gnd.n3196 gnd.n3195 585
R8846 gnd.n3197 gnd.n3196 585
R8847 gnd.n2827 gnd.n2826 585
R8848 gnd.n2826 gnd.n2822 585
R8849 gnd.n3186 gnd.n3185 585
R8850 gnd.n3187 gnd.n3186 585
R8851 gnd.n2837 gnd.n2836 585
R8852 gnd.n2842 gnd.n2836 585
R8853 gnd.n3164 gnd.n2855 585
R8854 gnd.n2855 gnd.n2841 585
R8855 gnd.n3166 gnd.n3165 585
R8856 gnd.n3167 gnd.n3166 585
R8857 gnd.n2856 gnd.n2854 585
R8858 gnd.n2854 gnd.n2850 585
R8859 gnd.n3155 gnd.n3154 585
R8860 gnd.n3156 gnd.n3155 585
R8861 gnd.n2863 gnd.n2862 585
R8862 gnd.n2867 gnd.n2862 585
R8863 gnd.n3132 gnd.n2884 585
R8864 gnd.n2884 gnd.n2866 585
R8865 gnd.n3134 gnd.n3133 585
R8866 gnd.n3135 gnd.n3134 585
R8867 gnd.n2885 gnd.n2883 585
R8868 gnd.n2883 gnd.n2874 585
R8869 gnd.n3127 gnd.n3126 585
R8870 gnd.n3126 gnd.n3125 585
R8871 gnd.n2932 gnd.n2931 585
R8872 gnd.n2933 gnd.n2932 585
R8873 gnd.n3086 gnd.n3085 585
R8874 gnd.n3087 gnd.n3086 585
R8875 gnd.n2942 gnd.n2941 585
R8876 gnd.n2941 gnd.n2940 585
R8877 gnd.n3081 gnd.n3080 585
R8878 gnd.n3080 gnd.n3079 585
R8879 gnd.n2945 gnd.n2944 585
R8880 gnd.n2946 gnd.n2945 585
R8881 gnd.n3070 gnd.n3069 585
R8882 gnd.n3071 gnd.n3070 585
R8883 gnd.n2953 gnd.n2952 585
R8884 gnd.n3062 gnd.n2952 585
R8885 gnd.n3065 gnd.n3064 585
R8886 gnd.n3064 gnd.n3063 585
R8887 gnd.n2956 gnd.n2955 585
R8888 gnd.n2957 gnd.n2956 585
R8889 gnd.n3051 gnd.n3050 585
R8890 gnd.n3049 gnd.n2975 585
R8891 gnd.n3048 gnd.n2974 585
R8892 gnd.n3053 gnd.n2974 585
R8893 gnd.n3047 gnd.n3046 585
R8894 gnd.n3045 gnd.n3044 585
R8895 gnd.n3043 gnd.n3042 585
R8896 gnd.n3041 gnd.n3040 585
R8897 gnd.n3039 gnd.n3038 585
R8898 gnd.n3037 gnd.n3036 585
R8899 gnd.n3035 gnd.n3034 585
R8900 gnd.n3033 gnd.n3032 585
R8901 gnd.n3031 gnd.n3030 585
R8902 gnd.n3029 gnd.n3028 585
R8903 gnd.n3027 gnd.n3026 585
R8904 gnd.n3025 gnd.n3024 585
R8905 gnd.n3023 gnd.n3022 585
R8906 gnd.n3021 gnd.n3020 585
R8907 gnd.n3019 gnd.n3018 585
R8908 gnd.n3017 gnd.n3016 585
R8909 gnd.n3015 gnd.n3014 585
R8910 gnd.n3013 gnd.n3012 585
R8911 gnd.n3011 gnd.n3010 585
R8912 gnd.n3009 gnd.n3008 585
R8913 gnd.n3007 gnd.n3006 585
R8914 gnd.n3005 gnd.n3004 585
R8915 gnd.n2962 gnd.n2961 585
R8916 gnd.n3056 gnd.n3055 585
R8917 gnd.n3817 gnd.n3816 585
R8918 gnd.n3819 gnd.n3818 585
R8919 gnd.n3821 gnd.n3820 585
R8920 gnd.n3823 gnd.n3822 585
R8921 gnd.n3825 gnd.n3824 585
R8922 gnd.n3827 gnd.n3826 585
R8923 gnd.n3829 gnd.n3828 585
R8924 gnd.n3831 gnd.n3830 585
R8925 gnd.n3833 gnd.n3832 585
R8926 gnd.n3835 gnd.n3834 585
R8927 gnd.n3837 gnd.n3836 585
R8928 gnd.n3839 gnd.n3838 585
R8929 gnd.n3841 gnd.n3840 585
R8930 gnd.n3843 gnd.n3842 585
R8931 gnd.n3845 gnd.n3844 585
R8932 gnd.n3847 gnd.n3846 585
R8933 gnd.n3849 gnd.n3848 585
R8934 gnd.n3851 gnd.n3850 585
R8935 gnd.n3853 gnd.n3852 585
R8936 gnd.n3855 gnd.n3854 585
R8937 gnd.n3857 gnd.n3856 585
R8938 gnd.n3859 gnd.n3858 585
R8939 gnd.n3861 gnd.n3860 585
R8940 gnd.n3863 gnd.n3862 585
R8941 gnd.n3865 gnd.n3864 585
R8942 gnd.n3866 gnd.n2455 585
R8943 gnd.n3867 gnd.n2413 585
R8944 gnd.n3905 gnd.n2413 585
R8945 gnd.n3815 gnd.n2485 585
R8946 gnd.n3815 gnd.n3814 585
R8947 gnd.n3484 gnd.n2484 585
R8948 gnd.n2494 gnd.n2484 585
R8949 gnd.n3486 gnd.n3485 585
R8950 gnd.n3485 gnd.n2493 585
R8951 gnd.n3487 gnd.n2503 585
R8952 gnd.n3791 gnd.n2503 585
R8953 gnd.n3489 gnd.n3488 585
R8954 gnd.n3488 gnd.n2501 585
R8955 gnd.n3490 gnd.n2514 585
R8956 gnd.n3520 gnd.n2514 585
R8957 gnd.n3493 gnd.n3492 585
R8958 gnd.n3492 gnd.n3491 585
R8959 gnd.n3494 gnd.n2521 585
R8960 gnd.n3509 gnd.n2521 585
R8961 gnd.n3496 gnd.n3495 585
R8962 gnd.n3497 gnd.n3496 585
R8963 gnd.n2531 gnd.n2530 585
R8964 gnd.n2538 gnd.n2530 585
R8965 gnd.n3472 gnd.n3471 585
R8966 gnd.n3471 gnd.n3470 585
R8967 gnd.n2534 gnd.n2533 585
R8968 gnd.n2548 gnd.n2534 585
R8969 gnd.n3398 gnd.n3397 585
R8970 gnd.n3397 gnd.n2547 585
R8971 gnd.n3399 gnd.n2557 585
R8972 gnd.n3448 gnd.n2557 585
R8973 gnd.n3401 gnd.n3400 585
R8974 gnd.n3400 gnd.n2555 585
R8975 gnd.n3402 gnd.n2568 585
R8976 gnd.n3431 gnd.n2568 585
R8977 gnd.n3404 gnd.n3403 585
R8978 gnd.n3403 gnd.n2576 585
R8979 gnd.n3405 gnd.n2575 585
R8980 gnd.n3420 gnd.n2575 585
R8981 gnd.n3407 gnd.n3406 585
R8982 gnd.n3408 gnd.n3407 585
R8983 gnd.n2587 gnd.n2586 585
R8984 gnd.n2586 gnd.n2583 585
R8985 gnd.n3387 gnd.n3386 585
R8986 gnd.n3386 gnd.n3385 585
R8987 gnd.n2590 gnd.n2589 585
R8988 gnd.n2603 gnd.n2590 585
R8989 gnd.n3311 gnd.n3310 585
R8990 gnd.n3310 gnd.n2602 585
R8991 gnd.n3312 gnd.n2612 585
R8992 gnd.n3363 gnd.n2612 585
R8993 gnd.n3314 gnd.n3313 585
R8994 gnd.n3313 gnd.n2610 585
R8995 gnd.n3315 gnd.n2623 585
R8996 gnd.n3346 gnd.n2623 585
R8997 gnd.n3317 gnd.n3316 585
R8998 gnd.n3316 gnd.n2630 585
R8999 gnd.n3318 gnd.n2629 585
R9000 gnd.n3335 gnd.n2629 585
R9001 gnd.n3320 gnd.n3319 585
R9002 gnd.n3323 gnd.n3320 585
R9003 gnd.n2640 gnd.n2639 585
R9004 gnd.n2639 gnd.n2637 585
R9005 gnd.n2763 gnd.n2762 585
R9006 gnd.n3278 gnd.n2762 585
R9007 gnd.n2765 gnd.n2764 585
R9008 gnd.n2766 gnd.n2765 585
R9009 gnd.n2776 gnd.n2752 585
R9010 gnd.n3284 gnd.n2752 585
R9011 gnd.n2778 gnd.n2777 585
R9012 gnd.n2779 gnd.n2778 585
R9013 gnd.n2775 gnd.n2774 585
R9014 gnd.n2775 gnd.n2742 585
R9015 gnd.n2773 gnd.n2740 585
R9016 gnd.n3292 gnd.n2740 585
R9017 gnd.n2729 gnd.n2727 585
R9018 gnd.n3254 gnd.n2729 585
R9019 gnd.n3300 gnd.n3299 585
R9020 gnd.n3299 gnd.n3298 585
R9021 gnd.n2728 gnd.n2726 585
R9022 gnd.n2793 gnd.n2728 585
R9023 gnd.n3225 gnd.n2792 585
R9024 gnd.n3244 gnd.n2792 585
R9025 gnd.n3227 gnd.n3226 585
R9026 gnd.n3228 gnd.n3227 585
R9027 gnd.n2802 gnd.n2801 585
R9028 gnd.n2808 gnd.n2801 585
R9029 gnd.n3220 gnd.n3219 585
R9030 gnd.n3219 gnd.n3218 585
R9031 gnd.n2805 gnd.n2804 585
R9032 gnd.n2816 gnd.n2805 585
R9033 gnd.n3105 gnd.n2824 585
R9034 gnd.n3197 gnd.n2824 585
R9035 gnd.n3107 gnd.n3106 585
R9036 gnd.n3106 gnd.n2822 585
R9037 gnd.n3108 gnd.n2835 585
R9038 gnd.n3187 gnd.n2835 585
R9039 gnd.n3110 gnd.n3109 585
R9040 gnd.n3110 gnd.n2842 585
R9041 gnd.n3112 gnd.n3111 585
R9042 gnd.n3111 gnd.n2841 585
R9043 gnd.n3113 gnd.n2852 585
R9044 gnd.n3167 gnd.n2852 585
R9045 gnd.n3115 gnd.n3114 585
R9046 gnd.n3114 gnd.n2850 585
R9047 gnd.n3116 gnd.n2861 585
R9048 gnd.n3156 gnd.n2861 585
R9049 gnd.n3118 gnd.n3117 585
R9050 gnd.n3118 gnd.n2867 585
R9051 gnd.n3120 gnd.n3119 585
R9052 gnd.n3119 gnd.n2866 585
R9053 gnd.n3121 gnd.n2882 585
R9054 gnd.n3135 gnd.n2882 585
R9055 gnd.n3122 gnd.n2935 585
R9056 gnd.n2935 gnd.n2874 585
R9057 gnd.n3124 gnd.n3123 585
R9058 gnd.n3125 gnd.n3124 585
R9059 gnd.n2936 gnd.n2934 585
R9060 gnd.n2934 gnd.n2933 585
R9061 gnd.n3089 gnd.n3088 585
R9062 gnd.n3088 gnd.n3087 585
R9063 gnd.n2939 gnd.n2938 585
R9064 gnd.n2940 gnd.n2939 585
R9065 gnd.n3078 gnd.n3077 585
R9066 gnd.n3079 gnd.n3078 585
R9067 gnd.n2948 gnd.n2947 585
R9068 gnd.n2947 gnd.n2946 585
R9069 gnd.n3073 gnd.n3072 585
R9070 gnd.n3072 gnd.n3071 585
R9071 gnd.n2951 gnd.n2950 585
R9072 gnd.n3062 gnd.n2951 585
R9073 gnd.n3061 gnd.n3060 585
R9074 gnd.n3063 gnd.n3061 585
R9075 gnd.n2959 gnd.n2958 585
R9076 gnd.n2958 gnd.n2957 585
R9077 gnd.n3800 gnd.n2435 585
R9078 gnd.n2435 gnd.n2412 585
R9079 gnd.n3801 gnd.n2496 585
R9080 gnd.n2496 gnd.n2486 585
R9081 gnd.n3803 gnd.n3802 585
R9082 gnd.n3804 gnd.n3803 585
R9083 gnd.n2497 gnd.n2495 585
R9084 gnd.n2504 gnd.n2495 585
R9085 gnd.n3794 gnd.n3793 585
R9086 gnd.n3793 gnd.n3792 585
R9087 gnd.n2500 gnd.n2499 585
R9088 gnd.n3519 gnd.n2500 585
R9089 gnd.n3505 gnd.n2523 585
R9090 gnd.n2523 gnd.n2513 585
R9091 gnd.n3507 gnd.n3506 585
R9092 gnd.n3508 gnd.n3507 585
R9093 gnd.n2524 gnd.n2522 585
R9094 gnd.n2522 gnd.n2520 585
R9095 gnd.n3500 gnd.n3499 585
R9096 gnd.n3499 gnd.n3498 585
R9097 gnd.n2527 gnd.n2526 585
R9098 gnd.n2536 gnd.n2527 585
R9099 gnd.n3456 gnd.n2550 585
R9100 gnd.n2550 gnd.n2535 585
R9101 gnd.n3458 gnd.n3457 585
R9102 gnd.n3459 gnd.n3458 585
R9103 gnd.n2551 gnd.n2549 585
R9104 gnd.n2558 gnd.n2549 585
R9105 gnd.n3451 gnd.n3450 585
R9106 gnd.n3450 gnd.n3449 585
R9107 gnd.n2554 gnd.n2553 585
R9108 gnd.n3430 gnd.n2554 585
R9109 gnd.n3416 gnd.n2578 585
R9110 gnd.n2578 gnd.n2567 585
R9111 gnd.n3418 gnd.n3417 585
R9112 gnd.n3419 gnd.n3418 585
R9113 gnd.n2579 gnd.n2577 585
R9114 gnd.n2577 gnd.n2574 585
R9115 gnd.n3411 gnd.n3410 585
R9116 gnd.n3410 gnd.n3409 585
R9117 gnd.n2582 gnd.n2581 585
R9118 gnd.n2592 gnd.n2582 585
R9119 gnd.n3371 gnd.n2605 585
R9120 gnd.n2605 gnd.n2591 585
R9121 gnd.n3373 gnd.n3372 585
R9122 gnd.n3374 gnd.n3373 585
R9123 gnd.n2606 gnd.n2604 585
R9124 gnd.n2613 gnd.n2604 585
R9125 gnd.n3366 gnd.n3365 585
R9126 gnd.n3365 gnd.n3364 585
R9127 gnd.n2609 gnd.n2608 585
R9128 gnd.n3345 gnd.n2609 585
R9129 gnd.n3331 gnd.n2632 585
R9130 gnd.n2632 gnd.n2622 585
R9131 gnd.n3333 gnd.n3332 585
R9132 gnd.n3334 gnd.n3333 585
R9133 gnd.n2633 gnd.n2631 585
R9134 gnd.n3322 gnd.n2631 585
R9135 gnd.n3326 gnd.n3325 585
R9136 gnd.n3325 gnd.n3324 585
R9137 gnd.n2636 gnd.n2635 585
R9138 gnd.n3277 gnd.n2636 585
R9139 gnd.n2770 gnd.n2769 585
R9140 gnd.n2771 gnd.n2770 585
R9141 gnd.n2750 gnd.n2749 585
R9142 gnd.n2753 gnd.n2750 585
R9143 gnd.n3287 gnd.n3286 585
R9144 gnd.n3286 gnd.n3285 585
R9145 gnd.n3288 gnd.n2744 585
R9146 gnd.n2780 gnd.n2744 585
R9147 gnd.n3290 gnd.n3289 585
R9148 gnd.n3291 gnd.n3290 585
R9149 gnd.n2745 gnd.n2743 585
R9150 gnd.n3255 gnd.n2743 585
R9151 gnd.n3239 gnd.n3238 585
R9152 gnd.n3238 gnd.n2731 585
R9153 gnd.n3240 gnd.n2795 585
R9154 gnd.n2795 gnd.n2730 585
R9155 gnd.n3242 gnd.n3241 585
R9156 gnd.n3243 gnd.n3242 585
R9157 gnd.n2796 gnd.n2794 585
R9158 gnd.n2794 gnd.n2791 585
R9159 gnd.n3231 gnd.n3230 585
R9160 gnd.n3230 gnd.n3229 585
R9161 gnd.n2799 gnd.n2798 585
R9162 gnd.n2806 gnd.n2799 585
R9163 gnd.n3205 gnd.n3204 585
R9164 gnd.n3206 gnd.n3205 585
R9165 gnd.n2818 gnd.n2817 585
R9166 gnd.n2825 gnd.n2817 585
R9167 gnd.n3200 gnd.n3199 585
R9168 gnd.n3199 gnd.n3198 585
R9169 gnd.n2821 gnd.n2820 585
R9170 gnd.n3188 gnd.n2821 585
R9171 gnd.n3175 gnd.n2845 585
R9172 gnd.n2845 gnd.n2844 585
R9173 gnd.n3177 gnd.n3176 585
R9174 gnd.n3178 gnd.n3177 585
R9175 gnd.n2846 gnd.n2843 585
R9176 gnd.n2853 gnd.n2843 585
R9177 gnd.n3170 gnd.n3169 585
R9178 gnd.n3169 gnd.n3168 585
R9179 gnd.n2849 gnd.n2848 585
R9180 gnd.n3157 gnd.n2849 585
R9181 gnd.n3144 gnd.n2870 585
R9182 gnd.n2870 gnd.n2869 585
R9183 gnd.n3146 gnd.n3145 585
R9184 gnd.n3147 gnd.n3146 585
R9185 gnd.n3140 gnd.n2868 585
R9186 gnd.n3139 gnd.n3138 585
R9187 gnd.n2873 gnd.n2872 585
R9188 gnd.n3136 gnd.n2873 585
R9189 gnd.n2895 gnd.n2894 585
R9190 gnd.n2898 gnd.n2897 585
R9191 gnd.n2896 gnd.n2891 585
R9192 gnd.n2903 gnd.n2902 585
R9193 gnd.n2905 gnd.n2904 585
R9194 gnd.n2908 gnd.n2907 585
R9195 gnd.n2906 gnd.n2889 585
R9196 gnd.n2913 gnd.n2912 585
R9197 gnd.n2915 gnd.n2914 585
R9198 gnd.n2918 gnd.n2917 585
R9199 gnd.n2916 gnd.n2887 585
R9200 gnd.n2923 gnd.n2922 585
R9201 gnd.n2927 gnd.n2924 585
R9202 gnd.n2928 gnd.n2865 585
R9203 gnd.n3806 gnd.n2450 585
R9204 gnd.n3873 gnd.n3872 585
R9205 gnd.n3875 gnd.n3874 585
R9206 gnd.n3877 gnd.n3876 585
R9207 gnd.n3879 gnd.n3878 585
R9208 gnd.n3881 gnd.n3880 585
R9209 gnd.n3883 gnd.n3882 585
R9210 gnd.n3885 gnd.n3884 585
R9211 gnd.n3887 gnd.n3886 585
R9212 gnd.n3889 gnd.n3888 585
R9213 gnd.n3891 gnd.n3890 585
R9214 gnd.n3893 gnd.n3892 585
R9215 gnd.n3895 gnd.n3894 585
R9216 gnd.n3898 gnd.n3897 585
R9217 gnd.n3896 gnd.n2438 585
R9218 gnd.n3902 gnd.n2436 585
R9219 gnd.n3904 gnd.n3903 585
R9220 gnd.n3905 gnd.n3904 585
R9221 gnd.n3807 gnd.n2491 585
R9222 gnd.n3807 gnd.n2412 585
R9223 gnd.n3809 gnd.n3808 585
R9224 gnd.n3808 gnd.n2486 585
R9225 gnd.n3805 gnd.n2490 585
R9226 gnd.n3805 gnd.n3804 585
R9227 gnd.n3784 gnd.n2492 585
R9228 gnd.n2504 gnd.n2492 585
R9229 gnd.n3783 gnd.n2502 585
R9230 gnd.n3792 gnd.n2502 585
R9231 gnd.n3518 gnd.n2509 585
R9232 gnd.n3519 gnd.n3518 585
R9233 gnd.n3517 gnd.n3516 585
R9234 gnd.n3517 gnd.n2513 585
R9235 gnd.n3515 gnd.n2515 585
R9236 gnd.n3508 gnd.n2515 585
R9237 gnd.n2528 gnd.n2516 585
R9238 gnd.n2528 gnd.n2520 585
R9239 gnd.n3464 gnd.n2529 585
R9240 gnd.n3498 gnd.n2529 585
R9241 gnd.n3463 gnd.n3462 585
R9242 gnd.n3462 gnd.n2536 585
R9243 gnd.n3461 gnd.n2544 585
R9244 gnd.n3461 gnd.n2535 585
R9245 gnd.n3460 gnd.n2546 585
R9246 gnd.n3460 gnd.n3459 585
R9247 gnd.n3439 gnd.n2545 585
R9248 gnd.n2558 gnd.n2545 585
R9249 gnd.n3438 gnd.n2556 585
R9250 gnd.n3449 gnd.n2556 585
R9251 gnd.n3429 gnd.n2563 585
R9252 gnd.n3430 gnd.n3429 585
R9253 gnd.n3428 gnd.n3427 585
R9254 gnd.n3428 gnd.n2567 585
R9255 gnd.n3426 gnd.n2569 585
R9256 gnd.n3419 gnd.n2569 585
R9257 gnd.n2584 gnd.n2570 585
R9258 gnd.n2584 gnd.n2574 585
R9259 gnd.n3379 gnd.n2585 585
R9260 gnd.n3409 gnd.n2585 585
R9261 gnd.n3378 gnd.n3377 585
R9262 gnd.n3377 gnd.n2592 585
R9263 gnd.n3376 gnd.n2599 585
R9264 gnd.n3376 gnd.n2591 585
R9265 gnd.n3375 gnd.n2601 585
R9266 gnd.n3375 gnd.n3374 585
R9267 gnd.n3354 gnd.n2600 585
R9268 gnd.n2613 gnd.n2600 585
R9269 gnd.n3353 gnd.n2611 585
R9270 gnd.n3364 gnd.n2611 585
R9271 gnd.n3344 gnd.n2618 585
R9272 gnd.n3345 gnd.n3344 585
R9273 gnd.n3343 gnd.n3342 585
R9274 gnd.n3343 gnd.n2622 585
R9275 gnd.n3341 gnd.n2624 585
R9276 gnd.n3334 gnd.n2624 585
R9277 gnd.n3321 gnd.n2625 585
R9278 gnd.n3322 gnd.n3321 585
R9279 gnd.n3274 gnd.n2638 585
R9280 gnd.n3324 gnd.n2638 585
R9281 gnd.n3276 gnd.n3275 585
R9282 gnd.n3277 gnd.n3276 585
R9283 gnd.n3269 gnd.n2772 585
R9284 gnd.n2772 gnd.n2771 585
R9285 gnd.n3267 gnd.n3266 585
R9286 gnd.n3266 gnd.n2753 585
R9287 gnd.n3264 gnd.n2751 585
R9288 gnd.n3285 gnd.n2751 585
R9289 gnd.n2782 gnd.n2781 585
R9290 gnd.n2781 gnd.n2780 585
R9291 gnd.n3258 gnd.n2741 585
R9292 gnd.n3291 gnd.n2741 585
R9293 gnd.n3257 gnd.n3256 585
R9294 gnd.n3256 gnd.n3255 585
R9295 gnd.n3253 gnd.n2784 585
R9296 gnd.n3253 gnd.n2731 585
R9297 gnd.n3252 gnd.n3251 585
R9298 gnd.n3252 gnd.n2730 585
R9299 gnd.n2787 gnd.n2786 585
R9300 gnd.n3243 gnd.n2786 585
R9301 gnd.n3211 gnd.n3210 585
R9302 gnd.n3210 gnd.n2791 585
R9303 gnd.n3212 gnd.n2800 585
R9304 gnd.n3229 gnd.n2800 585
R9305 gnd.n3209 gnd.n3208 585
R9306 gnd.n3208 gnd.n2806 585
R9307 gnd.n3207 gnd.n2814 585
R9308 gnd.n3207 gnd.n3206 585
R9309 gnd.n3192 gnd.n2815 585
R9310 gnd.n2825 gnd.n2815 585
R9311 gnd.n3191 gnd.n2823 585
R9312 gnd.n3198 gnd.n2823 585
R9313 gnd.n3190 gnd.n3189 585
R9314 gnd.n3189 gnd.n3188 585
R9315 gnd.n2834 gnd.n2831 585
R9316 gnd.n2844 gnd.n2834 585
R9317 gnd.n3180 gnd.n3179 585
R9318 gnd.n3179 gnd.n3178 585
R9319 gnd.n2840 gnd.n2839 585
R9320 gnd.n2853 gnd.n2840 585
R9321 gnd.n3160 gnd.n2851 585
R9322 gnd.n3168 gnd.n2851 585
R9323 gnd.n3159 gnd.n3158 585
R9324 gnd.n3158 gnd.n3157 585
R9325 gnd.n2860 gnd.n2858 585
R9326 gnd.n2869 gnd.n2860 585
R9327 gnd.n3149 gnd.n3148 585
R9328 gnd.n3148 gnd.n3147 585
R9329 gnd.n6451 gnd.n6450 585
R9330 gnd.n6452 gnd.n6451 585
R9331 gnd.n759 gnd.n757 585
R9332 gnd.n4547 gnd.n757 585
R9333 gnd.n4532 gnd.n2197 585
R9334 gnd.n2197 gnd.n2185 585
R9335 gnd.n4534 gnd.n4533 585
R9336 gnd.n4535 gnd.n4534 585
R9337 gnd.n2198 gnd.n2196 585
R9338 gnd.n2196 gnd.n2193 585
R9339 gnd.n4526 gnd.n4525 585
R9340 gnd.n4525 gnd.n4524 585
R9341 gnd.n2201 gnd.n2200 585
R9342 gnd.n4508 gnd.n2201 585
R9343 gnd.n4496 gnd.n2223 585
R9344 gnd.n2223 gnd.n2212 585
R9345 gnd.n4498 gnd.n4497 585
R9346 gnd.n4499 gnd.n4498 585
R9347 gnd.n2224 gnd.n2222 585
R9348 gnd.n2222 gnd.n2219 585
R9349 gnd.n4491 gnd.n4490 585
R9350 gnd.n4490 gnd.n4489 585
R9351 gnd.n2227 gnd.n2226 585
R9352 gnd.n4474 gnd.n2227 585
R9353 gnd.n4462 gnd.n2248 585
R9354 gnd.n2248 gnd.n2238 585
R9355 gnd.n4464 gnd.n4463 585
R9356 gnd.n4465 gnd.n4464 585
R9357 gnd.n2249 gnd.n2247 585
R9358 gnd.n2255 gnd.n2247 585
R9359 gnd.n4457 gnd.n4456 585
R9360 gnd.n4456 gnd.n4455 585
R9361 gnd.n2252 gnd.n2251 585
R9362 gnd.n4440 gnd.n2252 585
R9363 gnd.n4428 gnd.n2274 585
R9364 gnd.n2274 gnd.n2264 585
R9365 gnd.n4430 gnd.n4429 585
R9366 gnd.n4431 gnd.n4430 585
R9367 gnd.n2275 gnd.n2273 585
R9368 gnd.n2281 gnd.n2273 585
R9369 gnd.n4423 gnd.n4422 585
R9370 gnd.n4422 gnd.n4421 585
R9371 gnd.n2278 gnd.n2277 585
R9372 gnd.n4406 gnd.n2278 585
R9373 gnd.n4393 gnd.n2299 585
R9374 gnd.n2299 gnd.n2290 585
R9375 gnd.n4395 gnd.n4394 585
R9376 gnd.n4396 gnd.n4395 585
R9377 gnd.n2300 gnd.n2298 585
R9378 gnd.n2307 gnd.n2298 585
R9379 gnd.n4388 gnd.n4387 585
R9380 gnd.n4387 gnd.n4386 585
R9381 gnd.n2303 gnd.n2302 585
R9382 gnd.n2304 gnd.n2303 585
R9383 gnd.n4369 gnd.n4368 585
R9384 gnd.n4370 gnd.n4369 585
R9385 gnd.n2320 gnd.n2319 585
R9386 gnd.n2319 gnd.n2316 585
R9387 gnd.n4364 gnd.n4363 585
R9388 gnd.n4363 gnd.n4362 585
R9389 gnd.n2323 gnd.n2322 585
R9390 gnd.n2324 gnd.n2323 585
R9391 gnd.n4349 gnd.n4348 585
R9392 gnd.n4350 gnd.n4349 585
R9393 gnd.n2337 gnd.n2336 585
R9394 gnd.n2344 gnd.n2336 585
R9395 gnd.n4344 gnd.n4343 585
R9396 gnd.n4343 gnd.n4342 585
R9397 gnd.n2340 gnd.n2339 585
R9398 gnd.n2341 gnd.n2340 585
R9399 gnd.n4329 gnd.n4328 585
R9400 gnd.n4330 gnd.n4329 585
R9401 gnd.n2356 gnd.n2355 585
R9402 gnd.n2355 gnd.n2352 585
R9403 gnd.n4324 gnd.n4323 585
R9404 gnd.n4323 gnd.n4322 585
R9405 gnd.n2359 gnd.n2358 585
R9406 gnd.n2360 gnd.n2359 585
R9407 gnd.n4309 gnd.n4308 585
R9408 gnd.n4310 gnd.n4309 585
R9409 gnd.n2373 gnd.n2372 585
R9410 gnd.n2380 gnd.n2372 585
R9411 gnd.n4304 gnd.n4303 585
R9412 gnd.n4303 gnd.n4302 585
R9413 gnd.n2376 gnd.n2375 585
R9414 gnd.n2377 gnd.n2376 585
R9415 gnd.n4289 gnd.n4288 585
R9416 gnd.n4290 gnd.n4289 585
R9417 gnd.n2392 gnd.n2391 585
R9418 gnd.n2391 gnd.n2388 585
R9419 gnd.n4284 gnd.n4283 585
R9420 gnd.n4283 gnd.n4282 585
R9421 gnd.n2395 gnd.n2394 585
R9422 gnd.n2396 gnd.n2395 585
R9423 gnd.n4269 gnd.n4268 585
R9424 gnd.n4270 gnd.n4269 585
R9425 gnd.n2409 gnd.n2408 585
R9426 gnd.n3909 gnd.n2408 585
R9427 gnd.n4264 gnd.n4263 585
R9428 gnd.n4263 gnd.n4262 585
R9429 gnd.n3974 gnd.n2411 585
R9430 gnd.n3977 gnd.n3976 585
R9431 gnd.n3973 gnd.n3972 585
R9432 gnd.n3972 gnd.n3906 585
R9433 gnd.n3982 gnd.n3981 585
R9434 gnd.n3984 gnd.n3971 585
R9435 gnd.n3987 gnd.n3986 585
R9436 gnd.n3969 gnd.n3968 585
R9437 gnd.n3992 gnd.n3991 585
R9438 gnd.n3994 gnd.n3967 585
R9439 gnd.n3997 gnd.n3996 585
R9440 gnd.n3965 gnd.n3964 585
R9441 gnd.n4002 gnd.n4001 585
R9442 gnd.n4004 gnd.n3963 585
R9443 gnd.n4007 gnd.n4006 585
R9444 gnd.n3961 gnd.n3960 585
R9445 gnd.n4012 gnd.n4011 585
R9446 gnd.n4014 gnd.n3956 585
R9447 gnd.n4017 gnd.n4016 585
R9448 gnd.n3954 gnd.n3953 585
R9449 gnd.n4022 gnd.n4021 585
R9450 gnd.n4024 gnd.n3952 585
R9451 gnd.n4027 gnd.n4026 585
R9452 gnd.n3950 gnd.n3949 585
R9453 gnd.n4032 gnd.n4031 585
R9454 gnd.n4034 gnd.n3948 585
R9455 gnd.n4037 gnd.n4036 585
R9456 gnd.n3946 gnd.n3945 585
R9457 gnd.n4042 gnd.n4041 585
R9458 gnd.n4044 gnd.n3944 585
R9459 gnd.n4047 gnd.n4046 585
R9460 gnd.n3942 gnd.n3941 585
R9461 gnd.n4052 gnd.n4051 585
R9462 gnd.n4054 gnd.n3940 585
R9463 gnd.n4057 gnd.n4056 585
R9464 gnd.n3938 gnd.n3937 585
R9465 gnd.n4062 gnd.n4061 585
R9466 gnd.n4064 gnd.n3936 585
R9467 gnd.n4069 gnd.n4066 585
R9468 gnd.n3934 gnd.n3933 585
R9469 gnd.n4074 gnd.n4073 585
R9470 gnd.n4076 gnd.n3932 585
R9471 gnd.n4079 gnd.n4078 585
R9472 gnd.n3930 gnd.n3929 585
R9473 gnd.n4084 gnd.n4083 585
R9474 gnd.n4086 gnd.n3928 585
R9475 gnd.n4089 gnd.n4088 585
R9476 gnd.n3926 gnd.n3925 585
R9477 gnd.n4094 gnd.n4093 585
R9478 gnd.n4096 gnd.n3924 585
R9479 gnd.n4099 gnd.n4098 585
R9480 gnd.n3922 gnd.n3921 585
R9481 gnd.n4104 gnd.n4103 585
R9482 gnd.n4106 gnd.n3920 585
R9483 gnd.n4109 gnd.n4108 585
R9484 gnd.n3918 gnd.n3917 585
R9485 gnd.n4115 gnd.n4114 585
R9486 gnd.n4117 gnd.n3916 585
R9487 gnd.n4118 gnd.n3915 585
R9488 gnd.n4121 gnd.n4120 585
R9489 gnd.n2181 gnd.n754 585
R9490 gnd.n6452 gnd.n754 585
R9491 gnd.n4515 gnd.n2186 585
R9492 gnd.n4547 gnd.n2186 585
R9493 gnd.n4517 gnd.n4516 585
R9494 gnd.n4516 gnd.n2185 585
R9495 gnd.n4514 gnd.n2194 585
R9496 gnd.n4535 gnd.n2194 585
R9497 gnd.n4513 gnd.n4512 585
R9498 gnd.n4512 gnd.n2193 585
R9499 gnd.n4511 gnd.n2202 585
R9500 gnd.n4524 gnd.n2202 585
R9501 gnd.n4510 gnd.n4509 585
R9502 gnd.n4509 gnd.n4508 585
R9503 gnd.n2211 gnd.n2209 585
R9504 gnd.n2212 gnd.n2211 585
R9505 gnd.n4480 gnd.n2220 585
R9506 gnd.n4499 gnd.n2220 585
R9507 gnd.n4479 gnd.n4478 585
R9508 gnd.n4478 gnd.n2219 585
R9509 gnd.n4477 gnd.n2228 585
R9510 gnd.n4489 gnd.n2228 585
R9511 gnd.n4476 gnd.n4475 585
R9512 gnd.n4475 gnd.n4474 585
R9513 gnd.n2237 gnd.n2235 585
R9514 gnd.n2238 gnd.n2237 585
R9515 gnd.n4446 gnd.n2245 585
R9516 gnd.n4465 gnd.n2245 585
R9517 gnd.n4445 gnd.n4444 585
R9518 gnd.n4444 gnd.n2255 585
R9519 gnd.n4443 gnd.n2253 585
R9520 gnd.n4455 gnd.n2253 585
R9521 gnd.n4442 gnd.n4441 585
R9522 gnd.n4441 gnd.n4440 585
R9523 gnd.n2263 gnd.n2261 585
R9524 gnd.n2264 gnd.n2263 585
R9525 gnd.n4412 gnd.n2271 585
R9526 gnd.n4431 gnd.n2271 585
R9527 gnd.n4411 gnd.n4410 585
R9528 gnd.n4410 gnd.n2281 585
R9529 gnd.n4409 gnd.n2279 585
R9530 gnd.n4421 gnd.n2279 585
R9531 gnd.n4408 gnd.n4407 585
R9532 gnd.n4407 gnd.n4406 585
R9533 gnd.n2289 gnd.n2287 585
R9534 gnd.n2290 gnd.n2289 585
R9535 gnd.n4377 gnd.n2296 585
R9536 gnd.n4396 gnd.n2296 585
R9537 gnd.n4376 gnd.n4375 585
R9538 gnd.n4375 gnd.n2307 585
R9539 gnd.n4374 gnd.n2305 585
R9540 gnd.n4386 gnd.n2305 585
R9541 gnd.n4373 gnd.n4372 585
R9542 gnd.n4372 gnd.n2304 585
R9543 gnd.n4371 gnd.n2313 585
R9544 gnd.n4371 gnd.n4370 585
R9545 gnd.n4355 gnd.n2315 585
R9546 gnd.n2316 gnd.n2315 585
R9547 gnd.n4354 gnd.n2325 585
R9548 gnd.n4362 gnd.n2325 585
R9549 gnd.n4353 gnd.n4352 585
R9550 gnd.n4352 gnd.n2324 585
R9551 gnd.n4351 gnd.n2331 585
R9552 gnd.n4351 gnd.n4350 585
R9553 gnd.n4335 gnd.n2333 585
R9554 gnd.n2344 gnd.n2333 585
R9555 gnd.n4334 gnd.n2342 585
R9556 gnd.n4342 gnd.n2342 585
R9557 gnd.n4333 gnd.n4332 585
R9558 gnd.n4332 gnd.n2341 585
R9559 gnd.n4331 gnd.n2349 585
R9560 gnd.n4331 gnd.n4330 585
R9561 gnd.n4315 gnd.n2351 585
R9562 gnd.n2352 gnd.n2351 585
R9563 gnd.n4314 gnd.n2361 585
R9564 gnd.n4322 gnd.n2361 585
R9565 gnd.n4313 gnd.n4312 585
R9566 gnd.n4312 gnd.n2360 585
R9567 gnd.n4311 gnd.n2367 585
R9568 gnd.n4311 gnd.n4310 585
R9569 gnd.n4295 gnd.n2369 585
R9570 gnd.n2380 gnd.n2369 585
R9571 gnd.n4294 gnd.n2378 585
R9572 gnd.n4302 gnd.n2378 585
R9573 gnd.n4293 gnd.n4292 585
R9574 gnd.n4292 gnd.n2377 585
R9575 gnd.n4291 gnd.n2385 585
R9576 gnd.n4291 gnd.n4290 585
R9577 gnd.n4275 gnd.n2387 585
R9578 gnd.n2388 gnd.n2387 585
R9579 gnd.n4274 gnd.n2397 585
R9580 gnd.n4282 gnd.n2397 585
R9581 gnd.n4273 gnd.n4272 585
R9582 gnd.n4272 gnd.n2396 585
R9583 gnd.n4271 gnd.n2403 585
R9584 gnd.n4271 gnd.n4270 585
R9585 gnd.n4255 gnd.n2405 585
R9586 gnd.n3909 gnd.n2405 585
R9587 gnd.n4254 gnd.n3907 585
R9588 gnd.n4262 gnd.n3907 585
R9589 gnd.n4654 gnd.n751 585
R9590 gnd.n4658 gnd.n4656 585
R9591 gnd.n4659 gnd.n4653 585
R9592 gnd.n4659 gnd.n753 585
R9593 gnd.n4662 gnd.n4661 585
R9594 gnd.n4651 gnd.n4650 585
R9595 gnd.n4667 gnd.n4666 585
R9596 gnd.n4669 gnd.n4649 585
R9597 gnd.n4672 gnd.n4671 585
R9598 gnd.n4647 gnd.n4646 585
R9599 gnd.n4677 gnd.n4676 585
R9600 gnd.n4679 gnd.n4645 585
R9601 gnd.n4682 gnd.n4681 585
R9602 gnd.n4643 gnd.n4642 585
R9603 gnd.n4687 gnd.n4686 585
R9604 gnd.n4689 gnd.n4641 585
R9605 gnd.n4692 gnd.n4691 585
R9606 gnd.n4639 gnd.n4638 585
R9607 gnd.n4697 gnd.n4696 585
R9608 gnd.n4699 gnd.n4637 585
R9609 gnd.n4702 gnd.n4701 585
R9610 gnd.n4635 gnd.n4634 585
R9611 gnd.n4707 gnd.n4706 585
R9612 gnd.n4709 gnd.n4633 585
R9613 gnd.n4712 gnd.n4711 585
R9614 gnd.n4631 gnd.n4630 585
R9615 gnd.n4717 gnd.n4716 585
R9616 gnd.n4719 gnd.n4629 585
R9617 gnd.n4722 gnd.n4721 585
R9618 gnd.n4627 gnd.n4626 585
R9619 gnd.n4727 gnd.n4726 585
R9620 gnd.n4729 gnd.n4625 585
R9621 gnd.n4732 gnd.n4731 585
R9622 gnd.n4623 gnd.n4622 585
R9623 gnd.n4737 gnd.n4736 585
R9624 gnd.n4739 gnd.n4621 585
R9625 gnd.n4742 gnd.n4741 585
R9626 gnd.n4619 gnd.n4618 585
R9627 gnd.n4747 gnd.n4746 585
R9628 gnd.n4749 gnd.n4617 585
R9629 gnd.n4752 gnd.n4751 585
R9630 gnd.n4615 gnd.n4614 585
R9631 gnd.n4757 gnd.n4756 585
R9632 gnd.n4759 gnd.n4613 585
R9633 gnd.n4762 gnd.n4761 585
R9634 gnd.n4611 gnd.n4610 585
R9635 gnd.n4767 gnd.n4766 585
R9636 gnd.n4769 gnd.n4609 585
R9637 gnd.n4772 gnd.n4771 585
R9638 gnd.n4607 gnd.n4606 585
R9639 gnd.n4777 gnd.n4776 585
R9640 gnd.n4779 gnd.n4605 585
R9641 gnd.n4782 gnd.n4781 585
R9642 gnd.n4603 gnd.n4602 585
R9643 gnd.n4787 gnd.n4786 585
R9644 gnd.n4789 gnd.n4601 585
R9645 gnd.n4792 gnd.n4791 585
R9646 gnd.n4599 gnd.n4598 585
R9647 gnd.n4797 gnd.n4796 585
R9648 gnd.n4799 gnd.n4597 585
R9649 gnd.n4802 gnd.n4801 585
R9650 gnd.n4595 gnd.n4594 585
R9651 gnd.n4807 gnd.n4806 585
R9652 gnd.n4809 gnd.n4593 585
R9653 gnd.n4812 gnd.n4811 585
R9654 gnd.n4591 gnd.n4590 585
R9655 gnd.n4817 gnd.n4816 585
R9656 gnd.n4819 gnd.n4589 585
R9657 gnd.n4822 gnd.n4821 585
R9658 gnd.n4587 gnd.n4586 585
R9659 gnd.n4827 gnd.n4826 585
R9660 gnd.n4829 gnd.n4585 585
R9661 gnd.n4832 gnd.n4831 585
R9662 gnd.n4583 gnd.n4582 585
R9663 gnd.n4837 gnd.n4836 585
R9664 gnd.n4839 gnd.n4581 585
R9665 gnd.n4842 gnd.n4841 585
R9666 gnd.n4579 gnd.n4578 585
R9667 gnd.n4847 gnd.n4846 585
R9668 gnd.n4849 gnd.n4577 585
R9669 gnd.n4852 gnd.n4851 585
R9670 gnd.n4575 gnd.n4574 585
R9671 gnd.n4858 gnd.n4857 585
R9672 gnd.n4860 gnd.n4573 585
R9673 gnd.n4863 gnd.n4862 585
R9674 gnd.n4864 gnd.n4571 585
R9675 gnd.n6456 gnd.n6455 585
R9676 gnd.n6455 gnd.n6454 585
R9677 gnd.n749 gnd.n748 585
R9678 gnd.n748 gnd.n747 585
R9679 gnd.n6461 gnd.n6460 585
R9680 gnd.n6462 gnd.n6461 585
R9681 gnd.n746 gnd.n745 585
R9682 gnd.n6463 gnd.n746 585
R9683 gnd.n6466 gnd.n6465 585
R9684 gnd.n6465 gnd.n6464 585
R9685 gnd.n743 gnd.n742 585
R9686 gnd.n742 gnd.n741 585
R9687 gnd.n6471 gnd.n6470 585
R9688 gnd.n6472 gnd.n6471 585
R9689 gnd.n740 gnd.n739 585
R9690 gnd.n6473 gnd.n740 585
R9691 gnd.n6476 gnd.n6475 585
R9692 gnd.n6475 gnd.n6474 585
R9693 gnd.n737 gnd.n736 585
R9694 gnd.n736 gnd.n735 585
R9695 gnd.n6481 gnd.n6480 585
R9696 gnd.n6482 gnd.n6481 585
R9697 gnd.n734 gnd.n733 585
R9698 gnd.n6483 gnd.n734 585
R9699 gnd.n6486 gnd.n6485 585
R9700 gnd.n6485 gnd.n6484 585
R9701 gnd.n731 gnd.n730 585
R9702 gnd.n730 gnd.n729 585
R9703 gnd.n6491 gnd.n6490 585
R9704 gnd.n6492 gnd.n6491 585
R9705 gnd.n728 gnd.n727 585
R9706 gnd.n6493 gnd.n728 585
R9707 gnd.n6496 gnd.n6495 585
R9708 gnd.n6495 gnd.n6494 585
R9709 gnd.n725 gnd.n724 585
R9710 gnd.n724 gnd.n723 585
R9711 gnd.n6501 gnd.n6500 585
R9712 gnd.n6502 gnd.n6501 585
R9713 gnd.n722 gnd.n721 585
R9714 gnd.n6503 gnd.n722 585
R9715 gnd.n6506 gnd.n6505 585
R9716 gnd.n6505 gnd.n6504 585
R9717 gnd.n719 gnd.n718 585
R9718 gnd.n718 gnd.n717 585
R9719 gnd.n6511 gnd.n6510 585
R9720 gnd.n6512 gnd.n6511 585
R9721 gnd.n716 gnd.n715 585
R9722 gnd.n6513 gnd.n716 585
R9723 gnd.n6516 gnd.n6515 585
R9724 gnd.n6515 gnd.n6514 585
R9725 gnd.n713 gnd.n712 585
R9726 gnd.n712 gnd.n711 585
R9727 gnd.n6521 gnd.n6520 585
R9728 gnd.n6522 gnd.n6521 585
R9729 gnd.n710 gnd.n709 585
R9730 gnd.n6523 gnd.n710 585
R9731 gnd.n6526 gnd.n6525 585
R9732 gnd.n6525 gnd.n6524 585
R9733 gnd.n707 gnd.n706 585
R9734 gnd.n706 gnd.n705 585
R9735 gnd.n6531 gnd.n6530 585
R9736 gnd.n6532 gnd.n6531 585
R9737 gnd.n704 gnd.n703 585
R9738 gnd.n6533 gnd.n704 585
R9739 gnd.n6536 gnd.n6535 585
R9740 gnd.n6535 gnd.n6534 585
R9741 gnd.n701 gnd.n700 585
R9742 gnd.n700 gnd.n699 585
R9743 gnd.n6541 gnd.n6540 585
R9744 gnd.n6542 gnd.n6541 585
R9745 gnd.n698 gnd.n697 585
R9746 gnd.n6543 gnd.n698 585
R9747 gnd.n6546 gnd.n6545 585
R9748 gnd.n6545 gnd.n6544 585
R9749 gnd.n695 gnd.n694 585
R9750 gnd.n694 gnd.n693 585
R9751 gnd.n6551 gnd.n6550 585
R9752 gnd.n6552 gnd.n6551 585
R9753 gnd.n692 gnd.n691 585
R9754 gnd.n6553 gnd.n692 585
R9755 gnd.n6556 gnd.n6555 585
R9756 gnd.n6555 gnd.n6554 585
R9757 gnd.n689 gnd.n688 585
R9758 gnd.n688 gnd.n687 585
R9759 gnd.n6561 gnd.n6560 585
R9760 gnd.n6562 gnd.n6561 585
R9761 gnd.n686 gnd.n685 585
R9762 gnd.n6563 gnd.n686 585
R9763 gnd.n6566 gnd.n6565 585
R9764 gnd.n6565 gnd.n6564 585
R9765 gnd.n683 gnd.n682 585
R9766 gnd.n682 gnd.n681 585
R9767 gnd.n6571 gnd.n6570 585
R9768 gnd.n6572 gnd.n6571 585
R9769 gnd.n680 gnd.n679 585
R9770 gnd.n6573 gnd.n680 585
R9771 gnd.n6576 gnd.n6575 585
R9772 gnd.n6575 gnd.n6574 585
R9773 gnd.n677 gnd.n676 585
R9774 gnd.n676 gnd.n675 585
R9775 gnd.n6581 gnd.n6580 585
R9776 gnd.n6582 gnd.n6581 585
R9777 gnd.n674 gnd.n673 585
R9778 gnd.n6583 gnd.n674 585
R9779 gnd.n6586 gnd.n6585 585
R9780 gnd.n6585 gnd.n6584 585
R9781 gnd.n671 gnd.n670 585
R9782 gnd.n670 gnd.n669 585
R9783 gnd.n6591 gnd.n6590 585
R9784 gnd.n6592 gnd.n6591 585
R9785 gnd.n668 gnd.n667 585
R9786 gnd.n6593 gnd.n668 585
R9787 gnd.n6596 gnd.n6595 585
R9788 gnd.n6595 gnd.n6594 585
R9789 gnd.n665 gnd.n664 585
R9790 gnd.n664 gnd.n663 585
R9791 gnd.n6601 gnd.n6600 585
R9792 gnd.n6602 gnd.n6601 585
R9793 gnd.n662 gnd.n661 585
R9794 gnd.n6603 gnd.n662 585
R9795 gnd.n6606 gnd.n6605 585
R9796 gnd.n6605 gnd.n6604 585
R9797 gnd.n659 gnd.n658 585
R9798 gnd.n658 gnd.n657 585
R9799 gnd.n6611 gnd.n6610 585
R9800 gnd.n6612 gnd.n6611 585
R9801 gnd.n656 gnd.n655 585
R9802 gnd.n6613 gnd.n656 585
R9803 gnd.n6616 gnd.n6615 585
R9804 gnd.n6615 gnd.n6614 585
R9805 gnd.n653 gnd.n652 585
R9806 gnd.n652 gnd.n651 585
R9807 gnd.n6621 gnd.n6620 585
R9808 gnd.n6622 gnd.n6621 585
R9809 gnd.n650 gnd.n649 585
R9810 gnd.n6623 gnd.n650 585
R9811 gnd.n6626 gnd.n6625 585
R9812 gnd.n6625 gnd.n6624 585
R9813 gnd.n647 gnd.n646 585
R9814 gnd.n646 gnd.n645 585
R9815 gnd.n6631 gnd.n6630 585
R9816 gnd.n6632 gnd.n6631 585
R9817 gnd.n644 gnd.n643 585
R9818 gnd.n6633 gnd.n644 585
R9819 gnd.n6636 gnd.n6635 585
R9820 gnd.n6635 gnd.n6634 585
R9821 gnd.n641 gnd.n640 585
R9822 gnd.n640 gnd.n639 585
R9823 gnd.n6641 gnd.n6640 585
R9824 gnd.n6642 gnd.n6641 585
R9825 gnd.n638 gnd.n637 585
R9826 gnd.n6643 gnd.n638 585
R9827 gnd.n6646 gnd.n6645 585
R9828 gnd.n6645 gnd.n6644 585
R9829 gnd.n635 gnd.n634 585
R9830 gnd.n634 gnd.n633 585
R9831 gnd.n6651 gnd.n6650 585
R9832 gnd.n6652 gnd.n6651 585
R9833 gnd.n632 gnd.n631 585
R9834 gnd.n6653 gnd.n632 585
R9835 gnd.n6656 gnd.n6655 585
R9836 gnd.n6655 gnd.n6654 585
R9837 gnd.n629 gnd.n628 585
R9838 gnd.n628 gnd.n627 585
R9839 gnd.n6661 gnd.n6660 585
R9840 gnd.n6662 gnd.n6661 585
R9841 gnd.n626 gnd.n625 585
R9842 gnd.n6663 gnd.n626 585
R9843 gnd.n6666 gnd.n6665 585
R9844 gnd.n6665 gnd.n6664 585
R9845 gnd.n623 gnd.n622 585
R9846 gnd.n622 gnd.n621 585
R9847 gnd.n6671 gnd.n6670 585
R9848 gnd.n6672 gnd.n6671 585
R9849 gnd.n620 gnd.n619 585
R9850 gnd.n6673 gnd.n620 585
R9851 gnd.n6676 gnd.n6675 585
R9852 gnd.n6675 gnd.n6674 585
R9853 gnd.n617 gnd.n616 585
R9854 gnd.n616 gnd.n615 585
R9855 gnd.n6681 gnd.n6680 585
R9856 gnd.n6682 gnd.n6681 585
R9857 gnd.n614 gnd.n613 585
R9858 gnd.n6683 gnd.n614 585
R9859 gnd.n6686 gnd.n6685 585
R9860 gnd.n6685 gnd.n6684 585
R9861 gnd.n611 gnd.n610 585
R9862 gnd.n610 gnd.n609 585
R9863 gnd.n6691 gnd.n6690 585
R9864 gnd.n6692 gnd.n6691 585
R9865 gnd.n608 gnd.n607 585
R9866 gnd.n6693 gnd.n608 585
R9867 gnd.n6696 gnd.n6695 585
R9868 gnd.n6695 gnd.n6694 585
R9869 gnd.n605 gnd.n604 585
R9870 gnd.n604 gnd.n603 585
R9871 gnd.n6701 gnd.n6700 585
R9872 gnd.n6702 gnd.n6701 585
R9873 gnd.n602 gnd.n601 585
R9874 gnd.n6703 gnd.n602 585
R9875 gnd.n6706 gnd.n6705 585
R9876 gnd.n6705 gnd.n6704 585
R9877 gnd.n599 gnd.n598 585
R9878 gnd.n598 gnd.n597 585
R9879 gnd.n6711 gnd.n6710 585
R9880 gnd.n6712 gnd.n6711 585
R9881 gnd.n596 gnd.n595 585
R9882 gnd.n6713 gnd.n596 585
R9883 gnd.n6716 gnd.n6715 585
R9884 gnd.n6715 gnd.n6714 585
R9885 gnd.n593 gnd.n592 585
R9886 gnd.n592 gnd.n591 585
R9887 gnd.n6721 gnd.n6720 585
R9888 gnd.n6722 gnd.n6721 585
R9889 gnd.n590 gnd.n589 585
R9890 gnd.n6723 gnd.n590 585
R9891 gnd.n6726 gnd.n6725 585
R9892 gnd.n6725 gnd.n6724 585
R9893 gnd.n587 gnd.n586 585
R9894 gnd.n586 gnd.n585 585
R9895 gnd.n6731 gnd.n6730 585
R9896 gnd.n6732 gnd.n6731 585
R9897 gnd.n584 gnd.n583 585
R9898 gnd.n6733 gnd.n584 585
R9899 gnd.n6736 gnd.n6735 585
R9900 gnd.n6735 gnd.n6734 585
R9901 gnd.n581 gnd.n580 585
R9902 gnd.n580 gnd.n579 585
R9903 gnd.n6741 gnd.n6740 585
R9904 gnd.n6742 gnd.n6741 585
R9905 gnd.n578 gnd.n577 585
R9906 gnd.n6743 gnd.n578 585
R9907 gnd.n6746 gnd.n6745 585
R9908 gnd.n6745 gnd.n6744 585
R9909 gnd.n575 gnd.n574 585
R9910 gnd.n574 gnd.n573 585
R9911 gnd.n6751 gnd.n6750 585
R9912 gnd.n6752 gnd.n6751 585
R9913 gnd.n572 gnd.n571 585
R9914 gnd.n6753 gnd.n572 585
R9915 gnd.n6756 gnd.n6755 585
R9916 gnd.n6755 gnd.n6754 585
R9917 gnd.n569 gnd.n568 585
R9918 gnd.n568 gnd.n567 585
R9919 gnd.n6761 gnd.n6760 585
R9920 gnd.n6762 gnd.n6761 585
R9921 gnd.n566 gnd.n565 585
R9922 gnd.n6763 gnd.n566 585
R9923 gnd.n6766 gnd.n6765 585
R9924 gnd.n6765 gnd.n6764 585
R9925 gnd.n563 gnd.n562 585
R9926 gnd.n562 gnd.n561 585
R9927 gnd.n6771 gnd.n6770 585
R9928 gnd.n6772 gnd.n6771 585
R9929 gnd.n560 gnd.n559 585
R9930 gnd.n6773 gnd.n560 585
R9931 gnd.n6776 gnd.n6775 585
R9932 gnd.n6775 gnd.n6774 585
R9933 gnd.n557 gnd.n556 585
R9934 gnd.n556 gnd.n555 585
R9935 gnd.n6781 gnd.n6780 585
R9936 gnd.n6782 gnd.n6781 585
R9937 gnd.n554 gnd.n553 585
R9938 gnd.n6783 gnd.n554 585
R9939 gnd.n6786 gnd.n6785 585
R9940 gnd.n6785 gnd.n6784 585
R9941 gnd.n551 gnd.n550 585
R9942 gnd.n550 gnd.n549 585
R9943 gnd.n6791 gnd.n6790 585
R9944 gnd.n6792 gnd.n6791 585
R9945 gnd.n548 gnd.n547 585
R9946 gnd.n6793 gnd.n548 585
R9947 gnd.n6796 gnd.n6795 585
R9948 gnd.n6795 gnd.n6794 585
R9949 gnd.n545 gnd.n544 585
R9950 gnd.n544 gnd.n543 585
R9951 gnd.n6802 gnd.n6801 585
R9952 gnd.n6803 gnd.n6802 585
R9953 gnd.n542 gnd.n541 585
R9954 gnd.n6804 gnd.n542 585
R9955 gnd.n6807 gnd.n6806 585
R9956 gnd.n6806 gnd.n6805 585
R9957 gnd.n6808 gnd.n539 585
R9958 gnd.n539 gnd.n538 585
R9959 gnd.n414 gnd.n413 585
R9960 gnd.n7015 gnd.n413 585
R9961 gnd.n7018 gnd.n7017 585
R9962 gnd.n7017 gnd.n7016 585
R9963 gnd.n417 gnd.n416 585
R9964 gnd.n7014 gnd.n417 585
R9965 gnd.n7012 gnd.n7011 585
R9966 gnd.n7013 gnd.n7012 585
R9967 gnd.n420 gnd.n419 585
R9968 gnd.n419 gnd.n418 585
R9969 gnd.n7007 gnd.n7006 585
R9970 gnd.n7006 gnd.n7005 585
R9971 gnd.n423 gnd.n422 585
R9972 gnd.n7004 gnd.n423 585
R9973 gnd.n7002 gnd.n7001 585
R9974 gnd.n7003 gnd.n7002 585
R9975 gnd.n426 gnd.n425 585
R9976 gnd.n425 gnd.n424 585
R9977 gnd.n6997 gnd.n6996 585
R9978 gnd.n6996 gnd.n6995 585
R9979 gnd.n429 gnd.n428 585
R9980 gnd.n6994 gnd.n429 585
R9981 gnd.n6992 gnd.n6991 585
R9982 gnd.n6993 gnd.n6992 585
R9983 gnd.n432 gnd.n431 585
R9984 gnd.n431 gnd.n430 585
R9985 gnd.n6987 gnd.n6986 585
R9986 gnd.n6986 gnd.n6985 585
R9987 gnd.n435 gnd.n434 585
R9988 gnd.n6984 gnd.n435 585
R9989 gnd.n6982 gnd.n6981 585
R9990 gnd.n6983 gnd.n6982 585
R9991 gnd.n438 gnd.n437 585
R9992 gnd.n437 gnd.n436 585
R9993 gnd.n6977 gnd.n6976 585
R9994 gnd.n6976 gnd.n6975 585
R9995 gnd.n441 gnd.n440 585
R9996 gnd.n6974 gnd.n441 585
R9997 gnd.n6972 gnd.n6971 585
R9998 gnd.n6973 gnd.n6972 585
R9999 gnd.n444 gnd.n443 585
R10000 gnd.n443 gnd.n442 585
R10001 gnd.n6967 gnd.n6966 585
R10002 gnd.n6966 gnd.n6965 585
R10003 gnd.n447 gnd.n446 585
R10004 gnd.n6964 gnd.n447 585
R10005 gnd.n6962 gnd.n6961 585
R10006 gnd.n6963 gnd.n6962 585
R10007 gnd.n450 gnd.n449 585
R10008 gnd.n449 gnd.n448 585
R10009 gnd.n6957 gnd.n6956 585
R10010 gnd.n6956 gnd.n6955 585
R10011 gnd.n453 gnd.n452 585
R10012 gnd.n6954 gnd.n453 585
R10013 gnd.n6952 gnd.n6951 585
R10014 gnd.n6953 gnd.n6952 585
R10015 gnd.n456 gnd.n455 585
R10016 gnd.n455 gnd.n454 585
R10017 gnd.n6947 gnd.n6946 585
R10018 gnd.n6946 gnd.n6945 585
R10019 gnd.n459 gnd.n458 585
R10020 gnd.n6944 gnd.n459 585
R10021 gnd.n6942 gnd.n6941 585
R10022 gnd.n6943 gnd.n6942 585
R10023 gnd.n462 gnd.n461 585
R10024 gnd.n461 gnd.n460 585
R10025 gnd.n6937 gnd.n6936 585
R10026 gnd.n6936 gnd.n6935 585
R10027 gnd.n465 gnd.n464 585
R10028 gnd.n6934 gnd.n465 585
R10029 gnd.n6932 gnd.n6931 585
R10030 gnd.n6933 gnd.n6932 585
R10031 gnd.n468 gnd.n467 585
R10032 gnd.n467 gnd.n466 585
R10033 gnd.n6927 gnd.n6926 585
R10034 gnd.n6926 gnd.n6925 585
R10035 gnd.n471 gnd.n470 585
R10036 gnd.n6924 gnd.n471 585
R10037 gnd.n6922 gnd.n6921 585
R10038 gnd.n6923 gnd.n6922 585
R10039 gnd.n474 gnd.n473 585
R10040 gnd.n473 gnd.n472 585
R10041 gnd.n6917 gnd.n6916 585
R10042 gnd.n6916 gnd.n6915 585
R10043 gnd.n477 gnd.n476 585
R10044 gnd.n6914 gnd.n477 585
R10045 gnd.n6912 gnd.n6911 585
R10046 gnd.n6913 gnd.n6912 585
R10047 gnd.n480 gnd.n479 585
R10048 gnd.n479 gnd.n478 585
R10049 gnd.n6907 gnd.n6906 585
R10050 gnd.n6906 gnd.n6905 585
R10051 gnd.n483 gnd.n482 585
R10052 gnd.n6904 gnd.n483 585
R10053 gnd.n6902 gnd.n6901 585
R10054 gnd.n6903 gnd.n6902 585
R10055 gnd.n486 gnd.n485 585
R10056 gnd.n485 gnd.n484 585
R10057 gnd.n6897 gnd.n6896 585
R10058 gnd.n6896 gnd.n6895 585
R10059 gnd.n489 gnd.n488 585
R10060 gnd.n6894 gnd.n489 585
R10061 gnd.n6892 gnd.n6891 585
R10062 gnd.n6893 gnd.n6892 585
R10063 gnd.n492 gnd.n491 585
R10064 gnd.n491 gnd.n490 585
R10065 gnd.n6887 gnd.n6886 585
R10066 gnd.n6886 gnd.n6885 585
R10067 gnd.n495 gnd.n494 585
R10068 gnd.n6884 gnd.n495 585
R10069 gnd.n6882 gnd.n6881 585
R10070 gnd.n6883 gnd.n6882 585
R10071 gnd.n498 gnd.n497 585
R10072 gnd.n497 gnd.n496 585
R10073 gnd.n6877 gnd.n6876 585
R10074 gnd.n6876 gnd.n6875 585
R10075 gnd.n501 gnd.n500 585
R10076 gnd.n6874 gnd.n501 585
R10077 gnd.n6872 gnd.n6871 585
R10078 gnd.n6873 gnd.n6872 585
R10079 gnd.n504 gnd.n503 585
R10080 gnd.n503 gnd.n502 585
R10081 gnd.n6867 gnd.n6866 585
R10082 gnd.n6866 gnd.n6865 585
R10083 gnd.n507 gnd.n506 585
R10084 gnd.n6864 gnd.n507 585
R10085 gnd.n6862 gnd.n6861 585
R10086 gnd.n6863 gnd.n6862 585
R10087 gnd.n510 gnd.n509 585
R10088 gnd.n509 gnd.n508 585
R10089 gnd.n6857 gnd.n6856 585
R10090 gnd.n6856 gnd.n6855 585
R10091 gnd.n513 gnd.n512 585
R10092 gnd.n6854 gnd.n513 585
R10093 gnd.n6852 gnd.n6851 585
R10094 gnd.n6853 gnd.n6852 585
R10095 gnd.n516 gnd.n515 585
R10096 gnd.n515 gnd.n514 585
R10097 gnd.n6847 gnd.n6846 585
R10098 gnd.n6846 gnd.n6845 585
R10099 gnd.n519 gnd.n518 585
R10100 gnd.n6844 gnd.n519 585
R10101 gnd.n6842 gnd.n6841 585
R10102 gnd.n6843 gnd.n6842 585
R10103 gnd.n522 gnd.n521 585
R10104 gnd.n521 gnd.n520 585
R10105 gnd.n6837 gnd.n6836 585
R10106 gnd.n6836 gnd.n6835 585
R10107 gnd.n525 gnd.n524 585
R10108 gnd.n6834 gnd.n525 585
R10109 gnd.n6832 gnd.n6831 585
R10110 gnd.n6833 gnd.n6832 585
R10111 gnd.n528 gnd.n527 585
R10112 gnd.n527 gnd.n526 585
R10113 gnd.n6827 gnd.n6826 585
R10114 gnd.n6826 gnd.n6825 585
R10115 gnd.n531 gnd.n530 585
R10116 gnd.n6824 gnd.n531 585
R10117 gnd.n6822 gnd.n6821 585
R10118 gnd.n6823 gnd.n6822 585
R10119 gnd.n534 gnd.n533 585
R10120 gnd.n533 gnd.n532 585
R10121 gnd.n6817 gnd.n6816 585
R10122 gnd.n6816 gnd.n6815 585
R10123 gnd.n537 gnd.n536 585
R10124 gnd.n6814 gnd.n537 585
R10125 gnd.n6812 gnd.n6811 585
R10126 gnd.n6813 gnd.n6812 585
R10127 gnd.n6407 gnd.n833 585
R10128 gnd.n6400 gnd.n833 585
R10129 gnd.n6409 gnd.n6408 585
R10130 gnd.n6410 gnd.n6409 585
R10131 gnd.n817 gnd.n816 585
R10132 gnd.n4922 gnd.n817 585
R10133 gnd.n6418 gnd.n6417 585
R10134 gnd.n6417 gnd.n6416 585
R10135 gnd.n6419 gnd.n812 585
R10136 gnd.n4928 gnd.n812 585
R10137 gnd.n6421 gnd.n6420 585
R10138 gnd.n6422 gnd.n6421 585
R10139 gnd.n796 gnd.n795 585
R10140 gnd.n4916 gnd.n796 585
R10141 gnd.n6430 gnd.n6429 585
R10142 gnd.n6429 gnd.n6428 585
R10143 gnd.n6431 gnd.n791 585
R10144 gnd.n4908 gnd.n791 585
R10145 gnd.n6433 gnd.n6432 585
R10146 gnd.n6434 gnd.n6433 585
R10147 gnd.n776 gnd.n775 585
R10148 gnd.n4902 gnd.n776 585
R10149 gnd.n6442 gnd.n6441 585
R10150 gnd.n6441 gnd.n6440 585
R10151 gnd.n6443 gnd.n770 585
R10152 gnd.n4558 gnd.n770 585
R10153 gnd.n6445 gnd.n6444 585
R10154 gnd.n6446 gnd.n6445 585
R10155 gnd.n771 gnd.n769 585
R10156 gnd.n769 gnd.n752 585
R10157 gnd.n4943 gnd.n4942 585
R10158 gnd.n4940 gnd.n2152 585
R10159 gnd.n4950 gnd.n2149 585
R10160 gnd.n4951 gnd.n2147 585
R10161 gnd.n2146 gnd.n2137 585
R10162 gnd.n4958 gnd.n2136 585
R10163 gnd.n4959 gnd.n2135 585
R10164 gnd.n2133 gnd.n2124 585
R10165 gnd.n4966 gnd.n2123 585
R10166 gnd.n4967 gnd.n2121 585
R10167 gnd.n2120 gnd.n2111 585
R10168 gnd.n4974 gnd.n2110 585
R10169 gnd.n4975 gnd.n2109 585
R10170 gnd.n2107 gnd.n2098 585
R10171 gnd.n4982 gnd.n2097 585
R10172 gnd.n4983 gnd.n2095 585
R10173 gnd.n2094 gnd.n2082 585
R10174 gnd.n4990 gnd.n2081 585
R10175 gnd.n4991 gnd.n2080 585
R10176 gnd.n2080 gnd.n852 585
R10177 gnd.n4936 gnd.n842 585
R10178 gnd.n6400 gnd.n842 585
R10179 gnd.n4935 gnd.n831 585
R10180 gnd.n6410 gnd.n831 585
R10181 gnd.n4934 gnd.n2168 585
R10182 gnd.n4922 gnd.n2168 585
R10183 gnd.n2167 gnd.n820 585
R10184 gnd.n6416 gnd.n820 585
R10185 gnd.n4930 gnd.n4929 585
R10186 gnd.n4929 gnd.n4928 585
R10187 gnd.n2170 gnd.n810 585
R10188 gnd.n6422 gnd.n810 585
R10189 gnd.n4915 gnd.n4914 585
R10190 gnd.n4916 gnd.n4915 585
R10191 gnd.n2173 gnd.n799 585
R10192 gnd.n6428 gnd.n799 585
R10193 gnd.n4910 gnd.n4909 585
R10194 gnd.n4909 gnd.n4908 585
R10195 gnd.n2175 gnd.n789 585
R10196 gnd.n6434 gnd.n789 585
R10197 gnd.n4565 gnd.n4564 585
R10198 gnd.n4902 gnd.n4565 585
R10199 gnd.n2178 gnd.n779 585
R10200 gnd.n6440 gnd.n779 585
R10201 gnd.n4560 gnd.n4559 585
R10202 gnd.n4559 gnd.n4558 585
R10203 gnd.n2180 gnd.n767 585
R10204 gnd.n6446 gnd.n767 585
R10205 gnd.n4541 gnd.n4540 585
R10206 gnd.n4540 gnd.n752 585
R10207 gnd.n7644 gnd.n7643 585
R10208 gnd.n7645 gnd.n7644 585
R10209 gnd.n241 gnd.n240 585
R10210 gnd.n250 gnd.n241 585
R10211 gnd.n7653 gnd.n7652 585
R10212 gnd.n7652 gnd.n7651 585
R10213 gnd.n7654 gnd.n236 585
R10214 gnd.n236 gnd.n235 585
R10215 gnd.n7656 gnd.n7655 585
R10216 gnd.n7657 gnd.n7656 585
R10217 gnd.n222 gnd.n221 585
R10218 gnd.n225 gnd.n222 585
R10219 gnd.n7665 gnd.n7664 585
R10220 gnd.n7664 gnd.n7663 585
R10221 gnd.n7666 gnd.n217 585
R10222 gnd.n217 gnd.n216 585
R10223 gnd.n7668 gnd.n7667 585
R10224 gnd.n7669 gnd.n7668 585
R10225 gnd.n203 gnd.n202 585
R10226 gnd.n213 gnd.n203 585
R10227 gnd.n7677 gnd.n7676 585
R10228 gnd.n7676 gnd.n7675 585
R10229 gnd.n7678 gnd.n198 585
R10230 gnd.n198 gnd.n197 585
R10231 gnd.n7680 gnd.n7679 585
R10232 gnd.n7681 gnd.n7680 585
R10233 gnd.n184 gnd.n183 585
R10234 gnd.n187 gnd.n184 585
R10235 gnd.n7689 gnd.n7688 585
R10236 gnd.n7688 gnd.n7687 585
R10237 gnd.n7690 gnd.n179 585
R10238 gnd.n179 gnd.n178 585
R10239 gnd.n7692 gnd.n7691 585
R10240 gnd.n7693 gnd.n7692 585
R10241 gnd.n164 gnd.n163 585
R10242 gnd.n175 gnd.n164 585
R10243 gnd.n7701 gnd.n7700 585
R10244 gnd.n7700 gnd.n7699 585
R10245 gnd.n7702 gnd.n159 585
R10246 gnd.n159 gnd.n158 585
R10247 gnd.n7704 gnd.n7703 585
R10248 gnd.n7705 gnd.n7704 585
R10249 gnd.n145 gnd.n144 585
R10250 gnd.n148 gnd.n145 585
R10251 gnd.n7713 gnd.n7712 585
R10252 gnd.n7712 gnd.n7711 585
R10253 gnd.n7714 gnd.n140 585
R10254 gnd.n140 gnd.n139 585
R10255 gnd.n7716 gnd.n7715 585
R10256 gnd.n7717 gnd.n7716 585
R10257 gnd.n126 gnd.n125 585
R10258 gnd.n136 gnd.n126 585
R10259 gnd.n7725 gnd.n7724 585
R10260 gnd.n7724 gnd.n7723 585
R10261 gnd.n7726 gnd.n120 585
R10262 gnd.n120 gnd.n118 585
R10263 gnd.n7728 gnd.n7727 585
R10264 gnd.n7729 gnd.n7728 585
R10265 gnd.n121 gnd.n119 585
R10266 gnd.n119 gnd.n106 585
R10267 gnd.n7235 gnd.n107 585
R10268 gnd.n7735 gnd.n107 585
R10269 gnd.n7234 gnd.n7233 585
R10270 gnd.n7233 gnd.n7232 585
R10271 gnd.n259 gnd.n258 585
R10272 gnd.n260 gnd.n259 585
R10273 gnd.n7226 gnd.n7225 585
R10274 gnd.n7225 gnd.n7224 585
R10275 gnd.n265 gnd.n264 585
R10276 gnd.n277 gnd.n265 585
R10277 gnd.n7212 gnd.n7211 585
R10278 gnd.n7213 gnd.n7212 585
R10279 gnd.n279 gnd.n278 585
R10280 gnd.n7204 gnd.n278 585
R10281 gnd.n7176 gnd.n7175 585
R10282 gnd.n7175 gnd.n283 585
R10283 gnd.n7177 gnd.n291 585
R10284 gnd.n7191 gnd.n291 585
R10285 gnd.n7178 gnd.n303 585
R10286 gnd.n303 gnd.n301 585
R10287 gnd.n7180 gnd.n7179 585
R10288 gnd.n7181 gnd.n7180 585
R10289 gnd.n304 gnd.n302 585
R10290 gnd.n302 gnd.n298 585
R10291 gnd.n7153 gnd.n312 585
R10292 gnd.n7165 gnd.n312 585
R10293 gnd.n7154 gnd.n322 585
R10294 gnd.n322 gnd.n310 585
R10295 gnd.n7156 gnd.n7155 585
R10296 gnd.n7157 gnd.n7156 585
R10297 gnd.n323 gnd.n321 585
R10298 gnd.n321 gnd.n318 585
R10299 gnd.n7133 gnd.n329 585
R10300 gnd.n7145 gnd.n329 585
R10301 gnd.n7134 gnd.n340 585
R10302 gnd.n340 gnd.n338 585
R10303 gnd.n7136 gnd.n7135 585
R10304 gnd.n7137 gnd.n7136 585
R10305 gnd.n341 gnd.n339 585
R10306 gnd.n7126 gnd.n339 585
R10307 gnd.n7082 gnd.n7081 585
R10308 gnd.n7081 gnd.n7080 585
R10309 gnd.n7083 gnd.n355 585
R10310 gnd.n7097 gnd.n355 585
R10311 gnd.n7084 gnd.n367 585
R10312 gnd.n7074 gnd.n367 585
R10313 gnd.n7086 gnd.n7085 585
R10314 gnd.n7087 gnd.n7086 585
R10315 gnd.n368 gnd.n366 585
R10316 gnd.n7070 gnd.n366 585
R10317 gnd.n7046 gnd.n7045 585
R10318 gnd.n7045 gnd.n7044 585
R10319 gnd.n7047 gnd.n384 585
R10320 gnd.n7061 gnd.n384 585
R10321 gnd.n7048 gnd.n395 585
R10322 gnd.n7038 gnd.n395 585
R10323 gnd.n7050 gnd.n7049 585
R10324 gnd.n7051 gnd.n7050 585
R10325 gnd.n396 gnd.n394 585
R10326 gnd.n5981 gnd.n394 585
R10327 gnd.n5987 gnd.n5986 585
R10328 gnd.n5988 gnd.n5987 585
R10329 gnd.n5950 gnd.n5940 585
R10330 gnd.n6002 gnd.n5940 585
R10331 gnd.n5957 gnd.n5956 585
R10332 gnd.n5956 gnd.n5936 585
R10333 gnd.n5955 gnd.n1149 585
R10334 gnd.n1155 gnd.n1149 585
R10335 gnd.n6011 gnd.n1150 585
R10336 gnd.n6011 gnd.n6010 585
R10337 gnd.n6013 gnd.n6012 585
R10338 gnd.n6091 gnd.n6014 585
R10339 gnd.n6090 gnd.n6015 585
R10340 gnd.n6022 gnd.n6016 585
R10341 gnd.n6083 gnd.n6023 585
R10342 gnd.n6082 gnd.n6024 585
R10343 gnd.n6026 gnd.n6025 585
R10344 gnd.n6075 gnd.n6034 585
R10345 gnd.n6074 gnd.n6035 585
R10346 gnd.n6042 gnd.n6036 585
R10347 gnd.n6067 gnd.n6043 585
R10348 gnd.n6066 gnd.n6044 585
R10349 gnd.n6046 gnd.n6045 585
R10350 gnd.n6059 gnd.n6054 585
R10351 gnd.n6058 gnd.n6055 585
R10352 gnd.n1067 gnd.n1020 585
R10353 gnd.n6221 gnd.n1021 585
R10354 gnd.n6220 gnd.n6217 585
R10355 gnd.n1030 gnd.n1022 585
R10356 gnd.n6215 gnd.n1030 585
R10357 gnd.n7320 gnd.n7319 585
R10358 gnd.n7398 gnd.n7315 585
R10359 gnd.n7400 gnd.n7399 585
R10360 gnd.n7402 gnd.n7313 585
R10361 gnd.n7404 gnd.n7403 585
R10362 gnd.n7405 gnd.n7308 585
R10363 gnd.n7407 gnd.n7406 585
R10364 gnd.n7409 gnd.n7306 585
R10365 gnd.n7411 gnd.n7410 585
R10366 gnd.n7412 gnd.n7301 585
R10367 gnd.n7414 gnd.n7413 585
R10368 gnd.n7416 gnd.n7299 585
R10369 gnd.n7418 gnd.n7417 585
R10370 gnd.n7419 gnd.n7294 585
R10371 gnd.n7421 gnd.n7420 585
R10372 gnd.n7423 gnd.n7292 585
R10373 gnd.n7425 gnd.n7424 585
R10374 gnd.n7426 gnd.n7290 585
R10375 gnd.n7427 gnd.n254 585
R10376 gnd.n254 gnd.n253 585
R10377 gnd.n7394 gnd.n252 585
R10378 gnd.n7645 gnd.n252 585
R10379 gnd.n7393 gnd.n7392 585
R10380 gnd.n7392 gnd.n250 585
R10381 gnd.n7391 gnd.n243 585
R10382 gnd.n7651 gnd.n243 585
R10383 gnd.n7325 gnd.n7324 585
R10384 gnd.n7324 gnd.n235 585
R10385 gnd.n7387 gnd.n234 585
R10386 gnd.n7657 gnd.n234 585
R10387 gnd.n7386 gnd.n7385 585
R10388 gnd.n7385 gnd.n225 585
R10389 gnd.n7384 gnd.n224 585
R10390 gnd.n7663 gnd.n224 585
R10391 gnd.n7328 gnd.n7327 585
R10392 gnd.n7327 gnd.n216 585
R10393 gnd.n7380 gnd.n215 585
R10394 gnd.n7669 gnd.n215 585
R10395 gnd.n7379 gnd.n7378 585
R10396 gnd.n7378 gnd.n213 585
R10397 gnd.n7377 gnd.n205 585
R10398 gnd.n7675 gnd.n205 585
R10399 gnd.n7331 gnd.n7330 585
R10400 gnd.n7330 gnd.n197 585
R10401 gnd.n7373 gnd.n196 585
R10402 gnd.n7681 gnd.n196 585
R10403 gnd.n7372 gnd.n7371 585
R10404 gnd.n7371 gnd.n187 585
R10405 gnd.n7370 gnd.n186 585
R10406 gnd.n7687 gnd.n186 585
R10407 gnd.n7334 gnd.n7333 585
R10408 gnd.n7333 gnd.n178 585
R10409 gnd.n7366 gnd.n177 585
R10410 gnd.n7693 gnd.n177 585
R10411 gnd.n7365 gnd.n7364 585
R10412 gnd.n7364 gnd.n175 585
R10413 gnd.n7363 gnd.n166 585
R10414 gnd.n7699 gnd.n166 585
R10415 gnd.n7337 gnd.n7336 585
R10416 gnd.n7336 gnd.n158 585
R10417 gnd.n7359 gnd.n157 585
R10418 gnd.n7705 gnd.n157 585
R10419 gnd.n7358 gnd.n7357 585
R10420 gnd.n7357 gnd.n148 585
R10421 gnd.n7356 gnd.n147 585
R10422 gnd.n7711 gnd.n147 585
R10423 gnd.n7340 gnd.n7339 585
R10424 gnd.n7339 gnd.n139 585
R10425 gnd.n7352 gnd.n138 585
R10426 gnd.n7717 gnd.n138 585
R10427 gnd.n7351 gnd.n7350 585
R10428 gnd.n7350 gnd.n136 585
R10429 gnd.n7349 gnd.n128 585
R10430 gnd.n7723 gnd.n128 585
R10431 gnd.n7343 gnd.n7342 585
R10432 gnd.n7342 gnd.n118 585
R10433 gnd.n7345 gnd.n117 585
R10434 gnd.n7729 gnd.n117 585
R10435 gnd.n104 gnd.n103 585
R10436 gnd.n106 gnd.n104 585
R10437 gnd.n7737 gnd.n7736 585
R10438 gnd.n7736 gnd.n7735 585
R10439 gnd.n7738 gnd.n102 585
R10440 gnd.n7232 gnd.n102 585
R10441 gnd.n267 gnd.n100 585
R10442 gnd.n267 gnd.n260 585
R10443 gnd.n7197 gnd.n268 585
R10444 gnd.n7224 gnd.n268 585
R10445 gnd.n7198 gnd.n7196 585
R10446 gnd.n7196 gnd.n277 585
R10447 gnd.n286 gnd.n276 585
R10448 gnd.n7213 gnd.n276 585
R10449 gnd.n7203 gnd.n7202 585
R10450 gnd.n7204 gnd.n7203 585
R10451 gnd.n285 gnd.n284 585
R10452 gnd.n284 gnd.n283 585
R10453 gnd.n7193 gnd.n7192 585
R10454 gnd.n7192 gnd.n7191 585
R10455 gnd.n289 gnd.n288 585
R10456 gnd.n301 gnd.n289 585
R10457 gnd.n7109 gnd.n300 585
R10458 gnd.n7181 gnd.n300 585
R10459 gnd.n7112 gnd.n7108 585
R10460 gnd.n7108 gnd.n298 585
R10461 gnd.n7113 gnd.n311 585
R10462 gnd.n7165 gnd.n311 585
R10463 gnd.n7114 gnd.n7107 585
R10464 gnd.n7107 gnd.n310 585
R10465 gnd.n7105 gnd.n320 585
R10466 gnd.n7157 gnd.n320 585
R10467 gnd.n7118 gnd.n7104 585
R10468 gnd.n7104 gnd.n318 585
R10469 gnd.n7119 gnd.n328 585
R10470 gnd.n7145 gnd.n328 585
R10471 gnd.n7120 gnd.n7103 585
R10472 gnd.n7103 gnd.n338 585
R10473 gnd.n348 gnd.n337 585
R10474 gnd.n7137 gnd.n337 585
R10475 gnd.n7125 gnd.n7124 585
R10476 gnd.n7126 gnd.n7125 585
R10477 gnd.n347 gnd.n346 585
R10478 gnd.n7080 gnd.n346 585
R10479 gnd.n7099 gnd.n7098 585
R10480 gnd.n7098 gnd.n7097 585
R10481 gnd.n351 gnd.n350 585
R10482 gnd.n7074 gnd.n351 585
R10483 gnd.n377 gnd.n364 585
R10484 gnd.n7087 gnd.n364 585
R10485 gnd.n7069 gnd.n7068 585
R10486 gnd.n7070 gnd.n7069 585
R10487 gnd.n376 gnd.n375 585
R10488 gnd.n7044 gnd.n375 585
R10489 gnd.n7063 gnd.n7062 585
R10490 gnd.n7062 gnd.n7061 585
R10491 gnd.n380 gnd.n379 585
R10492 gnd.n7038 gnd.n380 585
R10493 gnd.n5965 gnd.n393 585
R10494 gnd.n7051 gnd.n393 585
R10495 gnd.n5980 gnd.n5979 585
R10496 gnd.n5981 gnd.n5980 585
R10497 gnd.n5964 gnd.n5943 585
R10498 gnd.n5988 gnd.n5943 585
R10499 gnd.n5974 gnd.n5938 585
R10500 gnd.n6002 gnd.n5938 585
R10501 gnd.n5973 gnd.n5972 585
R10502 gnd.n5972 gnd.n5936 585
R10503 gnd.n5971 gnd.n5970 585
R10504 gnd.n5971 gnd.n1155 585
R10505 gnd.n5967 gnd.n1154 585
R10506 gnd.n6010 gnd.n1154 585
R10507 gnd.n5804 gnd.n5803 585
R10508 gnd.n5803 gnd.n1219 585
R10509 gnd.n5805 gnd.n1230 585
R10510 gnd.n5683 gnd.n1230 585
R10511 gnd.n5807 gnd.n5806 585
R10512 gnd.n5808 gnd.n5807 585
R10513 gnd.n1231 gnd.n1229 585
R10514 gnd.n5678 gnd.n1229 585
R10515 gnd.n5676 gnd.n5675 585
R10516 gnd.n5677 gnd.n5676 585
R10517 gnd.n5674 gnd.n1310 585
R10518 gnd.n5644 gnd.n1310 585
R10519 gnd.n5673 gnd.n5672 585
R10520 gnd.n5672 gnd.n5671 585
R10521 gnd.n1312 gnd.n1311 585
R10522 gnd.n1313 gnd.n1312 585
R10523 gnd.n5659 gnd.n5658 585
R10524 gnd.n5660 gnd.n5659 585
R10525 gnd.n5657 gnd.n1324 585
R10526 gnd.n1324 gnd.n1321 585
R10527 gnd.n5656 gnd.n5655 585
R10528 gnd.n5655 gnd.n5654 585
R10529 gnd.n1326 gnd.n1325 585
R10530 gnd.n1333 gnd.n1326 585
R10531 gnd.n5639 gnd.n5638 585
R10532 gnd.n5640 gnd.n5639 585
R10533 gnd.n5637 gnd.n1335 585
R10534 gnd.n5633 gnd.n1335 585
R10535 gnd.n5636 gnd.n5635 585
R10536 gnd.n5635 gnd.n5634 585
R10537 gnd.n1337 gnd.n1336 585
R10538 gnd.n1361 gnd.n1337 585
R10539 gnd.n5626 gnd.n5625 585
R10540 gnd.n5627 gnd.n5626 585
R10541 gnd.n5624 gnd.n1342 585
R10542 gnd.n1348 gnd.n1342 585
R10543 gnd.n5623 gnd.n5622 585
R10544 gnd.n5622 gnd.n5621 585
R10545 gnd.n1344 gnd.n1343 585
R10546 gnd.n5566 gnd.n1344 585
R10547 gnd.n5568 gnd.n1383 585
R10548 gnd.n5568 gnd.n5567 585
R10549 gnd.n5570 gnd.n5569 585
R10550 gnd.n5569 gnd.n1369 585
R10551 gnd.n5571 gnd.n1381 585
R10552 gnd.n1381 gnd.n1379 585
R10553 gnd.n5573 gnd.n5572 585
R10554 gnd.n5574 gnd.n5573 585
R10555 gnd.n1382 gnd.n1380 585
R10556 gnd.n5554 gnd.n1380 585
R10557 gnd.n1410 gnd.n1409 585
R10558 gnd.n1409 gnd.n1387 585
R10559 gnd.n5523 gnd.n1411 585
R10560 gnd.n5523 gnd.n5522 585
R10561 gnd.n5524 gnd.n1408 585
R10562 gnd.n5524 gnd.n1395 585
R10563 gnd.n5526 gnd.n5525 585
R10564 gnd.n5525 gnd.n1394 585
R10565 gnd.n5527 gnd.n1406 585
R10566 gnd.n5515 gnd.n1406 585
R10567 gnd.n5529 gnd.n5528 585
R10568 gnd.n5530 gnd.n5529 585
R10569 gnd.n1407 gnd.n1405 585
R10570 gnd.n1405 gnd.n1402 585
R10571 gnd.n5507 gnd.n5506 585
R10572 gnd.n5508 gnd.n5507 585
R10573 gnd.n5505 gnd.n1419 585
R10574 gnd.n1425 gnd.n1419 585
R10575 gnd.n5504 gnd.n5503 585
R10576 gnd.n5503 gnd.n5502 585
R10577 gnd.n1421 gnd.n1420 585
R10578 gnd.n1422 gnd.n1421 585
R10579 gnd.n5491 gnd.n5490 585
R10580 gnd.n5492 gnd.n5491 585
R10581 gnd.n5489 gnd.n1434 585
R10582 gnd.n1434 gnd.n1431 585
R10583 gnd.n5488 gnd.n5487 585
R10584 gnd.n5487 gnd.n5486 585
R10585 gnd.n1436 gnd.n1435 585
R10586 gnd.n5421 gnd.n1436 585
R10587 gnd.n5447 gnd.n5446 585
R10588 gnd.n5447 gnd.n1445 585
R10589 gnd.n5449 gnd.n5448 585
R10590 gnd.n5448 gnd.n1444 585
R10591 gnd.n5450 gnd.n1457 585
R10592 gnd.n5435 gnd.n1457 585
R10593 gnd.n5452 gnd.n5451 585
R10594 gnd.n5453 gnd.n5452 585
R10595 gnd.n5445 gnd.n1456 585
R10596 gnd.n1456 gnd.n1452 585
R10597 gnd.n5444 gnd.n5443 585
R10598 gnd.n5443 gnd.n5442 585
R10599 gnd.n1459 gnd.n1458 585
R10600 gnd.n1466 gnd.n1459 585
R10601 gnd.n5414 gnd.n5413 585
R10602 gnd.n5415 gnd.n5414 585
R10603 gnd.n5412 gnd.n1468 585
R10604 gnd.n1468 gnd.n1465 585
R10605 gnd.n5411 gnd.n5410 585
R10606 gnd.n5410 gnd.n5409 585
R10607 gnd.n1470 gnd.n1469 585
R10608 gnd.n5327 gnd.n1470 585
R10609 gnd.n5396 gnd.n5395 585
R10610 gnd.n5397 gnd.n5396 585
R10611 gnd.n5394 gnd.n1484 585
R10612 gnd.n1484 gnd.n1481 585
R10613 gnd.n5393 gnd.n5392 585
R10614 gnd.n5392 gnd.n5391 585
R10615 gnd.n1486 gnd.n1485 585
R10616 gnd.n5324 gnd.n1486 585
R10617 gnd.n5351 gnd.n5350 585
R10618 gnd.n5351 gnd.n1495 585
R10619 gnd.n5353 gnd.n5352 585
R10620 gnd.n5352 gnd.n1494 585
R10621 gnd.n5354 gnd.n1507 585
R10622 gnd.n5339 gnd.n1507 585
R10623 gnd.n5356 gnd.n5355 585
R10624 gnd.n5357 gnd.n5356 585
R10625 gnd.n5349 gnd.n1506 585
R10626 gnd.n1506 gnd.n1503 585
R10627 gnd.n5348 gnd.n5347 585
R10628 gnd.n5347 gnd.n5346 585
R10629 gnd.n1509 gnd.n1508 585
R10630 gnd.n1510 gnd.n1509 585
R10631 gnd.n5317 gnd.n5316 585
R10632 gnd.n5318 gnd.n5317 585
R10633 gnd.n5315 gnd.n1518 585
R10634 gnd.n5311 gnd.n1518 585
R10635 gnd.n5314 gnd.n5313 585
R10636 gnd.n5313 gnd.n5312 585
R10637 gnd.n1520 gnd.n1519 585
R10638 gnd.n5299 gnd.n1520 585
R10639 gnd.n5289 gnd.n1538 585
R10640 gnd.n1538 gnd.n1530 585
R10641 gnd.n5291 gnd.n5290 585
R10642 gnd.n5292 gnd.n5291 585
R10643 gnd.n5288 gnd.n1537 585
R10644 gnd.n1544 gnd.n1537 585
R10645 gnd.n5287 gnd.n5286 585
R10646 gnd.n5286 gnd.n5285 585
R10647 gnd.n1540 gnd.n1539 585
R10648 gnd.n1541 gnd.n1540 585
R10649 gnd.n5274 gnd.n5273 585
R10650 gnd.n5275 gnd.n5274 585
R10651 gnd.n5272 gnd.n1553 585
R10652 gnd.n5268 gnd.n1553 585
R10653 gnd.n5271 gnd.n5270 585
R10654 gnd.n5270 gnd.n5269 585
R10655 gnd.n1555 gnd.n1554 585
R10656 gnd.n5258 gnd.n1555 585
R10657 gnd.n5244 gnd.n5243 585
R10658 gnd.n5243 gnd.n5242 585
R10659 gnd.n5245 gnd.n1571 585
R10660 gnd.n5241 gnd.n1571 585
R10661 gnd.n5247 gnd.n5246 585
R10662 gnd.n5248 gnd.n5247 585
R10663 gnd.n1572 gnd.n1570 585
R10664 gnd.n5235 gnd.n1570 585
R10665 gnd.n5233 gnd.n5232 585
R10666 gnd.n5234 gnd.n5233 585
R10667 gnd.n5231 gnd.n1577 585
R10668 gnd.n1583 gnd.n1577 585
R10669 gnd.n5230 gnd.n5229 585
R10670 gnd.n5229 gnd.n5228 585
R10671 gnd.n1579 gnd.n1578 585
R10672 gnd.n1580 gnd.n1579 585
R10673 gnd.n5217 gnd.n5216 585
R10674 gnd.n5218 gnd.n5217 585
R10675 gnd.n5215 gnd.n1592 585
R10676 gnd.n1598 gnd.n1592 585
R10677 gnd.n5214 gnd.n5213 585
R10678 gnd.n5213 gnd.n5212 585
R10679 gnd.n1594 gnd.n1593 585
R10680 gnd.n1603 gnd.n1594 585
R10681 gnd.n5198 gnd.n5197 585
R10682 gnd.n5199 gnd.n5198 585
R10683 gnd.n5196 gnd.n1605 585
R10684 gnd.n5192 gnd.n1605 585
R10685 gnd.n5195 gnd.n5194 585
R10686 gnd.n5194 gnd.n5193 585
R10687 gnd.n1607 gnd.n1606 585
R10688 gnd.n1612 gnd.n1607 585
R10689 gnd.n5185 gnd.n5184 585
R10690 gnd.n5186 gnd.n5185 585
R10691 gnd.n5183 gnd.n1615 585
R10692 gnd.n1621 gnd.n1615 585
R10693 gnd.n5182 gnd.n5181 585
R10694 gnd.n5181 gnd.n5180 585
R10695 gnd.n1617 gnd.n1616 585
R10696 gnd.n1630 gnd.n1617 585
R10697 gnd.n5158 gnd.n5157 585
R10698 gnd.n5159 gnd.n5158 585
R10699 gnd.n5155 gnd.n1631 585
R10700 gnd.n5154 gnd.n5153 585
R10701 gnd.n1653 gnd.n1652 585
R10702 gnd.n5151 gnd.n1653 585
R10703 gnd.n1693 gnd.n1692 585
R10704 gnd.n1695 gnd.n1694 585
R10705 gnd.n1697 gnd.n1696 585
R10706 gnd.n1699 gnd.n1698 585
R10707 gnd.n1701 gnd.n1700 585
R10708 gnd.n1703 gnd.n1702 585
R10709 gnd.n1705 gnd.n1704 585
R10710 gnd.n1707 gnd.n1706 585
R10711 gnd.n1709 gnd.n1708 585
R10712 gnd.n1711 gnd.n1710 585
R10713 gnd.n1713 gnd.n1712 585
R10714 gnd.n1715 gnd.n1714 585
R10715 gnd.n1717 gnd.n1716 585
R10716 gnd.n1719 gnd.n1718 585
R10717 gnd.n1721 gnd.n1720 585
R10718 gnd.n1723 gnd.n1722 585
R10719 gnd.n1725 gnd.n1724 585
R10720 gnd.n1727 gnd.n1726 585
R10721 gnd.n1729 gnd.n1728 585
R10722 gnd.n1731 gnd.n1730 585
R10723 gnd.n1733 gnd.n1732 585
R10724 gnd.n1735 gnd.n1734 585
R10725 gnd.n1737 gnd.n1736 585
R10726 gnd.n1739 gnd.n1738 585
R10727 gnd.n1741 gnd.n1740 585
R10728 gnd.n1743 gnd.n1742 585
R10729 gnd.n1745 gnd.n1744 585
R10730 gnd.n1747 gnd.n1746 585
R10731 gnd.n1749 gnd.n1748 585
R10732 gnd.n1955 gnd.n1954 585
R10733 gnd.n1957 gnd.n1956 585
R10734 gnd.n1959 gnd.n1958 585
R10735 gnd.n1961 gnd.n1960 585
R10736 gnd.n1964 gnd.n1963 585
R10737 gnd.n1966 gnd.n1965 585
R10738 gnd.n1968 gnd.n1967 585
R10739 gnd.n1970 gnd.n1969 585
R10740 gnd.n1972 gnd.n1971 585
R10741 gnd.n1974 gnd.n1973 585
R10742 gnd.n1976 gnd.n1975 585
R10743 gnd.n1978 gnd.n1977 585
R10744 gnd.n1980 gnd.n1979 585
R10745 gnd.n1982 gnd.n1981 585
R10746 gnd.n1984 gnd.n1983 585
R10747 gnd.n1986 gnd.n1985 585
R10748 gnd.n1988 gnd.n1987 585
R10749 gnd.n1990 gnd.n1989 585
R10750 gnd.n1992 gnd.n1991 585
R10751 gnd.n1994 gnd.n1993 585
R10752 gnd.n1996 gnd.n1995 585
R10753 gnd.n1998 gnd.n1997 585
R10754 gnd.n2000 gnd.n1999 585
R10755 gnd.n2002 gnd.n2001 585
R10756 gnd.n2004 gnd.n2003 585
R10757 gnd.n2006 gnd.n2005 585
R10758 gnd.n2008 gnd.n2007 585
R10759 gnd.n2010 gnd.n2009 585
R10760 gnd.n2012 gnd.n2011 585
R10761 gnd.n2014 gnd.n2013 585
R10762 gnd.n2016 gnd.n2015 585
R10763 gnd.n2017 gnd.n1686 585
R10764 gnd.n2023 gnd.n2022 585
R10765 gnd.n5687 gnd.n5686 585
R10766 gnd.n5688 gnd.n1304 585
R10767 gnd.n5690 gnd.n5689 585
R10768 gnd.n5692 gnd.n1302 585
R10769 gnd.n5694 gnd.n5693 585
R10770 gnd.n5695 gnd.n1301 585
R10771 gnd.n5697 gnd.n5696 585
R10772 gnd.n5699 gnd.n1299 585
R10773 gnd.n5701 gnd.n5700 585
R10774 gnd.n5702 gnd.n1298 585
R10775 gnd.n5704 gnd.n5703 585
R10776 gnd.n5706 gnd.n1296 585
R10777 gnd.n5708 gnd.n5707 585
R10778 gnd.n5709 gnd.n1295 585
R10779 gnd.n5711 gnd.n5710 585
R10780 gnd.n5713 gnd.n1293 585
R10781 gnd.n5715 gnd.n5714 585
R10782 gnd.n5716 gnd.n1292 585
R10783 gnd.n5718 gnd.n5717 585
R10784 gnd.n5720 gnd.n1290 585
R10785 gnd.n5722 gnd.n5721 585
R10786 gnd.n5723 gnd.n1289 585
R10787 gnd.n5725 gnd.n5724 585
R10788 gnd.n5727 gnd.n1287 585
R10789 gnd.n5729 gnd.n5728 585
R10790 gnd.n5730 gnd.n1286 585
R10791 gnd.n5732 gnd.n5731 585
R10792 gnd.n5734 gnd.n1284 585
R10793 gnd.n5736 gnd.n5735 585
R10794 gnd.n5738 gnd.n1281 585
R10795 gnd.n5740 gnd.n5739 585
R10796 gnd.n5742 gnd.n1280 585
R10797 gnd.n5743 gnd.n1253 585
R10798 gnd.n5746 gnd.n1101 585
R10799 gnd.n5748 gnd.n5747 585
R10800 gnd.n5749 gnd.n1275 585
R10801 gnd.n5751 gnd.n5750 585
R10802 gnd.n5753 gnd.n1273 585
R10803 gnd.n5755 gnd.n5754 585
R10804 gnd.n5756 gnd.n1272 585
R10805 gnd.n5758 gnd.n5757 585
R10806 gnd.n5760 gnd.n1270 585
R10807 gnd.n5762 gnd.n5761 585
R10808 gnd.n5763 gnd.n1269 585
R10809 gnd.n5765 gnd.n5764 585
R10810 gnd.n5767 gnd.n1267 585
R10811 gnd.n5769 gnd.n5768 585
R10812 gnd.n5770 gnd.n1266 585
R10813 gnd.n5772 gnd.n5771 585
R10814 gnd.n5774 gnd.n1264 585
R10815 gnd.n5776 gnd.n5775 585
R10816 gnd.n5777 gnd.n1263 585
R10817 gnd.n5779 gnd.n5778 585
R10818 gnd.n5781 gnd.n1261 585
R10819 gnd.n5783 gnd.n5782 585
R10820 gnd.n5784 gnd.n1260 585
R10821 gnd.n5786 gnd.n5785 585
R10822 gnd.n5788 gnd.n1258 585
R10823 gnd.n5790 gnd.n5789 585
R10824 gnd.n5791 gnd.n1257 585
R10825 gnd.n5793 gnd.n5792 585
R10826 gnd.n5795 gnd.n1255 585
R10827 gnd.n5797 gnd.n5796 585
R10828 gnd.n5798 gnd.n1254 585
R10829 gnd.n5800 gnd.n5799 585
R10830 gnd.n5802 gnd.n1252 585
R10831 gnd.n5685 gnd.n1305 585
R10832 gnd.n5685 gnd.n1219 585
R10833 gnd.n5684 gnd.n5682 585
R10834 gnd.n5684 gnd.n5683 585
R10835 gnd.n5681 gnd.n1227 585
R10836 gnd.n5808 gnd.n1227 585
R10837 gnd.n5680 gnd.n5679 585
R10838 gnd.n5679 gnd.n5678 585
R10839 gnd.n1308 gnd.n1307 585
R10840 gnd.n5677 gnd.n1308 585
R10841 gnd.n5646 gnd.n5645 585
R10842 gnd.n5645 gnd.n5644 585
R10843 gnd.n5647 gnd.n1314 585
R10844 gnd.n5671 gnd.n1314 585
R10845 gnd.n5649 gnd.n5648 585
R10846 gnd.n5648 gnd.n1313 585
R10847 gnd.n5650 gnd.n1323 585
R10848 gnd.n5660 gnd.n1323 585
R10849 gnd.n5651 gnd.n1329 585
R10850 gnd.n1329 gnd.n1321 585
R10851 gnd.n5653 gnd.n5652 585
R10852 gnd.n5654 gnd.n5653 585
R10853 gnd.n5643 gnd.n1328 585
R10854 gnd.n1333 gnd.n1328 585
R10855 gnd.n5642 gnd.n5641 585
R10856 gnd.n5641 gnd.n5640 585
R10857 gnd.n1331 gnd.n1330 585
R10858 gnd.n5633 gnd.n1331 585
R10859 gnd.n5632 gnd.n5631 585
R10860 gnd.n5634 gnd.n5632 585
R10861 gnd.n5630 gnd.n1338 585
R10862 gnd.n1361 gnd.n1338 585
R10863 gnd.n5629 gnd.n5628 585
R10864 gnd.n5628 gnd.n5627 585
R10865 gnd.n1340 gnd.n1339 585
R10866 gnd.n1348 gnd.n1340 585
R10867 gnd.n5563 gnd.n1346 585
R10868 gnd.n5621 gnd.n1346 585
R10869 gnd.n5565 gnd.n5564 585
R10870 gnd.n5566 gnd.n5565 585
R10871 gnd.n5562 gnd.n1384 585
R10872 gnd.n5567 gnd.n1384 585
R10873 gnd.n5561 gnd.n5560 585
R10874 gnd.n5560 gnd.n1369 585
R10875 gnd.n5559 gnd.n5558 585
R10876 gnd.n5559 gnd.n1379 585
R10877 gnd.n5557 gnd.n1377 585
R10878 gnd.n5574 gnd.n1377 585
R10879 gnd.n5556 gnd.n5555 585
R10880 gnd.n5555 gnd.n5554 585
R10881 gnd.n1386 gnd.n1385 585
R10882 gnd.n1387 gnd.n1386 585
R10883 gnd.n5521 gnd.n5520 585
R10884 gnd.n5522 gnd.n5521 585
R10885 gnd.n5519 gnd.n1414 585
R10886 gnd.n1414 gnd.n1395 585
R10887 gnd.n5518 gnd.n5517 585
R10888 gnd.n5517 gnd.n1394 585
R10889 gnd.n5516 gnd.n5513 585
R10890 gnd.n5516 gnd.n5515 585
R10891 gnd.n5512 gnd.n1404 585
R10892 gnd.n5530 gnd.n1404 585
R10893 gnd.n5511 gnd.n5510 585
R10894 gnd.n5510 gnd.n1402 585
R10895 gnd.n5509 gnd.n1415 585
R10896 gnd.n5509 gnd.n5508 585
R10897 gnd.n5423 gnd.n1416 585
R10898 gnd.n1425 gnd.n1416 585
R10899 gnd.n5424 gnd.n1423 585
R10900 gnd.n5502 gnd.n1423 585
R10901 gnd.n5426 gnd.n5425 585
R10902 gnd.n5425 gnd.n1422 585
R10903 gnd.n5427 gnd.n1433 585
R10904 gnd.n5492 gnd.n1433 585
R10905 gnd.n5429 gnd.n5428 585
R10906 gnd.n5428 gnd.n1431 585
R10907 gnd.n5430 gnd.n1437 585
R10908 gnd.n5486 gnd.n1437 585
R10909 gnd.n5431 gnd.n5422 585
R10910 gnd.n5422 gnd.n5421 585
R10911 gnd.n5433 gnd.n5432 585
R10912 gnd.n5433 gnd.n1445 585
R10913 gnd.n5434 gnd.n5419 585
R10914 gnd.n5434 gnd.n1444 585
R10915 gnd.n5437 gnd.n5436 585
R10916 gnd.n5436 gnd.n5435 585
R10917 gnd.n5438 gnd.n1454 585
R10918 gnd.n5453 gnd.n1454 585
R10919 gnd.n5439 gnd.n1462 585
R10920 gnd.n1462 gnd.n1452 585
R10921 gnd.n5441 gnd.n5440 585
R10922 gnd.n5442 gnd.n5441 585
R10923 gnd.n5418 gnd.n1461 585
R10924 gnd.n1466 gnd.n1461 585
R10925 gnd.n5417 gnd.n5416 585
R10926 gnd.n5416 gnd.n5415 585
R10927 gnd.n1464 gnd.n1463 585
R10928 gnd.n1465 gnd.n1464 585
R10929 gnd.n5326 gnd.n1473 585
R10930 gnd.n5409 gnd.n1473 585
R10931 gnd.n5329 gnd.n5328 585
R10932 gnd.n5328 gnd.n5327 585
R10933 gnd.n5330 gnd.n1483 585
R10934 gnd.n5397 gnd.n1483 585
R10935 gnd.n5332 gnd.n5331 585
R10936 gnd.n5331 gnd.n1481 585
R10937 gnd.n5333 gnd.n1487 585
R10938 gnd.n5391 gnd.n1487 585
R10939 gnd.n5334 gnd.n5325 585
R10940 gnd.n5325 gnd.n5324 585
R10941 gnd.n5336 gnd.n5335 585
R10942 gnd.n5336 gnd.n1495 585
R10943 gnd.n5337 gnd.n5322 585
R10944 gnd.n5337 gnd.n1494 585
R10945 gnd.n5341 gnd.n5340 585
R10946 gnd.n5340 gnd.n5339 585
R10947 gnd.n5342 gnd.n1505 585
R10948 gnd.n5357 gnd.n1505 585
R10949 gnd.n5343 gnd.n1513 585
R10950 gnd.n1513 gnd.n1503 585
R10951 gnd.n5345 gnd.n5344 585
R10952 gnd.n5346 gnd.n5345 585
R10953 gnd.n5321 gnd.n1512 585
R10954 gnd.n1512 gnd.n1510 585
R10955 gnd.n5320 gnd.n5319 585
R10956 gnd.n5319 gnd.n5318 585
R10957 gnd.n1515 gnd.n1514 585
R10958 gnd.n5311 gnd.n1515 585
R10959 gnd.n5296 gnd.n1522 585
R10960 gnd.n5312 gnd.n1522 585
R10961 gnd.n5298 gnd.n5297 585
R10962 gnd.n5299 gnd.n5298 585
R10963 gnd.n5295 gnd.n1532 585
R10964 gnd.n1532 gnd.n1530 585
R10965 gnd.n5294 gnd.n5293 585
R10966 gnd.n5293 gnd.n5292 585
R10967 gnd.n1534 gnd.n1533 585
R10968 gnd.n1544 gnd.n1534 585
R10969 gnd.n5262 gnd.n1542 585
R10970 gnd.n5285 gnd.n1542 585
R10971 gnd.n5264 gnd.n5263 585
R10972 gnd.n5263 gnd.n1541 585
R10973 gnd.n5265 gnd.n1551 585
R10974 gnd.n5275 gnd.n1551 585
R10975 gnd.n5267 gnd.n5266 585
R10976 gnd.n5268 gnd.n5267 585
R10977 gnd.n5261 gnd.n1558 585
R10978 gnd.n5269 gnd.n1558 585
R10979 gnd.n5260 gnd.n5259 585
R10980 gnd.n5259 gnd.n5258 585
R10981 gnd.n1560 gnd.n1559 585
R10982 gnd.n5242 gnd.n1560 585
R10983 gnd.n5240 gnd.n5239 585
R10984 gnd.n5241 gnd.n5240 585
R10985 gnd.n5238 gnd.n1568 585
R10986 gnd.n5248 gnd.n1568 585
R10987 gnd.n5237 gnd.n5236 585
R10988 gnd.n5236 gnd.n5235 585
R10989 gnd.n1574 gnd.n1573 585
R10990 gnd.n5234 gnd.n1574 585
R10991 gnd.n5204 gnd.n5203 585
R10992 gnd.n5203 gnd.n1583 585
R10993 gnd.n5205 gnd.n1581 585
R10994 gnd.n5228 gnd.n1581 585
R10995 gnd.n5207 gnd.n5206 585
R10996 gnd.n5206 gnd.n1580 585
R10997 gnd.n5208 gnd.n1590 585
R10998 gnd.n5218 gnd.n1590 585
R10999 gnd.n5209 gnd.n1599 585
R11000 gnd.n1599 gnd.n1598 585
R11001 gnd.n5211 gnd.n5210 585
R11002 gnd.n5212 gnd.n5211 585
R11003 gnd.n5202 gnd.n1597 585
R11004 gnd.n1603 gnd.n1597 585
R11005 gnd.n5201 gnd.n5200 585
R11006 gnd.n5200 gnd.n5199 585
R11007 gnd.n1601 gnd.n1600 585
R11008 gnd.n5192 gnd.n1601 585
R11009 gnd.n5191 gnd.n5190 585
R11010 gnd.n5193 gnd.n5191 585
R11011 gnd.n5189 gnd.n1609 585
R11012 gnd.n1612 gnd.n1609 585
R11013 gnd.n5188 gnd.n5187 585
R11014 gnd.n5187 gnd.n5186 585
R11015 gnd.n1611 gnd.n1610 585
R11016 gnd.n1621 gnd.n1611 585
R11017 gnd.n2018 gnd.n1619 585
R11018 gnd.n5180 gnd.n1619 585
R11019 gnd.n2020 gnd.n2019 585
R11020 gnd.n2019 gnd.n1630 585
R11021 gnd.n2021 gnd.n1629 585
R11022 gnd.n5159 gnd.n1629 585
R11023 gnd.n828 gnd.n827 585
R11024 gnd.n6400 gnd.n828 585
R11025 gnd.n6412 gnd.n6411 585
R11026 gnd.n6411 gnd.n6410 585
R11027 gnd.n6413 gnd.n822 585
R11028 gnd.n4922 gnd.n822 585
R11029 gnd.n6415 gnd.n6414 585
R11030 gnd.n6416 gnd.n6415 585
R11031 gnd.n807 gnd.n806 585
R11032 gnd.n4928 gnd.n807 585
R11033 gnd.n6424 gnd.n6423 585
R11034 gnd.n6423 gnd.n6422 585
R11035 gnd.n6425 gnd.n801 585
R11036 gnd.n4916 gnd.n801 585
R11037 gnd.n6427 gnd.n6426 585
R11038 gnd.n6428 gnd.n6427 585
R11039 gnd.n787 gnd.n786 585
R11040 gnd.n4908 gnd.n787 585
R11041 gnd.n6436 gnd.n6435 585
R11042 gnd.n6435 gnd.n6434 585
R11043 gnd.n6437 gnd.n781 585
R11044 gnd.n4902 gnd.n781 585
R11045 gnd.n6439 gnd.n6438 585
R11046 gnd.n6440 gnd.n6439 585
R11047 gnd.n764 gnd.n763 585
R11048 gnd.n4558 gnd.n764 585
R11049 gnd.n6448 gnd.n6447 585
R11050 gnd.n6447 gnd.n6446 585
R11051 gnd.n6449 gnd.n758 585
R11052 gnd.n758 gnd.n752 585
R11053 gnd.n6403 gnd.n6402 585
R11054 gnd.n1897 gnd.n840 585
R11055 gnd.n1899 gnd.n1898 585
R11056 gnd.n1900 gnd.n1891 585
R11057 gnd.n1902 gnd.n1901 585
R11058 gnd.n1904 gnd.n1889 585
R11059 gnd.n1906 gnd.n1905 585
R11060 gnd.n1907 gnd.n1884 585
R11061 gnd.n1909 gnd.n1908 585
R11062 gnd.n1911 gnd.n1882 585
R11063 gnd.n1913 gnd.n1912 585
R11064 gnd.n1914 gnd.n1877 585
R11065 gnd.n1916 gnd.n1915 585
R11066 gnd.n1918 gnd.n1875 585
R11067 gnd.n1920 gnd.n1919 585
R11068 gnd.n1921 gnd.n1870 585
R11069 gnd.n1923 gnd.n1922 585
R11070 gnd.n1925 gnd.n1869 585
R11071 gnd.n1926 gnd.n1866 585
R11072 gnd.n1929 gnd.n1928 585
R11073 gnd.n1868 gnd.n1862 585
R11074 gnd.n1933 gnd.n1859 585
R11075 gnd.n1935 gnd.n1934 585
R11076 gnd.n1937 gnd.n1857 585
R11077 gnd.n1939 gnd.n1938 585
R11078 gnd.n1940 gnd.n1852 585
R11079 gnd.n1942 gnd.n1941 585
R11080 gnd.n1944 gnd.n1851 585
R11081 gnd.n1945 gnd.n1848 585
R11082 gnd.n1948 gnd.n1947 585
R11083 gnd.n1850 gnd.n1750 585
R11084 gnd.n1842 gnd.n1751 585
R11085 gnd.n1844 gnd.n1843 585
R11086 gnd.n1839 gnd.n1754 585
R11087 gnd.n1838 gnd.n1837 585
R11088 gnd.n1831 gnd.n1756 585
R11089 gnd.n1833 gnd.n1832 585
R11090 gnd.n1829 gnd.n1758 585
R11091 gnd.n1828 gnd.n1827 585
R11092 gnd.n1824 gnd.n1823 585
R11093 gnd.n1822 gnd.n1764 585
R11094 gnd.n1820 gnd.n1819 585
R11095 gnd.n1766 gnd.n1765 585
R11096 gnd.n1815 gnd.n1814 585
R11097 gnd.n1812 gnd.n1768 585
R11098 gnd.n1810 gnd.n1809 585
R11099 gnd.n1770 gnd.n1769 585
R11100 gnd.n1805 gnd.n1804 585
R11101 gnd.n1802 gnd.n1772 585
R11102 gnd.n1800 gnd.n1799 585
R11103 gnd.n1774 gnd.n1773 585
R11104 gnd.n1795 gnd.n1794 585
R11105 gnd.n1792 gnd.n1776 585
R11106 gnd.n1790 gnd.n1789 585
R11107 gnd.n1778 gnd.n1777 585
R11108 gnd.n1785 gnd.n1784 585
R11109 gnd.n1782 gnd.n1781 585
R11110 gnd.n1782 gnd.n852 585
R11111 gnd.n6401 gnd.n835 585
R11112 gnd.n6401 gnd.n6400 585
R11113 gnd.n4921 gnd.n830 585
R11114 gnd.n6410 gnd.n830 585
R11115 gnd.n4924 gnd.n4923 585
R11116 gnd.n4923 gnd.n4922 585
R11117 gnd.n4925 gnd.n819 585
R11118 gnd.n6416 gnd.n819 585
R11119 gnd.n4927 gnd.n4926 585
R11120 gnd.n4928 gnd.n4927 585
R11121 gnd.n4919 gnd.n809 585
R11122 gnd.n6422 gnd.n809 585
R11123 gnd.n4918 gnd.n4917 585
R11124 gnd.n4917 gnd.n4916 585
R11125 gnd.n2171 gnd.n798 585
R11126 gnd.n6428 gnd.n798 585
R11127 gnd.n4907 gnd.n4906 585
R11128 gnd.n4908 gnd.n4907 585
R11129 gnd.n4905 gnd.n788 585
R11130 gnd.n6434 gnd.n788 585
R11131 gnd.n4904 gnd.n4903 585
R11132 gnd.n4903 gnd.n4902 585
R11133 gnd.n2176 gnd.n778 585
R11134 gnd.n6440 gnd.n778 585
R11135 gnd.n4557 gnd.n4556 585
R11136 gnd.n4558 gnd.n4557 585
R11137 gnd.n4555 gnd.n766 585
R11138 gnd.n6446 gnd.n766 585
R11139 gnd.n4554 gnd.n4553 585
R11140 gnd.n4553 gnd.n752 585
R11141 gnd.n7647 gnd.n7646 585
R11142 gnd.n7646 gnd.n7645 585
R11143 gnd.n7648 gnd.n244 585
R11144 gnd.n250 gnd.n244 585
R11145 gnd.n7650 gnd.n7649 585
R11146 gnd.n7651 gnd.n7650 585
R11147 gnd.n232 gnd.n231 585
R11148 gnd.n235 gnd.n232 585
R11149 gnd.n7659 gnd.n7658 585
R11150 gnd.n7658 gnd.n7657 585
R11151 gnd.n7660 gnd.n226 585
R11152 gnd.n226 gnd.n225 585
R11153 gnd.n7662 gnd.n7661 585
R11154 gnd.n7663 gnd.n7662 585
R11155 gnd.n212 gnd.n211 585
R11156 gnd.n216 gnd.n212 585
R11157 gnd.n7671 gnd.n7670 585
R11158 gnd.n7670 gnd.n7669 585
R11159 gnd.n7672 gnd.n206 585
R11160 gnd.n213 gnd.n206 585
R11161 gnd.n7674 gnd.n7673 585
R11162 gnd.n7675 gnd.n7674 585
R11163 gnd.n194 gnd.n193 585
R11164 gnd.n197 gnd.n194 585
R11165 gnd.n7683 gnd.n7682 585
R11166 gnd.n7682 gnd.n7681 585
R11167 gnd.n7684 gnd.n188 585
R11168 gnd.n188 gnd.n187 585
R11169 gnd.n7686 gnd.n7685 585
R11170 gnd.n7687 gnd.n7686 585
R11171 gnd.n174 gnd.n173 585
R11172 gnd.n178 gnd.n174 585
R11173 gnd.n7695 gnd.n7694 585
R11174 gnd.n7694 gnd.n7693 585
R11175 gnd.n7696 gnd.n168 585
R11176 gnd.n175 gnd.n168 585
R11177 gnd.n7698 gnd.n7697 585
R11178 gnd.n7699 gnd.n7698 585
R11179 gnd.n155 gnd.n154 585
R11180 gnd.n158 gnd.n155 585
R11181 gnd.n7707 gnd.n7706 585
R11182 gnd.n7706 gnd.n7705 585
R11183 gnd.n7708 gnd.n149 585
R11184 gnd.n149 gnd.n148 585
R11185 gnd.n7710 gnd.n7709 585
R11186 gnd.n7711 gnd.n7710 585
R11187 gnd.n135 gnd.n134 585
R11188 gnd.n139 gnd.n135 585
R11189 gnd.n7719 gnd.n7718 585
R11190 gnd.n7718 gnd.n7717 585
R11191 gnd.n7720 gnd.n129 585
R11192 gnd.n136 gnd.n129 585
R11193 gnd.n7722 gnd.n7721 585
R11194 gnd.n7723 gnd.n7722 585
R11195 gnd.n115 gnd.n114 585
R11196 gnd.n118 gnd.n115 585
R11197 gnd.n7731 gnd.n7730 585
R11198 gnd.n7730 gnd.n7729 585
R11199 gnd.n7732 gnd.n109 585
R11200 gnd.n109 gnd.n106 585
R11201 gnd.n7734 gnd.n7733 585
R11202 gnd.n7735 gnd.n7734 585
R11203 gnd.n110 gnd.n108 585
R11204 gnd.n7232 gnd.n108 585
R11205 gnd.n7221 gnd.n270 585
R11206 gnd.n270 gnd.n260 585
R11207 gnd.n7223 gnd.n7222 585
R11208 gnd.n7224 gnd.n7223 585
R11209 gnd.n271 gnd.n269 585
R11210 gnd.n277 gnd.n269 585
R11211 gnd.n7215 gnd.n7214 585
R11212 gnd.n7214 gnd.n7213 585
R11213 gnd.n274 gnd.n273 585
R11214 gnd.n7204 gnd.n274 585
R11215 gnd.n7188 gnd.n293 585
R11216 gnd.n293 gnd.n283 585
R11217 gnd.n7190 gnd.n7189 585
R11218 gnd.n7191 gnd.n7190 585
R11219 gnd.n294 gnd.n292 585
R11220 gnd.n301 gnd.n292 585
R11221 gnd.n7183 gnd.n7182 585
R11222 gnd.n7182 gnd.n7181 585
R11223 gnd.n297 gnd.n296 585
R11224 gnd.n298 gnd.n297 585
R11225 gnd.n7164 gnd.n7163 585
R11226 gnd.n7165 gnd.n7164 585
R11227 gnd.n314 gnd.n313 585
R11228 gnd.n313 gnd.n310 585
R11229 gnd.n7159 gnd.n7158 585
R11230 gnd.n7158 gnd.n7157 585
R11231 gnd.n317 gnd.n316 585
R11232 gnd.n318 gnd.n317 585
R11233 gnd.n7144 gnd.n7143 585
R11234 gnd.n7145 gnd.n7144 585
R11235 gnd.n331 gnd.n330 585
R11236 gnd.n338 gnd.n330 585
R11237 gnd.n7139 gnd.n7138 585
R11238 gnd.n7138 gnd.n7137 585
R11239 gnd.n334 gnd.n333 585
R11240 gnd.n7126 gnd.n334 585
R11241 gnd.n7094 gnd.n357 585
R11242 gnd.n7080 gnd.n357 585
R11243 gnd.n7096 gnd.n7095 585
R11244 gnd.n7097 gnd.n7096 585
R11245 gnd.n358 gnd.n356 585
R11246 gnd.n7074 gnd.n356 585
R11247 gnd.n7089 gnd.n7088 585
R11248 gnd.n7088 gnd.n7087 585
R11249 gnd.n361 gnd.n360 585
R11250 gnd.n7070 gnd.n361 585
R11251 gnd.n7058 gnd.n386 585
R11252 gnd.n7044 gnd.n386 585
R11253 gnd.n7060 gnd.n7059 585
R11254 gnd.n7061 gnd.n7060 585
R11255 gnd.n387 gnd.n385 585
R11256 gnd.n7038 gnd.n385 585
R11257 gnd.n7053 gnd.n7052 585
R11258 gnd.n7052 gnd.n7051 585
R11259 gnd.n390 gnd.n389 585
R11260 gnd.n5981 gnd.n390 585
R11261 gnd.n5999 gnd.n5989 585
R11262 gnd.n5989 gnd.n5988 585
R11263 gnd.n6001 gnd.n6000 585
R11264 gnd.n6002 gnd.n6001 585
R11265 gnd.n5990 gnd.n5941 585
R11266 gnd.n5941 gnd.n5936 585
R11267 gnd.n5994 gnd.n5993 585
R11268 gnd.n5993 gnd.n1155 585
R11269 gnd.n5992 gnd.n1072 585
R11270 gnd.n6010 gnd.n1072 585
R11271 gnd.n6213 gnd.n6212 585
R11272 gnd.n6211 gnd.n1071 585
R11273 gnd.n6210 gnd.n1070 585
R11274 gnd.n6215 gnd.n1070 585
R11275 gnd.n6209 gnd.n6208 585
R11276 gnd.n6207 gnd.n6206 585
R11277 gnd.n6205 gnd.n6204 585
R11278 gnd.n6203 gnd.n6202 585
R11279 gnd.n6201 gnd.n6200 585
R11280 gnd.n6199 gnd.n6198 585
R11281 gnd.n6197 gnd.n6196 585
R11282 gnd.n6195 gnd.n6194 585
R11283 gnd.n6193 gnd.n6192 585
R11284 gnd.n6191 gnd.n6190 585
R11285 gnd.n6189 gnd.n6188 585
R11286 gnd.n6187 gnd.n6186 585
R11287 gnd.n6185 gnd.n6184 585
R11288 gnd.n6183 gnd.n6182 585
R11289 gnd.n6181 gnd.n6180 585
R11290 gnd.n6178 gnd.n6177 585
R11291 gnd.n6176 gnd.n6175 585
R11292 gnd.n6174 gnd.n6173 585
R11293 gnd.n6172 gnd.n6171 585
R11294 gnd.n6170 gnd.n6169 585
R11295 gnd.n6168 gnd.n6167 585
R11296 gnd.n6166 gnd.n6165 585
R11297 gnd.n6164 gnd.n6163 585
R11298 gnd.n6161 gnd.n6160 585
R11299 gnd.n6159 gnd.n6158 585
R11300 gnd.n6157 gnd.n6156 585
R11301 gnd.n6155 gnd.n6154 585
R11302 gnd.n6153 gnd.n6152 585
R11303 gnd.n6151 gnd.n6150 585
R11304 gnd.n6149 gnd.n6148 585
R11305 gnd.n6147 gnd.n6146 585
R11306 gnd.n6145 gnd.n6144 585
R11307 gnd.n6143 gnd.n6142 585
R11308 gnd.n6141 gnd.n6140 585
R11309 gnd.n6139 gnd.n6138 585
R11310 gnd.n6137 gnd.n6136 585
R11311 gnd.n6135 gnd.n6134 585
R11312 gnd.n6133 gnd.n6132 585
R11313 gnd.n6131 gnd.n6130 585
R11314 gnd.n6129 gnd.n6128 585
R11315 gnd.n6127 gnd.n6126 585
R11316 gnd.n6125 gnd.n6124 585
R11317 gnd.n6123 gnd.n6122 585
R11318 gnd.n6121 gnd.n6120 585
R11319 gnd.n6119 gnd.n6118 585
R11320 gnd.n6117 gnd.n6116 585
R11321 gnd.n6115 gnd.n6114 585
R11322 gnd.n6113 gnd.n6112 585
R11323 gnd.n6111 gnd.n6110 585
R11324 gnd.n6109 gnd.n6108 585
R11325 gnd.n6107 gnd.n6106 585
R11326 gnd.n6105 gnd.n6104 585
R11327 gnd.n6103 gnd.n6102 585
R11328 gnd.n1152 gnd.n1135 585
R11329 gnd.n7639 gnd.n7638 585
R11330 gnd.n7636 gnd.n7432 585
R11331 gnd.n7635 gnd.n7634 585
R11332 gnd.n7628 gnd.n7434 585
R11333 gnd.n7630 gnd.n7629 585
R11334 gnd.n7626 gnd.n7436 585
R11335 gnd.n7625 gnd.n7624 585
R11336 gnd.n7618 gnd.n7438 585
R11337 gnd.n7620 gnd.n7619 585
R11338 gnd.n7616 gnd.n7440 585
R11339 gnd.n7615 gnd.n7614 585
R11340 gnd.n7608 gnd.n7442 585
R11341 gnd.n7610 gnd.n7609 585
R11342 gnd.n7606 gnd.n7444 585
R11343 gnd.n7605 gnd.n7604 585
R11344 gnd.n7598 gnd.n7446 585
R11345 gnd.n7600 gnd.n7599 585
R11346 gnd.n7596 gnd.n7448 585
R11347 gnd.n7595 gnd.n7594 585
R11348 gnd.n7588 gnd.n7450 585
R11349 gnd.n7590 gnd.n7589 585
R11350 gnd.n7586 gnd.n7454 585
R11351 gnd.n7585 gnd.n7584 585
R11352 gnd.n7578 gnd.n7456 585
R11353 gnd.n7580 gnd.n7579 585
R11354 gnd.n7576 gnd.n7458 585
R11355 gnd.n7575 gnd.n7574 585
R11356 gnd.n7568 gnd.n7460 585
R11357 gnd.n7570 gnd.n7569 585
R11358 gnd.n7566 gnd.n7462 585
R11359 gnd.n7565 gnd.n7564 585
R11360 gnd.n7558 gnd.n7464 585
R11361 gnd.n7560 gnd.n7559 585
R11362 gnd.n7556 gnd.n7466 585
R11363 gnd.n7555 gnd.n7554 585
R11364 gnd.n7548 gnd.n7468 585
R11365 gnd.n7550 gnd.n7549 585
R11366 gnd.n7546 gnd.n7470 585
R11367 gnd.n7545 gnd.n7544 585
R11368 gnd.n7538 gnd.n7472 585
R11369 gnd.n7540 gnd.n7539 585
R11370 gnd.n7536 gnd.n7535 585
R11371 gnd.n7534 gnd.n7477 585
R11372 gnd.n7528 gnd.n7478 585
R11373 gnd.n7530 gnd.n7529 585
R11374 gnd.n7525 gnd.n7480 585
R11375 gnd.n7524 gnd.n7523 585
R11376 gnd.n7517 gnd.n7482 585
R11377 gnd.n7519 gnd.n7518 585
R11378 gnd.n7515 gnd.n7484 585
R11379 gnd.n7514 gnd.n7513 585
R11380 gnd.n7507 gnd.n7486 585
R11381 gnd.n7509 gnd.n7508 585
R11382 gnd.n7505 gnd.n7488 585
R11383 gnd.n7504 gnd.n7503 585
R11384 gnd.n7497 gnd.n7490 585
R11385 gnd.n7499 gnd.n7498 585
R11386 gnd.n7495 gnd.n7494 585
R11387 gnd.n7493 gnd.n249 585
R11388 gnd.n253 gnd.n249 585
R11389 gnd.n7288 gnd.n251 585
R11390 gnd.n7645 gnd.n251 585
R11391 gnd.n7287 gnd.n7286 585
R11392 gnd.n7286 gnd.n250 585
R11393 gnd.n7285 gnd.n242 585
R11394 gnd.n7651 gnd.n242 585
R11395 gnd.n7284 gnd.n7283 585
R11396 gnd.n7283 gnd.n235 585
R11397 gnd.n7282 gnd.n233 585
R11398 gnd.n7657 gnd.n233 585
R11399 gnd.n7281 gnd.n7280 585
R11400 gnd.n7280 gnd.n225 585
R11401 gnd.n7278 gnd.n223 585
R11402 gnd.n7663 gnd.n223 585
R11403 gnd.n7277 gnd.n7276 585
R11404 gnd.n7276 gnd.n216 585
R11405 gnd.n7275 gnd.n214 585
R11406 gnd.n7669 gnd.n214 585
R11407 gnd.n7274 gnd.n7273 585
R11408 gnd.n7273 gnd.n213 585
R11409 gnd.n7271 gnd.n204 585
R11410 gnd.n7675 gnd.n204 585
R11411 gnd.n7270 gnd.n7269 585
R11412 gnd.n7269 gnd.n197 585
R11413 gnd.n7268 gnd.n195 585
R11414 gnd.n7681 gnd.n195 585
R11415 gnd.n7267 gnd.n7266 585
R11416 gnd.n7266 gnd.n187 585
R11417 gnd.n7264 gnd.n185 585
R11418 gnd.n7687 gnd.n185 585
R11419 gnd.n7263 gnd.n7262 585
R11420 gnd.n7262 gnd.n178 585
R11421 gnd.n7261 gnd.n176 585
R11422 gnd.n7693 gnd.n176 585
R11423 gnd.n7260 gnd.n7259 585
R11424 gnd.n7259 gnd.n175 585
R11425 gnd.n7257 gnd.n165 585
R11426 gnd.n7699 gnd.n165 585
R11427 gnd.n7256 gnd.n7255 585
R11428 gnd.n7255 gnd.n158 585
R11429 gnd.n7254 gnd.n156 585
R11430 gnd.n7705 gnd.n156 585
R11431 gnd.n7253 gnd.n7252 585
R11432 gnd.n7252 gnd.n148 585
R11433 gnd.n7250 gnd.n146 585
R11434 gnd.n7711 gnd.n146 585
R11435 gnd.n7249 gnd.n7248 585
R11436 gnd.n7248 gnd.n139 585
R11437 gnd.n7247 gnd.n137 585
R11438 gnd.n7717 gnd.n137 585
R11439 gnd.n7246 gnd.n7245 585
R11440 gnd.n7245 gnd.n136 585
R11441 gnd.n7243 gnd.n127 585
R11442 gnd.n7723 gnd.n127 585
R11443 gnd.n7242 gnd.n7241 585
R11444 gnd.n7241 gnd.n118 585
R11445 gnd.n7240 gnd.n116 585
R11446 gnd.n7729 gnd.n116 585
R11447 gnd.n7239 gnd.n7238 585
R11448 gnd.n7238 gnd.n106 585
R11449 gnd.n256 gnd.n105 585
R11450 gnd.n7735 gnd.n105 585
R11451 gnd.n7231 gnd.n7230 585
R11452 gnd.n7232 gnd.n7231 585
R11453 gnd.n7229 gnd.n261 585
R11454 gnd.n261 gnd.n260 585
R11455 gnd.n266 gnd.n262 585
R11456 gnd.n7224 gnd.n266 585
R11457 gnd.n7208 gnd.n7207 585
R11458 gnd.n7207 gnd.n277 585
R11459 gnd.n7209 gnd.n275 585
R11460 gnd.n7213 gnd.n275 585
R11461 gnd.n7206 gnd.n7205 585
R11462 gnd.n7205 gnd.n7204 585
R11463 gnd.n282 gnd.n281 585
R11464 gnd.n283 gnd.n282 585
R11465 gnd.n7172 gnd.n290 585
R11466 gnd.n7191 gnd.n290 585
R11467 gnd.n7171 gnd.n7170 585
R11468 gnd.n7170 gnd.n301 585
R11469 gnd.n7169 gnd.n299 585
R11470 gnd.n7181 gnd.n299 585
R11471 gnd.n7168 gnd.n7167 585
R11472 gnd.n7167 gnd.n298 585
R11473 gnd.n7166 gnd.n307 585
R11474 gnd.n7166 gnd.n7165 585
R11475 gnd.n7150 gnd.n309 585
R11476 gnd.n310 gnd.n309 585
R11477 gnd.n7149 gnd.n319 585
R11478 gnd.n7157 gnd.n319 585
R11479 gnd.n7148 gnd.n7147 585
R11480 gnd.n7147 gnd.n318 585
R11481 gnd.n7146 gnd.n325 585
R11482 gnd.n7146 gnd.n7145 585
R11483 gnd.n7130 gnd.n327 585
R11484 gnd.n338 gnd.n327 585
R11485 gnd.n7129 gnd.n336 585
R11486 gnd.n7137 gnd.n336 585
R11487 gnd.n7128 gnd.n7127 585
R11488 gnd.n7127 gnd.n7126 585
R11489 gnd.n345 gnd.n343 585
R11490 gnd.n7080 gnd.n345 585
R11491 gnd.n7077 gnd.n353 585
R11492 gnd.n7097 gnd.n353 585
R11493 gnd.n7076 gnd.n7075 585
R11494 gnd.n7075 gnd.n7074 585
R11495 gnd.n7073 gnd.n363 585
R11496 gnd.n7087 gnd.n363 585
R11497 gnd.n7072 gnd.n7071 585
R11498 gnd.n7071 gnd.n7070 585
R11499 gnd.n373 gnd.n371 585
R11500 gnd.n7044 gnd.n373 585
R11501 gnd.n7041 gnd.n382 585
R11502 gnd.n7061 gnd.n382 585
R11503 gnd.n7040 gnd.n7039 585
R11504 gnd.n7039 gnd.n7038 585
R11505 gnd.n399 gnd.n392 585
R11506 gnd.n7051 gnd.n392 585
R11507 gnd.n5983 gnd.n5982 585
R11508 gnd.n5982 gnd.n5981 585
R11509 gnd.n5963 gnd.n5942 585
R11510 gnd.n5988 gnd.n5942 585
R11511 gnd.n5962 gnd.n5937 585
R11512 gnd.n6002 gnd.n5937 585
R11513 gnd.n5961 gnd.n5960 585
R11514 gnd.n5960 gnd.n5936 585
R11515 gnd.n5959 gnd.n5953 585
R11516 gnd.n5959 gnd.n1155 585
R11517 gnd.n5952 gnd.n1153 585
R11518 gnd.n6010 gnd.n1153 585
R11519 gnd.n7024 gnd.n7023 585
R11520 gnd.n7024 gnd.n335 585
R11521 gnd.n7025 gnd.n412 585
R11522 gnd.n7025 gnd.n354 585
R11523 gnd.n7027 gnd.n7026 585
R11524 gnd.n7026 gnd.n352 585
R11525 gnd.n7028 gnd.n407 585
R11526 gnd.n407 gnd.n365 585
R11527 gnd.n7030 gnd.n7029 585
R11528 gnd.n7030 gnd.n362 585
R11529 gnd.n7031 gnd.n406 585
R11530 gnd.n7031 gnd.n374 585
R11531 gnd.n7033 gnd.n7032 585
R11532 gnd.n7032 gnd.n383 585
R11533 gnd.n7034 gnd.n401 585
R11534 gnd.n401 gnd.n381 585
R11535 gnd.n7036 gnd.n7035 585
R11536 gnd.n7037 gnd.n7036 585
R11537 gnd.n402 gnd.n400 585
R11538 gnd.n400 gnd.n391 585
R11539 gnd.n5948 gnd.n5947 585
R11540 gnd.n5949 gnd.n5948 585
R11541 gnd.n5934 gnd.n5933 585
R11542 gnd.n5939 gnd.n5934 585
R11543 gnd.n6005 gnd.n6004 585
R11544 gnd.n6004 gnd.n6003 585
R11545 gnd.n6006 gnd.n1157 585
R11546 gnd.n5935 gnd.n1157 585
R11547 gnd.n6008 gnd.n6007 585
R11548 gnd.n6009 gnd.n6008 585
R11549 gnd.n1158 gnd.n1156 585
R11550 gnd.n1156 gnd.n1151 585
R11551 gnd.n5927 gnd.n5926 585
R11552 gnd.n5926 gnd.n1069 585
R11553 gnd.n5925 gnd.n1160 585
R11554 gnd.n5925 gnd.n1031 585
R11555 gnd.n5924 gnd.n5922 585
R11556 gnd.n5924 gnd.n5923 585
R11557 gnd.n1162 gnd.n1161 585
R11558 gnd.n1161 gnd.n1011 585
R11559 gnd.n5918 gnd.n5917 585
R11560 gnd.n5917 gnd.n997 585
R11561 gnd.n5916 gnd.n1164 585
R11562 gnd.n5916 gnd.n5915 585
R11563 gnd.n5886 gnd.n1165 585
R11564 gnd.n1166 gnd.n1165 585
R11565 gnd.n5888 gnd.n5887 585
R11566 gnd.n5889 gnd.n5888 585
R11567 gnd.n1175 gnd.n1174 585
R11568 gnd.n1174 gnd.n1173 585
R11569 gnd.n5881 gnd.n5880 585
R11570 gnd.n5880 gnd.n5879 585
R11571 gnd.n1178 gnd.n1177 585
R11572 gnd.n1179 gnd.n1178 585
R11573 gnd.n5869 gnd.n5868 585
R11574 gnd.n5870 gnd.n5869 585
R11575 gnd.n1186 gnd.n1185 585
R11576 gnd.n5860 gnd.n1185 585
R11577 gnd.n5864 gnd.n5863 585
R11578 gnd.n5863 gnd.n5862 585
R11579 gnd.n1189 gnd.n1188 585
R11580 gnd.n1190 gnd.n1189 585
R11581 gnd.n5851 gnd.n5850 585
R11582 gnd.n5852 gnd.n5851 585
R11583 gnd.n1198 gnd.n1197 585
R11584 gnd.n1197 gnd.n1196 585
R11585 gnd.n5846 gnd.n5845 585
R11586 gnd.n5845 gnd.n5844 585
R11587 gnd.n1201 gnd.n1200 585
R11588 gnd.n1202 gnd.n1201 585
R11589 gnd.n5834 gnd.n5833 585
R11590 gnd.n5835 gnd.n5834 585
R11591 gnd.n1210 gnd.n1209 585
R11592 gnd.n1209 gnd.n1208 585
R11593 gnd.n5829 gnd.n5828 585
R11594 gnd.n5828 gnd.n5827 585
R11595 gnd.n1213 gnd.n1212 585
R11596 gnd.n1220 gnd.n1213 585
R11597 gnd.n5817 gnd.n5816 585
R11598 gnd.n5818 gnd.n5817 585
R11599 gnd.n1222 gnd.n1221 585
R11600 gnd.n1228 gnd.n1221 585
R11601 gnd.n5812 gnd.n5811 585
R11602 gnd.n5811 gnd.n5810 585
R11603 gnd.n1225 gnd.n1224 585
R11604 gnd.n1309 gnd.n1225 585
R11605 gnd.n5669 gnd.n5668 585
R11606 gnd.n5670 gnd.n5669 585
R11607 gnd.n1317 gnd.n1316 585
R11608 gnd.n5593 gnd.n1316 585
R11609 gnd.n5664 gnd.n5663 585
R11610 gnd.n5663 gnd.n5662 585
R11611 gnd.n1320 gnd.n1319 585
R11612 gnd.n5654 gnd.n1320 585
R11613 gnd.n1359 gnd.n1358 585
R11614 gnd.n1359 gnd.n1334 585
R11615 gnd.n1360 gnd.n1355 585
R11616 gnd.n1360 gnd.n1332 585
R11617 gnd.n5616 gnd.n5615 585
R11618 gnd.n5615 gnd.n5614 585
R11619 gnd.n5617 gnd.n1350 585
R11620 gnd.n1350 gnd.n1341 585
R11621 gnd.n5619 gnd.n5618 585
R11622 gnd.n5620 gnd.n5619 585
R11623 gnd.n1351 gnd.n1349 585
R11624 gnd.n1349 gnd.n1345 585
R11625 gnd.n5583 gnd.n5582 585
R11626 gnd.n5584 gnd.n5583 585
R11627 gnd.n1372 gnd.n1371 585
R11628 gnd.n1378 gnd.n1371 585
R11629 gnd.n5577 gnd.n5576 585
R11630 gnd.n5576 gnd.n5575 585
R11631 gnd.n1375 gnd.n1374 585
R11632 gnd.n5553 gnd.n1375 585
R11633 gnd.n5538 gnd.n1397 585
R11634 gnd.n1413 gnd.n1397 585
R11635 gnd.n5540 gnd.n5539 585
R11636 gnd.n5541 gnd.n5540 585
R11637 gnd.n1398 gnd.n1396 585
R11638 gnd.n5514 gnd.n1396 585
R11639 gnd.n5533 gnd.n5532 585
R11640 gnd.n5532 gnd.n5531 585
R11641 gnd.n1401 gnd.n1400 585
R11642 gnd.n1418 gnd.n1401 585
R11643 gnd.n5500 gnd.n5499 585
R11644 gnd.n5501 gnd.n5500 585
R11645 gnd.n1427 gnd.n1426 585
R11646 gnd.n1426 gnd.n1422 585
R11647 gnd.n5495 gnd.n5494 585
R11648 gnd.n5494 gnd.n5493 585
R11649 gnd.n1430 gnd.n1429 585
R11650 gnd.n5485 gnd.n1430 585
R11651 gnd.n5462 gnd.n1447 585
R11652 gnd.n5420 gnd.n1447 585
R11653 gnd.n5464 gnd.n5463 585
R11654 gnd.n5465 gnd.n5464 585
R11655 gnd.n1448 gnd.n1446 585
R11656 gnd.n1455 gnd.n1446 585
R11657 gnd.n5457 gnd.n5456 585
R11658 gnd.n5456 gnd.n5455 585
R11659 gnd.n1451 gnd.n1450 585
R11660 gnd.n1460 gnd.n1451 585
R11661 gnd.n5405 gnd.n1476 585
R11662 gnd.n1476 gnd.n1467 585
R11663 gnd.n5407 gnd.n5406 585
R11664 gnd.n5408 gnd.n5407 585
R11665 gnd.n1477 gnd.n1475 585
R11666 gnd.n1475 gnd.n1472 585
R11667 gnd.n5400 gnd.n5399 585
R11668 gnd.n5399 gnd.n5398 585
R11669 gnd.n1480 gnd.n1479 585
R11670 gnd.n5390 gnd.n1480 585
R11671 gnd.n5365 gnd.n1498 585
R11672 gnd.n5323 gnd.n1498 585
R11673 gnd.n5367 gnd.n5366 585
R11674 gnd.n5368 gnd.n5367 585
R11675 gnd.n1499 gnd.n1497 585
R11676 gnd.n5338 gnd.n1497 585
R11677 gnd.n5360 gnd.n5359 585
R11678 gnd.n5359 gnd.n5358 585
R11679 gnd.n1502 gnd.n1501 585
R11680 gnd.n5346 gnd.n1502 585
R11681 gnd.n5307 gnd.n1525 585
R11682 gnd.n1525 gnd.n1517 585
R11683 gnd.n5309 gnd.n5308 585
R11684 gnd.n5310 gnd.n5309 585
R11685 gnd.n1526 gnd.n1524 585
R11686 gnd.n1524 gnd.n1521 585
R11687 gnd.n5302 gnd.n5301 585
R11688 gnd.n5301 gnd.n5300 585
R11689 gnd.n1529 gnd.n1528 585
R11690 gnd.n1536 gnd.n1529 585
R11691 gnd.n5283 gnd.n5282 585
R11692 gnd.n5284 gnd.n5283 585
R11693 gnd.n1546 gnd.n1545 585
R11694 gnd.n1552 gnd.n1545 585
R11695 gnd.n5278 gnd.n5277 585
R11696 gnd.n5277 gnd.n5276 585
R11697 gnd.n1549 gnd.n1548 585
R11698 gnd.n1557 gnd.n1549 585
R11699 gnd.n5256 gnd.n5255 585
R11700 gnd.n5257 gnd.n5256 585
R11701 gnd.n1563 gnd.n1562 585
R11702 gnd.n1569 gnd.n1562 585
R11703 gnd.n5251 gnd.n5250 585
R11704 gnd.n5250 gnd.n5249 585
R11705 gnd.n1566 gnd.n1565 585
R11706 gnd.n1576 gnd.n1566 585
R11707 gnd.n5226 gnd.n5225 585
R11708 gnd.n5227 gnd.n5226 585
R11709 gnd.n1585 gnd.n1584 585
R11710 gnd.n1591 gnd.n1584 585
R11711 gnd.n5221 gnd.n5220 585
R11712 gnd.n5220 gnd.n5219 585
R11713 gnd.n1588 gnd.n1587 585
R11714 gnd.n5212 gnd.n1588 585
R11715 gnd.n5172 gnd.n5171 585
R11716 gnd.n5172 gnd.n1604 585
R11717 gnd.n5173 gnd.n5168 585
R11718 gnd.n5173 gnd.n1602 585
R11719 gnd.n5175 gnd.n5174 585
R11720 gnd.n5174 gnd.n1608 585
R11721 gnd.n5176 gnd.n1623 585
R11722 gnd.n1623 gnd.n1614 585
R11723 gnd.n5178 gnd.n5177 585
R11724 gnd.n5179 gnd.n5178 585
R11725 gnd.n1624 gnd.n1622 585
R11726 gnd.n1622 gnd.n1618 585
R11727 gnd.n5162 gnd.n5161 585
R11728 gnd.n5161 gnd.n5160 585
R11729 gnd.n1627 gnd.n1626 585
R11730 gnd.n5150 gnd.n1627 585
R11731 gnd.n5074 gnd.n2033 585
R11732 gnd.n2033 gnd.n1654 585
R11733 gnd.n5076 gnd.n5075 585
R11734 gnd.n5077 gnd.n5076 585
R11735 gnd.n2034 gnd.n2032 585
R11736 gnd.n2032 gnd.n2031 585
R11737 gnd.n5069 gnd.n5068 585
R11738 gnd.n5068 gnd.n5067 585
R11739 gnd.n2037 gnd.n2036 585
R11740 gnd.n2038 gnd.n2037 585
R11741 gnd.n5057 gnd.n5056 585
R11742 gnd.n5058 gnd.n5057 585
R11743 gnd.n2046 gnd.n2045 585
R11744 gnd.n2045 gnd.n2044 585
R11745 gnd.n5052 gnd.n5051 585
R11746 gnd.n5051 gnd.n5050 585
R11747 gnd.n2049 gnd.n2048 585
R11748 gnd.n2050 gnd.n2049 585
R11749 gnd.n5040 gnd.n5039 585
R11750 gnd.n5041 gnd.n5040 585
R11751 gnd.n2057 gnd.n2056 585
R11752 gnd.n5031 gnd.n2056 585
R11753 gnd.n5035 gnd.n5034 585
R11754 gnd.n5034 gnd.n5033 585
R11755 gnd.n2060 gnd.n2059 585
R11756 gnd.n2061 gnd.n2060 585
R11757 gnd.n5022 gnd.n5021 585
R11758 gnd.n5023 gnd.n5022 585
R11759 gnd.n5017 gnd.n5016 585
R11760 gnd.n5016 gnd.n5015 585
R11761 gnd.n860 gnd.n859 585
R11762 gnd.n863 gnd.n860 585
R11763 gnd.n6387 gnd.n6386 585
R11764 gnd.n6386 gnd.n6385 585
R11765 gnd.n6388 gnd.n854 585
R11766 gnd.n861 gnd.n854 585
R11767 gnd.n6390 gnd.n6389 585
R11768 gnd.n6391 gnd.n6390 585
R11769 gnd.n851 gnd.n850 585
R11770 gnd.n6392 gnd.n851 585
R11771 gnd.n6395 gnd.n6394 585
R11772 gnd.n6394 gnd.n6393 585
R11773 gnd.n6396 gnd.n845 585
R11774 gnd.n845 gnd.n843 585
R11775 gnd.n6398 gnd.n6397 585
R11776 gnd.n6399 gnd.n6398 585
R11777 gnd.n846 gnd.n844 585
R11778 gnd.n844 gnd.n832 585
R11779 gnd.n4888 gnd.n4887 585
R11780 gnd.n4888 gnd.n829 585
R11781 gnd.n4889 gnd.n4883 585
R11782 gnd.n4889 gnd.n821 585
R11783 gnd.n4891 gnd.n4890 585
R11784 gnd.n4890 gnd.n818 585
R11785 gnd.n4892 gnd.n4878 585
R11786 gnd.n4878 gnd.n811 585
R11787 gnd.n4894 gnd.n4893 585
R11788 gnd.n4894 gnd.n808 585
R11789 gnd.n4895 gnd.n4877 585
R11790 gnd.n4895 gnd.n800 585
R11791 gnd.n4897 gnd.n4896 585
R11792 gnd.n4896 gnd.n797 585
R11793 gnd.n4898 gnd.n4567 585
R11794 gnd.n4567 gnd.n790 585
R11795 gnd.n4900 gnd.n4899 585
R11796 gnd.n4901 gnd.n4900 585
R11797 gnd.n4568 gnd.n4566 585
R11798 gnd.n4566 gnd.n780 585
R11799 gnd.n4871 gnd.n4870 585
R11800 gnd.n4870 gnd.n777 585
R11801 gnd.n4869 gnd.n4570 585
R11802 gnd.n4869 gnd.n768 585
R11803 gnd.n4868 gnd.n4867 585
R11804 gnd.n4868 gnd.n765 585
R11805 gnd.n5914 gnd.n5913 585
R11806 gnd.n5915 gnd.n5914 585
R11807 gnd.n1169 gnd.n1167 585
R11808 gnd.n1167 gnd.n1166 585
R11809 gnd.n5891 gnd.n5890 585
R11810 gnd.n5890 gnd.n5889 585
R11811 gnd.n1172 gnd.n1171 585
R11812 gnd.n1173 gnd.n1172 585
R11813 gnd.n5877 gnd.n5876 585
R11814 gnd.n5879 gnd.n5877 585
R11815 gnd.n1181 gnd.n1180 585
R11816 gnd.n1180 gnd.n1179 585
R11817 gnd.n5872 gnd.n5871 585
R11818 gnd.n5871 gnd.n5870 585
R11819 gnd.n1184 gnd.n1183 585
R11820 gnd.n5860 gnd.n1184 585
R11821 gnd.n5859 gnd.n5858 585
R11822 gnd.n5862 gnd.n5859 585
R11823 gnd.n1192 gnd.n1191 585
R11824 gnd.n1191 gnd.n1190 585
R11825 gnd.n5854 gnd.n5853 585
R11826 gnd.n5853 gnd.n5852 585
R11827 gnd.n1195 gnd.n1194 585
R11828 gnd.n1196 gnd.n1195 585
R11829 gnd.n5842 gnd.n5841 585
R11830 gnd.n5844 gnd.n5842 585
R11831 gnd.n1204 gnd.n1203 585
R11832 gnd.n1203 gnd.n1202 585
R11833 gnd.n5837 gnd.n5836 585
R11834 gnd.n5836 gnd.n5835 585
R11835 gnd.n1207 gnd.n1206 585
R11836 gnd.n1208 gnd.n1207 585
R11837 gnd.n5825 gnd.n5824 585
R11838 gnd.n5827 gnd.n5825 585
R11839 gnd.n1215 gnd.n1214 585
R11840 gnd.n1220 gnd.n1214 585
R11841 gnd.n5820 gnd.n5819 585
R11842 gnd.n5819 gnd.n5818 585
R11843 gnd.n1218 gnd.n1217 585
R11844 gnd.n1228 gnd.n1218 585
R11845 gnd.n5599 gnd.n1226 585
R11846 gnd.n5810 gnd.n1226 585
R11847 gnd.n5600 gnd.n5597 585
R11848 gnd.n5597 gnd.n1309 585
R11849 gnd.n5601 gnd.n1315 585
R11850 gnd.n5670 gnd.n1315 585
R11851 gnd.n5595 gnd.n5594 585
R11852 gnd.n5594 gnd.n5593 585
R11853 gnd.n5605 gnd.n1322 585
R11854 gnd.n5662 gnd.n1322 585
R11855 gnd.n5606 gnd.n1327 585
R11856 gnd.n5654 gnd.n1327 585
R11857 gnd.n5607 gnd.n5592 585
R11858 gnd.n5592 gnd.n1334 585
R11859 gnd.n1365 gnd.n1363 585
R11860 gnd.n1363 gnd.n1332 585
R11861 gnd.n5612 gnd.n5611 585
R11862 gnd.n5614 gnd.n5612 585
R11863 gnd.n1364 gnd.n1362 585
R11864 gnd.n1362 gnd.n1341 585
R11865 gnd.n5588 gnd.n1347 585
R11866 gnd.n5620 gnd.n1347 585
R11867 gnd.n5587 gnd.n5586 585
R11868 gnd.n5586 gnd.n1345 585
R11869 gnd.n5585 gnd.n1367 585
R11870 gnd.n5585 gnd.n5584 585
R11871 gnd.n5547 gnd.n1368 585
R11872 gnd.n1378 gnd.n1368 585
R11873 gnd.n1390 gnd.n1376 585
R11874 gnd.n5575 gnd.n1376 585
R11875 gnd.n5552 gnd.n5551 585
R11876 gnd.n5553 gnd.n5552 585
R11877 gnd.n1389 gnd.n1388 585
R11878 gnd.n1413 gnd.n1388 585
R11879 gnd.n5543 gnd.n5542 585
R11880 gnd.n5542 gnd.n5541 585
R11881 gnd.n1393 gnd.n1392 585
R11882 gnd.n5514 gnd.n1393 585
R11883 gnd.n5473 gnd.n1403 585
R11884 gnd.n5531 gnd.n1403 585
R11885 gnd.n5476 gnd.n5472 585
R11886 gnd.n5472 gnd.n1418 585
R11887 gnd.n5477 gnd.n1424 585
R11888 gnd.n5501 gnd.n1424 585
R11889 gnd.n5478 gnd.n5471 585
R11890 gnd.n5471 gnd.n1422 585
R11891 gnd.n1440 gnd.n1432 585
R11892 gnd.n5493 gnd.n1432 585
R11893 gnd.n5483 gnd.n5482 585
R11894 gnd.n5485 gnd.n5483 585
R11895 gnd.n1439 gnd.n1438 585
R11896 gnd.n5420 gnd.n1438 585
R11897 gnd.n5467 gnd.n5466 585
R11898 gnd.n5466 gnd.n5465 585
R11899 gnd.n1443 gnd.n1442 585
R11900 gnd.n1455 gnd.n1443 585
R11901 gnd.n5378 gnd.n1453 585
R11902 gnd.n5455 gnd.n1453 585
R11903 gnd.n5377 gnd.n5376 585
R11904 gnd.n5376 gnd.n1460 585
R11905 gnd.n5382 gnd.n5375 585
R11906 gnd.n5375 gnd.n1467 585
R11907 gnd.n5383 gnd.n1474 585
R11908 gnd.n5408 gnd.n1474 585
R11909 gnd.n5384 gnd.n5374 585
R11910 gnd.n5374 gnd.n1472 585
R11911 gnd.n1490 gnd.n1482 585
R11912 gnd.n5398 gnd.n1482 585
R11913 gnd.n5389 gnd.n5388 585
R11914 gnd.n5390 gnd.n5389 585
R11915 gnd.n1489 gnd.n1488 585
R11916 gnd.n5323 gnd.n1488 585
R11917 gnd.n5370 gnd.n5369 585
R11918 gnd.n5369 gnd.n5368 585
R11919 gnd.n1493 gnd.n1492 585
R11920 gnd.n5338 gnd.n1493 585
R11921 gnd.n5107 gnd.n1504 585
R11922 gnd.n5358 gnd.n1504 585
R11923 gnd.n5106 gnd.n1511 585
R11924 gnd.n5346 gnd.n1511 585
R11925 gnd.n5111 gnd.n5105 585
R11926 gnd.n5105 gnd.n1517 585
R11927 gnd.n5112 gnd.n1523 585
R11928 gnd.n5310 gnd.n1523 585
R11929 gnd.n5113 gnd.n5104 585
R11930 gnd.n5104 gnd.n1521 585
R11931 gnd.n5102 gnd.n1531 585
R11932 gnd.n5300 gnd.n1531 585
R11933 gnd.n5117 gnd.n5101 585
R11934 gnd.n5101 gnd.n1536 585
R11935 gnd.n5118 gnd.n1543 585
R11936 gnd.n5284 gnd.n1543 585
R11937 gnd.n5119 gnd.n5100 585
R11938 gnd.n5100 gnd.n1552 585
R11939 gnd.n5098 gnd.n1550 585
R11940 gnd.n5276 gnd.n1550 585
R11941 gnd.n5123 gnd.n5097 585
R11942 gnd.n5097 gnd.n1557 585
R11943 gnd.n5124 gnd.n1561 585
R11944 gnd.n5257 gnd.n1561 585
R11945 gnd.n5125 gnd.n5096 585
R11946 gnd.n5096 gnd.n1569 585
R11947 gnd.n5094 gnd.n1567 585
R11948 gnd.n5249 gnd.n1567 585
R11949 gnd.n5129 gnd.n5093 585
R11950 gnd.n5093 gnd.n1576 585
R11951 gnd.n5130 gnd.n1582 585
R11952 gnd.n5227 gnd.n1582 585
R11953 gnd.n5131 gnd.n5092 585
R11954 gnd.n5092 gnd.n1591 585
R11955 gnd.n5090 gnd.n1589 585
R11956 gnd.n5219 gnd.n1589 585
R11957 gnd.n5135 gnd.n1595 585
R11958 gnd.n5212 gnd.n1595 585
R11959 gnd.n5136 gnd.n5089 585
R11960 gnd.n5089 gnd.n1604 585
R11961 gnd.n5137 gnd.n5088 585
R11962 gnd.n5088 gnd.n1602 585
R11963 gnd.n5087 gnd.n5085 585
R11964 gnd.n5087 gnd.n1608 585
R11965 gnd.n5141 gnd.n5084 585
R11966 gnd.n5084 gnd.n1614 585
R11967 gnd.n5142 gnd.n1620 585
R11968 gnd.n5179 gnd.n1620 585
R11969 gnd.n5143 gnd.n5083 585
R11970 gnd.n5083 gnd.n1618 585
R11971 gnd.n2027 gnd.n1628 585
R11972 gnd.n5160 gnd.n1628 585
R11973 gnd.n5148 gnd.n5147 585
R11974 gnd.n5150 gnd.n5148 585
R11975 gnd.n2026 gnd.n2025 585
R11976 gnd.n2025 gnd.n1654 585
R11977 gnd.n5079 gnd.n5078 585
R11978 gnd.n5078 gnd.n5077 585
R11979 gnd.n2030 gnd.n2029 585
R11980 gnd.n2031 gnd.n2030 585
R11981 gnd.n5065 gnd.n5064 585
R11982 gnd.n5067 gnd.n5065 585
R11983 gnd.n2040 gnd.n2039 585
R11984 gnd.n2039 gnd.n2038 585
R11985 gnd.n5060 gnd.n5059 585
R11986 gnd.n5059 gnd.n5058 585
R11987 gnd.n2043 gnd.n2042 585
R11988 gnd.n2044 gnd.n2043 585
R11989 gnd.n5048 gnd.n5047 585
R11990 gnd.n5050 gnd.n5048 585
R11991 gnd.n2052 gnd.n2051 585
R11992 gnd.n2051 gnd.n2050 585
R11993 gnd.n5043 gnd.n5042 585
R11994 gnd.n5042 gnd.n5041 585
R11995 gnd.n2055 gnd.n2054 585
R11996 gnd.n5031 gnd.n2055 585
R11997 gnd.n5030 gnd.n5029 585
R11998 gnd.n5033 gnd.n5030 585
R11999 gnd.n2063 gnd.n2062 585
R12000 gnd.n2062 gnd.n2061 585
R12001 gnd.n5025 gnd.n5024 585
R12002 gnd.n5024 gnd.n5023 585
R12003 gnd.n5014 gnd.n2065 585
R12004 gnd.n5015 gnd.n5014 585
R12005 gnd.n5013 gnd.n5012 585
R12006 gnd.n5013 gnd.n863 585
R12007 gnd.n2066 gnd.n862 585
R12008 gnd.n6385 gnd.n862 585
R12009 gnd.n5008 gnd.n5007 585
R12010 gnd.n5005 gnd.n2068 585
R12011 gnd.n5004 gnd.n5003 585
R12012 gnd.n5004 gnd.n853 585
R12013 gnd.n2070 gnd.n2069 585
R12014 gnd.n4999 gnd.n2073 585
R12015 gnd.n4998 gnd.n2074 585
R12016 gnd.n4997 gnd.n2076 585
R12017 gnd.n4995 gnd.n2077 585
R12018 gnd.n2086 gnd.n2078 585
R12019 gnd.n2087 gnd.n2084 585
R12020 gnd.n4987 gnd.n2089 585
R12021 gnd.n4986 gnd.n2090 585
R12022 gnd.n2101 gnd.n2091 585
R12023 gnd.n4979 gnd.n2102 585
R12024 gnd.n4978 gnd.n2104 585
R12025 gnd.n2113 gnd.n2105 585
R12026 gnd.n4971 gnd.n2115 585
R12027 gnd.n4970 gnd.n2116 585
R12028 gnd.n2127 gnd.n2117 585
R12029 gnd.n4963 gnd.n2128 585
R12030 gnd.n4962 gnd.n2130 585
R12031 gnd.n2139 gnd.n2131 585
R12032 gnd.n4955 gnd.n2141 585
R12033 gnd.n4954 gnd.n2142 585
R12034 gnd.n2158 gnd.n2143 585
R12035 gnd.n4947 gnd.n2159 585
R12036 gnd.n4946 gnd.n2161 585
R12037 gnd.n2165 gnd.n2163 585
R12038 gnd.n2164 gnd.n864 585
R12039 gnd.n995 gnd.n992 585
R12040 gnd.n5915 gnd.n995 585
R12041 gnd.n6233 gnd.n991 585
R12042 gnd.n1166 gnd.n991 585
R12043 gnd.n6234 gnd.n990 585
R12044 gnd.n5889 gnd.n990 585
R12045 gnd.n6235 gnd.n989 585
R12046 gnd.n1173 gnd.n989 585
R12047 gnd.n5878 gnd.n987 585
R12048 gnd.n5879 gnd.n5878 585
R12049 gnd.n6239 gnd.n986 585
R12050 gnd.n1179 gnd.n986 585
R12051 gnd.n6240 gnd.n985 585
R12052 gnd.n5870 gnd.n985 585
R12053 gnd.n6241 gnd.n984 585
R12054 gnd.n5860 gnd.n984 585
R12055 gnd.n5861 gnd.n982 585
R12056 gnd.n5862 gnd.n5861 585
R12057 gnd.n6245 gnd.n981 585
R12058 gnd.n1190 gnd.n981 585
R12059 gnd.n6246 gnd.n980 585
R12060 gnd.n5852 gnd.n980 585
R12061 gnd.n6247 gnd.n979 585
R12062 gnd.n1196 gnd.n979 585
R12063 gnd.n5843 gnd.n977 585
R12064 gnd.n5844 gnd.n5843 585
R12065 gnd.n6251 gnd.n976 585
R12066 gnd.n1202 gnd.n976 585
R12067 gnd.n6252 gnd.n975 585
R12068 gnd.n5835 gnd.n975 585
R12069 gnd.n6253 gnd.n974 585
R12070 gnd.n1208 gnd.n974 585
R12071 gnd.n5826 gnd.n972 585
R12072 gnd.n5827 gnd.n5826 585
R12073 gnd.n6257 gnd.n971 585
R12074 gnd.n1220 gnd.n971 585
R12075 gnd.n6258 gnd.n970 585
R12076 gnd.n5818 gnd.n970 585
R12077 gnd.n6259 gnd.n969 585
R12078 gnd.n1228 gnd.n969 585
R12079 gnd.n5809 gnd.n967 585
R12080 gnd.n5810 gnd.n5809 585
R12081 gnd.n6263 gnd.n966 585
R12082 gnd.n1309 gnd.n966 585
R12083 gnd.n6264 gnd.n965 585
R12084 gnd.n5670 gnd.n965 585
R12085 gnd.n6265 gnd.n964 585
R12086 gnd.n5593 gnd.n964 585
R12087 gnd.n5661 gnd.n962 585
R12088 gnd.n5662 gnd.n5661 585
R12089 gnd.n6269 gnd.n961 585
R12090 gnd.n5654 gnd.n961 585
R12091 gnd.n6270 gnd.n960 585
R12092 gnd.n1334 gnd.n960 585
R12093 gnd.n6271 gnd.n959 585
R12094 gnd.n1332 gnd.n959 585
R12095 gnd.n5613 gnd.n957 585
R12096 gnd.n5614 gnd.n5613 585
R12097 gnd.n6275 gnd.n956 585
R12098 gnd.n1341 gnd.n956 585
R12099 gnd.n6276 gnd.n955 585
R12100 gnd.n5620 gnd.n955 585
R12101 gnd.n6277 gnd.n954 585
R12102 gnd.n1345 gnd.n954 585
R12103 gnd.n1370 gnd.n952 585
R12104 gnd.n5584 gnd.n1370 585
R12105 gnd.n6281 gnd.n951 585
R12106 gnd.n1378 gnd.n951 585
R12107 gnd.n6282 gnd.n950 585
R12108 gnd.n5575 gnd.n950 585
R12109 gnd.n6283 gnd.n949 585
R12110 gnd.n5553 gnd.n949 585
R12111 gnd.n1412 gnd.n947 585
R12112 gnd.n1413 gnd.n1412 585
R12113 gnd.n6287 gnd.n946 585
R12114 gnd.n5541 gnd.n946 585
R12115 gnd.n6288 gnd.n945 585
R12116 gnd.n5514 gnd.n945 585
R12117 gnd.n6289 gnd.n944 585
R12118 gnd.n5531 gnd.n944 585
R12119 gnd.n1417 gnd.n942 585
R12120 gnd.n1418 gnd.n1417 585
R12121 gnd.n6293 gnd.n941 585
R12122 gnd.n5501 gnd.n941 585
R12123 gnd.n6294 gnd.n940 585
R12124 gnd.n1422 gnd.n940 585
R12125 gnd.n6295 gnd.n939 585
R12126 gnd.n5493 gnd.n939 585
R12127 gnd.n5484 gnd.n937 585
R12128 gnd.n5485 gnd.n5484 585
R12129 gnd.n6299 gnd.n936 585
R12130 gnd.n5420 gnd.n936 585
R12131 gnd.n6300 gnd.n935 585
R12132 gnd.n5465 gnd.n935 585
R12133 gnd.n6301 gnd.n934 585
R12134 gnd.n1455 gnd.n934 585
R12135 gnd.n5454 gnd.n932 585
R12136 gnd.n5455 gnd.n5454 585
R12137 gnd.n6305 gnd.n931 585
R12138 gnd.n1460 gnd.n931 585
R12139 gnd.n6306 gnd.n930 585
R12140 gnd.n1467 gnd.n930 585
R12141 gnd.n6307 gnd.n929 585
R12142 gnd.n5408 gnd.n929 585
R12143 gnd.n1471 gnd.n927 585
R12144 gnd.n1472 gnd.n1471 585
R12145 gnd.n6311 gnd.n926 585
R12146 gnd.n5398 gnd.n926 585
R12147 gnd.n6312 gnd.n925 585
R12148 gnd.n5390 gnd.n925 585
R12149 gnd.n6313 gnd.n924 585
R12150 gnd.n5323 gnd.n924 585
R12151 gnd.n1496 gnd.n922 585
R12152 gnd.n5368 gnd.n1496 585
R12153 gnd.n6317 gnd.n921 585
R12154 gnd.n5338 gnd.n921 585
R12155 gnd.n6318 gnd.n920 585
R12156 gnd.n5358 gnd.n920 585
R12157 gnd.n6319 gnd.n919 585
R12158 gnd.n5346 gnd.n919 585
R12159 gnd.n1516 gnd.n917 585
R12160 gnd.n1517 gnd.n1516 585
R12161 gnd.n6323 gnd.n916 585
R12162 gnd.n5310 gnd.n916 585
R12163 gnd.n6324 gnd.n915 585
R12164 gnd.n1521 gnd.n915 585
R12165 gnd.n6325 gnd.n914 585
R12166 gnd.n5300 gnd.n914 585
R12167 gnd.n1535 gnd.n912 585
R12168 gnd.n1536 gnd.n1535 585
R12169 gnd.n6329 gnd.n911 585
R12170 gnd.n5284 gnd.n911 585
R12171 gnd.n6330 gnd.n910 585
R12172 gnd.n1552 gnd.n910 585
R12173 gnd.n6331 gnd.n909 585
R12174 gnd.n5276 gnd.n909 585
R12175 gnd.n1556 gnd.n907 585
R12176 gnd.n1557 gnd.n1556 585
R12177 gnd.n6335 gnd.n906 585
R12178 gnd.n5257 gnd.n906 585
R12179 gnd.n6336 gnd.n905 585
R12180 gnd.n1569 gnd.n905 585
R12181 gnd.n6337 gnd.n904 585
R12182 gnd.n5249 gnd.n904 585
R12183 gnd.n1575 gnd.n902 585
R12184 gnd.n1576 gnd.n1575 585
R12185 gnd.n6341 gnd.n901 585
R12186 gnd.n5227 gnd.n901 585
R12187 gnd.n6342 gnd.n900 585
R12188 gnd.n1591 gnd.n900 585
R12189 gnd.n6343 gnd.n899 585
R12190 gnd.n5219 gnd.n899 585
R12191 gnd.n1596 gnd.n897 585
R12192 gnd.n5212 gnd.n1596 585
R12193 gnd.n6347 gnd.n896 585
R12194 gnd.n1604 gnd.n896 585
R12195 gnd.n6348 gnd.n895 585
R12196 gnd.n1602 gnd.n895 585
R12197 gnd.n6349 gnd.n894 585
R12198 gnd.n1608 gnd.n894 585
R12199 gnd.n1613 gnd.n892 585
R12200 gnd.n1614 gnd.n1613 585
R12201 gnd.n6353 gnd.n891 585
R12202 gnd.n5179 gnd.n891 585
R12203 gnd.n6354 gnd.n890 585
R12204 gnd.n1618 gnd.n890 585
R12205 gnd.n6355 gnd.n889 585
R12206 gnd.n5160 gnd.n889 585
R12207 gnd.n5149 gnd.n887 585
R12208 gnd.n5150 gnd.n5149 585
R12209 gnd.n6359 gnd.n886 585
R12210 gnd.n1654 gnd.n886 585
R12211 gnd.n6360 gnd.n885 585
R12212 gnd.n5077 gnd.n885 585
R12213 gnd.n6361 gnd.n884 585
R12214 gnd.n2031 gnd.n884 585
R12215 gnd.n5066 gnd.n882 585
R12216 gnd.n5067 gnd.n5066 585
R12217 gnd.n6365 gnd.n881 585
R12218 gnd.n2038 gnd.n881 585
R12219 gnd.n6366 gnd.n880 585
R12220 gnd.n5058 gnd.n880 585
R12221 gnd.n6367 gnd.n879 585
R12222 gnd.n2044 gnd.n879 585
R12223 gnd.n5049 gnd.n877 585
R12224 gnd.n5050 gnd.n5049 585
R12225 gnd.n6371 gnd.n876 585
R12226 gnd.n2050 gnd.n876 585
R12227 gnd.n6372 gnd.n875 585
R12228 gnd.n5041 gnd.n875 585
R12229 gnd.n6373 gnd.n874 585
R12230 gnd.n5031 gnd.n874 585
R12231 gnd.n5032 gnd.n872 585
R12232 gnd.n5033 gnd.n5032 585
R12233 gnd.n6377 gnd.n871 585
R12234 gnd.n2061 gnd.n871 585
R12235 gnd.n6378 gnd.n870 585
R12236 gnd.n5023 gnd.n870 585
R12237 gnd.n6379 gnd.n869 585
R12238 gnd.n5015 gnd.n869 585
R12239 gnd.n866 gnd.n865 585
R12240 gnd.n865 gnd.n863 585
R12241 gnd.n6384 gnd.n6383 585
R12242 gnd.n6385 gnd.n6384 585
R12243 gnd.n6225 gnd.n6224 585
R12244 gnd.n6226 gnd.n6225 585
R12245 gnd.n1014 gnd.n1012 585
R12246 gnd.n6052 gnd.n6051 585
R12247 gnd.n6062 gnd.n6050 585
R12248 gnd.n6063 gnd.n6049 585
R12249 gnd.n6048 gnd.n6040 585
R12250 gnd.n6070 gnd.n6039 585
R12251 gnd.n6071 gnd.n6038 585
R12252 gnd.n6032 gnd.n6031 585
R12253 gnd.n6078 gnd.n6030 585
R12254 gnd.n6079 gnd.n6029 585
R12255 gnd.n6028 gnd.n6020 585
R12256 gnd.n6086 gnd.n6019 585
R12257 gnd.n6087 gnd.n6018 585
R12258 gnd.n1146 gnd.n1145 585
R12259 gnd.n6094 gnd.n1144 585
R12260 gnd.n6095 gnd.n1143 585
R12261 gnd.n6096 gnd.n1142 585
R12262 gnd.n5901 gnd.n1141 585
R12263 gnd.n5903 gnd.n5902 585
R12264 gnd.n5904 gnd.n5900 585
R12265 gnd.n5899 gnd.n5897 585
R12266 gnd.n5908 gnd.n5896 585
R12267 gnd.n5909 gnd.n5895 585
R12268 gnd.n5910 gnd.n1168 585
R12269 gnd.n6229 gnd.n6228 585
R12270 gnd.n996 gnd.n994 585
R12271 gnd.n1027 gnd.n1026 585
R12272 gnd.n1025 gnd.n1013 585
R12273 gnd.n3906 gnd.n3905 537.605
R12274 gnd.n5803 gnd.n5802 482.89
R12275 gnd.n5686 gnd.n5685 482.89
R12276 gnd.n2023 gnd.n1629 482.89
R12277 gnd.n5158 gnd.n1631 482.89
R12278 gnd.n1687 gnd.t96 443.966
R12279 gnd.n1282 gnd.t116 443.966
R12280 gnd.n1689 gnd.t144 443.966
R12281 gnd.n1276 gnd.t45 443.966
R12282 gnd.n2154 gnd.t74 371.625
R12283 gnd.n6218 gnd.t34 371.625
R12284 gnd.n7430 gnd.t52 371.625
R12285 gnd.n7452 gnd.t60 371.625
R12286 gnd.n7474 gnd.t84 371.625
R12287 gnd.n1091 gnd.t122 371.625
R12288 gnd.n1114 gnd.t125 371.625
R12289 gnd.n1136 gnd.t87 371.625
R12290 gnd.n7321 gnd.t131 371.625
R12291 gnd.n2150 gnd.t63 371.625
R12292 gnd.n4146 gnd.t70 371.625
R12293 gnd.n3957 gnd.t78 371.625
R12294 gnd.n4067 gnd.t100 371.625
R12295 gnd.n3913 gnd.t119 371.625
R12296 gnd.n1760 gnd.t93 371.625
R12297 gnd.n838 gnd.t110 371.625
R12298 gnd.n1863 gnd.t138 371.625
R12299 gnd.n1015 gnd.t38 371.625
R12300 gnd.n2925 gnd.t56 323.425
R12301 gnd.n2451 gnd.t106 323.425
R12302 gnd.n3773 gnd.n3747 289.615
R12303 gnd.n3741 gnd.n3715 289.615
R12304 gnd.n3709 gnd.n3683 289.615
R12305 gnd.n3678 gnd.n3652 289.615
R12306 gnd.n3646 gnd.n3620 289.615
R12307 gnd.n3614 gnd.n3588 289.615
R12308 gnd.n3582 gnd.n3556 289.615
R12309 gnd.n3551 gnd.n3525 289.615
R12310 gnd.n2999 gnd.t30 279.217
R12311 gnd.n2477 gnd.t134 279.217
R12312 gnd.n1638 gnd.t130 260.649
R12313 gnd.n1243 gnd.t44 260.649
R12314 gnd.n5152 gnd.n5151 256.663
R12315 gnd.n5151 gnd.n1655 256.663
R12316 gnd.n5151 gnd.n1656 256.663
R12317 gnd.n5151 gnd.n1657 256.663
R12318 gnd.n5151 gnd.n1658 256.663
R12319 gnd.n5151 gnd.n1659 256.663
R12320 gnd.n5151 gnd.n1660 256.663
R12321 gnd.n5151 gnd.n1661 256.663
R12322 gnd.n5151 gnd.n1662 256.663
R12323 gnd.n5151 gnd.n1663 256.663
R12324 gnd.n5151 gnd.n1664 256.663
R12325 gnd.n5151 gnd.n1665 256.663
R12326 gnd.n5151 gnd.n1666 256.663
R12327 gnd.n5151 gnd.n1667 256.663
R12328 gnd.n5151 gnd.n1668 256.663
R12329 gnd.n5151 gnd.n1669 256.663
R12330 gnd.n1954 gnd.n1953 256.663
R12331 gnd.n5151 gnd.n1670 256.663
R12332 gnd.n5151 gnd.n1671 256.663
R12333 gnd.n5151 gnd.n1672 256.663
R12334 gnd.n5151 gnd.n1673 256.663
R12335 gnd.n5151 gnd.n1674 256.663
R12336 gnd.n5151 gnd.n1675 256.663
R12337 gnd.n5151 gnd.n1676 256.663
R12338 gnd.n5151 gnd.n1677 256.663
R12339 gnd.n5151 gnd.n1678 256.663
R12340 gnd.n5151 gnd.n1679 256.663
R12341 gnd.n5151 gnd.n1680 256.663
R12342 gnd.n5151 gnd.n1681 256.663
R12343 gnd.n5151 gnd.n1682 256.663
R12344 gnd.n5151 gnd.n1683 256.663
R12345 gnd.n5151 gnd.n1684 256.663
R12346 gnd.n5151 gnd.n1685 256.663
R12347 gnd.n5151 gnd.n2024 256.663
R12348 gnd.n1306 gnd.n1253 256.663
R12349 gnd.n5691 gnd.n1253 256.663
R12350 gnd.n1303 gnd.n1253 256.663
R12351 gnd.n5698 gnd.n1253 256.663
R12352 gnd.n1300 gnd.n1253 256.663
R12353 gnd.n5705 gnd.n1253 256.663
R12354 gnd.n1297 gnd.n1253 256.663
R12355 gnd.n5712 gnd.n1253 256.663
R12356 gnd.n1294 gnd.n1253 256.663
R12357 gnd.n5719 gnd.n1253 256.663
R12358 gnd.n1291 gnd.n1253 256.663
R12359 gnd.n5726 gnd.n1253 256.663
R12360 gnd.n1288 gnd.n1253 256.663
R12361 gnd.n5733 gnd.n1253 256.663
R12362 gnd.n1285 gnd.n1253 256.663
R12363 gnd.n5741 gnd.n1253 256.663
R12364 gnd.n5744 gnd.n1101 256.663
R12365 gnd.n5745 gnd.n1253 256.663
R12366 gnd.n1279 gnd.n1253 256.663
R12367 gnd.n5752 gnd.n1253 256.663
R12368 gnd.n1274 gnd.n1253 256.663
R12369 gnd.n5759 gnd.n1253 256.663
R12370 gnd.n1271 gnd.n1253 256.663
R12371 gnd.n5766 gnd.n1253 256.663
R12372 gnd.n1268 gnd.n1253 256.663
R12373 gnd.n5773 gnd.n1253 256.663
R12374 gnd.n1265 gnd.n1253 256.663
R12375 gnd.n5780 gnd.n1253 256.663
R12376 gnd.n1262 gnd.n1253 256.663
R12377 gnd.n5787 gnd.n1253 256.663
R12378 gnd.n1259 gnd.n1253 256.663
R12379 gnd.n5794 gnd.n1253 256.663
R12380 gnd.n1256 gnd.n1253 256.663
R12381 gnd.n5801 gnd.n1253 256.663
R12382 gnd.n4247 gnd.n3906 242.672
R12383 gnd.n4245 gnd.n3906 242.672
R12384 gnd.n4239 gnd.n3906 242.672
R12385 gnd.n4237 gnd.n3906 242.672
R12386 gnd.n4231 gnd.n3906 242.672
R12387 gnd.n4229 gnd.n3906 242.672
R12388 gnd.n4223 gnd.n3906 242.672
R12389 gnd.n4221 gnd.n3906 242.672
R12390 gnd.n4211 gnd.n3906 242.672
R12391 gnd.n3053 gnd.n3052 242.672
R12392 gnd.n3053 gnd.n2963 242.672
R12393 gnd.n3053 gnd.n2964 242.672
R12394 gnd.n3053 gnd.n2965 242.672
R12395 gnd.n3053 gnd.n2966 242.672
R12396 gnd.n3053 gnd.n2967 242.672
R12397 gnd.n3053 gnd.n2968 242.672
R12398 gnd.n3053 gnd.n2969 242.672
R12399 gnd.n3053 gnd.n2970 242.672
R12400 gnd.n3053 gnd.n2971 242.672
R12401 gnd.n3053 gnd.n2972 242.672
R12402 gnd.n3053 gnd.n2973 242.672
R12403 gnd.n3054 gnd.n3053 242.672
R12404 gnd.n3905 gnd.n2426 242.672
R12405 gnd.n3905 gnd.n2425 242.672
R12406 gnd.n3905 gnd.n2424 242.672
R12407 gnd.n3905 gnd.n2423 242.672
R12408 gnd.n3905 gnd.n2422 242.672
R12409 gnd.n3905 gnd.n2421 242.672
R12410 gnd.n3905 gnd.n2420 242.672
R12411 gnd.n3905 gnd.n2419 242.672
R12412 gnd.n3905 gnd.n2418 242.672
R12413 gnd.n3905 gnd.n2417 242.672
R12414 gnd.n3905 gnd.n2416 242.672
R12415 gnd.n3905 gnd.n2415 242.672
R12416 gnd.n3905 gnd.n2414 242.672
R12417 gnd.n3137 gnd.n3136 242.672
R12418 gnd.n3136 gnd.n2875 242.672
R12419 gnd.n3136 gnd.n2876 242.672
R12420 gnd.n3136 gnd.n2877 242.672
R12421 gnd.n3136 gnd.n2878 242.672
R12422 gnd.n3136 gnd.n2879 242.672
R12423 gnd.n3136 gnd.n2880 242.672
R12424 gnd.n3136 gnd.n2881 242.672
R12425 gnd.n3905 gnd.n2427 242.672
R12426 gnd.n3905 gnd.n2428 242.672
R12427 gnd.n3905 gnd.n2429 242.672
R12428 gnd.n3905 gnd.n2430 242.672
R12429 gnd.n3905 gnd.n2431 242.672
R12430 gnd.n3905 gnd.n2432 242.672
R12431 gnd.n3905 gnd.n2433 242.672
R12432 gnd.n3905 gnd.n2434 242.672
R12433 gnd.n3975 gnd.n3906 242.672
R12434 gnd.n3983 gnd.n3906 242.672
R12435 gnd.n3985 gnd.n3906 242.672
R12436 gnd.n3993 gnd.n3906 242.672
R12437 gnd.n3995 gnd.n3906 242.672
R12438 gnd.n4003 gnd.n3906 242.672
R12439 gnd.n4005 gnd.n3906 242.672
R12440 gnd.n4013 gnd.n3906 242.672
R12441 gnd.n4015 gnd.n3906 242.672
R12442 gnd.n4023 gnd.n3906 242.672
R12443 gnd.n4025 gnd.n3906 242.672
R12444 gnd.n4033 gnd.n3906 242.672
R12445 gnd.n4035 gnd.n3906 242.672
R12446 gnd.n4043 gnd.n3906 242.672
R12447 gnd.n4045 gnd.n3906 242.672
R12448 gnd.n4053 gnd.n3906 242.672
R12449 gnd.n4055 gnd.n3906 242.672
R12450 gnd.n4063 gnd.n3906 242.672
R12451 gnd.n4065 gnd.n3906 242.672
R12452 gnd.n4075 gnd.n3906 242.672
R12453 gnd.n4077 gnd.n3906 242.672
R12454 gnd.n4085 gnd.n3906 242.672
R12455 gnd.n4087 gnd.n3906 242.672
R12456 gnd.n4095 gnd.n3906 242.672
R12457 gnd.n4097 gnd.n3906 242.672
R12458 gnd.n4105 gnd.n3906 242.672
R12459 gnd.n4107 gnd.n3906 242.672
R12460 gnd.n4116 gnd.n3906 242.672
R12461 gnd.n4119 gnd.n3906 242.672
R12462 gnd.n4657 gnd.n753 242.672
R12463 gnd.n4660 gnd.n753 242.672
R12464 gnd.n4668 gnd.n753 242.672
R12465 gnd.n4670 gnd.n753 242.672
R12466 gnd.n4678 gnd.n753 242.672
R12467 gnd.n4680 gnd.n753 242.672
R12468 gnd.n4688 gnd.n753 242.672
R12469 gnd.n4690 gnd.n753 242.672
R12470 gnd.n4698 gnd.n753 242.672
R12471 gnd.n4700 gnd.n753 242.672
R12472 gnd.n4708 gnd.n753 242.672
R12473 gnd.n4710 gnd.n753 242.672
R12474 gnd.n4718 gnd.n753 242.672
R12475 gnd.n4720 gnd.n753 242.672
R12476 gnd.n4728 gnd.n753 242.672
R12477 gnd.n4730 gnd.n753 242.672
R12478 gnd.n4738 gnd.n753 242.672
R12479 gnd.n4740 gnd.n753 242.672
R12480 gnd.n4748 gnd.n753 242.672
R12481 gnd.n4750 gnd.n753 242.672
R12482 gnd.n4758 gnd.n753 242.672
R12483 gnd.n4760 gnd.n753 242.672
R12484 gnd.n4768 gnd.n753 242.672
R12485 gnd.n4770 gnd.n753 242.672
R12486 gnd.n4778 gnd.n753 242.672
R12487 gnd.n4780 gnd.n753 242.672
R12488 gnd.n4788 gnd.n753 242.672
R12489 gnd.n4790 gnd.n753 242.672
R12490 gnd.n4798 gnd.n753 242.672
R12491 gnd.n4800 gnd.n753 242.672
R12492 gnd.n4808 gnd.n753 242.672
R12493 gnd.n4810 gnd.n753 242.672
R12494 gnd.n4818 gnd.n753 242.672
R12495 gnd.n4820 gnd.n753 242.672
R12496 gnd.n4828 gnd.n753 242.672
R12497 gnd.n4830 gnd.n753 242.672
R12498 gnd.n4838 gnd.n753 242.672
R12499 gnd.n4840 gnd.n753 242.672
R12500 gnd.n4848 gnd.n753 242.672
R12501 gnd.n4850 gnd.n753 242.672
R12502 gnd.n4859 gnd.n753 242.672
R12503 gnd.n4861 gnd.n753 242.672
R12504 gnd.n4941 gnd.n852 242.672
R12505 gnd.n2148 gnd.n852 242.672
R12506 gnd.n2145 gnd.n852 242.672
R12507 gnd.n2134 gnd.n852 242.672
R12508 gnd.n2122 gnd.n852 242.672
R12509 gnd.n2119 gnd.n852 242.672
R12510 gnd.n2108 gnd.n852 242.672
R12511 gnd.n2096 gnd.n852 242.672
R12512 gnd.n2093 gnd.n852 242.672
R12513 gnd.n6215 gnd.n1060 242.672
R12514 gnd.n6215 gnd.n1061 242.672
R12515 gnd.n6215 gnd.n1062 242.672
R12516 gnd.n6215 gnd.n1063 242.672
R12517 gnd.n6215 gnd.n1064 242.672
R12518 gnd.n6215 gnd.n1065 242.672
R12519 gnd.n6215 gnd.n1066 242.672
R12520 gnd.n6215 gnd.n1068 242.672
R12521 gnd.n6216 gnd.n6215 242.672
R12522 gnd.n7318 gnd.n253 242.672
R12523 gnd.n7401 gnd.n253 242.672
R12524 gnd.n7314 gnd.n253 242.672
R12525 gnd.n7408 gnd.n253 242.672
R12526 gnd.n7307 gnd.n253 242.672
R12527 gnd.n7415 gnd.n253 242.672
R12528 gnd.n7300 gnd.n253 242.672
R12529 gnd.n7422 gnd.n253 242.672
R12530 gnd.n7293 gnd.n253 242.672
R12531 gnd.n852 gnd.n841 242.672
R12532 gnd.n1896 gnd.n852 242.672
R12533 gnd.n1903 gnd.n852 242.672
R12534 gnd.n1890 gnd.n852 242.672
R12535 gnd.n1910 gnd.n852 242.672
R12536 gnd.n1883 gnd.n852 242.672
R12537 gnd.n1917 gnd.n852 242.672
R12538 gnd.n1876 gnd.n852 242.672
R12539 gnd.n1924 gnd.n852 242.672
R12540 gnd.n1927 gnd.n852 242.672
R12541 gnd.n1867 gnd.n852 242.672
R12542 gnd.n1936 gnd.n852 242.672
R12543 gnd.n1858 gnd.n852 242.672
R12544 gnd.n1943 gnd.n852 242.672
R12545 gnd.n1946 gnd.n852 242.672
R12546 gnd.n1849 gnd.n852 242.672
R12547 gnd.n1952 gnd.n1752 242.672
R12548 gnd.n1841 gnd.n852 242.672
R12549 gnd.n1840 gnd.n852 242.672
R12550 gnd.n1755 gnd.n852 242.672
R12551 gnd.n1830 gnd.n852 242.672
R12552 gnd.n1759 gnd.n852 242.672
R12553 gnd.n1821 gnd.n852 242.672
R12554 gnd.n1813 gnd.n852 242.672
R12555 gnd.n1811 gnd.n852 242.672
R12556 gnd.n1803 gnd.n852 242.672
R12557 gnd.n1801 gnd.n852 242.672
R12558 gnd.n1793 gnd.n852 242.672
R12559 gnd.n1791 gnd.n852 242.672
R12560 gnd.n1783 gnd.n852 242.672
R12561 gnd.n6215 gnd.n6214 242.672
R12562 gnd.n6215 gnd.n1032 242.672
R12563 gnd.n6215 gnd.n1033 242.672
R12564 gnd.n6215 gnd.n1034 242.672
R12565 gnd.n6215 gnd.n1035 242.672
R12566 gnd.n6215 gnd.n1036 242.672
R12567 gnd.n6215 gnd.n1037 242.672
R12568 gnd.n6215 gnd.n1038 242.672
R12569 gnd.n6215 gnd.n1039 242.672
R12570 gnd.n6215 gnd.n1040 242.672
R12571 gnd.n6215 gnd.n1041 242.672
R12572 gnd.n6215 gnd.n1042 242.672
R12573 gnd.n6215 gnd.n1043 242.672
R12574 gnd.n6162 gnd.n1102 242.672
R12575 gnd.n6215 gnd.n1044 242.672
R12576 gnd.n6215 gnd.n1045 242.672
R12577 gnd.n6215 gnd.n1046 242.672
R12578 gnd.n6215 gnd.n1047 242.672
R12579 gnd.n6215 gnd.n1048 242.672
R12580 gnd.n6215 gnd.n1049 242.672
R12581 gnd.n6215 gnd.n1050 242.672
R12582 gnd.n6215 gnd.n1051 242.672
R12583 gnd.n6215 gnd.n1052 242.672
R12584 gnd.n6215 gnd.n1053 242.672
R12585 gnd.n6215 gnd.n1054 242.672
R12586 gnd.n6215 gnd.n1055 242.672
R12587 gnd.n6215 gnd.n1056 242.672
R12588 gnd.n6215 gnd.n1057 242.672
R12589 gnd.n6215 gnd.n1058 242.672
R12590 gnd.n6215 gnd.n1059 242.672
R12591 gnd.n7637 gnd.n253 242.672
R12592 gnd.n7433 gnd.n253 242.672
R12593 gnd.n7627 gnd.n253 242.672
R12594 gnd.n7437 gnd.n253 242.672
R12595 gnd.n7617 gnd.n253 242.672
R12596 gnd.n7441 gnd.n253 242.672
R12597 gnd.n7607 gnd.n253 242.672
R12598 gnd.n7445 gnd.n253 242.672
R12599 gnd.n7597 gnd.n253 242.672
R12600 gnd.n7449 gnd.n253 242.672
R12601 gnd.n7587 gnd.n253 242.672
R12602 gnd.n7455 gnd.n253 242.672
R12603 gnd.n7577 gnd.n253 242.672
R12604 gnd.n7459 gnd.n253 242.672
R12605 gnd.n7567 gnd.n253 242.672
R12606 gnd.n7463 gnd.n253 242.672
R12607 gnd.n7557 gnd.n253 242.672
R12608 gnd.n7467 gnd.n253 242.672
R12609 gnd.n7547 gnd.n253 242.672
R12610 gnd.n7471 gnd.n253 242.672
R12611 gnd.n7537 gnd.n253 242.672
R12612 gnd.n7527 gnd.n253 242.672
R12613 gnd.n7526 gnd.n253 242.672
R12614 gnd.n7481 gnd.n253 242.672
R12615 gnd.n7516 gnd.n253 242.672
R12616 gnd.n7485 gnd.n253 242.672
R12617 gnd.n7506 gnd.n253 242.672
R12618 gnd.n7489 gnd.n253 242.672
R12619 gnd.n7496 gnd.n253 242.672
R12620 gnd.n5006 gnd.n853 242.672
R12621 gnd.n2072 gnd.n853 242.672
R12622 gnd.n2075 gnd.n853 242.672
R12623 gnd.n2085 gnd.n853 242.672
R12624 gnd.n2088 gnd.n853 242.672
R12625 gnd.n2100 gnd.n853 242.672
R12626 gnd.n2103 gnd.n853 242.672
R12627 gnd.n2114 gnd.n853 242.672
R12628 gnd.n2126 gnd.n853 242.672
R12629 gnd.n2129 gnd.n853 242.672
R12630 gnd.n2140 gnd.n853 242.672
R12631 gnd.n2157 gnd.n853 242.672
R12632 gnd.n2160 gnd.n853 242.672
R12633 gnd.n2162 gnd.n853 242.672
R12634 gnd.n6226 gnd.n1009 242.672
R12635 gnd.n6226 gnd.n1008 242.672
R12636 gnd.n6226 gnd.n1007 242.672
R12637 gnd.n6226 gnd.n1006 242.672
R12638 gnd.n6226 gnd.n1005 242.672
R12639 gnd.n6226 gnd.n1004 242.672
R12640 gnd.n6226 gnd.n1003 242.672
R12641 gnd.n6226 gnd.n1002 242.672
R12642 gnd.n6226 gnd.n1001 242.672
R12643 gnd.n6226 gnd.n1000 242.672
R12644 gnd.n6226 gnd.n999 242.672
R12645 gnd.n6226 gnd.n998 242.672
R12646 gnd.n6227 gnd.n6226 242.672
R12647 gnd.n6226 gnd.n1010 242.672
R12648 gnd.n7495 gnd.n249 240.244
R12649 gnd.n7498 gnd.n7497 240.244
R12650 gnd.n7505 gnd.n7504 240.244
R12651 gnd.n7508 gnd.n7507 240.244
R12652 gnd.n7515 gnd.n7514 240.244
R12653 gnd.n7518 gnd.n7517 240.244
R12654 gnd.n7525 gnd.n7524 240.244
R12655 gnd.n7529 gnd.n7528 240.244
R12656 gnd.n7536 gnd.n7477 240.244
R12657 gnd.n7539 gnd.n7538 240.244
R12658 gnd.n7546 gnd.n7545 240.244
R12659 gnd.n7549 gnd.n7548 240.244
R12660 gnd.n7556 gnd.n7555 240.244
R12661 gnd.n7559 gnd.n7558 240.244
R12662 gnd.n7566 gnd.n7565 240.244
R12663 gnd.n7569 gnd.n7568 240.244
R12664 gnd.n7576 gnd.n7575 240.244
R12665 gnd.n7579 gnd.n7578 240.244
R12666 gnd.n7586 gnd.n7585 240.244
R12667 gnd.n7589 gnd.n7588 240.244
R12668 gnd.n7596 gnd.n7595 240.244
R12669 gnd.n7599 gnd.n7598 240.244
R12670 gnd.n7606 gnd.n7605 240.244
R12671 gnd.n7609 gnd.n7608 240.244
R12672 gnd.n7616 gnd.n7615 240.244
R12673 gnd.n7619 gnd.n7618 240.244
R12674 gnd.n7626 gnd.n7625 240.244
R12675 gnd.n7629 gnd.n7628 240.244
R12676 gnd.n7636 gnd.n7635 240.244
R12677 gnd.n5959 gnd.n1153 240.244
R12678 gnd.n5960 gnd.n5959 240.244
R12679 gnd.n5960 gnd.n5937 240.244
R12680 gnd.n5942 gnd.n5937 240.244
R12681 gnd.n5982 gnd.n5942 240.244
R12682 gnd.n5982 gnd.n392 240.244
R12683 gnd.n7039 gnd.n392 240.244
R12684 gnd.n7039 gnd.n382 240.244
R12685 gnd.n382 gnd.n373 240.244
R12686 gnd.n7071 gnd.n373 240.244
R12687 gnd.n7071 gnd.n363 240.244
R12688 gnd.n7075 gnd.n363 240.244
R12689 gnd.n7075 gnd.n353 240.244
R12690 gnd.n353 gnd.n345 240.244
R12691 gnd.n7127 gnd.n345 240.244
R12692 gnd.n7127 gnd.n336 240.244
R12693 gnd.n336 gnd.n327 240.244
R12694 gnd.n7146 gnd.n327 240.244
R12695 gnd.n7147 gnd.n7146 240.244
R12696 gnd.n7147 gnd.n319 240.244
R12697 gnd.n319 gnd.n309 240.244
R12698 gnd.n7166 gnd.n309 240.244
R12699 gnd.n7167 gnd.n7166 240.244
R12700 gnd.n7167 gnd.n299 240.244
R12701 gnd.n7170 gnd.n299 240.244
R12702 gnd.n7170 gnd.n290 240.244
R12703 gnd.n290 gnd.n282 240.244
R12704 gnd.n7205 gnd.n282 240.244
R12705 gnd.n7205 gnd.n275 240.244
R12706 gnd.n7207 gnd.n275 240.244
R12707 gnd.n7207 gnd.n266 240.244
R12708 gnd.n266 gnd.n261 240.244
R12709 gnd.n7231 gnd.n261 240.244
R12710 gnd.n7231 gnd.n105 240.244
R12711 gnd.n7238 gnd.n105 240.244
R12712 gnd.n7238 gnd.n116 240.244
R12713 gnd.n7241 gnd.n116 240.244
R12714 gnd.n7241 gnd.n127 240.244
R12715 gnd.n7245 gnd.n127 240.244
R12716 gnd.n7245 gnd.n137 240.244
R12717 gnd.n7248 gnd.n137 240.244
R12718 gnd.n7248 gnd.n146 240.244
R12719 gnd.n7252 gnd.n146 240.244
R12720 gnd.n7252 gnd.n156 240.244
R12721 gnd.n7255 gnd.n156 240.244
R12722 gnd.n7255 gnd.n165 240.244
R12723 gnd.n7259 gnd.n165 240.244
R12724 gnd.n7259 gnd.n176 240.244
R12725 gnd.n7262 gnd.n176 240.244
R12726 gnd.n7262 gnd.n185 240.244
R12727 gnd.n7266 gnd.n185 240.244
R12728 gnd.n7266 gnd.n195 240.244
R12729 gnd.n7269 gnd.n195 240.244
R12730 gnd.n7269 gnd.n204 240.244
R12731 gnd.n7273 gnd.n204 240.244
R12732 gnd.n7273 gnd.n214 240.244
R12733 gnd.n7276 gnd.n214 240.244
R12734 gnd.n7276 gnd.n223 240.244
R12735 gnd.n7280 gnd.n223 240.244
R12736 gnd.n7280 gnd.n233 240.244
R12737 gnd.n7283 gnd.n233 240.244
R12738 gnd.n7283 gnd.n242 240.244
R12739 gnd.n7286 gnd.n242 240.244
R12740 gnd.n7286 gnd.n251 240.244
R12741 gnd.n1071 gnd.n1070 240.244
R12742 gnd.n6208 gnd.n1070 240.244
R12743 gnd.n6206 gnd.n6205 240.244
R12744 gnd.n6202 gnd.n6201 240.244
R12745 gnd.n6198 gnd.n6197 240.244
R12746 gnd.n6194 gnd.n6193 240.244
R12747 gnd.n6190 gnd.n6189 240.244
R12748 gnd.n6186 gnd.n6185 240.244
R12749 gnd.n6182 gnd.n6181 240.244
R12750 gnd.n6177 gnd.n6176 240.244
R12751 gnd.n6173 gnd.n6172 240.244
R12752 gnd.n6169 gnd.n6168 240.244
R12753 gnd.n6165 gnd.n6164 240.244
R12754 gnd.n6160 gnd.n6159 240.244
R12755 gnd.n6156 gnd.n6155 240.244
R12756 gnd.n6152 gnd.n6151 240.244
R12757 gnd.n6148 gnd.n6147 240.244
R12758 gnd.n6144 gnd.n6143 240.244
R12759 gnd.n6140 gnd.n6139 240.244
R12760 gnd.n6136 gnd.n6135 240.244
R12761 gnd.n6132 gnd.n6131 240.244
R12762 gnd.n6128 gnd.n6127 240.244
R12763 gnd.n6124 gnd.n6123 240.244
R12764 gnd.n6120 gnd.n6119 240.244
R12765 gnd.n6116 gnd.n6115 240.244
R12766 gnd.n6112 gnd.n6111 240.244
R12767 gnd.n6108 gnd.n6107 240.244
R12768 gnd.n6104 gnd.n6103 240.244
R12769 gnd.n5993 gnd.n1072 240.244
R12770 gnd.n5993 gnd.n5941 240.244
R12771 gnd.n6001 gnd.n5941 240.244
R12772 gnd.n6001 gnd.n5989 240.244
R12773 gnd.n5989 gnd.n390 240.244
R12774 gnd.n7052 gnd.n390 240.244
R12775 gnd.n7052 gnd.n385 240.244
R12776 gnd.n7060 gnd.n385 240.244
R12777 gnd.n7060 gnd.n386 240.244
R12778 gnd.n386 gnd.n361 240.244
R12779 gnd.n7088 gnd.n361 240.244
R12780 gnd.n7088 gnd.n356 240.244
R12781 gnd.n7096 gnd.n356 240.244
R12782 gnd.n7096 gnd.n357 240.244
R12783 gnd.n357 gnd.n334 240.244
R12784 gnd.n7138 gnd.n334 240.244
R12785 gnd.n7138 gnd.n330 240.244
R12786 gnd.n7144 gnd.n330 240.244
R12787 gnd.n7144 gnd.n317 240.244
R12788 gnd.n7158 gnd.n317 240.244
R12789 gnd.n7158 gnd.n313 240.244
R12790 gnd.n7164 gnd.n313 240.244
R12791 gnd.n7164 gnd.n297 240.244
R12792 gnd.n7182 gnd.n297 240.244
R12793 gnd.n7182 gnd.n292 240.244
R12794 gnd.n7190 gnd.n292 240.244
R12795 gnd.n7190 gnd.n293 240.244
R12796 gnd.n293 gnd.n274 240.244
R12797 gnd.n7214 gnd.n274 240.244
R12798 gnd.n7214 gnd.n269 240.244
R12799 gnd.n7223 gnd.n269 240.244
R12800 gnd.n7223 gnd.n270 240.244
R12801 gnd.n270 gnd.n108 240.244
R12802 gnd.n7734 gnd.n108 240.244
R12803 gnd.n7734 gnd.n109 240.244
R12804 gnd.n7730 gnd.n109 240.244
R12805 gnd.n7730 gnd.n115 240.244
R12806 gnd.n7722 gnd.n115 240.244
R12807 gnd.n7722 gnd.n129 240.244
R12808 gnd.n7718 gnd.n129 240.244
R12809 gnd.n7718 gnd.n135 240.244
R12810 gnd.n7710 gnd.n135 240.244
R12811 gnd.n7710 gnd.n149 240.244
R12812 gnd.n7706 gnd.n149 240.244
R12813 gnd.n7706 gnd.n155 240.244
R12814 gnd.n7698 gnd.n155 240.244
R12815 gnd.n7698 gnd.n168 240.244
R12816 gnd.n7694 gnd.n168 240.244
R12817 gnd.n7694 gnd.n174 240.244
R12818 gnd.n7686 gnd.n174 240.244
R12819 gnd.n7686 gnd.n188 240.244
R12820 gnd.n7682 gnd.n188 240.244
R12821 gnd.n7682 gnd.n194 240.244
R12822 gnd.n7674 gnd.n194 240.244
R12823 gnd.n7674 gnd.n206 240.244
R12824 gnd.n7670 gnd.n206 240.244
R12825 gnd.n7670 gnd.n212 240.244
R12826 gnd.n7662 gnd.n212 240.244
R12827 gnd.n7662 gnd.n226 240.244
R12828 gnd.n7658 gnd.n226 240.244
R12829 gnd.n7658 gnd.n232 240.244
R12830 gnd.n7650 gnd.n232 240.244
R12831 gnd.n7650 gnd.n244 240.244
R12832 gnd.n7646 gnd.n244 240.244
R12833 gnd.n7290 gnd.n254 240.244
R12834 gnd.n7424 gnd.n7423 240.244
R12835 gnd.n7421 gnd.n7294 240.244
R12836 gnd.n7417 gnd.n7416 240.244
R12837 gnd.n7414 gnd.n7301 240.244
R12838 gnd.n7410 gnd.n7409 240.244
R12839 gnd.n7407 gnd.n7308 240.244
R12840 gnd.n7403 gnd.n7402 240.244
R12841 gnd.n7400 gnd.n7315 240.244
R12842 gnd.n5971 gnd.n1154 240.244
R12843 gnd.n5972 gnd.n5971 240.244
R12844 gnd.n5972 gnd.n5938 240.244
R12845 gnd.n5943 gnd.n5938 240.244
R12846 gnd.n5980 gnd.n5943 240.244
R12847 gnd.n5980 gnd.n393 240.244
R12848 gnd.n393 gnd.n380 240.244
R12849 gnd.n7062 gnd.n380 240.244
R12850 gnd.n7062 gnd.n375 240.244
R12851 gnd.n7069 gnd.n375 240.244
R12852 gnd.n7069 gnd.n364 240.244
R12853 gnd.n364 gnd.n351 240.244
R12854 gnd.n7098 gnd.n351 240.244
R12855 gnd.n7098 gnd.n346 240.244
R12856 gnd.n7125 gnd.n346 240.244
R12857 gnd.n7125 gnd.n337 240.244
R12858 gnd.n7103 gnd.n337 240.244
R12859 gnd.n7103 gnd.n328 240.244
R12860 gnd.n7104 gnd.n328 240.244
R12861 gnd.n7104 gnd.n320 240.244
R12862 gnd.n7107 gnd.n320 240.244
R12863 gnd.n7107 gnd.n311 240.244
R12864 gnd.n7108 gnd.n311 240.244
R12865 gnd.n7108 gnd.n300 240.244
R12866 gnd.n300 gnd.n289 240.244
R12867 gnd.n7192 gnd.n289 240.244
R12868 gnd.n7192 gnd.n284 240.244
R12869 gnd.n7203 gnd.n284 240.244
R12870 gnd.n7203 gnd.n276 240.244
R12871 gnd.n7196 gnd.n276 240.244
R12872 gnd.n7196 gnd.n268 240.244
R12873 gnd.n268 gnd.n267 240.244
R12874 gnd.n267 gnd.n102 240.244
R12875 gnd.n7736 gnd.n102 240.244
R12876 gnd.n7736 gnd.n104 240.244
R12877 gnd.n117 gnd.n104 240.244
R12878 gnd.n7342 gnd.n117 240.244
R12879 gnd.n7342 gnd.n128 240.244
R12880 gnd.n7350 gnd.n128 240.244
R12881 gnd.n7350 gnd.n138 240.244
R12882 gnd.n7339 gnd.n138 240.244
R12883 gnd.n7339 gnd.n147 240.244
R12884 gnd.n7357 gnd.n147 240.244
R12885 gnd.n7357 gnd.n157 240.244
R12886 gnd.n7336 gnd.n157 240.244
R12887 gnd.n7336 gnd.n166 240.244
R12888 gnd.n7364 gnd.n166 240.244
R12889 gnd.n7364 gnd.n177 240.244
R12890 gnd.n7333 gnd.n177 240.244
R12891 gnd.n7333 gnd.n186 240.244
R12892 gnd.n7371 gnd.n186 240.244
R12893 gnd.n7371 gnd.n196 240.244
R12894 gnd.n7330 gnd.n196 240.244
R12895 gnd.n7330 gnd.n205 240.244
R12896 gnd.n7378 gnd.n205 240.244
R12897 gnd.n7378 gnd.n215 240.244
R12898 gnd.n7327 gnd.n215 240.244
R12899 gnd.n7327 gnd.n224 240.244
R12900 gnd.n7385 gnd.n224 240.244
R12901 gnd.n7385 gnd.n234 240.244
R12902 gnd.n7324 gnd.n234 240.244
R12903 gnd.n7324 gnd.n243 240.244
R12904 gnd.n7392 gnd.n243 240.244
R12905 gnd.n7392 gnd.n252 240.244
R12906 gnd.n6015 gnd.n6014 240.244
R12907 gnd.n6023 gnd.n6022 240.244
R12908 gnd.n6025 gnd.n6024 240.244
R12909 gnd.n6035 gnd.n6034 240.244
R12910 gnd.n6043 gnd.n6042 240.244
R12911 gnd.n6045 gnd.n6044 240.244
R12912 gnd.n6055 gnd.n6054 240.244
R12913 gnd.n1067 gnd.n1021 240.244
R12914 gnd.n6217 gnd.n1030 240.244
R12915 gnd.n6011 gnd.n1149 240.244
R12916 gnd.n5956 gnd.n1149 240.244
R12917 gnd.n5956 gnd.n5940 240.244
R12918 gnd.n5987 gnd.n5940 240.244
R12919 gnd.n5987 gnd.n394 240.244
R12920 gnd.n7050 gnd.n394 240.244
R12921 gnd.n7050 gnd.n395 240.244
R12922 gnd.n395 gnd.n384 240.244
R12923 gnd.n7045 gnd.n384 240.244
R12924 gnd.n7045 gnd.n366 240.244
R12925 gnd.n7086 gnd.n366 240.244
R12926 gnd.n7086 gnd.n367 240.244
R12927 gnd.n367 gnd.n355 240.244
R12928 gnd.n7081 gnd.n355 240.244
R12929 gnd.n7081 gnd.n339 240.244
R12930 gnd.n7136 gnd.n339 240.244
R12931 gnd.n7136 gnd.n340 240.244
R12932 gnd.n340 gnd.n329 240.244
R12933 gnd.n329 gnd.n321 240.244
R12934 gnd.n7156 gnd.n321 240.244
R12935 gnd.n7156 gnd.n322 240.244
R12936 gnd.n322 gnd.n312 240.244
R12937 gnd.n312 gnd.n302 240.244
R12938 gnd.n7180 gnd.n302 240.244
R12939 gnd.n7180 gnd.n303 240.244
R12940 gnd.n303 gnd.n291 240.244
R12941 gnd.n7175 gnd.n291 240.244
R12942 gnd.n7175 gnd.n278 240.244
R12943 gnd.n7212 gnd.n278 240.244
R12944 gnd.n7212 gnd.n265 240.244
R12945 gnd.n7225 gnd.n265 240.244
R12946 gnd.n7225 gnd.n259 240.244
R12947 gnd.n7233 gnd.n259 240.244
R12948 gnd.n7233 gnd.n107 240.244
R12949 gnd.n119 gnd.n107 240.244
R12950 gnd.n7728 gnd.n119 240.244
R12951 gnd.n7728 gnd.n120 240.244
R12952 gnd.n7724 gnd.n120 240.244
R12953 gnd.n7724 gnd.n126 240.244
R12954 gnd.n7716 gnd.n126 240.244
R12955 gnd.n7716 gnd.n140 240.244
R12956 gnd.n7712 gnd.n140 240.244
R12957 gnd.n7712 gnd.n145 240.244
R12958 gnd.n7704 gnd.n145 240.244
R12959 gnd.n7704 gnd.n159 240.244
R12960 gnd.n7700 gnd.n159 240.244
R12961 gnd.n7700 gnd.n164 240.244
R12962 gnd.n7692 gnd.n164 240.244
R12963 gnd.n7692 gnd.n179 240.244
R12964 gnd.n7688 gnd.n179 240.244
R12965 gnd.n7688 gnd.n184 240.244
R12966 gnd.n7680 gnd.n184 240.244
R12967 gnd.n7680 gnd.n198 240.244
R12968 gnd.n7676 gnd.n198 240.244
R12969 gnd.n7676 gnd.n203 240.244
R12970 gnd.n7668 gnd.n203 240.244
R12971 gnd.n7668 gnd.n217 240.244
R12972 gnd.n7664 gnd.n217 240.244
R12973 gnd.n7664 gnd.n222 240.244
R12974 gnd.n7656 gnd.n222 240.244
R12975 gnd.n7656 gnd.n236 240.244
R12976 gnd.n7652 gnd.n236 240.244
R12977 gnd.n7652 gnd.n241 240.244
R12978 gnd.n7644 gnd.n241 240.244
R12979 gnd.n6455 gnd.n748 240.244
R12980 gnd.n6461 gnd.n748 240.244
R12981 gnd.n6461 gnd.n746 240.244
R12982 gnd.n6465 gnd.n746 240.244
R12983 gnd.n6465 gnd.n742 240.244
R12984 gnd.n6471 gnd.n742 240.244
R12985 gnd.n6471 gnd.n740 240.244
R12986 gnd.n6475 gnd.n740 240.244
R12987 gnd.n6475 gnd.n736 240.244
R12988 gnd.n6481 gnd.n736 240.244
R12989 gnd.n6481 gnd.n734 240.244
R12990 gnd.n6485 gnd.n734 240.244
R12991 gnd.n6485 gnd.n730 240.244
R12992 gnd.n6491 gnd.n730 240.244
R12993 gnd.n6491 gnd.n728 240.244
R12994 gnd.n6495 gnd.n728 240.244
R12995 gnd.n6495 gnd.n724 240.244
R12996 gnd.n6501 gnd.n724 240.244
R12997 gnd.n6501 gnd.n722 240.244
R12998 gnd.n6505 gnd.n722 240.244
R12999 gnd.n6505 gnd.n718 240.244
R13000 gnd.n6511 gnd.n718 240.244
R13001 gnd.n6511 gnd.n716 240.244
R13002 gnd.n6515 gnd.n716 240.244
R13003 gnd.n6515 gnd.n712 240.244
R13004 gnd.n6521 gnd.n712 240.244
R13005 gnd.n6521 gnd.n710 240.244
R13006 gnd.n6525 gnd.n710 240.244
R13007 gnd.n6525 gnd.n706 240.244
R13008 gnd.n6531 gnd.n706 240.244
R13009 gnd.n6531 gnd.n704 240.244
R13010 gnd.n6535 gnd.n704 240.244
R13011 gnd.n6535 gnd.n700 240.244
R13012 gnd.n6541 gnd.n700 240.244
R13013 gnd.n6541 gnd.n698 240.244
R13014 gnd.n6545 gnd.n698 240.244
R13015 gnd.n6545 gnd.n694 240.244
R13016 gnd.n6551 gnd.n694 240.244
R13017 gnd.n6551 gnd.n692 240.244
R13018 gnd.n6555 gnd.n692 240.244
R13019 gnd.n6555 gnd.n688 240.244
R13020 gnd.n6561 gnd.n688 240.244
R13021 gnd.n6561 gnd.n686 240.244
R13022 gnd.n6565 gnd.n686 240.244
R13023 gnd.n6565 gnd.n682 240.244
R13024 gnd.n6571 gnd.n682 240.244
R13025 gnd.n6571 gnd.n680 240.244
R13026 gnd.n6575 gnd.n680 240.244
R13027 gnd.n6575 gnd.n676 240.244
R13028 gnd.n6581 gnd.n676 240.244
R13029 gnd.n6581 gnd.n674 240.244
R13030 gnd.n6585 gnd.n674 240.244
R13031 gnd.n6585 gnd.n670 240.244
R13032 gnd.n6591 gnd.n670 240.244
R13033 gnd.n6591 gnd.n668 240.244
R13034 gnd.n6595 gnd.n668 240.244
R13035 gnd.n6595 gnd.n664 240.244
R13036 gnd.n6601 gnd.n664 240.244
R13037 gnd.n6601 gnd.n662 240.244
R13038 gnd.n6605 gnd.n662 240.244
R13039 gnd.n6605 gnd.n658 240.244
R13040 gnd.n6611 gnd.n658 240.244
R13041 gnd.n6611 gnd.n656 240.244
R13042 gnd.n6615 gnd.n656 240.244
R13043 gnd.n6615 gnd.n652 240.244
R13044 gnd.n6621 gnd.n652 240.244
R13045 gnd.n6621 gnd.n650 240.244
R13046 gnd.n6625 gnd.n650 240.244
R13047 gnd.n6625 gnd.n646 240.244
R13048 gnd.n6631 gnd.n646 240.244
R13049 gnd.n6631 gnd.n644 240.244
R13050 gnd.n6635 gnd.n644 240.244
R13051 gnd.n6635 gnd.n640 240.244
R13052 gnd.n6641 gnd.n640 240.244
R13053 gnd.n6641 gnd.n638 240.244
R13054 gnd.n6645 gnd.n638 240.244
R13055 gnd.n6645 gnd.n634 240.244
R13056 gnd.n6651 gnd.n634 240.244
R13057 gnd.n6651 gnd.n632 240.244
R13058 gnd.n6655 gnd.n632 240.244
R13059 gnd.n6655 gnd.n628 240.244
R13060 gnd.n6661 gnd.n628 240.244
R13061 gnd.n6661 gnd.n626 240.244
R13062 gnd.n6665 gnd.n626 240.244
R13063 gnd.n6665 gnd.n622 240.244
R13064 gnd.n6671 gnd.n622 240.244
R13065 gnd.n6671 gnd.n620 240.244
R13066 gnd.n6675 gnd.n620 240.244
R13067 gnd.n6675 gnd.n616 240.244
R13068 gnd.n6681 gnd.n616 240.244
R13069 gnd.n6681 gnd.n614 240.244
R13070 gnd.n6685 gnd.n614 240.244
R13071 gnd.n6685 gnd.n610 240.244
R13072 gnd.n6691 gnd.n610 240.244
R13073 gnd.n6691 gnd.n608 240.244
R13074 gnd.n6695 gnd.n608 240.244
R13075 gnd.n6695 gnd.n604 240.244
R13076 gnd.n6701 gnd.n604 240.244
R13077 gnd.n6701 gnd.n602 240.244
R13078 gnd.n6705 gnd.n602 240.244
R13079 gnd.n6705 gnd.n598 240.244
R13080 gnd.n6711 gnd.n598 240.244
R13081 gnd.n6711 gnd.n596 240.244
R13082 gnd.n6715 gnd.n596 240.244
R13083 gnd.n6715 gnd.n592 240.244
R13084 gnd.n6721 gnd.n592 240.244
R13085 gnd.n6721 gnd.n590 240.244
R13086 gnd.n6725 gnd.n590 240.244
R13087 gnd.n6725 gnd.n586 240.244
R13088 gnd.n6731 gnd.n586 240.244
R13089 gnd.n6731 gnd.n584 240.244
R13090 gnd.n6735 gnd.n584 240.244
R13091 gnd.n6735 gnd.n580 240.244
R13092 gnd.n6741 gnd.n580 240.244
R13093 gnd.n6741 gnd.n578 240.244
R13094 gnd.n6745 gnd.n578 240.244
R13095 gnd.n6745 gnd.n574 240.244
R13096 gnd.n6751 gnd.n574 240.244
R13097 gnd.n6751 gnd.n572 240.244
R13098 gnd.n6755 gnd.n572 240.244
R13099 gnd.n6755 gnd.n568 240.244
R13100 gnd.n6761 gnd.n568 240.244
R13101 gnd.n6761 gnd.n566 240.244
R13102 gnd.n6765 gnd.n566 240.244
R13103 gnd.n6765 gnd.n562 240.244
R13104 gnd.n6771 gnd.n562 240.244
R13105 gnd.n6771 gnd.n560 240.244
R13106 gnd.n6775 gnd.n560 240.244
R13107 gnd.n6775 gnd.n556 240.244
R13108 gnd.n6781 gnd.n556 240.244
R13109 gnd.n6781 gnd.n554 240.244
R13110 gnd.n6785 gnd.n554 240.244
R13111 gnd.n6785 gnd.n550 240.244
R13112 gnd.n6791 gnd.n550 240.244
R13113 gnd.n6791 gnd.n548 240.244
R13114 gnd.n6795 gnd.n548 240.244
R13115 gnd.n6795 gnd.n544 240.244
R13116 gnd.n6802 gnd.n544 240.244
R13117 gnd.n6802 gnd.n542 240.244
R13118 gnd.n6806 gnd.n542 240.244
R13119 gnd.n6806 gnd.n539 240.244
R13120 gnd.n6812 gnd.n537 240.244
R13121 gnd.n6816 gnd.n537 240.244
R13122 gnd.n6816 gnd.n533 240.244
R13123 gnd.n6822 gnd.n533 240.244
R13124 gnd.n6822 gnd.n531 240.244
R13125 gnd.n6826 gnd.n531 240.244
R13126 gnd.n6826 gnd.n527 240.244
R13127 gnd.n6832 gnd.n527 240.244
R13128 gnd.n6832 gnd.n525 240.244
R13129 gnd.n6836 gnd.n525 240.244
R13130 gnd.n6836 gnd.n521 240.244
R13131 gnd.n6842 gnd.n521 240.244
R13132 gnd.n6842 gnd.n519 240.244
R13133 gnd.n6846 gnd.n519 240.244
R13134 gnd.n6846 gnd.n515 240.244
R13135 gnd.n6852 gnd.n515 240.244
R13136 gnd.n6852 gnd.n513 240.244
R13137 gnd.n6856 gnd.n513 240.244
R13138 gnd.n6856 gnd.n509 240.244
R13139 gnd.n6862 gnd.n509 240.244
R13140 gnd.n6862 gnd.n507 240.244
R13141 gnd.n6866 gnd.n507 240.244
R13142 gnd.n6866 gnd.n503 240.244
R13143 gnd.n6872 gnd.n503 240.244
R13144 gnd.n6872 gnd.n501 240.244
R13145 gnd.n6876 gnd.n501 240.244
R13146 gnd.n6876 gnd.n497 240.244
R13147 gnd.n6882 gnd.n497 240.244
R13148 gnd.n6882 gnd.n495 240.244
R13149 gnd.n6886 gnd.n495 240.244
R13150 gnd.n6886 gnd.n491 240.244
R13151 gnd.n6892 gnd.n491 240.244
R13152 gnd.n6892 gnd.n489 240.244
R13153 gnd.n6896 gnd.n489 240.244
R13154 gnd.n6896 gnd.n485 240.244
R13155 gnd.n6902 gnd.n485 240.244
R13156 gnd.n6902 gnd.n483 240.244
R13157 gnd.n6906 gnd.n483 240.244
R13158 gnd.n6906 gnd.n479 240.244
R13159 gnd.n6912 gnd.n479 240.244
R13160 gnd.n6912 gnd.n477 240.244
R13161 gnd.n6916 gnd.n477 240.244
R13162 gnd.n6916 gnd.n473 240.244
R13163 gnd.n6922 gnd.n473 240.244
R13164 gnd.n6922 gnd.n471 240.244
R13165 gnd.n6926 gnd.n471 240.244
R13166 gnd.n6926 gnd.n467 240.244
R13167 gnd.n6932 gnd.n467 240.244
R13168 gnd.n6932 gnd.n465 240.244
R13169 gnd.n6936 gnd.n465 240.244
R13170 gnd.n6936 gnd.n461 240.244
R13171 gnd.n6942 gnd.n461 240.244
R13172 gnd.n6942 gnd.n459 240.244
R13173 gnd.n6946 gnd.n459 240.244
R13174 gnd.n6946 gnd.n455 240.244
R13175 gnd.n6952 gnd.n455 240.244
R13176 gnd.n6952 gnd.n453 240.244
R13177 gnd.n6956 gnd.n453 240.244
R13178 gnd.n6956 gnd.n449 240.244
R13179 gnd.n6962 gnd.n449 240.244
R13180 gnd.n6962 gnd.n447 240.244
R13181 gnd.n6966 gnd.n447 240.244
R13182 gnd.n6966 gnd.n443 240.244
R13183 gnd.n6972 gnd.n443 240.244
R13184 gnd.n6972 gnd.n441 240.244
R13185 gnd.n6976 gnd.n441 240.244
R13186 gnd.n6976 gnd.n437 240.244
R13187 gnd.n6982 gnd.n437 240.244
R13188 gnd.n6982 gnd.n435 240.244
R13189 gnd.n6986 gnd.n435 240.244
R13190 gnd.n6986 gnd.n431 240.244
R13191 gnd.n6992 gnd.n431 240.244
R13192 gnd.n6992 gnd.n429 240.244
R13193 gnd.n6996 gnd.n429 240.244
R13194 gnd.n6996 gnd.n425 240.244
R13195 gnd.n7002 gnd.n425 240.244
R13196 gnd.n7002 gnd.n423 240.244
R13197 gnd.n7006 gnd.n423 240.244
R13198 gnd.n7006 gnd.n419 240.244
R13199 gnd.n7012 gnd.n419 240.244
R13200 gnd.n7012 gnd.n417 240.244
R13201 gnd.n7017 gnd.n417 240.244
R13202 gnd.n7017 gnd.n413 240.244
R13203 gnd.n7024 gnd.n413 240.244
R13204 gnd.n4869 gnd.n4868 240.244
R13205 gnd.n4870 gnd.n4869 240.244
R13206 gnd.n4870 gnd.n4566 240.244
R13207 gnd.n4900 gnd.n4566 240.244
R13208 gnd.n4900 gnd.n4567 240.244
R13209 gnd.n4896 gnd.n4567 240.244
R13210 gnd.n4896 gnd.n4895 240.244
R13211 gnd.n4895 gnd.n4894 240.244
R13212 gnd.n4894 gnd.n4878 240.244
R13213 gnd.n4890 gnd.n4878 240.244
R13214 gnd.n4890 gnd.n4889 240.244
R13215 gnd.n4889 gnd.n4888 240.244
R13216 gnd.n4888 gnd.n844 240.244
R13217 gnd.n6398 gnd.n844 240.244
R13218 gnd.n6398 gnd.n845 240.244
R13219 gnd.n6394 gnd.n845 240.244
R13220 gnd.n6394 gnd.n851 240.244
R13221 gnd.n6390 gnd.n851 240.244
R13222 gnd.n6390 gnd.n854 240.244
R13223 gnd.n6386 gnd.n854 240.244
R13224 gnd.n6386 gnd.n860 240.244
R13225 gnd.n5016 gnd.n860 240.244
R13226 gnd.n5022 gnd.n5016 240.244
R13227 gnd.n5022 gnd.n2060 240.244
R13228 gnd.n5034 gnd.n2060 240.244
R13229 gnd.n5034 gnd.n2056 240.244
R13230 gnd.n5040 gnd.n2056 240.244
R13231 gnd.n5040 gnd.n2049 240.244
R13232 gnd.n5051 gnd.n2049 240.244
R13233 gnd.n5051 gnd.n2045 240.244
R13234 gnd.n5057 gnd.n2045 240.244
R13235 gnd.n5057 gnd.n2037 240.244
R13236 gnd.n5068 gnd.n2037 240.244
R13237 gnd.n5068 gnd.n2032 240.244
R13238 gnd.n5076 gnd.n2032 240.244
R13239 gnd.n5076 gnd.n2033 240.244
R13240 gnd.n2033 gnd.n1627 240.244
R13241 gnd.n5161 gnd.n1627 240.244
R13242 gnd.n5161 gnd.n1622 240.244
R13243 gnd.n5178 gnd.n1622 240.244
R13244 gnd.n5178 gnd.n1623 240.244
R13245 gnd.n5174 gnd.n1623 240.244
R13246 gnd.n5174 gnd.n5173 240.244
R13247 gnd.n5173 gnd.n5172 240.244
R13248 gnd.n5172 gnd.n1588 240.244
R13249 gnd.n5220 gnd.n1588 240.244
R13250 gnd.n5220 gnd.n1584 240.244
R13251 gnd.n5226 gnd.n1584 240.244
R13252 gnd.n5226 gnd.n1566 240.244
R13253 gnd.n5250 gnd.n1566 240.244
R13254 gnd.n5250 gnd.n1562 240.244
R13255 gnd.n5256 gnd.n1562 240.244
R13256 gnd.n5256 gnd.n1549 240.244
R13257 gnd.n5277 gnd.n1549 240.244
R13258 gnd.n5277 gnd.n1545 240.244
R13259 gnd.n5283 gnd.n1545 240.244
R13260 gnd.n5283 gnd.n1529 240.244
R13261 gnd.n5301 gnd.n1529 240.244
R13262 gnd.n5301 gnd.n1524 240.244
R13263 gnd.n5309 gnd.n1524 240.244
R13264 gnd.n5309 gnd.n1525 240.244
R13265 gnd.n1525 gnd.n1502 240.244
R13266 gnd.n5359 gnd.n1502 240.244
R13267 gnd.n5359 gnd.n1497 240.244
R13268 gnd.n5367 gnd.n1497 240.244
R13269 gnd.n5367 gnd.n1498 240.244
R13270 gnd.n1498 gnd.n1480 240.244
R13271 gnd.n5399 gnd.n1480 240.244
R13272 gnd.n5399 gnd.n1475 240.244
R13273 gnd.n5407 gnd.n1475 240.244
R13274 gnd.n5407 gnd.n1476 240.244
R13275 gnd.n1476 gnd.n1451 240.244
R13276 gnd.n5456 gnd.n1451 240.244
R13277 gnd.n5456 gnd.n1446 240.244
R13278 gnd.n5464 gnd.n1446 240.244
R13279 gnd.n5464 gnd.n1447 240.244
R13280 gnd.n1447 gnd.n1430 240.244
R13281 gnd.n5494 gnd.n1430 240.244
R13282 gnd.n5494 gnd.n1426 240.244
R13283 gnd.n5500 gnd.n1426 240.244
R13284 gnd.n5500 gnd.n1401 240.244
R13285 gnd.n5532 gnd.n1401 240.244
R13286 gnd.n5532 gnd.n1396 240.244
R13287 gnd.n5540 gnd.n1396 240.244
R13288 gnd.n5540 gnd.n1397 240.244
R13289 gnd.n1397 gnd.n1375 240.244
R13290 gnd.n5576 gnd.n1375 240.244
R13291 gnd.n5576 gnd.n1371 240.244
R13292 gnd.n5583 gnd.n1371 240.244
R13293 gnd.n5583 gnd.n1349 240.244
R13294 gnd.n5619 gnd.n1349 240.244
R13295 gnd.n5619 gnd.n1350 240.244
R13296 gnd.n5615 gnd.n1350 240.244
R13297 gnd.n5615 gnd.n1360 240.244
R13298 gnd.n1360 gnd.n1359 240.244
R13299 gnd.n1359 gnd.n1320 240.244
R13300 gnd.n5663 gnd.n1320 240.244
R13301 gnd.n5663 gnd.n1316 240.244
R13302 gnd.n5669 gnd.n1316 240.244
R13303 gnd.n5669 gnd.n1225 240.244
R13304 gnd.n5811 gnd.n1225 240.244
R13305 gnd.n5811 gnd.n1221 240.244
R13306 gnd.n5817 gnd.n1221 240.244
R13307 gnd.n5817 gnd.n1213 240.244
R13308 gnd.n5828 gnd.n1213 240.244
R13309 gnd.n5828 gnd.n1209 240.244
R13310 gnd.n5834 gnd.n1209 240.244
R13311 gnd.n5834 gnd.n1201 240.244
R13312 gnd.n5845 gnd.n1201 240.244
R13313 gnd.n5845 gnd.n1197 240.244
R13314 gnd.n5851 gnd.n1197 240.244
R13315 gnd.n5851 gnd.n1189 240.244
R13316 gnd.n5863 gnd.n1189 240.244
R13317 gnd.n5863 gnd.n1185 240.244
R13318 gnd.n5869 gnd.n1185 240.244
R13319 gnd.n5869 gnd.n1178 240.244
R13320 gnd.n5880 gnd.n1178 240.244
R13321 gnd.n5880 gnd.n1174 240.244
R13322 gnd.n5888 gnd.n1174 240.244
R13323 gnd.n5888 gnd.n1165 240.244
R13324 gnd.n5916 gnd.n1165 240.244
R13325 gnd.n5917 gnd.n5916 240.244
R13326 gnd.n5917 gnd.n1161 240.244
R13327 gnd.n5924 gnd.n1161 240.244
R13328 gnd.n5925 gnd.n5924 240.244
R13329 gnd.n5926 gnd.n5925 240.244
R13330 gnd.n5926 gnd.n1156 240.244
R13331 gnd.n6008 gnd.n1156 240.244
R13332 gnd.n6008 gnd.n1157 240.244
R13333 gnd.n6004 gnd.n1157 240.244
R13334 gnd.n6004 gnd.n5934 240.244
R13335 gnd.n5948 gnd.n5934 240.244
R13336 gnd.n5948 gnd.n400 240.244
R13337 gnd.n7036 gnd.n400 240.244
R13338 gnd.n7036 gnd.n401 240.244
R13339 gnd.n7032 gnd.n401 240.244
R13340 gnd.n7032 gnd.n7031 240.244
R13341 gnd.n7031 gnd.n7030 240.244
R13342 gnd.n7030 gnd.n407 240.244
R13343 gnd.n7026 gnd.n407 240.244
R13344 gnd.n7026 gnd.n7025 240.244
R13345 gnd.n4659 gnd.n4658 240.244
R13346 gnd.n4661 gnd.n4659 240.244
R13347 gnd.n4667 gnd.n4650 240.244
R13348 gnd.n4671 gnd.n4669 240.244
R13349 gnd.n4677 gnd.n4646 240.244
R13350 gnd.n4681 gnd.n4679 240.244
R13351 gnd.n4687 gnd.n4642 240.244
R13352 gnd.n4691 gnd.n4689 240.244
R13353 gnd.n4697 gnd.n4638 240.244
R13354 gnd.n4701 gnd.n4699 240.244
R13355 gnd.n4707 gnd.n4634 240.244
R13356 gnd.n4711 gnd.n4709 240.244
R13357 gnd.n4717 gnd.n4630 240.244
R13358 gnd.n4721 gnd.n4719 240.244
R13359 gnd.n4727 gnd.n4626 240.244
R13360 gnd.n4731 gnd.n4729 240.244
R13361 gnd.n4737 gnd.n4622 240.244
R13362 gnd.n4741 gnd.n4739 240.244
R13363 gnd.n4747 gnd.n4618 240.244
R13364 gnd.n4751 gnd.n4749 240.244
R13365 gnd.n4757 gnd.n4614 240.244
R13366 gnd.n4761 gnd.n4759 240.244
R13367 gnd.n4767 gnd.n4610 240.244
R13368 gnd.n4771 gnd.n4769 240.244
R13369 gnd.n4777 gnd.n4606 240.244
R13370 gnd.n4781 gnd.n4779 240.244
R13371 gnd.n4787 gnd.n4602 240.244
R13372 gnd.n4791 gnd.n4789 240.244
R13373 gnd.n4797 gnd.n4598 240.244
R13374 gnd.n4801 gnd.n4799 240.244
R13375 gnd.n4807 gnd.n4594 240.244
R13376 gnd.n4811 gnd.n4809 240.244
R13377 gnd.n4817 gnd.n4590 240.244
R13378 gnd.n4821 gnd.n4819 240.244
R13379 gnd.n4827 gnd.n4586 240.244
R13380 gnd.n4831 gnd.n4829 240.244
R13381 gnd.n4837 gnd.n4582 240.244
R13382 gnd.n4841 gnd.n4839 240.244
R13383 gnd.n4847 gnd.n4578 240.244
R13384 gnd.n4851 gnd.n4849 240.244
R13385 gnd.n4858 gnd.n4574 240.244
R13386 gnd.n4862 gnd.n4860 240.244
R13387 gnd.n1784 gnd.n1782 240.244
R13388 gnd.n1790 gnd.n1777 240.244
R13389 gnd.n1794 gnd.n1792 240.244
R13390 gnd.n1800 gnd.n1773 240.244
R13391 gnd.n1804 gnd.n1802 240.244
R13392 gnd.n1810 gnd.n1769 240.244
R13393 gnd.n1814 gnd.n1812 240.244
R13394 gnd.n1820 gnd.n1765 240.244
R13395 gnd.n1823 gnd.n1822 240.244
R13396 gnd.n1829 gnd.n1828 240.244
R13397 gnd.n1832 gnd.n1831 240.244
R13398 gnd.n1839 gnd.n1838 240.244
R13399 gnd.n1843 gnd.n1842 240.244
R13400 gnd.n1947 gnd.n1850 240.244
R13401 gnd.n1945 gnd.n1944 240.244
R13402 gnd.n1942 gnd.n1852 240.244
R13403 gnd.n1938 gnd.n1937 240.244
R13404 gnd.n1935 gnd.n1859 240.244
R13405 gnd.n1928 gnd.n1868 240.244
R13406 gnd.n1926 gnd.n1925 240.244
R13407 gnd.n1923 gnd.n1870 240.244
R13408 gnd.n1919 gnd.n1918 240.244
R13409 gnd.n1916 gnd.n1877 240.244
R13410 gnd.n1912 gnd.n1911 240.244
R13411 gnd.n1909 gnd.n1884 240.244
R13412 gnd.n1905 gnd.n1904 240.244
R13413 gnd.n1902 gnd.n1891 240.244
R13414 gnd.n1898 gnd.n1897 240.244
R13415 gnd.n3907 gnd.n2405 240.244
R13416 gnd.n4271 gnd.n2405 240.244
R13417 gnd.n4272 gnd.n4271 240.244
R13418 gnd.n4272 gnd.n2397 240.244
R13419 gnd.n2397 gnd.n2387 240.244
R13420 gnd.n4291 gnd.n2387 240.244
R13421 gnd.n4292 gnd.n4291 240.244
R13422 gnd.n4292 gnd.n2378 240.244
R13423 gnd.n2378 gnd.n2369 240.244
R13424 gnd.n4311 gnd.n2369 240.244
R13425 gnd.n4312 gnd.n4311 240.244
R13426 gnd.n4312 gnd.n2361 240.244
R13427 gnd.n2361 gnd.n2351 240.244
R13428 gnd.n4331 gnd.n2351 240.244
R13429 gnd.n4332 gnd.n4331 240.244
R13430 gnd.n4332 gnd.n2342 240.244
R13431 gnd.n2342 gnd.n2333 240.244
R13432 gnd.n4351 gnd.n2333 240.244
R13433 gnd.n4352 gnd.n4351 240.244
R13434 gnd.n4352 gnd.n2325 240.244
R13435 gnd.n2325 gnd.n2315 240.244
R13436 gnd.n4371 gnd.n2315 240.244
R13437 gnd.n4372 gnd.n4371 240.244
R13438 gnd.n4372 gnd.n2305 240.244
R13439 gnd.n4375 gnd.n2305 240.244
R13440 gnd.n4375 gnd.n2296 240.244
R13441 gnd.n2296 gnd.n2289 240.244
R13442 gnd.n4407 gnd.n2289 240.244
R13443 gnd.n4407 gnd.n2279 240.244
R13444 gnd.n4410 gnd.n2279 240.244
R13445 gnd.n4410 gnd.n2271 240.244
R13446 gnd.n2271 gnd.n2263 240.244
R13447 gnd.n4441 gnd.n2263 240.244
R13448 gnd.n4441 gnd.n2253 240.244
R13449 gnd.n4444 gnd.n2253 240.244
R13450 gnd.n4444 gnd.n2245 240.244
R13451 gnd.n2245 gnd.n2237 240.244
R13452 gnd.n4475 gnd.n2237 240.244
R13453 gnd.n4475 gnd.n2228 240.244
R13454 gnd.n4478 gnd.n2228 240.244
R13455 gnd.n4478 gnd.n2220 240.244
R13456 gnd.n2220 gnd.n2211 240.244
R13457 gnd.n4509 gnd.n2211 240.244
R13458 gnd.n4509 gnd.n2202 240.244
R13459 gnd.n4512 gnd.n2202 240.244
R13460 gnd.n4512 gnd.n2194 240.244
R13461 gnd.n4516 gnd.n2194 240.244
R13462 gnd.n4516 gnd.n2186 240.244
R13463 gnd.n2186 gnd.n754 240.244
R13464 gnd.n4553 gnd.n754 240.244
R13465 gnd.n4553 gnd.n766 240.244
R13466 gnd.n4557 gnd.n766 240.244
R13467 gnd.n4557 gnd.n778 240.244
R13468 gnd.n4903 gnd.n778 240.244
R13469 gnd.n4903 gnd.n788 240.244
R13470 gnd.n4907 gnd.n788 240.244
R13471 gnd.n4907 gnd.n798 240.244
R13472 gnd.n4917 gnd.n798 240.244
R13473 gnd.n4917 gnd.n809 240.244
R13474 gnd.n4927 gnd.n809 240.244
R13475 gnd.n4927 gnd.n819 240.244
R13476 gnd.n4923 gnd.n819 240.244
R13477 gnd.n4923 gnd.n830 240.244
R13478 gnd.n6401 gnd.n830 240.244
R13479 gnd.n3976 gnd.n3972 240.244
R13480 gnd.n3982 gnd.n3972 240.244
R13481 gnd.n3986 gnd.n3984 240.244
R13482 gnd.n3992 gnd.n3968 240.244
R13483 gnd.n3996 gnd.n3994 240.244
R13484 gnd.n4002 gnd.n3964 240.244
R13485 gnd.n4006 gnd.n4004 240.244
R13486 gnd.n4012 gnd.n3960 240.244
R13487 gnd.n4016 gnd.n4014 240.244
R13488 gnd.n4022 gnd.n3953 240.244
R13489 gnd.n4026 gnd.n4024 240.244
R13490 gnd.n4032 gnd.n3949 240.244
R13491 gnd.n4036 gnd.n4034 240.244
R13492 gnd.n4042 gnd.n3945 240.244
R13493 gnd.n4046 gnd.n4044 240.244
R13494 gnd.n4052 gnd.n3941 240.244
R13495 gnd.n4056 gnd.n4054 240.244
R13496 gnd.n4062 gnd.n3937 240.244
R13497 gnd.n4066 gnd.n4064 240.244
R13498 gnd.n4074 gnd.n3933 240.244
R13499 gnd.n4078 gnd.n4076 240.244
R13500 gnd.n4084 gnd.n3929 240.244
R13501 gnd.n4088 gnd.n4086 240.244
R13502 gnd.n4094 gnd.n3925 240.244
R13503 gnd.n4098 gnd.n4096 240.244
R13504 gnd.n4104 gnd.n3921 240.244
R13505 gnd.n4108 gnd.n4106 240.244
R13506 gnd.n4115 gnd.n3917 240.244
R13507 gnd.n4118 gnd.n4117 240.244
R13508 gnd.n4263 gnd.n2408 240.244
R13509 gnd.n4269 gnd.n2408 240.244
R13510 gnd.n4269 gnd.n2395 240.244
R13511 gnd.n4283 gnd.n2395 240.244
R13512 gnd.n4283 gnd.n2391 240.244
R13513 gnd.n4289 gnd.n2391 240.244
R13514 gnd.n4289 gnd.n2376 240.244
R13515 gnd.n4303 gnd.n2376 240.244
R13516 gnd.n4303 gnd.n2372 240.244
R13517 gnd.n4309 gnd.n2372 240.244
R13518 gnd.n4309 gnd.n2359 240.244
R13519 gnd.n4323 gnd.n2359 240.244
R13520 gnd.n4323 gnd.n2355 240.244
R13521 gnd.n4329 gnd.n2355 240.244
R13522 gnd.n4329 gnd.n2340 240.244
R13523 gnd.n4343 gnd.n2340 240.244
R13524 gnd.n4343 gnd.n2336 240.244
R13525 gnd.n4349 gnd.n2336 240.244
R13526 gnd.n4349 gnd.n2323 240.244
R13527 gnd.n4363 gnd.n2323 240.244
R13528 gnd.n4363 gnd.n2319 240.244
R13529 gnd.n4369 gnd.n2319 240.244
R13530 gnd.n4369 gnd.n2303 240.244
R13531 gnd.n4387 gnd.n2303 240.244
R13532 gnd.n4387 gnd.n2298 240.244
R13533 gnd.n4395 gnd.n2298 240.244
R13534 gnd.n4395 gnd.n2299 240.244
R13535 gnd.n2299 gnd.n2278 240.244
R13536 gnd.n4422 gnd.n2278 240.244
R13537 gnd.n4422 gnd.n2273 240.244
R13538 gnd.n4430 gnd.n2273 240.244
R13539 gnd.n4430 gnd.n2274 240.244
R13540 gnd.n2274 gnd.n2252 240.244
R13541 gnd.n4456 gnd.n2252 240.244
R13542 gnd.n4456 gnd.n2247 240.244
R13543 gnd.n4464 gnd.n2247 240.244
R13544 gnd.n4464 gnd.n2248 240.244
R13545 gnd.n2248 gnd.n2227 240.244
R13546 gnd.n4490 gnd.n2227 240.244
R13547 gnd.n4490 gnd.n2222 240.244
R13548 gnd.n4498 gnd.n2222 240.244
R13549 gnd.n4498 gnd.n2223 240.244
R13550 gnd.n2223 gnd.n2201 240.244
R13551 gnd.n4525 gnd.n2201 240.244
R13552 gnd.n4525 gnd.n2196 240.244
R13553 gnd.n4534 gnd.n2196 240.244
R13554 gnd.n4534 gnd.n2197 240.244
R13555 gnd.n2197 gnd.n757 240.244
R13556 gnd.n6451 gnd.n757 240.244
R13557 gnd.n6451 gnd.n758 240.244
R13558 gnd.n6447 gnd.n758 240.244
R13559 gnd.n6447 gnd.n764 240.244
R13560 gnd.n6439 gnd.n764 240.244
R13561 gnd.n6439 gnd.n781 240.244
R13562 gnd.n6435 gnd.n781 240.244
R13563 gnd.n6435 gnd.n787 240.244
R13564 gnd.n6427 gnd.n787 240.244
R13565 gnd.n6427 gnd.n801 240.244
R13566 gnd.n6423 gnd.n801 240.244
R13567 gnd.n6423 gnd.n807 240.244
R13568 gnd.n6415 gnd.n807 240.244
R13569 gnd.n6415 gnd.n822 240.244
R13570 gnd.n6411 gnd.n822 240.244
R13571 gnd.n6411 gnd.n828 240.244
R13572 gnd.n3904 gnd.n2436 240.244
R13573 gnd.n3897 gnd.n3896 240.244
R13574 gnd.n3894 gnd.n3893 240.244
R13575 gnd.n3890 gnd.n3889 240.244
R13576 gnd.n3886 gnd.n3885 240.244
R13577 gnd.n3882 gnd.n3881 240.244
R13578 gnd.n3878 gnd.n3877 240.244
R13579 gnd.n3874 gnd.n3873 240.244
R13580 gnd.n3148 gnd.n2860 240.244
R13581 gnd.n3158 gnd.n2860 240.244
R13582 gnd.n3158 gnd.n2851 240.244
R13583 gnd.n2851 gnd.n2840 240.244
R13584 gnd.n3179 gnd.n2840 240.244
R13585 gnd.n3179 gnd.n2834 240.244
R13586 gnd.n3189 gnd.n2834 240.244
R13587 gnd.n3189 gnd.n2823 240.244
R13588 gnd.n2823 gnd.n2815 240.244
R13589 gnd.n3207 gnd.n2815 240.244
R13590 gnd.n3208 gnd.n3207 240.244
R13591 gnd.n3208 gnd.n2800 240.244
R13592 gnd.n3210 gnd.n2800 240.244
R13593 gnd.n3210 gnd.n2786 240.244
R13594 gnd.n3252 gnd.n2786 240.244
R13595 gnd.n3253 gnd.n3252 240.244
R13596 gnd.n3256 gnd.n3253 240.244
R13597 gnd.n3256 gnd.n2741 240.244
R13598 gnd.n2781 gnd.n2741 240.244
R13599 gnd.n2781 gnd.n2751 240.244
R13600 gnd.n3266 gnd.n2751 240.244
R13601 gnd.n3266 gnd.n2772 240.244
R13602 gnd.n3276 gnd.n2772 240.244
R13603 gnd.n3276 gnd.n2638 240.244
R13604 gnd.n3321 gnd.n2638 240.244
R13605 gnd.n3321 gnd.n2624 240.244
R13606 gnd.n3343 gnd.n2624 240.244
R13607 gnd.n3344 gnd.n3343 240.244
R13608 gnd.n3344 gnd.n2611 240.244
R13609 gnd.n2611 gnd.n2600 240.244
R13610 gnd.n3375 gnd.n2600 240.244
R13611 gnd.n3376 gnd.n3375 240.244
R13612 gnd.n3377 gnd.n3376 240.244
R13613 gnd.n3377 gnd.n2585 240.244
R13614 gnd.n2585 gnd.n2584 240.244
R13615 gnd.n2584 gnd.n2569 240.244
R13616 gnd.n3428 gnd.n2569 240.244
R13617 gnd.n3429 gnd.n3428 240.244
R13618 gnd.n3429 gnd.n2556 240.244
R13619 gnd.n2556 gnd.n2545 240.244
R13620 gnd.n3460 gnd.n2545 240.244
R13621 gnd.n3461 gnd.n3460 240.244
R13622 gnd.n3462 gnd.n3461 240.244
R13623 gnd.n3462 gnd.n2529 240.244
R13624 gnd.n2529 gnd.n2528 240.244
R13625 gnd.n2528 gnd.n2515 240.244
R13626 gnd.n3517 gnd.n2515 240.244
R13627 gnd.n3518 gnd.n3517 240.244
R13628 gnd.n3518 gnd.n2502 240.244
R13629 gnd.n2502 gnd.n2492 240.244
R13630 gnd.n3805 gnd.n2492 240.244
R13631 gnd.n3808 gnd.n3805 240.244
R13632 gnd.n3808 gnd.n3807 240.244
R13633 gnd.n3138 gnd.n2873 240.244
R13634 gnd.n2894 gnd.n2873 240.244
R13635 gnd.n2897 gnd.n2896 240.244
R13636 gnd.n2904 gnd.n2903 240.244
R13637 gnd.n2907 gnd.n2906 240.244
R13638 gnd.n2914 gnd.n2913 240.244
R13639 gnd.n2917 gnd.n2916 240.244
R13640 gnd.n2924 gnd.n2923 240.244
R13641 gnd.n3146 gnd.n2870 240.244
R13642 gnd.n2870 gnd.n2849 240.244
R13643 gnd.n3169 gnd.n2849 240.244
R13644 gnd.n3169 gnd.n2843 240.244
R13645 gnd.n3177 gnd.n2843 240.244
R13646 gnd.n3177 gnd.n2845 240.244
R13647 gnd.n2845 gnd.n2821 240.244
R13648 gnd.n3199 gnd.n2821 240.244
R13649 gnd.n3199 gnd.n2817 240.244
R13650 gnd.n3205 gnd.n2817 240.244
R13651 gnd.n3205 gnd.n2799 240.244
R13652 gnd.n3230 gnd.n2799 240.244
R13653 gnd.n3230 gnd.n2794 240.244
R13654 gnd.n3242 gnd.n2794 240.244
R13655 gnd.n3242 gnd.n2795 240.244
R13656 gnd.n3238 gnd.n2795 240.244
R13657 gnd.n3238 gnd.n2743 240.244
R13658 gnd.n3290 gnd.n2743 240.244
R13659 gnd.n3290 gnd.n2744 240.244
R13660 gnd.n3286 gnd.n2744 240.244
R13661 gnd.n3286 gnd.n2750 240.244
R13662 gnd.n2770 gnd.n2750 240.244
R13663 gnd.n2770 gnd.n2636 240.244
R13664 gnd.n3325 gnd.n2636 240.244
R13665 gnd.n3325 gnd.n2631 240.244
R13666 gnd.n3333 gnd.n2631 240.244
R13667 gnd.n3333 gnd.n2632 240.244
R13668 gnd.n2632 gnd.n2609 240.244
R13669 gnd.n3365 gnd.n2609 240.244
R13670 gnd.n3365 gnd.n2604 240.244
R13671 gnd.n3373 gnd.n2604 240.244
R13672 gnd.n3373 gnd.n2605 240.244
R13673 gnd.n2605 gnd.n2582 240.244
R13674 gnd.n3410 gnd.n2582 240.244
R13675 gnd.n3410 gnd.n2577 240.244
R13676 gnd.n3418 gnd.n2577 240.244
R13677 gnd.n3418 gnd.n2578 240.244
R13678 gnd.n2578 gnd.n2554 240.244
R13679 gnd.n3450 gnd.n2554 240.244
R13680 gnd.n3450 gnd.n2549 240.244
R13681 gnd.n3458 gnd.n2549 240.244
R13682 gnd.n3458 gnd.n2550 240.244
R13683 gnd.n2550 gnd.n2527 240.244
R13684 gnd.n3499 gnd.n2527 240.244
R13685 gnd.n3499 gnd.n2522 240.244
R13686 gnd.n3507 gnd.n2522 240.244
R13687 gnd.n3507 gnd.n2523 240.244
R13688 gnd.n2523 gnd.n2500 240.244
R13689 gnd.n3793 gnd.n2500 240.244
R13690 gnd.n3793 gnd.n2495 240.244
R13691 gnd.n3803 gnd.n2495 240.244
R13692 gnd.n3803 gnd.n2496 240.244
R13693 gnd.n2496 gnd.n2435 240.244
R13694 gnd.n2455 gnd.n2413 240.244
R13695 gnd.n3864 gnd.n3863 240.244
R13696 gnd.n3860 gnd.n3859 240.244
R13697 gnd.n3856 gnd.n3855 240.244
R13698 gnd.n3852 gnd.n3851 240.244
R13699 gnd.n3848 gnd.n3847 240.244
R13700 gnd.n3844 gnd.n3843 240.244
R13701 gnd.n3840 gnd.n3839 240.244
R13702 gnd.n3836 gnd.n3835 240.244
R13703 gnd.n3832 gnd.n3831 240.244
R13704 gnd.n3828 gnd.n3827 240.244
R13705 gnd.n3824 gnd.n3823 240.244
R13706 gnd.n3820 gnd.n3819 240.244
R13707 gnd.n3061 gnd.n2958 240.244
R13708 gnd.n3061 gnd.n2951 240.244
R13709 gnd.n3072 gnd.n2951 240.244
R13710 gnd.n3072 gnd.n2947 240.244
R13711 gnd.n3078 gnd.n2947 240.244
R13712 gnd.n3078 gnd.n2939 240.244
R13713 gnd.n3088 gnd.n2939 240.244
R13714 gnd.n3088 gnd.n2934 240.244
R13715 gnd.n3124 gnd.n2934 240.244
R13716 gnd.n3124 gnd.n2935 240.244
R13717 gnd.n2935 gnd.n2882 240.244
R13718 gnd.n3119 gnd.n2882 240.244
R13719 gnd.n3119 gnd.n3118 240.244
R13720 gnd.n3118 gnd.n2861 240.244
R13721 gnd.n3114 gnd.n2861 240.244
R13722 gnd.n3114 gnd.n2852 240.244
R13723 gnd.n3111 gnd.n2852 240.244
R13724 gnd.n3111 gnd.n3110 240.244
R13725 gnd.n3110 gnd.n2835 240.244
R13726 gnd.n3106 gnd.n2835 240.244
R13727 gnd.n3106 gnd.n2824 240.244
R13728 gnd.n2824 gnd.n2805 240.244
R13729 gnd.n3219 gnd.n2805 240.244
R13730 gnd.n3219 gnd.n2801 240.244
R13731 gnd.n3227 gnd.n2801 240.244
R13732 gnd.n3227 gnd.n2792 240.244
R13733 gnd.n2792 gnd.n2728 240.244
R13734 gnd.n3299 gnd.n2728 240.244
R13735 gnd.n3299 gnd.n2729 240.244
R13736 gnd.n2740 gnd.n2729 240.244
R13737 gnd.n2775 gnd.n2740 240.244
R13738 gnd.n2778 gnd.n2775 240.244
R13739 gnd.n2778 gnd.n2752 240.244
R13740 gnd.n2765 gnd.n2752 240.244
R13741 gnd.n2765 gnd.n2762 240.244
R13742 gnd.n2762 gnd.n2639 240.244
R13743 gnd.n3320 gnd.n2639 240.244
R13744 gnd.n3320 gnd.n2629 240.244
R13745 gnd.n3316 gnd.n2629 240.244
R13746 gnd.n3316 gnd.n2623 240.244
R13747 gnd.n3313 gnd.n2623 240.244
R13748 gnd.n3313 gnd.n2612 240.244
R13749 gnd.n3310 gnd.n2612 240.244
R13750 gnd.n3310 gnd.n2590 240.244
R13751 gnd.n3386 gnd.n2590 240.244
R13752 gnd.n3386 gnd.n2586 240.244
R13753 gnd.n3407 gnd.n2586 240.244
R13754 gnd.n3407 gnd.n2575 240.244
R13755 gnd.n3403 gnd.n2575 240.244
R13756 gnd.n3403 gnd.n2568 240.244
R13757 gnd.n3400 gnd.n2568 240.244
R13758 gnd.n3400 gnd.n2557 240.244
R13759 gnd.n3397 gnd.n2557 240.244
R13760 gnd.n3397 gnd.n2534 240.244
R13761 gnd.n3471 gnd.n2534 240.244
R13762 gnd.n3471 gnd.n2530 240.244
R13763 gnd.n3496 gnd.n2530 240.244
R13764 gnd.n3496 gnd.n2521 240.244
R13765 gnd.n3492 gnd.n2521 240.244
R13766 gnd.n3492 gnd.n2514 240.244
R13767 gnd.n3488 gnd.n2514 240.244
R13768 gnd.n3488 gnd.n2503 240.244
R13769 gnd.n3485 gnd.n2503 240.244
R13770 gnd.n3485 gnd.n2484 240.244
R13771 gnd.n3815 gnd.n2484 240.244
R13772 gnd.n2975 gnd.n2974 240.244
R13773 gnd.n3046 gnd.n2974 240.244
R13774 gnd.n3044 gnd.n3043 240.244
R13775 gnd.n3040 gnd.n3039 240.244
R13776 gnd.n3036 gnd.n3035 240.244
R13777 gnd.n3032 gnd.n3031 240.244
R13778 gnd.n3028 gnd.n3027 240.244
R13779 gnd.n3024 gnd.n3023 240.244
R13780 gnd.n3020 gnd.n3019 240.244
R13781 gnd.n3016 gnd.n3015 240.244
R13782 gnd.n3012 gnd.n3011 240.244
R13783 gnd.n3008 gnd.n3007 240.244
R13784 gnd.n3004 gnd.n2962 240.244
R13785 gnd.n3064 gnd.n2956 240.244
R13786 gnd.n3064 gnd.n2952 240.244
R13787 gnd.n3070 gnd.n2952 240.244
R13788 gnd.n3070 gnd.n2945 240.244
R13789 gnd.n3080 gnd.n2945 240.244
R13790 gnd.n3080 gnd.n2941 240.244
R13791 gnd.n3086 gnd.n2941 240.244
R13792 gnd.n3086 gnd.n2932 240.244
R13793 gnd.n3126 gnd.n2932 240.244
R13794 gnd.n3126 gnd.n2883 240.244
R13795 gnd.n3134 gnd.n2883 240.244
R13796 gnd.n3134 gnd.n2884 240.244
R13797 gnd.n2884 gnd.n2862 240.244
R13798 gnd.n3155 gnd.n2862 240.244
R13799 gnd.n3155 gnd.n2854 240.244
R13800 gnd.n3166 gnd.n2854 240.244
R13801 gnd.n3166 gnd.n2855 240.244
R13802 gnd.n2855 gnd.n2836 240.244
R13803 gnd.n3186 gnd.n2836 240.244
R13804 gnd.n3186 gnd.n2826 240.244
R13805 gnd.n3196 gnd.n2826 240.244
R13806 gnd.n3196 gnd.n2807 240.244
R13807 gnd.n3217 gnd.n2807 240.244
R13808 gnd.n3217 gnd.n2809 240.244
R13809 gnd.n2809 gnd.n2790 240.244
R13810 gnd.n3245 gnd.n2790 240.244
R13811 gnd.n3245 gnd.n2732 240.244
R13812 gnd.n3297 gnd.n2732 240.244
R13813 gnd.n3297 gnd.n2733 240.244
R13814 gnd.n3293 gnd.n2733 240.244
R13815 gnd.n3293 gnd.n2739 240.244
R13816 gnd.n2754 gnd.n2739 240.244
R13817 gnd.n3283 gnd.n2754 240.244
R13818 gnd.n3283 gnd.n2755 240.244
R13819 gnd.n3279 gnd.n2755 240.244
R13820 gnd.n3279 gnd.n2761 240.244
R13821 gnd.n2761 gnd.n2628 240.244
R13822 gnd.n3336 gnd.n2628 240.244
R13823 gnd.n3336 gnd.n2621 240.244
R13824 gnd.n3347 gnd.n2621 240.244
R13825 gnd.n3347 gnd.n2614 240.244
R13826 gnd.n3362 gnd.n2614 240.244
R13827 gnd.n3362 gnd.n2615 240.244
R13828 gnd.n2615 gnd.n2593 240.244
R13829 gnd.n3384 gnd.n2593 240.244
R13830 gnd.n3384 gnd.n2594 240.244
R13831 gnd.n2594 gnd.n2573 240.244
R13832 gnd.n3421 gnd.n2573 240.244
R13833 gnd.n3421 gnd.n2566 240.244
R13834 gnd.n3432 gnd.n2566 240.244
R13835 gnd.n3432 gnd.n2559 240.244
R13836 gnd.n3447 gnd.n2559 240.244
R13837 gnd.n3447 gnd.n2560 240.244
R13838 gnd.n2560 gnd.n2537 240.244
R13839 gnd.n3469 gnd.n2537 240.244
R13840 gnd.n3469 gnd.n2539 240.244
R13841 gnd.n2539 gnd.n2519 240.244
R13842 gnd.n3510 gnd.n2519 240.244
R13843 gnd.n3510 gnd.n2512 240.244
R13844 gnd.n3521 gnd.n2512 240.244
R13845 gnd.n3521 gnd.n2505 240.244
R13846 gnd.n3790 gnd.n2505 240.244
R13847 gnd.n3790 gnd.n2506 240.244
R13848 gnd.n2506 gnd.n2487 240.244
R13849 gnd.n3813 gnd.n2487 240.244
R13850 gnd.n2081 gnd.n2080 240.244
R13851 gnd.n2095 gnd.n2094 240.244
R13852 gnd.n2107 gnd.n2097 240.244
R13853 gnd.n2110 gnd.n2109 240.244
R13854 gnd.n2121 gnd.n2120 240.244
R13855 gnd.n2133 gnd.n2123 240.244
R13856 gnd.n2136 gnd.n2135 240.244
R13857 gnd.n2147 gnd.n2146 240.244
R13858 gnd.n4940 gnd.n2149 240.244
R13859 gnd.n4207 gnd.n3908 240.244
R13860 gnd.n4207 gnd.n2406 240.244
R13861 gnd.n4204 gnd.n2406 240.244
R13862 gnd.n4204 gnd.n2398 240.244
R13863 gnd.n4201 gnd.n2398 240.244
R13864 gnd.n4201 gnd.n2389 240.244
R13865 gnd.n4198 gnd.n2389 240.244
R13866 gnd.n4198 gnd.n2379 240.244
R13867 gnd.n4195 gnd.n2379 240.244
R13868 gnd.n4195 gnd.n2370 240.244
R13869 gnd.n4192 gnd.n2370 240.244
R13870 gnd.n4192 gnd.n2362 240.244
R13871 gnd.n4189 gnd.n2362 240.244
R13872 gnd.n4189 gnd.n2353 240.244
R13873 gnd.n4186 gnd.n2353 240.244
R13874 gnd.n4186 gnd.n2343 240.244
R13875 gnd.n4183 gnd.n2343 240.244
R13876 gnd.n4183 gnd.n2334 240.244
R13877 gnd.n4180 gnd.n2334 240.244
R13878 gnd.n4180 gnd.n2326 240.244
R13879 gnd.n4177 gnd.n2326 240.244
R13880 gnd.n4177 gnd.n2317 240.244
R13881 gnd.n4174 gnd.n2317 240.244
R13882 gnd.n4174 gnd.n2306 240.244
R13883 gnd.n2306 gnd.n2295 240.244
R13884 gnd.n4397 gnd.n2295 240.244
R13885 gnd.n4397 gnd.n2291 240.244
R13886 gnd.n4405 gnd.n2291 240.244
R13887 gnd.n4405 gnd.n2280 240.244
R13888 gnd.n2280 gnd.n2270 240.244
R13889 gnd.n4432 gnd.n2270 240.244
R13890 gnd.n4432 gnd.n2265 240.244
R13891 gnd.n4439 gnd.n2265 240.244
R13892 gnd.n4439 gnd.n2254 240.244
R13893 gnd.n2254 gnd.n2244 240.244
R13894 gnd.n4466 gnd.n2244 240.244
R13895 gnd.n4466 gnd.n2239 240.244
R13896 gnd.n4473 gnd.n2239 240.244
R13897 gnd.n4473 gnd.n2229 240.244
R13898 gnd.n2229 gnd.n2218 240.244
R13899 gnd.n4500 gnd.n2218 240.244
R13900 gnd.n4500 gnd.n2213 240.244
R13901 gnd.n4507 gnd.n2213 240.244
R13902 gnd.n4507 gnd.n2203 240.244
R13903 gnd.n2203 gnd.n2192 240.244
R13904 gnd.n4536 gnd.n2192 240.244
R13905 gnd.n4536 gnd.n2187 240.244
R13906 gnd.n4546 gnd.n2187 240.244
R13907 gnd.n4546 gnd.n755 240.244
R13908 gnd.n4540 gnd.n755 240.244
R13909 gnd.n4540 gnd.n767 240.244
R13910 gnd.n4559 gnd.n767 240.244
R13911 gnd.n4559 gnd.n779 240.244
R13912 gnd.n4565 gnd.n779 240.244
R13913 gnd.n4565 gnd.n789 240.244
R13914 gnd.n4909 gnd.n789 240.244
R13915 gnd.n4909 gnd.n799 240.244
R13916 gnd.n4915 gnd.n799 240.244
R13917 gnd.n4915 gnd.n810 240.244
R13918 gnd.n4929 gnd.n810 240.244
R13919 gnd.n4929 gnd.n820 240.244
R13920 gnd.n2168 gnd.n820 240.244
R13921 gnd.n2168 gnd.n831 240.244
R13922 gnd.n842 gnd.n831 240.244
R13923 gnd.n4248 gnd.n4246 240.244
R13924 gnd.n4244 gnd.n4125 240.244
R13925 gnd.n4240 gnd.n4238 240.244
R13926 gnd.n4236 gnd.n4131 240.244
R13927 gnd.n4232 gnd.n4230 240.244
R13928 gnd.n4228 gnd.n4137 240.244
R13929 gnd.n4224 gnd.n4222 240.244
R13930 gnd.n4220 gnd.n4143 240.244
R13931 gnd.n4213 gnd.n4212 240.244
R13932 gnd.n4261 gnd.n3911 240.244
R13933 gnd.n3911 gnd.n2407 240.244
R13934 gnd.n2407 gnd.n2399 240.244
R13935 gnd.n4281 gnd.n2399 240.244
R13936 gnd.n4281 gnd.n2400 240.244
R13937 gnd.n2400 gnd.n2390 240.244
R13938 gnd.n2390 gnd.n2381 240.244
R13939 gnd.n4301 gnd.n2381 240.244
R13940 gnd.n4301 gnd.n2382 240.244
R13941 gnd.n2382 gnd.n2371 240.244
R13942 gnd.n2371 gnd.n2363 240.244
R13943 gnd.n4321 gnd.n2363 240.244
R13944 gnd.n4321 gnd.n2364 240.244
R13945 gnd.n2364 gnd.n2354 240.244
R13946 gnd.n2354 gnd.n2345 240.244
R13947 gnd.n4341 gnd.n2345 240.244
R13948 gnd.n4341 gnd.n2346 240.244
R13949 gnd.n2346 gnd.n2335 240.244
R13950 gnd.n2335 gnd.n2327 240.244
R13951 gnd.n4361 gnd.n2327 240.244
R13952 gnd.n4361 gnd.n2328 240.244
R13953 gnd.n2328 gnd.n2318 240.244
R13954 gnd.n2318 gnd.n2308 240.244
R13955 gnd.n4385 gnd.n2308 240.244
R13956 gnd.n4385 gnd.n2309 240.244
R13957 gnd.n2309 gnd.n2297 240.244
R13958 gnd.n4380 gnd.n2297 240.244
R13959 gnd.n4380 gnd.n2282 240.244
R13960 gnd.n4420 gnd.n2282 240.244
R13961 gnd.n4420 gnd.n2283 240.244
R13962 gnd.n2283 gnd.n2272 240.244
R13963 gnd.n4415 gnd.n2272 240.244
R13964 gnd.n4415 gnd.n2256 240.244
R13965 gnd.n4454 gnd.n2256 240.244
R13966 gnd.n4454 gnd.n2257 240.244
R13967 gnd.n2257 gnd.n2246 240.244
R13968 gnd.n4449 gnd.n2246 240.244
R13969 gnd.n4449 gnd.n2230 240.244
R13970 gnd.n4488 gnd.n2230 240.244
R13971 gnd.n4488 gnd.n2231 240.244
R13972 gnd.n2231 gnd.n2221 240.244
R13973 gnd.n4483 gnd.n2221 240.244
R13974 gnd.n4483 gnd.n2204 240.244
R13975 gnd.n4523 gnd.n2204 240.244
R13976 gnd.n4523 gnd.n2205 240.244
R13977 gnd.n2205 gnd.n2195 240.244
R13978 gnd.n2195 gnd.n2184 240.244
R13979 gnd.n4548 gnd.n2184 240.244
R13980 gnd.n4548 gnd.n756 240.244
R13981 gnd.n769 gnd.n756 240.244
R13982 gnd.n6445 gnd.n769 240.244
R13983 gnd.n6445 gnd.n770 240.244
R13984 gnd.n6441 gnd.n770 240.244
R13985 gnd.n6441 gnd.n776 240.244
R13986 gnd.n6433 gnd.n776 240.244
R13987 gnd.n6433 gnd.n791 240.244
R13988 gnd.n6429 gnd.n791 240.244
R13989 gnd.n6429 gnd.n796 240.244
R13990 gnd.n6421 gnd.n796 240.244
R13991 gnd.n6421 gnd.n812 240.244
R13992 gnd.n6417 gnd.n812 240.244
R13993 gnd.n6417 gnd.n817 240.244
R13994 gnd.n6409 gnd.n817 240.244
R13995 gnd.n6409 gnd.n833 240.244
R13996 gnd.n5013 gnd.n862 240.244
R13997 gnd.n5014 gnd.n5013 240.244
R13998 gnd.n5024 gnd.n5014 240.244
R13999 gnd.n5024 gnd.n2062 240.244
R14000 gnd.n5030 gnd.n2062 240.244
R14001 gnd.n5030 gnd.n2055 240.244
R14002 gnd.n5042 gnd.n2055 240.244
R14003 gnd.n5042 gnd.n2051 240.244
R14004 gnd.n5048 gnd.n2051 240.244
R14005 gnd.n5048 gnd.n2043 240.244
R14006 gnd.n5059 gnd.n2043 240.244
R14007 gnd.n5059 gnd.n2039 240.244
R14008 gnd.n5065 gnd.n2039 240.244
R14009 gnd.n5065 gnd.n2030 240.244
R14010 gnd.n5078 gnd.n2030 240.244
R14011 gnd.n5078 gnd.n2025 240.244
R14012 gnd.n5148 gnd.n2025 240.244
R14013 gnd.n5148 gnd.n1628 240.244
R14014 gnd.n5083 gnd.n1628 240.244
R14015 gnd.n5083 gnd.n1620 240.244
R14016 gnd.n5084 gnd.n1620 240.244
R14017 gnd.n5087 gnd.n5084 240.244
R14018 gnd.n5088 gnd.n5087 240.244
R14019 gnd.n5089 gnd.n5088 240.244
R14020 gnd.n5089 gnd.n1595 240.244
R14021 gnd.n1595 gnd.n1589 240.244
R14022 gnd.n5092 gnd.n1589 240.244
R14023 gnd.n5092 gnd.n1582 240.244
R14024 gnd.n5093 gnd.n1582 240.244
R14025 gnd.n5093 gnd.n1567 240.244
R14026 gnd.n5096 gnd.n1567 240.244
R14027 gnd.n5096 gnd.n1561 240.244
R14028 gnd.n5097 gnd.n1561 240.244
R14029 gnd.n5097 gnd.n1550 240.244
R14030 gnd.n5100 gnd.n1550 240.244
R14031 gnd.n5100 gnd.n1543 240.244
R14032 gnd.n5101 gnd.n1543 240.244
R14033 gnd.n5101 gnd.n1531 240.244
R14034 gnd.n5104 gnd.n1531 240.244
R14035 gnd.n5104 gnd.n1523 240.244
R14036 gnd.n5105 gnd.n1523 240.244
R14037 gnd.n5105 gnd.n1511 240.244
R14038 gnd.n1511 gnd.n1504 240.244
R14039 gnd.n1504 gnd.n1493 240.244
R14040 gnd.n5369 gnd.n1493 240.244
R14041 gnd.n5369 gnd.n1488 240.244
R14042 gnd.n5389 gnd.n1488 240.244
R14043 gnd.n5389 gnd.n1482 240.244
R14044 gnd.n5374 gnd.n1482 240.244
R14045 gnd.n5374 gnd.n1474 240.244
R14046 gnd.n5375 gnd.n1474 240.244
R14047 gnd.n5376 gnd.n5375 240.244
R14048 gnd.n5376 gnd.n1453 240.244
R14049 gnd.n1453 gnd.n1443 240.244
R14050 gnd.n5466 gnd.n1443 240.244
R14051 gnd.n5466 gnd.n1438 240.244
R14052 gnd.n5483 gnd.n1438 240.244
R14053 gnd.n5483 gnd.n1432 240.244
R14054 gnd.n5471 gnd.n1432 240.244
R14055 gnd.n5471 gnd.n1424 240.244
R14056 gnd.n5472 gnd.n1424 240.244
R14057 gnd.n5472 gnd.n1403 240.244
R14058 gnd.n1403 gnd.n1393 240.244
R14059 gnd.n5542 gnd.n1393 240.244
R14060 gnd.n5542 gnd.n1388 240.244
R14061 gnd.n5552 gnd.n1388 240.244
R14062 gnd.n5552 gnd.n1376 240.244
R14063 gnd.n1376 gnd.n1368 240.244
R14064 gnd.n5585 gnd.n1368 240.244
R14065 gnd.n5586 gnd.n5585 240.244
R14066 gnd.n5586 gnd.n1347 240.244
R14067 gnd.n1362 gnd.n1347 240.244
R14068 gnd.n5612 gnd.n1362 240.244
R14069 gnd.n5612 gnd.n1363 240.244
R14070 gnd.n5592 gnd.n1363 240.244
R14071 gnd.n5592 gnd.n1327 240.244
R14072 gnd.n1327 gnd.n1322 240.244
R14073 gnd.n5594 gnd.n1322 240.244
R14074 gnd.n5594 gnd.n1315 240.244
R14075 gnd.n5597 gnd.n1315 240.244
R14076 gnd.n5597 gnd.n1226 240.244
R14077 gnd.n1226 gnd.n1218 240.244
R14078 gnd.n5819 gnd.n1218 240.244
R14079 gnd.n5819 gnd.n1214 240.244
R14080 gnd.n5825 gnd.n1214 240.244
R14081 gnd.n5825 gnd.n1207 240.244
R14082 gnd.n5836 gnd.n1207 240.244
R14083 gnd.n5836 gnd.n1203 240.244
R14084 gnd.n5842 gnd.n1203 240.244
R14085 gnd.n5842 gnd.n1195 240.244
R14086 gnd.n5853 gnd.n1195 240.244
R14087 gnd.n5853 gnd.n1191 240.244
R14088 gnd.n5859 gnd.n1191 240.244
R14089 gnd.n5859 gnd.n1184 240.244
R14090 gnd.n5871 gnd.n1184 240.244
R14091 gnd.n5871 gnd.n1180 240.244
R14092 gnd.n5877 gnd.n1180 240.244
R14093 gnd.n5877 gnd.n1172 240.244
R14094 gnd.n5890 gnd.n1172 240.244
R14095 gnd.n5890 gnd.n1167 240.244
R14096 gnd.n5914 gnd.n1167 240.244
R14097 gnd.n5005 gnd.n5004 240.244
R14098 gnd.n5004 gnd.n2069 240.244
R14099 gnd.n2074 gnd.n2073 240.244
R14100 gnd.n2077 gnd.n2076 240.244
R14101 gnd.n2087 gnd.n2086 240.244
R14102 gnd.n2090 gnd.n2089 240.244
R14103 gnd.n2102 gnd.n2101 240.244
R14104 gnd.n2113 gnd.n2104 240.244
R14105 gnd.n2116 gnd.n2115 240.244
R14106 gnd.n2128 gnd.n2127 240.244
R14107 gnd.n2139 gnd.n2130 240.244
R14108 gnd.n2142 gnd.n2141 240.244
R14109 gnd.n2159 gnd.n2158 240.244
R14110 gnd.n2163 gnd.n2161 240.244
R14111 gnd.n6384 gnd.n865 240.244
R14112 gnd.n869 gnd.n865 240.244
R14113 gnd.n870 gnd.n869 240.244
R14114 gnd.n871 gnd.n870 240.244
R14115 gnd.n5032 gnd.n871 240.244
R14116 gnd.n5032 gnd.n874 240.244
R14117 gnd.n875 gnd.n874 240.244
R14118 gnd.n876 gnd.n875 240.244
R14119 gnd.n5049 gnd.n876 240.244
R14120 gnd.n5049 gnd.n879 240.244
R14121 gnd.n880 gnd.n879 240.244
R14122 gnd.n881 gnd.n880 240.244
R14123 gnd.n5066 gnd.n881 240.244
R14124 gnd.n5066 gnd.n884 240.244
R14125 gnd.n885 gnd.n884 240.244
R14126 gnd.n886 gnd.n885 240.244
R14127 gnd.n5149 gnd.n886 240.244
R14128 gnd.n5149 gnd.n889 240.244
R14129 gnd.n890 gnd.n889 240.244
R14130 gnd.n891 gnd.n890 240.244
R14131 gnd.n1613 gnd.n891 240.244
R14132 gnd.n1613 gnd.n894 240.244
R14133 gnd.n895 gnd.n894 240.244
R14134 gnd.n896 gnd.n895 240.244
R14135 gnd.n1596 gnd.n896 240.244
R14136 gnd.n1596 gnd.n899 240.244
R14137 gnd.n900 gnd.n899 240.244
R14138 gnd.n901 gnd.n900 240.244
R14139 gnd.n1575 gnd.n901 240.244
R14140 gnd.n1575 gnd.n904 240.244
R14141 gnd.n905 gnd.n904 240.244
R14142 gnd.n906 gnd.n905 240.244
R14143 gnd.n1556 gnd.n906 240.244
R14144 gnd.n1556 gnd.n909 240.244
R14145 gnd.n910 gnd.n909 240.244
R14146 gnd.n911 gnd.n910 240.244
R14147 gnd.n1535 gnd.n911 240.244
R14148 gnd.n1535 gnd.n914 240.244
R14149 gnd.n915 gnd.n914 240.244
R14150 gnd.n916 gnd.n915 240.244
R14151 gnd.n1516 gnd.n916 240.244
R14152 gnd.n1516 gnd.n919 240.244
R14153 gnd.n920 gnd.n919 240.244
R14154 gnd.n921 gnd.n920 240.244
R14155 gnd.n1496 gnd.n921 240.244
R14156 gnd.n1496 gnd.n924 240.244
R14157 gnd.n925 gnd.n924 240.244
R14158 gnd.n926 gnd.n925 240.244
R14159 gnd.n1471 gnd.n926 240.244
R14160 gnd.n1471 gnd.n929 240.244
R14161 gnd.n930 gnd.n929 240.244
R14162 gnd.n931 gnd.n930 240.244
R14163 gnd.n5454 gnd.n931 240.244
R14164 gnd.n5454 gnd.n934 240.244
R14165 gnd.n935 gnd.n934 240.244
R14166 gnd.n936 gnd.n935 240.244
R14167 gnd.n5484 gnd.n936 240.244
R14168 gnd.n5484 gnd.n939 240.244
R14169 gnd.n940 gnd.n939 240.244
R14170 gnd.n941 gnd.n940 240.244
R14171 gnd.n1417 gnd.n941 240.244
R14172 gnd.n1417 gnd.n944 240.244
R14173 gnd.n945 gnd.n944 240.244
R14174 gnd.n946 gnd.n945 240.244
R14175 gnd.n1412 gnd.n946 240.244
R14176 gnd.n1412 gnd.n949 240.244
R14177 gnd.n950 gnd.n949 240.244
R14178 gnd.n951 gnd.n950 240.244
R14179 gnd.n1370 gnd.n951 240.244
R14180 gnd.n1370 gnd.n954 240.244
R14181 gnd.n955 gnd.n954 240.244
R14182 gnd.n956 gnd.n955 240.244
R14183 gnd.n5613 gnd.n956 240.244
R14184 gnd.n5613 gnd.n959 240.244
R14185 gnd.n960 gnd.n959 240.244
R14186 gnd.n961 gnd.n960 240.244
R14187 gnd.n5661 gnd.n961 240.244
R14188 gnd.n5661 gnd.n964 240.244
R14189 gnd.n965 gnd.n964 240.244
R14190 gnd.n966 gnd.n965 240.244
R14191 gnd.n5809 gnd.n966 240.244
R14192 gnd.n5809 gnd.n969 240.244
R14193 gnd.n970 gnd.n969 240.244
R14194 gnd.n971 gnd.n970 240.244
R14195 gnd.n5826 gnd.n971 240.244
R14196 gnd.n5826 gnd.n974 240.244
R14197 gnd.n975 gnd.n974 240.244
R14198 gnd.n976 gnd.n975 240.244
R14199 gnd.n5843 gnd.n976 240.244
R14200 gnd.n5843 gnd.n979 240.244
R14201 gnd.n980 gnd.n979 240.244
R14202 gnd.n981 gnd.n980 240.244
R14203 gnd.n5861 gnd.n981 240.244
R14204 gnd.n5861 gnd.n984 240.244
R14205 gnd.n985 gnd.n984 240.244
R14206 gnd.n986 gnd.n985 240.244
R14207 gnd.n5878 gnd.n986 240.244
R14208 gnd.n5878 gnd.n989 240.244
R14209 gnd.n990 gnd.n989 240.244
R14210 gnd.n991 gnd.n990 240.244
R14211 gnd.n995 gnd.n991 240.244
R14212 gnd.n5896 gnd.n5895 240.244
R14213 gnd.n5900 gnd.n5899 240.244
R14214 gnd.n5902 gnd.n5901 240.244
R14215 gnd.n1143 gnd.n1142 240.244
R14216 gnd.n1145 gnd.n1144 240.244
R14217 gnd.n6019 gnd.n6018 240.244
R14218 gnd.n6029 gnd.n6028 240.244
R14219 gnd.n6031 gnd.n6030 240.244
R14220 gnd.n6039 gnd.n6038 240.244
R14221 gnd.n6049 gnd.n6048 240.244
R14222 gnd.n6051 gnd.n6050 240.244
R14223 gnd.n6225 gnd.n1012 240.244
R14224 gnd.n6225 gnd.n1013 240.244
R14225 gnd.n1026 gnd.n996 240.244
R14226 gnd.n1638 gnd.n1637 240.132
R14227 gnd.n1243 gnd.n1242 240.132
R14228 gnd.n6454 gnd.n747 225.874
R14229 gnd.n6462 gnd.n747 225.874
R14230 gnd.n6463 gnd.n6462 225.874
R14231 gnd.n6464 gnd.n6463 225.874
R14232 gnd.n6464 gnd.n741 225.874
R14233 gnd.n6472 gnd.n741 225.874
R14234 gnd.n6473 gnd.n6472 225.874
R14235 gnd.n6474 gnd.n6473 225.874
R14236 gnd.n6474 gnd.n735 225.874
R14237 gnd.n6482 gnd.n735 225.874
R14238 gnd.n6483 gnd.n6482 225.874
R14239 gnd.n6484 gnd.n6483 225.874
R14240 gnd.n6484 gnd.n729 225.874
R14241 gnd.n6492 gnd.n729 225.874
R14242 gnd.n6493 gnd.n6492 225.874
R14243 gnd.n6494 gnd.n6493 225.874
R14244 gnd.n6494 gnd.n723 225.874
R14245 gnd.n6502 gnd.n723 225.874
R14246 gnd.n6503 gnd.n6502 225.874
R14247 gnd.n6504 gnd.n6503 225.874
R14248 gnd.n6504 gnd.n717 225.874
R14249 gnd.n6512 gnd.n717 225.874
R14250 gnd.n6513 gnd.n6512 225.874
R14251 gnd.n6514 gnd.n6513 225.874
R14252 gnd.n6514 gnd.n711 225.874
R14253 gnd.n6522 gnd.n711 225.874
R14254 gnd.n6523 gnd.n6522 225.874
R14255 gnd.n6524 gnd.n6523 225.874
R14256 gnd.n6524 gnd.n705 225.874
R14257 gnd.n6532 gnd.n705 225.874
R14258 gnd.n6533 gnd.n6532 225.874
R14259 gnd.n6534 gnd.n6533 225.874
R14260 gnd.n6534 gnd.n699 225.874
R14261 gnd.n6542 gnd.n699 225.874
R14262 gnd.n6543 gnd.n6542 225.874
R14263 gnd.n6544 gnd.n6543 225.874
R14264 gnd.n6544 gnd.n693 225.874
R14265 gnd.n6552 gnd.n693 225.874
R14266 gnd.n6553 gnd.n6552 225.874
R14267 gnd.n6554 gnd.n6553 225.874
R14268 gnd.n6554 gnd.n687 225.874
R14269 gnd.n6562 gnd.n687 225.874
R14270 gnd.n6563 gnd.n6562 225.874
R14271 gnd.n6564 gnd.n6563 225.874
R14272 gnd.n6564 gnd.n681 225.874
R14273 gnd.n6572 gnd.n681 225.874
R14274 gnd.n6573 gnd.n6572 225.874
R14275 gnd.n6574 gnd.n6573 225.874
R14276 gnd.n6574 gnd.n675 225.874
R14277 gnd.n6582 gnd.n675 225.874
R14278 gnd.n6583 gnd.n6582 225.874
R14279 gnd.n6584 gnd.n6583 225.874
R14280 gnd.n6584 gnd.n669 225.874
R14281 gnd.n6592 gnd.n669 225.874
R14282 gnd.n6593 gnd.n6592 225.874
R14283 gnd.n6594 gnd.n6593 225.874
R14284 gnd.n6594 gnd.n663 225.874
R14285 gnd.n6602 gnd.n663 225.874
R14286 gnd.n6603 gnd.n6602 225.874
R14287 gnd.n6604 gnd.n6603 225.874
R14288 gnd.n6604 gnd.n657 225.874
R14289 gnd.n6612 gnd.n657 225.874
R14290 gnd.n6613 gnd.n6612 225.874
R14291 gnd.n6614 gnd.n6613 225.874
R14292 gnd.n6614 gnd.n651 225.874
R14293 gnd.n6622 gnd.n651 225.874
R14294 gnd.n6623 gnd.n6622 225.874
R14295 gnd.n6624 gnd.n6623 225.874
R14296 gnd.n6624 gnd.n645 225.874
R14297 gnd.n6632 gnd.n645 225.874
R14298 gnd.n6633 gnd.n6632 225.874
R14299 gnd.n6634 gnd.n6633 225.874
R14300 gnd.n6634 gnd.n639 225.874
R14301 gnd.n6642 gnd.n639 225.874
R14302 gnd.n6643 gnd.n6642 225.874
R14303 gnd.n6644 gnd.n6643 225.874
R14304 gnd.n6644 gnd.n633 225.874
R14305 gnd.n6652 gnd.n633 225.874
R14306 gnd.n6653 gnd.n6652 225.874
R14307 gnd.n6654 gnd.n6653 225.874
R14308 gnd.n6654 gnd.n627 225.874
R14309 gnd.n6662 gnd.n627 225.874
R14310 gnd.n6663 gnd.n6662 225.874
R14311 gnd.n6664 gnd.n6663 225.874
R14312 gnd.n6664 gnd.n621 225.874
R14313 gnd.n6672 gnd.n621 225.874
R14314 gnd.n6673 gnd.n6672 225.874
R14315 gnd.n6674 gnd.n6673 225.874
R14316 gnd.n6674 gnd.n615 225.874
R14317 gnd.n6682 gnd.n615 225.874
R14318 gnd.n6683 gnd.n6682 225.874
R14319 gnd.n6684 gnd.n6683 225.874
R14320 gnd.n6684 gnd.n609 225.874
R14321 gnd.n6692 gnd.n609 225.874
R14322 gnd.n6693 gnd.n6692 225.874
R14323 gnd.n6694 gnd.n6693 225.874
R14324 gnd.n6694 gnd.n603 225.874
R14325 gnd.n6702 gnd.n603 225.874
R14326 gnd.n6703 gnd.n6702 225.874
R14327 gnd.n6704 gnd.n6703 225.874
R14328 gnd.n6704 gnd.n597 225.874
R14329 gnd.n6712 gnd.n597 225.874
R14330 gnd.n6713 gnd.n6712 225.874
R14331 gnd.n6714 gnd.n6713 225.874
R14332 gnd.n6714 gnd.n591 225.874
R14333 gnd.n6722 gnd.n591 225.874
R14334 gnd.n6723 gnd.n6722 225.874
R14335 gnd.n6724 gnd.n6723 225.874
R14336 gnd.n6724 gnd.n585 225.874
R14337 gnd.n6732 gnd.n585 225.874
R14338 gnd.n6733 gnd.n6732 225.874
R14339 gnd.n6734 gnd.n6733 225.874
R14340 gnd.n6734 gnd.n579 225.874
R14341 gnd.n6742 gnd.n579 225.874
R14342 gnd.n6743 gnd.n6742 225.874
R14343 gnd.n6744 gnd.n6743 225.874
R14344 gnd.n6744 gnd.n573 225.874
R14345 gnd.n6752 gnd.n573 225.874
R14346 gnd.n6753 gnd.n6752 225.874
R14347 gnd.n6754 gnd.n6753 225.874
R14348 gnd.n6754 gnd.n567 225.874
R14349 gnd.n6762 gnd.n567 225.874
R14350 gnd.n6763 gnd.n6762 225.874
R14351 gnd.n6764 gnd.n6763 225.874
R14352 gnd.n6764 gnd.n561 225.874
R14353 gnd.n6772 gnd.n561 225.874
R14354 gnd.n6773 gnd.n6772 225.874
R14355 gnd.n6774 gnd.n6773 225.874
R14356 gnd.n6774 gnd.n555 225.874
R14357 gnd.n6782 gnd.n555 225.874
R14358 gnd.n6783 gnd.n6782 225.874
R14359 gnd.n6784 gnd.n6783 225.874
R14360 gnd.n6784 gnd.n549 225.874
R14361 gnd.n6792 gnd.n549 225.874
R14362 gnd.n6793 gnd.n6792 225.874
R14363 gnd.n6794 gnd.n6793 225.874
R14364 gnd.n6794 gnd.n543 225.874
R14365 gnd.n6803 gnd.n543 225.874
R14366 gnd.n6804 gnd.n6803 225.874
R14367 gnd.n6805 gnd.n6804 225.874
R14368 gnd.n6805 gnd.n538 225.874
R14369 gnd.n2999 gnd.t33 224.174
R14370 gnd.n2477 gnd.t136 224.174
R14371 gnd.n1102 gnd.n1043 199.319
R14372 gnd.n1102 gnd.n1044 199.319
R14373 gnd.n1841 gnd.n1752 199.319
R14374 gnd.n1849 gnd.n1752 199.319
R14375 gnd.n1639 gnd.n1636 186.49
R14376 gnd.n1244 gnd.n1241 186.49
R14377 gnd.n3774 gnd.n3773 185
R14378 gnd.n3772 gnd.n3771 185
R14379 gnd.n3751 gnd.n3750 185
R14380 gnd.n3766 gnd.n3765 185
R14381 gnd.n3764 gnd.n3763 185
R14382 gnd.n3755 gnd.n3754 185
R14383 gnd.n3758 gnd.n3757 185
R14384 gnd.n3742 gnd.n3741 185
R14385 gnd.n3740 gnd.n3739 185
R14386 gnd.n3719 gnd.n3718 185
R14387 gnd.n3734 gnd.n3733 185
R14388 gnd.n3732 gnd.n3731 185
R14389 gnd.n3723 gnd.n3722 185
R14390 gnd.n3726 gnd.n3725 185
R14391 gnd.n3710 gnd.n3709 185
R14392 gnd.n3708 gnd.n3707 185
R14393 gnd.n3687 gnd.n3686 185
R14394 gnd.n3702 gnd.n3701 185
R14395 gnd.n3700 gnd.n3699 185
R14396 gnd.n3691 gnd.n3690 185
R14397 gnd.n3694 gnd.n3693 185
R14398 gnd.n3679 gnd.n3678 185
R14399 gnd.n3677 gnd.n3676 185
R14400 gnd.n3656 gnd.n3655 185
R14401 gnd.n3671 gnd.n3670 185
R14402 gnd.n3669 gnd.n3668 185
R14403 gnd.n3660 gnd.n3659 185
R14404 gnd.n3663 gnd.n3662 185
R14405 gnd.n3647 gnd.n3646 185
R14406 gnd.n3645 gnd.n3644 185
R14407 gnd.n3624 gnd.n3623 185
R14408 gnd.n3639 gnd.n3638 185
R14409 gnd.n3637 gnd.n3636 185
R14410 gnd.n3628 gnd.n3627 185
R14411 gnd.n3631 gnd.n3630 185
R14412 gnd.n3615 gnd.n3614 185
R14413 gnd.n3613 gnd.n3612 185
R14414 gnd.n3592 gnd.n3591 185
R14415 gnd.n3607 gnd.n3606 185
R14416 gnd.n3605 gnd.n3604 185
R14417 gnd.n3596 gnd.n3595 185
R14418 gnd.n3599 gnd.n3598 185
R14419 gnd.n3583 gnd.n3582 185
R14420 gnd.n3581 gnd.n3580 185
R14421 gnd.n3560 gnd.n3559 185
R14422 gnd.n3575 gnd.n3574 185
R14423 gnd.n3573 gnd.n3572 185
R14424 gnd.n3564 gnd.n3563 185
R14425 gnd.n3567 gnd.n3566 185
R14426 gnd.n3552 gnd.n3551 185
R14427 gnd.n3550 gnd.n3549 185
R14428 gnd.n3529 gnd.n3528 185
R14429 gnd.n3544 gnd.n3543 185
R14430 gnd.n3542 gnd.n3541 185
R14431 gnd.n3533 gnd.n3532 185
R14432 gnd.n3536 gnd.n3535 185
R14433 gnd.n3000 gnd.t32 178.987
R14434 gnd.n2478 gnd.t137 178.987
R14435 gnd.n1 gnd.t205 170.774
R14436 gnd.n9 gnd.t162 170.103
R14437 gnd.n8 gnd.t168 170.103
R14438 gnd.n7 gnd.t201 170.103
R14439 gnd.n6 gnd.t148 170.103
R14440 gnd.n5 gnd.t211 170.103
R14441 gnd.n4 gnd.t199 170.103
R14442 gnd.n3 gnd.t16 170.103
R14443 gnd.n2 gnd.t203 170.103
R14444 gnd.n1 gnd.t22 170.103
R14445 gnd.n5800 gnd.n1254 163.367
R14446 gnd.n5796 gnd.n5795 163.367
R14447 gnd.n5793 gnd.n1257 163.367
R14448 gnd.n5789 gnd.n5788 163.367
R14449 gnd.n5786 gnd.n1260 163.367
R14450 gnd.n5782 gnd.n5781 163.367
R14451 gnd.n5779 gnd.n1263 163.367
R14452 gnd.n5775 gnd.n5774 163.367
R14453 gnd.n5772 gnd.n1266 163.367
R14454 gnd.n5768 gnd.n5767 163.367
R14455 gnd.n5765 gnd.n1269 163.367
R14456 gnd.n5761 gnd.n5760 163.367
R14457 gnd.n5758 gnd.n1272 163.367
R14458 gnd.n5754 gnd.n5753 163.367
R14459 gnd.n5751 gnd.n1275 163.367
R14460 gnd.n5747 gnd.n5746 163.367
R14461 gnd.n5743 gnd.n5742 163.367
R14462 gnd.n5740 gnd.n1281 163.367
R14463 gnd.n5735 gnd.n5734 163.367
R14464 gnd.n5732 gnd.n1286 163.367
R14465 gnd.n5728 gnd.n5727 163.367
R14466 gnd.n5725 gnd.n1289 163.367
R14467 gnd.n5721 gnd.n5720 163.367
R14468 gnd.n5718 gnd.n1292 163.367
R14469 gnd.n5714 gnd.n5713 163.367
R14470 gnd.n5711 gnd.n1295 163.367
R14471 gnd.n5707 gnd.n5706 163.367
R14472 gnd.n5704 gnd.n1298 163.367
R14473 gnd.n5700 gnd.n5699 163.367
R14474 gnd.n5697 gnd.n1301 163.367
R14475 gnd.n5693 gnd.n5692 163.367
R14476 gnd.n5690 gnd.n1304 163.367
R14477 gnd.n2019 gnd.n1629 163.367
R14478 gnd.n2019 gnd.n1619 163.367
R14479 gnd.n1619 gnd.n1611 163.367
R14480 gnd.n5187 gnd.n1611 163.367
R14481 gnd.n5187 gnd.n1609 163.367
R14482 gnd.n5191 gnd.n1609 163.367
R14483 gnd.n5191 gnd.n1601 163.367
R14484 gnd.n5200 gnd.n1601 163.367
R14485 gnd.n5200 gnd.n1597 163.367
R14486 gnd.n5211 gnd.n1597 163.367
R14487 gnd.n5211 gnd.n1599 163.367
R14488 gnd.n1599 gnd.n1590 163.367
R14489 gnd.n5206 gnd.n1590 163.367
R14490 gnd.n5206 gnd.n1581 163.367
R14491 gnd.n5203 gnd.n1581 163.367
R14492 gnd.n5203 gnd.n1574 163.367
R14493 gnd.n5236 gnd.n1574 163.367
R14494 gnd.n5236 gnd.n1568 163.367
R14495 gnd.n5240 gnd.n1568 163.367
R14496 gnd.n5240 gnd.n1560 163.367
R14497 gnd.n5259 gnd.n1560 163.367
R14498 gnd.n5259 gnd.n1558 163.367
R14499 gnd.n5267 gnd.n1558 163.367
R14500 gnd.n5267 gnd.n1551 163.367
R14501 gnd.n5263 gnd.n1551 163.367
R14502 gnd.n5263 gnd.n1542 163.367
R14503 gnd.n1542 gnd.n1534 163.367
R14504 gnd.n5293 gnd.n1534 163.367
R14505 gnd.n5293 gnd.n1532 163.367
R14506 gnd.n5298 gnd.n1532 163.367
R14507 gnd.n5298 gnd.n1522 163.367
R14508 gnd.n1522 gnd.n1515 163.367
R14509 gnd.n5319 gnd.n1515 163.367
R14510 gnd.n5319 gnd.n1512 163.367
R14511 gnd.n5345 gnd.n1512 163.367
R14512 gnd.n5345 gnd.n1513 163.367
R14513 gnd.n1513 gnd.n1505 163.367
R14514 gnd.n5340 gnd.n1505 163.367
R14515 gnd.n5340 gnd.n5337 163.367
R14516 gnd.n5337 gnd.n5336 163.367
R14517 gnd.n5336 gnd.n5325 163.367
R14518 gnd.n5325 gnd.n1487 163.367
R14519 gnd.n5331 gnd.n1487 163.367
R14520 gnd.n5331 gnd.n1483 163.367
R14521 gnd.n5328 gnd.n1483 163.367
R14522 gnd.n5328 gnd.n1473 163.367
R14523 gnd.n1473 gnd.n1464 163.367
R14524 gnd.n5416 gnd.n1464 163.367
R14525 gnd.n5416 gnd.n1461 163.367
R14526 gnd.n5441 gnd.n1461 163.367
R14527 gnd.n5441 gnd.n1462 163.367
R14528 gnd.n1462 gnd.n1454 163.367
R14529 gnd.n5436 gnd.n1454 163.367
R14530 gnd.n5436 gnd.n5434 163.367
R14531 gnd.n5434 gnd.n5433 163.367
R14532 gnd.n5433 gnd.n5422 163.367
R14533 gnd.n5422 gnd.n1437 163.367
R14534 gnd.n5428 gnd.n1437 163.367
R14535 gnd.n5428 gnd.n1433 163.367
R14536 gnd.n5425 gnd.n1433 163.367
R14537 gnd.n5425 gnd.n1423 163.367
R14538 gnd.n1423 gnd.n1416 163.367
R14539 gnd.n5509 gnd.n1416 163.367
R14540 gnd.n5510 gnd.n5509 163.367
R14541 gnd.n5510 gnd.n1404 163.367
R14542 gnd.n5516 gnd.n1404 163.367
R14543 gnd.n5517 gnd.n5516 163.367
R14544 gnd.n5517 gnd.n1414 163.367
R14545 gnd.n5521 gnd.n1414 163.367
R14546 gnd.n5521 gnd.n1386 163.367
R14547 gnd.n5555 gnd.n1386 163.367
R14548 gnd.n5555 gnd.n1377 163.367
R14549 gnd.n5559 gnd.n1377 163.367
R14550 gnd.n5560 gnd.n5559 163.367
R14551 gnd.n5560 gnd.n1384 163.367
R14552 gnd.n5565 gnd.n1384 163.367
R14553 gnd.n5565 gnd.n1346 163.367
R14554 gnd.n1346 gnd.n1340 163.367
R14555 gnd.n5628 gnd.n1340 163.367
R14556 gnd.n5628 gnd.n1338 163.367
R14557 gnd.n5632 gnd.n1338 163.367
R14558 gnd.n5632 gnd.n1331 163.367
R14559 gnd.n5641 gnd.n1331 163.367
R14560 gnd.n5641 gnd.n1328 163.367
R14561 gnd.n5653 gnd.n1328 163.367
R14562 gnd.n5653 gnd.n1329 163.367
R14563 gnd.n1329 gnd.n1323 163.367
R14564 gnd.n5648 gnd.n1323 163.367
R14565 gnd.n5648 gnd.n1314 163.367
R14566 gnd.n5645 gnd.n1314 163.367
R14567 gnd.n5645 gnd.n1308 163.367
R14568 gnd.n5679 gnd.n1308 163.367
R14569 gnd.n5679 gnd.n1227 163.367
R14570 gnd.n5684 gnd.n1227 163.367
R14571 gnd.n5685 gnd.n5684 163.367
R14572 gnd.n5153 gnd.n1653 163.367
R14573 gnd.n1692 gnd.n1653 163.367
R14574 gnd.n1696 gnd.n1695 163.367
R14575 gnd.n1700 gnd.n1699 163.367
R14576 gnd.n1704 gnd.n1703 163.367
R14577 gnd.n1708 gnd.n1707 163.367
R14578 gnd.n1712 gnd.n1711 163.367
R14579 gnd.n1716 gnd.n1715 163.367
R14580 gnd.n1720 gnd.n1719 163.367
R14581 gnd.n1724 gnd.n1723 163.367
R14582 gnd.n1728 gnd.n1727 163.367
R14583 gnd.n1732 gnd.n1731 163.367
R14584 gnd.n1736 gnd.n1735 163.367
R14585 gnd.n1740 gnd.n1739 163.367
R14586 gnd.n1744 gnd.n1743 163.367
R14587 gnd.n1748 gnd.n1747 163.367
R14588 gnd.n1956 gnd.n1955 163.367
R14589 gnd.n1960 gnd.n1959 163.367
R14590 gnd.n1965 gnd.n1964 163.367
R14591 gnd.n1969 gnd.n1968 163.367
R14592 gnd.n1973 gnd.n1972 163.367
R14593 gnd.n1977 gnd.n1976 163.367
R14594 gnd.n1981 gnd.n1980 163.367
R14595 gnd.n1985 gnd.n1984 163.367
R14596 gnd.n1989 gnd.n1988 163.367
R14597 gnd.n1993 gnd.n1992 163.367
R14598 gnd.n1997 gnd.n1996 163.367
R14599 gnd.n2001 gnd.n2000 163.367
R14600 gnd.n2005 gnd.n2004 163.367
R14601 gnd.n2009 gnd.n2008 163.367
R14602 gnd.n2013 gnd.n2012 163.367
R14603 gnd.n2015 gnd.n1686 163.367
R14604 gnd.n5158 gnd.n1617 163.367
R14605 gnd.n5181 gnd.n1617 163.367
R14606 gnd.n5181 gnd.n1615 163.367
R14607 gnd.n5185 gnd.n1615 163.367
R14608 gnd.n5185 gnd.n1607 163.367
R14609 gnd.n5194 gnd.n1607 163.367
R14610 gnd.n5194 gnd.n1605 163.367
R14611 gnd.n5198 gnd.n1605 163.367
R14612 gnd.n5198 gnd.n1594 163.367
R14613 gnd.n5213 gnd.n1594 163.367
R14614 gnd.n5213 gnd.n1592 163.367
R14615 gnd.n5217 gnd.n1592 163.367
R14616 gnd.n5217 gnd.n1579 163.367
R14617 gnd.n5229 gnd.n1579 163.367
R14618 gnd.n5229 gnd.n1577 163.367
R14619 gnd.n5233 gnd.n1577 163.367
R14620 gnd.n5233 gnd.n1570 163.367
R14621 gnd.n5247 gnd.n1570 163.367
R14622 gnd.n5247 gnd.n1571 163.367
R14623 gnd.n5243 gnd.n1571 163.367
R14624 gnd.n5243 gnd.n1555 163.367
R14625 gnd.n5270 gnd.n1555 163.367
R14626 gnd.n5270 gnd.n1553 163.367
R14627 gnd.n5274 gnd.n1553 163.367
R14628 gnd.n5274 gnd.n1540 163.367
R14629 gnd.n5286 gnd.n1540 163.367
R14630 gnd.n5286 gnd.n1537 163.367
R14631 gnd.n5291 gnd.n1537 163.367
R14632 gnd.n5291 gnd.n1538 163.367
R14633 gnd.n1538 gnd.n1520 163.367
R14634 gnd.n5313 gnd.n1520 163.367
R14635 gnd.n5313 gnd.n1518 163.367
R14636 gnd.n5317 gnd.n1518 163.367
R14637 gnd.n5317 gnd.n1509 163.367
R14638 gnd.n5347 gnd.n1509 163.367
R14639 gnd.n5347 gnd.n1506 163.367
R14640 gnd.n5356 gnd.n1506 163.367
R14641 gnd.n5356 gnd.n1507 163.367
R14642 gnd.n5352 gnd.n1507 163.367
R14643 gnd.n5352 gnd.n5351 163.367
R14644 gnd.n5351 gnd.n1486 163.367
R14645 gnd.n5392 gnd.n1486 163.367
R14646 gnd.n5392 gnd.n1484 163.367
R14647 gnd.n5396 gnd.n1484 163.367
R14648 gnd.n5396 gnd.n1470 163.367
R14649 gnd.n5410 gnd.n1470 163.367
R14650 gnd.n5410 gnd.n1468 163.367
R14651 gnd.n5414 gnd.n1468 163.367
R14652 gnd.n5414 gnd.n1459 163.367
R14653 gnd.n5443 gnd.n1459 163.367
R14654 gnd.n5443 gnd.n1456 163.367
R14655 gnd.n5452 gnd.n1456 163.367
R14656 gnd.n5452 gnd.n1457 163.367
R14657 gnd.n5448 gnd.n1457 163.367
R14658 gnd.n5448 gnd.n5447 163.367
R14659 gnd.n5447 gnd.n1436 163.367
R14660 gnd.n5487 gnd.n1436 163.367
R14661 gnd.n5487 gnd.n1434 163.367
R14662 gnd.n5491 gnd.n1434 163.367
R14663 gnd.n5491 gnd.n1421 163.367
R14664 gnd.n5503 gnd.n1421 163.367
R14665 gnd.n5503 gnd.n1419 163.367
R14666 gnd.n5507 gnd.n1419 163.367
R14667 gnd.n5507 gnd.n1405 163.367
R14668 gnd.n5529 gnd.n1405 163.367
R14669 gnd.n5529 gnd.n1406 163.367
R14670 gnd.n5525 gnd.n1406 163.367
R14671 gnd.n5525 gnd.n5524 163.367
R14672 gnd.n5524 gnd.n5523 163.367
R14673 gnd.n5523 gnd.n1409 163.367
R14674 gnd.n1409 gnd.n1380 163.367
R14675 gnd.n5573 gnd.n1380 163.367
R14676 gnd.n5573 gnd.n1381 163.367
R14677 gnd.n5569 gnd.n1381 163.367
R14678 gnd.n5569 gnd.n5568 163.367
R14679 gnd.n5568 gnd.n1344 163.367
R14680 gnd.n5622 gnd.n1344 163.367
R14681 gnd.n5622 gnd.n1342 163.367
R14682 gnd.n5626 gnd.n1342 163.367
R14683 gnd.n5626 gnd.n1337 163.367
R14684 gnd.n5635 gnd.n1337 163.367
R14685 gnd.n5635 gnd.n1335 163.367
R14686 gnd.n5639 gnd.n1335 163.367
R14687 gnd.n5639 gnd.n1326 163.367
R14688 gnd.n5655 gnd.n1326 163.367
R14689 gnd.n5655 gnd.n1324 163.367
R14690 gnd.n5659 gnd.n1324 163.367
R14691 gnd.n5659 gnd.n1312 163.367
R14692 gnd.n5672 gnd.n1312 163.367
R14693 gnd.n5672 gnd.n1310 163.367
R14694 gnd.n5676 gnd.n1310 163.367
R14695 gnd.n5676 gnd.n1229 163.367
R14696 gnd.n5807 gnd.n1229 163.367
R14697 gnd.n5807 gnd.n1230 163.367
R14698 gnd.n5803 gnd.n1230 163.367
R14699 gnd.n1250 gnd.n1249 156.462
R14700 gnd.n3714 gnd.n3682 153.042
R14701 gnd.n3778 gnd.n3777 152.079
R14702 gnd.n3746 gnd.n3745 152.079
R14703 gnd.n3714 gnd.n3713 152.079
R14704 gnd.n1644 gnd.n1643 152
R14705 gnd.n1645 gnd.n1634 152
R14706 gnd.n1647 gnd.n1646 152
R14707 gnd.n1649 gnd.n1632 152
R14708 gnd.n1651 gnd.n1650 152
R14709 gnd.n1248 gnd.n1232 152
R14710 gnd.n1240 gnd.n1233 152
R14711 gnd.n1239 gnd.n1238 152
R14712 gnd.n1237 gnd.n1234 152
R14713 gnd.n1235 gnd.t42 150.546
R14714 gnd.t213 gnd.n3756 147.661
R14715 gnd.t25 gnd.n3724 147.661
R14716 gnd.t150 gnd.n3692 147.661
R14717 gnd.t174 gnd.n3661 147.661
R14718 gnd.t181 gnd.n3629 147.661
R14719 gnd.t157 gnd.n3597 147.661
R14720 gnd.t176 gnd.n3565 147.661
R14721 gnd.t207 gnd.n3534 147.661
R14722 gnd.n5745 gnd.n5744 143.351
R14723 gnd.n1953 gnd.n1669 143.351
R14724 gnd.n1953 gnd.n1670 143.351
R14725 gnd.n6162 gnd.n1101 138.177
R14726 gnd.n1954 gnd.n1952 138.177
R14727 gnd.n1641 gnd.t103 130.484
R14728 gnd.n1650 gnd.t128 126.766
R14729 gnd.n1648 gnd.t49 126.766
R14730 gnd.n1634 gnd.t113 126.766
R14731 gnd.n1642 gnd.t81 126.766
R14732 gnd.n1236 gnd.t27 126.766
R14733 gnd.n1238 gnd.t141 126.766
R14734 gnd.n1247 gnd.t90 126.766
R14735 gnd.n1249 gnd.t67 126.766
R14736 gnd.n3773 gnd.n3772 104.615
R14737 gnd.n3772 gnd.n3750 104.615
R14738 gnd.n3765 gnd.n3750 104.615
R14739 gnd.n3765 gnd.n3764 104.615
R14740 gnd.n3764 gnd.n3754 104.615
R14741 gnd.n3757 gnd.n3754 104.615
R14742 gnd.n3741 gnd.n3740 104.615
R14743 gnd.n3740 gnd.n3718 104.615
R14744 gnd.n3733 gnd.n3718 104.615
R14745 gnd.n3733 gnd.n3732 104.615
R14746 gnd.n3732 gnd.n3722 104.615
R14747 gnd.n3725 gnd.n3722 104.615
R14748 gnd.n3709 gnd.n3708 104.615
R14749 gnd.n3708 gnd.n3686 104.615
R14750 gnd.n3701 gnd.n3686 104.615
R14751 gnd.n3701 gnd.n3700 104.615
R14752 gnd.n3700 gnd.n3690 104.615
R14753 gnd.n3693 gnd.n3690 104.615
R14754 gnd.n3678 gnd.n3677 104.615
R14755 gnd.n3677 gnd.n3655 104.615
R14756 gnd.n3670 gnd.n3655 104.615
R14757 gnd.n3670 gnd.n3669 104.615
R14758 gnd.n3669 gnd.n3659 104.615
R14759 gnd.n3662 gnd.n3659 104.615
R14760 gnd.n3646 gnd.n3645 104.615
R14761 gnd.n3645 gnd.n3623 104.615
R14762 gnd.n3638 gnd.n3623 104.615
R14763 gnd.n3638 gnd.n3637 104.615
R14764 gnd.n3637 gnd.n3627 104.615
R14765 gnd.n3630 gnd.n3627 104.615
R14766 gnd.n3614 gnd.n3613 104.615
R14767 gnd.n3613 gnd.n3591 104.615
R14768 gnd.n3606 gnd.n3591 104.615
R14769 gnd.n3606 gnd.n3605 104.615
R14770 gnd.n3605 gnd.n3595 104.615
R14771 gnd.n3598 gnd.n3595 104.615
R14772 gnd.n3582 gnd.n3581 104.615
R14773 gnd.n3581 gnd.n3559 104.615
R14774 gnd.n3574 gnd.n3559 104.615
R14775 gnd.n3574 gnd.n3573 104.615
R14776 gnd.n3573 gnd.n3563 104.615
R14777 gnd.n3566 gnd.n3563 104.615
R14778 gnd.n3551 gnd.n3550 104.615
R14779 gnd.n3550 gnd.n3528 104.615
R14780 gnd.n3543 gnd.n3528 104.615
R14781 gnd.n3543 gnd.n3542 104.615
R14782 gnd.n3542 gnd.n3532 104.615
R14783 gnd.n3535 gnd.n3532 104.615
R14784 gnd.n2925 gnd.t59 100.632
R14785 gnd.n2451 gnd.t108 100.632
R14786 gnd.n7498 gnd.n7496 99.6594
R14787 gnd.n7504 gnd.n7489 99.6594
R14788 gnd.n7508 gnd.n7506 99.6594
R14789 gnd.n7514 gnd.n7485 99.6594
R14790 gnd.n7518 gnd.n7516 99.6594
R14791 gnd.n7524 gnd.n7481 99.6594
R14792 gnd.n7529 gnd.n7526 99.6594
R14793 gnd.n7527 gnd.n7477 99.6594
R14794 gnd.n7539 gnd.n7537 99.6594
R14795 gnd.n7545 gnd.n7471 99.6594
R14796 gnd.n7549 gnd.n7547 99.6594
R14797 gnd.n7555 gnd.n7467 99.6594
R14798 gnd.n7559 gnd.n7557 99.6594
R14799 gnd.n7565 gnd.n7463 99.6594
R14800 gnd.n7569 gnd.n7567 99.6594
R14801 gnd.n7575 gnd.n7459 99.6594
R14802 gnd.n7579 gnd.n7577 99.6594
R14803 gnd.n7585 gnd.n7455 99.6594
R14804 gnd.n7589 gnd.n7587 99.6594
R14805 gnd.n7595 gnd.n7449 99.6594
R14806 gnd.n7599 gnd.n7597 99.6594
R14807 gnd.n7605 gnd.n7445 99.6594
R14808 gnd.n7609 gnd.n7607 99.6594
R14809 gnd.n7615 gnd.n7441 99.6594
R14810 gnd.n7619 gnd.n7617 99.6594
R14811 gnd.n7625 gnd.n7437 99.6594
R14812 gnd.n7629 gnd.n7627 99.6594
R14813 gnd.n7635 gnd.n7433 99.6594
R14814 gnd.n7638 gnd.n7637 99.6594
R14815 gnd.n6214 gnd.n6213 99.6594
R14816 gnd.n6208 gnd.n1032 99.6594
R14817 gnd.n6205 gnd.n1033 99.6594
R14818 gnd.n6201 gnd.n1034 99.6594
R14819 gnd.n6197 gnd.n1035 99.6594
R14820 gnd.n6193 gnd.n1036 99.6594
R14821 gnd.n6189 gnd.n1037 99.6594
R14822 gnd.n6185 gnd.n1038 99.6594
R14823 gnd.n6181 gnd.n1039 99.6594
R14824 gnd.n6176 gnd.n1040 99.6594
R14825 gnd.n6172 gnd.n1041 99.6594
R14826 gnd.n6168 gnd.n1042 99.6594
R14827 gnd.n6164 gnd.n1043 99.6594
R14828 gnd.n6159 gnd.n1045 99.6594
R14829 gnd.n6155 gnd.n1046 99.6594
R14830 gnd.n6151 gnd.n1047 99.6594
R14831 gnd.n6147 gnd.n1048 99.6594
R14832 gnd.n6143 gnd.n1049 99.6594
R14833 gnd.n6139 gnd.n1050 99.6594
R14834 gnd.n6135 gnd.n1051 99.6594
R14835 gnd.n6131 gnd.n1052 99.6594
R14836 gnd.n6127 gnd.n1053 99.6594
R14837 gnd.n6123 gnd.n1054 99.6594
R14838 gnd.n6119 gnd.n1055 99.6594
R14839 gnd.n6115 gnd.n1056 99.6594
R14840 gnd.n6111 gnd.n1057 99.6594
R14841 gnd.n6107 gnd.n1058 99.6594
R14842 gnd.n6103 gnd.n1059 99.6594
R14843 gnd.n7424 gnd.n7293 99.6594
R14844 gnd.n7422 gnd.n7421 99.6594
R14845 gnd.n7417 gnd.n7300 99.6594
R14846 gnd.n7415 gnd.n7414 99.6594
R14847 gnd.n7410 gnd.n7307 99.6594
R14848 gnd.n7408 gnd.n7407 99.6594
R14849 gnd.n7403 gnd.n7314 99.6594
R14850 gnd.n7401 gnd.n7400 99.6594
R14851 gnd.n7319 gnd.n7318 99.6594
R14852 gnd.n6012 gnd.n1060 99.6594
R14853 gnd.n6015 gnd.n1061 99.6594
R14854 gnd.n6023 gnd.n1062 99.6594
R14855 gnd.n6025 gnd.n1063 99.6594
R14856 gnd.n6035 gnd.n1064 99.6594
R14857 gnd.n6043 gnd.n1065 99.6594
R14858 gnd.n6045 gnd.n1066 99.6594
R14859 gnd.n6055 gnd.n1068 99.6594
R14860 gnd.n6216 gnd.n1021 99.6594
R14861 gnd.n4657 gnd.n751 99.6594
R14862 gnd.n4661 gnd.n4660 99.6594
R14863 gnd.n4668 gnd.n4667 99.6594
R14864 gnd.n4671 gnd.n4670 99.6594
R14865 gnd.n4678 gnd.n4677 99.6594
R14866 gnd.n4681 gnd.n4680 99.6594
R14867 gnd.n4688 gnd.n4687 99.6594
R14868 gnd.n4691 gnd.n4690 99.6594
R14869 gnd.n4698 gnd.n4697 99.6594
R14870 gnd.n4701 gnd.n4700 99.6594
R14871 gnd.n4708 gnd.n4707 99.6594
R14872 gnd.n4711 gnd.n4710 99.6594
R14873 gnd.n4718 gnd.n4717 99.6594
R14874 gnd.n4721 gnd.n4720 99.6594
R14875 gnd.n4728 gnd.n4727 99.6594
R14876 gnd.n4731 gnd.n4730 99.6594
R14877 gnd.n4738 gnd.n4737 99.6594
R14878 gnd.n4741 gnd.n4740 99.6594
R14879 gnd.n4748 gnd.n4747 99.6594
R14880 gnd.n4751 gnd.n4750 99.6594
R14881 gnd.n4758 gnd.n4757 99.6594
R14882 gnd.n4761 gnd.n4760 99.6594
R14883 gnd.n4768 gnd.n4767 99.6594
R14884 gnd.n4771 gnd.n4770 99.6594
R14885 gnd.n4778 gnd.n4777 99.6594
R14886 gnd.n4781 gnd.n4780 99.6594
R14887 gnd.n4788 gnd.n4787 99.6594
R14888 gnd.n4791 gnd.n4790 99.6594
R14889 gnd.n4798 gnd.n4797 99.6594
R14890 gnd.n4801 gnd.n4800 99.6594
R14891 gnd.n4808 gnd.n4807 99.6594
R14892 gnd.n4811 gnd.n4810 99.6594
R14893 gnd.n4818 gnd.n4817 99.6594
R14894 gnd.n4821 gnd.n4820 99.6594
R14895 gnd.n4828 gnd.n4827 99.6594
R14896 gnd.n4831 gnd.n4830 99.6594
R14897 gnd.n4838 gnd.n4837 99.6594
R14898 gnd.n4841 gnd.n4840 99.6594
R14899 gnd.n4848 gnd.n4847 99.6594
R14900 gnd.n4851 gnd.n4850 99.6594
R14901 gnd.n4859 gnd.n4858 99.6594
R14902 gnd.n4862 gnd.n4861 99.6594
R14903 gnd.n1783 gnd.n1777 99.6594
R14904 gnd.n1792 gnd.n1791 99.6594
R14905 gnd.n1793 gnd.n1773 99.6594
R14906 gnd.n1802 gnd.n1801 99.6594
R14907 gnd.n1803 gnd.n1769 99.6594
R14908 gnd.n1812 gnd.n1811 99.6594
R14909 gnd.n1813 gnd.n1765 99.6594
R14910 gnd.n1822 gnd.n1821 99.6594
R14911 gnd.n1828 gnd.n1759 99.6594
R14912 gnd.n1832 gnd.n1830 99.6594
R14913 gnd.n1838 gnd.n1755 99.6594
R14914 gnd.n1843 gnd.n1840 99.6594
R14915 gnd.n1850 gnd.n1849 99.6594
R14916 gnd.n1946 gnd.n1945 99.6594
R14917 gnd.n1943 gnd.n1942 99.6594
R14918 gnd.n1938 gnd.n1858 99.6594
R14919 gnd.n1936 gnd.n1935 99.6594
R14920 gnd.n1868 gnd.n1867 99.6594
R14921 gnd.n1927 gnd.n1926 99.6594
R14922 gnd.n1924 gnd.n1923 99.6594
R14923 gnd.n1919 gnd.n1876 99.6594
R14924 gnd.n1917 gnd.n1916 99.6594
R14925 gnd.n1912 gnd.n1883 99.6594
R14926 gnd.n1910 gnd.n1909 99.6594
R14927 gnd.n1905 gnd.n1890 99.6594
R14928 gnd.n1903 gnd.n1902 99.6594
R14929 gnd.n1898 gnd.n1896 99.6594
R14930 gnd.n6402 gnd.n841 99.6594
R14931 gnd.n3975 gnd.n2411 99.6594
R14932 gnd.n3983 gnd.n3982 99.6594
R14933 gnd.n3986 gnd.n3985 99.6594
R14934 gnd.n3993 gnd.n3992 99.6594
R14935 gnd.n3996 gnd.n3995 99.6594
R14936 gnd.n4003 gnd.n4002 99.6594
R14937 gnd.n4006 gnd.n4005 99.6594
R14938 gnd.n4013 gnd.n4012 99.6594
R14939 gnd.n4016 gnd.n4015 99.6594
R14940 gnd.n4023 gnd.n4022 99.6594
R14941 gnd.n4026 gnd.n4025 99.6594
R14942 gnd.n4033 gnd.n4032 99.6594
R14943 gnd.n4036 gnd.n4035 99.6594
R14944 gnd.n4043 gnd.n4042 99.6594
R14945 gnd.n4046 gnd.n4045 99.6594
R14946 gnd.n4053 gnd.n4052 99.6594
R14947 gnd.n4056 gnd.n4055 99.6594
R14948 gnd.n4063 gnd.n4062 99.6594
R14949 gnd.n4066 gnd.n4065 99.6594
R14950 gnd.n4075 gnd.n4074 99.6594
R14951 gnd.n4078 gnd.n4077 99.6594
R14952 gnd.n4085 gnd.n4084 99.6594
R14953 gnd.n4088 gnd.n4087 99.6594
R14954 gnd.n4095 gnd.n4094 99.6594
R14955 gnd.n4098 gnd.n4097 99.6594
R14956 gnd.n4105 gnd.n4104 99.6594
R14957 gnd.n4108 gnd.n4107 99.6594
R14958 gnd.n4116 gnd.n4115 99.6594
R14959 gnd.n4119 gnd.n4118 99.6594
R14960 gnd.n3896 gnd.n2434 99.6594
R14961 gnd.n3894 gnd.n2433 99.6594
R14962 gnd.n3890 gnd.n2432 99.6594
R14963 gnd.n3886 gnd.n2431 99.6594
R14964 gnd.n3882 gnd.n2430 99.6594
R14965 gnd.n3878 gnd.n2429 99.6594
R14966 gnd.n3874 gnd.n2428 99.6594
R14967 gnd.n3806 gnd.n2427 99.6594
R14968 gnd.n3137 gnd.n2868 99.6594
R14969 gnd.n2894 gnd.n2875 99.6594
R14970 gnd.n2896 gnd.n2876 99.6594
R14971 gnd.n2904 gnd.n2877 99.6594
R14972 gnd.n2906 gnd.n2878 99.6594
R14973 gnd.n2914 gnd.n2879 99.6594
R14974 gnd.n2916 gnd.n2880 99.6594
R14975 gnd.n2924 gnd.n2881 99.6594
R14976 gnd.n3864 gnd.n2414 99.6594
R14977 gnd.n3860 gnd.n2415 99.6594
R14978 gnd.n3856 gnd.n2416 99.6594
R14979 gnd.n3852 gnd.n2417 99.6594
R14980 gnd.n3848 gnd.n2418 99.6594
R14981 gnd.n3844 gnd.n2419 99.6594
R14982 gnd.n3840 gnd.n2420 99.6594
R14983 gnd.n3836 gnd.n2421 99.6594
R14984 gnd.n3832 gnd.n2422 99.6594
R14985 gnd.n3828 gnd.n2423 99.6594
R14986 gnd.n3824 gnd.n2424 99.6594
R14987 gnd.n3820 gnd.n2425 99.6594
R14988 gnd.n3816 gnd.n2426 99.6594
R14989 gnd.n3052 gnd.n3051 99.6594
R14990 gnd.n3046 gnd.n2963 99.6594
R14991 gnd.n3043 gnd.n2964 99.6594
R14992 gnd.n3039 gnd.n2965 99.6594
R14993 gnd.n3035 gnd.n2966 99.6594
R14994 gnd.n3031 gnd.n2967 99.6594
R14995 gnd.n3027 gnd.n2968 99.6594
R14996 gnd.n3023 gnd.n2969 99.6594
R14997 gnd.n3019 gnd.n2970 99.6594
R14998 gnd.n3015 gnd.n2971 99.6594
R14999 gnd.n3011 gnd.n2972 99.6594
R15000 gnd.n3007 gnd.n2973 99.6594
R15001 gnd.n3054 gnd.n2962 99.6594
R15002 gnd.n2094 gnd.n2093 99.6594
R15003 gnd.n2097 gnd.n2096 99.6594
R15004 gnd.n2109 gnd.n2108 99.6594
R15005 gnd.n2120 gnd.n2119 99.6594
R15006 gnd.n2123 gnd.n2122 99.6594
R15007 gnd.n2135 gnd.n2134 99.6594
R15008 gnd.n2146 gnd.n2145 99.6594
R15009 gnd.n2149 gnd.n2148 99.6594
R15010 gnd.n4942 gnd.n4941 99.6594
R15011 gnd.n4247 gnd.n3910 99.6594
R15012 gnd.n4246 gnd.n4245 99.6594
R15013 gnd.n4239 gnd.n4125 99.6594
R15014 gnd.n4238 gnd.n4237 99.6594
R15015 gnd.n4231 gnd.n4131 99.6594
R15016 gnd.n4230 gnd.n4229 99.6594
R15017 gnd.n4223 gnd.n4137 99.6594
R15018 gnd.n4222 gnd.n4221 99.6594
R15019 gnd.n4211 gnd.n4143 99.6594
R15020 gnd.n4248 gnd.n4247 99.6594
R15021 gnd.n4245 gnd.n4244 99.6594
R15022 gnd.n4240 gnd.n4239 99.6594
R15023 gnd.n4237 gnd.n4236 99.6594
R15024 gnd.n4232 gnd.n4231 99.6594
R15025 gnd.n4229 gnd.n4228 99.6594
R15026 gnd.n4224 gnd.n4223 99.6594
R15027 gnd.n4221 gnd.n4220 99.6594
R15028 gnd.n4212 gnd.n4211 99.6594
R15029 gnd.n3052 gnd.n2975 99.6594
R15030 gnd.n3044 gnd.n2963 99.6594
R15031 gnd.n3040 gnd.n2964 99.6594
R15032 gnd.n3036 gnd.n2965 99.6594
R15033 gnd.n3032 gnd.n2966 99.6594
R15034 gnd.n3028 gnd.n2967 99.6594
R15035 gnd.n3024 gnd.n2968 99.6594
R15036 gnd.n3020 gnd.n2969 99.6594
R15037 gnd.n3016 gnd.n2970 99.6594
R15038 gnd.n3012 gnd.n2971 99.6594
R15039 gnd.n3008 gnd.n2972 99.6594
R15040 gnd.n3004 gnd.n2973 99.6594
R15041 gnd.n3055 gnd.n3054 99.6594
R15042 gnd.n3819 gnd.n2426 99.6594
R15043 gnd.n3823 gnd.n2425 99.6594
R15044 gnd.n3827 gnd.n2424 99.6594
R15045 gnd.n3831 gnd.n2423 99.6594
R15046 gnd.n3835 gnd.n2422 99.6594
R15047 gnd.n3839 gnd.n2421 99.6594
R15048 gnd.n3843 gnd.n2420 99.6594
R15049 gnd.n3847 gnd.n2419 99.6594
R15050 gnd.n3851 gnd.n2418 99.6594
R15051 gnd.n3855 gnd.n2417 99.6594
R15052 gnd.n3859 gnd.n2416 99.6594
R15053 gnd.n3863 gnd.n2415 99.6594
R15054 gnd.n2455 gnd.n2414 99.6594
R15055 gnd.n3138 gnd.n3137 99.6594
R15056 gnd.n2897 gnd.n2875 99.6594
R15057 gnd.n2903 gnd.n2876 99.6594
R15058 gnd.n2907 gnd.n2877 99.6594
R15059 gnd.n2913 gnd.n2878 99.6594
R15060 gnd.n2917 gnd.n2879 99.6594
R15061 gnd.n2923 gnd.n2880 99.6594
R15062 gnd.n2881 gnd.n2865 99.6594
R15063 gnd.n3873 gnd.n2427 99.6594
R15064 gnd.n3877 gnd.n2428 99.6594
R15065 gnd.n3881 gnd.n2429 99.6594
R15066 gnd.n3885 gnd.n2430 99.6594
R15067 gnd.n3889 gnd.n2431 99.6594
R15068 gnd.n3893 gnd.n2432 99.6594
R15069 gnd.n3897 gnd.n2433 99.6594
R15070 gnd.n2436 gnd.n2434 99.6594
R15071 gnd.n3976 gnd.n3975 99.6594
R15072 gnd.n3984 gnd.n3983 99.6594
R15073 gnd.n3985 gnd.n3968 99.6594
R15074 gnd.n3994 gnd.n3993 99.6594
R15075 gnd.n3995 gnd.n3964 99.6594
R15076 gnd.n4004 gnd.n4003 99.6594
R15077 gnd.n4005 gnd.n3960 99.6594
R15078 gnd.n4014 gnd.n4013 99.6594
R15079 gnd.n4015 gnd.n3953 99.6594
R15080 gnd.n4024 gnd.n4023 99.6594
R15081 gnd.n4025 gnd.n3949 99.6594
R15082 gnd.n4034 gnd.n4033 99.6594
R15083 gnd.n4035 gnd.n3945 99.6594
R15084 gnd.n4044 gnd.n4043 99.6594
R15085 gnd.n4045 gnd.n3941 99.6594
R15086 gnd.n4054 gnd.n4053 99.6594
R15087 gnd.n4055 gnd.n3937 99.6594
R15088 gnd.n4064 gnd.n4063 99.6594
R15089 gnd.n4065 gnd.n3933 99.6594
R15090 gnd.n4076 gnd.n4075 99.6594
R15091 gnd.n4077 gnd.n3929 99.6594
R15092 gnd.n4086 gnd.n4085 99.6594
R15093 gnd.n4087 gnd.n3925 99.6594
R15094 gnd.n4096 gnd.n4095 99.6594
R15095 gnd.n4097 gnd.n3921 99.6594
R15096 gnd.n4106 gnd.n4105 99.6594
R15097 gnd.n4107 gnd.n3917 99.6594
R15098 gnd.n4117 gnd.n4116 99.6594
R15099 gnd.n4120 gnd.n4119 99.6594
R15100 gnd.n4658 gnd.n4657 99.6594
R15101 gnd.n4660 gnd.n4650 99.6594
R15102 gnd.n4669 gnd.n4668 99.6594
R15103 gnd.n4670 gnd.n4646 99.6594
R15104 gnd.n4679 gnd.n4678 99.6594
R15105 gnd.n4680 gnd.n4642 99.6594
R15106 gnd.n4689 gnd.n4688 99.6594
R15107 gnd.n4690 gnd.n4638 99.6594
R15108 gnd.n4699 gnd.n4698 99.6594
R15109 gnd.n4700 gnd.n4634 99.6594
R15110 gnd.n4709 gnd.n4708 99.6594
R15111 gnd.n4710 gnd.n4630 99.6594
R15112 gnd.n4719 gnd.n4718 99.6594
R15113 gnd.n4720 gnd.n4626 99.6594
R15114 gnd.n4729 gnd.n4728 99.6594
R15115 gnd.n4730 gnd.n4622 99.6594
R15116 gnd.n4739 gnd.n4738 99.6594
R15117 gnd.n4740 gnd.n4618 99.6594
R15118 gnd.n4749 gnd.n4748 99.6594
R15119 gnd.n4750 gnd.n4614 99.6594
R15120 gnd.n4759 gnd.n4758 99.6594
R15121 gnd.n4760 gnd.n4610 99.6594
R15122 gnd.n4769 gnd.n4768 99.6594
R15123 gnd.n4770 gnd.n4606 99.6594
R15124 gnd.n4779 gnd.n4778 99.6594
R15125 gnd.n4780 gnd.n4602 99.6594
R15126 gnd.n4789 gnd.n4788 99.6594
R15127 gnd.n4790 gnd.n4598 99.6594
R15128 gnd.n4799 gnd.n4798 99.6594
R15129 gnd.n4800 gnd.n4594 99.6594
R15130 gnd.n4809 gnd.n4808 99.6594
R15131 gnd.n4810 gnd.n4590 99.6594
R15132 gnd.n4819 gnd.n4818 99.6594
R15133 gnd.n4820 gnd.n4586 99.6594
R15134 gnd.n4829 gnd.n4828 99.6594
R15135 gnd.n4830 gnd.n4582 99.6594
R15136 gnd.n4839 gnd.n4838 99.6594
R15137 gnd.n4840 gnd.n4578 99.6594
R15138 gnd.n4849 gnd.n4848 99.6594
R15139 gnd.n4850 gnd.n4574 99.6594
R15140 gnd.n4860 gnd.n4859 99.6594
R15141 gnd.n4861 gnd.n4571 99.6594
R15142 gnd.n4941 gnd.n4940 99.6594
R15143 gnd.n2148 gnd.n2147 99.6594
R15144 gnd.n2145 gnd.n2136 99.6594
R15145 gnd.n2134 gnd.n2133 99.6594
R15146 gnd.n2122 gnd.n2121 99.6594
R15147 gnd.n2119 gnd.n2110 99.6594
R15148 gnd.n2108 gnd.n2107 99.6594
R15149 gnd.n2096 gnd.n2095 99.6594
R15150 gnd.n2093 gnd.n2081 99.6594
R15151 gnd.n6014 gnd.n1060 99.6594
R15152 gnd.n6022 gnd.n1061 99.6594
R15153 gnd.n6024 gnd.n1062 99.6594
R15154 gnd.n6034 gnd.n1063 99.6594
R15155 gnd.n6042 gnd.n1064 99.6594
R15156 gnd.n6044 gnd.n1065 99.6594
R15157 gnd.n6054 gnd.n1066 99.6594
R15158 gnd.n1068 gnd.n1067 99.6594
R15159 gnd.n6217 gnd.n6216 99.6594
R15160 gnd.n7318 gnd.n7315 99.6594
R15161 gnd.n7402 gnd.n7401 99.6594
R15162 gnd.n7314 gnd.n7308 99.6594
R15163 gnd.n7409 gnd.n7408 99.6594
R15164 gnd.n7307 gnd.n7301 99.6594
R15165 gnd.n7416 gnd.n7415 99.6594
R15166 gnd.n7300 gnd.n7294 99.6594
R15167 gnd.n7423 gnd.n7422 99.6594
R15168 gnd.n7293 gnd.n7290 99.6594
R15169 gnd.n1897 gnd.n841 99.6594
R15170 gnd.n1896 gnd.n1891 99.6594
R15171 gnd.n1904 gnd.n1903 99.6594
R15172 gnd.n1890 gnd.n1884 99.6594
R15173 gnd.n1911 gnd.n1910 99.6594
R15174 gnd.n1883 gnd.n1877 99.6594
R15175 gnd.n1918 gnd.n1917 99.6594
R15176 gnd.n1876 gnd.n1870 99.6594
R15177 gnd.n1925 gnd.n1924 99.6594
R15178 gnd.n1928 gnd.n1927 99.6594
R15179 gnd.n1867 gnd.n1859 99.6594
R15180 gnd.n1937 gnd.n1936 99.6594
R15181 gnd.n1858 gnd.n1852 99.6594
R15182 gnd.n1944 gnd.n1943 99.6594
R15183 gnd.n1947 gnd.n1946 99.6594
R15184 gnd.n1842 gnd.n1841 99.6594
R15185 gnd.n1840 gnd.n1839 99.6594
R15186 gnd.n1831 gnd.n1755 99.6594
R15187 gnd.n1830 gnd.n1829 99.6594
R15188 gnd.n1823 gnd.n1759 99.6594
R15189 gnd.n1821 gnd.n1820 99.6594
R15190 gnd.n1814 gnd.n1813 99.6594
R15191 gnd.n1811 gnd.n1810 99.6594
R15192 gnd.n1804 gnd.n1803 99.6594
R15193 gnd.n1801 gnd.n1800 99.6594
R15194 gnd.n1794 gnd.n1793 99.6594
R15195 gnd.n1791 gnd.n1790 99.6594
R15196 gnd.n1784 gnd.n1783 99.6594
R15197 gnd.n6214 gnd.n1071 99.6594
R15198 gnd.n6206 gnd.n1032 99.6594
R15199 gnd.n6202 gnd.n1033 99.6594
R15200 gnd.n6198 gnd.n1034 99.6594
R15201 gnd.n6194 gnd.n1035 99.6594
R15202 gnd.n6190 gnd.n1036 99.6594
R15203 gnd.n6186 gnd.n1037 99.6594
R15204 gnd.n6182 gnd.n1038 99.6594
R15205 gnd.n6177 gnd.n1039 99.6594
R15206 gnd.n6173 gnd.n1040 99.6594
R15207 gnd.n6169 gnd.n1041 99.6594
R15208 gnd.n6165 gnd.n1042 99.6594
R15209 gnd.n6160 gnd.n1044 99.6594
R15210 gnd.n6156 gnd.n1045 99.6594
R15211 gnd.n6152 gnd.n1046 99.6594
R15212 gnd.n6148 gnd.n1047 99.6594
R15213 gnd.n6144 gnd.n1048 99.6594
R15214 gnd.n6140 gnd.n1049 99.6594
R15215 gnd.n6136 gnd.n1050 99.6594
R15216 gnd.n6132 gnd.n1051 99.6594
R15217 gnd.n6128 gnd.n1052 99.6594
R15218 gnd.n6124 gnd.n1053 99.6594
R15219 gnd.n6120 gnd.n1054 99.6594
R15220 gnd.n6116 gnd.n1055 99.6594
R15221 gnd.n6112 gnd.n1056 99.6594
R15222 gnd.n6108 gnd.n1057 99.6594
R15223 gnd.n6104 gnd.n1058 99.6594
R15224 gnd.n1152 gnd.n1059 99.6594
R15225 gnd.n7637 gnd.n7636 99.6594
R15226 gnd.n7628 gnd.n7433 99.6594
R15227 gnd.n7627 gnd.n7626 99.6594
R15228 gnd.n7618 gnd.n7437 99.6594
R15229 gnd.n7617 gnd.n7616 99.6594
R15230 gnd.n7608 gnd.n7441 99.6594
R15231 gnd.n7607 gnd.n7606 99.6594
R15232 gnd.n7598 gnd.n7445 99.6594
R15233 gnd.n7597 gnd.n7596 99.6594
R15234 gnd.n7588 gnd.n7449 99.6594
R15235 gnd.n7587 gnd.n7586 99.6594
R15236 gnd.n7578 gnd.n7455 99.6594
R15237 gnd.n7577 gnd.n7576 99.6594
R15238 gnd.n7568 gnd.n7459 99.6594
R15239 gnd.n7567 gnd.n7566 99.6594
R15240 gnd.n7558 gnd.n7463 99.6594
R15241 gnd.n7557 gnd.n7556 99.6594
R15242 gnd.n7548 gnd.n7467 99.6594
R15243 gnd.n7547 gnd.n7546 99.6594
R15244 gnd.n7538 gnd.n7471 99.6594
R15245 gnd.n7537 gnd.n7536 99.6594
R15246 gnd.n7528 gnd.n7527 99.6594
R15247 gnd.n7526 gnd.n7525 99.6594
R15248 gnd.n7517 gnd.n7481 99.6594
R15249 gnd.n7516 gnd.n7515 99.6594
R15250 gnd.n7507 gnd.n7485 99.6594
R15251 gnd.n7506 gnd.n7505 99.6594
R15252 gnd.n7497 gnd.n7489 99.6594
R15253 gnd.n7496 gnd.n7495 99.6594
R15254 gnd.n5007 gnd.n5006 99.6594
R15255 gnd.n2072 gnd.n2069 99.6594
R15256 gnd.n2075 gnd.n2074 99.6594
R15257 gnd.n2085 gnd.n2077 99.6594
R15258 gnd.n2088 gnd.n2087 99.6594
R15259 gnd.n2100 gnd.n2090 99.6594
R15260 gnd.n2103 gnd.n2102 99.6594
R15261 gnd.n2114 gnd.n2113 99.6594
R15262 gnd.n2126 gnd.n2116 99.6594
R15263 gnd.n2129 gnd.n2128 99.6594
R15264 gnd.n2140 gnd.n2139 99.6594
R15265 gnd.n2157 gnd.n2142 99.6594
R15266 gnd.n2160 gnd.n2159 99.6594
R15267 gnd.n2163 gnd.n2162 99.6594
R15268 gnd.n5006 gnd.n5005 99.6594
R15269 gnd.n2073 gnd.n2072 99.6594
R15270 gnd.n2076 gnd.n2075 99.6594
R15271 gnd.n2086 gnd.n2085 99.6594
R15272 gnd.n2089 gnd.n2088 99.6594
R15273 gnd.n2101 gnd.n2100 99.6594
R15274 gnd.n2104 gnd.n2103 99.6594
R15275 gnd.n2115 gnd.n2114 99.6594
R15276 gnd.n2127 gnd.n2126 99.6594
R15277 gnd.n2130 gnd.n2129 99.6594
R15278 gnd.n2141 gnd.n2140 99.6594
R15279 gnd.n2158 gnd.n2157 99.6594
R15280 gnd.n2161 gnd.n2160 99.6594
R15281 gnd.n2162 gnd.n864 99.6594
R15282 gnd.n5895 gnd.n998 99.6594
R15283 gnd.n5899 gnd.n999 99.6594
R15284 gnd.n5902 gnd.n1000 99.6594
R15285 gnd.n1142 gnd.n1001 99.6594
R15286 gnd.n1144 gnd.n1002 99.6594
R15287 gnd.n6018 gnd.n1003 99.6594
R15288 gnd.n6028 gnd.n1004 99.6594
R15289 gnd.n6030 gnd.n1005 99.6594
R15290 gnd.n6038 gnd.n1006 99.6594
R15291 gnd.n6048 gnd.n1007 99.6594
R15292 gnd.n6050 gnd.n1008 99.6594
R15293 gnd.n1012 gnd.n1009 99.6594
R15294 gnd.n1013 gnd.n1010 99.6594
R15295 gnd.n6227 gnd.n996 99.6594
R15296 gnd.n6051 gnd.n1009 99.6594
R15297 gnd.n6049 gnd.n1008 99.6594
R15298 gnd.n6039 gnd.n1007 99.6594
R15299 gnd.n6031 gnd.n1006 99.6594
R15300 gnd.n6029 gnd.n1005 99.6594
R15301 gnd.n6019 gnd.n1004 99.6594
R15302 gnd.n1145 gnd.n1003 99.6594
R15303 gnd.n1143 gnd.n1002 99.6594
R15304 gnd.n5901 gnd.n1001 99.6594
R15305 gnd.n5900 gnd.n1000 99.6594
R15306 gnd.n5896 gnd.n999 99.6594
R15307 gnd.n1168 gnd.n998 99.6594
R15308 gnd.n6228 gnd.n6227 99.6594
R15309 gnd.n1026 gnd.n1010 99.6594
R15310 gnd.n2154 gnd.t77 98.63
R15311 gnd.n6218 gnd.t37 98.63
R15312 gnd.n7430 gnd.t54 98.63
R15313 gnd.n7452 gnd.t61 98.63
R15314 gnd.n7474 gnd.t85 98.63
R15315 gnd.n1091 gnd.t124 98.63
R15316 gnd.n1114 gnd.t127 98.63
R15317 gnd.n1136 gnd.t89 98.63
R15318 gnd.n7321 gnd.t132 98.63
R15319 gnd.n2150 gnd.t65 98.63
R15320 gnd.n4146 gnd.t73 98.63
R15321 gnd.n3957 gnd.t80 98.63
R15322 gnd.n4067 gnd.t102 98.63
R15323 gnd.n3913 gnd.t121 98.63
R15324 gnd.n1760 gnd.t94 98.63
R15325 gnd.n838 gnd.t111 98.63
R15326 gnd.n1863 gnd.t139 98.63
R15327 gnd.n1015 gnd.t40 98.63
R15328 gnd.n1687 gnd.t99 92.8196
R15329 gnd.n1282 gnd.t117 92.8196
R15330 gnd.n1689 gnd.t146 92.8118
R15331 gnd.n1276 gnd.t47 92.8118
R15332 gnd.n1641 gnd.n1640 81.8399
R15333 gnd.n2926 gnd.t58 74.8376
R15334 gnd.n2452 gnd.t109 74.8376
R15335 gnd.n1688 gnd.t98 72.8438
R15336 gnd.n1283 gnd.t118 72.8438
R15337 gnd.n1642 gnd.n1635 72.8411
R15338 gnd.n1648 gnd.n1633 72.8411
R15339 gnd.n1247 gnd.n1246 72.8411
R15340 gnd.n2155 gnd.t76 72.836
R15341 gnd.n1690 gnd.t145 72.836
R15342 gnd.n1277 gnd.t48 72.836
R15343 gnd.n6219 gnd.t36 72.836
R15344 gnd.n7431 gnd.t55 72.836
R15345 gnd.n7453 gnd.t62 72.836
R15346 gnd.n7475 gnd.t86 72.836
R15347 gnd.n1092 gnd.t123 72.836
R15348 gnd.n1115 gnd.t126 72.836
R15349 gnd.n1137 gnd.t88 72.836
R15350 gnd.n7322 gnd.t133 72.836
R15351 gnd.n2151 gnd.t66 72.836
R15352 gnd.n4147 gnd.t72 72.836
R15353 gnd.n3958 gnd.t79 72.836
R15354 gnd.n4068 gnd.t101 72.836
R15355 gnd.n3914 gnd.t120 72.836
R15356 gnd.n1761 gnd.t95 72.836
R15357 gnd.n839 gnd.t112 72.836
R15358 gnd.n1864 gnd.t140 72.836
R15359 gnd.n1016 gnd.t41 72.836
R15360 gnd.n5801 gnd.n5800 71.676
R15361 gnd.n5796 gnd.n1256 71.676
R15362 gnd.n5794 gnd.n5793 71.676
R15363 gnd.n5789 gnd.n1259 71.676
R15364 gnd.n5787 gnd.n5786 71.676
R15365 gnd.n5782 gnd.n1262 71.676
R15366 gnd.n5780 gnd.n5779 71.676
R15367 gnd.n5775 gnd.n1265 71.676
R15368 gnd.n5773 gnd.n5772 71.676
R15369 gnd.n5768 gnd.n1268 71.676
R15370 gnd.n5766 gnd.n5765 71.676
R15371 gnd.n5761 gnd.n1271 71.676
R15372 gnd.n5759 gnd.n5758 71.676
R15373 gnd.n5754 gnd.n1274 71.676
R15374 gnd.n5752 gnd.n5751 71.676
R15375 gnd.n5747 gnd.n1279 71.676
R15376 gnd.n5744 gnd.n5743 71.676
R15377 gnd.n5741 gnd.n5740 71.676
R15378 gnd.n5735 gnd.n1285 71.676
R15379 gnd.n5733 gnd.n5732 71.676
R15380 gnd.n5728 gnd.n1288 71.676
R15381 gnd.n5726 gnd.n5725 71.676
R15382 gnd.n5721 gnd.n1291 71.676
R15383 gnd.n5719 gnd.n5718 71.676
R15384 gnd.n5714 gnd.n1294 71.676
R15385 gnd.n5712 gnd.n5711 71.676
R15386 gnd.n5707 gnd.n1297 71.676
R15387 gnd.n5705 gnd.n5704 71.676
R15388 gnd.n5700 gnd.n1300 71.676
R15389 gnd.n5698 gnd.n5697 71.676
R15390 gnd.n5693 gnd.n1303 71.676
R15391 gnd.n5691 gnd.n5690 71.676
R15392 gnd.n5686 gnd.n1306 71.676
R15393 gnd.n5152 gnd.n1631 71.676
R15394 gnd.n1692 gnd.n1655 71.676
R15395 gnd.n1696 gnd.n1656 71.676
R15396 gnd.n1700 gnd.n1657 71.676
R15397 gnd.n1704 gnd.n1658 71.676
R15398 gnd.n1708 gnd.n1659 71.676
R15399 gnd.n1712 gnd.n1660 71.676
R15400 gnd.n1716 gnd.n1661 71.676
R15401 gnd.n1720 gnd.n1662 71.676
R15402 gnd.n1724 gnd.n1663 71.676
R15403 gnd.n1728 gnd.n1664 71.676
R15404 gnd.n1732 gnd.n1665 71.676
R15405 gnd.n1736 gnd.n1666 71.676
R15406 gnd.n1740 gnd.n1667 71.676
R15407 gnd.n1744 gnd.n1668 71.676
R15408 gnd.n1748 gnd.n1669 71.676
R15409 gnd.n1956 gnd.n1671 71.676
R15410 gnd.n1960 gnd.n1672 71.676
R15411 gnd.n1965 gnd.n1673 71.676
R15412 gnd.n1969 gnd.n1674 71.676
R15413 gnd.n1973 gnd.n1675 71.676
R15414 gnd.n1977 gnd.n1676 71.676
R15415 gnd.n1981 gnd.n1677 71.676
R15416 gnd.n1985 gnd.n1678 71.676
R15417 gnd.n1989 gnd.n1679 71.676
R15418 gnd.n1993 gnd.n1680 71.676
R15419 gnd.n1997 gnd.n1681 71.676
R15420 gnd.n2001 gnd.n1682 71.676
R15421 gnd.n2005 gnd.n1683 71.676
R15422 gnd.n2009 gnd.n1684 71.676
R15423 gnd.n2013 gnd.n1685 71.676
R15424 gnd.n2024 gnd.n1686 71.676
R15425 gnd.n5153 gnd.n5152 71.676
R15426 gnd.n1695 gnd.n1655 71.676
R15427 gnd.n1699 gnd.n1656 71.676
R15428 gnd.n1703 gnd.n1657 71.676
R15429 gnd.n1707 gnd.n1658 71.676
R15430 gnd.n1711 gnd.n1659 71.676
R15431 gnd.n1715 gnd.n1660 71.676
R15432 gnd.n1719 gnd.n1661 71.676
R15433 gnd.n1723 gnd.n1662 71.676
R15434 gnd.n1727 gnd.n1663 71.676
R15435 gnd.n1731 gnd.n1664 71.676
R15436 gnd.n1735 gnd.n1665 71.676
R15437 gnd.n1739 gnd.n1666 71.676
R15438 gnd.n1743 gnd.n1667 71.676
R15439 gnd.n1747 gnd.n1668 71.676
R15440 gnd.n1955 gnd.n1670 71.676
R15441 gnd.n1959 gnd.n1671 71.676
R15442 gnd.n1964 gnd.n1672 71.676
R15443 gnd.n1968 gnd.n1673 71.676
R15444 gnd.n1972 gnd.n1674 71.676
R15445 gnd.n1976 gnd.n1675 71.676
R15446 gnd.n1980 gnd.n1676 71.676
R15447 gnd.n1984 gnd.n1677 71.676
R15448 gnd.n1988 gnd.n1678 71.676
R15449 gnd.n1992 gnd.n1679 71.676
R15450 gnd.n1996 gnd.n1680 71.676
R15451 gnd.n2000 gnd.n1681 71.676
R15452 gnd.n2004 gnd.n1682 71.676
R15453 gnd.n2008 gnd.n1683 71.676
R15454 gnd.n2012 gnd.n1684 71.676
R15455 gnd.n2015 gnd.n1685 71.676
R15456 gnd.n2024 gnd.n2023 71.676
R15457 gnd.n1306 gnd.n1304 71.676
R15458 gnd.n5692 gnd.n5691 71.676
R15459 gnd.n1303 gnd.n1301 71.676
R15460 gnd.n5699 gnd.n5698 71.676
R15461 gnd.n1300 gnd.n1298 71.676
R15462 gnd.n5706 gnd.n5705 71.676
R15463 gnd.n1297 gnd.n1295 71.676
R15464 gnd.n5713 gnd.n5712 71.676
R15465 gnd.n1294 gnd.n1292 71.676
R15466 gnd.n5720 gnd.n5719 71.676
R15467 gnd.n1291 gnd.n1289 71.676
R15468 gnd.n5727 gnd.n5726 71.676
R15469 gnd.n1288 gnd.n1286 71.676
R15470 gnd.n5734 gnd.n5733 71.676
R15471 gnd.n1285 gnd.n1281 71.676
R15472 gnd.n5742 gnd.n5741 71.676
R15473 gnd.n5746 gnd.n5745 71.676
R15474 gnd.n1279 gnd.n1275 71.676
R15475 gnd.n5753 gnd.n5752 71.676
R15476 gnd.n1274 gnd.n1272 71.676
R15477 gnd.n5760 gnd.n5759 71.676
R15478 gnd.n1271 gnd.n1269 71.676
R15479 gnd.n5767 gnd.n5766 71.676
R15480 gnd.n1268 gnd.n1266 71.676
R15481 gnd.n5774 gnd.n5773 71.676
R15482 gnd.n1265 gnd.n1263 71.676
R15483 gnd.n5781 gnd.n5780 71.676
R15484 gnd.n1262 gnd.n1260 71.676
R15485 gnd.n5788 gnd.n5787 71.676
R15486 gnd.n1259 gnd.n1257 71.676
R15487 gnd.n5795 gnd.n5794 71.676
R15488 gnd.n1256 gnd.n1254 71.676
R15489 gnd.n5802 gnd.n5801 71.676
R15490 gnd.n10 gnd.t159 69.1507
R15491 gnd.n18 gnd.t155 68.4792
R15492 gnd.n17 gnd.t18 68.4792
R15493 gnd.n16 gnd.t166 68.4792
R15494 gnd.n15 gnd.t164 68.4792
R15495 gnd.n14 gnd.t209 68.4792
R15496 gnd.n13 gnd.t14 68.4792
R15497 gnd.n12 gnd.t172 68.4792
R15498 gnd.n11 gnd.t415 68.4792
R15499 gnd.n10 gnd.t179 68.4792
R15500 gnd.n6814 gnd.n6813 67.5577
R15501 gnd.n6815 gnd.n6814 67.5577
R15502 gnd.n6815 gnd.n532 67.5577
R15503 gnd.n6823 gnd.n532 67.5577
R15504 gnd.n6824 gnd.n6823 67.5577
R15505 gnd.n6825 gnd.n6824 67.5577
R15506 gnd.n6825 gnd.n526 67.5577
R15507 gnd.n6833 gnd.n526 67.5577
R15508 gnd.n6834 gnd.n6833 67.5577
R15509 gnd.n6835 gnd.n6834 67.5577
R15510 gnd.n6835 gnd.n520 67.5577
R15511 gnd.n6843 gnd.n520 67.5577
R15512 gnd.n6844 gnd.n6843 67.5577
R15513 gnd.n6845 gnd.n6844 67.5577
R15514 gnd.n6845 gnd.n514 67.5577
R15515 gnd.n6853 gnd.n514 67.5577
R15516 gnd.n6854 gnd.n6853 67.5577
R15517 gnd.n6855 gnd.n6854 67.5577
R15518 gnd.n6855 gnd.n508 67.5577
R15519 gnd.n6863 gnd.n508 67.5577
R15520 gnd.n6864 gnd.n6863 67.5577
R15521 gnd.n6865 gnd.n6864 67.5577
R15522 gnd.n6865 gnd.n502 67.5577
R15523 gnd.n6873 gnd.n502 67.5577
R15524 gnd.n6874 gnd.n6873 67.5577
R15525 gnd.n6875 gnd.n6874 67.5577
R15526 gnd.n6875 gnd.n496 67.5577
R15527 gnd.n6883 gnd.n496 67.5577
R15528 gnd.n6884 gnd.n6883 67.5577
R15529 gnd.n6885 gnd.n6884 67.5577
R15530 gnd.n6885 gnd.n490 67.5577
R15531 gnd.n6893 gnd.n490 67.5577
R15532 gnd.n6894 gnd.n6893 67.5577
R15533 gnd.n6895 gnd.n6894 67.5577
R15534 gnd.n6895 gnd.n484 67.5577
R15535 gnd.n6903 gnd.n484 67.5577
R15536 gnd.n6904 gnd.n6903 67.5577
R15537 gnd.n6905 gnd.n6904 67.5577
R15538 gnd.n6905 gnd.n478 67.5577
R15539 gnd.n6913 gnd.n478 67.5577
R15540 gnd.n6914 gnd.n6913 67.5577
R15541 gnd.n6915 gnd.n6914 67.5577
R15542 gnd.n6915 gnd.n472 67.5577
R15543 gnd.n6923 gnd.n472 67.5577
R15544 gnd.n6924 gnd.n6923 67.5577
R15545 gnd.n6925 gnd.n6924 67.5577
R15546 gnd.n6925 gnd.n466 67.5577
R15547 gnd.n6933 gnd.n466 67.5577
R15548 gnd.n6934 gnd.n6933 67.5577
R15549 gnd.n6935 gnd.n6934 67.5577
R15550 gnd.n6935 gnd.n460 67.5577
R15551 gnd.n6943 gnd.n460 67.5577
R15552 gnd.n6944 gnd.n6943 67.5577
R15553 gnd.n6945 gnd.n6944 67.5577
R15554 gnd.n6945 gnd.n454 67.5577
R15555 gnd.n6953 gnd.n454 67.5577
R15556 gnd.n6954 gnd.n6953 67.5577
R15557 gnd.n6955 gnd.n6954 67.5577
R15558 gnd.n6955 gnd.n448 67.5577
R15559 gnd.n6963 gnd.n448 67.5577
R15560 gnd.n6964 gnd.n6963 67.5577
R15561 gnd.n6965 gnd.n6964 67.5577
R15562 gnd.n6965 gnd.n442 67.5577
R15563 gnd.n6973 gnd.n442 67.5577
R15564 gnd.n6974 gnd.n6973 67.5577
R15565 gnd.n6975 gnd.n6974 67.5577
R15566 gnd.n6975 gnd.n436 67.5577
R15567 gnd.n6983 gnd.n436 67.5577
R15568 gnd.n6984 gnd.n6983 67.5577
R15569 gnd.n6985 gnd.n6984 67.5577
R15570 gnd.n6985 gnd.n430 67.5577
R15571 gnd.n6993 gnd.n430 67.5577
R15572 gnd.n6994 gnd.n6993 67.5577
R15573 gnd.n6995 gnd.n6994 67.5577
R15574 gnd.n6995 gnd.n424 67.5577
R15575 gnd.n7003 gnd.n424 67.5577
R15576 gnd.n7004 gnd.n7003 67.5577
R15577 gnd.n7005 gnd.n7004 67.5577
R15578 gnd.n7005 gnd.n418 67.5577
R15579 gnd.n7013 gnd.n418 67.5577
R15580 gnd.n7014 gnd.n7013 67.5577
R15581 gnd.n7016 gnd.n7014 67.5577
R15582 gnd.n7016 gnd.n7015 67.5577
R15583 gnd.n1962 gnd.n1688 59.5399
R15584 gnd.n5737 gnd.n1283 59.5399
R15585 gnd.n1691 gnd.n1690 59.5399
R15586 gnd.n1278 gnd.n1277 59.5399
R15587 gnd.n5156 gnd.n1651 59.1804
R15588 gnd.n6454 gnd.n6453 58.7274
R15589 gnd.n2704 gnd.t365 56.407
R15590 gnd.n2645 gnd.t391 56.407
R15591 gnd.n2664 gnd.t342 56.407
R15592 gnd.n2684 gnd.t235 56.407
R15593 gnd.n80 gnd.t335 56.407
R15594 gnd.n21 gnd.t252 56.407
R15595 gnd.n40 gnd.t321 56.407
R15596 gnd.n60 gnd.t378 56.407
R15597 gnd.n2721 gnd.t395 55.8337
R15598 gnd.n2662 gnd.t221 55.8337
R15599 gnd.n2681 gnd.t239 55.8337
R15600 gnd.n2701 gnd.t307 55.8337
R15601 gnd.n97 gnd.t338 55.8337
R15602 gnd.n38 gnd.t250 55.8337
R15603 gnd.n57 gnd.t390 55.8337
R15604 gnd.n77 gnd.t382 55.8337
R15605 gnd.n1639 gnd.n1638 54.358
R15606 gnd.n1244 gnd.n1243 54.358
R15607 gnd.n2704 gnd.n2703 53.0052
R15608 gnd.n2706 gnd.n2705 53.0052
R15609 gnd.n2708 gnd.n2707 53.0052
R15610 gnd.n2710 gnd.n2709 53.0052
R15611 gnd.n2712 gnd.n2711 53.0052
R15612 gnd.n2714 gnd.n2713 53.0052
R15613 gnd.n2716 gnd.n2715 53.0052
R15614 gnd.n2718 gnd.n2717 53.0052
R15615 gnd.n2720 gnd.n2719 53.0052
R15616 gnd.n2645 gnd.n2644 53.0052
R15617 gnd.n2647 gnd.n2646 53.0052
R15618 gnd.n2649 gnd.n2648 53.0052
R15619 gnd.n2651 gnd.n2650 53.0052
R15620 gnd.n2653 gnd.n2652 53.0052
R15621 gnd.n2655 gnd.n2654 53.0052
R15622 gnd.n2657 gnd.n2656 53.0052
R15623 gnd.n2659 gnd.n2658 53.0052
R15624 gnd.n2661 gnd.n2660 53.0052
R15625 gnd.n2664 gnd.n2663 53.0052
R15626 gnd.n2666 gnd.n2665 53.0052
R15627 gnd.n2668 gnd.n2667 53.0052
R15628 gnd.n2670 gnd.n2669 53.0052
R15629 gnd.n2672 gnd.n2671 53.0052
R15630 gnd.n2674 gnd.n2673 53.0052
R15631 gnd.n2676 gnd.n2675 53.0052
R15632 gnd.n2678 gnd.n2677 53.0052
R15633 gnd.n2680 gnd.n2679 53.0052
R15634 gnd.n2684 gnd.n2683 53.0052
R15635 gnd.n2686 gnd.n2685 53.0052
R15636 gnd.n2688 gnd.n2687 53.0052
R15637 gnd.n2690 gnd.n2689 53.0052
R15638 gnd.n2692 gnd.n2691 53.0052
R15639 gnd.n2694 gnd.n2693 53.0052
R15640 gnd.n2696 gnd.n2695 53.0052
R15641 gnd.n2698 gnd.n2697 53.0052
R15642 gnd.n2700 gnd.n2699 53.0052
R15643 gnd.n96 gnd.n95 53.0052
R15644 gnd.n94 gnd.n93 53.0052
R15645 gnd.n92 gnd.n91 53.0052
R15646 gnd.n90 gnd.n89 53.0052
R15647 gnd.n88 gnd.n87 53.0052
R15648 gnd.n86 gnd.n85 53.0052
R15649 gnd.n84 gnd.n83 53.0052
R15650 gnd.n82 gnd.n81 53.0052
R15651 gnd.n80 gnd.n79 53.0052
R15652 gnd.n37 gnd.n36 53.0052
R15653 gnd.n35 gnd.n34 53.0052
R15654 gnd.n33 gnd.n32 53.0052
R15655 gnd.n31 gnd.n30 53.0052
R15656 gnd.n29 gnd.n28 53.0052
R15657 gnd.n27 gnd.n26 53.0052
R15658 gnd.n25 gnd.n24 53.0052
R15659 gnd.n23 gnd.n22 53.0052
R15660 gnd.n21 gnd.n20 53.0052
R15661 gnd.n56 gnd.n55 53.0052
R15662 gnd.n54 gnd.n53 53.0052
R15663 gnd.n52 gnd.n51 53.0052
R15664 gnd.n50 gnd.n49 53.0052
R15665 gnd.n48 gnd.n47 53.0052
R15666 gnd.n46 gnd.n45 53.0052
R15667 gnd.n44 gnd.n43 53.0052
R15668 gnd.n42 gnd.n41 53.0052
R15669 gnd.n40 gnd.n39 53.0052
R15670 gnd.n76 gnd.n75 53.0052
R15671 gnd.n74 gnd.n73 53.0052
R15672 gnd.n72 gnd.n71 53.0052
R15673 gnd.n70 gnd.n69 53.0052
R15674 gnd.n68 gnd.n67 53.0052
R15675 gnd.n66 gnd.n65 53.0052
R15676 gnd.n64 gnd.n63 53.0052
R15677 gnd.n62 gnd.n61 53.0052
R15678 gnd.n60 gnd.n59 53.0052
R15679 gnd.n1235 gnd.n1234 52.4801
R15680 gnd.n3757 gnd.t213 52.3082
R15681 gnd.n3725 gnd.t25 52.3082
R15682 gnd.n3693 gnd.t150 52.3082
R15683 gnd.n3662 gnd.t174 52.3082
R15684 gnd.n3630 gnd.t181 52.3082
R15685 gnd.n3598 gnd.t157 52.3082
R15686 gnd.n3566 gnd.t176 52.3082
R15687 gnd.n3535 gnd.t207 52.3082
R15688 gnd.n7645 gnd.n253 51.6227
R15689 gnd.n3587 gnd.n3555 51.4173
R15690 gnd.n3651 gnd.n3650 50.455
R15691 gnd.n3619 gnd.n3618 50.455
R15692 gnd.n3587 gnd.n3586 50.455
R15693 gnd.n3000 gnd.n2999 45.1884
R15694 gnd.n2478 gnd.n2477 45.1884
R15695 gnd.n1251 gnd.n1250 44.3322
R15696 gnd.n1642 gnd.n1641 44.3189
R15697 gnd.n2156 gnd.n2155 42.4732
R15698 gnd.n1017 gnd.n1016 42.4732
R15699 gnd.n6220 gnd.n6219 42.2793
R15700 gnd.n7432 gnd.n7431 42.2793
R15701 gnd.n7454 gnd.n7453 42.2793
R15702 gnd.n7476 gnd.n7475 42.2793
R15703 gnd.n6179 gnd.n1092 42.2793
R15704 gnd.n6142 gnd.n1115 42.2793
R15705 gnd.n6102 gnd.n1137 42.2793
R15706 gnd.n7398 gnd.n7322 42.2793
R15707 gnd.n2152 gnd.n2151 42.2793
R15708 gnd.n3001 gnd.n3000 42.2793
R15709 gnd.n2479 gnd.n2478 42.2793
R15710 gnd.n2927 gnd.n2926 42.2793
R15711 gnd.n3872 gnd.n2452 42.2793
R15712 gnd.n4148 gnd.n4147 42.2793
R15713 gnd.n3959 gnd.n3958 42.2793
R15714 gnd.n4069 gnd.n4068 42.2793
R15715 gnd.n3915 gnd.n3914 42.2793
R15716 gnd.n1762 gnd.n1761 42.2793
R15717 gnd.n840 gnd.n839 42.2793
R15718 gnd.n1933 gnd.n1864 42.2793
R15719 gnd.n1640 gnd.n1639 41.6274
R15720 gnd.n1245 gnd.n1244 41.6274
R15721 gnd.n1649 gnd.n1648 40.8975
R15722 gnd.n1248 gnd.n1247 40.8975
R15723 gnd.n7015 gnd.n167 40.5348
R15724 gnd.n3053 gnd.n2957 36.8252
R15725 gnd.n1648 gnd.n1647 35.055
R15726 gnd.n1643 gnd.n1642 35.055
R15727 gnd.n1237 gnd.n1236 35.055
R15728 gnd.n1247 gnd.n1233 35.055
R15729 gnd.n3905 gnd.n2412 32.8146
R15730 gnd.n6399 gnd.n843 31.8661
R15731 gnd.n6393 gnd.n6392 31.8661
R15732 gnd.n6392 gnd.n6391 31.8661
R15733 gnd.n6385 gnd.n861 31.8661
R15734 gnd.n6385 gnd.n863 31.8661
R15735 gnd.n5023 gnd.n5015 31.8661
R15736 gnd.n5023 gnd.n2061 31.8661
R15737 gnd.n5033 gnd.n2061 31.8661
R15738 gnd.n5033 gnd.n5031 31.8661
R15739 gnd.n5041 gnd.n2050 31.8661
R15740 gnd.n5050 gnd.n2050 31.8661
R15741 gnd.n5050 gnd.n2044 31.8661
R15742 gnd.n5058 gnd.n2044 31.8661
R15743 gnd.n5067 gnd.n2038 31.8661
R15744 gnd.n5067 gnd.n2031 31.8661
R15745 gnd.n5077 gnd.n2031 31.8661
R15746 gnd.n5818 gnd.n1220 31.8661
R15747 gnd.n5835 gnd.n1208 31.8661
R15748 gnd.n5835 gnd.n1202 31.8661
R15749 gnd.n5844 gnd.n1202 31.8661
R15750 gnd.n5852 gnd.n1196 31.8661
R15751 gnd.n5852 gnd.n1190 31.8661
R15752 gnd.n5862 gnd.n1190 31.8661
R15753 gnd.n5862 gnd.n5860 31.8661
R15754 gnd.n5870 gnd.n1179 31.8661
R15755 gnd.n5879 gnd.n1179 31.8661
R15756 gnd.n5879 gnd.n1173 31.8661
R15757 gnd.n5889 gnd.n1173 31.8661
R15758 gnd.n5915 gnd.n1166 31.8661
R15759 gnd.n5915 gnd.n997 31.8661
R15760 gnd.n5923 gnd.n1011 31.8661
R15761 gnd.n5923 gnd.n1031 31.8661
R15762 gnd.n1151 gnd.n1069 31.8661
R15763 gnd.n7137 gnd.n338 31.8661
R15764 gnd.n7145 gnd.n318 31.8661
R15765 gnd.n7157 gnd.n318 31.8661
R15766 gnd.n7165 gnd.n310 31.8661
R15767 gnd.n7181 gnd.n298 31.8661
R15768 gnd.n7181 gnd.n301 31.8661
R15769 gnd.n7191 gnd.n283 31.8661
R15770 gnd.n7204 gnd.n283 31.8661
R15771 gnd.n7213 gnd.n277 31.8661
R15772 gnd.n7224 gnd.n260 31.8661
R15773 gnd.n7232 gnd.n260 31.8661
R15774 gnd.n7735 gnd.n106 31.8661
R15775 gnd.n7729 gnd.n118 31.8661
R15776 gnd.n7723 gnd.n118 31.8661
R15777 gnd.n7717 gnd.n136 31.8661
R15778 gnd.n7717 gnd.n139 31.8661
R15779 gnd.n7711 gnd.n148 31.8661
R15780 gnd.n7705 gnd.n158 31.8661
R15781 gnd.n7699 gnd.n158 31.8661
R15782 gnd.n7693 gnd.n175 31.8661
R15783 gnd.n7693 gnd.n178 31.8661
R15784 gnd.n7687 gnd.n187 31.8661
R15785 gnd.n7681 gnd.n197 31.8661
R15786 gnd.n7675 gnd.n197 31.8661
R15787 gnd.n7669 gnd.n213 31.8661
R15788 gnd.n7669 gnd.n216 31.8661
R15789 gnd.n7663 gnd.n225 31.8661
R15790 gnd.n7657 gnd.n225 31.8661
R15791 gnd.n7657 gnd.n235 31.8661
R15792 gnd.n7651 gnd.n235 31.8661
R15793 gnd.n7645 gnd.n250 31.8661
R15794 gnd.n7213 gnd.t228 31.5474
R15795 gnd.t216 gnd.n106 31.5474
R15796 gnd.n5687 gnd.n1305 31.3761
R15797 gnd.n2022 gnd.n2021 31.3761
R15798 gnd.n5151 gnd.n1654 30.9101
R15799 gnd.t298 gnd.n310 30.9101
R15800 gnd.t253 gnd.n148 30.9101
R15801 gnd.n5150 gnd.t129 30.5915
R15802 gnd.t354 gnd.n187 30.2728
R15803 gnd.n4262 gnd.n3906 29.5331
R15804 gnd.n250 gnd.t53 28.3609
R15805 gnd.n5077 gnd.t21 27.0862
R15806 gnd.t17 gnd.n1208 27.0862
R15807 gnd.n5827 gnd.t68 26.1303
R15808 gnd.n2155 gnd.n2154 25.7944
R15809 gnd.n6219 gnd.n6218 25.7944
R15810 gnd.n7431 gnd.n7430 25.7944
R15811 gnd.n7453 gnd.n7452 25.7944
R15812 gnd.n7475 gnd.n7474 25.7944
R15813 gnd.n1092 gnd.n1091 25.7944
R15814 gnd.n1115 gnd.n1114 25.7944
R15815 gnd.n1137 gnd.n1136 25.7944
R15816 gnd.n7322 gnd.n7321 25.7944
R15817 gnd.n2151 gnd.n2150 25.7944
R15818 gnd.n2926 gnd.n2925 25.7944
R15819 gnd.n2452 gnd.n2451 25.7944
R15820 gnd.n4147 gnd.n4146 25.7944
R15821 gnd.n3958 gnd.n3957 25.7944
R15822 gnd.n4068 gnd.n4067 25.7944
R15823 gnd.n3914 gnd.n3913 25.7944
R15824 gnd.n1761 gnd.n1760 25.7944
R15825 gnd.n839 gnd.n838 25.7944
R15826 gnd.n1864 gnd.n1863 25.7944
R15827 gnd.n1016 gnd.n1015 25.7944
R15828 gnd.t75 gnd.n863 24.537
R15829 gnd.t158 gnd.n2038 24.537
R15830 gnd.n5844 gnd.t161 24.537
R15831 gnd.t39 gnd.n1166 24.537
R15832 gnd.n6446 gnd.n765 24.2183
R15833 gnd.n6440 gnd.n777 24.2183
R15834 gnd.n4902 gnd.n780 24.2183
R15835 gnd.n4908 gnd.n790 24.2183
R15836 gnd.n6428 gnd.n797 24.2183
R15837 gnd.n6422 gnd.n808 24.2183
R15838 gnd.n4928 gnd.n811 24.2183
R15839 gnd.n6416 gnd.n818 24.2183
R15840 gnd.n4922 gnd.n821 24.2183
R15841 gnd.n6410 gnd.n829 24.2183
R15842 gnd.n6400 gnd.n832 24.2183
R15843 gnd.n6010 gnd.n6009 24.2183
R15844 gnd.n5935 gnd.n1155 24.2183
R15845 gnd.n6003 gnd.n5936 24.2183
R15846 gnd.n6002 gnd.n5939 24.2183
R15847 gnd.n5988 gnd.n5949 24.2183
R15848 gnd.n5981 gnd.n391 24.2183
R15849 gnd.n7038 gnd.n381 24.2183
R15850 gnd.n7061 gnd.n383 24.2183
R15851 gnd.n7070 gnd.n362 24.2183
R15852 gnd.n7087 gnd.n365 24.2183
R15853 gnd.n7097 gnd.n354 24.2183
R15854 gnd.n861 gnd.n853 23.8997
R15855 gnd.n6226 gnd.n997 23.8997
R15856 gnd.n4916 gnd.t234 23.2624
R15857 gnd.n7051 gnd.t251 23.2624
R15858 gnd.n7663 gnd.t249 23.2624
R15859 gnd.t329 gnd.n768 22.6251
R15860 gnd.t268 gnd.n352 22.6251
R15861 gnd.n7080 gnd.t218 22.6251
R15862 gnd.n7687 gnd.t270 22.6251
R15863 gnd.n7165 gnd.t301 21.9878
R15864 gnd.n7711 gnd.t318 21.9878
R15865 gnd.n5159 gnd.n1630 21.6691
R15866 gnd.n5228 gnd.n1580 21.6691
R15867 gnd.n5242 gnd.n5241 21.6691
R15868 gnd.n5269 gnd.n5268 21.6691
R15869 gnd.n5285 gnd.n1541 21.6691
R15870 gnd.n5292 gnd.n1530 21.6691
R15871 gnd.n5312 gnd.n5311 21.6691
R15872 gnd.n5346 gnd.n1510 21.6691
R15873 gnd.n5415 gnd.n1465 21.6691
R15874 gnd.n5502 gnd.n1422 21.6691
R15875 gnd.n5508 gnd.n1402 21.6691
R15876 gnd.n5515 gnd.n1394 21.6691
R15877 gnd.n5522 gnd.n1387 21.6691
R15878 gnd.n5574 gnd.n1379 21.6691
R15879 gnd.n5567 gnd.n5566 21.6691
R15880 gnd.n5634 gnd.n5633 21.6691
R15881 gnd.n5654 gnd.n1321 21.6691
R15882 gnd.n5671 gnd.n1313 21.6691
R15883 gnd.n277 gnd.t247 21.3504
R15884 gnd.n7735 gnd.t230 21.3504
R15885 gnd.n5193 gnd.t82 21.0318
R15886 gnd.n7191 gnd.t266 20.7131
R15887 gnd.n7723 gnd.t236 20.7131
R15888 gnd.n5199 gnd.n1602 20.3945
R15889 gnd.n5218 gnd.n1591 20.3945
R15890 gnd.n5640 gnd.n1332 20.3945
R15891 gnd.t414 gnd.n5234 20.0758
R15892 gnd.n5627 gnd.t200 20.0758
R15893 gnd.n7145 gnd.t214 20.0758
R15894 gnd.n1688 gnd.n1687 19.9763
R15895 gnd.n1283 gnd.n1282 19.9763
R15896 gnd.n1690 gnd.n1689 19.9763
R15897 gnd.n1277 gnd.n1276 19.9763
R15898 gnd.n1637 gnd.t51 19.8005
R15899 gnd.n1637 gnd.t115 19.8005
R15900 gnd.n1636 gnd.t83 19.8005
R15901 gnd.n1636 gnd.t105 19.8005
R15902 gnd.n1242 gnd.t29 19.8005
R15903 gnd.n1242 gnd.t143 19.8005
R15904 gnd.n1241 gnd.t92 19.8005
R15905 gnd.n1241 gnd.t69 19.8005
R15906 gnd.n6393 gnd.n852 19.7572
R15907 gnd.n6215 gnd.n1031 19.7572
R15908 gnd.n1633 gnd.n1632 19.5087
R15909 gnd.n1646 gnd.n1633 19.5087
R15910 gnd.n1644 gnd.n1635 19.5087
R15911 gnd.n1246 gnd.n1240 19.5087
R15912 gnd.n5031 gnd.t204 19.4385
R15913 gnd.n5870 gnd.t154 19.4385
R15914 gnd.n7675 gnd.t240 19.4385
R15915 gnd.n6383 gnd.n866 19.3944
R15916 gnd.n6379 gnd.n866 19.3944
R15917 gnd.n6379 gnd.n6378 19.3944
R15918 gnd.n6378 gnd.n6377 19.3944
R15919 gnd.n6377 gnd.n872 19.3944
R15920 gnd.n6373 gnd.n872 19.3944
R15921 gnd.n6373 gnd.n6372 19.3944
R15922 gnd.n6372 gnd.n6371 19.3944
R15923 gnd.n6371 gnd.n877 19.3944
R15924 gnd.n6367 gnd.n877 19.3944
R15925 gnd.n6367 gnd.n6366 19.3944
R15926 gnd.n6366 gnd.n6365 19.3944
R15927 gnd.n6365 gnd.n882 19.3944
R15928 gnd.n6361 gnd.n882 19.3944
R15929 gnd.n6361 gnd.n6360 19.3944
R15930 gnd.n6360 gnd.n6359 19.3944
R15931 gnd.n6359 gnd.n887 19.3944
R15932 gnd.n6355 gnd.n887 19.3944
R15933 gnd.n6355 gnd.n6354 19.3944
R15934 gnd.n6354 gnd.n6353 19.3944
R15935 gnd.n6353 gnd.n892 19.3944
R15936 gnd.n6349 gnd.n892 19.3944
R15937 gnd.n6349 gnd.n6348 19.3944
R15938 gnd.n6348 gnd.n6347 19.3944
R15939 gnd.n6347 gnd.n897 19.3944
R15940 gnd.n6343 gnd.n897 19.3944
R15941 gnd.n6343 gnd.n6342 19.3944
R15942 gnd.n6342 gnd.n6341 19.3944
R15943 gnd.n6341 gnd.n902 19.3944
R15944 gnd.n6337 gnd.n902 19.3944
R15945 gnd.n6337 gnd.n6336 19.3944
R15946 gnd.n6336 gnd.n6335 19.3944
R15947 gnd.n6335 gnd.n907 19.3944
R15948 gnd.n6331 gnd.n907 19.3944
R15949 gnd.n6331 gnd.n6330 19.3944
R15950 gnd.n6330 gnd.n6329 19.3944
R15951 gnd.n6329 gnd.n912 19.3944
R15952 gnd.n6325 gnd.n912 19.3944
R15953 gnd.n6325 gnd.n6324 19.3944
R15954 gnd.n6324 gnd.n6323 19.3944
R15955 gnd.n6323 gnd.n917 19.3944
R15956 gnd.n6319 gnd.n917 19.3944
R15957 gnd.n6319 gnd.n6318 19.3944
R15958 gnd.n6318 gnd.n6317 19.3944
R15959 gnd.n6317 gnd.n922 19.3944
R15960 gnd.n6313 gnd.n922 19.3944
R15961 gnd.n6313 gnd.n6312 19.3944
R15962 gnd.n6312 gnd.n6311 19.3944
R15963 gnd.n6311 gnd.n927 19.3944
R15964 gnd.n6307 gnd.n927 19.3944
R15965 gnd.n6307 gnd.n6306 19.3944
R15966 gnd.n6306 gnd.n6305 19.3944
R15967 gnd.n6305 gnd.n932 19.3944
R15968 gnd.n6301 gnd.n932 19.3944
R15969 gnd.n6301 gnd.n6300 19.3944
R15970 gnd.n6300 gnd.n6299 19.3944
R15971 gnd.n6299 gnd.n937 19.3944
R15972 gnd.n6295 gnd.n937 19.3944
R15973 gnd.n6295 gnd.n6294 19.3944
R15974 gnd.n6294 gnd.n6293 19.3944
R15975 gnd.n6293 gnd.n942 19.3944
R15976 gnd.n6289 gnd.n942 19.3944
R15977 gnd.n6289 gnd.n6288 19.3944
R15978 gnd.n6288 gnd.n6287 19.3944
R15979 gnd.n6287 gnd.n947 19.3944
R15980 gnd.n6283 gnd.n947 19.3944
R15981 gnd.n6283 gnd.n6282 19.3944
R15982 gnd.n6282 gnd.n6281 19.3944
R15983 gnd.n6281 gnd.n952 19.3944
R15984 gnd.n6277 gnd.n952 19.3944
R15985 gnd.n6277 gnd.n6276 19.3944
R15986 gnd.n6276 gnd.n6275 19.3944
R15987 gnd.n6275 gnd.n957 19.3944
R15988 gnd.n6271 gnd.n957 19.3944
R15989 gnd.n6271 gnd.n6270 19.3944
R15990 gnd.n6270 gnd.n6269 19.3944
R15991 gnd.n6269 gnd.n962 19.3944
R15992 gnd.n6265 gnd.n962 19.3944
R15993 gnd.n6265 gnd.n6264 19.3944
R15994 gnd.n6264 gnd.n6263 19.3944
R15995 gnd.n6263 gnd.n967 19.3944
R15996 gnd.n6259 gnd.n967 19.3944
R15997 gnd.n6259 gnd.n6258 19.3944
R15998 gnd.n6258 gnd.n6257 19.3944
R15999 gnd.n6257 gnd.n972 19.3944
R16000 gnd.n6253 gnd.n972 19.3944
R16001 gnd.n6253 gnd.n6252 19.3944
R16002 gnd.n6252 gnd.n6251 19.3944
R16003 gnd.n6251 gnd.n977 19.3944
R16004 gnd.n6247 gnd.n977 19.3944
R16005 gnd.n6247 gnd.n6246 19.3944
R16006 gnd.n6246 gnd.n6245 19.3944
R16007 gnd.n6245 gnd.n982 19.3944
R16008 gnd.n6241 gnd.n982 19.3944
R16009 gnd.n6241 gnd.n6240 19.3944
R16010 gnd.n6240 gnd.n6239 19.3944
R16011 gnd.n6239 gnd.n987 19.3944
R16012 gnd.n6235 gnd.n987 19.3944
R16013 gnd.n6235 gnd.n6234 19.3944
R16014 gnd.n6234 gnd.n6233 19.3944
R16015 gnd.n6233 gnd.n992 19.3944
R16016 gnd.n4947 gnd.n4946 19.3944
R16017 gnd.n4946 gnd.n2165 19.3944
R16018 gnd.n2165 gnd.n2164 19.3944
R16019 gnd.n5008 gnd.n2068 19.3944
R16020 gnd.n5003 gnd.n2068 19.3944
R16021 gnd.n5003 gnd.n2070 19.3944
R16022 gnd.n4999 gnd.n2070 19.3944
R16023 gnd.n4999 gnd.n4998 19.3944
R16024 gnd.n4998 gnd.n4997 19.3944
R16025 gnd.n4997 gnd.n4995 19.3944
R16026 gnd.n4995 gnd.n2078 19.3944
R16027 gnd.n2084 gnd.n2078 19.3944
R16028 gnd.n4987 gnd.n2084 19.3944
R16029 gnd.n4987 gnd.n4986 19.3944
R16030 gnd.n4986 gnd.n2091 19.3944
R16031 gnd.n4979 gnd.n2091 19.3944
R16032 gnd.n4979 gnd.n4978 19.3944
R16033 gnd.n4978 gnd.n2105 19.3944
R16034 gnd.n4971 gnd.n2105 19.3944
R16035 gnd.n4971 gnd.n4970 19.3944
R16036 gnd.n4970 gnd.n2117 19.3944
R16037 gnd.n4963 gnd.n2117 19.3944
R16038 gnd.n4963 gnd.n4962 19.3944
R16039 gnd.n4962 gnd.n2131 19.3944
R16040 gnd.n4955 gnd.n2131 19.3944
R16041 gnd.n4955 gnd.n4954 19.3944
R16042 gnd.n4954 gnd.n2143 19.3944
R16043 gnd.n6091 gnd.n6013 19.3944
R16044 gnd.n6091 gnd.n6090 19.3944
R16045 gnd.n6090 gnd.n6016 19.3944
R16046 gnd.n6083 gnd.n6016 19.3944
R16047 gnd.n6083 gnd.n6082 19.3944
R16048 gnd.n6082 gnd.n6026 19.3944
R16049 gnd.n6075 gnd.n6026 19.3944
R16050 gnd.n6075 gnd.n6074 19.3944
R16051 gnd.n6074 gnd.n6036 19.3944
R16052 gnd.n6067 gnd.n6036 19.3944
R16053 gnd.n6067 gnd.n6066 19.3944
R16054 gnd.n6066 gnd.n6046 19.3944
R16055 gnd.n6059 gnd.n6046 19.3944
R16056 gnd.n6059 gnd.n6058 19.3944
R16057 gnd.n6058 gnd.n1020 19.3944
R16058 gnd.n6221 gnd.n1020 19.3944
R16059 gnd.n5953 gnd.n5952 19.3944
R16060 gnd.n5961 gnd.n5953 19.3944
R16061 gnd.n5962 gnd.n5961 19.3944
R16062 gnd.n5963 gnd.n5962 19.3944
R16063 gnd.n5983 gnd.n5963 19.3944
R16064 gnd.n5983 gnd.n399 19.3944
R16065 gnd.n7040 gnd.n399 19.3944
R16066 gnd.n7041 gnd.n7040 19.3944
R16067 gnd.n7041 gnd.n371 19.3944
R16068 gnd.n7072 gnd.n371 19.3944
R16069 gnd.n7073 gnd.n7072 19.3944
R16070 gnd.n7076 gnd.n7073 19.3944
R16071 gnd.n7077 gnd.n7076 19.3944
R16072 gnd.n7077 gnd.n343 19.3944
R16073 gnd.n7128 gnd.n343 19.3944
R16074 gnd.n7129 gnd.n7128 19.3944
R16075 gnd.n7130 gnd.n7129 19.3944
R16076 gnd.n7130 gnd.n325 19.3944
R16077 gnd.n7148 gnd.n325 19.3944
R16078 gnd.n7149 gnd.n7148 19.3944
R16079 gnd.n7150 gnd.n7149 19.3944
R16080 gnd.n7150 gnd.n307 19.3944
R16081 gnd.n7168 gnd.n307 19.3944
R16082 gnd.n7169 gnd.n7168 19.3944
R16083 gnd.n7171 gnd.n7169 19.3944
R16084 gnd.n7172 gnd.n7171 19.3944
R16085 gnd.n7172 gnd.n281 19.3944
R16086 gnd.n7206 gnd.n281 19.3944
R16087 gnd.n7209 gnd.n7206 19.3944
R16088 gnd.n7209 gnd.n7208 19.3944
R16089 gnd.n7208 gnd.n262 19.3944
R16090 gnd.n7229 gnd.n262 19.3944
R16091 gnd.n7230 gnd.n7229 19.3944
R16092 gnd.n7230 gnd.n256 19.3944
R16093 gnd.n7239 gnd.n256 19.3944
R16094 gnd.n7240 gnd.n7239 19.3944
R16095 gnd.n7242 gnd.n7240 19.3944
R16096 gnd.n7243 gnd.n7242 19.3944
R16097 gnd.n7246 gnd.n7243 19.3944
R16098 gnd.n7247 gnd.n7246 19.3944
R16099 gnd.n7249 gnd.n7247 19.3944
R16100 gnd.n7250 gnd.n7249 19.3944
R16101 gnd.n7253 gnd.n7250 19.3944
R16102 gnd.n7254 gnd.n7253 19.3944
R16103 gnd.n7256 gnd.n7254 19.3944
R16104 gnd.n7257 gnd.n7256 19.3944
R16105 gnd.n7260 gnd.n7257 19.3944
R16106 gnd.n7261 gnd.n7260 19.3944
R16107 gnd.n7263 gnd.n7261 19.3944
R16108 gnd.n7264 gnd.n7263 19.3944
R16109 gnd.n7267 gnd.n7264 19.3944
R16110 gnd.n7268 gnd.n7267 19.3944
R16111 gnd.n7270 gnd.n7268 19.3944
R16112 gnd.n7271 gnd.n7270 19.3944
R16113 gnd.n7274 gnd.n7271 19.3944
R16114 gnd.n7275 gnd.n7274 19.3944
R16115 gnd.n7277 gnd.n7275 19.3944
R16116 gnd.n7278 gnd.n7277 19.3944
R16117 gnd.n7281 gnd.n7278 19.3944
R16118 gnd.n7282 gnd.n7281 19.3944
R16119 gnd.n7284 gnd.n7282 19.3944
R16120 gnd.n7285 gnd.n7284 19.3944
R16121 gnd.n7287 gnd.n7285 19.3944
R16122 gnd.n7288 gnd.n7287 19.3944
R16123 gnd.n7590 gnd.n7450 19.3944
R16124 gnd.n7594 gnd.n7450 19.3944
R16125 gnd.n7594 gnd.n7448 19.3944
R16126 gnd.n7600 gnd.n7448 19.3944
R16127 gnd.n7600 gnd.n7446 19.3944
R16128 gnd.n7604 gnd.n7446 19.3944
R16129 gnd.n7604 gnd.n7444 19.3944
R16130 gnd.n7610 gnd.n7444 19.3944
R16131 gnd.n7610 gnd.n7442 19.3944
R16132 gnd.n7614 gnd.n7442 19.3944
R16133 gnd.n7614 gnd.n7440 19.3944
R16134 gnd.n7620 gnd.n7440 19.3944
R16135 gnd.n7620 gnd.n7438 19.3944
R16136 gnd.n7624 gnd.n7438 19.3944
R16137 gnd.n7624 gnd.n7436 19.3944
R16138 gnd.n7630 gnd.n7436 19.3944
R16139 gnd.n7630 gnd.n7434 19.3944
R16140 gnd.n7634 gnd.n7434 19.3944
R16141 gnd.n7540 gnd.n7472 19.3944
R16142 gnd.n7544 gnd.n7472 19.3944
R16143 gnd.n7544 gnd.n7470 19.3944
R16144 gnd.n7550 gnd.n7470 19.3944
R16145 gnd.n7550 gnd.n7468 19.3944
R16146 gnd.n7554 gnd.n7468 19.3944
R16147 gnd.n7554 gnd.n7466 19.3944
R16148 gnd.n7560 gnd.n7466 19.3944
R16149 gnd.n7560 gnd.n7464 19.3944
R16150 gnd.n7564 gnd.n7464 19.3944
R16151 gnd.n7564 gnd.n7462 19.3944
R16152 gnd.n7570 gnd.n7462 19.3944
R16153 gnd.n7570 gnd.n7460 19.3944
R16154 gnd.n7574 gnd.n7460 19.3944
R16155 gnd.n7574 gnd.n7458 19.3944
R16156 gnd.n7580 gnd.n7458 19.3944
R16157 gnd.n7580 gnd.n7456 19.3944
R16158 gnd.n7584 gnd.n7456 19.3944
R16159 gnd.n7494 gnd.n7493 19.3944
R16160 gnd.n7499 gnd.n7494 19.3944
R16161 gnd.n7499 gnd.n7490 19.3944
R16162 gnd.n7503 gnd.n7490 19.3944
R16163 gnd.n7503 gnd.n7488 19.3944
R16164 gnd.n7509 gnd.n7488 19.3944
R16165 gnd.n7509 gnd.n7486 19.3944
R16166 gnd.n7513 gnd.n7486 19.3944
R16167 gnd.n7513 gnd.n7484 19.3944
R16168 gnd.n7519 gnd.n7484 19.3944
R16169 gnd.n7519 gnd.n7482 19.3944
R16170 gnd.n7523 gnd.n7482 19.3944
R16171 gnd.n7523 gnd.n7480 19.3944
R16172 gnd.n7530 gnd.n7480 19.3944
R16173 gnd.n7530 gnd.n7478 19.3944
R16174 gnd.n7534 gnd.n7478 19.3944
R16175 gnd.n7535 gnd.n7534 19.3944
R16176 gnd.n5994 gnd.n5992 19.3944
R16177 gnd.n5994 gnd.n5990 19.3944
R16178 gnd.n6000 gnd.n5990 19.3944
R16179 gnd.n6000 gnd.n5999 19.3944
R16180 gnd.n5999 gnd.n389 19.3944
R16181 gnd.n7053 gnd.n389 19.3944
R16182 gnd.n7053 gnd.n387 19.3944
R16183 gnd.n7059 gnd.n387 19.3944
R16184 gnd.n7059 gnd.n7058 19.3944
R16185 gnd.n7058 gnd.n360 19.3944
R16186 gnd.n7089 gnd.n360 19.3944
R16187 gnd.n7089 gnd.n358 19.3944
R16188 gnd.n7095 gnd.n358 19.3944
R16189 gnd.n7095 gnd.n7094 19.3944
R16190 gnd.n7094 gnd.n333 19.3944
R16191 gnd.n7139 gnd.n333 19.3944
R16192 gnd.n7139 gnd.n331 19.3944
R16193 gnd.n7143 gnd.n331 19.3944
R16194 gnd.n7143 gnd.n316 19.3944
R16195 gnd.n7159 gnd.n316 19.3944
R16196 gnd.n7159 gnd.n314 19.3944
R16197 gnd.n7163 gnd.n314 19.3944
R16198 gnd.n7163 gnd.n296 19.3944
R16199 gnd.n7183 gnd.n296 19.3944
R16200 gnd.n7183 gnd.n294 19.3944
R16201 gnd.n7189 gnd.n294 19.3944
R16202 gnd.n7189 gnd.n7188 19.3944
R16203 gnd.n7188 gnd.n273 19.3944
R16204 gnd.n7215 gnd.n273 19.3944
R16205 gnd.n7215 gnd.n271 19.3944
R16206 gnd.n7222 gnd.n271 19.3944
R16207 gnd.n7222 gnd.n7221 19.3944
R16208 gnd.n7221 gnd.n110 19.3944
R16209 gnd.n7733 gnd.n110 19.3944
R16210 gnd.n7733 gnd.n7732 19.3944
R16211 gnd.n7732 gnd.n7731 19.3944
R16212 gnd.n7731 gnd.n114 19.3944
R16213 gnd.n7721 gnd.n114 19.3944
R16214 gnd.n7721 gnd.n7720 19.3944
R16215 gnd.n7720 gnd.n7719 19.3944
R16216 gnd.n7719 gnd.n134 19.3944
R16217 gnd.n7709 gnd.n134 19.3944
R16218 gnd.n7709 gnd.n7708 19.3944
R16219 gnd.n7708 gnd.n7707 19.3944
R16220 gnd.n7707 gnd.n154 19.3944
R16221 gnd.n7697 gnd.n154 19.3944
R16222 gnd.n7697 gnd.n7696 19.3944
R16223 gnd.n7696 gnd.n7695 19.3944
R16224 gnd.n7695 gnd.n173 19.3944
R16225 gnd.n7685 gnd.n173 19.3944
R16226 gnd.n7685 gnd.n7684 19.3944
R16227 gnd.n7684 gnd.n7683 19.3944
R16228 gnd.n7683 gnd.n193 19.3944
R16229 gnd.n7673 gnd.n193 19.3944
R16230 gnd.n7673 gnd.n7672 19.3944
R16231 gnd.n7672 gnd.n7671 19.3944
R16232 gnd.n7671 gnd.n211 19.3944
R16233 gnd.n7661 gnd.n211 19.3944
R16234 gnd.n7661 gnd.n7660 19.3944
R16235 gnd.n7660 gnd.n7659 19.3944
R16236 gnd.n7659 gnd.n231 19.3944
R16237 gnd.n7649 gnd.n231 19.3944
R16238 gnd.n7649 gnd.n7648 19.3944
R16239 gnd.n7648 gnd.n7647 19.3944
R16240 gnd.n6212 gnd.n6211 19.3944
R16241 gnd.n6211 gnd.n6210 19.3944
R16242 gnd.n6210 gnd.n6209 19.3944
R16243 gnd.n6209 gnd.n6207 19.3944
R16244 gnd.n6207 gnd.n6204 19.3944
R16245 gnd.n6204 gnd.n6203 19.3944
R16246 gnd.n6203 gnd.n6200 19.3944
R16247 gnd.n6200 gnd.n6199 19.3944
R16248 gnd.n6199 gnd.n6196 19.3944
R16249 gnd.n6196 gnd.n6195 19.3944
R16250 gnd.n6195 gnd.n6192 19.3944
R16251 gnd.n6192 gnd.n6191 19.3944
R16252 gnd.n6191 gnd.n6188 19.3944
R16253 gnd.n6188 gnd.n6187 19.3944
R16254 gnd.n6187 gnd.n6184 19.3944
R16255 gnd.n6184 gnd.n6183 19.3944
R16256 gnd.n6183 gnd.n6180 19.3944
R16257 gnd.n6178 gnd.n6175 19.3944
R16258 gnd.n6175 gnd.n6174 19.3944
R16259 gnd.n6174 gnd.n6171 19.3944
R16260 gnd.n6171 gnd.n6170 19.3944
R16261 gnd.n6170 gnd.n6167 19.3944
R16262 gnd.n6167 gnd.n6166 19.3944
R16263 gnd.n6166 gnd.n6163 19.3944
R16264 gnd.n6161 gnd.n6158 19.3944
R16265 gnd.n6158 gnd.n6157 19.3944
R16266 gnd.n6157 gnd.n6154 19.3944
R16267 gnd.n6154 gnd.n6153 19.3944
R16268 gnd.n6153 gnd.n6150 19.3944
R16269 gnd.n6150 gnd.n6149 19.3944
R16270 gnd.n6149 gnd.n6146 19.3944
R16271 gnd.n6146 gnd.n6145 19.3944
R16272 gnd.n6141 gnd.n6138 19.3944
R16273 gnd.n6138 gnd.n6137 19.3944
R16274 gnd.n6137 gnd.n6134 19.3944
R16275 gnd.n6134 gnd.n6133 19.3944
R16276 gnd.n6133 gnd.n6130 19.3944
R16277 gnd.n6130 gnd.n6129 19.3944
R16278 gnd.n6129 gnd.n6126 19.3944
R16279 gnd.n6126 gnd.n6125 19.3944
R16280 gnd.n6125 gnd.n6122 19.3944
R16281 gnd.n6122 gnd.n6121 19.3944
R16282 gnd.n6121 gnd.n6118 19.3944
R16283 gnd.n6118 gnd.n6117 19.3944
R16284 gnd.n6117 gnd.n6114 19.3944
R16285 gnd.n6114 gnd.n6113 19.3944
R16286 gnd.n6113 gnd.n6110 19.3944
R16287 gnd.n6110 gnd.n6109 19.3944
R16288 gnd.n6109 gnd.n6106 19.3944
R16289 gnd.n6106 gnd.n6105 19.3944
R16290 gnd.n7427 gnd.n7426 19.3944
R16291 gnd.n7426 gnd.n7425 19.3944
R16292 gnd.n7425 gnd.n7292 19.3944
R16293 gnd.n7420 gnd.n7292 19.3944
R16294 gnd.n7420 gnd.n7419 19.3944
R16295 gnd.n7419 gnd.n7418 19.3944
R16296 gnd.n7418 gnd.n7299 19.3944
R16297 gnd.n7413 gnd.n7299 19.3944
R16298 gnd.n7413 gnd.n7412 19.3944
R16299 gnd.n7412 gnd.n7411 19.3944
R16300 gnd.n7411 gnd.n7306 19.3944
R16301 gnd.n7406 gnd.n7306 19.3944
R16302 gnd.n7406 gnd.n7405 19.3944
R16303 gnd.n7405 gnd.n7404 19.3944
R16304 gnd.n7404 gnd.n7313 19.3944
R16305 gnd.n7399 gnd.n7313 19.3944
R16306 gnd.n5970 gnd.n5967 19.3944
R16307 gnd.n5973 gnd.n5970 19.3944
R16308 gnd.n5974 gnd.n5973 19.3944
R16309 gnd.n5974 gnd.n5964 19.3944
R16310 gnd.n5979 gnd.n5964 19.3944
R16311 gnd.n5979 gnd.n5965 19.3944
R16312 gnd.n5965 gnd.n379 19.3944
R16313 gnd.n7063 gnd.n379 19.3944
R16314 gnd.n7063 gnd.n376 19.3944
R16315 gnd.n7068 gnd.n376 19.3944
R16316 gnd.n7068 gnd.n377 19.3944
R16317 gnd.n377 gnd.n350 19.3944
R16318 gnd.n7099 gnd.n350 19.3944
R16319 gnd.n7099 gnd.n347 19.3944
R16320 gnd.n7124 gnd.n347 19.3944
R16321 gnd.n7124 gnd.n348 19.3944
R16322 gnd.n7120 gnd.n348 19.3944
R16323 gnd.n7120 gnd.n7119 19.3944
R16324 gnd.n7119 gnd.n7118 19.3944
R16325 gnd.n7118 gnd.n7105 19.3944
R16326 gnd.n7114 gnd.n7105 19.3944
R16327 gnd.n7114 gnd.n7113 19.3944
R16328 gnd.n7113 gnd.n7112 19.3944
R16329 gnd.n7112 gnd.n7109 19.3944
R16330 gnd.n7109 gnd.n288 19.3944
R16331 gnd.n7193 gnd.n288 19.3944
R16332 gnd.n7193 gnd.n285 19.3944
R16333 gnd.n7202 gnd.n285 19.3944
R16334 gnd.n7202 gnd.n286 19.3944
R16335 gnd.n7198 gnd.n286 19.3944
R16336 gnd.n7198 gnd.n7197 19.3944
R16337 gnd.n7197 gnd.n100 19.3944
R16338 gnd.n7738 gnd.n100 19.3944
R16339 gnd.n7738 gnd.n7737 19.3944
R16340 gnd.n7737 gnd.n103 19.3944
R16341 gnd.n7345 gnd.n103 19.3944
R16342 gnd.n7345 gnd.n7343 19.3944
R16343 gnd.n7349 gnd.n7343 19.3944
R16344 gnd.n7351 gnd.n7349 19.3944
R16345 gnd.n7352 gnd.n7351 19.3944
R16346 gnd.n7352 gnd.n7340 19.3944
R16347 gnd.n7356 gnd.n7340 19.3944
R16348 gnd.n7358 gnd.n7356 19.3944
R16349 gnd.n7359 gnd.n7358 19.3944
R16350 gnd.n7359 gnd.n7337 19.3944
R16351 gnd.n7363 gnd.n7337 19.3944
R16352 gnd.n7365 gnd.n7363 19.3944
R16353 gnd.n7366 gnd.n7365 19.3944
R16354 gnd.n7366 gnd.n7334 19.3944
R16355 gnd.n7370 gnd.n7334 19.3944
R16356 gnd.n7372 gnd.n7370 19.3944
R16357 gnd.n7373 gnd.n7372 19.3944
R16358 gnd.n7373 gnd.n7331 19.3944
R16359 gnd.n7377 gnd.n7331 19.3944
R16360 gnd.n7379 gnd.n7377 19.3944
R16361 gnd.n7380 gnd.n7379 19.3944
R16362 gnd.n7380 gnd.n7328 19.3944
R16363 gnd.n7384 gnd.n7328 19.3944
R16364 gnd.n7386 gnd.n7384 19.3944
R16365 gnd.n7387 gnd.n7386 19.3944
R16366 gnd.n7387 gnd.n7325 19.3944
R16367 gnd.n7391 gnd.n7325 19.3944
R16368 gnd.n7393 gnd.n7391 19.3944
R16369 gnd.n7394 gnd.n7393 19.3944
R16370 gnd.n5955 gnd.n1150 19.3944
R16371 gnd.n5957 gnd.n5955 19.3944
R16372 gnd.n5957 gnd.n5950 19.3944
R16373 gnd.n5986 gnd.n5950 19.3944
R16374 gnd.n5986 gnd.n396 19.3944
R16375 gnd.n7049 gnd.n396 19.3944
R16376 gnd.n7049 gnd.n7048 19.3944
R16377 gnd.n7048 gnd.n7047 19.3944
R16378 gnd.n7047 gnd.n7046 19.3944
R16379 gnd.n7046 gnd.n368 19.3944
R16380 gnd.n7085 gnd.n368 19.3944
R16381 gnd.n7085 gnd.n7084 19.3944
R16382 gnd.n7084 gnd.n7083 19.3944
R16383 gnd.n7083 gnd.n7082 19.3944
R16384 gnd.n7082 gnd.n341 19.3944
R16385 gnd.n7135 gnd.n341 19.3944
R16386 gnd.n7135 gnd.n7134 19.3944
R16387 gnd.n7134 gnd.n7133 19.3944
R16388 gnd.n7133 gnd.n323 19.3944
R16389 gnd.n7155 gnd.n323 19.3944
R16390 gnd.n7155 gnd.n7154 19.3944
R16391 gnd.n7154 gnd.n7153 19.3944
R16392 gnd.n7153 gnd.n304 19.3944
R16393 gnd.n7179 gnd.n304 19.3944
R16394 gnd.n7179 gnd.n7178 19.3944
R16395 gnd.n7178 gnd.n7177 19.3944
R16396 gnd.n7177 gnd.n7176 19.3944
R16397 gnd.n7176 gnd.n279 19.3944
R16398 gnd.n7211 gnd.n279 19.3944
R16399 gnd.n7211 gnd.n264 19.3944
R16400 gnd.n7226 gnd.n264 19.3944
R16401 gnd.n7226 gnd.n258 19.3944
R16402 gnd.n7234 gnd.n258 19.3944
R16403 gnd.n7235 gnd.n7234 19.3944
R16404 gnd.n7235 gnd.n121 19.3944
R16405 gnd.n7727 gnd.n121 19.3944
R16406 gnd.n7727 gnd.n7726 19.3944
R16407 gnd.n7726 gnd.n7725 19.3944
R16408 gnd.n7725 gnd.n125 19.3944
R16409 gnd.n7715 gnd.n125 19.3944
R16410 gnd.n7715 gnd.n7714 19.3944
R16411 gnd.n7714 gnd.n7713 19.3944
R16412 gnd.n7713 gnd.n144 19.3944
R16413 gnd.n7703 gnd.n144 19.3944
R16414 gnd.n7703 gnd.n7702 19.3944
R16415 gnd.n7702 gnd.n7701 19.3944
R16416 gnd.n7701 gnd.n163 19.3944
R16417 gnd.n7691 gnd.n163 19.3944
R16418 gnd.n7691 gnd.n7690 19.3944
R16419 gnd.n7690 gnd.n7689 19.3944
R16420 gnd.n7689 gnd.n183 19.3944
R16421 gnd.n7679 gnd.n183 19.3944
R16422 gnd.n7679 gnd.n7678 19.3944
R16423 gnd.n7678 gnd.n7677 19.3944
R16424 gnd.n7677 gnd.n202 19.3944
R16425 gnd.n7667 gnd.n202 19.3944
R16426 gnd.n7667 gnd.n7666 19.3944
R16427 gnd.n7666 gnd.n7665 19.3944
R16428 gnd.n7665 gnd.n221 19.3944
R16429 gnd.n7655 gnd.n221 19.3944
R16430 gnd.n7655 gnd.n7654 19.3944
R16431 gnd.n7654 gnd.n7653 19.3944
R16432 gnd.n7653 gnd.n240 19.3944
R16433 gnd.n7643 gnd.n240 19.3944
R16434 gnd.n4991 gnd.n4990 19.3944
R16435 gnd.n4990 gnd.n2082 19.3944
R16436 gnd.n4983 gnd.n2082 19.3944
R16437 gnd.n4983 gnd.n4982 19.3944
R16438 gnd.n4982 gnd.n2098 19.3944
R16439 gnd.n4975 gnd.n2098 19.3944
R16440 gnd.n4975 gnd.n4974 19.3944
R16441 gnd.n4974 gnd.n2111 19.3944
R16442 gnd.n4967 gnd.n2111 19.3944
R16443 gnd.n4967 gnd.n4966 19.3944
R16444 gnd.n4966 gnd.n2124 19.3944
R16445 gnd.n4959 gnd.n2124 19.3944
R16446 gnd.n4959 gnd.n4958 19.3944
R16447 gnd.n4958 gnd.n2137 19.3944
R16448 gnd.n4951 gnd.n2137 19.3944
R16449 gnd.n4951 gnd.n4950 19.3944
R16450 gnd.n4867 gnd.n4570 19.3944
R16451 gnd.n4871 gnd.n4570 19.3944
R16452 gnd.n4871 gnd.n4568 19.3944
R16453 gnd.n4899 gnd.n4568 19.3944
R16454 gnd.n4899 gnd.n4898 19.3944
R16455 gnd.n4898 gnd.n4897 19.3944
R16456 gnd.n4897 gnd.n4877 19.3944
R16457 gnd.n4893 gnd.n4877 19.3944
R16458 gnd.n4893 gnd.n4892 19.3944
R16459 gnd.n4892 gnd.n4891 19.3944
R16460 gnd.n4891 gnd.n4883 19.3944
R16461 gnd.n4887 gnd.n4883 19.3944
R16462 gnd.n4887 gnd.n846 19.3944
R16463 gnd.n6397 gnd.n846 19.3944
R16464 gnd.n6397 gnd.n6396 19.3944
R16465 gnd.n6396 gnd.n6395 19.3944
R16466 gnd.n6395 gnd.n850 19.3944
R16467 gnd.n6389 gnd.n850 19.3944
R16468 gnd.n6389 gnd.n6388 19.3944
R16469 gnd.n6388 gnd.n6387 19.3944
R16470 gnd.n6387 gnd.n859 19.3944
R16471 gnd.n5017 gnd.n859 19.3944
R16472 gnd.n5021 gnd.n5017 19.3944
R16473 gnd.n5021 gnd.n2059 19.3944
R16474 gnd.n5035 gnd.n2059 19.3944
R16475 gnd.n5035 gnd.n2057 19.3944
R16476 gnd.n5039 gnd.n2057 19.3944
R16477 gnd.n5039 gnd.n2048 19.3944
R16478 gnd.n5052 gnd.n2048 19.3944
R16479 gnd.n5052 gnd.n2046 19.3944
R16480 gnd.n5056 gnd.n2046 19.3944
R16481 gnd.n5056 gnd.n2036 19.3944
R16482 gnd.n5069 gnd.n2036 19.3944
R16483 gnd.n5069 gnd.n2034 19.3944
R16484 gnd.n5075 gnd.n2034 19.3944
R16485 gnd.n5075 gnd.n5074 19.3944
R16486 gnd.n5074 gnd.n1626 19.3944
R16487 gnd.n5162 gnd.n1626 19.3944
R16488 gnd.n5162 gnd.n1624 19.3944
R16489 gnd.n5177 gnd.n1624 19.3944
R16490 gnd.n5177 gnd.n5176 19.3944
R16491 gnd.n5176 gnd.n5175 19.3944
R16492 gnd.n5175 gnd.n5168 19.3944
R16493 gnd.n5171 gnd.n5168 19.3944
R16494 gnd.n5171 gnd.n1587 19.3944
R16495 gnd.n5221 gnd.n1587 19.3944
R16496 gnd.n5221 gnd.n1585 19.3944
R16497 gnd.n5225 gnd.n1585 19.3944
R16498 gnd.n5225 gnd.n1565 19.3944
R16499 gnd.n5251 gnd.n1565 19.3944
R16500 gnd.n5251 gnd.n1563 19.3944
R16501 gnd.n5255 gnd.n1563 19.3944
R16502 gnd.n5255 gnd.n1548 19.3944
R16503 gnd.n5278 gnd.n1548 19.3944
R16504 gnd.n5278 gnd.n1546 19.3944
R16505 gnd.n5282 gnd.n1546 19.3944
R16506 gnd.n5282 gnd.n1528 19.3944
R16507 gnd.n5302 gnd.n1528 19.3944
R16508 gnd.n5302 gnd.n1526 19.3944
R16509 gnd.n5308 gnd.n1526 19.3944
R16510 gnd.n5308 gnd.n5307 19.3944
R16511 gnd.n5307 gnd.n1501 19.3944
R16512 gnd.n5360 gnd.n1501 19.3944
R16513 gnd.n5360 gnd.n1499 19.3944
R16514 gnd.n5366 gnd.n1499 19.3944
R16515 gnd.n5366 gnd.n5365 19.3944
R16516 gnd.n5365 gnd.n1479 19.3944
R16517 gnd.n5400 gnd.n1479 19.3944
R16518 gnd.n5400 gnd.n1477 19.3944
R16519 gnd.n5406 gnd.n1477 19.3944
R16520 gnd.n5406 gnd.n5405 19.3944
R16521 gnd.n5405 gnd.n1450 19.3944
R16522 gnd.n5457 gnd.n1450 19.3944
R16523 gnd.n5457 gnd.n1448 19.3944
R16524 gnd.n5463 gnd.n1448 19.3944
R16525 gnd.n5463 gnd.n5462 19.3944
R16526 gnd.n5462 gnd.n1429 19.3944
R16527 gnd.n5495 gnd.n1429 19.3944
R16528 gnd.n5495 gnd.n1427 19.3944
R16529 gnd.n5499 gnd.n1427 19.3944
R16530 gnd.n5499 gnd.n1400 19.3944
R16531 gnd.n5533 gnd.n1400 19.3944
R16532 gnd.n5533 gnd.n1398 19.3944
R16533 gnd.n5539 gnd.n1398 19.3944
R16534 gnd.n5539 gnd.n5538 19.3944
R16535 gnd.n5538 gnd.n1374 19.3944
R16536 gnd.n5577 gnd.n1374 19.3944
R16537 gnd.n5577 gnd.n1372 19.3944
R16538 gnd.n5582 gnd.n1372 19.3944
R16539 gnd.n5582 gnd.n1351 19.3944
R16540 gnd.n5618 gnd.n1351 19.3944
R16541 gnd.n5618 gnd.n5617 19.3944
R16542 gnd.n5617 gnd.n5616 19.3944
R16543 gnd.n5616 gnd.n1355 19.3944
R16544 gnd.n1358 gnd.n1355 19.3944
R16545 gnd.n1358 gnd.n1319 19.3944
R16546 gnd.n5664 gnd.n1319 19.3944
R16547 gnd.n5664 gnd.n1317 19.3944
R16548 gnd.n5668 gnd.n1317 19.3944
R16549 gnd.n5668 gnd.n1224 19.3944
R16550 gnd.n5812 gnd.n1224 19.3944
R16551 gnd.n5812 gnd.n1222 19.3944
R16552 gnd.n5816 gnd.n1222 19.3944
R16553 gnd.n5816 gnd.n1212 19.3944
R16554 gnd.n5829 gnd.n1212 19.3944
R16555 gnd.n5829 gnd.n1210 19.3944
R16556 gnd.n5833 gnd.n1210 19.3944
R16557 gnd.n5833 gnd.n1200 19.3944
R16558 gnd.n5846 gnd.n1200 19.3944
R16559 gnd.n5846 gnd.n1198 19.3944
R16560 gnd.n5850 gnd.n1198 19.3944
R16561 gnd.n5850 gnd.n1188 19.3944
R16562 gnd.n5864 gnd.n1188 19.3944
R16563 gnd.n5864 gnd.n1186 19.3944
R16564 gnd.n5868 gnd.n1186 19.3944
R16565 gnd.n5868 gnd.n1177 19.3944
R16566 gnd.n5881 gnd.n1177 19.3944
R16567 gnd.n5881 gnd.n1175 19.3944
R16568 gnd.n5887 gnd.n1175 19.3944
R16569 gnd.n5887 gnd.n5886 19.3944
R16570 gnd.n5886 gnd.n1164 19.3944
R16571 gnd.n5918 gnd.n1164 19.3944
R16572 gnd.n5918 gnd.n1162 19.3944
R16573 gnd.n5922 gnd.n1162 19.3944
R16574 gnd.n5922 gnd.n1160 19.3944
R16575 gnd.n5927 gnd.n1160 19.3944
R16576 gnd.n5927 gnd.n1158 19.3944
R16577 gnd.n6007 gnd.n1158 19.3944
R16578 gnd.n6007 gnd.n6006 19.3944
R16579 gnd.n6006 gnd.n6005 19.3944
R16580 gnd.n6005 gnd.n5933 19.3944
R16581 gnd.n5947 gnd.n5933 19.3944
R16582 gnd.n5947 gnd.n402 19.3944
R16583 gnd.n7035 gnd.n402 19.3944
R16584 gnd.n7035 gnd.n7034 19.3944
R16585 gnd.n7034 gnd.n7033 19.3944
R16586 gnd.n7033 gnd.n406 19.3944
R16587 gnd.n7029 gnd.n406 19.3944
R16588 gnd.n7029 gnd.n7028 19.3944
R16589 gnd.n7028 gnd.n7027 19.3944
R16590 gnd.n7027 gnd.n412 19.3944
R16591 gnd.n6811 gnd.n536 19.3944
R16592 gnd.n6817 gnd.n536 19.3944
R16593 gnd.n6817 gnd.n534 19.3944
R16594 gnd.n6821 gnd.n534 19.3944
R16595 gnd.n6821 gnd.n530 19.3944
R16596 gnd.n6827 gnd.n530 19.3944
R16597 gnd.n6827 gnd.n528 19.3944
R16598 gnd.n6831 gnd.n528 19.3944
R16599 gnd.n6831 gnd.n524 19.3944
R16600 gnd.n6837 gnd.n524 19.3944
R16601 gnd.n6837 gnd.n522 19.3944
R16602 gnd.n6841 gnd.n522 19.3944
R16603 gnd.n6841 gnd.n518 19.3944
R16604 gnd.n6847 gnd.n518 19.3944
R16605 gnd.n6847 gnd.n516 19.3944
R16606 gnd.n6851 gnd.n516 19.3944
R16607 gnd.n6851 gnd.n512 19.3944
R16608 gnd.n6857 gnd.n512 19.3944
R16609 gnd.n6857 gnd.n510 19.3944
R16610 gnd.n6861 gnd.n510 19.3944
R16611 gnd.n6861 gnd.n506 19.3944
R16612 gnd.n6867 gnd.n506 19.3944
R16613 gnd.n6867 gnd.n504 19.3944
R16614 gnd.n6871 gnd.n504 19.3944
R16615 gnd.n6871 gnd.n500 19.3944
R16616 gnd.n6877 gnd.n500 19.3944
R16617 gnd.n6877 gnd.n498 19.3944
R16618 gnd.n6881 gnd.n498 19.3944
R16619 gnd.n6881 gnd.n494 19.3944
R16620 gnd.n6887 gnd.n494 19.3944
R16621 gnd.n6887 gnd.n492 19.3944
R16622 gnd.n6891 gnd.n492 19.3944
R16623 gnd.n6891 gnd.n488 19.3944
R16624 gnd.n6897 gnd.n488 19.3944
R16625 gnd.n6897 gnd.n486 19.3944
R16626 gnd.n6901 gnd.n486 19.3944
R16627 gnd.n6901 gnd.n482 19.3944
R16628 gnd.n6907 gnd.n482 19.3944
R16629 gnd.n6907 gnd.n480 19.3944
R16630 gnd.n6911 gnd.n480 19.3944
R16631 gnd.n6911 gnd.n476 19.3944
R16632 gnd.n6917 gnd.n476 19.3944
R16633 gnd.n6917 gnd.n474 19.3944
R16634 gnd.n6921 gnd.n474 19.3944
R16635 gnd.n6921 gnd.n470 19.3944
R16636 gnd.n6927 gnd.n470 19.3944
R16637 gnd.n6927 gnd.n468 19.3944
R16638 gnd.n6931 gnd.n468 19.3944
R16639 gnd.n6931 gnd.n464 19.3944
R16640 gnd.n6937 gnd.n464 19.3944
R16641 gnd.n6937 gnd.n462 19.3944
R16642 gnd.n6941 gnd.n462 19.3944
R16643 gnd.n6941 gnd.n458 19.3944
R16644 gnd.n6947 gnd.n458 19.3944
R16645 gnd.n6947 gnd.n456 19.3944
R16646 gnd.n6951 gnd.n456 19.3944
R16647 gnd.n6951 gnd.n452 19.3944
R16648 gnd.n6957 gnd.n452 19.3944
R16649 gnd.n6957 gnd.n450 19.3944
R16650 gnd.n6961 gnd.n450 19.3944
R16651 gnd.n6961 gnd.n446 19.3944
R16652 gnd.n6967 gnd.n446 19.3944
R16653 gnd.n6967 gnd.n444 19.3944
R16654 gnd.n6971 gnd.n444 19.3944
R16655 gnd.n6971 gnd.n440 19.3944
R16656 gnd.n6977 gnd.n440 19.3944
R16657 gnd.n6977 gnd.n438 19.3944
R16658 gnd.n6981 gnd.n438 19.3944
R16659 gnd.n6981 gnd.n434 19.3944
R16660 gnd.n6987 gnd.n434 19.3944
R16661 gnd.n6987 gnd.n432 19.3944
R16662 gnd.n6991 gnd.n432 19.3944
R16663 gnd.n6991 gnd.n428 19.3944
R16664 gnd.n6997 gnd.n428 19.3944
R16665 gnd.n6997 gnd.n426 19.3944
R16666 gnd.n7001 gnd.n426 19.3944
R16667 gnd.n7001 gnd.n422 19.3944
R16668 gnd.n7007 gnd.n422 19.3944
R16669 gnd.n7007 gnd.n420 19.3944
R16670 gnd.n7011 gnd.n420 19.3944
R16671 gnd.n7011 gnd.n416 19.3944
R16672 gnd.n7018 gnd.n416 19.3944
R16673 gnd.n7018 gnd.n414 19.3944
R16674 gnd.n7023 gnd.n414 19.3944
R16675 gnd.n6456 gnd.n749 19.3944
R16676 gnd.n6460 gnd.n749 19.3944
R16677 gnd.n6460 gnd.n745 19.3944
R16678 gnd.n6466 gnd.n745 19.3944
R16679 gnd.n6466 gnd.n743 19.3944
R16680 gnd.n6470 gnd.n743 19.3944
R16681 gnd.n6470 gnd.n739 19.3944
R16682 gnd.n6476 gnd.n739 19.3944
R16683 gnd.n6476 gnd.n737 19.3944
R16684 gnd.n6480 gnd.n737 19.3944
R16685 gnd.n6480 gnd.n733 19.3944
R16686 gnd.n6486 gnd.n733 19.3944
R16687 gnd.n6486 gnd.n731 19.3944
R16688 gnd.n6490 gnd.n731 19.3944
R16689 gnd.n6490 gnd.n727 19.3944
R16690 gnd.n6496 gnd.n727 19.3944
R16691 gnd.n6496 gnd.n725 19.3944
R16692 gnd.n6500 gnd.n725 19.3944
R16693 gnd.n6500 gnd.n721 19.3944
R16694 gnd.n6506 gnd.n721 19.3944
R16695 gnd.n6506 gnd.n719 19.3944
R16696 gnd.n6510 gnd.n719 19.3944
R16697 gnd.n6510 gnd.n715 19.3944
R16698 gnd.n6516 gnd.n715 19.3944
R16699 gnd.n6516 gnd.n713 19.3944
R16700 gnd.n6520 gnd.n713 19.3944
R16701 gnd.n6520 gnd.n709 19.3944
R16702 gnd.n6526 gnd.n709 19.3944
R16703 gnd.n6526 gnd.n707 19.3944
R16704 gnd.n6530 gnd.n707 19.3944
R16705 gnd.n6530 gnd.n703 19.3944
R16706 gnd.n6536 gnd.n703 19.3944
R16707 gnd.n6536 gnd.n701 19.3944
R16708 gnd.n6540 gnd.n701 19.3944
R16709 gnd.n6540 gnd.n697 19.3944
R16710 gnd.n6546 gnd.n697 19.3944
R16711 gnd.n6546 gnd.n695 19.3944
R16712 gnd.n6550 gnd.n695 19.3944
R16713 gnd.n6550 gnd.n691 19.3944
R16714 gnd.n6556 gnd.n691 19.3944
R16715 gnd.n6556 gnd.n689 19.3944
R16716 gnd.n6560 gnd.n689 19.3944
R16717 gnd.n6560 gnd.n685 19.3944
R16718 gnd.n6566 gnd.n685 19.3944
R16719 gnd.n6566 gnd.n683 19.3944
R16720 gnd.n6570 gnd.n683 19.3944
R16721 gnd.n6570 gnd.n679 19.3944
R16722 gnd.n6576 gnd.n679 19.3944
R16723 gnd.n6576 gnd.n677 19.3944
R16724 gnd.n6580 gnd.n677 19.3944
R16725 gnd.n6580 gnd.n673 19.3944
R16726 gnd.n6586 gnd.n673 19.3944
R16727 gnd.n6586 gnd.n671 19.3944
R16728 gnd.n6590 gnd.n671 19.3944
R16729 gnd.n6590 gnd.n667 19.3944
R16730 gnd.n6596 gnd.n667 19.3944
R16731 gnd.n6596 gnd.n665 19.3944
R16732 gnd.n6600 gnd.n665 19.3944
R16733 gnd.n6600 gnd.n661 19.3944
R16734 gnd.n6606 gnd.n661 19.3944
R16735 gnd.n6606 gnd.n659 19.3944
R16736 gnd.n6610 gnd.n659 19.3944
R16737 gnd.n6610 gnd.n655 19.3944
R16738 gnd.n6616 gnd.n655 19.3944
R16739 gnd.n6616 gnd.n653 19.3944
R16740 gnd.n6620 gnd.n653 19.3944
R16741 gnd.n6620 gnd.n649 19.3944
R16742 gnd.n6626 gnd.n649 19.3944
R16743 gnd.n6626 gnd.n647 19.3944
R16744 gnd.n6630 gnd.n647 19.3944
R16745 gnd.n6630 gnd.n643 19.3944
R16746 gnd.n6636 gnd.n643 19.3944
R16747 gnd.n6636 gnd.n641 19.3944
R16748 gnd.n6640 gnd.n641 19.3944
R16749 gnd.n6640 gnd.n637 19.3944
R16750 gnd.n6646 gnd.n637 19.3944
R16751 gnd.n6646 gnd.n635 19.3944
R16752 gnd.n6650 gnd.n635 19.3944
R16753 gnd.n6650 gnd.n631 19.3944
R16754 gnd.n6656 gnd.n631 19.3944
R16755 gnd.n6656 gnd.n629 19.3944
R16756 gnd.n6660 gnd.n629 19.3944
R16757 gnd.n6660 gnd.n625 19.3944
R16758 gnd.n6666 gnd.n625 19.3944
R16759 gnd.n6666 gnd.n623 19.3944
R16760 gnd.n6670 gnd.n623 19.3944
R16761 gnd.n6670 gnd.n619 19.3944
R16762 gnd.n6676 gnd.n619 19.3944
R16763 gnd.n6676 gnd.n617 19.3944
R16764 gnd.n6680 gnd.n617 19.3944
R16765 gnd.n6680 gnd.n613 19.3944
R16766 gnd.n6686 gnd.n613 19.3944
R16767 gnd.n6686 gnd.n611 19.3944
R16768 gnd.n6690 gnd.n611 19.3944
R16769 gnd.n6690 gnd.n607 19.3944
R16770 gnd.n6696 gnd.n607 19.3944
R16771 gnd.n6696 gnd.n605 19.3944
R16772 gnd.n6700 gnd.n605 19.3944
R16773 gnd.n6700 gnd.n601 19.3944
R16774 gnd.n6706 gnd.n601 19.3944
R16775 gnd.n6706 gnd.n599 19.3944
R16776 gnd.n6710 gnd.n599 19.3944
R16777 gnd.n6710 gnd.n595 19.3944
R16778 gnd.n6716 gnd.n595 19.3944
R16779 gnd.n6716 gnd.n593 19.3944
R16780 gnd.n6720 gnd.n593 19.3944
R16781 gnd.n6720 gnd.n589 19.3944
R16782 gnd.n6726 gnd.n589 19.3944
R16783 gnd.n6726 gnd.n587 19.3944
R16784 gnd.n6730 gnd.n587 19.3944
R16785 gnd.n6730 gnd.n583 19.3944
R16786 gnd.n6736 gnd.n583 19.3944
R16787 gnd.n6736 gnd.n581 19.3944
R16788 gnd.n6740 gnd.n581 19.3944
R16789 gnd.n6740 gnd.n577 19.3944
R16790 gnd.n6746 gnd.n577 19.3944
R16791 gnd.n6746 gnd.n575 19.3944
R16792 gnd.n6750 gnd.n575 19.3944
R16793 gnd.n6750 gnd.n571 19.3944
R16794 gnd.n6756 gnd.n571 19.3944
R16795 gnd.n6756 gnd.n569 19.3944
R16796 gnd.n6760 gnd.n569 19.3944
R16797 gnd.n6760 gnd.n565 19.3944
R16798 gnd.n6766 gnd.n565 19.3944
R16799 gnd.n6766 gnd.n563 19.3944
R16800 gnd.n6770 gnd.n563 19.3944
R16801 gnd.n6770 gnd.n559 19.3944
R16802 gnd.n6776 gnd.n559 19.3944
R16803 gnd.n6776 gnd.n557 19.3944
R16804 gnd.n6780 gnd.n557 19.3944
R16805 gnd.n6780 gnd.n553 19.3944
R16806 gnd.n6786 gnd.n553 19.3944
R16807 gnd.n6786 gnd.n551 19.3944
R16808 gnd.n6790 gnd.n551 19.3944
R16809 gnd.n6790 gnd.n547 19.3944
R16810 gnd.n6796 gnd.n547 19.3944
R16811 gnd.n6796 gnd.n545 19.3944
R16812 gnd.n6801 gnd.n545 19.3944
R16813 gnd.n6801 gnd.n541 19.3944
R16814 gnd.n6807 gnd.n541 19.3944
R16815 gnd.n6808 gnd.n6807 19.3944
R16816 gnd.n4656 gnd.n4654 19.3944
R16817 gnd.n4656 gnd.n4653 19.3944
R16818 gnd.n4662 gnd.n4653 19.3944
R16819 gnd.n4662 gnd.n4651 19.3944
R16820 gnd.n4666 gnd.n4651 19.3944
R16821 gnd.n4666 gnd.n4649 19.3944
R16822 gnd.n4672 gnd.n4649 19.3944
R16823 gnd.n4672 gnd.n4647 19.3944
R16824 gnd.n4676 gnd.n4647 19.3944
R16825 gnd.n4676 gnd.n4645 19.3944
R16826 gnd.n4682 gnd.n4645 19.3944
R16827 gnd.n4682 gnd.n4643 19.3944
R16828 gnd.n4686 gnd.n4643 19.3944
R16829 gnd.n4686 gnd.n4641 19.3944
R16830 gnd.n4692 gnd.n4641 19.3944
R16831 gnd.n4692 gnd.n4639 19.3944
R16832 gnd.n4696 gnd.n4639 19.3944
R16833 gnd.n4696 gnd.n4637 19.3944
R16834 gnd.n4702 gnd.n4637 19.3944
R16835 gnd.n4702 gnd.n4635 19.3944
R16836 gnd.n4706 gnd.n4635 19.3944
R16837 gnd.n4706 gnd.n4633 19.3944
R16838 gnd.n4712 gnd.n4633 19.3944
R16839 gnd.n4712 gnd.n4631 19.3944
R16840 gnd.n4716 gnd.n4631 19.3944
R16841 gnd.n4716 gnd.n4629 19.3944
R16842 gnd.n4722 gnd.n4629 19.3944
R16843 gnd.n4722 gnd.n4627 19.3944
R16844 gnd.n4726 gnd.n4627 19.3944
R16845 gnd.n4726 gnd.n4625 19.3944
R16846 gnd.n4732 gnd.n4625 19.3944
R16847 gnd.n4732 gnd.n4623 19.3944
R16848 gnd.n4736 gnd.n4623 19.3944
R16849 gnd.n4736 gnd.n4621 19.3944
R16850 gnd.n4742 gnd.n4621 19.3944
R16851 gnd.n4742 gnd.n4619 19.3944
R16852 gnd.n4746 gnd.n4619 19.3944
R16853 gnd.n4746 gnd.n4617 19.3944
R16854 gnd.n4752 gnd.n4617 19.3944
R16855 gnd.n4752 gnd.n4615 19.3944
R16856 gnd.n4756 gnd.n4615 19.3944
R16857 gnd.n4756 gnd.n4613 19.3944
R16858 gnd.n4762 gnd.n4613 19.3944
R16859 gnd.n4762 gnd.n4611 19.3944
R16860 gnd.n4766 gnd.n4611 19.3944
R16861 gnd.n4766 gnd.n4609 19.3944
R16862 gnd.n4772 gnd.n4609 19.3944
R16863 gnd.n4772 gnd.n4607 19.3944
R16864 gnd.n4776 gnd.n4607 19.3944
R16865 gnd.n4776 gnd.n4605 19.3944
R16866 gnd.n4782 gnd.n4605 19.3944
R16867 gnd.n4782 gnd.n4603 19.3944
R16868 gnd.n4786 gnd.n4603 19.3944
R16869 gnd.n4786 gnd.n4601 19.3944
R16870 gnd.n4792 gnd.n4601 19.3944
R16871 gnd.n4792 gnd.n4599 19.3944
R16872 gnd.n4796 gnd.n4599 19.3944
R16873 gnd.n4796 gnd.n4597 19.3944
R16874 gnd.n4802 gnd.n4597 19.3944
R16875 gnd.n4802 gnd.n4595 19.3944
R16876 gnd.n4806 gnd.n4595 19.3944
R16877 gnd.n4806 gnd.n4593 19.3944
R16878 gnd.n4812 gnd.n4593 19.3944
R16879 gnd.n4812 gnd.n4591 19.3944
R16880 gnd.n4816 gnd.n4591 19.3944
R16881 gnd.n4816 gnd.n4589 19.3944
R16882 gnd.n4822 gnd.n4589 19.3944
R16883 gnd.n4822 gnd.n4587 19.3944
R16884 gnd.n4826 gnd.n4587 19.3944
R16885 gnd.n4826 gnd.n4585 19.3944
R16886 gnd.n4832 gnd.n4585 19.3944
R16887 gnd.n4832 gnd.n4583 19.3944
R16888 gnd.n4836 gnd.n4583 19.3944
R16889 gnd.n4836 gnd.n4581 19.3944
R16890 gnd.n4842 gnd.n4581 19.3944
R16891 gnd.n4842 gnd.n4579 19.3944
R16892 gnd.n4846 gnd.n4579 19.3944
R16893 gnd.n4846 gnd.n4577 19.3944
R16894 gnd.n4852 gnd.n4577 19.3944
R16895 gnd.n4852 gnd.n4575 19.3944
R16896 gnd.n4857 gnd.n4575 19.3944
R16897 gnd.n4857 gnd.n4573 19.3944
R16898 gnd.n4863 gnd.n4573 19.3944
R16899 gnd.n4864 gnd.n4863 19.3944
R16900 gnd.n3050 gnd.n3049 19.3944
R16901 gnd.n3049 gnd.n3048 19.3944
R16902 gnd.n3048 gnd.n3047 19.3944
R16903 gnd.n3047 gnd.n3045 19.3944
R16904 gnd.n3045 gnd.n3042 19.3944
R16905 gnd.n3042 gnd.n3041 19.3944
R16906 gnd.n3041 gnd.n3038 19.3944
R16907 gnd.n3038 gnd.n3037 19.3944
R16908 gnd.n3037 gnd.n3034 19.3944
R16909 gnd.n3034 gnd.n3033 19.3944
R16910 gnd.n3033 gnd.n3030 19.3944
R16911 gnd.n3030 gnd.n3029 19.3944
R16912 gnd.n3029 gnd.n3026 19.3944
R16913 gnd.n3026 gnd.n3025 19.3944
R16914 gnd.n3025 gnd.n3022 19.3944
R16915 gnd.n3022 gnd.n3021 19.3944
R16916 gnd.n3021 gnd.n3018 19.3944
R16917 gnd.n3018 gnd.n3017 19.3944
R16918 gnd.n3017 gnd.n3014 19.3944
R16919 gnd.n3014 gnd.n3013 19.3944
R16920 gnd.n3013 gnd.n3010 19.3944
R16921 gnd.n3010 gnd.n3009 19.3944
R16922 gnd.n3006 gnd.n3005 19.3944
R16923 gnd.n3005 gnd.n2961 19.3944
R16924 gnd.n3056 gnd.n2961 19.3944
R16925 gnd.n3822 gnd.n3821 19.3944
R16926 gnd.n3821 gnd.n3818 19.3944
R16927 gnd.n3818 gnd.n3817 19.3944
R16928 gnd.n3867 gnd.n3866 19.3944
R16929 gnd.n3866 gnd.n3865 19.3944
R16930 gnd.n3865 gnd.n3862 19.3944
R16931 gnd.n3862 gnd.n3861 19.3944
R16932 gnd.n3861 gnd.n3858 19.3944
R16933 gnd.n3858 gnd.n3857 19.3944
R16934 gnd.n3857 gnd.n3854 19.3944
R16935 gnd.n3854 gnd.n3853 19.3944
R16936 gnd.n3853 gnd.n3850 19.3944
R16937 gnd.n3850 gnd.n3849 19.3944
R16938 gnd.n3849 gnd.n3846 19.3944
R16939 gnd.n3846 gnd.n3845 19.3944
R16940 gnd.n3845 gnd.n3842 19.3944
R16941 gnd.n3842 gnd.n3841 19.3944
R16942 gnd.n3841 gnd.n3838 19.3944
R16943 gnd.n3838 gnd.n3837 19.3944
R16944 gnd.n3837 gnd.n3834 19.3944
R16945 gnd.n3834 gnd.n3833 19.3944
R16946 gnd.n3833 gnd.n3830 19.3944
R16947 gnd.n3830 gnd.n3829 19.3944
R16948 gnd.n3829 gnd.n3826 19.3944
R16949 gnd.n3826 gnd.n3825 19.3944
R16950 gnd.n3149 gnd.n2858 19.3944
R16951 gnd.n3159 gnd.n2858 19.3944
R16952 gnd.n3160 gnd.n3159 19.3944
R16953 gnd.n3160 gnd.n2839 19.3944
R16954 gnd.n3180 gnd.n2839 19.3944
R16955 gnd.n3180 gnd.n2831 19.3944
R16956 gnd.n3190 gnd.n2831 19.3944
R16957 gnd.n3191 gnd.n3190 19.3944
R16958 gnd.n3192 gnd.n3191 19.3944
R16959 gnd.n3192 gnd.n2814 19.3944
R16960 gnd.n3209 gnd.n2814 19.3944
R16961 gnd.n3212 gnd.n3209 19.3944
R16962 gnd.n3212 gnd.n3211 19.3944
R16963 gnd.n3211 gnd.n2787 19.3944
R16964 gnd.n3251 gnd.n2787 19.3944
R16965 gnd.n3251 gnd.n2784 19.3944
R16966 gnd.n3257 gnd.n2784 19.3944
R16967 gnd.n3258 gnd.n3257 19.3944
R16968 gnd.n3258 gnd.n2782 19.3944
R16969 gnd.n3264 gnd.n2782 19.3944
R16970 gnd.n3267 gnd.n3264 19.3944
R16971 gnd.n3269 gnd.n3267 19.3944
R16972 gnd.n3275 gnd.n3269 19.3944
R16973 gnd.n3275 gnd.n3274 19.3944
R16974 gnd.n3274 gnd.n2625 19.3944
R16975 gnd.n3341 gnd.n2625 19.3944
R16976 gnd.n3342 gnd.n3341 19.3944
R16977 gnd.n3342 gnd.n2618 19.3944
R16978 gnd.n3353 gnd.n2618 19.3944
R16979 gnd.n3354 gnd.n3353 19.3944
R16980 gnd.n3354 gnd.n2601 19.3944
R16981 gnd.n2601 gnd.n2599 19.3944
R16982 gnd.n3378 gnd.n2599 19.3944
R16983 gnd.n3379 gnd.n3378 19.3944
R16984 gnd.n3379 gnd.n2570 19.3944
R16985 gnd.n3426 gnd.n2570 19.3944
R16986 gnd.n3427 gnd.n3426 19.3944
R16987 gnd.n3427 gnd.n2563 19.3944
R16988 gnd.n3438 gnd.n2563 19.3944
R16989 gnd.n3439 gnd.n3438 19.3944
R16990 gnd.n3439 gnd.n2546 19.3944
R16991 gnd.n2546 gnd.n2544 19.3944
R16992 gnd.n3463 gnd.n2544 19.3944
R16993 gnd.n3464 gnd.n3463 19.3944
R16994 gnd.n3464 gnd.n2516 19.3944
R16995 gnd.n3515 gnd.n2516 19.3944
R16996 gnd.n3516 gnd.n3515 19.3944
R16997 gnd.n3516 gnd.n2509 19.3944
R16998 gnd.n3783 gnd.n2509 19.3944
R16999 gnd.n3784 gnd.n3783 19.3944
R17000 gnd.n3784 gnd.n2490 19.3944
R17001 gnd.n3809 gnd.n2490 19.3944
R17002 gnd.n3809 gnd.n2491 19.3944
R17003 gnd.n3140 gnd.n3139 19.3944
R17004 gnd.n3139 gnd.n2872 19.3944
R17005 gnd.n2895 gnd.n2872 19.3944
R17006 gnd.n2898 gnd.n2895 19.3944
R17007 gnd.n2898 gnd.n2891 19.3944
R17008 gnd.n2902 gnd.n2891 19.3944
R17009 gnd.n2905 gnd.n2902 19.3944
R17010 gnd.n2908 gnd.n2905 19.3944
R17011 gnd.n2908 gnd.n2889 19.3944
R17012 gnd.n2912 gnd.n2889 19.3944
R17013 gnd.n2915 gnd.n2912 19.3944
R17014 gnd.n2918 gnd.n2915 19.3944
R17015 gnd.n2918 gnd.n2887 19.3944
R17016 gnd.n2922 gnd.n2887 19.3944
R17017 gnd.n3145 gnd.n3144 19.3944
R17018 gnd.n3144 gnd.n2848 19.3944
R17019 gnd.n3170 gnd.n2848 19.3944
R17020 gnd.n3170 gnd.n2846 19.3944
R17021 gnd.n3176 gnd.n2846 19.3944
R17022 gnd.n3176 gnd.n3175 19.3944
R17023 gnd.n3175 gnd.n2820 19.3944
R17024 gnd.n3200 gnd.n2820 19.3944
R17025 gnd.n3200 gnd.n2818 19.3944
R17026 gnd.n3204 gnd.n2818 19.3944
R17027 gnd.n3204 gnd.n2798 19.3944
R17028 gnd.n3231 gnd.n2798 19.3944
R17029 gnd.n3231 gnd.n2796 19.3944
R17030 gnd.n3241 gnd.n2796 19.3944
R17031 gnd.n3241 gnd.n3240 19.3944
R17032 gnd.n3240 gnd.n3239 19.3944
R17033 gnd.n3239 gnd.n2745 19.3944
R17034 gnd.n3289 gnd.n2745 19.3944
R17035 gnd.n3289 gnd.n3288 19.3944
R17036 gnd.n3288 gnd.n3287 19.3944
R17037 gnd.n3287 gnd.n2749 19.3944
R17038 gnd.n2769 gnd.n2749 19.3944
R17039 gnd.n2769 gnd.n2635 19.3944
R17040 gnd.n3326 gnd.n2635 19.3944
R17041 gnd.n3326 gnd.n2633 19.3944
R17042 gnd.n3332 gnd.n2633 19.3944
R17043 gnd.n3332 gnd.n3331 19.3944
R17044 gnd.n3331 gnd.n2608 19.3944
R17045 gnd.n3366 gnd.n2608 19.3944
R17046 gnd.n3366 gnd.n2606 19.3944
R17047 gnd.n3372 gnd.n2606 19.3944
R17048 gnd.n3372 gnd.n3371 19.3944
R17049 gnd.n3371 gnd.n2581 19.3944
R17050 gnd.n3411 gnd.n2581 19.3944
R17051 gnd.n3411 gnd.n2579 19.3944
R17052 gnd.n3417 gnd.n2579 19.3944
R17053 gnd.n3417 gnd.n3416 19.3944
R17054 gnd.n3416 gnd.n2553 19.3944
R17055 gnd.n3451 gnd.n2553 19.3944
R17056 gnd.n3451 gnd.n2551 19.3944
R17057 gnd.n3457 gnd.n2551 19.3944
R17058 gnd.n3457 gnd.n3456 19.3944
R17059 gnd.n3456 gnd.n2526 19.3944
R17060 gnd.n3500 gnd.n2526 19.3944
R17061 gnd.n3500 gnd.n2524 19.3944
R17062 gnd.n3506 gnd.n2524 19.3944
R17063 gnd.n3506 gnd.n3505 19.3944
R17064 gnd.n3505 gnd.n2499 19.3944
R17065 gnd.n3794 gnd.n2499 19.3944
R17066 gnd.n3794 gnd.n2497 19.3944
R17067 gnd.n3802 gnd.n2497 19.3944
R17068 gnd.n3802 gnd.n3801 19.3944
R17069 gnd.n3801 gnd.n3800 19.3944
R17070 gnd.n3903 gnd.n3902 19.3944
R17071 gnd.n3902 gnd.n2438 19.3944
R17072 gnd.n3898 gnd.n2438 19.3944
R17073 gnd.n3898 gnd.n3895 19.3944
R17074 gnd.n3895 gnd.n3892 19.3944
R17075 gnd.n3892 gnd.n3891 19.3944
R17076 gnd.n3891 gnd.n3888 19.3944
R17077 gnd.n3888 gnd.n3887 19.3944
R17078 gnd.n3887 gnd.n3884 19.3944
R17079 gnd.n3884 gnd.n3883 19.3944
R17080 gnd.n3883 gnd.n3880 19.3944
R17081 gnd.n3880 gnd.n3879 19.3944
R17082 gnd.n3879 gnd.n3876 19.3944
R17083 gnd.n3876 gnd.n3875 19.3944
R17084 gnd.n3060 gnd.n2959 19.3944
R17085 gnd.n3060 gnd.n2950 19.3944
R17086 gnd.n3073 gnd.n2950 19.3944
R17087 gnd.n3073 gnd.n2948 19.3944
R17088 gnd.n3077 gnd.n2948 19.3944
R17089 gnd.n3077 gnd.n2938 19.3944
R17090 gnd.n3089 gnd.n2938 19.3944
R17091 gnd.n3089 gnd.n2936 19.3944
R17092 gnd.n3123 gnd.n2936 19.3944
R17093 gnd.n3123 gnd.n3122 19.3944
R17094 gnd.n3122 gnd.n3121 19.3944
R17095 gnd.n3121 gnd.n3120 19.3944
R17096 gnd.n3120 gnd.n3117 19.3944
R17097 gnd.n3117 gnd.n3116 19.3944
R17098 gnd.n3116 gnd.n3115 19.3944
R17099 gnd.n3115 gnd.n3113 19.3944
R17100 gnd.n3113 gnd.n3112 19.3944
R17101 gnd.n3112 gnd.n3109 19.3944
R17102 gnd.n3109 gnd.n3108 19.3944
R17103 gnd.n3108 gnd.n3107 19.3944
R17104 gnd.n3107 gnd.n3105 19.3944
R17105 gnd.n3105 gnd.n2804 19.3944
R17106 gnd.n3220 gnd.n2804 19.3944
R17107 gnd.n3220 gnd.n2802 19.3944
R17108 gnd.n3226 gnd.n2802 19.3944
R17109 gnd.n3226 gnd.n3225 19.3944
R17110 gnd.n3225 gnd.n2726 19.3944
R17111 gnd.n3300 gnd.n2726 19.3944
R17112 gnd.n3300 gnd.n2727 19.3944
R17113 gnd.n2774 gnd.n2773 19.3944
R17114 gnd.n2777 gnd.n2776 19.3944
R17115 gnd.n2764 gnd.n2763 19.3944
R17116 gnd.n3319 gnd.n2640 19.3944
R17117 gnd.n3319 gnd.n3318 19.3944
R17118 gnd.n3318 gnd.n3317 19.3944
R17119 gnd.n3317 gnd.n3315 19.3944
R17120 gnd.n3315 gnd.n3314 19.3944
R17121 gnd.n3314 gnd.n3312 19.3944
R17122 gnd.n3312 gnd.n3311 19.3944
R17123 gnd.n3311 gnd.n2589 19.3944
R17124 gnd.n3387 gnd.n2589 19.3944
R17125 gnd.n3387 gnd.n2587 19.3944
R17126 gnd.n3406 gnd.n2587 19.3944
R17127 gnd.n3406 gnd.n3405 19.3944
R17128 gnd.n3405 gnd.n3404 19.3944
R17129 gnd.n3404 gnd.n3402 19.3944
R17130 gnd.n3402 gnd.n3401 19.3944
R17131 gnd.n3401 gnd.n3399 19.3944
R17132 gnd.n3399 gnd.n3398 19.3944
R17133 gnd.n3398 gnd.n2533 19.3944
R17134 gnd.n3472 gnd.n2533 19.3944
R17135 gnd.n3472 gnd.n2531 19.3944
R17136 gnd.n3495 gnd.n2531 19.3944
R17137 gnd.n3495 gnd.n3494 19.3944
R17138 gnd.n3494 gnd.n3493 19.3944
R17139 gnd.n3493 gnd.n3490 19.3944
R17140 gnd.n3490 gnd.n3489 19.3944
R17141 gnd.n3489 gnd.n3487 19.3944
R17142 gnd.n3487 gnd.n3486 19.3944
R17143 gnd.n3486 gnd.n3484 19.3944
R17144 gnd.n3484 gnd.n2485 19.3944
R17145 gnd.n3065 gnd.n2955 19.3944
R17146 gnd.n3065 gnd.n2953 19.3944
R17147 gnd.n3069 gnd.n2953 19.3944
R17148 gnd.n3069 gnd.n2944 19.3944
R17149 gnd.n3081 gnd.n2944 19.3944
R17150 gnd.n3081 gnd.n2942 19.3944
R17151 gnd.n3085 gnd.n2942 19.3944
R17152 gnd.n3085 gnd.n2931 19.3944
R17153 gnd.n3127 gnd.n2931 19.3944
R17154 gnd.n3127 gnd.n2885 19.3944
R17155 gnd.n3133 gnd.n2885 19.3944
R17156 gnd.n3133 gnd.n3132 19.3944
R17157 gnd.n3132 gnd.n2863 19.3944
R17158 gnd.n3154 gnd.n2863 19.3944
R17159 gnd.n3154 gnd.n2856 19.3944
R17160 gnd.n3165 gnd.n2856 19.3944
R17161 gnd.n3165 gnd.n3164 19.3944
R17162 gnd.n3164 gnd.n2837 19.3944
R17163 gnd.n3185 gnd.n2837 19.3944
R17164 gnd.n3185 gnd.n2827 19.3944
R17165 gnd.n3195 gnd.n2827 19.3944
R17166 gnd.n3195 gnd.n2810 19.3944
R17167 gnd.n3216 gnd.n2810 19.3944
R17168 gnd.n3216 gnd.n3215 19.3944
R17169 gnd.n3215 gnd.n2789 19.3944
R17170 gnd.n3246 gnd.n2789 19.3944
R17171 gnd.n3246 gnd.n2734 19.3944
R17172 gnd.n3296 gnd.n2734 19.3944
R17173 gnd.n3296 gnd.n3295 19.3944
R17174 gnd.n3295 gnd.n3294 19.3944
R17175 gnd.n3294 gnd.n2738 19.3944
R17176 gnd.n2756 gnd.n2738 19.3944
R17177 gnd.n3282 gnd.n2756 19.3944
R17178 gnd.n3282 gnd.n3281 19.3944
R17179 gnd.n3281 gnd.n3280 19.3944
R17180 gnd.n3280 gnd.n2760 19.3944
R17181 gnd.n2760 gnd.n2627 19.3944
R17182 gnd.n3337 gnd.n2627 19.3944
R17183 gnd.n3337 gnd.n2620 19.3944
R17184 gnd.n3348 gnd.n2620 19.3944
R17185 gnd.n3348 gnd.n2616 19.3944
R17186 gnd.n3361 gnd.n2616 19.3944
R17187 gnd.n3361 gnd.n3360 19.3944
R17188 gnd.n3360 gnd.n2595 19.3944
R17189 gnd.n3383 gnd.n2595 19.3944
R17190 gnd.n3383 gnd.n3382 19.3944
R17191 gnd.n3382 gnd.n2572 19.3944
R17192 gnd.n3422 gnd.n2572 19.3944
R17193 gnd.n3422 gnd.n2565 19.3944
R17194 gnd.n3433 gnd.n2565 19.3944
R17195 gnd.n3433 gnd.n2561 19.3944
R17196 gnd.n3446 gnd.n2561 19.3944
R17197 gnd.n3446 gnd.n3445 19.3944
R17198 gnd.n3445 gnd.n2540 19.3944
R17199 gnd.n3468 gnd.n2540 19.3944
R17200 gnd.n3468 gnd.n3467 19.3944
R17201 gnd.n3467 gnd.n2518 19.3944
R17202 gnd.n3511 gnd.n2518 19.3944
R17203 gnd.n3511 gnd.n2511 19.3944
R17204 gnd.n3522 gnd.n2511 19.3944
R17205 gnd.n3522 gnd.n2507 19.3944
R17206 gnd.n3789 gnd.n2507 19.3944
R17207 gnd.n3789 gnd.n3788 19.3944
R17208 gnd.n3788 gnd.n2488 19.3944
R17209 gnd.n3812 gnd.n2488 19.3944
R17210 gnd.n4255 gnd.n4254 19.3944
R17211 gnd.n4255 gnd.n2403 19.3944
R17212 gnd.n4273 gnd.n2403 19.3944
R17213 gnd.n4274 gnd.n4273 19.3944
R17214 gnd.n4275 gnd.n4274 19.3944
R17215 gnd.n4275 gnd.n2385 19.3944
R17216 gnd.n4293 gnd.n2385 19.3944
R17217 gnd.n4294 gnd.n4293 19.3944
R17218 gnd.n4295 gnd.n4294 19.3944
R17219 gnd.n4295 gnd.n2367 19.3944
R17220 gnd.n4313 gnd.n2367 19.3944
R17221 gnd.n4314 gnd.n4313 19.3944
R17222 gnd.n4315 gnd.n4314 19.3944
R17223 gnd.n4315 gnd.n2349 19.3944
R17224 gnd.n4333 gnd.n2349 19.3944
R17225 gnd.n4334 gnd.n4333 19.3944
R17226 gnd.n4335 gnd.n4334 19.3944
R17227 gnd.n4335 gnd.n2331 19.3944
R17228 gnd.n4353 gnd.n2331 19.3944
R17229 gnd.n4354 gnd.n4353 19.3944
R17230 gnd.n4355 gnd.n4354 19.3944
R17231 gnd.n4355 gnd.n2313 19.3944
R17232 gnd.n4373 gnd.n2313 19.3944
R17233 gnd.n4374 gnd.n4373 19.3944
R17234 gnd.n4376 gnd.n4374 19.3944
R17235 gnd.n4377 gnd.n4376 19.3944
R17236 gnd.n4377 gnd.n2287 19.3944
R17237 gnd.n4408 gnd.n2287 19.3944
R17238 gnd.n4409 gnd.n4408 19.3944
R17239 gnd.n4411 gnd.n4409 19.3944
R17240 gnd.n4412 gnd.n4411 19.3944
R17241 gnd.n4412 gnd.n2261 19.3944
R17242 gnd.n4442 gnd.n2261 19.3944
R17243 gnd.n4443 gnd.n4442 19.3944
R17244 gnd.n4445 gnd.n4443 19.3944
R17245 gnd.n4446 gnd.n4445 19.3944
R17246 gnd.n4446 gnd.n2235 19.3944
R17247 gnd.n4476 gnd.n2235 19.3944
R17248 gnd.n4477 gnd.n4476 19.3944
R17249 gnd.n4479 gnd.n4477 19.3944
R17250 gnd.n4480 gnd.n4479 19.3944
R17251 gnd.n4480 gnd.n2209 19.3944
R17252 gnd.n4510 gnd.n2209 19.3944
R17253 gnd.n4511 gnd.n4510 19.3944
R17254 gnd.n4513 gnd.n4511 19.3944
R17255 gnd.n4514 gnd.n4513 19.3944
R17256 gnd.n4517 gnd.n4514 19.3944
R17257 gnd.n4517 gnd.n4515 19.3944
R17258 gnd.n4515 gnd.n2181 19.3944
R17259 gnd.n4554 gnd.n2181 19.3944
R17260 gnd.n4555 gnd.n4554 19.3944
R17261 gnd.n4556 gnd.n4555 19.3944
R17262 gnd.n4556 gnd.n2176 19.3944
R17263 gnd.n4904 gnd.n2176 19.3944
R17264 gnd.n4905 gnd.n4904 19.3944
R17265 gnd.n4906 gnd.n4905 19.3944
R17266 gnd.n4906 gnd.n2171 19.3944
R17267 gnd.n4918 gnd.n2171 19.3944
R17268 gnd.n4919 gnd.n4918 19.3944
R17269 gnd.n4926 gnd.n4919 19.3944
R17270 gnd.n4926 gnd.n4925 19.3944
R17271 gnd.n4925 gnd.n4924 19.3944
R17272 gnd.n4924 gnd.n4921 19.3944
R17273 gnd.n4921 gnd.n835 19.3944
R17274 gnd.n4250 gnd.n4249 19.3944
R17275 gnd.n4249 gnd.n4124 19.3944
R17276 gnd.n4243 gnd.n4124 19.3944
R17277 gnd.n4243 gnd.n4242 19.3944
R17278 gnd.n4242 gnd.n4241 19.3944
R17279 gnd.n4241 gnd.n4130 19.3944
R17280 gnd.n4235 gnd.n4130 19.3944
R17281 gnd.n4235 gnd.n4234 19.3944
R17282 gnd.n4234 gnd.n4233 19.3944
R17283 gnd.n4233 gnd.n4136 19.3944
R17284 gnd.n4227 gnd.n4136 19.3944
R17285 gnd.n4227 gnd.n4226 19.3944
R17286 gnd.n4226 gnd.n4225 19.3944
R17287 gnd.n4225 gnd.n4142 19.3944
R17288 gnd.n4219 gnd.n4142 19.3944
R17289 gnd.n4219 gnd.n4218 19.3944
R17290 gnd.n4209 gnd.n4208 19.3944
R17291 gnd.n4208 gnd.n4206 19.3944
R17292 gnd.n4206 gnd.n4205 19.3944
R17293 gnd.n4205 gnd.n4203 19.3944
R17294 gnd.n4203 gnd.n4202 19.3944
R17295 gnd.n4202 gnd.n4200 19.3944
R17296 gnd.n4200 gnd.n4199 19.3944
R17297 gnd.n4199 gnd.n4197 19.3944
R17298 gnd.n4197 gnd.n4196 19.3944
R17299 gnd.n4196 gnd.n4194 19.3944
R17300 gnd.n4194 gnd.n4193 19.3944
R17301 gnd.n4193 gnd.n4191 19.3944
R17302 gnd.n4191 gnd.n4190 19.3944
R17303 gnd.n4190 gnd.n4188 19.3944
R17304 gnd.n4188 gnd.n4187 19.3944
R17305 gnd.n4187 gnd.n4185 19.3944
R17306 gnd.n4185 gnd.n4184 19.3944
R17307 gnd.n4184 gnd.n4182 19.3944
R17308 gnd.n4182 gnd.n4181 19.3944
R17309 gnd.n4181 gnd.n4179 19.3944
R17310 gnd.n4179 gnd.n4178 19.3944
R17311 gnd.n4178 gnd.n4176 19.3944
R17312 gnd.n4176 gnd.n4175 19.3944
R17313 gnd.n4175 gnd.n4173 19.3944
R17314 gnd.n4173 gnd.n2294 19.3944
R17315 gnd.n4398 gnd.n2294 19.3944
R17316 gnd.n4398 gnd.n2292 19.3944
R17317 gnd.n4404 gnd.n2292 19.3944
R17318 gnd.n4404 gnd.n4403 19.3944
R17319 gnd.n4403 gnd.n2269 19.3944
R17320 gnd.n4433 gnd.n2269 19.3944
R17321 gnd.n4433 gnd.n2266 19.3944
R17322 gnd.n4438 gnd.n2266 19.3944
R17323 gnd.n4438 gnd.n2267 19.3944
R17324 gnd.n2267 gnd.n2243 19.3944
R17325 gnd.n4467 gnd.n2243 19.3944
R17326 gnd.n4467 gnd.n2240 19.3944
R17327 gnd.n4472 gnd.n2240 19.3944
R17328 gnd.n4472 gnd.n2241 19.3944
R17329 gnd.n2241 gnd.n2217 19.3944
R17330 gnd.n4501 gnd.n2217 19.3944
R17331 gnd.n4501 gnd.n2214 19.3944
R17332 gnd.n4506 gnd.n2214 19.3944
R17333 gnd.n4506 gnd.n2215 19.3944
R17334 gnd.n2215 gnd.n2191 19.3944
R17335 gnd.n4537 gnd.n2191 19.3944
R17336 gnd.n4537 gnd.n2188 19.3944
R17337 gnd.n4545 gnd.n2188 19.3944
R17338 gnd.n4545 gnd.n2189 19.3944
R17339 gnd.n4541 gnd.n2189 19.3944
R17340 gnd.n4541 gnd.n2180 19.3944
R17341 gnd.n4560 gnd.n2180 19.3944
R17342 gnd.n4560 gnd.n2178 19.3944
R17343 gnd.n4564 gnd.n2178 19.3944
R17344 gnd.n4564 gnd.n2175 19.3944
R17345 gnd.n4910 gnd.n2175 19.3944
R17346 gnd.n4910 gnd.n2173 19.3944
R17347 gnd.n4914 gnd.n2173 19.3944
R17348 gnd.n4914 gnd.n2170 19.3944
R17349 gnd.n4930 gnd.n2170 19.3944
R17350 gnd.n4930 gnd.n2167 19.3944
R17351 gnd.n4934 gnd.n2167 19.3944
R17352 gnd.n4935 gnd.n4934 19.3944
R17353 gnd.n4936 gnd.n4935 19.3944
R17354 gnd.n3977 gnd.n3974 19.3944
R17355 gnd.n3977 gnd.n3973 19.3944
R17356 gnd.n3981 gnd.n3973 19.3944
R17357 gnd.n3981 gnd.n3971 19.3944
R17358 gnd.n3987 gnd.n3971 19.3944
R17359 gnd.n3987 gnd.n3969 19.3944
R17360 gnd.n3991 gnd.n3969 19.3944
R17361 gnd.n3991 gnd.n3967 19.3944
R17362 gnd.n3997 gnd.n3967 19.3944
R17363 gnd.n3997 gnd.n3965 19.3944
R17364 gnd.n4001 gnd.n3965 19.3944
R17365 gnd.n4001 gnd.n3963 19.3944
R17366 gnd.n4007 gnd.n3963 19.3944
R17367 gnd.n4007 gnd.n3961 19.3944
R17368 gnd.n4011 gnd.n3961 19.3944
R17369 gnd.n4011 gnd.n3956 19.3944
R17370 gnd.n4017 gnd.n3956 19.3944
R17371 gnd.n4021 gnd.n3954 19.3944
R17372 gnd.n4021 gnd.n3952 19.3944
R17373 gnd.n4027 gnd.n3952 19.3944
R17374 gnd.n4027 gnd.n3950 19.3944
R17375 gnd.n4031 gnd.n3950 19.3944
R17376 gnd.n4031 gnd.n3948 19.3944
R17377 gnd.n4037 gnd.n3948 19.3944
R17378 gnd.n4037 gnd.n3946 19.3944
R17379 gnd.n4041 gnd.n3946 19.3944
R17380 gnd.n4041 gnd.n3944 19.3944
R17381 gnd.n4047 gnd.n3944 19.3944
R17382 gnd.n4047 gnd.n3942 19.3944
R17383 gnd.n4051 gnd.n3942 19.3944
R17384 gnd.n4051 gnd.n3940 19.3944
R17385 gnd.n4057 gnd.n3940 19.3944
R17386 gnd.n4057 gnd.n3938 19.3944
R17387 gnd.n4061 gnd.n3938 19.3944
R17388 gnd.n4061 gnd.n3936 19.3944
R17389 gnd.n4073 gnd.n3934 19.3944
R17390 gnd.n4073 gnd.n3932 19.3944
R17391 gnd.n4079 gnd.n3932 19.3944
R17392 gnd.n4079 gnd.n3930 19.3944
R17393 gnd.n4083 gnd.n3930 19.3944
R17394 gnd.n4083 gnd.n3928 19.3944
R17395 gnd.n4089 gnd.n3928 19.3944
R17396 gnd.n4089 gnd.n3926 19.3944
R17397 gnd.n4093 gnd.n3926 19.3944
R17398 gnd.n4093 gnd.n3924 19.3944
R17399 gnd.n4099 gnd.n3924 19.3944
R17400 gnd.n4099 gnd.n3922 19.3944
R17401 gnd.n4103 gnd.n3922 19.3944
R17402 gnd.n4103 gnd.n3920 19.3944
R17403 gnd.n4109 gnd.n3920 19.3944
R17404 gnd.n4109 gnd.n3918 19.3944
R17405 gnd.n4114 gnd.n3918 19.3944
R17406 gnd.n4114 gnd.n3916 19.3944
R17407 gnd.n1785 gnd.n1781 19.3944
R17408 gnd.n1785 gnd.n1778 19.3944
R17409 gnd.n1789 gnd.n1778 19.3944
R17410 gnd.n1789 gnd.n1776 19.3944
R17411 gnd.n1795 gnd.n1776 19.3944
R17412 gnd.n1795 gnd.n1774 19.3944
R17413 gnd.n1799 gnd.n1774 19.3944
R17414 gnd.n1799 gnd.n1772 19.3944
R17415 gnd.n1805 gnd.n1772 19.3944
R17416 gnd.n1805 gnd.n1770 19.3944
R17417 gnd.n1809 gnd.n1770 19.3944
R17418 gnd.n1809 gnd.n1768 19.3944
R17419 gnd.n1815 gnd.n1768 19.3944
R17420 gnd.n1815 gnd.n1766 19.3944
R17421 gnd.n1819 gnd.n1766 19.3944
R17422 gnd.n1819 gnd.n1764 19.3944
R17423 gnd.n1824 gnd.n1764 19.3944
R17424 gnd.n1929 gnd.n1862 19.3944
R17425 gnd.n1929 gnd.n1866 19.3944
R17426 gnd.n1869 gnd.n1866 19.3944
R17427 gnd.n1922 gnd.n1869 19.3944
R17428 gnd.n1922 gnd.n1921 19.3944
R17429 gnd.n1921 gnd.n1920 19.3944
R17430 gnd.n1920 gnd.n1875 19.3944
R17431 gnd.n1915 gnd.n1875 19.3944
R17432 gnd.n1915 gnd.n1914 19.3944
R17433 gnd.n1914 gnd.n1913 19.3944
R17434 gnd.n1913 gnd.n1882 19.3944
R17435 gnd.n1908 gnd.n1882 19.3944
R17436 gnd.n1908 gnd.n1907 19.3944
R17437 gnd.n1907 gnd.n1906 19.3944
R17438 gnd.n1906 gnd.n1889 19.3944
R17439 gnd.n1901 gnd.n1889 19.3944
R17440 gnd.n1901 gnd.n1900 19.3944
R17441 gnd.n1900 gnd.n1899 19.3944
R17442 gnd.n1948 gnd.n1750 19.3944
R17443 gnd.n1948 gnd.n1848 19.3944
R17444 gnd.n1851 gnd.n1848 19.3944
R17445 gnd.n1941 gnd.n1851 19.3944
R17446 gnd.n1941 gnd.n1940 19.3944
R17447 gnd.n1940 gnd.n1939 19.3944
R17448 gnd.n1939 gnd.n1857 19.3944
R17449 gnd.n1934 gnd.n1857 19.3944
R17450 gnd.n1827 gnd.n1758 19.3944
R17451 gnd.n1833 gnd.n1758 19.3944
R17452 gnd.n1833 gnd.n1756 19.3944
R17453 gnd.n1837 gnd.n1756 19.3944
R17454 gnd.n1837 gnd.n1754 19.3944
R17455 gnd.n1844 gnd.n1754 19.3944
R17456 gnd.n1844 gnd.n1751 19.3944
R17457 gnd.n4264 gnd.n2409 19.3944
R17458 gnd.n4268 gnd.n2409 19.3944
R17459 gnd.n4268 gnd.n2394 19.3944
R17460 gnd.n4284 gnd.n2394 19.3944
R17461 gnd.n4284 gnd.n2392 19.3944
R17462 gnd.n4288 gnd.n2392 19.3944
R17463 gnd.n4288 gnd.n2375 19.3944
R17464 gnd.n4304 gnd.n2375 19.3944
R17465 gnd.n4304 gnd.n2373 19.3944
R17466 gnd.n4308 gnd.n2373 19.3944
R17467 gnd.n4308 gnd.n2358 19.3944
R17468 gnd.n4324 gnd.n2358 19.3944
R17469 gnd.n4324 gnd.n2356 19.3944
R17470 gnd.n4328 gnd.n2356 19.3944
R17471 gnd.n4328 gnd.n2339 19.3944
R17472 gnd.n4344 gnd.n2339 19.3944
R17473 gnd.n4344 gnd.n2337 19.3944
R17474 gnd.n4348 gnd.n2337 19.3944
R17475 gnd.n4348 gnd.n2322 19.3944
R17476 gnd.n4364 gnd.n2322 19.3944
R17477 gnd.n4364 gnd.n2320 19.3944
R17478 gnd.n4368 gnd.n2320 19.3944
R17479 gnd.n4368 gnd.n2302 19.3944
R17480 gnd.n4388 gnd.n2302 19.3944
R17481 gnd.n4388 gnd.n2300 19.3944
R17482 gnd.n4394 gnd.n2300 19.3944
R17483 gnd.n4394 gnd.n4393 19.3944
R17484 gnd.n4393 gnd.n2277 19.3944
R17485 gnd.n4423 gnd.n2277 19.3944
R17486 gnd.n4423 gnd.n2275 19.3944
R17487 gnd.n4429 gnd.n2275 19.3944
R17488 gnd.n4429 gnd.n4428 19.3944
R17489 gnd.n4428 gnd.n2251 19.3944
R17490 gnd.n4457 gnd.n2251 19.3944
R17491 gnd.n4457 gnd.n2249 19.3944
R17492 gnd.n4463 gnd.n2249 19.3944
R17493 gnd.n4463 gnd.n4462 19.3944
R17494 gnd.n4462 gnd.n2226 19.3944
R17495 gnd.n4491 gnd.n2226 19.3944
R17496 gnd.n4491 gnd.n2224 19.3944
R17497 gnd.n4497 gnd.n2224 19.3944
R17498 gnd.n4497 gnd.n4496 19.3944
R17499 gnd.n4496 gnd.n2200 19.3944
R17500 gnd.n4526 gnd.n2200 19.3944
R17501 gnd.n4526 gnd.n2198 19.3944
R17502 gnd.n4533 gnd.n2198 19.3944
R17503 gnd.n4533 gnd.n4532 19.3944
R17504 gnd.n4532 gnd.n759 19.3944
R17505 gnd.n6450 gnd.n759 19.3944
R17506 gnd.n6450 gnd.n6449 19.3944
R17507 gnd.n6449 gnd.n6448 19.3944
R17508 gnd.n6448 gnd.n763 19.3944
R17509 gnd.n6438 gnd.n763 19.3944
R17510 gnd.n6438 gnd.n6437 19.3944
R17511 gnd.n6437 gnd.n6436 19.3944
R17512 gnd.n6436 gnd.n786 19.3944
R17513 gnd.n6426 gnd.n786 19.3944
R17514 gnd.n6426 gnd.n6425 19.3944
R17515 gnd.n6425 gnd.n6424 19.3944
R17516 gnd.n6424 gnd.n806 19.3944
R17517 gnd.n6414 gnd.n806 19.3944
R17518 gnd.n6414 gnd.n6413 19.3944
R17519 gnd.n6413 gnd.n6412 19.3944
R17520 gnd.n6412 gnd.n827 19.3944
R17521 gnd.n4260 gnd.n4259 19.3944
R17522 gnd.n4259 gnd.n4258 19.3944
R17523 gnd.n4258 gnd.n2401 19.3944
R17524 gnd.n4280 gnd.n2401 19.3944
R17525 gnd.n4280 gnd.n4279 19.3944
R17526 gnd.n4279 gnd.n4278 19.3944
R17527 gnd.n4278 gnd.n2383 19.3944
R17528 gnd.n4300 gnd.n2383 19.3944
R17529 gnd.n4300 gnd.n4299 19.3944
R17530 gnd.n4299 gnd.n4298 19.3944
R17531 gnd.n4298 gnd.n2365 19.3944
R17532 gnd.n4320 gnd.n2365 19.3944
R17533 gnd.n4320 gnd.n4319 19.3944
R17534 gnd.n4319 gnd.n4318 19.3944
R17535 gnd.n4318 gnd.n2347 19.3944
R17536 gnd.n4340 gnd.n2347 19.3944
R17537 gnd.n4340 gnd.n4339 19.3944
R17538 gnd.n4339 gnd.n4338 19.3944
R17539 gnd.n4338 gnd.n2329 19.3944
R17540 gnd.n4360 gnd.n2329 19.3944
R17541 gnd.n4360 gnd.n4359 19.3944
R17542 gnd.n4359 gnd.n4358 19.3944
R17543 gnd.n4358 gnd.n2310 19.3944
R17544 gnd.n4384 gnd.n2310 19.3944
R17545 gnd.n4384 gnd.n4383 19.3944
R17546 gnd.n4383 gnd.n4382 19.3944
R17547 gnd.n4382 gnd.n4381 19.3944
R17548 gnd.n4381 gnd.n2284 19.3944
R17549 gnd.n4419 gnd.n2284 19.3944
R17550 gnd.n4419 gnd.n4418 19.3944
R17551 gnd.n4418 gnd.n4417 19.3944
R17552 gnd.n4417 gnd.n4416 19.3944
R17553 gnd.n4416 gnd.n2258 19.3944
R17554 gnd.n4453 gnd.n2258 19.3944
R17555 gnd.n4453 gnd.n4452 19.3944
R17556 gnd.n4452 gnd.n4451 19.3944
R17557 gnd.n4451 gnd.n4450 19.3944
R17558 gnd.n4450 gnd.n2232 19.3944
R17559 gnd.n4487 gnd.n2232 19.3944
R17560 gnd.n4487 gnd.n4486 19.3944
R17561 gnd.n4486 gnd.n4485 19.3944
R17562 gnd.n4485 gnd.n4484 19.3944
R17563 gnd.n4484 gnd.n2206 19.3944
R17564 gnd.n4522 gnd.n2206 19.3944
R17565 gnd.n4522 gnd.n4521 19.3944
R17566 gnd.n4521 gnd.n4520 19.3944
R17567 gnd.n4520 gnd.n2183 19.3944
R17568 gnd.n4549 gnd.n2183 19.3944
R17569 gnd.n4550 gnd.n4549 19.3944
R17570 gnd.n4550 gnd.n771 19.3944
R17571 gnd.n6444 gnd.n771 19.3944
R17572 gnd.n6444 gnd.n6443 19.3944
R17573 gnd.n6443 gnd.n6442 19.3944
R17574 gnd.n6442 gnd.n775 19.3944
R17575 gnd.n6432 gnd.n775 19.3944
R17576 gnd.n6432 gnd.n6431 19.3944
R17577 gnd.n6431 gnd.n6430 19.3944
R17578 gnd.n6430 gnd.n795 19.3944
R17579 gnd.n6420 gnd.n795 19.3944
R17580 gnd.n6420 gnd.n6419 19.3944
R17581 gnd.n6419 gnd.n6418 19.3944
R17582 gnd.n6418 gnd.n816 19.3944
R17583 gnd.n6408 gnd.n816 19.3944
R17584 gnd.n6408 gnd.n6407 19.3944
R17585 gnd.n5012 gnd.n2066 19.3944
R17586 gnd.n5012 gnd.n2065 19.3944
R17587 gnd.n5025 gnd.n2065 19.3944
R17588 gnd.n5025 gnd.n2063 19.3944
R17589 gnd.n5029 gnd.n2063 19.3944
R17590 gnd.n5029 gnd.n2054 19.3944
R17591 gnd.n5043 gnd.n2054 19.3944
R17592 gnd.n5043 gnd.n2052 19.3944
R17593 gnd.n5047 gnd.n2052 19.3944
R17594 gnd.n5047 gnd.n2042 19.3944
R17595 gnd.n5060 gnd.n2042 19.3944
R17596 gnd.n5060 gnd.n2040 19.3944
R17597 gnd.n5064 gnd.n2040 19.3944
R17598 gnd.n5064 gnd.n2029 19.3944
R17599 gnd.n5079 gnd.n2029 19.3944
R17600 gnd.n5079 gnd.n2026 19.3944
R17601 gnd.n5147 gnd.n2026 19.3944
R17602 gnd.n5147 gnd.n2027 19.3944
R17603 gnd.n5143 gnd.n2027 19.3944
R17604 gnd.n5143 gnd.n5142 19.3944
R17605 gnd.n5142 gnd.n5141 19.3944
R17606 gnd.n5141 gnd.n5085 19.3944
R17607 gnd.n5137 gnd.n5085 19.3944
R17608 gnd.n5137 gnd.n5136 19.3944
R17609 gnd.n5136 gnd.n5135 19.3944
R17610 gnd.n5135 gnd.n5090 19.3944
R17611 gnd.n5131 gnd.n5090 19.3944
R17612 gnd.n5131 gnd.n5130 19.3944
R17613 gnd.n5130 gnd.n5129 19.3944
R17614 gnd.n5129 gnd.n5094 19.3944
R17615 gnd.n5125 gnd.n5094 19.3944
R17616 gnd.n5125 gnd.n5124 19.3944
R17617 gnd.n5124 gnd.n5123 19.3944
R17618 gnd.n5123 gnd.n5098 19.3944
R17619 gnd.n5119 gnd.n5098 19.3944
R17620 gnd.n5119 gnd.n5118 19.3944
R17621 gnd.n5118 gnd.n5117 19.3944
R17622 gnd.n5117 gnd.n5102 19.3944
R17623 gnd.n5113 gnd.n5102 19.3944
R17624 gnd.n5113 gnd.n5112 19.3944
R17625 gnd.n5112 gnd.n5111 19.3944
R17626 gnd.n5111 gnd.n5106 19.3944
R17627 gnd.n5107 gnd.n5106 19.3944
R17628 gnd.n5107 gnd.n1492 19.3944
R17629 gnd.n5370 gnd.n1492 19.3944
R17630 gnd.n5370 gnd.n1489 19.3944
R17631 gnd.n5388 gnd.n1489 19.3944
R17632 gnd.n5388 gnd.n1490 19.3944
R17633 gnd.n5384 gnd.n1490 19.3944
R17634 gnd.n5384 gnd.n5383 19.3944
R17635 gnd.n5383 gnd.n5382 19.3944
R17636 gnd.n5382 gnd.n5377 19.3944
R17637 gnd.n5378 gnd.n5377 19.3944
R17638 gnd.n5378 gnd.n1442 19.3944
R17639 gnd.n5467 gnd.n1442 19.3944
R17640 gnd.n5467 gnd.n1439 19.3944
R17641 gnd.n5482 gnd.n1439 19.3944
R17642 gnd.n5482 gnd.n1440 19.3944
R17643 gnd.n5478 gnd.n1440 19.3944
R17644 gnd.n5478 gnd.n5477 19.3944
R17645 gnd.n5477 gnd.n5476 19.3944
R17646 gnd.n5476 gnd.n5473 19.3944
R17647 gnd.n5473 gnd.n1392 19.3944
R17648 gnd.n5543 gnd.n1392 19.3944
R17649 gnd.n5543 gnd.n1389 19.3944
R17650 gnd.n5551 gnd.n1389 19.3944
R17651 gnd.n5551 gnd.n1390 19.3944
R17652 gnd.n5547 gnd.n1390 19.3944
R17653 gnd.n5547 gnd.n1367 19.3944
R17654 gnd.n5587 gnd.n1367 19.3944
R17655 gnd.n5588 gnd.n5587 19.3944
R17656 gnd.n5588 gnd.n1364 19.3944
R17657 gnd.n5611 gnd.n1364 19.3944
R17658 gnd.n5611 gnd.n1365 19.3944
R17659 gnd.n5607 gnd.n1365 19.3944
R17660 gnd.n5607 gnd.n5606 19.3944
R17661 gnd.n5606 gnd.n5605 19.3944
R17662 gnd.n5605 gnd.n5595 19.3944
R17663 gnd.n5601 gnd.n5595 19.3944
R17664 gnd.n5601 gnd.n5600 19.3944
R17665 gnd.n5600 gnd.n5599 19.3944
R17666 gnd.n5599 gnd.n1217 19.3944
R17667 gnd.n5820 gnd.n1217 19.3944
R17668 gnd.n5820 gnd.n1215 19.3944
R17669 gnd.n5824 gnd.n1215 19.3944
R17670 gnd.n5824 gnd.n1206 19.3944
R17671 gnd.n5837 gnd.n1206 19.3944
R17672 gnd.n5837 gnd.n1204 19.3944
R17673 gnd.n5841 gnd.n1204 19.3944
R17674 gnd.n5841 gnd.n1194 19.3944
R17675 gnd.n5854 gnd.n1194 19.3944
R17676 gnd.n5854 gnd.n1192 19.3944
R17677 gnd.n5858 gnd.n1192 19.3944
R17678 gnd.n5858 gnd.n1183 19.3944
R17679 gnd.n5872 gnd.n1183 19.3944
R17680 gnd.n5872 gnd.n1181 19.3944
R17681 gnd.n5876 gnd.n1181 19.3944
R17682 gnd.n5876 gnd.n1171 19.3944
R17683 gnd.n5891 gnd.n1171 19.3944
R17684 gnd.n5891 gnd.n1169 19.3944
R17685 gnd.n5913 gnd.n1169 19.3944
R17686 gnd.n5910 gnd.n5909 19.3944
R17687 gnd.n5909 gnd.n5908 19.3944
R17688 gnd.n5908 gnd.n5897 19.3944
R17689 gnd.n5904 gnd.n5897 19.3944
R17690 gnd.n5904 gnd.n5903 19.3944
R17691 gnd.n5903 gnd.n1141 19.3944
R17692 gnd.n6096 gnd.n1141 19.3944
R17693 gnd.n6096 gnd.n6095 19.3944
R17694 gnd.n6095 gnd.n6094 19.3944
R17695 gnd.n6094 gnd.n1146 19.3944
R17696 gnd.n6087 gnd.n1146 19.3944
R17697 gnd.n6087 gnd.n6086 19.3944
R17698 gnd.n6086 gnd.n6020 19.3944
R17699 gnd.n6079 gnd.n6020 19.3944
R17700 gnd.n6079 gnd.n6078 19.3944
R17701 gnd.n6078 gnd.n6032 19.3944
R17702 gnd.n6071 gnd.n6032 19.3944
R17703 gnd.n6071 gnd.n6070 19.3944
R17704 gnd.n6070 gnd.n6040 19.3944
R17705 gnd.n6063 gnd.n6040 19.3944
R17706 gnd.n6063 gnd.n6062 19.3944
R17707 gnd.n6062 gnd.n6052 19.3944
R17708 gnd.n6052 gnd.n1014 19.3944
R17709 gnd.n6224 gnd.n1014 19.3944
R17710 gnd.n1027 gnd.n1025 19.3944
R17711 gnd.n1027 gnd.n994 19.3944
R17712 gnd.n6229 gnd.n994 19.3944
R17713 gnd.n5157 gnd.n5156 19.2005
R17714 gnd.n5804 gnd.n1251 19.2005
R17715 gnd.n1583 gnd.n1576 19.1199
R17716 gnd.n5323 gnd.n1495 19.1199
R17717 gnd.n5465 gnd.n1445 19.1199
R17718 gnd.n1361 gnd.n1341 19.1199
R17719 gnd.n1598 gnd.t202 18.8012
R17720 gnd.n1333 gnd.t165 18.8012
R17721 gnd.n7699 gnd.n167 18.8012
R17722 gnd.n6163 gnd.n6162 18.4247
R17723 gnd.n1952 gnd.n1751 18.4247
R17724 gnd.n6221 gnd.n6220 18.2308
R17725 gnd.n7399 gnd.n7398 18.2308
R17726 gnd.n4950 gnd.n2152 18.2308
R17727 gnd.n4218 gnd.n4148 18.2308
R17728 gnd.n3063 gnd.n2957 18.2305
R17729 gnd.n3063 gnd.n3062 18.2305
R17730 gnd.n3071 gnd.n2946 18.2305
R17731 gnd.n3079 gnd.n2946 18.2305
R17732 gnd.n3079 gnd.n2940 18.2305
R17733 gnd.n3087 gnd.n2940 18.2305
R17734 gnd.n3087 gnd.n2933 18.2305
R17735 gnd.n3125 gnd.n2933 18.2305
R17736 gnd.n3135 gnd.n2866 18.2305
R17737 gnd.n4262 gnd.n3909 18.2305
R17738 gnd.n4270 gnd.n2396 18.2305
R17739 gnd.n4282 gnd.n2396 18.2305
R17740 gnd.n4282 gnd.n2388 18.2305
R17741 gnd.n4290 gnd.n2388 18.2305
R17742 gnd.n4302 gnd.n2377 18.2305
R17743 gnd.n4302 gnd.n2380 18.2305
R17744 gnd.n4310 gnd.n2360 18.2305
R17745 gnd.n4322 gnd.n2360 18.2305
R17746 gnd.n4330 gnd.n2352 18.2305
R17747 gnd.n4342 gnd.n2341 18.2305
R17748 gnd.n4342 gnd.n2344 18.2305
R17749 gnd.n4350 gnd.n2324 18.2305
R17750 gnd.n4362 gnd.n2324 18.2305
R17751 gnd.n4370 gnd.n2316 18.2305
R17752 gnd.n4386 gnd.n2304 18.2305
R17753 gnd.n4386 gnd.n2307 18.2305
R17754 gnd.n4396 gnd.n2290 18.2305
R17755 gnd.n4406 gnd.n2290 18.2305
R17756 gnd.n4421 gnd.n2281 18.2305
R17757 gnd.n4431 gnd.n2264 18.2305
R17758 gnd.n4440 gnd.n2264 18.2305
R17759 gnd.n4455 gnd.n2255 18.2305
R17760 gnd.n4465 gnd.n2238 18.2305
R17761 gnd.n4474 gnd.n2238 18.2305
R17762 gnd.n4489 gnd.n2219 18.2305
R17763 gnd.n4499 gnd.n2219 18.2305
R17764 gnd.n4508 gnd.n2212 18.2305
R17765 gnd.n4524 gnd.n2193 18.2305
R17766 gnd.n4535 gnd.n2193 18.2305
R17767 gnd.n4547 gnd.n2185 18.2305
R17768 gnd.n7137 gnd.n335 18.1639
R17769 gnd.n4421 gnd.t272 18.0482
R17770 gnd.n2255 gnd.t314 18.0482
R17771 gnd.n5180 gnd.n1618 17.8452
R17772 gnd.n5248 gnd.n1569 17.8452
R17773 gnd.n5398 gnd.n1481 17.8452
R17774 gnd.n5455 gnd.n5453 17.8452
R17775 gnd.n5621 gnd.n1345 17.8452
R17776 gnd.n5808 gnd.n1228 17.8452
R17777 gnd.t263 gnd.n2316 17.6836
R17778 gnd.n4508 gnd.t242 17.6836
R17779 gnd.t245 gnd.n2352 17.319
R17780 gnd.t26 gnd.n1544 17.2079
R17781 gnd.t169 gnd.n1395 17.2079
R17782 gnd.n7584 gnd.n7454 16.6793
R17783 gnd.n6145 gnd.n6142 16.6793
R17784 gnd.n4069 gnd.n3936 16.6793
R17785 gnd.n1934 gnd.n1933 16.6793
R17786 gnd.n5258 gnd.n1557 16.5706
R17787 gnd.t5 gnd.n5299 16.5706
R17788 gnd.n5409 gnd.n5408 16.5706
R17789 gnd.n1467 gnd.n1466 16.5706
R17790 gnd.n5530 gnd.t153 16.5706
R17791 gnd.n1378 gnd.n1369 16.5706
R17792 gnd.n3909 gnd.t71 16.2252
R17793 gnd.n5318 gnd.t1 15.9333
R17794 gnd.n1425 gnd.t4 15.9333
R17795 gnd.n3758 gnd.n3756 15.6674
R17796 gnd.n3726 gnd.n3724 15.6674
R17797 gnd.n3694 gnd.n3692 15.6674
R17798 gnd.n3663 gnd.n3661 15.6674
R17799 gnd.n3631 gnd.n3629 15.6674
R17800 gnd.n3599 gnd.n3597 15.6674
R17801 gnd.n3567 gnd.n3565 15.6674
R17802 gnd.n3536 gnd.n3534 15.6674
R17803 gnd.n7639 gnd.n7432 15.3217
R17804 gnd.n6102 gnd.n1135 15.3217
R17805 gnd.n4121 gnd.n3915 15.3217
R17806 gnd.n6403 gnd.n840 15.3217
R17807 gnd.n5258 gnd.n5257 15.296
R17808 gnd.n5275 gnd.n1552 15.296
R17809 gnd.t12 gnd.n1503 15.296
R17810 gnd.n5409 gnd.n1472 15.296
R17811 gnd.n1466 gnd.n1460 15.296
R17812 gnd.n5492 gnd.t177 15.296
R17813 gnd.n5554 gnd.n5553 15.296
R17814 gnd.n5584 gnd.n1369 15.296
R17815 gnd.t46 gnd.n1309 15.296
R17816 gnd.n1236 gnd.n1235 15.0827
R17817 gnd.n1640 gnd.n1635 15.0481
R17818 gnd.n1246 gnd.n1245 15.0481
R17819 gnd.t19 gnd.n1494 14.6587
R17820 gnd.n5421 gnd.t170 14.6587
R17821 gnd.n5593 gnd.t43 14.6587
R17822 gnd.n5186 gnd.t178 14.34
R17823 gnd.t167 gnd.n5677 14.34
R17824 gnd.n3147 gnd.n2867 14.2199
R17825 gnd.n3157 gnd.n2850 14.2199
R17826 gnd.n2853 gnd.n2841 14.2199
R17827 gnd.n3178 gnd.n2842 14.2199
R17828 gnd.n3188 gnd.n2822 14.2199
R17829 gnd.n3198 gnd.n3197 14.2199
R17830 gnd.n2808 gnd.n2806 14.2199
R17831 gnd.n3229 gnd.n3228 14.2199
R17832 gnd.n3244 gnd.n2791 14.2199
R17833 gnd.n3298 gnd.n2730 14.2199
R17834 gnd.n3254 gnd.n2731 14.2199
R17835 gnd.n3291 gnd.n2742 14.2199
R17836 gnd.n2780 gnd.n2779 14.2199
R17837 gnd.n3285 gnd.n3284 14.2199
R17838 gnd.n2766 gnd.n2753 14.2199
R17839 gnd.n3324 gnd.n3323 14.2199
R17840 gnd.n3334 gnd.n2630 14.2199
R17841 gnd.n3346 gnd.n2622 14.2199
R17842 gnd.n3345 gnd.n2610 14.2199
R17843 gnd.n3364 gnd.n3363 14.2199
R17844 gnd.n3374 gnd.n2603 14.2199
R17845 gnd.n3385 gnd.n2591 14.2199
R17846 gnd.n3409 gnd.n3408 14.2199
R17847 gnd.n3420 gnd.n2574 14.2199
R17848 gnd.n3419 gnd.n2576 14.2199
R17849 gnd.n3431 gnd.n2567 14.2199
R17850 gnd.n3449 gnd.n3448 14.2199
R17851 gnd.n2558 gnd.n2547 14.2199
R17852 gnd.n3470 gnd.n2535 14.2199
R17853 gnd.n3498 gnd.n3497 14.2199
R17854 gnd.n3509 gnd.n2520 14.2199
R17855 gnd.n3520 gnd.n2513 14.2199
R17856 gnd.n3519 gnd.n2501 14.2199
R17857 gnd.n3792 gnd.n3791 14.2199
R17858 gnd.n3814 gnd.n2486 14.2199
R17859 gnd.n5249 gnd.n5248 14.0214
R17860 gnd.n1544 gnd.n1536 14.0214
R17861 gnd.n5391 gnd.t23 14.0214
R17862 gnd.n5390 gnd.n1481 14.0214
R17863 gnd.n5453 gnd.n1455 14.0214
R17864 gnd.n5435 gnd.t7 14.0214
R17865 gnd.n5541 gnd.n1395 14.0214
R17866 gnd.n5621 gnd.n5620 14.0214
R17867 gnd.n5810 gnd.n5808 14.0214
R17868 gnd.n5338 gnd.t198 13.7027
R17869 gnd.n5485 gnd.t208 13.7027
R17870 gnd.n7126 gnd.n335 13.7027
R17871 gnd.n2928 gnd.n2927 13.5763
R17872 gnd.n3872 gnd.n2450 13.5763
R17873 gnd.n5327 gnd.t151 13.384
R17874 gnd.n5442 gnd.t2 13.384
R17875 gnd.n3168 gnd.t206 13.3084
R17876 gnd.n4290 gnd.t220 13.3084
R17877 gnd.n1651 gnd.n1632 13.1884
R17878 gnd.n1646 gnd.n1645 13.1884
R17879 gnd.n1645 gnd.n1644 13.1884
R17880 gnd.n1239 gnd.n1234 13.1884
R17881 gnd.n1240 gnd.n1239 13.1884
R17882 gnd.n1647 gnd.n1634 13.146
R17883 gnd.n1643 gnd.n1634 13.146
R17884 gnd.n1238 gnd.n1237 13.146
R17885 gnd.n1238 gnd.n1233 13.146
R17886 gnd.n2869 gnd.t57 12.9438
R17887 gnd.n4330 gnd.t232 12.9438
R17888 gnd.n3759 gnd.n3755 12.8005
R17889 gnd.n3727 gnd.n3723 12.8005
R17890 gnd.n3695 gnd.n3691 12.8005
R17891 gnd.n3664 gnd.n3660 12.8005
R17892 gnd.n3632 gnd.n3628 12.8005
R17893 gnd.n3600 gnd.n3596 12.8005
R17894 gnd.n3568 gnd.n3564 12.8005
R17895 gnd.n3537 gnd.n3533 12.8005
R17896 gnd.n1612 gnd.n1608 12.7467
R17897 gnd.n5212 gnd.t104 12.7467
R17898 gnd.n5227 gnd.n1583 12.7467
R17899 gnd.n5368 gnd.n1495 12.7467
R17900 gnd.n5420 gnd.n1445 12.7467
R17901 gnd.n5614 gnd.n1361 12.7467
R17902 gnd.n5683 gnd.t91 12.7467
R17903 gnd.n4370 gnd.t224 12.5792
R17904 gnd.t226 gnd.n2212 12.5792
R17905 gnd.n6434 gnd.t316 12.4281
R17906 gnd.n5041 gnd.t204 12.4281
R17907 gnd.n5860 gnd.t154 12.4281
R17908 gnd.n7044 gnd.t255 12.4281
R17909 gnd.n213 gnd.t240 12.4281
R17910 gnd.n2927 gnd.n2922 12.4126
R17911 gnd.n3875 gnd.n3872 12.4126
R17912 gnd.t173 gnd.n2874 12.2146
R17913 gnd.n2281 gnd.t222 12.2146
R17914 gnd.n4455 gnd.t290 12.2146
R17915 gnd.n5156 gnd.n5155 12.1761
R17916 gnd.n1252 gnd.n1251 12.1761
R17917 gnd.n852 gnd.n843 12.1094
R17918 gnd.t50 gnd.n5179 12.1094
R17919 gnd.n6215 gnd.n1069 12.1094
R17920 gnd.n3763 gnd.n3762 12.0247
R17921 gnd.n3731 gnd.n3730 12.0247
R17922 gnd.n3699 gnd.n3698 12.0247
R17923 gnd.n3668 gnd.n3667 12.0247
R17924 gnd.n3636 gnd.n3635 12.0247
R17925 gnd.n3604 gnd.n3603 12.0247
R17926 gnd.n3572 gnd.n3571 12.0247
R17927 gnd.n3541 gnd.n3540 12.0247
R17928 gnd.t189 gnd.n2548 11.85
R17929 gnd.n4396 gnd.t276 11.85
R17930 gnd.n4474 gnd.t258 11.85
R17931 gnd.n4901 gnd.t316 11.7908
R17932 gnd.t255 gnd.n374 11.7908
R17933 gnd.n338 gnd.t214 11.7908
R17934 gnd.n175 gnd.t278 11.7908
R17935 gnd.t191 gnd.n2583 11.4854
R17936 gnd.n4350 gnd.t260 11.4854
R17937 gnd.n4535 gnd.t294 11.4854
R17938 gnd.n5199 gnd.n1604 11.4721
R17939 gnd.n5219 gnd.n5218 11.4721
R17940 gnd.n5318 gnd.n1517 11.4721
R17941 gnd.n5358 gnd.n5357 11.4721
R17942 gnd.n5493 gnd.n1431 11.4721
R17943 gnd.n5501 gnd.n1425 11.4721
R17944 gnd.n5640 gnd.n1334 11.4721
R17945 gnd.n5662 gnd.n5660 11.4721
R17946 gnd.n3766 gnd.n3753 11.249
R17947 gnd.n3734 gnd.n3721 11.249
R17948 gnd.n3702 gnd.n3689 11.249
R17949 gnd.n3671 gnd.n3658 11.249
R17950 gnd.n3639 gnd.n3626 11.249
R17951 gnd.n3607 gnd.n3594 11.249
R17952 gnd.n3575 gnd.n3562 11.249
R17953 gnd.n3544 gnd.n3531 11.249
R17954 gnd.n5299 gnd.t171 11.1535
R17955 gnd.t147 gnd.n5530 11.1535
R17956 gnd.n301 gnd.t266 11.1535
R17957 gnd.n136 gnd.t236 11.1535
R17958 gnd.n3335 gnd.t197 11.1208
R17959 gnd.n4310 gnd.t285 11.1208
R17960 gnd.n3292 gnd.t187 10.7562
R17961 gnd.n3277 gnd.t24 10.7562
R17962 gnd.n7634 gnd.n7432 10.6672
R17963 gnd.n6105 gnd.n6102 10.6672
R17964 gnd.n3916 gnd.n3915 10.6672
R17965 gnd.n1899 gnd.n840 10.6672
R17966 gnd.n5739 gnd.n1280 10.6151
R17967 gnd.n5739 gnd.n5738 10.6151
R17968 gnd.n5736 gnd.n1284 10.6151
R17969 gnd.n5731 gnd.n1284 10.6151
R17970 gnd.n5731 gnd.n5730 10.6151
R17971 gnd.n5730 gnd.n5729 10.6151
R17972 gnd.n5729 gnd.n1287 10.6151
R17973 gnd.n5724 gnd.n1287 10.6151
R17974 gnd.n5724 gnd.n5723 10.6151
R17975 gnd.n5723 gnd.n5722 10.6151
R17976 gnd.n5722 gnd.n1290 10.6151
R17977 gnd.n5717 gnd.n1290 10.6151
R17978 gnd.n5717 gnd.n5716 10.6151
R17979 gnd.n5716 gnd.n5715 10.6151
R17980 gnd.n5715 gnd.n1293 10.6151
R17981 gnd.n5710 gnd.n1293 10.6151
R17982 gnd.n5710 gnd.n5709 10.6151
R17983 gnd.n5709 gnd.n5708 10.6151
R17984 gnd.n5708 gnd.n1296 10.6151
R17985 gnd.n5703 gnd.n1296 10.6151
R17986 gnd.n5703 gnd.n5702 10.6151
R17987 gnd.n5702 gnd.n5701 10.6151
R17988 gnd.n5701 gnd.n1299 10.6151
R17989 gnd.n5696 gnd.n1299 10.6151
R17990 gnd.n5696 gnd.n5695 10.6151
R17991 gnd.n5695 gnd.n5694 10.6151
R17992 gnd.n5694 gnd.n1302 10.6151
R17993 gnd.n5689 gnd.n1302 10.6151
R17994 gnd.n5689 gnd.n5688 10.6151
R17995 gnd.n5688 gnd.n5687 10.6151
R17996 gnd.n2021 gnd.n2020 10.6151
R17997 gnd.n2020 gnd.n2018 10.6151
R17998 gnd.n2018 gnd.n1610 10.6151
R17999 gnd.n5188 gnd.n1610 10.6151
R18000 gnd.n5189 gnd.n5188 10.6151
R18001 gnd.n5190 gnd.n5189 10.6151
R18002 gnd.n5190 gnd.n1600 10.6151
R18003 gnd.n5201 gnd.n1600 10.6151
R18004 gnd.n5202 gnd.n5201 10.6151
R18005 gnd.n5210 gnd.n5202 10.6151
R18006 gnd.n5210 gnd.n5209 10.6151
R18007 gnd.n5209 gnd.n5208 10.6151
R18008 gnd.n5208 gnd.n5207 10.6151
R18009 gnd.n5207 gnd.n5205 10.6151
R18010 gnd.n5205 gnd.n5204 10.6151
R18011 gnd.n5204 gnd.n1573 10.6151
R18012 gnd.n5237 gnd.n1573 10.6151
R18013 gnd.n5238 gnd.n5237 10.6151
R18014 gnd.n5239 gnd.n5238 10.6151
R18015 gnd.n5239 gnd.n1559 10.6151
R18016 gnd.n5260 gnd.n1559 10.6151
R18017 gnd.n5261 gnd.n5260 10.6151
R18018 gnd.n5266 gnd.n5261 10.6151
R18019 gnd.n5266 gnd.n5265 10.6151
R18020 gnd.n5265 gnd.n5264 10.6151
R18021 gnd.n5264 gnd.n5262 10.6151
R18022 gnd.n5262 gnd.n1533 10.6151
R18023 gnd.n5294 gnd.n1533 10.6151
R18024 gnd.n5295 gnd.n5294 10.6151
R18025 gnd.n5297 gnd.n5295 10.6151
R18026 gnd.n5297 gnd.n5296 10.6151
R18027 gnd.n5296 gnd.n1514 10.6151
R18028 gnd.n5320 gnd.n1514 10.6151
R18029 gnd.n5321 gnd.n5320 10.6151
R18030 gnd.n5344 gnd.n5321 10.6151
R18031 gnd.n5344 gnd.n5343 10.6151
R18032 gnd.n5343 gnd.n5342 10.6151
R18033 gnd.n5342 gnd.n5341 10.6151
R18034 gnd.n5341 gnd.n5322 10.6151
R18035 gnd.n5335 gnd.n5322 10.6151
R18036 gnd.n5335 gnd.n5334 10.6151
R18037 gnd.n5334 gnd.n5333 10.6151
R18038 gnd.n5333 gnd.n5332 10.6151
R18039 gnd.n5332 gnd.n5330 10.6151
R18040 gnd.n5330 gnd.n5329 10.6151
R18041 gnd.n5329 gnd.n5326 10.6151
R18042 gnd.n5326 gnd.n1463 10.6151
R18043 gnd.n5417 gnd.n1463 10.6151
R18044 gnd.n5418 gnd.n5417 10.6151
R18045 gnd.n5440 gnd.n5418 10.6151
R18046 gnd.n5440 gnd.n5439 10.6151
R18047 gnd.n5439 gnd.n5438 10.6151
R18048 gnd.n5438 gnd.n5437 10.6151
R18049 gnd.n5437 gnd.n5419 10.6151
R18050 gnd.n5432 gnd.n5419 10.6151
R18051 gnd.n5432 gnd.n5431 10.6151
R18052 gnd.n5431 gnd.n5430 10.6151
R18053 gnd.n5430 gnd.n5429 10.6151
R18054 gnd.n5429 gnd.n5427 10.6151
R18055 gnd.n5427 gnd.n5426 10.6151
R18056 gnd.n5426 gnd.n5424 10.6151
R18057 gnd.n5424 gnd.n5423 10.6151
R18058 gnd.n5423 gnd.n1415 10.6151
R18059 gnd.n5511 gnd.n1415 10.6151
R18060 gnd.n5512 gnd.n5511 10.6151
R18061 gnd.n5513 gnd.n5512 10.6151
R18062 gnd.n5518 gnd.n5513 10.6151
R18063 gnd.n5519 gnd.n5518 10.6151
R18064 gnd.n5520 gnd.n5519 10.6151
R18065 gnd.n5520 gnd.n1385 10.6151
R18066 gnd.n5556 gnd.n1385 10.6151
R18067 gnd.n5557 gnd.n5556 10.6151
R18068 gnd.n5558 gnd.n5557 10.6151
R18069 gnd.n5561 gnd.n5558 10.6151
R18070 gnd.n5562 gnd.n5561 10.6151
R18071 gnd.n5564 gnd.n5562 10.6151
R18072 gnd.n5564 gnd.n5563 10.6151
R18073 gnd.n5563 gnd.n1339 10.6151
R18074 gnd.n5629 gnd.n1339 10.6151
R18075 gnd.n5630 gnd.n5629 10.6151
R18076 gnd.n5631 gnd.n5630 10.6151
R18077 gnd.n5631 gnd.n1330 10.6151
R18078 gnd.n5642 gnd.n1330 10.6151
R18079 gnd.n5643 gnd.n5642 10.6151
R18080 gnd.n5652 gnd.n5643 10.6151
R18081 gnd.n5652 gnd.n5651 10.6151
R18082 gnd.n5651 gnd.n5650 10.6151
R18083 gnd.n5650 gnd.n5649 10.6151
R18084 gnd.n5649 gnd.n5647 10.6151
R18085 gnd.n5647 gnd.n5646 10.6151
R18086 gnd.n5646 gnd.n1307 10.6151
R18087 gnd.n5680 gnd.n1307 10.6151
R18088 gnd.n5681 gnd.n5680 10.6151
R18089 gnd.n5682 gnd.n5681 10.6151
R18090 gnd.n5682 gnd.n1305 10.6151
R18091 gnd.n1958 gnd.n1957 10.6151
R18092 gnd.n1961 gnd.n1958 10.6151
R18093 gnd.n1966 gnd.n1963 10.6151
R18094 gnd.n1967 gnd.n1966 10.6151
R18095 gnd.n1970 gnd.n1967 10.6151
R18096 gnd.n1971 gnd.n1970 10.6151
R18097 gnd.n1974 gnd.n1971 10.6151
R18098 gnd.n1975 gnd.n1974 10.6151
R18099 gnd.n1978 gnd.n1975 10.6151
R18100 gnd.n1979 gnd.n1978 10.6151
R18101 gnd.n1982 gnd.n1979 10.6151
R18102 gnd.n1983 gnd.n1982 10.6151
R18103 gnd.n1986 gnd.n1983 10.6151
R18104 gnd.n1987 gnd.n1986 10.6151
R18105 gnd.n1990 gnd.n1987 10.6151
R18106 gnd.n1991 gnd.n1990 10.6151
R18107 gnd.n1994 gnd.n1991 10.6151
R18108 gnd.n1995 gnd.n1994 10.6151
R18109 gnd.n1998 gnd.n1995 10.6151
R18110 gnd.n1999 gnd.n1998 10.6151
R18111 gnd.n2002 gnd.n1999 10.6151
R18112 gnd.n2003 gnd.n2002 10.6151
R18113 gnd.n2006 gnd.n2003 10.6151
R18114 gnd.n2007 gnd.n2006 10.6151
R18115 gnd.n2010 gnd.n2007 10.6151
R18116 gnd.n2011 gnd.n2010 10.6151
R18117 gnd.n2014 gnd.n2011 10.6151
R18118 gnd.n2016 gnd.n2014 10.6151
R18119 gnd.n2017 gnd.n2016 10.6151
R18120 gnd.n2022 gnd.n2017 10.6151
R18121 gnd.n5155 gnd.n5154 10.6151
R18122 gnd.n5154 gnd.n1652 10.6151
R18123 gnd.n1693 gnd.n1652 10.6151
R18124 gnd.n1694 gnd.n1693 10.6151
R18125 gnd.n1697 gnd.n1694 10.6151
R18126 gnd.n1698 gnd.n1697 10.6151
R18127 gnd.n1701 gnd.n1698 10.6151
R18128 gnd.n1702 gnd.n1701 10.6151
R18129 gnd.n1705 gnd.n1702 10.6151
R18130 gnd.n1706 gnd.n1705 10.6151
R18131 gnd.n1709 gnd.n1706 10.6151
R18132 gnd.n1710 gnd.n1709 10.6151
R18133 gnd.n1713 gnd.n1710 10.6151
R18134 gnd.n1714 gnd.n1713 10.6151
R18135 gnd.n1717 gnd.n1714 10.6151
R18136 gnd.n1718 gnd.n1717 10.6151
R18137 gnd.n1721 gnd.n1718 10.6151
R18138 gnd.n1722 gnd.n1721 10.6151
R18139 gnd.n1725 gnd.n1722 10.6151
R18140 gnd.n1726 gnd.n1725 10.6151
R18141 gnd.n1729 gnd.n1726 10.6151
R18142 gnd.n1730 gnd.n1729 10.6151
R18143 gnd.n1733 gnd.n1730 10.6151
R18144 gnd.n1734 gnd.n1733 10.6151
R18145 gnd.n1737 gnd.n1734 10.6151
R18146 gnd.n1738 gnd.n1737 10.6151
R18147 gnd.n1741 gnd.n1738 10.6151
R18148 gnd.n1742 gnd.n1741 10.6151
R18149 gnd.n1746 gnd.n1745 10.6151
R18150 gnd.n1749 gnd.n1746 10.6151
R18151 gnd.n5799 gnd.n1252 10.6151
R18152 gnd.n5799 gnd.n5798 10.6151
R18153 gnd.n5798 gnd.n5797 10.6151
R18154 gnd.n5797 gnd.n1255 10.6151
R18155 gnd.n5792 gnd.n1255 10.6151
R18156 gnd.n5792 gnd.n5791 10.6151
R18157 gnd.n5791 gnd.n5790 10.6151
R18158 gnd.n5790 gnd.n1258 10.6151
R18159 gnd.n5785 gnd.n1258 10.6151
R18160 gnd.n5785 gnd.n5784 10.6151
R18161 gnd.n5784 gnd.n5783 10.6151
R18162 gnd.n5783 gnd.n1261 10.6151
R18163 gnd.n5778 gnd.n1261 10.6151
R18164 gnd.n5778 gnd.n5777 10.6151
R18165 gnd.n5777 gnd.n5776 10.6151
R18166 gnd.n5776 gnd.n1264 10.6151
R18167 gnd.n5771 gnd.n1264 10.6151
R18168 gnd.n5771 gnd.n5770 10.6151
R18169 gnd.n5770 gnd.n5769 10.6151
R18170 gnd.n5769 gnd.n1267 10.6151
R18171 gnd.n5764 gnd.n1267 10.6151
R18172 gnd.n5764 gnd.n5763 10.6151
R18173 gnd.n5763 gnd.n5762 10.6151
R18174 gnd.n5762 gnd.n1270 10.6151
R18175 gnd.n5757 gnd.n1270 10.6151
R18176 gnd.n5757 gnd.n5756 10.6151
R18177 gnd.n5756 gnd.n5755 10.6151
R18178 gnd.n5755 gnd.n1273 10.6151
R18179 gnd.n5750 gnd.n5749 10.6151
R18180 gnd.n5749 gnd.n5748 10.6151
R18181 gnd.n5157 gnd.n1616 10.6151
R18182 gnd.n5182 gnd.n1616 10.6151
R18183 gnd.n5183 gnd.n5182 10.6151
R18184 gnd.n5184 gnd.n5183 10.6151
R18185 gnd.n5184 gnd.n1606 10.6151
R18186 gnd.n5195 gnd.n1606 10.6151
R18187 gnd.n5196 gnd.n5195 10.6151
R18188 gnd.n5197 gnd.n5196 10.6151
R18189 gnd.n5197 gnd.n1593 10.6151
R18190 gnd.n5214 gnd.n1593 10.6151
R18191 gnd.n5215 gnd.n5214 10.6151
R18192 gnd.n5216 gnd.n5215 10.6151
R18193 gnd.n5216 gnd.n1578 10.6151
R18194 gnd.n5230 gnd.n1578 10.6151
R18195 gnd.n5231 gnd.n5230 10.6151
R18196 gnd.n5232 gnd.n5231 10.6151
R18197 gnd.n5232 gnd.n1572 10.6151
R18198 gnd.n5246 gnd.n1572 10.6151
R18199 gnd.n5246 gnd.n5245 10.6151
R18200 gnd.n5245 gnd.n5244 10.6151
R18201 gnd.n5244 gnd.n1554 10.6151
R18202 gnd.n5271 gnd.n1554 10.6151
R18203 gnd.n5272 gnd.n5271 10.6151
R18204 gnd.n5273 gnd.n5272 10.6151
R18205 gnd.n5273 gnd.n1539 10.6151
R18206 gnd.n5287 gnd.n1539 10.6151
R18207 gnd.n5288 gnd.n5287 10.6151
R18208 gnd.n5290 gnd.n5288 10.6151
R18209 gnd.n5290 gnd.n5289 10.6151
R18210 gnd.n5289 gnd.n1519 10.6151
R18211 gnd.n5314 gnd.n1519 10.6151
R18212 gnd.n5315 gnd.n5314 10.6151
R18213 gnd.n5316 gnd.n5315 10.6151
R18214 gnd.n5316 gnd.n1508 10.6151
R18215 gnd.n5348 gnd.n1508 10.6151
R18216 gnd.n5349 gnd.n5348 10.6151
R18217 gnd.n5355 gnd.n5349 10.6151
R18218 gnd.n5355 gnd.n5354 10.6151
R18219 gnd.n5354 gnd.n5353 10.6151
R18220 gnd.n5353 gnd.n5350 10.6151
R18221 gnd.n5350 gnd.n1485 10.6151
R18222 gnd.n5393 gnd.n1485 10.6151
R18223 gnd.n5394 gnd.n5393 10.6151
R18224 gnd.n5395 gnd.n5394 10.6151
R18225 gnd.n5395 gnd.n1469 10.6151
R18226 gnd.n5411 gnd.n1469 10.6151
R18227 gnd.n5412 gnd.n5411 10.6151
R18228 gnd.n5413 gnd.n5412 10.6151
R18229 gnd.n5413 gnd.n1458 10.6151
R18230 gnd.n5444 gnd.n1458 10.6151
R18231 gnd.n5445 gnd.n5444 10.6151
R18232 gnd.n5451 gnd.n5445 10.6151
R18233 gnd.n5451 gnd.n5450 10.6151
R18234 gnd.n5450 gnd.n5449 10.6151
R18235 gnd.n5449 gnd.n5446 10.6151
R18236 gnd.n5446 gnd.n1435 10.6151
R18237 gnd.n5488 gnd.n1435 10.6151
R18238 gnd.n5489 gnd.n5488 10.6151
R18239 gnd.n5490 gnd.n5489 10.6151
R18240 gnd.n5490 gnd.n1420 10.6151
R18241 gnd.n5504 gnd.n1420 10.6151
R18242 gnd.n5505 gnd.n5504 10.6151
R18243 gnd.n5506 gnd.n5505 10.6151
R18244 gnd.n5506 gnd.n1407 10.6151
R18245 gnd.n5528 gnd.n1407 10.6151
R18246 gnd.n5528 gnd.n5527 10.6151
R18247 gnd.n5527 gnd.n5526 10.6151
R18248 gnd.n5526 gnd.n1408 10.6151
R18249 gnd.n1411 gnd.n1408 10.6151
R18250 gnd.n1411 gnd.n1410 10.6151
R18251 gnd.n1410 gnd.n1382 10.6151
R18252 gnd.n5572 gnd.n1382 10.6151
R18253 gnd.n5572 gnd.n5571 10.6151
R18254 gnd.n5571 gnd.n5570 10.6151
R18255 gnd.n5570 gnd.n1383 10.6151
R18256 gnd.n1383 gnd.n1343 10.6151
R18257 gnd.n5623 gnd.n1343 10.6151
R18258 gnd.n5624 gnd.n5623 10.6151
R18259 gnd.n5625 gnd.n5624 10.6151
R18260 gnd.n5625 gnd.n1336 10.6151
R18261 gnd.n5636 gnd.n1336 10.6151
R18262 gnd.n5637 gnd.n5636 10.6151
R18263 gnd.n5638 gnd.n5637 10.6151
R18264 gnd.n5638 gnd.n1325 10.6151
R18265 gnd.n5656 gnd.n1325 10.6151
R18266 gnd.n5657 gnd.n5656 10.6151
R18267 gnd.n5658 gnd.n5657 10.6151
R18268 gnd.n5658 gnd.n1311 10.6151
R18269 gnd.n5673 gnd.n1311 10.6151
R18270 gnd.n5674 gnd.n5673 10.6151
R18271 gnd.n5675 gnd.n5674 10.6151
R18272 gnd.n5675 gnd.n1231 10.6151
R18273 gnd.n5806 gnd.n1231 10.6151
R18274 gnd.n5806 gnd.n5805 10.6151
R18275 gnd.n5805 gnd.n5804 10.6151
R18276 gnd.n3136 gnd.n3135 10.5739
R18277 gnd.n5276 gnd.t15 10.5161
R18278 gnd.n5575 gnd.t163 10.5161
R18279 gnd.n7224 gnd.t247 10.5161
R18280 gnd.n7232 gnd.t230 10.5161
R18281 gnd.n3767 gnd.n3751 10.4732
R18282 gnd.n3735 gnd.n3719 10.4732
R18283 gnd.n3703 gnd.n3687 10.4732
R18284 gnd.n3672 gnd.n3656 10.4732
R18285 gnd.n3640 gnd.n3624 10.4732
R18286 gnd.n3608 gnd.n3592 10.4732
R18287 gnd.n3576 gnd.n3560 10.4732
R18288 gnd.n3545 gnd.n3529 10.4732
R18289 gnd.t188 gnd.n2816 10.3916
R18290 gnd.n4547 gnd.n753 10.3916
R18291 gnd.n1604 gnd.n1603 10.1975
R18292 gnd.n1517 gnd.n1510 10.1975
R18293 gnd.n5358 gnd.n1503 10.1975
R18294 gnd.n5493 gnd.n5492 10.1975
R18295 gnd.n5502 gnd.n5501 10.1975
R18296 gnd.n5662 gnd.n1321 10.1975
R18297 gnd.n2844 gnd.t185 10.027
R18298 gnd.t301 gnd.n298 9.87883
R18299 gnd.t318 gnd.n139 9.87883
R18300 gnd.n3771 gnd.n3770 9.69747
R18301 gnd.n3739 gnd.n3738 9.69747
R18302 gnd.n3707 gnd.n3706 9.69747
R18303 gnd.n3676 gnd.n3675 9.69747
R18304 gnd.n3644 gnd.n3643 9.69747
R18305 gnd.n3612 gnd.n3611 9.69747
R18306 gnd.n3580 gnd.n3579 9.69747
R18307 gnd.n3549 gnd.n3548 9.69747
R18308 gnd.n3243 gnd.t196 9.66242
R18309 gnd.n3777 gnd.n3776 9.45567
R18310 gnd.n3745 gnd.n3744 9.45567
R18311 gnd.n3713 gnd.n3712 9.45567
R18312 gnd.n3682 gnd.n3681 9.45567
R18313 gnd.n3650 gnd.n3649 9.45567
R18314 gnd.n3618 gnd.n3617 9.45567
R18315 gnd.n3586 gnd.n3585 9.45567
R18316 gnd.n3555 gnd.n3554 9.45567
R18317 gnd.n7590 gnd.n7454 9.30959
R18318 gnd.n6142 gnd.n6141 9.30959
R18319 gnd.n4069 gnd.n3934 9.30959
R18320 gnd.n1933 gnd.n1862 9.30959
R18321 gnd.n6102 gnd.n6101 9.3005
R18322 gnd.n6105 gnd.n1134 9.3005
R18323 gnd.n6106 gnd.n1133 9.3005
R18324 gnd.n6109 gnd.n1132 9.3005
R18325 gnd.n6110 gnd.n1131 9.3005
R18326 gnd.n6113 gnd.n1130 9.3005
R18327 gnd.n6114 gnd.n1129 9.3005
R18328 gnd.n6117 gnd.n1128 9.3005
R18329 gnd.n6118 gnd.n1127 9.3005
R18330 gnd.n6121 gnd.n1126 9.3005
R18331 gnd.n6122 gnd.n1125 9.3005
R18332 gnd.n6125 gnd.n1124 9.3005
R18333 gnd.n6126 gnd.n1123 9.3005
R18334 gnd.n6129 gnd.n1122 9.3005
R18335 gnd.n6130 gnd.n1121 9.3005
R18336 gnd.n6133 gnd.n1120 9.3005
R18337 gnd.n6134 gnd.n1119 9.3005
R18338 gnd.n6137 gnd.n1118 9.3005
R18339 gnd.n6138 gnd.n1117 9.3005
R18340 gnd.n6141 gnd.n1116 9.3005
R18341 gnd.n6145 gnd.n1112 9.3005
R18342 gnd.n6146 gnd.n1111 9.3005
R18343 gnd.n6149 gnd.n1110 9.3005
R18344 gnd.n6150 gnd.n1109 9.3005
R18345 gnd.n6153 gnd.n1108 9.3005
R18346 gnd.n6154 gnd.n1107 9.3005
R18347 gnd.n6157 gnd.n1106 9.3005
R18348 gnd.n6158 gnd.n1105 9.3005
R18349 gnd.n6161 gnd.n1104 9.3005
R18350 gnd.n6163 gnd.n1100 9.3005
R18351 gnd.n6166 gnd.n1099 9.3005
R18352 gnd.n6167 gnd.n1098 9.3005
R18353 gnd.n6170 gnd.n1097 9.3005
R18354 gnd.n6171 gnd.n1096 9.3005
R18355 gnd.n6174 gnd.n1095 9.3005
R18356 gnd.n6175 gnd.n1094 9.3005
R18357 gnd.n6178 gnd.n1093 9.3005
R18358 gnd.n6180 gnd.n1090 9.3005
R18359 gnd.n6183 gnd.n1089 9.3005
R18360 gnd.n6184 gnd.n1088 9.3005
R18361 gnd.n6187 gnd.n1087 9.3005
R18362 gnd.n6188 gnd.n1086 9.3005
R18363 gnd.n6191 gnd.n1085 9.3005
R18364 gnd.n6192 gnd.n1084 9.3005
R18365 gnd.n6195 gnd.n1083 9.3005
R18366 gnd.n6196 gnd.n1082 9.3005
R18367 gnd.n6199 gnd.n1081 9.3005
R18368 gnd.n6200 gnd.n1080 9.3005
R18369 gnd.n6203 gnd.n1079 9.3005
R18370 gnd.n6204 gnd.n1078 9.3005
R18371 gnd.n6207 gnd.n1077 9.3005
R18372 gnd.n6209 gnd.n1076 9.3005
R18373 gnd.n6210 gnd.n1075 9.3005
R18374 gnd.n6211 gnd.n1074 9.3005
R18375 gnd.n6212 gnd.n1073 9.3005
R18376 gnd.n6142 gnd.n1113 9.3005
R18377 gnd.n6100 gnd.n1135 9.3005
R18378 gnd.n5995 gnd.n5994 9.3005
R18379 gnd.n5996 gnd.n5990 9.3005
R18380 gnd.n6000 gnd.n5997 9.3005
R18381 gnd.n5999 gnd.n5998 9.3005
R18382 gnd.n389 gnd.n388 9.3005
R18383 gnd.n7054 gnd.n7053 9.3005
R18384 gnd.n7055 gnd.n387 9.3005
R18385 gnd.n7059 gnd.n7056 9.3005
R18386 gnd.n7058 gnd.n7057 9.3005
R18387 gnd.n360 gnd.n359 9.3005
R18388 gnd.n7090 gnd.n7089 9.3005
R18389 gnd.n7091 gnd.n358 9.3005
R18390 gnd.n7095 gnd.n7092 9.3005
R18391 gnd.n7094 gnd.n7093 9.3005
R18392 gnd.n333 gnd.n332 9.3005
R18393 gnd.n7140 gnd.n7139 9.3005
R18394 gnd.n7141 gnd.n331 9.3005
R18395 gnd.n7143 gnd.n7142 9.3005
R18396 gnd.n316 gnd.n315 9.3005
R18397 gnd.n7160 gnd.n7159 9.3005
R18398 gnd.n7161 gnd.n314 9.3005
R18399 gnd.n7163 gnd.n7162 9.3005
R18400 gnd.n296 gnd.n295 9.3005
R18401 gnd.n7184 gnd.n7183 9.3005
R18402 gnd.n7185 gnd.n294 9.3005
R18403 gnd.n7189 gnd.n7186 9.3005
R18404 gnd.n7188 gnd.n7187 9.3005
R18405 gnd.n5992 gnd.n5991 9.3005
R18406 gnd.n273 gnd.n272 9.3005
R18407 gnd.n7216 gnd.n7215 9.3005
R18408 gnd.n7217 gnd.n271 9.3005
R18409 gnd.n7222 gnd.n7218 9.3005
R18410 gnd.n7221 gnd.n7220 9.3005
R18411 gnd.n7219 gnd.n110 9.3005
R18412 gnd.n7733 gnd.n111 9.3005
R18413 gnd.n7732 gnd.n112 9.3005
R18414 gnd.n7731 gnd.n113 9.3005
R18415 gnd.n130 gnd.n114 9.3005
R18416 gnd.n7721 gnd.n131 9.3005
R18417 gnd.n7720 gnd.n132 9.3005
R18418 gnd.n7719 gnd.n133 9.3005
R18419 gnd.n150 gnd.n134 9.3005
R18420 gnd.n7709 gnd.n151 9.3005
R18421 gnd.n7708 gnd.n152 9.3005
R18422 gnd.n7707 gnd.n153 9.3005
R18423 gnd.n169 gnd.n154 9.3005
R18424 gnd.n7697 gnd.n170 9.3005
R18425 gnd.n7696 gnd.n171 9.3005
R18426 gnd.n7695 gnd.n172 9.3005
R18427 gnd.n189 gnd.n173 9.3005
R18428 gnd.n7685 gnd.n190 9.3005
R18429 gnd.n7684 gnd.n191 9.3005
R18430 gnd.n7683 gnd.n192 9.3005
R18431 gnd.n207 gnd.n193 9.3005
R18432 gnd.n7673 gnd.n208 9.3005
R18433 gnd.n7672 gnd.n209 9.3005
R18434 gnd.n7671 gnd.n210 9.3005
R18435 gnd.n227 gnd.n211 9.3005
R18436 gnd.n7661 gnd.n228 9.3005
R18437 gnd.n7660 gnd.n229 9.3005
R18438 gnd.n7659 gnd.n230 9.3005
R18439 gnd.n245 gnd.n231 9.3005
R18440 gnd.n7649 gnd.n246 9.3005
R18441 gnd.n7648 gnd.n247 9.3005
R18442 gnd.n7647 gnd.n248 9.3005
R18443 gnd.n7739 gnd.n7738 9.3005
R18444 gnd.n7737 gnd.n101 9.3005
R18445 gnd.n7344 gnd.n103 9.3005
R18446 gnd.n7346 gnd.n7345 9.3005
R18447 gnd.n7347 gnd.n7343 9.3005
R18448 gnd.n7349 gnd.n7348 9.3005
R18449 gnd.n7351 gnd.n7341 9.3005
R18450 gnd.n7353 gnd.n7352 9.3005
R18451 gnd.n7354 gnd.n7340 9.3005
R18452 gnd.n7356 gnd.n7355 9.3005
R18453 gnd.n7358 gnd.n7338 9.3005
R18454 gnd.n7360 gnd.n7359 9.3005
R18455 gnd.n7361 gnd.n7337 9.3005
R18456 gnd.n7363 gnd.n7362 9.3005
R18457 gnd.n7365 gnd.n7335 9.3005
R18458 gnd.n7367 gnd.n7366 9.3005
R18459 gnd.n7368 gnd.n7334 9.3005
R18460 gnd.n7370 gnd.n7369 9.3005
R18461 gnd.n7372 gnd.n7332 9.3005
R18462 gnd.n7374 gnd.n7373 9.3005
R18463 gnd.n7375 gnd.n7331 9.3005
R18464 gnd.n7377 gnd.n7376 9.3005
R18465 gnd.n7379 gnd.n7329 9.3005
R18466 gnd.n7381 gnd.n7380 9.3005
R18467 gnd.n7382 gnd.n7328 9.3005
R18468 gnd.n7384 gnd.n7383 9.3005
R18469 gnd.n7386 gnd.n7326 9.3005
R18470 gnd.n7388 gnd.n7387 9.3005
R18471 gnd.n7389 gnd.n7325 9.3005
R18472 gnd.n7391 gnd.n7390 9.3005
R18473 gnd.n7393 gnd.n7323 9.3005
R18474 gnd.n7395 gnd.n7394 9.3005
R18475 gnd.n7426 gnd.n7289 9.3005
R18476 gnd.n7425 gnd.n7291 9.3005
R18477 gnd.n7295 gnd.n7292 9.3005
R18478 gnd.n7420 gnd.n7296 9.3005
R18479 gnd.n7419 gnd.n7297 9.3005
R18480 gnd.n7418 gnd.n7298 9.3005
R18481 gnd.n7302 gnd.n7299 9.3005
R18482 gnd.n7413 gnd.n7303 9.3005
R18483 gnd.n7412 gnd.n7304 9.3005
R18484 gnd.n7411 gnd.n7305 9.3005
R18485 gnd.n7309 gnd.n7306 9.3005
R18486 gnd.n7406 gnd.n7310 9.3005
R18487 gnd.n7405 gnd.n7311 9.3005
R18488 gnd.n7404 gnd.n7312 9.3005
R18489 gnd.n7316 gnd.n7313 9.3005
R18490 gnd.n7399 gnd.n7317 9.3005
R18491 gnd.n7398 gnd.n7397 9.3005
R18492 gnd.n7396 gnd.n7320 9.3005
R18493 gnd.n7428 gnd.n7427 9.3005
R18494 gnd.n7494 gnd.n7491 9.3005
R18495 gnd.n7500 gnd.n7499 9.3005
R18496 gnd.n7501 gnd.n7490 9.3005
R18497 gnd.n7503 gnd.n7502 9.3005
R18498 gnd.n7488 gnd.n7487 9.3005
R18499 gnd.n7510 gnd.n7509 9.3005
R18500 gnd.n7511 gnd.n7486 9.3005
R18501 gnd.n7513 gnd.n7512 9.3005
R18502 gnd.n7484 gnd.n7483 9.3005
R18503 gnd.n7520 gnd.n7519 9.3005
R18504 gnd.n7521 gnd.n7482 9.3005
R18505 gnd.n7523 gnd.n7522 9.3005
R18506 gnd.n7480 gnd.n7479 9.3005
R18507 gnd.n7531 gnd.n7530 9.3005
R18508 gnd.n7532 gnd.n7478 9.3005
R18509 gnd.n7534 gnd.n7533 9.3005
R18510 gnd.n7535 gnd.n7473 9.3005
R18511 gnd.n7541 gnd.n7540 9.3005
R18512 gnd.n7542 gnd.n7472 9.3005
R18513 gnd.n7544 gnd.n7543 9.3005
R18514 gnd.n7470 gnd.n7469 9.3005
R18515 gnd.n7551 gnd.n7550 9.3005
R18516 gnd.n7552 gnd.n7468 9.3005
R18517 gnd.n7554 gnd.n7553 9.3005
R18518 gnd.n7466 gnd.n7465 9.3005
R18519 gnd.n7561 gnd.n7560 9.3005
R18520 gnd.n7562 gnd.n7464 9.3005
R18521 gnd.n7564 gnd.n7563 9.3005
R18522 gnd.n7462 gnd.n7461 9.3005
R18523 gnd.n7571 gnd.n7570 9.3005
R18524 gnd.n7572 gnd.n7460 9.3005
R18525 gnd.n7574 gnd.n7573 9.3005
R18526 gnd.n7458 gnd.n7457 9.3005
R18527 gnd.n7581 gnd.n7580 9.3005
R18528 gnd.n7582 gnd.n7456 9.3005
R18529 gnd.n7584 gnd.n7583 9.3005
R18530 gnd.n7454 gnd.n7451 9.3005
R18531 gnd.n7591 gnd.n7590 9.3005
R18532 gnd.n7592 gnd.n7450 9.3005
R18533 gnd.n7594 gnd.n7593 9.3005
R18534 gnd.n7448 gnd.n7447 9.3005
R18535 gnd.n7601 gnd.n7600 9.3005
R18536 gnd.n7602 gnd.n7446 9.3005
R18537 gnd.n7604 gnd.n7603 9.3005
R18538 gnd.n7444 gnd.n7443 9.3005
R18539 gnd.n7611 gnd.n7610 9.3005
R18540 gnd.n7612 gnd.n7442 9.3005
R18541 gnd.n7614 gnd.n7613 9.3005
R18542 gnd.n7440 gnd.n7439 9.3005
R18543 gnd.n7621 gnd.n7620 9.3005
R18544 gnd.n7622 gnd.n7438 9.3005
R18545 gnd.n7624 gnd.n7623 9.3005
R18546 gnd.n7436 gnd.n7435 9.3005
R18547 gnd.n7631 gnd.n7630 9.3005
R18548 gnd.n7632 gnd.n7434 9.3005
R18549 gnd.n7634 gnd.n7633 9.3005
R18550 gnd.n7432 gnd.n7429 9.3005
R18551 gnd.n7640 gnd.n7639 9.3005
R18552 gnd.n7493 gnd.n7492 9.3005
R18553 gnd.n5954 gnd.n5953 9.3005
R18554 gnd.n5961 gnd.n5958 9.3005
R18555 gnd.n5962 gnd.n5951 9.3005
R18556 gnd.n5985 gnd.n5963 9.3005
R18557 gnd.n5984 gnd.n5983 9.3005
R18558 gnd.n399 gnd.n397 9.3005
R18559 gnd.n7040 gnd.n398 9.3005
R18560 gnd.n7042 gnd.n7041 9.3005
R18561 gnd.n7043 gnd.n371 9.3005
R18562 gnd.n7072 gnd.n372 9.3005
R18563 gnd.n7073 gnd.n369 9.3005
R18564 gnd.n7076 gnd.n370 9.3005
R18565 gnd.n7078 gnd.n7077 9.3005
R18566 gnd.n7079 gnd.n343 9.3005
R18567 gnd.n7128 gnd.n344 9.3005
R18568 gnd.n7129 gnd.n342 9.3005
R18569 gnd.n7131 gnd.n7130 9.3005
R18570 gnd.n7132 gnd.n325 9.3005
R18571 gnd.n7148 gnd.n326 9.3005
R18572 gnd.n7149 gnd.n324 9.3005
R18573 gnd.n7151 gnd.n7150 9.3005
R18574 gnd.n7152 gnd.n307 9.3005
R18575 gnd.n7168 gnd.n308 9.3005
R18576 gnd.n7169 gnd.n305 9.3005
R18577 gnd.n7171 gnd.n306 9.3005
R18578 gnd.n7173 gnd.n7172 9.3005
R18579 gnd.n7174 gnd.n281 9.3005
R18580 gnd.n7206 gnd.n280 9.3005
R18581 gnd.n7210 gnd.n7209 9.3005
R18582 gnd.n7208 gnd.n263 9.3005
R18583 gnd.n7227 gnd.n262 9.3005
R18584 gnd.n7229 gnd.n7228 9.3005
R18585 gnd.n7230 gnd.n257 9.3005
R18586 gnd.n7236 gnd.n256 9.3005
R18587 gnd.n7239 gnd.n7237 9.3005
R18588 gnd.n7240 gnd.n122 9.3005
R18589 gnd.n7242 gnd.n123 9.3005
R18590 gnd.n7243 gnd.n124 9.3005
R18591 gnd.n7246 gnd.n7244 9.3005
R18592 gnd.n7247 gnd.n141 9.3005
R18593 gnd.n7249 gnd.n142 9.3005
R18594 gnd.n7250 gnd.n143 9.3005
R18595 gnd.n7253 gnd.n7251 9.3005
R18596 gnd.n7254 gnd.n160 9.3005
R18597 gnd.n7256 gnd.n161 9.3005
R18598 gnd.n7257 gnd.n162 9.3005
R18599 gnd.n7260 gnd.n7258 9.3005
R18600 gnd.n7261 gnd.n180 9.3005
R18601 gnd.n7263 gnd.n181 9.3005
R18602 gnd.n7264 gnd.n182 9.3005
R18603 gnd.n7267 gnd.n7265 9.3005
R18604 gnd.n7268 gnd.n199 9.3005
R18605 gnd.n7270 gnd.n200 9.3005
R18606 gnd.n7271 gnd.n201 9.3005
R18607 gnd.n7274 gnd.n7272 9.3005
R18608 gnd.n7275 gnd.n218 9.3005
R18609 gnd.n7277 gnd.n219 9.3005
R18610 gnd.n7278 gnd.n220 9.3005
R18611 gnd.n7281 gnd.n7279 9.3005
R18612 gnd.n7282 gnd.n237 9.3005
R18613 gnd.n7284 gnd.n238 9.3005
R18614 gnd.n7285 gnd.n239 9.3005
R18615 gnd.n7287 gnd.n255 9.3005
R18616 gnd.n7642 gnd.n7288 9.3005
R18617 gnd.n5952 gnd.n1138 9.3005
R18618 gnd.n5955 gnd.n5954 9.3005
R18619 gnd.n5958 gnd.n5957 9.3005
R18620 gnd.n5951 gnd.n5950 9.3005
R18621 gnd.n5986 gnd.n5985 9.3005
R18622 gnd.n5984 gnd.n396 9.3005
R18623 gnd.n7049 gnd.n397 9.3005
R18624 gnd.n7048 gnd.n398 9.3005
R18625 gnd.n7047 gnd.n7042 9.3005
R18626 gnd.n7046 gnd.n7043 9.3005
R18627 gnd.n372 gnd.n368 9.3005
R18628 gnd.n7085 gnd.n369 9.3005
R18629 gnd.n7084 gnd.n370 9.3005
R18630 gnd.n7083 gnd.n7078 9.3005
R18631 gnd.n7082 gnd.n7079 9.3005
R18632 gnd.n344 gnd.n341 9.3005
R18633 gnd.n7135 gnd.n342 9.3005
R18634 gnd.n7134 gnd.n7131 9.3005
R18635 gnd.n7133 gnd.n7132 9.3005
R18636 gnd.n326 gnd.n323 9.3005
R18637 gnd.n7155 gnd.n324 9.3005
R18638 gnd.n7154 gnd.n7151 9.3005
R18639 gnd.n7153 gnd.n7152 9.3005
R18640 gnd.n308 gnd.n304 9.3005
R18641 gnd.n7179 gnd.n305 9.3005
R18642 gnd.n7178 gnd.n306 9.3005
R18643 gnd.n7177 gnd.n7173 9.3005
R18644 gnd.n7176 gnd.n7174 9.3005
R18645 gnd.n280 gnd.n279 9.3005
R18646 gnd.n7211 gnd.n7210 9.3005
R18647 gnd.n264 gnd.n263 9.3005
R18648 gnd.n7227 gnd.n7226 9.3005
R18649 gnd.n7228 gnd.n258 9.3005
R18650 gnd.n7234 gnd.n257 9.3005
R18651 gnd.n7236 gnd.n7235 9.3005
R18652 gnd.n7237 gnd.n121 9.3005
R18653 gnd.n7727 gnd.n122 9.3005
R18654 gnd.n7726 gnd.n123 9.3005
R18655 gnd.n7725 gnd.n124 9.3005
R18656 gnd.n7244 gnd.n125 9.3005
R18657 gnd.n7715 gnd.n141 9.3005
R18658 gnd.n7714 gnd.n142 9.3005
R18659 gnd.n7713 gnd.n143 9.3005
R18660 gnd.n7251 gnd.n144 9.3005
R18661 gnd.n7703 gnd.n160 9.3005
R18662 gnd.n7702 gnd.n161 9.3005
R18663 gnd.n7701 gnd.n162 9.3005
R18664 gnd.n7258 gnd.n163 9.3005
R18665 gnd.n7691 gnd.n180 9.3005
R18666 gnd.n7690 gnd.n181 9.3005
R18667 gnd.n7689 gnd.n182 9.3005
R18668 gnd.n7265 gnd.n183 9.3005
R18669 gnd.n7679 gnd.n199 9.3005
R18670 gnd.n7678 gnd.n200 9.3005
R18671 gnd.n7677 gnd.n201 9.3005
R18672 gnd.n7272 gnd.n202 9.3005
R18673 gnd.n7667 gnd.n218 9.3005
R18674 gnd.n7666 gnd.n219 9.3005
R18675 gnd.n7665 gnd.n220 9.3005
R18676 gnd.n7279 gnd.n221 9.3005
R18677 gnd.n7655 gnd.n237 9.3005
R18678 gnd.n7654 gnd.n238 9.3005
R18679 gnd.n7653 gnd.n239 9.3005
R18680 gnd.n255 gnd.n240 9.3005
R18681 gnd.n7643 gnd.n7642 9.3005
R18682 gnd.n1150 gnd.n1138 9.3005
R18683 gnd.n6457 gnd.n6456 9.3005
R18684 gnd.n6458 gnd.n749 9.3005
R18685 gnd.n6460 gnd.n6459 9.3005
R18686 gnd.n745 gnd.n744 9.3005
R18687 gnd.n6467 gnd.n6466 9.3005
R18688 gnd.n6468 gnd.n743 9.3005
R18689 gnd.n6470 gnd.n6469 9.3005
R18690 gnd.n739 gnd.n738 9.3005
R18691 gnd.n6477 gnd.n6476 9.3005
R18692 gnd.n6478 gnd.n737 9.3005
R18693 gnd.n6480 gnd.n6479 9.3005
R18694 gnd.n733 gnd.n732 9.3005
R18695 gnd.n6487 gnd.n6486 9.3005
R18696 gnd.n6488 gnd.n731 9.3005
R18697 gnd.n6490 gnd.n6489 9.3005
R18698 gnd.n727 gnd.n726 9.3005
R18699 gnd.n6497 gnd.n6496 9.3005
R18700 gnd.n6498 gnd.n725 9.3005
R18701 gnd.n6500 gnd.n6499 9.3005
R18702 gnd.n721 gnd.n720 9.3005
R18703 gnd.n6507 gnd.n6506 9.3005
R18704 gnd.n6508 gnd.n719 9.3005
R18705 gnd.n6510 gnd.n6509 9.3005
R18706 gnd.n715 gnd.n714 9.3005
R18707 gnd.n6517 gnd.n6516 9.3005
R18708 gnd.n6518 gnd.n713 9.3005
R18709 gnd.n6520 gnd.n6519 9.3005
R18710 gnd.n709 gnd.n708 9.3005
R18711 gnd.n6527 gnd.n6526 9.3005
R18712 gnd.n6528 gnd.n707 9.3005
R18713 gnd.n6530 gnd.n6529 9.3005
R18714 gnd.n703 gnd.n702 9.3005
R18715 gnd.n6537 gnd.n6536 9.3005
R18716 gnd.n6538 gnd.n701 9.3005
R18717 gnd.n6540 gnd.n6539 9.3005
R18718 gnd.n697 gnd.n696 9.3005
R18719 gnd.n6547 gnd.n6546 9.3005
R18720 gnd.n6548 gnd.n695 9.3005
R18721 gnd.n6550 gnd.n6549 9.3005
R18722 gnd.n691 gnd.n690 9.3005
R18723 gnd.n6557 gnd.n6556 9.3005
R18724 gnd.n6558 gnd.n689 9.3005
R18725 gnd.n6560 gnd.n6559 9.3005
R18726 gnd.n685 gnd.n684 9.3005
R18727 gnd.n6567 gnd.n6566 9.3005
R18728 gnd.n6568 gnd.n683 9.3005
R18729 gnd.n6570 gnd.n6569 9.3005
R18730 gnd.n679 gnd.n678 9.3005
R18731 gnd.n6577 gnd.n6576 9.3005
R18732 gnd.n6578 gnd.n677 9.3005
R18733 gnd.n6580 gnd.n6579 9.3005
R18734 gnd.n673 gnd.n672 9.3005
R18735 gnd.n6587 gnd.n6586 9.3005
R18736 gnd.n6588 gnd.n671 9.3005
R18737 gnd.n6590 gnd.n6589 9.3005
R18738 gnd.n667 gnd.n666 9.3005
R18739 gnd.n6597 gnd.n6596 9.3005
R18740 gnd.n6598 gnd.n665 9.3005
R18741 gnd.n6600 gnd.n6599 9.3005
R18742 gnd.n661 gnd.n660 9.3005
R18743 gnd.n6607 gnd.n6606 9.3005
R18744 gnd.n6608 gnd.n659 9.3005
R18745 gnd.n6610 gnd.n6609 9.3005
R18746 gnd.n655 gnd.n654 9.3005
R18747 gnd.n6617 gnd.n6616 9.3005
R18748 gnd.n6618 gnd.n653 9.3005
R18749 gnd.n6620 gnd.n6619 9.3005
R18750 gnd.n649 gnd.n648 9.3005
R18751 gnd.n6627 gnd.n6626 9.3005
R18752 gnd.n6628 gnd.n647 9.3005
R18753 gnd.n6630 gnd.n6629 9.3005
R18754 gnd.n643 gnd.n642 9.3005
R18755 gnd.n6637 gnd.n6636 9.3005
R18756 gnd.n6638 gnd.n641 9.3005
R18757 gnd.n6640 gnd.n6639 9.3005
R18758 gnd.n637 gnd.n636 9.3005
R18759 gnd.n6647 gnd.n6646 9.3005
R18760 gnd.n6648 gnd.n635 9.3005
R18761 gnd.n6650 gnd.n6649 9.3005
R18762 gnd.n631 gnd.n630 9.3005
R18763 gnd.n6657 gnd.n6656 9.3005
R18764 gnd.n6658 gnd.n629 9.3005
R18765 gnd.n6660 gnd.n6659 9.3005
R18766 gnd.n625 gnd.n624 9.3005
R18767 gnd.n6667 gnd.n6666 9.3005
R18768 gnd.n6668 gnd.n623 9.3005
R18769 gnd.n6670 gnd.n6669 9.3005
R18770 gnd.n619 gnd.n618 9.3005
R18771 gnd.n6677 gnd.n6676 9.3005
R18772 gnd.n6678 gnd.n617 9.3005
R18773 gnd.n6680 gnd.n6679 9.3005
R18774 gnd.n613 gnd.n612 9.3005
R18775 gnd.n6687 gnd.n6686 9.3005
R18776 gnd.n6688 gnd.n611 9.3005
R18777 gnd.n6690 gnd.n6689 9.3005
R18778 gnd.n607 gnd.n606 9.3005
R18779 gnd.n6697 gnd.n6696 9.3005
R18780 gnd.n6698 gnd.n605 9.3005
R18781 gnd.n6700 gnd.n6699 9.3005
R18782 gnd.n601 gnd.n600 9.3005
R18783 gnd.n6707 gnd.n6706 9.3005
R18784 gnd.n6708 gnd.n599 9.3005
R18785 gnd.n6710 gnd.n6709 9.3005
R18786 gnd.n595 gnd.n594 9.3005
R18787 gnd.n6717 gnd.n6716 9.3005
R18788 gnd.n6718 gnd.n593 9.3005
R18789 gnd.n6720 gnd.n6719 9.3005
R18790 gnd.n589 gnd.n588 9.3005
R18791 gnd.n6727 gnd.n6726 9.3005
R18792 gnd.n6728 gnd.n587 9.3005
R18793 gnd.n6730 gnd.n6729 9.3005
R18794 gnd.n583 gnd.n582 9.3005
R18795 gnd.n6737 gnd.n6736 9.3005
R18796 gnd.n6738 gnd.n581 9.3005
R18797 gnd.n6740 gnd.n6739 9.3005
R18798 gnd.n577 gnd.n576 9.3005
R18799 gnd.n6747 gnd.n6746 9.3005
R18800 gnd.n6748 gnd.n575 9.3005
R18801 gnd.n6750 gnd.n6749 9.3005
R18802 gnd.n571 gnd.n570 9.3005
R18803 gnd.n6757 gnd.n6756 9.3005
R18804 gnd.n6758 gnd.n569 9.3005
R18805 gnd.n6760 gnd.n6759 9.3005
R18806 gnd.n565 gnd.n564 9.3005
R18807 gnd.n6767 gnd.n6766 9.3005
R18808 gnd.n6768 gnd.n563 9.3005
R18809 gnd.n6770 gnd.n6769 9.3005
R18810 gnd.n559 gnd.n558 9.3005
R18811 gnd.n6777 gnd.n6776 9.3005
R18812 gnd.n6778 gnd.n557 9.3005
R18813 gnd.n6780 gnd.n6779 9.3005
R18814 gnd.n553 gnd.n552 9.3005
R18815 gnd.n6787 gnd.n6786 9.3005
R18816 gnd.n6788 gnd.n551 9.3005
R18817 gnd.n6790 gnd.n6789 9.3005
R18818 gnd.n547 gnd.n546 9.3005
R18819 gnd.n6797 gnd.n6796 9.3005
R18820 gnd.n6798 gnd.n545 9.3005
R18821 gnd.n6801 gnd.n6800 9.3005
R18822 gnd.n6799 gnd.n541 9.3005
R18823 gnd.n6807 gnd.n540 9.3005
R18824 gnd.n6809 gnd.n6808 9.3005
R18825 gnd.n536 gnd.n535 9.3005
R18826 gnd.n6818 gnd.n6817 9.3005
R18827 gnd.n6819 gnd.n534 9.3005
R18828 gnd.n6821 gnd.n6820 9.3005
R18829 gnd.n530 gnd.n529 9.3005
R18830 gnd.n6828 gnd.n6827 9.3005
R18831 gnd.n6829 gnd.n528 9.3005
R18832 gnd.n6831 gnd.n6830 9.3005
R18833 gnd.n524 gnd.n523 9.3005
R18834 gnd.n6838 gnd.n6837 9.3005
R18835 gnd.n6839 gnd.n522 9.3005
R18836 gnd.n6841 gnd.n6840 9.3005
R18837 gnd.n518 gnd.n517 9.3005
R18838 gnd.n6848 gnd.n6847 9.3005
R18839 gnd.n6849 gnd.n516 9.3005
R18840 gnd.n6851 gnd.n6850 9.3005
R18841 gnd.n512 gnd.n511 9.3005
R18842 gnd.n6858 gnd.n6857 9.3005
R18843 gnd.n6859 gnd.n510 9.3005
R18844 gnd.n6861 gnd.n6860 9.3005
R18845 gnd.n506 gnd.n505 9.3005
R18846 gnd.n6868 gnd.n6867 9.3005
R18847 gnd.n6869 gnd.n504 9.3005
R18848 gnd.n6871 gnd.n6870 9.3005
R18849 gnd.n500 gnd.n499 9.3005
R18850 gnd.n6878 gnd.n6877 9.3005
R18851 gnd.n6879 gnd.n498 9.3005
R18852 gnd.n6881 gnd.n6880 9.3005
R18853 gnd.n494 gnd.n493 9.3005
R18854 gnd.n6888 gnd.n6887 9.3005
R18855 gnd.n6889 gnd.n492 9.3005
R18856 gnd.n6891 gnd.n6890 9.3005
R18857 gnd.n488 gnd.n487 9.3005
R18858 gnd.n6898 gnd.n6897 9.3005
R18859 gnd.n6899 gnd.n486 9.3005
R18860 gnd.n6901 gnd.n6900 9.3005
R18861 gnd.n482 gnd.n481 9.3005
R18862 gnd.n6908 gnd.n6907 9.3005
R18863 gnd.n6909 gnd.n480 9.3005
R18864 gnd.n6911 gnd.n6910 9.3005
R18865 gnd.n476 gnd.n475 9.3005
R18866 gnd.n6918 gnd.n6917 9.3005
R18867 gnd.n6919 gnd.n474 9.3005
R18868 gnd.n6921 gnd.n6920 9.3005
R18869 gnd.n470 gnd.n469 9.3005
R18870 gnd.n6928 gnd.n6927 9.3005
R18871 gnd.n6929 gnd.n468 9.3005
R18872 gnd.n6931 gnd.n6930 9.3005
R18873 gnd.n464 gnd.n463 9.3005
R18874 gnd.n6938 gnd.n6937 9.3005
R18875 gnd.n6939 gnd.n462 9.3005
R18876 gnd.n6941 gnd.n6940 9.3005
R18877 gnd.n458 gnd.n457 9.3005
R18878 gnd.n6948 gnd.n6947 9.3005
R18879 gnd.n6949 gnd.n456 9.3005
R18880 gnd.n6951 gnd.n6950 9.3005
R18881 gnd.n452 gnd.n451 9.3005
R18882 gnd.n6958 gnd.n6957 9.3005
R18883 gnd.n6959 gnd.n450 9.3005
R18884 gnd.n6961 gnd.n6960 9.3005
R18885 gnd.n446 gnd.n445 9.3005
R18886 gnd.n6968 gnd.n6967 9.3005
R18887 gnd.n6969 gnd.n444 9.3005
R18888 gnd.n6971 gnd.n6970 9.3005
R18889 gnd.n440 gnd.n439 9.3005
R18890 gnd.n6978 gnd.n6977 9.3005
R18891 gnd.n6979 gnd.n438 9.3005
R18892 gnd.n6981 gnd.n6980 9.3005
R18893 gnd.n434 gnd.n433 9.3005
R18894 gnd.n6988 gnd.n6987 9.3005
R18895 gnd.n6989 gnd.n432 9.3005
R18896 gnd.n6991 gnd.n6990 9.3005
R18897 gnd.n428 gnd.n427 9.3005
R18898 gnd.n6998 gnd.n6997 9.3005
R18899 gnd.n6999 gnd.n426 9.3005
R18900 gnd.n7001 gnd.n7000 9.3005
R18901 gnd.n422 gnd.n421 9.3005
R18902 gnd.n7008 gnd.n7007 9.3005
R18903 gnd.n7009 gnd.n420 9.3005
R18904 gnd.n7011 gnd.n7010 9.3005
R18905 gnd.n416 gnd.n415 9.3005
R18906 gnd.n7019 gnd.n7018 9.3005
R18907 gnd.n7020 gnd.n414 9.3005
R18908 gnd.n7023 gnd.n7022 9.3005
R18909 gnd.n6811 gnd.n6810 9.3005
R18910 gnd.n4570 gnd.n4569 9.3005
R18911 gnd.n4872 gnd.n4871 9.3005
R18912 gnd.n4873 gnd.n4568 9.3005
R18913 gnd.n4899 gnd.n4874 9.3005
R18914 gnd.n4898 gnd.n4875 9.3005
R18915 gnd.n4897 gnd.n4876 9.3005
R18916 gnd.n4879 gnd.n4877 9.3005
R18917 gnd.n4893 gnd.n4880 9.3005
R18918 gnd.n4892 gnd.n4881 9.3005
R18919 gnd.n4891 gnd.n4882 9.3005
R18920 gnd.n4884 gnd.n4883 9.3005
R18921 gnd.n4887 gnd.n4886 9.3005
R18922 gnd.n4885 gnd.n846 9.3005
R18923 gnd.n6397 gnd.n847 9.3005
R18924 gnd.n6396 gnd.n848 9.3005
R18925 gnd.n6395 gnd.n849 9.3005
R18926 gnd.n855 gnd.n850 9.3005
R18927 gnd.n6389 gnd.n856 9.3005
R18928 gnd.n6388 gnd.n857 9.3005
R18929 gnd.n6387 gnd.n858 9.3005
R18930 gnd.n5018 gnd.n859 9.3005
R18931 gnd.n5019 gnd.n5017 9.3005
R18932 gnd.n5021 gnd.n5020 9.3005
R18933 gnd.n2059 gnd.n2058 9.3005
R18934 gnd.n5036 gnd.n5035 9.3005
R18935 gnd.n5037 gnd.n2057 9.3005
R18936 gnd.n5039 gnd.n5038 9.3005
R18937 gnd.n2048 gnd.n2047 9.3005
R18938 gnd.n5053 gnd.n5052 9.3005
R18939 gnd.n5054 gnd.n2046 9.3005
R18940 gnd.n5056 gnd.n5055 9.3005
R18941 gnd.n2036 gnd.n2035 9.3005
R18942 gnd.n5070 gnd.n5069 9.3005
R18943 gnd.n5071 gnd.n2034 9.3005
R18944 gnd.n5075 gnd.n5072 9.3005
R18945 gnd.n5074 gnd.n5073 9.3005
R18946 gnd.n1626 gnd.n1625 9.3005
R18947 gnd.n5163 gnd.n5162 9.3005
R18948 gnd.n5164 gnd.n1624 9.3005
R18949 gnd.n5177 gnd.n5165 9.3005
R18950 gnd.n5176 gnd.n5166 9.3005
R18951 gnd.n5175 gnd.n5167 9.3005
R18952 gnd.n5169 gnd.n5168 9.3005
R18953 gnd.n5171 gnd.n5170 9.3005
R18954 gnd.n1587 gnd.n1586 9.3005
R18955 gnd.n5222 gnd.n5221 9.3005
R18956 gnd.n5223 gnd.n1585 9.3005
R18957 gnd.n5225 gnd.n5224 9.3005
R18958 gnd.n1565 gnd.n1564 9.3005
R18959 gnd.n5252 gnd.n5251 9.3005
R18960 gnd.n5253 gnd.n1563 9.3005
R18961 gnd.n5255 gnd.n5254 9.3005
R18962 gnd.n1548 gnd.n1547 9.3005
R18963 gnd.n5279 gnd.n5278 9.3005
R18964 gnd.n5280 gnd.n1546 9.3005
R18965 gnd.n5282 gnd.n5281 9.3005
R18966 gnd.n1528 gnd.n1527 9.3005
R18967 gnd.n5303 gnd.n5302 9.3005
R18968 gnd.n5304 gnd.n1526 9.3005
R18969 gnd.n5308 gnd.n5305 9.3005
R18970 gnd.n5307 gnd.n5306 9.3005
R18971 gnd.n1501 gnd.n1500 9.3005
R18972 gnd.n5361 gnd.n5360 9.3005
R18973 gnd.n5362 gnd.n1499 9.3005
R18974 gnd.n5366 gnd.n5363 9.3005
R18975 gnd.n5365 gnd.n5364 9.3005
R18976 gnd.n1479 gnd.n1478 9.3005
R18977 gnd.n5401 gnd.n5400 9.3005
R18978 gnd.n5402 gnd.n1477 9.3005
R18979 gnd.n5406 gnd.n5403 9.3005
R18980 gnd.n5405 gnd.n5404 9.3005
R18981 gnd.n1450 gnd.n1449 9.3005
R18982 gnd.n5458 gnd.n5457 9.3005
R18983 gnd.n5459 gnd.n1448 9.3005
R18984 gnd.n5463 gnd.n5460 9.3005
R18985 gnd.n5462 gnd.n5461 9.3005
R18986 gnd.n1429 gnd.n1428 9.3005
R18987 gnd.n5496 gnd.n5495 9.3005
R18988 gnd.n5497 gnd.n1427 9.3005
R18989 gnd.n5499 gnd.n5498 9.3005
R18990 gnd.n1400 gnd.n1399 9.3005
R18991 gnd.n5534 gnd.n5533 9.3005
R18992 gnd.n5535 gnd.n1398 9.3005
R18993 gnd.n5539 gnd.n5536 9.3005
R18994 gnd.n5538 gnd.n5537 9.3005
R18995 gnd.n1374 gnd.n1373 9.3005
R18996 gnd.n5578 gnd.n5577 9.3005
R18997 gnd.n5579 gnd.n1372 9.3005
R18998 gnd.n5582 gnd.n5581 9.3005
R18999 gnd.n5580 gnd.n1351 9.3005
R19000 gnd.n5618 gnd.n1352 9.3005
R19001 gnd.n5617 gnd.n1353 9.3005
R19002 gnd.n5616 gnd.n1354 9.3005
R19003 gnd.n1356 gnd.n1355 9.3005
R19004 gnd.n1358 gnd.n1357 9.3005
R19005 gnd.n1319 gnd.n1318 9.3005
R19006 gnd.n5665 gnd.n5664 9.3005
R19007 gnd.n5666 gnd.n1317 9.3005
R19008 gnd.n5668 gnd.n5667 9.3005
R19009 gnd.n1224 gnd.n1223 9.3005
R19010 gnd.n5813 gnd.n5812 9.3005
R19011 gnd.n5814 gnd.n1222 9.3005
R19012 gnd.n5816 gnd.n5815 9.3005
R19013 gnd.n1212 gnd.n1211 9.3005
R19014 gnd.n5830 gnd.n5829 9.3005
R19015 gnd.n5831 gnd.n1210 9.3005
R19016 gnd.n5833 gnd.n5832 9.3005
R19017 gnd.n1200 gnd.n1199 9.3005
R19018 gnd.n5847 gnd.n5846 9.3005
R19019 gnd.n5848 gnd.n1198 9.3005
R19020 gnd.n5850 gnd.n5849 9.3005
R19021 gnd.n1188 gnd.n1187 9.3005
R19022 gnd.n5865 gnd.n5864 9.3005
R19023 gnd.n5866 gnd.n1186 9.3005
R19024 gnd.n5868 gnd.n5867 9.3005
R19025 gnd.n1177 gnd.n1176 9.3005
R19026 gnd.n5882 gnd.n5881 9.3005
R19027 gnd.n5883 gnd.n1175 9.3005
R19028 gnd.n5887 gnd.n5884 9.3005
R19029 gnd.n5886 gnd.n5885 9.3005
R19030 gnd.n1164 gnd.n1163 9.3005
R19031 gnd.n5919 gnd.n5918 9.3005
R19032 gnd.n5920 gnd.n1162 9.3005
R19033 gnd.n5922 gnd.n5921 9.3005
R19034 gnd.n1160 gnd.n1159 9.3005
R19035 gnd.n5928 gnd.n5927 9.3005
R19036 gnd.n5929 gnd.n1158 9.3005
R19037 gnd.n6007 gnd.n5930 9.3005
R19038 gnd.n6006 gnd.n5931 9.3005
R19039 gnd.n6005 gnd.n5932 9.3005
R19040 gnd.n5944 gnd.n5933 9.3005
R19041 gnd.n5947 gnd.n5946 9.3005
R19042 gnd.n5945 gnd.n402 9.3005
R19043 gnd.n7035 gnd.n403 9.3005
R19044 gnd.n7034 gnd.n404 9.3005
R19045 gnd.n7033 gnd.n405 9.3005
R19046 gnd.n408 gnd.n406 9.3005
R19047 gnd.n7029 gnd.n409 9.3005
R19048 gnd.n7028 gnd.n410 9.3005
R19049 gnd.n7027 gnd.n411 9.3005
R19050 gnd.n7021 gnd.n412 9.3005
R19051 gnd.n4867 gnd.n4866 9.3005
R19052 gnd.n4863 gnd.n4572 9.3005
R19053 gnd.n4855 gnd.n4573 9.3005
R19054 gnd.n4857 gnd.n4856 9.3005
R19055 gnd.n4854 gnd.n4575 9.3005
R19056 gnd.n4853 gnd.n4852 9.3005
R19057 gnd.n4577 gnd.n4576 9.3005
R19058 gnd.n4846 gnd.n4845 9.3005
R19059 gnd.n4844 gnd.n4579 9.3005
R19060 gnd.n4843 gnd.n4842 9.3005
R19061 gnd.n4581 gnd.n4580 9.3005
R19062 gnd.n4836 gnd.n4835 9.3005
R19063 gnd.n4834 gnd.n4583 9.3005
R19064 gnd.n4833 gnd.n4832 9.3005
R19065 gnd.n4585 gnd.n4584 9.3005
R19066 gnd.n4826 gnd.n4825 9.3005
R19067 gnd.n4824 gnd.n4587 9.3005
R19068 gnd.n4823 gnd.n4822 9.3005
R19069 gnd.n4589 gnd.n4588 9.3005
R19070 gnd.n4816 gnd.n4815 9.3005
R19071 gnd.n4814 gnd.n4591 9.3005
R19072 gnd.n4813 gnd.n4812 9.3005
R19073 gnd.n4593 gnd.n4592 9.3005
R19074 gnd.n4806 gnd.n4805 9.3005
R19075 gnd.n4804 gnd.n4595 9.3005
R19076 gnd.n4803 gnd.n4802 9.3005
R19077 gnd.n4597 gnd.n4596 9.3005
R19078 gnd.n4796 gnd.n4795 9.3005
R19079 gnd.n4794 gnd.n4599 9.3005
R19080 gnd.n4793 gnd.n4792 9.3005
R19081 gnd.n4601 gnd.n4600 9.3005
R19082 gnd.n4786 gnd.n4785 9.3005
R19083 gnd.n4784 gnd.n4603 9.3005
R19084 gnd.n4783 gnd.n4782 9.3005
R19085 gnd.n4605 gnd.n4604 9.3005
R19086 gnd.n4776 gnd.n4775 9.3005
R19087 gnd.n4774 gnd.n4607 9.3005
R19088 gnd.n4773 gnd.n4772 9.3005
R19089 gnd.n4609 gnd.n4608 9.3005
R19090 gnd.n4766 gnd.n4765 9.3005
R19091 gnd.n4764 gnd.n4611 9.3005
R19092 gnd.n4763 gnd.n4762 9.3005
R19093 gnd.n4613 gnd.n4612 9.3005
R19094 gnd.n4756 gnd.n4755 9.3005
R19095 gnd.n4754 gnd.n4615 9.3005
R19096 gnd.n4753 gnd.n4752 9.3005
R19097 gnd.n4617 gnd.n4616 9.3005
R19098 gnd.n4746 gnd.n4745 9.3005
R19099 gnd.n4744 gnd.n4619 9.3005
R19100 gnd.n4743 gnd.n4742 9.3005
R19101 gnd.n4621 gnd.n4620 9.3005
R19102 gnd.n4736 gnd.n4735 9.3005
R19103 gnd.n4734 gnd.n4623 9.3005
R19104 gnd.n4733 gnd.n4732 9.3005
R19105 gnd.n4625 gnd.n4624 9.3005
R19106 gnd.n4726 gnd.n4725 9.3005
R19107 gnd.n4724 gnd.n4627 9.3005
R19108 gnd.n4723 gnd.n4722 9.3005
R19109 gnd.n4629 gnd.n4628 9.3005
R19110 gnd.n4716 gnd.n4715 9.3005
R19111 gnd.n4714 gnd.n4631 9.3005
R19112 gnd.n4713 gnd.n4712 9.3005
R19113 gnd.n4633 gnd.n4632 9.3005
R19114 gnd.n4706 gnd.n4705 9.3005
R19115 gnd.n4704 gnd.n4635 9.3005
R19116 gnd.n4703 gnd.n4702 9.3005
R19117 gnd.n4637 gnd.n4636 9.3005
R19118 gnd.n4696 gnd.n4695 9.3005
R19119 gnd.n4694 gnd.n4639 9.3005
R19120 gnd.n4693 gnd.n4692 9.3005
R19121 gnd.n4641 gnd.n4640 9.3005
R19122 gnd.n4686 gnd.n4685 9.3005
R19123 gnd.n4684 gnd.n4643 9.3005
R19124 gnd.n4683 gnd.n4682 9.3005
R19125 gnd.n4645 gnd.n4644 9.3005
R19126 gnd.n4676 gnd.n4675 9.3005
R19127 gnd.n4674 gnd.n4647 9.3005
R19128 gnd.n4673 gnd.n4672 9.3005
R19129 gnd.n4649 gnd.n4648 9.3005
R19130 gnd.n4666 gnd.n4665 9.3005
R19131 gnd.n4664 gnd.n4651 9.3005
R19132 gnd.n4663 gnd.n4662 9.3005
R19133 gnd.n4653 gnd.n4652 9.3005
R19134 gnd.n4656 gnd.n4655 9.3005
R19135 gnd.n4654 gnd.n750 9.3005
R19136 gnd.n4865 gnd.n4864 9.3005
R19137 gnd.n3776 gnd.n3775 9.3005
R19138 gnd.n3749 gnd.n3748 9.3005
R19139 gnd.n3770 gnd.n3769 9.3005
R19140 gnd.n3768 gnd.n3767 9.3005
R19141 gnd.n3753 gnd.n3752 9.3005
R19142 gnd.n3762 gnd.n3761 9.3005
R19143 gnd.n3760 gnd.n3759 9.3005
R19144 gnd.n3744 gnd.n3743 9.3005
R19145 gnd.n3717 gnd.n3716 9.3005
R19146 gnd.n3738 gnd.n3737 9.3005
R19147 gnd.n3736 gnd.n3735 9.3005
R19148 gnd.n3721 gnd.n3720 9.3005
R19149 gnd.n3730 gnd.n3729 9.3005
R19150 gnd.n3728 gnd.n3727 9.3005
R19151 gnd.n3712 gnd.n3711 9.3005
R19152 gnd.n3685 gnd.n3684 9.3005
R19153 gnd.n3706 gnd.n3705 9.3005
R19154 gnd.n3704 gnd.n3703 9.3005
R19155 gnd.n3689 gnd.n3688 9.3005
R19156 gnd.n3698 gnd.n3697 9.3005
R19157 gnd.n3696 gnd.n3695 9.3005
R19158 gnd.n3681 gnd.n3680 9.3005
R19159 gnd.n3654 gnd.n3653 9.3005
R19160 gnd.n3675 gnd.n3674 9.3005
R19161 gnd.n3673 gnd.n3672 9.3005
R19162 gnd.n3658 gnd.n3657 9.3005
R19163 gnd.n3667 gnd.n3666 9.3005
R19164 gnd.n3665 gnd.n3664 9.3005
R19165 gnd.n3649 gnd.n3648 9.3005
R19166 gnd.n3622 gnd.n3621 9.3005
R19167 gnd.n3643 gnd.n3642 9.3005
R19168 gnd.n3641 gnd.n3640 9.3005
R19169 gnd.n3626 gnd.n3625 9.3005
R19170 gnd.n3635 gnd.n3634 9.3005
R19171 gnd.n3633 gnd.n3632 9.3005
R19172 gnd.n3617 gnd.n3616 9.3005
R19173 gnd.n3590 gnd.n3589 9.3005
R19174 gnd.n3611 gnd.n3610 9.3005
R19175 gnd.n3609 gnd.n3608 9.3005
R19176 gnd.n3594 gnd.n3593 9.3005
R19177 gnd.n3603 gnd.n3602 9.3005
R19178 gnd.n3601 gnd.n3600 9.3005
R19179 gnd.n3585 gnd.n3584 9.3005
R19180 gnd.n3558 gnd.n3557 9.3005
R19181 gnd.n3579 gnd.n3578 9.3005
R19182 gnd.n3577 gnd.n3576 9.3005
R19183 gnd.n3562 gnd.n3561 9.3005
R19184 gnd.n3571 gnd.n3570 9.3005
R19185 gnd.n3569 gnd.n3568 9.3005
R19186 gnd.n3554 gnd.n3553 9.3005
R19187 gnd.n3527 gnd.n3526 9.3005
R19188 gnd.n3548 gnd.n3547 9.3005
R19189 gnd.n3546 gnd.n3545 9.3005
R19190 gnd.n3531 gnd.n3530 9.3005
R19191 gnd.n3540 gnd.n3539 9.3005
R19192 gnd.n3538 gnd.n3537 9.3005
R19193 gnd.n3902 gnd.n3901 9.3005
R19194 gnd.n3900 gnd.n2438 9.3005
R19195 gnd.n3899 gnd.n3898 9.3005
R19196 gnd.n3895 gnd.n2439 9.3005
R19197 gnd.n3892 gnd.n2440 9.3005
R19198 gnd.n3891 gnd.n2441 9.3005
R19199 gnd.n3888 gnd.n2442 9.3005
R19200 gnd.n3887 gnd.n2443 9.3005
R19201 gnd.n3884 gnd.n2444 9.3005
R19202 gnd.n3883 gnd.n2445 9.3005
R19203 gnd.n3880 gnd.n2446 9.3005
R19204 gnd.n3879 gnd.n2447 9.3005
R19205 gnd.n3876 gnd.n2448 9.3005
R19206 gnd.n3875 gnd.n2449 9.3005
R19207 gnd.n3872 gnd.n3871 9.3005
R19208 gnd.n3870 gnd.n2450 9.3005
R19209 gnd.n3903 gnd.n2437 9.3005
R19210 gnd.n3144 gnd.n3143 9.3005
R19211 gnd.n2848 gnd.n2847 9.3005
R19212 gnd.n3171 gnd.n3170 9.3005
R19213 gnd.n3172 gnd.n2846 9.3005
R19214 gnd.n3176 gnd.n3173 9.3005
R19215 gnd.n3175 gnd.n3174 9.3005
R19216 gnd.n2820 gnd.n2819 9.3005
R19217 gnd.n3201 gnd.n3200 9.3005
R19218 gnd.n3202 gnd.n2818 9.3005
R19219 gnd.n3204 gnd.n3203 9.3005
R19220 gnd.n2798 gnd.n2797 9.3005
R19221 gnd.n3232 gnd.n3231 9.3005
R19222 gnd.n3233 gnd.n2796 9.3005
R19223 gnd.n3241 gnd.n3234 9.3005
R19224 gnd.n3240 gnd.n3235 9.3005
R19225 gnd.n3239 gnd.n3237 9.3005
R19226 gnd.n3236 gnd.n2745 9.3005
R19227 gnd.n3289 gnd.n2746 9.3005
R19228 gnd.n3288 gnd.n2747 9.3005
R19229 gnd.n3287 gnd.n2748 9.3005
R19230 gnd.n2767 gnd.n2749 9.3005
R19231 gnd.n2769 gnd.n2768 9.3005
R19232 gnd.n2635 gnd.n2634 9.3005
R19233 gnd.n3327 gnd.n3326 9.3005
R19234 gnd.n3328 gnd.n2633 9.3005
R19235 gnd.n3332 gnd.n3329 9.3005
R19236 gnd.n3331 gnd.n3330 9.3005
R19237 gnd.n2608 gnd.n2607 9.3005
R19238 gnd.n3367 gnd.n3366 9.3005
R19239 gnd.n3368 gnd.n2606 9.3005
R19240 gnd.n3372 gnd.n3369 9.3005
R19241 gnd.n3371 gnd.n3370 9.3005
R19242 gnd.n2581 gnd.n2580 9.3005
R19243 gnd.n3412 gnd.n3411 9.3005
R19244 gnd.n3413 gnd.n2579 9.3005
R19245 gnd.n3417 gnd.n3414 9.3005
R19246 gnd.n3416 gnd.n3415 9.3005
R19247 gnd.n2553 gnd.n2552 9.3005
R19248 gnd.n3452 gnd.n3451 9.3005
R19249 gnd.n3453 gnd.n2551 9.3005
R19250 gnd.n3457 gnd.n3454 9.3005
R19251 gnd.n3456 gnd.n3455 9.3005
R19252 gnd.n2526 gnd.n2525 9.3005
R19253 gnd.n3501 gnd.n3500 9.3005
R19254 gnd.n3502 gnd.n2524 9.3005
R19255 gnd.n3506 gnd.n3503 9.3005
R19256 gnd.n3505 gnd.n3504 9.3005
R19257 gnd.n2499 gnd.n2498 9.3005
R19258 gnd.n3795 gnd.n3794 9.3005
R19259 gnd.n3796 gnd.n2497 9.3005
R19260 gnd.n3802 gnd.n3797 9.3005
R19261 gnd.n3801 gnd.n3798 9.3005
R19262 gnd.n3800 gnd.n3799 9.3005
R19263 gnd.n3145 gnd.n3142 9.3005
R19264 gnd.n2927 gnd.n2886 9.3005
R19265 gnd.n2922 gnd.n2921 9.3005
R19266 gnd.n2920 gnd.n2887 9.3005
R19267 gnd.n2919 gnd.n2918 9.3005
R19268 gnd.n2915 gnd.n2888 9.3005
R19269 gnd.n2912 gnd.n2911 9.3005
R19270 gnd.n2910 gnd.n2889 9.3005
R19271 gnd.n2909 gnd.n2908 9.3005
R19272 gnd.n2905 gnd.n2890 9.3005
R19273 gnd.n2902 gnd.n2901 9.3005
R19274 gnd.n2900 gnd.n2891 9.3005
R19275 gnd.n2899 gnd.n2898 9.3005
R19276 gnd.n2895 gnd.n2893 9.3005
R19277 gnd.n2892 gnd.n2872 9.3005
R19278 gnd.n3139 gnd.n2871 9.3005
R19279 gnd.n3141 gnd.n3140 9.3005
R19280 gnd.n2929 gnd.n2928 9.3005
R19281 gnd.n3152 gnd.n2858 9.3005
R19282 gnd.n3159 gnd.n2859 9.3005
R19283 gnd.n3161 gnd.n3160 9.3005
R19284 gnd.n3162 gnd.n2839 9.3005
R19285 gnd.n3181 gnd.n3180 9.3005
R19286 gnd.n3183 gnd.n2831 9.3005
R19287 gnd.n3190 gnd.n2833 9.3005
R19288 gnd.n3191 gnd.n2828 9.3005
R19289 gnd.n3193 gnd.n3192 9.3005
R19290 gnd.n2829 gnd.n2814 9.3005
R19291 gnd.n3209 gnd.n2812 9.3005
R19292 gnd.n3213 gnd.n3212 9.3005
R19293 gnd.n3211 gnd.n2788 9.3005
R19294 gnd.n3248 gnd.n2787 9.3005
R19295 gnd.n3251 gnd.n3250 9.3005
R19296 gnd.n2784 gnd.n2783 9.3005
R19297 gnd.n3257 gnd.n2785 9.3005
R19298 gnd.n3259 gnd.n3258 9.3005
R19299 gnd.n3261 gnd.n2782 9.3005
R19300 gnd.n3264 gnd.n3263 9.3005
R19301 gnd.n3267 gnd.n3265 9.3005
R19302 gnd.n3269 gnd.n3268 9.3005
R19303 gnd.n3275 gnd.n3270 9.3005
R19304 gnd.n3274 gnd.n3273 9.3005
R19305 gnd.n2626 gnd.n2625 9.3005
R19306 gnd.n3341 gnd.n3340 9.3005
R19307 gnd.n3342 gnd.n2619 9.3005
R19308 gnd.n3350 gnd.n2618 9.3005
R19309 gnd.n3353 gnd.n3352 9.3005
R19310 gnd.n3355 gnd.n3354 9.3005
R19311 gnd.n3358 gnd.n2601 9.3005
R19312 gnd.n3356 gnd.n2599 9.3005
R19313 gnd.n3378 gnd.n2597 9.3005
R19314 gnd.n3380 gnd.n3379 9.3005
R19315 gnd.n2571 gnd.n2570 9.3005
R19316 gnd.n3426 gnd.n3425 9.3005
R19317 gnd.n3427 gnd.n2564 9.3005
R19318 gnd.n3435 gnd.n2563 9.3005
R19319 gnd.n3438 gnd.n3437 9.3005
R19320 gnd.n3440 gnd.n3439 9.3005
R19321 gnd.n3443 gnd.n2546 9.3005
R19322 gnd.n3441 gnd.n2544 9.3005
R19323 gnd.n3463 gnd.n2542 9.3005
R19324 gnd.n3465 gnd.n3464 9.3005
R19325 gnd.n2517 gnd.n2516 9.3005
R19326 gnd.n3515 gnd.n3514 9.3005
R19327 gnd.n3516 gnd.n2510 9.3005
R19328 gnd.n3524 gnd.n2509 9.3005
R19329 gnd.n3783 gnd.n3782 9.3005
R19330 gnd.n3785 gnd.n3784 9.3005
R19331 gnd.n3786 gnd.n2490 9.3005
R19332 gnd.n3810 gnd.n3809 9.3005
R19333 gnd.n2491 gnd.n2453 9.3005
R19334 gnd.n3150 gnd.n3149 9.3005
R19335 gnd.n3866 gnd.n2454 9.3005
R19336 gnd.n3865 gnd.n2456 9.3005
R19337 gnd.n3862 gnd.n2457 9.3005
R19338 gnd.n3861 gnd.n2458 9.3005
R19339 gnd.n3858 gnd.n2459 9.3005
R19340 gnd.n3857 gnd.n2460 9.3005
R19341 gnd.n3854 gnd.n2461 9.3005
R19342 gnd.n3853 gnd.n2462 9.3005
R19343 gnd.n3850 gnd.n2463 9.3005
R19344 gnd.n3849 gnd.n2464 9.3005
R19345 gnd.n3846 gnd.n2465 9.3005
R19346 gnd.n3845 gnd.n2466 9.3005
R19347 gnd.n3842 gnd.n2467 9.3005
R19348 gnd.n3841 gnd.n2468 9.3005
R19349 gnd.n3838 gnd.n2469 9.3005
R19350 gnd.n3837 gnd.n2470 9.3005
R19351 gnd.n3834 gnd.n2471 9.3005
R19352 gnd.n3833 gnd.n2472 9.3005
R19353 gnd.n3830 gnd.n2473 9.3005
R19354 gnd.n3829 gnd.n2474 9.3005
R19355 gnd.n3826 gnd.n2475 9.3005
R19356 gnd.n3825 gnd.n2476 9.3005
R19357 gnd.n3822 gnd.n2480 9.3005
R19358 gnd.n3821 gnd.n2481 9.3005
R19359 gnd.n3818 gnd.n2482 9.3005
R19360 gnd.n3817 gnd.n2483 9.3005
R19361 gnd.n3868 gnd.n3867 9.3005
R19362 gnd.n3319 gnd.n3303 9.3005
R19363 gnd.n3318 gnd.n3304 9.3005
R19364 gnd.n3317 gnd.n3305 9.3005
R19365 gnd.n3315 gnd.n3306 9.3005
R19366 gnd.n3314 gnd.n3307 9.3005
R19367 gnd.n3312 gnd.n3308 9.3005
R19368 gnd.n3311 gnd.n3309 9.3005
R19369 gnd.n2589 gnd.n2588 9.3005
R19370 gnd.n3388 gnd.n3387 9.3005
R19371 gnd.n3389 gnd.n2587 9.3005
R19372 gnd.n3406 gnd.n3390 9.3005
R19373 gnd.n3405 gnd.n3391 9.3005
R19374 gnd.n3404 gnd.n3392 9.3005
R19375 gnd.n3402 gnd.n3393 9.3005
R19376 gnd.n3401 gnd.n3394 9.3005
R19377 gnd.n3399 gnd.n3395 9.3005
R19378 gnd.n3398 gnd.n3396 9.3005
R19379 gnd.n2533 gnd.n2532 9.3005
R19380 gnd.n3473 gnd.n3472 9.3005
R19381 gnd.n3474 gnd.n2531 9.3005
R19382 gnd.n3495 gnd.n3475 9.3005
R19383 gnd.n3494 gnd.n3476 9.3005
R19384 gnd.n3493 gnd.n3477 9.3005
R19385 gnd.n3490 gnd.n3478 9.3005
R19386 gnd.n3489 gnd.n3479 9.3005
R19387 gnd.n3487 gnd.n3480 9.3005
R19388 gnd.n3486 gnd.n3481 9.3005
R19389 gnd.n3484 gnd.n3483 9.3005
R19390 gnd.n3482 gnd.n2485 9.3005
R19391 gnd.n3060 gnd.n3059 9.3005
R19392 gnd.n2950 gnd.n2949 9.3005
R19393 gnd.n3074 gnd.n3073 9.3005
R19394 gnd.n3075 gnd.n2948 9.3005
R19395 gnd.n3077 gnd.n3076 9.3005
R19396 gnd.n2938 gnd.n2937 9.3005
R19397 gnd.n3090 gnd.n3089 9.3005
R19398 gnd.n3091 gnd.n2936 9.3005
R19399 gnd.n3123 gnd.n3092 9.3005
R19400 gnd.n3122 gnd.n3093 9.3005
R19401 gnd.n3121 gnd.n3094 9.3005
R19402 gnd.n3120 gnd.n3095 9.3005
R19403 gnd.n3117 gnd.n3096 9.3005
R19404 gnd.n3116 gnd.n3097 9.3005
R19405 gnd.n3115 gnd.n3098 9.3005
R19406 gnd.n3113 gnd.n3099 9.3005
R19407 gnd.n3112 gnd.n3100 9.3005
R19408 gnd.n3109 gnd.n3101 9.3005
R19409 gnd.n3108 gnd.n3102 9.3005
R19410 gnd.n3107 gnd.n3103 9.3005
R19411 gnd.n3105 gnd.n3104 9.3005
R19412 gnd.n2804 gnd.n2803 9.3005
R19413 gnd.n3221 gnd.n3220 9.3005
R19414 gnd.n3222 gnd.n2802 9.3005
R19415 gnd.n3226 gnd.n3223 9.3005
R19416 gnd.n3225 gnd.n3224 9.3005
R19417 gnd.n2726 gnd.n2725 9.3005
R19418 gnd.n3301 gnd.n3300 9.3005
R19419 gnd.n3058 gnd.n2959 9.3005
R19420 gnd.n2961 gnd.n2960 9.3005
R19421 gnd.n3005 gnd.n3003 9.3005
R19422 gnd.n3006 gnd.n3002 9.3005
R19423 gnd.n3009 gnd.n2998 9.3005
R19424 gnd.n3010 gnd.n2997 9.3005
R19425 gnd.n3013 gnd.n2996 9.3005
R19426 gnd.n3014 gnd.n2995 9.3005
R19427 gnd.n3017 gnd.n2994 9.3005
R19428 gnd.n3018 gnd.n2993 9.3005
R19429 gnd.n3021 gnd.n2992 9.3005
R19430 gnd.n3022 gnd.n2991 9.3005
R19431 gnd.n3025 gnd.n2990 9.3005
R19432 gnd.n3026 gnd.n2989 9.3005
R19433 gnd.n3029 gnd.n2988 9.3005
R19434 gnd.n3030 gnd.n2987 9.3005
R19435 gnd.n3033 gnd.n2986 9.3005
R19436 gnd.n3034 gnd.n2985 9.3005
R19437 gnd.n3037 gnd.n2984 9.3005
R19438 gnd.n3038 gnd.n2983 9.3005
R19439 gnd.n3041 gnd.n2982 9.3005
R19440 gnd.n3042 gnd.n2981 9.3005
R19441 gnd.n3045 gnd.n2980 9.3005
R19442 gnd.n3047 gnd.n2979 9.3005
R19443 gnd.n3048 gnd.n2978 9.3005
R19444 gnd.n3049 gnd.n2977 9.3005
R19445 gnd.n3050 gnd.n2976 9.3005
R19446 gnd.n3057 gnd.n3056 9.3005
R19447 gnd.n3066 gnd.n3065 9.3005
R19448 gnd.n3067 gnd.n2953 9.3005
R19449 gnd.n3069 gnd.n3068 9.3005
R19450 gnd.n2944 gnd.n2943 9.3005
R19451 gnd.n3082 gnd.n3081 9.3005
R19452 gnd.n3083 gnd.n2942 9.3005
R19453 gnd.n3085 gnd.n3084 9.3005
R19454 gnd.n2931 gnd.n2930 9.3005
R19455 gnd.n3128 gnd.n3127 9.3005
R19456 gnd.n3129 gnd.n2885 9.3005
R19457 gnd.n3133 gnd.n3131 9.3005
R19458 gnd.n3132 gnd.n2864 9.3005
R19459 gnd.n3151 gnd.n2863 9.3005
R19460 gnd.n3154 gnd.n3153 9.3005
R19461 gnd.n2857 gnd.n2856 9.3005
R19462 gnd.n3165 gnd.n3163 9.3005
R19463 gnd.n3164 gnd.n2838 9.3005
R19464 gnd.n3182 gnd.n2837 9.3005
R19465 gnd.n3185 gnd.n3184 9.3005
R19466 gnd.n2832 gnd.n2827 9.3005
R19467 gnd.n3195 gnd.n3194 9.3005
R19468 gnd.n2830 gnd.n2810 9.3005
R19469 gnd.n3216 gnd.n2811 9.3005
R19470 gnd.n3215 gnd.n3214 9.3005
R19471 gnd.n2813 gnd.n2789 9.3005
R19472 gnd.n3247 gnd.n3246 9.3005
R19473 gnd.n3249 gnd.n2734 9.3005
R19474 gnd.n3296 gnd.n2735 9.3005
R19475 gnd.n3295 gnd.n2736 9.3005
R19476 gnd.n3294 gnd.n2737 9.3005
R19477 gnd.n3260 gnd.n2738 9.3005
R19478 gnd.n3262 gnd.n2756 9.3005
R19479 gnd.n3282 gnd.n2757 9.3005
R19480 gnd.n3281 gnd.n2758 9.3005
R19481 gnd.n3280 gnd.n2759 9.3005
R19482 gnd.n3271 gnd.n2760 9.3005
R19483 gnd.n3272 gnd.n2627 9.3005
R19484 gnd.n3338 gnd.n3337 9.3005
R19485 gnd.n3339 gnd.n2620 9.3005
R19486 gnd.n3349 gnd.n3348 9.3005
R19487 gnd.n3351 gnd.n2616 9.3005
R19488 gnd.n3361 gnd.n2617 9.3005
R19489 gnd.n3360 gnd.n3359 9.3005
R19490 gnd.n3357 gnd.n2595 9.3005
R19491 gnd.n3383 gnd.n2596 9.3005
R19492 gnd.n3382 gnd.n3381 9.3005
R19493 gnd.n2598 gnd.n2572 9.3005
R19494 gnd.n3423 gnd.n3422 9.3005
R19495 gnd.n3424 gnd.n2565 9.3005
R19496 gnd.n3434 gnd.n3433 9.3005
R19497 gnd.n3436 gnd.n2561 9.3005
R19498 gnd.n3446 gnd.n2562 9.3005
R19499 gnd.n3445 gnd.n3444 9.3005
R19500 gnd.n3442 gnd.n2540 9.3005
R19501 gnd.n3468 gnd.n2541 9.3005
R19502 gnd.n3467 gnd.n3466 9.3005
R19503 gnd.n2543 gnd.n2518 9.3005
R19504 gnd.n3512 gnd.n3511 9.3005
R19505 gnd.n3513 gnd.n2511 9.3005
R19506 gnd.n3523 gnd.n3522 9.3005
R19507 gnd.n3781 gnd.n2507 9.3005
R19508 gnd.n3789 gnd.n2508 9.3005
R19509 gnd.n3788 gnd.n3787 9.3005
R19510 gnd.n2489 gnd.n2488 9.3005
R19511 gnd.n3812 gnd.n3811 9.3005
R19512 gnd.n2955 gnd.n2954 9.3005
R19513 gnd.n4435 gnd.n2266 9.3005
R19514 gnd.n4208 gnd.n4149 9.3005
R19515 gnd.n4206 gnd.n4150 9.3005
R19516 gnd.n4205 gnd.n4151 9.3005
R19517 gnd.n4203 gnd.n4152 9.3005
R19518 gnd.n4202 gnd.n4153 9.3005
R19519 gnd.n4200 gnd.n4154 9.3005
R19520 gnd.n4199 gnd.n4155 9.3005
R19521 gnd.n4197 gnd.n4156 9.3005
R19522 gnd.n4196 gnd.n4157 9.3005
R19523 gnd.n4194 gnd.n4158 9.3005
R19524 gnd.n4193 gnd.n4159 9.3005
R19525 gnd.n4191 gnd.n4160 9.3005
R19526 gnd.n4190 gnd.n4161 9.3005
R19527 gnd.n4188 gnd.n4162 9.3005
R19528 gnd.n4187 gnd.n4163 9.3005
R19529 gnd.n4185 gnd.n4164 9.3005
R19530 gnd.n4184 gnd.n4165 9.3005
R19531 gnd.n4182 gnd.n4166 9.3005
R19532 gnd.n4181 gnd.n4167 9.3005
R19533 gnd.n4179 gnd.n4168 9.3005
R19534 gnd.n4178 gnd.n4169 9.3005
R19535 gnd.n4176 gnd.n4170 9.3005
R19536 gnd.n4175 gnd.n4171 9.3005
R19537 gnd.n4173 gnd.n4172 9.3005
R19538 gnd.n2294 gnd.n2293 9.3005
R19539 gnd.n4399 gnd.n4398 9.3005
R19540 gnd.n4400 gnd.n2292 9.3005
R19541 gnd.n4404 gnd.n4401 9.3005
R19542 gnd.n4403 gnd.n4402 9.3005
R19543 gnd.n2269 gnd.n2268 9.3005
R19544 gnd.n4434 gnd.n4433 9.3005
R19545 gnd.n4210 gnd.n4209 9.3005
R19546 gnd.n1846 gnd.n1751 9.3005
R19547 gnd.n1845 gnd.n1844 9.3005
R19548 gnd.n1754 gnd.n1753 9.3005
R19549 gnd.n1837 gnd.n1836 9.3005
R19550 gnd.n1835 gnd.n1756 9.3005
R19551 gnd.n1834 gnd.n1833 9.3005
R19552 gnd.n1758 gnd.n1757 9.3005
R19553 gnd.n1827 gnd.n1826 9.3005
R19554 gnd.n1825 gnd.n1824 9.3005
R19555 gnd.n1764 gnd.n1763 9.3005
R19556 gnd.n1819 gnd.n1818 9.3005
R19557 gnd.n1817 gnd.n1766 9.3005
R19558 gnd.n1816 gnd.n1815 9.3005
R19559 gnd.n1768 gnd.n1767 9.3005
R19560 gnd.n1809 gnd.n1808 9.3005
R19561 gnd.n1807 gnd.n1770 9.3005
R19562 gnd.n1806 gnd.n1805 9.3005
R19563 gnd.n1772 gnd.n1771 9.3005
R19564 gnd.n1799 gnd.n1798 9.3005
R19565 gnd.n1797 gnd.n1774 9.3005
R19566 gnd.n1796 gnd.n1795 9.3005
R19567 gnd.n1776 gnd.n1775 9.3005
R19568 gnd.n1789 gnd.n1788 9.3005
R19569 gnd.n1787 gnd.n1778 9.3005
R19570 gnd.n1786 gnd.n1785 9.3005
R19571 gnd.n1781 gnd.n1780 9.3005
R19572 gnd.n1949 gnd.n1948 9.3005
R19573 gnd.n1848 gnd.n1847 9.3005
R19574 gnd.n1853 gnd.n1851 9.3005
R19575 gnd.n1941 gnd.n1854 9.3005
R19576 gnd.n1940 gnd.n1855 9.3005
R19577 gnd.n1939 gnd.n1856 9.3005
R19578 gnd.n1860 gnd.n1857 9.3005
R19579 gnd.n1934 gnd.n1861 9.3005
R19580 gnd.n1933 gnd.n1932 9.3005
R19581 gnd.n1931 gnd.n1862 9.3005
R19582 gnd.n1930 gnd.n1929 9.3005
R19583 gnd.n1866 gnd.n1865 9.3005
R19584 gnd.n1871 gnd.n1869 9.3005
R19585 gnd.n1922 gnd.n1872 9.3005
R19586 gnd.n1921 gnd.n1873 9.3005
R19587 gnd.n1920 gnd.n1874 9.3005
R19588 gnd.n1878 gnd.n1875 9.3005
R19589 gnd.n1915 gnd.n1879 9.3005
R19590 gnd.n1914 gnd.n1880 9.3005
R19591 gnd.n1913 gnd.n1881 9.3005
R19592 gnd.n1885 gnd.n1882 9.3005
R19593 gnd.n1908 gnd.n1886 9.3005
R19594 gnd.n1907 gnd.n1887 9.3005
R19595 gnd.n1906 gnd.n1888 9.3005
R19596 gnd.n1892 gnd.n1889 9.3005
R19597 gnd.n1901 gnd.n1893 9.3005
R19598 gnd.n1900 gnd.n1894 9.3005
R19599 gnd.n1899 gnd.n1895 9.3005
R19600 gnd.n840 gnd.n837 9.3005
R19601 gnd.n6404 gnd.n6403 9.3005
R19602 gnd.n1950 gnd.n1750 9.3005
R19603 gnd.n2277 gnd.n2276 9.3005
R19604 gnd.n4424 gnd.n4423 9.3005
R19605 gnd.n4425 gnd.n2275 9.3005
R19606 gnd.n4429 gnd.n4426 9.3005
R19607 gnd.n4428 gnd.n4427 9.3005
R19608 gnd.n2251 gnd.n2250 9.3005
R19609 gnd.n4458 gnd.n4457 9.3005
R19610 gnd.n4459 gnd.n2249 9.3005
R19611 gnd.n4463 gnd.n4460 9.3005
R19612 gnd.n4462 gnd.n4461 9.3005
R19613 gnd.n2226 gnd.n2225 9.3005
R19614 gnd.n4492 gnd.n4491 9.3005
R19615 gnd.n4493 gnd.n2224 9.3005
R19616 gnd.n4497 gnd.n4494 9.3005
R19617 gnd.n4496 gnd.n4495 9.3005
R19618 gnd.n2200 gnd.n2199 9.3005
R19619 gnd.n4527 gnd.n4526 9.3005
R19620 gnd.n4528 gnd.n2198 9.3005
R19621 gnd.n4533 gnd.n4529 9.3005
R19622 gnd.n4532 gnd.n4531 9.3005
R19623 gnd.n4530 gnd.n759 9.3005
R19624 gnd.n6450 gnd.n760 9.3005
R19625 gnd.n6449 gnd.n761 9.3005
R19626 gnd.n6448 gnd.n762 9.3005
R19627 gnd.n782 gnd.n763 9.3005
R19628 gnd.n6438 gnd.n783 9.3005
R19629 gnd.n6437 gnd.n784 9.3005
R19630 gnd.n6436 gnd.n785 9.3005
R19631 gnd.n802 gnd.n786 9.3005
R19632 gnd.n6426 gnd.n803 9.3005
R19633 gnd.n6425 gnd.n804 9.3005
R19634 gnd.n6424 gnd.n805 9.3005
R19635 gnd.n823 gnd.n806 9.3005
R19636 gnd.n6414 gnd.n824 9.3005
R19637 gnd.n6413 gnd.n825 9.3005
R19638 gnd.n6412 gnd.n826 9.3005
R19639 gnd.n1779 gnd.n827 9.3005
R19640 gnd.n4266 gnd.n2409 9.3005
R19641 gnd.n4268 gnd.n4267 9.3005
R19642 gnd.n2394 gnd.n2393 9.3005
R19643 gnd.n4285 gnd.n4284 9.3005
R19644 gnd.n4286 gnd.n2392 9.3005
R19645 gnd.n4288 gnd.n4287 9.3005
R19646 gnd.n2375 gnd.n2374 9.3005
R19647 gnd.n4305 gnd.n4304 9.3005
R19648 gnd.n4306 gnd.n2373 9.3005
R19649 gnd.n4308 gnd.n4307 9.3005
R19650 gnd.n2358 gnd.n2357 9.3005
R19651 gnd.n4325 gnd.n4324 9.3005
R19652 gnd.n4326 gnd.n2356 9.3005
R19653 gnd.n4328 gnd.n4327 9.3005
R19654 gnd.n2339 gnd.n2338 9.3005
R19655 gnd.n4345 gnd.n4344 9.3005
R19656 gnd.n4346 gnd.n2337 9.3005
R19657 gnd.n4348 gnd.n4347 9.3005
R19658 gnd.n2322 gnd.n2321 9.3005
R19659 gnd.n4365 gnd.n4364 9.3005
R19660 gnd.n4366 gnd.n2320 9.3005
R19661 gnd.n4368 gnd.n4367 9.3005
R19662 gnd.n2302 gnd.n2301 9.3005
R19663 gnd.n4389 gnd.n4388 9.3005
R19664 gnd.n4390 gnd.n2300 9.3005
R19665 gnd.n4394 gnd.n4391 9.3005
R19666 gnd.n4393 gnd.n4392 9.3005
R19667 gnd.n4265 gnd.n4264 9.3005
R19668 gnd.n3915 gnd.n3912 9.3005
R19669 gnd.n4112 gnd.n3916 9.3005
R19670 gnd.n4114 gnd.n4113 9.3005
R19671 gnd.n4111 gnd.n3918 9.3005
R19672 gnd.n4110 gnd.n4109 9.3005
R19673 gnd.n3920 gnd.n3919 9.3005
R19674 gnd.n4103 gnd.n4102 9.3005
R19675 gnd.n4101 gnd.n3922 9.3005
R19676 gnd.n4100 gnd.n4099 9.3005
R19677 gnd.n3924 gnd.n3923 9.3005
R19678 gnd.n4093 gnd.n4092 9.3005
R19679 gnd.n4091 gnd.n3926 9.3005
R19680 gnd.n4090 gnd.n4089 9.3005
R19681 gnd.n3928 gnd.n3927 9.3005
R19682 gnd.n4083 gnd.n4082 9.3005
R19683 gnd.n4081 gnd.n3930 9.3005
R19684 gnd.n4080 gnd.n4079 9.3005
R19685 gnd.n3932 gnd.n3931 9.3005
R19686 gnd.n4073 gnd.n4072 9.3005
R19687 gnd.n4071 gnd.n3934 9.3005
R19688 gnd.n3936 gnd.n3935 9.3005
R19689 gnd.n4061 gnd.n4060 9.3005
R19690 gnd.n4059 gnd.n3938 9.3005
R19691 gnd.n4058 gnd.n4057 9.3005
R19692 gnd.n3940 gnd.n3939 9.3005
R19693 gnd.n4051 gnd.n4050 9.3005
R19694 gnd.n4049 gnd.n3942 9.3005
R19695 gnd.n4048 gnd.n4047 9.3005
R19696 gnd.n3944 gnd.n3943 9.3005
R19697 gnd.n4041 gnd.n4040 9.3005
R19698 gnd.n4039 gnd.n3946 9.3005
R19699 gnd.n4038 gnd.n4037 9.3005
R19700 gnd.n3948 gnd.n3947 9.3005
R19701 gnd.n4031 gnd.n4030 9.3005
R19702 gnd.n4029 gnd.n3950 9.3005
R19703 gnd.n4028 gnd.n4027 9.3005
R19704 gnd.n3952 gnd.n3951 9.3005
R19705 gnd.n4021 gnd.n4020 9.3005
R19706 gnd.n4019 gnd.n3954 9.3005
R19707 gnd.n4018 gnd.n4017 9.3005
R19708 gnd.n3956 gnd.n3955 9.3005
R19709 gnd.n4011 gnd.n4010 9.3005
R19710 gnd.n4009 gnd.n3961 9.3005
R19711 gnd.n4008 gnd.n4007 9.3005
R19712 gnd.n3963 gnd.n3962 9.3005
R19713 gnd.n4001 gnd.n4000 9.3005
R19714 gnd.n3999 gnd.n3965 9.3005
R19715 gnd.n3998 gnd.n3997 9.3005
R19716 gnd.n3967 gnd.n3966 9.3005
R19717 gnd.n3991 gnd.n3990 9.3005
R19718 gnd.n3989 gnd.n3969 9.3005
R19719 gnd.n3988 gnd.n3987 9.3005
R19720 gnd.n3971 gnd.n3970 9.3005
R19721 gnd.n3981 gnd.n3980 9.3005
R19722 gnd.n3979 gnd.n3973 9.3005
R19723 gnd.n3978 gnd.n3977 9.3005
R19724 gnd.n3974 gnd.n2410 9.3005
R19725 gnd.n4070 gnd.n4069 9.3005
R19726 gnd.n4122 gnd.n4121 9.3005
R19727 gnd.n4218 gnd.n4217 9.3005
R19728 gnd.n4219 gnd.n4145 9.3005
R19729 gnd.n4144 gnd.n4142 9.3005
R19730 gnd.n4225 gnd.n4141 9.3005
R19731 gnd.n4226 gnd.n4140 9.3005
R19732 gnd.n4227 gnd.n4139 9.3005
R19733 gnd.n4138 gnd.n4136 9.3005
R19734 gnd.n4233 gnd.n4135 9.3005
R19735 gnd.n4234 gnd.n4134 9.3005
R19736 gnd.n4235 gnd.n4133 9.3005
R19737 gnd.n4132 gnd.n4130 9.3005
R19738 gnd.n4241 gnd.n4129 9.3005
R19739 gnd.n4242 gnd.n4128 9.3005
R19740 gnd.n4243 gnd.n4127 9.3005
R19741 gnd.n4126 gnd.n4124 9.3005
R19742 gnd.n4249 gnd.n4123 9.3005
R19743 gnd.n4251 gnd.n4250 9.3005
R19744 gnd.n4216 gnd.n4148 9.3005
R19745 gnd.n4215 gnd.n4214 9.3005
R19746 gnd.n4256 gnd.n4255 9.3005
R19747 gnd.n4257 gnd.n2403 9.3005
R19748 gnd.n4273 gnd.n2404 9.3005
R19749 gnd.n4274 gnd.n2402 9.3005
R19750 gnd.n4276 gnd.n4275 9.3005
R19751 gnd.n4277 gnd.n2385 9.3005
R19752 gnd.n4293 gnd.n2386 9.3005
R19753 gnd.n4294 gnd.n2384 9.3005
R19754 gnd.n4296 gnd.n4295 9.3005
R19755 gnd.n4297 gnd.n2367 9.3005
R19756 gnd.n4313 gnd.n2368 9.3005
R19757 gnd.n4314 gnd.n2366 9.3005
R19758 gnd.n4316 gnd.n4315 9.3005
R19759 gnd.n4317 gnd.n2349 9.3005
R19760 gnd.n4333 gnd.n2350 9.3005
R19761 gnd.n4334 gnd.n2348 9.3005
R19762 gnd.n4336 gnd.n4335 9.3005
R19763 gnd.n4337 gnd.n2331 9.3005
R19764 gnd.n4353 gnd.n2332 9.3005
R19765 gnd.n4354 gnd.n2330 9.3005
R19766 gnd.n4356 gnd.n4355 9.3005
R19767 gnd.n4357 gnd.n2313 9.3005
R19768 gnd.n4373 gnd.n2314 9.3005
R19769 gnd.n4374 gnd.n2311 9.3005
R19770 gnd.n4376 gnd.n2312 9.3005
R19771 gnd.n4378 gnd.n4377 9.3005
R19772 gnd.n4379 gnd.n2287 9.3005
R19773 gnd.n4408 gnd.n2288 9.3005
R19774 gnd.n4409 gnd.n2285 9.3005
R19775 gnd.n4411 gnd.n2286 9.3005
R19776 gnd.n4413 gnd.n4412 9.3005
R19777 gnd.n4414 gnd.n2261 9.3005
R19778 gnd.n4442 gnd.n2262 9.3005
R19779 gnd.n4443 gnd.n2259 9.3005
R19780 gnd.n4445 gnd.n2260 9.3005
R19781 gnd.n4447 gnd.n4446 9.3005
R19782 gnd.n4448 gnd.n2235 9.3005
R19783 gnd.n4476 gnd.n2236 9.3005
R19784 gnd.n4477 gnd.n2233 9.3005
R19785 gnd.n4479 gnd.n2234 9.3005
R19786 gnd.n4481 gnd.n4480 9.3005
R19787 gnd.n4482 gnd.n2209 9.3005
R19788 gnd.n4510 gnd.n2210 9.3005
R19789 gnd.n4511 gnd.n2207 9.3005
R19790 gnd.n4513 gnd.n2208 9.3005
R19791 gnd.n4519 gnd.n4514 9.3005
R19792 gnd.n4518 gnd.n4517 9.3005
R19793 gnd.n4515 gnd.n2182 9.3005
R19794 gnd.n4551 gnd.n2181 9.3005
R19795 gnd.n4554 gnd.n4552 9.3005
R19796 gnd.n4555 gnd.n772 9.3005
R19797 gnd.n4556 gnd.n773 9.3005
R19798 gnd.n2176 gnd.n774 9.3005
R19799 gnd.n4904 gnd.n2177 9.3005
R19800 gnd.n4905 gnd.n792 9.3005
R19801 gnd.n4906 gnd.n793 9.3005
R19802 gnd.n2171 gnd.n794 9.3005
R19803 gnd.n4918 gnd.n2172 9.3005
R19804 gnd.n4919 gnd.n813 9.3005
R19805 gnd.n4926 gnd.n814 9.3005
R19806 gnd.n4925 gnd.n815 9.3005
R19807 gnd.n4924 gnd.n4920 9.3005
R19808 gnd.n4921 gnd.n834 9.3005
R19809 gnd.n6406 gnd.n835 9.3005
R19810 gnd.n4254 gnd.n4253 9.3005
R19811 gnd.n4259 gnd.n4256 9.3005
R19812 gnd.n4258 gnd.n4257 9.3005
R19813 gnd.n2404 gnd.n2401 9.3005
R19814 gnd.n4280 gnd.n2402 9.3005
R19815 gnd.n4279 gnd.n4276 9.3005
R19816 gnd.n4278 gnd.n4277 9.3005
R19817 gnd.n2386 gnd.n2383 9.3005
R19818 gnd.n4300 gnd.n2384 9.3005
R19819 gnd.n4299 gnd.n4296 9.3005
R19820 gnd.n4298 gnd.n4297 9.3005
R19821 gnd.n2368 gnd.n2365 9.3005
R19822 gnd.n4320 gnd.n2366 9.3005
R19823 gnd.n4319 gnd.n4316 9.3005
R19824 gnd.n4318 gnd.n4317 9.3005
R19825 gnd.n2350 gnd.n2347 9.3005
R19826 gnd.n4340 gnd.n2348 9.3005
R19827 gnd.n4339 gnd.n4336 9.3005
R19828 gnd.n4338 gnd.n4337 9.3005
R19829 gnd.n2332 gnd.n2329 9.3005
R19830 gnd.n4360 gnd.n2330 9.3005
R19831 gnd.n4359 gnd.n4356 9.3005
R19832 gnd.n4358 gnd.n4357 9.3005
R19833 gnd.n2314 gnd.n2310 9.3005
R19834 gnd.n4384 gnd.n2311 9.3005
R19835 gnd.n4383 gnd.n2312 9.3005
R19836 gnd.n4382 gnd.n4378 9.3005
R19837 gnd.n4381 gnd.n4379 9.3005
R19838 gnd.n2288 gnd.n2284 9.3005
R19839 gnd.n4419 gnd.n2285 9.3005
R19840 gnd.n4418 gnd.n2286 9.3005
R19841 gnd.n4417 gnd.n4413 9.3005
R19842 gnd.n4416 gnd.n4414 9.3005
R19843 gnd.n2262 gnd.n2258 9.3005
R19844 gnd.n4453 gnd.n2259 9.3005
R19845 gnd.n4452 gnd.n2260 9.3005
R19846 gnd.n4451 gnd.n4447 9.3005
R19847 gnd.n4450 gnd.n4448 9.3005
R19848 gnd.n2236 gnd.n2232 9.3005
R19849 gnd.n4487 gnd.n2233 9.3005
R19850 gnd.n4486 gnd.n2234 9.3005
R19851 gnd.n4485 gnd.n4481 9.3005
R19852 gnd.n4484 gnd.n4482 9.3005
R19853 gnd.n2210 gnd.n2206 9.3005
R19854 gnd.n4522 gnd.n2207 9.3005
R19855 gnd.n4521 gnd.n2208 9.3005
R19856 gnd.n4520 gnd.n4519 9.3005
R19857 gnd.n4518 gnd.n2183 9.3005
R19858 gnd.n4549 gnd.n2182 9.3005
R19859 gnd.n4551 gnd.n4550 9.3005
R19860 gnd.n4552 gnd.n771 9.3005
R19861 gnd.n6444 gnd.n772 9.3005
R19862 gnd.n6443 gnd.n773 9.3005
R19863 gnd.n6442 gnd.n774 9.3005
R19864 gnd.n2177 gnd.n775 9.3005
R19865 gnd.n6432 gnd.n792 9.3005
R19866 gnd.n6431 gnd.n793 9.3005
R19867 gnd.n6430 gnd.n794 9.3005
R19868 gnd.n2172 gnd.n795 9.3005
R19869 gnd.n6420 gnd.n813 9.3005
R19870 gnd.n6419 gnd.n814 9.3005
R19871 gnd.n6418 gnd.n815 9.3005
R19872 gnd.n4920 gnd.n816 9.3005
R19873 gnd.n6408 gnd.n834 9.3005
R19874 gnd.n6407 gnd.n6406 9.3005
R19875 gnd.n4260 gnd.n4253 9.3005
R19876 gnd.n6230 gnd.n6229 9.3005
R19877 gnd.n6381 gnd.n866 9.3005
R19878 gnd.n6380 gnd.n6379 9.3005
R19879 gnd.n6378 gnd.n868 9.3005
R19880 gnd.n6377 gnd.n6376 9.3005
R19881 gnd.n6375 gnd.n872 9.3005
R19882 gnd.n6374 gnd.n6373 9.3005
R19883 gnd.n6372 gnd.n873 9.3005
R19884 gnd.n6371 gnd.n6370 9.3005
R19885 gnd.n6369 gnd.n877 9.3005
R19886 gnd.n6368 gnd.n6367 9.3005
R19887 gnd.n6366 gnd.n878 9.3005
R19888 gnd.n6365 gnd.n6364 9.3005
R19889 gnd.n6363 gnd.n882 9.3005
R19890 gnd.n6362 gnd.n6361 9.3005
R19891 gnd.n6360 gnd.n883 9.3005
R19892 gnd.n6359 gnd.n6358 9.3005
R19893 gnd.n6357 gnd.n887 9.3005
R19894 gnd.n6356 gnd.n6355 9.3005
R19895 gnd.n6354 gnd.n888 9.3005
R19896 gnd.n6353 gnd.n6352 9.3005
R19897 gnd.n6351 gnd.n892 9.3005
R19898 gnd.n6350 gnd.n6349 9.3005
R19899 gnd.n6348 gnd.n893 9.3005
R19900 gnd.n6347 gnd.n6346 9.3005
R19901 gnd.n6345 gnd.n897 9.3005
R19902 gnd.n6344 gnd.n6343 9.3005
R19903 gnd.n6342 gnd.n898 9.3005
R19904 gnd.n6341 gnd.n6340 9.3005
R19905 gnd.n6339 gnd.n902 9.3005
R19906 gnd.n6338 gnd.n6337 9.3005
R19907 gnd.n6336 gnd.n903 9.3005
R19908 gnd.n6335 gnd.n6334 9.3005
R19909 gnd.n6333 gnd.n907 9.3005
R19910 gnd.n6332 gnd.n6331 9.3005
R19911 gnd.n6330 gnd.n908 9.3005
R19912 gnd.n6329 gnd.n6328 9.3005
R19913 gnd.n6327 gnd.n912 9.3005
R19914 gnd.n6326 gnd.n6325 9.3005
R19915 gnd.n6324 gnd.n913 9.3005
R19916 gnd.n6323 gnd.n6322 9.3005
R19917 gnd.n6321 gnd.n917 9.3005
R19918 gnd.n6320 gnd.n6319 9.3005
R19919 gnd.n6318 gnd.n918 9.3005
R19920 gnd.n6317 gnd.n6316 9.3005
R19921 gnd.n6315 gnd.n922 9.3005
R19922 gnd.n6314 gnd.n6313 9.3005
R19923 gnd.n6312 gnd.n923 9.3005
R19924 gnd.n6311 gnd.n6310 9.3005
R19925 gnd.n6309 gnd.n927 9.3005
R19926 gnd.n6308 gnd.n6307 9.3005
R19927 gnd.n6306 gnd.n928 9.3005
R19928 gnd.n6305 gnd.n6304 9.3005
R19929 gnd.n6303 gnd.n932 9.3005
R19930 gnd.n6302 gnd.n6301 9.3005
R19931 gnd.n6300 gnd.n933 9.3005
R19932 gnd.n6299 gnd.n6298 9.3005
R19933 gnd.n6297 gnd.n937 9.3005
R19934 gnd.n6296 gnd.n6295 9.3005
R19935 gnd.n6294 gnd.n938 9.3005
R19936 gnd.n6293 gnd.n6292 9.3005
R19937 gnd.n6291 gnd.n942 9.3005
R19938 gnd.n6290 gnd.n6289 9.3005
R19939 gnd.n6288 gnd.n943 9.3005
R19940 gnd.n6287 gnd.n6286 9.3005
R19941 gnd.n6285 gnd.n947 9.3005
R19942 gnd.n6284 gnd.n6283 9.3005
R19943 gnd.n6282 gnd.n948 9.3005
R19944 gnd.n6281 gnd.n6280 9.3005
R19945 gnd.n6279 gnd.n952 9.3005
R19946 gnd.n6278 gnd.n6277 9.3005
R19947 gnd.n6276 gnd.n953 9.3005
R19948 gnd.n6275 gnd.n6274 9.3005
R19949 gnd.n6273 gnd.n957 9.3005
R19950 gnd.n6272 gnd.n6271 9.3005
R19951 gnd.n6270 gnd.n958 9.3005
R19952 gnd.n6269 gnd.n6268 9.3005
R19953 gnd.n6267 gnd.n962 9.3005
R19954 gnd.n6266 gnd.n6265 9.3005
R19955 gnd.n6264 gnd.n963 9.3005
R19956 gnd.n6263 gnd.n6262 9.3005
R19957 gnd.n6261 gnd.n967 9.3005
R19958 gnd.n6260 gnd.n6259 9.3005
R19959 gnd.n6258 gnd.n968 9.3005
R19960 gnd.n6257 gnd.n6256 9.3005
R19961 gnd.n6255 gnd.n972 9.3005
R19962 gnd.n6254 gnd.n6253 9.3005
R19963 gnd.n6252 gnd.n973 9.3005
R19964 gnd.n6251 gnd.n6250 9.3005
R19965 gnd.n6249 gnd.n977 9.3005
R19966 gnd.n6248 gnd.n6247 9.3005
R19967 gnd.n6246 gnd.n978 9.3005
R19968 gnd.n6245 gnd.n6244 9.3005
R19969 gnd.n6243 gnd.n982 9.3005
R19970 gnd.n6242 gnd.n6241 9.3005
R19971 gnd.n6240 gnd.n983 9.3005
R19972 gnd.n6239 gnd.n6238 9.3005
R19973 gnd.n6237 gnd.n987 9.3005
R19974 gnd.n6236 gnd.n6235 9.3005
R19975 gnd.n6234 gnd.n988 9.3005
R19976 gnd.n6233 gnd.n6232 9.3005
R19977 gnd.n6231 gnd.n992 9.3005
R19978 gnd.n6383 gnd.n6382 9.3005
R19979 gnd.n2164 gnd.n867 9.3005
R19980 gnd.n4438 gnd.n4437 9.3005
R19981 gnd.n4436 gnd.n2267 9.3005
R19982 gnd.n2243 gnd.n2242 9.3005
R19983 gnd.n4468 gnd.n4467 9.3005
R19984 gnd.n4469 gnd.n2240 9.3005
R19985 gnd.n4472 gnd.n4471 9.3005
R19986 gnd.n4470 gnd.n2241 9.3005
R19987 gnd.n2217 gnd.n2216 9.3005
R19988 gnd.n4502 gnd.n4501 9.3005
R19989 gnd.n4503 gnd.n2214 9.3005
R19990 gnd.n4506 gnd.n4505 9.3005
R19991 gnd.n4504 gnd.n2215 9.3005
R19992 gnd.n2191 gnd.n2190 9.3005
R19993 gnd.n4538 gnd.n4537 9.3005
R19994 gnd.n4539 gnd.n2188 9.3005
R19995 gnd.n4545 gnd.n4544 9.3005
R19996 gnd.n4543 gnd.n2189 9.3005
R19997 gnd.n4542 gnd.n4541 9.3005
R19998 gnd.n2180 gnd.n2179 9.3005
R19999 gnd.n4561 gnd.n4560 9.3005
R20000 gnd.n4562 gnd.n2178 9.3005
R20001 gnd.n4564 gnd.n4563 9.3005
R20002 gnd.n2175 gnd.n2174 9.3005
R20003 gnd.n4911 gnd.n4910 9.3005
R20004 gnd.n4912 gnd.n2173 9.3005
R20005 gnd.n4914 gnd.n4913 9.3005
R20006 gnd.n2170 gnd.n2169 9.3005
R20007 gnd.n4931 gnd.n4930 9.3005
R20008 gnd.n4932 gnd.n2167 9.3005
R20009 gnd.n4934 gnd.n4933 9.3005
R20010 gnd.n4935 gnd.n2166 9.3005
R20011 gnd.n4937 gnd.n4936 9.3005
R20012 gnd.n4990 gnd.n4989 9.3005
R20013 gnd.n2083 gnd.n2082 9.3005
R20014 gnd.n4984 gnd.n4983 9.3005
R20015 gnd.n4982 gnd.n4981 9.3005
R20016 gnd.n2099 gnd.n2098 9.3005
R20017 gnd.n4976 gnd.n4975 9.3005
R20018 gnd.n4974 gnd.n4973 9.3005
R20019 gnd.n2112 gnd.n2111 9.3005
R20020 gnd.n4968 gnd.n4967 9.3005
R20021 gnd.n4966 gnd.n4965 9.3005
R20022 gnd.n2125 gnd.n2124 9.3005
R20023 gnd.n4960 gnd.n4959 9.3005
R20024 gnd.n4958 gnd.n4957 9.3005
R20025 gnd.n2138 gnd.n2137 9.3005
R20026 gnd.n4952 gnd.n4951 9.3005
R20027 gnd.n4950 gnd.n4949 9.3005
R20028 gnd.n2153 gnd.n2152 9.3005
R20029 gnd.n4944 gnd.n4943 9.3005
R20030 gnd.n4992 gnd.n4991 9.3005
R20031 gnd.n4939 gnd.n2165 9.3005
R20032 gnd.n4946 gnd.n4945 9.3005
R20033 gnd.n4948 gnd.n4947 9.3005
R20034 gnd.n2144 gnd.n2143 9.3005
R20035 gnd.n4954 gnd.n4953 9.3005
R20036 gnd.n4956 gnd.n4955 9.3005
R20037 gnd.n2132 gnd.n2131 9.3005
R20038 gnd.n4962 gnd.n4961 9.3005
R20039 gnd.n4964 gnd.n4963 9.3005
R20040 gnd.n2118 gnd.n2117 9.3005
R20041 gnd.n4970 gnd.n4969 9.3005
R20042 gnd.n4972 gnd.n4971 9.3005
R20043 gnd.n2106 gnd.n2105 9.3005
R20044 gnd.n4978 gnd.n4977 9.3005
R20045 gnd.n4980 gnd.n4979 9.3005
R20046 gnd.n2092 gnd.n2091 9.3005
R20047 gnd.n4986 gnd.n4985 9.3005
R20048 gnd.n4988 gnd.n4987 9.3005
R20049 gnd.n2084 gnd.n2079 9.3005
R20050 gnd.n4993 gnd.n2078 9.3005
R20051 gnd.n4995 gnd.n4994 9.3005
R20052 gnd.n4997 gnd.n4996 9.3005
R20053 gnd.n4998 gnd.n2071 9.3005
R20054 gnd.n5000 gnd.n4999 9.3005
R20055 gnd.n5001 gnd.n2070 9.3005
R20056 gnd.n5003 gnd.n5002 9.3005
R20057 gnd.n2068 gnd.n2067 9.3005
R20058 gnd.n5009 gnd.n5008 9.3005
R20059 gnd.n5012 gnd.n5011 9.3005
R20060 gnd.n2065 gnd.n2064 9.3005
R20061 gnd.n5026 gnd.n5025 9.3005
R20062 gnd.n5027 gnd.n2063 9.3005
R20063 gnd.n5029 gnd.n5028 9.3005
R20064 gnd.n2054 gnd.n2053 9.3005
R20065 gnd.n5044 gnd.n5043 9.3005
R20066 gnd.n5045 gnd.n2052 9.3005
R20067 gnd.n5047 gnd.n5046 9.3005
R20068 gnd.n2042 gnd.n2041 9.3005
R20069 gnd.n5061 gnd.n5060 9.3005
R20070 gnd.n5062 gnd.n2040 9.3005
R20071 gnd.n5064 gnd.n5063 9.3005
R20072 gnd.n2029 gnd.n2028 9.3005
R20073 gnd.n5080 gnd.n5079 9.3005
R20074 gnd.n5081 gnd.n2026 9.3005
R20075 gnd.n5147 gnd.n5146 9.3005
R20076 gnd.n5145 gnd.n2027 9.3005
R20077 gnd.n5144 gnd.n5143 9.3005
R20078 gnd.n5142 gnd.n5082 9.3005
R20079 gnd.n5141 gnd.n5140 9.3005
R20080 gnd.n5139 gnd.n5085 9.3005
R20081 gnd.n5138 gnd.n5137 9.3005
R20082 gnd.n5136 gnd.n5086 9.3005
R20083 gnd.n5135 gnd.n5134 9.3005
R20084 gnd.n5133 gnd.n5090 9.3005
R20085 gnd.n5132 gnd.n5131 9.3005
R20086 gnd.n5130 gnd.n5091 9.3005
R20087 gnd.n5129 gnd.n5128 9.3005
R20088 gnd.n5127 gnd.n5094 9.3005
R20089 gnd.n5126 gnd.n5125 9.3005
R20090 gnd.n5124 gnd.n5095 9.3005
R20091 gnd.n5123 gnd.n5122 9.3005
R20092 gnd.n5121 gnd.n5098 9.3005
R20093 gnd.n5120 gnd.n5119 9.3005
R20094 gnd.n5118 gnd.n5099 9.3005
R20095 gnd.n5117 gnd.n5116 9.3005
R20096 gnd.n5115 gnd.n5102 9.3005
R20097 gnd.n5114 gnd.n5113 9.3005
R20098 gnd.n5112 gnd.n5103 9.3005
R20099 gnd.n5111 gnd.n5110 9.3005
R20100 gnd.n5109 gnd.n5106 9.3005
R20101 gnd.n5108 gnd.n5107 9.3005
R20102 gnd.n1492 gnd.n1491 9.3005
R20103 gnd.n5371 gnd.n5370 9.3005
R20104 gnd.n5372 gnd.n1489 9.3005
R20105 gnd.n5388 gnd.n5387 9.3005
R20106 gnd.n5386 gnd.n1490 9.3005
R20107 gnd.n5385 gnd.n5384 9.3005
R20108 gnd.n5383 gnd.n5373 9.3005
R20109 gnd.n5382 gnd.n5381 9.3005
R20110 gnd.n5380 gnd.n5377 9.3005
R20111 gnd.n5379 gnd.n5378 9.3005
R20112 gnd.n1442 gnd.n1441 9.3005
R20113 gnd.n5468 gnd.n5467 9.3005
R20114 gnd.n5469 gnd.n1439 9.3005
R20115 gnd.n5482 gnd.n5481 9.3005
R20116 gnd.n5480 gnd.n1440 9.3005
R20117 gnd.n5479 gnd.n5478 9.3005
R20118 gnd.n5477 gnd.n5470 9.3005
R20119 gnd.n5476 gnd.n5475 9.3005
R20120 gnd.n5474 gnd.n5473 9.3005
R20121 gnd.n1392 gnd.n1391 9.3005
R20122 gnd.n5544 gnd.n5543 9.3005
R20123 gnd.n5545 gnd.n1389 9.3005
R20124 gnd.n5551 gnd.n5550 9.3005
R20125 gnd.n5549 gnd.n1390 9.3005
R20126 gnd.n5548 gnd.n5547 9.3005
R20127 gnd.n5546 gnd.n1367 9.3005
R20128 gnd.n5587 gnd.n1366 9.3005
R20129 gnd.n5589 gnd.n5588 9.3005
R20130 gnd.n5590 gnd.n1364 9.3005
R20131 gnd.n5611 gnd.n5610 9.3005
R20132 gnd.n5609 gnd.n1365 9.3005
R20133 gnd.n5608 gnd.n5607 9.3005
R20134 gnd.n5606 gnd.n5591 9.3005
R20135 gnd.n5605 gnd.n5604 9.3005
R20136 gnd.n5603 gnd.n5595 9.3005
R20137 gnd.n5602 gnd.n5601 9.3005
R20138 gnd.n5600 gnd.n5596 9.3005
R20139 gnd.n5599 gnd.n5598 9.3005
R20140 gnd.n1217 gnd.n1216 9.3005
R20141 gnd.n5821 gnd.n5820 9.3005
R20142 gnd.n5822 gnd.n1215 9.3005
R20143 gnd.n5824 gnd.n5823 9.3005
R20144 gnd.n1206 gnd.n1205 9.3005
R20145 gnd.n5838 gnd.n5837 9.3005
R20146 gnd.n5839 gnd.n1204 9.3005
R20147 gnd.n5841 gnd.n5840 9.3005
R20148 gnd.n1194 gnd.n1193 9.3005
R20149 gnd.n5855 gnd.n5854 9.3005
R20150 gnd.n5856 gnd.n1192 9.3005
R20151 gnd.n5858 gnd.n5857 9.3005
R20152 gnd.n1183 gnd.n1182 9.3005
R20153 gnd.n5873 gnd.n5872 9.3005
R20154 gnd.n5874 gnd.n1181 9.3005
R20155 gnd.n5876 gnd.n5875 9.3005
R20156 gnd.n1171 gnd.n1170 9.3005
R20157 gnd.n5892 gnd.n5891 9.3005
R20158 gnd.n5893 gnd.n1169 9.3005
R20159 gnd.n5913 gnd.n5912 9.3005
R20160 gnd.n5010 gnd.n2066 9.3005
R20161 gnd.n5909 gnd.n5894 9.3005
R20162 gnd.n5908 gnd.n5907 9.3005
R20163 gnd.n5906 gnd.n5897 9.3005
R20164 gnd.n5905 gnd.n5904 9.3005
R20165 gnd.n5903 gnd.n5898 9.3005
R20166 gnd.n1141 gnd.n1139 9.3005
R20167 gnd.n5911 gnd.n5910 9.3005
R20168 gnd.n6222 gnd.n6221 9.3005
R20169 gnd.n1020 gnd.n1018 9.3005
R20170 gnd.n6058 gnd.n6057 9.3005
R20171 gnd.n6060 gnd.n6059 9.3005
R20172 gnd.n6047 gnd.n6046 9.3005
R20173 gnd.n6066 gnd.n6065 9.3005
R20174 gnd.n6068 gnd.n6067 9.3005
R20175 gnd.n6037 gnd.n6036 9.3005
R20176 gnd.n6074 gnd.n6073 9.3005
R20177 gnd.n6076 gnd.n6075 9.3005
R20178 gnd.n6027 gnd.n6026 9.3005
R20179 gnd.n6082 gnd.n6081 9.3005
R20180 gnd.n6084 gnd.n6083 9.3005
R20181 gnd.n6017 gnd.n6016 9.3005
R20182 gnd.n6090 gnd.n6089 9.3005
R20183 gnd.n6092 gnd.n6091 9.3005
R20184 gnd.n6013 gnd.n1147 9.3005
R20185 gnd.n6220 gnd.n1029 9.3005
R20186 gnd.n1024 gnd.n1022 9.3005
R20187 gnd.n6097 gnd.n6096 9.3005
R20188 gnd.n6095 gnd.n1140 9.3005
R20189 gnd.n6094 gnd.n6093 9.3005
R20190 gnd.n1148 gnd.n1146 9.3005
R20191 gnd.n6088 gnd.n6087 9.3005
R20192 gnd.n6086 gnd.n6085 9.3005
R20193 gnd.n6021 gnd.n6020 9.3005
R20194 gnd.n6080 gnd.n6079 9.3005
R20195 gnd.n6078 gnd.n6077 9.3005
R20196 gnd.n6033 gnd.n6032 9.3005
R20197 gnd.n6072 gnd.n6071 9.3005
R20198 gnd.n6070 gnd.n6069 9.3005
R20199 gnd.n6041 gnd.n6040 9.3005
R20200 gnd.n6064 gnd.n6063 9.3005
R20201 gnd.n6062 gnd.n6061 9.3005
R20202 gnd.n6053 gnd.n6052 9.3005
R20203 gnd.n6056 gnd.n1014 9.3005
R20204 gnd.n6224 gnd.n6223 9.3005
R20205 gnd.n1025 gnd.n1019 9.3005
R20206 gnd.n1028 gnd.n1027 9.3005
R20207 gnd.n1023 gnd.n994 9.3005
R20208 gnd.n5970 gnd.n5969 9.3005
R20209 gnd.n5973 gnd.n5966 9.3005
R20210 gnd.n5975 gnd.n5974 9.3005
R20211 gnd.n5976 gnd.n5964 9.3005
R20212 gnd.n5979 gnd.n5978 9.3005
R20213 gnd.n5977 gnd.n5965 9.3005
R20214 gnd.n379 gnd.n378 9.3005
R20215 gnd.n7064 gnd.n7063 9.3005
R20216 gnd.n7065 gnd.n376 9.3005
R20217 gnd.n7068 gnd.n7067 9.3005
R20218 gnd.n7066 gnd.n377 9.3005
R20219 gnd.n350 gnd.n349 9.3005
R20220 gnd.n7100 gnd.n7099 9.3005
R20221 gnd.n7101 gnd.n347 9.3005
R20222 gnd.n7124 gnd.n7123 9.3005
R20223 gnd.n7122 gnd.n348 9.3005
R20224 gnd.n7121 gnd.n7120 9.3005
R20225 gnd.n7119 gnd.n7102 9.3005
R20226 gnd.n7118 gnd.n7117 9.3005
R20227 gnd.n7116 gnd.n7105 9.3005
R20228 gnd.n7115 gnd.n7114 9.3005
R20229 gnd.n7113 gnd.n7106 9.3005
R20230 gnd.n7112 gnd.n7111 9.3005
R20231 gnd.n7110 gnd.n7109 9.3005
R20232 gnd.n288 gnd.n287 9.3005
R20233 gnd.n7194 gnd.n7193 9.3005
R20234 gnd.n7195 gnd.n285 9.3005
R20235 gnd.n7202 gnd.n7201 9.3005
R20236 gnd.n7200 gnd.n286 9.3005
R20237 gnd.n7199 gnd.n7198 9.3005
R20238 gnd.n7197 gnd.n99 9.3005
R20239 gnd.n5968 gnd.n5967 9.3005
R20240 gnd.n7740 gnd.n100 9.3005
R20241 gnd.n3071 gnd.t31 9.29782
R20242 gnd.n2771 gnd.t195 9.29782
R20243 gnd.n7126 gnd.t218 9.24152
R20244 gnd.t270 gnd.n178 9.24152
R20245 gnd.n3062 gnd.t31 8.93321
R20246 gnd.t135 gnd.n2493 8.93321
R20247 gnd.t107 gnd.n2494 8.93321
R20248 gnd.n1614 gnd.t114 8.92286
R20249 gnd.n5193 gnd.n1608 8.92286
R20250 gnd.n1603 gnd.t104 8.92286
R20251 gnd.n5219 gnd.t9 8.92286
R20252 gnd.n5312 gnd.n1521 8.92286
R20253 gnd.n5368 gnd.n1494 8.92286
R20254 gnd.n5421 gnd.n5420 8.92286
R20255 gnd.n5531 gnd.n1402 8.92286
R20256 gnd.n1334 gnd.t160 8.92286
R20257 gnd.n5671 gnd.n5670 8.92286
R20258 gnd.t91 gnd.n1219 8.92286
R20259 gnd.n3774 gnd.n3749 8.92171
R20260 gnd.n3742 gnd.n3717 8.92171
R20261 gnd.n3710 gnd.n3685 8.92171
R20262 gnd.n3679 gnd.n3654 8.92171
R20263 gnd.n3647 gnd.n3622 8.92171
R20264 gnd.n3615 gnd.n3590 8.92171
R20265 gnd.n3583 gnd.n3558 8.92171
R20266 gnd.n3552 gnd.n3527 8.92171
R20267 gnd.n1250 gnd.n1232 8.72777
R20268 gnd.t249 gnd.n216 8.60421
R20269 gnd.n3430 gnd.t190 8.56861
R20270 gnd.n2682 gnd.n2662 8.43656
R20271 gnd.n58 gnd.n38 8.43656
R20272 gnd.t180 gnd.n2536 8.20401
R20273 gnd.n3508 gnd.t183 8.20401
R20274 gnd.n3775 gnd.n3747 8.14595
R20275 gnd.n3743 gnd.n3715 8.14595
R20276 gnd.n3711 gnd.n3683 8.14595
R20277 gnd.n3680 gnd.n3652 8.14595
R20278 gnd.n3648 gnd.n3620 8.14595
R20279 gnd.n3616 gnd.n3588 8.14595
R20280 gnd.n3584 gnd.n3556 8.14595
R20281 gnd.n3553 gnd.n3525 8.14595
R20282 gnd.n4435 gnd.n0 8.10675
R20283 gnd.n7741 gnd.n7740 8.10675
R20284 gnd.n6453 gnd.t308 8.00176
R20285 gnd.n3780 gnd.n3779 7.97301
R20286 gnd.n6391 gnd.n853 7.9669
R20287 gnd.n6226 gnd.n1011 7.9669
R20288 gnd.n7741 gnd.n98 7.95236
R20289 gnd.n3218 gnd.t149 7.83941
R20290 gnd.n6452 gnd.n753 7.83941
R20291 gnd.n6220 gnd.n1022 7.75808
R20292 gnd.n7398 gnd.n7320 7.75808
R20293 gnd.n4943 gnd.n2152 7.75808
R20294 gnd.n4214 gnd.n4148 7.75808
R20295 gnd.n3136 gnd.n2874 7.65711
R20296 gnd.n765 gnd.n752 7.64824
R20297 gnd.n6446 gnd.n768 7.64824
R20298 gnd.n4558 gnd.n777 7.64824
R20299 gnd.n6440 gnd.n780 7.64824
R20300 gnd.n4902 gnd.n4901 7.64824
R20301 gnd.n6434 gnd.n790 7.64824
R20302 gnd.n4908 gnd.n797 7.64824
R20303 gnd.n6428 gnd.n800 7.64824
R20304 gnd.n4916 gnd.n808 7.64824
R20305 gnd.n6422 gnd.n811 7.64824
R20306 gnd.n4928 gnd.n818 7.64824
R20307 gnd.n6416 gnd.n821 7.64824
R20308 gnd.n6410 gnd.n832 7.64824
R20309 gnd.n6400 gnd.n6399 7.64824
R20310 gnd.n5179 gnd.n1621 7.64824
R20311 gnd.n5292 gnd.n1536 7.64824
R20312 gnd.n5324 gnd.t23 7.64824
R20313 gnd.n5391 gnd.n5390 7.64824
R20314 gnd.n5435 gnd.n1455 7.64824
R20315 gnd.t7 gnd.n1444 7.64824
R20316 gnd.n5541 gnd.n1394 7.64824
R20317 gnd.n6010 gnd.n1151 7.64824
R20318 gnd.n6009 gnd.n1155 7.64824
R20319 gnd.n6003 gnd.n6002 7.64824
R20320 gnd.n5988 gnd.n5939 7.64824
R20321 gnd.n5981 gnd.n5949 7.64824
R20322 gnd.n7051 gnd.n391 7.64824
R20323 gnd.n7038 gnd.n7037 7.64824
R20324 gnd.n7061 gnd.n381 7.64824
R20325 gnd.n7044 gnd.n383 7.64824
R20326 gnd.n7070 gnd.n374 7.64824
R20327 gnd.n7087 gnd.n362 7.64824
R20328 gnd.n7074 gnd.n365 7.64824
R20329 gnd.n7097 gnd.n352 7.64824
R20330 gnd.n7080 gnd.n354 7.64824
R20331 gnd.n2723 gnd.n2722 7.53171
R20332 gnd.n5015 gnd.t75 7.32958
R20333 gnd.n5058 gnd.t158 7.32958
R20334 gnd.n1621 gnd.t178 7.32958
R20335 gnd.n5678 gnd.t167 7.32958
R20336 gnd.t161 gnd.n1196 7.32958
R20337 gnd.n5889 gnd.t39 7.32958
R20338 gnd.n1650 gnd.n1649 7.30353
R20339 gnd.n1249 gnd.n1248 7.30353
R20340 gnd.n2380 gnd.t285 7.11021
R20341 gnd.t8 gnd.n5227 7.01093
R20342 gnd.n5339 gnd.t19 7.01093
R20343 gnd.n5486 gnd.t170 7.01093
R20344 gnd.n5614 gnd.t6 7.01093
R20345 gnd.n2344 gnd.t260 6.74561
R20346 gnd.t294 gnd.n2185 6.74561
R20347 gnd.n5357 gnd.t198 6.69227
R20348 gnd.t208 gnd.n1431 6.69227
R20349 gnd.n5738 gnd.n5737 6.5566
R20350 gnd.n1962 gnd.n1961 6.5566
R20351 gnd.n1745 gnd.n1691 6.5566
R20352 gnd.n5750 gnd.n1278 6.5566
R20353 gnd.n3206 gnd.t149 6.38101
R20354 gnd.n2307 gnd.t276 6.38101
R20355 gnd.n4489 gnd.t258 6.38101
R20356 gnd.n5160 gnd.n5159 6.37362
R20357 gnd.t114 gnd.t97 6.37362
R20358 gnd.n1552 gnd.n1541 6.37362
R20359 gnd.n5346 gnd.t12 6.37362
R20360 gnd.n5327 gnd.n1472 6.37362
R20361 gnd.n5442 gnd.n1460 6.37362
R20362 gnd.t177 gnd.n1422 6.37362
R20363 gnd.n5553 gnd.n1387 6.37362
R20364 gnd.n5670 gnd.t28 6.37362
R20365 gnd.n5644 gnd.t28 6.37362
R20366 gnd.n5818 gnd.n1219 6.37362
R20367 gnd.n4947 gnd.n2156 6.20656
R20368 gnd.n1025 gnd.n1017 6.20656
R20369 gnd.t15 gnd.n5275 6.05496
R20370 gnd.t151 gnd.t13 6.05496
R20371 gnd.t2 gnd.t210 6.05496
R20372 gnd.n5554 gnd.t163 6.05496
R20373 gnd.n3125 gnd.t173 6.01641
R20374 gnd.n2538 gnd.t180 6.01641
R20375 gnd.n3491 gnd.t183 6.01641
R20376 gnd.n4431 gnd.t222 6.01641
R20377 gnd.n4440 gnd.t290 6.01641
R20378 gnd.n3777 gnd.n3747 5.81868
R20379 gnd.n3745 gnd.n3715 5.81868
R20380 gnd.n3713 gnd.n3683 5.81868
R20381 gnd.n3682 gnd.n3652 5.81868
R20382 gnd.n3650 gnd.n3620 5.81868
R20383 gnd.n3618 gnd.n3588 5.81868
R20384 gnd.n3586 gnd.n3556 5.81868
R20385 gnd.n3555 gnd.n3525 5.81868
R20386 gnd.n5660 gnd.t43 5.73631
R20387 gnd.t190 gnd.n2555 5.65181
R20388 gnd.t224 gnd.n2304 5.65181
R20389 gnd.n4499 gnd.t226 5.65181
R20390 gnd.n1280 gnd.n1101 5.62001
R20391 gnd.n1957 gnd.n1954 5.62001
R20392 gnd.n1954 gnd.n1749 5.62001
R20393 gnd.n5748 gnd.n1101 5.62001
R20394 gnd.n3006 gnd.n3001 5.4308
R20395 gnd.n3822 gnd.n2479 5.4308
R20396 gnd.t192 gnd.n2602 5.28721
R20397 gnd.n2504 gnd.t135 5.28721
R20398 gnd.n3804 gnd.t107 5.28721
R20399 gnd.t232 gnd.n2341 5.28721
R20400 gnd.t308 gnd.n6452 5.28721
R20401 gnd.t156 gnd.t192 5.10491
R20402 gnd.n5249 gnd.t11 5.09899
R20403 gnd.n5269 gnd.n1557 5.09899
R20404 gnd.n5408 gnd.n1465 5.09899
R20405 gnd.n5415 gnd.n1467 5.09899
R20406 gnd.n1379 gnd.n1378 5.09899
R20407 gnd.n5620 gnd.t3 5.09899
R20408 gnd.n3775 gnd.n3774 5.04292
R20409 gnd.n3743 gnd.n3742 5.04292
R20410 gnd.n3711 gnd.n3710 5.04292
R20411 gnd.n3680 gnd.n3679 5.04292
R20412 gnd.n3648 gnd.n3647 5.04292
R20413 gnd.n3616 gnd.n3615 5.04292
R20414 gnd.n3584 gnd.n3583 5.04292
R20415 gnd.n3553 gnd.n3552 5.04292
R20416 gnd.n3278 gnd.t195 4.92261
R20417 gnd.t220 gnd.n2377 4.92261
R20418 gnd.t21 gnd.n1654 4.78034
R20419 gnd.n1253 gnd.t68 4.78034
R20420 gnd.n5827 gnd.t17 4.78034
R20421 gnd.n2727 gnd.n2724 4.74817
R20422 gnd.n2777 gnd.n2643 4.74817
R20423 gnd.n2764 gnd.n2642 4.74817
R20424 gnd.n2641 gnd.n2640 4.74817
R20425 gnd.n2773 gnd.n2724 4.74817
R20426 gnd.n2774 gnd.n2643 4.74817
R20427 gnd.n2776 gnd.n2642 4.74817
R20428 gnd.n2763 gnd.n2641 4.74817
R20429 gnd.n2722 gnd.n2721 4.74296
R20430 gnd.n98 gnd.n97 4.74296
R20431 gnd.n2682 gnd.n2681 4.7074
R20432 gnd.n2702 gnd.n2701 4.7074
R20433 gnd.n58 gnd.n57 4.7074
R20434 gnd.n78 gnd.n77 4.7074
R20435 gnd.n2722 gnd.n2702 4.65959
R20436 gnd.n98 gnd.n78 4.65959
R20437 gnd.n6162 gnd.n1103 4.6132
R20438 gnd.n1952 gnd.n1951 4.6132
R20439 gnd.t196 gnd.n2793 4.55801
R20440 gnd.n5310 gnd.t1 4.46168
R20441 gnd.t4 gnd.n1418 4.46168
R20442 gnd.n5810 gnd.t142 4.46168
R20443 gnd.n1245 gnd.n1232 4.46111
R20444 gnd.n3760 gnd.n3756 4.38594
R20445 gnd.n3728 gnd.n3724 4.38594
R20446 gnd.n3696 gnd.n3692 4.38594
R20447 gnd.n3665 gnd.n3661 4.38594
R20448 gnd.n3633 gnd.n3629 4.38594
R20449 gnd.n3601 gnd.n3597 4.38594
R20450 gnd.n3569 gnd.n3565 4.38594
R20451 gnd.n3538 gnd.n3534 4.38594
R20452 gnd.n3771 gnd.n3749 4.26717
R20453 gnd.n3739 gnd.n3717 4.26717
R20454 gnd.n3707 gnd.n3685 4.26717
R20455 gnd.n3676 gnd.n3654 4.26717
R20456 gnd.n3644 gnd.n3622 4.26717
R20457 gnd.n3612 gnd.n3590 4.26717
R20458 gnd.n3580 gnd.n3558 4.26717
R20459 gnd.n3549 gnd.n3527 4.26717
R20460 gnd.n3187 gnd.t185 4.19341
R20461 gnd.t64 gnd.n829 4.14303
R20462 gnd.t35 gnd.n5935 4.14303
R20463 gnd.n3779 gnd.n3778 4.08274
R20464 gnd.n5737 gnd.n5736 4.05904
R20465 gnd.n1963 gnd.n1962 4.05904
R20466 gnd.n1742 gnd.n1691 4.05904
R20467 gnd.n1278 gnd.n1273 4.05904
R20468 gnd.n3147 gnd.n2866 4.01111
R20469 gnd.n2869 gnd.n2867 4.01111
R20470 gnd.n3157 gnd.n3156 4.01111
R20471 gnd.n3168 gnd.n2850 4.01111
R20472 gnd.n3167 gnd.n2853 4.01111
R20473 gnd.n3178 gnd.n2841 4.01111
R20474 gnd.n2844 gnd.n2842 4.01111
R20475 gnd.n3188 gnd.n3187 4.01111
R20476 gnd.n3198 gnd.n2822 4.01111
R20477 gnd.n3197 gnd.n2825 4.01111
R20478 gnd.n3206 gnd.n2816 4.01111
R20479 gnd.n3218 gnd.n2806 4.01111
R20480 gnd.n3228 gnd.n2791 4.01111
R20481 gnd.n3244 gnd.n3243 4.01111
R20482 gnd.n2793 gnd.n2730 4.01111
R20483 gnd.n3298 gnd.n2731 4.01111
R20484 gnd.n3292 gnd.n3291 4.01111
R20485 gnd.n2780 gnd.n2742 4.01111
R20486 gnd.n3284 gnd.n2753 4.01111
R20487 gnd.n2771 gnd.n2766 4.01111
R20488 gnd.n3278 gnd.n3277 4.01111
R20489 gnd.n3324 gnd.n2637 4.01111
R20490 gnd.n3323 gnd.n3322 4.01111
R20491 gnd.n3335 gnd.n3334 4.01111
R20492 gnd.n2630 gnd.n2622 4.01111
R20493 gnd.n3364 gnd.n2610 4.01111
R20494 gnd.n3363 gnd.n2613 4.01111
R20495 gnd.n3374 gnd.n2602 4.01111
R20496 gnd.n2603 gnd.n2591 4.01111
R20497 gnd.n3385 gnd.n2592 4.01111
R20498 gnd.n3409 gnd.n2583 4.01111
R20499 gnd.n3408 gnd.n2574 4.01111
R20500 gnd.n3431 gnd.n3430 4.01111
R20501 gnd.n3449 gnd.n2555 4.01111
R20502 gnd.n3448 gnd.n2558 4.01111
R20503 gnd.n3459 gnd.n2547 4.01111
R20504 gnd.n2548 gnd.n2535 4.01111
R20505 gnd.n3470 gnd.n2536 4.01111
R20506 gnd.n3497 gnd.n2520 4.01111
R20507 gnd.n3509 gnd.n3508 4.01111
R20508 gnd.n3491 gnd.n2513 4.01111
R20509 gnd.n3520 gnd.n3519 4.01111
R20510 gnd.n3792 gnd.n2501 4.01111
R20511 gnd.n3791 gnd.n2504 4.01111
R20512 gnd.n3804 gnd.n2493 4.01111
R20513 gnd.n2494 gnd.n2486 4.01111
R20514 gnd.n3814 gnd.n2412 4.01111
R20515 gnd.n19 gnd.n9 3.99943
R20516 gnd.n2825 gnd.t188 3.82881
R20517 gnd.n2613 gnd.t156 3.82881
R20518 gnd.n3498 gnd.t194 3.82881
R20519 gnd.n1630 gnd.n1618 3.82437
R20520 gnd.t97 gnd.n1612 3.82437
R20521 gnd.n5241 gnd.n1569 3.82437
R20522 gnd.n5268 gnd.t10 3.82437
R20523 gnd.n5285 gnd.n5284 3.82437
R20524 gnd.n5398 gnd.n5397 3.82437
R20525 gnd.n5455 gnd.n1452 3.82437
R20526 gnd.n5522 gnd.n1413 3.82437
R20527 gnd.t152 gnd.n5574 3.82437
R20528 gnd.n5566 gnd.n1345 3.82437
R20529 gnd.n5644 gnd.t46 3.82437
R20530 gnd.n5683 gnd.n1228 3.82437
R20531 gnd.n3302 gnd.n2723 3.81325
R20532 gnd.n2702 gnd.n2682 3.72967
R20533 gnd.n78 gnd.n58 3.72967
R20534 gnd.n3779 gnd.n3651 3.70378
R20535 gnd.n19 gnd.n18 3.60163
R20536 gnd.n4922 gnd.t64 3.50571
R20537 gnd.n5936 gnd.t35 3.50571
R20538 gnd.n7651 gnd.t53 3.50571
R20539 gnd.n3770 gnd.n3751 3.49141
R20540 gnd.n3738 gnd.n3719 3.49141
R20541 gnd.n3706 gnd.n3687 3.49141
R20542 gnd.n3675 gnd.n3656 3.49141
R20543 gnd.n3643 gnd.n3624 3.49141
R20544 gnd.n3611 gnd.n3592 3.49141
R20545 gnd.n3579 gnd.n3560 3.49141
R20546 gnd.n3548 gnd.n3529 3.49141
R20547 gnd.t175 gnd.n3254 3.46421
R20548 gnd.n3255 gnd.t187 3.46421
R20549 gnd.t24 gnd.n2637 3.46421
R20550 gnd.t182 gnd.n3419 3.46421
R20551 gnd.n7540 gnd.n7476 3.29747
R20552 gnd.n7535 gnd.n7476 3.29747
R20553 gnd.n6180 gnd.n6179 3.29747
R20554 gnd.n6179 gnd.n6178 3.29747
R20555 gnd.n4017 gnd.n3959 3.29747
R20556 gnd.n3959 gnd.n3954 3.29747
R20557 gnd.n1824 gnd.n1762 3.29747
R20558 gnd.n1827 gnd.n1762 3.29747
R20559 gnd.n5242 gnd.t20 3.18706
R20560 gnd.n5257 gnd.t20 3.18706
R20561 gnd.n5584 gnd.t0 3.18706
R20562 gnd.n5567 gnd.t0 3.18706
R20563 gnd.n5678 gnd.t142 3.18706
R20564 gnd.n3322 gnd.t197 3.0996
R20565 gnd.t184 gnd.n3345 3.0996
R20566 gnd.t212 gnd.n2567 3.0996
R20567 gnd.n5212 gnd.t202 2.8684
R20568 gnd.n5654 gnd.t165 2.8684
R20569 gnd.n2703 gnd.t340 2.82907
R20570 gnd.n2703 gnd.t413 2.82907
R20571 gnd.n2705 gnd.t295 2.82907
R20572 gnd.n2705 gnd.t396 2.82907
R20573 gnd.n2707 gnd.t227 2.82907
R20574 gnd.n2707 gnd.t369 2.82907
R20575 gnd.n2709 gnd.t400 2.82907
R20576 gnd.n2709 gnd.t292 2.82907
R20577 gnd.n2711 gnd.t326 2.82907
R20578 gnd.n2711 gnd.t304 2.82907
R20579 gnd.n2713 gnd.t303 2.82907
R20580 gnd.n2713 gnd.t273 2.82907
R20581 gnd.n2715 gnd.t312 2.82907
R20582 gnd.n2715 gnd.t356 2.82907
R20583 gnd.n2717 gnd.t363 2.82907
R20584 gnd.n2717 gnd.t313 2.82907
R20585 gnd.n2719 gnd.t349 2.82907
R20586 gnd.n2719 gnd.t246 2.82907
R20587 gnd.n2644 gnd.t346 2.82907
R20588 gnd.n2644 gnd.t366 2.82907
R20589 gnd.n2646 gnd.t379 2.82907
R20590 gnd.n2646 gnd.t403 2.82907
R20591 gnd.n2648 gnd.t336 2.82907
R20592 gnd.n2648 gnd.t352 2.82907
R20593 gnd.n2650 gnd.t367 2.82907
R20594 gnd.n2650 gnd.t259 2.82907
R20595 gnd.n2652 gnd.t351 2.82907
R20596 gnd.n2652 gnd.t345 2.82907
R20597 gnd.n2654 gnd.t385 2.82907
R20598 gnd.n2654 gnd.t380 2.82907
R20599 gnd.n2656 gnd.t282 2.82907
R20600 gnd.n2656 gnd.t360 2.82907
R20601 gnd.n2658 gnd.t401 2.82907
R20602 gnd.n2658 gnd.t261 2.82907
R20603 gnd.n2660 gnd.t286 2.82907
R20604 gnd.n2660 gnd.t376 2.82907
R20605 gnd.n2663 gnd.t330 2.82907
R20606 gnd.n2663 gnd.t317 2.82907
R20607 gnd.n2665 gnd.t297 2.82907
R20608 gnd.n2665 gnd.t343 2.82907
R20609 gnd.n2667 gnd.t289 2.82907
R20610 gnd.n2667 gnd.t331 2.82907
R20611 gnd.n2669 gnd.t332 2.82907
R20612 gnd.n2669 gnd.t306 2.82907
R20613 gnd.n2671 gnd.t223 2.82907
R20614 gnd.n2671 gnd.t291 2.82907
R20615 gnd.n2673 gnd.t277 2.82907
R20616 gnd.n2673 gnd.t334 2.82907
R20617 gnd.n2675 gnd.t264 2.82907
R20618 gnd.n2675 gnd.t225 2.82907
R20619 gnd.n2677 gnd.t238 2.82907
R20620 gnd.n2677 gnd.t287 2.82907
R20621 gnd.n2679 gnd.t288 2.82907
R20622 gnd.n2679 gnd.t257 2.82907
R20623 gnd.n2683 gnd.t388 2.82907
R20624 gnd.n2683 gnd.t328 2.82907
R20625 gnd.n2685 gnd.t359 2.82907
R20626 gnd.n2685 gnd.t309 2.82907
R20627 gnd.n2687 gnd.t339 2.82907
R20628 gnd.n2687 gnd.t243 2.82907
R20629 gnd.n2689 gnd.t315 2.82907
R20630 gnd.n2689 gnd.t357 2.82907
R20631 gnd.n2691 gnd.t377 2.82907
R20632 gnd.n2691 gnd.t364 2.82907
R20633 gnd.n2693 gnd.t361 2.82907
R20634 gnd.n2693 gnd.t350 2.82907
R20635 gnd.n2695 gnd.t368 2.82907
R20636 gnd.n2695 gnd.t408 2.82907
R20637 gnd.n2697 gnd.t233 2.82907
R20638 gnd.n2697 gnd.t370 2.82907
R20639 gnd.n2699 gnd.t402 2.82907
R20640 gnd.n2699 gnd.t344 2.82907
R20641 gnd.n95 gnd.t355 2.82907
R20642 gnd.n95 gnd.t241 2.82907
R20643 gnd.n93 gnd.t384 2.82907
R20644 gnd.n93 gnd.t271 2.82907
R20645 gnd.n91 gnd.t319 2.82907
R20646 gnd.n91 gnd.t372 2.82907
R20647 gnd.n89 gnd.t394 2.82907
R20648 gnd.n89 gnd.t407 2.82907
R20649 gnd.n87 gnd.t409 2.82907
R20650 gnd.n87 gnd.t284 2.82907
R20651 gnd.n85 gnd.t404 2.82907
R20652 gnd.n85 gnd.t362 2.82907
R20653 gnd.n83 gnd.t337 2.82907
R20654 gnd.n83 gnd.t392 2.82907
R20655 gnd.n81 gnd.t358 2.82907
R20656 gnd.n81 gnd.t405 2.82907
R20657 gnd.n79 gnd.t375 2.82907
R20658 gnd.n79 gnd.t269 2.82907
R20659 gnd.n36 gnd.t383 2.82907
R20660 gnd.n36 gnd.t310 2.82907
R20661 gnd.n34 gnd.t279 2.82907
R20662 gnd.n34 gnd.t411 2.82907
R20663 gnd.n32 gnd.t393 2.82907
R20664 gnd.n32 gnd.t262 2.82907
R20665 gnd.n30 gnd.t217 2.82907
R20666 gnd.n30 gnd.t244 2.82907
R20667 gnd.n28 gnd.t373 2.82907
R20668 gnd.n28 gnd.t231 2.82907
R20669 gnd.n26 gnd.t325 2.82907
R20670 gnd.n26 gnd.t399 2.82907
R20671 gnd.n24 gnd.t387 2.82907
R20672 gnd.n24 gnd.t311 2.82907
R20673 gnd.n22 gnd.t281 2.82907
R20674 gnd.n22 gnd.t215 2.82907
R20675 gnd.n20 gnd.t398 2.82907
R20676 gnd.n20 gnd.t374 2.82907
R20677 gnd.n55 gnd.t397 2.82907
R20678 gnd.n55 gnd.t412 2.82907
R20679 gnd.n53 gnd.t410 2.82907
R20680 gnd.n53 gnd.t389 2.82907
R20681 gnd.n51 gnd.t386 2.82907
R20682 gnd.n51 gnd.t280 2.82907
R20683 gnd.n49 gnd.t300 2.82907
R20684 gnd.n49 gnd.t237 2.82907
R20685 gnd.n47 gnd.t248 2.82907
R20686 gnd.n47 gnd.t265 2.82907
R20687 gnd.n45 gnd.t267 2.82907
R20688 gnd.n45 gnd.t296 2.82907
R20689 gnd.n43 gnd.t299 2.82907
R20690 gnd.n43 gnd.t322 2.82907
R20691 gnd.n41 gnd.t320 2.82907
R20692 gnd.n41 gnd.t274 2.82907
R20693 gnd.n39 gnd.t275 2.82907
R20694 gnd.n39 gnd.t293 2.82907
R20695 gnd.n75 gnd.t406 2.82907
R20696 gnd.n75 gnd.t341 2.82907
R20697 gnd.n73 gnd.t283 2.82907
R20698 gnd.n73 gnd.t348 2.82907
R20699 gnd.n71 gnd.t371 2.82907
R20700 gnd.n71 gnd.t254 2.82907
R20701 gnd.n69 gnd.t305 2.82907
R20702 gnd.n69 gnd.t327 2.82907
R20703 gnd.n67 gnd.t333 2.82907
R20704 gnd.n67 gnd.t353 2.82907
R20705 gnd.n65 gnd.t323 2.82907
R20706 gnd.n65 gnd.t229 2.82907
R20707 gnd.n63 gnd.t381 2.82907
R20708 gnd.n63 gnd.t302 2.82907
R20709 gnd.n61 gnd.t219 2.82907
R20710 gnd.n61 gnd.t324 2.82907
R20711 gnd.n59 gnd.t256 2.82907
R20712 gnd.n59 gnd.t347 2.82907
R20713 gnd.n3285 gnd.t186 2.735
R20714 gnd.n2592 gnd.t191 2.735
R20715 gnd.n3767 gnd.n3766 2.71565
R20716 gnd.n3735 gnd.n3734 2.71565
R20717 gnd.n3703 gnd.n3702 2.71565
R20718 gnd.n3672 gnd.n3671 2.71565
R20719 gnd.n3640 gnd.n3639 2.71565
R20720 gnd.n3608 gnd.n3607 2.71565
R20721 gnd.n3576 gnd.n3575 2.71565
R20722 gnd.n3545 gnd.n3544 2.71565
R20723 gnd.n5186 gnd.n1614 2.54975
R20724 gnd.n5234 gnd.n1576 2.54975
R20725 gnd.n5235 gnd.t11 2.54975
R20726 gnd.n5300 gnd.n1530 2.54975
R20727 gnd.n5300 gnd.t5 2.54975
R20728 gnd.n5324 gnd.n5323 2.54975
R20729 gnd.n5465 gnd.n1444 2.54975
R20730 gnd.n5514 gnd.t153 2.54975
R20731 gnd.n5515 gnd.n5514 2.54975
R20732 gnd.t3 gnd.n1348 2.54975
R20733 gnd.n5627 gnd.n1341 2.54975
R20734 gnd.n5677 gnd.n1309 2.54975
R20735 gnd.n3229 gnd.t193 2.3704
R20736 gnd.n3459 gnd.t189 2.3704
R20737 gnd.n3302 gnd.n2724 2.27742
R20738 gnd.n3302 gnd.n2643 2.27742
R20739 gnd.n3302 gnd.n2642 2.27742
R20740 gnd.n3302 gnd.n2641 2.27742
R20741 gnd.n5397 gnd.t13 2.23109
R20742 gnd.t210 gnd.n1452 2.23109
R20743 gnd.n4270 gnd.t71 2.0058
R20744 gnd.n3763 gnd.n3753 1.93989
R20745 gnd.n3731 gnd.n3721 1.93989
R20746 gnd.n3699 gnd.n3689 1.93989
R20747 gnd.n3668 gnd.n3658 1.93989
R20748 gnd.n3636 gnd.n3626 1.93989
R20749 gnd.n3604 gnd.n3594 1.93989
R20750 gnd.n3572 gnd.n3562 1.93989
R20751 gnd.n3541 gnd.n3531 1.93989
R20752 gnd.n5180 gnd.t50 1.91244
R20753 gnd.n5228 gnd.t8 1.91244
R20754 gnd.n5634 gnd.t6 1.91244
R20755 gnd.n2808 gnd.t193 1.6412
R20756 gnd.n4558 gnd.t329 1.59378
R20757 gnd.n5235 gnd.t414 1.59378
R20758 gnd.t171 gnd.n1521 1.59378
R20759 gnd.n5531 gnd.t147 1.59378
R20760 gnd.n1348 gnd.t200 1.59378
R20761 gnd.n7074 gnd.t268 1.59378
R20762 gnd.n7681 gnd.t354 1.59378
R20763 gnd.n3156 gnd.t57 1.2766
R20764 gnd.n2779 gnd.t186 1.2766
R20765 gnd.n5160 gnd.t129 1.27512
R20766 gnd.n5192 gnd.n1602 1.27512
R20767 gnd.n1598 gnd.t9 1.27512
R20768 gnd.n1591 gnd.n1580 1.27512
R20769 gnd.n5276 gnd.t10 1.27512
R20770 gnd.n5311 gnd.n5310 1.27512
R20771 gnd.n5339 gnd.n5338 1.27512
R20772 gnd.n5486 gnd.n5485 1.27512
R20773 gnd.n5508 gnd.n1418 1.27512
R20774 gnd.n5575 gnd.t152 1.27512
R20775 gnd.n5633 gnd.n1332 1.27512
R20776 gnd.t160 gnd.n1333 1.27512
R20777 gnd.n5593 gnd.n1313 1.27512
R20778 gnd.t278 gnd.n167 1.27512
R20779 gnd.n3009 gnd.n3001 1.16414
R20780 gnd.n3825 gnd.n2479 1.16414
R20781 gnd.n3762 gnd.n3755 1.16414
R20782 gnd.n3730 gnd.n3723 1.16414
R20783 gnd.n3698 gnd.n3691 1.16414
R20784 gnd.n3667 gnd.n3660 1.16414
R20785 gnd.n3635 gnd.n3628 1.16414
R20786 gnd.n3603 gnd.n3596 1.16414
R20787 gnd.n3571 gnd.n3564 1.16414
R20788 gnd.n3540 gnd.n3533 1.16414
R20789 gnd.n6162 gnd.n6161 0.970197
R20790 gnd.n1952 gnd.n1750 0.970197
R20791 gnd.n3746 gnd.n3714 0.962709
R20792 gnd.n3778 gnd.n3746 0.962709
R20793 gnd.n3619 gnd.n3587 0.962709
R20794 gnd.n3651 gnd.n3619 0.962709
R20795 gnd.t234 gnd.n800 0.956468
R20796 gnd.n5151 gnd.n5150 0.956468
R20797 gnd.n1253 gnd.n1220 0.956468
R20798 gnd.n7037 gnd.t251 0.956468
R20799 gnd.n7157 gnd.t298 0.956468
R20800 gnd.n7705 gnd.t253 0.956468
R20801 gnd.t206 gnd.n3167 0.912001
R20802 gnd.n3346 gnd.t184 0.912001
R20803 gnd.n2576 gnd.t212 0.912001
R20804 gnd.n4322 gnd.t245 0.912001
R20805 gnd gnd.n0 0.70738
R20806 gnd.n2 gnd.n1 0.672012
R20807 gnd.n3 gnd.n2 0.672012
R20808 gnd.n4 gnd.n3 0.672012
R20809 gnd.n5 gnd.n4 0.672012
R20810 gnd.n6 gnd.n5 0.672012
R20811 gnd.n7 gnd.n6 0.672012
R20812 gnd.n8 gnd.n7 0.672012
R20813 gnd.n9 gnd.n8 0.672012
R20814 gnd.n11 gnd.n10 0.672012
R20815 gnd.n12 gnd.n11 0.672012
R20816 gnd.n13 gnd.n12 0.672012
R20817 gnd.n14 gnd.n13 0.672012
R20818 gnd.n15 gnd.n14 0.672012
R20819 gnd.n16 gnd.n15 0.672012
R20820 gnd.n17 gnd.n16 0.672012
R20821 gnd.n18 gnd.n17 0.672012
R20822 gnd.n6453 gnd.n752 0.637812
R20823 gnd.t82 gnd.n5192 0.637812
R20824 gnd.n5284 gnd.t26 0.637812
R20825 gnd.n1413 gnd.t169 0.637812
R20826 gnd.n7742 gnd.n7741 0.637193
R20827 gnd.n2721 gnd.n2720 0.573776
R20828 gnd.n2720 gnd.n2718 0.573776
R20829 gnd.n2718 gnd.n2716 0.573776
R20830 gnd.n2716 gnd.n2714 0.573776
R20831 gnd.n2714 gnd.n2712 0.573776
R20832 gnd.n2712 gnd.n2710 0.573776
R20833 gnd.n2710 gnd.n2708 0.573776
R20834 gnd.n2708 gnd.n2706 0.573776
R20835 gnd.n2706 gnd.n2704 0.573776
R20836 gnd.n2662 gnd.n2661 0.573776
R20837 gnd.n2661 gnd.n2659 0.573776
R20838 gnd.n2659 gnd.n2657 0.573776
R20839 gnd.n2657 gnd.n2655 0.573776
R20840 gnd.n2655 gnd.n2653 0.573776
R20841 gnd.n2653 gnd.n2651 0.573776
R20842 gnd.n2651 gnd.n2649 0.573776
R20843 gnd.n2649 gnd.n2647 0.573776
R20844 gnd.n2647 gnd.n2645 0.573776
R20845 gnd.n2681 gnd.n2680 0.573776
R20846 gnd.n2680 gnd.n2678 0.573776
R20847 gnd.n2678 gnd.n2676 0.573776
R20848 gnd.n2676 gnd.n2674 0.573776
R20849 gnd.n2674 gnd.n2672 0.573776
R20850 gnd.n2672 gnd.n2670 0.573776
R20851 gnd.n2670 gnd.n2668 0.573776
R20852 gnd.n2668 gnd.n2666 0.573776
R20853 gnd.n2666 gnd.n2664 0.573776
R20854 gnd.n2701 gnd.n2700 0.573776
R20855 gnd.n2700 gnd.n2698 0.573776
R20856 gnd.n2698 gnd.n2696 0.573776
R20857 gnd.n2696 gnd.n2694 0.573776
R20858 gnd.n2694 gnd.n2692 0.573776
R20859 gnd.n2692 gnd.n2690 0.573776
R20860 gnd.n2690 gnd.n2688 0.573776
R20861 gnd.n2688 gnd.n2686 0.573776
R20862 gnd.n2686 gnd.n2684 0.573776
R20863 gnd.n82 gnd.n80 0.573776
R20864 gnd.n84 gnd.n82 0.573776
R20865 gnd.n86 gnd.n84 0.573776
R20866 gnd.n88 gnd.n86 0.573776
R20867 gnd.n90 gnd.n88 0.573776
R20868 gnd.n92 gnd.n90 0.573776
R20869 gnd.n94 gnd.n92 0.573776
R20870 gnd.n96 gnd.n94 0.573776
R20871 gnd.n97 gnd.n96 0.573776
R20872 gnd.n23 gnd.n21 0.573776
R20873 gnd.n25 gnd.n23 0.573776
R20874 gnd.n27 gnd.n25 0.573776
R20875 gnd.n29 gnd.n27 0.573776
R20876 gnd.n31 gnd.n29 0.573776
R20877 gnd.n33 gnd.n31 0.573776
R20878 gnd.n35 gnd.n33 0.573776
R20879 gnd.n37 gnd.n35 0.573776
R20880 gnd.n38 gnd.n37 0.573776
R20881 gnd.n42 gnd.n40 0.573776
R20882 gnd.n44 gnd.n42 0.573776
R20883 gnd.n46 gnd.n44 0.573776
R20884 gnd.n48 gnd.n46 0.573776
R20885 gnd.n50 gnd.n48 0.573776
R20886 gnd.n52 gnd.n50 0.573776
R20887 gnd.n54 gnd.n52 0.573776
R20888 gnd.n56 gnd.n54 0.573776
R20889 gnd.n57 gnd.n56 0.573776
R20890 gnd.n62 gnd.n60 0.573776
R20891 gnd.n64 gnd.n62 0.573776
R20892 gnd.n66 gnd.n64 0.573776
R20893 gnd.n68 gnd.n66 0.573776
R20894 gnd.n70 gnd.n68 0.573776
R20895 gnd.n72 gnd.n70 0.573776
R20896 gnd.n74 gnd.n72 0.573776
R20897 gnd.n76 gnd.n74 0.573776
R20898 gnd.n77 gnd.n76 0.573776
R20899 gnd.n3255 gnd.t175 0.547401
R20900 gnd.n3420 gnd.t182 0.547401
R20901 gnd.n4362 gnd.t263 0.547401
R20902 gnd.n4524 gnd.t242 0.547401
R20903 gnd.n3482 gnd.n2483 0.486781
R20904 gnd.n3058 gnd.n3057 0.48678
R20905 gnd.n3799 gnd.n2437 0.480683
R20906 gnd.n3142 gnd.n3141 0.480683
R20907 gnd.n7396 gnd.n7395 0.477634
R20908 gnd.n4215 gnd.n4210 0.477634
R20909 gnd.n6231 gnd.n6230 0.451719
R20910 gnd.n6382 gnd.n867 0.451719
R20911 gnd.n5010 gnd.n5009 0.451719
R20912 gnd.n5912 gnd.n5911 0.451719
R20913 gnd.n5991 gnd.n1073 0.442573
R20914 gnd.n7492 gnd.n248 0.442573
R20915 gnd.n1780 gnd.n1779 0.442573
R20916 gnd.n4265 gnd.n2410 0.442573
R20917 gnd.n6457 gnd.n750 0.438
R20918 gnd.n6810 gnd.n6809 0.438
R20919 gnd.n7022 gnd.n7021 0.438
R20920 gnd.n4866 gnd.n4865 0.438
R20921 gnd.n2156 gnd.n2143 0.388379
R20922 gnd.n3759 gnd.n3758 0.388379
R20923 gnd.n3727 gnd.n3726 0.388379
R20924 gnd.n3695 gnd.n3694 0.388379
R20925 gnd.n3664 gnd.n3663 0.388379
R20926 gnd.n3632 gnd.n3631 0.388379
R20927 gnd.n3600 gnd.n3599 0.388379
R20928 gnd.n3568 gnd.n3567 0.388379
R20929 gnd.n3537 gnd.n3536 0.388379
R20930 gnd.n6224 gnd.n1017 0.388379
R20931 gnd.n7742 gnd.n19 0.374463
R20932 gnd gnd.n7742 0.367492
R20933 gnd.n7204 gnd.t228 0.319156
R20934 gnd.n7729 gnd.t216 0.319156
R20935 gnd.n2976 gnd.n2954 0.311721
R20936 gnd.n7641 gnd.n7428 0.293183
R20937 gnd.n4252 gnd.n4251 0.293183
R20938 gnd.n3870 gnd.n3869 0.268793
R20939 gnd.n6100 gnd.n6099 0.258122
R20940 gnd.n7641 gnd.n7640 0.258122
R20941 gnd.n6405 gnd.n6404 0.258122
R20942 gnd.n4252 gnd.n4122 0.258122
R20943 gnd.n4938 gnd.n4937 0.247451
R20944 gnd.n5968 gnd.n993 0.247451
R20945 gnd.n3869 gnd.n3868 0.241354
R20946 gnd.n1103 gnd.n1100 0.229039
R20947 gnd.n1104 gnd.n1103 0.229039
R20948 gnd.n1951 gnd.n1846 0.229039
R20949 gnd.n1951 gnd.n1950 0.229039
R20950 gnd.n2723 gnd.n0 0.210825
R20951 gnd.n3130 gnd.n2929 0.206293
R20952 gnd.n2538 gnd.t194 0.1828
R20953 gnd.n4406 gnd.t272 0.1828
R20954 gnd.n4465 gnd.t314 0.1828
R20955 gnd.n3776 gnd.n3748 0.155672
R20956 gnd.n3769 gnd.n3748 0.155672
R20957 gnd.n3769 gnd.n3768 0.155672
R20958 gnd.n3768 gnd.n3752 0.155672
R20959 gnd.n3761 gnd.n3752 0.155672
R20960 gnd.n3761 gnd.n3760 0.155672
R20961 gnd.n3744 gnd.n3716 0.155672
R20962 gnd.n3737 gnd.n3716 0.155672
R20963 gnd.n3737 gnd.n3736 0.155672
R20964 gnd.n3736 gnd.n3720 0.155672
R20965 gnd.n3729 gnd.n3720 0.155672
R20966 gnd.n3729 gnd.n3728 0.155672
R20967 gnd.n3712 gnd.n3684 0.155672
R20968 gnd.n3705 gnd.n3684 0.155672
R20969 gnd.n3705 gnd.n3704 0.155672
R20970 gnd.n3704 gnd.n3688 0.155672
R20971 gnd.n3697 gnd.n3688 0.155672
R20972 gnd.n3697 gnd.n3696 0.155672
R20973 gnd.n3681 gnd.n3653 0.155672
R20974 gnd.n3674 gnd.n3653 0.155672
R20975 gnd.n3674 gnd.n3673 0.155672
R20976 gnd.n3673 gnd.n3657 0.155672
R20977 gnd.n3666 gnd.n3657 0.155672
R20978 gnd.n3666 gnd.n3665 0.155672
R20979 gnd.n3649 gnd.n3621 0.155672
R20980 gnd.n3642 gnd.n3621 0.155672
R20981 gnd.n3642 gnd.n3641 0.155672
R20982 gnd.n3641 gnd.n3625 0.155672
R20983 gnd.n3634 gnd.n3625 0.155672
R20984 gnd.n3634 gnd.n3633 0.155672
R20985 gnd.n3617 gnd.n3589 0.155672
R20986 gnd.n3610 gnd.n3589 0.155672
R20987 gnd.n3610 gnd.n3609 0.155672
R20988 gnd.n3609 gnd.n3593 0.155672
R20989 gnd.n3602 gnd.n3593 0.155672
R20990 gnd.n3602 gnd.n3601 0.155672
R20991 gnd.n3585 gnd.n3557 0.155672
R20992 gnd.n3578 gnd.n3557 0.155672
R20993 gnd.n3578 gnd.n3577 0.155672
R20994 gnd.n3577 gnd.n3561 0.155672
R20995 gnd.n3570 gnd.n3561 0.155672
R20996 gnd.n3570 gnd.n3569 0.155672
R20997 gnd.n3554 gnd.n3526 0.155672
R20998 gnd.n3547 gnd.n3526 0.155672
R20999 gnd.n3547 gnd.n3546 0.155672
R21000 gnd.n3546 gnd.n3530 0.155672
R21001 gnd.n3539 gnd.n3530 0.155672
R21002 gnd.n3539 gnd.n3538 0.155672
R21003 gnd.n1074 gnd.n1073 0.152939
R21004 gnd.n1075 gnd.n1074 0.152939
R21005 gnd.n1076 gnd.n1075 0.152939
R21006 gnd.n1077 gnd.n1076 0.152939
R21007 gnd.n1078 gnd.n1077 0.152939
R21008 gnd.n1079 gnd.n1078 0.152939
R21009 gnd.n1080 gnd.n1079 0.152939
R21010 gnd.n1081 gnd.n1080 0.152939
R21011 gnd.n1082 gnd.n1081 0.152939
R21012 gnd.n1083 gnd.n1082 0.152939
R21013 gnd.n1084 gnd.n1083 0.152939
R21014 gnd.n1085 gnd.n1084 0.152939
R21015 gnd.n1086 gnd.n1085 0.152939
R21016 gnd.n1087 gnd.n1086 0.152939
R21017 gnd.n1088 gnd.n1087 0.152939
R21018 gnd.n1089 gnd.n1088 0.152939
R21019 gnd.n1090 gnd.n1089 0.152939
R21020 gnd.n1093 gnd.n1090 0.152939
R21021 gnd.n1094 gnd.n1093 0.152939
R21022 gnd.n1095 gnd.n1094 0.152939
R21023 gnd.n1096 gnd.n1095 0.152939
R21024 gnd.n1097 gnd.n1096 0.152939
R21025 gnd.n1098 gnd.n1097 0.152939
R21026 gnd.n1099 gnd.n1098 0.152939
R21027 gnd.n1100 gnd.n1099 0.152939
R21028 gnd.n1105 gnd.n1104 0.152939
R21029 gnd.n1106 gnd.n1105 0.152939
R21030 gnd.n1107 gnd.n1106 0.152939
R21031 gnd.n1108 gnd.n1107 0.152939
R21032 gnd.n1109 gnd.n1108 0.152939
R21033 gnd.n1110 gnd.n1109 0.152939
R21034 gnd.n1111 gnd.n1110 0.152939
R21035 gnd.n1112 gnd.n1111 0.152939
R21036 gnd.n1113 gnd.n1112 0.152939
R21037 gnd.n1116 gnd.n1113 0.152939
R21038 gnd.n1117 gnd.n1116 0.152939
R21039 gnd.n1118 gnd.n1117 0.152939
R21040 gnd.n1119 gnd.n1118 0.152939
R21041 gnd.n1120 gnd.n1119 0.152939
R21042 gnd.n1121 gnd.n1120 0.152939
R21043 gnd.n1122 gnd.n1121 0.152939
R21044 gnd.n1123 gnd.n1122 0.152939
R21045 gnd.n1124 gnd.n1123 0.152939
R21046 gnd.n1125 gnd.n1124 0.152939
R21047 gnd.n1126 gnd.n1125 0.152939
R21048 gnd.n1127 gnd.n1126 0.152939
R21049 gnd.n1128 gnd.n1127 0.152939
R21050 gnd.n1129 gnd.n1128 0.152939
R21051 gnd.n1130 gnd.n1129 0.152939
R21052 gnd.n1131 gnd.n1130 0.152939
R21053 gnd.n1132 gnd.n1131 0.152939
R21054 gnd.n1133 gnd.n1132 0.152939
R21055 gnd.n1134 gnd.n1133 0.152939
R21056 gnd.n6101 gnd.n1134 0.152939
R21057 gnd.n6101 gnd.n6100 0.152939
R21058 gnd.n5995 gnd.n5991 0.152939
R21059 gnd.n5996 gnd.n5995 0.152939
R21060 gnd.n5997 gnd.n5996 0.152939
R21061 gnd.n5998 gnd.n5997 0.152939
R21062 gnd.n5998 gnd.n388 0.152939
R21063 gnd.n7054 gnd.n388 0.152939
R21064 gnd.n7055 gnd.n7054 0.152939
R21065 gnd.n7056 gnd.n7055 0.152939
R21066 gnd.n7057 gnd.n7056 0.152939
R21067 gnd.n7057 gnd.n359 0.152939
R21068 gnd.n7090 gnd.n359 0.152939
R21069 gnd.n7091 gnd.n7090 0.152939
R21070 gnd.n7092 gnd.n7091 0.152939
R21071 gnd.n7093 gnd.n7092 0.152939
R21072 gnd.n7093 gnd.n332 0.152939
R21073 gnd.n7140 gnd.n332 0.152939
R21074 gnd.n7141 gnd.n7140 0.152939
R21075 gnd.n7142 gnd.n7141 0.152939
R21076 gnd.n7142 gnd.n315 0.152939
R21077 gnd.n7160 gnd.n315 0.152939
R21078 gnd.n7161 gnd.n7160 0.152939
R21079 gnd.n7162 gnd.n7161 0.152939
R21080 gnd.n7162 gnd.n295 0.152939
R21081 gnd.n7184 gnd.n295 0.152939
R21082 gnd.n7185 gnd.n7184 0.152939
R21083 gnd.n7186 gnd.n7185 0.152939
R21084 gnd.n7187 gnd.n7186 0.152939
R21085 gnd.n131 gnd.n130 0.152939
R21086 gnd.n132 gnd.n131 0.152939
R21087 gnd.n133 gnd.n132 0.152939
R21088 gnd.n150 gnd.n133 0.152939
R21089 gnd.n151 gnd.n150 0.152939
R21090 gnd.n152 gnd.n151 0.152939
R21091 gnd.n153 gnd.n152 0.152939
R21092 gnd.n169 gnd.n153 0.152939
R21093 gnd.n170 gnd.n169 0.152939
R21094 gnd.n171 gnd.n170 0.152939
R21095 gnd.n172 gnd.n171 0.152939
R21096 gnd.n189 gnd.n172 0.152939
R21097 gnd.n190 gnd.n189 0.152939
R21098 gnd.n191 gnd.n190 0.152939
R21099 gnd.n192 gnd.n191 0.152939
R21100 gnd.n207 gnd.n192 0.152939
R21101 gnd.n208 gnd.n207 0.152939
R21102 gnd.n209 gnd.n208 0.152939
R21103 gnd.n210 gnd.n209 0.152939
R21104 gnd.n227 gnd.n210 0.152939
R21105 gnd.n228 gnd.n227 0.152939
R21106 gnd.n229 gnd.n228 0.152939
R21107 gnd.n230 gnd.n229 0.152939
R21108 gnd.n245 gnd.n230 0.152939
R21109 gnd.n246 gnd.n245 0.152939
R21110 gnd.n247 gnd.n246 0.152939
R21111 gnd.n248 gnd.n247 0.152939
R21112 gnd.n7739 gnd.n101 0.152939
R21113 gnd.n7344 gnd.n101 0.152939
R21114 gnd.n7346 gnd.n7344 0.152939
R21115 gnd.n7347 gnd.n7346 0.152939
R21116 gnd.n7348 gnd.n7347 0.152939
R21117 gnd.n7348 gnd.n7341 0.152939
R21118 gnd.n7353 gnd.n7341 0.152939
R21119 gnd.n7354 gnd.n7353 0.152939
R21120 gnd.n7355 gnd.n7354 0.152939
R21121 gnd.n7355 gnd.n7338 0.152939
R21122 gnd.n7360 gnd.n7338 0.152939
R21123 gnd.n7361 gnd.n7360 0.152939
R21124 gnd.n7362 gnd.n7361 0.152939
R21125 gnd.n7362 gnd.n7335 0.152939
R21126 gnd.n7367 gnd.n7335 0.152939
R21127 gnd.n7368 gnd.n7367 0.152939
R21128 gnd.n7369 gnd.n7368 0.152939
R21129 gnd.n7369 gnd.n7332 0.152939
R21130 gnd.n7374 gnd.n7332 0.152939
R21131 gnd.n7375 gnd.n7374 0.152939
R21132 gnd.n7376 gnd.n7375 0.152939
R21133 gnd.n7376 gnd.n7329 0.152939
R21134 gnd.n7381 gnd.n7329 0.152939
R21135 gnd.n7382 gnd.n7381 0.152939
R21136 gnd.n7383 gnd.n7382 0.152939
R21137 gnd.n7383 gnd.n7326 0.152939
R21138 gnd.n7388 gnd.n7326 0.152939
R21139 gnd.n7389 gnd.n7388 0.152939
R21140 gnd.n7390 gnd.n7389 0.152939
R21141 gnd.n7390 gnd.n7323 0.152939
R21142 gnd.n7395 gnd.n7323 0.152939
R21143 gnd.n7428 gnd.n7289 0.152939
R21144 gnd.n7291 gnd.n7289 0.152939
R21145 gnd.n7295 gnd.n7291 0.152939
R21146 gnd.n7296 gnd.n7295 0.152939
R21147 gnd.n7297 gnd.n7296 0.152939
R21148 gnd.n7298 gnd.n7297 0.152939
R21149 gnd.n7302 gnd.n7298 0.152939
R21150 gnd.n7303 gnd.n7302 0.152939
R21151 gnd.n7304 gnd.n7303 0.152939
R21152 gnd.n7305 gnd.n7304 0.152939
R21153 gnd.n7309 gnd.n7305 0.152939
R21154 gnd.n7310 gnd.n7309 0.152939
R21155 gnd.n7311 gnd.n7310 0.152939
R21156 gnd.n7312 gnd.n7311 0.152939
R21157 gnd.n7316 gnd.n7312 0.152939
R21158 gnd.n7317 gnd.n7316 0.152939
R21159 gnd.n7397 gnd.n7317 0.152939
R21160 gnd.n7397 gnd.n7396 0.152939
R21161 gnd.n7492 gnd.n7491 0.152939
R21162 gnd.n7500 gnd.n7491 0.152939
R21163 gnd.n7501 gnd.n7500 0.152939
R21164 gnd.n7502 gnd.n7501 0.152939
R21165 gnd.n7502 gnd.n7487 0.152939
R21166 gnd.n7510 gnd.n7487 0.152939
R21167 gnd.n7511 gnd.n7510 0.152939
R21168 gnd.n7512 gnd.n7511 0.152939
R21169 gnd.n7512 gnd.n7483 0.152939
R21170 gnd.n7520 gnd.n7483 0.152939
R21171 gnd.n7521 gnd.n7520 0.152939
R21172 gnd.n7522 gnd.n7521 0.152939
R21173 gnd.n7522 gnd.n7479 0.152939
R21174 gnd.n7531 gnd.n7479 0.152939
R21175 gnd.n7532 gnd.n7531 0.152939
R21176 gnd.n7533 gnd.n7532 0.152939
R21177 gnd.n7533 gnd.n7473 0.152939
R21178 gnd.n7541 gnd.n7473 0.152939
R21179 gnd.n7542 gnd.n7541 0.152939
R21180 gnd.n7543 gnd.n7542 0.152939
R21181 gnd.n7543 gnd.n7469 0.152939
R21182 gnd.n7551 gnd.n7469 0.152939
R21183 gnd.n7552 gnd.n7551 0.152939
R21184 gnd.n7553 gnd.n7552 0.152939
R21185 gnd.n7553 gnd.n7465 0.152939
R21186 gnd.n7561 gnd.n7465 0.152939
R21187 gnd.n7562 gnd.n7561 0.152939
R21188 gnd.n7563 gnd.n7562 0.152939
R21189 gnd.n7563 gnd.n7461 0.152939
R21190 gnd.n7571 gnd.n7461 0.152939
R21191 gnd.n7572 gnd.n7571 0.152939
R21192 gnd.n7573 gnd.n7572 0.152939
R21193 gnd.n7573 gnd.n7457 0.152939
R21194 gnd.n7581 gnd.n7457 0.152939
R21195 gnd.n7582 gnd.n7581 0.152939
R21196 gnd.n7583 gnd.n7582 0.152939
R21197 gnd.n7583 gnd.n7451 0.152939
R21198 gnd.n7591 gnd.n7451 0.152939
R21199 gnd.n7592 gnd.n7591 0.152939
R21200 gnd.n7593 gnd.n7592 0.152939
R21201 gnd.n7593 gnd.n7447 0.152939
R21202 gnd.n7601 gnd.n7447 0.152939
R21203 gnd.n7602 gnd.n7601 0.152939
R21204 gnd.n7603 gnd.n7602 0.152939
R21205 gnd.n7603 gnd.n7443 0.152939
R21206 gnd.n7611 gnd.n7443 0.152939
R21207 gnd.n7612 gnd.n7611 0.152939
R21208 gnd.n7613 gnd.n7612 0.152939
R21209 gnd.n7613 gnd.n7439 0.152939
R21210 gnd.n7621 gnd.n7439 0.152939
R21211 gnd.n7622 gnd.n7621 0.152939
R21212 gnd.n7623 gnd.n7622 0.152939
R21213 gnd.n7623 gnd.n7435 0.152939
R21214 gnd.n7631 gnd.n7435 0.152939
R21215 gnd.n7632 gnd.n7631 0.152939
R21216 gnd.n7633 gnd.n7632 0.152939
R21217 gnd.n7633 gnd.n7429 0.152939
R21218 gnd.n7640 gnd.n7429 0.152939
R21219 gnd.n6458 gnd.n6457 0.152939
R21220 gnd.n6459 gnd.n6458 0.152939
R21221 gnd.n6459 gnd.n744 0.152939
R21222 gnd.n6467 gnd.n744 0.152939
R21223 gnd.n6468 gnd.n6467 0.152939
R21224 gnd.n6469 gnd.n6468 0.152939
R21225 gnd.n6469 gnd.n738 0.152939
R21226 gnd.n6477 gnd.n738 0.152939
R21227 gnd.n6478 gnd.n6477 0.152939
R21228 gnd.n6479 gnd.n6478 0.152939
R21229 gnd.n6479 gnd.n732 0.152939
R21230 gnd.n6487 gnd.n732 0.152939
R21231 gnd.n6488 gnd.n6487 0.152939
R21232 gnd.n6489 gnd.n6488 0.152939
R21233 gnd.n6489 gnd.n726 0.152939
R21234 gnd.n6497 gnd.n726 0.152939
R21235 gnd.n6498 gnd.n6497 0.152939
R21236 gnd.n6499 gnd.n6498 0.152939
R21237 gnd.n6499 gnd.n720 0.152939
R21238 gnd.n6507 gnd.n720 0.152939
R21239 gnd.n6508 gnd.n6507 0.152939
R21240 gnd.n6509 gnd.n6508 0.152939
R21241 gnd.n6509 gnd.n714 0.152939
R21242 gnd.n6517 gnd.n714 0.152939
R21243 gnd.n6518 gnd.n6517 0.152939
R21244 gnd.n6519 gnd.n6518 0.152939
R21245 gnd.n6519 gnd.n708 0.152939
R21246 gnd.n6527 gnd.n708 0.152939
R21247 gnd.n6528 gnd.n6527 0.152939
R21248 gnd.n6529 gnd.n6528 0.152939
R21249 gnd.n6529 gnd.n702 0.152939
R21250 gnd.n6537 gnd.n702 0.152939
R21251 gnd.n6538 gnd.n6537 0.152939
R21252 gnd.n6539 gnd.n6538 0.152939
R21253 gnd.n6539 gnd.n696 0.152939
R21254 gnd.n6547 gnd.n696 0.152939
R21255 gnd.n6548 gnd.n6547 0.152939
R21256 gnd.n6549 gnd.n6548 0.152939
R21257 gnd.n6549 gnd.n690 0.152939
R21258 gnd.n6557 gnd.n690 0.152939
R21259 gnd.n6558 gnd.n6557 0.152939
R21260 gnd.n6559 gnd.n6558 0.152939
R21261 gnd.n6559 gnd.n684 0.152939
R21262 gnd.n6567 gnd.n684 0.152939
R21263 gnd.n6568 gnd.n6567 0.152939
R21264 gnd.n6569 gnd.n6568 0.152939
R21265 gnd.n6569 gnd.n678 0.152939
R21266 gnd.n6577 gnd.n678 0.152939
R21267 gnd.n6578 gnd.n6577 0.152939
R21268 gnd.n6579 gnd.n6578 0.152939
R21269 gnd.n6579 gnd.n672 0.152939
R21270 gnd.n6587 gnd.n672 0.152939
R21271 gnd.n6588 gnd.n6587 0.152939
R21272 gnd.n6589 gnd.n6588 0.152939
R21273 gnd.n6589 gnd.n666 0.152939
R21274 gnd.n6597 gnd.n666 0.152939
R21275 gnd.n6598 gnd.n6597 0.152939
R21276 gnd.n6599 gnd.n6598 0.152939
R21277 gnd.n6599 gnd.n660 0.152939
R21278 gnd.n6607 gnd.n660 0.152939
R21279 gnd.n6608 gnd.n6607 0.152939
R21280 gnd.n6609 gnd.n6608 0.152939
R21281 gnd.n6609 gnd.n654 0.152939
R21282 gnd.n6617 gnd.n654 0.152939
R21283 gnd.n6618 gnd.n6617 0.152939
R21284 gnd.n6619 gnd.n6618 0.152939
R21285 gnd.n6619 gnd.n648 0.152939
R21286 gnd.n6627 gnd.n648 0.152939
R21287 gnd.n6628 gnd.n6627 0.152939
R21288 gnd.n6629 gnd.n6628 0.152939
R21289 gnd.n6629 gnd.n642 0.152939
R21290 gnd.n6637 gnd.n642 0.152939
R21291 gnd.n6638 gnd.n6637 0.152939
R21292 gnd.n6639 gnd.n6638 0.152939
R21293 gnd.n6639 gnd.n636 0.152939
R21294 gnd.n6647 gnd.n636 0.152939
R21295 gnd.n6648 gnd.n6647 0.152939
R21296 gnd.n6649 gnd.n6648 0.152939
R21297 gnd.n6649 gnd.n630 0.152939
R21298 gnd.n6657 gnd.n630 0.152939
R21299 gnd.n6658 gnd.n6657 0.152939
R21300 gnd.n6659 gnd.n6658 0.152939
R21301 gnd.n6659 gnd.n624 0.152939
R21302 gnd.n6667 gnd.n624 0.152939
R21303 gnd.n6668 gnd.n6667 0.152939
R21304 gnd.n6669 gnd.n6668 0.152939
R21305 gnd.n6669 gnd.n618 0.152939
R21306 gnd.n6677 gnd.n618 0.152939
R21307 gnd.n6678 gnd.n6677 0.152939
R21308 gnd.n6679 gnd.n6678 0.152939
R21309 gnd.n6679 gnd.n612 0.152939
R21310 gnd.n6687 gnd.n612 0.152939
R21311 gnd.n6688 gnd.n6687 0.152939
R21312 gnd.n6689 gnd.n6688 0.152939
R21313 gnd.n6689 gnd.n606 0.152939
R21314 gnd.n6697 gnd.n606 0.152939
R21315 gnd.n6698 gnd.n6697 0.152939
R21316 gnd.n6699 gnd.n6698 0.152939
R21317 gnd.n6699 gnd.n600 0.152939
R21318 gnd.n6707 gnd.n600 0.152939
R21319 gnd.n6708 gnd.n6707 0.152939
R21320 gnd.n6709 gnd.n6708 0.152939
R21321 gnd.n6709 gnd.n594 0.152939
R21322 gnd.n6717 gnd.n594 0.152939
R21323 gnd.n6718 gnd.n6717 0.152939
R21324 gnd.n6719 gnd.n6718 0.152939
R21325 gnd.n6719 gnd.n588 0.152939
R21326 gnd.n6727 gnd.n588 0.152939
R21327 gnd.n6728 gnd.n6727 0.152939
R21328 gnd.n6729 gnd.n6728 0.152939
R21329 gnd.n6729 gnd.n582 0.152939
R21330 gnd.n6737 gnd.n582 0.152939
R21331 gnd.n6738 gnd.n6737 0.152939
R21332 gnd.n6739 gnd.n6738 0.152939
R21333 gnd.n6739 gnd.n576 0.152939
R21334 gnd.n6747 gnd.n576 0.152939
R21335 gnd.n6748 gnd.n6747 0.152939
R21336 gnd.n6749 gnd.n6748 0.152939
R21337 gnd.n6749 gnd.n570 0.152939
R21338 gnd.n6757 gnd.n570 0.152939
R21339 gnd.n6758 gnd.n6757 0.152939
R21340 gnd.n6759 gnd.n6758 0.152939
R21341 gnd.n6759 gnd.n564 0.152939
R21342 gnd.n6767 gnd.n564 0.152939
R21343 gnd.n6768 gnd.n6767 0.152939
R21344 gnd.n6769 gnd.n6768 0.152939
R21345 gnd.n6769 gnd.n558 0.152939
R21346 gnd.n6777 gnd.n558 0.152939
R21347 gnd.n6778 gnd.n6777 0.152939
R21348 gnd.n6779 gnd.n6778 0.152939
R21349 gnd.n6779 gnd.n552 0.152939
R21350 gnd.n6787 gnd.n552 0.152939
R21351 gnd.n6788 gnd.n6787 0.152939
R21352 gnd.n6789 gnd.n6788 0.152939
R21353 gnd.n6789 gnd.n546 0.152939
R21354 gnd.n6797 gnd.n546 0.152939
R21355 gnd.n6798 gnd.n6797 0.152939
R21356 gnd.n6800 gnd.n6798 0.152939
R21357 gnd.n6800 gnd.n6799 0.152939
R21358 gnd.n6799 gnd.n540 0.152939
R21359 gnd.n6809 gnd.n540 0.152939
R21360 gnd.n6810 gnd.n535 0.152939
R21361 gnd.n6818 gnd.n535 0.152939
R21362 gnd.n6819 gnd.n6818 0.152939
R21363 gnd.n6820 gnd.n6819 0.152939
R21364 gnd.n6820 gnd.n529 0.152939
R21365 gnd.n6828 gnd.n529 0.152939
R21366 gnd.n6829 gnd.n6828 0.152939
R21367 gnd.n6830 gnd.n6829 0.152939
R21368 gnd.n6830 gnd.n523 0.152939
R21369 gnd.n6838 gnd.n523 0.152939
R21370 gnd.n6839 gnd.n6838 0.152939
R21371 gnd.n6840 gnd.n6839 0.152939
R21372 gnd.n6840 gnd.n517 0.152939
R21373 gnd.n6848 gnd.n517 0.152939
R21374 gnd.n6849 gnd.n6848 0.152939
R21375 gnd.n6850 gnd.n6849 0.152939
R21376 gnd.n6850 gnd.n511 0.152939
R21377 gnd.n6858 gnd.n511 0.152939
R21378 gnd.n6859 gnd.n6858 0.152939
R21379 gnd.n6860 gnd.n6859 0.152939
R21380 gnd.n6860 gnd.n505 0.152939
R21381 gnd.n6868 gnd.n505 0.152939
R21382 gnd.n6869 gnd.n6868 0.152939
R21383 gnd.n6870 gnd.n6869 0.152939
R21384 gnd.n6870 gnd.n499 0.152939
R21385 gnd.n6878 gnd.n499 0.152939
R21386 gnd.n6879 gnd.n6878 0.152939
R21387 gnd.n6880 gnd.n6879 0.152939
R21388 gnd.n6880 gnd.n493 0.152939
R21389 gnd.n6888 gnd.n493 0.152939
R21390 gnd.n6889 gnd.n6888 0.152939
R21391 gnd.n6890 gnd.n6889 0.152939
R21392 gnd.n6890 gnd.n487 0.152939
R21393 gnd.n6898 gnd.n487 0.152939
R21394 gnd.n6899 gnd.n6898 0.152939
R21395 gnd.n6900 gnd.n6899 0.152939
R21396 gnd.n6900 gnd.n481 0.152939
R21397 gnd.n6908 gnd.n481 0.152939
R21398 gnd.n6909 gnd.n6908 0.152939
R21399 gnd.n6910 gnd.n6909 0.152939
R21400 gnd.n6910 gnd.n475 0.152939
R21401 gnd.n6918 gnd.n475 0.152939
R21402 gnd.n6919 gnd.n6918 0.152939
R21403 gnd.n6920 gnd.n6919 0.152939
R21404 gnd.n6920 gnd.n469 0.152939
R21405 gnd.n6928 gnd.n469 0.152939
R21406 gnd.n6929 gnd.n6928 0.152939
R21407 gnd.n6930 gnd.n6929 0.152939
R21408 gnd.n6930 gnd.n463 0.152939
R21409 gnd.n6938 gnd.n463 0.152939
R21410 gnd.n6939 gnd.n6938 0.152939
R21411 gnd.n6940 gnd.n6939 0.152939
R21412 gnd.n6940 gnd.n457 0.152939
R21413 gnd.n6948 gnd.n457 0.152939
R21414 gnd.n6949 gnd.n6948 0.152939
R21415 gnd.n6950 gnd.n6949 0.152939
R21416 gnd.n6950 gnd.n451 0.152939
R21417 gnd.n6958 gnd.n451 0.152939
R21418 gnd.n6959 gnd.n6958 0.152939
R21419 gnd.n6960 gnd.n6959 0.152939
R21420 gnd.n6960 gnd.n445 0.152939
R21421 gnd.n6968 gnd.n445 0.152939
R21422 gnd.n6969 gnd.n6968 0.152939
R21423 gnd.n6970 gnd.n6969 0.152939
R21424 gnd.n6970 gnd.n439 0.152939
R21425 gnd.n6978 gnd.n439 0.152939
R21426 gnd.n6979 gnd.n6978 0.152939
R21427 gnd.n6980 gnd.n6979 0.152939
R21428 gnd.n6980 gnd.n433 0.152939
R21429 gnd.n6988 gnd.n433 0.152939
R21430 gnd.n6989 gnd.n6988 0.152939
R21431 gnd.n6990 gnd.n6989 0.152939
R21432 gnd.n6990 gnd.n427 0.152939
R21433 gnd.n6998 gnd.n427 0.152939
R21434 gnd.n6999 gnd.n6998 0.152939
R21435 gnd.n7000 gnd.n6999 0.152939
R21436 gnd.n7000 gnd.n421 0.152939
R21437 gnd.n7008 gnd.n421 0.152939
R21438 gnd.n7009 gnd.n7008 0.152939
R21439 gnd.n7010 gnd.n7009 0.152939
R21440 gnd.n7010 gnd.n415 0.152939
R21441 gnd.n7019 gnd.n415 0.152939
R21442 gnd.n7020 gnd.n7019 0.152939
R21443 gnd.n7022 gnd.n7020 0.152939
R21444 gnd.n4866 gnd.n4569 0.152939
R21445 gnd.n4872 gnd.n4569 0.152939
R21446 gnd.n4873 gnd.n4872 0.152939
R21447 gnd.n4874 gnd.n4873 0.152939
R21448 gnd.n4875 gnd.n4874 0.152939
R21449 gnd.n4876 gnd.n4875 0.152939
R21450 gnd.n4879 gnd.n4876 0.152939
R21451 gnd.n4880 gnd.n4879 0.152939
R21452 gnd.n4881 gnd.n4880 0.152939
R21453 gnd.n4882 gnd.n4881 0.152939
R21454 gnd.n4884 gnd.n4882 0.152939
R21455 gnd.n4886 gnd.n4884 0.152939
R21456 gnd.n4886 gnd.n4885 0.152939
R21457 gnd.n4885 gnd.n847 0.152939
R21458 gnd.n848 gnd.n847 0.152939
R21459 gnd.n849 gnd.n848 0.152939
R21460 gnd.n855 gnd.n849 0.152939
R21461 gnd.n856 gnd.n855 0.152939
R21462 gnd.n857 gnd.n856 0.152939
R21463 gnd.n858 gnd.n857 0.152939
R21464 gnd.n5018 gnd.n858 0.152939
R21465 gnd.n5019 gnd.n5018 0.152939
R21466 gnd.n5020 gnd.n5019 0.152939
R21467 gnd.n5020 gnd.n2058 0.152939
R21468 gnd.n5036 gnd.n2058 0.152939
R21469 gnd.n5037 gnd.n5036 0.152939
R21470 gnd.n5038 gnd.n5037 0.152939
R21471 gnd.n5038 gnd.n2047 0.152939
R21472 gnd.n5053 gnd.n2047 0.152939
R21473 gnd.n5054 gnd.n5053 0.152939
R21474 gnd.n5055 gnd.n5054 0.152939
R21475 gnd.n5055 gnd.n2035 0.152939
R21476 gnd.n5070 gnd.n2035 0.152939
R21477 gnd.n5071 gnd.n5070 0.152939
R21478 gnd.n5072 gnd.n5071 0.152939
R21479 gnd.n5073 gnd.n5072 0.152939
R21480 gnd.n5073 gnd.n1625 0.152939
R21481 gnd.n5163 gnd.n1625 0.152939
R21482 gnd.n5164 gnd.n5163 0.152939
R21483 gnd.n5165 gnd.n5164 0.152939
R21484 gnd.n5166 gnd.n5165 0.152939
R21485 gnd.n5167 gnd.n5166 0.152939
R21486 gnd.n5169 gnd.n5167 0.152939
R21487 gnd.n5170 gnd.n5169 0.152939
R21488 gnd.n5170 gnd.n1586 0.152939
R21489 gnd.n5222 gnd.n1586 0.152939
R21490 gnd.n5223 gnd.n5222 0.152939
R21491 gnd.n5224 gnd.n5223 0.152939
R21492 gnd.n5224 gnd.n1564 0.152939
R21493 gnd.n5252 gnd.n1564 0.152939
R21494 gnd.n5253 gnd.n5252 0.152939
R21495 gnd.n5254 gnd.n5253 0.152939
R21496 gnd.n5254 gnd.n1547 0.152939
R21497 gnd.n5279 gnd.n1547 0.152939
R21498 gnd.n5280 gnd.n5279 0.152939
R21499 gnd.n5281 gnd.n5280 0.152939
R21500 gnd.n5281 gnd.n1527 0.152939
R21501 gnd.n5303 gnd.n1527 0.152939
R21502 gnd.n5304 gnd.n5303 0.152939
R21503 gnd.n5305 gnd.n5304 0.152939
R21504 gnd.n5306 gnd.n5305 0.152939
R21505 gnd.n5306 gnd.n1500 0.152939
R21506 gnd.n5361 gnd.n1500 0.152939
R21507 gnd.n5362 gnd.n5361 0.152939
R21508 gnd.n5363 gnd.n5362 0.152939
R21509 gnd.n5364 gnd.n5363 0.152939
R21510 gnd.n5364 gnd.n1478 0.152939
R21511 gnd.n5401 gnd.n1478 0.152939
R21512 gnd.n5402 gnd.n5401 0.152939
R21513 gnd.n5403 gnd.n5402 0.152939
R21514 gnd.n5404 gnd.n5403 0.152939
R21515 gnd.n5404 gnd.n1449 0.152939
R21516 gnd.n5458 gnd.n1449 0.152939
R21517 gnd.n5459 gnd.n5458 0.152939
R21518 gnd.n5460 gnd.n5459 0.152939
R21519 gnd.n5461 gnd.n5460 0.152939
R21520 gnd.n5461 gnd.n1428 0.152939
R21521 gnd.n5496 gnd.n1428 0.152939
R21522 gnd.n5497 gnd.n5496 0.152939
R21523 gnd.n5498 gnd.n5497 0.152939
R21524 gnd.n5498 gnd.n1399 0.152939
R21525 gnd.n5534 gnd.n1399 0.152939
R21526 gnd.n5535 gnd.n5534 0.152939
R21527 gnd.n5536 gnd.n5535 0.152939
R21528 gnd.n5537 gnd.n5536 0.152939
R21529 gnd.n5537 gnd.n1373 0.152939
R21530 gnd.n5578 gnd.n1373 0.152939
R21531 gnd.n5579 gnd.n5578 0.152939
R21532 gnd.n5581 gnd.n5579 0.152939
R21533 gnd.n5581 gnd.n5580 0.152939
R21534 gnd.n5580 gnd.n1352 0.152939
R21535 gnd.n1353 gnd.n1352 0.152939
R21536 gnd.n1354 gnd.n1353 0.152939
R21537 gnd.n1356 gnd.n1354 0.152939
R21538 gnd.n1357 gnd.n1356 0.152939
R21539 gnd.n1357 gnd.n1318 0.152939
R21540 gnd.n5665 gnd.n1318 0.152939
R21541 gnd.n5666 gnd.n5665 0.152939
R21542 gnd.n5667 gnd.n5666 0.152939
R21543 gnd.n5667 gnd.n1223 0.152939
R21544 gnd.n5813 gnd.n1223 0.152939
R21545 gnd.n5814 gnd.n5813 0.152939
R21546 gnd.n5815 gnd.n5814 0.152939
R21547 gnd.n5815 gnd.n1211 0.152939
R21548 gnd.n5830 gnd.n1211 0.152939
R21549 gnd.n5831 gnd.n5830 0.152939
R21550 gnd.n5832 gnd.n5831 0.152939
R21551 gnd.n5832 gnd.n1199 0.152939
R21552 gnd.n5847 gnd.n1199 0.152939
R21553 gnd.n5848 gnd.n5847 0.152939
R21554 gnd.n5849 gnd.n5848 0.152939
R21555 gnd.n5849 gnd.n1187 0.152939
R21556 gnd.n5865 gnd.n1187 0.152939
R21557 gnd.n5866 gnd.n5865 0.152939
R21558 gnd.n5867 gnd.n5866 0.152939
R21559 gnd.n5867 gnd.n1176 0.152939
R21560 gnd.n5882 gnd.n1176 0.152939
R21561 gnd.n5883 gnd.n5882 0.152939
R21562 gnd.n5884 gnd.n5883 0.152939
R21563 gnd.n5885 gnd.n5884 0.152939
R21564 gnd.n5885 gnd.n1163 0.152939
R21565 gnd.n5919 gnd.n1163 0.152939
R21566 gnd.n5920 gnd.n5919 0.152939
R21567 gnd.n5921 gnd.n5920 0.152939
R21568 gnd.n5921 gnd.n1159 0.152939
R21569 gnd.n5928 gnd.n1159 0.152939
R21570 gnd.n5929 gnd.n5928 0.152939
R21571 gnd.n5930 gnd.n5929 0.152939
R21572 gnd.n5931 gnd.n5930 0.152939
R21573 gnd.n5932 gnd.n5931 0.152939
R21574 gnd.n5944 gnd.n5932 0.152939
R21575 gnd.n5946 gnd.n5944 0.152939
R21576 gnd.n5946 gnd.n5945 0.152939
R21577 gnd.n5945 gnd.n403 0.152939
R21578 gnd.n404 gnd.n403 0.152939
R21579 gnd.n405 gnd.n404 0.152939
R21580 gnd.n408 gnd.n405 0.152939
R21581 gnd.n409 gnd.n408 0.152939
R21582 gnd.n410 gnd.n409 0.152939
R21583 gnd.n411 gnd.n410 0.152939
R21584 gnd.n7021 gnd.n411 0.152939
R21585 gnd.n4655 gnd.n750 0.152939
R21586 gnd.n4655 gnd.n4652 0.152939
R21587 gnd.n4663 gnd.n4652 0.152939
R21588 gnd.n4664 gnd.n4663 0.152939
R21589 gnd.n4665 gnd.n4664 0.152939
R21590 gnd.n4665 gnd.n4648 0.152939
R21591 gnd.n4673 gnd.n4648 0.152939
R21592 gnd.n4674 gnd.n4673 0.152939
R21593 gnd.n4675 gnd.n4674 0.152939
R21594 gnd.n4675 gnd.n4644 0.152939
R21595 gnd.n4683 gnd.n4644 0.152939
R21596 gnd.n4684 gnd.n4683 0.152939
R21597 gnd.n4685 gnd.n4684 0.152939
R21598 gnd.n4685 gnd.n4640 0.152939
R21599 gnd.n4693 gnd.n4640 0.152939
R21600 gnd.n4694 gnd.n4693 0.152939
R21601 gnd.n4695 gnd.n4694 0.152939
R21602 gnd.n4695 gnd.n4636 0.152939
R21603 gnd.n4703 gnd.n4636 0.152939
R21604 gnd.n4704 gnd.n4703 0.152939
R21605 gnd.n4705 gnd.n4704 0.152939
R21606 gnd.n4705 gnd.n4632 0.152939
R21607 gnd.n4713 gnd.n4632 0.152939
R21608 gnd.n4714 gnd.n4713 0.152939
R21609 gnd.n4715 gnd.n4714 0.152939
R21610 gnd.n4715 gnd.n4628 0.152939
R21611 gnd.n4723 gnd.n4628 0.152939
R21612 gnd.n4724 gnd.n4723 0.152939
R21613 gnd.n4725 gnd.n4724 0.152939
R21614 gnd.n4725 gnd.n4624 0.152939
R21615 gnd.n4733 gnd.n4624 0.152939
R21616 gnd.n4734 gnd.n4733 0.152939
R21617 gnd.n4735 gnd.n4734 0.152939
R21618 gnd.n4735 gnd.n4620 0.152939
R21619 gnd.n4743 gnd.n4620 0.152939
R21620 gnd.n4744 gnd.n4743 0.152939
R21621 gnd.n4745 gnd.n4744 0.152939
R21622 gnd.n4745 gnd.n4616 0.152939
R21623 gnd.n4753 gnd.n4616 0.152939
R21624 gnd.n4754 gnd.n4753 0.152939
R21625 gnd.n4755 gnd.n4754 0.152939
R21626 gnd.n4755 gnd.n4612 0.152939
R21627 gnd.n4763 gnd.n4612 0.152939
R21628 gnd.n4764 gnd.n4763 0.152939
R21629 gnd.n4765 gnd.n4764 0.152939
R21630 gnd.n4765 gnd.n4608 0.152939
R21631 gnd.n4773 gnd.n4608 0.152939
R21632 gnd.n4774 gnd.n4773 0.152939
R21633 gnd.n4775 gnd.n4774 0.152939
R21634 gnd.n4775 gnd.n4604 0.152939
R21635 gnd.n4783 gnd.n4604 0.152939
R21636 gnd.n4784 gnd.n4783 0.152939
R21637 gnd.n4785 gnd.n4784 0.152939
R21638 gnd.n4785 gnd.n4600 0.152939
R21639 gnd.n4793 gnd.n4600 0.152939
R21640 gnd.n4794 gnd.n4793 0.152939
R21641 gnd.n4795 gnd.n4794 0.152939
R21642 gnd.n4795 gnd.n4596 0.152939
R21643 gnd.n4803 gnd.n4596 0.152939
R21644 gnd.n4804 gnd.n4803 0.152939
R21645 gnd.n4805 gnd.n4804 0.152939
R21646 gnd.n4805 gnd.n4592 0.152939
R21647 gnd.n4813 gnd.n4592 0.152939
R21648 gnd.n4814 gnd.n4813 0.152939
R21649 gnd.n4815 gnd.n4814 0.152939
R21650 gnd.n4815 gnd.n4588 0.152939
R21651 gnd.n4823 gnd.n4588 0.152939
R21652 gnd.n4824 gnd.n4823 0.152939
R21653 gnd.n4825 gnd.n4824 0.152939
R21654 gnd.n4825 gnd.n4584 0.152939
R21655 gnd.n4833 gnd.n4584 0.152939
R21656 gnd.n4834 gnd.n4833 0.152939
R21657 gnd.n4835 gnd.n4834 0.152939
R21658 gnd.n4835 gnd.n4580 0.152939
R21659 gnd.n4843 gnd.n4580 0.152939
R21660 gnd.n4844 gnd.n4843 0.152939
R21661 gnd.n4845 gnd.n4844 0.152939
R21662 gnd.n4845 gnd.n4576 0.152939
R21663 gnd.n4853 gnd.n4576 0.152939
R21664 gnd.n4854 gnd.n4853 0.152939
R21665 gnd.n4856 gnd.n4854 0.152939
R21666 gnd.n4856 gnd.n4855 0.152939
R21667 gnd.n4855 gnd.n4572 0.152939
R21668 gnd.n4865 gnd.n4572 0.152939
R21669 gnd.n3901 gnd.n2437 0.152939
R21670 gnd.n3901 gnd.n3900 0.152939
R21671 gnd.n3900 gnd.n3899 0.152939
R21672 gnd.n3899 gnd.n2439 0.152939
R21673 gnd.n2440 gnd.n2439 0.152939
R21674 gnd.n2441 gnd.n2440 0.152939
R21675 gnd.n2442 gnd.n2441 0.152939
R21676 gnd.n2443 gnd.n2442 0.152939
R21677 gnd.n2444 gnd.n2443 0.152939
R21678 gnd.n2445 gnd.n2444 0.152939
R21679 gnd.n2446 gnd.n2445 0.152939
R21680 gnd.n2447 gnd.n2446 0.152939
R21681 gnd.n2448 gnd.n2447 0.152939
R21682 gnd.n2449 gnd.n2448 0.152939
R21683 gnd.n3871 gnd.n2449 0.152939
R21684 gnd.n3871 gnd.n3870 0.152939
R21685 gnd.n3143 gnd.n3142 0.152939
R21686 gnd.n3143 gnd.n2847 0.152939
R21687 gnd.n3171 gnd.n2847 0.152939
R21688 gnd.n3172 gnd.n3171 0.152939
R21689 gnd.n3173 gnd.n3172 0.152939
R21690 gnd.n3174 gnd.n3173 0.152939
R21691 gnd.n3174 gnd.n2819 0.152939
R21692 gnd.n3201 gnd.n2819 0.152939
R21693 gnd.n3202 gnd.n3201 0.152939
R21694 gnd.n3203 gnd.n3202 0.152939
R21695 gnd.n3203 gnd.n2797 0.152939
R21696 gnd.n3232 gnd.n2797 0.152939
R21697 gnd.n3233 gnd.n3232 0.152939
R21698 gnd.n3234 gnd.n3233 0.152939
R21699 gnd.n3235 gnd.n3234 0.152939
R21700 gnd.n3237 gnd.n3235 0.152939
R21701 gnd.n3237 gnd.n3236 0.152939
R21702 gnd.n3236 gnd.n2746 0.152939
R21703 gnd.n2747 gnd.n2746 0.152939
R21704 gnd.n2748 gnd.n2747 0.152939
R21705 gnd.n2767 gnd.n2748 0.152939
R21706 gnd.n2768 gnd.n2767 0.152939
R21707 gnd.n2768 gnd.n2634 0.152939
R21708 gnd.n3327 gnd.n2634 0.152939
R21709 gnd.n3328 gnd.n3327 0.152939
R21710 gnd.n3329 gnd.n3328 0.152939
R21711 gnd.n3330 gnd.n3329 0.152939
R21712 gnd.n3330 gnd.n2607 0.152939
R21713 gnd.n3367 gnd.n2607 0.152939
R21714 gnd.n3368 gnd.n3367 0.152939
R21715 gnd.n3369 gnd.n3368 0.152939
R21716 gnd.n3370 gnd.n3369 0.152939
R21717 gnd.n3370 gnd.n2580 0.152939
R21718 gnd.n3412 gnd.n2580 0.152939
R21719 gnd.n3413 gnd.n3412 0.152939
R21720 gnd.n3414 gnd.n3413 0.152939
R21721 gnd.n3415 gnd.n3414 0.152939
R21722 gnd.n3415 gnd.n2552 0.152939
R21723 gnd.n3452 gnd.n2552 0.152939
R21724 gnd.n3453 gnd.n3452 0.152939
R21725 gnd.n3454 gnd.n3453 0.152939
R21726 gnd.n3455 gnd.n3454 0.152939
R21727 gnd.n3455 gnd.n2525 0.152939
R21728 gnd.n3501 gnd.n2525 0.152939
R21729 gnd.n3502 gnd.n3501 0.152939
R21730 gnd.n3503 gnd.n3502 0.152939
R21731 gnd.n3504 gnd.n3503 0.152939
R21732 gnd.n3504 gnd.n2498 0.152939
R21733 gnd.n3795 gnd.n2498 0.152939
R21734 gnd.n3796 gnd.n3795 0.152939
R21735 gnd.n3797 gnd.n3796 0.152939
R21736 gnd.n3798 gnd.n3797 0.152939
R21737 gnd.n3799 gnd.n3798 0.152939
R21738 gnd.n3141 gnd.n2871 0.152939
R21739 gnd.n2892 gnd.n2871 0.152939
R21740 gnd.n2893 gnd.n2892 0.152939
R21741 gnd.n2899 gnd.n2893 0.152939
R21742 gnd.n2900 gnd.n2899 0.152939
R21743 gnd.n2901 gnd.n2900 0.152939
R21744 gnd.n2901 gnd.n2890 0.152939
R21745 gnd.n2909 gnd.n2890 0.152939
R21746 gnd.n2910 gnd.n2909 0.152939
R21747 gnd.n2911 gnd.n2910 0.152939
R21748 gnd.n2911 gnd.n2888 0.152939
R21749 gnd.n2919 gnd.n2888 0.152939
R21750 gnd.n2920 gnd.n2919 0.152939
R21751 gnd.n2921 gnd.n2920 0.152939
R21752 gnd.n2921 gnd.n2886 0.152939
R21753 gnd.n2929 gnd.n2886 0.152939
R21754 gnd.n3868 gnd.n2454 0.152939
R21755 gnd.n2456 gnd.n2454 0.152939
R21756 gnd.n2457 gnd.n2456 0.152939
R21757 gnd.n2458 gnd.n2457 0.152939
R21758 gnd.n2459 gnd.n2458 0.152939
R21759 gnd.n2460 gnd.n2459 0.152939
R21760 gnd.n2461 gnd.n2460 0.152939
R21761 gnd.n2462 gnd.n2461 0.152939
R21762 gnd.n2463 gnd.n2462 0.152939
R21763 gnd.n2464 gnd.n2463 0.152939
R21764 gnd.n2465 gnd.n2464 0.152939
R21765 gnd.n2466 gnd.n2465 0.152939
R21766 gnd.n2467 gnd.n2466 0.152939
R21767 gnd.n2468 gnd.n2467 0.152939
R21768 gnd.n2469 gnd.n2468 0.152939
R21769 gnd.n2470 gnd.n2469 0.152939
R21770 gnd.n2471 gnd.n2470 0.152939
R21771 gnd.n2472 gnd.n2471 0.152939
R21772 gnd.n2473 gnd.n2472 0.152939
R21773 gnd.n2474 gnd.n2473 0.152939
R21774 gnd.n2475 gnd.n2474 0.152939
R21775 gnd.n2476 gnd.n2475 0.152939
R21776 gnd.n2480 gnd.n2476 0.152939
R21777 gnd.n2481 gnd.n2480 0.152939
R21778 gnd.n2482 gnd.n2481 0.152939
R21779 gnd.n2483 gnd.n2482 0.152939
R21780 gnd.n3304 gnd.n3303 0.152939
R21781 gnd.n3305 gnd.n3304 0.152939
R21782 gnd.n3306 gnd.n3305 0.152939
R21783 gnd.n3307 gnd.n3306 0.152939
R21784 gnd.n3308 gnd.n3307 0.152939
R21785 gnd.n3309 gnd.n3308 0.152939
R21786 gnd.n3309 gnd.n2588 0.152939
R21787 gnd.n3388 gnd.n2588 0.152939
R21788 gnd.n3389 gnd.n3388 0.152939
R21789 gnd.n3390 gnd.n3389 0.152939
R21790 gnd.n3391 gnd.n3390 0.152939
R21791 gnd.n3392 gnd.n3391 0.152939
R21792 gnd.n3393 gnd.n3392 0.152939
R21793 gnd.n3394 gnd.n3393 0.152939
R21794 gnd.n3395 gnd.n3394 0.152939
R21795 gnd.n3396 gnd.n3395 0.152939
R21796 gnd.n3396 gnd.n2532 0.152939
R21797 gnd.n3473 gnd.n2532 0.152939
R21798 gnd.n3474 gnd.n3473 0.152939
R21799 gnd.n3475 gnd.n3474 0.152939
R21800 gnd.n3476 gnd.n3475 0.152939
R21801 gnd.n3477 gnd.n3476 0.152939
R21802 gnd.n3478 gnd.n3477 0.152939
R21803 gnd.n3479 gnd.n3478 0.152939
R21804 gnd.n3480 gnd.n3479 0.152939
R21805 gnd.n3481 gnd.n3480 0.152939
R21806 gnd.n3483 gnd.n3481 0.152939
R21807 gnd.n3483 gnd.n3482 0.152939
R21808 gnd.n3059 gnd.n3058 0.152939
R21809 gnd.n3059 gnd.n2949 0.152939
R21810 gnd.n3074 gnd.n2949 0.152939
R21811 gnd.n3075 gnd.n3074 0.152939
R21812 gnd.n3076 gnd.n3075 0.152939
R21813 gnd.n3076 gnd.n2937 0.152939
R21814 gnd.n3090 gnd.n2937 0.152939
R21815 gnd.n3091 gnd.n3090 0.152939
R21816 gnd.n3092 gnd.n3091 0.152939
R21817 gnd.n3093 gnd.n3092 0.152939
R21818 gnd.n3094 gnd.n3093 0.152939
R21819 gnd.n3095 gnd.n3094 0.152939
R21820 gnd.n3096 gnd.n3095 0.152939
R21821 gnd.n3097 gnd.n3096 0.152939
R21822 gnd.n3098 gnd.n3097 0.152939
R21823 gnd.n3099 gnd.n3098 0.152939
R21824 gnd.n3100 gnd.n3099 0.152939
R21825 gnd.n3101 gnd.n3100 0.152939
R21826 gnd.n3102 gnd.n3101 0.152939
R21827 gnd.n3103 gnd.n3102 0.152939
R21828 gnd.n3104 gnd.n3103 0.152939
R21829 gnd.n3104 gnd.n2803 0.152939
R21830 gnd.n3221 gnd.n2803 0.152939
R21831 gnd.n3222 gnd.n3221 0.152939
R21832 gnd.n3223 gnd.n3222 0.152939
R21833 gnd.n3224 gnd.n3223 0.152939
R21834 gnd.n3224 gnd.n2725 0.152939
R21835 gnd.n3301 gnd.n2725 0.152939
R21836 gnd.n2977 gnd.n2976 0.152939
R21837 gnd.n2978 gnd.n2977 0.152939
R21838 gnd.n2979 gnd.n2978 0.152939
R21839 gnd.n2980 gnd.n2979 0.152939
R21840 gnd.n2981 gnd.n2980 0.152939
R21841 gnd.n2982 gnd.n2981 0.152939
R21842 gnd.n2983 gnd.n2982 0.152939
R21843 gnd.n2984 gnd.n2983 0.152939
R21844 gnd.n2985 gnd.n2984 0.152939
R21845 gnd.n2986 gnd.n2985 0.152939
R21846 gnd.n2987 gnd.n2986 0.152939
R21847 gnd.n2988 gnd.n2987 0.152939
R21848 gnd.n2989 gnd.n2988 0.152939
R21849 gnd.n2990 gnd.n2989 0.152939
R21850 gnd.n2991 gnd.n2990 0.152939
R21851 gnd.n2992 gnd.n2991 0.152939
R21852 gnd.n2993 gnd.n2992 0.152939
R21853 gnd.n2994 gnd.n2993 0.152939
R21854 gnd.n2995 gnd.n2994 0.152939
R21855 gnd.n2996 gnd.n2995 0.152939
R21856 gnd.n2997 gnd.n2996 0.152939
R21857 gnd.n2998 gnd.n2997 0.152939
R21858 gnd.n3002 gnd.n2998 0.152939
R21859 gnd.n3003 gnd.n3002 0.152939
R21860 gnd.n3003 gnd.n2960 0.152939
R21861 gnd.n3057 gnd.n2960 0.152939
R21862 gnd.n4210 gnd.n4149 0.152939
R21863 gnd.n4150 gnd.n4149 0.152939
R21864 gnd.n4151 gnd.n4150 0.152939
R21865 gnd.n4152 gnd.n4151 0.152939
R21866 gnd.n4153 gnd.n4152 0.152939
R21867 gnd.n4154 gnd.n4153 0.152939
R21868 gnd.n4155 gnd.n4154 0.152939
R21869 gnd.n4156 gnd.n4155 0.152939
R21870 gnd.n4157 gnd.n4156 0.152939
R21871 gnd.n4158 gnd.n4157 0.152939
R21872 gnd.n4159 gnd.n4158 0.152939
R21873 gnd.n4160 gnd.n4159 0.152939
R21874 gnd.n4161 gnd.n4160 0.152939
R21875 gnd.n4162 gnd.n4161 0.152939
R21876 gnd.n4163 gnd.n4162 0.152939
R21877 gnd.n4164 gnd.n4163 0.152939
R21878 gnd.n4165 gnd.n4164 0.152939
R21879 gnd.n4166 gnd.n4165 0.152939
R21880 gnd.n4167 gnd.n4166 0.152939
R21881 gnd.n4168 gnd.n4167 0.152939
R21882 gnd.n4169 gnd.n4168 0.152939
R21883 gnd.n4170 gnd.n4169 0.152939
R21884 gnd.n4171 gnd.n4170 0.152939
R21885 gnd.n4172 gnd.n4171 0.152939
R21886 gnd.n4172 gnd.n2293 0.152939
R21887 gnd.n4399 gnd.n2293 0.152939
R21888 gnd.n4400 gnd.n4399 0.152939
R21889 gnd.n4401 gnd.n4400 0.152939
R21890 gnd.n4402 gnd.n4401 0.152939
R21891 gnd.n4402 gnd.n2268 0.152939
R21892 gnd.n4434 gnd.n2268 0.152939
R21893 gnd.n1786 gnd.n1780 0.152939
R21894 gnd.n1787 gnd.n1786 0.152939
R21895 gnd.n1788 gnd.n1787 0.152939
R21896 gnd.n1788 gnd.n1775 0.152939
R21897 gnd.n1796 gnd.n1775 0.152939
R21898 gnd.n1797 gnd.n1796 0.152939
R21899 gnd.n1798 gnd.n1797 0.152939
R21900 gnd.n1798 gnd.n1771 0.152939
R21901 gnd.n1806 gnd.n1771 0.152939
R21902 gnd.n1807 gnd.n1806 0.152939
R21903 gnd.n1808 gnd.n1807 0.152939
R21904 gnd.n1808 gnd.n1767 0.152939
R21905 gnd.n1816 gnd.n1767 0.152939
R21906 gnd.n1817 gnd.n1816 0.152939
R21907 gnd.n1818 gnd.n1817 0.152939
R21908 gnd.n1818 gnd.n1763 0.152939
R21909 gnd.n1825 gnd.n1763 0.152939
R21910 gnd.n1826 gnd.n1825 0.152939
R21911 gnd.n1826 gnd.n1757 0.152939
R21912 gnd.n1834 gnd.n1757 0.152939
R21913 gnd.n1835 gnd.n1834 0.152939
R21914 gnd.n1836 gnd.n1835 0.152939
R21915 gnd.n1836 gnd.n1753 0.152939
R21916 gnd.n1845 gnd.n1753 0.152939
R21917 gnd.n1846 gnd.n1845 0.152939
R21918 gnd.n1950 gnd.n1949 0.152939
R21919 gnd.n1949 gnd.n1847 0.152939
R21920 gnd.n1853 gnd.n1847 0.152939
R21921 gnd.n1854 gnd.n1853 0.152939
R21922 gnd.n1855 gnd.n1854 0.152939
R21923 gnd.n1856 gnd.n1855 0.152939
R21924 gnd.n1860 gnd.n1856 0.152939
R21925 gnd.n1861 gnd.n1860 0.152939
R21926 gnd.n1932 gnd.n1861 0.152939
R21927 gnd.n1932 gnd.n1931 0.152939
R21928 gnd.n1931 gnd.n1930 0.152939
R21929 gnd.n1930 gnd.n1865 0.152939
R21930 gnd.n1871 gnd.n1865 0.152939
R21931 gnd.n1872 gnd.n1871 0.152939
R21932 gnd.n1873 gnd.n1872 0.152939
R21933 gnd.n1874 gnd.n1873 0.152939
R21934 gnd.n1878 gnd.n1874 0.152939
R21935 gnd.n1879 gnd.n1878 0.152939
R21936 gnd.n1880 gnd.n1879 0.152939
R21937 gnd.n1881 gnd.n1880 0.152939
R21938 gnd.n1885 gnd.n1881 0.152939
R21939 gnd.n1886 gnd.n1885 0.152939
R21940 gnd.n1887 gnd.n1886 0.152939
R21941 gnd.n1888 gnd.n1887 0.152939
R21942 gnd.n1892 gnd.n1888 0.152939
R21943 gnd.n1893 gnd.n1892 0.152939
R21944 gnd.n1894 gnd.n1893 0.152939
R21945 gnd.n1895 gnd.n1894 0.152939
R21946 gnd.n1895 gnd.n837 0.152939
R21947 gnd.n6404 gnd.n837 0.152939
R21948 gnd.n4461 gnd.n2225 0.152939
R21949 gnd.n4492 gnd.n2225 0.152939
R21950 gnd.n4493 gnd.n4492 0.152939
R21951 gnd.n4494 gnd.n4493 0.152939
R21952 gnd.n4495 gnd.n4494 0.152939
R21953 gnd.n4495 gnd.n2199 0.152939
R21954 gnd.n4527 gnd.n2199 0.152939
R21955 gnd.n4528 gnd.n4527 0.152939
R21956 gnd.n4529 gnd.n4528 0.152939
R21957 gnd.n4531 gnd.n4529 0.152939
R21958 gnd.n4531 gnd.n4530 0.152939
R21959 gnd.n4530 gnd.n760 0.152939
R21960 gnd.n761 gnd.n760 0.152939
R21961 gnd.n762 gnd.n761 0.152939
R21962 gnd.n782 gnd.n762 0.152939
R21963 gnd.n783 gnd.n782 0.152939
R21964 gnd.n784 gnd.n783 0.152939
R21965 gnd.n785 gnd.n784 0.152939
R21966 gnd.n802 gnd.n785 0.152939
R21967 gnd.n803 gnd.n802 0.152939
R21968 gnd.n804 gnd.n803 0.152939
R21969 gnd.n805 gnd.n804 0.152939
R21970 gnd.n823 gnd.n805 0.152939
R21971 gnd.n824 gnd.n823 0.152939
R21972 gnd.n825 gnd.n824 0.152939
R21973 gnd.n826 gnd.n825 0.152939
R21974 gnd.n1779 gnd.n826 0.152939
R21975 gnd.n4266 gnd.n4265 0.152939
R21976 gnd.n4267 gnd.n4266 0.152939
R21977 gnd.n4267 gnd.n2393 0.152939
R21978 gnd.n4285 gnd.n2393 0.152939
R21979 gnd.n4286 gnd.n4285 0.152939
R21980 gnd.n4287 gnd.n4286 0.152939
R21981 gnd.n4287 gnd.n2374 0.152939
R21982 gnd.n4305 gnd.n2374 0.152939
R21983 gnd.n4306 gnd.n4305 0.152939
R21984 gnd.n4307 gnd.n4306 0.152939
R21985 gnd.n4307 gnd.n2357 0.152939
R21986 gnd.n4325 gnd.n2357 0.152939
R21987 gnd.n4326 gnd.n4325 0.152939
R21988 gnd.n4327 gnd.n4326 0.152939
R21989 gnd.n4327 gnd.n2338 0.152939
R21990 gnd.n4345 gnd.n2338 0.152939
R21991 gnd.n4346 gnd.n4345 0.152939
R21992 gnd.n4347 gnd.n4346 0.152939
R21993 gnd.n4347 gnd.n2321 0.152939
R21994 gnd.n4365 gnd.n2321 0.152939
R21995 gnd.n4366 gnd.n4365 0.152939
R21996 gnd.n4367 gnd.n4366 0.152939
R21997 gnd.n4367 gnd.n2301 0.152939
R21998 gnd.n4389 gnd.n2301 0.152939
R21999 gnd.n4390 gnd.n4389 0.152939
R22000 gnd.n4391 gnd.n4390 0.152939
R22001 gnd.n4392 gnd.n4391 0.152939
R22002 gnd.n3978 gnd.n2410 0.152939
R22003 gnd.n3979 gnd.n3978 0.152939
R22004 gnd.n3980 gnd.n3979 0.152939
R22005 gnd.n3980 gnd.n3970 0.152939
R22006 gnd.n3988 gnd.n3970 0.152939
R22007 gnd.n3989 gnd.n3988 0.152939
R22008 gnd.n3990 gnd.n3989 0.152939
R22009 gnd.n3990 gnd.n3966 0.152939
R22010 gnd.n3998 gnd.n3966 0.152939
R22011 gnd.n3999 gnd.n3998 0.152939
R22012 gnd.n4000 gnd.n3999 0.152939
R22013 gnd.n4000 gnd.n3962 0.152939
R22014 gnd.n4008 gnd.n3962 0.152939
R22015 gnd.n4009 gnd.n4008 0.152939
R22016 gnd.n4010 gnd.n4009 0.152939
R22017 gnd.n4010 gnd.n3955 0.152939
R22018 gnd.n4018 gnd.n3955 0.152939
R22019 gnd.n4019 gnd.n4018 0.152939
R22020 gnd.n4020 gnd.n4019 0.152939
R22021 gnd.n4020 gnd.n3951 0.152939
R22022 gnd.n4028 gnd.n3951 0.152939
R22023 gnd.n4029 gnd.n4028 0.152939
R22024 gnd.n4030 gnd.n4029 0.152939
R22025 gnd.n4030 gnd.n3947 0.152939
R22026 gnd.n4038 gnd.n3947 0.152939
R22027 gnd.n4039 gnd.n4038 0.152939
R22028 gnd.n4040 gnd.n4039 0.152939
R22029 gnd.n4040 gnd.n3943 0.152939
R22030 gnd.n4048 gnd.n3943 0.152939
R22031 gnd.n4049 gnd.n4048 0.152939
R22032 gnd.n4050 gnd.n4049 0.152939
R22033 gnd.n4050 gnd.n3939 0.152939
R22034 gnd.n4058 gnd.n3939 0.152939
R22035 gnd.n4059 gnd.n4058 0.152939
R22036 gnd.n4060 gnd.n4059 0.152939
R22037 gnd.n4060 gnd.n3935 0.152939
R22038 gnd.n4070 gnd.n3935 0.152939
R22039 gnd.n4071 gnd.n4070 0.152939
R22040 gnd.n4072 gnd.n4071 0.152939
R22041 gnd.n4072 gnd.n3931 0.152939
R22042 gnd.n4080 gnd.n3931 0.152939
R22043 gnd.n4081 gnd.n4080 0.152939
R22044 gnd.n4082 gnd.n4081 0.152939
R22045 gnd.n4082 gnd.n3927 0.152939
R22046 gnd.n4090 gnd.n3927 0.152939
R22047 gnd.n4091 gnd.n4090 0.152939
R22048 gnd.n4092 gnd.n4091 0.152939
R22049 gnd.n4092 gnd.n3923 0.152939
R22050 gnd.n4100 gnd.n3923 0.152939
R22051 gnd.n4101 gnd.n4100 0.152939
R22052 gnd.n4102 gnd.n4101 0.152939
R22053 gnd.n4102 gnd.n3919 0.152939
R22054 gnd.n4110 gnd.n3919 0.152939
R22055 gnd.n4111 gnd.n4110 0.152939
R22056 gnd.n4113 gnd.n4111 0.152939
R22057 gnd.n4113 gnd.n4112 0.152939
R22058 gnd.n4112 gnd.n3912 0.152939
R22059 gnd.n4122 gnd.n3912 0.152939
R22060 gnd.n4251 gnd.n4123 0.152939
R22061 gnd.n4126 gnd.n4123 0.152939
R22062 gnd.n4127 gnd.n4126 0.152939
R22063 gnd.n4128 gnd.n4127 0.152939
R22064 gnd.n4129 gnd.n4128 0.152939
R22065 gnd.n4132 gnd.n4129 0.152939
R22066 gnd.n4133 gnd.n4132 0.152939
R22067 gnd.n4134 gnd.n4133 0.152939
R22068 gnd.n4135 gnd.n4134 0.152939
R22069 gnd.n4138 gnd.n4135 0.152939
R22070 gnd.n4139 gnd.n4138 0.152939
R22071 gnd.n4140 gnd.n4139 0.152939
R22072 gnd.n4141 gnd.n4140 0.152939
R22073 gnd.n4144 gnd.n4141 0.152939
R22074 gnd.n4145 gnd.n4144 0.152939
R22075 gnd.n4217 gnd.n4145 0.152939
R22076 gnd.n4217 gnd.n4216 0.152939
R22077 gnd.n4216 gnd.n4215 0.152939
R22078 gnd.n6382 gnd.n6381 0.152939
R22079 gnd.n6381 gnd.n6380 0.152939
R22080 gnd.n6380 gnd.n868 0.152939
R22081 gnd.n6376 gnd.n868 0.152939
R22082 gnd.n6376 gnd.n6375 0.152939
R22083 gnd.n6375 gnd.n6374 0.152939
R22084 gnd.n6374 gnd.n873 0.152939
R22085 gnd.n6370 gnd.n873 0.152939
R22086 gnd.n6370 gnd.n6369 0.152939
R22087 gnd.n6369 gnd.n6368 0.152939
R22088 gnd.n6368 gnd.n878 0.152939
R22089 gnd.n6364 gnd.n878 0.152939
R22090 gnd.n6364 gnd.n6363 0.152939
R22091 gnd.n6363 gnd.n6362 0.152939
R22092 gnd.n6362 gnd.n883 0.152939
R22093 gnd.n6358 gnd.n883 0.152939
R22094 gnd.n6358 gnd.n6357 0.152939
R22095 gnd.n6357 gnd.n6356 0.152939
R22096 gnd.n6356 gnd.n888 0.152939
R22097 gnd.n6352 gnd.n888 0.152939
R22098 gnd.n6352 gnd.n6351 0.152939
R22099 gnd.n6351 gnd.n6350 0.152939
R22100 gnd.n6350 gnd.n893 0.152939
R22101 gnd.n6346 gnd.n893 0.152939
R22102 gnd.n6346 gnd.n6345 0.152939
R22103 gnd.n6345 gnd.n6344 0.152939
R22104 gnd.n6344 gnd.n898 0.152939
R22105 gnd.n6340 gnd.n898 0.152939
R22106 gnd.n6340 gnd.n6339 0.152939
R22107 gnd.n6339 gnd.n6338 0.152939
R22108 gnd.n6338 gnd.n903 0.152939
R22109 gnd.n6334 gnd.n903 0.152939
R22110 gnd.n6334 gnd.n6333 0.152939
R22111 gnd.n6333 gnd.n6332 0.152939
R22112 gnd.n6332 gnd.n908 0.152939
R22113 gnd.n6328 gnd.n908 0.152939
R22114 gnd.n6328 gnd.n6327 0.152939
R22115 gnd.n6327 gnd.n6326 0.152939
R22116 gnd.n6326 gnd.n913 0.152939
R22117 gnd.n6322 gnd.n913 0.152939
R22118 gnd.n6322 gnd.n6321 0.152939
R22119 gnd.n6321 gnd.n6320 0.152939
R22120 gnd.n6320 gnd.n918 0.152939
R22121 gnd.n6316 gnd.n918 0.152939
R22122 gnd.n6316 gnd.n6315 0.152939
R22123 gnd.n6315 gnd.n6314 0.152939
R22124 gnd.n6314 gnd.n923 0.152939
R22125 gnd.n6310 gnd.n923 0.152939
R22126 gnd.n6310 gnd.n6309 0.152939
R22127 gnd.n6309 gnd.n6308 0.152939
R22128 gnd.n6308 gnd.n928 0.152939
R22129 gnd.n6304 gnd.n928 0.152939
R22130 gnd.n6304 gnd.n6303 0.152939
R22131 gnd.n6303 gnd.n6302 0.152939
R22132 gnd.n6302 gnd.n933 0.152939
R22133 gnd.n6298 gnd.n933 0.152939
R22134 gnd.n6298 gnd.n6297 0.152939
R22135 gnd.n6297 gnd.n6296 0.152939
R22136 gnd.n6296 gnd.n938 0.152939
R22137 gnd.n6292 gnd.n938 0.152939
R22138 gnd.n6292 gnd.n6291 0.152939
R22139 gnd.n6291 gnd.n6290 0.152939
R22140 gnd.n6290 gnd.n943 0.152939
R22141 gnd.n6286 gnd.n943 0.152939
R22142 gnd.n6286 gnd.n6285 0.152939
R22143 gnd.n6285 gnd.n6284 0.152939
R22144 gnd.n6284 gnd.n948 0.152939
R22145 gnd.n6280 gnd.n948 0.152939
R22146 gnd.n6280 gnd.n6279 0.152939
R22147 gnd.n6279 gnd.n6278 0.152939
R22148 gnd.n6278 gnd.n953 0.152939
R22149 gnd.n6274 gnd.n953 0.152939
R22150 gnd.n6274 gnd.n6273 0.152939
R22151 gnd.n6273 gnd.n6272 0.152939
R22152 gnd.n6272 gnd.n958 0.152939
R22153 gnd.n6268 gnd.n958 0.152939
R22154 gnd.n6268 gnd.n6267 0.152939
R22155 gnd.n6267 gnd.n6266 0.152939
R22156 gnd.n6266 gnd.n963 0.152939
R22157 gnd.n6262 gnd.n963 0.152939
R22158 gnd.n6262 gnd.n6261 0.152939
R22159 gnd.n6261 gnd.n6260 0.152939
R22160 gnd.n6260 gnd.n968 0.152939
R22161 gnd.n6256 gnd.n968 0.152939
R22162 gnd.n6256 gnd.n6255 0.152939
R22163 gnd.n6255 gnd.n6254 0.152939
R22164 gnd.n6254 gnd.n973 0.152939
R22165 gnd.n6250 gnd.n973 0.152939
R22166 gnd.n6250 gnd.n6249 0.152939
R22167 gnd.n6249 gnd.n6248 0.152939
R22168 gnd.n6248 gnd.n978 0.152939
R22169 gnd.n6244 gnd.n978 0.152939
R22170 gnd.n6244 gnd.n6243 0.152939
R22171 gnd.n6243 gnd.n6242 0.152939
R22172 gnd.n6242 gnd.n983 0.152939
R22173 gnd.n6238 gnd.n983 0.152939
R22174 gnd.n6238 gnd.n6237 0.152939
R22175 gnd.n6237 gnd.n6236 0.152939
R22176 gnd.n6236 gnd.n988 0.152939
R22177 gnd.n6232 gnd.n988 0.152939
R22178 gnd.n6232 gnd.n6231 0.152939
R22179 gnd.n4437 gnd.n4436 0.152939
R22180 gnd.n4436 gnd.n2242 0.152939
R22181 gnd.n4468 gnd.n2242 0.152939
R22182 gnd.n4469 gnd.n4468 0.152939
R22183 gnd.n4471 gnd.n4469 0.152939
R22184 gnd.n4471 gnd.n4470 0.152939
R22185 gnd.n4470 gnd.n2216 0.152939
R22186 gnd.n4502 gnd.n2216 0.152939
R22187 gnd.n4503 gnd.n4502 0.152939
R22188 gnd.n4505 gnd.n4503 0.152939
R22189 gnd.n4505 gnd.n4504 0.152939
R22190 gnd.n4504 gnd.n2190 0.152939
R22191 gnd.n4538 gnd.n2190 0.152939
R22192 gnd.n4539 gnd.n4538 0.152939
R22193 gnd.n4544 gnd.n4539 0.152939
R22194 gnd.n4544 gnd.n4543 0.152939
R22195 gnd.n4543 gnd.n4542 0.152939
R22196 gnd.n4542 gnd.n2179 0.152939
R22197 gnd.n4561 gnd.n2179 0.152939
R22198 gnd.n4562 gnd.n4561 0.152939
R22199 gnd.n4563 gnd.n4562 0.152939
R22200 gnd.n4563 gnd.n2174 0.152939
R22201 gnd.n4911 gnd.n2174 0.152939
R22202 gnd.n4912 gnd.n4911 0.152939
R22203 gnd.n4913 gnd.n4912 0.152939
R22204 gnd.n4913 gnd.n2169 0.152939
R22205 gnd.n4931 gnd.n2169 0.152939
R22206 gnd.n4932 gnd.n4931 0.152939
R22207 gnd.n4933 gnd.n4932 0.152939
R22208 gnd.n4933 gnd.n2166 0.152939
R22209 gnd.n4937 gnd.n2166 0.152939
R22210 gnd.n5009 gnd.n2067 0.152939
R22211 gnd.n5002 gnd.n2067 0.152939
R22212 gnd.n5002 gnd.n5001 0.152939
R22213 gnd.n5001 gnd.n5000 0.152939
R22214 gnd.n5000 gnd.n2071 0.152939
R22215 gnd.n4996 gnd.n2071 0.152939
R22216 gnd.n5011 gnd.n5010 0.152939
R22217 gnd.n5011 gnd.n2064 0.152939
R22218 gnd.n5026 gnd.n2064 0.152939
R22219 gnd.n5027 gnd.n5026 0.152939
R22220 gnd.n5028 gnd.n5027 0.152939
R22221 gnd.n5028 gnd.n2053 0.152939
R22222 gnd.n5044 gnd.n2053 0.152939
R22223 gnd.n5045 gnd.n5044 0.152939
R22224 gnd.n5046 gnd.n5045 0.152939
R22225 gnd.n5046 gnd.n2041 0.152939
R22226 gnd.n5061 gnd.n2041 0.152939
R22227 gnd.n5062 gnd.n5061 0.152939
R22228 gnd.n5063 gnd.n5062 0.152939
R22229 gnd.n5063 gnd.n2028 0.152939
R22230 gnd.n5080 gnd.n2028 0.152939
R22231 gnd.n5081 gnd.n5080 0.152939
R22232 gnd.n5146 gnd.n5081 0.152939
R22233 gnd.n5146 gnd.n5145 0.152939
R22234 gnd.n5145 gnd.n5144 0.152939
R22235 gnd.n5144 gnd.n5082 0.152939
R22236 gnd.n5140 gnd.n5082 0.152939
R22237 gnd.n5140 gnd.n5139 0.152939
R22238 gnd.n5139 gnd.n5138 0.152939
R22239 gnd.n5138 gnd.n5086 0.152939
R22240 gnd.n5134 gnd.n5086 0.152939
R22241 gnd.n5134 gnd.n5133 0.152939
R22242 gnd.n5133 gnd.n5132 0.152939
R22243 gnd.n5132 gnd.n5091 0.152939
R22244 gnd.n5128 gnd.n5091 0.152939
R22245 gnd.n5128 gnd.n5127 0.152939
R22246 gnd.n5127 gnd.n5126 0.152939
R22247 gnd.n5126 gnd.n5095 0.152939
R22248 gnd.n5122 gnd.n5095 0.152939
R22249 gnd.n5122 gnd.n5121 0.152939
R22250 gnd.n5121 gnd.n5120 0.152939
R22251 gnd.n5120 gnd.n5099 0.152939
R22252 gnd.n5116 gnd.n5099 0.152939
R22253 gnd.n5116 gnd.n5115 0.152939
R22254 gnd.n5115 gnd.n5114 0.152939
R22255 gnd.n5114 gnd.n5103 0.152939
R22256 gnd.n5110 gnd.n5103 0.152939
R22257 gnd.n5110 gnd.n5109 0.152939
R22258 gnd.n5109 gnd.n5108 0.152939
R22259 gnd.n5108 gnd.n1491 0.152939
R22260 gnd.n5371 gnd.n1491 0.152939
R22261 gnd.n5372 gnd.n5371 0.152939
R22262 gnd.n5387 gnd.n5372 0.152939
R22263 gnd.n5387 gnd.n5386 0.152939
R22264 gnd.n5386 gnd.n5385 0.152939
R22265 gnd.n5385 gnd.n5373 0.152939
R22266 gnd.n5381 gnd.n5373 0.152939
R22267 gnd.n5381 gnd.n5380 0.152939
R22268 gnd.n5380 gnd.n5379 0.152939
R22269 gnd.n5379 gnd.n1441 0.152939
R22270 gnd.n5468 gnd.n1441 0.152939
R22271 gnd.n5469 gnd.n5468 0.152939
R22272 gnd.n5481 gnd.n5469 0.152939
R22273 gnd.n5481 gnd.n5480 0.152939
R22274 gnd.n5480 gnd.n5479 0.152939
R22275 gnd.n5479 gnd.n5470 0.152939
R22276 gnd.n5475 gnd.n5470 0.152939
R22277 gnd.n5475 gnd.n5474 0.152939
R22278 gnd.n5474 gnd.n1391 0.152939
R22279 gnd.n5544 gnd.n1391 0.152939
R22280 gnd.n5545 gnd.n5544 0.152939
R22281 gnd.n5550 gnd.n5545 0.152939
R22282 gnd.n5550 gnd.n5549 0.152939
R22283 gnd.n5549 gnd.n5548 0.152939
R22284 gnd.n5548 gnd.n5546 0.152939
R22285 gnd.n5546 gnd.n1366 0.152939
R22286 gnd.n5589 gnd.n1366 0.152939
R22287 gnd.n5590 gnd.n5589 0.152939
R22288 gnd.n5610 gnd.n5590 0.152939
R22289 gnd.n5610 gnd.n5609 0.152939
R22290 gnd.n5609 gnd.n5608 0.152939
R22291 gnd.n5608 gnd.n5591 0.152939
R22292 gnd.n5604 gnd.n5591 0.152939
R22293 gnd.n5604 gnd.n5603 0.152939
R22294 gnd.n5603 gnd.n5602 0.152939
R22295 gnd.n5602 gnd.n5596 0.152939
R22296 gnd.n5598 gnd.n5596 0.152939
R22297 gnd.n5598 gnd.n1216 0.152939
R22298 gnd.n5821 gnd.n1216 0.152939
R22299 gnd.n5822 gnd.n5821 0.152939
R22300 gnd.n5823 gnd.n5822 0.152939
R22301 gnd.n5823 gnd.n1205 0.152939
R22302 gnd.n5838 gnd.n1205 0.152939
R22303 gnd.n5839 gnd.n5838 0.152939
R22304 gnd.n5840 gnd.n5839 0.152939
R22305 gnd.n5840 gnd.n1193 0.152939
R22306 gnd.n5855 gnd.n1193 0.152939
R22307 gnd.n5856 gnd.n5855 0.152939
R22308 gnd.n5857 gnd.n5856 0.152939
R22309 gnd.n5857 gnd.n1182 0.152939
R22310 gnd.n5873 gnd.n1182 0.152939
R22311 gnd.n5874 gnd.n5873 0.152939
R22312 gnd.n5875 gnd.n5874 0.152939
R22313 gnd.n5875 gnd.n1170 0.152939
R22314 gnd.n5892 gnd.n1170 0.152939
R22315 gnd.n5893 gnd.n5892 0.152939
R22316 gnd.n5912 gnd.n5893 0.152939
R22317 gnd.n5911 gnd.n5894 0.152939
R22318 gnd.n5907 gnd.n5894 0.152939
R22319 gnd.n5907 gnd.n5906 0.152939
R22320 gnd.n5906 gnd.n5905 0.152939
R22321 gnd.n5905 gnd.n5898 0.152939
R22322 gnd.n5898 gnd.n1139 0.152939
R22323 gnd.n5969 gnd.n5968 0.152939
R22324 gnd.n5969 gnd.n5966 0.152939
R22325 gnd.n5975 gnd.n5966 0.152939
R22326 gnd.n5976 gnd.n5975 0.152939
R22327 gnd.n5978 gnd.n5976 0.152939
R22328 gnd.n5978 gnd.n5977 0.152939
R22329 gnd.n5977 gnd.n378 0.152939
R22330 gnd.n7064 gnd.n378 0.152939
R22331 gnd.n7065 gnd.n7064 0.152939
R22332 gnd.n7067 gnd.n7065 0.152939
R22333 gnd.n7067 gnd.n7066 0.152939
R22334 gnd.n7066 gnd.n349 0.152939
R22335 gnd.n7100 gnd.n349 0.152939
R22336 gnd.n7101 gnd.n7100 0.152939
R22337 gnd.n7123 gnd.n7101 0.152939
R22338 gnd.n7123 gnd.n7122 0.152939
R22339 gnd.n7122 gnd.n7121 0.152939
R22340 gnd.n7121 gnd.n7102 0.152939
R22341 gnd.n7117 gnd.n7102 0.152939
R22342 gnd.n7117 gnd.n7116 0.152939
R22343 gnd.n7116 gnd.n7115 0.152939
R22344 gnd.n7115 gnd.n7106 0.152939
R22345 gnd.n7111 gnd.n7106 0.152939
R22346 gnd.n7111 gnd.n7110 0.152939
R22347 gnd.n7110 gnd.n287 0.152939
R22348 gnd.n7194 gnd.n287 0.152939
R22349 gnd.n7195 gnd.n7194 0.152939
R22350 gnd.n7201 gnd.n7195 0.152939
R22351 gnd.n7201 gnd.n7200 0.152939
R22352 gnd.n7200 gnd.n7199 0.152939
R22353 gnd.n7199 gnd.n99 0.152939
R22354 gnd.n7740 gnd.n7739 0.145814
R22355 gnd.n4435 gnd.n4434 0.145814
R22356 gnd.n4437 gnd.n4435 0.145814
R22357 gnd.n7740 gnd.n99 0.145814
R22358 gnd.n4996 gnd.n836 0.128549
R22359 gnd.n6098 gnd.n1139 0.128549
R22360 gnd.n3303 gnd.n3302 0.0767195
R22361 gnd.n3302 gnd.n3301 0.0767195
R22362 gnd.n6405 gnd.n836 0.063
R22363 gnd.n6099 gnd.n6098 0.063
R22364 gnd.n3869 gnd.n2453 0.0477147
R22365 gnd.n3066 gnd.n2954 0.0442063
R22366 gnd.n3067 gnd.n3066 0.0442063
R22367 gnd.n3068 gnd.n3067 0.0442063
R22368 gnd.n3068 gnd.n2943 0.0442063
R22369 gnd.n3082 gnd.n2943 0.0442063
R22370 gnd.n3083 gnd.n3082 0.0442063
R22371 gnd.n3084 gnd.n3083 0.0442063
R22372 gnd.n3084 gnd.n2930 0.0442063
R22373 gnd.n3128 gnd.n2930 0.0442063
R22374 gnd.n3129 gnd.n3128 0.0442063
R22375 gnd.n6099 gnd.n1138 0.0416005
R22376 gnd.n7642 gnd.n7641 0.0416005
R22377 gnd.n4253 gnd.n4252 0.0416005
R22378 gnd.n6406 gnd.n6405 0.0416005
R22379 gnd.n5954 gnd.n1138 0.0344674
R22380 gnd.n5958 gnd.n5954 0.0344674
R22381 gnd.n5958 gnd.n5951 0.0344674
R22382 gnd.n5985 gnd.n5951 0.0344674
R22383 gnd.n5985 gnd.n5984 0.0344674
R22384 gnd.n5984 gnd.n397 0.0344674
R22385 gnd.n398 gnd.n397 0.0344674
R22386 gnd.n7042 gnd.n398 0.0344674
R22387 gnd.n7043 gnd.n7042 0.0344674
R22388 gnd.n7043 gnd.n372 0.0344674
R22389 gnd.n372 gnd.n369 0.0344674
R22390 gnd.n370 gnd.n369 0.0344674
R22391 gnd.n7078 gnd.n370 0.0344674
R22392 gnd.n7079 gnd.n7078 0.0344674
R22393 gnd.n7079 gnd.n344 0.0344674
R22394 gnd.n344 gnd.n342 0.0344674
R22395 gnd.n7131 gnd.n342 0.0344674
R22396 gnd.n7132 gnd.n7131 0.0344674
R22397 gnd.n7132 gnd.n326 0.0344674
R22398 gnd.n326 gnd.n324 0.0344674
R22399 gnd.n7151 gnd.n324 0.0344674
R22400 gnd.n7152 gnd.n7151 0.0344674
R22401 gnd.n7152 gnd.n308 0.0344674
R22402 gnd.n308 gnd.n305 0.0344674
R22403 gnd.n306 gnd.n305 0.0344674
R22404 gnd.n7173 gnd.n306 0.0344674
R22405 gnd.n7174 gnd.n7173 0.0344674
R22406 gnd.n7174 gnd.n280 0.0344674
R22407 gnd.n7210 gnd.n280 0.0344674
R22408 gnd.n7210 gnd.n263 0.0344674
R22409 gnd.n7227 gnd.n263 0.0344674
R22410 gnd.n7228 gnd.n7227 0.0344674
R22411 gnd.n7228 gnd.n257 0.0344674
R22412 gnd.n7236 gnd.n257 0.0344674
R22413 gnd.n7237 gnd.n7236 0.0344674
R22414 gnd.n7237 gnd.n122 0.0344674
R22415 gnd.n123 gnd.n122 0.0344674
R22416 gnd.n124 gnd.n123 0.0344674
R22417 gnd.n7244 gnd.n124 0.0344674
R22418 gnd.n7244 gnd.n141 0.0344674
R22419 gnd.n142 gnd.n141 0.0344674
R22420 gnd.n143 gnd.n142 0.0344674
R22421 gnd.n7251 gnd.n143 0.0344674
R22422 gnd.n7251 gnd.n160 0.0344674
R22423 gnd.n161 gnd.n160 0.0344674
R22424 gnd.n162 gnd.n161 0.0344674
R22425 gnd.n7258 gnd.n162 0.0344674
R22426 gnd.n7258 gnd.n180 0.0344674
R22427 gnd.n181 gnd.n180 0.0344674
R22428 gnd.n182 gnd.n181 0.0344674
R22429 gnd.n7265 gnd.n182 0.0344674
R22430 gnd.n7265 gnd.n199 0.0344674
R22431 gnd.n200 gnd.n199 0.0344674
R22432 gnd.n201 gnd.n200 0.0344674
R22433 gnd.n7272 gnd.n201 0.0344674
R22434 gnd.n7272 gnd.n218 0.0344674
R22435 gnd.n219 gnd.n218 0.0344674
R22436 gnd.n220 gnd.n219 0.0344674
R22437 gnd.n7279 gnd.n220 0.0344674
R22438 gnd.n7279 gnd.n237 0.0344674
R22439 gnd.n238 gnd.n237 0.0344674
R22440 gnd.n239 gnd.n238 0.0344674
R22441 gnd.n255 gnd.n239 0.0344674
R22442 gnd.n7642 gnd.n255 0.0344674
R22443 gnd.n3131 gnd.n2864 0.0344674
R22444 gnd.n4256 gnd.n4253 0.0344674
R22445 gnd.n4257 gnd.n4256 0.0344674
R22446 gnd.n4257 gnd.n2404 0.0344674
R22447 gnd.n2404 gnd.n2402 0.0344674
R22448 gnd.n4276 gnd.n2402 0.0344674
R22449 gnd.n4277 gnd.n4276 0.0344674
R22450 gnd.n4277 gnd.n2386 0.0344674
R22451 gnd.n2386 gnd.n2384 0.0344674
R22452 gnd.n4296 gnd.n2384 0.0344674
R22453 gnd.n4297 gnd.n4296 0.0344674
R22454 gnd.n4297 gnd.n2368 0.0344674
R22455 gnd.n2368 gnd.n2366 0.0344674
R22456 gnd.n4316 gnd.n2366 0.0344674
R22457 gnd.n4317 gnd.n4316 0.0344674
R22458 gnd.n4317 gnd.n2350 0.0344674
R22459 gnd.n2350 gnd.n2348 0.0344674
R22460 gnd.n4336 gnd.n2348 0.0344674
R22461 gnd.n4337 gnd.n4336 0.0344674
R22462 gnd.n4337 gnd.n2332 0.0344674
R22463 gnd.n2332 gnd.n2330 0.0344674
R22464 gnd.n4356 gnd.n2330 0.0344674
R22465 gnd.n4357 gnd.n4356 0.0344674
R22466 gnd.n4357 gnd.n2314 0.0344674
R22467 gnd.n2314 gnd.n2311 0.0344674
R22468 gnd.n2312 gnd.n2311 0.0344674
R22469 gnd.n4378 gnd.n2312 0.0344674
R22470 gnd.n4379 gnd.n4378 0.0344674
R22471 gnd.n4379 gnd.n2288 0.0344674
R22472 gnd.n2288 gnd.n2285 0.0344674
R22473 gnd.n2286 gnd.n2285 0.0344674
R22474 gnd.n4413 gnd.n2286 0.0344674
R22475 gnd.n4414 gnd.n4413 0.0344674
R22476 gnd.n4414 gnd.n2262 0.0344674
R22477 gnd.n2262 gnd.n2259 0.0344674
R22478 gnd.n2260 gnd.n2259 0.0344674
R22479 gnd.n4447 gnd.n2260 0.0344674
R22480 gnd.n4448 gnd.n4447 0.0344674
R22481 gnd.n4448 gnd.n2236 0.0344674
R22482 gnd.n2236 gnd.n2233 0.0344674
R22483 gnd.n2234 gnd.n2233 0.0344674
R22484 gnd.n4481 gnd.n2234 0.0344674
R22485 gnd.n4482 gnd.n4481 0.0344674
R22486 gnd.n4482 gnd.n2210 0.0344674
R22487 gnd.n2210 gnd.n2207 0.0344674
R22488 gnd.n2208 gnd.n2207 0.0344674
R22489 gnd.n4519 gnd.n2208 0.0344674
R22490 gnd.n4519 gnd.n4518 0.0344674
R22491 gnd.n4518 gnd.n2182 0.0344674
R22492 gnd.n4551 gnd.n2182 0.0344674
R22493 gnd.n4552 gnd.n4551 0.0344674
R22494 gnd.n4552 gnd.n772 0.0344674
R22495 gnd.n773 gnd.n772 0.0344674
R22496 gnd.n774 gnd.n773 0.0344674
R22497 gnd.n2177 gnd.n774 0.0344674
R22498 gnd.n2177 gnd.n792 0.0344674
R22499 gnd.n793 gnd.n792 0.0344674
R22500 gnd.n794 gnd.n793 0.0344674
R22501 gnd.n2172 gnd.n794 0.0344674
R22502 gnd.n2172 gnd.n813 0.0344674
R22503 gnd.n814 gnd.n813 0.0344674
R22504 gnd.n815 gnd.n814 0.0344674
R22505 gnd.n4920 gnd.n815 0.0344674
R22506 gnd.n4920 gnd.n834 0.0344674
R22507 gnd.n6406 gnd.n834 0.0344674
R22508 gnd.n4994 gnd.n4993 0.0343753
R22509 gnd.n6097 gnd.n1140 0.0343753
R22510 gnd.n4939 gnd.n4938 0.0296328
R22511 gnd.n1023 gnd.n993 0.0296328
R22512 gnd.n3151 gnd.n3150 0.0269946
R22513 gnd.n3153 gnd.n3152 0.0269946
R22514 gnd.n2859 gnd.n2857 0.0269946
R22515 gnd.n3163 gnd.n3161 0.0269946
R22516 gnd.n3162 gnd.n2838 0.0269946
R22517 gnd.n3182 gnd.n3181 0.0269946
R22518 gnd.n3184 gnd.n3183 0.0269946
R22519 gnd.n2833 gnd.n2832 0.0269946
R22520 gnd.n3194 gnd.n2828 0.0269946
R22521 gnd.n3193 gnd.n2830 0.0269946
R22522 gnd.n2829 gnd.n2811 0.0269946
R22523 gnd.n3214 gnd.n2812 0.0269946
R22524 gnd.n3213 gnd.n2813 0.0269946
R22525 gnd.n3247 gnd.n2788 0.0269946
R22526 gnd.n3249 gnd.n3248 0.0269946
R22527 gnd.n3250 gnd.n2735 0.0269946
R22528 gnd.n2783 gnd.n2736 0.0269946
R22529 gnd.n2785 gnd.n2737 0.0269946
R22530 gnd.n3260 gnd.n3259 0.0269946
R22531 gnd.n3262 gnd.n3261 0.0269946
R22532 gnd.n3263 gnd.n2757 0.0269946
R22533 gnd.n3265 gnd.n2758 0.0269946
R22534 gnd.n3268 gnd.n2759 0.0269946
R22535 gnd.n3271 gnd.n3270 0.0269946
R22536 gnd.n3273 gnd.n3272 0.0269946
R22537 gnd.n3338 gnd.n2626 0.0269946
R22538 gnd.n3340 gnd.n3339 0.0269946
R22539 gnd.n3349 gnd.n2619 0.0269946
R22540 gnd.n3351 gnd.n3350 0.0269946
R22541 gnd.n3352 gnd.n2617 0.0269946
R22542 gnd.n3359 gnd.n3355 0.0269946
R22543 gnd.n3358 gnd.n3357 0.0269946
R22544 gnd.n3356 gnd.n2596 0.0269946
R22545 gnd.n3381 gnd.n2597 0.0269946
R22546 gnd.n3380 gnd.n2598 0.0269946
R22547 gnd.n3423 gnd.n2571 0.0269946
R22548 gnd.n3425 gnd.n3424 0.0269946
R22549 gnd.n3434 gnd.n2564 0.0269946
R22550 gnd.n3436 gnd.n3435 0.0269946
R22551 gnd.n3437 gnd.n2562 0.0269946
R22552 gnd.n3444 gnd.n3440 0.0269946
R22553 gnd.n3443 gnd.n3442 0.0269946
R22554 gnd.n3441 gnd.n2541 0.0269946
R22555 gnd.n3466 gnd.n2542 0.0269946
R22556 gnd.n3465 gnd.n2543 0.0269946
R22557 gnd.n3512 gnd.n2517 0.0269946
R22558 gnd.n3514 gnd.n3513 0.0269946
R22559 gnd.n3523 gnd.n2510 0.0269946
R22560 gnd.n3782 gnd.n2508 0.0269946
R22561 gnd.n3787 gnd.n3785 0.0269946
R22562 gnd.n3786 gnd.n2489 0.0269946
R22563 gnd.n3811 gnd.n3810 0.0269946
R22564 gnd.n4992 gnd.n2079 0.022519
R22565 gnd.n4989 gnd.n4988 0.022519
R22566 gnd.n4985 gnd.n2083 0.022519
R22567 gnd.n4984 gnd.n2092 0.022519
R22568 gnd.n4981 gnd.n4980 0.022519
R22569 gnd.n4977 gnd.n2099 0.022519
R22570 gnd.n4976 gnd.n2106 0.022519
R22571 gnd.n4973 gnd.n4972 0.022519
R22572 gnd.n4969 gnd.n2112 0.022519
R22573 gnd.n4968 gnd.n2118 0.022519
R22574 gnd.n4965 gnd.n4964 0.022519
R22575 gnd.n4961 gnd.n2125 0.022519
R22576 gnd.n4960 gnd.n2132 0.022519
R22577 gnd.n4957 gnd.n4956 0.022519
R22578 gnd.n4953 gnd.n2138 0.022519
R22579 gnd.n4952 gnd.n2144 0.022519
R22580 gnd.n4949 gnd.n4948 0.022519
R22581 gnd.n4945 gnd.n2153 0.022519
R22582 gnd.n4944 gnd.n4939 0.022519
R22583 gnd.n6093 gnd.n1147 0.022519
R22584 gnd.n6092 gnd.n1148 0.022519
R22585 gnd.n6089 gnd.n6088 0.022519
R22586 gnd.n6085 gnd.n6017 0.022519
R22587 gnd.n6084 gnd.n6021 0.022519
R22588 gnd.n6081 gnd.n6080 0.022519
R22589 gnd.n6077 gnd.n6027 0.022519
R22590 gnd.n6076 gnd.n6033 0.022519
R22591 gnd.n6073 gnd.n6072 0.022519
R22592 gnd.n6069 gnd.n6037 0.022519
R22593 gnd.n6068 gnd.n6041 0.022519
R22594 gnd.n6065 gnd.n6064 0.022519
R22595 gnd.n6061 gnd.n6047 0.022519
R22596 gnd.n6060 gnd.n6053 0.022519
R22597 gnd.n6057 gnd.n6056 0.022519
R22598 gnd.n6223 gnd.n1018 0.022519
R22599 gnd.n6222 gnd.n1019 0.022519
R22600 gnd.n1029 gnd.n1028 0.022519
R22601 gnd.n1024 gnd.n1023 0.022519
R22602 gnd.n6230 gnd.n993 0.0218415
R22603 gnd.n4938 gnd.n867 0.0218415
R22604 gnd.n3131 gnd.n3130 0.0202011
R22605 gnd.n3130 gnd.n3129 0.0148637
R22606 gnd.n3780 gnd.n3524 0.0144266
R22607 gnd.n3781 gnd.n3780 0.0130679
R22608 gnd.n4993 gnd.n4992 0.0123564
R22609 gnd.n4989 gnd.n2079 0.0123564
R22610 gnd.n4988 gnd.n2083 0.0123564
R22611 gnd.n4985 gnd.n4984 0.0123564
R22612 gnd.n4981 gnd.n2092 0.0123564
R22613 gnd.n4980 gnd.n2099 0.0123564
R22614 gnd.n4977 gnd.n4976 0.0123564
R22615 gnd.n4973 gnd.n2106 0.0123564
R22616 gnd.n4972 gnd.n2112 0.0123564
R22617 gnd.n4969 gnd.n4968 0.0123564
R22618 gnd.n4965 gnd.n2118 0.0123564
R22619 gnd.n4964 gnd.n2125 0.0123564
R22620 gnd.n4961 gnd.n4960 0.0123564
R22621 gnd.n4957 gnd.n2132 0.0123564
R22622 gnd.n4956 gnd.n2138 0.0123564
R22623 gnd.n4953 gnd.n4952 0.0123564
R22624 gnd.n4949 gnd.n2144 0.0123564
R22625 gnd.n4948 gnd.n2153 0.0123564
R22626 gnd.n4945 gnd.n4944 0.0123564
R22627 gnd.n1147 gnd.n1140 0.0123564
R22628 gnd.n6093 gnd.n6092 0.0123564
R22629 gnd.n6089 gnd.n1148 0.0123564
R22630 gnd.n6088 gnd.n6017 0.0123564
R22631 gnd.n6085 gnd.n6084 0.0123564
R22632 gnd.n6081 gnd.n6021 0.0123564
R22633 gnd.n6080 gnd.n6027 0.0123564
R22634 gnd.n6077 gnd.n6076 0.0123564
R22635 gnd.n6073 gnd.n6033 0.0123564
R22636 gnd.n6072 gnd.n6037 0.0123564
R22637 gnd.n6069 gnd.n6068 0.0123564
R22638 gnd.n6065 gnd.n6041 0.0123564
R22639 gnd.n6064 gnd.n6047 0.0123564
R22640 gnd.n6061 gnd.n6060 0.0123564
R22641 gnd.n6057 gnd.n6053 0.0123564
R22642 gnd.n6056 gnd.n1018 0.0123564
R22643 gnd.n6223 gnd.n6222 0.0123564
R22644 gnd.n1029 gnd.n1019 0.0123564
R22645 gnd.n1028 gnd.n1024 0.0123564
R22646 gnd.n3150 gnd.n2864 0.00797283
R22647 gnd.n3152 gnd.n3151 0.00797283
R22648 gnd.n3153 gnd.n2859 0.00797283
R22649 gnd.n3161 gnd.n2857 0.00797283
R22650 gnd.n3163 gnd.n3162 0.00797283
R22651 gnd.n3181 gnd.n2838 0.00797283
R22652 gnd.n3183 gnd.n3182 0.00797283
R22653 gnd.n3184 gnd.n2833 0.00797283
R22654 gnd.n2832 gnd.n2828 0.00797283
R22655 gnd.n3194 gnd.n3193 0.00797283
R22656 gnd.n2830 gnd.n2829 0.00797283
R22657 gnd.n2812 gnd.n2811 0.00797283
R22658 gnd.n3214 gnd.n3213 0.00797283
R22659 gnd.n2813 gnd.n2788 0.00797283
R22660 gnd.n3248 gnd.n3247 0.00797283
R22661 gnd.n3250 gnd.n3249 0.00797283
R22662 gnd.n2783 gnd.n2735 0.00797283
R22663 gnd.n2785 gnd.n2736 0.00797283
R22664 gnd.n3259 gnd.n2737 0.00797283
R22665 gnd.n3261 gnd.n3260 0.00797283
R22666 gnd.n3263 gnd.n3262 0.00797283
R22667 gnd.n3265 gnd.n2757 0.00797283
R22668 gnd.n3268 gnd.n2758 0.00797283
R22669 gnd.n3270 gnd.n2759 0.00797283
R22670 gnd.n3273 gnd.n3271 0.00797283
R22671 gnd.n3272 gnd.n2626 0.00797283
R22672 gnd.n3340 gnd.n3338 0.00797283
R22673 gnd.n3339 gnd.n2619 0.00797283
R22674 gnd.n3350 gnd.n3349 0.00797283
R22675 gnd.n3352 gnd.n3351 0.00797283
R22676 gnd.n3355 gnd.n2617 0.00797283
R22677 gnd.n3359 gnd.n3358 0.00797283
R22678 gnd.n3357 gnd.n3356 0.00797283
R22679 gnd.n2597 gnd.n2596 0.00797283
R22680 gnd.n3381 gnd.n3380 0.00797283
R22681 gnd.n2598 gnd.n2571 0.00797283
R22682 gnd.n3425 gnd.n3423 0.00797283
R22683 gnd.n3424 gnd.n2564 0.00797283
R22684 gnd.n3435 gnd.n3434 0.00797283
R22685 gnd.n3437 gnd.n3436 0.00797283
R22686 gnd.n3440 gnd.n2562 0.00797283
R22687 gnd.n3444 gnd.n3443 0.00797283
R22688 gnd.n3442 gnd.n3441 0.00797283
R22689 gnd.n2542 gnd.n2541 0.00797283
R22690 gnd.n3466 gnd.n3465 0.00797283
R22691 gnd.n2543 gnd.n2517 0.00797283
R22692 gnd.n3514 gnd.n3512 0.00797283
R22693 gnd.n3513 gnd.n2510 0.00797283
R22694 gnd.n3524 gnd.n3523 0.00797283
R22695 gnd.n3782 gnd.n3781 0.00797283
R22696 gnd.n3785 gnd.n2508 0.00797283
R22697 gnd.n3787 gnd.n3786 0.00797283
R22698 gnd.n3810 gnd.n2489 0.00797283
R22699 gnd.n3811 gnd.n2453 0.00797283
R22700 gnd.n4994 gnd.n836 0.00592005
R22701 gnd.n6098 gnd.n6097 0.00592005
R22702 gnd.n7187 gnd.n272 0.00417647
R22703 gnd.n7216 gnd.n272 0.00417647
R22704 gnd.n7217 gnd.n7216 0.00417647
R22705 gnd.n7218 gnd.n7217 0.00417647
R22706 gnd.n7220 gnd.n7218 0.00417647
R22707 gnd.n7220 gnd.n7219 0.00417647
R22708 gnd.n7219 gnd.n111 0.00417647
R22709 gnd.n112 gnd.n111 0.00417647
R22710 gnd.n113 gnd.n112 0.00417647
R22711 gnd.n130 gnd.n113 0.00417647
R22712 gnd.n4392 gnd.n2276 0.00417647
R22713 gnd.n4424 gnd.n2276 0.00417647
R22714 gnd.n4425 gnd.n4424 0.00417647
R22715 gnd.n4426 gnd.n4425 0.00417647
R22716 gnd.n4427 gnd.n4426 0.00417647
R22717 gnd.n4427 gnd.n2250 0.00417647
R22718 gnd.n4458 gnd.n2250 0.00417647
R22719 gnd.n4459 gnd.n4458 0.00417647
R22720 gnd.n4460 gnd.n4459 0.00417647
R22721 gnd.n4461 gnd.n4460 0.00417647
R22722 plus.n53 plus.t20 323.478
R22723 plus.n11 plus.t15 323.478
R22724 plus.n52 plus.t19 297.12
R22725 plus.n56 plus.t26 297.12
R22726 plus.n58 plus.t25 297.12
R22727 plus.n62 plus.t27 297.12
R22728 plus.n64 plus.t9 297.12
R22729 plus.n68 plus.t7 297.12
R22730 plus.n70 plus.t14 297.12
R22731 plus.n74 plus.t12 297.12
R22732 plus.n76 plus.t28 297.12
R22733 plus.n80 plus.t10 297.12
R22734 plus.n82 plus.t8 297.12
R22735 plus.n40 plus.t21 297.12
R22736 plus.n38 plus.t22 297.12
R22737 plus.n2 plus.t16 297.12
R22738 plus.n32 plus.t17 297.12
R22739 plus.n4 plus.t11 297.12
R22740 plus.n26 plus.t5 297.12
R22741 plus.n6 plus.t6 297.12
R22742 plus.n20 plus.t23 297.12
R22743 plus.n8 plus.t24 297.12
R22744 plus.n14 plus.t18 297.12
R22745 plus.n10 plus.t13 297.12
R22746 plus.n86 plus.t2 243.97
R22747 plus.n86 plus.n85 223.454
R22748 plus.n88 plus.n87 223.454
R22749 plus.n83 plus.n82 161.3
R22750 plus.n81 plus.n42 161.3
R22751 plus.n80 plus.n79 161.3
R22752 plus.n78 plus.n43 161.3
R22753 plus.n77 plus.n76 161.3
R22754 plus.n75 plus.n44 161.3
R22755 plus.n74 plus.n73 161.3
R22756 plus.n72 plus.n45 161.3
R22757 plus.n71 plus.n70 161.3
R22758 plus.n69 plus.n46 161.3
R22759 plus.n68 plus.n67 161.3
R22760 plus.n66 plus.n47 161.3
R22761 plus.n65 plus.n64 161.3
R22762 plus.n63 plus.n48 161.3
R22763 plus.n62 plus.n61 161.3
R22764 plus.n60 plus.n49 161.3
R22765 plus.n59 plus.n58 161.3
R22766 plus.n57 plus.n50 161.3
R22767 plus.n56 plus.n55 161.3
R22768 plus.n54 plus.n51 161.3
R22769 plus.n13 plus.n12 161.3
R22770 plus.n14 plus.n9 161.3
R22771 plus.n16 plus.n15 161.3
R22772 plus.n17 plus.n8 161.3
R22773 plus.n19 plus.n18 161.3
R22774 plus.n20 plus.n7 161.3
R22775 plus.n22 plus.n21 161.3
R22776 plus.n23 plus.n6 161.3
R22777 plus.n25 plus.n24 161.3
R22778 plus.n26 plus.n5 161.3
R22779 plus.n28 plus.n27 161.3
R22780 plus.n29 plus.n4 161.3
R22781 plus.n31 plus.n30 161.3
R22782 plus.n32 plus.n3 161.3
R22783 plus.n34 plus.n33 161.3
R22784 plus.n35 plus.n2 161.3
R22785 plus.n37 plus.n36 161.3
R22786 plus.n38 plus.n1 161.3
R22787 plus.n39 plus.n0 161.3
R22788 plus.n41 plus.n40 161.3
R22789 plus.n82 plus.n81 46.0096
R22790 plus.n40 plus.n39 46.0096
R22791 plus.n54 plus.n53 45.0871
R22792 plus.n12 plus.n11 45.0871
R22793 plus.n52 plus.n51 41.6278
R22794 plus.n80 plus.n43 41.6278
R22795 plus.n38 plus.n37 41.6278
R22796 plus.n13 plus.n10 41.6278
R22797 plus.n57 plus.n56 37.246
R22798 plus.n76 plus.n75 37.246
R22799 plus.n33 plus.n2 37.246
R22800 plus.n15 plus.n14 37.246
R22801 plus.n84 plus.n83 33.1766
R22802 plus.n58 plus.n49 32.8641
R22803 plus.n74 plus.n45 32.8641
R22804 plus.n32 plus.n31 32.8641
R22805 plus.n19 plus.n8 32.8641
R22806 plus.n63 plus.n62 28.4823
R22807 plus.n70 plus.n69 28.4823
R22808 plus.n27 plus.n4 28.4823
R22809 plus.n21 plus.n20 28.4823
R22810 plus.n64 plus.n47 24.1005
R22811 plus.n68 plus.n47 24.1005
R22812 plus.n26 plus.n25 24.1005
R22813 plus.n25 plus.n6 24.1005
R22814 plus.n85 plus.t3 19.8005
R22815 plus.n85 plus.t1 19.8005
R22816 plus.n87 plus.t4 19.8005
R22817 plus.n87 plus.t0 19.8005
R22818 plus.n64 plus.n63 19.7187
R22819 plus.n69 plus.n68 19.7187
R22820 plus.n27 plus.n26 19.7187
R22821 plus.n21 plus.n6 19.7187
R22822 plus.n62 plus.n49 15.3369
R22823 plus.n70 plus.n45 15.3369
R22824 plus.n31 plus.n4 15.3369
R22825 plus.n20 plus.n19 15.3369
R22826 plus plus.n89 15.1953
R22827 plus.n53 plus.n52 14.1472
R22828 plus.n11 plus.n10 14.1472
R22829 plus.n84 plus.n41 11.8774
R22830 plus.n58 plus.n57 10.955
R22831 plus.n75 plus.n74 10.955
R22832 plus.n33 plus.n32 10.955
R22833 plus.n15 plus.n8 10.955
R22834 plus.n56 plus.n51 6.57323
R22835 plus.n76 plus.n43 6.57323
R22836 plus.n37 plus.n2 6.57323
R22837 plus.n14 plus.n13 6.57323
R22838 plus.n89 plus.n88 5.40567
R22839 plus.n81 plus.n80 2.19141
R22840 plus.n39 plus.n38 2.19141
R22841 plus.n89 plus.n84 1.188
R22842 plus.n88 plus.n86 0.716017
R22843 plus.n55 plus.n54 0.189894
R22844 plus.n55 plus.n50 0.189894
R22845 plus.n59 plus.n50 0.189894
R22846 plus.n60 plus.n59 0.189894
R22847 plus.n61 plus.n60 0.189894
R22848 plus.n61 plus.n48 0.189894
R22849 plus.n65 plus.n48 0.189894
R22850 plus.n66 plus.n65 0.189894
R22851 plus.n67 plus.n66 0.189894
R22852 plus.n67 plus.n46 0.189894
R22853 plus.n71 plus.n46 0.189894
R22854 plus.n72 plus.n71 0.189894
R22855 plus.n73 plus.n72 0.189894
R22856 plus.n73 plus.n44 0.189894
R22857 plus.n77 plus.n44 0.189894
R22858 plus.n78 plus.n77 0.189894
R22859 plus.n79 plus.n78 0.189894
R22860 plus.n79 plus.n42 0.189894
R22861 plus.n83 plus.n42 0.189894
R22862 plus.n41 plus.n0 0.189894
R22863 plus.n1 plus.n0 0.189894
R22864 plus.n36 plus.n1 0.189894
R22865 plus.n36 plus.n35 0.189894
R22866 plus.n35 plus.n34 0.189894
R22867 plus.n34 plus.n3 0.189894
R22868 plus.n30 plus.n3 0.189894
R22869 plus.n30 plus.n29 0.189894
R22870 plus.n29 plus.n28 0.189894
R22871 plus.n28 plus.n5 0.189894
R22872 plus.n24 plus.n5 0.189894
R22873 plus.n24 plus.n23 0.189894
R22874 plus.n23 plus.n22 0.189894
R22875 plus.n22 plus.n7 0.189894
R22876 plus.n18 plus.n7 0.189894
R22877 plus.n18 plus.n17 0.189894
R22878 plus.n17 plus.n16 0.189894
R22879 plus.n16 plus.n9 0.189894
R22880 plus.n12 plus.n9 0.189894
R22881 a_n3827_n3924.n30 a_n3827_n3924.t55 214.994
R22882 a_n3827_n3924.n39 a_n3827_n3924.t22 214.786
R22883 a_n3827_n3924.n38 a_n3827_n3924.t23 214.321
R22884 a_n3827_n3924.n37 a_n3827_n3924.t53 214.321
R22885 a_n3827_n3924.n36 a_n3827_n3924.t17 214.321
R22886 a_n3827_n3924.n35 a_n3827_n3924.t57 214.321
R22887 a_n3827_n3924.n34 a_n3827_n3924.t52 214.321
R22888 a_n3827_n3924.n33 a_n3827_n3924.t11 214.321
R22889 a_n3827_n3924.n32 a_n3827_n3924.t54 214.321
R22890 a_n3827_n3924.n30 a_n3827_n3924.t14 214.321
R22891 a_n3827_n3924.n13 a_n3827_n3924.t36 55.8337
R22892 a_n3827_n3924.n14 a_n3827_n3924.t18 55.8337
R22893 a_n3827_n3924.n25 a_n3827_n3924.t8 55.8337
R22894 a_n3827_n3924.n2 a_n3827_n3924.t48 55.8335
R22895 a_n3827_n3924.n41 a_n3827_n3924.t21 55.8335
R22896 a_n3827_n3924.n52 a_n3827_n3924.t2 55.8335
R22897 a_n3827_n3924.n53 a_n3827_n3924.t41 55.8335
R22898 a_n3827_n3924.n28 a_n3827_n3924.t35 55.8335
R22899 a_n3827_n3924.n59 a_n3827_n3924.n58 53.0054
R22900 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R22901 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R22902 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R22903 a_n3827_n3924.n10 a_n3827_n3924.n9 53.0052
R22904 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R22905 a_n3827_n3924.n16 a_n3827_n3924.n15 53.0052
R22906 a_n3827_n3924.n18 a_n3827_n3924.n17 53.0052
R22907 a_n3827_n3924.n20 a_n3827_n3924.n19 53.0052
R22908 a_n3827_n3924.n22 a_n3827_n3924.n21 53.0052
R22909 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0052
R22910 a_n3827_n3924.n43 a_n3827_n3924.n42 53.0051
R22911 a_n3827_n3924.n45 a_n3827_n3924.n44 53.0051
R22912 a_n3827_n3924.n47 a_n3827_n3924.n46 53.0051
R22913 a_n3827_n3924.n49 a_n3827_n3924.n48 53.0051
R22914 a_n3827_n3924.n51 a_n3827_n3924.n50 53.0051
R22915 a_n3827_n3924.n55 a_n3827_n3924.n54 53.0051
R22916 a_n3827_n3924.n57 a_n3827_n3924.n56 53.0051
R22917 a_n3827_n3924.n1 a_n3827_n3924.n0 53.0051
R22918 a_n3827_n3924.n27 a_n3827_n3924.n26 53.0051
R22919 a_n3827_n3924.n29 a_n3827_n3924.n25 12.1986
R22920 a_n3827_n3924.n40 a_n3827_n3924.n2 12.1986
R22921 a_n3827_n3924.n29 a_n3827_n3924.n28 5.11903
R22922 a_n3827_n3924.n41 a_n3827_n3924.n40 5.11903
R22923 a_n3827_n3924.n42 a_n3827_n3924.t3 2.82907
R22924 a_n3827_n3924.n42 a_n3827_n3924.t6 2.82907
R22925 a_n3827_n3924.n44 a_n3827_n3924.t19 2.82907
R22926 a_n3827_n3924.n44 a_n3827_n3924.t0 2.82907
R22927 a_n3827_n3924.n46 a_n3827_n3924.t20 2.82907
R22928 a_n3827_n3924.n46 a_n3827_n3924.t56 2.82907
R22929 a_n3827_n3924.n48 a_n3827_n3924.t26 2.82907
R22930 a_n3827_n3924.n48 a_n3827_n3924.t4 2.82907
R22931 a_n3827_n3924.n50 a_n3827_n3924.t7 2.82907
R22932 a_n3827_n3924.n50 a_n3827_n3924.t25 2.82907
R22933 a_n3827_n3924.n54 a_n3827_n3924.t38 2.82907
R22934 a_n3827_n3924.n54 a_n3827_n3924.t43 2.82907
R22935 a_n3827_n3924.n56 a_n3827_n3924.t33 2.82907
R22936 a_n3827_n3924.n56 a_n3827_n3924.t32 2.82907
R22937 a_n3827_n3924.n0 a_n3827_n3924.t39 2.82907
R22938 a_n3827_n3924.n0 a_n3827_n3924.t45 2.82907
R22939 a_n3827_n3924.n26 a_n3827_n3924.t34 2.82907
R22940 a_n3827_n3924.n26 a_n3827_n3924.t40 2.82907
R22941 a_n3827_n3924.n3 a_n3827_n3924.t28 2.82907
R22942 a_n3827_n3924.n3 a_n3827_n3924.t46 2.82907
R22943 a_n3827_n3924.n5 a_n3827_n3924.t42 2.82907
R22944 a_n3827_n3924.n5 a_n3827_n3924.t44 2.82907
R22945 a_n3827_n3924.n7 a_n3827_n3924.t47 2.82907
R22946 a_n3827_n3924.n7 a_n3827_n3924.t49 2.82907
R22947 a_n3827_n3924.n9 a_n3827_n3924.t31 2.82907
R22948 a_n3827_n3924.n9 a_n3827_n3924.t29 2.82907
R22949 a_n3827_n3924.n11 a_n3827_n3924.t37 2.82907
R22950 a_n3827_n3924.n11 a_n3827_n3924.t30 2.82907
R22951 a_n3827_n3924.n15 a_n3827_n3924.t12 2.82907
R22952 a_n3827_n3924.n15 a_n3827_n3924.t15 2.82907
R22953 a_n3827_n3924.n17 a_n3827_n3924.t1 2.82907
R22954 a_n3827_n3924.n17 a_n3827_n3924.t27 2.82907
R22955 a_n3827_n3924.n19 a_n3827_n3924.t16 2.82907
R22956 a_n3827_n3924.n19 a_n3827_n3924.t5 2.82907
R22957 a_n3827_n3924.n21 a_n3827_n3924.t13 2.82907
R22958 a_n3827_n3924.n21 a_n3827_n3924.t9 2.82907
R22959 a_n3827_n3924.n23 a_n3827_n3924.t24 2.82907
R22960 a_n3827_n3924.n23 a_n3827_n3924.t10 2.82907
R22961 a_n3827_n3924.t51 a_n3827_n3924.n59 2.82907
R22962 a_n3827_n3924.n59 a_n3827_n3924.t50 2.82907
R22963 a_n3827_n3924.n31 a_n3827_n3924.n29 1.95694
R22964 a_n3827_n3924.n40 a_n3827_n3924.n39 1.95694
R22965 a_n3827_n3924.n33 a_n3827_n3924.n32 0.672012
R22966 a_n3827_n3924.n34 a_n3827_n3924.n33 0.672012
R22967 a_n3827_n3924.n35 a_n3827_n3924.n34 0.672012
R22968 a_n3827_n3924.n36 a_n3827_n3924.n35 0.672012
R22969 a_n3827_n3924.n37 a_n3827_n3924.n36 0.672012
R22970 a_n3827_n3924.n38 a_n3827_n3924.n37 0.672012
R22971 a_n3827_n3924.n25 a_n3827_n3924.n24 0.444466
R22972 a_n3827_n3924.n24 a_n3827_n3924.n22 0.444466
R22973 a_n3827_n3924.n22 a_n3827_n3924.n20 0.444466
R22974 a_n3827_n3924.n20 a_n3827_n3924.n18 0.444466
R22975 a_n3827_n3924.n18 a_n3827_n3924.n16 0.444466
R22976 a_n3827_n3924.n16 a_n3827_n3924.n14 0.444466
R22977 a_n3827_n3924.n13 a_n3827_n3924.n12 0.444466
R22978 a_n3827_n3924.n12 a_n3827_n3924.n10 0.444466
R22979 a_n3827_n3924.n10 a_n3827_n3924.n8 0.444466
R22980 a_n3827_n3924.n8 a_n3827_n3924.n6 0.444466
R22981 a_n3827_n3924.n6 a_n3827_n3924.n4 0.444466
R22982 a_n3827_n3924.n4 a_n3827_n3924.n2 0.444466
R22983 a_n3827_n3924.n28 a_n3827_n3924.n27 0.444466
R22984 a_n3827_n3924.n27 a_n3827_n3924.n1 0.444466
R22985 a_n3827_n3924.n58 a_n3827_n3924.n1 0.444466
R22986 a_n3827_n3924.n58 a_n3827_n3924.n57 0.444466
R22987 a_n3827_n3924.n57 a_n3827_n3924.n55 0.444466
R22988 a_n3827_n3924.n55 a_n3827_n3924.n53 0.444466
R22989 a_n3827_n3924.n52 a_n3827_n3924.n51 0.444466
R22990 a_n3827_n3924.n51 a_n3827_n3924.n49 0.444466
R22991 a_n3827_n3924.n49 a_n3827_n3924.n47 0.444466
R22992 a_n3827_n3924.n47 a_n3827_n3924.n45 0.444466
R22993 a_n3827_n3924.n45 a_n3827_n3924.n43 0.444466
R22994 a_n3827_n3924.n43 a_n3827_n3924.n41 0.444466
R22995 a_n3827_n3924.n32 a_n3827_n3924.n31 0.350064
R22996 a_n3827_n3924.n31 a_n3827_n3924.n30 0.322448
R22997 a_n3827_n3924.n14 a_n3827_n3924.n13 0.235414
R22998 a_n3827_n3924.n53 a_n3827_n3924.n52 0.235414
R22999 a_n3827_n3924.n39 a_n3827_n3924.n38 0.207622
R23000 a_n2408_n452.n81 a_n2408_n452.t63 512.366
R23001 a_n2408_n452.n80 a_n2408_n452.t54 512.366
R23002 a_n2408_n452.n79 a_n2408_n452.t48 512.366
R23003 a_n2408_n452.n83 a_n2408_n452.t71 512.366
R23004 a_n2408_n452.n82 a_n2408_n452.t60 512.366
R23005 a_n2408_n452.n78 a_n2408_n452.t59 512.366
R23006 a_n2408_n452.n85 a_n2408_n452.t67 512.366
R23007 a_n2408_n452.n84 a_n2408_n452.t52 512.366
R23008 a_n2408_n452.n77 a_n2408_n452.t53 512.366
R23009 a_n2408_n452.n87 a_n2408_n452.t55 512.366
R23010 a_n2408_n452.n86 a_n2408_n452.t65 512.366
R23011 a_n2408_n452.n76 a_n2408_n452.t75 512.366
R23012 a_n2408_n452.n26 a_n2408_n452.t74 539.01
R23013 a_n2408_n452.n56 a_n2408_n452.t57 512.366
R23014 a_n2408_n452.n55 a_n2408_n452.t61 512.366
R23015 a_n2408_n452.n53 a_n2408_n452.t51 512.366
R23016 a_n2408_n452.n54 a_n2408_n452.t66 512.366
R23017 a_n2408_n452.n22 a_n2408_n452.t33 539.01
R23018 a_n2408_n452.n71 a_n2408_n452.t35 512.366
R23019 a_n2408_n452.n70 a_n2408_n452.t41 512.366
R23020 a_n2408_n452.n50 a_n2408_n452.t23 512.366
R23021 a_n2408_n452.n57 a_n2408_n452.t39 512.366
R23022 a_n2408_n452.n16 a_n2408_n452.t25 539.01
R23023 a_n2408_n452.n92 a_n2408_n452.t21 512.366
R23024 a_n2408_n452.n93 a_n2408_n452.t19 512.366
R23025 a_n2408_n452.n51 a_n2408_n452.t37 512.366
R23026 a_n2408_n452.n94 a_n2408_n452.t29 512.366
R23027 a_n2408_n452.n20 a_n2408_n452.t69 539.01
R23028 a_n2408_n452.n89 a_n2408_n452.t70 512.366
R23029 a_n2408_n452.n90 a_n2408_n452.t49 512.366
R23030 a_n2408_n452.n52 a_n2408_n452.t56 512.366
R23031 a_n2408_n452.n91 a_n2408_n452.t64 512.366
R23032 a_n2408_n452.n5 a_n2408_n452.n49 70.1674
R23033 a_n2408_n452.n7 a_n2408_n452.n47 70.1674
R23034 a_n2408_n452.n9 a_n2408_n452.n45 70.1674
R23035 a_n2408_n452.n11 a_n2408_n452.n43 70.1674
R23036 a_n2408_n452.n34 a_n2408_n452.n24 70.3058
R23037 a_n2408_n452.n28 a_n2408_n452.n27 44.8194
R23038 a_n2408_n452.n28 a_n2408_n452.n57 13.6566
R23039 a_n2408_n452.n25 a_n2408_n452.n32 70.1674
R23040 a_n2408_n452.n32 a_n2408_n452.n53 20.9683
R23041 a_n2408_n452.n31 a_n2408_n452.n25 75.0448
R23042 a_n2408_n452.n55 a_n2408_n452.n31 11.2134
R23043 a_n2408_n452.n23 a_n2408_n452.n26 44.8194
R23044 a_n2408_n452.n35 a_n2408_n452.n27 44.5595
R23045 a_n2408_n452.n70 a_n2408_n452.n35 20.9685
R23046 a_n2408_n452.n21 a_n2408_n452.n22 44.8194
R23047 a_n2408_n452.n13 a_n2408_n452.n41 70.3058
R23048 a_n2408_n452.n17 a_n2408_n452.n38 70.3058
R23049 a_n2408_n452.n37 a_n2408_n452.n18 70.1674
R23050 a_n2408_n452.n37 a_n2408_n452.n52 20.9683
R23051 a_n2408_n452.n18 a_n2408_n452.n36 75.0448
R23052 a_n2408_n452.n90 a_n2408_n452.n36 11.2134
R23053 a_n2408_n452.n19 a_n2408_n452.n20 44.8194
R23054 a_n2408_n452.n40 a_n2408_n452.n14 70.1674
R23055 a_n2408_n452.n40 a_n2408_n452.n51 20.9683
R23056 a_n2408_n452.n14 a_n2408_n452.n39 75.0448
R23057 a_n2408_n452.n93 a_n2408_n452.n39 11.2134
R23058 a_n2408_n452.n15 a_n2408_n452.n16 44.8194
R23059 a_n2408_n452.n43 a_n2408_n452.n76 20.9683
R23060 a_n2408_n452.n42 a_n2408_n452.n12 75.0448
R23061 a_n2408_n452.n86 a_n2408_n452.n42 11.2134
R23062 a_n2408_n452.n12 a_n2408_n452.n87 161.3
R23063 a_n2408_n452.n45 a_n2408_n452.n77 20.9683
R23064 a_n2408_n452.n44 a_n2408_n452.n10 75.0448
R23065 a_n2408_n452.n84 a_n2408_n452.n44 11.2134
R23066 a_n2408_n452.n10 a_n2408_n452.n85 161.3
R23067 a_n2408_n452.n47 a_n2408_n452.n78 20.9683
R23068 a_n2408_n452.n46 a_n2408_n452.n8 75.0448
R23069 a_n2408_n452.n82 a_n2408_n452.n46 11.2134
R23070 a_n2408_n452.n8 a_n2408_n452.n83 161.3
R23071 a_n2408_n452.n49 a_n2408_n452.n79 20.9683
R23072 a_n2408_n452.n48 a_n2408_n452.n6 75.0448
R23073 a_n2408_n452.n80 a_n2408_n452.n48 11.2134
R23074 a_n2408_n452.n6 a_n2408_n452.n81 161.3
R23075 a_n2408_n452.n3 a_n2408_n452.n67 81.3764
R23076 a_n2408_n452.n4 a_n2408_n452.n61 81.3764
R23077 a_n2408_n452.n0 a_n2408_n452.n58 81.3764
R23078 a_n2408_n452.n3 a_n2408_n452.n68 80.9324
R23079 a_n2408_n452.n2 a_n2408_n452.n69 80.9324
R23080 a_n2408_n452.n2 a_n2408_n452.n66 80.9324
R23081 a_n2408_n452.n2 a_n2408_n452.n65 80.9324
R23082 a_n2408_n452.n1 a_n2408_n452.n64 80.9324
R23083 a_n2408_n452.n4 a_n2408_n452.n62 80.9324
R23084 a_n2408_n452.n0 a_n2408_n452.n63 80.9324
R23085 a_n2408_n452.n0 a_n2408_n452.n60 80.9324
R23086 a_n2408_n452.n0 a_n2408_n452.n59 80.9324
R23087 a_n2408_n452.n97 a_n2408_n452.t26 74.6477
R23088 a_n2408_n452.n29 a_n2408_n452.t28 74.6477
R23089 a_n2408_n452.n74 a_n2408_n452.t34 74.2899
R23090 a_n2408_n452.n30 a_n2408_n452.t32 74.2897
R23091 a_n2408_n452.n30 a_n2408_n452.n96 70.6783
R23092 a_n2408_n452.n29 a_n2408_n452.n72 70.6783
R23093 a_n2408_n452.n29 a_n2408_n452.n73 70.6783
R23094 a_n2408_n452.n98 a_n2408_n452.n97 70.6782
R23095 a_n2408_n452.n81 a_n2408_n452.n80 48.2005
R23096 a_n2408_n452.t68 a_n2408_n452.n49 533.335
R23097 a_n2408_n452.n83 a_n2408_n452.n82 48.2005
R23098 a_n2408_n452.t73 a_n2408_n452.n47 533.335
R23099 a_n2408_n452.n85 a_n2408_n452.n84 48.2005
R23100 a_n2408_n452.t62 a_n2408_n452.n45 533.335
R23101 a_n2408_n452.n87 a_n2408_n452.n86 48.2005
R23102 a_n2408_n452.t58 a_n2408_n452.n43 533.335
R23103 a_n2408_n452.n56 a_n2408_n452.n55 48.2005
R23104 a_n2408_n452.n54 a_n2408_n452.n32 20.9683
R23105 a_n2408_n452.n71 a_n2408_n452.n70 48.2005
R23106 a_n2408_n452.n57 a_n2408_n452.n50 48.2005
R23107 a_n2408_n452.n93 a_n2408_n452.n92 48.2005
R23108 a_n2408_n452.n94 a_n2408_n452.n40 20.9683
R23109 a_n2408_n452.n90 a_n2408_n452.n89 48.2005
R23110 a_n2408_n452.n91 a_n2408_n452.n37 20.9683
R23111 a_n2408_n452.n34 a_n2408_n452.t72 533.058
R23112 a_n2408_n452.n28 a_n2408_n452.t27 539.01
R23113 a_n2408_n452.t31 a_n2408_n452.n41 533.058
R23114 a_n2408_n452.t50 a_n2408_n452.n38 533.058
R23115 a_n2408_n452.n1 a_n2408_n452.n0 32.6799
R23116 a_n2408_n452.n48 a_n2408_n452.n79 35.3134
R23117 a_n2408_n452.n46 a_n2408_n452.n78 35.3134
R23118 a_n2408_n452.n44 a_n2408_n452.n77 35.3134
R23119 a_n2408_n452.n42 a_n2408_n452.n76 35.3134
R23120 a_n2408_n452.n31 a_n2408_n452.n53 35.3134
R23121 a_n2408_n452.n35 a_n2408_n452.n50 20.9689
R23122 a_n2408_n452.n51 a_n2408_n452.n39 35.3134
R23123 a_n2408_n452.n52 a_n2408_n452.n36 35.3134
R23124 a_n2408_n452.n27 a_n2408_n452.n2 23.891
R23125 a_n2408_n452.n19 a_n2408_n452.n88 12.046
R23126 a_n2408_n452.n24 a_n2408_n452.n33 11.8414
R23127 a_n2408_n452.n75 a_n2408_n452.n21 10.5365
R23128 a_n2408_n452.n30 a_n2408_n452.n95 9.50122
R23129 a_n2408_n452.n88 a_n2408_n452.n12 7.47588
R23130 a_n2408_n452.n5 a_n2408_n452.n33 7.47588
R23131 a_n2408_n452.n95 a_n2408_n452.n13 6.70126
R23132 a_n2408_n452.n75 a_n2408_n452.n74 5.65783
R23133 a_n2408_n452.n95 a_n2408_n452.n33 5.3452
R23134 a_n2408_n452.n27 a_n2408_n452.n23 3.95126
R23135 a_n2408_n452.n15 a_n2408_n452.n17 3.95126
R23136 a_n2408_n452.n96 a_n2408_n452.t38 3.61217
R23137 a_n2408_n452.n96 a_n2408_n452.t30 3.61217
R23138 a_n2408_n452.n72 a_n2408_n452.t24 3.61217
R23139 a_n2408_n452.n72 a_n2408_n452.t40 3.61217
R23140 a_n2408_n452.n73 a_n2408_n452.t36 3.61217
R23141 a_n2408_n452.n73 a_n2408_n452.t42 3.61217
R23142 a_n2408_n452.n98 a_n2408_n452.t22 3.61217
R23143 a_n2408_n452.t20 a_n2408_n452.n98 3.61217
R23144 a_n2408_n452.n67 a_n2408_n452.t13 2.82907
R23145 a_n2408_n452.n67 a_n2408_n452.t15 2.82907
R23146 a_n2408_n452.n68 a_n2408_n452.t46 2.82907
R23147 a_n2408_n452.n68 a_n2408_n452.t11 2.82907
R23148 a_n2408_n452.n69 a_n2408_n452.t5 2.82907
R23149 a_n2408_n452.n69 a_n2408_n452.t1 2.82907
R23150 a_n2408_n452.n66 a_n2408_n452.t9 2.82907
R23151 a_n2408_n452.n66 a_n2408_n452.t14 2.82907
R23152 a_n2408_n452.n65 a_n2408_n452.t10 2.82907
R23153 a_n2408_n452.n65 a_n2408_n452.t12 2.82907
R23154 a_n2408_n452.n64 a_n2408_n452.t8 2.82907
R23155 a_n2408_n452.n64 a_n2408_n452.t43 2.82907
R23156 a_n2408_n452.n61 a_n2408_n452.t6 2.82907
R23157 a_n2408_n452.n61 a_n2408_n452.t18 2.82907
R23158 a_n2408_n452.n62 a_n2408_n452.t0 2.82907
R23159 a_n2408_n452.n62 a_n2408_n452.t3 2.82907
R23160 a_n2408_n452.n63 a_n2408_n452.t47 2.82907
R23161 a_n2408_n452.n63 a_n2408_n452.t16 2.82907
R23162 a_n2408_n452.n60 a_n2408_n452.t4 2.82907
R23163 a_n2408_n452.n60 a_n2408_n452.t17 2.82907
R23164 a_n2408_n452.n59 a_n2408_n452.t44 2.82907
R23165 a_n2408_n452.n59 a_n2408_n452.t45 2.82907
R23166 a_n2408_n452.n58 a_n2408_n452.t2 2.82907
R23167 a_n2408_n452.n58 a_n2408_n452.t7 2.82907
R23168 a_n2408_n452.n88 a_n2408_n452.n75 1.30542
R23169 a_n2408_n452.n9 a_n2408_n452.n8 1.04595
R23170 a_n2408_n452.n26 a_n2408_n452.n56 13.657
R23171 a_n2408_n452.n54 a_n2408_n452.n34 21.4216
R23172 a_n2408_n452.n22 a_n2408_n452.n71 13.657
R23173 a_n2408_n452.n92 a_n2408_n452.n16 13.657
R23174 a_n2408_n452.n41 a_n2408_n452.n94 21.4216
R23175 a_n2408_n452.n89 a_n2408_n452.n20 13.657
R23176 a_n2408_n452.n38 a_n2408_n452.n91 21.4216
R23177 a_n2408_n452.n27 a_n2408_n452.n21 1.47777
R23178 a_n2408_n452.n0 a_n2408_n452.n4 1.3324
R23179 a_n2408_n452.n2 a_n2408_n452.n3 0.888431
R23180 a_n2408_n452.n2 a_n2408_n452.n1 0.888431
R23181 a_n2408_n452.n25 a_n2408_n452.n23 0.758076
R23182 a_n2408_n452.n25 a_n2408_n452.n24 0.758076
R23183 a_n2408_n452.n19 a_n2408_n452.n18 0.758076
R23184 a_n2408_n452.n18 a_n2408_n452.n17 0.758076
R23185 a_n2408_n452.n15 a_n2408_n452.n14 0.758076
R23186 a_n2408_n452.n14 a_n2408_n452.n13 0.758076
R23187 a_n2408_n452.n12 a_n2408_n452.n11 0.758076
R23188 a_n2408_n452.n10 a_n2408_n452.n9 0.758076
R23189 a_n2408_n452.n8 a_n2408_n452.n7 0.758076
R23190 a_n2408_n452.n6 a_n2408_n452.n5 0.758076
R23191 a_n2408_n452.n97 a_n2408_n452.n30 0.716017
R23192 a_n2408_n452.n74 a_n2408_n452.n29 0.716017
R23193 a_n2408_n452.n11 a_n2408_n452.n10 0.67853
R23194 a_n2408_n452.n7 a_n2408_n452.n6 0.67853
R23195 a_n1808_13878.n2 a_n1808_13878.n0 98.9633
R23196 a_n1808_13878.n5 a_n1808_13878.n3 98.7517
R23197 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R23198 a_n1808_13878.n7 a_n1808_13878.n6 98.6055
R23199 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R23200 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R23201 a_n1808_13878.n9 a_n1808_13878.t1 74.6477
R23202 a_n1808_13878.n14 a_n1808_13878.t2 74.2899
R23203 a_n1808_13878.n11 a_n1808_13878.t3 74.2899
R23204 a_n1808_13878.n10 a_n1808_13878.t0 74.2899
R23205 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R23206 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R23207 a_n1808_13878.n15 a_n1808_13878.n7 13.5694
R23208 a_n1808_13878.n16 a_n1808_13878.n15 11.5762
R23209 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R23210 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R23211 a_n1808_13878.n1 a_n1808_13878.t13 3.61217
R23212 a_n1808_13878.n0 a_n1808_13878.t15 3.61217
R23213 a_n1808_13878.n0 a_n1808_13878.t19 3.61217
R23214 a_n1808_13878.n12 a_n1808_13878.t6 3.61217
R23215 a_n1808_13878.n12 a_n1808_13878.t7 3.61217
R23216 a_n1808_13878.n8 a_n1808_13878.t4 3.61217
R23217 a_n1808_13878.n8 a_n1808_13878.t5 3.61217
R23218 a_n1808_13878.n6 a_n1808_13878.t14 3.61217
R23219 a_n1808_13878.n6 a_n1808_13878.t9 3.61217
R23220 a_n1808_13878.n4 a_n1808_13878.t16 3.61217
R23221 a_n1808_13878.n4 a_n1808_13878.t11 3.61217
R23222 a_n1808_13878.n3 a_n1808_13878.t10 3.61217
R23223 a_n1808_13878.n3 a_n1808_13878.t12 3.61217
R23224 a_n1808_13878.n17 a_n1808_13878.t17 3.61217
R23225 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R23226 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R23227 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R23228 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R23229 a_n1808_13878.n16 a_n1808_13878.n2 0.358259
R23230 a_n1808_13878.n7 a_n1808_13878.n5 0.146627
R23231 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R23232 minus.n53 minus.t28 323.478
R23233 minus.n11 minus.t8 323.478
R23234 minus.n82 minus.t13 297.12
R23235 minus.n80 minus.t15 297.12
R23236 minus.n44 minus.t5 297.12
R23237 minus.n74 minus.t6 297.12
R23238 minus.n46 minus.t26 297.12
R23239 minus.n68 minus.t21 297.12
R23240 minus.n48 minus.t23 297.12
R23241 minus.n62 minus.t16 297.12
R23242 minus.n50 minus.t17 297.12
R23243 minus.n56 minus.t9 297.12
R23244 minus.n52 minus.t27 297.12
R23245 minus.n10 minus.t7 297.12
R23246 minus.n14 minus.t11 297.12
R23247 minus.n16 minus.t10 297.12
R23248 minus.n20 minus.t12 297.12
R23249 minus.n22 minus.t20 297.12
R23250 minus.n26 minus.t18 297.12
R23251 minus.n28 minus.t25 297.12
R23252 minus.n32 minus.t24 297.12
R23253 minus.n34 minus.t14 297.12
R23254 minus.n38 minus.t22 297.12
R23255 minus.n40 minus.t19 297.12
R23256 minus.n88 minus.t2 243.255
R23257 minus.n87 minus.n85 224.169
R23258 minus.n87 minus.n86 223.454
R23259 minus.n55 minus.n54 161.3
R23260 minus.n56 minus.n51 161.3
R23261 minus.n58 minus.n57 161.3
R23262 minus.n59 minus.n50 161.3
R23263 minus.n61 minus.n60 161.3
R23264 minus.n62 minus.n49 161.3
R23265 minus.n64 minus.n63 161.3
R23266 minus.n65 minus.n48 161.3
R23267 minus.n67 minus.n66 161.3
R23268 minus.n68 minus.n47 161.3
R23269 minus.n70 minus.n69 161.3
R23270 minus.n71 minus.n46 161.3
R23271 minus.n73 minus.n72 161.3
R23272 minus.n74 minus.n45 161.3
R23273 minus.n76 minus.n75 161.3
R23274 minus.n77 minus.n44 161.3
R23275 minus.n79 minus.n78 161.3
R23276 minus.n80 minus.n43 161.3
R23277 minus.n81 minus.n42 161.3
R23278 minus.n83 minus.n82 161.3
R23279 minus.n41 minus.n40 161.3
R23280 minus.n39 minus.n0 161.3
R23281 minus.n38 minus.n37 161.3
R23282 minus.n36 minus.n1 161.3
R23283 minus.n35 minus.n34 161.3
R23284 minus.n33 minus.n2 161.3
R23285 minus.n32 minus.n31 161.3
R23286 minus.n30 minus.n3 161.3
R23287 minus.n29 minus.n28 161.3
R23288 minus.n27 minus.n4 161.3
R23289 minus.n26 minus.n25 161.3
R23290 minus.n24 minus.n5 161.3
R23291 minus.n23 minus.n22 161.3
R23292 minus.n21 minus.n6 161.3
R23293 minus.n20 minus.n19 161.3
R23294 minus.n18 minus.n7 161.3
R23295 minus.n17 minus.n16 161.3
R23296 minus.n15 minus.n8 161.3
R23297 minus.n14 minus.n13 161.3
R23298 minus.n12 minus.n9 161.3
R23299 minus.n82 minus.n81 46.0096
R23300 minus.n40 minus.n39 46.0096
R23301 minus.n12 minus.n11 45.0871
R23302 minus.n54 minus.n53 45.0871
R23303 minus.n80 minus.n79 41.6278
R23304 minus.n55 minus.n52 41.6278
R23305 minus.n10 minus.n9 41.6278
R23306 minus.n38 minus.n1 41.6278
R23307 minus.n75 minus.n44 37.246
R23308 minus.n57 minus.n56 37.246
R23309 minus.n15 minus.n14 37.246
R23310 minus.n34 minus.n33 37.246
R23311 minus.n84 minus.n83 33.3925
R23312 minus.n74 minus.n73 32.8641
R23313 minus.n61 minus.n50 32.8641
R23314 minus.n16 minus.n7 32.8641
R23315 minus.n32 minus.n3 32.8641
R23316 minus.n69 minus.n46 28.4823
R23317 minus.n63 minus.n62 28.4823
R23318 minus.n21 minus.n20 28.4823
R23319 minus.n28 minus.n27 28.4823
R23320 minus.n68 minus.n67 24.1005
R23321 minus.n67 minus.n48 24.1005
R23322 minus.n22 minus.n5 24.1005
R23323 minus.n26 minus.n5 24.1005
R23324 minus.n86 minus.t4 19.8005
R23325 minus.n86 minus.t3 19.8005
R23326 minus.n85 minus.t1 19.8005
R23327 minus.n85 minus.t0 19.8005
R23328 minus.n69 minus.n68 19.7187
R23329 minus.n63 minus.n48 19.7187
R23330 minus.n22 minus.n21 19.7187
R23331 minus.n27 minus.n26 19.7187
R23332 minus.n73 minus.n46 15.3369
R23333 minus.n62 minus.n61 15.3369
R23334 minus.n20 minus.n7 15.3369
R23335 minus.n28 minus.n3 15.3369
R23336 minus.n53 minus.n52 14.1472
R23337 minus.n11 minus.n10 14.1472
R23338 minus.n84 minus.n41 12.0933
R23339 minus minus.n89 12.0331
R23340 minus.n75 minus.n74 10.955
R23341 minus.n57 minus.n50 10.955
R23342 minus.n16 minus.n15 10.955
R23343 minus.n33 minus.n32 10.955
R23344 minus.n79 minus.n44 6.57323
R23345 minus.n56 minus.n55 6.57323
R23346 minus.n14 minus.n9 6.57323
R23347 minus.n34 minus.n1 6.57323
R23348 minus.n89 minus.n88 4.80222
R23349 minus.n81 minus.n80 2.19141
R23350 minus.n39 minus.n38 2.19141
R23351 minus.n89 minus.n84 0.972091
R23352 minus.n88 minus.n87 0.716017
R23353 minus.n83 minus.n42 0.189894
R23354 minus.n43 minus.n42 0.189894
R23355 minus.n78 minus.n43 0.189894
R23356 minus.n78 minus.n77 0.189894
R23357 minus.n77 minus.n76 0.189894
R23358 minus.n76 minus.n45 0.189894
R23359 minus.n72 minus.n45 0.189894
R23360 minus.n72 minus.n71 0.189894
R23361 minus.n71 minus.n70 0.189894
R23362 minus.n70 minus.n47 0.189894
R23363 minus.n66 minus.n47 0.189894
R23364 minus.n66 minus.n65 0.189894
R23365 minus.n65 minus.n64 0.189894
R23366 minus.n64 minus.n49 0.189894
R23367 minus.n60 minus.n49 0.189894
R23368 minus.n60 minus.n59 0.189894
R23369 minus.n59 minus.n58 0.189894
R23370 minus.n58 minus.n51 0.189894
R23371 minus.n54 minus.n51 0.189894
R23372 minus.n13 minus.n12 0.189894
R23373 minus.n13 minus.n8 0.189894
R23374 minus.n17 minus.n8 0.189894
R23375 minus.n18 minus.n17 0.189894
R23376 minus.n19 minus.n18 0.189894
R23377 minus.n19 minus.n6 0.189894
R23378 minus.n23 minus.n6 0.189894
R23379 minus.n24 minus.n23 0.189894
R23380 minus.n25 minus.n24 0.189894
R23381 minus.n25 minus.n4 0.189894
R23382 minus.n29 minus.n4 0.189894
R23383 minus.n30 minus.n29 0.189894
R23384 minus.n31 minus.n30 0.189894
R23385 minus.n31 minus.n2 0.189894
R23386 minus.n35 minus.n2 0.189894
R23387 minus.n36 minus.n35 0.189894
R23388 minus.n37 minus.n36 0.189894
R23389 minus.n37 minus.n0 0.189894
R23390 minus.n41 minus.n0 0.189894
R23391 diffpairibias.n0 diffpairibias.t27 436.822
R23392 diffpairibias.n27 diffpairibias.t24 435.479
R23393 diffpairibias.n26 diffpairibias.t21 435.479
R23394 diffpairibias.n25 diffpairibias.t22 435.479
R23395 diffpairibias.n24 diffpairibias.t26 435.479
R23396 diffpairibias.n23 diffpairibias.t20 435.479
R23397 diffpairibias.n0 diffpairibias.t23 435.479
R23398 diffpairibias.n1 diffpairibias.t28 435.479
R23399 diffpairibias.n2 diffpairibias.t25 435.479
R23400 diffpairibias.n3 diffpairibias.t29 435.479
R23401 diffpairibias.n13 diffpairibias.t14 377.536
R23402 diffpairibias.n13 diffpairibias.t0 376.193
R23403 diffpairibias.n14 diffpairibias.t10 376.193
R23404 diffpairibias.n15 diffpairibias.t12 376.193
R23405 diffpairibias.n16 diffpairibias.t6 376.193
R23406 diffpairibias.n17 diffpairibias.t2 376.193
R23407 diffpairibias.n18 diffpairibias.t16 376.193
R23408 diffpairibias.n19 diffpairibias.t4 376.193
R23409 diffpairibias.n20 diffpairibias.t18 376.193
R23410 diffpairibias.n21 diffpairibias.t8 376.193
R23411 diffpairibias.n4 diffpairibias.t15 113.368
R23412 diffpairibias.n4 diffpairibias.t1 112.698
R23413 diffpairibias.n5 diffpairibias.t11 112.698
R23414 diffpairibias.n6 diffpairibias.t13 112.698
R23415 diffpairibias.n7 diffpairibias.t7 112.698
R23416 diffpairibias.n8 diffpairibias.t3 112.698
R23417 diffpairibias.n9 diffpairibias.t17 112.698
R23418 diffpairibias.n10 diffpairibias.t5 112.698
R23419 diffpairibias.n11 diffpairibias.t19 112.698
R23420 diffpairibias.n12 diffpairibias.t9 112.698
R23421 diffpairibias.n22 diffpairibias.n21 4.77242
R23422 diffpairibias.n22 diffpairibias.n12 4.30807
R23423 diffpairibias.n23 diffpairibias.n22 4.13945
R23424 diffpairibias.n21 diffpairibias.n20 1.34352
R23425 diffpairibias.n20 diffpairibias.n19 1.34352
R23426 diffpairibias.n19 diffpairibias.n18 1.34352
R23427 diffpairibias.n18 diffpairibias.n17 1.34352
R23428 diffpairibias.n17 diffpairibias.n16 1.34352
R23429 diffpairibias.n16 diffpairibias.n15 1.34352
R23430 diffpairibias.n15 diffpairibias.n14 1.34352
R23431 diffpairibias.n14 diffpairibias.n13 1.34352
R23432 diffpairibias.n3 diffpairibias.n2 1.34352
R23433 diffpairibias.n2 diffpairibias.n1 1.34352
R23434 diffpairibias.n1 diffpairibias.n0 1.34352
R23435 diffpairibias.n24 diffpairibias.n23 1.34352
R23436 diffpairibias.n25 diffpairibias.n24 1.34352
R23437 diffpairibias.n26 diffpairibias.n25 1.34352
R23438 diffpairibias.n27 diffpairibias.n26 1.34352
R23439 diffpairibias.n28 diffpairibias.n27 0.862419
R23440 diffpairibias diffpairibias.n28 0.684875
R23441 diffpairibias.n12 diffpairibias.n11 0.672012
R23442 diffpairibias.n11 diffpairibias.n10 0.672012
R23443 diffpairibias.n10 diffpairibias.n9 0.672012
R23444 diffpairibias.n9 diffpairibias.n8 0.672012
R23445 diffpairibias.n8 diffpairibias.n7 0.672012
R23446 diffpairibias.n7 diffpairibias.n6 0.672012
R23447 diffpairibias.n6 diffpairibias.n5 0.672012
R23448 diffpairibias.n5 diffpairibias.n4 0.672012
R23449 diffpairibias.n28 diffpairibias.n3 0.190907
R23450 a_n1986_8322.n6 a_n1986_8322.t3 74.6477
R23451 a_n1986_8322.n1 a_n1986_8322.t9 74.6477
R23452 a_n1986_8322.n16 a_n1986_8322.t18 74.6474
R23453 a_n1986_8322.n14 a_n1986_8322.t11 74.2899
R23454 a_n1986_8322.n7 a_n1986_8322.t1 74.2899
R23455 a_n1986_8322.n8 a_n1986_8322.t4 74.2899
R23456 a_n1986_8322.n11 a_n1986_8322.t5 74.2899
R23457 a_n1986_8322.n4 a_n1986_8322.t8 74.2899
R23458 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R23459 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R23460 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R23461 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R23462 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R23463 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R23464 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R23465 a_n1986_8322.n13 a_n1986_8322.t20 10.2757
R23466 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R23467 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R23468 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R23469 a_n1986_8322.n15 a_n1986_8322.t16 3.61217
R23470 a_n1986_8322.n15 a_n1986_8322.t13 3.61217
R23471 a_n1986_8322.n5 a_n1986_8322.t7 3.61217
R23472 a_n1986_8322.n5 a_n1986_8322.t6 3.61217
R23473 a_n1986_8322.n9 a_n1986_8322.t2 3.61217
R23474 a_n1986_8322.n9 a_n1986_8322.t0 3.61217
R23475 a_n1986_8322.n0 a_n1986_8322.t17 3.61217
R23476 a_n1986_8322.n0 a_n1986_8322.t12 3.61217
R23477 a_n1986_8322.n2 a_n1986_8322.t15 3.61217
R23478 a_n1986_8322.n2 a_n1986_8322.t14 3.61217
R23479 a_n1986_8322.n18 a_n1986_8322.t10 3.61217
R23480 a_n1986_8322.t19 a_n1986_8322.n18 3.61217
R23481 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R23482 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R23483 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R23484 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R23485 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R23486 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R23487 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R23488 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R23489 a_n1986_8322.t20 a_n1986_8322.t21 0.057021
R23490 outputibias.n27 outputibias.n1 289.615
R23491 outputibias.n58 outputibias.n32 289.615
R23492 outputibias.n90 outputibias.n64 289.615
R23493 outputibias.n122 outputibias.n96 289.615
R23494 outputibias.n28 outputibias.n27 185
R23495 outputibias.n26 outputibias.n25 185
R23496 outputibias.n5 outputibias.n4 185
R23497 outputibias.n20 outputibias.n19 185
R23498 outputibias.n18 outputibias.n17 185
R23499 outputibias.n9 outputibias.n8 185
R23500 outputibias.n12 outputibias.n11 185
R23501 outputibias.n59 outputibias.n58 185
R23502 outputibias.n57 outputibias.n56 185
R23503 outputibias.n36 outputibias.n35 185
R23504 outputibias.n51 outputibias.n50 185
R23505 outputibias.n49 outputibias.n48 185
R23506 outputibias.n40 outputibias.n39 185
R23507 outputibias.n43 outputibias.n42 185
R23508 outputibias.n91 outputibias.n90 185
R23509 outputibias.n89 outputibias.n88 185
R23510 outputibias.n68 outputibias.n67 185
R23511 outputibias.n83 outputibias.n82 185
R23512 outputibias.n81 outputibias.n80 185
R23513 outputibias.n72 outputibias.n71 185
R23514 outputibias.n75 outputibias.n74 185
R23515 outputibias.n123 outputibias.n122 185
R23516 outputibias.n121 outputibias.n120 185
R23517 outputibias.n100 outputibias.n99 185
R23518 outputibias.n115 outputibias.n114 185
R23519 outputibias.n113 outputibias.n112 185
R23520 outputibias.n104 outputibias.n103 185
R23521 outputibias.n107 outputibias.n106 185
R23522 outputibias.n0 outputibias.t11 178.945
R23523 outputibias.n133 outputibias.t8 177.018
R23524 outputibias.n132 outputibias.t10 177.018
R23525 outputibias.n0 outputibias.t9 177.018
R23526 outputibias.t5 outputibias.n10 147.661
R23527 outputibias.t7 outputibias.n41 147.661
R23528 outputibias.t3 outputibias.n73 147.661
R23529 outputibias.t1 outputibias.n105 147.661
R23530 outputibias.n128 outputibias.t4 132.363
R23531 outputibias.n128 outputibias.t6 130.436
R23532 outputibias.n129 outputibias.t2 130.436
R23533 outputibias.n130 outputibias.t0 130.436
R23534 outputibias.n27 outputibias.n26 104.615
R23535 outputibias.n26 outputibias.n4 104.615
R23536 outputibias.n19 outputibias.n4 104.615
R23537 outputibias.n19 outputibias.n18 104.615
R23538 outputibias.n18 outputibias.n8 104.615
R23539 outputibias.n11 outputibias.n8 104.615
R23540 outputibias.n58 outputibias.n57 104.615
R23541 outputibias.n57 outputibias.n35 104.615
R23542 outputibias.n50 outputibias.n35 104.615
R23543 outputibias.n50 outputibias.n49 104.615
R23544 outputibias.n49 outputibias.n39 104.615
R23545 outputibias.n42 outputibias.n39 104.615
R23546 outputibias.n90 outputibias.n89 104.615
R23547 outputibias.n89 outputibias.n67 104.615
R23548 outputibias.n82 outputibias.n67 104.615
R23549 outputibias.n82 outputibias.n81 104.615
R23550 outputibias.n81 outputibias.n71 104.615
R23551 outputibias.n74 outputibias.n71 104.615
R23552 outputibias.n122 outputibias.n121 104.615
R23553 outputibias.n121 outputibias.n99 104.615
R23554 outputibias.n114 outputibias.n99 104.615
R23555 outputibias.n114 outputibias.n113 104.615
R23556 outputibias.n113 outputibias.n103 104.615
R23557 outputibias.n106 outputibias.n103 104.615
R23558 outputibias.n63 outputibias.n31 95.6354
R23559 outputibias.n63 outputibias.n62 94.6732
R23560 outputibias.n95 outputibias.n94 94.6732
R23561 outputibias.n127 outputibias.n126 94.6732
R23562 outputibias.n11 outputibias.t5 52.3082
R23563 outputibias.n42 outputibias.t7 52.3082
R23564 outputibias.n74 outputibias.t3 52.3082
R23565 outputibias.n106 outputibias.t1 52.3082
R23566 outputibias.n12 outputibias.n10 15.6674
R23567 outputibias.n43 outputibias.n41 15.6674
R23568 outputibias.n75 outputibias.n73 15.6674
R23569 outputibias.n107 outputibias.n105 15.6674
R23570 outputibias.n13 outputibias.n9 12.8005
R23571 outputibias.n44 outputibias.n40 12.8005
R23572 outputibias.n76 outputibias.n72 12.8005
R23573 outputibias.n108 outputibias.n104 12.8005
R23574 outputibias.n17 outputibias.n16 12.0247
R23575 outputibias.n48 outputibias.n47 12.0247
R23576 outputibias.n80 outputibias.n79 12.0247
R23577 outputibias.n112 outputibias.n111 12.0247
R23578 outputibias.n20 outputibias.n7 11.249
R23579 outputibias.n51 outputibias.n38 11.249
R23580 outputibias.n83 outputibias.n70 11.249
R23581 outputibias.n115 outputibias.n102 11.249
R23582 outputibias.n21 outputibias.n5 10.4732
R23583 outputibias.n52 outputibias.n36 10.4732
R23584 outputibias.n84 outputibias.n68 10.4732
R23585 outputibias.n116 outputibias.n100 10.4732
R23586 outputibias.n25 outputibias.n24 9.69747
R23587 outputibias.n56 outputibias.n55 9.69747
R23588 outputibias.n88 outputibias.n87 9.69747
R23589 outputibias.n120 outputibias.n119 9.69747
R23590 outputibias.n31 outputibias.n30 9.45567
R23591 outputibias.n62 outputibias.n61 9.45567
R23592 outputibias.n94 outputibias.n93 9.45567
R23593 outputibias.n126 outputibias.n125 9.45567
R23594 outputibias.n30 outputibias.n29 9.3005
R23595 outputibias.n3 outputibias.n2 9.3005
R23596 outputibias.n24 outputibias.n23 9.3005
R23597 outputibias.n22 outputibias.n21 9.3005
R23598 outputibias.n7 outputibias.n6 9.3005
R23599 outputibias.n16 outputibias.n15 9.3005
R23600 outputibias.n14 outputibias.n13 9.3005
R23601 outputibias.n61 outputibias.n60 9.3005
R23602 outputibias.n34 outputibias.n33 9.3005
R23603 outputibias.n55 outputibias.n54 9.3005
R23604 outputibias.n53 outputibias.n52 9.3005
R23605 outputibias.n38 outputibias.n37 9.3005
R23606 outputibias.n47 outputibias.n46 9.3005
R23607 outputibias.n45 outputibias.n44 9.3005
R23608 outputibias.n93 outputibias.n92 9.3005
R23609 outputibias.n66 outputibias.n65 9.3005
R23610 outputibias.n87 outputibias.n86 9.3005
R23611 outputibias.n85 outputibias.n84 9.3005
R23612 outputibias.n70 outputibias.n69 9.3005
R23613 outputibias.n79 outputibias.n78 9.3005
R23614 outputibias.n77 outputibias.n76 9.3005
R23615 outputibias.n125 outputibias.n124 9.3005
R23616 outputibias.n98 outputibias.n97 9.3005
R23617 outputibias.n119 outputibias.n118 9.3005
R23618 outputibias.n117 outputibias.n116 9.3005
R23619 outputibias.n102 outputibias.n101 9.3005
R23620 outputibias.n111 outputibias.n110 9.3005
R23621 outputibias.n109 outputibias.n108 9.3005
R23622 outputibias.n28 outputibias.n3 8.92171
R23623 outputibias.n59 outputibias.n34 8.92171
R23624 outputibias.n91 outputibias.n66 8.92171
R23625 outputibias.n123 outputibias.n98 8.92171
R23626 outputibias.n29 outputibias.n1 8.14595
R23627 outputibias.n60 outputibias.n32 8.14595
R23628 outputibias.n92 outputibias.n64 8.14595
R23629 outputibias.n124 outputibias.n96 8.14595
R23630 outputibias.n31 outputibias.n1 5.81868
R23631 outputibias.n62 outputibias.n32 5.81868
R23632 outputibias.n94 outputibias.n64 5.81868
R23633 outputibias.n126 outputibias.n96 5.81868
R23634 outputibias.n131 outputibias.n130 5.20947
R23635 outputibias.n29 outputibias.n28 5.04292
R23636 outputibias.n60 outputibias.n59 5.04292
R23637 outputibias.n92 outputibias.n91 5.04292
R23638 outputibias.n124 outputibias.n123 5.04292
R23639 outputibias.n131 outputibias.n127 4.42209
R23640 outputibias.n14 outputibias.n10 4.38594
R23641 outputibias.n45 outputibias.n41 4.38594
R23642 outputibias.n77 outputibias.n73 4.38594
R23643 outputibias.n109 outputibias.n105 4.38594
R23644 outputibias.n132 outputibias.n131 4.28454
R23645 outputibias.n25 outputibias.n3 4.26717
R23646 outputibias.n56 outputibias.n34 4.26717
R23647 outputibias.n88 outputibias.n66 4.26717
R23648 outputibias.n120 outputibias.n98 4.26717
R23649 outputibias.n24 outputibias.n5 3.49141
R23650 outputibias.n55 outputibias.n36 3.49141
R23651 outputibias.n87 outputibias.n68 3.49141
R23652 outputibias.n119 outputibias.n100 3.49141
R23653 outputibias.n21 outputibias.n20 2.71565
R23654 outputibias.n52 outputibias.n51 2.71565
R23655 outputibias.n84 outputibias.n83 2.71565
R23656 outputibias.n116 outputibias.n115 2.71565
R23657 outputibias.n17 outputibias.n7 1.93989
R23658 outputibias.n48 outputibias.n38 1.93989
R23659 outputibias.n80 outputibias.n70 1.93989
R23660 outputibias.n112 outputibias.n102 1.93989
R23661 outputibias.n130 outputibias.n129 1.9266
R23662 outputibias.n129 outputibias.n128 1.9266
R23663 outputibias.n133 outputibias.n132 1.92658
R23664 outputibias.n134 outputibias.n133 1.29913
R23665 outputibias.n16 outputibias.n9 1.16414
R23666 outputibias.n47 outputibias.n40 1.16414
R23667 outputibias.n79 outputibias.n72 1.16414
R23668 outputibias.n111 outputibias.n104 1.16414
R23669 outputibias.n127 outputibias.n95 0.962709
R23670 outputibias.n95 outputibias.n63 0.962709
R23671 outputibias.n13 outputibias.n12 0.388379
R23672 outputibias.n44 outputibias.n43 0.388379
R23673 outputibias.n76 outputibias.n75 0.388379
R23674 outputibias.n108 outputibias.n107 0.388379
R23675 outputibias.n134 outputibias.n0 0.337251
R23676 outputibias outputibias.n134 0.302375
R23677 outputibias.n30 outputibias.n2 0.155672
R23678 outputibias.n23 outputibias.n2 0.155672
R23679 outputibias.n23 outputibias.n22 0.155672
R23680 outputibias.n22 outputibias.n6 0.155672
R23681 outputibias.n15 outputibias.n6 0.155672
R23682 outputibias.n15 outputibias.n14 0.155672
R23683 outputibias.n61 outputibias.n33 0.155672
R23684 outputibias.n54 outputibias.n33 0.155672
R23685 outputibias.n54 outputibias.n53 0.155672
R23686 outputibias.n53 outputibias.n37 0.155672
R23687 outputibias.n46 outputibias.n37 0.155672
R23688 outputibias.n46 outputibias.n45 0.155672
R23689 outputibias.n93 outputibias.n65 0.155672
R23690 outputibias.n86 outputibias.n65 0.155672
R23691 outputibias.n86 outputibias.n85 0.155672
R23692 outputibias.n85 outputibias.n69 0.155672
R23693 outputibias.n78 outputibias.n69 0.155672
R23694 outputibias.n78 outputibias.n77 0.155672
R23695 outputibias.n125 outputibias.n97 0.155672
R23696 outputibias.n118 outputibias.n97 0.155672
R23697 outputibias.n118 outputibias.n117 0.155672
R23698 outputibias.n117 outputibias.n101 0.155672
R23699 outputibias.n110 outputibias.n101 0.155672
R23700 outputibias.n110 outputibias.n109 0.155672
R23701 output.n41 output.n15 289.615
R23702 output.n72 output.n46 289.615
R23703 output.n104 output.n78 289.615
R23704 output.n136 output.n110 289.615
R23705 output.n77 output.n45 197.26
R23706 output.n77 output.n76 196.298
R23707 output.n109 output.n108 196.298
R23708 output.n141 output.n140 196.298
R23709 output.n42 output.n41 185
R23710 output.n40 output.n39 185
R23711 output.n19 output.n18 185
R23712 output.n34 output.n33 185
R23713 output.n32 output.n31 185
R23714 output.n23 output.n22 185
R23715 output.n26 output.n25 185
R23716 output.n73 output.n72 185
R23717 output.n71 output.n70 185
R23718 output.n50 output.n49 185
R23719 output.n65 output.n64 185
R23720 output.n63 output.n62 185
R23721 output.n54 output.n53 185
R23722 output.n57 output.n56 185
R23723 output.n105 output.n104 185
R23724 output.n103 output.n102 185
R23725 output.n82 output.n81 185
R23726 output.n97 output.n96 185
R23727 output.n95 output.n94 185
R23728 output.n86 output.n85 185
R23729 output.n89 output.n88 185
R23730 output.n137 output.n136 185
R23731 output.n135 output.n134 185
R23732 output.n114 output.n113 185
R23733 output.n129 output.n128 185
R23734 output.n127 output.n126 185
R23735 output.n118 output.n117 185
R23736 output.n121 output.n120 185
R23737 output.t0 output.n24 147.661
R23738 output.t2 output.n55 147.661
R23739 output.t3 output.n87 147.661
R23740 output.t1 output.n119 147.661
R23741 output.n41 output.n40 104.615
R23742 output.n40 output.n18 104.615
R23743 output.n33 output.n18 104.615
R23744 output.n33 output.n32 104.615
R23745 output.n32 output.n22 104.615
R23746 output.n25 output.n22 104.615
R23747 output.n72 output.n71 104.615
R23748 output.n71 output.n49 104.615
R23749 output.n64 output.n49 104.615
R23750 output.n64 output.n63 104.615
R23751 output.n63 output.n53 104.615
R23752 output.n56 output.n53 104.615
R23753 output.n104 output.n103 104.615
R23754 output.n103 output.n81 104.615
R23755 output.n96 output.n81 104.615
R23756 output.n96 output.n95 104.615
R23757 output.n95 output.n85 104.615
R23758 output.n88 output.n85 104.615
R23759 output.n136 output.n135 104.615
R23760 output.n135 output.n113 104.615
R23761 output.n128 output.n113 104.615
R23762 output.n128 output.n127 104.615
R23763 output.n127 output.n117 104.615
R23764 output.n120 output.n117 104.615
R23765 output.n1 output.t5 77.056
R23766 output.n14 output.t7 76.6694
R23767 output.n1 output.n0 72.7095
R23768 output.n3 output.n2 72.7095
R23769 output.n5 output.n4 72.7095
R23770 output.n7 output.n6 72.7095
R23771 output.n9 output.n8 72.7095
R23772 output.n11 output.n10 72.7095
R23773 output.n13 output.n12 72.7095
R23774 output.n25 output.t0 52.3082
R23775 output.n56 output.t2 52.3082
R23776 output.n88 output.t3 52.3082
R23777 output.n120 output.t1 52.3082
R23778 output.n26 output.n24 15.6674
R23779 output.n57 output.n55 15.6674
R23780 output.n89 output.n87 15.6674
R23781 output.n121 output.n119 15.6674
R23782 output.n27 output.n23 12.8005
R23783 output.n58 output.n54 12.8005
R23784 output.n90 output.n86 12.8005
R23785 output.n122 output.n118 12.8005
R23786 output.n31 output.n30 12.0247
R23787 output.n62 output.n61 12.0247
R23788 output.n94 output.n93 12.0247
R23789 output.n126 output.n125 12.0247
R23790 output.n34 output.n21 11.249
R23791 output.n65 output.n52 11.249
R23792 output.n97 output.n84 11.249
R23793 output.n129 output.n116 11.249
R23794 output.n35 output.n19 10.4732
R23795 output.n66 output.n50 10.4732
R23796 output.n98 output.n82 10.4732
R23797 output.n130 output.n114 10.4732
R23798 output.n39 output.n38 9.69747
R23799 output.n70 output.n69 9.69747
R23800 output.n102 output.n101 9.69747
R23801 output.n134 output.n133 9.69747
R23802 output.n45 output.n44 9.45567
R23803 output.n76 output.n75 9.45567
R23804 output.n108 output.n107 9.45567
R23805 output.n140 output.n139 9.45567
R23806 output.n44 output.n43 9.3005
R23807 output.n17 output.n16 9.3005
R23808 output.n38 output.n37 9.3005
R23809 output.n36 output.n35 9.3005
R23810 output.n21 output.n20 9.3005
R23811 output.n30 output.n29 9.3005
R23812 output.n28 output.n27 9.3005
R23813 output.n75 output.n74 9.3005
R23814 output.n48 output.n47 9.3005
R23815 output.n69 output.n68 9.3005
R23816 output.n67 output.n66 9.3005
R23817 output.n52 output.n51 9.3005
R23818 output.n61 output.n60 9.3005
R23819 output.n59 output.n58 9.3005
R23820 output.n107 output.n106 9.3005
R23821 output.n80 output.n79 9.3005
R23822 output.n101 output.n100 9.3005
R23823 output.n99 output.n98 9.3005
R23824 output.n84 output.n83 9.3005
R23825 output.n93 output.n92 9.3005
R23826 output.n91 output.n90 9.3005
R23827 output.n139 output.n138 9.3005
R23828 output.n112 output.n111 9.3005
R23829 output.n133 output.n132 9.3005
R23830 output.n131 output.n130 9.3005
R23831 output.n116 output.n115 9.3005
R23832 output.n125 output.n124 9.3005
R23833 output.n123 output.n122 9.3005
R23834 output.n42 output.n17 8.92171
R23835 output.n73 output.n48 8.92171
R23836 output.n105 output.n80 8.92171
R23837 output.n137 output.n112 8.92171
R23838 output output.n141 8.15037
R23839 output.n43 output.n15 8.14595
R23840 output.n74 output.n46 8.14595
R23841 output.n106 output.n78 8.14595
R23842 output.n138 output.n110 8.14595
R23843 output.n45 output.n15 5.81868
R23844 output.n76 output.n46 5.81868
R23845 output.n108 output.n78 5.81868
R23846 output.n140 output.n110 5.81868
R23847 output.n43 output.n42 5.04292
R23848 output.n74 output.n73 5.04292
R23849 output.n106 output.n105 5.04292
R23850 output.n138 output.n137 5.04292
R23851 output.n28 output.n24 4.38594
R23852 output.n59 output.n55 4.38594
R23853 output.n91 output.n87 4.38594
R23854 output.n123 output.n119 4.38594
R23855 output.n39 output.n17 4.26717
R23856 output.n70 output.n48 4.26717
R23857 output.n102 output.n80 4.26717
R23858 output.n134 output.n112 4.26717
R23859 output.n0 output.t11 3.9605
R23860 output.n0 output.t16 3.9605
R23861 output.n2 output.t4 3.9605
R23862 output.n2 output.t12 3.9605
R23863 output.n4 output.t14 3.9605
R23864 output.n4 output.t13 3.9605
R23865 output.n6 output.t19 3.9605
R23866 output.n6 output.t6 3.9605
R23867 output.n8 output.t8 3.9605
R23868 output.n8 output.t17 3.9605
R23869 output.n10 output.t18 3.9605
R23870 output.n10 output.t9 3.9605
R23871 output.n12 output.t10 3.9605
R23872 output.n12 output.t15 3.9605
R23873 output.n38 output.n19 3.49141
R23874 output.n69 output.n50 3.49141
R23875 output.n101 output.n82 3.49141
R23876 output.n133 output.n114 3.49141
R23877 output.n35 output.n34 2.71565
R23878 output.n66 output.n65 2.71565
R23879 output.n98 output.n97 2.71565
R23880 output.n130 output.n129 2.71565
R23881 output.n31 output.n21 1.93989
R23882 output.n62 output.n52 1.93989
R23883 output.n94 output.n84 1.93989
R23884 output.n126 output.n116 1.93989
R23885 output.n30 output.n23 1.16414
R23886 output.n61 output.n54 1.16414
R23887 output.n93 output.n86 1.16414
R23888 output.n125 output.n118 1.16414
R23889 output.n141 output.n109 0.962709
R23890 output.n109 output.n77 0.962709
R23891 output.n27 output.n26 0.388379
R23892 output.n58 output.n57 0.388379
R23893 output.n90 output.n89 0.388379
R23894 output.n122 output.n121 0.388379
R23895 output.n14 output.n13 0.387128
R23896 output.n13 output.n11 0.387128
R23897 output.n11 output.n9 0.387128
R23898 output.n9 output.n7 0.387128
R23899 output.n7 output.n5 0.387128
R23900 output.n5 output.n3 0.387128
R23901 output.n3 output.n1 0.387128
R23902 output.n44 output.n16 0.155672
R23903 output.n37 output.n16 0.155672
R23904 output.n37 output.n36 0.155672
R23905 output.n36 output.n20 0.155672
R23906 output.n29 output.n20 0.155672
R23907 output.n29 output.n28 0.155672
R23908 output.n75 output.n47 0.155672
R23909 output.n68 output.n47 0.155672
R23910 output.n68 output.n67 0.155672
R23911 output.n67 output.n51 0.155672
R23912 output.n60 output.n51 0.155672
R23913 output.n60 output.n59 0.155672
R23914 output.n107 output.n79 0.155672
R23915 output.n100 output.n79 0.155672
R23916 output.n100 output.n99 0.155672
R23917 output.n99 output.n83 0.155672
R23918 output.n92 output.n83 0.155672
R23919 output.n92 output.n91 0.155672
R23920 output.n139 output.n111 0.155672
R23921 output.n132 output.n111 0.155672
R23922 output.n132 output.n131 0.155672
R23923 output.n131 output.n115 0.155672
R23924 output.n124 output.n115 0.155672
R23925 output.n124 output.n123 0.155672
R23926 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13881f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 91.9904f
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 4.33e-19
C7 CSoutput minus 3.17016f
C8 vdd plus 0.077622f
C9 plus diffpairibias 4.56e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.91196f
C13 commonsourceibias diffpairibias 0.064336f
C14 CSoutput commonsourceibias 66.8263f
C15 minus plus 10.303599f
C16 minus commonsourceibias 0.337549f
C17 plus commonsourceibias 0.283677f
C18 diffpairibias gnd 60.00273f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.223205p
C22 plus gnd 37.739304f
C23 minus gnd 31.372768f
C24 CSoutput gnd 0.145127p
C25 vdd gnd 0.377108p
C26 output.t5 gnd 0.464308f
C27 output.t11 gnd 0.044422f
C28 output.t16 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t4 gnd 0.044422f
C32 output.t12 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t14 gnd 0.044422f
C36 output.t13 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t19 gnd 0.044422f
C40 output.t6 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t8 gnd 0.044422f
C44 output.t17 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t18 gnd 0.044422f
C48 output.t9 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t10 gnd 0.044422f
C52 output.t15 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t7 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t0 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t2 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t3 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t1 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 outputibias.t9 gnd 0.11477f
C189 outputibias.t11 gnd 0.115567f
C190 outputibias.n0 gnd 0.130108f
C191 outputibias.n1 gnd 0.001372f
C192 outputibias.n2 gnd 9.76e-19
C193 outputibias.n3 gnd 5.24e-19
C194 outputibias.n4 gnd 0.001239f
C195 outputibias.n5 gnd 5.55e-19
C196 outputibias.n6 gnd 9.76e-19
C197 outputibias.n7 gnd 5.24e-19
C198 outputibias.n8 gnd 0.001239f
C199 outputibias.n9 gnd 5.55e-19
C200 outputibias.n10 gnd 0.004176f
C201 outputibias.t5 gnd 0.00202f
C202 outputibias.n11 gnd 9.3e-19
C203 outputibias.n12 gnd 7.32e-19
C204 outputibias.n13 gnd 5.24e-19
C205 outputibias.n14 gnd 0.02322f
C206 outputibias.n15 gnd 9.76e-19
C207 outputibias.n16 gnd 5.24e-19
C208 outputibias.n17 gnd 5.55e-19
C209 outputibias.n18 gnd 0.001239f
C210 outputibias.n19 gnd 0.001239f
C211 outputibias.n20 gnd 5.55e-19
C212 outputibias.n21 gnd 5.24e-19
C213 outputibias.n22 gnd 9.76e-19
C214 outputibias.n23 gnd 9.76e-19
C215 outputibias.n24 gnd 5.24e-19
C216 outputibias.n25 gnd 5.55e-19
C217 outputibias.n26 gnd 0.001239f
C218 outputibias.n27 gnd 0.002683f
C219 outputibias.n28 gnd 5.55e-19
C220 outputibias.n29 gnd 5.24e-19
C221 outputibias.n30 gnd 0.002256f
C222 outputibias.n31 gnd 0.005781f
C223 outputibias.n32 gnd 0.001372f
C224 outputibias.n33 gnd 9.76e-19
C225 outputibias.n34 gnd 5.24e-19
C226 outputibias.n35 gnd 0.001239f
C227 outputibias.n36 gnd 5.55e-19
C228 outputibias.n37 gnd 9.76e-19
C229 outputibias.n38 gnd 5.24e-19
C230 outputibias.n39 gnd 0.001239f
C231 outputibias.n40 gnd 5.55e-19
C232 outputibias.n41 gnd 0.004176f
C233 outputibias.t7 gnd 0.00202f
C234 outputibias.n42 gnd 9.3e-19
C235 outputibias.n43 gnd 7.32e-19
C236 outputibias.n44 gnd 5.24e-19
C237 outputibias.n45 gnd 0.02322f
C238 outputibias.n46 gnd 9.76e-19
C239 outputibias.n47 gnd 5.24e-19
C240 outputibias.n48 gnd 5.55e-19
C241 outputibias.n49 gnd 0.001239f
C242 outputibias.n50 gnd 0.001239f
C243 outputibias.n51 gnd 5.55e-19
C244 outputibias.n52 gnd 5.24e-19
C245 outputibias.n53 gnd 9.76e-19
C246 outputibias.n54 gnd 9.76e-19
C247 outputibias.n55 gnd 5.24e-19
C248 outputibias.n56 gnd 5.55e-19
C249 outputibias.n57 gnd 0.001239f
C250 outputibias.n58 gnd 0.002683f
C251 outputibias.n59 gnd 5.55e-19
C252 outputibias.n60 gnd 5.24e-19
C253 outputibias.n61 gnd 0.002256f
C254 outputibias.n62 gnd 0.005197f
C255 outputibias.n63 gnd 0.121892f
C256 outputibias.n64 gnd 0.001372f
C257 outputibias.n65 gnd 9.76e-19
C258 outputibias.n66 gnd 5.24e-19
C259 outputibias.n67 gnd 0.001239f
C260 outputibias.n68 gnd 5.55e-19
C261 outputibias.n69 gnd 9.76e-19
C262 outputibias.n70 gnd 5.24e-19
C263 outputibias.n71 gnd 0.001239f
C264 outputibias.n72 gnd 5.55e-19
C265 outputibias.n73 gnd 0.004176f
C266 outputibias.t3 gnd 0.00202f
C267 outputibias.n74 gnd 9.3e-19
C268 outputibias.n75 gnd 7.32e-19
C269 outputibias.n76 gnd 5.24e-19
C270 outputibias.n77 gnd 0.02322f
C271 outputibias.n78 gnd 9.76e-19
C272 outputibias.n79 gnd 5.24e-19
C273 outputibias.n80 gnd 5.55e-19
C274 outputibias.n81 gnd 0.001239f
C275 outputibias.n82 gnd 0.001239f
C276 outputibias.n83 gnd 5.55e-19
C277 outputibias.n84 gnd 5.24e-19
C278 outputibias.n85 gnd 9.76e-19
C279 outputibias.n86 gnd 9.76e-19
C280 outputibias.n87 gnd 5.24e-19
C281 outputibias.n88 gnd 5.55e-19
C282 outputibias.n89 gnd 0.001239f
C283 outputibias.n90 gnd 0.002683f
C284 outputibias.n91 gnd 5.55e-19
C285 outputibias.n92 gnd 5.24e-19
C286 outputibias.n93 gnd 0.002256f
C287 outputibias.n94 gnd 0.005197f
C288 outputibias.n95 gnd 0.064513f
C289 outputibias.n96 gnd 0.001372f
C290 outputibias.n97 gnd 9.76e-19
C291 outputibias.n98 gnd 5.24e-19
C292 outputibias.n99 gnd 0.001239f
C293 outputibias.n100 gnd 5.55e-19
C294 outputibias.n101 gnd 9.76e-19
C295 outputibias.n102 gnd 5.24e-19
C296 outputibias.n103 gnd 0.001239f
C297 outputibias.n104 gnd 5.55e-19
C298 outputibias.n105 gnd 0.004176f
C299 outputibias.t1 gnd 0.00202f
C300 outputibias.n106 gnd 9.3e-19
C301 outputibias.n107 gnd 7.32e-19
C302 outputibias.n108 gnd 5.24e-19
C303 outputibias.n109 gnd 0.02322f
C304 outputibias.n110 gnd 9.76e-19
C305 outputibias.n111 gnd 5.24e-19
C306 outputibias.n112 gnd 5.55e-19
C307 outputibias.n113 gnd 0.001239f
C308 outputibias.n114 gnd 0.001239f
C309 outputibias.n115 gnd 5.55e-19
C310 outputibias.n116 gnd 5.24e-19
C311 outputibias.n117 gnd 9.76e-19
C312 outputibias.n118 gnd 9.76e-19
C313 outputibias.n119 gnd 5.24e-19
C314 outputibias.n120 gnd 5.55e-19
C315 outputibias.n121 gnd 0.001239f
C316 outputibias.n122 gnd 0.002683f
C317 outputibias.n123 gnd 5.55e-19
C318 outputibias.n124 gnd 5.24e-19
C319 outputibias.n125 gnd 0.002256f
C320 outputibias.n126 gnd 0.005197f
C321 outputibias.n127 gnd 0.084814f
C322 outputibias.t0 gnd 0.108319f
C323 outputibias.t2 gnd 0.108319f
C324 outputibias.t6 gnd 0.108319f
C325 outputibias.t4 gnd 0.109238f
C326 outputibias.n128 gnd 0.134674f
C327 outputibias.n129 gnd 0.07244f
C328 outputibias.n130 gnd 0.079818f
C329 outputibias.n131 gnd 0.164901f
C330 outputibias.t10 gnd 0.11477f
C331 outputibias.n132 gnd 0.067481f
C332 outputibias.t8 gnd 0.11477f
C333 outputibias.n133 gnd 0.065115f
C334 outputibias.n134 gnd 0.029159f
C335 a_n1986_8322.t21 gnd 49.329998f
C336 a_n1986_8322.t20 gnd 76.771f
C337 a_n1986_8322.t10 gnd 0.09348f
C338 a_n1986_8322.t9 gnd 0.875297f
C339 a_n1986_8322.t17 gnd 0.09348f
C340 a_n1986_8322.t12 gnd 0.09348f
C341 a_n1986_8322.n0 gnd 0.658471f
C342 a_n1986_8322.n1 gnd 0.735745f
C343 a_n1986_8322.t15 gnd 0.09348f
C344 a_n1986_8322.t14 gnd 0.09348f
C345 a_n1986_8322.n2 gnd 0.658471f
C346 a_n1986_8322.n3 gnd 0.373822f
C347 a_n1986_8322.t8 gnd 0.873554f
C348 a_n1986_8322.n4 gnd 1.39817f
C349 a_n1986_8322.t3 gnd 0.875297f
C350 a_n1986_8322.t7 gnd 0.09348f
C351 a_n1986_8322.t6 gnd 0.09348f
C352 a_n1986_8322.n5 gnd 0.658471f
C353 a_n1986_8322.n6 gnd 0.735745f
C354 a_n1986_8322.t1 gnd 0.873554f
C355 a_n1986_8322.n7 gnd 0.370237f
C356 a_n1986_8322.t4 gnd 0.873554f
C357 a_n1986_8322.n8 gnd 0.370237f
C358 a_n1986_8322.t2 gnd 0.09348f
C359 a_n1986_8322.t0 gnd 0.09348f
C360 a_n1986_8322.n9 gnd 0.658471f
C361 a_n1986_8322.n10 gnd 0.373822f
C362 a_n1986_8322.t5 gnd 0.873554f
C363 a_n1986_8322.n11 gnd 0.871824f
C364 a_n1986_8322.n12 gnd 1.58981f
C365 a_n1986_8322.n13 gnd 4.0376f
C366 a_n1986_8322.t11 gnd 0.873554f
C367 a_n1986_8322.n14 gnd 0.766087f
C368 a_n1986_8322.t18 gnd 0.875294f
C369 a_n1986_8322.t16 gnd 0.09348f
C370 a_n1986_8322.t13 gnd 0.09348f
C371 a_n1986_8322.n15 gnd 0.658471f
C372 a_n1986_8322.n16 gnd 0.735747f
C373 a_n1986_8322.n17 gnd 0.373821f
C374 a_n1986_8322.n18 gnd 0.658473f
C375 a_n1986_8322.t19 gnd 0.09348f
C376 diffpairibias.t27 gnd 0.090128f
C377 diffpairibias.t23 gnd 0.08996f
C378 diffpairibias.n0 gnd 0.105991f
C379 diffpairibias.t28 gnd 0.08996f
C380 diffpairibias.n1 gnd 0.051736f
C381 diffpairibias.t25 gnd 0.08996f
C382 diffpairibias.n2 gnd 0.051736f
C383 diffpairibias.t29 gnd 0.08996f
C384 diffpairibias.n3 gnd 0.041084f
C385 diffpairibias.t15 gnd 0.086371f
C386 diffpairibias.t1 gnd 0.085993f
C387 diffpairibias.n4 gnd 0.13579f
C388 diffpairibias.t11 gnd 0.085993f
C389 diffpairibias.n5 gnd 0.072463f
C390 diffpairibias.t13 gnd 0.085993f
C391 diffpairibias.n6 gnd 0.072463f
C392 diffpairibias.t7 gnd 0.085993f
C393 diffpairibias.n7 gnd 0.072463f
C394 diffpairibias.t3 gnd 0.085993f
C395 diffpairibias.n8 gnd 0.072463f
C396 diffpairibias.t17 gnd 0.085993f
C397 diffpairibias.n9 gnd 0.072463f
C398 diffpairibias.t5 gnd 0.085993f
C399 diffpairibias.n10 gnd 0.072463f
C400 diffpairibias.t19 gnd 0.085993f
C401 diffpairibias.n11 gnd 0.072463f
C402 diffpairibias.t9 gnd 0.085993f
C403 diffpairibias.n12 gnd 0.102883f
C404 diffpairibias.t14 gnd 0.086899f
C405 diffpairibias.t0 gnd 0.086748f
C406 diffpairibias.n13 gnd 0.094648f
C407 diffpairibias.t10 gnd 0.086748f
C408 diffpairibias.n14 gnd 0.052262f
C409 diffpairibias.t12 gnd 0.086748f
C410 diffpairibias.n15 gnd 0.052262f
C411 diffpairibias.t6 gnd 0.086748f
C412 diffpairibias.n16 gnd 0.052262f
C413 diffpairibias.t2 gnd 0.086748f
C414 diffpairibias.n17 gnd 0.052262f
C415 diffpairibias.t16 gnd 0.086748f
C416 diffpairibias.n18 gnd 0.052262f
C417 diffpairibias.t4 gnd 0.086748f
C418 diffpairibias.n19 gnd 0.052262f
C419 diffpairibias.t18 gnd 0.086748f
C420 diffpairibias.n20 gnd 0.052262f
C421 diffpairibias.t8 gnd 0.086748f
C422 diffpairibias.n21 gnd 0.061849f
C423 diffpairibias.n22 gnd 0.233513f
C424 diffpairibias.t20 gnd 0.08996f
C425 diffpairibias.n23 gnd 0.051747f
C426 diffpairibias.t26 gnd 0.08996f
C427 diffpairibias.n24 gnd 0.051736f
C428 diffpairibias.t22 gnd 0.08996f
C429 diffpairibias.n25 gnd 0.051736f
C430 diffpairibias.t21 gnd 0.08996f
C431 diffpairibias.n26 gnd 0.051736f
C432 diffpairibias.t24 gnd 0.08996f
C433 diffpairibias.n27 gnd 0.04729f
C434 diffpairibias.n28 gnd 0.047711f
C435 minus.n0 gnd 0.031253f
C436 minus.n1 gnd 0.007092f
C437 minus.n2 gnd 0.031253f
C438 minus.n3 gnd 0.007092f
C439 minus.n4 gnd 0.031253f
C440 minus.n5 gnd 0.007092f
C441 minus.n6 gnd 0.031253f
C442 minus.n7 gnd 0.007092f
C443 minus.n8 gnd 0.031253f
C444 minus.n9 gnd 0.007092f
C445 minus.t8 gnd 0.458091f
C446 minus.t7 gnd 0.442045f
C447 minus.n10 gnd 0.202766f
C448 minus.n11 gnd 0.181989f
C449 minus.n12 gnd 0.134546f
C450 minus.n13 gnd 0.031253f
C451 minus.t11 gnd 0.442045f
C452 minus.n14 gnd 0.196371f
C453 minus.n15 gnd 0.007092f
C454 minus.t10 gnd 0.442045f
C455 minus.n16 gnd 0.196371f
C456 minus.n17 gnd 0.031253f
C457 minus.n18 gnd 0.031253f
C458 minus.n19 gnd 0.031253f
C459 minus.t12 gnd 0.442045f
C460 minus.n20 gnd 0.196371f
C461 minus.n21 gnd 0.007092f
C462 minus.t20 gnd 0.442045f
C463 minus.n22 gnd 0.196371f
C464 minus.n23 gnd 0.031253f
C465 minus.n24 gnd 0.031253f
C466 minus.n25 gnd 0.031253f
C467 minus.t18 gnd 0.442045f
C468 minus.n26 gnd 0.196371f
C469 minus.n27 gnd 0.007092f
C470 minus.t25 gnd 0.442045f
C471 minus.n28 gnd 0.196371f
C472 minus.n29 gnd 0.031253f
C473 minus.n30 gnd 0.031253f
C474 minus.n31 gnd 0.031253f
C475 minus.t24 gnd 0.442045f
C476 minus.n32 gnd 0.196371f
C477 minus.n33 gnd 0.007092f
C478 minus.t14 gnd 0.442045f
C479 minus.n34 gnd 0.196371f
C480 minus.n35 gnd 0.031253f
C481 minus.n36 gnd 0.031253f
C482 minus.n37 gnd 0.031253f
C483 minus.t22 gnd 0.442045f
C484 minus.n38 gnd 0.196371f
C485 minus.n39 gnd 0.007092f
C486 minus.t19 gnd 0.442045f
C487 minus.n40 gnd 0.19666f
C488 minus.n41 gnd 0.361941f
C489 minus.n42 gnd 0.031253f
C490 minus.t13 gnd 0.442045f
C491 minus.t15 gnd 0.442045f
C492 minus.n43 gnd 0.031253f
C493 minus.t5 gnd 0.442045f
C494 minus.n44 gnd 0.196371f
C495 minus.n45 gnd 0.031253f
C496 minus.t6 gnd 0.442045f
C497 minus.t26 gnd 0.442045f
C498 minus.n46 gnd 0.196371f
C499 minus.n47 gnd 0.031253f
C500 minus.t21 gnd 0.442045f
C501 minus.t23 gnd 0.442045f
C502 minus.n48 gnd 0.196371f
C503 minus.n49 gnd 0.031253f
C504 minus.t16 gnd 0.442045f
C505 minus.t17 gnd 0.442045f
C506 minus.n50 gnd 0.196371f
C507 minus.n51 gnd 0.031253f
C508 minus.t9 gnd 0.442045f
C509 minus.t27 gnd 0.442045f
C510 minus.n52 gnd 0.202766f
C511 minus.t28 gnd 0.458091f
C512 minus.n53 gnd 0.181989f
C513 minus.n54 gnd 0.134546f
C514 minus.n55 gnd 0.007092f
C515 minus.n56 gnd 0.196371f
C516 minus.n57 gnd 0.007092f
C517 minus.n58 gnd 0.031253f
C518 minus.n59 gnd 0.031253f
C519 minus.n60 gnd 0.031253f
C520 minus.n61 gnd 0.007092f
C521 minus.n62 gnd 0.196371f
C522 minus.n63 gnd 0.007092f
C523 minus.n64 gnd 0.031253f
C524 minus.n65 gnd 0.031253f
C525 minus.n66 gnd 0.031253f
C526 minus.n67 gnd 0.007092f
C527 minus.n68 gnd 0.196371f
C528 minus.n69 gnd 0.007092f
C529 minus.n70 gnd 0.031253f
C530 minus.n71 gnd 0.031253f
C531 minus.n72 gnd 0.031253f
C532 minus.n73 gnd 0.007092f
C533 minus.n74 gnd 0.196371f
C534 minus.n75 gnd 0.007092f
C535 minus.n76 gnd 0.031253f
C536 minus.n77 gnd 0.031253f
C537 minus.n78 gnd 0.031253f
C538 minus.n79 gnd 0.007092f
C539 minus.n80 gnd 0.196371f
C540 minus.n81 gnd 0.007092f
C541 minus.n82 gnd 0.19666f
C542 minus.n83 gnd 1.04701f
C543 minus.n84 gnd 1.56003f
C544 minus.t1 gnd 0.009634f
C545 minus.t0 gnd 0.009634f
C546 minus.n85 gnd 0.03168f
C547 minus.t4 gnd 0.009634f
C548 minus.t3 gnd 0.009634f
C549 minus.n86 gnd 0.031246f
C550 minus.n87 gnd 0.266671f
C551 minus.t2 gnd 0.053624f
C552 minus.n88 gnd 0.14552f
C553 minus.n89 gnd 2.31716f
C554 a_n1808_13878.t17 gnd 0.185195f
C555 a_n1808_13878.t15 gnd 0.185195f
C556 a_n1808_13878.t19 gnd 0.185195f
C557 a_n1808_13878.n0 gnd 1.46067f
C558 a_n1808_13878.t8 gnd 0.185195f
C559 a_n1808_13878.t13 gnd 0.185195f
C560 a_n1808_13878.n1 gnd 1.45825f
C561 a_n1808_13878.n2 gnd 1.31079f
C562 a_n1808_13878.t10 gnd 0.185195f
C563 a_n1808_13878.t12 gnd 0.185195f
C564 a_n1808_13878.n3 gnd 1.4598f
C565 a_n1808_13878.t16 gnd 0.185195f
C566 a_n1808_13878.t11 gnd 0.185195f
C567 a_n1808_13878.n4 gnd 1.45825f
C568 a_n1808_13878.n5 gnd 2.03762f
C569 a_n1808_13878.t14 gnd 0.185195f
C570 a_n1808_13878.t9 gnd 0.185195f
C571 a_n1808_13878.n6 gnd 1.45825f
C572 a_n1808_13878.n7 gnd 3.69301f
C573 a_n1808_13878.t1 gnd 1.73408f
C574 a_n1808_13878.t4 gnd 0.185195f
C575 a_n1808_13878.t5 gnd 0.185195f
C576 a_n1808_13878.n8 gnd 1.30452f
C577 a_n1808_13878.n9 gnd 1.4576f
C578 a_n1808_13878.t0 gnd 1.73062f
C579 a_n1808_13878.n10 gnd 0.733487f
C580 a_n1808_13878.t3 gnd 1.73062f
C581 a_n1808_13878.n11 gnd 0.733487f
C582 a_n1808_13878.t6 gnd 0.185195f
C583 a_n1808_13878.t7 gnd 0.185195f
C584 a_n1808_13878.n12 gnd 1.30452f
C585 a_n1808_13878.n13 gnd 0.74059f
C586 a_n1808_13878.t2 gnd 1.73062f
C587 a_n1808_13878.n14 gnd 1.7272f
C588 a_n1808_13878.n15 gnd 2.51438f
C589 a_n1808_13878.n16 gnd 1.80025f
C590 a_n1808_13878.n17 gnd 1.45826f
C591 a_n1808_13878.t18 gnd 0.185195f
C592 a_n2408_n452.n0 gnd 3.99939f
C593 a_n2408_n452.n1 gnd 2.94086f
C594 a_n2408_n452.n2 gnd 3.93642f
C595 a_n2408_n452.n3 gnd 0.830148f
C596 a_n2408_n452.n4 gnd 0.83015f
C597 a_n2408_n452.n5 gnd 0.532573f
C598 a_n2408_n452.n6 gnd 0.207439f
C599 a_n2408_n452.n7 gnd 0.152783f
C600 a_n2408_n452.n8 gnd 0.240126f
C601 a_n2408_n452.n9 gnd 0.18547f
C602 a_n2408_n452.n10 gnd 0.207439f
C603 a_n2408_n452.n11 gnd 0.152783f
C604 a_n2408_n452.n12 gnd 0.587229f
C605 a_n2408_n452.n13 gnd 0.437659f
C606 a_n2408_n452.n14 gnd 0.218625f
C607 a_n2408_n452.n15 gnd 0.49859f
C608 a_n2408_n452.n16 gnd 0.286021f
C609 a_n2408_n452.n17 gnd 0.443934f
C610 a_n2408_n452.n18 gnd 0.218625f
C611 a_n2408_n452.n19 gnd 0.740623f
C612 a_n2408_n452.n20 gnd 0.286021f
C613 a_n2408_n452.n21 gnd 0.647141f
C614 a_n2408_n452.n22 gnd 0.286021f
C615 a_n2408_n452.n23 gnd 0.49859f
C616 a_n2408_n452.n24 gnd 0.67269f
C617 a_n2408_n452.n25 gnd 0.218625f
C618 a_n2408_n452.n26 gnd 0.286021f
C619 a_n2408_n452.n27 gnd 3.36354f
C620 a_n2408_n452.n28 gnd 0.286021f
C621 a_n2408_n452.n29 gnd 1.79992f
C622 a_n2408_n452.n30 gnd 1.93948f
C623 a_n2408_n452.n31 gnd 0.008464f
C624 a_n2408_n452.n33 gnd 1.35508f
C625 a_n2408_n452.n34 gnd 0.289215f
C626 a_n2408_n452.n35 gnd 0.004526f
C627 a_n2408_n452.n36 gnd 0.008464f
C628 a_n2408_n452.n38 gnd 0.289215f
C629 a_n2408_n452.n39 gnd 0.008464f
C630 a_n2408_n452.n41 gnd 0.289215f
C631 a_n2408_n452.n42 gnd 0.008464f
C632 a_n2408_n452.n43 gnd 0.288804f
C633 a_n2408_n452.n44 gnd 0.008464f
C634 a_n2408_n452.n45 gnd 0.288804f
C635 a_n2408_n452.n46 gnd 0.008464f
C636 a_n2408_n452.n47 gnd 0.288804f
C637 a_n2408_n452.n48 gnd 0.008464f
C638 a_n2408_n452.n49 gnd 0.288804f
C639 a_n2408_n452.n50 gnd 0.310121f
C640 a_n2408_n452.t22 gnd 0.151641f
C641 a_n2408_n452.t26 gnd 1.41989f
C642 a_n2408_n452.t37 gnd 0.70536f
C643 a_n2408_n452.n51 gnd 0.310121f
C644 a_n2408_n452.t29 gnd 0.70536f
C645 a_n2408_n452.t21 gnd 0.70536f
C646 a_n2408_n452.t56 gnd 0.70536f
C647 a_n2408_n452.n52 gnd 0.310121f
C648 a_n2408_n452.t64 gnd 0.70536f
C649 a_n2408_n452.t70 gnd 0.70536f
C650 a_n2408_n452.t33 gnd 0.720216f
C651 a_n2408_n452.t35 gnd 0.70536f
C652 a_n2408_n452.t41 gnd 0.70536f
C653 a_n2408_n452.t23 gnd 0.70536f
C654 a_n2408_n452.t39 gnd 0.70536f
C655 a_n2408_n452.t27 gnd 0.720216f
C656 a_n2408_n452.t74 gnd 0.720216f
C657 a_n2408_n452.t57 gnd 0.70536f
C658 a_n2408_n452.t61 gnd 0.70536f
C659 a_n2408_n452.t51 gnd 0.70536f
C660 a_n2408_n452.n53 gnd 0.310121f
C661 a_n2408_n452.t66 gnd 0.70536f
C662 a_n2408_n452.t72 gnd 0.717022f
C663 a_n2408_n452.n54 gnd 0.312771f
C664 a_n2408_n452.n55 gnd 0.306183f
C665 a_n2408_n452.n56 gnd 0.31277f
C666 a_n2408_n452.n57 gnd 0.312771f
C667 a_n2408_n452.t2 gnd 0.117943f
C668 a_n2408_n452.t7 gnd 0.117943f
C669 a_n2408_n452.n58 gnd 1.0445f
C670 a_n2408_n452.t44 gnd 0.117943f
C671 a_n2408_n452.t45 gnd 0.117943f
C672 a_n2408_n452.n59 gnd 1.04218f
C673 a_n2408_n452.t4 gnd 0.117943f
C674 a_n2408_n452.t17 gnd 0.117943f
C675 a_n2408_n452.n60 gnd 1.04218f
C676 a_n2408_n452.t6 gnd 0.117943f
C677 a_n2408_n452.t18 gnd 0.117943f
C678 a_n2408_n452.n61 gnd 1.0445f
C679 a_n2408_n452.t0 gnd 0.117943f
C680 a_n2408_n452.t3 gnd 0.117943f
C681 a_n2408_n452.n62 gnd 1.04218f
C682 a_n2408_n452.t47 gnd 0.117943f
C683 a_n2408_n452.t16 gnd 0.117943f
C684 a_n2408_n452.n63 gnd 1.04218f
C685 a_n2408_n452.t8 gnd 0.117943f
C686 a_n2408_n452.t43 gnd 0.117943f
C687 a_n2408_n452.n64 gnd 1.04218f
C688 a_n2408_n452.t10 gnd 0.117943f
C689 a_n2408_n452.t12 gnd 0.117943f
C690 a_n2408_n452.n65 gnd 1.04218f
C691 a_n2408_n452.t9 gnd 0.117943f
C692 a_n2408_n452.t14 gnd 0.117943f
C693 a_n2408_n452.n66 gnd 1.04218f
C694 a_n2408_n452.t13 gnd 0.117943f
C695 a_n2408_n452.t15 gnd 0.117943f
C696 a_n2408_n452.n67 gnd 1.0445f
C697 a_n2408_n452.t46 gnd 0.117943f
C698 a_n2408_n452.t11 gnd 0.117943f
C699 a_n2408_n452.n68 gnd 1.04218f
C700 a_n2408_n452.t5 gnd 0.117943f
C701 a_n2408_n452.t1 gnd 0.117943f
C702 a_n2408_n452.n69 gnd 1.04218f
C703 a_n2408_n452.n70 gnd 0.310121f
C704 a_n2408_n452.n71 gnd 0.31277f
C705 a_n2408_n452.t28 gnd 1.41989f
C706 a_n2408_n452.t24 gnd 0.151641f
C707 a_n2408_n452.t40 gnd 0.151641f
C708 a_n2408_n452.n72 gnd 1.06816f
C709 a_n2408_n452.t36 gnd 0.151641f
C710 a_n2408_n452.t42 gnd 0.151641f
C711 a_n2408_n452.n73 gnd 1.06816f
C712 a_n2408_n452.t34 gnd 1.41706f
C713 a_n2408_n452.n74 gnd 1.1588f
C714 a_n2408_n452.n75 gnd 0.796711f
C715 a_n2408_n452.t55 gnd 0.70536f
C716 a_n2408_n452.t65 gnd 0.70536f
C717 a_n2408_n452.t75 gnd 0.70536f
C718 a_n2408_n452.n76 gnd 0.310121f
C719 a_n2408_n452.t67 gnd 0.70536f
C720 a_n2408_n452.t52 gnd 0.70536f
C721 a_n2408_n452.t53 gnd 0.70536f
C722 a_n2408_n452.n77 gnd 0.310121f
C723 a_n2408_n452.t71 gnd 0.70536f
C724 a_n2408_n452.t60 gnd 0.70536f
C725 a_n2408_n452.t59 gnd 0.70536f
C726 a_n2408_n452.n78 gnd 0.310121f
C727 a_n2408_n452.t63 gnd 0.70536f
C728 a_n2408_n452.t54 gnd 0.70536f
C729 a_n2408_n452.t48 gnd 0.70536f
C730 a_n2408_n452.n79 gnd 0.310121f
C731 a_n2408_n452.t68 gnd 0.717179f
C732 a_n2408_n452.n80 gnd 0.306183f
C733 a_n2408_n452.n81 gnd 0.300622f
C734 a_n2408_n452.t73 gnd 0.717179f
C735 a_n2408_n452.n82 gnd 0.306183f
C736 a_n2408_n452.n83 gnd 0.300622f
C737 a_n2408_n452.t62 gnd 0.717179f
C738 a_n2408_n452.n84 gnd 0.306183f
C739 a_n2408_n452.n85 gnd 0.300622f
C740 a_n2408_n452.t58 gnd 0.717179f
C741 a_n2408_n452.n86 gnd 0.306183f
C742 a_n2408_n452.n87 gnd 0.300622f
C743 a_n2408_n452.n88 gnd 1.0188f
C744 a_n2408_n452.t69 gnd 0.720216f
C745 a_n2408_n452.n89 gnd 0.31277f
C746 a_n2408_n452.t49 gnd 0.70536f
C747 a_n2408_n452.n90 gnd 0.306183f
C748 a_n2408_n452.n91 gnd 0.312771f
C749 a_n2408_n452.t50 gnd 0.717022f
C750 a_n2408_n452.t25 gnd 0.720216f
C751 a_n2408_n452.n92 gnd 0.31277f
C752 a_n2408_n452.t19 gnd 0.70536f
C753 a_n2408_n452.n93 gnd 0.306183f
C754 a_n2408_n452.n94 gnd 0.312771f
C755 a_n2408_n452.t31 gnd 0.717022f
C756 a_n2408_n452.n95 gnd 1.1461f
C757 a_n2408_n452.t32 gnd 1.41706f
C758 a_n2408_n452.t38 gnd 0.151641f
C759 a_n2408_n452.t30 gnd 0.151641f
C760 a_n2408_n452.n96 gnd 1.06816f
C761 a_n2408_n452.n97 gnd 1.19351f
C762 a_n2408_n452.n98 gnd 1.06816f
C763 a_n2408_n452.t20 gnd 0.151641f
C764 a_n3827_n3924.t39 gnd 0.097472f
C765 a_n3827_n3924.t45 gnd 0.097472f
C766 a_n3827_n3924.n0 gnd 0.796067f
C767 a_n3827_n3924.n1 gnd 0.362017f
C768 a_n3827_n3924.t48 gnd 1.01304f
C769 a_n3827_n3924.n2 gnd 0.911283f
C770 a_n3827_n3924.t28 gnd 0.097472f
C771 a_n3827_n3924.t46 gnd 0.097472f
C772 a_n3827_n3924.n3 gnd 0.796069f
C773 a_n3827_n3924.n4 gnd 0.362016f
C774 a_n3827_n3924.t42 gnd 0.097472f
C775 a_n3827_n3924.t44 gnd 0.097472f
C776 a_n3827_n3924.n5 gnd 0.796069f
C777 a_n3827_n3924.n6 gnd 0.362016f
C778 a_n3827_n3924.t47 gnd 0.097472f
C779 a_n3827_n3924.t49 gnd 0.097472f
C780 a_n3827_n3924.n7 gnd 0.796069f
C781 a_n3827_n3924.n8 gnd 0.362016f
C782 a_n3827_n3924.t31 gnd 0.097472f
C783 a_n3827_n3924.t29 gnd 0.097472f
C784 a_n3827_n3924.n9 gnd 0.796069f
C785 a_n3827_n3924.n10 gnd 0.362016f
C786 a_n3827_n3924.t37 gnd 0.097472f
C787 a_n3827_n3924.t30 gnd 0.097472f
C788 a_n3827_n3924.n11 gnd 0.796069f
C789 a_n3827_n3924.n12 gnd 0.362016f
C790 a_n3827_n3924.t36 gnd 1.01304f
C791 a_n3827_n3924.n13 gnd 0.363396f
C792 a_n3827_n3924.t18 gnd 1.01304f
C793 a_n3827_n3924.n14 gnd 0.363396f
C794 a_n3827_n3924.t12 gnd 0.097472f
C795 a_n3827_n3924.t15 gnd 0.097472f
C796 a_n3827_n3924.n15 gnd 0.796069f
C797 a_n3827_n3924.n16 gnd 0.362016f
C798 a_n3827_n3924.t1 gnd 0.097472f
C799 a_n3827_n3924.t27 gnd 0.097472f
C800 a_n3827_n3924.n17 gnd 0.796069f
C801 a_n3827_n3924.n18 gnd 0.362016f
C802 a_n3827_n3924.t16 gnd 0.097472f
C803 a_n3827_n3924.t5 gnd 0.097472f
C804 a_n3827_n3924.n19 gnd 0.796069f
C805 a_n3827_n3924.n20 gnd 0.362016f
C806 a_n3827_n3924.t13 gnd 0.097472f
C807 a_n3827_n3924.t9 gnd 0.097472f
C808 a_n3827_n3924.n21 gnd 0.796069f
C809 a_n3827_n3924.n22 gnd 0.362016f
C810 a_n3827_n3924.t24 gnd 0.097472f
C811 a_n3827_n3924.t10 gnd 0.097472f
C812 a_n3827_n3924.n23 gnd 0.796069f
C813 a_n3827_n3924.n24 gnd 0.362016f
C814 a_n3827_n3924.t8 gnd 1.01304f
C815 a_n3827_n3924.n25 gnd 0.911279f
C816 a_n3827_n3924.t34 gnd 0.097472f
C817 a_n3827_n3924.t40 gnd 0.097472f
C818 a_n3827_n3924.n26 gnd 0.796067f
C819 a_n3827_n3924.n27 gnd 0.362017f
C820 a_n3827_n3924.t35 gnd 1.01304f
C821 a_n3827_n3924.n28 gnd 0.592532f
C822 a_n3827_n3924.n29 gnd 0.914318f
C823 a_n3827_n3924.t55 gnd 1.26048f
C824 a_n3827_n3924.t14 gnd 1.25868f
C825 a_n3827_n3924.n30 gnd 1.28533f
C826 a_n3827_n3924.n31 gnd 0.479144f
C827 a_n3827_n3924.t54 gnd 1.25868f
C828 a_n3827_n3924.n32 gnd 0.725754f
C829 a_n3827_n3924.t11 gnd 1.25868f
C830 a_n3827_n3924.n33 gnd 0.886511f
C831 a_n3827_n3924.t52 gnd 1.25868f
C832 a_n3827_n3924.n34 gnd 0.886511f
C833 a_n3827_n3924.t57 gnd 1.25868f
C834 a_n3827_n3924.n35 gnd 0.886511f
C835 a_n3827_n3924.t17 gnd 1.25868f
C836 a_n3827_n3924.n36 gnd 0.886511f
C837 a_n3827_n3924.t53 gnd 1.25868f
C838 a_n3827_n3924.n37 gnd 0.886511f
C839 a_n3827_n3924.t23 gnd 1.25868f
C840 a_n3827_n3924.n38 gnd 0.654629f
C841 a_n3827_n3924.t22 gnd 1.26084f
C842 a_n3827_n3924.n39 gnd 1.47707f
C843 a_n3827_n3924.n40 gnd 0.914318f
C844 a_n3827_n3924.t21 gnd 1.01304f
C845 a_n3827_n3924.n41 gnd 0.592532f
C846 a_n3827_n3924.t3 gnd 0.097472f
C847 a_n3827_n3924.t6 gnd 0.097472f
C848 a_n3827_n3924.n42 gnd 0.796067f
C849 a_n3827_n3924.n43 gnd 0.362017f
C850 a_n3827_n3924.t19 gnd 0.097472f
C851 a_n3827_n3924.t0 gnd 0.097472f
C852 a_n3827_n3924.n44 gnd 0.796067f
C853 a_n3827_n3924.n45 gnd 0.362017f
C854 a_n3827_n3924.t20 gnd 0.097472f
C855 a_n3827_n3924.t56 gnd 0.097472f
C856 a_n3827_n3924.n46 gnd 0.796067f
C857 a_n3827_n3924.n47 gnd 0.362017f
C858 a_n3827_n3924.t26 gnd 0.097472f
C859 a_n3827_n3924.t4 gnd 0.097472f
C860 a_n3827_n3924.n48 gnd 0.796067f
C861 a_n3827_n3924.n49 gnd 0.362017f
C862 a_n3827_n3924.t7 gnd 0.097472f
C863 a_n3827_n3924.t25 gnd 0.097472f
C864 a_n3827_n3924.n50 gnd 0.796067f
C865 a_n3827_n3924.n51 gnd 0.362017f
C866 a_n3827_n3924.t2 gnd 1.01304f
C867 a_n3827_n3924.n52 gnd 0.3634f
C868 a_n3827_n3924.t41 gnd 1.01304f
C869 a_n3827_n3924.n53 gnd 0.3634f
C870 a_n3827_n3924.t38 gnd 0.097472f
C871 a_n3827_n3924.t43 gnd 0.097472f
C872 a_n3827_n3924.n54 gnd 0.796067f
C873 a_n3827_n3924.n55 gnd 0.362017f
C874 a_n3827_n3924.t33 gnd 0.097472f
C875 a_n3827_n3924.t32 gnd 0.097472f
C876 a_n3827_n3924.n56 gnd 0.796067f
C877 a_n3827_n3924.n57 gnd 0.362017f
C878 a_n3827_n3924.n58 gnd 0.36202f
C879 a_n3827_n3924.t50 gnd 0.097472f
C880 a_n3827_n3924.n59 gnd 0.796064f
C881 a_n3827_n3924.t51 gnd 0.097472f
C882 plus.n0 gnd 0.022995f
C883 plus.t21 gnd 0.325242f
C884 plus.n1 gnd 0.022995f
C885 plus.t22 gnd 0.325242f
C886 plus.t16 gnd 0.325242f
C887 plus.n2 gnd 0.144483f
C888 plus.n3 gnd 0.022995f
C889 plus.t17 gnd 0.325242f
C890 plus.t11 gnd 0.325242f
C891 plus.n4 gnd 0.144483f
C892 plus.n5 gnd 0.022995f
C893 plus.t5 gnd 0.325242f
C894 plus.t6 gnd 0.325242f
C895 plus.n6 gnd 0.144483f
C896 plus.n7 gnd 0.022995f
C897 plus.t23 gnd 0.325242f
C898 plus.t24 gnd 0.325242f
C899 plus.n8 gnd 0.144483f
C900 plus.n9 gnd 0.022995f
C901 plus.t18 gnd 0.325242f
C902 plus.t13 gnd 0.325242f
C903 plus.n10 gnd 0.149189f
C904 plus.t15 gnd 0.337048f
C905 plus.n11 gnd 0.133901f
C906 plus.n12 gnd 0.098995f
C907 plus.n13 gnd 0.005218f
C908 plus.n14 gnd 0.144483f
C909 plus.n15 gnd 0.005218f
C910 plus.n16 gnd 0.022995f
C911 plus.n17 gnd 0.022995f
C912 plus.n18 gnd 0.022995f
C913 plus.n19 gnd 0.005218f
C914 plus.n20 gnd 0.144483f
C915 plus.n21 gnd 0.005218f
C916 plus.n22 gnd 0.022995f
C917 plus.n23 gnd 0.022995f
C918 plus.n24 gnd 0.022995f
C919 plus.n25 gnd 0.005218f
C920 plus.n26 gnd 0.144483f
C921 plus.n27 gnd 0.005218f
C922 plus.n28 gnd 0.022995f
C923 plus.n29 gnd 0.022995f
C924 plus.n30 gnd 0.022995f
C925 plus.n31 gnd 0.005218f
C926 plus.n32 gnd 0.144483f
C927 plus.n33 gnd 0.005218f
C928 plus.n34 gnd 0.022995f
C929 plus.n35 gnd 0.022995f
C930 plus.n36 gnd 0.022995f
C931 plus.n37 gnd 0.005218f
C932 plus.n38 gnd 0.144483f
C933 plus.n39 gnd 0.005218f
C934 plus.n40 gnd 0.144696f
C935 plus.n41 gnd 0.260382f
C936 plus.n42 gnd 0.022995f
C937 plus.n43 gnd 0.005218f
C938 plus.t10 gnd 0.325242f
C939 plus.n44 gnd 0.022995f
C940 plus.n45 gnd 0.005218f
C941 plus.t12 gnd 0.325242f
C942 plus.n46 gnd 0.022995f
C943 plus.n47 gnd 0.005218f
C944 plus.t7 gnd 0.325242f
C945 plus.n48 gnd 0.022995f
C946 plus.n49 gnd 0.005218f
C947 plus.t27 gnd 0.325242f
C948 plus.n50 gnd 0.022995f
C949 plus.n51 gnd 0.005218f
C950 plus.t26 gnd 0.325242f
C951 plus.t20 gnd 0.337048f
C952 plus.t19 gnd 0.325242f
C953 plus.n52 gnd 0.149189f
C954 plus.n53 gnd 0.133901f
C955 plus.n54 gnd 0.098995f
C956 plus.n55 gnd 0.022995f
C957 plus.n56 gnd 0.144483f
C958 plus.n57 gnd 0.005218f
C959 plus.t25 gnd 0.325242f
C960 plus.n58 gnd 0.144483f
C961 plus.n59 gnd 0.022995f
C962 plus.n60 gnd 0.022995f
C963 plus.n61 gnd 0.022995f
C964 plus.n62 gnd 0.144483f
C965 plus.n63 gnd 0.005218f
C966 plus.t9 gnd 0.325242f
C967 plus.n64 gnd 0.144483f
C968 plus.n65 gnd 0.022995f
C969 plus.n66 gnd 0.022995f
C970 plus.n67 gnd 0.022995f
C971 plus.n68 gnd 0.144483f
C972 plus.n69 gnd 0.005218f
C973 plus.t14 gnd 0.325242f
C974 plus.n70 gnd 0.144483f
C975 plus.n71 gnd 0.022995f
C976 plus.n72 gnd 0.022995f
C977 plus.n73 gnd 0.022995f
C978 plus.n74 gnd 0.144483f
C979 plus.n75 gnd 0.005218f
C980 plus.t28 gnd 0.325242f
C981 plus.n76 gnd 0.144483f
C982 plus.n77 gnd 0.022995f
C983 plus.n78 gnd 0.022995f
C984 plus.n79 gnd 0.022995f
C985 plus.n80 gnd 0.144483f
C986 plus.n81 gnd 0.005218f
C987 plus.t8 gnd 0.325242f
C988 plus.n82 gnd 0.144696f
C989 plus.n83 gnd 0.761135f
C990 plus.n84 gnd 1.13871f
C991 plus.t2 gnd 0.039696f
C992 plus.t3 gnd 0.007089f
C993 plus.t1 gnd 0.007089f
C994 plus.n85 gnd 0.02299f
C995 plus.n86 gnd 0.178472f
C996 plus.t4 gnd 0.007089f
C997 plus.t0 gnd 0.007089f
C998 plus.n87 gnd 0.02299f
C999 plus.n88 gnd 0.133965f
C1000 plus.n89 gnd 3.14792f
C1001 commonsourceibias.n0 gnd 0.012818f
C1002 commonsourceibias.t104 gnd 0.19409f
C1003 commonsourceibias.t181 gnd 0.179464f
C1004 commonsourceibias.n1 gnd 0.00935f
C1005 commonsourceibias.n2 gnd 0.009606f
C1006 commonsourceibias.t124 gnd 0.179464f
C1007 commonsourceibias.n3 gnd 0.012358f
C1008 commonsourceibias.n4 gnd 0.009606f
C1009 commonsourceibias.t197 gnd 0.179464f
C1010 commonsourceibias.n5 gnd 0.071606f
C1011 commonsourceibias.t142 gnd 0.179464f
C1012 commonsourceibias.n6 gnd 0.009057f
C1013 commonsourceibias.n7 gnd 0.009606f
C1014 commonsourceibias.t101 gnd 0.179464f
C1015 commonsourceibias.n8 gnd 0.012175f
C1016 commonsourceibias.n9 gnd 0.009606f
C1017 commonsourceibias.t156 gnd 0.179464f
C1018 commonsourceibias.n10 gnd 0.071606f
C1019 commonsourceibias.t143 gnd 0.179464f
C1020 commonsourceibias.n11 gnd 0.008798f
C1021 commonsourceibias.n12 gnd 0.009606f
C1022 commonsourceibias.t193 gnd 0.179464f
C1023 commonsourceibias.n13 gnd 0.01197f
C1024 commonsourceibias.n14 gnd 0.012818f
C1025 commonsourceibias.t50 gnd 0.19409f
C1026 commonsourceibias.t40 gnd 0.179464f
C1027 commonsourceibias.n15 gnd 0.00935f
C1028 commonsourceibias.n16 gnd 0.009606f
C1029 commonsourceibias.t0 gnd 0.179464f
C1030 commonsourceibias.n17 gnd 0.012358f
C1031 commonsourceibias.n18 gnd 0.009606f
C1032 commonsourceibias.t74 gnd 0.179464f
C1033 commonsourceibias.n19 gnd 0.071606f
C1034 commonsourceibias.t34 gnd 0.179464f
C1035 commonsourceibias.n20 gnd 0.009057f
C1036 commonsourceibias.n21 gnd 0.009606f
C1037 commonsourceibias.t6 gnd 0.179464f
C1038 commonsourceibias.n22 gnd 0.012175f
C1039 commonsourceibias.n23 gnd 0.009606f
C1040 commonsourceibias.t12 gnd 0.179464f
C1041 commonsourceibias.n24 gnd 0.071606f
C1042 commonsourceibias.t32 gnd 0.179464f
C1043 commonsourceibias.n25 gnd 0.008798f
C1044 commonsourceibias.n26 gnd 0.009606f
C1045 commonsourceibias.t76 gnd 0.179464f
C1046 commonsourceibias.n27 gnd 0.01197f
C1047 commonsourceibias.n28 gnd 0.009606f
C1048 commonsourceibias.t26 gnd 0.179464f
C1049 commonsourceibias.n29 gnd 0.071606f
C1050 commonsourceibias.t64 gnd 0.179464f
C1051 commonsourceibias.n30 gnd 0.008572f
C1052 commonsourceibias.n31 gnd 0.009606f
C1053 commonsourceibias.t14 gnd 0.179464f
C1054 commonsourceibias.n32 gnd 0.011742f
C1055 commonsourceibias.n33 gnd 0.009606f
C1056 commonsourceibias.t36 gnd 0.179464f
C1057 commonsourceibias.n34 gnd 0.071606f
C1058 commonsourceibias.t52 gnd 0.179464f
C1059 commonsourceibias.n35 gnd 0.008375f
C1060 commonsourceibias.n36 gnd 0.009606f
C1061 commonsourceibias.t46 gnd 0.179464f
C1062 commonsourceibias.n37 gnd 0.011489f
C1063 commonsourceibias.n38 gnd 0.009606f
C1064 commonsourceibias.t38 gnd 0.179464f
C1065 commonsourceibias.n39 gnd 0.071606f
C1066 commonsourceibias.t2 gnd 0.179464f
C1067 commonsourceibias.n40 gnd 0.008208f
C1068 commonsourceibias.n41 gnd 0.009606f
C1069 commonsourceibias.t70 gnd 0.179464f
C1070 commonsourceibias.n42 gnd 0.011208f
C1071 commonsourceibias.t8 gnd 0.199531f
C1072 commonsourceibias.t66 gnd 0.179464f
C1073 commonsourceibias.n43 gnd 0.078223f
C1074 commonsourceibias.n44 gnd 0.08584f
C1075 commonsourceibias.n45 gnd 0.039831f
C1076 commonsourceibias.n46 gnd 0.009606f
C1077 commonsourceibias.n47 gnd 0.00935f
C1078 commonsourceibias.n48 gnd 0.013398f
C1079 commonsourceibias.n49 gnd 0.071606f
C1080 commonsourceibias.n50 gnd 0.013389f
C1081 commonsourceibias.n51 gnd 0.009606f
C1082 commonsourceibias.n52 gnd 0.009606f
C1083 commonsourceibias.n53 gnd 0.009606f
C1084 commonsourceibias.n54 gnd 0.012358f
C1085 commonsourceibias.n55 gnd 0.071606f
C1086 commonsourceibias.n56 gnd 0.012648f
C1087 commonsourceibias.n57 gnd 0.012289f
C1088 commonsourceibias.n58 gnd 0.009606f
C1089 commonsourceibias.n59 gnd 0.009606f
C1090 commonsourceibias.n60 gnd 0.009606f
C1091 commonsourceibias.n61 gnd 0.009057f
C1092 commonsourceibias.n62 gnd 0.01341f
C1093 commonsourceibias.n63 gnd 0.071606f
C1094 commonsourceibias.n64 gnd 0.013406f
C1095 commonsourceibias.n65 gnd 0.009606f
C1096 commonsourceibias.n66 gnd 0.009606f
C1097 commonsourceibias.n67 gnd 0.009606f
C1098 commonsourceibias.n68 gnd 0.012175f
C1099 commonsourceibias.n69 gnd 0.071606f
C1100 commonsourceibias.n70 gnd 0.012558f
C1101 commonsourceibias.n71 gnd 0.012378f
C1102 commonsourceibias.n72 gnd 0.009606f
C1103 commonsourceibias.n73 gnd 0.009606f
C1104 commonsourceibias.n74 gnd 0.009606f
C1105 commonsourceibias.n75 gnd 0.008798f
C1106 commonsourceibias.n76 gnd 0.013416f
C1107 commonsourceibias.n77 gnd 0.071606f
C1108 commonsourceibias.n78 gnd 0.013414f
C1109 commonsourceibias.n79 gnd 0.009606f
C1110 commonsourceibias.n80 gnd 0.009606f
C1111 commonsourceibias.n81 gnd 0.009606f
C1112 commonsourceibias.n82 gnd 0.01197f
C1113 commonsourceibias.n83 gnd 0.071606f
C1114 commonsourceibias.n84 gnd 0.012468f
C1115 commonsourceibias.n85 gnd 0.012468f
C1116 commonsourceibias.n86 gnd 0.009606f
C1117 commonsourceibias.n87 gnd 0.009606f
C1118 commonsourceibias.n88 gnd 0.009606f
C1119 commonsourceibias.n89 gnd 0.008572f
C1120 commonsourceibias.n90 gnd 0.013414f
C1121 commonsourceibias.n91 gnd 0.071606f
C1122 commonsourceibias.n92 gnd 0.013416f
C1123 commonsourceibias.n93 gnd 0.009606f
C1124 commonsourceibias.n94 gnd 0.009606f
C1125 commonsourceibias.n95 gnd 0.009606f
C1126 commonsourceibias.n96 gnd 0.011742f
C1127 commonsourceibias.n97 gnd 0.071606f
C1128 commonsourceibias.n98 gnd 0.012378f
C1129 commonsourceibias.n99 gnd 0.012558f
C1130 commonsourceibias.n100 gnd 0.009606f
C1131 commonsourceibias.n101 gnd 0.009606f
C1132 commonsourceibias.n102 gnd 0.009606f
C1133 commonsourceibias.n103 gnd 0.008375f
C1134 commonsourceibias.n104 gnd 0.013406f
C1135 commonsourceibias.n105 gnd 0.071606f
C1136 commonsourceibias.n106 gnd 0.01341f
C1137 commonsourceibias.n107 gnd 0.009606f
C1138 commonsourceibias.n108 gnd 0.009606f
C1139 commonsourceibias.n109 gnd 0.009606f
C1140 commonsourceibias.n110 gnd 0.011489f
C1141 commonsourceibias.n111 gnd 0.071606f
C1142 commonsourceibias.n112 gnd 0.012289f
C1143 commonsourceibias.n113 gnd 0.012648f
C1144 commonsourceibias.n114 gnd 0.009606f
C1145 commonsourceibias.n115 gnd 0.009606f
C1146 commonsourceibias.n116 gnd 0.009606f
C1147 commonsourceibias.n117 gnd 0.008208f
C1148 commonsourceibias.n118 gnd 0.013389f
C1149 commonsourceibias.n119 gnd 0.071606f
C1150 commonsourceibias.n120 gnd 0.013398f
C1151 commonsourceibias.n121 gnd 0.009606f
C1152 commonsourceibias.n122 gnd 0.009606f
C1153 commonsourceibias.n123 gnd 0.009606f
C1154 commonsourceibias.n124 gnd 0.011208f
C1155 commonsourceibias.n125 gnd 0.071606f
C1156 commonsourceibias.n126 gnd 0.011785f
C1157 commonsourceibias.n127 gnd 0.085921f
C1158 commonsourceibias.n128 gnd 0.095704f
C1159 commonsourceibias.t51 gnd 0.020728f
C1160 commonsourceibias.t41 gnd 0.020728f
C1161 commonsourceibias.n129 gnd 0.183161f
C1162 commonsourceibias.n130 gnd 0.158435f
C1163 commonsourceibias.t1 gnd 0.020728f
C1164 commonsourceibias.t75 gnd 0.020728f
C1165 commonsourceibias.n131 gnd 0.183161f
C1166 commonsourceibias.n132 gnd 0.084133f
C1167 commonsourceibias.t35 gnd 0.020728f
C1168 commonsourceibias.t7 gnd 0.020728f
C1169 commonsourceibias.n133 gnd 0.183161f
C1170 commonsourceibias.n134 gnd 0.084133f
C1171 commonsourceibias.t13 gnd 0.020728f
C1172 commonsourceibias.t33 gnd 0.020728f
C1173 commonsourceibias.n135 gnd 0.183161f
C1174 commonsourceibias.n136 gnd 0.084133f
C1175 commonsourceibias.t77 gnd 0.020728f
C1176 commonsourceibias.t27 gnd 0.020728f
C1177 commonsourceibias.n137 gnd 0.183161f
C1178 commonsourceibias.n138 gnd 0.070289f
C1179 commonsourceibias.t67 gnd 0.020728f
C1180 commonsourceibias.t9 gnd 0.020728f
C1181 commonsourceibias.n139 gnd 0.183774f
C1182 commonsourceibias.t3 gnd 0.020728f
C1183 commonsourceibias.t71 gnd 0.020728f
C1184 commonsourceibias.n140 gnd 0.183161f
C1185 commonsourceibias.n141 gnd 0.170671f
C1186 commonsourceibias.t47 gnd 0.020728f
C1187 commonsourceibias.t39 gnd 0.020728f
C1188 commonsourceibias.n142 gnd 0.183161f
C1189 commonsourceibias.n143 gnd 0.084133f
C1190 commonsourceibias.t37 gnd 0.020728f
C1191 commonsourceibias.t53 gnd 0.020728f
C1192 commonsourceibias.n144 gnd 0.183161f
C1193 commonsourceibias.n145 gnd 0.084133f
C1194 commonsourceibias.t65 gnd 0.020728f
C1195 commonsourceibias.t15 gnd 0.020728f
C1196 commonsourceibias.n146 gnd 0.183161f
C1197 commonsourceibias.n147 gnd 0.070289f
C1198 commonsourceibias.n148 gnd 0.085113f
C1199 commonsourceibias.n149 gnd 0.062168f
C1200 commonsourceibias.t136 gnd 0.179464f
C1201 commonsourceibias.n150 gnd 0.071606f
C1202 commonsourceibias.t119 gnd 0.179464f
C1203 commonsourceibias.n151 gnd 0.071606f
C1204 commonsourceibias.n152 gnd 0.009606f
C1205 commonsourceibias.t155 gnd 0.179464f
C1206 commonsourceibias.n153 gnd 0.071606f
C1207 commonsourceibias.n154 gnd 0.009606f
C1208 commonsourceibias.t140 gnd 0.179464f
C1209 commonsourceibias.n155 gnd 0.071606f
C1210 commonsourceibias.n156 gnd 0.009606f
C1211 commonsourceibias.t109 gnd 0.179464f
C1212 commonsourceibias.n157 gnd 0.008375f
C1213 commonsourceibias.n158 gnd 0.009606f
C1214 commonsourceibias.t182 gnd 0.179464f
C1215 commonsourceibias.n159 gnd 0.011489f
C1216 commonsourceibias.n160 gnd 0.009606f
C1217 commonsourceibias.t166 gnd 0.179464f
C1218 commonsourceibias.n161 gnd 0.071606f
C1219 commonsourceibias.t123 gnd 0.179464f
C1220 commonsourceibias.n162 gnd 0.008208f
C1221 commonsourceibias.n163 gnd 0.009606f
C1222 commonsourceibias.t84 gnd 0.179464f
C1223 commonsourceibias.n164 gnd 0.011208f
C1224 commonsourceibias.t100 gnd 0.199531f
C1225 commonsourceibias.t131 gnd 0.179464f
C1226 commonsourceibias.n165 gnd 0.078223f
C1227 commonsourceibias.n166 gnd 0.08584f
C1228 commonsourceibias.n167 gnd 0.039831f
C1229 commonsourceibias.n168 gnd 0.009606f
C1230 commonsourceibias.n169 gnd 0.00935f
C1231 commonsourceibias.n170 gnd 0.013398f
C1232 commonsourceibias.n171 gnd 0.071606f
C1233 commonsourceibias.n172 gnd 0.013389f
C1234 commonsourceibias.n173 gnd 0.009606f
C1235 commonsourceibias.n174 gnd 0.009606f
C1236 commonsourceibias.n175 gnd 0.009606f
C1237 commonsourceibias.n176 gnd 0.012358f
C1238 commonsourceibias.n177 gnd 0.071606f
C1239 commonsourceibias.n178 gnd 0.012648f
C1240 commonsourceibias.n179 gnd 0.012289f
C1241 commonsourceibias.n180 gnd 0.009606f
C1242 commonsourceibias.n181 gnd 0.009606f
C1243 commonsourceibias.n182 gnd 0.009606f
C1244 commonsourceibias.n183 gnd 0.009057f
C1245 commonsourceibias.n184 gnd 0.01341f
C1246 commonsourceibias.n185 gnd 0.071606f
C1247 commonsourceibias.n186 gnd 0.013406f
C1248 commonsourceibias.n187 gnd 0.009606f
C1249 commonsourceibias.n188 gnd 0.009606f
C1250 commonsourceibias.n189 gnd 0.009606f
C1251 commonsourceibias.n190 gnd 0.012175f
C1252 commonsourceibias.n191 gnd 0.071606f
C1253 commonsourceibias.n192 gnd 0.012558f
C1254 commonsourceibias.n193 gnd 0.012378f
C1255 commonsourceibias.n194 gnd 0.009606f
C1256 commonsourceibias.n195 gnd 0.009606f
C1257 commonsourceibias.n196 gnd 0.011742f
C1258 commonsourceibias.n197 gnd 0.008798f
C1259 commonsourceibias.n198 gnd 0.013416f
C1260 commonsourceibias.n199 gnd 0.009606f
C1261 commonsourceibias.n200 gnd 0.009606f
C1262 commonsourceibias.n201 gnd 0.013414f
C1263 commonsourceibias.n202 gnd 0.008572f
C1264 commonsourceibias.n203 gnd 0.01197f
C1265 commonsourceibias.n204 gnd 0.009606f
C1266 commonsourceibias.n205 gnd 0.008392f
C1267 commonsourceibias.n206 gnd 0.012468f
C1268 commonsourceibias.n207 gnd 0.012468f
C1269 commonsourceibias.n208 gnd 0.008392f
C1270 commonsourceibias.n209 gnd 0.009606f
C1271 commonsourceibias.n210 gnd 0.009606f
C1272 commonsourceibias.n211 gnd 0.008572f
C1273 commonsourceibias.n212 gnd 0.013414f
C1274 commonsourceibias.n213 gnd 0.071606f
C1275 commonsourceibias.n214 gnd 0.013416f
C1276 commonsourceibias.n215 gnd 0.009606f
C1277 commonsourceibias.n216 gnd 0.009606f
C1278 commonsourceibias.n217 gnd 0.009606f
C1279 commonsourceibias.n218 gnd 0.011742f
C1280 commonsourceibias.n219 gnd 0.071606f
C1281 commonsourceibias.n220 gnd 0.012378f
C1282 commonsourceibias.n221 gnd 0.012558f
C1283 commonsourceibias.n222 gnd 0.009606f
C1284 commonsourceibias.n223 gnd 0.009606f
C1285 commonsourceibias.n224 gnd 0.009606f
C1286 commonsourceibias.n225 gnd 0.008375f
C1287 commonsourceibias.n226 gnd 0.013406f
C1288 commonsourceibias.n227 gnd 0.071606f
C1289 commonsourceibias.n228 gnd 0.01341f
C1290 commonsourceibias.n229 gnd 0.009606f
C1291 commonsourceibias.n230 gnd 0.009606f
C1292 commonsourceibias.n231 gnd 0.009606f
C1293 commonsourceibias.n232 gnd 0.011489f
C1294 commonsourceibias.n233 gnd 0.071606f
C1295 commonsourceibias.n234 gnd 0.012289f
C1296 commonsourceibias.n235 gnd 0.012648f
C1297 commonsourceibias.n236 gnd 0.009606f
C1298 commonsourceibias.n237 gnd 0.009606f
C1299 commonsourceibias.n238 gnd 0.009606f
C1300 commonsourceibias.n239 gnd 0.008208f
C1301 commonsourceibias.n240 gnd 0.013389f
C1302 commonsourceibias.n241 gnd 0.071606f
C1303 commonsourceibias.n242 gnd 0.013398f
C1304 commonsourceibias.n243 gnd 0.009606f
C1305 commonsourceibias.n244 gnd 0.009606f
C1306 commonsourceibias.n245 gnd 0.009606f
C1307 commonsourceibias.n246 gnd 0.011208f
C1308 commonsourceibias.n247 gnd 0.071606f
C1309 commonsourceibias.n248 gnd 0.011785f
C1310 commonsourceibias.n249 gnd 0.085921f
C1311 commonsourceibias.n250 gnd 0.056157f
C1312 commonsourceibias.n251 gnd 0.012818f
C1313 commonsourceibias.t145 gnd 0.19409f
C1314 commonsourceibias.t172 gnd 0.179464f
C1315 commonsourceibias.n252 gnd 0.00935f
C1316 commonsourceibias.n253 gnd 0.009606f
C1317 commonsourceibias.t160 gnd 0.179464f
C1318 commonsourceibias.n254 gnd 0.012358f
C1319 commonsourceibias.n255 gnd 0.009606f
C1320 commonsourceibias.t146 gnd 0.179464f
C1321 commonsourceibias.n256 gnd 0.071606f
C1322 commonsourceibias.t173 gnd 0.179464f
C1323 commonsourceibias.n257 gnd 0.009057f
C1324 commonsourceibias.n258 gnd 0.009606f
C1325 commonsourceibias.t158 gnd 0.179464f
C1326 commonsourceibias.n259 gnd 0.012175f
C1327 commonsourceibias.n260 gnd 0.009606f
C1328 commonsourceibias.t144 gnd 0.179464f
C1329 commonsourceibias.n261 gnd 0.071606f
C1330 commonsourceibias.t174 gnd 0.179464f
C1331 commonsourceibias.n262 gnd 0.008798f
C1332 commonsourceibias.n263 gnd 0.009606f
C1333 commonsourceibias.t159 gnd 0.179464f
C1334 commonsourceibias.n264 gnd 0.01197f
C1335 commonsourceibias.n265 gnd 0.009606f
C1336 commonsourceibias.t185 gnd 0.179464f
C1337 commonsourceibias.n266 gnd 0.071606f
C1338 commonsourceibias.t175 gnd 0.179464f
C1339 commonsourceibias.n267 gnd 0.008572f
C1340 commonsourceibias.n268 gnd 0.009606f
C1341 commonsourceibias.t157 gnd 0.179464f
C1342 commonsourceibias.n269 gnd 0.011742f
C1343 commonsourceibias.n270 gnd 0.009606f
C1344 commonsourceibias.t190 gnd 0.179464f
C1345 commonsourceibias.n271 gnd 0.071606f
C1346 commonsourceibias.t91 gnd 0.179464f
C1347 commonsourceibias.n272 gnd 0.008375f
C1348 commonsourceibias.n273 gnd 0.009606f
C1349 commonsourceibias.t169 gnd 0.179464f
C1350 commonsourceibias.n274 gnd 0.011489f
C1351 commonsourceibias.n275 gnd 0.009606f
C1352 commonsourceibias.t82 gnd 0.179464f
C1353 commonsourceibias.n276 gnd 0.071606f
C1354 commonsourceibias.t95 gnd 0.179464f
C1355 commonsourceibias.n277 gnd 0.008208f
C1356 commonsourceibias.n278 gnd 0.009606f
C1357 commonsourceibias.t90 gnd 0.179464f
C1358 commonsourceibias.n279 gnd 0.011208f
C1359 commonsourceibias.t94 gnd 0.199531f
C1360 commonsourceibias.t80 gnd 0.179464f
C1361 commonsourceibias.n280 gnd 0.078223f
C1362 commonsourceibias.n281 gnd 0.08584f
C1363 commonsourceibias.n282 gnd 0.039831f
C1364 commonsourceibias.n283 gnd 0.009606f
C1365 commonsourceibias.n284 gnd 0.00935f
C1366 commonsourceibias.n285 gnd 0.013398f
C1367 commonsourceibias.n286 gnd 0.071606f
C1368 commonsourceibias.n287 gnd 0.013389f
C1369 commonsourceibias.n288 gnd 0.009606f
C1370 commonsourceibias.n289 gnd 0.009606f
C1371 commonsourceibias.n290 gnd 0.009606f
C1372 commonsourceibias.n291 gnd 0.012358f
C1373 commonsourceibias.n292 gnd 0.071606f
C1374 commonsourceibias.n293 gnd 0.012648f
C1375 commonsourceibias.n294 gnd 0.012289f
C1376 commonsourceibias.n295 gnd 0.009606f
C1377 commonsourceibias.n296 gnd 0.009606f
C1378 commonsourceibias.n297 gnd 0.009606f
C1379 commonsourceibias.n298 gnd 0.009057f
C1380 commonsourceibias.n299 gnd 0.01341f
C1381 commonsourceibias.n300 gnd 0.071606f
C1382 commonsourceibias.n301 gnd 0.013406f
C1383 commonsourceibias.n302 gnd 0.009606f
C1384 commonsourceibias.n303 gnd 0.009606f
C1385 commonsourceibias.n304 gnd 0.009606f
C1386 commonsourceibias.n305 gnd 0.012175f
C1387 commonsourceibias.n306 gnd 0.071606f
C1388 commonsourceibias.n307 gnd 0.012558f
C1389 commonsourceibias.n308 gnd 0.012378f
C1390 commonsourceibias.n309 gnd 0.009606f
C1391 commonsourceibias.n310 gnd 0.009606f
C1392 commonsourceibias.n311 gnd 0.009606f
C1393 commonsourceibias.n312 gnd 0.008798f
C1394 commonsourceibias.n313 gnd 0.013416f
C1395 commonsourceibias.n314 gnd 0.071606f
C1396 commonsourceibias.n315 gnd 0.013414f
C1397 commonsourceibias.n316 gnd 0.009606f
C1398 commonsourceibias.n317 gnd 0.009606f
C1399 commonsourceibias.n318 gnd 0.009606f
C1400 commonsourceibias.n319 gnd 0.01197f
C1401 commonsourceibias.n320 gnd 0.071606f
C1402 commonsourceibias.n321 gnd 0.012468f
C1403 commonsourceibias.n322 gnd 0.012468f
C1404 commonsourceibias.n323 gnd 0.009606f
C1405 commonsourceibias.n324 gnd 0.009606f
C1406 commonsourceibias.n325 gnd 0.009606f
C1407 commonsourceibias.n326 gnd 0.008572f
C1408 commonsourceibias.n327 gnd 0.013414f
C1409 commonsourceibias.n328 gnd 0.071606f
C1410 commonsourceibias.n329 gnd 0.013416f
C1411 commonsourceibias.n330 gnd 0.009606f
C1412 commonsourceibias.n331 gnd 0.009606f
C1413 commonsourceibias.n332 gnd 0.009606f
C1414 commonsourceibias.n333 gnd 0.011742f
C1415 commonsourceibias.n334 gnd 0.071606f
C1416 commonsourceibias.n335 gnd 0.012378f
C1417 commonsourceibias.n336 gnd 0.012558f
C1418 commonsourceibias.n337 gnd 0.009606f
C1419 commonsourceibias.n338 gnd 0.009606f
C1420 commonsourceibias.n339 gnd 0.009606f
C1421 commonsourceibias.n340 gnd 0.008375f
C1422 commonsourceibias.n341 gnd 0.013406f
C1423 commonsourceibias.n342 gnd 0.071606f
C1424 commonsourceibias.n343 gnd 0.01341f
C1425 commonsourceibias.n344 gnd 0.009606f
C1426 commonsourceibias.n345 gnd 0.009606f
C1427 commonsourceibias.n346 gnd 0.009606f
C1428 commonsourceibias.n347 gnd 0.011489f
C1429 commonsourceibias.n348 gnd 0.071606f
C1430 commonsourceibias.n349 gnd 0.012289f
C1431 commonsourceibias.n350 gnd 0.012648f
C1432 commonsourceibias.n351 gnd 0.009606f
C1433 commonsourceibias.n352 gnd 0.009606f
C1434 commonsourceibias.n353 gnd 0.009606f
C1435 commonsourceibias.n354 gnd 0.008208f
C1436 commonsourceibias.n355 gnd 0.013389f
C1437 commonsourceibias.n356 gnd 0.071606f
C1438 commonsourceibias.n357 gnd 0.013398f
C1439 commonsourceibias.n358 gnd 0.009606f
C1440 commonsourceibias.n359 gnd 0.009606f
C1441 commonsourceibias.n360 gnd 0.009606f
C1442 commonsourceibias.n361 gnd 0.011208f
C1443 commonsourceibias.n362 gnd 0.071606f
C1444 commonsourceibias.n363 gnd 0.011785f
C1445 commonsourceibias.n364 gnd 0.085921f
C1446 commonsourceibias.n365 gnd 0.029883f
C1447 commonsourceibias.n366 gnd 0.153513f
C1448 commonsourceibias.n367 gnd 0.012818f
C1449 commonsourceibias.t89 gnd 0.179464f
C1450 commonsourceibias.n368 gnd 0.00935f
C1451 commonsourceibias.n369 gnd 0.009606f
C1452 commonsourceibias.t107 gnd 0.179464f
C1453 commonsourceibias.n370 gnd 0.012358f
C1454 commonsourceibias.n371 gnd 0.009606f
C1455 commonsourceibias.t168 gnd 0.179464f
C1456 commonsourceibias.n372 gnd 0.071606f
C1457 commonsourceibias.t199 gnd 0.179464f
C1458 commonsourceibias.n373 gnd 0.009057f
C1459 commonsourceibias.n374 gnd 0.009606f
C1460 commonsourceibias.t98 gnd 0.179464f
C1461 commonsourceibias.n375 gnd 0.012175f
C1462 commonsourceibias.n376 gnd 0.009606f
C1463 commonsourceibias.t150 gnd 0.179464f
C1464 commonsourceibias.n377 gnd 0.071606f
C1465 commonsourceibias.t141 gnd 0.179464f
C1466 commonsourceibias.n378 gnd 0.008798f
C1467 commonsourceibias.n379 gnd 0.009606f
C1468 commonsourceibias.t88 gnd 0.179464f
C1469 commonsourceibias.n380 gnd 0.01197f
C1470 commonsourceibias.n381 gnd 0.009606f
C1471 commonsourceibias.t108 gnd 0.179464f
C1472 commonsourceibias.n382 gnd 0.071606f
C1473 commonsourceibias.t130 gnd 0.179464f
C1474 commonsourceibias.n383 gnd 0.008572f
C1475 commonsourceibias.n384 gnd 0.009606f
C1476 commonsourceibias.t198 gnd 0.179464f
C1477 commonsourceibias.n385 gnd 0.011742f
C1478 commonsourceibias.n386 gnd 0.009606f
C1479 commonsourceibias.t186 gnd 0.179464f
C1480 commonsourceibias.n387 gnd 0.071606f
C1481 commonsourceibias.t92 gnd 0.179464f
C1482 commonsourceibias.n388 gnd 0.008375f
C1483 commonsourceibias.n389 gnd 0.009606f
C1484 commonsourceibias.t177 gnd 0.179464f
C1485 commonsourceibias.n390 gnd 0.011489f
C1486 commonsourceibias.n391 gnd 0.009606f
C1487 commonsourceibias.t170 gnd 0.179464f
C1488 commonsourceibias.n392 gnd 0.071606f
C1489 commonsourceibias.t81 gnd 0.179464f
C1490 commonsourceibias.n393 gnd 0.008208f
C1491 commonsourceibias.n394 gnd 0.009606f
C1492 commonsourceibias.t99 gnd 0.179464f
C1493 commonsourceibias.n395 gnd 0.011208f
C1494 commonsourceibias.t184 gnd 0.199531f
C1495 commonsourceibias.t151 gnd 0.179464f
C1496 commonsourceibias.n396 gnd 0.078223f
C1497 commonsourceibias.n397 gnd 0.08584f
C1498 commonsourceibias.n398 gnd 0.039831f
C1499 commonsourceibias.n399 gnd 0.009606f
C1500 commonsourceibias.n400 gnd 0.00935f
C1501 commonsourceibias.n401 gnd 0.013398f
C1502 commonsourceibias.n402 gnd 0.071606f
C1503 commonsourceibias.n403 gnd 0.013389f
C1504 commonsourceibias.n404 gnd 0.009606f
C1505 commonsourceibias.n405 gnd 0.009606f
C1506 commonsourceibias.n406 gnd 0.009606f
C1507 commonsourceibias.n407 gnd 0.012358f
C1508 commonsourceibias.n408 gnd 0.071606f
C1509 commonsourceibias.n409 gnd 0.012648f
C1510 commonsourceibias.n410 gnd 0.012289f
C1511 commonsourceibias.n411 gnd 0.009606f
C1512 commonsourceibias.n412 gnd 0.009606f
C1513 commonsourceibias.n413 gnd 0.009606f
C1514 commonsourceibias.n414 gnd 0.009057f
C1515 commonsourceibias.n415 gnd 0.01341f
C1516 commonsourceibias.n416 gnd 0.071606f
C1517 commonsourceibias.n417 gnd 0.013406f
C1518 commonsourceibias.n418 gnd 0.009606f
C1519 commonsourceibias.n419 gnd 0.009606f
C1520 commonsourceibias.n420 gnd 0.009606f
C1521 commonsourceibias.n421 gnd 0.012175f
C1522 commonsourceibias.n422 gnd 0.071606f
C1523 commonsourceibias.n423 gnd 0.012558f
C1524 commonsourceibias.n424 gnd 0.012378f
C1525 commonsourceibias.n425 gnd 0.009606f
C1526 commonsourceibias.n426 gnd 0.009606f
C1527 commonsourceibias.n427 gnd 0.009606f
C1528 commonsourceibias.n428 gnd 0.008798f
C1529 commonsourceibias.n429 gnd 0.013416f
C1530 commonsourceibias.n430 gnd 0.071606f
C1531 commonsourceibias.n431 gnd 0.013414f
C1532 commonsourceibias.n432 gnd 0.009606f
C1533 commonsourceibias.n433 gnd 0.009606f
C1534 commonsourceibias.n434 gnd 0.009606f
C1535 commonsourceibias.n435 gnd 0.01197f
C1536 commonsourceibias.n436 gnd 0.071606f
C1537 commonsourceibias.n437 gnd 0.012468f
C1538 commonsourceibias.n438 gnd 0.012468f
C1539 commonsourceibias.n439 gnd 0.009606f
C1540 commonsourceibias.n440 gnd 0.009606f
C1541 commonsourceibias.n441 gnd 0.009606f
C1542 commonsourceibias.n442 gnd 0.008572f
C1543 commonsourceibias.n443 gnd 0.013414f
C1544 commonsourceibias.n444 gnd 0.071606f
C1545 commonsourceibias.n445 gnd 0.013416f
C1546 commonsourceibias.n446 gnd 0.009606f
C1547 commonsourceibias.n447 gnd 0.009606f
C1548 commonsourceibias.n448 gnd 0.009606f
C1549 commonsourceibias.n449 gnd 0.011742f
C1550 commonsourceibias.n450 gnd 0.071606f
C1551 commonsourceibias.n451 gnd 0.012378f
C1552 commonsourceibias.n452 gnd 0.012558f
C1553 commonsourceibias.n453 gnd 0.009606f
C1554 commonsourceibias.n454 gnd 0.009606f
C1555 commonsourceibias.n455 gnd 0.009606f
C1556 commonsourceibias.n456 gnd 0.008375f
C1557 commonsourceibias.n457 gnd 0.013406f
C1558 commonsourceibias.n458 gnd 0.071606f
C1559 commonsourceibias.n459 gnd 0.01341f
C1560 commonsourceibias.n460 gnd 0.009606f
C1561 commonsourceibias.n461 gnd 0.009606f
C1562 commonsourceibias.n462 gnd 0.009606f
C1563 commonsourceibias.n463 gnd 0.011489f
C1564 commonsourceibias.n464 gnd 0.071606f
C1565 commonsourceibias.n465 gnd 0.012289f
C1566 commonsourceibias.n466 gnd 0.012648f
C1567 commonsourceibias.n467 gnd 0.009606f
C1568 commonsourceibias.n468 gnd 0.009606f
C1569 commonsourceibias.n469 gnd 0.009606f
C1570 commonsourceibias.n470 gnd 0.008208f
C1571 commonsourceibias.n471 gnd 0.013389f
C1572 commonsourceibias.n472 gnd 0.071606f
C1573 commonsourceibias.n473 gnd 0.013398f
C1574 commonsourceibias.n474 gnd 0.009606f
C1575 commonsourceibias.n475 gnd 0.009606f
C1576 commonsourceibias.n476 gnd 0.009606f
C1577 commonsourceibias.n477 gnd 0.011208f
C1578 commonsourceibias.n478 gnd 0.071606f
C1579 commonsourceibias.n479 gnd 0.011785f
C1580 commonsourceibias.t183 gnd 0.19409f
C1581 commonsourceibias.n480 gnd 0.085921f
C1582 commonsourceibias.n481 gnd 0.029883f
C1583 commonsourceibias.n482 gnd 0.5392f
C1584 commonsourceibias.n483 gnd 0.012818f
C1585 commonsourceibias.t191 gnd 0.19409f
C1586 commonsourceibias.t134 gnd 0.179464f
C1587 commonsourceibias.n484 gnd 0.00935f
C1588 commonsourceibias.n485 gnd 0.009606f
C1589 commonsourceibias.t97 gnd 0.179464f
C1590 commonsourceibias.n486 gnd 0.012358f
C1591 commonsourceibias.n487 gnd 0.009606f
C1592 commonsourceibias.t117 gnd 0.179464f
C1593 commonsourceibias.n488 gnd 0.009057f
C1594 commonsourceibias.n489 gnd 0.009606f
C1595 commonsourceibias.t187 gnd 0.179464f
C1596 commonsourceibias.n490 gnd 0.012175f
C1597 commonsourceibias.n491 gnd 0.009606f
C1598 commonsourceibias.t118 gnd 0.179464f
C1599 commonsourceibias.n492 gnd 0.008798f
C1600 commonsourceibias.n493 gnd 0.009606f
C1601 commonsourceibias.t149 gnd 0.179464f
C1602 commonsourceibias.n494 gnd 0.01197f
C1603 commonsourceibias.t17 gnd 0.020728f
C1604 commonsourceibias.t49 gnd 0.020728f
C1605 commonsourceibias.n495 gnd 0.183774f
C1606 commonsourceibias.t25 gnd 0.020728f
C1607 commonsourceibias.t79 gnd 0.020728f
C1608 commonsourceibias.n496 gnd 0.183161f
C1609 commonsourceibias.n497 gnd 0.170671f
C1610 commonsourceibias.t59 gnd 0.020728f
C1611 commonsourceibias.t57 gnd 0.020728f
C1612 commonsourceibias.n498 gnd 0.183161f
C1613 commonsourceibias.n499 gnd 0.084133f
C1614 commonsourceibias.t73 gnd 0.020728f
C1615 commonsourceibias.t61 gnd 0.020728f
C1616 commonsourceibias.n500 gnd 0.183161f
C1617 commonsourceibias.n501 gnd 0.084133f
C1618 commonsourceibias.t5 gnd 0.020728f
C1619 commonsourceibias.t55 gnd 0.020728f
C1620 commonsourceibias.n502 gnd 0.183161f
C1621 commonsourceibias.n503 gnd 0.070289f
C1622 commonsourceibias.n504 gnd 0.012818f
C1623 commonsourceibias.t28 gnd 0.179464f
C1624 commonsourceibias.n505 gnd 0.00935f
C1625 commonsourceibias.n506 gnd 0.009606f
C1626 commonsourceibias.t10 gnd 0.179464f
C1627 commonsourceibias.n507 gnd 0.012358f
C1628 commonsourceibias.n508 gnd 0.009606f
C1629 commonsourceibias.t22 gnd 0.179464f
C1630 commonsourceibias.n509 gnd 0.009057f
C1631 commonsourceibias.n510 gnd 0.009606f
C1632 commonsourceibias.t44 gnd 0.179464f
C1633 commonsourceibias.n511 gnd 0.012175f
C1634 commonsourceibias.n512 gnd 0.009606f
C1635 commonsourceibias.t20 gnd 0.179464f
C1636 commonsourceibias.n513 gnd 0.008798f
C1637 commonsourceibias.n514 gnd 0.009606f
C1638 commonsourceibias.t30 gnd 0.179464f
C1639 commonsourceibias.n515 gnd 0.01197f
C1640 commonsourceibias.n516 gnd 0.009606f
C1641 commonsourceibias.t54 gnd 0.179464f
C1642 commonsourceibias.n517 gnd 0.008572f
C1643 commonsourceibias.n518 gnd 0.009606f
C1644 commonsourceibias.t4 gnd 0.179464f
C1645 commonsourceibias.n519 gnd 0.011742f
C1646 commonsourceibias.n520 gnd 0.009606f
C1647 commonsourceibias.t72 gnd 0.179464f
C1648 commonsourceibias.n521 gnd 0.008375f
C1649 commonsourceibias.n522 gnd 0.009606f
C1650 commonsourceibias.t56 gnd 0.179464f
C1651 commonsourceibias.n523 gnd 0.011489f
C1652 commonsourceibias.n524 gnd 0.009606f
C1653 commonsourceibias.t78 gnd 0.179464f
C1654 commonsourceibias.n525 gnd 0.008208f
C1655 commonsourceibias.n526 gnd 0.009606f
C1656 commonsourceibias.t24 gnd 0.179464f
C1657 commonsourceibias.n527 gnd 0.011208f
C1658 commonsourceibias.t16 gnd 0.199531f
C1659 commonsourceibias.t48 gnd 0.179464f
C1660 commonsourceibias.n528 gnd 0.078223f
C1661 commonsourceibias.n529 gnd 0.08584f
C1662 commonsourceibias.n530 gnd 0.039831f
C1663 commonsourceibias.n531 gnd 0.009606f
C1664 commonsourceibias.n532 gnd 0.00935f
C1665 commonsourceibias.n533 gnd 0.013398f
C1666 commonsourceibias.n534 gnd 0.071606f
C1667 commonsourceibias.n535 gnd 0.013389f
C1668 commonsourceibias.n536 gnd 0.009606f
C1669 commonsourceibias.n537 gnd 0.009606f
C1670 commonsourceibias.n538 gnd 0.009606f
C1671 commonsourceibias.n539 gnd 0.012358f
C1672 commonsourceibias.n540 gnd 0.071606f
C1673 commonsourceibias.n541 gnd 0.012648f
C1674 commonsourceibias.t58 gnd 0.179464f
C1675 commonsourceibias.n542 gnd 0.071606f
C1676 commonsourceibias.n543 gnd 0.012289f
C1677 commonsourceibias.n544 gnd 0.009606f
C1678 commonsourceibias.n545 gnd 0.009606f
C1679 commonsourceibias.n546 gnd 0.009606f
C1680 commonsourceibias.n547 gnd 0.009057f
C1681 commonsourceibias.n548 gnd 0.01341f
C1682 commonsourceibias.n549 gnd 0.071606f
C1683 commonsourceibias.n550 gnd 0.013406f
C1684 commonsourceibias.n551 gnd 0.009606f
C1685 commonsourceibias.n552 gnd 0.009606f
C1686 commonsourceibias.n553 gnd 0.009606f
C1687 commonsourceibias.n554 gnd 0.012175f
C1688 commonsourceibias.n555 gnd 0.071606f
C1689 commonsourceibias.n556 gnd 0.012558f
C1690 commonsourceibias.t60 gnd 0.179464f
C1691 commonsourceibias.n557 gnd 0.071606f
C1692 commonsourceibias.n558 gnd 0.012378f
C1693 commonsourceibias.n559 gnd 0.009606f
C1694 commonsourceibias.n560 gnd 0.009606f
C1695 commonsourceibias.n561 gnd 0.009606f
C1696 commonsourceibias.n562 gnd 0.008798f
C1697 commonsourceibias.n563 gnd 0.013416f
C1698 commonsourceibias.n564 gnd 0.071606f
C1699 commonsourceibias.n565 gnd 0.013414f
C1700 commonsourceibias.n566 gnd 0.009606f
C1701 commonsourceibias.n567 gnd 0.009606f
C1702 commonsourceibias.n568 gnd 0.009606f
C1703 commonsourceibias.n569 gnd 0.01197f
C1704 commonsourceibias.n570 gnd 0.071606f
C1705 commonsourceibias.n571 gnd 0.012468f
C1706 commonsourceibias.t62 gnd 0.179464f
C1707 commonsourceibias.n572 gnd 0.071606f
C1708 commonsourceibias.n573 gnd 0.012468f
C1709 commonsourceibias.n574 gnd 0.009606f
C1710 commonsourceibias.n575 gnd 0.009606f
C1711 commonsourceibias.n576 gnd 0.009606f
C1712 commonsourceibias.n577 gnd 0.008572f
C1713 commonsourceibias.n578 gnd 0.013414f
C1714 commonsourceibias.n579 gnd 0.071606f
C1715 commonsourceibias.n580 gnd 0.013416f
C1716 commonsourceibias.n581 gnd 0.009606f
C1717 commonsourceibias.n582 gnd 0.009606f
C1718 commonsourceibias.n583 gnd 0.009606f
C1719 commonsourceibias.n584 gnd 0.011742f
C1720 commonsourceibias.n585 gnd 0.071606f
C1721 commonsourceibias.n586 gnd 0.012378f
C1722 commonsourceibias.t68 gnd 0.179464f
C1723 commonsourceibias.n587 gnd 0.071606f
C1724 commonsourceibias.n588 gnd 0.012558f
C1725 commonsourceibias.n589 gnd 0.009606f
C1726 commonsourceibias.n590 gnd 0.009606f
C1727 commonsourceibias.n591 gnd 0.009606f
C1728 commonsourceibias.n592 gnd 0.008375f
C1729 commonsourceibias.n593 gnd 0.013406f
C1730 commonsourceibias.n594 gnd 0.071606f
C1731 commonsourceibias.n595 gnd 0.01341f
C1732 commonsourceibias.n596 gnd 0.009606f
C1733 commonsourceibias.n597 gnd 0.009606f
C1734 commonsourceibias.n598 gnd 0.009606f
C1735 commonsourceibias.n599 gnd 0.011489f
C1736 commonsourceibias.n600 gnd 0.071606f
C1737 commonsourceibias.n601 gnd 0.012289f
C1738 commonsourceibias.t18 gnd 0.179464f
C1739 commonsourceibias.n602 gnd 0.071606f
C1740 commonsourceibias.n603 gnd 0.012648f
C1741 commonsourceibias.n604 gnd 0.009606f
C1742 commonsourceibias.n605 gnd 0.009606f
C1743 commonsourceibias.n606 gnd 0.009606f
C1744 commonsourceibias.n607 gnd 0.008208f
C1745 commonsourceibias.n608 gnd 0.013389f
C1746 commonsourceibias.n609 gnd 0.071606f
C1747 commonsourceibias.n610 gnd 0.013398f
C1748 commonsourceibias.n611 gnd 0.009606f
C1749 commonsourceibias.n612 gnd 0.009606f
C1750 commonsourceibias.n613 gnd 0.009606f
C1751 commonsourceibias.n614 gnd 0.011208f
C1752 commonsourceibias.n615 gnd 0.071606f
C1753 commonsourceibias.n616 gnd 0.011785f
C1754 commonsourceibias.t42 gnd 0.19409f
C1755 commonsourceibias.n617 gnd 0.085921f
C1756 commonsourceibias.n618 gnd 0.095704f
C1757 commonsourceibias.t29 gnd 0.020728f
C1758 commonsourceibias.t43 gnd 0.020728f
C1759 commonsourceibias.n619 gnd 0.183161f
C1760 commonsourceibias.n620 gnd 0.158435f
C1761 commonsourceibias.t19 gnd 0.020728f
C1762 commonsourceibias.t11 gnd 0.020728f
C1763 commonsourceibias.n621 gnd 0.183161f
C1764 commonsourceibias.n622 gnd 0.084133f
C1765 commonsourceibias.t45 gnd 0.020728f
C1766 commonsourceibias.t23 gnd 0.020728f
C1767 commonsourceibias.n623 gnd 0.183161f
C1768 commonsourceibias.n624 gnd 0.084133f
C1769 commonsourceibias.t21 gnd 0.020728f
C1770 commonsourceibias.t69 gnd 0.020728f
C1771 commonsourceibias.n625 gnd 0.183161f
C1772 commonsourceibias.n626 gnd 0.084133f
C1773 commonsourceibias.t63 gnd 0.020728f
C1774 commonsourceibias.t31 gnd 0.020728f
C1775 commonsourceibias.n627 gnd 0.183161f
C1776 commonsourceibias.n628 gnd 0.070289f
C1777 commonsourceibias.n629 gnd 0.085113f
C1778 commonsourceibias.n630 gnd 0.062168f
C1779 commonsourceibias.t105 gnd 0.179464f
C1780 commonsourceibias.n631 gnd 0.071606f
C1781 commonsourceibias.n632 gnd 0.009606f
C1782 commonsourceibias.t122 gnd 0.179464f
C1783 commonsourceibias.n633 gnd 0.071606f
C1784 commonsourceibias.n634 gnd 0.009606f
C1785 commonsourceibias.t115 gnd 0.179464f
C1786 commonsourceibias.n635 gnd 0.071606f
C1787 commonsourceibias.n636 gnd 0.009606f
C1788 commonsourceibias.t83 gnd 0.179464f
C1789 commonsourceibias.n637 gnd 0.008375f
C1790 commonsourceibias.n638 gnd 0.009606f
C1791 commonsourceibias.t111 gnd 0.179464f
C1792 commonsourceibias.n639 gnd 0.011489f
C1793 commonsourceibias.n640 gnd 0.009606f
C1794 commonsourceibias.t192 gnd 0.179464f
C1795 commonsourceibias.n641 gnd 0.008208f
C1796 commonsourceibias.n642 gnd 0.009606f
C1797 commonsourceibias.t127 gnd 0.179464f
C1798 commonsourceibias.n643 gnd 0.011208f
C1799 commonsourceibias.t153 gnd 0.199531f
C1800 commonsourceibias.t86 gnd 0.179464f
C1801 commonsourceibias.n644 gnd 0.078223f
C1802 commonsourceibias.n645 gnd 0.08584f
C1803 commonsourceibias.n646 gnd 0.039831f
C1804 commonsourceibias.n647 gnd 0.009606f
C1805 commonsourceibias.n648 gnd 0.00935f
C1806 commonsourceibias.n649 gnd 0.013398f
C1807 commonsourceibias.n650 gnd 0.071606f
C1808 commonsourceibias.n651 gnd 0.013389f
C1809 commonsourceibias.n652 gnd 0.009606f
C1810 commonsourceibias.n653 gnd 0.009606f
C1811 commonsourceibias.n654 gnd 0.009606f
C1812 commonsourceibias.n655 gnd 0.012358f
C1813 commonsourceibias.n656 gnd 0.071606f
C1814 commonsourceibias.n657 gnd 0.012648f
C1815 commonsourceibias.t110 gnd 0.179464f
C1816 commonsourceibias.n658 gnd 0.071606f
C1817 commonsourceibias.n659 gnd 0.012289f
C1818 commonsourceibias.n660 gnd 0.009606f
C1819 commonsourceibias.n661 gnd 0.009606f
C1820 commonsourceibias.n662 gnd 0.009606f
C1821 commonsourceibias.n663 gnd 0.009057f
C1822 commonsourceibias.n664 gnd 0.01341f
C1823 commonsourceibias.n665 gnd 0.071606f
C1824 commonsourceibias.n666 gnd 0.013406f
C1825 commonsourceibias.n667 gnd 0.009606f
C1826 commonsourceibias.n668 gnd 0.009606f
C1827 commonsourceibias.n669 gnd 0.009606f
C1828 commonsourceibias.n670 gnd 0.012175f
C1829 commonsourceibias.n671 gnd 0.071606f
C1830 commonsourceibias.n672 gnd 0.012558f
C1831 commonsourceibias.n673 gnd 0.012378f
C1832 commonsourceibias.n674 gnd 0.009606f
C1833 commonsourceibias.n675 gnd 0.009606f
C1834 commonsourceibias.n676 gnd 0.011742f
C1835 commonsourceibias.n677 gnd 0.008798f
C1836 commonsourceibias.n678 gnd 0.013416f
C1837 commonsourceibias.n679 gnd 0.009606f
C1838 commonsourceibias.n680 gnd 0.009606f
C1839 commonsourceibias.n681 gnd 0.013414f
C1840 commonsourceibias.n682 gnd 0.008572f
C1841 commonsourceibias.n683 gnd 0.01197f
C1842 commonsourceibias.n684 gnd 0.009606f
C1843 commonsourceibias.n685 gnd 0.008392f
C1844 commonsourceibias.n686 gnd 0.012468f
C1845 commonsourceibias.t114 gnd 0.179464f
C1846 commonsourceibias.n687 gnd 0.071606f
C1847 commonsourceibias.n688 gnd 0.012468f
C1848 commonsourceibias.n689 gnd 0.008392f
C1849 commonsourceibias.n690 gnd 0.009606f
C1850 commonsourceibias.n691 gnd 0.009606f
C1851 commonsourceibias.n692 gnd 0.008572f
C1852 commonsourceibias.n693 gnd 0.013414f
C1853 commonsourceibias.n694 gnd 0.071606f
C1854 commonsourceibias.n695 gnd 0.013416f
C1855 commonsourceibias.n696 gnd 0.009606f
C1856 commonsourceibias.n697 gnd 0.009606f
C1857 commonsourceibias.n698 gnd 0.009606f
C1858 commonsourceibias.n699 gnd 0.011742f
C1859 commonsourceibias.n700 gnd 0.071606f
C1860 commonsourceibias.n701 gnd 0.012378f
C1861 commonsourceibias.t132 gnd 0.179464f
C1862 commonsourceibias.n702 gnd 0.071606f
C1863 commonsourceibias.n703 gnd 0.012558f
C1864 commonsourceibias.n704 gnd 0.009606f
C1865 commonsourceibias.n705 gnd 0.009606f
C1866 commonsourceibias.n706 gnd 0.009606f
C1867 commonsourceibias.n707 gnd 0.008375f
C1868 commonsourceibias.n708 gnd 0.013406f
C1869 commonsourceibias.n709 gnd 0.071606f
C1870 commonsourceibias.n710 gnd 0.01341f
C1871 commonsourceibias.n711 gnd 0.009606f
C1872 commonsourceibias.n712 gnd 0.009606f
C1873 commonsourceibias.n713 gnd 0.009606f
C1874 commonsourceibias.n714 gnd 0.011489f
C1875 commonsourceibias.n715 gnd 0.071606f
C1876 commonsourceibias.n716 gnd 0.012289f
C1877 commonsourceibias.t152 gnd 0.179464f
C1878 commonsourceibias.n717 gnd 0.071606f
C1879 commonsourceibias.n718 gnd 0.012648f
C1880 commonsourceibias.n719 gnd 0.009606f
C1881 commonsourceibias.n720 gnd 0.009606f
C1882 commonsourceibias.n721 gnd 0.009606f
C1883 commonsourceibias.n722 gnd 0.008208f
C1884 commonsourceibias.n723 gnd 0.013389f
C1885 commonsourceibias.n724 gnd 0.071606f
C1886 commonsourceibias.n725 gnd 0.013398f
C1887 commonsourceibias.n726 gnd 0.009606f
C1888 commonsourceibias.n727 gnd 0.009606f
C1889 commonsourceibias.n728 gnd 0.009606f
C1890 commonsourceibias.n729 gnd 0.011208f
C1891 commonsourceibias.n730 gnd 0.071606f
C1892 commonsourceibias.n731 gnd 0.011785f
C1893 commonsourceibias.n732 gnd 0.085921f
C1894 commonsourceibias.n733 gnd 0.056157f
C1895 commonsourceibias.n734 gnd 0.012818f
C1896 commonsourceibias.t148 gnd 0.179464f
C1897 commonsourceibias.n735 gnd 0.00935f
C1898 commonsourceibias.n736 gnd 0.009606f
C1899 commonsourceibias.t139 gnd 0.179464f
C1900 commonsourceibias.n737 gnd 0.012358f
C1901 commonsourceibias.n738 gnd 0.009606f
C1902 commonsourceibias.t147 gnd 0.179464f
C1903 commonsourceibias.n739 gnd 0.009057f
C1904 commonsourceibias.n740 gnd 0.009606f
C1905 commonsourceibias.t138 gnd 0.179464f
C1906 commonsourceibias.n741 gnd 0.012175f
C1907 commonsourceibias.n742 gnd 0.009606f
C1908 commonsourceibias.t154 gnd 0.179464f
C1909 commonsourceibias.n743 gnd 0.008798f
C1910 commonsourceibias.n744 gnd 0.009606f
C1911 commonsourceibias.t137 gnd 0.179464f
C1912 commonsourceibias.n745 gnd 0.01197f
C1913 commonsourceibias.n746 gnd 0.009606f
C1914 commonsourceibias.t195 gnd 0.179464f
C1915 commonsourceibias.n747 gnd 0.008572f
C1916 commonsourceibias.n748 gnd 0.009606f
C1917 commonsourceibias.t135 gnd 0.179464f
C1918 commonsourceibias.n749 gnd 0.011742f
C1919 commonsourceibias.n750 gnd 0.009606f
C1920 commonsourceibias.t194 gnd 0.179464f
C1921 commonsourceibias.n751 gnd 0.008375f
C1922 commonsourceibias.n752 gnd 0.009606f
C1923 commonsourceibias.t176 gnd 0.179464f
C1924 commonsourceibias.n753 gnd 0.011489f
C1925 commonsourceibias.n754 gnd 0.009606f
C1926 commonsourceibias.t189 gnd 0.179464f
C1927 commonsourceibias.n755 gnd 0.008208f
C1928 commonsourceibias.n756 gnd 0.009606f
C1929 commonsourceibias.t180 gnd 0.179464f
C1930 commonsourceibias.n757 gnd 0.011208f
C1931 commonsourceibias.t188 gnd 0.199531f
C1932 commonsourceibias.t163 gnd 0.179464f
C1933 commonsourceibias.n758 gnd 0.078223f
C1934 commonsourceibias.n759 gnd 0.08584f
C1935 commonsourceibias.n760 gnd 0.039831f
C1936 commonsourceibias.n761 gnd 0.009606f
C1937 commonsourceibias.n762 gnd 0.00935f
C1938 commonsourceibias.n763 gnd 0.013398f
C1939 commonsourceibias.n764 gnd 0.071606f
C1940 commonsourceibias.n765 gnd 0.013389f
C1941 commonsourceibias.n766 gnd 0.009606f
C1942 commonsourceibias.n767 gnd 0.009606f
C1943 commonsourceibias.n768 gnd 0.009606f
C1944 commonsourceibias.n769 gnd 0.012358f
C1945 commonsourceibias.n770 gnd 0.071606f
C1946 commonsourceibias.n771 gnd 0.012648f
C1947 commonsourceibias.t164 gnd 0.179464f
C1948 commonsourceibias.n772 gnd 0.071606f
C1949 commonsourceibias.n773 gnd 0.012289f
C1950 commonsourceibias.n774 gnd 0.009606f
C1951 commonsourceibias.n775 gnd 0.009606f
C1952 commonsourceibias.n776 gnd 0.009606f
C1953 commonsourceibias.n777 gnd 0.009057f
C1954 commonsourceibias.n778 gnd 0.01341f
C1955 commonsourceibias.n779 gnd 0.071606f
C1956 commonsourceibias.n780 gnd 0.013406f
C1957 commonsourceibias.n781 gnd 0.009606f
C1958 commonsourceibias.n782 gnd 0.009606f
C1959 commonsourceibias.n783 gnd 0.009606f
C1960 commonsourceibias.n784 gnd 0.012175f
C1961 commonsourceibias.n785 gnd 0.071606f
C1962 commonsourceibias.n786 gnd 0.012558f
C1963 commonsourceibias.t171 gnd 0.179464f
C1964 commonsourceibias.n787 gnd 0.071606f
C1965 commonsourceibias.n788 gnd 0.012378f
C1966 commonsourceibias.n789 gnd 0.009606f
C1967 commonsourceibias.n790 gnd 0.009606f
C1968 commonsourceibias.n791 gnd 0.009606f
C1969 commonsourceibias.n792 gnd 0.008798f
C1970 commonsourceibias.n793 gnd 0.013416f
C1971 commonsourceibias.n794 gnd 0.071606f
C1972 commonsourceibias.n795 gnd 0.013414f
C1973 commonsourceibias.n796 gnd 0.009606f
C1974 commonsourceibias.n797 gnd 0.009606f
C1975 commonsourceibias.n798 gnd 0.009606f
C1976 commonsourceibias.n799 gnd 0.01197f
C1977 commonsourceibias.n800 gnd 0.071606f
C1978 commonsourceibias.n801 gnd 0.012468f
C1979 commonsourceibias.t161 gnd 0.179464f
C1980 commonsourceibias.n802 gnd 0.071606f
C1981 commonsourceibias.n803 gnd 0.012468f
C1982 commonsourceibias.n804 gnd 0.009606f
C1983 commonsourceibias.n805 gnd 0.009606f
C1984 commonsourceibias.n806 gnd 0.009606f
C1985 commonsourceibias.n807 gnd 0.008572f
C1986 commonsourceibias.n808 gnd 0.013414f
C1987 commonsourceibias.n809 gnd 0.071606f
C1988 commonsourceibias.n810 gnd 0.013416f
C1989 commonsourceibias.n811 gnd 0.009606f
C1990 commonsourceibias.n812 gnd 0.009606f
C1991 commonsourceibias.n813 gnd 0.009606f
C1992 commonsourceibias.n814 gnd 0.011742f
C1993 commonsourceibias.n815 gnd 0.071606f
C1994 commonsourceibias.n816 gnd 0.012378f
C1995 commonsourceibias.t162 gnd 0.179464f
C1996 commonsourceibias.n817 gnd 0.071606f
C1997 commonsourceibias.n818 gnd 0.012558f
C1998 commonsourceibias.n819 gnd 0.009606f
C1999 commonsourceibias.n820 gnd 0.009606f
C2000 commonsourceibias.n821 gnd 0.009606f
C2001 commonsourceibias.n822 gnd 0.008375f
C2002 commonsourceibias.n823 gnd 0.013406f
C2003 commonsourceibias.n824 gnd 0.071606f
C2004 commonsourceibias.n825 gnd 0.01341f
C2005 commonsourceibias.n826 gnd 0.009606f
C2006 commonsourceibias.n827 gnd 0.009606f
C2007 commonsourceibias.n828 gnd 0.009606f
C2008 commonsourceibias.n829 gnd 0.011489f
C2009 commonsourceibias.n830 gnd 0.071606f
C2010 commonsourceibias.n831 gnd 0.012289f
C2011 commonsourceibias.t128 gnd 0.179464f
C2012 commonsourceibias.n832 gnd 0.071606f
C2013 commonsourceibias.n833 gnd 0.012648f
C2014 commonsourceibias.n834 gnd 0.009606f
C2015 commonsourceibias.n835 gnd 0.009606f
C2016 commonsourceibias.n836 gnd 0.009606f
C2017 commonsourceibias.n837 gnd 0.008208f
C2018 commonsourceibias.n838 gnd 0.013389f
C2019 commonsourceibias.n839 gnd 0.071606f
C2020 commonsourceibias.n840 gnd 0.013398f
C2021 commonsourceibias.n841 gnd 0.009606f
C2022 commonsourceibias.n842 gnd 0.009606f
C2023 commonsourceibias.n843 gnd 0.009606f
C2024 commonsourceibias.n844 gnd 0.011208f
C2025 commonsourceibias.n845 gnd 0.071606f
C2026 commonsourceibias.n846 gnd 0.011785f
C2027 commonsourceibias.t129 gnd 0.19409f
C2028 commonsourceibias.n847 gnd 0.085921f
C2029 commonsourceibias.n848 gnd 0.029883f
C2030 commonsourceibias.n849 gnd 0.153513f
C2031 commonsourceibias.n850 gnd 0.012818f
C2032 commonsourceibias.t113 gnd 0.179464f
C2033 commonsourceibias.n851 gnd 0.00935f
C2034 commonsourceibias.n852 gnd 0.009606f
C2035 commonsourceibias.t125 gnd 0.179464f
C2036 commonsourceibias.n853 gnd 0.012358f
C2037 commonsourceibias.n854 gnd 0.009606f
C2038 commonsourceibias.t103 gnd 0.179464f
C2039 commonsourceibias.n855 gnd 0.009057f
C2040 commonsourceibias.n856 gnd 0.009606f
C2041 commonsourceibias.t120 gnd 0.179464f
C2042 commonsourceibias.n857 gnd 0.012175f
C2043 commonsourceibias.n858 gnd 0.009606f
C2044 commonsourceibias.t179 gnd 0.179464f
C2045 commonsourceibias.n859 gnd 0.008798f
C2046 commonsourceibias.n860 gnd 0.009606f
C2047 commonsourceibias.t112 gnd 0.179464f
C2048 commonsourceibias.n861 gnd 0.01197f
C2049 commonsourceibias.n862 gnd 0.009606f
C2050 commonsourceibias.t121 gnd 0.179464f
C2051 commonsourceibias.n863 gnd 0.008572f
C2052 commonsourceibias.n864 gnd 0.009606f
C2053 commonsourceibias.t102 gnd 0.179464f
C2054 commonsourceibias.n865 gnd 0.011742f
C2055 commonsourceibias.n866 gnd 0.009606f
C2056 commonsourceibias.t116 gnd 0.179464f
C2057 commonsourceibias.n867 gnd 0.008375f
C2058 commonsourceibias.n868 gnd 0.009606f
C2059 commonsourceibias.t167 gnd 0.179464f
C2060 commonsourceibias.n869 gnd 0.011489f
C2061 commonsourceibias.n870 gnd 0.009606f
C2062 commonsourceibias.t87 gnd 0.179464f
C2063 commonsourceibias.n871 gnd 0.008208f
C2064 commonsourceibias.n872 gnd 0.009606f
C2065 commonsourceibias.t106 gnd 0.179464f
C2066 commonsourceibias.n873 gnd 0.011208f
C2067 commonsourceibias.t196 gnd 0.199531f
C2068 commonsourceibias.t165 gnd 0.179464f
C2069 commonsourceibias.n874 gnd 0.078223f
C2070 commonsourceibias.n875 gnd 0.08584f
C2071 commonsourceibias.n876 gnd 0.039831f
C2072 commonsourceibias.n877 gnd 0.009606f
C2073 commonsourceibias.n878 gnd 0.00935f
C2074 commonsourceibias.n879 gnd 0.013398f
C2075 commonsourceibias.n880 gnd 0.071606f
C2076 commonsourceibias.n881 gnd 0.013389f
C2077 commonsourceibias.n882 gnd 0.009606f
C2078 commonsourceibias.n883 gnd 0.009606f
C2079 commonsourceibias.n884 gnd 0.009606f
C2080 commonsourceibias.n885 gnd 0.012358f
C2081 commonsourceibias.n886 gnd 0.071606f
C2082 commonsourceibias.n887 gnd 0.012648f
C2083 commonsourceibias.t178 gnd 0.179464f
C2084 commonsourceibias.n888 gnd 0.071606f
C2085 commonsourceibias.n889 gnd 0.012289f
C2086 commonsourceibias.n890 gnd 0.009606f
C2087 commonsourceibias.n891 gnd 0.009606f
C2088 commonsourceibias.n892 gnd 0.009606f
C2089 commonsourceibias.n893 gnd 0.009057f
C2090 commonsourceibias.n894 gnd 0.01341f
C2091 commonsourceibias.n895 gnd 0.071606f
C2092 commonsourceibias.n896 gnd 0.013406f
C2093 commonsourceibias.n897 gnd 0.009606f
C2094 commonsourceibias.n898 gnd 0.009606f
C2095 commonsourceibias.n899 gnd 0.009606f
C2096 commonsourceibias.n900 gnd 0.012175f
C2097 commonsourceibias.n901 gnd 0.071606f
C2098 commonsourceibias.n902 gnd 0.012558f
C2099 commonsourceibias.t96 gnd 0.179464f
C2100 commonsourceibias.n903 gnd 0.071606f
C2101 commonsourceibias.n904 gnd 0.012378f
C2102 commonsourceibias.n905 gnd 0.009606f
C2103 commonsourceibias.n906 gnd 0.009606f
C2104 commonsourceibias.n907 gnd 0.009606f
C2105 commonsourceibias.n908 gnd 0.008798f
C2106 commonsourceibias.n909 gnd 0.013416f
C2107 commonsourceibias.n910 gnd 0.071606f
C2108 commonsourceibias.n911 gnd 0.013414f
C2109 commonsourceibias.n912 gnd 0.009606f
C2110 commonsourceibias.n913 gnd 0.009606f
C2111 commonsourceibias.n914 gnd 0.009606f
C2112 commonsourceibias.n915 gnd 0.01197f
C2113 commonsourceibias.n916 gnd 0.071606f
C2114 commonsourceibias.n917 gnd 0.012468f
C2115 commonsourceibias.t126 gnd 0.179464f
C2116 commonsourceibias.n918 gnd 0.071606f
C2117 commonsourceibias.n919 gnd 0.012468f
C2118 commonsourceibias.n920 gnd 0.009606f
C2119 commonsourceibias.n921 gnd 0.009606f
C2120 commonsourceibias.n922 gnd 0.009606f
C2121 commonsourceibias.n923 gnd 0.008572f
C2122 commonsourceibias.n924 gnd 0.013414f
C2123 commonsourceibias.n925 gnd 0.071606f
C2124 commonsourceibias.n926 gnd 0.013416f
C2125 commonsourceibias.n927 gnd 0.009606f
C2126 commonsourceibias.n928 gnd 0.009606f
C2127 commonsourceibias.n929 gnd 0.009606f
C2128 commonsourceibias.n930 gnd 0.011742f
C2129 commonsourceibias.n931 gnd 0.071606f
C2130 commonsourceibias.n932 gnd 0.012378f
C2131 commonsourceibias.t133 gnd 0.179464f
C2132 commonsourceibias.n933 gnd 0.071606f
C2133 commonsourceibias.n934 gnd 0.012558f
C2134 commonsourceibias.n935 gnd 0.009606f
C2135 commonsourceibias.n936 gnd 0.009606f
C2136 commonsourceibias.n937 gnd 0.009606f
C2137 commonsourceibias.n938 gnd 0.008375f
C2138 commonsourceibias.n939 gnd 0.013406f
C2139 commonsourceibias.n940 gnd 0.071606f
C2140 commonsourceibias.n941 gnd 0.01341f
C2141 commonsourceibias.n942 gnd 0.009606f
C2142 commonsourceibias.n943 gnd 0.009606f
C2143 commonsourceibias.n944 gnd 0.009606f
C2144 commonsourceibias.n945 gnd 0.011489f
C2145 commonsourceibias.n946 gnd 0.071606f
C2146 commonsourceibias.n947 gnd 0.012289f
C2147 commonsourceibias.t85 gnd 0.179464f
C2148 commonsourceibias.n948 gnd 0.071606f
C2149 commonsourceibias.n949 gnd 0.012648f
C2150 commonsourceibias.n950 gnd 0.009606f
C2151 commonsourceibias.n951 gnd 0.009606f
C2152 commonsourceibias.n952 gnd 0.009606f
C2153 commonsourceibias.n953 gnd 0.008208f
C2154 commonsourceibias.n954 gnd 0.013389f
C2155 commonsourceibias.n955 gnd 0.071606f
C2156 commonsourceibias.n956 gnd 0.013398f
C2157 commonsourceibias.n957 gnd 0.009606f
C2158 commonsourceibias.n958 gnd 0.009606f
C2159 commonsourceibias.n959 gnd 0.009606f
C2160 commonsourceibias.n960 gnd 0.011208f
C2161 commonsourceibias.n961 gnd 0.071606f
C2162 commonsourceibias.n962 gnd 0.011785f
C2163 commonsourceibias.t93 gnd 0.19409f
C2164 commonsourceibias.n963 gnd 0.085921f
C2165 commonsourceibias.n964 gnd 0.029883f
C2166 commonsourceibias.n965 gnd 0.202576f
C2167 commonsourceibias.n966 gnd 5.69738f
C2168 CSoutput.n0 gnd 0.042058f
C2169 CSoutput.t197 gnd 0.278203f
C2170 CSoutput.n1 gnd 0.125622f
C2171 CSoutput.n2 gnd 0.042058f
C2172 CSoutput.t204 gnd 0.278203f
C2173 CSoutput.n3 gnd 0.033334f
C2174 CSoutput.n4 gnd 0.042058f
C2175 CSoutput.t213 gnd 0.278203f
C2176 CSoutput.n5 gnd 0.028744f
C2177 CSoutput.n6 gnd 0.042058f
C2178 CSoutput.t202 gnd 0.278203f
C2179 CSoutput.t199 gnd 0.278203f
C2180 CSoutput.n7 gnd 0.124253f
C2181 CSoutput.n8 gnd 0.042058f
C2182 CSoutput.t211 gnd 0.278203f
C2183 CSoutput.n9 gnd 0.027406f
C2184 CSoutput.n10 gnd 0.042058f
C2185 CSoutput.t192 gnd 0.278203f
C2186 CSoutput.t195 gnd 0.278203f
C2187 CSoutput.n11 gnd 0.124253f
C2188 CSoutput.n12 gnd 0.042058f
C2189 CSoutput.t208 gnd 0.278203f
C2190 CSoutput.n13 gnd 0.028744f
C2191 CSoutput.n14 gnd 0.042058f
C2192 CSoutput.t207 gnd 0.278203f
C2193 CSoutput.t193 gnd 0.278203f
C2194 CSoutput.n15 gnd 0.124253f
C2195 CSoutput.n16 gnd 0.042058f
C2196 CSoutput.t198 gnd 0.278203f
C2197 CSoutput.n17 gnd 0.0307f
C2198 CSoutput.t209 gnd 0.33246f
C2199 CSoutput.t205 gnd 0.278203f
C2200 CSoutput.n18 gnd 0.158623f
C2201 CSoutput.n19 gnd 0.153919f
C2202 CSoutput.n20 gnd 0.178565f
C2203 CSoutput.n21 gnd 0.042058f
C2204 CSoutput.n22 gnd 0.035102f
C2205 CSoutput.n23 gnd 0.124253f
C2206 CSoutput.n24 gnd 0.033837f
C2207 CSoutput.n25 gnd 0.033334f
C2208 CSoutput.n26 gnd 0.042058f
C2209 CSoutput.n27 gnd 0.042058f
C2210 CSoutput.n28 gnd 0.034832f
C2211 CSoutput.n29 gnd 0.029573f
C2212 CSoutput.n30 gnd 0.127019f
C2213 CSoutput.n31 gnd 0.029981f
C2214 CSoutput.n32 gnd 0.042058f
C2215 CSoutput.n33 gnd 0.042058f
C2216 CSoutput.n34 gnd 0.042058f
C2217 CSoutput.n35 gnd 0.034461f
C2218 CSoutput.n36 gnd 0.124253f
C2219 CSoutput.n37 gnd 0.032957f
C2220 CSoutput.n38 gnd 0.034214f
C2221 CSoutput.n39 gnd 0.042058f
C2222 CSoutput.n40 gnd 0.042058f
C2223 CSoutput.n41 gnd 0.035095f
C2224 CSoutput.n42 gnd 0.032077f
C2225 CSoutput.n43 gnd 0.124253f
C2226 CSoutput.n44 gnd 0.03289f
C2227 CSoutput.n45 gnd 0.042058f
C2228 CSoutput.n46 gnd 0.042058f
C2229 CSoutput.n47 gnd 0.042058f
C2230 CSoutput.n48 gnd 0.03289f
C2231 CSoutput.n49 gnd 0.124253f
C2232 CSoutput.n50 gnd 0.032077f
C2233 CSoutput.n51 gnd 0.035095f
C2234 CSoutput.n52 gnd 0.042058f
C2235 CSoutput.n53 gnd 0.042058f
C2236 CSoutput.n54 gnd 0.034214f
C2237 CSoutput.n55 gnd 0.032957f
C2238 CSoutput.n56 gnd 0.124253f
C2239 CSoutput.n57 gnd 0.034461f
C2240 CSoutput.n58 gnd 0.042058f
C2241 CSoutput.n59 gnd 0.042058f
C2242 CSoutput.n60 gnd 0.042058f
C2243 CSoutput.n61 gnd 0.029981f
C2244 CSoutput.n62 gnd 0.127019f
C2245 CSoutput.n63 gnd 0.029573f
C2246 CSoutput.t203 gnd 0.278203f
C2247 CSoutput.n64 gnd 0.124253f
C2248 CSoutput.n65 gnd 0.034832f
C2249 CSoutput.n66 gnd 0.042058f
C2250 CSoutput.n67 gnd 0.042058f
C2251 CSoutput.n68 gnd 0.042058f
C2252 CSoutput.n69 gnd 0.033837f
C2253 CSoutput.n70 gnd 0.124253f
C2254 CSoutput.n71 gnd 0.035102f
C2255 CSoutput.n72 gnd 0.0307f
C2256 CSoutput.n73 gnd 0.042058f
C2257 CSoutput.n74 gnd 0.042058f
C2258 CSoutput.n75 gnd 0.031838f
C2259 CSoutput.n76 gnd 0.018909f
C2260 CSoutput.t212 gnd 0.312581f
C2261 CSoutput.n77 gnd 0.155278f
C2262 CSoutput.n78 gnd 0.635233f
C2263 CSoutput.t159 gnd 0.052461f
C2264 CSoutput.t100 gnd 0.052461f
C2265 CSoutput.n79 gnd 0.406172f
C2266 CSoutput.t147 gnd 0.052461f
C2267 CSoutput.t131 gnd 0.052461f
C2268 CSoutput.n80 gnd 0.405447f
C2269 CSoutput.n81 gnd 0.411529f
C2270 CSoutput.t154 gnd 0.052461f
C2271 CSoutput.t113 gnd 0.052461f
C2272 CSoutput.n82 gnd 0.405447f
C2273 CSoutput.n83 gnd 0.202784f
C2274 CSoutput.t166 gnd 0.052461f
C2275 CSoutput.t125 gnd 0.052461f
C2276 CSoutput.n84 gnd 0.405447f
C2277 CSoutput.n85 gnd 0.202784f
C2278 CSoutput.t104 gnd 0.052461f
C2279 CSoutput.t135 gnd 0.052461f
C2280 CSoutput.n86 gnd 0.405447f
C2281 CSoutput.n87 gnd 0.202784f
C2282 CSoutput.t107 gnd 0.052461f
C2283 CSoutput.t120 gnd 0.052461f
C2284 CSoutput.n88 gnd 0.405447f
C2285 CSoutput.n89 gnd 0.371859f
C2286 CSoutput.t157 gnd 0.052461f
C2287 CSoutput.t155 gnd 0.052461f
C2288 CSoutput.n90 gnd 0.406172f
C2289 CSoutput.t142 gnd 0.052461f
C2290 CSoutput.t105 gnd 0.052461f
C2291 CSoutput.n91 gnd 0.405447f
C2292 CSoutput.n92 gnd 0.411529f
C2293 CSoutput.t101 gnd 0.052461f
C2294 CSoutput.t152 gnd 0.052461f
C2295 CSoutput.n93 gnd 0.405447f
C2296 CSoutput.n94 gnd 0.202784f
C2297 CSoutput.t141 gnd 0.052461f
C2298 CSoutput.t127 gnd 0.052461f
C2299 CSoutput.n95 gnd 0.405447f
C2300 CSoutput.n96 gnd 0.202784f
C2301 CSoutput.t114 gnd 0.052461f
C2302 CSoutput.t162 gnd 0.052461f
C2303 CSoutput.n97 gnd 0.405447f
C2304 CSoutput.n98 gnd 0.202784f
C2305 CSoutput.t140 gnd 0.052461f
C2306 CSoutput.t139 gnd 0.052461f
C2307 CSoutput.n99 gnd 0.405447f
C2308 CSoutput.n100 gnd 0.302402f
C2309 CSoutput.n101 gnd 0.381327f
C2310 CSoutput.t164 gnd 0.052461f
C2311 CSoutput.t163 gnd 0.052461f
C2312 CSoutput.n102 gnd 0.406172f
C2313 CSoutput.t150 gnd 0.052461f
C2314 CSoutput.t111 gnd 0.052461f
C2315 CSoutput.n103 gnd 0.405447f
C2316 CSoutput.n104 gnd 0.411529f
C2317 CSoutput.t109 gnd 0.052461f
C2318 CSoutput.t161 gnd 0.052461f
C2319 CSoutput.n105 gnd 0.405447f
C2320 CSoutput.n106 gnd 0.202784f
C2321 CSoutput.t148 gnd 0.052461f
C2322 CSoutput.t134 gnd 0.052461f
C2323 CSoutput.n107 gnd 0.405447f
C2324 CSoutput.n108 gnd 0.202784f
C2325 CSoutput.t121 gnd 0.052461f
C2326 CSoutput.t169 gnd 0.052461f
C2327 CSoutput.n109 gnd 0.405447f
C2328 CSoutput.n110 gnd 0.202784f
C2329 CSoutput.t146 gnd 0.052461f
C2330 CSoutput.t145 gnd 0.052461f
C2331 CSoutput.n111 gnd 0.405447f
C2332 CSoutput.n112 gnd 0.302402f
C2333 CSoutput.n113 gnd 0.426226f
C2334 CSoutput.n114 gnd 8.723889f
C2335 CSoutput.n116 gnd 0.743994f
C2336 CSoutput.n117 gnd 0.557996f
C2337 CSoutput.n118 gnd 0.743994f
C2338 CSoutput.n119 gnd 0.743994f
C2339 CSoutput.n120 gnd 2.00306f
C2340 CSoutput.n121 gnd 0.743994f
C2341 CSoutput.n122 gnd 0.743994f
C2342 CSoutput.t201 gnd 0.929993f
C2343 CSoutput.n123 gnd 0.743994f
C2344 CSoutput.n124 gnd 0.743994f
C2345 CSoutput.n128 gnd 0.743994f
C2346 CSoutput.n132 gnd 0.743994f
C2347 CSoutput.n133 gnd 0.743994f
C2348 CSoutput.n135 gnd 0.743994f
C2349 CSoutput.n140 gnd 0.743994f
C2350 CSoutput.n142 gnd 0.743994f
C2351 CSoutput.n143 gnd 0.743994f
C2352 CSoutput.n145 gnd 0.743994f
C2353 CSoutput.n146 gnd 0.743994f
C2354 CSoutput.n148 gnd 0.743994f
C2355 CSoutput.t194 gnd 12.4321f
C2356 CSoutput.n150 gnd 0.743994f
C2357 CSoutput.n151 gnd 0.557996f
C2358 CSoutput.n152 gnd 0.743994f
C2359 CSoutput.n153 gnd 0.743994f
C2360 CSoutput.n154 gnd 2.00306f
C2361 CSoutput.n155 gnd 0.743994f
C2362 CSoutput.n156 gnd 0.743994f
C2363 CSoutput.t196 gnd 0.929993f
C2364 CSoutput.n157 gnd 0.743994f
C2365 CSoutput.n158 gnd 0.743994f
C2366 CSoutput.n162 gnd 0.743994f
C2367 CSoutput.n166 gnd 0.743994f
C2368 CSoutput.n167 gnd 0.743994f
C2369 CSoutput.n169 gnd 0.743994f
C2370 CSoutput.n174 gnd 0.743994f
C2371 CSoutput.n176 gnd 0.743994f
C2372 CSoutput.n177 gnd 0.743994f
C2373 CSoutput.n179 gnd 0.743994f
C2374 CSoutput.n180 gnd 0.743994f
C2375 CSoutput.n182 gnd 0.743994f
C2376 CSoutput.n183 gnd 0.557996f
C2377 CSoutput.n185 gnd 0.743994f
C2378 CSoutput.n186 gnd 0.557996f
C2379 CSoutput.n187 gnd 0.743994f
C2380 CSoutput.n188 gnd 0.743994f
C2381 CSoutput.n189 gnd 2.00306f
C2382 CSoutput.n190 gnd 0.743994f
C2383 CSoutput.n191 gnd 0.743994f
C2384 CSoutput.t200 gnd 0.929993f
C2385 CSoutput.n192 gnd 0.743994f
C2386 CSoutput.n193 gnd 2.00306f
C2387 CSoutput.n195 gnd 0.743994f
C2388 CSoutput.n196 gnd 0.743994f
C2389 CSoutput.n198 gnd 0.743994f
C2390 CSoutput.n199 gnd 0.743994f
C2391 CSoutput.t210 gnd 12.2295f
C2392 CSoutput.t206 gnd 12.4321f
C2393 CSoutput.n205 gnd 2.33402f
C2394 CSoutput.n206 gnd 9.50795f
C2395 CSoutput.n207 gnd 9.9058f
C2396 CSoutput.n212 gnd 2.52837f
C2397 CSoutput.n218 gnd 0.743994f
C2398 CSoutput.n220 gnd 0.743994f
C2399 CSoutput.n222 gnd 0.743994f
C2400 CSoutput.n224 gnd 0.743994f
C2401 CSoutput.n226 gnd 0.743994f
C2402 CSoutput.n232 gnd 0.743994f
C2403 CSoutput.n239 gnd 1.36494f
C2404 CSoutput.n240 gnd 1.36494f
C2405 CSoutput.n241 gnd 0.743994f
C2406 CSoutput.n242 gnd 0.743994f
C2407 CSoutput.n244 gnd 0.557996f
C2408 CSoutput.n245 gnd 0.477873f
C2409 CSoutput.n247 gnd 0.557996f
C2410 CSoutput.n248 gnd 0.477873f
C2411 CSoutput.n249 gnd 0.557996f
C2412 CSoutput.n251 gnd 0.743994f
C2413 CSoutput.n253 gnd 2.00306f
C2414 CSoutput.n254 gnd 2.33402f
C2415 CSoutput.n255 gnd 8.74487f
C2416 CSoutput.n257 gnd 0.557996f
C2417 CSoutput.n258 gnd 1.43576f
C2418 CSoutput.n259 gnd 0.557996f
C2419 CSoutput.n261 gnd 0.743994f
C2420 CSoutput.n263 gnd 2.00306f
C2421 CSoutput.n264 gnd 4.36299f
C2422 CSoutput.t99 gnd 0.052461f
C2423 CSoutput.t158 gnd 0.052461f
C2424 CSoutput.n265 gnd 0.406172f
C2425 CSoutput.t130 gnd 0.052461f
C2426 CSoutput.t168 gnd 0.052461f
C2427 CSoutput.n266 gnd 0.405447f
C2428 CSoutput.n267 gnd 0.411529f
C2429 CSoutput.t112 gnd 0.052461f
C2430 CSoutput.t153 gnd 0.052461f
C2431 CSoutput.n268 gnd 0.405447f
C2432 CSoutput.n269 gnd 0.202784f
C2433 CSoutput.t124 gnd 0.052461f
C2434 CSoutput.t165 gnd 0.052461f
C2435 CSoutput.n270 gnd 0.405447f
C2436 CSoutput.n271 gnd 0.202784f
C2437 CSoutput.t149 gnd 0.052461f
C2438 CSoutput.t103 gnd 0.052461f
C2439 CSoutput.n272 gnd 0.405447f
C2440 CSoutput.n273 gnd 0.202784f
C2441 CSoutput.t119 gnd 0.052461f
C2442 CSoutput.t106 gnd 0.052461f
C2443 CSoutput.n274 gnd 0.405447f
C2444 CSoutput.n275 gnd 0.371859f
C2445 CSoutput.t132 gnd 0.052461f
C2446 CSoutput.t133 gnd 0.052461f
C2447 CSoutput.n276 gnd 0.406172f
C2448 CSoutput.t144 gnd 0.052461f
C2449 CSoutput.t102 gnd 0.052461f
C2450 CSoutput.n277 gnd 0.405447f
C2451 CSoutput.n278 gnd 0.411529f
C2452 CSoutput.t129 gnd 0.052461f
C2453 CSoutput.t143 gnd 0.052461f
C2454 CSoutput.n279 gnd 0.405447f
C2455 CSoutput.n280 gnd 0.202784f
C2456 CSoutput.t98 gnd 0.052461f
C2457 CSoutput.t117 gnd 0.052461f
C2458 CSoutput.n281 gnd 0.405447f
C2459 CSoutput.n282 gnd 0.202784f
C2460 CSoutput.t118 gnd 0.052461f
C2461 CSoutput.t160 gnd 0.052461f
C2462 CSoutput.n283 gnd 0.405447f
C2463 CSoutput.n284 gnd 0.202784f
C2464 CSoutput.t115 gnd 0.052461f
C2465 CSoutput.t116 gnd 0.052461f
C2466 CSoutput.n285 gnd 0.405447f
C2467 CSoutput.n286 gnd 0.302402f
C2468 CSoutput.n287 gnd 0.381327f
C2469 CSoutput.t137 gnd 0.052461f
C2470 CSoutput.t138 gnd 0.052461f
C2471 CSoutput.n288 gnd 0.406172f
C2472 CSoutput.t156 gnd 0.052461f
C2473 CSoutput.t110 gnd 0.052461f
C2474 CSoutput.n289 gnd 0.405447f
C2475 CSoutput.n290 gnd 0.411529f
C2476 CSoutput.t136 gnd 0.052461f
C2477 CSoutput.t151 gnd 0.052461f
C2478 CSoutput.n291 gnd 0.405447f
C2479 CSoutput.n292 gnd 0.202784f
C2480 CSoutput.t108 gnd 0.052461f
C2481 CSoutput.t126 gnd 0.052461f
C2482 CSoutput.n293 gnd 0.405447f
C2483 CSoutput.n294 gnd 0.202784f
C2484 CSoutput.t128 gnd 0.052461f
C2485 CSoutput.t167 gnd 0.052461f
C2486 CSoutput.n295 gnd 0.405447f
C2487 CSoutput.n296 gnd 0.202784f
C2488 CSoutput.t122 gnd 0.052461f
C2489 CSoutput.t123 gnd 0.052461f
C2490 CSoutput.n297 gnd 0.405446f
C2491 CSoutput.n298 gnd 0.302403f
C2492 CSoutput.n299 gnd 0.426226f
C2493 CSoutput.n300 gnd 12.0492f
C2494 CSoutput.t46 gnd 0.045903f
C2495 CSoutput.t88 gnd 0.045903f
C2496 CSoutput.n301 gnd 0.406977f
C2497 CSoutput.t93 gnd 0.045903f
C2498 CSoutput.t186 gnd 0.045903f
C2499 CSoutput.n302 gnd 0.405619f
C2500 CSoutput.n303 gnd 0.377962f
C2501 CSoutput.t74 gnd 0.045903f
C2502 CSoutput.t31 gnd 0.045903f
C2503 CSoutput.n304 gnd 0.405619f
C2504 CSoutput.n305 gnd 0.186317f
C2505 CSoutput.t86 gnd 0.045903f
C2506 CSoutput.t92 gnd 0.045903f
C2507 CSoutput.n306 gnd 0.405619f
C2508 CSoutput.n307 gnd 0.186317f
C2509 CSoutput.t41 gnd 0.045903f
C2510 CSoutput.t51 gnd 0.045903f
C2511 CSoutput.n308 gnd 0.405619f
C2512 CSoutput.n309 gnd 0.186317f
C2513 CSoutput.t65 gnd 0.045903f
C2514 CSoutput.t181 gnd 0.045903f
C2515 CSoutput.n310 gnd 0.405619f
C2516 CSoutput.n311 gnd 0.186317f
C2517 CSoutput.t19 gnd 0.045903f
C2518 CSoutput.t58 gnd 0.045903f
C2519 CSoutput.n312 gnd 0.405619f
C2520 CSoutput.n313 gnd 0.186317f
C2521 CSoutput.t176 gnd 0.045903f
C2522 CSoutput.t87 gnd 0.045903f
C2523 CSoutput.n314 gnd 0.405619f
C2524 CSoutput.n315 gnd 0.186317f
C2525 CSoutput.t45 gnd 0.045903f
C2526 CSoutput.t82 gnd 0.045903f
C2527 CSoutput.n316 gnd 0.405619f
C2528 CSoutput.n317 gnd 0.186317f
C2529 CSoutput.t66 gnd 0.045903f
C2530 CSoutput.t85 gnd 0.045903f
C2531 CSoutput.n318 gnd 0.405619f
C2532 CSoutput.n319 gnd 0.343652f
C2533 CSoutput.t50 gnd 0.045903f
C2534 CSoutput.t36 gnd 0.045903f
C2535 CSoutput.n320 gnd 0.406977f
C2536 CSoutput.t0 gnd 0.045903f
C2537 CSoutput.t170 gnd 0.045903f
C2538 CSoutput.n321 gnd 0.405619f
C2539 CSoutput.n322 gnd 0.377962f
C2540 CSoutput.t184 gnd 0.045903f
C2541 CSoutput.t59 gnd 0.045903f
C2542 CSoutput.n323 gnd 0.405619f
C2543 CSoutput.n324 gnd 0.186317f
C2544 CSoutput.t38 gnd 0.045903f
C2545 CSoutput.t15 gnd 0.045903f
C2546 CSoutput.n325 gnd 0.405619f
C2547 CSoutput.n326 gnd 0.186317f
C2548 CSoutput.t71 gnd 0.045903f
C2549 CSoutput.t20 gnd 0.045903f
C2550 CSoutput.n327 gnd 0.405619f
C2551 CSoutput.n328 gnd 0.186317f
C2552 CSoutput.t90 gnd 0.045903f
C2553 CSoutput.t84 gnd 0.045903f
C2554 CSoutput.n329 gnd 0.405619f
C2555 CSoutput.n330 gnd 0.186317f
C2556 CSoutput.t189 gnd 0.045903f
C2557 CSoutput.t190 gnd 0.045903f
C2558 CSoutput.n331 gnd 0.405619f
C2559 CSoutput.n332 gnd 0.186317f
C2560 CSoutput.t35 gnd 0.045903f
C2561 CSoutput.t64 gnd 0.045903f
C2562 CSoutput.n333 gnd 0.405619f
C2563 CSoutput.n334 gnd 0.186317f
C2564 CSoutput.t73 gnd 0.045903f
C2565 CSoutput.t182 gnd 0.045903f
C2566 CSoutput.n335 gnd 0.405619f
C2567 CSoutput.n336 gnd 0.186317f
C2568 CSoutput.t56 gnd 0.045903f
C2569 CSoutput.t30 gnd 0.045903f
C2570 CSoutput.n337 gnd 0.405619f
C2571 CSoutput.n338 gnd 0.28287f
C2572 CSoutput.n339 gnd 0.356786f
C2573 CSoutput.t171 gnd 0.045903f
C2574 CSoutput.t44 gnd 0.045903f
C2575 CSoutput.n340 gnd 0.406977f
C2576 CSoutput.t22 gnd 0.045903f
C2577 CSoutput.t25 gnd 0.045903f
C2578 CSoutput.n341 gnd 0.405619f
C2579 CSoutput.n342 gnd 0.377962f
C2580 CSoutput.t1 gnd 0.045903f
C2581 CSoutput.t95 gnd 0.045903f
C2582 CSoutput.n343 gnd 0.405619f
C2583 CSoutput.n344 gnd 0.186317f
C2584 CSoutput.t81 gnd 0.045903f
C2585 CSoutput.t21 gnd 0.045903f
C2586 CSoutput.n345 gnd 0.405619f
C2587 CSoutput.n346 gnd 0.186317f
C2588 CSoutput.t96 gnd 0.045903f
C2589 CSoutput.t43 gnd 0.045903f
C2590 CSoutput.n347 gnd 0.405619f
C2591 CSoutput.n348 gnd 0.186317f
C2592 CSoutput.t61 gnd 0.045903f
C2593 CSoutput.t69 gnd 0.045903f
C2594 CSoutput.n349 gnd 0.405619f
C2595 CSoutput.n350 gnd 0.186317f
C2596 CSoutput.t33 gnd 0.045903f
C2597 CSoutput.t187 gnd 0.045903f
C2598 CSoutput.n351 gnd 0.405619f
C2599 CSoutput.n352 gnd 0.186317f
C2600 CSoutput.t55 gnd 0.045903f
C2601 CSoutput.t97 gnd 0.045903f
C2602 CSoutput.n353 gnd 0.405619f
C2603 CSoutput.n354 gnd 0.186317f
C2604 CSoutput.t191 gnd 0.045903f
C2605 CSoutput.t7 gnd 0.045903f
C2606 CSoutput.n355 gnd 0.405619f
C2607 CSoutput.n356 gnd 0.186317f
C2608 CSoutput.t9 gnd 0.045903f
C2609 CSoutput.t52 gnd 0.045903f
C2610 CSoutput.n357 gnd 0.405619f
C2611 CSoutput.n358 gnd 0.28287f
C2612 CSoutput.n359 gnd 0.383132f
C2613 CSoutput.n360 gnd 13.1554f
C2614 CSoutput.t4 gnd 0.045903f
C2615 CSoutput.t68 gnd 0.045903f
C2616 CSoutput.n361 gnd 0.406977f
C2617 CSoutput.t34 gnd 0.045903f
C2618 CSoutput.t91 gnd 0.045903f
C2619 CSoutput.n362 gnd 0.405619f
C2620 CSoutput.n363 gnd 0.377962f
C2621 CSoutput.t27 gnd 0.045903f
C2622 CSoutput.t49 gnd 0.045903f
C2623 CSoutput.n364 gnd 0.405619f
C2624 CSoutput.n365 gnd 0.186317f
C2625 CSoutput.t83 gnd 0.045903f
C2626 CSoutput.t89 gnd 0.045903f
C2627 CSoutput.n366 gnd 0.405619f
C2628 CSoutput.n367 gnd 0.186317f
C2629 CSoutput.t23 gnd 0.045903f
C2630 CSoutput.t188 gnd 0.045903f
C2631 CSoutput.n368 gnd 0.405619f
C2632 CSoutput.n369 gnd 0.186317f
C2633 CSoutput.t174 gnd 0.045903f
C2634 CSoutput.t183 gnd 0.045903f
C2635 CSoutput.n370 gnd 0.405619f
C2636 CSoutput.n371 gnd 0.186317f
C2637 CSoutput.t62 gnd 0.045903f
C2638 CSoutput.t60 gnd 0.045903f
C2639 CSoutput.n372 gnd 0.405619f
C2640 CSoutput.n373 gnd 0.186317f
C2641 CSoutput.t40 gnd 0.045903f
C2642 CSoutput.t26 gnd 0.045903f
C2643 CSoutput.n374 gnd 0.405619f
C2644 CSoutput.n375 gnd 0.186317f
C2645 CSoutput.t72 gnd 0.045903f
C2646 CSoutput.t70 gnd 0.045903f
C2647 CSoutput.n376 gnd 0.405619f
C2648 CSoutput.n377 gnd 0.186317f
C2649 CSoutput.t57 gnd 0.045903f
C2650 CSoutput.t67 gnd 0.045903f
C2651 CSoutput.n378 gnd 0.405619f
C2652 CSoutput.n379 gnd 0.343652f
C2653 CSoutput.t179 gnd 0.045903f
C2654 CSoutput.t10 gnd 0.045903f
C2655 CSoutput.n380 gnd 0.406977f
C2656 CSoutput.t48 gnd 0.045903f
C2657 CSoutput.t80 gnd 0.045903f
C2658 CSoutput.n381 gnd 0.405619f
C2659 CSoutput.n382 gnd 0.377962f
C2660 CSoutput.t8 gnd 0.045903f
C2661 CSoutput.t32 gnd 0.045903f
C2662 CSoutput.n383 gnd 0.405619f
C2663 CSoutput.n384 gnd 0.186317f
C2664 CSoutput.t39 gnd 0.045903f
C2665 CSoutput.t6 gnd 0.045903f
C2666 CSoutput.n385 gnd 0.405619f
C2667 CSoutput.n386 gnd 0.186317f
C2668 CSoutput.t63 gnd 0.045903f
C2669 CSoutput.t16 gnd 0.045903f
C2670 CSoutput.n387 gnd 0.405619f
C2671 CSoutput.n388 gnd 0.186317f
C2672 CSoutput.t175 gnd 0.045903f
C2673 CSoutput.t24 gnd 0.045903f
C2674 CSoutput.n389 gnd 0.405619f
C2675 CSoutput.n390 gnd 0.186317f
C2676 CSoutput.t76 gnd 0.045903f
C2677 CSoutput.t47 gnd 0.045903f
C2678 CSoutput.n391 gnd 0.405619f
C2679 CSoutput.n392 gnd 0.186317f
C2680 CSoutput.t18 gnd 0.045903f
C2681 CSoutput.t28 gnd 0.045903f
C2682 CSoutput.n393 gnd 0.405619f
C2683 CSoutput.n394 gnd 0.186317f
C2684 CSoutput.t173 gnd 0.045903f
C2685 CSoutput.t178 gnd 0.045903f
C2686 CSoutput.n395 gnd 0.405619f
C2687 CSoutput.n396 gnd 0.186317f
C2688 CSoutput.t77 gnd 0.045903f
C2689 CSoutput.t12 gnd 0.045903f
C2690 CSoutput.n397 gnd 0.405619f
C2691 CSoutput.n398 gnd 0.28287f
C2692 CSoutput.n399 gnd 0.356786f
C2693 CSoutput.t29 gnd 0.045903f
C2694 CSoutput.t177 gnd 0.045903f
C2695 CSoutput.n400 gnd 0.406977f
C2696 CSoutput.t11 gnd 0.045903f
C2697 CSoutput.t79 gnd 0.045903f
C2698 CSoutput.n401 gnd 0.405619f
C2699 CSoutput.n402 gnd 0.377962f
C2700 CSoutput.t78 gnd 0.045903f
C2701 CSoutput.t37 gnd 0.045903f
C2702 CSoutput.n403 gnd 0.405619f
C2703 CSoutput.n404 gnd 0.186317f
C2704 CSoutput.t180 gnd 0.045903f
C2705 CSoutput.t5 gnd 0.045903f
C2706 CSoutput.n405 gnd 0.405619f
C2707 CSoutput.n406 gnd 0.186317f
C2708 CSoutput.t17 gnd 0.045903f
C2709 CSoutput.t14 gnd 0.045903f
C2710 CSoutput.n407 gnd 0.405619f
C2711 CSoutput.n408 gnd 0.186317f
C2712 CSoutput.t53 gnd 0.045903f
C2713 CSoutput.t54 gnd 0.045903f
C2714 CSoutput.n409 gnd 0.405619f
C2715 CSoutput.n410 gnd 0.186317f
C2716 CSoutput.t172 gnd 0.045903f
C2717 CSoutput.t94 gnd 0.045903f
C2718 CSoutput.n411 gnd 0.405619f
C2719 CSoutput.n412 gnd 0.186317f
C2720 CSoutput.t13 gnd 0.045903f
C2721 CSoutput.t2 gnd 0.045903f
C2722 CSoutput.n413 gnd 0.405619f
C2723 CSoutput.n414 gnd 0.186317f
C2724 CSoutput.t75 gnd 0.045903f
C2725 CSoutput.t3 gnd 0.045903f
C2726 CSoutput.n415 gnd 0.405619f
C2727 CSoutput.n416 gnd 0.186317f
C2728 CSoutput.t185 gnd 0.045903f
C2729 CSoutput.t42 gnd 0.045903f
C2730 CSoutput.n417 gnd 0.405619f
C2731 CSoutput.n418 gnd 0.28287f
C2732 CSoutput.n419 gnd 0.383132f
C2733 CSoutput.n420 gnd 7.86968f
C2734 CSoutput.n421 gnd 13.1099f
C2735 vdd.t106 gnd 0.035972f
C2736 vdd.t102 gnd 0.035972f
C2737 vdd.n0 gnd 0.283719f
C2738 vdd.t99 gnd 0.035972f
C2739 vdd.t86 gnd 0.035972f
C2740 vdd.n1 gnd 0.283251f
C2741 vdd.n2 gnd 0.261211f
C2742 vdd.t84 gnd 0.035972f
C2743 vdd.t120 gnd 0.035972f
C2744 vdd.n3 gnd 0.283251f
C2745 vdd.n4 gnd 0.132104f
C2746 vdd.t122 gnd 0.035972f
C2747 vdd.t229 gnd 0.035972f
C2748 vdd.n5 gnd 0.283251f
C2749 vdd.n6 gnd 0.123956f
C2750 vdd.t80 gnd 0.035972f
C2751 vdd.t108 gnd 0.035972f
C2752 vdd.n7 gnd 0.283719f
C2753 vdd.t231 gnd 0.035972f
C2754 vdd.t104 gnd 0.035972f
C2755 vdd.n8 gnd 0.283251f
C2756 vdd.n9 gnd 0.261212f
C2757 vdd.t88 gnd 0.035972f
C2758 vdd.t125 gnd 0.035972f
C2759 vdd.n10 gnd 0.283251f
C2760 vdd.n11 gnd 0.132104f
C2761 vdd.t112 gnd 0.035972f
C2762 vdd.t95 gnd 0.035972f
C2763 vdd.n12 gnd 0.283251f
C2764 vdd.n13 gnd 0.123956f
C2765 vdd.n14 gnd 0.087634f
C2766 vdd.t91 gnd 0.019985f
C2767 vdd.t131 gnd 0.019985f
C2768 vdd.n15 gnd 0.18395f
C2769 vdd.t1 gnd 0.019985f
C2770 vdd.t2 gnd 0.019985f
C2771 vdd.n16 gnd 0.183412f
C2772 vdd.n17 gnd 0.319194f
C2773 vdd.t0 gnd 0.019985f
C2774 vdd.t116 gnd 0.019985f
C2775 vdd.n18 gnd 0.183412f
C2776 vdd.n19 gnd 0.132055f
C2777 vdd.t129 gnd 0.019985f
C2778 vdd.t126 gnd 0.019985f
C2779 vdd.n20 gnd 0.18395f
C2780 vdd.t92 gnd 0.019985f
C2781 vdd.t89 gnd 0.019985f
C2782 vdd.n21 gnd 0.183412f
C2783 vdd.n22 gnd 0.319194f
C2784 vdd.t127 gnd 0.019985f
C2785 vdd.t128 gnd 0.019985f
C2786 vdd.n23 gnd 0.183412f
C2787 vdd.n24 gnd 0.132055f
C2788 vdd.t90 gnd 0.019985f
C2789 vdd.t123 gnd 0.019985f
C2790 vdd.n25 gnd 0.183412f
C2791 vdd.t130 gnd 0.019985f
C2792 vdd.t93 gnd 0.019985f
C2793 vdd.n26 gnd 0.183412f
C2794 vdd.n27 gnd 20.5189f
C2795 vdd.n28 gnd 7.8839f
C2796 vdd.n29 gnd 0.005451f
C2797 vdd.n30 gnd 0.005058f
C2798 vdd.n31 gnd 0.002798f
C2799 vdd.n32 gnd 0.006424f
C2800 vdd.n33 gnd 0.002718f
C2801 vdd.n34 gnd 0.002878f
C2802 vdd.n35 gnd 0.005058f
C2803 vdd.n36 gnd 0.002718f
C2804 vdd.n37 gnd 0.006424f
C2805 vdd.n38 gnd 0.002878f
C2806 vdd.n39 gnd 0.005058f
C2807 vdd.n40 gnd 0.002718f
C2808 vdd.n41 gnd 0.004818f
C2809 vdd.n42 gnd 0.004833f
C2810 vdd.t135 gnd 0.013802f
C2811 vdd.n43 gnd 0.030709f
C2812 vdd.n44 gnd 0.159815f
C2813 vdd.n45 gnd 0.002718f
C2814 vdd.n46 gnd 0.002878f
C2815 vdd.n47 gnd 0.006424f
C2816 vdd.n48 gnd 0.006424f
C2817 vdd.n49 gnd 0.002878f
C2818 vdd.n50 gnd 0.002718f
C2819 vdd.n51 gnd 0.005058f
C2820 vdd.n52 gnd 0.005058f
C2821 vdd.n53 gnd 0.002718f
C2822 vdd.n54 gnd 0.002878f
C2823 vdd.n55 gnd 0.006424f
C2824 vdd.n56 gnd 0.006424f
C2825 vdd.n57 gnd 0.002878f
C2826 vdd.n58 gnd 0.002718f
C2827 vdd.n59 gnd 0.005058f
C2828 vdd.n60 gnd 0.005058f
C2829 vdd.n61 gnd 0.002718f
C2830 vdd.n62 gnd 0.002878f
C2831 vdd.n63 gnd 0.006424f
C2832 vdd.n64 gnd 0.006424f
C2833 vdd.n65 gnd 0.015188f
C2834 vdd.n66 gnd 0.002798f
C2835 vdd.n67 gnd 0.002718f
C2836 vdd.n68 gnd 0.013073f
C2837 vdd.n69 gnd 0.009127f
C2838 vdd.t216 gnd 0.031975f
C2839 vdd.t184 gnd 0.031975f
C2840 vdd.n70 gnd 0.219757f
C2841 vdd.n71 gnd 0.172805f
C2842 vdd.t222 gnd 0.031975f
C2843 vdd.t162 gnd 0.031975f
C2844 vdd.n72 gnd 0.219757f
C2845 vdd.n73 gnd 0.139453f
C2846 vdd.t204 gnd 0.031975f
C2847 vdd.t174 gnd 0.031975f
C2848 vdd.n74 gnd 0.219757f
C2849 vdd.n75 gnd 0.139453f
C2850 vdd.t220 gnd 0.031975f
C2851 vdd.t207 gnd 0.031975f
C2852 vdd.n76 gnd 0.219757f
C2853 vdd.n77 gnd 0.139453f
C2854 vdd.t149 gnd 0.031975f
C2855 vdd.t143 gnd 0.031975f
C2856 vdd.n78 gnd 0.219757f
C2857 vdd.n79 gnd 0.139453f
C2858 vdd.n80 gnd 0.005451f
C2859 vdd.n81 gnd 0.005058f
C2860 vdd.n82 gnd 0.002798f
C2861 vdd.n83 gnd 0.006424f
C2862 vdd.n84 gnd 0.002718f
C2863 vdd.n85 gnd 0.002878f
C2864 vdd.n86 gnd 0.005058f
C2865 vdd.n87 gnd 0.002718f
C2866 vdd.n88 gnd 0.006424f
C2867 vdd.n89 gnd 0.002878f
C2868 vdd.n90 gnd 0.005058f
C2869 vdd.n91 gnd 0.002718f
C2870 vdd.n92 gnd 0.004818f
C2871 vdd.n93 gnd 0.004833f
C2872 vdd.t154 gnd 0.013802f
C2873 vdd.n94 gnd 0.030709f
C2874 vdd.n95 gnd 0.159815f
C2875 vdd.n96 gnd 0.002718f
C2876 vdd.n97 gnd 0.002878f
C2877 vdd.n98 gnd 0.006424f
C2878 vdd.n99 gnd 0.006424f
C2879 vdd.n100 gnd 0.002878f
C2880 vdd.n101 gnd 0.002718f
C2881 vdd.n102 gnd 0.005058f
C2882 vdd.n103 gnd 0.005058f
C2883 vdd.n104 gnd 0.002718f
C2884 vdd.n105 gnd 0.002878f
C2885 vdd.n106 gnd 0.006424f
C2886 vdd.n107 gnd 0.006424f
C2887 vdd.n108 gnd 0.002878f
C2888 vdd.n109 gnd 0.002718f
C2889 vdd.n110 gnd 0.005058f
C2890 vdd.n111 gnd 0.005058f
C2891 vdd.n112 gnd 0.002718f
C2892 vdd.n113 gnd 0.002878f
C2893 vdd.n114 gnd 0.006424f
C2894 vdd.n115 gnd 0.006424f
C2895 vdd.n116 gnd 0.015188f
C2896 vdd.n117 gnd 0.002798f
C2897 vdd.n118 gnd 0.002718f
C2898 vdd.n119 gnd 0.013073f
C2899 vdd.n120 gnd 0.008841f
C2900 vdd.n121 gnd 0.103754f
C2901 vdd.n122 gnd 0.005451f
C2902 vdd.n123 gnd 0.005058f
C2903 vdd.n124 gnd 0.002798f
C2904 vdd.n125 gnd 0.006424f
C2905 vdd.n126 gnd 0.002718f
C2906 vdd.n127 gnd 0.002878f
C2907 vdd.n128 gnd 0.005058f
C2908 vdd.n129 gnd 0.002718f
C2909 vdd.n130 gnd 0.006424f
C2910 vdd.n131 gnd 0.002878f
C2911 vdd.n132 gnd 0.005058f
C2912 vdd.n133 gnd 0.002718f
C2913 vdd.n134 gnd 0.004818f
C2914 vdd.n135 gnd 0.004833f
C2915 vdd.t186 gnd 0.013802f
C2916 vdd.n136 gnd 0.030709f
C2917 vdd.n137 gnd 0.159815f
C2918 vdd.n138 gnd 0.002718f
C2919 vdd.n139 gnd 0.002878f
C2920 vdd.n140 gnd 0.006424f
C2921 vdd.n141 gnd 0.006424f
C2922 vdd.n142 gnd 0.002878f
C2923 vdd.n143 gnd 0.002718f
C2924 vdd.n144 gnd 0.005058f
C2925 vdd.n145 gnd 0.005058f
C2926 vdd.n146 gnd 0.002718f
C2927 vdd.n147 gnd 0.002878f
C2928 vdd.n148 gnd 0.006424f
C2929 vdd.n149 gnd 0.006424f
C2930 vdd.n150 gnd 0.002878f
C2931 vdd.n151 gnd 0.002718f
C2932 vdd.n152 gnd 0.005058f
C2933 vdd.n153 gnd 0.005058f
C2934 vdd.n154 gnd 0.002718f
C2935 vdd.n155 gnd 0.002878f
C2936 vdd.n156 gnd 0.006424f
C2937 vdd.n157 gnd 0.006424f
C2938 vdd.n158 gnd 0.015188f
C2939 vdd.n159 gnd 0.002798f
C2940 vdd.n160 gnd 0.002718f
C2941 vdd.n161 gnd 0.013073f
C2942 vdd.n162 gnd 0.009127f
C2943 vdd.t182 gnd 0.031975f
C2944 vdd.t201 gnd 0.031975f
C2945 vdd.n163 gnd 0.219757f
C2946 vdd.n164 gnd 0.172805f
C2947 vdd.t147 gnd 0.031975f
C2948 vdd.t180 gnd 0.031975f
C2949 vdd.n165 gnd 0.219757f
C2950 vdd.n166 gnd 0.139453f
C2951 vdd.t200 gnd 0.031975f
C2952 vdd.t133 gnd 0.031975f
C2953 vdd.n167 gnd 0.219757f
C2954 vdd.n168 gnd 0.139453f
C2955 vdd.t141 gnd 0.031975f
C2956 vdd.t168 gnd 0.031975f
C2957 vdd.n169 gnd 0.219757f
C2958 vdd.n170 gnd 0.139453f
C2959 vdd.t218 gnd 0.031975f
C2960 vdd.t165 gnd 0.031975f
C2961 vdd.n171 gnd 0.219757f
C2962 vdd.n172 gnd 0.139453f
C2963 vdd.n173 gnd 0.005451f
C2964 vdd.n174 gnd 0.005058f
C2965 vdd.n175 gnd 0.002798f
C2966 vdd.n176 gnd 0.006424f
C2967 vdd.n177 gnd 0.002718f
C2968 vdd.n178 gnd 0.002878f
C2969 vdd.n179 gnd 0.005058f
C2970 vdd.n180 gnd 0.002718f
C2971 vdd.n181 gnd 0.006424f
C2972 vdd.n182 gnd 0.002878f
C2973 vdd.n183 gnd 0.005058f
C2974 vdd.n184 gnd 0.002718f
C2975 vdd.n185 gnd 0.004818f
C2976 vdd.n186 gnd 0.004833f
C2977 vdd.t166 gnd 0.013802f
C2978 vdd.n187 gnd 0.030709f
C2979 vdd.n188 gnd 0.159815f
C2980 vdd.n189 gnd 0.002718f
C2981 vdd.n190 gnd 0.002878f
C2982 vdd.n191 gnd 0.006424f
C2983 vdd.n192 gnd 0.006424f
C2984 vdd.n193 gnd 0.002878f
C2985 vdd.n194 gnd 0.002718f
C2986 vdd.n195 gnd 0.005058f
C2987 vdd.n196 gnd 0.005058f
C2988 vdd.n197 gnd 0.002718f
C2989 vdd.n198 gnd 0.002878f
C2990 vdd.n199 gnd 0.006424f
C2991 vdd.n200 gnd 0.006424f
C2992 vdd.n201 gnd 0.002878f
C2993 vdd.n202 gnd 0.002718f
C2994 vdd.n203 gnd 0.005058f
C2995 vdd.n204 gnd 0.005058f
C2996 vdd.n205 gnd 0.002718f
C2997 vdd.n206 gnd 0.002878f
C2998 vdd.n207 gnd 0.006424f
C2999 vdd.n208 gnd 0.006424f
C3000 vdd.n209 gnd 0.015188f
C3001 vdd.n210 gnd 0.002798f
C3002 vdd.n211 gnd 0.002718f
C3003 vdd.n212 gnd 0.013073f
C3004 vdd.n213 gnd 0.008841f
C3005 vdd.n214 gnd 0.061723f
C3006 vdd.n215 gnd 0.222404f
C3007 vdd.n216 gnd 0.005451f
C3008 vdd.n217 gnd 0.005058f
C3009 vdd.n218 gnd 0.002798f
C3010 vdd.n219 gnd 0.006424f
C3011 vdd.n220 gnd 0.002718f
C3012 vdd.n221 gnd 0.002878f
C3013 vdd.n222 gnd 0.005058f
C3014 vdd.n223 gnd 0.002718f
C3015 vdd.n224 gnd 0.006424f
C3016 vdd.n225 gnd 0.002878f
C3017 vdd.n226 gnd 0.005058f
C3018 vdd.n227 gnd 0.002718f
C3019 vdd.n228 gnd 0.004818f
C3020 vdd.n229 gnd 0.004833f
C3021 vdd.t191 gnd 0.013802f
C3022 vdd.n230 gnd 0.030709f
C3023 vdd.n231 gnd 0.159815f
C3024 vdd.n232 gnd 0.002718f
C3025 vdd.n233 gnd 0.002878f
C3026 vdd.n234 gnd 0.006424f
C3027 vdd.n235 gnd 0.006424f
C3028 vdd.n236 gnd 0.002878f
C3029 vdd.n237 gnd 0.002718f
C3030 vdd.n238 gnd 0.005058f
C3031 vdd.n239 gnd 0.005058f
C3032 vdd.n240 gnd 0.002718f
C3033 vdd.n241 gnd 0.002878f
C3034 vdd.n242 gnd 0.006424f
C3035 vdd.n243 gnd 0.006424f
C3036 vdd.n244 gnd 0.002878f
C3037 vdd.n245 gnd 0.002718f
C3038 vdd.n246 gnd 0.005058f
C3039 vdd.n247 gnd 0.005058f
C3040 vdd.n248 gnd 0.002718f
C3041 vdd.n249 gnd 0.002878f
C3042 vdd.n250 gnd 0.006424f
C3043 vdd.n251 gnd 0.006424f
C3044 vdd.n252 gnd 0.015188f
C3045 vdd.n253 gnd 0.002798f
C3046 vdd.n254 gnd 0.002718f
C3047 vdd.n255 gnd 0.013073f
C3048 vdd.n256 gnd 0.009127f
C3049 vdd.t192 gnd 0.031975f
C3050 vdd.t213 gnd 0.031975f
C3051 vdd.n257 gnd 0.219757f
C3052 vdd.n258 gnd 0.172805f
C3053 vdd.t159 gnd 0.031975f
C3054 vdd.t190 gnd 0.031975f
C3055 vdd.n259 gnd 0.219757f
C3056 vdd.n260 gnd 0.139453f
C3057 vdd.t209 gnd 0.031975f
C3058 vdd.t157 gnd 0.031975f
C3059 vdd.n261 gnd 0.219757f
C3060 vdd.n262 gnd 0.139453f
C3061 vdd.t177 gnd 0.031975f
C3062 vdd.t179 gnd 0.031975f
C3063 vdd.n263 gnd 0.219757f
C3064 vdd.n264 gnd 0.139453f
C3065 vdd.t226 gnd 0.031975f
C3066 vdd.t172 gnd 0.031975f
C3067 vdd.n265 gnd 0.219757f
C3068 vdd.n266 gnd 0.139453f
C3069 vdd.n267 gnd 0.005451f
C3070 vdd.n268 gnd 0.005058f
C3071 vdd.n269 gnd 0.002798f
C3072 vdd.n270 gnd 0.006424f
C3073 vdd.n271 gnd 0.002718f
C3074 vdd.n272 gnd 0.002878f
C3075 vdd.n273 gnd 0.005058f
C3076 vdd.n274 gnd 0.002718f
C3077 vdd.n275 gnd 0.006424f
C3078 vdd.n276 gnd 0.002878f
C3079 vdd.n277 gnd 0.005058f
C3080 vdd.n278 gnd 0.002718f
C3081 vdd.n279 gnd 0.004818f
C3082 vdd.n280 gnd 0.004833f
C3083 vdd.t173 gnd 0.013802f
C3084 vdd.n281 gnd 0.030709f
C3085 vdd.n282 gnd 0.159815f
C3086 vdd.n283 gnd 0.002718f
C3087 vdd.n284 gnd 0.002878f
C3088 vdd.n285 gnd 0.006424f
C3089 vdd.n286 gnd 0.006424f
C3090 vdd.n287 gnd 0.002878f
C3091 vdd.n288 gnd 0.002718f
C3092 vdd.n289 gnd 0.005058f
C3093 vdd.n290 gnd 0.005058f
C3094 vdd.n291 gnd 0.002718f
C3095 vdd.n292 gnd 0.002878f
C3096 vdd.n293 gnd 0.006424f
C3097 vdd.n294 gnd 0.006424f
C3098 vdd.n295 gnd 0.002878f
C3099 vdd.n296 gnd 0.002718f
C3100 vdd.n297 gnd 0.005058f
C3101 vdd.n298 gnd 0.005058f
C3102 vdd.n299 gnd 0.002718f
C3103 vdd.n300 gnd 0.002878f
C3104 vdd.n301 gnd 0.006424f
C3105 vdd.n302 gnd 0.006424f
C3106 vdd.n303 gnd 0.015188f
C3107 vdd.n304 gnd 0.002798f
C3108 vdd.n305 gnd 0.002718f
C3109 vdd.n306 gnd 0.013073f
C3110 vdd.n307 gnd 0.008841f
C3111 vdd.n308 gnd 0.061723f
C3112 vdd.n309 gnd 0.244429f
C3113 vdd.n310 gnd 0.009898f
C3114 vdd.n311 gnd 0.009898f
C3115 vdd.n312 gnd 0.007994f
C3116 vdd.n313 gnd 0.007994f
C3117 vdd.n314 gnd 0.009932f
C3118 vdd.n315 gnd 0.009932f
C3119 vdd.t199 gnd 0.507488f
C3120 vdd.n316 gnd 0.009932f
C3121 vdd.n317 gnd 0.009932f
C3122 vdd.n318 gnd 0.009932f
C3123 vdd.t140 gnd 0.507488f
C3124 vdd.n319 gnd 0.009932f
C3125 vdd.n320 gnd 0.009932f
C3126 vdd.n321 gnd 0.009932f
C3127 vdd.n322 gnd 0.009932f
C3128 vdd.n323 gnd 0.007994f
C3129 vdd.n324 gnd 0.009932f
C3130 vdd.n325 gnd 0.817056f
C3131 vdd.n326 gnd 0.009932f
C3132 vdd.n327 gnd 0.009932f
C3133 vdd.n328 gnd 0.009932f
C3134 vdd.n329 gnd 0.695259f
C3135 vdd.n330 gnd 0.009932f
C3136 vdd.n331 gnd 0.009932f
C3137 vdd.n332 gnd 0.009932f
C3138 vdd.n333 gnd 0.009932f
C3139 vdd.n334 gnd 0.009932f
C3140 vdd.n335 gnd 0.007994f
C3141 vdd.n336 gnd 0.009932f
C3142 vdd.t142 gnd 0.507488f
C3143 vdd.n337 gnd 0.009932f
C3144 vdd.n338 gnd 0.009932f
C3145 vdd.n339 gnd 0.009932f
C3146 vdd.n340 gnd 1.01498f
C3147 vdd.n341 gnd 0.009932f
C3148 vdd.n342 gnd 0.009932f
C3149 vdd.n343 gnd 0.009932f
C3150 vdd.n344 gnd 0.009932f
C3151 vdd.n345 gnd 0.009932f
C3152 vdd.n346 gnd 0.007994f
C3153 vdd.n347 gnd 0.009932f
C3154 vdd.n348 gnd 0.009932f
C3155 vdd.n349 gnd 0.009932f
C3156 vdd.n350 gnd 0.023405f
C3157 vdd.n351 gnd 2.33445f
C3158 vdd.n352 gnd 0.023771f
C3159 vdd.n353 gnd 0.009932f
C3160 vdd.n354 gnd 0.009932f
C3161 vdd.n356 gnd 0.009932f
C3162 vdd.n357 gnd 0.009932f
C3163 vdd.n358 gnd 0.007994f
C3164 vdd.n359 gnd 0.007994f
C3165 vdd.n360 gnd 0.009932f
C3166 vdd.n361 gnd 0.009932f
C3167 vdd.n362 gnd 0.009932f
C3168 vdd.n363 gnd 0.009932f
C3169 vdd.n364 gnd 0.009932f
C3170 vdd.n365 gnd 0.009932f
C3171 vdd.n366 gnd 0.007994f
C3172 vdd.n368 gnd 0.009932f
C3173 vdd.n369 gnd 0.009932f
C3174 vdd.n370 gnd 0.009932f
C3175 vdd.n371 gnd 0.009932f
C3176 vdd.n372 gnd 0.009932f
C3177 vdd.n373 gnd 0.007994f
C3178 vdd.n375 gnd 0.009932f
C3179 vdd.n376 gnd 0.009932f
C3180 vdd.n377 gnd 0.009932f
C3181 vdd.n378 gnd 0.009932f
C3182 vdd.n379 gnd 0.009932f
C3183 vdd.n380 gnd 0.007994f
C3184 vdd.n382 gnd 0.009932f
C3185 vdd.n383 gnd 0.009932f
C3186 vdd.n384 gnd 0.009932f
C3187 vdd.n385 gnd 0.009932f
C3188 vdd.n386 gnd 0.006675f
C3189 vdd.t14 gnd 0.122186f
C3190 vdd.t13 gnd 0.130584f
C3191 vdd.t11 gnd 0.159574f
C3192 vdd.n387 gnd 0.204551f
C3193 vdd.n388 gnd 0.172659f
C3194 vdd.n390 gnd 0.009932f
C3195 vdd.n391 gnd 0.009932f
C3196 vdd.n392 gnd 0.007994f
C3197 vdd.n393 gnd 0.009932f
C3198 vdd.n395 gnd 0.009932f
C3199 vdd.n396 gnd 0.009932f
C3200 vdd.n397 gnd 0.009932f
C3201 vdd.n398 gnd 0.009932f
C3202 vdd.n399 gnd 0.007994f
C3203 vdd.n401 gnd 0.009932f
C3204 vdd.n402 gnd 0.009932f
C3205 vdd.n403 gnd 0.009932f
C3206 vdd.n404 gnd 0.009932f
C3207 vdd.n405 gnd 0.009932f
C3208 vdd.n406 gnd 0.007994f
C3209 vdd.n408 gnd 0.009932f
C3210 vdd.n409 gnd 0.009932f
C3211 vdd.n410 gnd 0.009932f
C3212 vdd.n411 gnd 0.009932f
C3213 vdd.n412 gnd 0.009932f
C3214 vdd.n413 gnd 0.007994f
C3215 vdd.n415 gnd 0.009932f
C3216 vdd.n416 gnd 0.009932f
C3217 vdd.n417 gnd 0.009932f
C3218 vdd.n418 gnd 0.009932f
C3219 vdd.n419 gnd 0.009932f
C3220 vdd.n420 gnd 0.007994f
C3221 vdd.n422 gnd 0.009932f
C3222 vdd.n423 gnd 0.009932f
C3223 vdd.n424 gnd 0.009932f
C3224 vdd.n425 gnd 0.009932f
C3225 vdd.n426 gnd 0.007914f
C3226 vdd.t75 gnd 0.122186f
C3227 vdd.t74 gnd 0.130584f
C3228 vdd.t73 gnd 0.159574f
C3229 vdd.n427 gnd 0.204551f
C3230 vdd.n428 gnd 0.172659f
C3231 vdd.n430 gnd 0.009932f
C3232 vdd.n431 gnd 0.009932f
C3233 vdd.n432 gnd 0.007994f
C3234 vdd.n433 gnd 0.009932f
C3235 vdd.n435 gnd 0.009932f
C3236 vdd.n436 gnd 0.009932f
C3237 vdd.n437 gnd 0.009932f
C3238 vdd.n438 gnd 0.009932f
C3239 vdd.n439 gnd 0.007994f
C3240 vdd.n441 gnd 0.009932f
C3241 vdd.n442 gnd 0.009932f
C3242 vdd.n443 gnd 0.009932f
C3243 vdd.n444 gnd 0.009932f
C3244 vdd.n445 gnd 0.009932f
C3245 vdd.n446 gnd 0.007994f
C3246 vdd.n448 gnd 0.009932f
C3247 vdd.n449 gnd 0.009932f
C3248 vdd.n450 gnd 0.009932f
C3249 vdd.n451 gnd 0.009932f
C3250 vdd.n452 gnd 0.009932f
C3251 vdd.n453 gnd 0.007994f
C3252 vdd.n455 gnd 0.009932f
C3253 vdd.n456 gnd 0.009932f
C3254 vdd.n457 gnd 0.009932f
C3255 vdd.n458 gnd 0.009932f
C3256 vdd.n459 gnd 0.009932f
C3257 vdd.n460 gnd 0.007994f
C3258 vdd.n462 gnd 0.009932f
C3259 vdd.n463 gnd 0.009932f
C3260 vdd.n464 gnd 0.009932f
C3261 vdd.n465 gnd 0.009932f
C3262 vdd.n466 gnd 0.009932f
C3263 vdd.n467 gnd 0.009932f
C3264 vdd.n468 gnd 0.007994f
C3265 vdd.n469 gnd 0.009932f
C3266 vdd.n470 gnd 0.009932f
C3267 vdd.n471 gnd 0.007994f
C3268 vdd.n472 gnd 0.009932f
C3269 vdd.n473 gnd 0.009932f
C3270 vdd.n474 gnd 0.007994f
C3271 vdd.n475 gnd 0.009932f
C3272 vdd.n476 gnd 0.007994f
C3273 vdd.n477 gnd 0.009932f
C3274 vdd.n478 gnd 0.007994f
C3275 vdd.n479 gnd 0.009932f
C3276 vdd.n480 gnd 0.009932f
C3277 vdd.t161 gnd 0.507488f
C3278 vdd.n481 gnd 0.543012f
C3279 vdd.n482 gnd 0.009932f
C3280 vdd.n483 gnd 0.007994f
C3281 vdd.n484 gnd 0.009932f
C3282 vdd.n485 gnd 0.007994f
C3283 vdd.n486 gnd 0.009932f
C3284 vdd.t146 gnd 0.507488f
C3285 vdd.n487 gnd 0.009932f
C3286 vdd.n488 gnd 0.007994f
C3287 vdd.n489 gnd 0.009932f
C3288 vdd.n490 gnd 0.007994f
C3289 vdd.n491 gnd 0.009932f
C3290 vdd.n492 gnd 0.796757f
C3291 vdd.n493 gnd 0.84243f
C3292 vdd.t183 gnd 0.507488f
C3293 vdd.n494 gnd 0.009932f
C3294 vdd.n495 gnd 0.007994f
C3295 vdd.n496 gnd 0.009932f
C3296 vdd.n497 gnd 0.007994f
C3297 vdd.n498 gnd 0.009932f
C3298 vdd.n499 gnd 0.624211f
C3299 vdd.n500 gnd 0.009932f
C3300 vdd.n501 gnd 0.007994f
C3301 vdd.n502 gnd 0.009932f
C3302 vdd.n503 gnd 0.007994f
C3303 vdd.n504 gnd 0.009932f
C3304 vdd.n505 gnd 1.01498f
C3305 vdd.t134 gnd 0.507488f
C3306 vdd.n506 gnd 0.009932f
C3307 vdd.n507 gnd 0.007994f
C3308 vdd.n508 gnd 0.009932f
C3309 vdd.n509 gnd 0.007994f
C3310 vdd.n510 gnd 0.009932f
C3311 vdd.n511 gnd 0.543012f
C3312 vdd.n512 gnd 0.009932f
C3313 vdd.n513 gnd 0.007994f
C3314 vdd.n514 gnd 0.023771f
C3315 vdd.n515 gnd 0.023771f
C3316 vdd.n516 gnd 7.26723f
C3317 vdd.t16 gnd 0.507488f
C3318 vdd.n517 gnd 0.023771f
C3319 vdd.n518 gnd 0.008541f
C3320 vdd.n519 gnd 0.007994f
C3321 vdd.n524 gnd 0.006356f
C3322 vdd.n525 gnd 0.007994f
C3323 vdd.n526 gnd 0.009932f
C3324 vdd.n527 gnd 0.009932f
C3325 vdd.n528 gnd 0.009932f
C3326 vdd.n529 gnd 0.009932f
C3327 vdd.n530 gnd 0.009932f
C3328 vdd.n531 gnd 0.007994f
C3329 vdd.n532 gnd 0.009932f
C3330 vdd.n533 gnd 0.009932f
C3331 vdd.n534 gnd 0.009932f
C3332 vdd.n535 gnd 0.009932f
C3333 vdd.n536 gnd 0.009932f
C3334 vdd.n537 gnd 0.007994f
C3335 vdd.n538 gnd 0.009932f
C3336 vdd.n539 gnd 0.009932f
C3337 vdd.n540 gnd 0.009932f
C3338 vdd.n541 gnd 0.009932f
C3339 vdd.n542 gnd 0.009932f
C3340 vdd.t20 gnd 0.122186f
C3341 vdd.t21 gnd 0.130584f
C3342 vdd.t19 gnd 0.159574f
C3343 vdd.n543 gnd 0.204551f
C3344 vdd.n544 gnd 0.17186f
C3345 vdd.n545 gnd 0.016307f
C3346 vdd.n546 gnd 0.009932f
C3347 vdd.n547 gnd 0.009932f
C3348 vdd.n548 gnd 0.009932f
C3349 vdd.n549 gnd 0.009932f
C3350 vdd.n550 gnd 0.009932f
C3351 vdd.n551 gnd 0.007994f
C3352 vdd.n552 gnd 0.009932f
C3353 vdd.n553 gnd 0.009932f
C3354 vdd.n554 gnd 0.009932f
C3355 vdd.n555 gnd 0.009932f
C3356 vdd.n556 gnd 0.009932f
C3357 vdd.n557 gnd 0.007994f
C3358 vdd.n558 gnd 0.009932f
C3359 vdd.n559 gnd 0.009932f
C3360 vdd.n560 gnd 0.009932f
C3361 vdd.n561 gnd 0.009932f
C3362 vdd.n562 gnd 0.009932f
C3363 vdd.n563 gnd 0.007994f
C3364 vdd.n564 gnd 0.009932f
C3365 vdd.n565 gnd 0.009932f
C3366 vdd.n566 gnd 0.009932f
C3367 vdd.n567 gnd 0.009932f
C3368 vdd.n568 gnd 0.009932f
C3369 vdd.n569 gnd 0.007994f
C3370 vdd.n570 gnd 0.009932f
C3371 vdd.n571 gnd 0.009932f
C3372 vdd.n572 gnd 0.009932f
C3373 vdd.n573 gnd 0.009932f
C3374 vdd.n574 gnd 0.009932f
C3375 vdd.n575 gnd 0.007994f
C3376 vdd.n576 gnd 0.009932f
C3377 vdd.n577 gnd 0.009932f
C3378 vdd.n578 gnd 0.009932f
C3379 vdd.n579 gnd 0.007914f
C3380 vdd.t17 gnd 0.122186f
C3381 vdd.t18 gnd 0.130584f
C3382 vdd.t15 gnd 0.159574f
C3383 vdd.n580 gnd 0.204551f
C3384 vdd.n581 gnd 0.17186f
C3385 vdd.n582 gnd 0.009932f
C3386 vdd.n583 gnd 0.007994f
C3387 vdd.n585 gnd 0.009932f
C3388 vdd.n587 gnd 0.009932f
C3389 vdd.n588 gnd 0.009932f
C3390 vdd.n589 gnd 0.007994f
C3391 vdd.n590 gnd 0.009932f
C3392 vdd.n591 gnd 0.009932f
C3393 vdd.n592 gnd 0.009932f
C3394 vdd.n593 gnd 0.009932f
C3395 vdd.n594 gnd 0.009932f
C3396 vdd.n595 gnd 0.007994f
C3397 vdd.n596 gnd 0.009932f
C3398 vdd.n597 gnd 0.009932f
C3399 vdd.n598 gnd 0.009932f
C3400 vdd.n599 gnd 0.009932f
C3401 vdd.n600 gnd 0.009932f
C3402 vdd.n601 gnd 0.007994f
C3403 vdd.n602 gnd 0.009932f
C3404 vdd.n603 gnd 0.009932f
C3405 vdd.n604 gnd 0.009932f
C3406 vdd.n605 gnd 0.006356f
C3407 vdd.n610 gnd 0.006754f
C3408 vdd.n611 gnd 0.006754f
C3409 vdd.n612 gnd 0.006754f
C3410 vdd.n613 gnd 6.99319f
C3411 vdd.n614 gnd 0.006754f
C3412 vdd.n615 gnd 0.006754f
C3413 vdd.n616 gnd 0.006754f
C3414 vdd.n618 gnd 0.006754f
C3415 vdd.n619 gnd 0.006754f
C3416 vdd.n621 gnd 0.006754f
C3417 vdd.n622 gnd 0.004916f
C3418 vdd.n624 gnd 0.006754f
C3419 vdd.t56 gnd 0.272911f
C3420 vdd.t55 gnd 0.279359f
C3421 vdd.t54 gnd 0.178167f
C3422 vdd.n625 gnd 0.096289f
C3423 vdd.n626 gnd 0.054619f
C3424 vdd.n627 gnd 0.009652f
C3425 vdd.n628 gnd 0.015784f
C3426 vdd.n630 gnd 0.006754f
C3427 vdd.n631 gnd 0.690184f
C3428 vdd.n632 gnd 0.014962f
C3429 vdd.n633 gnd 0.014962f
C3430 vdd.n634 gnd 0.006754f
C3431 vdd.n635 gnd 0.016025f
C3432 vdd.n636 gnd 0.006754f
C3433 vdd.n637 gnd 0.006754f
C3434 vdd.n638 gnd 0.006754f
C3435 vdd.n639 gnd 0.006754f
C3436 vdd.n640 gnd 0.006754f
C3437 vdd.n642 gnd 0.006754f
C3438 vdd.n643 gnd 0.006754f
C3439 vdd.n645 gnd 0.006754f
C3440 vdd.n646 gnd 0.006754f
C3441 vdd.n648 gnd 0.006754f
C3442 vdd.n649 gnd 0.006754f
C3443 vdd.n651 gnd 0.006754f
C3444 vdd.n652 gnd 0.006754f
C3445 vdd.n654 gnd 0.006754f
C3446 vdd.n655 gnd 0.006754f
C3447 vdd.n657 gnd 0.006754f
C3448 vdd.n658 gnd 0.004916f
C3449 vdd.n660 gnd 0.006754f
C3450 vdd.t49 gnd 0.272911f
C3451 vdd.t48 gnd 0.279359f
C3452 vdd.t46 gnd 0.178167f
C3453 vdd.n661 gnd 0.096289f
C3454 vdd.n662 gnd 0.054619f
C3455 vdd.n663 gnd 0.009652f
C3456 vdd.n664 gnd 0.006754f
C3457 vdd.n665 gnd 0.006754f
C3458 vdd.t47 gnd 0.345092f
C3459 vdd.n666 gnd 0.006754f
C3460 vdd.n667 gnd 0.006754f
C3461 vdd.n668 gnd 0.006754f
C3462 vdd.n669 gnd 0.006754f
C3463 vdd.n670 gnd 0.006754f
C3464 vdd.n671 gnd 0.690184f
C3465 vdd.n672 gnd 0.006754f
C3466 vdd.n673 gnd 0.006754f
C3467 vdd.n674 gnd 0.603911f
C3468 vdd.n675 gnd 0.006754f
C3469 vdd.n676 gnd 0.006754f
C3470 vdd.n677 gnd 0.005959f
C3471 vdd.n678 gnd 0.006754f
C3472 vdd.n679 gnd 0.608986f
C3473 vdd.n680 gnd 0.006754f
C3474 vdd.n681 gnd 0.006754f
C3475 vdd.n682 gnd 0.006754f
C3476 vdd.n683 gnd 0.006754f
C3477 vdd.n684 gnd 0.006754f
C3478 vdd.n685 gnd 0.690184f
C3479 vdd.n686 gnd 0.006754f
C3480 vdd.n687 gnd 0.006754f
C3481 vdd.t30 gnd 0.309568f
C3482 vdd.t114 gnd 0.081198f
C3483 vdd.n688 gnd 0.006754f
C3484 vdd.n689 gnd 0.006754f
C3485 vdd.n690 gnd 0.006754f
C3486 vdd.t82 gnd 0.345092f
C3487 vdd.n691 gnd 0.006754f
C3488 vdd.n692 gnd 0.006754f
C3489 vdd.n693 gnd 0.006754f
C3490 vdd.n694 gnd 0.006754f
C3491 vdd.n695 gnd 0.006754f
C3492 vdd.t113 gnd 0.345092f
C3493 vdd.n696 gnd 0.006754f
C3494 vdd.n697 gnd 0.006754f
C3495 vdd.n698 gnd 0.573462f
C3496 vdd.n699 gnd 0.006754f
C3497 vdd.n700 gnd 0.006754f
C3498 vdd.n701 gnd 0.006754f
C3499 vdd.n702 gnd 0.421215f
C3500 vdd.n703 gnd 0.006754f
C3501 vdd.n704 gnd 0.006754f
C3502 vdd.t107 gnd 0.345092f
C3503 vdd.n705 gnd 0.006754f
C3504 vdd.n706 gnd 0.006754f
C3505 vdd.n707 gnd 0.006754f
C3506 vdd.n708 gnd 0.573462f
C3507 vdd.n709 gnd 0.006754f
C3508 vdd.n710 gnd 0.006754f
C3509 vdd.t96 gnd 0.294343f
C3510 vdd.t79 gnd 0.268969f
C3511 vdd.n711 gnd 0.006754f
C3512 vdd.n712 gnd 0.006754f
C3513 vdd.n713 gnd 0.006754f
C3514 vdd.t103 gnd 0.345092f
C3515 vdd.n714 gnd 0.006754f
C3516 vdd.n715 gnd 0.006754f
C3517 vdd.t118 gnd 0.345092f
C3518 vdd.n716 gnd 0.006754f
C3519 vdd.n717 gnd 0.006754f
C3520 vdd.n718 gnd 0.006754f
C3521 vdd.t97 gnd 0.253744f
C3522 vdd.n719 gnd 0.006754f
C3523 vdd.n720 gnd 0.006754f
C3524 vdd.n721 gnd 0.588686f
C3525 vdd.n722 gnd 0.006754f
C3526 vdd.n723 gnd 0.006754f
C3527 vdd.n724 gnd 0.006754f
C3528 vdd.n725 gnd 0.690184f
C3529 vdd.n726 gnd 0.006754f
C3530 vdd.n727 gnd 0.006754f
C3531 vdd.t230 gnd 0.309568f
C3532 vdd.n728 gnd 0.43644f
C3533 vdd.n729 gnd 0.006754f
C3534 vdd.n730 gnd 0.006754f
C3535 vdd.n731 gnd 0.006754f
C3536 vdd.t124 gnd 0.345092f
C3537 vdd.n732 gnd 0.006754f
C3538 vdd.n733 gnd 0.006754f
C3539 vdd.n734 gnd 0.006754f
C3540 vdd.n735 gnd 0.006754f
C3541 vdd.n736 gnd 0.006754f
C3542 vdd.t87 gnd 0.690184f
C3543 vdd.n737 gnd 0.006754f
C3544 vdd.n738 gnd 0.006754f
C3545 vdd.t51 gnd 0.345092f
C3546 vdd.n739 gnd 0.006754f
C3547 vdd.n740 gnd 0.016025f
C3548 vdd.n741 gnd 0.016025f
C3549 vdd.t94 gnd 0.649585f
C3550 vdd.n742 gnd 0.014962f
C3551 vdd.n743 gnd 0.014962f
C3552 vdd.n744 gnd 0.016025f
C3553 vdd.n745 gnd 0.006754f
C3554 vdd.n746 gnd 0.006754f
C3555 vdd.t121 gnd 0.649585f
C3556 vdd.n764 gnd 0.016025f
C3557 vdd.n782 gnd 0.014962f
C3558 vdd.n783 gnd 0.006754f
C3559 vdd.n784 gnd 0.014962f
C3560 vdd.t69 gnd 0.272911f
C3561 vdd.t68 gnd 0.279359f
C3562 vdd.t67 gnd 0.178167f
C3563 vdd.n785 gnd 0.096289f
C3564 vdd.n786 gnd 0.054619f
C3565 vdd.n787 gnd 0.015784f
C3566 vdd.n788 gnd 0.006754f
C3567 vdd.t119 gnd 0.690184f
C3568 vdd.n789 gnd 0.014962f
C3569 vdd.n790 gnd 0.006754f
C3570 vdd.n791 gnd 0.016025f
C3571 vdd.n792 gnd 0.006754f
C3572 vdd.t45 gnd 0.272911f
C3573 vdd.t44 gnd 0.279359f
C3574 vdd.t42 gnd 0.178167f
C3575 vdd.n793 gnd 0.096289f
C3576 vdd.n794 gnd 0.054619f
C3577 vdd.n795 gnd 0.009652f
C3578 vdd.n796 gnd 0.006754f
C3579 vdd.n797 gnd 0.006754f
C3580 vdd.t43 gnd 0.345092f
C3581 vdd.n798 gnd 0.006754f
C3582 vdd.n799 gnd 0.006754f
C3583 vdd.n800 gnd 0.006754f
C3584 vdd.n801 gnd 0.006754f
C3585 vdd.n802 gnd 0.006754f
C3586 vdd.n803 gnd 0.006754f
C3587 vdd.n804 gnd 0.690184f
C3588 vdd.n805 gnd 0.006754f
C3589 vdd.n806 gnd 0.006754f
C3590 vdd.t83 gnd 0.345092f
C3591 vdd.n807 gnd 0.006754f
C3592 vdd.n808 gnd 0.006754f
C3593 vdd.n809 gnd 0.006754f
C3594 vdd.n810 gnd 0.006754f
C3595 vdd.n811 gnd 0.43644f
C3596 vdd.n812 gnd 0.006754f
C3597 vdd.n813 gnd 0.006754f
C3598 vdd.n814 gnd 0.006754f
C3599 vdd.n815 gnd 0.006754f
C3600 vdd.n816 gnd 0.006754f
C3601 vdd.n817 gnd 0.588686f
C3602 vdd.n818 gnd 0.006754f
C3603 vdd.n819 gnd 0.006754f
C3604 vdd.t85 gnd 0.309568f
C3605 vdd.t115 gnd 0.253744f
C3606 vdd.n820 gnd 0.006754f
C3607 vdd.n821 gnd 0.006754f
C3608 vdd.n822 gnd 0.006754f
C3609 vdd.t100 gnd 0.345092f
C3610 vdd.n823 gnd 0.006754f
C3611 vdd.n824 gnd 0.006754f
C3612 vdd.t98 gnd 0.345092f
C3613 vdd.n825 gnd 0.006754f
C3614 vdd.n826 gnd 0.006754f
C3615 vdd.n827 gnd 0.006754f
C3616 vdd.t101 gnd 0.268969f
C3617 vdd.n828 gnd 0.006754f
C3618 vdd.n829 gnd 0.006754f
C3619 vdd.n830 gnd 0.573462f
C3620 vdd.n831 gnd 0.006754f
C3621 vdd.n832 gnd 0.006754f
C3622 vdd.n833 gnd 0.006754f
C3623 vdd.t105 gnd 0.345092f
C3624 vdd.n834 gnd 0.006754f
C3625 vdd.n835 gnd 0.006754f
C3626 vdd.t117 gnd 0.294343f
C3627 vdd.n836 gnd 0.421215f
C3628 vdd.n837 gnd 0.006754f
C3629 vdd.n838 gnd 0.006754f
C3630 vdd.n839 gnd 0.006754f
C3631 vdd.n840 gnd 0.573462f
C3632 vdd.n841 gnd 0.006754f
C3633 vdd.n842 gnd 0.006754f
C3634 vdd.t81 gnd 0.345092f
C3635 vdd.n843 gnd 0.006754f
C3636 vdd.n844 gnd 0.006754f
C3637 vdd.n845 gnd 0.006754f
C3638 vdd.n846 gnd 0.690184f
C3639 vdd.n847 gnd 0.006754f
C3640 vdd.n848 gnd 0.006754f
C3641 vdd.t110 gnd 0.345092f
C3642 vdd.n849 gnd 0.006754f
C3643 vdd.n850 gnd 0.006754f
C3644 vdd.n851 gnd 0.006754f
C3645 vdd.t109 gnd 0.081198f
C3646 vdd.n852 gnd 0.006754f
C3647 vdd.n853 gnd 0.006754f
C3648 vdd.n854 gnd 0.006754f
C3649 vdd.t62 gnd 0.279359f
C3650 vdd.t60 gnd 0.178167f
C3651 vdd.t63 gnd 0.279359f
C3652 vdd.n855 gnd 0.157011f
C3653 vdd.n856 gnd 0.006754f
C3654 vdd.n857 gnd 0.006754f
C3655 vdd.n858 gnd 0.690184f
C3656 vdd.n859 gnd 0.006754f
C3657 vdd.n860 gnd 0.006754f
C3658 vdd.t61 gnd 0.309568f
C3659 vdd.n861 gnd 0.608986f
C3660 vdd.n862 gnd 0.006754f
C3661 vdd.n863 gnd 0.006754f
C3662 vdd.n864 gnd 0.006754f
C3663 vdd.n865 gnd 0.603911f
C3664 vdd.n866 gnd 0.006754f
C3665 vdd.n867 gnd 0.006754f
C3666 vdd.n868 gnd 0.006754f
C3667 vdd.n869 gnd 0.006754f
C3668 vdd.n870 gnd 0.006754f
C3669 vdd.n871 gnd 0.690184f
C3670 vdd.n872 gnd 0.006754f
C3671 vdd.n873 gnd 0.006754f
C3672 vdd.t8 gnd 0.345092f
C3673 vdd.n874 gnd 0.006754f
C3674 vdd.n875 gnd 0.016025f
C3675 vdd.n876 gnd 0.016025f
C3676 vdd.n877 gnd 6.99319f
C3677 vdd.n878 gnd 0.014962f
C3678 vdd.n879 gnd 0.014962f
C3679 vdd.n880 gnd 0.016025f
C3680 vdd.n881 gnd 0.006754f
C3681 vdd.n882 gnd 0.006754f
C3682 vdd.n883 gnd 0.006754f
C3683 vdd.n884 gnd 0.006754f
C3684 vdd.n885 gnd 0.006754f
C3685 vdd.n886 gnd 0.006754f
C3686 vdd.n887 gnd 0.006754f
C3687 vdd.n888 gnd 0.006754f
C3688 vdd.n890 gnd 0.006754f
C3689 vdd.n891 gnd 0.006754f
C3690 vdd.n892 gnd 0.006356f
C3691 vdd.n895 gnd 0.023771f
C3692 vdd.n896 gnd 0.007994f
C3693 vdd.n897 gnd 0.009932f
C3694 vdd.n899 gnd 0.009932f
C3695 vdd.n900 gnd 0.006635f
C3696 vdd.t23 gnd 0.507488f
C3697 vdd.n901 gnd 7.26723f
C3698 vdd.n902 gnd 0.009932f
C3699 vdd.n903 gnd 0.023771f
C3700 vdd.n904 gnd 0.007994f
C3701 vdd.n905 gnd 0.009932f
C3702 vdd.n906 gnd 0.007994f
C3703 vdd.n907 gnd 0.009932f
C3704 vdd.n908 gnd 1.01498f
C3705 vdd.n909 gnd 0.009932f
C3706 vdd.n910 gnd 0.007994f
C3707 vdd.n911 gnd 0.007994f
C3708 vdd.n912 gnd 0.009932f
C3709 vdd.n913 gnd 0.007994f
C3710 vdd.n914 gnd 0.009932f
C3711 vdd.t136 gnd 0.507488f
C3712 vdd.n915 gnd 0.009932f
C3713 vdd.n916 gnd 0.007994f
C3714 vdd.n917 gnd 0.009932f
C3715 vdd.n918 gnd 0.007994f
C3716 vdd.n919 gnd 0.009932f
C3717 vdd.t214 gnd 0.507488f
C3718 vdd.n920 gnd 0.009932f
C3719 vdd.n921 gnd 0.007994f
C3720 vdd.n922 gnd 0.009932f
C3721 vdd.n923 gnd 0.007994f
C3722 vdd.n924 gnd 0.009932f
C3723 vdd.t150 gnd 0.507488f
C3724 vdd.n925 gnd 0.796757f
C3725 vdd.n926 gnd 0.009932f
C3726 vdd.n927 gnd 0.007994f
C3727 vdd.n928 gnd 0.009932f
C3728 vdd.n929 gnd 0.007994f
C3729 vdd.n930 gnd 0.009932f
C3730 vdd.n931 gnd 0.715558f
C3731 vdd.n932 gnd 0.009932f
C3732 vdd.n933 gnd 0.007994f
C3733 vdd.n934 gnd 0.009932f
C3734 vdd.n935 gnd 0.007994f
C3735 vdd.n936 gnd 0.009932f
C3736 vdd.n937 gnd 0.543012f
C3737 vdd.t163 gnd 0.507488f
C3738 vdd.n938 gnd 0.009932f
C3739 vdd.n939 gnd 0.007994f
C3740 vdd.n940 gnd 0.009898f
C3741 vdd.n941 gnd 0.007994f
C3742 vdd.n942 gnd 0.009932f
C3743 vdd.t175 gnd 0.507488f
C3744 vdd.n943 gnd 0.009932f
C3745 vdd.n944 gnd 0.007994f
C3746 vdd.n945 gnd 0.009932f
C3747 vdd.n946 gnd 0.007994f
C3748 vdd.n947 gnd 0.009932f
C3749 vdd.t195 gnd 0.507488f
C3750 vdd.n948 gnd 0.64451f
C3751 vdd.n949 gnd 0.009932f
C3752 vdd.n950 gnd 0.007994f
C3753 vdd.n951 gnd 0.009932f
C3754 vdd.n952 gnd 0.007994f
C3755 vdd.n953 gnd 0.009932f
C3756 vdd.t188 gnd 0.507488f
C3757 vdd.n954 gnd 0.009932f
C3758 vdd.n955 gnd 0.007994f
C3759 vdd.n956 gnd 0.009932f
C3760 vdd.n957 gnd 0.007994f
C3761 vdd.n958 gnd 0.009932f
C3762 vdd.n959 gnd 0.695259f
C3763 vdd.n960 gnd 0.84243f
C3764 vdd.t144 gnd 0.507488f
C3765 vdd.n961 gnd 0.009932f
C3766 vdd.n962 gnd 0.007994f
C3767 vdd.n963 gnd 0.009932f
C3768 vdd.n964 gnd 0.007994f
C3769 vdd.n965 gnd 0.009932f
C3770 vdd.n966 gnd 0.522713f
C3771 vdd.n967 gnd 0.009932f
C3772 vdd.n968 gnd 0.007994f
C3773 vdd.n969 gnd 0.009932f
C3774 vdd.n970 gnd 0.007994f
C3775 vdd.n971 gnd 0.009932f
C3776 vdd.n972 gnd 1.01498f
C3777 vdd.t155 gnd 0.507488f
C3778 vdd.n973 gnd 0.009932f
C3779 vdd.n974 gnd 0.007994f
C3780 vdd.n975 gnd 0.009932f
C3781 vdd.n976 gnd 0.007994f
C3782 vdd.n977 gnd 0.009932f
C3783 vdd.t4 gnd 0.507488f
C3784 vdd.n978 gnd 0.009932f
C3785 vdd.n979 gnd 0.007994f
C3786 vdd.n980 gnd 0.023771f
C3787 vdd.n981 gnd 0.023771f
C3788 vdd.n982 gnd 2.33445f
C3789 vdd.n983 gnd 0.573462f
C3790 vdd.n984 gnd 0.023771f
C3791 vdd.n985 gnd 0.009932f
C3792 vdd.n987 gnd 0.009932f
C3793 vdd.n988 gnd 0.009932f
C3794 vdd.n989 gnd 0.007994f
C3795 vdd.n990 gnd 0.009932f
C3796 vdd.n991 gnd 0.009932f
C3797 vdd.n993 gnd 0.009932f
C3798 vdd.n994 gnd 0.009932f
C3799 vdd.n996 gnd 0.009932f
C3800 vdd.n997 gnd 0.007994f
C3801 vdd.n998 gnd 0.009932f
C3802 vdd.n999 gnd 0.009932f
C3803 vdd.n1001 gnd 0.009932f
C3804 vdd.n1002 gnd 0.009932f
C3805 vdd.n1004 gnd 0.009932f
C3806 vdd.n1005 gnd 0.007994f
C3807 vdd.n1006 gnd 0.009932f
C3808 vdd.n1007 gnd 0.009932f
C3809 vdd.n1009 gnd 0.009932f
C3810 vdd.n1010 gnd 0.009932f
C3811 vdd.n1012 gnd 0.009932f
C3812 vdd.n1013 gnd 0.007994f
C3813 vdd.n1014 gnd 0.009932f
C3814 vdd.n1015 gnd 0.009932f
C3815 vdd.n1017 gnd 0.009932f
C3816 vdd.n1018 gnd 0.009932f
C3817 vdd.n1020 gnd 0.009932f
C3818 vdd.t37 gnd 0.122186f
C3819 vdd.t38 gnd 0.130584f
C3820 vdd.t36 gnd 0.159574f
C3821 vdd.n1021 gnd 0.204551f
C3822 vdd.n1022 gnd 0.172659f
C3823 vdd.n1023 gnd 0.017107f
C3824 vdd.n1024 gnd 0.009932f
C3825 vdd.n1025 gnd 0.009932f
C3826 vdd.n1027 gnd 0.009932f
C3827 vdd.n1028 gnd 0.009932f
C3828 vdd.n1030 gnd 0.009932f
C3829 vdd.n1031 gnd 0.007994f
C3830 vdd.n1032 gnd 0.009932f
C3831 vdd.n1033 gnd 0.009932f
C3832 vdd.n1035 gnd 0.009932f
C3833 vdd.n1036 gnd 0.009932f
C3834 vdd.n1038 gnd 0.009932f
C3835 vdd.n1039 gnd 0.007994f
C3836 vdd.n1040 gnd 0.009932f
C3837 vdd.n1041 gnd 0.009932f
C3838 vdd.n1043 gnd 0.009932f
C3839 vdd.n1044 gnd 0.009932f
C3840 vdd.n1046 gnd 0.009932f
C3841 vdd.n1047 gnd 0.007994f
C3842 vdd.n1048 gnd 0.009932f
C3843 vdd.n1049 gnd 0.009932f
C3844 vdd.n1051 gnd 0.009932f
C3845 vdd.n1052 gnd 0.009932f
C3846 vdd.n1054 gnd 0.009932f
C3847 vdd.n1055 gnd 0.007994f
C3848 vdd.n1056 gnd 0.009932f
C3849 vdd.n1057 gnd 0.009932f
C3850 vdd.n1059 gnd 0.009932f
C3851 vdd.n1060 gnd 0.009932f
C3852 vdd.n1062 gnd 0.009932f
C3853 vdd.n1063 gnd 0.007994f
C3854 vdd.n1064 gnd 0.009932f
C3855 vdd.n1065 gnd 0.009932f
C3856 vdd.n1067 gnd 0.009932f
C3857 vdd.n1068 gnd 0.007914f
C3858 vdd.n1070 gnd 0.007994f
C3859 vdd.n1071 gnd 0.009932f
C3860 vdd.n1072 gnd 0.009932f
C3861 vdd.n1073 gnd 0.009932f
C3862 vdd.n1074 gnd 0.009932f
C3863 vdd.n1076 gnd 0.009932f
C3864 vdd.n1077 gnd 0.009932f
C3865 vdd.n1078 gnd 0.007994f
C3866 vdd.n1079 gnd 0.009932f
C3867 vdd.n1081 gnd 0.009932f
C3868 vdd.n1082 gnd 0.009932f
C3869 vdd.n1084 gnd 0.009932f
C3870 vdd.n1085 gnd 0.009932f
C3871 vdd.n1086 gnd 0.007994f
C3872 vdd.n1087 gnd 0.009932f
C3873 vdd.n1089 gnd 0.009932f
C3874 vdd.n1090 gnd 0.009932f
C3875 vdd.n1092 gnd 0.009932f
C3876 vdd.n1093 gnd 0.009932f
C3877 vdd.n1094 gnd 0.007994f
C3878 vdd.n1095 gnd 0.009932f
C3879 vdd.n1097 gnd 0.009932f
C3880 vdd.n1098 gnd 0.009932f
C3881 vdd.n1100 gnd 0.009932f
C3882 vdd.n1101 gnd 0.009932f
C3883 vdd.n1102 gnd 0.007994f
C3884 vdd.n1103 gnd 0.009932f
C3885 vdd.n1105 gnd 0.009932f
C3886 vdd.n1106 gnd 0.009932f
C3887 vdd.n1108 gnd 0.009932f
C3888 vdd.n1109 gnd 0.003797f
C3889 vdd.t5 gnd 0.122186f
C3890 vdd.t6 gnd 0.130584f
C3891 vdd.t3 gnd 0.159574f
C3892 vdd.n1110 gnd 0.204551f
C3893 vdd.n1111 gnd 0.172659f
C3894 vdd.n1112 gnd 0.01311f
C3895 vdd.n1113 gnd 0.004197f
C3896 vdd.n1114 gnd 0.007994f
C3897 vdd.n1115 gnd 0.009932f
C3898 vdd.n1116 gnd 0.009932f
C3899 vdd.n1117 gnd 0.009932f
C3900 vdd.n1118 gnd 0.007994f
C3901 vdd.n1119 gnd 0.007994f
C3902 vdd.n1120 gnd 0.007994f
C3903 vdd.n1121 gnd 0.009932f
C3904 vdd.n1122 gnd 0.009932f
C3905 vdd.n1123 gnd 0.009932f
C3906 vdd.n1124 gnd 0.007994f
C3907 vdd.n1125 gnd 0.007994f
C3908 vdd.n1126 gnd 0.007994f
C3909 vdd.n1127 gnd 0.009932f
C3910 vdd.n1128 gnd 0.009932f
C3911 vdd.n1129 gnd 0.009932f
C3912 vdd.n1130 gnd 0.007994f
C3913 vdd.n1131 gnd 0.007994f
C3914 vdd.n1132 gnd 0.007994f
C3915 vdd.n1133 gnd 0.009932f
C3916 vdd.n1134 gnd 0.009932f
C3917 vdd.n1135 gnd 0.009932f
C3918 vdd.n1136 gnd 0.007994f
C3919 vdd.n1137 gnd 0.007994f
C3920 vdd.n1138 gnd 0.007994f
C3921 vdd.n1139 gnd 0.009932f
C3922 vdd.n1140 gnd 0.009932f
C3923 vdd.n1141 gnd 0.009932f
C3924 vdd.n1142 gnd 0.007994f
C3925 vdd.n1143 gnd 0.009932f
C3926 vdd.n1144 gnd 0.009932f
C3927 vdd.n1146 gnd 0.009932f
C3928 vdd.t27 gnd 0.122186f
C3929 vdd.t28 gnd 0.130584f
C3930 vdd.t26 gnd 0.159574f
C3931 vdd.n1147 gnd 0.204551f
C3932 vdd.n1148 gnd 0.172659f
C3933 vdd.n1149 gnd 0.017107f
C3934 vdd.n1150 gnd 0.005436f
C3935 vdd.n1151 gnd 0.009932f
C3936 vdd.n1152 gnd 0.009932f
C3937 vdd.n1153 gnd 0.009932f
C3938 vdd.n1154 gnd 0.007994f
C3939 vdd.n1155 gnd 0.007994f
C3940 vdd.n1156 gnd 0.007994f
C3941 vdd.n1157 gnd 0.009932f
C3942 vdd.n1158 gnd 0.009932f
C3943 vdd.n1159 gnd 0.009932f
C3944 vdd.n1160 gnd 0.007994f
C3945 vdd.n1161 gnd 0.007994f
C3946 vdd.n1162 gnd 0.007994f
C3947 vdd.n1163 gnd 0.009932f
C3948 vdd.n1164 gnd 0.009932f
C3949 vdd.n1165 gnd 0.009932f
C3950 vdd.n1166 gnd 0.007994f
C3951 vdd.n1167 gnd 0.007994f
C3952 vdd.n1168 gnd 0.007994f
C3953 vdd.n1169 gnd 0.009932f
C3954 vdd.n1170 gnd 0.009932f
C3955 vdd.n1171 gnd 0.009932f
C3956 vdd.n1172 gnd 0.007994f
C3957 vdd.n1173 gnd 0.007994f
C3958 vdd.n1174 gnd 0.007994f
C3959 vdd.n1175 gnd 0.009932f
C3960 vdd.n1176 gnd 0.009932f
C3961 vdd.n1177 gnd 0.009932f
C3962 vdd.n1178 gnd 0.007994f
C3963 vdd.n1179 gnd 0.007994f
C3964 vdd.n1180 gnd 0.006675f
C3965 vdd.n1181 gnd 0.009932f
C3966 vdd.n1182 gnd 0.009932f
C3967 vdd.n1183 gnd 0.009932f
C3968 vdd.n1184 gnd 0.006675f
C3969 vdd.n1185 gnd 0.007994f
C3970 vdd.n1186 gnd 0.007994f
C3971 vdd.n1187 gnd 0.009932f
C3972 vdd.n1188 gnd 0.009932f
C3973 vdd.n1189 gnd 0.009932f
C3974 vdd.n1190 gnd 0.007994f
C3975 vdd.n1191 gnd 0.007994f
C3976 vdd.n1192 gnd 0.007994f
C3977 vdd.n1193 gnd 0.009932f
C3978 vdd.n1194 gnd 0.009932f
C3979 vdd.n1195 gnd 0.009932f
C3980 vdd.n1196 gnd 0.007994f
C3981 vdd.n1197 gnd 0.007994f
C3982 vdd.n1198 gnd 0.007994f
C3983 vdd.n1199 gnd 0.009932f
C3984 vdd.n1200 gnd 0.009932f
C3985 vdd.n1201 gnd 0.009932f
C3986 vdd.n1202 gnd 0.007994f
C3987 vdd.n1203 gnd 0.007994f
C3988 vdd.n1204 gnd 0.007994f
C3989 vdd.n1205 gnd 0.009932f
C3990 vdd.n1206 gnd 0.009932f
C3991 vdd.n1207 gnd 0.009932f
C3992 vdd.n1208 gnd 0.007994f
C3993 vdd.n1209 gnd 0.007994f
C3994 vdd.n1210 gnd 0.006635f
C3995 vdd.n1211 gnd 0.023771f
C3996 vdd.n1212 gnd 0.023405f
C3997 vdd.n1213 gnd 0.006635f
C3998 vdd.n1214 gnd 0.023405f
C3999 vdd.n1215 gnd 1.43112f
C4000 vdd.n1216 gnd 0.023405f
C4001 vdd.n1217 gnd 0.006635f
C4002 vdd.n1218 gnd 0.023405f
C4003 vdd.n1219 gnd 0.009932f
C4004 vdd.n1220 gnd 0.009932f
C4005 vdd.n1221 gnd 0.007994f
C4006 vdd.n1222 gnd 0.009932f
C4007 vdd.n1223 gnd 0.949003f
C4008 vdd.n1224 gnd 0.009932f
C4009 vdd.n1225 gnd 0.007994f
C4010 vdd.n1226 gnd 0.009932f
C4011 vdd.n1227 gnd 0.009932f
C4012 vdd.n1228 gnd 0.009932f
C4013 vdd.n1229 gnd 0.007994f
C4014 vdd.n1230 gnd 0.009932f
C4015 vdd.n1231 gnd 0.999752f
C4016 vdd.n1232 gnd 0.009932f
C4017 vdd.n1233 gnd 0.007994f
C4018 vdd.n1234 gnd 0.009932f
C4019 vdd.n1235 gnd 0.009932f
C4020 vdd.n1236 gnd 0.009932f
C4021 vdd.n1237 gnd 0.007994f
C4022 vdd.n1238 gnd 0.009932f
C4023 vdd.t169 gnd 0.507488f
C4024 vdd.n1239 gnd 0.827206f
C4025 vdd.n1240 gnd 0.009932f
C4026 vdd.n1241 gnd 0.007994f
C4027 vdd.n1242 gnd 0.009932f
C4028 vdd.n1243 gnd 0.009932f
C4029 vdd.n1244 gnd 0.009932f
C4030 vdd.n1245 gnd 0.007994f
C4031 vdd.n1246 gnd 0.009932f
C4032 vdd.n1247 gnd 0.65466f
C4033 vdd.n1248 gnd 0.009932f
C4034 vdd.n1249 gnd 0.007994f
C4035 vdd.n1250 gnd 0.009932f
C4036 vdd.n1251 gnd 0.009932f
C4037 vdd.n1252 gnd 0.009932f
C4038 vdd.n1253 gnd 0.007994f
C4039 vdd.n1254 gnd 0.009932f
C4040 vdd.n1255 gnd 0.817056f
C4041 vdd.n1256 gnd 0.532863f
C4042 vdd.n1257 gnd 0.009932f
C4043 vdd.n1258 gnd 0.007994f
C4044 vdd.n1259 gnd 0.009932f
C4045 vdd.n1260 gnd 0.009932f
C4046 vdd.n1261 gnd 0.009932f
C4047 vdd.n1262 gnd 0.007994f
C4048 vdd.n1263 gnd 0.009932f
C4049 vdd.n1264 gnd 0.705409f
C4050 vdd.n1265 gnd 0.009932f
C4051 vdd.n1266 gnd 0.007994f
C4052 vdd.n1267 gnd 0.009932f
C4053 vdd.n1268 gnd 0.009932f
C4054 vdd.n1269 gnd 0.009932f
C4055 vdd.n1270 gnd 0.007994f
C4056 vdd.n1271 gnd 0.009932f
C4057 vdd.t138 gnd 0.507488f
C4058 vdd.n1272 gnd 0.84243f
C4059 vdd.n1273 gnd 0.009932f
C4060 vdd.n1274 gnd 0.007994f
C4061 vdd.n1275 gnd 0.005451f
C4062 vdd.n1276 gnd 0.005058f
C4063 vdd.n1277 gnd 0.002798f
C4064 vdd.n1278 gnd 0.006424f
C4065 vdd.n1279 gnd 0.002718f
C4066 vdd.n1280 gnd 0.002878f
C4067 vdd.n1281 gnd 0.005058f
C4068 vdd.n1282 gnd 0.002718f
C4069 vdd.n1283 gnd 0.006424f
C4070 vdd.n1284 gnd 0.002878f
C4071 vdd.n1285 gnd 0.005058f
C4072 vdd.n1286 gnd 0.002718f
C4073 vdd.n1287 gnd 0.004818f
C4074 vdd.n1288 gnd 0.004833f
C4075 vdd.t137 gnd 0.013802f
C4076 vdd.n1289 gnd 0.030709f
C4077 vdd.n1290 gnd 0.159815f
C4078 vdd.n1291 gnd 0.002718f
C4079 vdd.n1292 gnd 0.002878f
C4080 vdd.n1293 gnd 0.006424f
C4081 vdd.n1294 gnd 0.006424f
C4082 vdd.n1295 gnd 0.002878f
C4083 vdd.n1296 gnd 0.002718f
C4084 vdd.n1297 gnd 0.005058f
C4085 vdd.n1298 gnd 0.005058f
C4086 vdd.n1299 gnd 0.002718f
C4087 vdd.n1300 gnd 0.002878f
C4088 vdd.n1301 gnd 0.006424f
C4089 vdd.n1302 gnd 0.006424f
C4090 vdd.n1303 gnd 0.002878f
C4091 vdd.n1304 gnd 0.002718f
C4092 vdd.n1305 gnd 0.005058f
C4093 vdd.n1306 gnd 0.005058f
C4094 vdd.n1307 gnd 0.002718f
C4095 vdd.n1308 gnd 0.002878f
C4096 vdd.n1309 gnd 0.006424f
C4097 vdd.n1310 gnd 0.006424f
C4098 vdd.n1311 gnd 0.015188f
C4099 vdd.n1312 gnd 0.002798f
C4100 vdd.n1313 gnd 0.002718f
C4101 vdd.n1314 gnd 0.013073f
C4102 vdd.n1315 gnd 0.009127f
C4103 vdd.t185 gnd 0.031975f
C4104 vdd.t217 gnd 0.031975f
C4105 vdd.n1316 gnd 0.219757f
C4106 vdd.n1317 gnd 0.172805f
C4107 vdd.t164 gnd 0.031975f
C4108 vdd.t205 gnd 0.031975f
C4109 vdd.n1318 gnd 0.219757f
C4110 vdd.n1319 gnd 0.139453f
C4111 vdd.t176 gnd 0.031975f
C4112 vdd.t211 gnd 0.031975f
C4113 vdd.n1320 gnd 0.219757f
C4114 vdd.n1321 gnd 0.139453f
C4115 vdd.t189 gnd 0.031975f
C4116 vdd.t221 gnd 0.031975f
C4117 vdd.n1322 gnd 0.219757f
C4118 vdd.n1323 gnd 0.139453f
C4119 vdd.t170 gnd 0.031975f
C4120 vdd.t152 gnd 0.031975f
C4121 vdd.n1324 gnd 0.219757f
C4122 vdd.n1325 gnd 0.139453f
C4123 vdd.n1326 gnd 0.005451f
C4124 vdd.n1327 gnd 0.005058f
C4125 vdd.n1328 gnd 0.002798f
C4126 vdd.n1329 gnd 0.006424f
C4127 vdd.n1330 gnd 0.002718f
C4128 vdd.n1331 gnd 0.002878f
C4129 vdd.n1332 gnd 0.005058f
C4130 vdd.n1333 gnd 0.002718f
C4131 vdd.n1334 gnd 0.006424f
C4132 vdd.n1335 gnd 0.002878f
C4133 vdd.n1336 gnd 0.005058f
C4134 vdd.n1337 gnd 0.002718f
C4135 vdd.n1338 gnd 0.004818f
C4136 vdd.n1339 gnd 0.004833f
C4137 vdd.t156 gnd 0.013802f
C4138 vdd.n1340 gnd 0.030709f
C4139 vdd.n1341 gnd 0.159815f
C4140 vdd.n1342 gnd 0.002718f
C4141 vdd.n1343 gnd 0.002878f
C4142 vdd.n1344 gnd 0.006424f
C4143 vdd.n1345 gnd 0.006424f
C4144 vdd.n1346 gnd 0.002878f
C4145 vdd.n1347 gnd 0.002718f
C4146 vdd.n1348 gnd 0.005058f
C4147 vdd.n1349 gnd 0.005058f
C4148 vdd.n1350 gnd 0.002718f
C4149 vdd.n1351 gnd 0.002878f
C4150 vdd.n1352 gnd 0.006424f
C4151 vdd.n1353 gnd 0.006424f
C4152 vdd.n1354 gnd 0.002878f
C4153 vdd.n1355 gnd 0.002718f
C4154 vdd.n1356 gnd 0.005058f
C4155 vdd.n1357 gnd 0.005058f
C4156 vdd.n1358 gnd 0.002718f
C4157 vdd.n1359 gnd 0.002878f
C4158 vdd.n1360 gnd 0.006424f
C4159 vdd.n1361 gnd 0.006424f
C4160 vdd.n1362 gnd 0.015188f
C4161 vdd.n1363 gnd 0.002798f
C4162 vdd.n1364 gnd 0.002718f
C4163 vdd.n1365 gnd 0.013073f
C4164 vdd.n1366 gnd 0.008841f
C4165 vdd.n1367 gnd 0.103754f
C4166 vdd.n1368 gnd 0.005451f
C4167 vdd.n1369 gnd 0.005058f
C4168 vdd.n1370 gnd 0.002798f
C4169 vdd.n1371 gnd 0.006424f
C4170 vdd.n1372 gnd 0.002718f
C4171 vdd.n1373 gnd 0.002878f
C4172 vdd.n1374 gnd 0.005058f
C4173 vdd.n1375 gnd 0.002718f
C4174 vdd.n1376 gnd 0.006424f
C4175 vdd.n1377 gnd 0.002878f
C4176 vdd.n1378 gnd 0.005058f
C4177 vdd.n1379 gnd 0.002718f
C4178 vdd.n1380 gnd 0.004818f
C4179 vdd.n1381 gnd 0.004833f
C4180 vdd.t212 gnd 0.013802f
C4181 vdd.n1382 gnd 0.030709f
C4182 vdd.n1383 gnd 0.159815f
C4183 vdd.n1384 gnd 0.002718f
C4184 vdd.n1385 gnd 0.002878f
C4185 vdd.n1386 gnd 0.006424f
C4186 vdd.n1387 gnd 0.006424f
C4187 vdd.n1388 gnd 0.002878f
C4188 vdd.n1389 gnd 0.002718f
C4189 vdd.n1390 gnd 0.005058f
C4190 vdd.n1391 gnd 0.005058f
C4191 vdd.n1392 gnd 0.002718f
C4192 vdd.n1393 gnd 0.002878f
C4193 vdd.n1394 gnd 0.006424f
C4194 vdd.n1395 gnd 0.006424f
C4195 vdd.n1396 gnd 0.002878f
C4196 vdd.n1397 gnd 0.002718f
C4197 vdd.n1398 gnd 0.005058f
C4198 vdd.n1399 gnd 0.005058f
C4199 vdd.n1400 gnd 0.002718f
C4200 vdd.n1401 gnd 0.002878f
C4201 vdd.n1402 gnd 0.006424f
C4202 vdd.n1403 gnd 0.006424f
C4203 vdd.n1404 gnd 0.015188f
C4204 vdd.n1405 gnd 0.002798f
C4205 vdd.n1406 gnd 0.002718f
C4206 vdd.n1407 gnd 0.013073f
C4207 vdd.n1408 gnd 0.009127f
C4208 vdd.t151 gnd 0.031975f
C4209 vdd.t215 gnd 0.031975f
C4210 vdd.n1409 gnd 0.219757f
C4211 vdd.n1410 gnd 0.172805f
C4212 vdd.t210 gnd 0.031975f
C4213 vdd.t198 gnd 0.031975f
C4214 vdd.n1411 gnd 0.219757f
C4215 vdd.n1412 gnd 0.139453f
C4216 vdd.t178 gnd 0.031975f
C4217 vdd.t139 gnd 0.031975f
C4218 vdd.n1413 gnd 0.219757f
C4219 vdd.n1414 gnd 0.139453f
C4220 vdd.t223 gnd 0.031975f
C4221 vdd.t196 gnd 0.031975f
C4222 vdd.n1415 gnd 0.219757f
C4223 vdd.n1416 gnd 0.139453f
C4224 vdd.t193 gnd 0.031975f
C4225 vdd.t145 gnd 0.031975f
C4226 vdd.n1417 gnd 0.219757f
C4227 vdd.n1418 gnd 0.139453f
C4228 vdd.n1419 gnd 0.005451f
C4229 vdd.n1420 gnd 0.005058f
C4230 vdd.n1421 gnd 0.002798f
C4231 vdd.n1422 gnd 0.006424f
C4232 vdd.n1423 gnd 0.002718f
C4233 vdd.n1424 gnd 0.002878f
C4234 vdd.n1425 gnd 0.005058f
C4235 vdd.n1426 gnd 0.002718f
C4236 vdd.n1427 gnd 0.006424f
C4237 vdd.n1428 gnd 0.002878f
C4238 vdd.n1429 gnd 0.005058f
C4239 vdd.n1430 gnd 0.002718f
C4240 vdd.n1431 gnd 0.004818f
C4241 vdd.n1432 gnd 0.004833f
C4242 vdd.t194 gnd 0.013802f
C4243 vdd.n1433 gnd 0.030709f
C4244 vdd.n1434 gnd 0.159815f
C4245 vdd.n1435 gnd 0.002718f
C4246 vdd.n1436 gnd 0.002878f
C4247 vdd.n1437 gnd 0.006424f
C4248 vdd.n1438 gnd 0.006424f
C4249 vdd.n1439 gnd 0.002878f
C4250 vdd.n1440 gnd 0.002718f
C4251 vdd.n1441 gnd 0.005058f
C4252 vdd.n1442 gnd 0.005058f
C4253 vdd.n1443 gnd 0.002718f
C4254 vdd.n1444 gnd 0.002878f
C4255 vdd.n1445 gnd 0.006424f
C4256 vdd.n1446 gnd 0.006424f
C4257 vdd.n1447 gnd 0.002878f
C4258 vdd.n1448 gnd 0.002718f
C4259 vdd.n1449 gnd 0.005058f
C4260 vdd.n1450 gnd 0.005058f
C4261 vdd.n1451 gnd 0.002718f
C4262 vdd.n1452 gnd 0.002878f
C4263 vdd.n1453 gnd 0.006424f
C4264 vdd.n1454 gnd 0.006424f
C4265 vdd.n1455 gnd 0.015188f
C4266 vdd.n1456 gnd 0.002798f
C4267 vdd.n1457 gnd 0.002718f
C4268 vdd.n1458 gnd 0.013073f
C4269 vdd.n1459 gnd 0.008841f
C4270 vdd.n1460 gnd 0.061723f
C4271 vdd.n1461 gnd 0.222404f
C4272 vdd.n1462 gnd 0.005451f
C4273 vdd.n1463 gnd 0.005058f
C4274 vdd.n1464 gnd 0.002798f
C4275 vdd.n1465 gnd 0.006424f
C4276 vdd.n1466 gnd 0.002718f
C4277 vdd.n1467 gnd 0.002878f
C4278 vdd.n1468 gnd 0.005058f
C4279 vdd.n1469 gnd 0.002718f
C4280 vdd.n1470 gnd 0.006424f
C4281 vdd.n1471 gnd 0.002878f
C4282 vdd.n1472 gnd 0.005058f
C4283 vdd.n1473 gnd 0.002718f
C4284 vdd.n1474 gnd 0.004818f
C4285 vdd.n1475 gnd 0.004833f
C4286 vdd.t224 gnd 0.013802f
C4287 vdd.n1476 gnd 0.030709f
C4288 vdd.n1477 gnd 0.159815f
C4289 vdd.n1478 gnd 0.002718f
C4290 vdd.n1479 gnd 0.002878f
C4291 vdd.n1480 gnd 0.006424f
C4292 vdd.n1481 gnd 0.006424f
C4293 vdd.n1482 gnd 0.002878f
C4294 vdd.n1483 gnd 0.002718f
C4295 vdd.n1484 gnd 0.005058f
C4296 vdd.n1485 gnd 0.005058f
C4297 vdd.n1486 gnd 0.002718f
C4298 vdd.n1487 gnd 0.002878f
C4299 vdd.n1488 gnd 0.006424f
C4300 vdd.n1489 gnd 0.006424f
C4301 vdd.n1490 gnd 0.002878f
C4302 vdd.n1491 gnd 0.002718f
C4303 vdd.n1492 gnd 0.005058f
C4304 vdd.n1493 gnd 0.005058f
C4305 vdd.n1494 gnd 0.002718f
C4306 vdd.n1495 gnd 0.002878f
C4307 vdd.n1496 gnd 0.006424f
C4308 vdd.n1497 gnd 0.006424f
C4309 vdd.n1498 gnd 0.015188f
C4310 vdd.n1499 gnd 0.002798f
C4311 vdd.n1500 gnd 0.002718f
C4312 vdd.n1501 gnd 0.013073f
C4313 vdd.n1502 gnd 0.009127f
C4314 vdd.t160 gnd 0.031975f
C4315 vdd.t225 gnd 0.031975f
C4316 vdd.n1503 gnd 0.219757f
C4317 vdd.n1504 gnd 0.172805f
C4318 vdd.t219 gnd 0.031975f
C4319 vdd.t208 gnd 0.031975f
C4320 vdd.n1505 gnd 0.219757f
C4321 vdd.n1506 gnd 0.139453f
C4322 vdd.t187 gnd 0.031975f
C4323 vdd.t158 gnd 0.031975f
C4324 vdd.n1507 gnd 0.219757f
C4325 vdd.n1508 gnd 0.139453f
C4326 vdd.t227 gnd 0.031975f
C4327 vdd.t206 gnd 0.031975f
C4328 vdd.n1509 gnd 0.219757f
C4329 vdd.n1510 gnd 0.139453f
C4330 vdd.t202 gnd 0.031975f
C4331 vdd.t171 gnd 0.031975f
C4332 vdd.n1511 gnd 0.219757f
C4333 vdd.n1512 gnd 0.139453f
C4334 vdd.n1513 gnd 0.005451f
C4335 vdd.n1514 gnd 0.005058f
C4336 vdd.n1515 gnd 0.002798f
C4337 vdd.n1516 gnd 0.006424f
C4338 vdd.n1517 gnd 0.002718f
C4339 vdd.n1518 gnd 0.002878f
C4340 vdd.n1519 gnd 0.005058f
C4341 vdd.n1520 gnd 0.002718f
C4342 vdd.n1521 gnd 0.006424f
C4343 vdd.n1522 gnd 0.002878f
C4344 vdd.n1523 gnd 0.005058f
C4345 vdd.n1524 gnd 0.002718f
C4346 vdd.n1525 gnd 0.004818f
C4347 vdd.n1526 gnd 0.004833f
C4348 vdd.t203 gnd 0.013802f
C4349 vdd.n1527 gnd 0.030709f
C4350 vdd.n1528 gnd 0.159815f
C4351 vdd.n1529 gnd 0.002718f
C4352 vdd.n1530 gnd 0.002878f
C4353 vdd.n1531 gnd 0.006424f
C4354 vdd.n1532 gnd 0.006424f
C4355 vdd.n1533 gnd 0.002878f
C4356 vdd.n1534 gnd 0.002718f
C4357 vdd.n1535 gnd 0.005058f
C4358 vdd.n1536 gnd 0.005058f
C4359 vdd.n1537 gnd 0.002718f
C4360 vdd.n1538 gnd 0.002878f
C4361 vdd.n1539 gnd 0.006424f
C4362 vdd.n1540 gnd 0.006424f
C4363 vdd.n1541 gnd 0.002878f
C4364 vdd.n1542 gnd 0.002718f
C4365 vdd.n1543 gnd 0.005058f
C4366 vdd.n1544 gnd 0.005058f
C4367 vdd.n1545 gnd 0.002718f
C4368 vdd.n1546 gnd 0.002878f
C4369 vdd.n1547 gnd 0.006424f
C4370 vdd.n1548 gnd 0.006424f
C4371 vdd.n1549 gnd 0.015188f
C4372 vdd.n1550 gnd 0.002798f
C4373 vdd.n1551 gnd 0.002718f
C4374 vdd.n1552 gnd 0.013073f
C4375 vdd.n1553 gnd 0.008841f
C4376 vdd.n1554 gnd 0.061723f
C4377 vdd.n1555 gnd 0.244429f
C4378 vdd.n1556 gnd 2.19991f
C4379 vdd.n1557 gnd 0.591214f
C4380 vdd.n1558 gnd 0.009898f
C4381 vdd.n1559 gnd 0.009932f
C4382 vdd.n1560 gnd 0.007994f
C4383 vdd.n1561 gnd 0.009932f
C4384 vdd.n1562 gnd 0.806906f
C4385 vdd.n1563 gnd 0.009932f
C4386 vdd.n1564 gnd 0.007994f
C4387 vdd.n1565 gnd 0.009932f
C4388 vdd.n1566 gnd 0.009932f
C4389 vdd.n1567 gnd 0.009932f
C4390 vdd.n1568 gnd 0.007994f
C4391 vdd.n1569 gnd 0.009932f
C4392 vdd.n1570 gnd 0.84243f
C4393 vdd.t197 gnd 0.507488f
C4394 vdd.n1571 gnd 0.63436f
C4395 vdd.n1572 gnd 0.009932f
C4396 vdd.n1573 gnd 0.007994f
C4397 vdd.n1574 gnd 0.009932f
C4398 vdd.n1575 gnd 0.009932f
C4399 vdd.n1576 gnd 0.009932f
C4400 vdd.n1577 gnd 0.007994f
C4401 vdd.n1578 gnd 0.009932f
C4402 vdd.n1579 gnd 0.553162f
C4403 vdd.n1580 gnd 0.009932f
C4404 vdd.n1581 gnd 0.007994f
C4405 vdd.n1582 gnd 0.009932f
C4406 vdd.n1583 gnd 0.009932f
C4407 vdd.n1584 gnd 0.009932f
C4408 vdd.n1585 gnd 0.007994f
C4409 vdd.n1586 gnd 0.009932f
C4410 vdd.n1587 gnd 0.624211f
C4411 vdd.n1588 gnd 0.725708f
C4412 vdd.n1589 gnd 0.009932f
C4413 vdd.n1590 gnd 0.007994f
C4414 vdd.n1591 gnd 0.009932f
C4415 vdd.n1592 gnd 0.009932f
C4416 vdd.n1593 gnd 0.009932f
C4417 vdd.n1594 gnd 0.007994f
C4418 vdd.n1595 gnd 0.009932f
C4419 vdd.n1596 gnd 0.898254f
C4420 vdd.n1597 gnd 0.009932f
C4421 vdd.n1598 gnd 0.007994f
C4422 vdd.n1599 gnd 0.009932f
C4423 vdd.n1600 gnd 0.009932f
C4424 vdd.n1601 gnd 0.023405f
C4425 vdd.n1602 gnd 0.009932f
C4426 vdd.n1603 gnd 0.009932f
C4427 vdd.n1604 gnd 0.007994f
C4428 vdd.n1605 gnd 0.009932f
C4429 vdd.n1606 gnd 0.543012f
C4430 vdd.n1607 gnd 1.01498f
C4431 vdd.n1608 gnd 0.009932f
C4432 vdd.n1609 gnd 0.007994f
C4433 vdd.n1610 gnd 0.009932f
C4434 vdd.n1611 gnd 0.009932f
C4435 vdd.n1612 gnd 0.008541f
C4436 vdd.n1613 gnd 0.007994f
C4437 vdd.n1615 gnd 0.009932f
C4438 vdd.n1617 gnd 0.007994f
C4439 vdd.n1618 gnd 0.009932f
C4440 vdd.n1619 gnd 0.007994f
C4441 vdd.n1621 gnd 0.009932f
C4442 vdd.n1622 gnd 0.007994f
C4443 vdd.n1623 gnd 0.009932f
C4444 vdd.n1624 gnd 0.009932f
C4445 vdd.n1625 gnd 0.009932f
C4446 vdd.n1626 gnd 0.009932f
C4447 vdd.n1627 gnd 0.009932f
C4448 vdd.n1628 gnd 0.007994f
C4449 vdd.n1630 gnd 0.009932f
C4450 vdd.n1631 gnd 0.009932f
C4451 vdd.n1632 gnd 0.009932f
C4452 vdd.n1633 gnd 0.009932f
C4453 vdd.n1634 gnd 0.009932f
C4454 vdd.n1635 gnd 0.007994f
C4455 vdd.n1637 gnd 0.009932f
C4456 vdd.n1638 gnd 0.009932f
C4457 vdd.n1639 gnd 0.009932f
C4458 vdd.n1640 gnd 0.009932f
C4459 vdd.n1641 gnd 0.006675f
C4460 vdd.t41 gnd 0.122186f
C4461 vdd.t40 gnd 0.130584f
C4462 vdd.t39 gnd 0.159574f
C4463 vdd.n1642 gnd 0.204551f
C4464 vdd.n1643 gnd 0.17186f
C4465 vdd.n1645 gnd 0.009932f
C4466 vdd.n1646 gnd 0.009932f
C4467 vdd.n1647 gnd 0.007994f
C4468 vdd.n1648 gnd 0.009932f
C4469 vdd.n1650 gnd 0.009932f
C4470 vdd.n1651 gnd 0.009932f
C4471 vdd.n1652 gnd 0.009932f
C4472 vdd.n1653 gnd 0.009932f
C4473 vdd.n1654 gnd 0.007994f
C4474 vdd.n1656 gnd 0.009932f
C4475 vdd.n1657 gnd 0.009932f
C4476 vdd.n1658 gnd 0.009932f
C4477 vdd.n1659 gnd 0.009932f
C4478 vdd.n1660 gnd 0.009932f
C4479 vdd.n1661 gnd 0.007994f
C4480 vdd.n1663 gnd 0.009932f
C4481 vdd.n1664 gnd 0.009932f
C4482 vdd.n1665 gnd 0.009932f
C4483 vdd.n1666 gnd 0.009932f
C4484 vdd.n1667 gnd 0.009932f
C4485 vdd.n1668 gnd 0.007994f
C4486 vdd.n1670 gnd 0.009932f
C4487 vdd.n1671 gnd 0.009932f
C4488 vdd.n1672 gnd 0.009932f
C4489 vdd.n1673 gnd 0.009932f
C4490 vdd.n1674 gnd 0.009932f
C4491 vdd.n1675 gnd 0.007994f
C4492 vdd.n1677 gnd 0.009932f
C4493 vdd.n1678 gnd 0.009932f
C4494 vdd.n1679 gnd 0.009932f
C4495 vdd.n1680 gnd 0.009932f
C4496 vdd.n1681 gnd 0.007914f
C4497 vdd.t35 gnd 0.122186f
C4498 vdd.t34 gnd 0.130584f
C4499 vdd.t33 gnd 0.159574f
C4500 vdd.n1682 gnd 0.204551f
C4501 vdd.n1683 gnd 0.17186f
C4502 vdd.n1685 gnd 0.009932f
C4503 vdd.n1686 gnd 0.009932f
C4504 vdd.n1687 gnd 0.007994f
C4505 vdd.n1688 gnd 0.009932f
C4506 vdd.n1690 gnd 0.009932f
C4507 vdd.n1691 gnd 0.009932f
C4508 vdd.n1692 gnd 0.009932f
C4509 vdd.n1693 gnd 0.009932f
C4510 vdd.n1694 gnd 0.007994f
C4511 vdd.n1696 gnd 0.009932f
C4512 vdd.n1697 gnd 0.009932f
C4513 vdd.n1698 gnd 0.009932f
C4514 vdd.n1699 gnd 0.009932f
C4515 vdd.n1700 gnd 0.009932f
C4516 vdd.n1701 gnd 0.007994f
C4517 vdd.n1703 gnd 0.009932f
C4518 vdd.n1704 gnd 0.009932f
C4519 vdd.n1705 gnd 0.009932f
C4520 vdd.n1706 gnd 0.009932f
C4521 vdd.n1707 gnd 0.009932f
C4522 vdd.n1708 gnd 0.009932f
C4523 vdd.n1709 gnd 0.007994f
C4524 vdd.n1711 gnd 0.009932f
C4525 vdd.n1713 gnd 0.009932f
C4526 vdd.n1714 gnd 0.007994f
C4527 vdd.n1715 gnd 0.007994f
C4528 vdd.n1716 gnd 0.009932f
C4529 vdd.n1718 gnd 0.009932f
C4530 vdd.n1719 gnd 0.007994f
C4531 vdd.n1720 gnd 0.007994f
C4532 vdd.n1721 gnd 0.009932f
C4533 vdd.n1723 gnd 0.009932f
C4534 vdd.n1724 gnd 0.009932f
C4535 vdd.n1725 gnd 0.007994f
C4536 vdd.n1726 gnd 0.007994f
C4537 vdd.n1727 gnd 0.007994f
C4538 vdd.n1728 gnd 0.009932f
C4539 vdd.n1730 gnd 0.009932f
C4540 vdd.n1731 gnd 0.009932f
C4541 vdd.n1732 gnd 0.007994f
C4542 vdd.n1733 gnd 0.007994f
C4543 vdd.n1734 gnd 0.007994f
C4544 vdd.n1735 gnd 0.009932f
C4545 vdd.n1737 gnd 0.009932f
C4546 vdd.n1738 gnd 0.009932f
C4547 vdd.n1739 gnd 0.007994f
C4548 vdd.n1740 gnd 0.007994f
C4549 vdd.n1741 gnd 0.007994f
C4550 vdd.n1742 gnd 0.009932f
C4551 vdd.n1744 gnd 0.009932f
C4552 vdd.n1745 gnd 0.009932f
C4553 vdd.n1746 gnd 0.007994f
C4554 vdd.n1747 gnd 0.009932f
C4555 vdd.n1748 gnd 0.009932f
C4556 vdd.n1749 gnd 0.009932f
C4557 vdd.n1750 gnd 0.016307f
C4558 vdd.n1751 gnd 0.005436f
C4559 vdd.n1752 gnd 0.007994f
C4560 vdd.n1753 gnd 0.009932f
C4561 vdd.n1755 gnd 0.009932f
C4562 vdd.n1756 gnd 0.009932f
C4563 vdd.n1757 gnd 0.007994f
C4564 vdd.n1758 gnd 0.007994f
C4565 vdd.n1759 gnd 0.007994f
C4566 vdd.n1760 gnd 0.009932f
C4567 vdd.n1762 gnd 0.009932f
C4568 vdd.n1763 gnd 0.009932f
C4569 vdd.n1764 gnd 0.007994f
C4570 vdd.n1765 gnd 0.007994f
C4571 vdd.n1766 gnd 0.007994f
C4572 vdd.n1767 gnd 0.009932f
C4573 vdd.n1769 gnd 0.009932f
C4574 vdd.n1770 gnd 0.009932f
C4575 vdd.n1771 gnd 0.007994f
C4576 vdd.n1772 gnd 0.007994f
C4577 vdd.n1773 gnd 0.007994f
C4578 vdd.n1774 gnd 0.009932f
C4579 vdd.n1776 gnd 0.009932f
C4580 vdd.n1777 gnd 0.009932f
C4581 vdd.n1778 gnd 0.007994f
C4582 vdd.n1779 gnd 0.007994f
C4583 vdd.n1780 gnd 0.007994f
C4584 vdd.n1781 gnd 0.009932f
C4585 vdd.n1783 gnd 0.009932f
C4586 vdd.n1784 gnd 0.009932f
C4587 vdd.n1785 gnd 0.007994f
C4588 vdd.n1786 gnd 0.009932f
C4589 vdd.n1787 gnd 0.009932f
C4590 vdd.n1788 gnd 0.009932f
C4591 vdd.n1789 gnd 0.016307f
C4592 vdd.n1790 gnd 0.006675f
C4593 vdd.n1791 gnd 0.007994f
C4594 vdd.n1792 gnd 0.009932f
C4595 vdd.n1794 gnd 0.009932f
C4596 vdd.n1795 gnd 0.009932f
C4597 vdd.n1796 gnd 0.007994f
C4598 vdd.n1797 gnd 0.007994f
C4599 vdd.n1798 gnd 0.007994f
C4600 vdd.n1799 gnd 0.009932f
C4601 vdd.n1801 gnd 0.009932f
C4602 vdd.n1802 gnd 0.009932f
C4603 vdd.n1803 gnd 0.007994f
C4604 vdd.n1804 gnd 0.007994f
C4605 vdd.n1805 gnd 0.007994f
C4606 vdd.n1806 gnd 0.009932f
C4607 vdd.n1808 gnd 0.009932f
C4608 vdd.n1809 gnd 0.009932f
C4609 vdd.n1811 gnd 0.009932f
C4610 vdd.n1812 gnd 0.007994f
C4611 vdd.n1813 gnd 0.006356f
C4612 vdd.n1814 gnd 0.006754f
C4613 vdd.n1815 gnd 0.006754f
C4614 vdd.n1816 gnd 0.006754f
C4615 vdd.n1817 gnd 0.006754f
C4616 vdd.n1818 gnd 0.006754f
C4617 vdd.n1819 gnd 0.006754f
C4618 vdd.n1820 gnd 0.006754f
C4619 vdd.n1821 gnd 0.006754f
C4620 vdd.n1823 gnd 0.006754f
C4621 vdd.n1824 gnd 0.006754f
C4622 vdd.n1825 gnd 0.006754f
C4623 vdd.n1826 gnd 0.006754f
C4624 vdd.n1827 gnd 0.006754f
C4625 vdd.n1829 gnd 0.006754f
C4626 vdd.n1831 gnd 0.006754f
C4627 vdd.n1832 gnd 0.006754f
C4628 vdd.n1833 gnd 0.006754f
C4629 vdd.n1834 gnd 0.006754f
C4630 vdd.n1835 gnd 0.006754f
C4631 vdd.n1837 gnd 0.006754f
C4632 vdd.n1839 gnd 0.006754f
C4633 vdd.n1840 gnd 0.006754f
C4634 vdd.n1841 gnd 0.006754f
C4635 vdd.n1842 gnd 0.006754f
C4636 vdd.n1843 gnd 0.006754f
C4637 vdd.n1845 gnd 0.006754f
C4638 vdd.n1847 gnd 0.006754f
C4639 vdd.n1848 gnd 0.006754f
C4640 vdd.n1849 gnd 0.006754f
C4641 vdd.n1850 gnd 0.006754f
C4642 vdd.n1851 gnd 0.006754f
C4643 vdd.n1853 gnd 0.006754f
C4644 vdd.n1854 gnd 0.006754f
C4645 vdd.n1855 gnd 0.006754f
C4646 vdd.n1856 gnd 0.006754f
C4647 vdd.n1857 gnd 0.006754f
C4648 vdd.n1858 gnd 0.006754f
C4649 vdd.n1859 gnd 0.006754f
C4650 vdd.n1860 gnd 0.006754f
C4651 vdd.n1861 gnd 0.004916f
C4652 vdd.n1862 gnd 0.006754f
C4653 vdd.t9 gnd 0.272911f
C4654 vdd.t10 gnd 0.279359f
C4655 vdd.t7 gnd 0.178167f
C4656 vdd.n1863 gnd 0.096289f
C4657 vdd.n1864 gnd 0.054619f
C4658 vdd.n1865 gnd 0.009652f
C4659 vdd.n1866 gnd 0.006754f
C4660 vdd.n1867 gnd 0.006754f
C4661 vdd.n1868 gnd 0.411065f
C4662 vdd.n1869 gnd 0.006754f
C4663 vdd.n1870 gnd 0.006754f
C4664 vdd.n1871 gnd 0.006754f
C4665 vdd.n1872 gnd 0.006754f
C4666 vdd.n1873 gnd 0.006754f
C4667 vdd.n1874 gnd 0.006754f
C4668 vdd.n1875 gnd 0.006754f
C4669 vdd.n1876 gnd 0.006754f
C4670 vdd.n1877 gnd 0.006754f
C4671 vdd.n1878 gnd 0.006754f
C4672 vdd.n1879 gnd 0.006754f
C4673 vdd.n1880 gnd 0.006754f
C4674 vdd.n1881 gnd 0.006754f
C4675 vdd.n1882 gnd 0.006754f
C4676 vdd.n1883 gnd 0.006754f
C4677 vdd.n1884 gnd 0.006754f
C4678 vdd.n1885 gnd 0.006754f
C4679 vdd.n1886 gnd 0.006754f
C4680 vdd.n1887 gnd 0.006754f
C4681 vdd.n1888 gnd 0.006754f
C4682 vdd.t58 gnd 0.272911f
C4683 vdd.t59 gnd 0.279359f
C4684 vdd.t57 gnd 0.178167f
C4685 vdd.n1889 gnd 0.096289f
C4686 vdd.n1890 gnd 0.054619f
C4687 vdd.n1891 gnd 0.006754f
C4688 vdd.n1892 gnd 0.006754f
C4689 vdd.n1893 gnd 0.006754f
C4690 vdd.n1894 gnd 0.006754f
C4691 vdd.n1895 gnd 0.006754f
C4692 vdd.n1896 gnd 0.006754f
C4693 vdd.n1898 gnd 0.006754f
C4694 vdd.n1899 gnd 0.006754f
C4695 vdd.n1900 gnd 0.006754f
C4696 vdd.n1901 gnd 0.006754f
C4697 vdd.n1903 gnd 0.006754f
C4698 vdd.n1905 gnd 0.006754f
C4699 vdd.n1906 gnd 0.006754f
C4700 vdd.n1907 gnd 0.006754f
C4701 vdd.n1908 gnd 0.006754f
C4702 vdd.n1909 gnd 0.006754f
C4703 vdd.n1911 gnd 0.006754f
C4704 vdd.n1913 gnd 0.006754f
C4705 vdd.n1914 gnd 0.006754f
C4706 vdd.n1915 gnd 0.006754f
C4707 vdd.n1916 gnd 0.006754f
C4708 vdd.n1917 gnd 0.006754f
C4709 vdd.n1919 gnd 0.006754f
C4710 vdd.n1921 gnd 0.006754f
C4711 vdd.n1922 gnd 0.006754f
C4712 vdd.n1923 gnd 0.004916f
C4713 vdd.n1924 gnd 0.009652f
C4714 vdd.n1925 gnd 0.005214f
C4715 vdd.n1926 gnd 0.006754f
C4716 vdd.n1928 gnd 0.006754f
C4717 vdd.n1929 gnd 0.016025f
C4718 vdd.n1930 gnd 0.016025f
C4719 vdd.n1931 gnd 0.014962f
C4720 vdd.n1932 gnd 0.006754f
C4721 vdd.n1933 gnd 0.006754f
C4722 vdd.n1934 gnd 0.006754f
C4723 vdd.n1935 gnd 0.006754f
C4724 vdd.n1936 gnd 0.006754f
C4725 vdd.n1937 gnd 0.006754f
C4726 vdd.n1938 gnd 0.006754f
C4727 vdd.n1939 gnd 0.006754f
C4728 vdd.n1940 gnd 0.006754f
C4729 vdd.n1941 gnd 0.006754f
C4730 vdd.n1942 gnd 0.006754f
C4731 vdd.n1943 gnd 0.006754f
C4732 vdd.n1944 gnd 0.006754f
C4733 vdd.n1945 gnd 0.006754f
C4734 vdd.n1946 gnd 0.006754f
C4735 vdd.n1947 gnd 0.006754f
C4736 vdd.n1948 gnd 0.006754f
C4737 vdd.n1949 gnd 0.006754f
C4738 vdd.n1950 gnd 0.006754f
C4739 vdd.n1951 gnd 0.006754f
C4740 vdd.n1952 gnd 0.006754f
C4741 vdd.n1953 gnd 0.006754f
C4742 vdd.n1954 gnd 0.006754f
C4743 vdd.n1955 gnd 0.006754f
C4744 vdd.n1956 gnd 0.006754f
C4745 vdd.n1957 gnd 0.006754f
C4746 vdd.n1958 gnd 0.006754f
C4747 vdd.n1959 gnd 0.006754f
C4748 vdd.n1960 gnd 0.006754f
C4749 vdd.n1961 gnd 0.006754f
C4750 vdd.n1962 gnd 0.006754f
C4751 vdd.n1963 gnd 0.006754f
C4752 vdd.n1964 gnd 0.006754f
C4753 vdd.n1965 gnd 0.006754f
C4754 vdd.n1966 gnd 0.006754f
C4755 vdd.n1967 gnd 0.006754f
C4756 vdd.n1968 gnd 0.006754f
C4757 vdd.n1969 gnd 0.21822f
C4758 vdd.n1970 gnd 0.006754f
C4759 vdd.n1971 gnd 0.006754f
C4760 vdd.n1972 gnd 0.006754f
C4761 vdd.n1973 gnd 0.006754f
C4762 vdd.n1974 gnd 0.006754f
C4763 vdd.n1975 gnd 0.006754f
C4764 vdd.n1976 gnd 0.006754f
C4765 vdd.n1977 gnd 0.006754f
C4766 vdd.n1978 gnd 0.006754f
C4767 vdd.n1979 gnd 0.006754f
C4768 vdd.n1980 gnd 0.006754f
C4769 vdd.n1981 gnd 0.006754f
C4770 vdd.n1982 gnd 0.006754f
C4771 vdd.n1983 gnd 0.006754f
C4772 vdd.n1984 gnd 0.006754f
C4773 vdd.n1985 gnd 0.006754f
C4774 vdd.n1986 gnd 0.006754f
C4775 vdd.n1987 gnd 0.006754f
C4776 vdd.n1988 gnd 0.006754f
C4777 vdd.n1989 gnd 0.006754f
C4778 vdd.n1990 gnd 0.014962f
C4779 vdd.n1992 gnd 0.016025f
C4780 vdd.n1993 gnd 0.016025f
C4781 vdd.n1994 gnd 0.006754f
C4782 vdd.n1995 gnd 0.005214f
C4783 vdd.n1996 gnd 0.006754f
C4784 vdd.n1998 gnd 0.006754f
C4785 vdd.n2000 gnd 0.006754f
C4786 vdd.n2001 gnd 0.006754f
C4787 vdd.n2002 gnd 0.006754f
C4788 vdd.n2003 gnd 0.006754f
C4789 vdd.n2004 gnd 0.006754f
C4790 vdd.n2006 gnd 0.006754f
C4791 vdd.n2008 gnd 0.006754f
C4792 vdd.n2009 gnd 0.006754f
C4793 vdd.n2010 gnd 0.006754f
C4794 vdd.n2011 gnd 0.006754f
C4795 vdd.n2012 gnd 0.006754f
C4796 vdd.n2014 gnd 0.006754f
C4797 vdd.n2016 gnd 0.006754f
C4798 vdd.n2017 gnd 0.006754f
C4799 vdd.n2018 gnd 0.006754f
C4800 vdd.n2019 gnd 0.006754f
C4801 vdd.n2020 gnd 0.006754f
C4802 vdd.n2022 gnd 0.006754f
C4803 vdd.n2024 gnd 0.006754f
C4804 vdd.n2025 gnd 0.006754f
C4805 vdd.n2026 gnd 0.020145f
C4806 vdd.n2027 gnd 0.59717f
C4807 vdd.n2029 gnd 0.007994f
C4808 vdd.n2030 gnd 0.007994f
C4809 vdd.n2031 gnd 0.009932f
C4810 vdd.n2033 gnd 0.009932f
C4811 vdd.n2034 gnd 0.009932f
C4812 vdd.n2035 gnd 0.007994f
C4813 vdd.n2036 gnd 0.006635f
C4814 vdd.n2037 gnd 0.023771f
C4815 vdd.n2038 gnd 0.023405f
C4816 vdd.n2039 gnd 0.006635f
C4817 vdd.n2040 gnd 0.023405f
C4818 vdd.n2041 gnd 1.39559f
C4819 vdd.n2042 gnd 0.023405f
C4820 vdd.n2043 gnd 0.023771f
C4821 vdd.n2044 gnd 0.003797f
C4822 vdd.t25 gnd 0.122186f
C4823 vdd.t24 gnd 0.130584f
C4824 vdd.t22 gnd 0.159574f
C4825 vdd.n2045 gnd 0.204551f
C4826 vdd.n2046 gnd 0.17186f
C4827 vdd.n2047 gnd 0.01231f
C4828 vdd.n2048 gnd 0.004197f
C4829 vdd.n2049 gnd 0.008541f
C4830 vdd.n2050 gnd 0.59717f
C4831 vdd.n2051 gnd 0.020145f
C4832 vdd.n2052 gnd 0.006754f
C4833 vdd.n2053 gnd 0.006754f
C4834 vdd.n2054 gnd 0.006754f
C4835 vdd.n2056 gnd 0.006754f
C4836 vdd.n2058 gnd 0.006754f
C4837 vdd.n2059 gnd 0.006754f
C4838 vdd.n2060 gnd 0.006754f
C4839 vdd.n2061 gnd 0.006754f
C4840 vdd.n2062 gnd 0.006754f
C4841 vdd.n2064 gnd 0.006754f
C4842 vdd.n2066 gnd 0.006754f
C4843 vdd.n2067 gnd 0.006754f
C4844 vdd.n2068 gnd 0.006754f
C4845 vdd.n2069 gnd 0.006754f
C4846 vdd.n2070 gnd 0.006754f
C4847 vdd.n2072 gnd 0.006754f
C4848 vdd.n2074 gnd 0.006754f
C4849 vdd.n2075 gnd 0.006754f
C4850 vdd.n2076 gnd 0.006754f
C4851 vdd.n2077 gnd 0.006754f
C4852 vdd.n2078 gnd 0.006754f
C4853 vdd.n2080 gnd 0.006754f
C4854 vdd.n2082 gnd 0.006754f
C4855 vdd.n2083 gnd 0.006754f
C4856 vdd.n2084 gnd 0.016025f
C4857 vdd.n2085 gnd 0.014962f
C4858 vdd.n2086 gnd 0.014962f
C4859 vdd.n2087 gnd 0.994677f
C4860 vdd.n2088 gnd 0.014962f
C4861 vdd.n2089 gnd 0.014962f
C4862 vdd.n2090 gnd 0.006754f
C4863 vdd.n2091 gnd 0.006754f
C4864 vdd.n2092 gnd 0.006754f
C4865 vdd.n2093 gnd 0.431365f
C4866 vdd.n2094 gnd 0.006754f
C4867 vdd.n2095 gnd 0.006754f
C4868 vdd.n2096 gnd 0.006754f
C4869 vdd.n2097 gnd 0.006754f
C4870 vdd.n2098 gnd 0.006754f
C4871 vdd.n2099 gnd 0.690184f
C4872 vdd.n2100 gnd 0.006754f
C4873 vdd.n2101 gnd 0.006754f
C4874 vdd.n2102 gnd 0.006754f
C4875 vdd.n2103 gnd 0.006754f
C4876 vdd.n2104 gnd 0.006754f
C4877 vdd.n2105 gnd 0.690184f
C4878 vdd.n2106 gnd 0.006754f
C4879 vdd.n2107 gnd 0.006754f
C4880 vdd.n2108 gnd 0.005959f
C4881 vdd.n2109 gnd 0.019564f
C4882 vdd.n2110 gnd 0.004171f
C4883 vdd.n2111 gnd 0.006754f
C4884 vdd.n2112 gnd 0.380616f
C4885 vdd.n2113 gnd 0.006754f
C4886 vdd.n2114 gnd 0.006754f
C4887 vdd.n2115 gnd 0.006754f
C4888 vdd.n2116 gnd 0.006754f
C4889 vdd.n2117 gnd 0.006754f
C4890 vdd.n2118 gnd 0.461814f
C4891 vdd.n2119 gnd 0.006754f
C4892 vdd.n2120 gnd 0.006754f
C4893 vdd.n2121 gnd 0.006754f
C4894 vdd.n2122 gnd 0.006754f
C4895 vdd.n2123 gnd 0.006754f
C4896 vdd.n2124 gnd 0.614061f
C4897 vdd.n2125 gnd 0.006754f
C4898 vdd.n2126 gnd 0.006754f
C4899 vdd.n2127 gnd 0.006754f
C4900 vdd.n2128 gnd 0.006754f
C4901 vdd.n2129 gnd 0.006754f
C4902 vdd.n2130 gnd 0.548087f
C4903 vdd.n2131 gnd 0.006754f
C4904 vdd.n2132 gnd 0.006754f
C4905 vdd.n2133 gnd 0.006754f
C4906 vdd.n2134 gnd 0.006754f
C4907 vdd.n2135 gnd 0.006754f
C4908 vdd.n2136 gnd 0.395841f
C4909 vdd.n2137 gnd 0.006754f
C4910 vdd.n2138 gnd 0.006754f
C4911 vdd.n2139 gnd 0.006754f
C4912 vdd.n2140 gnd 0.006754f
C4913 vdd.n2141 gnd 0.006754f
C4914 vdd.n2142 gnd 0.21822f
C4915 vdd.n2143 gnd 0.006754f
C4916 vdd.n2144 gnd 0.006754f
C4917 vdd.n2145 gnd 0.006754f
C4918 vdd.n2146 gnd 0.006754f
C4919 vdd.n2147 gnd 0.006754f
C4920 vdd.n2148 gnd 0.380616f
C4921 vdd.n2149 gnd 0.006754f
C4922 vdd.n2150 gnd 0.006754f
C4923 vdd.n2151 gnd 0.006754f
C4924 vdd.n2152 gnd 0.006754f
C4925 vdd.n2153 gnd 0.006754f
C4926 vdd.n2154 gnd 0.690184f
C4927 vdd.n2155 gnd 0.006754f
C4928 vdd.n2156 gnd 0.006754f
C4929 vdd.n2157 gnd 0.006754f
C4930 vdd.n2158 gnd 0.006754f
C4931 vdd.n2159 gnd 0.006754f
C4932 vdd.n2160 gnd 0.006754f
C4933 vdd.n2161 gnd 0.006754f
C4934 vdd.n2162 gnd 0.537938f
C4935 vdd.n2163 gnd 0.006754f
C4936 vdd.n2164 gnd 0.006754f
C4937 vdd.n2165 gnd 0.006754f
C4938 vdd.n2166 gnd 0.006754f
C4939 vdd.n2167 gnd 0.006754f
C4940 vdd.n2168 gnd 0.006754f
C4941 vdd.n2169 gnd 0.431365f
C4942 vdd.n2170 gnd 0.006754f
C4943 vdd.n2171 gnd 0.006754f
C4944 vdd.n2172 gnd 0.006754f
C4945 vdd.n2173 gnd 0.015784f
C4946 vdd.n2174 gnd 0.015203f
C4947 vdd.n2175 gnd 0.006754f
C4948 vdd.n2176 gnd 0.006754f
C4949 vdd.n2177 gnd 0.005214f
C4950 vdd.n2178 gnd 0.006754f
C4951 vdd.n2179 gnd 0.006754f
C4952 vdd.n2180 gnd 0.004916f
C4953 vdd.n2181 gnd 0.006754f
C4954 vdd.n2182 gnd 0.006754f
C4955 vdd.n2183 gnd 0.006754f
C4956 vdd.n2184 gnd 0.006754f
C4957 vdd.n2185 gnd 0.006754f
C4958 vdd.n2186 gnd 0.006754f
C4959 vdd.n2187 gnd 0.006754f
C4960 vdd.n2188 gnd 0.006754f
C4961 vdd.n2189 gnd 0.006754f
C4962 vdd.n2190 gnd 0.006754f
C4963 vdd.n2191 gnd 0.006754f
C4964 vdd.n2192 gnd 0.006754f
C4965 vdd.n2193 gnd 0.006754f
C4966 vdd.n2194 gnd 0.006754f
C4967 vdd.n2195 gnd 0.006754f
C4968 vdd.n2196 gnd 0.006754f
C4969 vdd.n2197 gnd 0.006754f
C4970 vdd.n2198 gnd 0.006754f
C4971 vdd.n2199 gnd 0.006754f
C4972 vdd.n2200 gnd 0.006754f
C4973 vdd.n2201 gnd 0.006754f
C4974 vdd.n2202 gnd 0.006754f
C4975 vdd.n2203 gnd 0.006754f
C4976 vdd.n2204 gnd 0.006754f
C4977 vdd.n2205 gnd 0.006754f
C4978 vdd.n2206 gnd 0.006754f
C4979 vdd.n2207 gnd 0.006754f
C4980 vdd.n2208 gnd 0.006754f
C4981 vdd.n2209 gnd 0.006754f
C4982 vdd.n2210 gnd 0.006754f
C4983 vdd.n2211 gnd 0.006754f
C4984 vdd.n2212 gnd 0.006754f
C4985 vdd.n2213 gnd 0.006754f
C4986 vdd.n2214 gnd 0.006754f
C4987 vdd.n2215 gnd 0.006754f
C4988 vdd.n2216 gnd 0.006754f
C4989 vdd.n2217 gnd 0.006754f
C4990 vdd.n2218 gnd 0.006754f
C4991 vdd.n2219 gnd 0.006754f
C4992 vdd.n2220 gnd 0.006754f
C4993 vdd.n2221 gnd 0.006754f
C4994 vdd.n2222 gnd 0.006754f
C4995 vdd.n2223 gnd 0.006754f
C4996 vdd.n2224 gnd 0.006754f
C4997 vdd.n2225 gnd 0.006754f
C4998 vdd.n2226 gnd 0.006754f
C4999 vdd.n2227 gnd 0.006754f
C5000 vdd.n2228 gnd 0.006754f
C5001 vdd.n2229 gnd 0.006754f
C5002 vdd.n2230 gnd 0.006754f
C5003 vdd.n2231 gnd 0.006754f
C5004 vdd.n2232 gnd 0.006754f
C5005 vdd.n2233 gnd 0.006754f
C5006 vdd.n2234 gnd 0.006754f
C5007 vdd.n2235 gnd 0.006754f
C5008 vdd.n2236 gnd 0.006754f
C5009 vdd.n2237 gnd 0.006754f
C5010 vdd.n2238 gnd 0.006754f
C5011 vdd.n2239 gnd 0.006754f
C5012 vdd.n2240 gnd 0.006754f
C5013 vdd.n2241 gnd 0.016025f
C5014 vdd.n2242 gnd 0.014962f
C5015 vdd.n2243 gnd 0.014962f
C5016 vdd.n2244 gnd 0.84243f
C5017 vdd.n2245 gnd 0.014962f
C5018 vdd.n2246 gnd 0.016025f
C5019 vdd.n2247 gnd 0.015203f
C5020 vdd.n2248 gnd 0.006754f
C5021 vdd.n2249 gnd 0.006754f
C5022 vdd.n2250 gnd 0.006754f
C5023 vdd.n2251 gnd 0.005214f
C5024 vdd.n2252 gnd 0.009652f
C5025 vdd.n2253 gnd 0.004916f
C5026 vdd.n2254 gnd 0.006754f
C5027 vdd.n2255 gnd 0.006754f
C5028 vdd.n2256 gnd 0.006754f
C5029 vdd.n2257 gnd 0.006754f
C5030 vdd.n2258 gnd 0.006754f
C5031 vdd.n2259 gnd 0.006754f
C5032 vdd.n2260 gnd 0.006754f
C5033 vdd.n2261 gnd 0.006754f
C5034 vdd.n2262 gnd 0.006754f
C5035 vdd.n2263 gnd 0.006754f
C5036 vdd.n2264 gnd 0.006754f
C5037 vdd.n2265 gnd 0.006754f
C5038 vdd.n2266 gnd 0.006754f
C5039 vdd.n2267 gnd 0.006754f
C5040 vdd.n2268 gnd 0.006754f
C5041 vdd.n2269 gnd 0.006754f
C5042 vdd.n2270 gnd 0.006754f
C5043 vdd.n2271 gnd 0.006754f
C5044 vdd.n2272 gnd 0.006754f
C5045 vdd.n2273 gnd 0.006754f
C5046 vdd.n2274 gnd 0.006754f
C5047 vdd.n2275 gnd 0.006754f
C5048 vdd.n2276 gnd 0.006754f
C5049 vdd.n2277 gnd 0.006754f
C5050 vdd.n2278 gnd 0.006754f
C5051 vdd.n2279 gnd 0.006754f
C5052 vdd.n2280 gnd 0.006754f
C5053 vdd.n2281 gnd 0.006754f
C5054 vdd.n2282 gnd 0.006754f
C5055 vdd.n2283 gnd 0.006754f
C5056 vdd.n2284 gnd 0.006754f
C5057 vdd.n2285 gnd 0.006754f
C5058 vdd.n2286 gnd 0.006754f
C5059 vdd.n2287 gnd 0.006754f
C5060 vdd.n2288 gnd 0.006754f
C5061 vdd.n2289 gnd 0.006754f
C5062 vdd.n2290 gnd 0.006754f
C5063 vdd.n2291 gnd 0.006754f
C5064 vdd.n2292 gnd 0.006754f
C5065 vdd.n2293 gnd 0.006754f
C5066 vdd.n2294 gnd 0.006754f
C5067 vdd.n2295 gnd 0.006754f
C5068 vdd.n2296 gnd 0.006754f
C5069 vdd.n2297 gnd 0.006754f
C5070 vdd.n2298 gnd 0.006754f
C5071 vdd.n2299 gnd 0.006754f
C5072 vdd.n2300 gnd 0.006754f
C5073 vdd.n2301 gnd 0.006754f
C5074 vdd.n2302 gnd 0.006754f
C5075 vdd.n2303 gnd 0.006754f
C5076 vdd.n2304 gnd 0.006754f
C5077 vdd.n2305 gnd 0.006754f
C5078 vdd.n2306 gnd 0.006754f
C5079 vdd.n2307 gnd 0.006754f
C5080 vdd.n2308 gnd 0.006754f
C5081 vdd.n2309 gnd 0.006754f
C5082 vdd.n2310 gnd 0.006754f
C5083 vdd.n2311 gnd 0.006754f
C5084 vdd.n2312 gnd 0.006754f
C5085 vdd.n2313 gnd 0.006754f
C5086 vdd.n2314 gnd 0.016025f
C5087 vdd.n2315 gnd 0.016025f
C5088 vdd.n2316 gnd 0.84243f
C5089 vdd.t228 gnd 2.99418f
C5090 vdd.t111 gnd 2.99418f
C5091 vdd.n2349 gnd 0.016025f
C5092 vdd.n2350 gnd 0.006754f
C5093 vdd.t52 gnd 0.272911f
C5094 vdd.t53 gnd 0.279359f
C5095 vdd.t50 gnd 0.178167f
C5096 vdd.n2351 gnd 0.096289f
C5097 vdd.n2352 gnd 0.054619f
C5098 vdd.n2353 gnd 0.006754f
C5099 vdd.t65 gnd 0.272911f
C5100 vdd.t66 gnd 0.279359f
C5101 vdd.t64 gnd 0.178167f
C5102 vdd.n2354 gnd 0.096289f
C5103 vdd.n2355 gnd 0.054619f
C5104 vdd.n2356 gnd 0.009652f
C5105 vdd.n2357 gnd 0.006754f
C5106 vdd.n2358 gnd 0.006754f
C5107 vdd.n2359 gnd 0.006754f
C5108 vdd.n2360 gnd 0.006754f
C5109 vdd.n2361 gnd 0.006754f
C5110 vdd.n2362 gnd 0.006754f
C5111 vdd.n2363 gnd 0.006754f
C5112 vdd.n2364 gnd 0.006754f
C5113 vdd.n2365 gnd 0.006754f
C5114 vdd.n2366 gnd 0.006754f
C5115 vdd.n2367 gnd 0.006754f
C5116 vdd.n2368 gnd 0.006754f
C5117 vdd.n2369 gnd 0.006754f
C5118 vdd.n2370 gnd 0.006754f
C5119 vdd.n2371 gnd 0.006754f
C5120 vdd.n2372 gnd 0.006754f
C5121 vdd.n2373 gnd 0.006754f
C5122 vdd.n2374 gnd 0.006754f
C5123 vdd.n2375 gnd 0.006754f
C5124 vdd.n2376 gnd 0.006754f
C5125 vdd.n2377 gnd 0.006754f
C5126 vdd.n2378 gnd 0.006754f
C5127 vdd.n2379 gnd 0.006754f
C5128 vdd.n2380 gnd 0.006754f
C5129 vdd.n2381 gnd 0.006754f
C5130 vdd.n2382 gnd 0.006754f
C5131 vdd.n2383 gnd 0.006754f
C5132 vdd.n2384 gnd 0.006754f
C5133 vdd.n2385 gnd 0.006754f
C5134 vdd.n2386 gnd 0.006754f
C5135 vdd.n2387 gnd 0.006754f
C5136 vdd.n2388 gnd 0.006754f
C5137 vdd.n2389 gnd 0.006754f
C5138 vdd.n2390 gnd 0.006754f
C5139 vdd.n2391 gnd 0.006754f
C5140 vdd.n2392 gnd 0.006754f
C5141 vdd.n2393 gnd 0.006754f
C5142 vdd.n2394 gnd 0.006754f
C5143 vdd.n2395 gnd 0.006754f
C5144 vdd.n2396 gnd 0.006754f
C5145 vdd.n2397 gnd 0.006754f
C5146 vdd.n2398 gnd 0.006754f
C5147 vdd.n2399 gnd 0.006754f
C5148 vdd.n2400 gnd 0.006754f
C5149 vdd.n2401 gnd 0.006754f
C5150 vdd.n2402 gnd 0.006754f
C5151 vdd.n2403 gnd 0.006754f
C5152 vdd.n2404 gnd 0.006754f
C5153 vdd.n2405 gnd 0.006754f
C5154 vdd.n2406 gnd 0.006754f
C5155 vdd.n2407 gnd 0.006754f
C5156 vdd.n2408 gnd 0.006754f
C5157 vdd.n2409 gnd 0.006754f
C5158 vdd.n2410 gnd 0.006754f
C5159 vdd.n2411 gnd 0.006754f
C5160 vdd.n2412 gnd 0.006754f
C5161 vdd.n2413 gnd 0.004916f
C5162 vdd.n2414 gnd 0.006754f
C5163 vdd.n2415 gnd 0.006754f
C5164 vdd.n2416 gnd 0.005214f
C5165 vdd.n2417 gnd 0.006754f
C5166 vdd.n2418 gnd 0.006754f
C5167 vdd.n2419 gnd 0.016025f
C5168 vdd.n2420 gnd 0.014962f
C5169 vdd.n2421 gnd 0.006754f
C5170 vdd.n2422 gnd 0.006754f
C5171 vdd.n2423 gnd 0.006754f
C5172 vdd.n2424 gnd 0.006754f
C5173 vdd.n2425 gnd 0.006754f
C5174 vdd.n2426 gnd 0.006754f
C5175 vdd.n2427 gnd 0.006754f
C5176 vdd.n2428 gnd 0.006754f
C5177 vdd.n2429 gnd 0.006754f
C5178 vdd.n2430 gnd 0.006754f
C5179 vdd.n2431 gnd 0.006754f
C5180 vdd.n2432 gnd 0.006754f
C5181 vdd.n2433 gnd 0.006754f
C5182 vdd.n2434 gnd 0.006754f
C5183 vdd.n2435 gnd 0.006754f
C5184 vdd.n2436 gnd 0.006754f
C5185 vdd.n2437 gnd 0.006754f
C5186 vdd.n2438 gnd 0.006754f
C5187 vdd.n2439 gnd 0.006754f
C5188 vdd.n2440 gnd 0.006754f
C5189 vdd.n2441 gnd 0.006754f
C5190 vdd.n2442 gnd 0.006754f
C5191 vdd.n2443 gnd 0.006754f
C5192 vdd.n2444 gnd 0.006754f
C5193 vdd.n2445 gnd 0.006754f
C5194 vdd.n2446 gnd 0.006754f
C5195 vdd.n2447 gnd 0.006754f
C5196 vdd.n2448 gnd 0.006754f
C5197 vdd.n2449 gnd 0.006754f
C5198 vdd.n2450 gnd 0.006754f
C5199 vdd.n2451 gnd 0.006754f
C5200 vdd.n2452 gnd 0.006754f
C5201 vdd.n2453 gnd 0.006754f
C5202 vdd.n2454 gnd 0.006754f
C5203 vdd.n2455 gnd 0.006754f
C5204 vdd.n2456 gnd 0.006754f
C5205 vdd.n2457 gnd 0.006754f
C5206 vdd.n2458 gnd 0.006754f
C5207 vdd.n2459 gnd 0.006754f
C5208 vdd.n2460 gnd 0.006754f
C5209 vdd.n2461 gnd 0.006754f
C5210 vdd.n2462 gnd 0.006754f
C5211 vdd.n2463 gnd 0.006754f
C5212 vdd.n2464 gnd 0.006754f
C5213 vdd.n2465 gnd 0.006754f
C5214 vdd.n2466 gnd 0.006754f
C5215 vdd.n2467 gnd 0.006754f
C5216 vdd.n2468 gnd 0.006754f
C5217 vdd.n2469 gnd 0.006754f
C5218 vdd.n2470 gnd 0.006754f
C5219 vdd.n2471 gnd 0.006754f
C5220 vdd.n2472 gnd 0.21822f
C5221 vdd.n2473 gnd 0.006754f
C5222 vdd.n2474 gnd 0.006754f
C5223 vdd.n2475 gnd 0.006754f
C5224 vdd.n2476 gnd 0.006754f
C5225 vdd.n2477 gnd 0.006754f
C5226 vdd.n2478 gnd 0.006754f
C5227 vdd.n2479 gnd 0.006754f
C5228 vdd.n2480 gnd 0.006754f
C5229 vdd.n2481 gnd 0.006754f
C5230 vdd.n2482 gnd 0.006754f
C5231 vdd.n2483 gnd 0.006754f
C5232 vdd.n2484 gnd 0.006754f
C5233 vdd.n2485 gnd 0.006754f
C5234 vdd.n2486 gnd 0.006754f
C5235 vdd.n2487 gnd 0.006754f
C5236 vdd.n2488 gnd 0.006754f
C5237 vdd.n2489 gnd 0.006754f
C5238 vdd.n2490 gnd 0.006754f
C5239 vdd.n2491 gnd 0.006754f
C5240 vdd.n2492 gnd 0.006754f
C5241 vdd.n2493 gnd 0.411065f
C5242 vdd.n2494 gnd 0.006754f
C5243 vdd.n2495 gnd 0.006754f
C5244 vdd.n2496 gnd 0.006754f
C5245 vdd.n2497 gnd 0.006754f
C5246 vdd.n2498 gnd 0.006754f
C5247 vdd.n2499 gnd 0.014962f
C5248 vdd.n2500 gnd 0.016025f
C5249 vdd.n2501 gnd 0.016025f
C5250 vdd.n2502 gnd 0.006754f
C5251 vdd.n2503 gnd 0.006754f
C5252 vdd.n2504 gnd 0.006754f
C5253 vdd.n2505 gnd 0.005214f
C5254 vdd.n2506 gnd 0.009652f
C5255 vdd.n2507 gnd 0.004916f
C5256 vdd.n2508 gnd 0.006754f
C5257 vdd.n2509 gnd 0.006754f
C5258 vdd.n2510 gnd 0.006754f
C5259 vdd.n2511 gnd 0.006754f
C5260 vdd.n2512 gnd 0.006754f
C5261 vdd.n2513 gnd 0.006754f
C5262 vdd.n2514 gnd 0.006754f
C5263 vdd.n2515 gnd 0.006754f
C5264 vdd.n2516 gnd 0.006754f
C5265 vdd.n2517 gnd 0.006754f
C5266 vdd.n2518 gnd 0.006754f
C5267 vdd.n2519 gnd 0.006754f
C5268 vdd.n2520 gnd 0.006754f
C5269 vdd.n2521 gnd 0.006754f
C5270 vdd.n2522 gnd 0.006754f
C5271 vdd.n2523 gnd 0.006754f
C5272 vdd.n2524 gnd 0.006754f
C5273 vdd.n2525 gnd 0.006754f
C5274 vdd.n2526 gnd 0.006754f
C5275 vdd.n2527 gnd 0.006754f
C5276 vdd.n2528 gnd 0.006754f
C5277 vdd.n2529 gnd 0.006754f
C5278 vdd.n2530 gnd 0.006754f
C5279 vdd.n2531 gnd 0.006754f
C5280 vdd.n2532 gnd 0.006754f
C5281 vdd.n2533 gnd 0.006754f
C5282 vdd.n2534 gnd 0.006754f
C5283 vdd.n2535 gnd 0.006754f
C5284 vdd.n2536 gnd 0.006754f
C5285 vdd.n2537 gnd 0.006754f
C5286 vdd.n2538 gnd 0.006754f
C5287 vdd.n2539 gnd 0.006754f
C5288 vdd.n2540 gnd 0.006754f
C5289 vdd.n2541 gnd 0.006754f
C5290 vdd.n2542 gnd 0.006754f
C5291 vdd.n2543 gnd 0.006754f
C5292 vdd.n2544 gnd 0.006754f
C5293 vdd.n2545 gnd 0.006754f
C5294 vdd.n2546 gnd 0.006754f
C5295 vdd.n2547 gnd 0.006754f
C5296 vdd.n2548 gnd 0.006754f
C5297 vdd.n2549 gnd 0.006754f
C5298 vdd.n2550 gnd 0.006754f
C5299 vdd.n2551 gnd 0.006754f
C5300 vdd.n2552 gnd 0.006754f
C5301 vdd.n2553 gnd 0.006754f
C5302 vdd.n2554 gnd 0.006754f
C5303 vdd.n2555 gnd 0.006754f
C5304 vdd.n2556 gnd 0.006754f
C5305 vdd.n2557 gnd 0.006754f
C5306 vdd.n2558 gnd 0.006754f
C5307 vdd.n2559 gnd 0.006754f
C5308 vdd.n2560 gnd 0.006754f
C5309 vdd.n2561 gnd 0.006754f
C5310 vdd.n2562 gnd 0.006754f
C5311 vdd.n2563 gnd 0.006754f
C5312 vdd.n2564 gnd 0.006754f
C5313 vdd.n2565 gnd 0.006754f
C5314 vdd.n2566 gnd 0.006754f
C5315 vdd.n2567 gnd 0.006754f
C5316 vdd.n2569 gnd 0.84243f
C5317 vdd.n2571 gnd 0.006754f
C5318 vdd.n2572 gnd 0.006754f
C5319 vdd.n2573 gnd 0.016025f
C5320 vdd.n2574 gnd 0.014962f
C5321 vdd.n2575 gnd 0.014962f
C5322 vdd.n2576 gnd 0.84243f
C5323 vdd.n2577 gnd 0.014962f
C5324 vdd.n2578 gnd 0.014962f
C5325 vdd.n2579 gnd 0.006754f
C5326 vdd.n2580 gnd 0.006754f
C5327 vdd.n2581 gnd 0.006754f
C5328 vdd.n2582 gnd 0.431365f
C5329 vdd.n2583 gnd 0.006754f
C5330 vdd.n2584 gnd 0.006754f
C5331 vdd.n2585 gnd 0.006754f
C5332 vdd.n2586 gnd 0.006754f
C5333 vdd.n2587 gnd 0.006754f
C5334 vdd.n2588 gnd 0.537938f
C5335 vdd.n2589 gnd 0.006754f
C5336 vdd.n2590 gnd 0.006754f
C5337 vdd.n2591 gnd 0.006754f
C5338 vdd.n2592 gnd 0.006754f
C5339 vdd.n2593 gnd 0.006754f
C5340 vdd.n2594 gnd 0.690184f
C5341 vdd.n2595 gnd 0.006754f
C5342 vdd.n2596 gnd 0.006754f
C5343 vdd.n2597 gnd 0.006754f
C5344 vdd.n2598 gnd 0.006754f
C5345 vdd.n2599 gnd 0.006754f
C5346 vdd.n2600 gnd 0.380616f
C5347 vdd.n2601 gnd 0.006754f
C5348 vdd.n2602 gnd 0.006754f
C5349 vdd.n2603 gnd 0.006754f
C5350 vdd.n2604 gnd 0.006754f
C5351 vdd.n2605 gnd 0.006754f
C5352 vdd.n2606 gnd 0.21822f
C5353 vdd.n2607 gnd 0.006754f
C5354 vdd.n2608 gnd 0.006754f
C5355 vdd.n2609 gnd 0.006754f
C5356 vdd.n2610 gnd 0.006754f
C5357 vdd.n2611 gnd 0.006754f
C5358 vdd.n2612 gnd 0.395841f
C5359 vdd.n2613 gnd 0.006754f
C5360 vdd.n2614 gnd 0.006754f
C5361 vdd.n2615 gnd 0.006754f
C5362 vdd.n2616 gnd 0.006754f
C5363 vdd.n2617 gnd 0.006754f
C5364 vdd.n2618 gnd 0.548087f
C5365 vdd.n2619 gnd 0.006754f
C5366 vdd.n2620 gnd 0.006754f
C5367 vdd.n2621 gnd 0.006754f
C5368 vdd.n2622 gnd 0.006754f
C5369 vdd.n2623 gnd 0.006754f
C5370 vdd.n2624 gnd 0.614061f
C5371 vdd.n2625 gnd 0.006754f
C5372 vdd.n2626 gnd 0.006754f
C5373 vdd.n2627 gnd 0.006754f
C5374 vdd.n2628 gnd 0.006754f
C5375 vdd.n2629 gnd 0.006754f
C5376 vdd.n2630 gnd 0.461814f
C5377 vdd.n2631 gnd 0.006754f
C5378 vdd.n2632 gnd 0.006754f
C5379 vdd.n2633 gnd 0.006754f
C5380 vdd.t31 gnd 0.279359f
C5381 vdd.t29 gnd 0.178167f
C5382 vdd.t32 gnd 0.279359f
C5383 vdd.n2634 gnd 0.157011f
C5384 vdd.n2635 gnd 0.019564f
C5385 vdd.n2636 gnd 0.004171f
C5386 vdd.n2637 gnd 0.006754f
C5387 vdd.n2638 gnd 0.380616f
C5388 vdd.n2639 gnd 0.006754f
C5389 vdd.n2640 gnd 0.006754f
C5390 vdd.n2641 gnd 0.006754f
C5391 vdd.n2642 gnd 0.006754f
C5392 vdd.n2643 gnd 0.006754f
C5393 vdd.n2644 gnd 0.690184f
C5394 vdd.n2645 gnd 0.006754f
C5395 vdd.n2646 gnd 0.006754f
C5396 vdd.n2647 gnd 0.006754f
C5397 vdd.n2648 gnd 0.006754f
C5398 vdd.n2649 gnd 0.006754f
C5399 vdd.n2650 gnd 0.006754f
C5400 vdd.n2652 gnd 0.006754f
C5401 vdd.n2653 gnd 0.006754f
C5402 vdd.n2655 gnd 0.006754f
C5403 vdd.n2656 gnd 0.006754f
C5404 vdd.n2659 gnd 0.006754f
C5405 vdd.n2660 gnd 0.006754f
C5406 vdd.n2661 gnd 0.006754f
C5407 vdd.n2662 gnd 0.006754f
C5408 vdd.n2664 gnd 0.006754f
C5409 vdd.n2665 gnd 0.006754f
C5410 vdd.n2666 gnd 0.006754f
C5411 vdd.n2667 gnd 0.006754f
C5412 vdd.n2668 gnd 0.006754f
C5413 vdd.n2669 gnd 0.006754f
C5414 vdd.n2671 gnd 0.006754f
C5415 vdd.n2672 gnd 0.006754f
C5416 vdd.n2673 gnd 0.006754f
C5417 vdd.n2674 gnd 0.006754f
C5418 vdd.n2675 gnd 0.006754f
C5419 vdd.n2676 gnd 0.006754f
C5420 vdd.n2678 gnd 0.006754f
C5421 vdd.n2679 gnd 0.006754f
C5422 vdd.n2680 gnd 0.006754f
C5423 vdd.n2681 gnd 0.006754f
C5424 vdd.n2682 gnd 0.006754f
C5425 vdd.n2683 gnd 0.006754f
C5426 vdd.n2685 gnd 0.006754f
C5427 vdd.n2686 gnd 0.016025f
C5428 vdd.n2687 gnd 0.016025f
C5429 vdd.n2688 gnd 0.014962f
C5430 vdd.n2689 gnd 0.006754f
C5431 vdd.n2690 gnd 0.006754f
C5432 vdd.n2691 gnd 0.006754f
C5433 vdd.n2692 gnd 0.006754f
C5434 vdd.n2693 gnd 0.006754f
C5435 vdd.n2694 gnd 0.006754f
C5436 vdd.n2695 gnd 0.690184f
C5437 vdd.n2696 gnd 0.006754f
C5438 vdd.n2697 gnd 0.006754f
C5439 vdd.n2698 gnd 0.006754f
C5440 vdd.n2699 gnd 0.006754f
C5441 vdd.n2700 gnd 0.006754f
C5442 vdd.n2701 gnd 0.431365f
C5443 vdd.n2702 gnd 0.006754f
C5444 vdd.n2703 gnd 0.006754f
C5445 vdd.n2704 gnd 0.006754f
C5446 vdd.n2705 gnd 0.015784f
C5447 vdd.n2707 gnd 0.016025f
C5448 vdd.n2708 gnd 0.015203f
C5449 vdd.n2709 gnd 0.006754f
C5450 vdd.n2710 gnd 0.005214f
C5451 vdd.n2711 gnd 0.006754f
C5452 vdd.n2713 gnd 0.006754f
C5453 vdd.n2714 gnd 0.006754f
C5454 vdd.n2715 gnd 0.006754f
C5455 vdd.n2716 gnd 0.006754f
C5456 vdd.n2717 gnd 0.006754f
C5457 vdd.n2718 gnd 0.006754f
C5458 vdd.n2720 gnd 0.006754f
C5459 vdd.n2721 gnd 0.006754f
C5460 vdd.n2722 gnd 0.006754f
C5461 vdd.n2723 gnd 0.006754f
C5462 vdd.n2724 gnd 0.006754f
C5463 vdd.n2725 gnd 0.006754f
C5464 vdd.n2727 gnd 0.006754f
C5465 vdd.n2728 gnd 0.006754f
C5466 vdd.n2729 gnd 0.006754f
C5467 vdd.n2730 gnd 0.006754f
C5468 vdd.n2731 gnd 0.006754f
C5469 vdd.n2732 gnd 0.006754f
C5470 vdd.n2734 gnd 0.006754f
C5471 vdd.n2735 gnd 0.006754f
C5472 vdd.n2736 gnd 0.006754f
C5473 vdd.n2737 gnd 0.601085f
C5474 vdd.n2738 gnd 0.016229f
C5475 vdd.n2739 gnd 0.006754f
C5476 vdd.n2740 gnd 0.006754f
C5477 vdd.n2742 gnd 0.006754f
C5478 vdd.n2743 gnd 0.006754f
C5479 vdd.n2744 gnd 0.006754f
C5480 vdd.n2745 gnd 0.006754f
C5481 vdd.n2746 gnd 0.006754f
C5482 vdd.n2747 gnd 0.006754f
C5483 vdd.n2749 gnd 0.006754f
C5484 vdd.n2750 gnd 0.006754f
C5485 vdd.n2751 gnd 0.006754f
C5486 vdd.n2752 gnd 0.006754f
C5487 vdd.n2753 gnd 0.006754f
C5488 vdd.n2754 gnd 0.006754f
C5489 vdd.n2756 gnd 0.006754f
C5490 vdd.n2757 gnd 0.006754f
C5491 vdd.n2758 gnd 0.006754f
C5492 vdd.n2759 gnd 0.006754f
C5493 vdd.n2760 gnd 0.006754f
C5494 vdd.n2761 gnd 0.006754f
C5495 vdd.n2763 gnd 0.006754f
C5496 vdd.n2764 gnd 0.006754f
C5497 vdd.n2766 gnd 0.006754f
C5498 vdd.n2767 gnd 0.006754f
C5499 vdd.n2768 gnd 0.016025f
C5500 vdd.n2769 gnd 0.014962f
C5501 vdd.n2770 gnd 0.014962f
C5502 vdd.n2771 gnd 0.994677f
C5503 vdd.n2772 gnd 0.014962f
C5504 vdd.n2773 gnd 0.016025f
C5505 vdd.n2774 gnd 0.015203f
C5506 vdd.n2775 gnd 0.006754f
C5507 vdd.n2776 gnd 0.005214f
C5508 vdd.n2777 gnd 0.006754f
C5509 vdd.n2779 gnd 0.006754f
C5510 vdd.n2780 gnd 0.006754f
C5511 vdd.n2781 gnd 0.006754f
C5512 vdd.n2782 gnd 0.006754f
C5513 vdd.n2783 gnd 0.006754f
C5514 vdd.n2784 gnd 0.006754f
C5515 vdd.n2786 gnd 0.006754f
C5516 vdd.n2787 gnd 0.006754f
C5517 vdd.n2788 gnd 0.006754f
C5518 vdd.n2789 gnd 0.006754f
C5519 vdd.n2790 gnd 0.006754f
C5520 vdd.n2791 gnd 0.006754f
C5521 vdd.n2793 gnd 0.006754f
C5522 vdd.n2794 gnd 0.006754f
C5523 vdd.n2795 gnd 0.006754f
C5524 vdd.n2796 gnd 0.006754f
C5525 vdd.n2797 gnd 0.006754f
C5526 vdd.n2798 gnd 0.006754f
C5527 vdd.n2800 gnd 0.006754f
C5528 vdd.n2801 gnd 0.006754f
C5529 vdd.n2803 gnd 0.006754f
C5530 vdd.n2804 gnd 0.016229f
C5531 vdd.n2805 gnd 0.601085f
C5532 vdd.n2806 gnd 0.008541f
C5533 vdd.n2807 gnd 0.003797f
C5534 vdd.t71 gnd 0.122186f
C5535 vdd.t72 gnd 0.130584f
C5536 vdd.t70 gnd 0.159574f
C5537 vdd.n2808 gnd 0.204551f
C5538 vdd.n2809 gnd 0.17186f
C5539 vdd.n2810 gnd 0.01231f
C5540 vdd.n2811 gnd 0.009932f
C5541 vdd.n2812 gnd 0.004197f
C5542 vdd.n2813 gnd 0.007994f
C5543 vdd.n2814 gnd 0.009932f
C5544 vdd.n2815 gnd 0.009932f
C5545 vdd.n2816 gnd 0.007994f
C5546 vdd.n2817 gnd 0.007994f
C5547 vdd.n2818 gnd 0.009932f
C5548 vdd.n2820 gnd 0.009932f
C5549 vdd.n2821 gnd 0.007994f
C5550 vdd.n2822 gnd 0.007994f
C5551 vdd.n2823 gnd 0.007994f
C5552 vdd.n2824 gnd 0.009932f
C5553 vdd.n2826 gnd 0.009932f
C5554 vdd.n2828 gnd 0.009932f
C5555 vdd.n2829 gnd 0.007994f
C5556 vdd.n2830 gnd 0.007994f
C5557 vdd.n2831 gnd 0.007994f
C5558 vdd.n2832 gnd 0.009932f
C5559 vdd.n2834 gnd 0.009932f
C5560 vdd.n2836 gnd 0.009932f
C5561 vdd.n2837 gnd 0.007994f
C5562 vdd.n2838 gnd 0.007994f
C5563 vdd.n2839 gnd 0.007994f
C5564 vdd.n2840 gnd 0.009932f
C5565 vdd.n2842 gnd 0.009932f
C5566 vdd.n2843 gnd 0.009932f
C5567 vdd.n2844 gnd 0.007994f
C5568 vdd.n2845 gnd 0.007994f
C5569 vdd.n2846 gnd 0.009932f
C5570 vdd.n2847 gnd 0.009932f
C5571 vdd.n2849 gnd 0.009932f
C5572 vdd.n2850 gnd 0.007994f
C5573 vdd.n2851 gnd 0.009932f
C5574 vdd.n2852 gnd 0.009932f
C5575 vdd.n2853 gnd 0.009932f
C5576 vdd.n2854 gnd 0.016307f
C5577 vdd.n2855 gnd 0.005436f
C5578 vdd.n2856 gnd 0.009932f
C5579 vdd.n2858 gnd 0.009932f
C5580 vdd.n2860 gnd 0.009932f
C5581 vdd.n2861 gnd 0.007994f
C5582 vdd.n2862 gnd 0.007994f
C5583 vdd.n2863 gnd 0.007994f
C5584 vdd.n2864 gnd 0.009932f
C5585 vdd.n2866 gnd 0.009932f
C5586 vdd.n2868 gnd 0.009932f
C5587 vdd.n2869 gnd 0.007994f
C5588 vdd.n2870 gnd 0.007994f
C5589 vdd.n2871 gnd 0.007994f
C5590 vdd.n2872 gnd 0.009932f
C5591 vdd.n2874 gnd 0.009932f
C5592 vdd.n2876 gnd 0.009932f
C5593 vdd.n2877 gnd 0.007994f
C5594 vdd.n2878 gnd 0.007994f
C5595 vdd.n2879 gnd 0.007994f
C5596 vdd.n2880 gnd 0.009932f
C5597 vdd.n2882 gnd 0.009932f
C5598 vdd.n2884 gnd 0.009932f
C5599 vdd.n2885 gnd 0.007994f
C5600 vdd.n2886 gnd 0.007994f
C5601 vdd.n2887 gnd 0.007994f
C5602 vdd.n2888 gnd 0.009932f
C5603 vdd.n2890 gnd 0.009932f
C5604 vdd.n2892 gnd 0.009932f
C5605 vdd.n2893 gnd 0.007994f
C5606 vdd.n2894 gnd 0.007994f
C5607 vdd.n2895 gnd 0.006675f
C5608 vdd.n2896 gnd 0.009932f
C5609 vdd.n2898 gnd 0.009932f
C5610 vdd.n2900 gnd 0.009932f
C5611 vdd.n2901 gnd 0.006675f
C5612 vdd.n2902 gnd 0.007994f
C5613 vdd.n2903 gnd 0.007994f
C5614 vdd.n2904 gnd 0.009932f
C5615 vdd.n2906 gnd 0.009932f
C5616 vdd.n2908 gnd 0.009932f
C5617 vdd.n2909 gnd 0.007994f
C5618 vdd.n2910 gnd 0.007994f
C5619 vdd.n2911 gnd 0.007994f
C5620 vdd.n2912 gnd 0.009932f
C5621 vdd.n2914 gnd 0.009932f
C5622 vdd.n2916 gnd 0.009932f
C5623 vdd.n2917 gnd 0.007994f
C5624 vdd.n2918 gnd 0.007994f
C5625 vdd.n2919 gnd 0.007994f
C5626 vdd.n2920 gnd 0.009932f
C5627 vdd.n2922 gnd 0.009932f
C5628 vdd.n2923 gnd 0.009932f
C5629 vdd.n2924 gnd 0.007994f
C5630 vdd.n2925 gnd 0.007994f
C5631 vdd.n2926 gnd 0.009932f
C5632 vdd.n2927 gnd 0.009932f
C5633 vdd.n2928 gnd 0.007994f
C5634 vdd.n2929 gnd 0.007994f
C5635 vdd.n2930 gnd 0.009932f
C5636 vdd.n2931 gnd 0.009932f
C5637 vdd.n2933 gnd 0.009932f
C5638 vdd.n2934 gnd 0.007994f
C5639 vdd.n2935 gnd 0.006635f
C5640 vdd.n2936 gnd 0.023771f
C5641 vdd.n2937 gnd 0.023405f
C5642 vdd.n2938 gnd 0.006635f
C5643 vdd.n2939 gnd 0.023405f
C5644 vdd.n2940 gnd 1.39559f
C5645 vdd.n2941 gnd 0.023405f
C5646 vdd.n2942 gnd 0.006635f
C5647 vdd.n2943 gnd 0.023405f
C5648 vdd.n2944 gnd 0.009932f
C5649 vdd.n2945 gnd 0.009932f
C5650 vdd.n2946 gnd 0.007994f
C5651 vdd.n2947 gnd 0.009932f
C5652 vdd.n2948 gnd 1.01498f
C5653 vdd.n2949 gnd 0.009932f
C5654 vdd.n2950 gnd 0.007994f
C5655 vdd.n2951 gnd 0.009932f
C5656 vdd.n2952 gnd 0.009932f
C5657 vdd.n2953 gnd 0.009932f
C5658 vdd.n2954 gnd 0.007994f
C5659 vdd.n2955 gnd 0.009932f
C5660 vdd.n2956 gnd 0.898254f
C5661 vdd.n2957 gnd 0.009932f
C5662 vdd.n2958 gnd 0.007994f
C5663 vdd.n2959 gnd 0.009932f
C5664 vdd.n2960 gnd 0.009932f
C5665 vdd.n2961 gnd 0.009932f
C5666 vdd.n2962 gnd 0.007994f
C5667 vdd.n2963 gnd 0.009932f
C5668 vdd.t181 gnd 0.507488f
C5669 vdd.n2964 gnd 0.725708f
C5670 vdd.n2965 gnd 0.009932f
C5671 vdd.n2966 gnd 0.007994f
C5672 vdd.n2967 gnd 0.009932f
C5673 vdd.n2968 gnd 0.009932f
C5674 vdd.n2969 gnd 0.009932f
C5675 vdd.n2970 gnd 0.007994f
C5676 vdd.n2971 gnd 0.009932f
C5677 vdd.n2972 gnd 0.553162f
C5678 vdd.n2973 gnd 0.009932f
C5679 vdd.n2974 gnd 0.007994f
C5680 vdd.n2975 gnd 0.009932f
C5681 vdd.n2976 gnd 0.009932f
C5682 vdd.n2977 gnd 0.009932f
C5683 vdd.n2978 gnd 0.007994f
C5684 vdd.n2979 gnd 0.009932f
C5685 vdd.n2980 gnd 0.715558f
C5686 vdd.n2981 gnd 0.63436f
C5687 vdd.n2982 gnd 0.009932f
C5688 vdd.n2983 gnd 0.007994f
C5689 vdd.n2984 gnd 0.009932f
C5690 vdd.n2985 gnd 0.009932f
C5691 vdd.n2986 gnd 0.009932f
C5692 vdd.n2987 gnd 0.007994f
C5693 vdd.n2988 gnd 0.009932f
C5694 vdd.n2989 gnd 0.806906f
C5695 vdd.n2990 gnd 0.009932f
C5696 vdd.n2991 gnd 0.007994f
C5697 vdd.n2992 gnd 0.009932f
C5698 vdd.n2993 gnd 0.009932f
C5699 vdd.n2994 gnd 0.009932f
C5700 vdd.n2995 gnd 0.007994f
C5701 vdd.n2996 gnd 0.007994f
C5702 vdd.n2997 gnd 0.007994f
C5703 vdd.n2998 gnd 0.009932f
C5704 vdd.n2999 gnd 0.009932f
C5705 vdd.n3000 gnd 0.009932f
C5706 vdd.n3001 gnd 0.007994f
C5707 vdd.n3002 gnd 0.007994f
C5708 vdd.n3003 gnd 0.007994f
C5709 vdd.n3004 gnd 0.009932f
C5710 vdd.n3005 gnd 0.009932f
C5711 vdd.n3006 gnd 0.009932f
C5712 vdd.n3007 gnd 0.007994f
C5713 vdd.n3008 gnd 0.007994f
C5714 vdd.n3009 gnd 0.007994f
C5715 vdd.n3010 gnd 0.009932f
C5716 vdd.n3011 gnd 0.009932f
C5717 vdd.n3012 gnd 0.009932f
C5718 vdd.n3013 gnd 0.007994f
C5719 vdd.n3014 gnd 0.007994f
C5720 vdd.n3015 gnd 0.006635f
C5721 vdd.n3016 gnd 0.023405f
C5722 vdd.n3017 gnd 0.023771f
C5723 vdd.n3019 gnd 0.023771f
C5724 vdd.n3020 gnd 0.003797f
C5725 vdd.t78 gnd 0.122186f
C5726 vdd.t77 gnd 0.130584f
C5727 vdd.t76 gnd 0.159574f
C5728 vdd.n3021 gnd 0.204551f
C5729 vdd.n3022 gnd 0.172659f
C5730 vdd.n3023 gnd 0.01311f
C5731 vdd.n3024 gnd 0.004197f
C5732 vdd.n3025 gnd 0.007994f
C5733 vdd.n3026 gnd 0.009932f
C5734 vdd.n3028 gnd 0.009932f
C5735 vdd.n3029 gnd 0.009932f
C5736 vdd.n3030 gnd 0.007994f
C5737 vdd.n3031 gnd 0.007994f
C5738 vdd.n3032 gnd 0.007994f
C5739 vdd.n3033 gnd 0.009932f
C5740 vdd.n3035 gnd 0.009932f
C5741 vdd.n3036 gnd 0.009932f
C5742 vdd.n3037 gnd 0.007994f
C5743 vdd.n3038 gnd 0.007994f
C5744 vdd.n3039 gnd 0.007994f
C5745 vdd.n3040 gnd 0.009932f
C5746 vdd.n3042 gnd 0.009932f
C5747 vdd.n3043 gnd 0.009932f
C5748 vdd.n3044 gnd 0.007994f
C5749 vdd.n3045 gnd 0.007994f
C5750 vdd.n3046 gnd 0.007994f
C5751 vdd.n3047 gnd 0.009932f
C5752 vdd.n3049 gnd 0.009932f
C5753 vdd.n3050 gnd 0.009932f
C5754 vdd.n3051 gnd 0.007994f
C5755 vdd.n3052 gnd 0.007994f
C5756 vdd.n3053 gnd 0.007994f
C5757 vdd.n3054 gnd 0.009932f
C5758 vdd.n3056 gnd 0.009932f
C5759 vdd.n3057 gnd 0.009932f
C5760 vdd.n3058 gnd 0.007994f
C5761 vdd.n3059 gnd 0.009932f
C5762 vdd.n3060 gnd 0.009932f
C5763 vdd.n3061 gnd 0.009932f
C5764 vdd.n3062 gnd 0.017107f
C5765 vdd.n3063 gnd 0.005436f
C5766 vdd.n3064 gnd 0.007994f
C5767 vdd.n3065 gnd 0.009932f
C5768 vdd.n3067 gnd 0.009932f
C5769 vdd.n3068 gnd 0.009932f
C5770 vdd.n3069 gnd 0.007994f
C5771 vdd.n3070 gnd 0.007994f
C5772 vdd.n3071 gnd 0.007994f
C5773 vdd.n3072 gnd 0.009932f
C5774 vdd.n3074 gnd 0.009932f
C5775 vdd.n3075 gnd 0.009932f
C5776 vdd.n3076 gnd 0.007994f
C5777 vdd.n3077 gnd 0.007994f
C5778 vdd.n3078 gnd 0.007994f
C5779 vdd.n3079 gnd 0.009932f
C5780 vdd.n3081 gnd 0.009932f
C5781 vdd.n3082 gnd 0.009932f
C5782 vdd.n3083 gnd 0.007994f
C5783 vdd.n3084 gnd 0.007994f
C5784 vdd.n3085 gnd 0.007994f
C5785 vdd.n3086 gnd 0.009932f
C5786 vdd.n3088 gnd 0.009932f
C5787 vdd.n3089 gnd 0.009932f
C5788 vdd.n3090 gnd 0.007994f
C5789 vdd.n3091 gnd 0.007994f
C5790 vdd.n3092 gnd 0.007994f
C5791 vdd.n3093 gnd 0.009932f
C5792 vdd.n3095 gnd 0.009932f
C5793 vdd.n3096 gnd 0.009932f
C5794 vdd.n3097 gnd 0.007994f
C5795 vdd.n3098 gnd 0.009932f
C5796 vdd.n3099 gnd 0.009932f
C5797 vdd.n3100 gnd 0.009932f
C5798 vdd.n3101 gnd 0.017107f
C5799 vdd.n3102 gnd 0.006675f
C5800 vdd.n3103 gnd 0.007994f
C5801 vdd.n3104 gnd 0.009932f
C5802 vdd.n3106 gnd 0.009932f
C5803 vdd.n3107 gnd 0.009932f
C5804 vdd.n3108 gnd 0.007994f
C5805 vdd.n3109 gnd 0.007994f
C5806 vdd.n3110 gnd 0.007994f
C5807 vdd.n3111 gnd 0.009932f
C5808 vdd.n3113 gnd 0.009932f
C5809 vdd.n3114 gnd 0.009932f
C5810 vdd.n3115 gnd 0.007994f
C5811 vdd.n3116 gnd 0.007994f
C5812 vdd.n3117 gnd 0.007994f
C5813 vdd.n3118 gnd 0.009932f
C5814 vdd.n3120 gnd 0.009932f
C5815 vdd.n3121 gnd 0.009932f
C5816 vdd.n3122 gnd 0.007994f
C5817 vdd.n3123 gnd 0.007994f
C5818 vdd.n3124 gnd 0.007994f
C5819 vdd.n3125 gnd 0.009932f
C5820 vdd.n3127 gnd 0.009932f
C5821 vdd.n3128 gnd 0.009932f
C5822 vdd.n3130 gnd 0.009932f
C5823 vdd.n3131 gnd 0.007994f
C5824 vdd.n3132 gnd 0.007994f
C5825 vdd.n3133 gnd 0.006635f
C5826 vdd.n3134 gnd 0.023771f
C5827 vdd.n3135 gnd 0.023405f
C5828 vdd.n3136 gnd 0.006635f
C5829 vdd.n3137 gnd 0.023405f
C5830 vdd.n3138 gnd 1.43112f
C5831 vdd.n3139 gnd 0.573462f
C5832 vdd.t12 gnd 0.507488f
C5833 vdd.n3140 gnd 0.949003f
C5834 vdd.n3141 gnd 0.009932f
C5835 vdd.n3142 gnd 0.007994f
C5836 vdd.n3143 gnd 0.007994f
C5837 vdd.n3144 gnd 0.007994f
C5838 vdd.n3145 gnd 0.009932f
C5839 vdd.n3146 gnd 0.999752f
C5840 vdd.t153 gnd 0.507488f
C5841 vdd.n3147 gnd 0.522713f
C5842 vdd.n3148 gnd 0.827206f
C5843 vdd.n3149 gnd 0.009932f
C5844 vdd.n3150 gnd 0.007994f
C5845 vdd.n3151 gnd 0.007994f
C5846 vdd.n3152 gnd 0.007994f
C5847 vdd.n3153 gnd 0.009932f
C5848 vdd.n3154 gnd 0.65466f
C5849 vdd.t148 gnd 0.507488f
C5850 vdd.n3155 gnd 0.84243f
C5851 vdd.t167 gnd 0.507488f
C5852 vdd.n3156 gnd 0.532863f
C5853 vdd.n3157 gnd 0.009932f
C5854 vdd.n3158 gnd 0.007994f
C5855 vdd.n3159 gnd 0.007994f
C5856 vdd.n3160 gnd 0.007994f
C5857 vdd.n3161 gnd 0.009932f
C5858 vdd.n3162 gnd 0.705409f
C5859 vdd.n3163 gnd 0.64451f
C5860 vdd.t132 gnd 0.507488f
C5861 vdd.n3164 gnd 0.84243f
C5862 vdd.n3165 gnd 0.009932f
C5863 vdd.n3166 gnd 0.007994f
C5864 vdd.n3167 gnd 0.591214f
C5865 vdd.n3168 gnd 2.18846f
C5866 a_n6308_8799.n0 gnd 3.87215f
C5867 a_n6308_8799.n1 gnd 1.93002f
C5868 a_n6308_8799.n2 gnd 3.25964f
C5869 a_n6308_8799.n3 gnd 0.793828f
C5870 a_n6308_8799.n4 gnd 0.178521f
C5871 a_n6308_8799.n5 gnd 0.20906f
C5872 a_n6308_8799.n6 gnd 0.20906f
C5873 a_n6308_8799.n7 gnd 0.20906f
C5874 a_n6308_8799.n8 gnd 0.178521f
C5875 a_n6308_8799.n9 gnd 0.20906f
C5876 a_n6308_8799.n10 gnd 0.20906f
C5877 a_n6308_8799.n11 gnd 0.20906f
C5878 a_n6308_8799.n12 gnd 0.344841f
C5879 a_n6308_8799.n13 gnd 0.20906f
C5880 a_n6308_8799.n14 gnd 0.20906f
C5881 a_n6308_8799.n15 gnd 0.20906f
C5882 a_n6308_8799.n16 gnd 0.20906f
C5883 a_n6308_8799.n17 gnd 0.20906f
C5884 a_n6308_8799.n18 gnd 0.178521f
C5885 a_n6308_8799.n19 gnd 0.20906f
C5886 a_n6308_8799.n20 gnd 0.20906f
C5887 a_n6308_8799.n21 gnd 0.20906f
C5888 a_n6308_8799.n22 gnd 0.178521f
C5889 a_n6308_8799.n23 gnd 0.20906f
C5890 a_n6308_8799.n24 gnd 0.20906f
C5891 a_n6308_8799.n25 gnd 0.20906f
C5892 a_n6308_8799.n26 gnd 0.344841f
C5893 a_n6308_8799.n27 gnd 0.20906f
C5894 a_n6308_8799.n28 gnd 2.82984f
C5895 a_n6308_8799.n29 gnd 4.02299f
C5896 a_n6308_8799.n30 gnd 0.252822f
C5897 a_n6308_8799.n32 gnd 0.007787f
C5898 a_n6308_8799.n33 gnd 0.011769f
C5899 a_n6308_8799.n34 gnd 0.008094f
C5900 a_n6308_8799.n36 gnd 4.04e-19
C5901 a_n6308_8799.n37 gnd 0.008389f
C5902 a_n6308_8799.n38 gnd 0.264482f
C5903 a_n6308_8799.n39 gnd 0.252822f
C5904 a_n6308_8799.n41 gnd 0.007787f
C5905 a_n6308_8799.n42 gnd 0.011769f
C5906 a_n6308_8799.n43 gnd 0.008094f
C5907 a_n6308_8799.n45 gnd 4.04e-19
C5908 a_n6308_8799.n46 gnd 0.008389f
C5909 a_n6308_8799.n47 gnd 0.264482f
C5910 a_n6308_8799.n48 gnd 0.252822f
C5911 a_n6308_8799.n50 gnd 0.007787f
C5912 a_n6308_8799.n51 gnd 0.011769f
C5913 a_n6308_8799.n52 gnd 0.008094f
C5914 a_n6308_8799.n54 gnd 4.04e-19
C5915 a_n6308_8799.n55 gnd 0.008389f
C5916 a_n6308_8799.n56 gnd 0.264482f
C5917 a_n6308_8799.n57 gnd 0.008389f
C5918 a_n6308_8799.n58 gnd 0.264482f
C5919 a_n6308_8799.n59 gnd 4.04e-19
C5920 a_n6308_8799.n61 gnd 0.008094f
C5921 a_n6308_8799.n62 gnd 0.011769f
C5922 a_n6308_8799.n63 gnd 0.007787f
C5923 a_n6308_8799.n65 gnd 0.252822f
C5924 a_n6308_8799.n66 gnd 0.008389f
C5925 a_n6308_8799.n67 gnd 0.264482f
C5926 a_n6308_8799.n68 gnd 4.04e-19
C5927 a_n6308_8799.n70 gnd 0.008094f
C5928 a_n6308_8799.n71 gnd 0.011769f
C5929 a_n6308_8799.n72 gnd 0.007787f
C5930 a_n6308_8799.n74 gnd 0.252822f
C5931 a_n6308_8799.n75 gnd 0.008389f
C5932 a_n6308_8799.n76 gnd 0.264482f
C5933 a_n6308_8799.n77 gnd 4.04e-19
C5934 a_n6308_8799.n79 gnd 0.008094f
C5935 a_n6308_8799.n80 gnd 0.011769f
C5936 a_n6308_8799.n81 gnd 0.007787f
C5937 a_n6308_8799.n83 gnd 0.252822f
C5938 a_n6308_8799.t22 gnd 0.145006f
C5939 a_n6308_8799.t8 gnd 0.145006f
C5940 a_n6308_8799.t23 gnd 0.145006f
C5941 a_n6308_8799.n84 gnd 1.14369f
C5942 a_n6308_8799.t6 gnd 0.145006f
C5943 a_n6308_8799.t28 gnd 0.145006f
C5944 a_n6308_8799.n85 gnd 1.1418f
C5945 a_n6308_8799.t5 gnd 0.145006f
C5946 a_n6308_8799.t29 gnd 0.145006f
C5947 a_n6308_8799.n86 gnd 1.1418f
C5948 a_n6308_8799.t25 gnd 0.112783f
C5949 a_n6308_8799.t2 gnd 0.112783f
C5950 a_n6308_8799.n87 gnd 0.998803f
C5951 a_n6308_8799.t17 gnd 0.112783f
C5952 a_n6308_8799.t34 gnd 0.112783f
C5953 a_n6308_8799.n88 gnd 0.996586f
C5954 a_n6308_8799.t30 gnd 0.112783f
C5955 a_n6308_8799.t11 gnd 0.112783f
C5956 a_n6308_8799.n89 gnd 0.996586f
C5957 a_n6308_8799.t18 gnd 0.112783f
C5958 a_n6308_8799.t1 gnd 0.112783f
C5959 a_n6308_8799.n90 gnd 0.998802f
C5960 a_n6308_8799.t10 gnd 0.112783f
C5961 a_n6308_8799.t9 gnd 0.112783f
C5962 a_n6308_8799.n91 gnd 0.996586f
C5963 a_n6308_8799.t15 gnd 0.112783f
C5964 a_n6308_8799.t21 gnd 0.112783f
C5965 a_n6308_8799.n92 gnd 0.996586f
C5966 a_n6308_8799.t32 gnd 0.112783f
C5967 a_n6308_8799.t19 gnd 0.112783f
C5968 a_n6308_8799.n93 gnd 0.998802f
C5969 a_n6308_8799.t3 gnd 0.112783f
C5970 a_n6308_8799.t33 gnd 0.112783f
C5971 a_n6308_8799.n94 gnd 0.996586f
C5972 a_n6308_8799.t24 gnd 0.112783f
C5973 a_n6308_8799.t35 gnd 0.112783f
C5974 a_n6308_8799.n95 gnd 0.996586f
C5975 a_n6308_8799.t20 gnd 0.112783f
C5976 a_n6308_8799.t31 gnd 0.112783f
C5977 a_n6308_8799.n96 gnd 0.996586f
C5978 a_n6308_8799.t0 gnd 0.112783f
C5979 a_n6308_8799.t7 gnd 0.112783f
C5980 a_n6308_8799.n97 gnd 0.996586f
C5981 a_n6308_8799.t16 gnd 0.112783f
C5982 a_n6308_8799.t26 gnd 0.112783f
C5983 a_n6308_8799.n98 gnd 0.996586f
C5984 a_n6308_8799.t94 gnd 0.601263f
C5985 a_n6308_8799.n99 gnd 0.272125f
C5986 a_n6308_8799.t41 gnd 0.601263f
C5987 a_n6308_8799.t44 gnd 0.601263f
C5988 a_n6308_8799.n100 gnd 0.263219f
C5989 a_n6308_8799.t57 gnd 0.601263f
C5990 a_n6308_8799.n101 gnd 0.274674f
C5991 a_n6308_8799.t71 gnd 0.601263f
C5992 a_n6308_8799.t84 gnd 0.601263f
C5993 a_n6308_8799.n102 gnd 0.268052f
C5994 a_n6308_8799.t59 gnd 0.615394f
C5995 a_n6308_8799.t60 gnd 0.601263f
C5996 a_n6308_8799.n103 gnd 0.274236f
C5997 a_n6308_8799.n104 gnd 0.250639f
C5998 a_n6308_8799.t36 gnd 0.601263f
C5999 a_n6308_8799.n105 gnd 0.272007f
C6000 a_n6308_8799.n106 gnd 0.27214f
C6001 a_n6308_8799.t96 gnd 0.601263f
C6002 a_n6308_8799.n107 gnd 0.268374f
C6003 a_n6308_8799.t55 gnd 0.601263f
C6004 a_n6308_8799.n108 gnd 0.268626f
C6005 a_n6308_8799.n109 gnd 0.274237f
C6006 a_n6308_8799.t42 gnd 0.612179f
C6007 a_n6308_8799.t100 gnd 0.601263f
C6008 a_n6308_8799.n110 gnd 0.272125f
C6009 a_n6308_8799.t48 gnd 0.601263f
C6010 a_n6308_8799.t53 gnd 0.601263f
C6011 a_n6308_8799.n111 gnd 0.263219f
C6012 a_n6308_8799.t64 gnd 0.601263f
C6013 a_n6308_8799.n112 gnd 0.274674f
C6014 a_n6308_8799.t78 gnd 0.601263f
C6015 a_n6308_8799.t91 gnd 0.601263f
C6016 a_n6308_8799.n113 gnd 0.268052f
C6017 a_n6308_8799.t65 gnd 0.615394f
C6018 a_n6308_8799.t66 gnd 0.601263f
C6019 a_n6308_8799.n114 gnd 0.274236f
C6020 a_n6308_8799.n115 gnd 0.250639f
C6021 a_n6308_8799.t43 gnd 0.601263f
C6022 a_n6308_8799.n116 gnd 0.272007f
C6023 a_n6308_8799.n117 gnd 0.27214f
C6024 a_n6308_8799.t104 gnd 0.601263f
C6025 a_n6308_8799.n118 gnd 0.268374f
C6026 a_n6308_8799.t63 gnd 0.601263f
C6027 a_n6308_8799.n119 gnd 0.268626f
C6028 a_n6308_8799.n120 gnd 0.274237f
C6029 a_n6308_8799.t50 gnd 0.612179f
C6030 a_n6308_8799.n121 gnd 0.902661f
C6031 a_n6308_8799.t74 gnd 0.601263f
C6032 a_n6308_8799.n122 gnd 0.272125f
C6033 a_n6308_8799.t46 gnd 0.601263f
C6034 a_n6308_8799.t92 gnd 0.601263f
C6035 a_n6308_8799.n123 gnd 0.263219f
C6036 a_n6308_8799.t39 gnd 0.601263f
C6037 a_n6308_8799.n124 gnd 0.274674f
C6038 a_n6308_8799.t80 gnd 0.601263f
C6039 a_n6308_8799.t101 gnd 0.601263f
C6040 a_n6308_8799.n125 gnd 0.268052f
C6041 a_n6308_8799.t98 gnd 0.615394f
C6042 a_n6308_8799.t85 gnd 0.601263f
C6043 a_n6308_8799.n126 gnd 0.274236f
C6044 a_n6308_8799.n127 gnd 0.250639f
C6045 a_n6308_8799.t70 gnd 0.601263f
C6046 a_n6308_8799.n128 gnd 0.272007f
C6047 a_n6308_8799.n129 gnd 0.27214f
C6048 a_n6308_8799.t51 gnd 0.601263f
C6049 a_n6308_8799.n130 gnd 0.268374f
C6050 a_n6308_8799.t58 gnd 0.601263f
C6051 a_n6308_8799.n131 gnd 0.268626f
C6052 a_n6308_8799.n132 gnd 0.274237f
C6053 a_n6308_8799.t105 gnd 0.612179f
C6054 a_n6308_8799.n133 gnd 1.50375f
C6055 a_n6308_8799.t68 gnd 0.612179f
C6056 a_n6308_8799.t67 gnd 0.601263f
C6057 a_n6308_8799.t49 gnd 0.601263f
C6058 a_n6308_8799.t95 gnd 0.601263f
C6059 a_n6308_8799.n134 gnd 0.268626f
C6060 a_n6308_8799.t69 gnd 0.601263f
C6061 a_n6308_8799.t54 gnd 0.601263f
C6062 a_n6308_8799.t97 gnd 0.601263f
C6063 a_n6308_8799.n135 gnd 0.27214f
C6064 a_n6308_8799.t79 gnd 0.601263f
C6065 a_n6308_8799.t77 gnd 0.601263f
C6066 a_n6308_8799.t38 gnd 0.601263f
C6067 a_n6308_8799.n136 gnd 0.268052f
C6068 a_n6308_8799.t82 gnd 0.615394f
C6069 a_n6308_8799.t83 gnd 0.601263f
C6070 a_n6308_8799.n137 gnd 0.274236f
C6071 a_n6308_8799.n138 gnd 0.250639f
C6072 a_n6308_8799.n139 gnd 0.272007f
C6073 a_n6308_8799.n140 gnd 0.274674f
C6074 a_n6308_8799.n141 gnd 0.268374f
C6075 a_n6308_8799.n142 gnd 0.263219f
C6076 a_n6308_8799.n143 gnd 0.272125f
C6077 a_n6308_8799.n144 gnd 0.274237f
C6078 a_n6308_8799.t73 gnd 0.612179f
C6079 a_n6308_8799.t72 gnd 0.601263f
C6080 a_n6308_8799.t61 gnd 0.601263f
C6081 a_n6308_8799.t103 gnd 0.601263f
C6082 a_n6308_8799.n145 gnd 0.268626f
C6083 a_n6308_8799.t76 gnd 0.601263f
C6084 a_n6308_8799.t62 gnd 0.601263f
C6085 a_n6308_8799.t107 gnd 0.601263f
C6086 a_n6308_8799.n146 gnd 0.27214f
C6087 a_n6308_8799.t88 gnd 0.601263f
C6088 a_n6308_8799.t87 gnd 0.601263f
C6089 a_n6308_8799.t45 gnd 0.601263f
C6090 a_n6308_8799.n147 gnd 0.268052f
C6091 a_n6308_8799.t89 gnd 0.615394f
C6092 a_n6308_8799.t90 gnd 0.601263f
C6093 a_n6308_8799.n148 gnd 0.274236f
C6094 a_n6308_8799.n149 gnd 0.250639f
C6095 a_n6308_8799.n150 gnd 0.272007f
C6096 a_n6308_8799.n151 gnd 0.274674f
C6097 a_n6308_8799.n152 gnd 0.268374f
C6098 a_n6308_8799.n153 gnd 0.263219f
C6099 a_n6308_8799.n154 gnd 0.272125f
C6100 a_n6308_8799.n155 gnd 0.274237f
C6101 a_n6308_8799.n156 gnd 0.902661f
C6102 a_n6308_8799.t106 gnd 0.612179f
C6103 a_n6308_8799.t47 gnd 0.601263f
C6104 a_n6308_8799.t75 gnd 0.601263f
C6105 a_n6308_8799.t37 gnd 0.601263f
C6106 a_n6308_8799.n157 gnd 0.268626f
C6107 a_n6308_8799.t93 gnd 0.601263f
C6108 a_n6308_8799.t52 gnd 0.601263f
C6109 a_n6308_8799.t81 gnd 0.601263f
C6110 a_n6308_8799.n158 gnd 0.27214f
C6111 a_n6308_8799.t40 gnd 0.601263f
C6112 a_n6308_8799.t56 gnd 0.601263f
C6113 a_n6308_8799.t102 gnd 0.601263f
C6114 a_n6308_8799.n159 gnd 0.268052f
C6115 a_n6308_8799.t99 gnd 0.615394f
C6116 a_n6308_8799.t86 gnd 0.601263f
C6117 a_n6308_8799.n160 gnd 0.274236f
C6118 a_n6308_8799.n161 gnd 0.250639f
C6119 a_n6308_8799.n162 gnd 0.272007f
C6120 a_n6308_8799.n163 gnd 0.274674f
C6121 a_n6308_8799.n164 gnd 0.268374f
C6122 a_n6308_8799.n165 gnd 0.263219f
C6123 a_n6308_8799.n166 gnd 0.272125f
C6124 a_n6308_8799.n167 gnd 0.274237f
C6125 a_n6308_8799.n168 gnd 1.11639f
C6126 a_n6308_8799.n169 gnd 12.2999f
C6127 a_n6308_8799.n170 gnd 4.40037f
C6128 a_n6308_8799.n171 gnd 5.7182f
C6129 a_n6308_8799.t13 gnd 0.145006f
C6130 a_n6308_8799.t14 gnd 0.145006f
C6131 a_n6308_8799.n172 gnd 1.1418f
C6132 a_n6308_8799.t12 gnd 0.145006f
C6133 a_n6308_8799.t27 gnd 0.145006f
C6134 a_n6308_8799.n173 gnd 1.14368f
C6135 a_n6308_8799.n174 gnd 1.1418f
C6136 a_n6308_8799.t4 gnd 0.145006f
.ends

