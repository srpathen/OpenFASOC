* NGSPICE file created from opamp0.ext - technology: sky130A

.subckt opamp0 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 gnd.t315 commonsourceibias.t18 commonsourceibias.t19 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t119 a_n7636_8799.t28 vdd.t173 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n1808_13878.t19 a_n1986_13878.t40 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n1808_13878.t11 a_n1986_13878.t20 a_n1986_13878.t21 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t172 a_n7636_8799.t29 CSoutput.t118 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 CSoutput.t117 a_n7636_8799.t30 vdd.t171 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 commonsourceibias.t17 commonsourceibias.t16 gnd.t314 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 a_n3827_n3924.t38 diffpairibias.t20 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X8 CSoutput.t116 a_n7636_8799.t31 vdd.t170 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X9 gnd.t313 commonsourceibias.t14 commonsourceibias.t15 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 vdd.t286 vdd.t284 vdd.t285 vdd.t238 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X11 a_n1986_8322.t13 a_n1986_13878.t41 a_n7636_8799.t0 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X12 commonsourceibias.t13 commonsourceibias.t12 gnd.t312 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t311 commonsourceibias.t48 CSoutput.t191 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 CSoutput.t115 a_n7636_8799.t32 vdd.t169 vdd.t71 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 a_n7636_8799.t23 plus.t5 a_n3827_n3924.t27 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X16 vdd.t160 a_n7636_8799.t33 CSoutput.t114 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 gnd.t120 gnd.t118 gnd.t119 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X18 output.t3 outputibias.t8 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X19 vdd.t168 a_n7636_8799.t34 CSoutput.t113 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 CSoutput.t112 a_n7636_8799.t35 vdd.t167 vdd.t73 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 vdd.t166 a_n7636_8799.t36 CSoutput.t111 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 commonsourceibias.t11 commonsourceibias.t10 gnd.t310 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t165 a_n7636_8799.t37 CSoutput.t110 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 a_n7636_8799.t4 a_n1986_13878.t42 a_n1986_8322.t12 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X25 gnd.t117 gnd.t114 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X26 gnd.t113 gnd.t110 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X27 CSoutput.t109 a_n7636_8799.t38 vdd.t164 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X28 a_n7636_8799.t18 plus.t6 a_n3827_n3924.t22 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X29 gnd.t309 commonsourceibias.t49 CSoutput.t190 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X30 CSoutput.t189 commonsourceibias.t50 gnd.t308 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X31 gnd.t307 commonsourceibias.t34 commonsourceibias.t35 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 CSoutput.t108 a_n7636_8799.t39 vdd.t163 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 vdd.t283 vdd.t281 vdd.t282 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X34 a_n3827_n3924.t37 diffpairibias.t21 gnd.t317 gnd.t316 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X35 a_n3827_n3924.t39 minus.t5 a_n1986_13878.t38 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X36 CSoutput.t107 a_n7636_8799.t40 vdd.t159 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 commonsourceibias.t33 commonsourceibias.t32 gnd.t306 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X38 gnd.t109 gnd.t107 plus.t4 gnd.t108 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X39 a_n3827_n3924.t16 plus.t7 a_n7636_8799.t12 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X40 a_n1986_13878.t39 minus.t6 a_n3827_n3924.t40 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X41 a_n3827_n3924.t5 minus.t7 a_n1986_13878.t5 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X42 CSoutput.t106 a_n7636_8799.t41 vdd.t162 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 gnd.t305 commonsourceibias.t30 commonsourceibias.t31 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 CSoutput.t188 commonsourceibias.t51 gnd.t304 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X45 vdd.t161 a_n7636_8799.t42 CSoutput.t105 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 vdd.t280 vdd.t278 vdd.t279 vdd.t238 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X47 a_n1808_13878.t10 a_n1986_13878.t28 a_n1986_13878.t29 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X48 CSoutput.t104 a_n7636_8799.t43 vdd.t158 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 a_n1986_13878.t33 a_n1986_13878.t32 a_n1808_13878.t9 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X50 output.t2 outputibias.t9 gnd.t182 gnd.t181 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X51 CSoutput.t103 a_n7636_8799.t44 vdd.t157 vdd.t71 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 a_n3827_n3924.t4 minus.t8 a_n1986_13878.t4 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X53 vdd.t277 vdd.t275 vdd.t276 vdd.t251 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X54 vdd.t156 a_n7636_8799.t45 CSoutput.t102 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 diffpairibias.t19 diffpairibias.t18 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X56 CSoutput.t187 commonsourceibias.t52 gnd.t303 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 CSoutput.t186 commonsourceibias.t53 gnd.t302 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 CSoutput.t101 a_n7636_8799.t46 vdd.t155 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X59 gnd.t106 gnd.t104 gnd.t105 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X60 gnd.t103 gnd.t101 plus.t3 gnd.t102 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X61 vdd.t154 a_n7636_8799.t47 CSoutput.t100 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X62 vdd.t153 a_n7636_8799.t48 CSoutput.t99 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 minus.t4 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X64 vdd.t152 a_n7636_8799.t49 CSoutput.t98 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X65 vdd.t150 a_n7636_8799.t50 CSoutput.t97 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 diffpairibias.t17 diffpairibias.t16 gnd.t174 gnd.t173 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X67 CSoutput.t96 a_n7636_8799.t51 vdd.t149 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X68 CSoutput.t95 a_n7636_8799.t52 vdd.t148 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 gnd.t97 gnd.t95 gnd.t96 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X70 CSoutput.t192 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X71 vdd.t147 a_n7636_8799.t53 CSoutput.t94 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 CSoutput.t185 commonsourceibias.t54 gnd.t301 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 CSoutput.t93 a_n7636_8799.t54 vdd.t146 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t92 a_n7636_8799.t55 vdd.t145 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 CSoutput.t91 a_n7636_8799.t56 vdd.t144 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X76 CSoutput.t90 a_n7636_8799.t57 vdd.t143 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 output.t19 CSoutput.t193 vdd.t291 gnd.t318 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X78 vdd.t142 a_n7636_8799.t58 CSoutput.t89 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 gnd.t300 commonsourceibias.t55 CSoutput.t184 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t194 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X81 CSoutput.t183 commonsourceibias.t56 gnd.t299 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 a_n7636_8799.t27 plus.t8 a_n3827_n3924.t41 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X83 gnd.t298 commonsourceibias.t57 CSoutput.t182 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X84 gnd.t94 gnd.t92 gnd.t93 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X85 a_n3827_n3924.t36 diffpairibias.t22 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X86 vdd.t141 a_n7636_8799.t59 CSoutput.t88 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 a_n3827_n3924.t19 minus.t9 a_n1986_13878.t35 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X88 CSoutput.t181 commonsourceibias.t58 gnd.t297 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 a_n1986_13878.t11 a_n1986_13878.t10 a_n1808_13878.t8 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X90 vdd.t140 a_n7636_8799.t60 CSoutput.t87 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X91 a_n7636_8799.t1 a_n1986_13878.t43 a_n1986_8322.t11 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X92 vdd.t139 a_n7636_8799.t61 CSoutput.t86 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X93 a_n1986_13878.t19 a_n1986_13878.t18 a_n1808_13878.t7 vdd.t179 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X94 a_n1986_13878.t1 minus.t10 a_n3827_n3924.t1 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X95 vdd.t138 a_n7636_8799.t62 CSoutput.t85 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 a_n3827_n3924.t23 plus.t9 a_n7636_8799.t20 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X97 outputibias.t7 outputibias.t6 gnd.t167 gnd.t166 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X98 commonsourceibias.t29 commonsourceibias.t28 gnd.t296 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X99 gnd.t295 commonsourceibias.t59 CSoutput.t180 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 CSoutput.t179 commonsourceibias.t60 gnd.t294 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 vdd.t137 a_n7636_8799.t63 CSoutput.t84 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 CSoutput.t83 a_n7636_8799.t64 vdd.t115 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 gnd.t73 gnd.t71 gnd.t72 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X104 outputibias.t5 outputibias.t4 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X105 diffpairibias.t15 diffpairibias.t14 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X106 a_n3827_n3924.t3 minus.t11 a_n1986_13878.t3 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X107 vdd.t274 vdd.t272 vdd.t273 vdd.t259 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X108 vdd.t136 a_n7636_8799.t65 CSoutput.t82 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 CSoutput.t81 a_n7636_8799.t66 vdd.t135 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X110 vdd.t271 vdd.t268 vdd.t270 vdd.t269 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X111 vdd.t267 vdd.t265 vdd.t266 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X112 vdd.t264 vdd.t262 vdd.t263 vdd.t255 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X113 vdd.t293 a_n1986_13878.t44 a_n1986_8322.t21 vdd.t292 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X114 gnd.t293 commonsourceibias.t42 commonsourceibias.t43 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X115 output.t18 CSoutput.t195 vdd.t174 gnd.t131 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X116 CSoutput.t178 commonsourceibias.t61 gnd.t292 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 a_n1986_8322.t20 a_n1986_13878.t45 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X118 a_n3827_n3924.t35 diffpairibias.t23 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X119 CSoutput.t80 a_n7636_8799.t67 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X120 CSoutput.t79 a_n7636_8799.t68 vdd.t134 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X121 gnd.t291 commonsourceibias.t62 CSoutput.t177 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 a_n1986_13878.t6 minus.t12 a_n3827_n3924.t6 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X123 vdd.t131 a_n7636_8799.t69 CSoutput.t78 vdd.t130 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 commonsourceibias.t41 commonsourceibias.t40 gnd.t290 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X125 a_n3827_n3924.t28 plus.t10 a_n7636_8799.t24 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X126 vdd.t13 a_n1986_13878.t46 a_n1808_13878.t18 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X127 gnd.t289 commonsourceibias.t63 CSoutput.t176 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 gnd.t91 gnd.t89 gnd.t90 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X129 gnd.t85 gnd.t83 gnd.t84 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X130 gnd.t288 commonsourceibias.t38 commonsourceibias.t39 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 vdd.t261 vdd.t258 vdd.t260 vdd.t259 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X132 vdd.t129 a_n7636_8799.t70 CSoutput.t77 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 vdd.t257 vdd.t254 vdd.t256 vdd.t255 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X134 CSoutput.t175 commonsourceibias.t64 gnd.t287 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 a_n7636_8799.t9 plus.t11 a_n3827_n3924.t13 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X136 commonsourceibias.t37 commonsourceibias.t36 gnd.t286 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 vdd.t253 vdd.t250 vdd.t252 vdd.t251 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X138 a_n1986_8322.t19 a_n1986_13878.t47 vdd.t288 vdd.t287 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X139 gnd.t285 commonsourceibias.t65 CSoutput.t174 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X140 a_n7636_8799.t25 a_n1986_13878.t48 a_n1986_8322.t10 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X141 CSoutput.t76 a_n7636_8799.t71 vdd.t127 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 diffpairibias.t13 diffpairibias.t12 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X143 vdd.t126 a_n7636_8799.t72 CSoutput.t75 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X144 a_n1986_13878.t27 a_n1986_13878.t26 a_n1808_13878.t6 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 vdd.t124 a_n7636_8799.t73 CSoutput.t74 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X146 a_n7636_8799.t5 a_n1986_13878.t49 a_n1986_8322.t9 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 CSoutput.t73 a_n7636_8799.t74 vdd.t123 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 a_n1808_13878.t5 a_n1986_13878.t16 a_n1986_13878.t17 vdd.t11 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 plus.t2 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X150 gnd.t284 commonsourceibias.t66 CSoutput.t173 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 output.t17 CSoutput.t196 vdd.t175 gnd.t132 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X152 vdd.t8 CSoutput.t197 output.t16 gnd.t121 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X153 gnd.t283 commonsourceibias.t67 CSoutput.t172 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 gnd.t82 gnd.t80 minus.t3 gnd.t81 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X155 CSoutput.t72 a_n7636_8799.t75 vdd.t122 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 a_n1986_13878.t37 minus.t13 a_n3827_n3924.t26 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X157 vdd.t290 a_n1986_13878.t50 a_n1986_8322.t18 vdd.t289 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X158 vdd.t120 a_n7636_8799.t76 CSoutput.t71 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 gnd.t79 gnd.t77 gnd.t78 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X160 vdd.t9 CSoutput.t198 output.t15 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X161 CSoutput.t70 a_n7636_8799.t77 vdd.t121 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X162 CSoutput.t171 commonsourceibias.t68 gnd.t282 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 vdd.t119 a_n7636_8799.t78 CSoutput.t69 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X164 gnd.t281 commonsourceibias.t69 CSoutput.t170 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X165 gnd.t280 commonsourceibias.t70 CSoutput.t169 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 vdd.t118 a_n7636_8799.t79 CSoutput.t68 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X167 a_n3827_n3924.t34 diffpairibias.t24 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X168 a_n3827_n3924.t33 diffpairibias.t25 gnd.t184 gnd.t183 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X169 a_n1986_13878.t2 minus.t14 a_n3827_n3924.t2 gnd.t128 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X170 vdd.t117 a_n7636_8799.t80 CSoutput.t67 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X171 vdd.t116 a_n7636_8799.t81 CSoutput.t66 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 gnd.t76 gnd.t74 gnd.t75 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X173 CSoutput.t65 a_n7636_8799.t82 vdd.t114 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 CSoutput.t64 a_n7636_8799.t83 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X175 vdd.t10 CSoutput.t199 output.t14 gnd.t123 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X176 a_n1986_13878.t36 minus.t15 a_n3827_n3924.t25 gnd.t163 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X177 CSoutput.t63 a_n7636_8799.t84 vdd.t111 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 CSoutput.t168 commonsourceibias.t71 gnd.t279 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X179 output.t13 CSoutput.t200 vdd.t180 gnd.t139 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X180 gnd.t70 gnd.t68 gnd.t69 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X181 gnd.t278 commonsourceibias.t72 CSoutput.t167 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 diffpairibias.t11 diffpairibias.t10 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X183 a_n1808_13878.t17 a_n1986_13878.t51 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X184 vdd.t194 a_n1986_13878.t52 a_n1808_13878.t16 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 vdd.t249 vdd.t247 vdd.t248 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X186 vdd.t246 vdd.t244 vdd.t245 vdd.t231 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X187 CSoutput.t62 a_n7636_8799.t85 vdd.t110 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 gnd.t277 commonsourceibias.t73 CSoutput.t166 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 a_n3827_n3924.t10 plus.t12 a_n7636_8799.t7 gnd.t146 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X190 CSoutput.t165 commonsourceibias.t74 gnd.t276 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X191 vdd.t108 a_n7636_8799.t86 CSoutput.t61 vdd.t107 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X192 output.t12 CSoutput.t201 vdd.t181 gnd.t140 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X193 vdd.t243 vdd.t241 vdd.t242 vdd.t231 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X194 gnd.t67 gnd.t65 gnd.t66 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X195 plus.t1 gnd.t62 gnd.t64 gnd.t63 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X196 diffpairibias.t9 diffpairibias.t8 gnd.t322 gnd.t321 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X197 a_n3827_n3924.t24 plus.t13 a_n7636_8799.t21 gnd.t135 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X198 gnd.t275 commonsourceibias.t75 CSoutput.t164 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 gnd.t12 gnd.t9 gnd.t11 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X200 gnd.t61 gnd.t59 minus.t2 gnd.t60 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X201 CSoutput.t202 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X202 CSoutput.t60 a_n7636_8799.t87 vdd.t106 vdd.t105 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 vdd.t104 a_n7636_8799.t88 CSoutput.t59 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X204 gnd.t58 gnd.t56 gnd.t57 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X205 vdd.t103 a_n7636_8799.t89 CSoutput.t58 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X206 commonsourceibias.t25 commonsourceibias.t24 gnd.t274 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 a_n1986_8322.t8 a_n1986_13878.t53 a_n7636_8799.t22 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X208 CSoutput.t57 a_n7636_8799.t90 vdd.t102 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 diffpairibias.t7 diffpairibias.t6 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X210 vdd.t101 a_n7636_8799.t91 CSoutput.t56 vdd.t100 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 CSoutput.t55 a_n7636_8799.t92 vdd.t99 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X212 vdd.t98 a_n7636_8799.t93 CSoutput.t54 vdd.t97 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 vdd.t197 a_n1986_13878.t54 a_n1986_8322.t17 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X214 vdd.t96 a_n7636_8799.t94 CSoutput.t53 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X215 vdd.t95 a_n7636_8799.t95 CSoutput.t52 vdd.t94 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X216 gnd.t55 gnd.t52 gnd.t54 gnd.t53 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X217 CSoutput.t163 commonsourceibias.t76 gnd.t273 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X218 CSoutput.t203 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X219 output.t1 outputibias.t10 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X220 gnd.t51 gnd.t49 gnd.t50 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X221 commonsourceibias.t23 commonsourceibias.t22 gnd.t272 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 gnd.t48 gnd.t45 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X223 a_n1808_13878.t15 a_n1986_13878.t55 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X224 vdd.t202 CSoutput.t204 output.t11 gnd.t175 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X225 CSoutput.t162 commonsourceibias.t77 gnd.t271 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X226 gnd.t269 commonsourceibias.t78 CSoutput.t161 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 output.t0 outputibias.t11 gnd.t134 gnd.t133 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X228 vdd.t93 a_n7636_8799.t96 CSoutput.t51 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X229 CSoutput.t50 a_n7636_8799.t97 vdd.t92 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 gnd.t270 commonsourceibias.t20 commonsourceibias.t21 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X231 CSoutput.t49 a_n7636_8799.t98 vdd.t91 vdd.t73 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 gnd.t268 commonsourceibias.t79 CSoutput.t160 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X233 CSoutput.t159 commonsourceibias.t80 gnd.t267 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X234 gnd.t44 gnd.t42 minus.t1 gnd.t43 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X235 CSoutput.t158 commonsourceibias.t81 gnd.t266 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 gnd.t41 gnd.t38 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X237 vdd.t240 vdd.t237 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X238 CSoutput.t157 commonsourceibias.t82 gnd.t265 gnd.t264 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 gnd.t263 commonsourceibias.t83 CSoutput.t156 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 vdd.t236 vdd.t234 vdd.t235 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X241 a_n3827_n3924.t32 diffpairibias.t26 gnd.t165 gnd.t164 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X242 commonsourceibias.t45 commonsourceibias.t44 gnd.t262 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X243 vdd.t233 vdd.t230 vdd.t232 vdd.t231 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X244 vdd.t207 a_n1986_13878.t56 a_n1986_8322.t16 vdd.t206 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X245 a_n1986_8322.t7 a_n1986_13878.t57 a_n7636_8799.t26 vdd.t198 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X246 CSoutput.t48 a_n7636_8799.t99 vdd.t90 vdd.t89 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X247 vdd.t88 a_n7636_8799.t100 CSoutput.t47 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t155 commonsourceibias.t84 gnd.t259 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X249 CSoutput.t46 a_n7636_8799.t101 vdd.t87 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 gnd.t261 commonsourceibias.t85 CSoutput.t154 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X251 vdd.t86 a_n7636_8799.t102 CSoutput.t45 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 vdd.t85 a_n7636_8799.t103 CSoutput.t44 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 CSoutput.t153 commonsourceibias.t86 gnd.t260 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t258 commonsourceibias.t87 CSoutput.t152 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 gnd.t257 commonsourceibias.t88 CSoutput.t151 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X256 CSoutput.t150 commonsourceibias.t89 gnd.t256 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 gnd.t37 gnd.t34 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X258 a_n3827_n3924.t17 plus.t14 a_n7636_8799.t13 gnd.t157 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X259 vdd.t229 vdd.t226 vdd.t228 vdd.t227 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X260 vdd.t84 a_n7636_8799.t104 CSoutput.t43 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X261 a_n7636_8799.t8 plus.t15 a_n3827_n3924.t12 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X262 CSoutput.t42 a_n7636_8799.t105 vdd.t83 vdd.t82 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X263 a_n3827_n3924.t8 minus.t16 a_n1986_13878.t8 gnd.t144 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X264 a_n1808_13878.t4 a_n1986_13878.t22 a_n1986_13878.t23 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X265 CSoutput.t41 a_n7636_8799.t106 vdd.t81 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X266 CSoutput.t149 commonsourceibias.t90 gnd.t255 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 a_n1986_8322.t6 a_n1986_13878.t58 a_n7636_8799.t15 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X268 gnd.t254 commonsourceibias.t91 CSoutput.t148 gnd.t253 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 diffpairibias.t5 diffpairibias.t4 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X270 CSoutput.t147 commonsourceibias.t92 gnd.t252 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 a_n3827_n3924.t7 minus.t17 a_n1986_13878.t7 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X272 a_n7636_8799.t6 plus.t16 a_n3827_n3924.t9 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X273 output.t10 CSoutput.t205 vdd.t203 gnd.t176 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X274 CSoutput.t40 a_n7636_8799.t107 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 gnd.t250 commonsourceibias.t93 CSoutput.t146 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 CSoutput.t39 a_n7636_8799.t108 vdd.t78 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 a_n3827_n3924.t31 diffpairibias.t27 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X278 vdd.t77 a_n7636_8799.t109 CSoutput.t38 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 gnd.t201 commonsourceibias.t94 CSoutput.t145 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 vdd.t76 a_n7636_8799.t110 CSoutput.t37 vdd.t75 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X281 a_n1986_8322.t15 a_n1986_13878.t59 vdd.t7 vdd.t6 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X282 gnd.t249 commonsourceibias.t95 CSoutput.t144 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X283 CSoutput.t143 commonsourceibias.t96 gnd.t248 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X284 CSoutput.t36 a_n7636_8799.t111 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 outputibias.t3 outputibias.t2 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X286 gnd.t247 commonsourceibias.t26 commonsourceibias.t27 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 a_n3827_n3924.t18 plus.t17 a_n7636_8799.t14 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X288 vdd.t191 a_n1986_13878.t60 a_n1808_13878.t14 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X289 CSoutput.t35 a_n7636_8799.t112 vdd.t72 vdd.t71 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 gnd.t246 commonsourceibias.t97 CSoutput.t142 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X291 CSoutput.t141 commonsourceibias.t98 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X292 CSoutput.t34 a_n7636_8799.t113 vdd.t70 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 CSoutput.t140 commonsourceibias.t99 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 gnd.t242 commonsourceibias.t100 CSoutput.t139 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 commonsourceibias.t9 commonsourceibias.t8 gnd.t241 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X296 gnd.t239 commonsourceibias.t101 CSoutput.t138 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X297 vdd.t69 a_n7636_8799.t114 CSoutput.t33 vdd.t68 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 vdd.t67 a_n7636_8799.t115 CSoutput.t32 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 vdd.t225 vdd.t222 vdd.t224 vdd.t223 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X300 gnd.t238 commonsourceibias.t6 commonsourceibias.t7 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 a_n3827_n3924.t14 minus.t18 a_n1986_13878.t34 gnd.t150 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X302 a_n1986_8322.t5 a_n1986_13878.t61 a_n7636_8799.t19 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X303 CSoutput.t31 a_n7636_8799.t116 vdd.t66 vdd.t65 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X304 vdd.t221 vdd.t219 vdd.t220 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X305 a_n7636_8799.t10 a_n1986_13878.t62 a_n1986_8322.t4 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X306 gnd.t237 commonsourceibias.t102 CSoutput.t137 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 vdd.t59 a_n7636_8799.t117 CSoutput.t30 vdd.t58 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 a_n1808_13878.t13 a_n1986_13878.t63 vdd.t295 vdd.t294 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X309 CSoutput.t136 commonsourceibias.t103 gnd.t235 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X310 vdd.t64 a_n7636_8799.t118 CSoutput.t29 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X311 CSoutput.t28 a_n7636_8799.t119 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X312 vdd.t208 CSoutput.t206 output.t9 gnd.t185 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X313 gnd.t234 commonsourceibias.t4 commonsourceibias.t5 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 CSoutput.t135 commonsourceibias.t104 gnd.t233 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X315 a_n1986_13878.t9 minus.t19 a_n3827_n3924.t11 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X316 vdd.t61 a_n7636_8799.t120 CSoutput.t27 vdd.t60 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 CSoutput.t26 a_n7636_8799.t121 vdd.t57 vdd.t56 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 CSoutput.t25 a_n7636_8799.t122 vdd.t55 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X319 CSoutput.t134 commonsourceibias.t105 gnd.t232 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 gnd.t231 commonsourceibias.t106 CSoutput.t133 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 CSoutput.t24 a_n7636_8799.t123 vdd.t54 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 a_n1808_13878.t3 a_n1986_13878.t12 a_n1986_13878.t13 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X323 CSoutput.t23 a_n7636_8799.t124 vdd.t53 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 vdd.t52 a_n7636_8799.t125 CSoutput.t22 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 gnd.t230 commonsourceibias.t2 commonsourceibias.t3 gnd.t229 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X326 gnd.t228 commonsourceibias.t0 commonsourceibias.t1 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 CSoutput.t21 a_n7636_8799.t126 vdd.t51 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 a_n7636_8799.t17 plus.t18 a_n3827_n3924.t21 gnd.t162 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X329 a_n3827_n3924.t30 diffpairibias.t28 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X330 vdd.t50 a_n7636_8799.t127 CSoutput.t20 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X331 vdd.t49 a_n7636_8799.t128 CSoutput.t19 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X332 CSoutput.t132 commonsourceibias.t107 gnd.t226 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 gnd.t224 commonsourceibias.t108 CSoutput.t131 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 CSoutput.t18 a_n7636_8799.t129 vdd.t48 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 a_n1986_13878.t31 a_n1986_13878.t30 a_n1808_13878.t2 vdd.t4 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X336 output.t8 CSoutput.t207 vdd.t209 gnd.t186 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X337 a_n7636_8799.t2 a_n1986_13878.t64 a_n1986_8322.t3 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X338 vdd.t47 a_n7636_8799.t130 CSoutput.t17 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 CSoutput.t16 a_n7636_8799.t131 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 a_n3827_n3924.t15 plus.t19 a_n7636_8799.t11 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X341 gnd.t33 gnd.t30 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X342 vdd.t16 a_n7636_8799.t132 CSoutput.t15 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 gnd.t222 commonsourceibias.t109 CSoutput.t130 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 gnd.t29 gnd.t26 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X345 diffpairibias.t3 diffpairibias.t2 gnd.t324 gnd.t323 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X346 vdd.t44 a_n7636_8799.t133 CSoutput.t14 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 vdd.t218 vdd.t215 vdd.t217 vdd.t216 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X348 CSoutput.t129 commonsourceibias.t110 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 CSoutput.t13 a_n7636_8799.t134 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 output.t7 CSoutput.t208 vdd.t210 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X351 vdd.t199 CSoutput.t209 output.t6 gnd.t168 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X352 gnd.t218 commonsourceibias.t111 CSoutput.t128 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X353 vdd.t40 a_n7636_8799.t135 CSoutput.t12 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X354 gnd.t25 gnd.t22 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X355 CSoutput.t210 a_n1986_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X356 diffpairibias.t1 diffpairibias.t0 gnd.t326 gnd.t325 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X357 a_n7636_8799.t16 plus.t20 a_n3827_n3924.t20 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X358 CSoutput.t127 commonsourceibias.t112 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 outputibias.t1 outputibias.t0 gnd.t178 gnd.t177 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X360 CSoutput.t211 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X361 vdd.t177 a_n1986_13878.t65 a_n1808_13878.t12 vdd.t176 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X362 CSoutput.t11 a_n7636_8799.t136 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 CSoutput.t10 a_n7636_8799.t137 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 vdd.t34 a_n7636_8799.t138 CSoutput.t9 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 gnd.t214 commonsourceibias.t113 CSoutput.t126 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 vdd.t32 a_n7636_8799.t139 CSoutput.t8 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 CSoutput.t7 a_n7636_8799.t140 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X368 gnd.t21 gnd.t18 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X369 a_n1986_13878.t0 minus.t20 a_n3827_n3924.t0 gnd.t124 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X370 CSoutput.t6 a_n7636_8799.t141 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X371 vdd.t188 CSoutput.t212 output.t5 gnd.t155 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X372 a_n1986_8322.t2 a_n1986_13878.t66 a_n7636_8799.t3 vdd.t179 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X373 CSoutput.t125 commonsourceibias.t114 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X374 vdd.t26 a_n7636_8799.t142 CSoutput.t5 vdd.t25 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X375 vdd.t24 a_n7636_8799.t143 CSoutput.t4 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 CSoutput.t3 a_n7636_8799.t144 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X377 CSoutput.t2 a_n7636_8799.t145 vdd.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 vdd.t18 a_n7636_8799.t146 CSoutput.t1 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X379 gnd.t8 gnd.t5 gnd.t7 gnd.t6 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X380 gnd.t210 commonsourceibias.t115 CSoutput.t124 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X381 commonsourceibias.t47 commonsourceibias.t46 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 gnd.t17 gnd.t15 gnd.t16 gnd.t10 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X383 gnd.t14 gnd.t13 plus.t0 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X384 CSoutput.t123 commonsourceibias.t116 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X385 a_n1986_8322.t14 a_n1986_13878.t67 vdd.t3 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X386 a_n1808_13878.t1 a_n1986_13878.t14 a_n1986_13878.t15 vdd.t182 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X387 vdd.t189 CSoutput.t213 output.t4 gnd.t156 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X388 vdd.t15 a_n7636_8799.t147 CSoutput.t0 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X389 minus.t0 gnd.t2 gnd.t4 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X390 a_n3827_n3924.t29 diffpairibias.t29 gnd.t127 gnd.t126 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X391 CSoutput.t122 commonsourceibias.t117 gnd.t206 gnd.t205 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 CSoutput.t121 commonsourceibias.t118 gnd.t204 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X393 gnd.t197 commonsourceibias.t119 CSoutput.t120 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 a_n1986_13878.t25 a_n1986_13878.t24 a_n1808_13878.t0 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X395 vdd.t214 vdd.t211 vdd.t213 vdd.t212 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
R0 commonsourceibias.n25 commonsourceibias.t32 230.006
R1 commonsourceibias.n91 commonsourceibias.t96 230.006
R2 commonsourceibias.n218 commonsourceibias.t118 230.006
R3 commonsourceibias.n154 commonsourceibias.t98 230.006
R4 commonsourceibias.n322 commonsourceibias.t2 230.006
R5 commonsourceibias.n281 commonsourceibias.t69 230.006
R6 commonsourceibias.n483 commonsourceibias.t55 230.006
R7 commonsourceibias.n419 commonsourceibias.t79 230.006
R8 commonsourceibias.n70 commonsourceibias.t20 207.983
R9 commonsourceibias.n136 commonsourceibias.t57 207.983
R10 commonsourceibias.n263 commonsourceibias.t111 207.983
R11 commonsourceibias.n199 commonsourceibias.t88 207.983
R12 commonsourceibias.n368 commonsourceibias.t40 207.983
R13 commonsourceibias.n402 commonsourceibias.t114 207.983
R14 commonsourceibias.n529 commonsourceibias.t51 207.983
R15 commonsourceibias.n465 commonsourceibias.t74 207.983
R16 commonsourceibias.n10 commonsourceibias.t28 168.701
R17 commonsourceibias.n63 commonsourceibias.t0 168.701
R18 commonsourceibias.n57 commonsourceibias.t36 168.701
R19 commonsourceibias.n16 commonsourceibias.t14 168.701
R20 commonsourceibias.n49 commonsourceibias.t22 168.701
R21 commonsourceibias.n43 commonsourceibias.t30 168.701
R22 commonsourceibias.n19 commonsourceibias.t12 168.701
R23 commonsourceibias.n21 commonsourceibias.t38 168.701
R24 commonsourceibias.n23 commonsourceibias.t16 168.701
R25 commonsourceibias.n26 commonsourceibias.t4 168.701
R26 commonsourceibias.n1 commonsourceibias.t110 168.701
R27 commonsourceibias.n129 commonsourceibias.t70 168.701
R28 commonsourceibias.n123 commonsourceibias.t117 168.701
R29 commonsourceibias.n7 commonsourceibias.t85 168.701
R30 commonsourceibias.n115 commonsourceibias.t54 168.701
R31 commonsourceibias.n109 commonsourceibias.t97 168.701
R32 commonsourceibias.n85 commonsourceibias.t86 168.701
R33 commonsourceibias.n87 commonsourceibias.t115 168.701
R34 commonsourceibias.n89 commonsourceibias.t80 168.701
R35 commonsourceibias.n92 commonsourceibias.t66 168.701
R36 commonsourceibias.n219 commonsourceibias.t75 168.701
R37 commonsourceibias.n216 commonsourceibias.t60 168.701
R38 commonsourceibias.n214 commonsourceibias.t49 168.701
R39 commonsourceibias.n212 commonsourceibias.t84 168.701
R40 commonsourceibias.n236 commonsourceibias.t93 168.701
R41 commonsourceibias.n242 commonsourceibias.t53 168.701
R42 commonsourceibias.n209 commonsourceibias.t119 168.701
R43 commonsourceibias.n250 commonsourceibias.t104 168.701
R44 commonsourceibias.n256 commonsourceibias.t59 168.701
R45 commonsourceibias.n203 commonsourceibias.t50 168.701
R46 commonsourceibias.n139 commonsourceibias.t105 168.701
R47 commonsourceibias.n192 commonsourceibias.t101 168.701
R48 commonsourceibias.n186 commonsourceibias.t89 168.701
R49 commonsourceibias.n145 commonsourceibias.t106 168.701
R50 commonsourceibias.n178 commonsourceibias.t99 168.701
R51 commonsourceibias.n172 commonsourceibias.t87 168.701
R52 commonsourceibias.n148 commonsourceibias.t107 168.701
R53 commonsourceibias.n150 commonsourceibias.t100 168.701
R54 commonsourceibias.n152 commonsourceibias.t112 168.701
R55 commonsourceibias.n155 commonsourceibias.t108 168.701
R56 commonsourceibias.n323 commonsourceibias.t44 168.701
R57 commonsourceibias.n320 commonsourceibias.t26 168.701
R58 commonsourceibias.n318 commonsourceibias.t10 168.701
R59 commonsourceibias.n316 commonsourceibias.t6 168.701
R60 commonsourceibias.n340 commonsourceibias.t46 168.701
R61 commonsourceibias.n346 commonsourceibias.t42 168.701
R62 commonsourceibias.n348 commonsourceibias.t8 168.701
R63 commonsourceibias.n355 commonsourceibias.t34 168.701
R64 commonsourceibias.n361 commonsourceibias.t24 168.701
R65 commonsourceibias.n308 commonsourceibias.t18 168.701
R66 commonsourceibias.n267 commonsourceibias.t78 168.701
R67 commonsourceibias.n395 commonsourceibias.t52 168.701
R68 commonsourceibias.n389 commonsourceibias.t94 168.701
R69 commonsourceibias.n382 commonsourceibias.t64 168.701
R70 commonsourceibias.n380 commonsourceibias.t113 168.701
R71 commonsourceibias.n282 commonsourceibias.t58 168.701
R72 commonsourceibias.n279 commonsourceibias.t63 168.701
R73 commonsourceibias.n277 commonsourceibias.t92 168.701
R74 commonsourceibias.n275 commonsourceibias.t65 168.701
R75 commonsourceibias.n299 commonsourceibias.t76 168.701
R76 commonsourceibias.n484 commonsourceibias.t68 168.701
R77 commonsourceibias.n481 commonsourceibias.t72 168.701
R78 commonsourceibias.n479 commonsourceibias.t61 168.701
R79 commonsourceibias.n477 commonsourceibias.t109 168.701
R80 commonsourceibias.n501 commonsourceibias.t77 168.701
R81 commonsourceibias.n507 commonsourceibias.t67 168.701
R82 commonsourceibias.n509 commonsourceibias.t56 168.701
R83 commonsourceibias.n516 commonsourceibias.t48 168.701
R84 commonsourceibias.n522 commonsourceibias.t71 168.701
R85 commonsourceibias.n469 commonsourceibias.t62 168.701
R86 commonsourceibias.n420 commonsourceibias.t116 168.701
R87 commonsourceibias.n417 commonsourceibias.t102 168.701
R88 commonsourceibias.n415 commonsourceibias.t81 168.701
R89 commonsourceibias.n413 commonsourceibias.t95 168.701
R90 commonsourceibias.n437 commonsourceibias.t103 168.701
R91 commonsourceibias.n443 commonsourceibias.t83 168.701
R92 commonsourceibias.n445 commonsourceibias.t90 168.701
R93 commonsourceibias.n452 commonsourceibias.t73 168.701
R94 commonsourceibias.n458 commonsourceibias.t82 168.701
R95 commonsourceibias.n405 commonsourceibias.t91 168.701
R96 commonsourceibias.n27 commonsourceibias.n24 161.3
R97 commonsourceibias.n29 commonsourceibias.n28 161.3
R98 commonsourceibias.n31 commonsourceibias.n30 161.3
R99 commonsourceibias.n32 commonsourceibias.n22 161.3
R100 commonsourceibias.n34 commonsourceibias.n33 161.3
R101 commonsourceibias.n36 commonsourceibias.n35 161.3
R102 commonsourceibias.n37 commonsourceibias.n20 161.3
R103 commonsourceibias.n39 commonsourceibias.n38 161.3
R104 commonsourceibias.n41 commonsourceibias.n40 161.3
R105 commonsourceibias.n42 commonsourceibias.n18 161.3
R106 commonsourceibias.n45 commonsourceibias.n44 161.3
R107 commonsourceibias.n46 commonsourceibias.n17 161.3
R108 commonsourceibias.n48 commonsourceibias.n47 161.3
R109 commonsourceibias.n50 commonsourceibias.n15 161.3
R110 commonsourceibias.n52 commonsourceibias.n51 161.3
R111 commonsourceibias.n53 commonsourceibias.n14 161.3
R112 commonsourceibias.n55 commonsourceibias.n54 161.3
R113 commonsourceibias.n56 commonsourceibias.n13 161.3
R114 commonsourceibias.n59 commonsourceibias.n58 161.3
R115 commonsourceibias.n60 commonsourceibias.n12 161.3
R116 commonsourceibias.n62 commonsourceibias.n61 161.3
R117 commonsourceibias.n64 commonsourceibias.n11 161.3
R118 commonsourceibias.n66 commonsourceibias.n65 161.3
R119 commonsourceibias.n68 commonsourceibias.n67 161.3
R120 commonsourceibias.n69 commonsourceibias.n9 161.3
R121 commonsourceibias.n93 commonsourceibias.n90 161.3
R122 commonsourceibias.n95 commonsourceibias.n94 161.3
R123 commonsourceibias.n97 commonsourceibias.n96 161.3
R124 commonsourceibias.n98 commonsourceibias.n88 161.3
R125 commonsourceibias.n100 commonsourceibias.n99 161.3
R126 commonsourceibias.n102 commonsourceibias.n101 161.3
R127 commonsourceibias.n103 commonsourceibias.n86 161.3
R128 commonsourceibias.n105 commonsourceibias.n104 161.3
R129 commonsourceibias.n107 commonsourceibias.n106 161.3
R130 commonsourceibias.n108 commonsourceibias.n84 161.3
R131 commonsourceibias.n111 commonsourceibias.n110 161.3
R132 commonsourceibias.n112 commonsourceibias.n8 161.3
R133 commonsourceibias.n114 commonsourceibias.n113 161.3
R134 commonsourceibias.n116 commonsourceibias.n6 161.3
R135 commonsourceibias.n118 commonsourceibias.n117 161.3
R136 commonsourceibias.n119 commonsourceibias.n5 161.3
R137 commonsourceibias.n121 commonsourceibias.n120 161.3
R138 commonsourceibias.n122 commonsourceibias.n4 161.3
R139 commonsourceibias.n125 commonsourceibias.n124 161.3
R140 commonsourceibias.n126 commonsourceibias.n3 161.3
R141 commonsourceibias.n128 commonsourceibias.n127 161.3
R142 commonsourceibias.n130 commonsourceibias.n2 161.3
R143 commonsourceibias.n132 commonsourceibias.n131 161.3
R144 commonsourceibias.n134 commonsourceibias.n133 161.3
R145 commonsourceibias.n135 commonsourceibias.n0 161.3
R146 commonsourceibias.n262 commonsourceibias.n202 161.3
R147 commonsourceibias.n261 commonsourceibias.n260 161.3
R148 commonsourceibias.n259 commonsourceibias.n258 161.3
R149 commonsourceibias.n257 commonsourceibias.n204 161.3
R150 commonsourceibias.n255 commonsourceibias.n254 161.3
R151 commonsourceibias.n253 commonsourceibias.n205 161.3
R152 commonsourceibias.n252 commonsourceibias.n251 161.3
R153 commonsourceibias.n249 commonsourceibias.n206 161.3
R154 commonsourceibias.n248 commonsourceibias.n247 161.3
R155 commonsourceibias.n246 commonsourceibias.n207 161.3
R156 commonsourceibias.n245 commonsourceibias.n244 161.3
R157 commonsourceibias.n243 commonsourceibias.n208 161.3
R158 commonsourceibias.n241 commonsourceibias.n240 161.3
R159 commonsourceibias.n239 commonsourceibias.n210 161.3
R160 commonsourceibias.n238 commonsourceibias.n237 161.3
R161 commonsourceibias.n235 commonsourceibias.n211 161.3
R162 commonsourceibias.n234 commonsourceibias.n233 161.3
R163 commonsourceibias.n232 commonsourceibias.n231 161.3
R164 commonsourceibias.n230 commonsourceibias.n213 161.3
R165 commonsourceibias.n229 commonsourceibias.n228 161.3
R166 commonsourceibias.n227 commonsourceibias.n226 161.3
R167 commonsourceibias.n225 commonsourceibias.n215 161.3
R168 commonsourceibias.n224 commonsourceibias.n223 161.3
R169 commonsourceibias.n222 commonsourceibias.n221 161.3
R170 commonsourceibias.n220 commonsourceibias.n217 161.3
R171 commonsourceibias.n156 commonsourceibias.n153 161.3
R172 commonsourceibias.n158 commonsourceibias.n157 161.3
R173 commonsourceibias.n160 commonsourceibias.n159 161.3
R174 commonsourceibias.n161 commonsourceibias.n151 161.3
R175 commonsourceibias.n163 commonsourceibias.n162 161.3
R176 commonsourceibias.n165 commonsourceibias.n164 161.3
R177 commonsourceibias.n166 commonsourceibias.n149 161.3
R178 commonsourceibias.n168 commonsourceibias.n167 161.3
R179 commonsourceibias.n170 commonsourceibias.n169 161.3
R180 commonsourceibias.n171 commonsourceibias.n147 161.3
R181 commonsourceibias.n174 commonsourceibias.n173 161.3
R182 commonsourceibias.n175 commonsourceibias.n146 161.3
R183 commonsourceibias.n177 commonsourceibias.n176 161.3
R184 commonsourceibias.n179 commonsourceibias.n144 161.3
R185 commonsourceibias.n181 commonsourceibias.n180 161.3
R186 commonsourceibias.n182 commonsourceibias.n143 161.3
R187 commonsourceibias.n184 commonsourceibias.n183 161.3
R188 commonsourceibias.n185 commonsourceibias.n142 161.3
R189 commonsourceibias.n188 commonsourceibias.n187 161.3
R190 commonsourceibias.n189 commonsourceibias.n141 161.3
R191 commonsourceibias.n191 commonsourceibias.n190 161.3
R192 commonsourceibias.n193 commonsourceibias.n140 161.3
R193 commonsourceibias.n195 commonsourceibias.n194 161.3
R194 commonsourceibias.n197 commonsourceibias.n196 161.3
R195 commonsourceibias.n198 commonsourceibias.n138 161.3
R196 commonsourceibias.n367 commonsourceibias.n307 161.3
R197 commonsourceibias.n366 commonsourceibias.n365 161.3
R198 commonsourceibias.n364 commonsourceibias.n363 161.3
R199 commonsourceibias.n362 commonsourceibias.n309 161.3
R200 commonsourceibias.n360 commonsourceibias.n359 161.3
R201 commonsourceibias.n358 commonsourceibias.n310 161.3
R202 commonsourceibias.n357 commonsourceibias.n356 161.3
R203 commonsourceibias.n354 commonsourceibias.n311 161.3
R204 commonsourceibias.n353 commonsourceibias.n352 161.3
R205 commonsourceibias.n351 commonsourceibias.n312 161.3
R206 commonsourceibias.n350 commonsourceibias.n349 161.3
R207 commonsourceibias.n347 commonsourceibias.n313 161.3
R208 commonsourceibias.n345 commonsourceibias.n344 161.3
R209 commonsourceibias.n343 commonsourceibias.n314 161.3
R210 commonsourceibias.n342 commonsourceibias.n341 161.3
R211 commonsourceibias.n339 commonsourceibias.n315 161.3
R212 commonsourceibias.n338 commonsourceibias.n337 161.3
R213 commonsourceibias.n336 commonsourceibias.n335 161.3
R214 commonsourceibias.n334 commonsourceibias.n317 161.3
R215 commonsourceibias.n333 commonsourceibias.n332 161.3
R216 commonsourceibias.n331 commonsourceibias.n330 161.3
R217 commonsourceibias.n329 commonsourceibias.n319 161.3
R218 commonsourceibias.n328 commonsourceibias.n327 161.3
R219 commonsourceibias.n326 commonsourceibias.n325 161.3
R220 commonsourceibias.n324 commonsourceibias.n321 161.3
R221 commonsourceibias.n301 commonsourceibias.n300 161.3
R222 commonsourceibias.n298 commonsourceibias.n274 161.3
R223 commonsourceibias.n297 commonsourceibias.n296 161.3
R224 commonsourceibias.n295 commonsourceibias.n294 161.3
R225 commonsourceibias.n293 commonsourceibias.n276 161.3
R226 commonsourceibias.n292 commonsourceibias.n291 161.3
R227 commonsourceibias.n290 commonsourceibias.n289 161.3
R228 commonsourceibias.n288 commonsourceibias.n278 161.3
R229 commonsourceibias.n287 commonsourceibias.n286 161.3
R230 commonsourceibias.n285 commonsourceibias.n284 161.3
R231 commonsourceibias.n283 commonsourceibias.n280 161.3
R232 commonsourceibias.n377 commonsourceibias.n273 161.3
R233 commonsourceibias.n401 commonsourceibias.n266 161.3
R234 commonsourceibias.n400 commonsourceibias.n399 161.3
R235 commonsourceibias.n398 commonsourceibias.n397 161.3
R236 commonsourceibias.n396 commonsourceibias.n268 161.3
R237 commonsourceibias.n394 commonsourceibias.n393 161.3
R238 commonsourceibias.n392 commonsourceibias.n269 161.3
R239 commonsourceibias.n391 commonsourceibias.n390 161.3
R240 commonsourceibias.n388 commonsourceibias.n270 161.3
R241 commonsourceibias.n387 commonsourceibias.n386 161.3
R242 commonsourceibias.n385 commonsourceibias.n271 161.3
R243 commonsourceibias.n384 commonsourceibias.n383 161.3
R244 commonsourceibias.n381 commonsourceibias.n272 161.3
R245 commonsourceibias.n379 commonsourceibias.n378 161.3
R246 commonsourceibias.n528 commonsourceibias.n468 161.3
R247 commonsourceibias.n527 commonsourceibias.n526 161.3
R248 commonsourceibias.n525 commonsourceibias.n524 161.3
R249 commonsourceibias.n523 commonsourceibias.n470 161.3
R250 commonsourceibias.n521 commonsourceibias.n520 161.3
R251 commonsourceibias.n519 commonsourceibias.n471 161.3
R252 commonsourceibias.n518 commonsourceibias.n517 161.3
R253 commonsourceibias.n515 commonsourceibias.n472 161.3
R254 commonsourceibias.n514 commonsourceibias.n513 161.3
R255 commonsourceibias.n512 commonsourceibias.n473 161.3
R256 commonsourceibias.n511 commonsourceibias.n510 161.3
R257 commonsourceibias.n508 commonsourceibias.n474 161.3
R258 commonsourceibias.n506 commonsourceibias.n505 161.3
R259 commonsourceibias.n504 commonsourceibias.n475 161.3
R260 commonsourceibias.n503 commonsourceibias.n502 161.3
R261 commonsourceibias.n500 commonsourceibias.n476 161.3
R262 commonsourceibias.n499 commonsourceibias.n498 161.3
R263 commonsourceibias.n497 commonsourceibias.n496 161.3
R264 commonsourceibias.n495 commonsourceibias.n478 161.3
R265 commonsourceibias.n494 commonsourceibias.n493 161.3
R266 commonsourceibias.n492 commonsourceibias.n491 161.3
R267 commonsourceibias.n490 commonsourceibias.n480 161.3
R268 commonsourceibias.n489 commonsourceibias.n488 161.3
R269 commonsourceibias.n487 commonsourceibias.n486 161.3
R270 commonsourceibias.n485 commonsourceibias.n482 161.3
R271 commonsourceibias.n464 commonsourceibias.n404 161.3
R272 commonsourceibias.n463 commonsourceibias.n462 161.3
R273 commonsourceibias.n461 commonsourceibias.n460 161.3
R274 commonsourceibias.n459 commonsourceibias.n406 161.3
R275 commonsourceibias.n457 commonsourceibias.n456 161.3
R276 commonsourceibias.n455 commonsourceibias.n407 161.3
R277 commonsourceibias.n454 commonsourceibias.n453 161.3
R278 commonsourceibias.n451 commonsourceibias.n408 161.3
R279 commonsourceibias.n450 commonsourceibias.n449 161.3
R280 commonsourceibias.n448 commonsourceibias.n409 161.3
R281 commonsourceibias.n447 commonsourceibias.n446 161.3
R282 commonsourceibias.n444 commonsourceibias.n410 161.3
R283 commonsourceibias.n442 commonsourceibias.n441 161.3
R284 commonsourceibias.n440 commonsourceibias.n411 161.3
R285 commonsourceibias.n439 commonsourceibias.n438 161.3
R286 commonsourceibias.n436 commonsourceibias.n412 161.3
R287 commonsourceibias.n435 commonsourceibias.n434 161.3
R288 commonsourceibias.n433 commonsourceibias.n432 161.3
R289 commonsourceibias.n431 commonsourceibias.n414 161.3
R290 commonsourceibias.n430 commonsourceibias.n429 161.3
R291 commonsourceibias.n428 commonsourceibias.n427 161.3
R292 commonsourceibias.n426 commonsourceibias.n416 161.3
R293 commonsourceibias.n425 commonsourceibias.n424 161.3
R294 commonsourceibias.n423 commonsourceibias.n422 161.3
R295 commonsourceibias.n421 commonsourceibias.n418 161.3
R296 commonsourceibias.n80 commonsourceibias.n78 81.5057
R297 commonsourceibias.n304 commonsourceibias.n302 81.5057
R298 commonsourceibias.n80 commonsourceibias.n79 80.9324
R299 commonsourceibias.n82 commonsourceibias.n81 80.9324
R300 commonsourceibias.n77 commonsourceibias.n76 80.9324
R301 commonsourceibias.n75 commonsourceibias.n74 80.9324
R302 commonsourceibias.n73 commonsourceibias.n72 80.9324
R303 commonsourceibias.n371 commonsourceibias.n370 80.9324
R304 commonsourceibias.n373 commonsourceibias.n372 80.9324
R305 commonsourceibias.n375 commonsourceibias.n374 80.9324
R306 commonsourceibias.n306 commonsourceibias.n305 80.9324
R307 commonsourceibias.n304 commonsourceibias.n303 80.9324
R308 commonsourceibias.n71 commonsourceibias.n70 80.6037
R309 commonsourceibias.n137 commonsourceibias.n136 80.6037
R310 commonsourceibias.n264 commonsourceibias.n263 80.6037
R311 commonsourceibias.n200 commonsourceibias.n199 80.6037
R312 commonsourceibias.n369 commonsourceibias.n368 80.6037
R313 commonsourceibias.n403 commonsourceibias.n402 80.6037
R314 commonsourceibias.n530 commonsourceibias.n529 80.6037
R315 commonsourceibias.n466 commonsourceibias.n465 80.6037
R316 commonsourceibias.n65 commonsourceibias.n64 56.5617
R317 commonsourceibias.n51 commonsourceibias.n50 56.5617
R318 commonsourceibias.n42 commonsourceibias.n41 56.5617
R319 commonsourceibias.n28 commonsourceibias.n27 56.5617
R320 commonsourceibias.n131 commonsourceibias.n130 56.5617
R321 commonsourceibias.n117 commonsourceibias.n116 56.5617
R322 commonsourceibias.n108 commonsourceibias.n107 56.5617
R323 commonsourceibias.n94 commonsourceibias.n93 56.5617
R324 commonsourceibias.n221 commonsourceibias.n220 56.5617
R325 commonsourceibias.n235 commonsourceibias.n234 56.5617
R326 commonsourceibias.n244 commonsourceibias.n243 56.5617
R327 commonsourceibias.n258 commonsourceibias.n257 56.5617
R328 commonsourceibias.n194 commonsourceibias.n193 56.5617
R329 commonsourceibias.n180 commonsourceibias.n179 56.5617
R330 commonsourceibias.n171 commonsourceibias.n170 56.5617
R331 commonsourceibias.n157 commonsourceibias.n156 56.5617
R332 commonsourceibias.n325 commonsourceibias.n324 56.5617
R333 commonsourceibias.n339 commonsourceibias.n338 56.5617
R334 commonsourceibias.n349 commonsourceibias.n347 56.5617
R335 commonsourceibias.n363 commonsourceibias.n362 56.5617
R336 commonsourceibias.n397 commonsourceibias.n396 56.5617
R337 commonsourceibias.n383 commonsourceibias.n381 56.5617
R338 commonsourceibias.n284 commonsourceibias.n283 56.5617
R339 commonsourceibias.n298 commonsourceibias.n297 56.5617
R340 commonsourceibias.n486 commonsourceibias.n485 56.5617
R341 commonsourceibias.n500 commonsourceibias.n499 56.5617
R342 commonsourceibias.n510 commonsourceibias.n508 56.5617
R343 commonsourceibias.n524 commonsourceibias.n523 56.5617
R344 commonsourceibias.n422 commonsourceibias.n421 56.5617
R345 commonsourceibias.n436 commonsourceibias.n435 56.5617
R346 commonsourceibias.n446 commonsourceibias.n444 56.5617
R347 commonsourceibias.n460 commonsourceibias.n459 56.5617
R348 commonsourceibias.n56 commonsourceibias.n55 56.0773
R349 commonsourceibias.n37 commonsourceibias.n36 56.0773
R350 commonsourceibias.n122 commonsourceibias.n121 56.0773
R351 commonsourceibias.n103 commonsourceibias.n102 56.0773
R352 commonsourceibias.n230 commonsourceibias.n229 56.0773
R353 commonsourceibias.n249 commonsourceibias.n248 56.0773
R354 commonsourceibias.n185 commonsourceibias.n184 56.0773
R355 commonsourceibias.n166 commonsourceibias.n165 56.0773
R356 commonsourceibias.n334 commonsourceibias.n333 56.0773
R357 commonsourceibias.n354 commonsourceibias.n353 56.0773
R358 commonsourceibias.n388 commonsourceibias.n387 56.0773
R359 commonsourceibias.n293 commonsourceibias.n292 56.0773
R360 commonsourceibias.n495 commonsourceibias.n494 56.0773
R361 commonsourceibias.n515 commonsourceibias.n514 56.0773
R362 commonsourceibias.n431 commonsourceibias.n430 56.0773
R363 commonsourceibias.n451 commonsourceibias.n450 56.0773
R364 commonsourceibias.n70 commonsourceibias.n69 46.0096
R365 commonsourceibias.n136 commonsourceibias.n135 46.0096
R366 commonsourceibias.n263 commonsourceibias.n262 46.0096
R367 commonsourceibias.n199 commonsourceibias.n198 46.0096
R368 commonsourceibias.n368 commonsourceibias.n367 46.0096
R369 commonsourceibias.n402 commonsourceibias.n401 46.0096
R370 commonsourceibias.n529 commonsourceibias.n528 46.0096
R371 commonsourceibias.n465 commonsourceibias.n464 46.0096
R372 commonsourceibias.n58 commonsourceibias.n12 41.5458
R373 commonsourceibias.n33 commonsourceibias.n32 41.5458
R374 commonsourceibias.n124 commonsourceibias.n3 41.5458
R375 commonsourceibias.n99 commonsourceibias.n98 41.5458
R376 commonsourceibias.n226 commonsourceibias.n225 41.5458
R377 commonsourceibias.n251 commonsourceibias.n205 41.5458
R378 commonsourceibias.n187 commonsourceibias.n141 41.5458
R379 commonsourceibias.n162 commonsourceibias.n161 41.5458
R380 commonsourceibias.n330 commonsourceibias.n329 41.5458
R381 commonsourceibias.n356 commonsourceibias.n310 41.5458
R382 commonsourceibias.n390 commonsourceibias.n269 41.5458
R383 commonsourceibias.n289 commonsourceibias.n288 41.5458
R384 commonsourceibias.n491 commonsourceibias.n490 41.5458
R385 commonsourceibias.n517 commonsourceibias.n471 41.5458
R386 commonsourceibias.n427 commonsourceibias.n426 41.5458
R387 commonsourceibias.n453 commonsourceibias.n407 41.5458
R388 commonsourceibias.n48 commonsourceibias.n17 40.577
R389 commonsourceibias.n44 commonsourceibias.n17 40.577
R390 commonsourceibias.n114 commonsourceibias.n8 40.577
R391 commonsourceibias.n110 commonsourceibias.n8 40.577
R392 commonsourceibias.n237 commonsourceibias.n210 40.577
R393 commonsourceibias.n241 commonsourceibias.n210 40.577
R394 commonsourceibias.n177 commonsourceibias.n146 40.577
R395 commonsourceibias.n173 commonsourceibias.n146 40.577
R396 commonsourceibias.n341 commonsourceibias.n314 40.577
R397 commonsourceibias.n345 commonsourceibias.n314 40.577
R398 commonsourceibias.n379 commonsourceibias.n273 40.577
R399 commonsourceibias.n300 commonsourceibias.n273 40.577
R400 commonsourceibias.n502 commonsourceibias.n475 40.577
R401 commonsourceibias.n506 commonsourceibias.n475 40.577
R402 commonsourceibias.n438 commonsourceibias.n411 40.577
R403 commonsourceibias.n442 commonsourceibias.n411 40.577
R404 commonsourceibias.n62 commonsourceibias.n12 39.6083
R405 commonsourceibias.n32 commonsourceibias.n31 39.6083
R406 commonsourceibias.n128 commonsourceibias.n3 39.6083
R407 commonsourceibias.n98 commonsourceibias.n97 39.6083
R408 commonsourceibias.n225 commonsourceibias.n224 39.6083
R409 commonsourceibias.n255 commonsourceibias.n205 39.6083
R410 commonsourceibias.n191 commonsourceibias.n141 39.6083
R411 commonsourceibias.n161 commonsourceibias.n160 39.6083
R412 commonsourceibias.n329 commonsourceibias.n328 39.6083
R413 commonsourceibias.n360 commonsourceibias.n310 39.6083
R414 commonsourceibias.n394 commonsourceibias.n269 39.6083
R415 commonsourceibias.n288 commonsourceibias.n287 39.6083
R416 commonsourceibias.n490 commonsourceibias.n489 39.6083
R417 commonsourceibias.n521 commonsourceibias.n471 39.6083
R418 commonsourceibias.n426 commonsourceibias.n425 39.6083
R419 commonsourceibias.n457 commonsourceibias.n407 39.6083
R420 commonsourceibias.n26 commonsourceibias.n25 33.0515
R421 commonsourceibias.n92 commonsourceibias.n91 33.0515
R422 commonsourceibias.n155 commonsourceibias.n154 33.0515
R423 commonsourceibias.n219 commonsourceibias.n218 33.0515
R424 commonsourceibias.n323 commonsourceibias.n322 33.0515
R425 commonsourceibias.n282 commonsourceibias.n281 33.0515
R426 commonsourceibias.n484 commonsourceibias.n483 33.0515
R427 commonsourceibias.n420 commonsourceibias.n419 33.0515
R428 commonsourceibias.n25 commonsourceibias.n24 28.5514
R429 commonsourceibias.n91 commonsourceibias.n90 28.5514
R430 commonsourceibias.n218 commonsourceibias.n217 28.5514
R431 commonsourceibias.n154 commonsourceibias.n153 28.5514
R432 commonsourceibias.n322 commonsourceibias.n321 28.5514
R433 commonsourceibias.n281 commonsourceibias.n280 28.5514
R434 commonsourceibias.n483 commonsourceibias.n482 28.5514
R435 commonsourceibias.n419 commonsourceibias.n418 28.5514
R436 commonsourceibias.n69 commonsourceibias.n68 26.0455
R437 commonsourceibias.n135 commonsourceibias.n134 26.0455
R438 commonsourceibias.n262 commonsourceibias.n261 26.0455
R439 commonsourceibias.n198 commonsourceibias.n197 26.0455
R440 commonsourceibias.n367 commonsourceibias.n366 26.0455
R441 commonsourceibias.n401 commonsourceibias.n400 26.0455
R442 commonsourceibias.n528 commonsourceibias.n527 26.0455
R443 commonsourceibias.n464 commonsourceibias.n463 26.0455
R444 commonsourceibias.n55 commonsourceibias.n14 25.0767
R445 commonsourceibias.n38 commonsourceibias.n37 25.0767
R446 commonsourceibias.n121 commonsourceibias.n5 25.0767
R447 commonsourceibias.n104 commonsourceibias.n103 25.0767
R448 commonsourceibias.n231 commonsourceibias.n230 25.0767
R449 commonsourceibias.n248 commonsourceibias.n207 25.0767
R450 commonsourceibias.n184 commonsourceibias.n143 25.0767
R451 commonsourceibias.n167 commonsourceibias.n166 25.0767
R452 commonsourceibias.n335 commonsourceibias.n334 25.0767
R453 commonsourceibias.n353 commonsourceibias.n312 25.0767
R454 commonsourceibias.n387 commonsourceibias.n271 25.0767
R455 commonsourceibias.n294 commonsourceibias.n293 25.0767
R456 commonsourceibias.n496 commonsourceibias.n495 25.0767
R457 commonsourceibias.n514 commonsourceibias.n473 25.0767
R458 commonsourceibias.n432 commonsourceibias.n431 25.0767
R459 commonsourceibias.n450 commonsourceibias.n409 25.0767
R460 commonsourceibias.n51 commonsourceibias.n16 24.3464
R461 commonsourceibias.n41 commonsourceibias.n19 24.3464
R462 commonsourceibias.n117 commonsourceibias.n7 24.3464
R463 commonsourceibias.n107 commonsourceibias.n85 24.3464
R464 commonsourceibias.n234 commonsourceibias.n212 24.3464
R465 commonsourceibias.n244 commonsourceibias.n209 24.3464
R466 commonsourceibias.n180 commonsourceibias.n145 24.3464
R467 commonsourceibias.n170 commonsourceibias.n148 24.3464
R468 commonsourceibias.n338 commonsourceibias.n316 24.3464
R469 commonsourceibias.n349 commonsourceibias.n348 24.3464
R470 commonsourceibias.n383 commonsourceibias.n382 24.3464
R471 commonsourceibias.n297 commonsourceibias.n275 24.3464
R472 commonsourceibias.n499 commonsourceibias.n477 24.3464
R473 commonsourceibias.n510 commonsourceibias.n509 24.3464
R474 commonsourceibias.n435 commonsourceibias.n413 24.3464
R475 commonsourceibias.n446 commonsourceibias.n445 24.3464
R476 commonsourceibias.n65 commonsourceibias.n10 23.8546
R477 commonsourceibias.n27 commonsourceibias.n26 23.8546
R478 commonsourceibias.n131 commonsourceibias.n1 23.8546
R479 commonsourceibias.n93 commonsourceibias.n92 23.8546
R480 commonsourceibias.n220 commonsourceibias.n219 23.8546
R481 commonsourceibias.n258 commonsourceibias.n203 23.8546
R482 commonsourceibias.n194 commonsourceibias.n139 23.8546
R483 commonsourceibias.n156 commonsourceibias.n155 23.8546
R484 commonsourceibias.n324 commonsourceibias.n323 23.8546
R485 commonsourceibias.n363 commonsourceibias.n308 23.8546
R486 commonsourceibias.n397 commonsourceibias.n267 23.8546
R487 commonsourceibias.n283 commonsourceibias.n282 23.8546
R488 commonsourceibias.n485 commonsourceibias.n484 23.8546
R489 commonsourceibias.n524 commonsourceibias.n469 23.8546
R490 commonsourceibias.n421 commonsourceibias.n420 23.8546
R491 commonsourceibias.n460 commonsourceibias.n405 23.8546
R492 commonsourceibias.n64 commonsourceibias.n63 16.9689
R493 commonsourceibias.n28 commonsourceibias.n23 16.9689
R494 commonsourceibias.n130 commonsourceibias.n129 16.9689
R495 commonsourceibias.n94 commonsourceibias.n89 16.9689
R496 commonsourceibias.n221 commonsourceibias.n216 16.9689
R497 commonsourceibias.n257 commonsourceibias.n256 16.9689
R498 commonsourceibias.n193 commonsourceibias.n192 16.9689
R499 commonsourceibias.n157 commonsourceibias.n152 16.9689
R500 commonsourceibias.n325 commonsourceibias.n320 16.9689
R501 commonsourceibias.n362 commonsourceibias.n361 16.9689
R502 commonsourceibias.n396 commonsourceibias.n395 16.9689
R503 commonsourceibias.n284 commonsourceibias.n279 16.9689
R504 commonsourceibias.n486 commonsourceibias.n481 16.9689
R505 commonsourceibias.n523 commonsourceibias.n522 16.9689
R506 commonsourceibias.n422 commonsourceibias.n417 16.9689
R507 commonsourceibias.n459 commonsourceibias.n458 16.9689
R508 commonsourceibias.n50 commonsourceibias.n49 16.477
R509 commonsourceibias.n43 commonsourceibias.n42 16.477
R510 commonsourceibias.n116 commonsourceibias.n115 16.477
R511 commonsourceibias.n109 commonsourceibias.n108 16.477
R512 commonsourceibias.n236 commonsourceibias.n235 16.477
R513 commonsourceibias.n243 commonsourceibias.n242 16.477
R514 commonsourceibias.n179 commonsourceibias.n178 16.477
R515 commonsourceibias.n172 commonsourceibias.n171 16.477
R516 commonsourceibias.n340 commonsourceibias.n339 16.477
R517 commonsourceibias.n347 commonsourceibias.n346 16.477
R518 commonsourceibias.n381 commonsourceibias.n380 16.477
R519 commonsourceibias.n299 commonsourceibias.n298 16.477
R520 commonsourceibias.n501 commonsourceibias.n500 16.477
R521 commonsourceibias.n508 commonsourceibias.n507 16.477
R522 commonsourceibias.n437 commonsourceibias.n436 16.477
R523 commonsourceibias.n444 commonsourceibias.n443 16.477
R524 commonsourceibias.n57 commonsourceibias.n56 15.9852
R525 commonsourceibias.n36 commonsourceibias.n21 15.9852
R526 commonsourceibias.n123 commonsourceibias.n122 15.9852
R527 commonsourceibias.n102 commonsourceibias.n87 15.9852
R528 commonsourceibias.n229 commonsourceibias.n214 15.9852
R529 commonsourceibias.n250 commonsourceibias.n249 15.9852
R530 commonsourceibias.n186 commonsourceibias.n185 15.9852
R531 commonsourceibias.n165 commonsourceibias.n150 15.9852
R532 commonsourceibias.n333 commonsourceibias.n318 15.9852
R533 commonsourceibias.n355 commonsourceibias.n354 15.9852
R534 commonsourceibias.n389 commonsourceibias.n388 15.9852
R535 commonsourceibias.n292 commonsourceibias.n277 15.9852
R536 commonsourceibias.n494 commonsourceibias.n479 15.9852
R537 commonsourceibias.n516 commonsourceibias.n515 15.9852
R538 commonsourceibias.n430 commonsourceibias.n415 15.9852
R539 commonsourceibias.n452 commonsourceibias.n451 15.9852
R540 commonsourceibias.n73 commonsourceibias.n71 13.2057
R541 commonsourceibias.n371 commonsourceibias.n369 13.2057
R542 commonsourceibias.n532 commonsourceibias.n265 10.4122
R543 commonsourceibias.n112 commonsourceibias.n83 9.50363
R544 commonsourceibias.n377 commonsourceibias.n376 9.50363
R545 commonsourceibias.n201 commonsourceibias.n137 8.7339
R546 commonsourceibias.n467 commonsourceibias.n403 8.7339
R547 commonsourceibias.n58 commonsourceibias.n57 8.60764
R548 commonsourceibias.n33 commonsourceibias.n21 8.60764
R549 commonsourceibias.n124 commonsourceibias.n123 8.60764
R550 commonsourceibias.n99 commonsourceibias.n87 8.60764
R551 commonsourceibias.n226 commonsourceibias.n214 8.60764
R552 commonsourceibias.n251 commonsourceibias.n250 8.60764
R553 commonsourceibias.n187 commonsourceibias.n186 8.60764
R554 commonsourceibias.n162 commonsourceibias.n150 8.60764
R555 commonsourceibias.n330 commonsourceibias.n318 8.60764
R556 commonsourceibias.n356 commonsourceibias.n355 8.60764
R557 commonsourceibias.n390 commonsourceibias.n389 8.60764
R558 commonsourceibias.n289 commonsourceibias.n277 8.60764
R559 commonsourceibias.n491 commonsourceibias.n479 8.60764
R560 commonsourceibias.n517 commonsourceibias.n516 8.60764
R561 commonsourceibias.n427 commonsourceibias.n415 8.60764
R562 commonsourceibias.n453 commonsourceibias.n452 8.60764
R563 commonsourceibias.n532 commonsourceibias.n531 8.46921
R564 commonsourceibias.n49 commonsourceibias.n48 8.11581
R565 commonsourceibias.n44 commonsourceibias.n43 8.11581
R566 commonsourceibias.n115 commonsourceibias.n114 8.11581
R567 commonsourceibias.n110 commonsourceibias.n109 8.11581
R568 commonsourceibias.n237 commonsourceibias.n236 8.11581
R569 commonsourceibias.n242 commonsourceibias.n241 8.11581
R570 commonsourceibias.n178 commonsourceibias.n177 8.11581
R571 commonsourceibias.n173 commonsourceibias.n172 8.11581
R572 commonsourceibias.n341 commonsourceibias.n340 8.11581
R573 commonsourceibias.n346 commonsourceibias.n345 8.11581
R574 commonsourceibias.n380 commonsourceibias.n379 8.11581
R575 commonsourceibias.n300 commonsourceibias.n299 8.11581
R576 commonsourceibias.n502 commonsourceibias.n501 8.11581
R577 commonsourceibias.n507 commonsourceibias.n506 8.11581
R578 commonsourceibias.n438 commonsourceibias.n437 8.11581
R579 commonsourceibias.n443 commonsourceibias.n442 8.11581
R580 commonsourceibias.n63 commonsourceibias.n62 7.62397
R581 commonsourceibias.n31 commonsourceibias.n23 7.62397
R582 commonsourceibias.n129 commonsourceibias.n128 7.62397
R583 commonsourceibias.n97 commonsourceibias.n89 7.62397
R584 commonsourceibias.n224 commonsourceibias.n216 7.62397
R585 commonsourceibias.n256 commonsourceibias.n255 7.62397
R586 commonsourceibias.n192 commonsourceibias.n191 7.62397
R587 commonsourceibias.n160 commonsourceibias.n152 7.62397
R588 commonsourceibias.n328 commonsourceibias.n320 7.62397
R589 commonsourceibias.n361 commonsourceibias.n360 7.62397
R590 commonsourceibias.n395 commonsourceibias.n394 7.62397
R591 commonsourceibias.n287 commonsourceibias.n279 7.62397
R592 commonsourceibias.n489 commonsourceibias.n481 7.62397
R593 commonsourceibias.n522 commonsourceibias.n521 7.62397
R594 commonsourceibias.n425 commonsourceibias.n417 7.62397
R595 commonsourceibias.n458 commonsourceibias.n457 7.62397
R596 commonsourceibias.n265 commonsourceibias.n264 5.00473
R597 commonsourceibias.n201 commonsourceibias.n200 5.00473
R598 commonsourceibias.n531 commonsourceibias.n530 5.00473
R599 commonsourceibias.n467 commonsourceibias.n466 5.00473
R600 commonsourceibias commonsourceibias.n532 3.87639
R601 commonsourceibias.n265 commonsourceibias.n201 3.72967
R602 commonsourceibias.n531 commonsourceibias.n467 3.72967
R603 commonsourceibias.n78 commonsourceibias.t5 2.82907
R604 commonsourceibias.n78 commonsourceibias.t33 2.82907
R605 commonsourceibias.n79 commonsourceibias.t39 2.82907
R606 commonsourceibias.n79 commonsourceibias.t17 2.82907
R607 commonsourceibias.n81 commonsourceibias.t31 2.82907
R608 commonsourceibias.n81 commonsourceibias.t13 2.82907
R609 commonsourceibias.n76 commonsourceibias.t15 2.82907
R610 commonsourceibias.n76 commonsourceibias.t23 2.82907
R611 commonsourceibias.n74 commonsourceibias.t1 2.82907
R612 commonsourceibias.n74 commonsourceibias.t37 2.82907
R613 commonsourceibias.n72 commonsourceibias.t21 2.82907
R614 commonsourceibias.n72 commonsourceibias.t29 2.82907
R615 commonsourceibias.n370 commonsourceibias.t19 2.82907
R616 commonsourceibias.n370 commonsourceibias.t41 2.82907
R617 commonsourceibias.n372 commonsourceibias.t35 2.82907
R618 commonsourceibias.n372 commonsourceibias.t25 2.82907
R619 commonsourceibias.n374 commonsourceibias.t43 2.82907
R620 commonsourceibias.n374 commonsourceibias.t9 2.82907
R621 commonsourceibias.n305 commonsourceibias.t7 2.82907
R622 commonsourceibias.n305 commonsourceibias.t47 2.82907
R623 commonsourceibias.n303 commonsourceibias.t27 2.82907
R624 commonsourceibias.n303 commonsourceibias.t11 2.82907
R625 commonsourceibias.n302 commonsourceibias.t3 2.82907
R626 commonsourceibias.n302 commonsourceibias.t45 2.82907
R627 commonsourceibias.n68 commonsourceibias.n10 0.738255
R628 commonsourceibias.n134 commonsourceibias.n1 0.738255
R629 commonsourceibias.n261 commonsourceibias.n203 0.738255
R630 commonsourceibias.n197 commonsourceibias.n139 0.738255
R631 commonsourceibias.n366 commonsourceibias.n308 0.738255
R632 commonsourceibias.n400 commonsourceibias.n267 0.738255
R633 commonsourceibias.n527 commonsourceibias.n469 0.738255
R634 commonsourceibias.n463 commonsourceibias.n405 0.738255
R635 commonsourceibias.n75 commonsourceibias.n73 0.573776
R636 commonsourceibias.n77 commonsourceibias.n75 0.573776
R637 commonsourceibias.n82 commonsourceibias.n80 0.573776
R638 commonsourceibias.n306 commonsourceibias.n304 0.573776
R639 commonsourceibias.n375 commonsourceibias.n373 0.573776
R640 commonsourceibias.n373 commonsourceibias.n371 0.573776
R641 commonsourceibias.n83 commonsourceibias.n77 0.287138
R642 commonsourceibias.n83 commonsourceibias.n82 0.287138
R643 commonsourceibias.n376 commonsourceibias.n306 0.287138
R644 commonsourceibias.n376 commonsourceibias.n375 0.287138
R645 commonsourceibias.n71 commonsourceibias.n9 0.285035
R646 commonsourceibias.n137 commonsourceibias.n0 0.285035
R647 commonsourceibias.n264 commonsourceibias.n202 0.285035
R648 commonsourceibias.n200 commonsourceibias.n138 0.285035
R649 commonsourceibias.n369 commonsourceibias.n307 0.285035
R650 commonsourceibias.n403 commonsourceibias.n266 0.285035
R651 commonsourceibias.n530 commonsourceibias.n468 0.285035
R652 commonsourceibias.n466 commonsourceibias.n404 0.285035
R653 commonsourceibias.n16 commonsourceibias.n14 0.246418
R654 commonsourceibias.n38 commonsourceibias.n19 0.246418
R655 commonsourceibias.n7 commonsourceibias.n5 0.246418
R656 commonsourceibias.n104 commonsourceibias.n85 0.246418
R657 commonsourceibias.n231 commonsourceibias.n212 0.246418
R658 commonsourceibias.n209 commonsourceibias.n207 0.246418
R659 commonsourceibias.n145 commonsourceibias.n143 0.246418
R660 commonsourceibias.n167 commonsourceibias.n148 0.246418
R661 commonsourceibias.n335 commonsourceibias.n316 0.246418
R662 commonsourceibias.n348 commonsourceibias.n312 0.246418
R663 commonsourceibias.n382 commonsourceibias.n271 0.246418
R664 commonsourceibias.n294 commonsourceibias.n275 0.246418
R665 commonsourceibias.n496 commonsourceibias.n477 0.246418
R666 commonsourceibias.n509 commonsourceibias.n473 0.246418
R667 commonsourceibias.n432 commonsourceibias.n413 0.246418
R668 commonsourceibias.n445 commonsourceibias.n409 0.246418
R669 commonsourceibias.n67 commonsourceibias.n9 0.189894
R670 commonsourceibias.n67 commonsourceibias.n66 0.189894
R671 commonsourceibias.n66 commonsourceibias.n11 0.189894
R672 commonsourceibias.n61 commonsourceibias.n11 0.189894
R673 commonsourceibias.n61 commonsourceibias.n60 0.189894
R674 commonsourceibias.n60 commonsourceibias.n59 0.189894
R675 commonsourceibias.n59 commonsourceibias.n13 0.189894
R676 commonsourceibias.n54 commonsourceibias.n13 0.189894
R677 commonsourceibias.n54 commonsourceibias.n53 0.189894
R678 commonsourceibias.n53 commonsourceibias.n52 0.189894
R679 commonsourceibias.n52 commonsourceibias.n15 0.189894
R680 commonsourceibias.n47 commonsourceibias.n15 0.189894
R681 commonsourceibias.n47 commonsourceibias.n46 0.189894
R682 commonsourceibias.n46 commonsourceibias.n45 0.189894
R683 commonsourceibias.n45 commonsourceibias.n18 0.189894
R684 commonsourceibias.n40 commonsourceibias.n18 0.189894
R685 commonsourceibias.n40 commonsourceibias.n39 0.189894
R686 commonsourceibias.n39 commonsourceibias.n20 0.189894
R687 commonsourceibias.n35 commonsourceibias.n20 0.189894
R688 commonsourceibias.n35 commonsourceibias.n34 0.189894
R689 commonsourceibias.n34 commonsourceibias.n22 0.189894
R690 commonsourceibias.n30 commonsourceibias.n22 0.189894
R691 commonsourceibias.n30 commonsourceibias.n29 0.189894
R692 commonsourceibias.n29 commonsourceibias.n24 0.189894
R693 commonsourceibias.n111 commonsourceibias.n84 0.189894
R694 commonsourceibias.n106 commonsourceibias.n84 0.189894
R695 commonsourceibias.n106 commonsourceibias.n105 0.189894
R696 commonsourceibias.n105 commonsourceibias.n86 0.189894
R697 commonsourceibias.n101 commonsourceibias.n86 0.189894
R698 commonsourceibias.n101 commonsourceibias.n100 0.189894
R699 commonsourceibias.n100 commonsourceibias.n88 0.189894
R700 commonsourceibias.n96 commonsourceibias.n88 0.189894
R701 commonsourceibias.n96 commonsourceibias.n95 0.189894
R702 commonsourceibias.n95 commonsourceibias.n90 0.189894
R703 commonsourceibias.n133 commonsourceibias.n0 0.189894
R704 commonsourceibias.n133 commonsourceibias.n132 0.189894
R705 commonsourceibias.n132 commonsourceibias.n2 0.189894
R706 commonsourceibias.n127 commonsourceibias.n2 0.189894
R707 commonsourceibias.n127 commonsourceibias.n126 0.189894
R708 commonsourceibias.n126 commonsourceibias.n125 0.189894
R709 commonsourceibias.n125 commonsourceibias.n4 0.189894
R710 commonsourceibias.n120 commonsourceibias.n4 0.189894
R711 commonsourceibias.n120 commonsourceibias.n119 0.189894
R712 commonsourceibias.n119 commonsourceibias.n118 0.189894
R713 commonsourceibias.n118 commonsourceibias.n6 0.189894
R714 commonsourceibias.n113 commonsourceibias.n6 0.189894
R715 commonsourceibias.n260 commonsourceibias.n202 0.189894
R716 commonsourceibias.n260 commonsourceibias.n259 0.189894
R717 commonsourceibias.n259 commonsourceibias.n204 0.189894
R718 commonsourceibias.n254 commonsourceibias.n204 0.189894
R719 commonsourceibias.n254 commonsourceibias.n253 0.189894
R720 commonsourceibias.n253 commonsourceibias.n252 0.189894
R721 commonsourceibias.n252 commonsourceibias.n206 0.189894
R722 commonsourceibias.n247 commonsourceibias.n206 0.189894
R723 commonsourceibias.n247 commonsourceibias.n246 0.189894
R724 commonsourceibias.n246 commonsourceibias.n245 0.189894
R725 commonsourceibias.n245 commonsourceibias.n208 0.189894
R726 commonsourceibias.n240 commonsourceibias.n208 0.189894
R727 commonsourceibias.n240 commonsourceibias.n239 0.189894
R728 commonsourceibias.n239 commonsourceibias.n238 0.189894
R729 commonsourceibias.n238 commonsourceibias.n211 0.189894
R730 commonsourceibias.n233 commonsourceibias.n211 0.189894
R731 commonsourceibias.n233 commonsourceibias.n232 0.189894
R732 commonsourceibias.n232 commonsourceibias.n213 0.189894
R733 commonsourceibias.n228 commonsourceibias.n213 0.189894
R734 commonsourceibias.n228 commonsourceibias.n227 0.189894
R735 commonsourceibias.n227 commonsourceibias.n215 0.189894
R736 commonsourceibias.n223 commonsourceibias.n215 0.189894
R737 commonsourceibias.n223 commonsourceibias.n222 0.189894
R738 commonsourceibias.n222 commonsourceibias.n217 0.189894
R739 commonsourceibias.n196 commonsourceibias.n138 0.189894
R740 commonsourceibias.n196 commonsourceibias.n195 0.189894
R741 commonsourceibias.n195 commonsourceibias.n140 0.189894
R742 commonsourceibias.n190 commonsourceibias.n140 0.189894
R743 commonsourceibias.n190 commonsourceibias.n189 0.189894
R744 commonsourceibias.n189 commonsourceibias.n188 0.189894
R745 commonsourceibias.n188 commonsourceibias.n142 0.189894
R746 commonsourceibias.n183 commonsourceibias.n142 0.189894
R747 commonsourceibias.n183 commonsourceibias.n182 0.189894
R748 commonsourceibias.n182 commonsourceibias.n181 0.189894
R749 commonsourceibias.n181 commonsourceibias.n144 0.189894
R750 commonsourceibias.n176 commonsourceibias.n144 0.189894
R751 commonsourceibias.n176 commonsourceibias.n175 0.189894
R752 commonsourceibias.n175 commonsourceibias.n174 0.189894
R753 commonsourceibias.n174 commonsourceibias.n147 0.189894
R754 commonsourceibias.n169 commonsourceibias.n147 0.189894
R755 commonsourceibias.n169 commonsourceibias.n168 0.189894
R756 commonsourceibias.n168 commonsourceibias.n149 0.189894
R757 commonsourceibias.n164 commonsourceibias.n149 0.189894
R758 commonsourceibias.n164 commonsourceibias.n163 0.189894
R759 commonsourceibias.n163 commonsourceibias.n151 0.189894
R760 commonsourceibias.n159 commonsourceibias.n151 0.189894
R761 commonsourceibias.n159 commonsourceibias.n158 0.189894
R762 commonsourceibias.n158 commonsourceibias.n153 0.189894
R763 commonsourceibias.n326 commonsourceibias.n321 0.189894
R764 commonsourceibias.n327 commonsourceibias.n326 0.189894
R765 commonsourceibias.n327 commonsourceibias.n319 0.189894
R766 commonsourceibias.n331 commonsourceibias.n319 0.189894
R767 commonsourceibias.n332 commonsourceibias.n331 0.189894
R768 commonsourceibias.n332 commonsourceibias.n317 0.189894
R769 commonsourceibias.n336 commonsourceibias.n317 0.189894
R770 commonsourceibias.n337 commonsourceibias.n336 0.189894
R771 commonsourceibias.n337 commonsourceibias.n315 0.189894
R772 commonsourceibias.n342 commonsourceibias.n315 0.189894
R773 commonsourceibias.n343 commonsourceibias.n342 0.189894
R774 commonsourceibias.n344 commonsourceibias.n343 0.189894
R775 commonsourceibias.n344 commonsourceibias.n313 0.189894
R776 commonsourceibias.n350 commonsourceibias.n313 0.189894
R777 commonsourceibias.n351 commonsourceibias.n350 0.189894
R778 commonsourceibias.n352 commonsourceibias.n351 0.189894
R779 commonsourceibias.n352 commonsourceibias.n311 0.189894
R780 commonsourceibias.n357 commonsourceibias.n311 0.189894
R781 commonsourceibias.n358 commonsourceibias.n357 0.189894
R782 commonsourceibias.n359 commonsourceibias.n358 0.189894
R783 commonsourceibias.n359 commonsourceibias.n309 0.189894
R784 commonsourceibias.n364 commonsourceibias.n309 0.189894
R785 commonsourceibias.n365 commonsourceibias.n364 0.189894
R786 commonsourceibias.n365 commonsourceibias.n307 0.189894
R787 commonsourceibias.n285 commonsourceibias.n280 0.189894
R788 commonsourceibias.n286 commonsourceibias.n285 0.189894
R789 commonsourceibias.n286 commonsourceibias.n278 0.189894
R790 commonsourceibias.n290 commonsourceibias.n278 0.189894
R791 commonsourceibias.n291 commonsourceibias.n290 0.189894
R792 commonsourceibias.n291 commonsourceibias.n276 0.189894
R793 commonsourceibias.n295 commonsourceibias.n276 0.189894
R794 commonsourceibias.n296 commonsourceibias.n295 0.189894
R795 commonsourceibias.n296 commonsourceibias.n274 0.189894
R796 commonsourceibias.n301 commonsourceibias.n274 0.189894
R797 commonsourceibias.n378 commonsourceibias.n272 0.189894
R798 commonsourceibias.n384 commonsourceibias.n272 0.189894
R799 commonsourceibias.n385 commonsourceibias.n384 0.189894
R800 commonsourceibias.n386 commonsourceibias.n385 0.189894
R801 commonsourceibias.n386 commonsourceibias.n270 0.189894
R802 commonsourceibias.n391 commonsourceibias.n270 0.189894
R803 commonsourceibias.n392 commonsourceibias.n391 0.189894
R804 commonsourceibias.n393 commonsourceibias.n392 0.189894
R805 commonsourceibias.n393 commonsourceibias.n268 0.189894
R806 commonsourceibias.n398 commonsourceibias.n268 0.189894
R807 commonsourceibias.n399 commonsourceibias.n398 0.189894
R808 commonsourceibias.n399 commonsourceibias.n266 0.189894
R809 commonsourceibias.n487 commonsourceibias.n482 0.189894
R810 commonsourceibias.n488 commonsourceibias.n487 0.189894
R811 commonsourceibias.n488 commonsourceibias.n480 0.189894
R812 commonsourceibias.n492 commonsourceibias.n480 0.189894
R813 commonsourceibias.n493 commonsourceibias.n492 0.189894
R814 commonsourceibias.n493 commonsourceibias.n478 0.189894
R815 commonsourceibias.n497 commonsourceibias.n478 0.189894
R816 commonsourceibias.n498 commonsourceibias.n497 0.189894
R817 commonsourceibias.n498 commonsourceibias.n476 0.189894
R818 commonsourceibias.n503 commonsourceibias.n476 0.189894
R819 commonsourceibias.n504 commonsourceibias.n503 0.189894
R820 commonsourceibias.n505 commonsourceibias.n504 0.189894
R821 commonsourceibias.n505 commonsourceibias.n474 0.189894
R822 commonsourceibias.n511 commonsourceibias.n474 0.189894
R823 commonsourceibias.n512 commonsourceibias.n511 0.189894
R824 commonsourceibias.n513 commonsourceibias.n512 0.189894
R825 commonsourceibias.n513 commonsourceibias.n472 0.189894
R826 commonsourceibias.n518 commonsourceibias.n472 0.189894
R827 commonsourceibias.n519 commonsourceibias.n518 0.189894
R828 commonsourceibias.n520 commonsourceibias.n519 0.189894
R829 commonsourceibias.n520 commonsourceibias.n470 0.189894
R830 commonsourceibias.n525 commonsourceibias.n470 0.189894
R831 commonsourceibias.n526 commonsourceibias.n525 0.189894
R832 commonsourceibias.n526 commonsourceibias.n468 0.189894
R833 commonsourceibias.n423 commonsourceibias.n418 0.189894
R834 commonsourceibias.n424 commonsourceibias.n423 0.189894
R835 commonsourceibias.n424 commonsourceibias.n416 0.189894
R836 commonsourceibias.n428 commonsourceibias.n416 0.189894
R837 commonsourceibias.n429 commonsourceibias.n428 0.189894
R838 commonsourceibias.n429 commonsourceibias.n414 0.189894
R839 commonsourceibias.n433 commonsourceibias.n414 0.189894
R840 commonsourceibias.n434 commonsourceibias.n433 0.189894
R841 commonsourceibias.n434 commonsourceibias.n412 0.189894
R842 commonsourceibias.n439 commonsourceibias.n412 0.189894
R843 commonsourceibias.n440 commonsourceibias.n439 0.189894
R844 commonsourceibias.n441 commonsourceibias.n440 0.189894
R845 commonsourceibias.n441 commonsourceibias.n410 0.189894
R846 commonsourceibias.n447 commonsourceibias.n410 0.189894
R847 commonsourceibias.n448 commonsourceibias.n447 0.189894
R848 commonsourceibias.n449 commonsourceibias.n448 0.189894
R849 commonsourceibias.n449 commonsourceibias.n408 0.189894
R850 commonsourceibias.n454 commonsourceibias.n408 0.189894
R851 commonsourceibias.n455 commonsourceibias.n454 0.189894
R852 commonsourceibias.n456 commonsourceibias.n455 0.189894
R853 commonsourceibias.n456 commonsourceibias.n406 0.189894
R854 commonsourceibias.n461 commonsourceibias.n406 0.189894
R855 commonsourceibias.n462 commonsourceibias.n461 0.189894
R856 commonsourceibias.n462 commonsourceibias.n404 0.189894
R857 commonsourceibias.n112 commonsourceibias.n111 0.170955
R858 commonsourceibias.n113 commonsourceibias.n112 0.170955
R859 commonsourceibias.n377 commonsourceibias.n301 0.170955
R860 commonsourceibias.n378 commonsourceibias.n377 0.170955
R861 gnd.n6566 gnd.n310 1552.66
R862 gnd.n3667 gnd.n3666 939.716
R863 gnd.n7146 gnd.n171 838.452
R864 gnd.n7088 gnd.n169 838.452
R865 gnd.n1485 gnd.n1373 838.452
R866 gnd.n5375 gnd.n1487 838.452
R867 gnd.n5884 gnd.n863 838.452
R868 gnd.n5804 gnd.n861 838.452
R869 gnd.n3735 gnd.n3669 838.452
R870 gnd.n3962 gnd.n2204 838.452
R871 gnd.n7148 gnd.n166 783.196
R872 gnd.n6963 gnd.n168 783.196
R873 gnd.n5378 gnd.n5377 783.196
R874 gnd.n5495 gnd.n1419 783.196
R875 gnd.n5886 gnd.n858 783.196
R876 gnd.n1069 gnd.n860 783.196
R877 gnd.n3841 gnd.n3668 783.196
R878 gnd.n3960 gnd.n3745 783.196
R879 gnd.n3574 gnd.n2206 766.379
R880 gnd.n3577 gnd.n3576 766.379
R881 gnd.n2816 gnd.n2719 766.379
R882 gnd.n2812 gnd.n2717 766.379
R883 gnd.n3665 gnd.n2228 756.769
R884 gnd.n3568 gnd.n3567 756.769
R885 gnd.n2909 gnd.n2626 756.769
R886 gnd.n2907 gnd.n2629 756.769
R887 gnd.n6144 gnd.n562 756.769
R888 gnd.n6565 gnd.n311 756.769
R889 gnd.n6777 gnd.n6776 756.769
R890 gnd.n5968 gnd.n727 756.769
R891 gnd.n5865 gnd.n893 711.122
R892 gnd.n5564 gnd.n1309 711.122
R893 gnd.n5869 gnd.n875 711.122
R894 gnd.n5566 gnd.n1304 711.122
R895 gnd.n6140 gnd.n562 585
R896 gnd.n562 gnd.n561 585
R897 gnd.n6139 gnd.n6138 585
R898 gnd.n6138 gnd.n6137 585
R899 gnd.n565 gnd.n564 585
R900 gnd.n6136 gnd.n565 585
R901 gnd.n6134 gnd.n6133 585
R902 gnd.n6135 gnd.n6134 585
R903 gnd.n6132 gnd.n567 585
R904 gnd.n567 gnd.n566 585
R905 gnd.n6131 gnd.n6130 585
R906 gnd.n6130 gnd.n6129 585
R907 gnd.n573 gnd.n572 585
R908 gnd.n6128 gnd.n573 585
R909 gnd.n6126 gnd.n6125 585
R910 gnd.n6127 gnd.n6126 585
R911 gnd.n6124 gnd.n575 585
R912 gnd.n575 gnd.n574 585
R913 gnd.n6123 gnd.n6122 585
R914 gnd.n6122 gnd.n6121 585
R915 gnd.n581 gnd.n580 585
R916 gnd.n6120 gnd.n581 585
R917 gnd.n6118 gnd.n6117 585
R918 gnd.n6119 gnd.n6118 585
R919 gnd.n6116 gnd.n583 585
R920 gnd.n583 gnd.n582 585
R921 gnd.n6115 gnd.n6114 585
R922 gnd.n6114 gnd.n6113 585
R923 gnd.n589 gnd.n588 585
R924 gnd.n6112 gnd.n589 585
R925 gnd.n6110 gnd.n6109 585
R926 gnd.n6111 gnd.n6110 585
R927 gnd.n6108 gnd.n591 585
R928 gnd.n591 gnd.n590 585
R929 gnd.n6107 gnd.n6106 585
R930 gnd.n6106 gnd.n6105 585
R931 gnd.n597 gnd.n596 585
R932 gnd.n6104 gnd.n597 585
R933 gnd.n6102 gnd.n6101 585
R934 gnd.n6103 gnd.n6102 585
R935 gnd.n6100 gnd.n599 585
R936 gnd.n599 gnd.n598 585
R937 gnd.n6099 gnd.n6098 585
R938 gnd.n6098 gnd.n6097 585
R939 gnd.n605 gnd.n604 585
R940 gnd.n6096 gnd.n605 585
R941 gnd.n6094 gnd.n6093 585
R942 gnd.n6095 gnd.n6094 585
R943 gnd.n6092 gnd.n607 585
R944 gnd.n607 gnd.n606 585
R945 gnd.n6091 gnd.n6090 585
R946 gnd.n6090 gnd.n6089 585
R947 gnd.n613 gnd.n612 585
R948 gnd.n6088 gnd.n613 585
R949 gnd.n6086 gnd.n6085 585
R950 gnd.n6087 gnd.n6086 585
R951 gnd.n6084 gnd.n615 585
R952 gnd.n615 gnd.n614 585
R953 gnd.n6083 gnd.n6082 585
R954 gnd.n6082 gnd.n6081 585
R955 gnd.n621 gnd.n620 585
R956 gnd.n6080 gnd.n621 585
R957 gnd.n6078 gnd.n6077 585
R958 gnd.n6079 gnd.n6078 585
R959 gnd.n6076 gnd.n623 585
R960 gnd.n623 gnd.n622 585
R961 gnd.n6075 gnd.n6074 585
R962 gnd.n6074 gnd.n6073 585
R963 gnd.n629 gnd.n628 585
R964 gnd.n6072 gnd.n629 585
R965 gnd.n6070 gnd.n6069 585
R966 gnd.n6071 gnd.n6070 585
R967 gnd.n6068 gnd.n631 585
R968 gnd.n631 gnd.n630 585
R969 gnd.n6067 gnd.n6066 585
R970 gnd.n6066 gnd.n6065 585
R971 gnd.n637 gnd.n636 585
R972 gnd.n6064 gnd.n637 585
R973 gnd.n6062 gnd.n6061 585
R974 gnd.n6063 gnd.n6062 585
R975 gnd.n6060 gnd.n639 585
R976 gnd.n639 gnd.n638 585
R977 gnd.n6059 gnd.n6058 585
R978 gnd.n6058 gnd.n6057 585
R979 gnd.n645 gnd.n644 585
R980 gnd.n6056 gnd.n645 585
R981 gnd.n6054 gnd.n6053 585
R982 gnd.n6055 gnd.n6054 585
R983 gnd.n6052 gnd.n647 585
R984 gnd.n647 gnd.n646 585
R985 gnd.n6051 gnd.n6050 585
R986 gnd.n6050 gnd.n6049 585
R987 gnd.n653 gnd.n652 585
R988 gnd.n6048 gnd.n653 585
R989 gnd.n6046 gnd.n6045 585
R990 gnd.n6047 gnd.n6046 585
R991 gnd.n6044 gnd.n655 585
R992 gnd.n655 gnd.n654 585
R993 gnd.n6043 gnd.n6042 585
R994 gnd.n6042 gnd.n6041 585
R995 gnd.n661 gnd.n660 585
R996 gnd.n6040 gnd.n661 585
R997 gnd.n6038 gnd.n6037 585
R998 gnd.n6039 gnd.n6038 585
R999 gnd.n6036 gnd.n663 585
R1000 gnd.n663 gnd.n662 585
R1001 gnd.n6035 gnd.n6034 585
R1002 gnd.n6034 gnd.n6033 585
R1003 gnd.n669 gnd.n668 585
R1004 gnd.n6032 gnd.n669 585
R1005 gnd.n6030 gnd.n6029 585
R1006 gnd.n6031 gnd.n6030 585
R1007 gnd.n6028 gnd.n671 585
R1008 gnd.n671 gnd.n670 585
R1009 gnd.n6027 gnd.n6026 585
R1010 gnd.n6026 gnd.n6025 585
R1011 gnd.n677 gnd.n676 585
R1012 gnd.n6024 gnd.n677 585
R1013 gnd.n6022 gnd.n6021 585
R1014 gnd.n6023 gnd.n6022 585
R1015 gnd.n6020 gnd.n679 585
R1016 gnd.n679 gnd.n678 585
R1017 gnd.n6019 gnd.n6018 585
R1018 gnd.n6018 gnd.n6017 585
R1019 gnd.n685 gnd.n684 585
R1020 gnd.n6016 gnd.n685 585
R1021 gnd.n6014 gnd.n6013 585
R1022 gnd.n6015 gnd.n6014 585
R1023 gnd.n6012 gnd.n687 585
R1024 gnd.n687 gnd.n686 585
R1025 gnd.n6011 gnd.n6010 585
R1026 gnd.n6010 gnd.n6009 585
R1027 gnd.n693 gnd.n692 585
R1028 gnd.n6008 gnd.n693 585
R1029 gnd.n6006 gnd.n6005 585
R1030 gnd.n6007 gnd.n6006 585
R1031 gnd.n6004 gnd.n695 585
R1032 gnd.n695 gnd.n694 585
R1033 gnd.n6003 gnd.n6002 585
R1034 gnd.n6002 gnd.n6001 585
R1035 gnd.n701 gnd.n700 585
R1036 gnd.n6000 gnd.n701 585
R1037 gnd.n5998 gnd.n5997 585
R1038 gnd.n5999 gnd.n5998 585
R1039 gnd.n5996 gnd.n703 585
R1040 gnd.n703 gnd.n702 585
R1041 gnd.n5995 gnd.n5994 585
R1042 gnd.n5994 gnd.n5993 585
R1043 gnd.n709 gnd.n708 585
R1044 gnd.n5992 gnd.n709 585
R1045 gnd.n5990 gnd.n5989 585
R1046 gnd.n5991 gnd.n5990 585
R1047 gnd.n5988 gnd.n711 585
R1048 gnd.n711 gnd.n710 585
R1049 gnd.n5987 gnd.n5986 585
R1050 gnd.n5986 gnd.n5985 585
R1051 gnd.n717 gnd.n716 585
R1052 gnd.n5984 gnd.n717 585
R1053 gnd.n5982 gnd.n5981 585
R1054 gnd.n5983 gnd.n5982 585
R1055 gnd.n5980 gnd.n719 585
R1056 gnd.n719 gnd.n718 585
R1057 gnd.n5979 gnd.n5978 585
R1058 gnd.n5978 gnd.n5977 585
R1059 gnd.n725 gnd.n724 585
R1060 gnd.n5976 gnd.n725 585
R1061 gnd.n5974 gnd.n5973 585
R1062 gnd.n5975 gnd.n5974 585
R1063 gnd.n6144 gnd.n6143 585
R1064 gnd.n6145 gnd.n6144 585
R1065 gnd.n560 gnd.n559 585
R1066 gnd.n6146 gnd.n560 585
R1067 gnd.n6149 gnd.n6148 585
R1068 gnd.n6148 gnd.n6147 585
R1069 gnd.n557 gnd.n556 585
R1070 gnd.n556 gnd.n555 585
R1071 gnd.n6154 gnd.n6153 585
R1072 gnd.n6155 gnd.n6154 585
R1073 gnd.n554 gnd.n553 585
R1074 gnd.n6156 gnd.n554 585
R1075 gnd.n6159 gnd.n6158 585
R1076 gnd.n6158 gnd.n6157 585
R1077 gnd.n551 gnd.n550 585
R1078 gnd.n550 gnd.n549 585
R1079 gnd.n6164 gnd.n6163 585
R1080 gnd.n6165 gnd.n6164 585
R1081 gnd.n548 gnd.n547 585
R1082 gnd.n6166 gnd.n548 585
R1083 gnd.n6169 gnd.n6168 585
R1084 gnd.n6168 gnd.n6167 585
R1085 gnd.n545 gnd.n544 585
R1086 gnd.n544 gnd.n543 585
R1087 gnd.n6174 gnd.n6173 585
R1088 gnd.n6175 gnd.n6174 585
R1089 gnd.n542 gnd.n541 585
R1090 gnd.n6176 gnd.n542 585
R1091 gnd.n6179 gnd.n6178 585
R1092 gnd.n6178 gnd.n6177 585
R1093 gnd.n539 gnd.n538 585
R1094 gnd.n538 gnd.n537 585
R1095 gnd.n6184 gnd.n6183 585
R1096 gnd.n6185 gnd.n6184 585
R1097 gnd.n536 gnd.n535 585
R1098 gnd.n6186 gnd.n536 585
R1099 gnd.n6189 gnd.n6188 585
R1100 gnd.n6188 gnd.n6187 585
R1101 gnd.n533 gnd.n532 585
R1102 gnd.n532 gnd.n531 585
R1103 gnd.n6194 gnd.n6193 585
R1104 gnd.n6195 gnd.n6194 585
R1105 gnd.n530 gnd.n529 585
R1106 gnd.n6196 gnd.n530 585
R1107 gnd.n6199 gnd.n6198 585
R1108 gnd.n6198 gnd.n6197 585
R1109 gnd.n527 gnd.n526 585
R1110 gnd.n526 gnd.n525 585
R1111 gnd.n6204 gnd.n6203 585
R1112 gnd.n6205 gnd.n6204 585
R1113 gnd.n524 gnd.n523 585
R1114 gnd.n6206 gnd.n524 585
R1115 gnd.n6209 gnd.n6208 585
R1116 gnd.n6208 gnd.n6207 585
R1117 gnd.n521 gnd.n520 585
R1118 gnd.n520 gnd.n519 585
R1119 gnd.n6214 gnd.n6213 585
R1120 gnd.n6215 gnd.n6214 585
R1121 gnd.n518 gnd.n517 585
R1122 gnd.n6216 gnd.n518 585
R1123 gnd.n6219 gnd.n6218 585
R1124 gnd.n6218 gnd.n6217 585
R1125 gnd.n515 gnd.n514 585
R1126 gnd.n514 gnd.n513 585
R1127 gnd.n6224 gnd.n6223 585
R1128 gnd.n6225 gnd.n6224 585
R1129 gnd.n512 gnd.n511 585
R1130 gnd.n6226 gnd.n512 585
R1131 gnd.n6229 gnd.n6228 585
R1132 gnd.n6228 gnd.n6227 585
R1133 gnd.n509 gnd.n508 585
R1134 gnd.n508 gnd.n507 585
R1135 gnd.n6234 gnd.n6233 585
R1136 gnd.n6235 gnd.n6234 585
R1137 gnd.n506 gnd.n505 585
R1138 gnd.n6236 gnd.n506 585
R1139 gnd.n6239 gnd.n6238 585
R1140 gnd.n6238 gnd.n6237 585
R1141 gnd.n503 gnd.n502 585
R1142 gnd.n502 gnd.n501 585
R1143 gnd.n6244 gnd.n6243 585
R1144 gnd.n6245 gnd.n6244 585
R1145 gnd.n500 gnd.n499 585
R1146 gnd.n6246 gnd.n500 585
R1147 gnd.n6249 gnd.n6248 585
R1148 gnd.n6248 gnd.n6247 585
R1149 gnd.n497 gnd.n496 585
R1150 gnd.n496 gnd.n495 585
R1151 gnd.n6254 gnd.n6253 585
R1152 gnd.n6255 gnd.n6254 585
R1153 gnd.n494 gnd.n493 585
R1154 gnd.n6256 gnd.n494 585
R1155 gnd.n6259 gnd.n6258 585
R1156 gnd.n6258 gnd.n6257 585
R1157 gnd.n491 gnd.n490 585
R1158 gnd.n490 gnd.n489 585
R1159 gnd.n6264 gnd.n6263 585
R1160 gnd.n6265 gnd.n6264 585
R1161 gnd.n488 gnd.n487 585
R1162 gnd.n6266 gnd.n488 585
R1163 gnd.n6269 gnd.n6268 585
R1164 gnd.n6268 gnd.n6267 585
R1165 gnd.n485 gnd.n484 585
R1166 gnd.n484 gnd.n483 585
R1167 gnd.n6274 gnd.n6273 585
R1168 gnd.n6275 gnd.n6274 585
R1169 gnd.n482 gnd.n481 585
R1170 gnd.n6276 gnd.n482 585
R1171 gnd.n6279 gnd.n6278 585
R1172 gnd.n6278 gnd.n6277 585
R1173 gnd.n479 gnd.n478 585
R1174 gnd.n478 gnd.n477 585
R1175 gnd.n6284 gnd.n6283 585
R1176 gnd.n6285 gnd.n6284 585
R1177 gnd.n476 gnd.n475 585
R1178 gnd.n6286 gnd.n476 585
R1179 gnd.n6289 gnd.n6288 585
R1180 gnd.n6288 gnd.n6287 585
R1181 gnd.n473 gnd.n472 585
R1182 gnd.n472 gnd.n471 585
R1183 gnd.n6294 gnd.n6293 585
R1184 gnd.n6295 gnd.n6294 585
R1185 gnd.n470 gnd.n469 585
R1186 gnd.n6296 gnd.n470 585
R1187 gnd.n6299 gnd.n6298 585
R1188 gnd.n6298 gnd.n6297 585
R1189 gnd.n467 gnd.n466 585
R1190 gnd.n466 gnd.n465 585
R1191 gnd.n6304 gnd.n6303 585
R1192 gnd.n6305 gnd.n6304 585
R1193 gnd.n464 gnd.n463 585
R1194 gnd.n6306 gnd.n464 585
R1195 gnd.n6309 gnd.n6308 585
R1196 gnd.n6308 gnd.n6307 585
R1197 gnd.n461 gnd.n460 585
R1198 gnd.n460 gnd.n459 585
R1199 gnd.n6314 gnd.n6313 585
R1200 gnd.n6315 gnd.n6314 585
R1201 gnd.n458 gnd.n457 585
R1202 gnd.n6316 gnd.n458 585
R1203 gnd.n6319 gnd.n6318 585
R1204 gnd.n6318 gnd.n6317 585
R1205 gnd.n455 gnd.n454 585
R1206 gnd.n454 gnd.n453 585
R1207 gnd.n6324 gnd.n6323 585
R1208 gnd.n6325 gnd.n6324 585
R1209 gnd.n452 gnd.n451 585
R1210 gnd.n6326 gnd.n452 585
R1211 gnd.n6329 gnd.n6328 585
R1212 gnd.n6328 gnd.n6327 585
R1213 gnd.n449 gnd.n448 585
R1214 gnd.n448 gnd.n447 585
R1215 gnd.n6334 gnd.n6333 585
R1216 gnd.n6335 gnd.n6334 585
R1217 gnd.n446 gnd.n445 585
R1218 gnd.n6336 gnd.n446 585
R1219 gnd.n6339 gnd.n6338 585
R1220 gnd.n6338 gnd.n6337 585
R1221 gnd.n443 gnd.n442 585
R1222 gnd.n442 gnd.n441 585
R1223 gnd.n6344 gnd.n6343 585
R1224 gnd.n6345 gnd.n6344 585
R1225 gnd.n440 gnd.n439 585
R1226 gnd.n6346 gnd.n440 585
R1227 gnd.n6349 gnd.n6348 585
R1228 gnd.n6348 gnd.n6347 585
R1229 gnd.n437 gnd.n436 585
R1230 gnd.n436 gnd.n435 585
R1231 gnd.n6354 gnd.n6353 585
R1232 gnd.n6355 gnd.n6354 585
R1233 gnd.n434 gnd.n433 585
R1234 gnd.n6356 gnd.n434 585
R1235 gnd.n6359 gnd.n6358 585
R1236 gnd.n6358 gnd.n6357 585
R1237 gnd.n431 gnd.n430 585
R1238 gnd.n430 gnd.n429 585
R1239 gnd.n6364 gnd.n6363 585
R1240 gnd.n6365 gnd.n6364 585
R1241 gnd.n428 gnd.n427 585
R1242 gnd.n6366 gnd.n428 585
R1243 gnd.n6369 gnd.n6368 585
R1244 gnd.n6368 gnd.n6367 585
R1245 gnd.n425 gnd.n424 585
R1246 gnd.n424 gnd.n423 585
R1247 gnd.n6374 gnd.n6373 585
R1248 gnd.n6375 gnd.n6374 585
R1249 gnd.n422 gnd.n421 585
R1250 gnd.n6376 gnd.n422 585
R1251 gnd.n6379 gnd.n6378 585
R1252 gnd.n6378 gnd.n6377 585
R1253 gnd.n419 gnd.n418 585
R1254 gnd.n418 gnd.n417 585
R1255 gnd.n6384 gnd.n6383 585
R1256 gnd.n6385 gnd.n6384 585
R1257 gnd.n416 gnd.n415 585
R1258 gnd.n6386 gnd.n416 585
R1259 gnd.n6389 gnd.n6388 585
R1260 gnd.n6388 gnd.n6387 585
R1261 gnd.n413 gnd.n412 585
R1262 gnd.n412 gnd.n411 585
R1263 gnd.n6394 gnd.n6393 585
R1264 gnd.n6395 gnd.n6394 585
R1265 gnd.n410 gnd.n409 585
R1266 gnd.n6396 gnd.n410 585
R1267 gnd.n6399 gnd.n6398 585
R1268 gnd.n6398 gnd.n6397 585
R1269 gnd.n407 gnd.n406 585
R1270 gnd.n406 gnd.n405 585
R1271 gnd.n6404 gnd.n6403 585
R1272 gnd.n6405 gnd.n6404 585
R1273 gnd.n404 gnd.n403 585
R1274 gnd.n6406 gnd.n404 585
R1275 gnd.n6409 gnd.n6408 585
R1276 gnd.n6408 gnd.n6407 585
R1277 gnd.n401 gnd.n400 585
R1278 gnd.n400 gnd.n399 585
R1279 gnd.n6414 gnd.n6413 585
R1280 gnd.n6415 gnd.n6414 585
R1281 gnd.n398 gnd.n397 585
R1282 gnd.n6416 gnd.n398 585
R1283 gnd.n6419 gnd.n6418 585
R1284 gnd.n6418 gnd.n6417 585
R1285 gnd.n395 gnd.n394 585
R1286 gnd.n394 gnd.n393 585
R1287 gnd.n6424 gnd.n6423 585
R1288 gnd.n6425 gnd.n6424 585
R1289 gnd.n392 gnd.n391 585
R1290 gnd.n6426 gnd.n392 585
R1291 gnd.n6429 gnd.n6428 585
R1292 gnd.n6428 gnd.n6427 585
R1293 gnd.n389 gnd.n388 585
R1294 gnd.n388 gnd.n387 585
R1295 gnd.n6434 gnd.n6433 585
R1296 gnd.n6435 gnd.n6434 585
R1297 gnd.n386 gnd.n385 585
R1298 gnd.n6436 gnd.n386 585
R1299 gnd.n6439 gnd.n6438 585
R1300 gnd.n6438 gnd.n6437 585
R1301 gnd.n383 gnd.n382 585
R1302 gnd.n382 gnd.n381 585
R1303 gnd.n6444 gnd.n6443 585
R1304 gnd.n6445 gnd.n6444 585
R1305 gnd.n380 gnd.n379 585
R1306 gnd.n6446 gnd.n380 585
R1307 gnd.n6449 gnd.n6448 585
R1308 gnd.n6448 gnd.n6447 585
R1309 gnd.n377 gnd.n376 585
R1310 gnd.n376 gnd.n375 585
R1311 gnd.n6454 gnd.n6453 585
R1312 gnd.n6455 gnd.n6454 585
R1313 gnd.n374 gnd.n373 585
R1314 gnd.n6456 gnd.n374 585
R1315 gnd.n6459 gnd.n6458 585
R1316 gnd.n6458 gnd.n6457 585
R1317 gnd.n371 gnd.n370 585
R1318 gnd.n370 gnd.n369 585
R1319 gnd.n6464 gnd.n6463 585
R1320 gnd.n6465 gnd.n6464 585
R1321 gnd.n368 gnd.n367 585
R1322 gnd.n6466 gnd.n368 585
R1323 gnd.n6469 gnd.n6468 585
R1324 gnd.n6468 gnd.n6467 585
R1325 gnd.n365 gnd.n364 585
R1326 gnd.n364 gnd.n363 585
R1327 gnd.n6474 gnd.n6473 585
R1328 gnd.n6475 gnd.n6474 585
R1329 gnd.n362 gnd.n361 585
R1330 gnd.n6476 gnd.n362 585
R1331 gnd.n6479 gnd.n6478 585
R1332 gnd.n6478 gnd.n6477 585
R1333 gnd.n359 gnd.n358 585
R1334 gnd.n358 gnd.n357 585
R1335 gnd.n6484 gnd.n6483 585
R1336 gnd.n6485 gnd.n6484 585
R1337 gnd.n356 gnd.n355 585
R1338 gnd.n6486 gnd.n356 585
R1339 gnd.n6489 gnd.n6488 585
R1340 gnd.n6488 gnd.n6487 585
R1341 gnd.n353 gnd.n352 585
R1342 gnd.n352 gnd.n351 585
R1343 gnd.n6494 gnd.n6493 585
R1344 gnd.n6495 gnd.n6494 585
R1345 gnd.n350 gnd.n349 585
R1346 gnd.n6496 gnd.n350 585
R1347 gnd.n6499 gnd.n6498 585
R1348 gnd.n6498 gnd.n6497 585
R1349 gnd.n347 gnd.n346 585
R1350 gnd.n346 gnd.n345 585
R1351 gnd.n6504 gnd.n6503 585
R1352 gnd.n6505 gnd.n6504 585
R1353 gnd.n344 gnd.n343 585
R1354 gnd.n6506 gnd.n344 585
R1355 gnd.n6509 gnd.n6508 585
R1356 gnd.n6508 gnd.n6507 585
R1357 gnd.n341 gnd.n340 585
R1358 gnd.n340 gnd.n339 585
R1359 gnd.n6514 gnd.n6513 585
R1360 gnd.n6515 gnd.n6514 585
R1361 gnd.n338 gnd.n337 585
R1362 gnd.n6516 gnd.n338 585
R1363 gnd.n6519 gnd.n6518 585
R1364 gnd.n6518 gnd.n6517 585
R1365 gnd.n335 gnd.n334 585
R1366 gnd.n334 gnd.n333 585
R1367 gnd.n6524 gnd.n6523 585
R1368 gnd.n6525 gnd.n6524 585
R1369 gnd.n332 gnd.n331 585
R1370 gnd.n6526 gnd.n332 585
R1371 gnd.n6529 gnd.n6528 585
R1372 gnd.n6528 gnd.n6527 585
R1373 gnd.n329 gnd.n328 585
R1374 gnd.n328 gnd.n327 585
R1375 gnd.n6534 gnd.n6533 585
R1376 gnd.n6535 gnd.n6534 585
R1377 gnd.n326 gnd.n325 585
R1378 gnd.n6536 gnd.n326 585
R1379 gnd.n6539 gnd.n6538 585
R1380 gnd.n6538 gnd.n6537 585
R1381 gnd.n323 gnd.n322 585
R1382 gnd.n322 gnd.n321 585
R1383 gnd.n6544 gnd.n6543 585
R1384 gnd.n6545 gnd.n6544 585
R1385 gnd.n320 gnd.n319 585
R1386 gnd.n6546 gnd.n320 585
R1387 gnd.n6549 gnd.n6548 585
R1388 gnd.n6548 gnd.n6547 585
R1389 gnd.n317 gnd.n316 585
R1390 gnd.n316 gnd.n315 585
R1391 gnd.n6555 gnd.n6554 585
R1392 gnd.n6556 gnd.n6555 585
R1393 gnd.n314 gnd.n313 585
R1394 gnd.n6557 gnd.n314 585
R1395 gnd.n6560 gnd.n6559 585
R1396 gnd.n6559 gnd.n6558 585
R1397 gnd.n6561 gnd.n311 585
R1398 gnd.n311 gnd.n310 585
R1399 gnd.n186 gnd.n185 585
R1400 gnd.n6768 gnd.n185 585
R1401 gnd.n6771 gnd.n6770 585
R1402 gnd.n6770 gnd.n6769 585
R1403 gnd.n189 gnd.n188 585
R1404 gnd.n6767 gnd.n189 585
R1405 gnd.n6765 gnd.n6764 585
R1406 gnd.n6766 gnd.n6765 585
R1407 gnd.n192 gnd.n191 585
R1408 gnd.n191 gnd.n190 585
R1409 gnd.n6760 gnd.n6759 585
R1410 gnd.n6759 gnd.n6758 585
R1411 gnd.n195 gnd.n194 585
R1412 gnd.n6757 gnd.n195 585
R1413 gnd.n6755 gnd.n6754 585
R1414 gnd.n6756 gnd.n6755 585
R1415 gnd.n198 gnd.n197 585
R1416 gnd.n197 gnd.n196 585
R1417 gnd.n6750 gnd.n6749 585
R1418 gnd.n6749 gnd.n6748 585
R1419 gnd.n201 gnd.n200 585
R1420 gnd.n6747 gnd.n201 585
R1421 gnd.n6745 gnd.n6744 585
R1422 gnd.n6746 gnd.n6745 585
R1423 gnd.n204 gnd.n203 585
R1424 gnd.n203 gnd.n202 585
R1425 gnd.n6740 gnd.n6739 585
R1426 gnd.n6739 gnd.n6738 585
R1427 gnd.n207 gnd.n206 585
R1428 gnd.n6737 gnd.n207 585
R1429 gnd.n6735 gnd.n6734 585
R1430 gnd.n6736 gnd.n6735 585
R1431 gnd.n210 gnd.n209 585
R1432 gnd.n209 gnd.n208 585
R1433 gnd.n6730 gnd.n6729 585
R1434 gnd.n6729 gnd.n6728 585
R1435 gnd.n213 gnd.n212 585
R1436 gnd.n6727 gnd.n213 585
R1437 gnd.n6725 gnd.n6724 585
R1438 gnd.n6726 gnd.n6725 585
R1439 gnd.n216 gnd.n215 585
R1440 gnd.n215 gnd.n214 585
R1441 gnd.n6720 gnd.n6719 585
R1442 gnd.n6719 gnd.n6718 585
R1443 gnd.n219 gnd.n218 585
R1444 gnd.n6717 gnd.n219 585
R1445 gnd.n6715 gnd.n6714 585
R1446 gnd.n6716 gnd.n6715 585
R1447 gnd.n222 gnd.n221 585
R1448 gnd.n221 gnd.n220 585
R1449 gnd.n6710 gnd.n6709 585
R1450 gnd.n6709 gnd.n6708 585
R1451 gnd.n225 gnd.n224 585
R1452 gnd.n6707 gnd.n225 585
R1453 gnd.n6705 gnd.n6704 585
R1454 gnd.n6706 gnd.n6705 585
R1455 gnd.n228 gnd.n227 585
R1456 gnd.n227 gnd.n226 585
R1457 gnd.n6700 gnd.n6699 585
R1458 gnd.n6699 gnd.n6698 585
R1459 gnd.n231 gnd.n230 585
R1460 gnd.n6697 gnd.n231 585
R1461 gnd.n6695 gnd.n6694 585
R1462 gnd.n6696 gnd.n6695 585
R1463 gnd.n234 gnd.n233 585
R1464 gnd.n233 gnd.n232 585
R1465 gnd.n6690 gnd.n6689 585
R1466 gnd.n6689 gnd.n6688 585
R1467 gnd.n237 gnd.n236 585
R1468 gnd.n6687 gnd.n237 585
R1469 gnd.n6685 gnd.n6684 585
R1470 gnd.n6686 gnd.n6685 585
R1471 gnd.n240 gnd.n239 585
R1472 gnd.n239 gnd.n238 585
R1473 gnd.n6680 gnd.n6679 585
R1474 gnd.n6679 gnd.n6678 585
R1475 gnd.n243 gnd.n242 585
R1476 gnd.n6677 gnd.n243 585
R1477 gnd.n6675 gnd.n6674 585
R1478 gnd.n6676 gnd.n6675 585
R1479 gnd.n246 gnd.n245 585
R1480 gnd.n245 gnd.n244 585
R1481 gnd.n6670 gnd.n6669 585
R1482 gnd.n6669 gnd.n6668 585
R1483 gnd.n249 gnd.n248 585
R1484 gnd.n6667 gnd.n249 585
R1485 gnd.n6665 gnd.n6664 585
R1486 gnd.n6666 gnd.n6665 585
R1487 gnd.n252 gnd.n251 585
R1488 gnd.n251 gnd.n250 585
R1489 gnd.n6660 gnd.n6659 585
R1490 gnd.n6659 gnd.n6658 585
R1491 gnd.n255 gnd.n254 585
R1492 gnd.n6657 gnd.n255 585
R1493 gnd.n6655 gnd.n6654 585
R1494 gnd.n6656 gnd.n6655 585
R1495 gnd.n258 gnd.n257 585
R1496 gnd.n257 gnd.n256 585
R1497 gnd.n6650 gnd.n6649 585
R1498 gnd.n6649 gnd.n6648 585
R1499 gnd.n261 gnd.n260 585
R1500 gnd.n6647 gnd.n261 585
R1501 gnd.n6645 gnd.n6644 585
R1502 gnd.n6646 gnd.n6645 585
R1503 gnd.n264 gnd.n263 585
R1504 gnd.n263 gnd.n262 585
R1505 gnd.n6640 gnd.n6639 585
R1506 gnd.n6639 gnd.n6638 585
R1507 gnd.n267 gnd.n266 585
R1508 gnd.n6637 gnd.n267 585
R1509 gnd.n6635 gnd.n6634 585
R1510 gnd.n6636 gnd.n6635 585
R1511 gnd.n270 gnd.n269 585
R1512 gnd.n269 gnd.n268 585
R1513 gnd.n6630 gnd.n6629 585
R1514 gnd.n6629 gnd.n6628 585
R1515 gnd.n273 gnd.n272 585
R1516 gnd.n6627 gnd.n273 585
R1517 gnd.n6625 gnd.n6624 585
R1518 gnd.n6626 gnd.n6625 585
R1519 gnd.n276 gnd.n275 585
R1520 gnd.n275 gnd.n274 585
R1521 gnd.n6620 gnd.n6619 585
R1522 gnd.n6619 gnd.n6618 585
R1523 gnd.n279 gnd.n278 585
R1524 gnd.n6617 gnd.n279 585
R1525 gnd.n6615 gnd.n6614 585
R1526 gnd.n6616 gnd.n6615 585
R1527 gnd.n282 gnd.n281 585
R1528 gnd.n281 gnd.n280 585
R1529 gnd.n6610 gnd.n6609 585
R1530 gnd.n6609 gnd.n6608 585
R1531 gnd.n285 gnd.n284 585
R1532 gnd.n6607 gnd.n285 585
R1533 gnd.n6605 gnd.n6604 585
R1534 gnd.n6606 gnd.n6605 585
R1535 gnd.n288 gnd.n287 585
R1536 gnd.n287 gnd.n286 585
R1537 gnd.n6600 gnd.n6599 585
R1538 gnd.n6599 gnd.n6598 585
R1539 gnd.n291 gnd.n290 585
R1540 gnd.n6597 gnd.n291 585
R1541 gnd.n6595 gnd.n6594 585
R1542 gnd.n6596 gnd.n6595 585
R1543 gnd.n294 gnd.n293 585
R1544 gnd.n293 gnd.n292 585
R1545 gnd.n6590 gnd.n6589 585
R1546 gnd.n6589 gnd.n6588 585
R1547 gnd.n297 gnd.n296 585
R1548 gnd.n6587 gnd.n297 585
R1549 gnd.n6585 gnd.n6584 585
R1550 gnd.n6586 gnd.n6585 585
R1551 gnd.n300 gnd.n299 585
R1552 gnd.n299 gnd.n298 585
R1553 gnd.n6580 gnd.n6579 585
R1554 gnd.n6579 gnd.n6578 585
R1555 gnd.n303 gnd.n302 585
R1556 gnd.n6577 gnd.n303 585
R1557 gnd.n6575 gnd.n6574 585
R1558 gnd.n6576 gnd.n6575 585
R1559 gnd.n306 gnd.n305 585
R1560 gnd.n305 gnd.n304 585
R1561 gnd.n6570 gnd.n6569 585
R1562 gnd.n6569 gnd.n6568 585
R1563 gnd.n309 gnd.n308 585
R1564 gnd.n6567 gnd.n309 585
R1565 gnd.n6565 gnd.n6564 585
R1566 gnd.n6566 gnd.n6565 585
R1567 gnd.n5884 gnd.n5883 585
R1568 gnd.n5885 gnd.n5884 585
R1569 gnd.n849 gnd.n848 585
R1570 gnd.n5878 gnd.n849 585
R1571 gnd.n5893 gnd.n5892 585
R1572 gnd.n5892 gnd.n5891 585
R1573 gnd.n5894 gnd.n844 585
R1574 gnd.n4188 gnd.n844 585
R1575 gnd.n5896 gnd.n5895 585
R1576 gnd.n5897 gnd.n5896 585
R1577 gnd.n829 gnd.n828 585
R1578 gnd.n4182 gnd.n829 585
R1579 gnd.n5905 gnd.n5904 585
R1580 gnd.n5904 gnd.n5903 585
R1581 gnd.n5906 gnd.n824 585
R1582 gnd.n4199 gnd.n824 585
R1583 gnd.n5908 gnd.n5907 585
R1584 gnd.n5909 gnd.n5908 585
R1585 gnd.n808 gnd.n807 585
R1586 gnd.n4175 gnd.n808 585
R1587 gnd.n5917 gnd.n5916 585
R1588 gnd.n5916 gnd.n5915 585
R1589 gnd.n5918 gnd.n803 585
R1590 gnd.n4167 gnd.n803 585
R1591 gnd.n5920 gnd.n5919 585
R1592 gnd.n5921 gnd.n5920 585
R1593 gnd.n789 gnd.n788 585
R1594 gnd.n4161 gnd.n789 585
R1595 gnd.n5929 gnd.n5928 585
R1596 gnd.n5928 gnd.n5927 585
R1597 gnd.n5930 gnd.n784 585
R1598 gnd.n4153 gnd.n784 585
R1599 gnd.n5932 gnd.n5931 585
R1600 gnd.n5933 gnd.n5932 585
R1601 gnd.n771 gnd.n770 585
R1602 gnd.n4109 gnd.n771 585
R1603 gnd.n5942 gnd.n5941 585
R1604 gnd.n5941 gnd.n5940 585
R1605 gnd.n5943 gnd.n766 585
R1606 gnd.n4117 gnd.n766 585
R1607 gnd.n5945 gnd.n5944 585
R1608 gnd.n5946 gnd.n5945 585
R1609 gnd.n755 gnd.n754 585
R1610 gnd.n4098 gnd.n755 585
R1611 gnd.n5955 gnd.n5954 585
R1612 gnd.n5954 gnd.n5953 585
R1613 gnd.n5956 gnd.n749 585
R1614 gnd.n4090 gnd.n749 585
R1615 gnd.n5958 gnd.n5957 585
R1616 gnd.n5959 gnd.n5958 585
R1617 gnd.n750 gnd.n748 585
R1618 gnd.n4072 gnd.n748 585
R1619 gnd.n4047 gnd.n737 585
R1620 gnd.n5966 gnd.n737 585
R1621 gnd.n4049 gnd.n4048 585
R1622 gnd.n4048 gnd.n733 585
R1623 gnd.n4050 gnd.n2136 585
R1624 gnd.n4063 gnd.n2136 585
R1625 gnd.n4051 gnd.n2146 585
R1626 gnd.n2146 gnd.n2144 585
R1627 gnd.n4053 gnd.n4052 585
R1628 gnd.n4054 gnd.n4053 585
R1629 gnd.n2147 gnd.n2145 585
R1630 gnd.n4036 gnd.n2145 585
R1631 gnd.n4009 gnd.n4008 585
R1632 gnd.n4008 gnd.n2154 585
R1633 gnd.n4010 gnd.n2162 585
R1634 gnd.n4024 gnd.n2162 585
R1635 gnd.n4011 gnd.n2172 585
R1636 gnd.n2172 gnd.n2160 585
R1637 gnd.n4013 gnd.n4012 585
R1638 gnd.n4014 gnd.n4013 585
R1639 gnd.n2173 gnd.n2171 585
R1640 gnd.n3999 gnd.n2171 585
R1641 gnd.n3974 gnd.n3973 585
R1642 gnd.n3973 gnd.n2179 585
R1643 gnd.n3975 gnd.n2187 585
R1644 gnd.n3989 gnd.n2187 585
R1645 gnd.n3976 gnd.n2197 585
R1646 gnd.n2197 gnd.n2185 585
R1647 gnd.n3978 gnd.n3977 585
R1648 gnd.n3979 gnd.n3978 585
R1649 gnd.n2198 gnd.n2196 585
R1650 gnd.n3744 gnd.n2196 585
R1651 gnd.n3963 gnd.n3962 585
R1652 gnd.n3962 gnd.n3961 585
R1653 gnd.n3691 gnd.n2204 585
R1654 gnd.n3694 gnd.n3692 585
R1655 gnd.n3697 gnd.n3696 585
R1656 gnd.n3688 gnd.n3687 585
R1657 gnd.n3702 gnd.n3701 585
R1658 gnd.n3704 gnd.n3686 585
R1659 gnd.n3707 gnd.n3706 585
R1660 gnd.n3684 gnd.n3683 585
R1661 gnd.n3712 gnd.n3711 585
R1662 gnd.n3714 gnd.n3682 585
R1663 gnd.n3717 gnd.n3716 585
R1664 gnd.n3680 gnd.n3679 585
R1665 gnd.n3722 gnd.n3721 585
R1666 gnd.n3724 gnd.n3678 585
R1667 gnd.n3727 gnd.n3726 585
R1668 gnd.n3676 gnd.n3675 585
R1669 gnd.n3732 gnd.n3731 585
R1670 gnd.n3734 gnd.n3674 585
R1671 gnd.n3736 gnd.n3735 585
R1672 gnd.n3735 gnd.n3667 585
R1673 gnd.n5805 gnd.n5804 585
R1674 gnd.n5806 gnd.n964 585
R1675 gnd.n5807 gnd.n959 585
R1676 gnd.n977 gnd.n948 585
R1677 gnd.n5814 gnd.n947 585
R1678 gnd.n5815 gnd.n946 585
R1679 gnd.n974 gnd.n940 585
R1680 gnd.n5822 gnd.n939 585
R1681 gnd.n5823 gnd.n938 585
R1682 gnd.n972 gnd.n930 585
R1683 gnd.n5830 gnd.n929 585
R1684 gnd.n5831 gnd.n928 585
R1685 gnd.n969 gnd.n922 585
R1686 gnd.n5838 gnd.n921 585
R1687 gnd.n5839 gnd.n920 585
R1688 gnd.n967 gnd.n912 585
R1689 gnd.n5846 gnd.n911 585
R1690 gnd.n5847 gnd.n910 585
R1691 gnd.n909 gnd.n863 585
R1692 gnd.n5802 gnd.n863 585
R1693 gnd.n869 gnd.n861 585
R1694 gnd.n5885 gnd.n861 585
R1695 gnd.n5877 gnd.n5876 585
R1696 gnd.n5878 gnd.n5877 585
R1697 gnd.n868 gnd.n852 585
R1698 gnd.n5891 gnd.n852 585
R1699 gnd.n4191 gnd.n4189 585
R1700 gnd.n4189 gnd.n4188 585
R1701 gnd.n4192 gnd.n842 585
R1702 gnd.n5897 gnd.n842 585
R1703 gnd.n4193 gnd.n2100 585
R1704 gnd.n4182 gnd.n2100 585
R1705 gnd.n2097 gnd.n831 585
R1706 gnd.n5903 gnd.n831 585
R1707 gnd.n4198 gnd.n4197 585
R1708 gnd.n4199 gnd.n4198 585
R1709 gnd.n2096 gnd.n822 585
R1710 gnd.n5909 gnd.n822 585
R1711 gnd.n4174 gnd.n4173 585
R1712 gnd.n4175 gnd.n4174 585
R1713 gnd.n2103 gnd.n811 585
R1714 gnd.n5915 gnd.n811 585
R1715 gnd.n4169 gnd.n4168 585
R1716 gnd.n4168 gnd.n4167 585
R1717 gnd.n2105 gnd.n802 585
R1718 gnd.n5921 gnd.n802 585
R1719 gnd.n4160 gnd.n4159 585
R1720 gnd.n4161 gnd.n4160 585
R1721 gnd.n2109 gnd.n791 585
R1722 gnd.n5927 gnd.n791 585
R1723 gnd.n4155 gnd.n4154 585
R1724 gnd.n4154 gnd.n4153 585
R1725 gnd.n2111 gnd.n782 585
R1726 gnd.n5933 gnd.n782 585
R1727 gnd.n4111 gnd.n4110 585
R1728 gnd.n4110 gnd.n4109 585
R1729 gnd.n2121 gnd.n774 585
R1730 gnd.n5940 gnd.n774 585
R1731 gnd.n4116 gnd.n4115 585
R1732 gnd.n4117 gnd.n4116 585
R1733 gnd.n2120 gnd.n765 585
R1734 gnd.n5946 gnd.n765 585
R1735 gnd.n4097 gnd.n4096 585
R1736 gnd.n4098 gnd.n4097 585
R1737 gnd.n2125 gnd.n757 585
R1738 gnd.n5953 gnd.n757 585
R1739 gnd.n4092 gnd.n4091 585
R1740 gnd.n4091 gnd.n4090 585
R1741 gnd.n2127 gnd.n746 585
R1742 gnd.n5959 gnd.n746 585
R1743 gnd.n4071 gnd.n4070 585
R1744 gnd.n4072 gnd.n4071 585
R1745 gnd.n2130 gnd.n735 585
R1746 gnd.n5966 gnd.n735 585
R1747 gnd.n4066 gnd.n4065 585
R1748 gnd.n4065 gnd.n733 585
R1749 gnd.n4064 gnd.n2132 585
R1750 gnd.n4064 gnd.n4063 585
R1751 gnd.n4032 gnd.n2133 585
R1752 gnd.n2144 gnd.n2133 585
R1753 gnd.n4033 gnd.n2143 585
R1754 gnd.n4054 gnd.n2143 585
R1755 gnd.n4035 gnd.n4034 585
R1756 gnd.n4036 gnd.n4035 585
R1757 gnd.n2156 gnd.n2155 585
R1758 gnd.n2155 gnd.n2154 585
R1759 gnd.n4026 gnd.n4025 585
R1760 gnd.n4025 gnd.n4024 585
R1761 gnd.n2159 gnd.n2158 585
R1762 gnd.n2160 gnd.n2159 585
R1763 gnd.n3996 gnd.n2170 585
R1764 gnd.n4014 gnd.n2170 585
R1765 gnd.n3998 gnd.n3997 585
R1766 gnd.n3999 gnd.n3998 585
R1767 gnd.n2181 gnd.n2180 585
R1768 gnd.n2180 gnd.n2179 585
R1769 gnd.n3991 gnd.n3990 585
R1770 gnd.n3990 gnd.n3989 585
R1771 gnd.n2184 gnd.n2183 585
R1772 gnd.n2185 gnd.n2184 585
R1773 gnd.n3741 gnd.n2195 585
R1774 gnd.n3979 gnd.n2195 585
R1775 gnd.n3743 gnd.n3742 585
R1776 gnd.n3744 gnd.n3743 585
R1777 gnd.n3670 gnd.n3669 585
R1778 gnd.n3961 gnd.n3669 585
R1779 gnd.n3574 gnd.n3573 585
R1780 gnd.n3575 gnd.n3574 585
R1781 gnd.n2281 gnd.n2280 585
R1782 gnd.n2287 gnd.n2280 585
R1783 gnd.n3549 gnd.n2299 585
R1784 gnd.n2299 gnd.n2286 585
R1785 gnd.n3551 gnd.n3550 585
R1786 gnd.n3552 gnd.n3551 585
R1787 gnd.n2300 gnd.n2298 585
R1788 gnd.n2298 gnd.n2294 585
R1789 gnd.n3283 gnd.n3282 585
R1790 gnd.n3282 gnd.n3281 585
R1791 gnd.n2305 gnd.n2304 585
R1792 gnd.n3252 gnd.n2305 585
R1793 gnd.n3272 gnd.n3271 585
R1794 gnd.n3271 gnd.n3270 585
R1795 gnd.n2312 gnd.n2311 585
R1796 gnd.n3258 gnd.n2312 585
R1797 gnd.n3228 gnd.n2332 585
R1798 gnd.n2332 gnd.n2331 585
R1799 gnd.n3230 gnd.n3229 585
R1800 gnd.n3231 gnd.n3230 585
R1801 gnd.n2333 gnd.n2330 585
R1802 gnd.n2341 gnd.n2330 585
R1803 gnd.n3206 gnd.n2353 585
R1804 gnd.n2353 gnd.n2340 585
R1805 gnd.n3208 gnd.n3207 585
R1806 gnd.n3209 gnd.n3208 585
R1807 gnd.n2354 gnd.n2352 585
R1808 gnd.n2352 gnd.n2348 585
R1809 gnd.n3194 gnd.n3193 585
R1810 gnd.n3193 gnd.n3192 585
R1811 gnd.n2359 gnd.n2358 585
R1812 gnd.n2369 gnd.n2359 585
R1813 gnd.n3183 gnd.n3182 585
R1814 gnd.n3182 gnd.n3181 585
R1815 gnd.n2366 gnd.n2365 585
R1816 gnd.n3169 gnd.n2366 585
R1817 gnd.n3143 gnd.n2387 585
R1818 gnd.n2387 gnd.n2376 585
R1819 gnd.n3145 gnd.n3144 585
R1820 gnd.n3146 gnd.n3145 585
R1821 gnd.n2388 gnd.n2386 585
R1822 gnd.n2396 gnd.n2386 585
R1823 gnd.n3121 gnd.n2408 585
R1824 gnd.n2408 gnd.n2395 585
R1825 gnd.n3123 gnd.n3122 585
R1826 gnd.n3124 gnd.n3123 585
R1827 gnd.n2409 gnd.n2407 585
R1828 gnd.n2407 gnd.n2403 585
R1829 gnd.n3109 gnd.n3108 585
R1830 gnd.n3108 gnd.n3107 585
R1831 gnd.n2414 gnd.n2413 585
R1832 gnd.n2423 gnd.n2414 585
R1833 gnd.n3098 gnd.n3097 585
R1834 gnd.n3097 gnd.n3096 585
R1835 gnd.n2421 gnd.n2420 585
R1836 gnd.n3084 gnd.n2421 585
R1837 gnd.n2522 gnd.n2521 585
R1838 gnd.n2522 gnd.n2430 585
R1839 gnd.n3041 gnd.n3040 585
R1840 gnd.n3040 gnd.n3039 585
R1841 gnd.n3042 gnd.n2516 585
R1842 gnd.n2527 gnd.n2516 585
R1843 gnd.n3044 gnd.n3043 585
R1844 gnd.n3045 gnd.n3044 585
R1845 gnd.n2517 gnd.n2515 585
R1846 gnd.n2540 gnd.n2515 585
R1847 gnd.n2500 gnd.n2499 585
R1848 gnd.n2503 gnd.n2500 585
R1849 gnd.n3055 gnd.n3054 585
R1850 gnd.n3054 gnd.n3053 585
R1851 gnd.n3056 gnd.n2494 585
R1852 gnd.n3015 gnd.n2494 585
R1853 gnd.n3058 gnd.n3057 585
R1854 gnd.n3059 gnd.n3058 585
R1855 gnd.n2495 gnd.n2493 585
R1856 gnd.n2554 gnd.n2493 585
R1857 gnd.n3007 gnd.n3006 585
R1858 gnd.n3006 gnd.n3005 585
R1859 gnd.n2551 gnd.n2550 585
R1860 gnd.n2989 gnd.n2551 585
R1861 gnd.n2976 gnd.n2570 585
R1862 gnd.n2570 gnd.n2569 585
R1863 gnd.n2978 gnd.n2977 585
R1864 gnd.n2979 gnd.n2978 585
R1865 gnd.n2571 gnd.n2568 585
R1866 gnd.n2577 gnd.n2568 585
R1867 gnd.n2957 gnd.n2956 585
R1868 gnd.n2958 gnd.n2957 585
R1869 gnd.n2588 gnd.n2587 585
R1870 gnd.n2587 gnd.n2583 585
R1871 gnd.n2947 gnd.n2946 585
R1872 gnd.n2948 gnd.n2947 585
R1873 gnd.n2598 gnd.n2597 585
R1874 gnd.n2603 gnd.n2597 585
R1875 gnd.n2925 gnd.n2616 585
R1876 gnd.n2616 gnd.n2602 585
R1877 gnd.n2927 gnd.n2926 585
R1878 gnd.n2928 gnd.n2927 585
R1879 gnd.n2617 gnd.n2615 585
R1880 gnd.n2615 gnd.n2611 585
R1881 gnd.n2916 gnd.n2915 585
R1882 gnd.n2917 gnd.n2916 585
R1883 gnd.n2624 gnd.n2623 585
R1884 gnd.n2628 gnd.n2623 585
R1885 gnd.n2893 gnd.n2645 585
R1886 gnd.n2645 gnd.n2627 585
R1887 gnd.n2895 gnd.n2894 585
R1888 gnd.n2896 gnd.n2895 585
R1889 gnd.n2646 gnd.n2644 585
R1890 gnd.n2644 gnd.n2635 585
R1891 gnd.n2888 gnd.n2887 585
R1892 gnd.n2887 gnd.n2886 585
R1893 gnd.n2693 gnd.n2692 585
R1894 gnd.n2694 gnd.n2693 585
R1895 gnd.n2847 gnd.n2846 585
R1896 gnd.n2848 gnd.n2847 585
R1897 gnd.n2703 gnd.n2702 585
R1898 gnd.n2702 gnd.n2701 585
R1899 gnd.n2842 gnd.n2841 585
R1900 gnd.n2841 gnd.n2840 585
R1901 gnd.n2706 gnd.n2705 585
R1902 gnd.n2707 gnd.n2706 585
R1903 gnd.n2831 gnd.n2830 585
R1904 gnd.n2832 gnd.n2831 585
R1905 gnd.n2714 gnd.n2713 585
R1906 gnd.n2823 gnd.n2713 585
R1907 gnd.n2826 gnd.n2825 585
R1908 gnd.n2825 gnd.n2824 585
R1909 gnd.n2717 gnd.n2716 585
R1910 gnd.n2718 gnd.n2717 585
R1911 gnd.n2812 gnd.n2811 585
R1912 gnd.n2810 gnd.n2736 585
R1913 gnd.n2809 gnd.n2735 585
R1914 gnd.n2814 gnd.n2735 585
R1915 gnd.n2808 gnd.n2807 585
R1916 gnd.n2806 gnd.n2805 585
R1917 gnd.n2804 gnd.n2803 585
R1918 gnd.n2802 gnd.n2801 585
R1919 gnd.n2800 gnd.n2799 585
R1920 gnd.n2798 gnd.n2797 585
R1921 gnd.n2796 gnd.n2795 585
R1922 gnd.n2794 gnd.n2793 585
R1923 gnd.n2792 gnd.n2791 585
R1924 gnd.n2790 gnd.n2789 585
R1925 gnd.n2788 gnd.n2787 585
R1926 gnd.n2786 gnd.n2785 585
R1927 gnd.n2784 gnd.n2783 585
R1928 gnd.n2782 gnd.n2781 585
R1929 gnd.n2780 gnd.n2779 585
R1930 gnd.n2778 gnd.n2777 585
R1931 gnd.n2776 gnd.n2775 585
R1932 gnd.n2774 gnd.n2773 585
R1933 gnd.n2772 gnd.n2771 585
R1934 gnd.n2770 gnd.n2769 585
R1935 gnd.n2768 gnd.n2767 585
R1936 gnd.n2766 gnd.n2765 585
R1937 gnd.n2723 gnd.n2722 585
R1938 gnd.n2817 gnd.n2816 585
R1939 gnd.n3578 gnd.n3577 585
R1940 gnd.n3580 gnd.n3579 585
R1941 gnd.n3582 gnd.n3581 585
R1942 gnd.n3584 gnd.n3583 585
R1943 gnd.n3586 gnd.n3585 585
R1944 gnd.n3588 gnd.n3587 585
R1945 gnd.n3590 gnd.n3589 585
R1946 gnd.n3592 gnd.n3591 585
R1947 gnd.n3594 gnd.n3593 585
R1948 gnd.n3596 gnd.n3595 585
R1949 gnd.n3598 gnd.n3597 585
R1950 gnd.n3600 gnd.n3599 585
R1951 gnd.n3602 gnd.n3601 585
R1952 gnd.n3604 gnd.n3603 585
R1953 gnd.n3606 gnd.n3605 585
R1954 gnd.n3608 gnd.n3607 585
R1955 gnd.n3610 gnd.n3609 585
R1956 gnd.n3612 gnd.n3611 585
R1957 gnd.n3614 gnd.n3613 585
R1958 gnd.n3616 gnd.n3615 585
R1959 gnd.n3618 gnd.n3617 585
R1960 gnd.n3620 gnd.n3619 585
R1961 gnd.n3622 gnd.n3621 585
R1962 gnd.n3624 gnd.n3623 585
R1963 gnd.n3626 gnd.n3625 585
R1964 gnd.n3627 gnd.n2248 585
R1965 gnd.n3628 gnd.n2206 585
R1966 gnd.n3666 gnd.n2206 585
R1967 gnd.n3576 gnd.n2278 585
R1968 gnd.n3576 gnd.n3575 585
R1969 gnd.n3245 gnd.n2277 585
R1970 gnd.n2287 gnd.n2277 585
R1971 gnd.n3247 gnd.n3246 585
R1972 gnd.n3246 gnd.n2286 585
R1973 gnd.n3248 gnd.n2296 585
R1974 gnd.n3552 gnd.n2296 585
R1975 gnd.n3250 gnd.n3249 585
R1976 gnd.n3249 gnd.n2294 585
R1977 gnd.n3251 gnd.n2307 585
R1978 gnd.n3281 gnd.n2307 585
R1979 gnd.n3254 gnd.n3253 585
R1980 gnd.n3253 gnd.n3252 585
R1981 gnd.n3255 gnd.n2314 585
R1982 gnd.n3270 gnd.n2314 585
R1983 gnd.n3257 gnd.n3256 585
R1984 gnd.n3258 gnd.n3257 585
R1985 gnd.n2324 gnd.n2323 585
R1986 gnd.n2331 gnd.n2323 585
R1987 gnd.n3233 gnd.n3232 585
R1988 gnd.n3232 gnd.n3231 585
R1989 gnd.n2327 gnd.n2326 585
R1990 gnd.n2341 gnd.n2327 585
R1991 gnd.n3159 gnd.n3158 585
R1992 gnd.n3158 gnd.n2340 585
R1993 gnd.n3160 gnd.n2350 585
R1994 gnd.n3209 gnd.n2350 585
R1995 gnd.n3162 gnd.n3161 585
R1996 gnd.n3161 gnd.n2348 585
R1997 gnd.n3163 gnd.n2361 585
R1998 gnd.n3192 gnd.n2361 585
R1999 gnd.n3165 gnd.n3164 585
R2000 gnd.n3164 gnd.n2369 585
R2001 gnd.n3166 gnd.n2368 585
R2002 gnd.n3181 gnd.n2368 585
R2003 gnd.n3168 gnd.n3167 585
R2004 gnd.n3169 gnd.n3168 585
R2005 gnd.n2380 gnd.n2379 585
R2006 gnd.n2379 gnd.n2376 585
R2007 gnd.n3148 gnd.n3147 585
R2008 gnd.n3147 gnd.n3146 585
R2009 gnd.n2383 gnd.n2382 585
R2010 gnd.n2396 gnd.n2383 585
R2011 gnd.n3072 gnd.n3071 585
R2012 gnd.n3071 gnd.n2395 585
R2013 gnd.n3073 gnd.n2405 585
R2014 gnd.n3124 gnd.n2405 585
R2015 gnd.n3075 gnd.n3074 585
R2016 gnd.n3074 gnd.n2403 585
R2017 gnd.n3076 gnd.n2416 585
R2018 gnd.n3107 gnd.n2416 585
R2019 gnd.n3078 gnd.n3077 585
R2020 gnd.n3077 gnd.n2423 585
R2021 gnd.n3079 gnd.n2422 585
R2022 gnd.n3096 gnd.n2422 585
R2023 gnd.n3081 gnd.n3080 585
R2024 gnd.n3084 gnd.n3081 585
R2025 gnd.n2433 gnd.n2432 585
R2026 gnd.n2432 gnd.n2430 585
R2027 gnd.n2524 gnd.n2523 585
R2028 gnd.n3039 gnd.n2523 585
R2029 gnd.n2526 gnd.n2525 585
R2030 gnd.n2527 gnd.n2526 585
R2031 gnd.n2537 gnd.n2513 585
R2032 gnd.n3045 gnd.n2513 585
R2033 gnd.n2539 gnd.n2538 585
R2034 gnd.n2540 gnd.n2539 585
R2035 gnd.n2536 gnd.n2535 585
R2036 gnd.n2536 gnd.n2503 585
R2037 gnd.n2534 gnd.n2501 585
R2038 gnd.n3053 gnd.n2501 585
R2039 gnd.n2490 gnd.n2488 585
R2040 gnd.n3015 gnd.n2490 585
R2041 gnd.n3061 gnd.n3060 585
R2042 gnd.n3060 gnd.n3059 585
R2043 gnd.n2489 gnd.n2487 585
R2044 gnd.n2554 gnd.n2489 585
R2045 gnd.n2986 gnd.n2553 585
R2046 gnd.n3005 gnd.n2553 585
R2047 gnd.n2988 gnd.n2987 585
R2048 gnd.n2989 gnd.n2988 585
R2049 gnd.n2563 gnd.n2562 585
R2050 gnd.n2569 gnd.n2562 585
R2051 gnd.n2981 gnd.n2980 585
R2052 gnd.n2980 gnd.n2979 585
R2053 gnd.n2566 gnd.n2565 585
R2054 gnd.n2577 gnd.n2566 585
R2055 gnd.n2866 gnd.n2585 585
R2056 gnd.n2958 gnd.n2585 585
R2057 gnd.n2868 gnd.n2867 585
R2058 gnd.n2867 gnd.n2583 585
R2059 gnd.n2869 gnd.n2596 585
R2060 gnd.n2948 gnd.n2596 585
R2061 gnd.n2871 gnd.n2870 585
R2062 gnd.n2871 gnd.n2603 585
R2063 gnd.n2873 gnd.n2872 585
R2064 gnd.n2872 gnd.n2602 585
R2065 gnd.n2874 gnd.n2613 585
R2066 gnd.n2928 gnd.n2613 585
R2067 gnd.n2876 gnd.n2875 585
R2068 gnd.n2875 gnd.n2611 585
R2069 gnd.n2877 gnd.n2622 585
R2070 gnd.n2917 gnd.n2622 585
R2071 gnd.n2879 gnd.n2878 585
R2072 gnd.n2879 gnd.n2628 585
R2073 gnd.n2881 gnd.n2880 585
R2074 gnd.n2880 gnd.n2627 585
R2075 gnd.n2882 gnd.n2643 585
R2076 gnd.n2896 gnd.n2643 585
R2077 gnd.n2883 gnd.n2696 585
R2078 gnd.n2696 gnd.n2635 585
R2079 gnd.n2885 gnd.n2884 585
R2080 gnd.n2886 gnd.n2885 585
R2081 gnd.n2697 gnd.n2695 585
R2082 gnd.n2695 gnd.n2694 585
R2083 gnd.n2850 gnd.n2849 585
R2084 gnd.n2849 gnd.n2848 585
R2085 gnd.n2700 gnd.n2699 585
R2086 gnd.n2701 gnd.n2700 585
R2087 gnd.n2839 gnd.n2838 585
R2088 gnd.n2840 gnd.n2839 585
R2089 gnd.n2709 gnd.n2708 585
R2090 gnd.n2708 gnd.n2707 585
R2091 gnd.n2834 gnd.n2833 585
R2092 gnd.n2833 gnd.n2832 585
R2093 gnd.n2712 gnd.n2711 585
R2094 gnd.n2823 gnd.n2712 585
R2095 gnd.n2822 gnd.n2821 585
R2096 gnd.n2824 gnd.n2822 585
R2097 gnd.n2720 gnd.n2719 585
R2098 gnd.n2719 gnd.n2718 585
R2099 gnd.n7146 gnd.n7145 585
R2100 gnd.n7147 gnd.n7146 585
R2101 gnd.n158 gnd.n157 585
R2102 gnd.n167 gnd.n158 585
R2103 gnd.n7155 gnd.n7154 585
R2104 gnd.n7154 gnd.n7153 585
R2105 gnd.n7156 gnd.n153 585
R2106 gnd.n153 gnd.n152 585
R2107 gnd.n7158 gnd.n7157 585
R2108 gnd.n7159 gnd.n7158 585
R2109 gnd.n139 gnd.n138 585
R2110 gnd.n142 gnd.n139 585
R2111 gnd.n7167 gnd.n7166 585
R2112 gnd.n7166 gnd.n7165 585
R2113 gnd.n7168 gnd.n134 585
R2114 gnd.n134 gnd.n133 585
R2115 gnd.n7170 gnd.n7169 585
R2116 gnd.n7171 gnd.n7170 585
R2117 gnd.n119 gnd.n118 585
R2118 gnd.n130 gnd.n119 585
R2119 gnd.n7179 gnd.n7178 585
R2120 gnd.n7178 gnd.n7177 585
R2121 gnd.n7180 gnd.n114 585
R2122 gnd.n120 gnd.n114 585
R2123 gnd.n7182 gnd.n7181 585
R2124 gnd.n7183 gnd.n7182 585
R2125 gnd.n101 gnd.n100 585
R2126 gnd.n111 gnd.n101 585
R2127 gnd.n7191 gnd.n7190 585
R2128 gnd.n7190 gnd.n7189 585
R2129 gnd.n7192 gnd.n95 585
R2130 gnd.n7116 gnd.n95 585
R2131 gnd.n7194 gnd.n7193 585
R2132 gnd.n7195 gnd.n7194 585
R2133 gnd.n96 gnd.n94 585
R2134 gnd.n6791 gnd.n94 585
R2135 gnd.n6786 gnd.n6785 585
R2136 gnd.n6785 gnd.n6784 585
R2137 gnd.n180 gnd.n76 585
R2138 gnd.n7203 gnd.n76 585
R2139 gnd.n5305 gnd.n5304 585
R2140 gnd.n5306 gnd.n5305 585
R2141 gnd.n1599 gnd.n1598 585
R2142 gnd.n1598 gnd.n1596 585
R2143 gnd.n5296 gnd.n5295 585
R2144 gnd.n5297 gnd.n5296 585
R2145 gnd.n1577 gnd.n1576 585
R2146 gnd.n5315 gnd.n1577 585
R2147 gnd.n5322 gnd.n5321 585
R2148 gnd.n5321 gnd.n5320 585
R2149 gnd.n5323 gnd.n1572 585
R2150 gnd.n5288 gnd.n1572 585
R2151 gnd.n5325 gnd.n5324 585
R2152 gnd.n5326 gnd.n5325 585
R2153 gnd.n1560 gnd.n1559 585
R2154 gnd.n5276 gnd.n1560 585
R2155 gnd.n5334 gnd.n5333 585
R2156 gnd.n5333 gnd.n5332 585
R2157 gnd.n5335 gnd.n1555 585
R2158 gnd.n5269 gnd.n1555 585
R2159 gnd.n5337 gnd.n5336 585
R2160 gnd.n5338 gnd.n5337 585
R2161 gnd.n1540 gnd.n1539 585
R2162 gnd.n5261 gnd.n1540 585
R2163 gnd.n5346 gnd.n5345 585
R2164 gnd.n5345 gnd.n5344 585
R2165 gnd.n5347 gnd.n1535 585
R2166 gnd.n5201 gnd.n1535 585
R2167 gnd.n5349 gnd.n5348 585
R2168 gnd.n5350 gnd.n5349 585
R2169 gnd.n1520 gnd.n1519 585
R2170 gnd.n5192 gnd.n1520 585
R2171 gnd.n5358 gnd.n5357 585
R2172 gnd.n5357 gnd.n5356 585
R2173 gnd.n5359 gnd.n1513 585
R2174 gnd.n5186 gnd.n1513 585
R2175 gnd.n5361 gnd.n5360 585
R2176 gnd.n5362 gnd.n5361 585
R2177 gnd.n1514 gnd.n1512 585
R2178 gnd.n5179 gnd.n1512 585
R2179 gnd.n1496 gnd.n1490 585
R2180 gnd.n5368 gnd.n1496 585
R2181 gnd.n5373 gnd.n1488 585
R2182 gnd.n5218 gnd.n1488 585
R2183 gnd.n5375 gnd.n5374 585
R2184 gnd.n5376 gnd.n5375 585
R2185 gnd.n1487 gnd.n1327 585
R2186 gnd.n5543 gnd.n1328 585
R2187 gnd.n5542 gnd.n1329 585
R2188 gnd.n1404 gnd.n1330 585
R2189 gnd.n5535 gnd.n1336 585
R2190 gnd.n5534 gnd.n1337 585
R2191 gnd.n1407 gnd.n1338 585
R2192 gnd.n5527 gnd.n1344 585
R2193 gnd.n5526 gnd.n1345 585
R2194 gnd.n1409 gnd.n1346 585
R2195 gnd.n5519 gnd.n1352 585
R2196 gnd.n5518 gnd.n1353 585
R2197 gnd.n1412 gnd.n1354 585
R2198 gnd.n5511 gnd.n1360 585
R2199 gnd.n5510 gnd.n1361 585
R2200 gnd.n1414 gnd.n1362 585
R2201 gnd.n5503 gnd.n1370 585
R2202 gnd.n5502 gnd.n5499 585
R2203 gnd.n1373 gnd.n1371 585
R2204 gnd.n5497 gnd.n1373 585
R2205 gnd.n7089 gnd.n7088 585
R2206 gnd.n6815 gnd.n6814 585
R2207 gnd.n6872 gnd.n6871 585
R2208 gnd.n6824 gnd.n6823 585
R2209 gnd.n6867 gnd.n6866 585
R2210 gnd.n6865 gnd.n6864 585
R2211 gnd.n6863 gnd.n6862 585
R2212 gnd.n6856 gnd.n6826 585
R2213 gnd.n6858 gnd.n6857 585
R2214 gnd.n6855 gnd.n6854 585
R2215 gnd.n6853 gnd.n6852 585
R2216 gnd.n6846 gnd.n6828 585
R2217 gnd.n6848 gnd.n6847 585
R2218 gnd.n6845 gnd.n6844 585
R2219 gnd.n6843 gnd.n6842 585
R2220 gnd.n6836 gnd.n6830 585
R2221 gnd.n6838 gnd.n6837 585
R2222 gnd.n6835 gnd.n6834 585
R2223 gnd.n6833 gnd.n171 585
R2224 gnd.n7086 gnd.n171 585
R2225 gnd.n7092 gnd.n169 585
R2226 gnd.n7147 gnd.n169 585
R2227 gnd.n7094 gnd.n7093 585
R2228 gnd.n7093 gnd.n167 585
R2229 gnd.n7095 gnd.n160 585
R2230 gnd.n7153 gnd.n160 585
R2231 gnd.n7097 gnd.n7096 585
R2232 gnd.n7096 gnd.n152 585
R2233 gnd.n7098 gnd.n151 585
R2234 gnd.n7159 gnd.n151 585
R2235 gnd.n7100 gnd.n7099 585
R2236 gnd.n7099 gnd.n142 585
R2237 gnd.n7101 gnd.n141 585
R2238 gnd.n7165 gnd.n141 585
R2239 gnd.n7103 gnd.n7102 585
R2240 gnd.n7102 gnd.n133 585
R2241 gnd.n7104 gnd.n132 585
R2242 gnd.n7171 gnd.n132 585
R2243 gnd.n7106 gnd.n7105 585
R2244 gnd.n7105 gnd.n130 585
R2245 gnd.n7107 gnd.n122 585
R2246 gnd.n7177 gnd.n122 585
R2247 gnd.n7109 gnd.n7108 585
R2248 gnd.n7108 gnd.n120 585
R2249 gnd.n7110 gnd.n113 585
R2250 gnd.n7183 gnd.n113 585
R2251 gnd.n7112 gnd.n7111 585
R2252 gnd.n7111 gnd.n111 585
R2253 gnd.n7113 gnd.n103 585
R2254 gnd.n7189 gnd.n103 585
R2255 gnd.n7115 gnd.n7114 585
R2256 gnd.n7116 gnd.n7115 585
R2257 gnd.n175 gnd.n92 585
R2258 gnd.n7195 gnd.n92 585
R2259 gnd.n6793 gnd.n6792 585
R2260 gnd.n6792 gnd.n6791 585
R2261 gnd.n72 gnd.n71 585
R2262 gnd.n6784 gnd.n72 585
R2263 gnd.n7205 gnd.n7204 585
R2264 gnd.n7204 gnd.n7203 585
R2265 gnd.n7206 gnd.n70 585
R2266 gnd.n5306 gnd.n70 585
R2267 gnd.n1602 gnd.n68 585
R2268 gnd.n1602 gnd.n1596 585
R2269 gnd.n5281 gnd.n1603 585
R2270 gnd.n5297 gnd.n1603 585
R2271 gnd.n5282 gnd.n1586 585
R2272 gnd.n5315 gnd.n1586 585
R2273 gnd.n1607 gnd.n1580 585
R2274 gnd.n5320 gnd.n1580 585
R2275 gnd.n5287 gnd.n5286 585
R2276 gnd.n5288 gnd.n5287 585
R2277 gnd.n1606 gnd.n1570 585
R2278 gnd.n5326 gnd.n1570 585
R2279 gnd.n5278 gnd.n5277 585
R2280 gnd.n5277 gnd.n5276 585
R2281 gnd.n1609 gnd.n1563 585
R2282 gnd.n5332 gnd.n1563 585
R2283 gnd.n5268 gnd.n5267 585
R2284 gnd.n5269 gnd.n5268 585
R2285 gnd.n1612 gnd.n1553 585
R2286 gnd.n5338 gnd.n1553 585
R2287 gnd.n5263 gnd.n5262 585
R2288 gnd.n5262 gnd.n5261 585
R2289 gnd.n1614 gnd.n1543 585
R2290 gnd.n5344 gnd.n1543 585
R2291 gnd.n5204 gnd.n5202 585
R2292 gnd.n5202 gnd.n5201 585
R2293 gnd.n5205 gnd.n1533 585
R2294 gnd.n5350 gnd.n1533 585
R2295 gnd.n5206 gnd.n5184 585
R2296 gnd.n5192 gnd.n5184 585
R2297 gnd.n5182 gnd.n1523 585
R2298 gnd.n5356 gnd.n1523 585
R2299 gnd.n5210 gnd.n5181 585
R2300 gnd.n5186 gnd.n5181 585
R2301 gnd.n5211 gnd.n1510 585
R2302 gnd.n5362 gnd.n1510 585
R2303 gnd.n5212 gnd.n5180 585
R2304 gnd.n5180 gnd.n5179 585
R2305 gnd.n1631 gnd.n1494 585
R2306 gnd.n5368 gnd.n1494 585
R2307 gnd.n5217 gnd.n5216 585
R2308 gnd.n5218 gnd.n5217 585
R2309 gnd.n1630 gnd.n1485 585
R2310 gnd.n5376 gnd.n1485 585
R2311 gnd.n3561 gnd.n2228 585
R2312 gnd.n2228 gnd.n2205 585
R2313 gnd.n3562 gnd.n2289 585
R2314 gnd.n2289 gnd.n2279 585
R2315 gnd.n3564 gnd.n3563 585
R2316 gnd.n3565 gnd.n3564 585
R2317 gnd.n2290 gnd.n2288 585
R2318 gnd.n2297 gnd.n2288 585
R2319 gnd.n3555 gnd.n3554 585
R2320 gnd.n3554 gnd.n3553 585
R2321 gnd.n2293 gnd.n2292 585
R2322 gnd.n3280 gnd.n2293 585
R2323 gnd.n3266 gnd.n2316 585
R2324 gnd.n2316 gnd.n2306 585
R2325 gnd.n3268 gnd.n3267 585
R2326 gnd.n3269 gnd.n3268 585
R2327 gnd.n2317 gnd.n2315 585
R2328 gnd.n2315 gnd.n2313 585
R2329 gnd.n3261 gnd.n3260 585
R2330 gnd.n3260 gnd.n3259 585
R2331 gnd.n2320 gnd.n2319 585
R2332 gnd.n2329 gnd.n2320 585
R2333 gnd.n3217 gnd.n2343 585
R2334 gnd.n2343 gnd.n2328 585
R2335 gnd.n3219 gnd.n3218 585
R2336 gnd.n3220 gnd.n3219 585
R2337 gnd.n2344 gnd.n2342 585
R2338 gnd.n2351 gnd.n2342 585
R2339 gnd.n3212 gnd.n3211 585
R2340 gnd.n3211 gnd.n3210 585
R2341 gnd.n2347 gnd.n2346 585
R2342 gnd.n3191 gnd.n2347 585
R2343 gnd.n3177 gnd.n2371 585
R2344 gnd.n2371 gnd.n2360 585
R2345 gnd.n3179 gnd.n3178 585
R2346 gnd.n3180 gnd.n3179 585
R2347 gnd.n2372 gnd.n2370 585
R2348 gnd.n2370 gnd.n2367 585
R2349 gnd.n3172 gnd.n3171 585
R2350 gnd.n3171 gnd.n3170 585
R2351 gnd.n2375 gnd.n2374 585
R2352 gnd.n2385 gnd.n2375 585
R2353 gnd.n3132 gnd.n2398 585
R2354 gnd.n2398 gnd.n2384 585
R2355 gnd.n3134 gnd.n3133 585
R2356 gnd.n3135 gnd.n3134 585
R2357 gnd.n2399 gnd.n2397 585
R2358 gnd.n2406 gnd.n2397 585
R2359 gnd.n3127 gnd.n3126 585
R2360 gnd.n3126 gnd.n3125 585
R2361 gnd.n2402 gnd.n2401 585
R2362 gnd.n3106 gnd.n2402 585
R2363 gnd.n3092 gnd.n2425 585
R2364 gnd.n2425 gnd.n2415 585
R2365 gnd.n3094 gnd.n3093 585
R2366 gnd.n3095 gnd.n3094 585
R2367 gnd.n2426 gnd.n2424 585
R2368 gnd.n3083 gnd.n2424 585
R2369 gnd.n3087 gnd.n3086 585
R2370 gnd.n3086 gnd.n3085 585
R2371 gnd.n2429 gnd.n2428 585
R2372 gnd.n3038 gnd.n2429 585
R2373 gnd.n2531 gnd.n2530 585
R2374 gnd.n2532 gnd.n2531 585
R2375 gnd.n2511 gnd.n2510 585
R2376 gnd.n2514 gnd.n2511 585
R2377 gnd.n3048 gnd.n3047 585
R2378 gnd.n3047 gnd.n3046 585
R2379 gnd.n3049 gnd.n2505 585
R2380 gnd.n2541 gnd.n2505 585
R2381 gnd.n3051 gnd.n3050 585
R2382 gnd.n3052 gnd.n3051 585
R2383 gnd.n2506 gnd.n2504 585
R2384 gnd.n3016 gnd.n2504 585
R2385 gnd.n3000 gnd.n2999 585
R2386 gnd.n2999 gnd.n2492 585
R2387 gnd.n3001 gnd.n2556 585
R2388 gnd.n2556 gnd.n2491 585
R2389 gnd.n3003 gnd.n3002 585
R2390 gnd.n3004 gnd.n3003 585
R2391 gnd.n2557 gnd.n2555 585
R2392 gnd.n2555 gnd.n2552 585
R2393 gnd.n2992 gnd.n2991 585
R2394 gnd.n2991 gnd.n2990 585
R2395 gnd.n2560 gnd.n2559 585
R2396 gnd.n2567 gnd.n2560 585
R2397 gnd.n2966 gnd.n2965 585
R2398 gnd.n2967 gnd.n2966 585
R2399 gnd.n2579 gnd.n2578 585
R2400 gnd.n2586 gnd.n2578 585
R2401 gnd.n2961 gnd.n2960 585
R2402 gnd.n2960 gnd.n2959 585
R2403 gnd.n2582 gnd.n2581 585
R2404 gnd.n2949 gnd.n2582 585
R2405 gnd.n2936 gnd.n2606 585
R2406 gnd.n2606 gnd.n2605 585
R2407 gnd.n2938 gnd.n2937 585
R2408 gnd.n2939 gnd.n2938 585
R2409 gnd.n2607 gnd.n2604 585
R2410 gnd.n2614 gnd.n2604 585
R2411 gnd.n2931 gnd.n2930 585
R2412 gnd.n2930 gnd.n2929 585
R2413 gnd.n2610 gnd.n2609 585
R2414 gnd.n2918 gnd.n2610 585
R2415 gnd.n2905 gnd.n2631 585
R2416 gnd.n2631 gnd.n2630 585
R2417 gnd.n2907 gnd.n2906 585
R2418 gnd.n2908 gnd.n2907 585
R2419 gnd.n2901 gnd.n2629 585
R2420 gnd.n2900 gnd.n2899 585
R2421 gnd.n2634 gnd.n2633 585
R2422 gnd.n2897 gnd.n2634 585
R2423 gnd.n2656 gnd.n2655 585
R2424 gnd.n2659 gnd.n2658 585
R2425 gnd.n2657 gnd.n2652 585
R2426 gnd.n2664 gnd.n2663 585
R2427 gnd.n2666 gnd.n2665 585
R2428 gnd.n2669 gnd.n2668 585
R2429 gnd.n2667 gnd.n2650 585
R2430 gnd.n2674 gnd.n2673 585
R2431 gnd.n2676 gnd.n2675 585
R2432 gnd.n2679 gnd.n2678 585
R2433 gnd.n2677 gnd.n2648 585
R2434 gnd.n2684 gnd.n2683 585
R2435 gnd.n2688 gnd.n2685 585
R2436 gnd.n2689 gnd.n2626 585
R2437 gnd.n3567 gnd.n2243 585
R2438 gnd.n3634 gnd.n3633 585
R2439 gnd.n3636 gnd.n3635 585
R2440 gnd.n3638 gnd.n3637 585
R2441 gnd.n3640 gnd.n3639 585
R2442 gnd.n3642 gnd.n3641 585
R2443 gnd.n3644 gnd.n3643 585
R2444 gnd.n3646 gnd.n3645 585
R2445 gnd.n3648 gnd.n3647 585
R2446 gnd.n3650 gnd.n3649 585
R2447 gnd.n3652 gnd.n3651 585
R2448 gnd.n3654 gnd.n3653 585
R2449 gnd.n3656 gnd.n3655 585
R2450 gnd.n3659 gnd.n3658 585
R2451 gnd.n3657 gnd.n2231 585
R2452 gnd.n3663 gnd.n2229 585
R2453 gnd.n3665 gnd.n3664 585
R2454 gnd.n3666 gnd.n3665 585
R2455 gnd.n3568 gnd.n2284 585
R2456 gnd.n3568 gnd.n2205 585
R2457 gnd.n3570 gnd.n3569 585
R2458 gnd.n3569 gnd.n2279 585
R2459 gnd.n3566 gnd.n2283 585
R2460 gnd.n3566 gnd.n3565 585
R2461 gnd.n3545 gnd.n2285 585
R2462 gnd.n2297 gnd.n2285 585
R2463 gnd.n3544 gnd.n2295 585
R2464 gnd.n3553 gnd.n2295 585
R2465 gnd.n3279 gnd.n2302 585
R2466 gnd.n3280 gnd.n3279 585
R2467 gnd.n3278 gnd.n3277 585
R2468 gnd.n3278 gnd.n2306 585
R2469 gnd.n3276 gnd.n2308 585
R2470 gnd.n3269 gnd.n2308 585
R2471 gnd.n2321 gnd.n2309 585
R2472 gnd.n2321 gnd.n2313 585
R2473 gnd.n3225 gnd.n2322 585
R2474 gnd.n3259 gnd.n2322 585
R2475 gnd.n3224 gnd.n3223 585
R2476 gnd.n3223 gnd.n2329 585
R2477 gnd.n3222 gnd.n2337 585
R2478 gnd.n3222 gnd.n2328 585
R2479 gnd.n3221 gnd.n2339 585
R2480 gnd.n3221 gnd.n3220 585
R2481 gnd.n3200 gnd.n2338 585
R2482 gnd.n2351 gnd.n2338 585
R2483 gnd.n3199 gnd.n2349 585
R2484 gnd.n3210 gnd.n2349 585
R2485 gnd.n3190 gnd.n2356 585
R2486 gnd.n3191 gnd.n3190 585
R2487 gnd.n3189 gnd.n3188 585
R2488 gnd.n3189 gnd.n2360 585
R2489 gnd.n3187 gnd.n2362 585
R2490 gnd.n3180 gnd.n2362 585
R2491 gnd.n2377 gnd.n2363 585
R2492 gnd.n2377 gnd.n2367 585
R2493 gnd.n3140 gnd.n2378 585
R2494 gnd.n3170 gnd.n2378 585
R2495 gnd.n3139 gnd.n3138 585
R2496 gnd.n3138 gnd.n2385 585
R2497 gnd.n3137 gnd.n2392 585
R2498 gnd.n3137 gnd.n2384 585
R2499 gnd.n3136 gnd.n2394 585
R2500 gnd.n3136 gnd.n3135 585
R2501 gnd.n3115 gnd.n2393 585
R2502 gnd.n2406 gnd.n2393 585
R2503 gnd.n3114 gnd.n2404 585
R2504 gnd.n3125 gnd.n2404 585
R2505 gnd.n3105 gnd.n2411 585
R2506 gnd.n3106 gnd.n3105 585
R2507 gnd.n3104 gnd.n3103 585
R2508 gnd.n3104 gnd.n2415 585
R2509 gnd.n3102 gnd.n2417 585
R2510 gnd.n3095 gnd.n2417 585
R2511 gnd.n3082 gnd.n2418 585
R2512 gnd.n3083 gnd.n3082 585
R2513 gnd.n3035 gnd.n2431 585
R2514 gnd.n3085 gnd.n2431 585
R2515 gnd.n3037 gnd.n3036 585
R2516 gnd.n3038 gnd.n3037 585
R2517 gnd.n3030 gnd.n2533 585
R2518 gnd.n2533 gnd.n2532 585
R2519 gnd.n3028 gnd.n3027 585
R2520 gnd.n3027 gnd.n2514 585
R2521 gnd.n3025 gnd.n2512 585
R2522 gnd.n3046 gnd.n2512 585
R2523 gnd.n2543 gnd.n2542 585
R2524 gnd.n2542 gnd.n2541 585
R2525 gnd.n3019 gnd.n2502 585
R2526 gnd.n3052 gnd.n2502 585
R2527 gnd.n3018 gnd.n3017 585
R2528 gnd.n3017 gnd.n3016 585
R2529 gnd.n3014 gnd.n2545 585
R2530 gnd.n3014 gnd.n2492 585
R2531 gnd.n3013 gnd.n3012 585
R2532 gnd.n3013 gnd.n2491 585
R2533 gnd.n2548 gnd.n2547 585
R2534 gnd.n3004 gnd.n2547 585
R2535 gnd.n2972 gnd.n2971 585
R2536 gnd.n2971 gnd.n2552 585
R2537 gnd.n2973 gnd.n2561 585
R2538 gnd.n2990 gnd.n2561 585
R2539 gnd.n2970 gnd.n2969 585
R2540 gnd.n2969 gnd.n2567 585
R2541 gnd.n2968 gnd.n2575 585
R2542 gnd.n2968 gnd.n2967 585
R2543 gnd.n2953 gnd.n2576 585
R2544 gnd.n2586 gnd.n2576 585
R2545 gnd.n2952 gnd.n2584 585
R2546 gnd.n2959 gnd.n2584 585
R2547 gnd.n2951 gnd.n2950 585
R2548 gnd.n2950 gnd.n2949 585
R2549 gnd.n2595 gnd.n2592 585
R2550 gnd.n2605 gnd.n2595 585
R2551 gnd.n2941 gnd.n2940 585
R2552 gnd.n2940 gnd.n2939 585
R2553 gnd.n2601 gnd.n2600 585
R2554 gnd.n2614 gnd.n2601 585
R2555 gnd.n2921 gnd.n2612 585
R2556 gnd.n2929 gnd.n2612 585
R2557 gnd.n2920 gnd.n2919 585
R2558 gnd.n2919 gnd.n2918 585
R2559 gnd.n2621 gnd.n2619 585
R2560 gnd.n2630 gnd.n2621 585
R2561 gnd.n2910 gnd.n2909 585
R2562 gnd.n2909 gnd.n2908 585
R2563 gnd.n4958 gnd.n1799 585
R2564 gnd.n1799 gnd.n1755 585
R2565 gnd.n4960 gnd.n4959 585
R2566 gnd.n4961 gnd.n4960 585
R2567 gnd.n4869 gnd.n1798 585
R2568 gnd.n1805 gnd.n1798 585
R2569 gnd.n4868 gnd.n4867 585
R2570 gnd.n4867 gnd.n4866 585
R2571 gnd.n1801 gnd.n1800 585
R2572 gnd.n1802 gnd.n1801 585
R2573 gnd.n4855 gnd.n4854 585
R2574 gnd.n4856 gnd.n4855 585
R2575 gnd.n4853 gnd.n1814 585
R2576 gnd.n1814 gnd.n1811 585
R2577 gnd.n4852 gnd.n4851 585
R2578 gnd.n4851 gnd.n4850 585
R2579 gnd.n1816 gnd.n1815 585
R2580 gnd.n1824 gnd.n1816 585
R2581 gnd.n4837 gnd.n4836 585
R2582 gnd.n4838 gnd.n4837 585
R2583 gnd.n4835 gnd.n1826 585
R2584 gnd.n1826 gnd.n1823 585
R2585 gnd.n4834 gnd.n4833 585
R2586 gnd.n4833 gnd.n4832 585
R2587 gnd.n1828 gnd.n1827 585
R2588 gnd.n4750 gnd.n1828 585
R2589 gnd.n4818 gnd.n4817 585
R2590 gnd.n4819 gnd.n4818 585
R2591 gnd.n4816 gnd.n1841 585
R2592 gnd.n1841 gnd.n1838 585
R2593 gnd.n4815 gnd.n4814 585
R2594 gnd.n4814 gnd.n4813 585
R2595 gnd.n1843 gnd.n1842 585
R2596 gnd.n1844 gnd.n1843 585
R2597 gnd.n4762 gnd.n1865 585
R2598 gnd.n4762 gnd.n4761 585
R2599 gnd.n4764 gnd.n4763 585
R2600 gnd.n4763 gnd.n1852 585
R2601 gnd.n4765 gnd.n1863 585
R2602 gnd.n4745 gnd.n1863 585
R2603 gnd.n4767 gnd.n4766 585
R2604 gnd.n4768 gnd.n4767 585
R2605 gnd.n1864 gnd.n1862 585
R2606 gnd.n1862 gnd.n1859 585
R2607 gnd.n4737 gnd.n4736 585
R2608 gnd.n4738 gnd.n4737 585
R2609 gnd.n4735 gnd.n1871 585
R2610 gnd.n1876 gnd.n1871 585
R2611 gnd.n4734 gnd.n4733 585
R2612 gnd.n4733 gnd.n4732 585
R2613 gnd.n1873 gnd.n1872 585
R2614 gnd.n1884 gnd.n1873 585
R2615 gnd.n4721 gnd.n4720 585
R2616 gnd.n4722 gnd.n4721 585
R2617 gnd.n4719 gnd.n1885 585
R2618 gnd.n4714 gnd.n1885 585
R2619 gnd.n4718 gnd.n4717 585
R2620 gnd.n4717 gnd.n4716 585
R2621 gnd.n1887 gnd.n1886 585
R2622 gnd.n1888 gnd.n1887 585
R2623 gnd.n4701 gnd.n4700 585
R2624 gnd.n4702 gnd.n4701 585
R2625 gnd.n4699 gnd.n1896 585
R2626 gnd.n4695 gnd.n1896 585
R2627 gnd.n4698 gnd.n4697 585
R2628 gnd.n4697 gnd.n4696 585
R2629 gnd.n1898 gnd.n1897 585
R2630 gnd.n1904 gnd.n1898 585
R2631 gnd.n4687 gnd.n4686 585
R2632 gnd.n4688 gnd.n4687 585
R2633 gnd.n4685 gnd.n1906 585
R2634 gnd.n1906 gnd.n1903 585
R2635 gnd.n4684 gnd.n4683 585
R2636 gnd.n4683 gnd.n4682 585
R2637 gnd.n1908 gnd.n1907 585
R2638 gnd.n4581 gnd.n1908 585
R2639 gnd.n4660 gnd.n4659 585
R2640 gnd.n4661 gnd.n4660 585
R2641 gnd.n4658 gnd.n1922 585
R2642 gnd.n1922 gnd.n1919 585
R2643 gnd.n4657 gnd.n4656 585
R2644 gnd.n4656 gnd.n4655 585
R2645 gnd.n1924 gnd.n1923 585
R2646 gnd.n4589 gnd.n1924 585
R2647 gnd.n1948 gnd.n1947 585
R2648 gnd.n1948 gnd.n1932 585
R2649 gnd.n4597 gnd.n4596 585
R2650 gnd.n4596 gnd.n4595 585
R2651 gnd.n4598 gnd.n1945 585
R2652 gnd.n1945 gnd.n1943 585
R2653 gnd.n4600 gnd.n4599 585
R2654 gnd.n4601 gnd.n4600 585
R2655 gnd.n1946 gnd.n1944 585
R2656 gnd.n1944 gnd.n1940 585
R2657 gnd.n4573 gnd.n4572 585
R2658 gnd.n4574 gnd.n4573 585
R2659 gnd.n4571 gnd.n1954 585
R2660 gnd.n1960 gnd.n1954 585
R2661 gnd.n4570 gnd.n4569 585
R2662 gnd.n4569 gnd.n4568 585
R2663 gnd.n1956 gnd.n1955 585
R2664 gnd.n4512 gnd.n1956 585
R2665 gnd.n4557 gnd.n4556 585
R2666 gnd.n4558 gnd.n4557 585
R2667 gnd.n4555 gnd.n1971 585
R2668 gnd.n1971 gnd.n1968 585
R2669 gnd.n4554 gnd.n4553 585
R2670 gnd.n4553 gnd.n4552 585
R2671 gnd.n1973 gnd.n1972 585
R2672 gnd.n4521 gnd.n1973 585
R2673 gnd.n4525 gnd.n4524 585
R2674 gnd.n4524 gnd.n4523 585
R2675 gnd.n4526 gnd.n4434 585
R2676 gnd.n4434 gnd.n1213 585
R2677 gnd.n4528 gnd.n4527 585
R2678 gnd.n4529 gnd.n4528 585
R2679 gnd.n1200 gnd.n1199 585
R2680 gnd.t87 gnd.n1200 585
R2681 gnd.n5680 gnd.n5679 585
R2682 gnd.n5679 gnd.n5678 585
R2683 gnd.n5681 gnd.n1178 585
R2684 gnd.n1201 gnd.n1178 585
R2685 gnd.n5746 gnd.n5745 585
R2686 gnd.n5744 gnd.n1177 585
R2687 gnd.n5743 gnd.n1176 585
R2688 gnd.n5748 gnd.n1176 585
R2689 gnd.n5742 gnd.n5741 585
R2690 gnd.n5740 gnd.n5739 585
R2691 gnd.n5738 gnd.n5737 585
R2692 gnd.n5736 gnd.n5735 585
R2693 gnd.n5734 gnd.n5733 585
R2694 gnd.n5732 gnd.n5731 585
R2695 gnd.n5730 gnd.n5729 585
R2696 gnd.n5728 gnd.n5727 585
R2697 gnd.n5726 gnd.n5725 585
R2698 gnd.n5724 gnd.n5723 585
R2699 gnd.n5722 gnd.n5721 585
R2700 gnd.n5720 gnd.n5719 585
R2701 gnd.n5718 gnd.n5717 585
R2702 gnd.n5716 gnd.n5715 585
R2703 gnd.n5714 gnd.n5713 585
R2704 gnd.n5712 gnd.n5711 585
R2705 gnd.n5710 gnd.n5709 585
R2706 gnd.n5708 gnd.n5707 585
R2707 gnd.n5706 gnd.n5705 585
R2708 gnd.n5704 gnd.n5703 585
R2709 gnd.n5702 gnd.n5701 585
R2710 gnd.n5700 gnd.n5699 585
R2711 gnd.n5698 gnd.n5697 585
R2712 gnd.n5696 gnd.n5695 585
R2713 gnd.n5694 gnd.n5693 585
R2714 gnd.n5692 gnd.n5691 585
R2715 gnd.n5690 gnd.n5689 585
R2716 gnd.n5688 gnd.n5687 585
R2717 gnd.n5686 gnd.n1140 585
R2718 gnd.n5751 gnd.n5750 585
R2719 gnd.n1142 gnd.n1139 585
R2720 gnd.n4439 gnd.n4438 585
R2721 gnd.n4441 gnd.n4440 585
R2722 gnd.n4444 gnd.n4443 585
R2723 gnd.n4446 gnd.n4445 585
R2724 gnd.n4448 gnd.n4447 585
R2725 gnd.n4450 gnd.n4449 585
R2726 gnd.n4452 gnd.n4451 585
R2727 gnd.n4454 gnd.n4453 585
R2728 gnd.n4456 gnd.n4455 585
R2729 gnd.n4458 gnd.n4457 585
R2730 gnd.n4460 gnd.n4459 585
R2731 gnd.n4462 gnd.n4461 585
R2732 gnd.n4464 gnd.n4463 585
R2733 gnd.n4466 gnd.n4465 585
R2734 gnd.n4468 gnd.n4467 585
R2735 gnd.n4470 gnd.n4469 585
R2736 gnd.n4472 gnd.n4471 585
R2737 gnd.n4474 gnd.n4473 585
R2738 gnd.n4476 gnd.n4475 585
R2739 gnd.n4478 gnd.n4477 585
R2740 gnd.n4480 gnd.n4479 585
R2741 gnd.n4482 gnd.n4481 585
R2742 gnd.n4484 gnd.n4483 585
R2743 gnd.n4486 gnd.n4485 585
R2744 gnd.n4488 gnd.n4487 585
R2745 gnd.n4490 gnd.n4489 585
R2746 gnd.n4492 gnd.n4491 585
R2747 gnd.n4494 gnd.n4493 585
R2748 gnd.n4496 gnd.n4495 585
R2749 gnd.n4498 gnd.n4497 585
R2750 gnd.n4500 gnd.n4499 585
R2751 gnd.n4965 gnd.n4964 585
R2752 gnd.n4967 gnd.n4966 585
R2753 gnd.n4969 gnd.n4968 585
R2754 gnd.n4971 gnd.n4970 585
R2755 gnd.n4973 gnd.n4972 585
R2756 gnd.n4975 gnd.n4974 585
R2757 gnd.n4977 gnd.n4976 585
R2758 gnd.n4979 gnd.n4978 585
R2759 gnd.n4981 gnd.n4980 585
R2760 gnd.n4983 gnd.n4982 585
R2761 gnd.n4985 gnd.n4984 585
R2762 gnd.n4987 gnd.n4986 585
R2763 gnd.n4989 gnd.n4988 585
R2764 gnd.n4991 gnd.n4990 585
R2765 gnd.n4993 gnd.n4992 585
R2766 gnd.n4995 gnd.n4994 585
R2767 gnd.n4997 gnd.n4996 585
R2768 gnd.n4999 gnd.n4998 585
R2769 gnd.n5001 gnd.n5000 585
R2770 gnd.n5003 gnd.n5002 585
R2771 gnd.n5005 gnd.n5004 585
R2772 gnd.n5007 gnd.n5006 585
R2773 gnd.n5009 gnd.n5008 585
R2774 gnd.n5011 gnd.n5010 585
R2775 gnd.n5013 gnd.n5012 585
R2776 gnd.n5015 gnd.n5014 585
R2777 gnd.n5017 gnd.n5016 585
R2778 gnd.n5019 gnd.n5018 585
R2779 gnd.n5021 gnd.n5020 585
R2780 gnd.n5024 gnd.n5023 585
R2781 gnd.n5026 gnd.n5025 585
R2782 gnd.n5028 gnd.n5027 585
R2783 gnd.n5030 gnd.n5029 585
R2784 gnd.n4891 gnd.n1448 585
R2785 gnd.n4893 gnd.n4892 585
R2786 gnd.n4895 gnd.n4894 585
R2787 gnd.n4897 gnd.n4896 585
R2788 gnd.n4900 gnd.n4899 585
R2789 gnd.n4902 gnd.n4901 585
R2790 gnd.n4904 gnd.n4903 585
R2791 gnd.n4906 gnd.n4905 585
R2792 gnd.n4908 gnd.n4907 585
R2793 gnd.n4910 gnd.n4909 585
R2794 gnd.n4912 gnd.n4911 585
R2795 gnd.n4914 gnd.n4913 585
R2796 gnd.n4916 gnd.n4915 585
R2797 gnd.n4918 gnd.n4917 585
R2798 gnd.n4920 gnd.n4919 585
R2799 gnd.n4922 gnd.n4921 585
R2800 gnd.n4924 gnd.n4923 585
R2801 gnd.n4926 gnd.n4925 585
R2802 gnd.n4928 gnd.n4927 585
R2803 gnd.n4930 gnd.n4929 585
R2804 gnd.n4932 gnd.n4931 585
R2805 gnd.n4934 gnd.n4933 585
R2806 gnd.n4936 gnd.n4935 585
R2807 gnd.n4938 gnd.n4937 585
R2808 gnd.n4940 gnd.n4939 585
R2809 gnd.n4942 gnd.n4941 585
R2810 gnd.n4944 gnd.n4943 585
R2811 gnd.n4946 gnd.n4945 585
R2812 gnd.n4948 gnd.n4947 585
R2813 gnd.n4950 gnd.n4949 585
R2814 gnd.n4952 gnd.n4951 585
R2815 gnd.n4954 gnd.n4953 585
R2816 gnd.n4956 gnd.n4955 585
R2817 gnd.n4963 gnd.n1793 585
R2818 gnd.n4963 gnd.n1755 585
R2819 gnd.n4962 gnd.n1795 585
R2820 gnd.n4962 gnd.n4961 585
R2821 gnd.n4842 gnd.n1794 585
R2822 gnd.n1805 gnd.n1794 585
R2823 gnd.n4843 gnd.n1803 585
R2824 gnd.n4866 gnd.n1803 585
R2825 gnd.n4845 gnd.n4844 585
R2826 gnd.n4844 gnd.n1802 585
R2827 gnd.n4846 gnd.n1813 585
R2828 gnd.n4856 gnd.n1813 585
R2829 gnd.n4847 gnd.n1820 585
R2830 gnd.n1820 gnd.n1811 585
R2831 gnd.n4849 gnd.n4848 585
R2832 gnd.n4850 gnd.n4849 585
R2833 gnd.n4841 gnd.n1819 585
R2834 gnd.n1824 gnd.n1819 585
R2835 gnd.n4840 gnd.n4839 585
R2836 gnd.n4839 gnd.n4838 585
R2837 gnd.n1822 gnd.n1821 585
R2838 gnd.n1823 gnd.n1822 585
R2839 gnd.n4749 gnd.n1830 585
R2840 gnd.n4832 gnd.n1830 585
R2841 gnd.n4752 gnd.n4751 585
R2842 gnd.n4751 gnd.n4750 585
R2843 gnd.n4753 gnd.n1840 585
R2844 gnd.n4819 gnd.n1840 585
R2845 gnd.n4755 gnd.n4754 585
R2846 gnd.n4754 gnd.n1838 585
R2847 gnd.n4756 gnd.n1845 585
R2848 gnd.n4813 gnd.n1845 585
R2849 gnd.n4757 gnd.n1867 585
R2850 gnd.n1867 gnd.n1844 585
R2851 gnd.n4759 gnd.n4758 585
R2852 gnd.n4761 gnd.n4759 585
R2853 gnd.n4748 gnd.n1866 585
R2854 gnd.n1866 gnd.n1852 585
R2855 gnd.n4747 gnd.n4746 585
R2856 gnd.n4746 gnd.n4745 585
R2857 gnd.n4742 gnd.n1861 585
R2858 gnd.n4768 gnd.n1861 585
R2859 gnd.n4741 gnd.n4740 585
R2860 gnd.n4740 gnd.n1859 585
R2861 gnd.n4739 gnd.n1868 585
R2862 gnd.n4739 gnd.n4738 585
R2863 gnd.n4707 gnd.n1869 585
R2864 gnd.n1876 gnd.n1869 585
R2865 gnd.n4708 gnd.n1874 585
R2866 gnd.n4732 gnd.n1874 585
R2867 gnd.n4710 gnd.n4709 585
R2868 gnd.n4709 gnd.n1884 585
R2869 gnd.n4711 gnd.n1883 585
R2870 gnd.n4722 gnd.n1883 585
R2871 gnd.n4713 gnd.n4712 585
R2872 gnd.n4714 gnd.n4713 585
R2873 gnd.n4706 gnd.n1889 585
R2874 gnd.n4716 gnd.n1889 585
R2875 gnd.n4705 gnd.n4704 585
R2876 gnd.n4704 gnd.n1888 585
R2877 gnd.n4703 gnd.n1891 585
R2878 gnd.n4703 gnd.n4702 585
R2879 gnd.n4692 gnd.n1892 585
R2880 gnd.n4695 gnd.n1892 585
R2881 gnd.n4694 gnd.n4693 585
R2882 gnd.n4696 gnd.n4694 585
R2883 gnd.n4691 gnd.n1900 585
R2884 gnd.n1904 gnd.n1900 585
R2885 gnd.n4690 gnd.n4689 585
R2886 gnd.n4689 gnd.n4688 585
R2887 gnd.n1902 gnd.n1901 585
R2888 gnd.n1903 gnd.n1902 585
R2889 gnd.n4580 gnd.n1911 585
R2890 gnd.n4682 gnd.n1911 585
R2891 gnd.n4583 gnd.n4582 585
R2892 gnd.n4582 gnd.n4581 585
R2893 gnd.n4584 gnd.n1921 585
R2894 gnd.n4661 gnd.n1921 585
R2895 gnd.n4586 gnd.n4585 585
R2896 gnd.n4585 gnd.n1919 585
R2897 gnd.n4587 gnd.n1925 585
R2898 gnd.n4655 gnd.n1925 585
R2899 gnd.n4591 gnd.n4590 585
R2900 gnd.n4590 gnd.n4589 585
R2901 gnd.n4592 gnd.n1951 585
R2902 gnd.n1951 gnd.n1932 585
R2903 gnd.n4594 gnd.n4593 585
R2904 gnd.n4595 gnd.n4594 585
R2905 gnd.n4579 gnd.n1950 585
R2906 gnd.n1950 gnd.n1943 585
R2907 gnd.n4578 gnd.n1942 585
R2908 gnd.n4601 gnd.n1942 585
R2909 gnd.n4577 gnd.n4576 585
R2910 gnd.n4576 gnd.n1940 585
R2911 gnd.n4575 gnd.n1952 585
R2912 gnd.n4575 gnd.n4574 585
R2913 gnd.n4510 gnd.n1953 585
R2914 gnd.n1960 gnd.n1953 585
R2915 gnd.n4511 gnd.n1958 585
R2916 gnd.n4568 gnd.n1958 585
R2917 gnd.n4514 gnd.n4513 585
R2918 gnd.n4513 gnd.n4512 585
R2919 gnd.n4515 gnd.n1970 585
R2920 gnd.n4558 gnd.n1970 585
R2921 gnd.n4517 gnd.n4516 585
R2922 gnd.n4516 gnd.n1968 585
R2923 gnd.n4518 gnd.n1974 585
R2924 gnd.n4552 gnd.n1974 585
R2925 gnd.n4520 gnd.n4519 585
R2926 gnd.n4521 gnd.n4520 585
R2927 gnd.n4509 gnd.n4435 585
R2928 gnd.n4523 gnd.n4435 585
R2929 gnd.n4508 gnd.n4507 585
R2930 gnd.n4507 gnd.n1213 585
R2931 gnd.n4506 gnd.n4433 585
R2932 gnd.n4529 gnd.n4433 585
R2933 gnd.n4505 gnd.n4504 585
R2934 gnd.n4504 gnd.t87 585
R2935 gnd.n4503 gnd.n1202 585
R2936 gnd.n5678 gnd.n1202 585
R2937 gnd.n4502 gnd.n4501 585
R2938 gnd.n4501 gnd.n1201 585
R2939 gnd.n5887 gnd.n5886 585
R2940 gnd.n5886 gnd.n5885 585
R2941 gnd.n5888 gnd.n853 585
R2942 gnd.n5878 gnd.n853 585
R2943 gnd.n5890 gnd.n5889 585
R2944 gnd.n5891 gnd.n5890 585
R2945 gnd.n839 gnd.n838 585
R2946 gnd.n4188 gnd.n839 585
R2947 gnd.n5899 gnd.n5898 585
R2948 gnd.n5898 gnd.n5897 585
R2949 gnd.n5900 gnd.n833 585
R2950 gnd.n4182 gnd.n833 585
R2951 gnd.n5902 gnd.n5901 585
R2952 gnd.n5903 gnd.n5902 585
R2953 gnd.n819 gnd.n818 585
R2954 gnd.n4199 gnd.n819 585
R2955 gnd.n5911 gnd.n5910 585
R2956 gnd.n5910 gnd.n5909 585
R2957 gnd.n5912 gnd.n813 585
R2958 gnd.n4175 gnd.n813 585
R2959 gnd.n5914 gnd.n5913 585
R2960 gnd.n5915 gnd.n5914 585
R2961 gnd.n799 gnd.n798 585
R2962 gnd.n4167 gnd.n799 585
R2963 gnd.n5923 gnd.n5922 585
R2964 gnd.n5922 gnd.n5921 585
R2965 gnd.n5924 gnd.n793 585
R2966 gnd.n4161 gnd.n793 585
R2967 gnd.n5926 gnd.n5925 585
R2968 gnd.n5927 gnd.n5926 585
R2969 gnd.n779 gnd.n778 585
R2970 gnd.n4153 gnd.n779 585
R2971 gnd.n5935 gnd.n5934 585
R2972 gnd.n5934 gnd.n5933 585
R2973 gnd.n5936 gnd.n776 585
R2974 gnd.n4109 gnd.n776 585
R2975 gnd.n5939 gnd.n5938 585
R2976 gnd.n5940 gnd.n5939 585
R2977 gnd.n777 gnd.n762 585
R2978 gnd.n4117 gnd.n762 585
R2979 gnd.n5948 gnd.n5947 585
R2980 gnd.n5947 gnd.n5946 585
R2981 gnd.n5949 gnd.n759 585
R2982 gnd.n4098 gnd.n759 585
R2983 gnd.n5952 gnd.n5951 585
R2984 gnd.n5953 gnd.n5952 585
R2985 gnd.n760 gnd.n743 585
R2986 gnd.n4090 gnd.n743 585
R2987 gnd.n5961 gnd.n5960 585
R2988 gnd.n5960 gnd.n5959 585
R2989 gnd.n5962 gnd.n739 585
R2990 gnd.n4072 gnd.n739 585
R2991 gnd.n5965 gnd.n5964 585
R2992 gnd.n5966 gnd.n5965 585
R2993 gnd.n740 gnd.n738 585
R2994 gnd.n738 gnd.n733 585
R2995 gnd.n4062 gnd.n4061 585
R2996 gnd.n4063 gnd.n4062 585
R2997 gnd.n2138 gnd.n2137 585
R2998 gnd.n2144 gnd.n2137 585
R2999 gnd.n4056 gnd.n4055 585
R3000 gnd.n4055 gnd.n4054 585
R3001 gnd.n2141 gnd.n2140 585
R3002 gnd.n4036 gnd.n2141 585
R3003 gnd.n4021 gnd.n2164 585
R3004 gnd.n2164 gnd.n2154 585
R3005 gnd.n4023 gnd.n4022 585
R3006 gnd.n4024 gnd.n4023 585
R3007 gnd.n2165 gnd.n2163 585
R3008 gnd.n2163 gnd.n2160 585
R3009 gnd.n4016 gnd.n4015 585
R3010 gnd.n4015 gnd.n4014 585
R3011 gnd.n2168 gnd.n2167 585
R3012 gnd.n3999 gnd.n2168 585
R3013 gnd.n3986 gnd.n2189 585
R3014 gnd.n2189 gnd.n2179 585
R3015 gnd.n3988 gnd.n3987 585
R3016 gnd.n3989 gnd.n3988 585
R3017 gnd.n2190 gnd.n2188 585
R3018 gnd.n2188 gnd.n2185 585
R3019 gnd.n3981 gnd.n3980 585
R3020 gnd.n3980 gnd.n3979 585
R3021 gnd.n2193 gnd.n2192 585
R3022 gnd.n3744 gnd.n2193 585
R3023 gnd.n3960 gnd.n3959 585
R3024 gnd.n3961 gnd.n3960 585
R3025 gnd.n3956 gnd.n3745 585
R3026 gnd.n3955 gnd.n3954 585
R3027 gnd.n3952 gnd.n3747 585
R3028 gnd.n3952 gnd.n3667 585
R3029 gnd.n3951 gnd.n3950 585
R3030 gnd.n3949 gnd.n3948 585
R3031 gnd.n3947 gnd.n3752 585
R3032 gnd.n3945 gnd.n3944 585
R3033 gnd.n3943 gnd.n3753 585
R3034 gnd.n3942 gnd.n3941 585
R3035 gnd.n3939 gnd.n3758 585
R3036 gnd.n3937 gnd.n3936 585
R3037 gnd.n3935 gnd.n3759 585
R3038 gnd.n3934 gnd.n3933 585
R3039 gnd.n3931 gnd.n3764 585
R3040 gnd.n3929 gnd.n3928 585
R3041 gnd.n3927 gnd.n3765 585
R3042 gnd.n3926 gnd.n3925 585
R3043 gnd.n3923 gnd.n3770 585
R3044 gnd.n3921 gnd.n3920 585
R3045 gnd.n3919 gnd.n3771 585
R3046 gnd.n3918 gnd.n3917 585
R3047 gnd.n3915 gnd.n3779 585
R3048 gnd.n3913 gnd.n3912 585
R3049 gnd.n3911 gnd.n3780 585
R3050 gnd.n3910 gnd.n3909 585
R3051 gnd.n3907 gnd.n3785 585
R3052 gnd.n3905 gnd.n3904 585
R3053 gnd.n3903 gnd.n3786 585
R3054 gnd.n3902 gnd.n3901 585
R3055 gnd.n3899 gnd.n3791 585
R3056 gnd.n3897 gnd.n3896 585
R3057 gnd.n3895 gnd.n3792 585
R3058 gnd.n3894 gnd.n3893 585
R3059 gnd.n3891 gnd.n3797 585
R3060 gnd.n3889 gnd.n3888 585
R3061 gnd.n3887 gnd.n3798 585
R3062 gnd.n3886 gnd.n3885 585
R3063 gnd.n3883 gnd.n3805 585
R3064 gnd.n3881 gnd.n3880 585
R3065 gnd.n3879 gnd.n3806 585
R3066 gnd.n3878 gnd.n3877 585
R3067 gnd.n3875 gnd.n3811 585
R3068 gnd.n3873 gnd.n3872 585
R3069 gnd.n3871 gnd.n3812 585
R3070 gnd.n3870 gnd.n3869 585
R3071 gnd.n3867 gnd.n3817 585
R3072 gnd.n3865 gnd.n3864 585
R3073 gnd.n3863 gnd.n3818 585
R3074 gnd.n3862 gnd.n3861 585
R3075 gnd.n3859 gnd.n3823 585
R3076 gnd.n3857 gnd.n3856 585
R3077 gnd.n3855 gnd.n3824 585
R3078 gnd.n3854 gnd.n3853 585
R3079 gnd.n3851 gnd.n3829 585
R3080 gnd.n3849 gnd.n3848 585
R3081 gnd.n3847 gnd.n3830 585
R3082 gnd.n3846 gnd.n3845 585
R3083 gnd.n3843 gnd.n3837 585
R3084 gnd.n3841 gnd.n3840 585
R3085 gnd.n1070 gnd.n1069 585
R3086 gnd.n1076 gnd.n1075 585
R3087 gnd.n1078 gnd.n1077 585
R3088 gnd.n1080 gnd.n1079 585
R3089 gnd.n1082 gnd.n1081 585
R3090 gnd.n1084 gnd.n1083 585
R3091 gnd.n1086 gnd.n1085 585
R3092 gnd.n1088 gnd.n1087 585
R3093 gnd.n1090 gnd.n1089 585
R3094 gnd.n1092 gnd.n1091 585
R3095 gnd.n1094 gnd.n1093 585
R3096 gnd.n1096 gnd.n1095 585
R3097 gnd.n1098 gnd.n1097 585
R3098 gnd.n1100 gnd.n1099 585
R3099 gnd.n1102 gnd.n1101 585
R3100 gnd.n1104 gnd.n1103 585
R3101 gnd.n1106 gnd.n1105 585
R3102 gnd.n1108 gnd.n1107 585
R3103 gnd.n1110 gnd.n1109 585
R3104 gnd.n1113 gnd.n1112 585
R3105 gnd.n1111 gnd.n1049 585
R3106 gnd.n1118 gnd.n1117 585
R3107 gnd.n1120 gnd.n1119 585
R3108 gnd.n1122 gnd.n1121 585
R3109 gnd.n1124 gnd.n1123 585
R3110 gnd.n1126 gnd.n1125 585
R3111 gnd.n1128 gnd.n1127 585
R3112 gnd.n1130 gnd.n1129 585
R3113 gnd.n1132 gnd.n1131 585
R3114 gnd.n1135 gnd.n1134 585
R3115 gnd.n1133 gnd.n1040 585
R3116 gnd.n5754 gnd.n5753 585
R3117 gnd.n5756 gnd.n5755 585
R3118 gnd.n5758 gnd.n5757 585
R3119 gnd.n5760 gnd.n5759 585
R3120 gnd.n5762 gnd.n5761 585
R3121 gnd.n5764 gnd.n5763 585
R3122 gnd.n5766 gnd.n5765 585
R3123 gnd.n5768 gnd.n5767 585
R3124 gnd.n5771 gnd.n5770 585
R3125 gnd.n5773 gnd.n5772 585
R3126 gnd.n5775 gnd.n5774 585
R3127 gnd.n5777 gnd.n5776 585
R3128 gnd.n5779 gnd.n5778 585
R3129 gnd.n5781 gnd.n5780 585
R3130 gnd.n5783 gnd.n5782 585
R3131 gnd.n5785 gnd.n5784 585
R3132 gnd.n5787 gnd.n5786 585
R3133 gnd.n5789 gnd.n5788 585
R3134 gnd.n5791 gnd.n5790 585
R3135 gnd.n5793 gnd.n5792 585
R3136 gnd.n5795 gnd.n5794 585
R3137 gnd.n5797 gnd.n5796 585
R3138 gnd.n5798 gnd.n1009 585
R3139 gnd.n5800 gnd.n5799 585
R3140 gnd.n1010 gnd.n1008 585
R3141 gnd.n1011 gnd.n858 585
R3142 gnd.n5802 gnd.n858 585
R3143 gnd.n5881 gnd.n860 585
R3144 gnd.n5885 gnd.n860 585
R3145 gnd.n5880 gnd.n5879 585
R3146 gnd.n5879 gnd.n5878 585
R3147 gnd.n866 gnd.n851 585
R3148 gnd.n5891 gnd.n851 585
R3149 gnd.n4187 gnd.n4186 585
R3150 gnd.n4188 gnd.n4187 585
R3151 gnd.n4185 gnd.n841 585
R3152 gnd.n5897 gnd.n841 585
R3153 gnd.n4184 gnd.n4183 585
R3154 gnd.n4183 gnd.n4182 585
R3155 gnd.n4180 gnd.n830 585
R3156 gnd.n5903 gnd.n830 585
R3157 gnd.n4179 gnd.n2095 585
R3158 gnd.n4199 gnd.n2095 585
R3159 gnd.n4178 gnd.n821 585
R3160 gnd.n5909 gnd.n821 585
R3161 gnd.n4177 gnd.n4176 585
R3162 gnd.n4176 gnd.n4175 585
R3163 gnd.n2101 gnd.n810 585
R3164 gnd.n5915 gnd.n810 585
R3165 gnd.n4166 gnd.n4165 585
R3166 gnd.n4167 gnd.n4166 585
R3167 gnd.n4164 gnd.n801 585
R3168 gnd.n5921 gnd.n801 585
R3169 gnd.n4163 gnd.n4162 585
R3170 gnd.n4162 gnd.n4161 585
R3171 gnd.n2107 gnd.n790 585
R3172 gnd.n5927 gnd.n790 585
R3173 gnd.n4105 gnd.n2112 585
R3174 gnd.n4153 gnd.n2112 585
R3175 gnd.n4106 gnd.n781 585
R3176 gnd.n5933 gnd.n781 585
R3177 gnd.n4108 gnd.n4107 585
R3178 gnd.n4109 gnd.n4108 585
R3179 gnd.n4103 gnd.n773 585
R3180 gnd.n5940 gnd.n773 585
R3181 gnd.n4102 gnd.n2119 585
R3182 gnd.n4117 gnd.n2119 585
R3183 gnd.n4101 gnd.n764 585
R3184 gnd.n5946 gnd.n764 585
R3185 gnd.n4100 gnd.n4099 585
R3186 gnd.n4099 gnd.n4098 585
R3187 gnd.n2123 gnd.n756 585
R3188 gnd.n5953 gnd.n756 585
R3189 gnd.n4077 gnd.n4076 585
R3190 gnd.n4090 gnd.n4077 585
R3191 gnd.n4075 gnd.n745 585
R3192 gnd.n5959 gnd.n745 585
R3193 gnd.n4074 gnd.n4073 585
R3194 gnd.n4073 gnd.n4072 585
R3195 gnd.n2128 gnd.n734 585
R3196 gnd.n5966 gnd.n734 585
R3197 gnd.n4044 gnd.n4043 585
R3198 gnd.n4043 gnd.n733 585
R3199 gnd.n4042 gnd.n2135 585
R3200 gnd.n4063 gnd.n2135 585
R3201 gnd.n4041 gnd.n4040 585
R3202 gnd.n4040 gnd.n2144 585
R3203 gnd.n4039 gnd.n2142 585
R3204 gnd.n4054 gnd.n2142 585
R3205 gnd.n4038 gnd.n4037 585
R3206 gnd.n4037 gnd.n4036 585
R3207 gnd.n2153 gnd.n2151 585
R3208 gnd.n2154 gnd.n2153 585
R3209 gnd.n4005 gnd.n2161 585
R3210 gnd.n4024 gnd.n2161 585
R3211 gnd.n4004 gnd.n4003 585
R3212 gnd.n4003 gnd.n2160 585
R3213 gnd.n4002 gnd.n2169 585
R3214 gnd.n4014 gnd.n2169 585
R3215 gnd.n4001 gnd.n4000 585
R3216 gnd.n4000 gnd.n3999 585
R3217 gnd.n2178 gnd.n2176 585
R3218 gnd.n2179 gnd.n2178 585
R3219 gnd.n3970 gnd.n2186 585
R3220 gnd.n3989 gnd.n2186 585
R3221 gnd.n3969 gnd.n3968 585
R3222 gnd.n3968 gnd.n2185 585
R3223 gnd.n3967 gnd.n2194 585
R3224 gnd.n3979 gnd.n2194 585
R3225 gnd.n3966 gnd.n2202 585
R3226 gnd.n3744 gnd.n2202 585
R3227 gnd.n3668 gnd.n2201 585
R3228 gnd.n3961 gnd.n3668 585
R3229 gnd.n7149 gnd.n7148 585
R3230 gnd.n7148 gnd.n7147 585
R3231 gnd.n7150 gnd.n161 585
R3232 gnd.n167 gnd.n161 585
R3233 gnd.n7152 gnd.n7151 585
R3234 gnd.n7153 gnd.n7152 585
R3235 gnd.n149 gnd.n148 585
R3236 gnd.n152 gnd.n149 585
R3237 gnd.n7161 gnd.n7160 585
R3238 gnd.n7160 gnd.n7159 585
R3239 gnd.n7162 gnd.n143 585
R3240 gnd.n143 gnd.n142 585
R3241 gnd.n7164 gnd.n7163 585
R3242 gnd.n7165 gnd.n7164 585
R3243 gnd.n129 gnd.n128 585
R3244 gnd.n133 gnd.n129 585
R3245 gnd.n7173 gnd.n7172 585
R3246 gnd.n7172 gnd.n7171 585
R3247 gnd.n7174 gnd.n123 585
R3248 gnd.n130 gnd.n123 585
R3249 gnd.n7176 gnd.n7175 585
R3250 gnd.n7177 gnd.n7176 585
R3251 gnd.n110 gnd.n109 585
R3252 gnd.n120 gnd.n110 585
R3253 gnd.n7185 gnd.n7184 585
R3254 gnd.n7184 gnd.n7183 585
R3255 gnd.n7186 gnd.n105 585
R3256 gnd.n111 gnd.n105 585
R3257 gnd.n7188 gnd.n7187 585
R3258 gnd.n7189 gnd.n7188 585
R3259 gnd.n89 gnd.n87 585
R3260 gnd.n7116 gnd.n89 585
R3261 gnd.n7197 gnd.n7196 585
R3262 gnd.n7196 gnd.n7195 585
R3263 gnd.n88 gnd.n80 585
R3264 gnd.n6791 gnd.n88 585
R3265 gnd.n7200 gnd.n78 585
R3266 gnd.n6784 gnd.n78 585
R3267 gnd.n7202 gnd.n7201 585
R3268 gnd.n7203 gnd.n7202 585
R3269 gnd.n1593 gnd.n77 585
R3270 gnd.n5306 gnd.n77 585
R3271 gnd.n1595 gnd.n1594 585
R3272 gnd.n1596 gnd.n1595 585
R3273 gnd.n1583 gnd.n1582 585
R3274 gnd.n5297 gnd.n1582 585
R3275 gnd.n5316 gnd.n1584 585
R3276 gnd.n5316 gnd.n5315 585
R3277 gnd.n5319 gnd.n5318 585
R3278 gnd.n5320 gnd.n5319 585
R3279 gnd.n5317 gnd.n1567 585
R3280 gnd.n5288 gnd.n1567 585
R3281 gnd.n5328 gnd.n5327 585
R3282 gnd.n5327 gnd.n5326 585
R3283 gnd.n5329 gnd.n1564 585
R3284 gnd.n5276 gnd.n1564 585
R3285 gnd.n5331 gnd.n5330 585
R3286 gnd.n5332 gnd.n5331 585
R3287 gnd.n1551 gnd.n1550 585
R3288 gnd.n5269 gnd.n1551 585
R3289 gnd.n5340 gnd.n5339 585
R3290 gnd.n5339 gnd.n5338 585
R3291 gnd.n5341 gnd.n1545 585
R3292 gnd.n5261 gnd.n1545 585
R3293 gnd.n5343 gnd.n5342 585
R3294 gnd.n5344 gnd.n5343 585
R3295 gnd.n1530 gnd.n1529 585
R3296 gnd.n5201 gnd.n1530 585
R3297 gnd.n5352 gnd.n5351 585
R3298 gnd.n5351 gnd.n5350 585
R3299 gnd.n5353 gnd.n1524 585
R3300 gnd.n5192 gnd.n1524 585
R3301 gnd.n5355 gnd.n5354 585
R3302 gnd.n5356 gnd.n5355 585
R3303 gnd.n1507 gnd.n1506 585
R3304 gnd.n5186 gnd.n1507 585
R3305 gnd.n5364 gnd.n5363 585
R3306 gnd.n5363 gnd.n5362 585
R3307 gnd.n5365 gnd.n1498 585
R3308 gnd.n5179 gnd.n1498 585
R3309 gnd.n5367 gnd.n5366 585
R3310 gnd.n5368 gnd.n5367 585
R3311 gnd.n1499 gnd.n1497 585
R3312 gnd.n5218 gnd.n1497 585
R3313 gnd.n1500 gnd.n1419 585
R3314 gnd.n5376 gnd.n1419 585
R3315 gnd.n5495 gnd.n5494 585
R3316 gnd.n5493 gnd.n1418 585
R3317 gnd.n5492 gnd.n1417 585
R3318 gnd.n5497 gnd.n1417 585
R3319 gnd.n5491 gnd.n5490 585
R3320 gnd.n5489 gnd.n5488 585
R3321 gnd.n5487 gnd.n5486 585
R3322 gnd.n5485 gnd.n5484 585
R3323 gnd.n5483 gnd.n5482 585
R3324 gnd.n5481 gnd.n5480 585
R3325 gnd.n5479 gnd.n5478 585
R3326 gnd.n5477 gnd.n5476 585
R3327 gnd.n5475 gnd.n5474 585
R3328 gnd.n5473 gnd.n5472 585
R3329 gnd.n5471 gnd.n5470 585
R3330 gnd.n5469 gnd.n5468 585
R3331 gnd.n5467 gnd.n5466 585
R3332 gnd.n5465 gnd.n5464 585
R3333 gnd.n5463 gnd.n5462 585
R3334 gnd.n5460 gnd.n5459 585
R3335 gnd.n5458 gnd.n5457 585
R3336 gnd.n5456 gnd.n5455 585
R3337 gnd.n5454 gnd.n5453 585
R3338 gnd.n5452 gnd.n5451 585
R3339 gnd.n5450 gnd.n5449 585
R3340 gnd.n5448 gnd.n5447 585
R3341 gnd.n5446 gnd.n5445 585
R3342 gnd.n5443 gnd.n5442 585
R3343 gnd.n5441 gnd.n5440 585
R3344 gnd.n5439 gnd.n5438 585
R3345 gnd.n5437 gnd.n5436 585
R3346 gnd.n5435 gnd.n5434 585
R3347 gnd.n5433 gnd.n5432 585
R3348 gnd.n5431 gnd.n5430 585
R3349 gnd.n5429 gnd.n5428 585
R3350 gnd.n5427 gnd.n5426 585
R3351 gnd.n5425 gnd.n5424 585
R3352 gnd.n5423 gnd.n5422 585
R3353 gnd.n5421 gnd.n5420 585
R3354 gnd.n5419 gnd.n5418 585
R3355 gnd.n5417 gnd.n5416 585
R3356 gnd.n5415 gnd.n5414 585
R3357 gnd.n5413 gnd.n5412 585
R3358 gnd.n5411 gnd.n5410 585
R3359 gnd.n5409 gnd.n5408 585
R3360 gnd.n5407 gnd.n5406 585
R3361 gnd.n5405 gnd.n5404 585
R3362 gnd.n5403 gnd.n5402 585
R3363 gnd.n5401 gnd.n5400 585
R3364 gnd.n5399 gnd.n5398 585
R3365 gnd.n5397 gnd.n5396 585
R3366 gnd.n5395 gnd.n5394 585
R3367 gnd.n5393 gnd.n5392 585
R3368 gnd.n5391 gnd.n5390 585
R3369 gnd.n5389 gnd.n5388 585
R3370 gnd.n5387 gnd.n5386 585
R3371 gnd.n5385 gnd.n5384 585
R3372 gnd.n5379 gnd.n5378 585
R3373 gnd.n6964 gnd.n6963 585
R3374 gnd.n6970 gnd.n6969 585
R3375 gnd.n6972 gnd.n6971 585
R3376 gnd.n6974 gnd.n6973 585
R3377 gnd.n6976 gnd.n6975 585
R3378 gnd.n6978 gnd.n6977 585
R3379 gnd.n6980 gnd.n6979 585
R3380 gnd.n6982 gnd.n6981 585
R3381 gnd.n6984 gnd.n6983 585
R3382 gnd.n6986 gnd.n6985 585
R3383 gnd.n6988 gnd.n6987 585
R3384 gnd.n6990 gnd.n6989 585
R3385 gnd.n6992 gnd.n6991 585
R3386 gnd.n6994 gnd.n6993 585
R3387 gnd.n6996 gnd.n6995 585
R3388 gnd.n6998 gnd.n6997 585
R3389 gnd.n7000 gnd.n6999 585
R3390 gnd.n7002 gnd.n7001 585
R3391 gnd.n7004 gnd.n7003 585
R3392 gnd.n7007 gnd.n7006 585
R3393 gnd.n7005 gnd.n6943 585
R3394 gnd.n7012 gnd.n7011 585
R3395 gnd.n7014 gnd.n7013 585
R3396 gnd.n7016 gnd.n7015 585
R3397 gnd.n7018 gnd.n7017 585
R3398 gnd.n7020 gnd.n7019 585
R3399 gnd.n7022 gnd.n7021 585
R3400 gnd.n7024 gnd.n7023 585
R3401 gnd.n7026 gnd.n7025 585
R3402 gnd.n7028 gnd.n7027 585
R3403 gnd.n7030 gnd.n7029 585
R3404 gnd.n7032 gnd.n7031 585
R3405 gnd.n7034 gnd.n7033 585
R3406 gnd.n7036 gnd.n7035 585
R3407 gnd.n7038 gnd.n7037 585
R3408 gnd.n7040 gnd.n7039 585
R3409 gnd.n7042 gnd.n7041 585
R3410 gnd.n7044 gnd.n7043 585
R3411 gnd.n7046 gnd.n7045 585
R3412 gnd.n7048 gnd.n7047 585
R3413 gnd.n7050 gnd.n7049 585
R3414 gnd.n7055 gnd.n7054 585
R3415 gnd.n7057 gnd.n7056 585
R3416 gnd.n7059 gnd.n7058 585
R3417 gnd.n7061 gnd.n7060 585
R3418 gnd.n7063 gnd.n7062 585
R3419 gnd.n7065 gnd.n7064 585
R3420 gnd.n7067 gnd.n7066 585
R3421 gnd.n7069 gnd.n7068 585
R3422 gnd.n7071 gnd.n7070 585
R3423 gnd.n7073 gnd.n7072 585
R3424 gnd.n7075 gnd.n7074 585
R3425 gnd.n7077 gnd.n7076 585
R3426 gnd.n7079 gnd.n7078 585
R3427 gnd.n7081 gnd.n7080 585
R3428 gnd.n7082 gnd.n6903 585
R3429 gnd.n7084 gnd.n7083 585
R3430 gnd.n6904 gnd.n6902 585
R3431 gnd.n6905 gnd.n166 585
R3432 gnd.n7086 gnd.n166 585
R3433 gnd.n7143 gnd.n168 585
R3434 gnd.n7147 gnd.n168 585
R3435 gnd.n7142 gnd.n7141 585
R3436 gnd.n7141 gnd.n167 585
R3437 gnd.n7140 gnd.n159 585
R3438 gnd.n7153 gnd.n159 585
R3439 gnd.n7139 gnd.n7138 585
R3440 gnd.n7138 gnd.n152 585
R3441 gnd.n7137 gnd.n150 585
R3442 gnd.n7159 gnd.n150 585
R3443 gnd.n7136 gnd.n7135 585
R3444 gnd.n7135 gnd.n142 585
R3445 gnd.n7133 gnd.n140 585
R3446 gnd.n7165 gnd.n140 585
R3447 gnd.n7132 gnd.n7131 585
R3448 gnd.n7131 gnd.n133 585
R3449 gnd.n7130 gnd.n131 585
R3450 gnd.n7171 gnd.n131 585
R3451 gnd.n7129 gnd.n7128 585
R3452 gnd.n7128 gnd.n130 585
R3453 gnd.n7126 gnd.n121 585
R3454 gnd.n7177 gnd.n121 585
R3455 gnd.n7125 gnd.n7124 585
R3456 gnd.n7124 gnd.n120 585
R3457 gnd.n7123 gnd.n112 585
R3458 gnd.n7183 gnd.n112 585
R3459 gnd.n7122 gnd.n7121 585
R3460 gnd.n7121 gnd.n111 585
R3461 gnd.n7119 gnd.n102 585
R3462 gnd.n7189 gnd.n102 585
R3463 gnd.n7118 gnd.n7117 585
R3464 gnd.n7117 gnd.n7116 585
R3465 gnd.n174 gnd.n91 585
R3466 gnd.n7195 gnd.n91 585
R3467 gnd.n6790 gnd.n6789 585
R3468 gnd.n6791 gnd.n6790 585
R3469 gnd.n178 gnd.n177 585
R3470 gnd.n6784 gnd.n177 585
R3471 gnd.n5301 gnd.n74 585
R3472 gnd.n7203 gnd.n74 585
R3473 gnd.n5302 gnd.n1597 585
R3474 gnd.n5306 gnd.n1597 585
R3475 gnd.n5300 gnd.n5299 585
R3476 gnd.n5299 gnd.n1596 585
R3477 gnd.n5298 gnd.n1601 585
R3478 gnd.n5298 gnd.n5297 585
R3479 gnd.n5292 gnd.n1585 585
R3480 gnd.n5315 gnd.n1585 585
R3481 gnd.n5291 gnd.n1579 585
R3482 gnd.n5320 gnd.n1579 585
R3483 gnd.n5290 gnd.n5289 585
R3484 gnd.n5289 gnd.n5288 585
R3485 gnd.n1605 gnd.n1569 585
R3486 gnd.n5326 gnd.n1569 585
R3487 gnd.n5275 gnd.n5274 585
R3488 gnd.n5276 gnd.n5275 585
R3489 gnd.n5272 gnd.n1562 585
R3490 gnd.n5332 gnd.n1562 585
R3491 gnd.n5271 gnd.n5270 585
R3492 gnd.n5270 gnd.n5269 585
R3493 gnd.n1611 gnd.n1552 585
R3494 gnd.n5338 gnd.n1552 585
R3495 gnd.n5197 gnd.n1615 585
R3496 gnd.n5261 gnd.n1615 585
R3497 gnd.n5198 gnd.n1542 585
R3498 gnd.n5344 gnd.n1542 585
R3499 gnd.n5200 gnd.n5199 585
R3500 gnd.n5201 gnd.n5200 585
R3501 gnd.n5195 gnd.n1532 585
R3502 gnd.n5350 gnd.n1532 585
R3503 gnd.n5194 gnd.n5193 585
R3504 gnd.n5193 gnd.n5192 585
R3505 gnd.n5189 gnd.n1522 585
R3506 gnd.n5356 gnd.n1522 585
R3507 gnd.n5188 gnd.n5187 585
R3508 gnd.n5187 gnd.n5186 585
R3509 gnd.n5185 gnd.n1509 585
R3510 gnd.n5362 gnd.n1509 585
R3511 gnd.n1493 gnd.n1492 585
R3512 gnd.n5179 gnd.n1493 585
R3513 gnd.n5370 gnd.n5369 585
R3514 gnd.n5369 gnd.n5368 585
R3515 gnd.n5371 gnd.n1482 585
R3516 gnd.n5218 gnd.n1482 585
R3517 gnd.n5377 gnd.n1483 585
R3518 gnd.n5377 gnd.n5376 585
R3519 gnd.n5972 gnd.n727 585
R3520 gnd.n2134 gnd.n727 585
R3521 gnd.n6776 gnd.n6775 585
R3522 gnd.n6776 gnd.n104 585
R3523 gnd.n6778 gnd.n6777 585
R3524 gnd.n6777 gnd.n93 585
R3525 gnd.n6779 gnd.n182 585
R3526 gnd.n182 gnd.n90 585
R3527 gnd.n6782 gnd.n6781 585
R3528 gnd.n6783 gnd.n6782 585
R3529 gnd.n183 gnd.n181 585
R3530 gnd.n181 gnd.n75 585
R3531 gnd.n1592 gnd.n1591 585
R3532 gnd.n1592 gnd.n73 585
R3533 gnd.n5309 gnd.n5308 585
R3534 gnd.n5308 gnd.n5307 585
R3535 gnd.n5311 gnd.n1588 585
R3536 gnd.n1604 gnd.n1588 585
R3537 gnd.n5313 gnd.n5312 585
R3538 gnd.n5314 gnd.n5313 585
R3539 gnd.n5247 gnd.n1587 585
R3540 gnd.n1587 gnd.n1581 585
R3541 gnd.n5249 gnd.n5248 585
R3542 gnd.n5248 gnd.n1578 585
R3543 gnd.n5251 gnd.n5244 585
R3544 gnd.n5244 gnd.n1571 585
R3545 gnd.n5253 gnd.n5252 585
R3546 gnd.n5253 gnd.n1568 585
R3547 gnd.n5254 gnd.n5243 585
R3548 gnd.n5254 gnd.n1610 585
R3549 gnd.n5256 gnd.n5255 585
R3550 gnd.n5255 gnd.n1561 585
R3551 gnd.n5257 gnd.n1617 585
R3552 gnd.n1617 gnd.n1554 585
R3553 gnd.n5259 gnd.n5258 585
R3554 gnd.n5260 gnd.n5259 585
R3555 gnd.n1618 gnd.n1616 585
R3556 gnd.n1616 gnd.n1544 585
R3557 gnd.n5237 gnd.n5236 585
R3558 gnd.n5236 gnd.n1541 585
R3559 gnd.n5235 gnd.n1620 585
R3560 gnd.n5235 gnd.n1534 585
R3561 gnd.n5234 gnd.n5233 585
R3562 gnd.n5234 gnd.n1531 585
R3563 gnd.n1622 gnd.n1621 585
R3564 gnd.n5191 gnd.n1621 585
R3565 gnd.n5229 gnd.n5228 585
R3566 gnd.n5228 gnd.n1521 585
R3567 gnd.n5227 gnd.n1624 585
R3568 gnd.n5227 gnd.n1511 585
R3569 gnd.n5226 gnd.n5225 585
R3570 gnd.n5226 gnd.n1508 585
R3571 gnd.n1626 gnd.n1625 585
R3572 gnd.n1625 gnd.n1495 585
R3573 gnd.n5221 gnd.n5220 585
R3574 gnd.n5220 gnd.n5219 585
R3575 gnd.n1629 gnd.n1628 585
R3576 gnd.n1629 gnd.n1486 585
R3577 gnd.n5162 gnd.n5161 585
R3578 gnd.n5162 gnd.n1484 585
R3579 gnd.n5163 gnd.n5158 585
R3580 gnd.n5163 gnd.n1416 585
R3581 gnd.n5165 gnd.n5164 585
R3582 gnd.n5164 gnd.n1374 585
R3583 gnd.n5166 gnd.n1661 585
R3584 gnd.n1661 gnd.n1659 585
R3585 gnd.n5168 gnd.n5167 585
R3586 gnd.n5169 gnd.n5168 585
R3587 gnd.n1662 gnd.n1660 585
R3588 gnd.n1660 gnd.n1307 585
R3589 gnd.n5152 gnd.n1306 585
R3590 gnd.n5565 gnd.n1306 585
R3591 gnd.n5151 gnd.n5150 585
R3592 gnd.n5150 gnd.n1305 585
R3593 gnd.n5149 gnd.n1664 585
R3594 gnd.n5149 gnd.n5148 585
R3595 gnd.n5137 gnd.n1665 585
R3596 gnd.n1667 gnd.n1665 585
R3597 gnd.n5139 gnd.n5138 585
R3598 gnd.n5140 gnd.n5139 585
R3599 gnd.n1675 gnd.n1674 585
R3600 gnd.n1674 gnd.n1673 585
R3601 gnd.n5131 gnd.n5130 585
R3602 gnd.n5130 gnd.n5129 585
R3603 gnd.n1678 gnd.n1677 585
R3604 gnd.n1686 gnd.n1678 585
R3605 gnd.n5120 gnd.n5119 585
R3606 gnd.n5121 gnd.n5120 585
R3607 gnd.n1688 gnd.n1687 585
R3608 gnd.n1687 gnd.n1684 585
R3609 gnd.n5115 gnd.n5114 585
R3610 gnd.n5114 gnd.n5113 585
R3611 gnd.n1691 gnd.n1690 585
R3612 gnd.n1693 gnd.n1691 585
R3613 gnd.n5104 gnd.n5103 585
R3614 gnd.n5105 gnd.n5104 585
R3615 gnd.n1701 gnd.n1700 585
R3616 gnd.n1700 gnd.n1699 585
R3617 gnd.n5099 gnd.n5098 585
R3618 gnd.n5098 gnd.n5097 585
R3619 gnd.n1704 gnd.n1703 585
R3620 gnd.n1706 gnd.n1704 585
R3621 gnd.n5088 gnd.n5087 585
R3622 gnd.n5089 gnd.n5088 585
R3623 gnd.n1714 gnd.n1713 585
R3624 gnd.n1713 gnd.n1712 585
R3625 gnd.n5083 gnd.n5082 585
R3626 gnd.n5082 gnd.n5081 585
R3627 gnd.n1717 gnd.n1716 585
R3628 gnd.n1719 gnd.n1717 585
R3629 gnd.n5072 gnd.n5071 585
R3630 gnd.n5073 gnd.n5072 585
R3631 gnd.n1726 gnd.n1725 585
R3632 gnd.n5064 gnd.n1725 585
R3633 gnd.n5067 gnd.n5066 585
R3634 gnd.n5066 gnd.n5065 585
R3635 gnd.n1729 gnd.n1728 585
R3636 gnd.n1731 gnd.n1729 585
R3637 gnd.n5055 gnd.n5054 585
R3638 gnd.n5056 gnd.n5055 585
R3639 gnd.n1739 gnd.n1738 585
R3640 gnd.n1738 gnd.n1737 585
R3641 gnd.n5050 gnd.n5049 585
R3642 gnd.n5049 gnd.n5048 585
R3643 gnd.n1742 gnd.n1741 585
R3644 gnd.n1744 gnd.n1742 585
R3645 gnd.n5039 gnd.n5038 585
R3646 gnd.n5040 gnd.n5039 585
R3647 gnd.n1751 gnd.n1750 585
R3648 gnd.n5031 gnd.n1750 585
R3649 gnd.n5034 gnd.n5033 585
R3650 gnd.n5033 gnd.n5032 585
R3651 gnd.n1754 gnd.n1753 585
R3652 gnd.n1797 gnd.n1754 585
R3653 gnd.n4864 gnd.n4863 585
R3654 gnd.n4865 gnd.n4864 585
R3655 gnd.n1807 gnd.n1806 585
R3656 gnd.n4790 gnd.n1806 585
R3657 gnd.n4859 gnd.n4858 585
R3658 gnd.n4858 gnd.n4857 585
R3659 gnd.n1810 gnd.n1809 585
R3660 gnd.n1818 gnd.n1810 585
R3661 gnd.n4828 gnd.n1833 585
R3662 gnd.n1833 gnd.n1825 585
R3663 gnd.n4830 gnd.n4829 585
R3664 gnd.n4831 gnd.n4830 585
R3665 gnd.n1834 gnd.n1832 585
R3666 gnd.n1832 gnd.n1829 585
R3667 gnd.n4823 gnd.n4822 585
R3668 gnd.n4822 gnd.n4821 585
R3669 gnd.n1837 gnd.n1836 585
R3670 gnd.n4812 gnd.n1837 585
R3671 gnd.n4776 gnd.n1854 585
R3672 gnd.n4760 gnd.n1854 585
R3673 gnd.n4778 gnd.n4777 585
R3674 gnd.n4779 gnd.n4778 585
R3675 gnd.n1855 gnd.n1853 585
R3676 gnd.n4744 gnd.n1853 585
R3677 gnd.n4771 gnd.n4770 585
R3678 gnd.n4770 gnd.n4769 585
R3679 gnd.n1858 gnd.n1857 585
R3680 gnd.n1870 gnd.n1858 585
R3681 gnd.n4730 gnd.n4729 585
R3682 gnd.n4731 gnd.n4730 585
R3683 gnd.n1878 gnd.n1877 585
R3684 gnd.n4628 gnd.n1877 585
R3685 gnd.n4725 gnd.n4724 585
R3686 gnd.n4724 gnd.n4723 585
R3687 gnd.n1881 gnd.n1880 585
R3688 gnd.n4715 gnd.n1881 585
R3689 gnd.n4674 gnd.n4673 585
R3690 gnd.n4674 gnd.n1895 585
R3691 gnd.n4675 gnd.n4670 585
R3692 gnd.n4675 gnd.n1894 585
R3693 gnd.n4677 gnd.n4676 585
R3694 gnd.n4676 gnd.n1899 585
R3695 gnd.n4678 gnd.n1914 585
R3696 gnd.n1914 gnd.n1905 585
R3697 gnd.n4680 gnd.n4679 585
R3698 gnd.n4681 gnd.n4680 585
R3699 gnd.n1915 gnd.n1913 585
R3700 gnd.n1913 gnd.n1910 585
R3701 gnd.n4664 gnd.n4663 585
R3702 gnd.n4663 gnd.n4662 585
R3703 gnd.n1918 gnd.n1917 585
R3704 gnd.n4654 gnd.n1918 585
R3705 gnd.n4609 gnd.n1935 585
R3706 gnd.n4588 gnd.n1935 585
R3707 gnd.n4611 gnd.n4610 585
R3708 gnd.n4612 gnd.n4611 585
R3709 gnd.n1936 gnd.n1934 585
R3710 gnd.n1949 gnd.n1934 585
R3711 gnd.n4604 gnd.n4603 585
R3712 gnd.n4603 gnd.n4602 585
R3713 gnd.n1939 gnd.n1938 585
R3714 gnd.n4538 gnd.n1939 585
R3715 gnd.n4566 gnd.n4565 585
R3716 gnd.n4567 gnd.n4566 585
R3717 gnd.n1963 gnd.n1962 585
R3718 gnd.n1962 gnd.n1957 585
R3719 gnd.n4561 gnd.n4560 585
R3720 gnd.n4560 gnd.n4559 585
R3721 gnd.n1967 gnd.n1966 585
R3722 gnd.n4551 gnd.n1967 585
R3723 gnd.n1212 gnd.n1211 585
R3724 gnd.n4522 gnd.n1212 585
R3725 gnd.n5673 gnd.n5672 585
R3726 gnd.n5672 gnd.n5671 585
R3727 gnd.n5674 gnd.n1206 585
R3728 gnd.n4530 gnd.n1206 585
R3729 gnd.n5676 gnd.n5675 585
R3730 gnd.n5677 gnd.n5676 585
R3731 gnd.n1207 gnd.n1205 585
R3732 gnd.n4425 gnd.n1205 585
R3733 gnd.n4411 gnd.n4410 585
R3734 gnd.n4410 gnd.n1175 585
R3735 gnd.n4412 gnd.n1992 585
R3736 gnd.n1992 gnd.n1143 585
R3737 gnd.n4414 gnd.n4413 585
R3738 gnd.n4415 gnd.n4414 585
R3739 gnd.n1993 gnd.n1991 585
R3740 gnd.n1991 gnd.n1989 585
R3741 gnd.n4403 gnd.n4402 585
R3742 gnd.n4402 gnd.n4401 585
R3743 gnd.n1996 gnd.n1995 585
R3744 gnd.n1997 gnd.n1996 585
R3745 gnd.n4391 gnd.n4390 585
R3746 gnd.n4392 gnd.n4391 585
R3747 gnd.n2008 gnd.n2007 585
R3748 gnd.n2007 gnd.n2005 585
R3749 gnd.n4386 gnd.n4385 585
R3750 gnd.n4385 gnd.n4384 585
R3751 gnd.n2011 gnd.n2010 585
R3752 gnd.n2020 gnd.n2011 585
R3753 gnd.n4375 gnd.n4374 585
R3754 gnd.n4376 gnd.n4375 585
R3755 gnd.n2022 gnd.n2021 585
R3756 gnd.n2021 gnd.n2018 585
R3757 gnd.n4370 gnd.n4369 585
R3758 gnd.n4369 gnd.n4368 585
R3759 gnd.n2025 gnd.n2024 585
R3760 gnd.n2026 gnd.n2025 585
R3761 gnd.n4359 gnd.n4358 585
R3762 gnd.n4360 gnd.n4359 585
R3763 gnd.n2036 gnd.n2035 585
R3764 gnd.n2035 gnd.n2033 585
R3765 gnd.n4354 gnd.n4353 585
R3766 gnd.n4353 gnd.n4352 585
R3767 gnd.n2039 gnd.n2038 585
R3768 gnd.n2040 gnd.n2039 585
R3769 gnd.n4343 gnd.n4342 585
R3770 gnd.n4344 gnd.n4343 585
R3771 gnd.n2050 gnd.n2049 585
R3772 gnd.n2049 gnd.n2047 585
R3773 gnd.n4338 gnd.n4337 585
R3774 gnd.n4337 gnd.n4336 585
R3775 gnd.n2053 gnd.n2052 585
R3776 gnd.n2054 gnd.n2053 585
R3777 gnd.n4327 gnd.n4326 585
R3778 gnd.n4328 gnd.n4327 585
R3779 gnd.n2063 gnd.n2062 585
R3780 gnd.n2069 gnd.n2062 585
R3781 gnd.n4322 gnd.n4321 585
R3782 gnd.n4321 gnd.n4320 585
R3783 gnd.n2066 gnd.n2065 585
R3784 gnd.n2067 gnd.n2066 585
R3785 gnd.n4311 gnd.n4310 585
R3786 gnd.n4312 gnd.n4311 585
R3787 gnd.n2078 gnd.n2077 585
R3788 gnd.n2077 gnd.n2075 585
R3789 gnd.n4306 gnd.n4305 585
R3790 gnd.n4305 gnd.n4304 585
R3791 gnd.n4227 gnd.n2080 585
R3792 gnd.n4228 gnd.n4227 585
R3793 gnd.n4226 gnd.n4225 585
R3794 gnd.n4226 gnd.n890 585
R3795 gnd.n2082 gnd.n2081 585
R3796 gnd.n2081 gnd.n876 585
R3797 gnd.n4221 gnd.n4220 585
R3798 gnd.n4220 gnd.n4219 585
R3799 gnd.n4218 gnd.n2084 585
R3800 gnd.n4218 gnd.n979 585
R3801 gnd.n4217 gnd.n4216 585
R3802 gnd.n4217 gnd.n965 585
R3803 gnd.n2086 gnd.n2085 585
R3804 gnd.n2085 gnd.n862 585
R3805 gnd.n4212 gnd.n4211 585
R3806 gnd.n4211 gnd.n859 585
R3807 gnd.n4210 gnd.n2088 585
R3808 gnd.n4210 gnd.n867 585
R3809 gnd.n4209 gnd.n4208 585
R3810 gnd.n4209 gnd.n850 585
R3811 gnd.n2090 gnd.n2089 585
R3812 gnd.n2089 gnd.n843 585
R3813 gnd.n4204 gnd.n4203 585
R3814 gnd.n4203 gnd.n840 585
R3815 gnd.n4202 gnd.n2092 585
R3816 gnd.n4202 gnd.n832 585
R3817 gnd.n4201 gnd.n2094 585
R3818 gnd.n4201 gnd.n4200 585
R3819 gnd.n4140 gnd.n2093 585
R3820 gnd.n2093 gnd.n823 585
R3821 gnd.n4142 gnd.n4141 585
R3822 gnd.n4141 gnd.n820 585
R3823 gnd.n4143 gnd.n4133 585
R3824 gnd.n4133 gnd.n812 585
R3825 gnd.n4145 gnd.n4144 585
R3826 gnd.n4145 gnd.n809 585
R3827 gnd.n4146 gnd.n4132 585
R3828 gnd.n4146 gnd.n2106 585
R3829 gnd.n4148 gnd.n4147 585
R3830 gnd.n4147 gnd.n800 585
R3831 gnd.n4149 gnd.n2114 585
R3832 gnd.n2114 gnd.n792 585
R3833 gnd.n4151 gnd.n4150 585
R3834 gnd.n4152 gnd.n4151 585
R3835 gnd.n4127 gnd.n2113 585
R3836 gnd.n2113 gnd.n783 585
R3837 gnd.n4126 gnd.n4125 585
R3838 gnd.n4125 gnd.n780 585
R3839 gnd.n4124 gnd.n4123 585
R3840 gnd.n4124 gnd.n775 585
R3841 gnd.n4122 gnd.n2116 585
R3842 gnd.n2116 gnd.n772 585
R3843 gnd.n4120 gnd.n4119 585
R3844 gnd.n4119 gnd.n4118 585
R3845 gnd.n2118 gnd.n2117 585
R3846 gnd.n2118 gnd.n763 585
R3847 gnd.n4086 gnd.n4079 585
R3848 gnd.n4079 gnd.n758 585
R3849 gnd.n4088 gnd.n4087 585
R3850 gnd.n4089 gnd.n4088 585
R3851 gnd.n4083 gnd.n4078 585
R3852 gnd.n4078 gnd.n747 585
R3853 gnd.n4082 gnd.n4081 585
R3854 gnd.n4081 gnd.n744 585
R3855 gnd.n732 gnd.n731 585
R3856 gnd.n736 gnd.n732 585
R3857 gnd.n5969 gnd.n5968 585
R3858 gnd.n5968 gnd.n5967 585
R3859 gnd.n5564 gnd.n5563 585
R3860 gnd.n5565 gnd.n5564 585
R3861 gnd.n1310 gnd.n1308 585
R3862 gnd.n1308 gnd.n1305 585
R3863 gnd.n5147 gnd.n5146 585
R3864 gnd.n5148 gnd.n5147 585
R3865 gnd.n1669 gnd.n1668 585
R3866 gnd.n1668 gnd.n1667 585
R3867 gnd.n5142 gnd.n5141 585
R3868 gnd.n5141 gnd.n5140 585
R3869 gnd.n1672 gnd.n1671 585
R3870 gnd.n1673 gnd.n1672 585
R3871 gnd.n5128 gnd.n5127 585
R3872 gnd.n5129 gnd.n5128 585
R3873 gnd.n1680 gnd.n1679 585
R3874 gnd.n1686 gnd.n1679 585
R3875 gnd.n5123 gnd.n5122 585
R3876 gnd.n5122 gnd.n5121 585
R3877 gnd.n1683 gnd.n1682 585
R3878 gnd.n1684 gnd.n1683 585
R3879 gnd.n5112 gnd.n5111 585
R3880 gnd.n5113 gnd.n5112 585
R3881 gnd.n1695 gnd.n1694 585
R3882 gnd.n1694 gnd.n1693 585
R3883 gnd.n5107 gnd.n5106 585
R3884 gnd.n5106 gnd.n5105 585
R3885 gnd.n1698 gnd.n1697 585
R3886 gnd.n1699 gnd.n1698 585
R3887 gnd.n5096 gnd.n5095 585
R3888 gnd.n5097 gnd.n5096 585
R3889 gnd.n1708 gnd.n1707 585
R3890 gnd.n1707 gnd.n1706 585
R3891 gnd.n5091 gnd.n5090 585
R3892 gnd.n5090 gnd.n5089 585
R3893 gnd.n1711 gnd.n1710 585
R3894 gnd.n1712 gnd.n1711 585
R3895 gnd.n5080 gnd.n5079 585
R3896 gnd.n5081 gnd.n5080 585
R3897 gnd.n1721 gnd.n1720 585
R3898 gnd.n1720 gnd.n1719 585
R3899 gnd.n5075 gnd.n5074 585
R3900 gnd.n5074 gnd.n5073 585
R3901 gnd.n1724 gnd.n1723 585
R3902 gnd.n5064 gnd.n1724 585
R3903 gnd.n5063 gnd.n5062 585
R3904 gnd.n5065 gnd.n5063 585
R3905 gnd.n1733 gnd.n1732 585
R3906 gnd.n1732 gnd.n1731 585
R3907 gnd.n5058 gnd.n5057 585
R3908 gnd.n5057 gnd.n5056 585
R3909 gnd.n1736 gnd.n1735 585
R3910 gnd.n1737 gnd.n1736 585
R3911 gnd.n5047 gnd.n5046 585
R3912 gnd.n5048 gnd.n5047 585
R3913 gnd.n1746 gnd.n1745 585
R3914 gnd.n1745 gnd.n1744 585
R3915 gnd.n5042 gnd.n5041 585
R3916 gnd.n5041 gnd.n5040 585
R3917 gnd.n1749 gnd.n1748 585
R3918 gnd.n5031 gnd.n1749 585
R3919 gnd.n4794 gnd.n1756 585
R3920 gnd.n5032 gnd.n1756 585
R3921 gnd.n4793 gnd.n4792 585
R3922 gnd.n4792 gnd.n1797 585
R3923 gnd.n4798 gnd.n1804 585
R3924 gnd.n4865 gnd.n1804 585
R3925 gnd.n4799 gnd.n4791 585
R3926 gnd.n4791 gnd.n4790 585
R3927 gnd.n4800 gnd.n1812 585
R3928 gnd.n4857 gnd.n1812 585
R3929 gnd.n4788 gnd.n4787 585
R3930 gnd.n4787 gnd.n1818 585
R3931 gnd.n4804 gnd.n4786 585
R3932 gnd.n4786 gnd.n1825 585
R3933 gnd.n4805 gnd.n1831 585
R3934 gnd.n4831 gnd.n1831 585
R3935 gnd.n4806 gnd.n4785 585
R3936 gnd.n4785 gnd.n1829 585
R3937 gnd.n1848 gnd.n1839 585
R3938 gnd.n4821 gnd.n1839 585
R3939 gnd.n4811 gnd.n4810 585
R3940 gnd.n4812 gnd.n4811 585
R3941 gnd.n1847 gnd.n1846 585
R3942 gnd.n4760 gnd.n1846 585
R3943 gnd.n4781 gnd.n4780 585
R3944 gnd.n4780 gnd.n4779 585
R3945 gnd.n1851 gnd.n1850 585
R3946 gnd.n4744 gnd.n1851 585
R3947 gnd.n4631 gnd.n1860 585
R3948 gnd.n4769 gnd.n1860 585
R3949 gnd.n4634 gnd.n4630 585
R3950 gnd.n4630 gnd.n1870 585
R3951 gnd.n4635 gnd.n1875 585
R3952 gnd.n4731 gnd.n1875 585
R3953 gnd.n4636 gnd.n4629 585
R3954 gnd.n4629 gnd.n4628 585
R3955 gnd.n4625 gnd.n1882 585
R3956 gnd.n4723 gnd.n1882 585
R3957 gnd.n4640 gnd.n1890 585
R3958 gnd.n4715 gnd.n1890 585
R3959 gnd.n4641 gnd.n4624 585
R3960 gnd.n4624 gnd.n1895 585
R3961 gnd.n4642 gnd.n4623 585
R3962 gnd.n4623 gnd.n1894 585
R3963 gnd.n4622 gnd.n4620 585
R3964 gnd.n4622 gnd.n1899 585
R3965 gnd.n4646 gnd.n4619 585
R3966 gnd.n4619 gnd.n1905 585
R3967 gnd.n4647 gnd.n1912 585
R3968 gnd.n4681 gnd.n1912 585
R3969 gnd.n4648 gnd.n4618 585
R3970 gnd.n4618 gnd.n1910 585
R3971 gnd.n1928 gnd.n1920 585
R3972 gnd.n4662 gnd.n1920 585
R3973 gnd.n4653 gnd.n4652 585
R3974 gnd.n4654 gnd.n4653 585
R3975 gnd.n1927 gnd.n1926 585
R3976 gnd.n4588 gnd.n1926 585
R3977 gnd.n4614 gnd.n4613 585
R3978 gnd.n4613 gnd.n4612 585
R3979 gnd.n1931 gnd.n1930 585
R3980 gnd.n1949 gnd.n1931 585
R3981 gnd.n4540 gnd.n1941 585
R3982 gnd.n4602 gnd.n1941 585
R3983 gnd.n4543 gnd.n4539 585
R3984 gnd.n4539 gnd.n4538 585
R3985 gnd.n4544 gnd.n1959 585
R3986 gnd.n4567 gnd.n1959 585
R3987 gnd.n4545 gnd.n4537 585
R3988 gnd.n4537 gnd.n1957 585
R3989 gnd.n1977 gnd.n1969 585
R3990 gnd.n4559 gnd.n1969 585
R3991 gnd.n4550 gnd.n4549 585
R3992 gnd.n4551 gnd.n4550 585
R3993 gnd.n1976 gnd.n1975 585
R3994 gnd.n4522 gnd.n1975 585
R3995 gnd.n4533 gnd.n1214 585
R3996 gnd.n5671 gnd.n1214 585
R3997 gnd.n4532 gnd.n4531 585
R3998 gnd.n4531 gnd.n4530 585
R3999 gnd.n4432 gnd.n1203 585
R4000 gnd.n5677 gnd.n1203 585
R4001 gnd.n4426 gnd.n1979 585
R4002 gnd.n4426 gnd.n4425 585
R4003 gnd.n4428 gnd.n4427 585
R4004 gnd.n4427 gnd.n1175 585
R4005 gnd.n1982 gnd.n1981 585
R4006 gnd.n1982 gnd.n1143 585
R4007 gnd.n4257 gnd.n1990 585
R4008 gnd.n4415 gnd.n1990 585
R4009 gnd.n4256 gnd.n4255 585
R4010 gnd.n4255 gnd.n1989 585
R4011 gnd.n4261 gnd.n1998 585
R4012 gnd.n4401 gnd.n1998 585
R4013 gnd.n4262 gnd.n4254 585
R4014 gnd.n4254 gnd.n1997 585
R4015 gnd.n4263 gnd.n2006 585
R4016 gnd.n4392 gnd.n2006 585
R4017 gnd.n4252 gnd.n4251 585
R4018 gnd.n4251 gnd.n2005 585
R4019 gnd.n4267 gnd.n2012 585
R4020 gnd.n4384 gnd.n2012 585
R4021 gnd.n4268 gnd.n4250 585
R4022 gnd.n4250 gnd.n2020 585
R4023 gnd.n4269 gnd.n2019 585
R4024 gnd.n4376 gnd.n2019 585
R4025 gnd.n4248 gnd.n4247 585
R4026 gnd.n4247 gnd.n2018 585
R4027 gnd.n4273 gnd.n2027 585
R4028 gnd.n4368 gnd.n2027 585
R4029 gnd.n4274 gnd.n4246 585
R4030 gnd.n4246 gnd.n2026 585
R4031 gnd.n4275 gnd.n2034 585
R4032 gnd.n4360 gnd.n2034 585
R4033 gnd.n4244 gnd.n4243 585
R4034 gnd.n4243 gnd.n2033 585
R4035 gnd.n4279 gnd.n2041 585
R4036 gnd.n4352 gnd.n2041 585
R4037 gnd.n4280 gnd.n4242 585
R4038 gnd.n4242 gnd.n2040 585
R4039 gnd.n4281 gnd.n2048 585
R4040 gnd.n4344 gnd.n2048 585
R4041 gnd.n4240 gnd.n4239 585
R4042 gnd.n4239 gnd.n2047 585
R4043 gnd.n4285 gnd.n2055 585
R4044 gnd.n4336 gnd.n2055 585
R4045 gnd.n4286 gnd.n4238 585
R4046 gnd.n4238 gnd.n2054 585
R4047 gnd.n4287 gnd.n2061 585
R4048 gnd.n4328 gnd.n2061 585
R4049 gnd.n4236 gnd.n4235 585
R4050 gnd.n4235 gnd.n2069 585
R4051 gnd.n4291 gnd.n2068 585
R4052 gnd.n4320 gnd.n2068 585
R4053 gnd.n4292 gnd.n4234 585
R4054 gnd.n4234 gnd.n2067 585
R4055 gnd.n4293 gnd.n2076 585
R4056 gnd.n4312 gnd.n2076 585
R4057 gnd.n4231 gnd.n4229 585
R4058 gnd.n4229 gnd.n2075 585
R4059 gnd.n4298 gnd.n4297 585
R4060 gnd.n4304 gnd.n4298 585
R4061 gnd.n4230 gnd.n893 585
R4062 gnd.n4228 gnd.n893 585
R4063 gnd.n5865 gnd.n5864 585
R4064 gnd.n5863 gnd.n892 585
R4065 gnd.n895 gnd.n891 585
R4066 gnd.n5867 gnd.n891 585
R4067 gnd.n5859 gnd.n897 585
R4068 gnd.n5858 gnd.n898 585
R4069 gnd.n5857 gnd.n899 585
R4070 gnd.n902 gnd.n900 585
R4071 gnd.n5852 gnd.n903 585
R4072 gnd.n5851 gnd.n904 585
R4073 gnd.n5850 gnd.n905 585
R4074 gnd.n914 gnd.n906 585
R4075 gnd.n5843 gnd.n915 585
R4076 gnd.n5842 gnd.n916 585
R4077 gnd.n918 gnd.n917 585
R4078 gnd.n5835 gnd.n924 585
R4079 gnd.n5834 gnd.n925 585
R4080 gnd.n932 gnd.n926 585
R4081 gnd.n5827 gnd.n933 585
R4082 gnd.n5826 gnd.n934 585
R4083 gnd.n936 gnd.n935 585
R4084 gnd.n5819 gnd.n942 585
R4085 gnd.n5818 gnd.n943 585
R4086 gnd.n950 gnd.n944 585
R4087 gnd.n5811 gnd.n951 585
R4088 gnd.n5810 gnd.n952 585
R4089 gnd.n957 gnd.n956 585
R4090 gnd.n888 gnd.n873 585
R4091 gnd.n5871 gnd.n874 585
R4092 gnd.n5870 gnd.n5869 585
R4093 gnd.n5567 gnd.n5566 585
R4094 gnd.n5566 gnd.n5565 585
R4095 gnd.n5568 gnd.n1302 585
R4096 gnd.n1305 gnd.n1302 585
R4097 gnd.n5569 gnd.n1301 585
R4098 gnd.n5148 gnd.n1301 585
R4099 gnd.n1666 gnd.n1299 585
R4100 gnd.n1667 gnd.n1666 585
R4101 gnd.n5573 gnd.n1298 585
R4102 gnd.n5140 gnd.n1298 585
R4103 gnd.n5574 gnd.n1297 585
R4104 gnd.n1673 gnd.n1297 585
R4105 gnd.n5575 gnd.n1296 585
R4106 gnd.n5129 gnd.n1296 585
R4107 gnd.n1685 gnd.n1294 585
R4108 gnd.n1686 gnd.n1685 585
R4109 gnd.n5579 gnd.n1293 585
R4110 gnd.n5121 gnd.n1293 585
R4111 gnd.n5580 gnd.n1292 585
R4112 gnd.n1684 gnd.n1292 585
R4113 gnd.n5581 gnd.n1291 585
R4114 gnd.n5113 gnd.n1291 585
R4115 gnd.n1692 gnd.n1289 585
R4116 gnd.n1693 gnd.n1692 585
R4117 gnd.n5585 gnd.n1288 585
R4118 gnd.n5105 gnd.n1288 585
R4119 gnd.n5586 gnd.n1287 585
R4120 gnd.n1699 gnd.n1287 585
R4121 gnd.n5587 gnd.n1286 585
R4122 gnd.n5097 gnd.n1286 585
R4123 gnd.n1705 gnd.n1284 585
R4124 gnd.n1706 gnd.n1705 585
R4125 gnd.n5591 gnd.n1283 585
R4126 gnd.n5089 gnd.n1283 585
R4127 gnd.n5592 gnd.n1282 585
R4128 gnd.n1712 gnd.n1282 585
R4129 gnd.n5593 gnd.n1281 585
R4130 gnd.n5081 gnd.n1281 585
R4131 gnd.n1718 gnd.n1279 585
R4132 gnd.n1719 gnd.n1718 585
R4133 gnd.n5597 gnd.n1278 585
R4134 gnd.n5073 gnd.n1278 585
R4135 gnd.n5598 gnd.n1277 585
R4136 gnd.n5064 gnd.n1277 585
R4137 gnd.n5599 gnd.n1276 585
R4138 gnd.n5065 gnd.n1276 585
R4139 gnd.n1730 gnd.n1274 585
R4140 gnd.n1731 gnd.n1730 585
R4141 gnd.n5603 gnd.n1273 585
R4142 gnd.n5056 gnd.n1273 585
R4143 gnd.n5604 gnd.n1272 585
R4144 gnd.n1737 gnd.n1272 585
R4145 gnd.n5605 gnd.n1271 585
R4146 gnd.n5048 gnd.n1271 585
R4147 gnd.n1743 gnd.n1269 585
R4148 gnd.n1744 gnd.n1743 585
R4149 gnd.n5609 gnd.n1268 585
R4150 gnd.n5040 gnd.n1268 585
R4151 gnd.n5610 gnd.n1267 585
R4152 gnd.n5031 gnd.n1267 585
R4153 gnd.n5611 gnd.n1266 585
R4154 gnd.n5032 gnd.n1266 585
R4155 gnd.n1796 gnd.n1264 585
R4156 gnd.n1797 gnd.n1796 585
R4157 gnd.n5615 gnd.n1263 585
R4158 gnd.n4865 gnd.n1263 585
R4159 gnd.n5616 gnd.n1262 585
R4160 gnd.n4790 gnd.n1262 585
R4161 gnd.n5617 gnd.n1261 585
R4162 gnd.n4857 gnd.n1261 585
R4163 gnd.n1817 gnd.n1259 585
R4164 gnd.n1818 gnd.n1817 585
R4165 gnd.n5621 gnd.n1258 585
R4166 gnd.n1825 gnd.n1258 585
R4167 gnd.n5622 gnd.n1257 585
R4168 gnd.n4831 gnd.n1257 585
R4169 gnd.n5623 gnd.n1256 585
R4170 gnd.n1829 gnd.n1256 585
R4171 gnd.n4820 gnd.n1254 585
R4172 gnd.n4821 gnd.n4820 585
R4173 gnd.n5627 gnd.n1253 585
R4174 gnd.n4812 gnd.n1253 585
R4175 gnd.n5628 gnd.n1252 585
R4176 gnd.n4760 gnd.n1252 585
R4177 gnd.n5629 gnd.n1251 585
R4178 gnd.n4779 gnd.n1251 585
R4179 gnd.n4743 gnd.n1249 585
R4180 gnd.n4744 gnd.n4743 585
R4181 gnd.n5633 gnd.n1248 585
R4182 gnd.n4769 gnd.n1248 585
R4183 gnd.n5634 gnd.n1247 585
R4184 gnd.n1870 gnd.n1247 585
R4185 gnd.n5635 gnd.n1246 585
R4186 gnd.n4731 gnd.n1246 585
R4187 gnd.n4627 gnd.n1244 585
R4188 gnd.n4628 gnd.n4627 585
R4189 gnd.n5639 gnd.n1243 585
R4190 gnd.n4723 gnd.n1243 585
R4191 gnd.n5640 gnd.n1242 585
R4192 gnd.n4715 gnd.n1242 585
R4193 gnd.n5641 gnd.n1241 585
R4194 gnd.n1895 gnd.n1241 585
R4195 gnd.n1893 gnd.n1239 585
R4196 gnd.n1894 gnd.n1893 585
R4197 gnd.n5645 gnd.n1238 585
R4198 gnd.n1899 gnd.n1238 585
R4199 gnd.n5646 gnd.n1237 585
R4200 gnd.n1905 gnd.n1237 585
R4201 gnd.n5647 gnd.n1236 585
R4202 gnd.n4681 gnd.n1236 585
R4203 gnd.n1909 gnd.n1234 585
R4204 gnd.n1910 gnd.n1909 585
R4205 gnd.n5651 gnd.n1233 585
R4206 gnd.n4662 gnd.n1233 585
R4207 gnd.n5652 gnd.n1232 585
R4208 gnd.n4654 gnd.n1232 585
R4209 gnd.n5653 gnd.n1231 585
R4210 gnd.n4588 gnd.n1231 585
R4211 gnd.n1933 gnd.n1229 585
R4212 gnd.n4612 gnd.n1933 585
R4213 gnd.n5657 gnd.n1228 585
R4214 gnd.n1949 gnd.n1228 585
R4215 gnd.n5658 gnd.n1227 585
R4216 gnd.n4602 gnd.n1227 585
R4217 gnd.n5659 gnd.n1226 585
R4218 gnd.n4538 gnd.n1226 585
R4219 gnd.n1961 gnd.n1224 585
R4220 gnd.n4567 gnd.n1961 585
R4221 gnd.n5663 gnd.n1223 585
R4222 gnd.n1957 gnd.n1223 585
R4223 gnd.n5664 gnd.n1222 585
R4224 gnd.n4559 gnd.n1222 585
R4225 gnd.n5665 gnd.n1221 585
R4226 gnd.n4551 gnd.n1221 585
R4227 gnd.n1218 gnd.n1216 585
R4228 gnd.n4522 gnd.n1216 585
R4229 gnd.n5670 gnd.n5669 585
R4230 gnd.n5671 gnd.n5670 585
R4231 gnd.n1217 gnd.n1215 585
R4232 gnd.n4530 gnd.n1215 585
R4233 gnd.n1985 gnd.n1204 585
R4234 gnd.n5677 gnd.n1204 585
R4235 gnd.n4424 gnd.n4423 585
R4236 gnd.n4425 gnd.n4424 585
R4237 gnd.n1984 gnd.n1983 585
R4238 gnd.n1983 gnd.n1175 585
R4239 gnd.n4418 gnd.n4417 585
R4240 gnd.n4417 gnd.n1143 585
R4241 gnd.n4416 gnd.n1987 585
R4242 gnd.n4416 gnd.n4415 585
R4243 gnd.n2001 gnd.n1988 585
R4244 gnd.n1989 gnd.n1988 585
R4245 gnd.n4400 gnd.n4399 585
R4246 gnd.n4401 gnd.n4400 585
R4247 gnd.n2000 gnd.n1999 585
R4248 gnd.n1999 gnd.n1997 585
R4249 gnd.n4394 gnd.n4393 585
R4250 gnd.n4393 gnd.n4392 585
R4251 gnd.n2004 gnd.n2003 585
R4252 gnd.n2005 gnd.n2004 585
R4253 gnd.n4383 gnd.n4382 585
R4254 gnd.n4384 gnd.n4383 585
R4255 gnd.n2014 gnd.n2013 585
R4256 gnd.n2020 gnd.n2013 585
R4257 gnd.n4378 gnd.n4377 585
R4258 gnd.n4377 gnd.n4376 585
R4259 gnd.n2017 gnd.n2016 585
R4260 gnd.n2018 gnd.n2017 585
R4261 gnd.n4367 gnd.n4366 585
R4262 gnd.n4368 gnd.n4367 585
R4263 gnd.n2029 gnd.n2028 585
R4264 gnd.n2028 gnd.n2026 585
R4265 gnd.n4362 gnd.n4361 585
R4266 gnd.n4361 gnd.n4360 585
R4267 gnd.n2032 gnd.n2031 585
R4268 gnd.n2033 gnd.n2032 585
R4269 gnd.n4351 gnd.n4350 585
R4270 gnd.n4352 gnd.n4351 585
R4271 gnd.n2043 gnd.n2042 585
R4272 gnd.n2042 gnd.n2040 585
R4273 gnd.n4346 gnd.n4345 585
R4274 gnd.n4345 gnd.n4344 585
R4275 gnd.n2046 gnd.n2045 585
R4276 gnd.n2047 gnd.n2046 585
R4277 gnd.n4335 gnd.n4334 585
R4278 gnd.n4336 gnd.n4335 585
R4279 gnd.n2057 gnd.n2056 585
R4280 gnd.n2056 gnd.n2054 585
R4281 gnd.n4330 gnd.n4329 585
R4282 gnd.n4329 gnd.n4328 585
R4283 gnd.n2060 gnd.n2059 585
R4284 gnd.n2069 gnd.n2060 585
R4285 gnd.n4319 gnd.n4318 585
R4286 gnd.n4320 gnd.n4319 585
R4287 gnd.n2071 gnd.n2070 585
R4288 gnd.n2070 gnd.n2067 585
R4289 gnd.n4314 gnd.n4313 585
R4290 gnd.n4313 gnd.n4312 585
R4291 gnd.n2074 gnd.n2073 585
R4292 gnd.n2075 gnd.n2074 585
R4293 gnd.n4303 gnd.n4302 585
R4294 gnd.n4304 gnd.n4303 585
R4295 gnd.n4299 gnd.n875 585
R4296 gnd.n4228 gnd.n875 585
R4297 gnd.n5506 gnd.n1365 585
R4298 gnd.n5170 gnd.n1365 585
R4299 gnd.n5507 gnd.n1364 585
R4300 gnd.n1654 gnd.n1358 585
R4301 gnd.n5514 gnd.n1357 585
R4302 gnd.n5515 gnd.n1356 585
R4303 gnd.n1651 gnd.n1350 585
R4304 gnd.n5522 gnd.n1349 585
R4305 gnd.n5523 gnd.n1348 585
R4306 gnd.n1649 gnd.n1342 585
R4307 gnd.n5530 gnd.n1341 585
R4308 gnd.n5531 gnd.n1340 585
R4309 gnd.n1646 gnd.n1334 585
R4310 gnd.n5538 gnd.n1333 585
R4311 gnd.n5539 gnd.n1332 585
R4312 gnd.n1644 gnd.n1325 585
R4313 gnd.n5546 gnd.n1324 585
R4314 gnd.n5547 gnd.n1323 585
R4315 gnd.n1641 gnd.n1320 585
R4316 gnd.n5552 gnd.n1319 585
R4317 gnd.n5553 gnd.n1318 585
R4318 gnd.n5554 gnd.n1317 585
R4319 gnd.n1638 gnd.n1315 585
R4320 gnd.n5558 gnd.n1314 585
R4321 gnd.n5559 gnd.n1313 585
R4322 gnd.n5560 gnd.n1309 585
R4323 gnd.n5173 gnd.n1304 585
R4324 gnd.n5174 gnd.n5172 585
R4325 gnd.n1636 gnd.n1635 585
R4326 gnd.n1657 gnd.n1656 585
R4327 gnd.n4436 gnd.t5 543.808
R4328 gnd.n1791 gnd.t15 543.808
R4329 gnd.n5683 gnd.t65 543.808
R4330 gnd.n4889 gnd.t9 543.808
R4331 gnd.n6145 gnd.n561 498.228
R4332 gnd.n4955 gnd.n1799 497.305
R4333 gnd.n4964 gnd.n4963 497.305
R4334 gnd.n4501 gnd.n4500 497.305
R4335 gnd.n5746 gnd.n1178 497.305
R4336 gnd.n953 gnd.t45 371.625
R4337 gnd.n5500 gnd.t22 371.625
R4338 gnd.n960 gnd.t38 371.625
R4339 gnd.n1438 gnd.t95 371.625
R4340 gnd.n1461 gnd.t104 371.625
R4341 gnd.n5380 gnd.t68 371.625
R4342 gnd.n6965 gnd.t56 371.625
R4343 gnd.n6944 gnd.t74 371.625
R4344 gnd.n7051 gnd.t83 371.625
R4345 gnd.n6812 gnd.t18 371.625
R4346 gnd.n3772 gnd.t49 371.625
R4347 gnd.n3803 gnd.t89 371.625
R4348 gnd.n3835 gnd.t71 371.625
R4349 gnd.n3672 gnd.t34 371.625
R4350 gnd.n1030 gnd.t77 371.625
R4351 gnd.n1071 gnd.t92 371.625
R4352 gnd.n1050 gnd.t118 371.625
R4353 gnd.n1366 gnd.t30 371.625
R4354 gnd.n2686 gnd.t52 323.425
R4355 gnd.n2244 gnd.t110 323.425
R4356 gnd.n3534 gnd.n3508 289.615
R4357 gnd.n3502 gnd.n3476 289.615
R4358 gnd.n3470 gnd.n3444 289.615
R4359 gnd.n3439 gnd.n3413 289.615
R4360 gnd.n3407 gnd.n3381 289.615
R4361 gnd.n3375 gnd.n3349 289.615
R4362 gnd.n3343 gnd.n3317 289.615
R4363 gnd.n3312 gnd.n3286 289.615
R4364 gnd.n2760 gnd.t114 279.217
R4365 gnd.n2270 gnd.t26 279.217
R4366 gnd.n1185 gnd.t103 260.649
R4367 gnd.n4881 gnd.t61 260.649
R4368 gnd.n5748 gnd.n5747 256.663
R4369 gnd.n5748 gnd.n1144 256.663
R4370 gnd.n5748 gnd.n1145 256.663
R4371 gnd.n5748 gnd.n1146 256.663
R4372 gnd.n5748 gnd.n1147 256.663
R4373 gnd.n5748 gnd.n1148 256.663
R4374 gnd.n5748 gnd.n1149 256.663
R4375 gnd.n5748 gnd.n1150 256.663
R4376 gnd.n5748 gnd.n1151 256.663
R4377 gnd.n5748 gnd.n1152 256.663
R4378 gnd.n5748 gnd.n1153 256.663
R4379 gnd.n5748 gnd.n1154 256.663
R4380 gnd.n5748 gnd.n1155 256.663
R4381 gnd.n5748 gnd.n1156 256.663
R4382 gnd.n5748 gnd.n1157 256.663
R4383 gnd.n5748 gnd.n1158 256.663
R4384 gnd.n5751 gnd.n1141 256.663
R4385 gnd.n5749 gnd.n5748 256.663
R4386 gnd.n5748 gnd.n1159 256.663
R4387 gnd.n5748 gnd.n1160 256.663
R4388 gnd.n5748 gnd.n1161 256.663
R4389 gnd.n5748 gnd.n1162 256.663
R4390 gnd.n5748 gnd.n1163 256.663
R4391 gnd.n5748 gnd.n1164 256.663
R4392 gnd.n5748 gnd.n1165 256.663
R4393 gnd.n5748 gnd.n1166 256.663
R4394 gnd.n5748 gnd.n1167 256.663
R4395 gnd.n5748 gnd.n1168 256.663
R4396 gnd.n5748 gnd.n1169 256.663
R4397 gnd.n5748 gnd.n1170 256.663
R4398 gnd.n5748 gnd.n1171 256.663
R4399 gnd.n5748 gnd.n1172 256.663
R4400 gnd.n5748 gnd.n1173 256.663
R4401 gnd.n5748 gnd.n1174 256.663
R4402 gnd.n5030 gnd.n1774 256.663
R4403 gnd.n5030 gnd.n1775 256.663
R4404 gnd.n5030 gnd.n1776 256.663
R4405 gnd.n5030 gnd.n1777 256.663
R4406 gnd.n5030 gnd.n1778 256.663
R4407 gnd.n5030 gnd.n1779 256.663
R4408 gnd.n5030 gnd.n1780 256.663
R4409 gnd.n5030 gnd.n1781 256.663
R4410 gnd.n5030 gnd.n1782 256.663
R4411 gnd.n5030 gnd.n1783 256.663
R4412 gnd.n5030 gnd.n1784 256.663
R4413 gnd.n5030 gnd.n1785 256.663
R4414 gnd.n5030 gnd.n1786 256.663
R4415 gnd.n5030 gnd.n1787 256.663
R4416 gnd.n5030 gnd.n1788 256.663
R4417 gnd.n5030 gnd.n1789 256.663
R4418 gnd.n1790 gnd.n1448 256.663
R4419 gnd.n5030 gnd.n1773 256.663
R4420 gnd.n5030 gnd.n1772 256.663
R4421 gnd.n5030 gnd.n1771 256.663
R4422 gnd.n5030 gnd.n1770 256.663
R4423 gnd.n5030 gnd.n1769 256.663
R4424 gnd.n5030 gnd.n1768 256.663
R4425 gnd.n5030 gnd.n1767 256.663
R4426 gnd.n5030 gnd.n1766 256.663
R4427 gnd.n5030 gnd.n1765 256.663
R4428 gnd.n5030 gnd.n1764 256.663
R4429 gnd.n5030 gnd.n1763 256.663
R4430 gnd.n5030 gnd.n1762 256.663
R4431 gnd.n5030 gnd.n1761 256.663
R4432 gnd.n5030 gnd.n1760 256.663
R4433 gnd.n5030 gnd.n1759 256.663
R4434 gnd.n5030 gnd.n1758 256.663
R4435 gnd.n5030 gnd.n1757 256.663
R4436 gnd.n3693 gnd.n3667 242.672
R4437 gnd.n3695 gnd.n3667 242.672
R4438 gnd.n3703 gnd.n3667 242.672
R4439 gnd.n3705 gnd.n3667 242.672
R4440 gnd.n3713 gnd.n3667 242.672
R4441 gnd.n3715 gnd.n3667 242.672
R4442 gnd.n3723 gnd.n3667 242.672
R4443 gnd.n3725 gnd.n3667 242.672
R4444 gnd.n3733 gnd.n3667 242.672
R4445 gnd.n5803 gnd.n5802 242.672
R4446 gnd.n5802 gnd.n978 242.672
R4447 gnd.n5802 gnd.n976 242.672
R4448 gnd.n5802 gnd.n975 242.672
R4449 gnd.n5802 gnd.n973 242.672
R4450 gnd.n5802 gnd.n971 242.672
R4451 gnd.n5802 gnd.n970 242.672
R4452 gnd.n5802 gnd.n968 242.672
R4453 gnd.n5802 gnd.n966 242.672
R4454 gnd.n2814 gnd.n2813 242.672
R4455 gnd.n2814 gnd.n2724 242.672
R4456 gnd.n2814 gnd.n2725 242.672
R4457 gnd.n2814 gnd.n2726 242.672
R4458 gnd.n2814 gnd.n2727 242.672
R4459 gnd.n2814 gnd.n2728 242.672
R4460 gnd.n2814 gnd.n2729 242.672
R4461 gnd.n2814 gnd.n2730 242.672
R4462 gnd.n2814 gnd.n2731 242.672
R4463 gnd.n2814 gnd.n2732 242.672
R4464 gnd.n2814 gnd.n2733 242.672
R4465 gnd.n2814 gnd.n2734 242.672
R4466 gnd.n2815 gnd.n2814 242.672
R4467 gnd.n3666 gnd.n2219 242.672
R4468 gnd.n3666 gnd.n2218 242.672
R4469 gnd.n3666 gnd.n2217 242.672
R4470 gnd.n3666 gnd.n2216 242.672
R4471 gnd.n3666 gnd.n2215 242.672
R4472 gnd.n3666 gnd.n2214 242.672
R4473 gnd.n3666 gnd.n2213 242.672
R4474 gnd.n3666 gnd.n2212 242.672
R4475 gnd.n3666 gnd.n2211 242.672
R4476 gnd.n3666 gnd.n2210 242.672
R4477 gnd.n3666 gnd.n2209 242.672
R4478 gnd.n3666 gnd.n2208 242.672
R4479 gnd.n3666 gnd.n2207 242.672
R4480 gnd.n5497 gnd.n1403 242.672
R4481 gnd.n5497 gnd.n1405 242.672
R4482 gnd.n5497 gnd.n1406 242.672
R4483 gnd.n5497 gnd.n1408 242.672
R4484 gnd.n5497 gnd.n1410 242.672
R4485 gnd.n5497 gnd.n1411 242.672
R4486 gnd.n5497 gnd.n1413 242.672
R4487 gnd.n5497 gnd.n1415 242.672
R4488 gnd.n5498 gnd.n5497 242.672
R4489 gnd.n7087 gnd.n7086 242.672
R4490 gnd.n7086 gnd.n6873 242.672
R4491 gnd.n7086 gnd.n6822 242.672
R4492 gnd.n7086 gnd.n6821 242.672
R4493 gnd.n7086 gnd.n6820 242.672
R4494 gnd.n7086 gnd.n6819 242.672
R4495 gnd.n7086 gnd.n6818 242.672
R4496 gnd.n7086 gnd.n6817 242.672
R4497 gnd.n7086 gnd.n6816 242.672
R4498 gnd.n2898 gnd.n2897 242.672
R4499 gnd.n2897 gnd.n2636 242.672
R4500 gnd.n2897 gnd.n2637 242.672
R4501 gnd.n2897 gnd.n2638 242.672
R4502 gnd.n2897 gnd.n2639 242.672
R4503 gnd.n2897 gnd.n2640 242.672
R4504 gnd.n2897 gnd.n2641 242.672
R4505 gnd.n2897 gnd.n2642 242.672
R4506 gnd.n3666 gnd.n2220 242.672
R4507 gnd.n3666 gnd.n2221 242.672
R4508 gnd.n3666 gnd.n2222 242.672
R4509 gnd.n3666 gnd.n2223 242.672
R4510 gnd.n3666 gnd.n2224 242.672
R4511 gnd.n3666 gnd.n2225 242.672
R4512 gnd.n3666 gnd.n2226 242.672
R4513 gnd.n3666 gnd.n2227 242.672
R4514 gnd.n3953 gnd.n3667 242.672
R4515 gnd.n3748 gnd.n3667 242.672
R4516 gnd.n3946 gnd.n3667 242.672
R4517 gnd.n3940 gnd.n3667 242.672
R4518 gnd.n3938 gnd.n3667 242.672
R4519 gnd.n3932 gnd.n3667 242.672
R4520 gnd.n3930 gnd.n3667 242.672
R4521 gnd.n3924 gnd.n3667 242.672
R4522 gnd.n3922 gnd.n3667 242.672
R4523 gnd.n3916 gnd.n3667 242.672
R4524 gnd.n3914 gnd.n3667 242.672
R4525 gnd.n3908 gnd.n3667 242.672
R4526 gnd.n3906 gnd.n3667 242.672
R4527 gnd.n3900 gnd.n3667 242.672
R4528 gnd.n3898 gnd.n3667 242.672
R4529 gnd.n3892 gnd.n3667 242.672
R4530 gnd.n3890 gnd.n3667 242.672
R4531 gnd.n3884 gnd.n3667 242.672
R4532 gnd.n3882 gnd.n3667 242.672
R4533 gnd.n3876 gnd.n3667 242.672
R4534 gnd.n3874 gnd.n3667 242.672
R4535 gnd.n3868 gnd.n3667 242.672
R4536 gnd.n3866 gnd.n3667 242.672
R4537 gnd.n3860 gnd.n3667 242.672
R4538 gnd.n3858 gnd.n3667 242.672
R4539 gnd.n3852 gnd.n3667 242.672
R4540 gnd.n3850 gnd.n3667 242.672
R4541 gnd.n3844 gnd.n3667 242.672
R4542 gnd.n3842 gnd.n3667 242.672
R4543 gnd.n5802 gnd.n980 242.672
R4544 gnd.n5802 gnd.n981 242.672
R4545 gnd.n5802 gnd.n982 242.672
R4546 gnd.n5802 gnd.n983 242.672
R4547 gnd.n5802 gnd.n984 242.672
R4548 gnd.n5802 gnd.n985 242.672
R4549 gnd.n5802 gnd.n986 242.672
R4550 gnd.n5802 gnd.n987 242.672
R4551 gnd.n5802 gnd.n988 242.672
R4552 gnd.n5802 gnd.n989 242.672
R4553 gnd.n5802 gnd.n990 242.672
R4554 gnd.n5802 gnd.n991 242.672
R4555 gnd.n5802 gnd.n992 242.672
R4556 gnd.n5802 gnd.n993 242.672
R4557 gnd.n5802 gnd.n994 242.672
R4558 gnd.n5802 gnd.n995 242.672
R4559 gnd.n5752 gnd.n1041 242.672
R4560 gnd.n5802 gnd.n996 242.672
R4561 gnd.n5802 gnd.n997 242.672
R4562 gnd.n5802 gnd.n998 242.672
R4563 gnd.n5802 gnd.n999 242.672
R4564 gnd.n5802 gnd.n1000 242.672
R4565 gnd.n5802 gnd.n1001 242.672
R4566 gnd.n5802 gnd.n1002 242.672
R4567 gnd.n5802 gnd.n1003 242.672
R4568 gnd.n5802 gnd.n1004 242.672
R4569 gnd.n5802 gnd.n1005 242.672
R4570 gnd.n5802 gnd.n1006 242.672
R4571 gnd.n5802 gnd.n1007 242.672
R4572 gnd.n5802 gnd.n5801 242.672
R4573 gnd.n5497 gnd.n5496 242.672
R4574 gnd.n5497 gnd.n1375 242.672
R4575 gnd.n5497 gnd.n1376 242.672
R4576 gnd.n5497 gnd.n1377 242.672
R4577 gnd.n5497 gnd.n1378 242.672
R4578 gnd.n5497 gnd.n1379 242.672
R4579 gnd.n5497 gnd.n1380 242.672
R4580 gnd.n5497 gnd.n1381 242.672
R4581 gnd.n5497 gnd.n1382 242.672
R4582 gnd.n5497 gnd.n1383 242.672
R4583 gnd.n5497 gnd.n1384 242.672
R4584 gnd.n5497 gnd.n1385 242.672
R4585 gnd.n5497 gnd.n1386 242.672
R4586 gnd.n5444 gnd.n1449 242.672
R4587 gnd.n5497 gnd.n1387 242.672
R4588 gnd.n5497 gnd.n1388 242.672
R4589 gnd.n5497 gnd.n1389 242.672
R4590 gnd.n5497 gnd.n1390 242.672
R4591 gnd.n5497 gnd.n1391 242.672
R4592 gnd.n5497 gnd.n1392 242.672
R4593 gnd.n5497 gnd.n1393 242.672
R4594 gnd.n5497 gnd.n1394 242.672
R4595 gnd.n5497 gnd.n1395 242.672
R4596 gnd.n5497 gnd.n1396 242.672
R4597 gnd.n5497 gnd.n1397 242.672
R4598 gnd.n5497 gnd.n1398 242.672
R4599 gnd.n5497 gnd.n1399 242.672
R4600 gnd.n5497 gnd.n1400 242.672
R4601 gnd.n5497 gnd.n1401 242.672
R4602 gnd.n5497 gnd.n1402 242.672
R4603 gnd.n7086 gnd.n6874 242.672
R4604 gnd.n7086 gnd.n6875 242.672
R4605 gnd.n7086 gnd.n6876 242.672
R4606 gnd.n7086 gnd.n6877 242.672
R4607 gnd.n7086 gnd.n6878 242.672
R4608 gnd.n7086 gnd.n6879 242.672
R4609 gnd.n7086 gnd.n6880 242.672
R4610 gnd.n7086 gnd.n6881 242.672
R4611 gnd.n7086 gnd.n6882 242.672
R4612 gnd.n7086 gnd.n6883 242.672
R4613 gnd.n7086 gnd.n6884 242.672
R4614 gnd.n7086 gnd.n6885 242.672
R4615 gnd.n7086 gnd.n6886 242.672
R4616 gnd.n7086 gnd.n6887 242.672
R4617 gnd.n7086 gnd.n6888 242.672
R4618 gnd.n7086 gnd.n6889 242.672
R4619 gnd.n7086 gnd.n6890 242.672
R4620 gnd.n7086 gnd.n6891 242.672
R4621 gnd.n7086 gnd.n6892 242.672
R4622 gnd.n7086 gnd.n6893 242.672
R4623 gnd.n7086 gnd.n6894 242.672
R4624 gnd.n7086 gnd.n6895 242.672
R4625 gnd.n7086 gnd.n6896 242.672
R4626 gnd.n7086 gnd.n6897 242.672
R4627 gnd.n7086 gnd.n6898 242.672
R4628 gnd.n7086 gnd.n6899 242.672
R4629 gnd.n7086 gnd.n6900 242.672
R4630 gnd.n7086 gnd.n6901 242.672
R4631 gnd.n7086 gnd.n7085 242.672
R4632 gnd.n5867 gnd.n5866 242.672
R4633 gnd.n5867 gnd.n877 242.672
R4634 gnd.n5867 gnd.n878 242.672
R4635 gnd.n5867 gnd.n879 242.672
R4636 gnd.n5867 gnd.n880 242.672
R4637 gnd.n5867 gnd.n881 242.672
R4638 gnd.n5867 gnd.n882 242.672
R4639 gnd.n5867 gnd.n883 242.672
R4640 gnd.n5867 gnd.n884 242.672
R4641 gnd.n5867 gnd.n885 242.672
R4642 gnd.n5867 gnd.n886 242.672
R4643 gnd.n5867 gnd.n887 242.672
R4644 gnd.n5867 gnd.n889 242.672
R4645 gnd.n5868 gnd.n5867 242.672
R4646 gnd.n5170 gnd.n1655 242.672
R4647 gnd.n5170 gnd.n1653 242.672
R4648 gnd.n5170 gnd.n1652 242.672
R4649 gnd.n5170 gnd.n1650 242.672
R4650 gnd.n5170 gnd.n1648 242.672
R4651 gnd.n5170 gnd.n1647 242.672
R4652 gnd.n5170 gnd.n1645 242.672
R4653 gnd.n5170 gnd.n1643 242.672
R4654 gnd.n5170 gnd.n1642 242.672
R4655 gnd.n5170 gnd.n1640 242.672
R4656 gnd.n5170 gnd.n1639 242.672
R4657 gnd.n5170 gnd.n1637 242.672
R4658 gnd.n5171 gnd.n5170 242.672
R4659 gnd.n5170 gnd.n1658 242.672
R4660 gnd.n6902 gnd.n166 240.244
R4661 gnd.n7084 gnd.n6903 240.244
R4662 gnd.n7080 gnd.n7079 240.244
R4663 gnd.n7076 gnd.n7075 240.244
R4664 gnd.n7072 gnd.n7071 240.244
R4665 gnd.n7068 gnd.n7067 240.244
R4666 gnd.n7064 gnd.n7063 240.244
R4667 gnd.n7060 gnd.n7059 240.244
R4668 gnd.n7056 gnd.n7055 240.244
R4669 gnd.n7049 gnd.n7048 240.244
R4670 gnd.n7045 gnd.n7044 240.244
R4671 gnd.n7041 gnd.n7040 240.244
R4672 gnd.n7037 gnd.n7036 240.244
R4673 gnd.n7033 gnd.n7032 240.244
R4674 gnd.n7029 gnd.n7028 240.244
R4675 gnd.n7025 gnd.n7024 240.244
R4676 gnd.n7021 gnd.n7020 240.244
R4677 gnd.n7017 gnd.n7016 240.244
R4678 gnd.n7013 gnd.n7012 240.244
R4679 gnd.n7006 gnd.n7005 240.244
R4680 gnd.n7003 gnd.n7002 240.244
R4681 gnd.n6999 gnd.n6998 240.244
R4682 gnd.n6995 gnd.n6994 240.244
R4683 gnd.n6991 gnd.n6990 240.244
R4684 gnd.n6987 gnd.n6986 240.244
R4685 gnd.n6983 gnd.n6982 240.244
R4686 gnd.n6979 gnd.n6978 240.244
R4687 gnd.n6975 gnd.n6974 240.244
R4688 gnd.n6971 gnd.n6970 240.244
R4689 gnd.n5377 gnd.n1482 240.244
R4690 gnd.n5369 gnd.n1482 240.244
R4691 gnd.n5369 gnd.n1493 240.244
R4692 gnd.n1509 gnd.n1493 240.244
R4693 gnd.n5187 gnd.n1509 240.244
R4694 gnd.n5187 gnd.n1522 240.244
R4695 gnd.n5193 gnd.n1522 240.244
R4696 gnd.n5193 gnd.n1532 240.244
R4697 gnd.n5200 gnd.n1532 240.244
R4698 gnd.n5200 gnd.n1542 240.244
R4699 gnd.n1615 gnd.n1542 240.244
R4700 gnd.n1615 gnd.n1552 240.244
R4701 gnd.n5270 gnd.n1552 240.244
R4702 gnd.n5270 gnd.n1562 240.244
R4703 gnd.n5275 gnd.n1562 240.244
R4704 gnd.n5275 gnd.n1569 240.244
R4705 gnd.n5289 gnd.n1569 240.244
R4706 gnd.n5289 gnd.n1579 240.244
R4707 gnd.n1585 gnd.n1579 240.244
R4708 gnd.n5298 gnd.n1585 240.244
R4709 gnd.n5299 gnd.n5298 240.244
R4710 gnd.n5299 gnd.n1597 240.244
R4711 gnd.n1597 gnd.n74 240.244
R4712 gnd.n177 gnd.n74 240.244
R4713 gnd.n6790 gnd.n177 240.244
R4714 gnd.n6790 gnd.n91 240.244
R4715 gnd.n7117 gnd.n91 240.244
R4716 gnd.n7117 gnd.n102 240.244
R4717 gnd.n7121 gnd.n102 240.244
R4718 gnd.n7121 gnd.n112 240.244
R4719 gnd.n7124 gnd.n112 240.244
R4720 gnd.n7124 gnd.n121 240.244
R4721 gnd.n7128 gnd.n121 240.244
R4722 gnd.n7128 gnd.n131 240.244
R4723 gnd.n7131 gnd.n131 240.244
R4724 gnd.n7131 gnd.n140 240.244
R4725 gnd.n7135 gnd.n140 240.244
R4726 gnd.n7135 gnd.n150 240.244
R4727 gnd.n7138 gnd.n150 240.244
R4728 gnd.n7138 gnd.n159 240.244
R4729 gnd.n7141 gnd.n159 240.244
R4730 gnd.n7141 gnd.n168 240.244
R4731 gnd.n1418 gnd.n1417 240.244
R4732 gnd.n5490 gnd.n1417 240.244
R4733 gnd.n5488 gnd.n5487 240.244
R4734 gnd.n5484 gnd.n5483 240.244
R4735 gnd.n5480 gnd.n5479 240.244
R4736 gnd.n5476 gnd.n5475 240.244
R4737 gnd.n5472 gnd.n5471 240.244
R4738 gnd.n5468 gnd.n5467 240.244
R4739 gnd.n5464 gnd.n5463 240.244
R4740 gnd.n5459 gnd.n5458 240.244
R4741 gnd.n5455 gnd.n5454 240.244
R4742 gnd.n5451 gnd.n5450 240.244
R4743 gnd.n5447 gnd.n5446 240.244
R4744 gnd.n5442 gnd.n5441 240.244
R4745 gnd.n5438 gnd.n5437 240.244
R4746 gnd.n5434 gnd.n5433 240.244
R4747 gnd.n5430 gnd.n5429 240.244
R4748 gnd.n5426 gnd.n5425 240.244
R4749 gnd.n5422 gnd.n5421 240.244
R4750 gnd.n5418 gnd.n5417 240.244
R4751 gnd.n5414 gnd.n5413 240.244
R4752 gnd.n5410 gnd.n5409 240.244
R4753 gnd.n5406 gnd.n5405 240.244
R4754 gnd.n5402 gnd.n5401 240.244
R4755 gnd.n5398 gnd.n5397 240.244
R4756 gnd.n5394 gnd.n5393 240.244
R4757 gnd.n5390 gnd.n5389 240.244
R4758 gnd.n5386 gnd.n5385 240.244
R4759 gnd.n1497 gnd.n1419 240.244
R4760 gnd.n5367 gnd.n1497 240.244
R4761 gnd.n5367 gnd.n1498 240.244
R4762 gnd.n5363 gnd.n1498 240.244
R4763 gnd.n5363 gnd.n1507 240.244
R4764 gnd.n5355 gnd.n1507 240.244
R4765 gnd.n5355 gnd.n1524 240.244
R4766 gnd.n5351 gnd.n1524 240.244
R4767 gnd.n5351 gnd.n1530 240.244
R4768 gnd.n5343 gnd.n1530 240.244
R4769 gnd.n5343 gnd.n1545 240.244
R4770 gnd.n5339 gnd.n1545 240.244
R4771 gnd.n5339 gnd.n1551 240.244
R4772 gnd.n5331 gnd.n1551 240.244
R4773 gnd.n5331 gnd.n1564 240.244
R4774 gnd.n5327 gnd.n1564 240.244
R4775 gnd.n5327 gnd.n1567 240.244
R4776 gnd.n5319 gnd.n1567 240.244
R4777 gnd.n5319 gnd.n5316 240.244
R4778 gnd.n5316 gnd.n1582 240.244
R4779 gnd.n1595 gnd.n1582 240.244
R4780 gnd.n1595 gnd.n77 240.244
R4781 gnd.n7202 gnd.n77 240.244
R4782 gnd.n7202 gnd.n78 240.244
R4783 gnd.n88 gnd.n78 240.244
R4784 gnd.n7196 gnd.n88 240.244
R4785 gnd.n7196 gnd.n89 240.244
R4786 gnd.n7188 gnd.n89 240.244
R4787 gnd.n7188 gnd.n105 240.244
R4788 gnd.n7184 gnd.n105 240.244
R4789 gnd.n7184 gnd.n110 240.244
R4790 gnd.n7176 gnd.n110 240.244
R4791 gnd.n7176 gnd.n123 240.244
R4792 gnd.n7172 gnd.n123 240.244
R4793 gnd.n7172 gnd.n129 240.244
R4794 gnd.n7164 gnd.n129 240.244
R4795 gnd.n7164 gnd.n143 240.244
R4796 gnd.n7160 gnd.n143 240.244
R4797 gnd.n7160 gnd.n149 240.244
R4798 gnd.n7152 gnd.n149 240.244
R4799 gnd.n7152 gnd.n161 240.244
R4800 gnd.n7148 gnd.n161 240.244
R4801 gnd.n1008 gnd.n858 240.244
R4802 gnd.n5800 gnd.n1009 240.244
R4803 gnd.n5796 gnd.n5795 240.244
R4804 gnd.n5792 gnd.n5791 240.244
R4805 gnd.n5788 gnd.n5787 240.244
R4806 gnd.n5784 gnd.n5783 240.244
R4807 gnd.n5780 gnd.n5779 240.244
R4808 gnd.n5776 gnd.n5775 240.244
R4809 gnd.n5772 gnd.n5771 240.244
R4810 gnd.n5767 gnd.n5766 240.244
R4811 gnd.n5763 gnd.n5762 240.244
R4812 gnd.n5759 gnd.n5758 240.244
R4813 gnd.n5755 gnd.n5754 240.244
R4814 gnd.n1134 gnd.n1133 240.244
R4815 gnd.n1131 gnd.n1130 240.244
R4816 gnd.n1127 gnd.n1126 240.244
R4817 gnd.n1123 gnd.n1122 240.244
R4818 gnd.n1119 gnd.n1118 240.244
R4819 gnd.n1112 gnd.n1111 240.244
R4820 gnd.n1109 gnd.n1108 240.244
R4821 gnd.n1105 gnd.n1104 240.244
R4822 gnd.n1101 gnd.n1100 240.244
R4823 gnd.n1097 gnd.n1096 240.244
R4824 gnd.n1093 gnd.n1092 240.244
R4825 gnd.n1089 gnd.n1088 240.244
R4826 gnd.n1085 gnd.n1084 240.244
R4827 gnd.n1081 gnd.n1080 240.244
R4828 gnd.n1077 gnd.n1076 240.244
R4829 gnd.n3668 gnd.n2202 240.244
R4830 gnd.n2202 gnd.n2194 240.244
R4831 gnd.n3968 gnd.n2194 240.244
R4832 gnd.n3968 gnd.n2186 240.244
R4833 gnd.n2186 gnd.n2178 240.244
R4834 gnd.n4000 gnd.n2178 240.244
R4835 gnd.n4000 gnd.n2169 240.244
R4836 gnd.n4003 gnd.n2169 240.244
R4837 gnd.n4003 gnd.n2161 240.244
R4838 gnd.n2161 gnd.n2153 240.244
R4839 gnd.n4037 gnd.n2153 240.244
R4840 gnd.n4037 gnd.n2142 240.244
R4841 gnd.n4040 gnd.n2142 240.244
R4842 gnd.n4040 gnd.n2135 240.244
R4843 gnd.n4043 gnd.n2135 240.244
R4844 gnd.n4043 gnd.n734 240.244
R4845 gnd.n4073 gnd.n734 240.244
R4846 gnd.n4073 gnd.n745 240.244
R4847 gnd.n4077 gnd.n745 240.244
R4848 gnd.n4077 gnd.n756 240.244
R4849 gnd.n4099 gnd.n756 240.244
R4850 gnd.n4099 gnd.n764 240.244
R4851 gnd.n2119 gnd.n764 240.244
R4852 gnd.n2119 gnd.n773 240.244
R4853 gnd.n4108 gnd.n773 240.244
R4854 gnd.n4108 gnd.n781 240.244
R4855 gnd.n2112 gnd.n781 240.244
R4856 gnd.n2112 gnd.n790 240.244
R4857 gnd.n4162 gnd.n790 240.244
R4858 gnd.n4162 gnd.n801 240.244
R4859 gnd.n4166 gnd.n801 240.244
R4860 gnd.n4166 gnd.n810 240.244
R4861 gnd.n4176 gnd.n810 240.244
R4862 gnd.n4176 gnd.n821 240.244
R4863 gnd.n2095 gnd.n821 240.244
R4864 gnd.n2095 gnd.n830 240.244
R4865 gnd.n4183 gnd.n830 240.244
R4866 gnd.n4183 gnd.n841 240.244
R4867 gnd.n4187 gnd.n841 240.244
R4868 gnd.n4187 gnd.n851 240.244
R4869 gnd.n5879 gnd.n851 240.244
R4870 gnd.n5879 gnd.n860 240.244
R4871 gnd.n3954 gnd.n3952 240.244
R4872 gnd.n3952 gnd.n3951 240.244
R4873 gnd.n3948 gnd.n3947 240.244
R4874 gnd.n3945 gnd.n3753 240.244
R4875 gnd.n3941 gnd.n3939 240.244
R4876 gnd.n3937 gnd.n3759 240.244
R4877 gnd.n3933 gnd.n3931 240.244
R4878 gnd.n3929 gnd.n3765 240.244
R4879 gnd.n3925 gnd.n3923 240.244
R4880 gnd.n3921 gnd.n3771 240.244
R4881 gnd.n3917 gnd.n3915 240.244
R4882 gnd.n3913 gnd.n3780 240.244
R4883 gnd.n3909 gnd.n3907 240.244
R4884 gnd.n3905 gnd.n3786 240.244
R4885 gnd.n3901 gnd.n3899 240.244
R4886 gnd.n3897 gnd.n3792 240.244
R4887 gnd.n3893 gnd.n3891 240.244
R4888 gnd.n3889 gnd.n3798 240.244
R4889 gnd.n3885 gnd.n3883 240.244
R4890 gnd.n3881 gnd.n3806 240.244
R4891 gnd.n3877 gnd.n3875 240.244
R4892 gnd.n3873 gnd.n3812 240.244
R4893 gnd.n3869 gnd.n3867 240.244
R4894 gnd.n3865 gnd.n3818 240.244
R4895 gnd.n3861 gnd.n3859 240.244
R4896 gnd.n3857 gnd.n3824 240.244
R4897 gnd.n3853 gnd.n3851 240.244
R4898 gnd.n3849 gnd.n3830 240.244
R4899 gnd.n3845 gnd.n3843 240.244
R4900 gnd.n3960 gnd.n2193 240.244
R4901 gnd.n3980 gnd.n2193 240.244
R4902 gnd.n3980 gnd.n2188 240.244
R4903 gnd.n3988 gnd.n2188 240.244
R4904 gnd.n3988 gnd.n2189 240.244
R4905 gnd.n2189 gnd.n2168 240.244
R4906 gnd.n4015 gnd.n2168 240.244
R4907 gnd.n4015 gnd.n2163 240.244
R4908 gnd.n4023 gnd.n2163 240.244
R4909 gnd.n4023 gnd.n2164 240.244
R4910 gnd.n2164 gnd.n2141 240.244
R4911 gnd.n4055 gnd.n2141 240.244
R4912 gnd.n4055 gnd.n2137 240.244
R4913 gnd.n4062 gnd.n2137 240.244
R4914 gnd.n4062 gnd.n738 240.244
R4915 gnd.n5965 gnd.n738 240.244
R4916 gnd.n5965 gnd.n739 240.244
R4917 gnd.n5960 gnd.n739 240.244
R4918 gnd.n5960 gnd.n743 240.244
R4919 gnd.n5952 gnd.n743 240.244
R4920 gnd.n5952 gnd.n759 240.244
R4921 gnd.n5947 gnd.n759 240.244
R4922 gnd.n5947 gnd.n762 240.244
R4923 gnd.n5939 gnd.n762 240.244
R4924 gnd.n5939 gnd.n776 240.244
R4925 gnd.n5934 gnd.n776 240.244
R4926 gnd.n5934 gnd.n779 240.244
R4927 gnd.n5926 gnd.n779 240.244
R4928 gnd.n5926 gnd.n793 240.244
R4929 gnd.n5922 gnd.n793 240.244
R4930 gnd.n5922 gnd.n799 240.244
R4931 gnd.n5914 gnd.n799 240.244
R4932 gnd.n5914 gnd.n813 240.244
R4933 gnd.n5910 gnd.n813 240.244
R4934 gnd.n5910 gnd.n819 240.244
R4935 gnd.n5902 gnd.n819 240.244
R4936 gnd.n5902 gnd.n833 240.244
R4937 gnd.n5898 gnd.n833 240.244
R4938 gnd.n5898 gnd.n839 240.244
R4939 gnd.n5890 gnd.n839 240.244
R4940 gnd.n5890 gnd.n853 240.244
R4941 gnd.n5886 gnd.n853 240.244
R4942 gnd.n3665 gnd.n2229 240.244
R4943 gnd.n3658 gnd.n3657 240.244
R4944 gnd.n3655 gnd.n3654 240.244
R4945 gnd.n3651 gnd.n3650 240.244
R4946 gnd.n3647 gnd.n3646 240.244
R4947 gnd.n3643 gnd.n3642 240.244
R4948 gnd.n3639 gnd.n3638 240.244
R4949 gnd.n3635 gnd.n3634 240.244
R4950 gnd.n2909 gnd.n2621 240.244
R4951 gnd.n2919 gnd.n2621 240.244
R4952 gnd.n2919 gnd.n2612 240.244
R4953 gnd.n2612 gnd.n2601 240.244
R4954 gnd.n2940 gnd.n2601 240.244
R4955 gnd.n2940 gnd.n2595 240.244
R4956 gnd.n2950 gnd.n2595 240.244
R4957 gnd.n2950 gnd.n2584 240.244
R4958 gnd.n2584 gnd.n2576 240.244
R4959 gnd.n2968 gnd.n2576 240.244
R4960 gnd.n2969 gnd.n2968 240.244
R4961 gnd.n2969 gnd.n2561 240.244
R4962 gnd.n2971 gnd.n2561 240.244
R4963 gnd.n2971 gnd.n2547 240.244
R4964 gnd.n3013 gnd.n2547 240.244
R4965 gnd.n3014 gnd.n3013 240.244
R4966 gnd.n3017 gnd.n3014 240.244
R4967 gnd.n3017 gnd.n2502 240.244
R4968 gnd.n2542 gnd.n2502 240.244
R4969 gnd.n2542 gnd.n2512 240.244
R4970 gnd.n3027 gnd.n2512 240.244
R4971 gnd.n3027 gnd.n2533 240.244
R4972 gnd.n3037 gnd.n2533 240.244
R4973 gnd.n3037 gnd.n2431 240.244
R4974 gnd.n3082 gnd.n2431 240.244
R4975 gnd.n3082 gnd.n2417 240.244
R4976 gnd.n3104 gnd.n2417 240.244
R4977 gnd.n3105 gnd.n3104 240.244
R4978 gnd.n3105 gnd.n2404 240.244
R4979 gnd.n2404 gnd.n2393 240.244
R4980 gnd.n3136 gnd.n2393 240.244
R4981 gnd.n3137 gnd.n3136 240.244
R4982 gnd.n3138 gnd.n3137 240.244
R4983 gnd.n3138 gnd.n2378 240.244
R4984 gnd.n2378 gnd.n2377 240.244
R4985 gnd.n2377 gnd.n2362 240.244
R4986 gnd.n3189 gnd.n2362 240.244
R4987 gnd.n3190 gnd.n3189 240.244
R4988 gnd.n3190 gnd.n2349 240.244
R4989 gnd.n2349 gnd.n2338 240.244
R4990 gnd.n3221 gnd.n2338 240.244
R4991 gnd.n3222 gnd.n3221 240.244
R4992 gnd.n3223 gnd.n3222 240.244
R4993 gnd.n3223 gnd.n2322 240.244
R4994 gnd.n2322 gnd.n2321 240.244
R4995 gnd.n2321 gnd.n2308 240.244
R4996 gnd.n3278 gnd.n2308 240.244
R4997 gnd.n3279 gnd.n3278 240.244
R4998 gnd.n3279 gnd.n2295 240.244
R4999 gnd.n2295 gnd.n2285 240.244
R5000 gnd.n3566 gnd.n2285 240.244
R5001 gnd.n3569 gnd.n3566 240.244
R5002 gnd.n3569 gnd.n3568 240.244
R5003 gnd.n2899 gnd.n2634 240.244
R5004 gnd.n2655 gnd.n2634 240.244
R5005 gnd.n2658 gnd.n2657 240.244
R5006 gnd.n2665 gnd.n2664 240.244
R5007 gnd.n2668 gnd.n2667 240.244
R5008 gnd.n2675 gnd.n2674 240.244
R5009 gnd.n2678 gnd.n2677 240.244
R5010 gnd.n2685 gnd.n2684 240.244
R5011 gnd.n2907 gnd.n2631 240.244
R5012 gnd.n2631 gnd.n2610 240.244
R5013 gnd.n2930 gnd.n2610 240.244
R5014 gnd.n2930 gnd.n2604 240.244
R5015 gnd.n2938 gnd.n2604 240.244
R5016 gnd.n2938 gnd.n2606 240.244
R5017 gnd.n2606 gnd.n2582 240.244
R5018 gnd.n2960 gnd.n2582 240.244
R5019 gnd.n2960 gnd.n2578 240.244
R5020 gnd.n2966 gnd.n2578 240.244
R5021 gnd.n2966 gnd.n2560 240.244
R5022 gnd.n2991 gnd.n2560 240.244
R5023 gnd.n2991 gnd.n2555 240.244
R5024 gnd.n3003 gnd.n2555 240.244
R5025 gnd.n3003 gnd.n2556 240.244
R5026 gnd.n2999 gnd.n2556 240.244
R5027 gnd.n2999 gnd.n2504 240.244
R5028 gnd.n3051 gnd.n2504 240.244
R5029 gnd.n3051 gnd.n2505 240.244
R5030 gnd.n3047 gnd.n2505 240.244
R5031 gnd.n3047 gnd.n2511 240.244
R5032 gnd.n2531 gnd.n2511 240.244
R5033 gnd.n2531 gnd.n2429 240.244
R5034 gnd.n3086 gnd.n2429 240.244
R5035 gnd.n3086 gnd.n2424 240.244
R5036 gnd.n3094 gnd.n2424 240.244
R5037 gnd.n3094 gnd.n2425 240.244
R5038 gnd.n2425 gnd.n2402 240.244
R5039 gnd.n3126 gnd.n2402 240.244
R5040 gnd.n3126 gnd.n2397 240.244
R5041 gnd.n3134 gnd.n2397 240.244
R5042 gnd.n3134 gnd.n2398 240.244
R5043 gnd.n2398 gnd.n2375 240.244
R5044 gnd.n3171 gnd.n2375 240.244
R5045 gnd.n3171 gnd.n2370 240.244
R5046 gnd.n3179 gnd.n2370 240.244
R5047 gnd.n3179 gnd.n2371 240.244
R5048 gnd.n2371 gnd.n2347 240.244
R5049 gnd.n3211 gnd.n2347 240.244
R5050 gnd.n3211 gnd.n2342 240.244
R5051 gnd.n3219 gnd.n2342 240.244
R5052 gnd.n3219 gnd.n2343 240.244
R5053 gnd.n2343 gnd.n2320 240.244
R5054 gnd.n3260 gnd.n2320 240.244
R5055 gnd.n3260 gnd.n2315 240.244
R5056 gnd.n3268 gnd.n2315 240.244
R5057 gnd.n3268 gnd.n2316 240.244
R5058 gnd.n2316 gnd.n2293 240.244
R5059 gnd.n3554 gnd.n2293 240.244
R5060 gnd.n3554 gnd.n2288 240.244
R5061 gnd.n3564 gnd.n2288 240.244
R5062 gnd.n3564 gnd.n2289 240.244
R5063 gnd.n2289 gnd.n2228 240.244
R5064 gnd.n6834 gnd.n171 240.244
R5065 gnd.n6837 gnd.n6836 240.244
R5066 gnd.n6844 gnd.n6843 240.244
R5067 gnd.n6847 gnd.n6846 240.244
R5068 gnd.n6854 gnd.n6853 240.244
R5069 gnd.n6857 gnd.n6856 240.244
R5070 gnd.n6864 gnd.n6863 240.244
R5071 gnd.n6866 gnd.n6823 240.244
R5072 gnd.n6872 gnd.n6815 240.244
R5073 gnd.n5217 gnd.n1485 240.244
R5074 gnd.n5217 gnd.n1494 240.244
R5075 gnd.n5180 gnd.n1494 240.244
R5076 gnd.n5180 gnd.n1510 240.244
R5077 gnd.n5181 gnd.n1510 240.244
R5078 gnd.n5181 gnd.n1523 240.244
R5079 gnd.n5184 gnd.n1523 240.244
R5080 gnd.n5184 gnd.n1533 240.244
R5081 gnd.n5202 gnd.n1533 240.244
R5082 gnd.n5202 gnd.n1543 240.244
R5083 gnd.n5262 gnd.n1543 240.244
R5084 gnd.n5262 gnd.n1553 240.244
R5085 gnd.n5268 gnd.n1553 240.244
R5086 gnd.n5268 gnd.n1563 240.244
R5087 gnd.n5277 gnd.n1563 240.244
R5088 gnd.n5277 gnd.n1570 240.244
R5089 gnd.n5287 gnd.n1570 240.244
R5090 gnd.n5287 gnd.n1580 240.244
R5091 gnd.n1586 gnd.n1580 240.244
R5092 gnd.n1603 gnd.n1586 240.244
R5093 gnd.n1603 gnd.n1602 240.244
R5094 gnd.n1602 gnd.n70 240.244
R5095 gnd.n7204 gnd.n70 240.244
R5096 gnd.n7204 gnd.n72 240.244
R5097 gnd.n6792 gnd.n72 240.244
R5098 gnd.n6792 gnd.n92 240.244
R5099 gnd.n7115 gnd.n92 240.244
R5100 gnd.n7115 gnd.n103 240.244
R5101 gnd.n7111 gnd.n103 240.244
R5102 gnd.n7111 gnd.n113 240.244
R5103 gnd.n7108 gnd.n113 240.244
R5104 gnd.n7108 gnd.n122 240.244
R5105 gnd.n7105 gnd.n122 240.244
R5106 gnd.n7105 gnd.n132 240.244
R5107 gnd.n7102 gnd.n132 240.244
R5108 gnd.n7102 gnd.n141 240.244
R5109 gnd.n7099 gnd.n141 240.244
R5110 gnd.n7099 gnd.n151 240.244
R5111 gnd.n7096 gnd.n151 240.244
R5112 gnd.n7096 gnd.n160 240.244
R5113 gnd.n7093 gnd.n160 240.244
R5114 gnd.n7093 gnd.n169 240.244
R5115 gnd.n1329 gnd.n1328 240.244
R5116 gnd.n1404 gnd.n1336 240.244
R5117 gnd.n1407 gnd.n1337 240.244
R5118 gnd.n1345 gnd.n1344 240.244
R5119 gnd.n1409 gnd.n1352 240.244
R5120 gnd.n1412 gnd.n1353 240.244
R5121 gnd.n1361 gnd.n1360 240.244
R5122 gnd.n1414 gnd.n1370 240.244
R5123 gnd.n5499 gnd.n1373 240.244
R5124 gnd.n5375 gnd.n1488 240.244
R5125 gnd.n1496 gnd.n1488 240.244
R5126 gnd.n1512 gnd.n1496 240.244
R5127 gnd.n5361 gnd.n1512 240.244
R5128 gnd.n5361 gnd.n1513 240.244
R5129 gnd.n5357 gnd.n1513 240.244
R5130 gnd.n5357 gnd.n1520 240.244
R5131 gnd.n5349 gnd.n1520 240.244
R5132 gnd.n5349 gnd.n1535 240.244
R5133 gnd.n5345 gnd.n1535 240.244
R5134 gnd.n5345 gnd.n1540 240.244
R5135 gnd.n5337 gnd.n1540 240.244
R5136 gnd.n5337 gnd.n1555 240.244
R5137 gnd.n5333 gnd.n1555 240.244
R5138 gnd.n5333 gnd.n1560 240.244
R5139 gnd.n5325 gnd.n1560 240.244
R5140 gnd.n5325 gnd.n1572 240.244
R5141 gnd.n5321 gnd.n1572 240.244
R5142 gnd.n5321 gnd.n1577 240.244
R5143 gnd.n5296 gnd.n1577 240.244
R5144 gnd.n5296 gnd.n1598 240.244
R5145 gnd.n5305 gnd.n1598 240.244
R5146 gnd.n5305 gnd.n76 240.244
R5147 gnd.n6785 gnd.n76 240.244
R5148 gnd.n6785 gnd.n94 240.244
R5149 gnd.n7194 gnd.n94 240.244
R5150 gnd.n7194 gnd.n95 240.244
R5151 gnd.n7190 gnd.n95 240.244
R5152 gnd.n7190 gnd.n101 240.244
R5153 gnd.n7182 gnd.n101 240.244
R5154 gnd.n7182 gnd.n114 240.244
R5155 gnd.n7178 gnd.n114 240.244
R5156 gnd.n7178 gnd.n119 240.244
R5157 gnd.n7170 gnd.n119 240.244
R5158 gnd.n7170 gnd.n134 240.244
R5159 gnd.n7166 gnd.n134 240.244
R5160 gnd.n7166 gnd.n139 240.244
R5161 gnd.n7158 gnd.n139 240.244
R5162 gnd.n7158 gnd.n153 240.244
R5163 gnd.n7154 gnd.n153 240.244
R5164 gnd.n7154 gnd.n158 240.244
R5165 gnd.n7146 gnd.n158 240.244
R5166 gnd.n2248 gnd.n2206 240.244
R5167 gnd.n3625 gnd.n3624 240.244
R5168 gnd.n3621 gnd.n3620 240.244
R5169 gnd.n3617 gnd.n3616 240.244
R5170 gnd.n3613 gnd.n3612 240.244
R5171 gnd.n3609 gnd.n3608 240.244
R5172 gnd.n3605 gnd.n3604 240.244
R5173 gnd.n3601 gnd.n3600 240.244
R5174 gnd.n3597 gnd.n3596 240.244
R5175 gnd.n3593 gnd.n3592 240.244
R5176 gnd.n3589 gnd.n3588 240.244
R5177 gnd.n3585 gnd.n3584 240.244
R5178 gnd.n3581 gnd.n3580 240.244
R5179 gnd.n2822 gnd.n2719 240.244
R5180 gnd.n2822 gnd.n2712 240.244
R5181 gnd.n2833 gnd.n2712 240.244
R5182 gnd.n2833 gnd.n2708 240.244
R5183 gnd.n2839 gnd.n2708 240.244
R5184 gnd.n2839 gnd.n2700 240.244
R5185 gnd.n2849 gnd.n2700 240.244
R5186 gnd.n2849 gnd.n2695 240.244
R5187 gnd.n2885 gnd.n2695 240.244
R5188 gnd.n2885 gnd.n2696 240.244
R5189 gnd.n2696 gnd.n2643 240.244
R5190 gnd.n2880 gnd.n2643 240.244
R5191 gnd.n2880 gnd.n2879 240.244
R5192 gnd.n2879 gnd.n2622 240.244
R5193 gnd.n2875 gnd.n2622 240.244
R5194 gnd.n2875 gnd.n2613 240.244
R5195 gnd.n2872 gnd.n2613 240.244
R5196 gnd.n2872 gnd.n2871 240.244
R5197 gnd.n2871 gnd.n2596 240.244
R5198 gnd.n2867 gnd.n2596 240.244
R5199 gnd.n2867 gnd.n2585 240.244
R5200 gnd.n2585 gnd.n2566 240.244
R5201 gnd.n2980 gnd.n2566 240.244
R5202 gnd.n2980 gnd.n2562 240.244
R5203 gnd.n2988 gnd.n2562 240.244
R5204 gnd.n2988 gnd.n2553 240.244
R5205 gnd.n2553 gnd.n2489 240.244
R5206 gnd.n3060 gnd.n2489 240.244
R5207 gnd.n3060 gnd.n2490 240.244
R5208 gnd.n2501 gnd.n2490 240.244
R5209 gnd.n2536 gnd.n2501 240.244
R5210 gnd.n2539 gnd.n2536 240.244
R5211 gnd.n2539 gnd.n2513 240.244
R5212 gnd.n2526 gnd.n2513 240.244
R5213 gnd.n2526 gnd.n2523 240.244
R5214 gnd.n2523 gnd.n2432 240.244
R5215 gnd.n3081 gnd.n2432 240.244
R5216 gnd.n3081 gnd.n2422 240.244
R5217 gnd.n3077 gnd.n2422 240.244
R5218 gnd.n3077 gnd.n2416 240.244
R5219 gnd.n3074 gnd.n2416 240.244
R5220 gnd.n3074 gnd.n2405 240.244
R5221 gnd.n3071 gnd.n2405 240.244
R5222 gnd.n3071 gnd.n2383 240.244
R5223 gnd.n3147 gnd.n2383 240.244
R5224 gnd.n3147 gnd.n2379 240.244
R5225 gnd.n3168 gnd.n2379 240.244
R5226 gnd.n3168 gnd.n2368 240.244
R5227 gnd.n3164 gnd.n2368 240.244
R5228 gnd.n3164 gnd.n2361 240.244
R5229 gnd.n3161 gnd.n2361 240.244
R5230 gnd.n3161 gnd.n2350 240.244
R5231 gnd.n3158 gnd.n2350 240.244
R5232 gnd.n3158 gnd.n2327 240.244
R5233 gnd.n3232 gnd.n2327 240.244
R5234 gnd.n3232 gnd.n2323 240.244
R5235 gnd.n3257 gnd.n2323 240.244
R5236 gnd.n3257 gnd.n2314 240.244
R5237 gnd.n3253 gnd.n2314 240.244
R5238 gnd.n3253 gnd.n2307 240.244
R5239 gnd.n3249 gnd.n2307 240.244
R5240 gnd.n3249 gnd.n2296 240.244
R5241 gnd.n3246 gnd.n2296 240.244
R5242 gnd.n3246 gnd.n2277 240.244
R5243 gnd.n3576 gnd.n2277 240.244
R5244 gnd.n2736 gnd.n2735 240.244
R5245 gnd.n2807 gnd.n2735 240.244
R5246 gnd.n2805 gnd.n2804 240.244
R5247 gnd.n2801 gnd.n2800 240.244
R5248 gnd.n2797 gnd.n2796 240.244
R5249 gnd.n2793 gnd.n2792 240.244
R5250 gnd.n2789 gnd.n2788 240.244
R5251 gnd.n2785 gnd.n2784 240.244
R5252 gnd.n2781 gnd.n2780 240.244
R5253 gnd.n2777 gnd.n2776 240.244
R5254 gnd.n2773 gnd.n2772 240.244
R5255 gnd.n2769 gnd.n2768 240.244
R5256 gnd.n2765 gnd.n2723 240.244
R5257 gnd.n2825 gnd.n2717 240.244
R5258 gnd.n2825 gnd.n2713 240.244
R5259 gnd.n2831 gnd.n2713 240.244
R5260 gnd.n2831 gnd.n2706 240.244
R5261 gnd.n2841 gnd.n2706 240.244
R5262 gnd.n2841 gnd.n2702 240.244
R5263 gnd.n2847 gnd.n2702 240.244
R5264 gnd.n2847 gnd.n2693 240.244
R5265 gnd.n2887 gnd.n2693 240.244
R5266 gnd.n2887 gnd.n2644 240.244
R5267 gnd.n2895 gnd.n2644 240.244
R5268 gnd.n2895 gnd.n2645 240.244
R5269 gnd.n2645 gnd.n2623 240.244
R5270 gnd.n2916 gnd.n2623 240.244
R5271 gnd.n2916 gnd.n2615 240.244
R5272 gnd.n2927 gnd.n2615 240.244
R5273 gnd.n2927 gnd.n2616 240.244
R5274 gnd.n2616 gnd.n2597 240.244
R5275 gnd.n2947 gnd.n2597 240.244
R5276 gnd.n2947 gnd.n2587 240.244
R5277 gnd.n2957 gnd.n2587 240.244
R5278 gnd.n2957 gnd.n2568 240.244
R5279 gnd.n2978 gnd.n2568 240.244
R5280 gnd.n2978 gnd.n2570 240.244
R5281 gnd.n2570 gnd.n2551 240.244
R5282 gnd.n3006 gnd.n2551 240.244
R5283 gnd.n3006 gnd.n2493 240.244
R5284 gnd.n3058 gnd.n2493 240.244
R5285 gnd.n3058 gnd.n2494 240.244
R5286 gnd.n3054 gnd.n2494 240.244
R5287 gnd.n3054 gnd.n2500 240.244
R5288 gnd.n2515 gnd.n2500 240.244
R5289 gnd.n3044 gnd.n2515 240.244
R5290 gnd.n3044 gnd.n2516 240.244
R5291 gnd.n3040 gnd.n2516 240.244
R5292 gnd.n3040 gnd.n2522 240.244
R5293 gnd.n2522 gnd.n2421 240.244
R5294 gnd.n3097 gnd.n2421 240.244
R5295 gnd.n3097 gnd.n2414 240.244
R5296 gnd.n3108 gnd.n2414 240.244
R5297 gnd.n3108 gnd.n2407 240.244
R5298 gnd.n3123 gnd.n2407 240.244
R5299 gnd.n3123 gnd.n2408 240.244
R5300 gnd.n2408 gnd.n2386 240.244
R5301 gnd.n3145 gnd.n2386 240.244
R5302 gnd.n3145 gnd.n2387 240.244
R5303 gnd.n2387 gnd.n2366 240.244
R5304 gnd.n3182 gnd.n2366 240.244
R5305 gnd.n3182 gnd.n2359 240.244
R5306 gnd.n3193 gnd.n2359 240.244
R5307 gnd.n3193 gnd.n2352 240.244
R5308 gnd.n3208 gnd.n2352 240.244
R5309 gnd.n3208 gnd.n2353 240.244
R5310 gnd.n2353 gnd.n2330 240.244
R5311 gnd.n3230 gnd.n2330 240.244
R5312 gnd.n3230 gnd.n2332 240.244
R5313 gnd.n2332 gnd.n2312 240.244
R5314 gnd.n3271 gnd.n2312 240.244
R5315 gnd.n3271 gnd.n2305 240.244
R5316 gnd.n3282 gnd.n2305 240.244
R5317 gnd.n3282 gnd.n2298 240.244
R5318 gnd.n3551 gnd.n2298 240.244
R5319 gnd.n3551 gnd.n2299 240.244
R5320 gnd.n2299 gnd.n2280 240.244
R5321 gnd.n3574 gnd.n2280 240.244
R5322 gnd.n910 gnd.n863 240.244
R5323 gnd.n967 gnd.n911 240.244
R5324 gnd.n921 gnd.n920 240.244
R5325 gnd.n969 gnd.n928 240.244
R5326 gnd.n972 gnd.n929 240.244
R5327 gnd.n939 gnd.n938 240.244
R5328 gnd.n974 gnd.n946 240.244
R5329 gnd.n977 gnd.n947 240.244
R5330 gnd.n964 gnd.n959 240.244
R5331 gnd.n3743 gnd.n3669 240.244
R5332 gnd.n3743 gnd.n2195 240.244
R5333 gnd.n2195 gnd.n2184 240.244
R5334 gnd.n3990 gnd.n2184 240.244
R5335 gnd.n3990 gnd.n2180 240.244
R5336 gnd.n3998 gnd.n2180 240.244
R5337 gnd.n3998 gnd.n2170 240.244
R5338 gnd.n2170 gnd.n2159 240.244
R5339 gnd.n4025 gnd.n2159 240.244
R5340 gnd.n4025 gnd.n2155 240.244
R5341 gnd.n4035 gnd.n2155 240.244
R5342 gnd.n4035 gnd.n2143 240.244
R5343 gnd.n2143 gnd.n2133 240.244
R5344 gnd.n4064 gnd.n2133 240.244
R5345 gnd.n4065 gnd.n4064 240.244
R5346 gnd.n4065 gnd.n735 240.244
R5347 gnd.n4071 gnd.n735 240.244
R5348 gnd.n4071 gnd.n746 240.244
R5349 gnd.n4091 gnd.n746 240.244
R5350 gnd.n4091 gnd.n757 240.244
R5351 gnd.n4097 gnd.n757 240.244
R5352 gnd.n4097 gnd.n765 240.244
R5353 gnd.n4116 gnd.n765 240.244
R5354 gnd.n4116 gnd.n774 240.244
R5355 gnd.n4110 gnd.n774 240.244
R5356 gnd.n4110 gnd.n782 240.244
R5357 gnd.n4154 gnd.n782 240.244
R5358 gnd.n4154 gnd.n791 240.244
R5359 gnd.n4160 gnd.n791 240.244
R5360 gnd.n4160 gnd.n802 240.244
R5361 gnd.n4168 gnd.n802 240.244
R5362 gnd.n4168 gnd.n811 240.244
R5363 gnd.n4174 gnd.n811 240.244
R5364 gnd.n4174 gnd.n822 240.244
R5365 gnd.n4198 gnd.n822 240.244
R5366 gnd.n4198 gnd.n831 240.244
R5367 gnd.n2100 gnd.n831 240.244
R5368 gnd.n2100 gnd.n842 240.244
R5369 gnd.n4189 gnd.n842 240.244
R5370 gnd.n4189 gnd.n852 240.244
R5371 gnd.n5877 gnd.n852 240.244
R5372 gnd.n5877 gnd.n861 240.244
R5373 gnd.n3696 gnd.n3694 240.244
R5374 gnd.n3702 gnd.n3687 240.244
R5375 gnd.n3706 gnd.n3704 240.244
R5376 gnd.n3712 gnd.n3683 240.244
R5377 gnd.n3716 gnd.n3714 240.244
R5378 gnd.n3722 gnd.n3679 240.244
R5379 gnd.n3726 gnd.n3724 240.244
R5380 gnd.n3732 gnd.n3675 240.244
R5381 gnd.n3735 gnd.n3734 240.244
R5382 gnd.n3962 gnd.n2196 240.244
R5383 gnd.n3978 gnd.n2196 240.244
R5384 gnd.n3978 gnd.n2197 240.244
R5385 gnd.n2197 gnd.n2187 240.244
R5386 gnd.n3973 gnd.n2187 240.244
R5387 gnd.n3973 gnd.n2171 240.244
R5388 gnd.n4013 gnd.n2171 240.244
R5389 gnd.n4013 gnd.n2172 240.244
R5390 gnd.n2172 gnd.n2162 240.244
R5391 gnd.n4008 gnd.n2162 240.244
R5392 gnd.n4008 gnd.n2145 240.244
R5393 gnd.n4053 gnd.n2145 240.244
R5394 gnd.n4053 gnd.n2146 240.244
R5395 gnd.n2146 gnd.n2136 240.244
R5396 gnd.n4048 gnd.n2136 240.244
R5397 gnd.n4048 gnd.n737 240.244
R5398 gnd.n748 gnd.n737 240.244
R5399 gnd.n5958 gnd.n748 240.244
R5400 gnd.n5958 gnd.n749 240.244
R5401 gnd.n5954 gnd.n749 240.244
R5402 gnd.n5954 gnd.n755 240.244
R5403 gnd.n5945 gnd.n755 240.244
R5404 gnd.n5945 gnd.n766 240.244
R5405 gnd.n5941 gnd.n766 240.244
R5406 gnd.n5941 gnd.n771 240.244
R5407 gnd.n5932 gnd.n771 240.244
R5408 gnd.n5932 gnd.n784 240.244
R5409 gnd.n5928 gnd.n784 240.244
R5410 gnd.n5928 gnd.n789 240.244
R5411 gnd.n5920 gnd.n789 240.244
R5412 gnd.n5920 gnd.n803 240.244
R5413 gnd.n5916 gnd.n803 240.244
R5414 gnd.n5916 gnd.n808 240.244
R5415 gnd.n5908 gnd.n808 240.244
R5416 gnd.n5908 gnd.n824 240.244
R5417 gnd.n5904 gnd.n824 240.244
R5418 gnd.n5904 gnd.n829 240.244
R5419 gnd.n5896 gnd.n829 240.244
R5420 gnd.n5896 gnd.n844 240.244
R5421 gnd.n5892 gnd.n844 240.244
R5422 gnd.n5892 gnd.n849 240.244
R5423 gnd.n5884 gnd.n849 240.244
R5424 gnd.n6144 gnd.n560 240.244
R5425 gnd.n6148 gnd.n560 240.244
R5426 gnd.n6148 gnd.n556 240.244
R5427 gnd.n6154 gnd.n556 240.244
R5428 gnd.n6154 gnd.n554 240.244
R5429 gnd.n6158 gnd.n554 240.244
R5430 gnd.n6158 gnd.n550 240.244
R5431 gnd.n6164 gnd.n550 240.244
R5432 gnd.n6164 gnd.n548 240.244
R5433 gnd.n6168 gnd.n548 240.244
R5434 gnd.n6168 gnd.n544 240.244
R5435 gnd.n6174 gnd.n544 240.244
R5436 gnd.n6174 gnd.n542 240.244
R5437 gnd.n6178 gnd.n542 240.244
R5438 gnd.n6178 gnd.n538 240.244
R5439 gnd.n6184 gnd.n538 240.244
R5440 gnd.n6184 gnd.n536 240.244
R5441 gnd.n6188 gnd.n536 240.244
R5442 gnd.n6188 gnd.n532 240.244
R5443 gnd.n6194 gnd.n532 240.244
R5444 gnd.n6194 gnd.n530 240.244
R5445 gnd.n6198 gnd.n530 240.244
R5446 gnd.n6198 gnd.n526 240.244
R5447 gnd.n6204 gnd.n526 240.244
R5448 gnd.n6204 gnd.n524 240.244
R5449 gnd.n6208 gnd.n524 240.244
R5450 gnd.n6208 gnd.n520 240.244
R5451 gnd.n6214 gnd.n520 240.244
R5452 gnd.n6214 gnd.n518 240.244
R5453 gnd.n6218 gnd.n518 240.244
R5454 gnd.n6218 gnd.n514 240.244
R5455 gnd.n6224 gnd.n514 240.244
R5456 gnd.n6224 gnd.n512 240.244
R5457 gnd.n6228 gnd.n512 240.244
R5458 gnd.n6228 gnd.n508 240.244
R5459 gnd.n6234 gnd.n508 240.244
R5460 gnd.n6234 gnd.n506 240.244
R5461 gnd.n6238 gnd.n506 240.244
R5462 gnd.n6238 gnd.n502 240.244
R5463 gnd.n6244 gnd.n502 240.244
R5464 gnd.n6244 gnd.n500 240.244
R5465 gnd.n6248 gnd.n500 240.244
R5466 gnd.n6248 gnd.n496 240.244
R5467 gnd.n6254 gnd.n496 240.244
R5468 gnd.n6254 gnd.n494 240.244
R5469 gnd.n6258 gnd.n494 240.244
R5470 gnd.n6258 gnd.n490 240.244
R5471 gnd.n6264 gnd.n490 240.244
R5472 gnd.n6264 gnd.n488 240.244
R5473 gnd.n6268 gnd.n488 240.244
R5474 gnd.n6268 gnd.n484 240.244
R5475 gnd.n6274 gnd.n484 240.244
R5476 gnd.n6274 gnd.n482 240.244
R5477 gnd.n6278 gnd.n482 240.244
R5478 gnd.n6278 gnd.n478 240.244
R5479 gnd.n6284 gnd.n478 240.244
R5480 gnd.n6284 gnd.n476 240.244
R5481 gnd.n6288 gnd.n476 240.244
R5482 gnd.n6288 gnd.n472 240.244
R5483 gnd.n6294 gnd.n472 240.244
R5484 gnd.n6294 gnd.n470 240.244
R5485 gnd.n6298 gnd.n470 240.244
R5486 gnd.n6298 gnd.n466 240.244
R5487 gnd.n6304 gnd.n466 240.244
R5488 gnd.n6304 gnd.n464 240.244
R5489 gnd.n6308 gnd.n464 240.244
R5490 gnd.n6308 gnd.n460 240.244
R5491 gnd.n6314 gnd.n460 240.244
R5492 gnd.n6314 gnd.n458 240.244
R5493 gnd.n6318 gnd.n458 240.244
R5494 gnd.n6318 gnd.n454 240.244
R5495 gnd.n6324 gnd.n454 240.244
R5496 gnd.n6324 gnd.n452 240.244
R5497 gnd.n6328 gnd.n452 240.244
R5498 gnd.n6328 gnd.n448 240.244
R5499 gnd.n6334 gnd.n448 240.244
R5500 gnd.n6334 gnd.n446 240.244
R5501 gnd.n6338 gnd.n446 240.244
R5502 gnd.n6338 gnd.n442 240.244
R5503 gnd.n6344 gnd.n442 240.244
R5504 gnd.n6344 gnd.n440 240.244
R5505 gnd.n6348 gnd.n440 240.244
R5506 gnd.n6348 gnd.n436 240.244
R5507 gnd.n6354 gnd.n436 240.244
R5508 gnd.n6354 gnd.n434 240.244
R5509 gnd.n6358 gnd.n434 240.244
R5510 gnd.n6358 gnd.n430 240.244
R5511 gnd.n6364 gnd.n430 240.244
R5512 gnd.n6364 gnd.n428 240.244
R5513 gnd.n6368 gnd.n428 240.244
R5514 gnd.n6368 gnd.n424 240.244
R5515 gnd.n6374 gnd.n424 240.244
R5516 gnd.n6374 gnd.n422 240.244
R5517 gnd.n6378 gnd.n422 240.244
R5518 gnd.n6378 gnd.n418 240.244
R5519 gnd.n6384 gnd.n418 240.244
R5520 gnd.n6384 gnd.n416 240.244
R5521 gnd.n6388 gnd.n416 240.244
R5522 gnd.n6388 gnd.n412 240.244
R5523 gnd.n6394 gnd.n412 240.244
R5524 gnd.n6394 gnd.n410 240.244
R5525 gnd.n6398 gnd.n410 240.244
R5526 gnd.n6398 gnd.n406 240.244
R5527 gnd.n6404 gnd.n406 240.244
R5528 gnd.n6404 gnd.n404 240.244
R5529 gnd.n6408 gnd.n404 240.244
R5530 gnd.n6408 gnd.n400 240.244
R5531 gnd.n6414 gnd.n400 240.244
R5532 gnd.n6414 gnd.n398 240.244
R5533 gnd.n6418 gnd.n398 240.244
R5534 gnd.n6418 gnd.n394 240.244
R5535 gnd.n6424 gnd.n394 240.244
R5536 gnd.n6424 gnd.n392 240.244
R5537 gnd.n6428 gnd.n392 240.244
R5538 gnd.n6428 gnd.n388 240.244
R5539 gnd.n6434 gnd.n388 240.244
R5540 gnd.n6434 gnd.n386 240.244
R5541 gnd.n6438 gnd.n386 240.244
R5542 gnd.n6438 gnd.n382 240.244
R5543 gnd.n6444 gnd.n382 240.244
R5544 gnd.n6444 gnd.n380 240.244
R5545 gnd.n6448 gnd.n380 240.244
R5546 gnd.n6448 gnd.n376 240.244
R5547 gnd.n6454 gnd.n376 240.244
R5548 gnd.n6454 gnd.n374 240.244
R5549 gnd.n6458 gnd.n374 240.244
R5550 gnd.n6458 gnd.n370 240.244
R5551 gnd.n6464 gnd.n370 240.244
R5552 gnd.n6464 gnd.n368 240.244
R5553 gnd.n6468 gnd.n368 240.244
R5554 gnd.n6468 gnd.n364 240.244
R5555 gnd.n6474 gnd.n364 240.244
R5556 gnd.n6474 gnd.n362 240.244
R5557 gnd.n6478 gnd.n362 240.244
R5558 gnd.n6478 gnd.n358 240.244
R5559 gnd.n6484 gnd.n358 240.244
R5560 gnd.n6484 gnd.n356 240.244
R5561 gnd.n6488 gnd.n356 240.244
R5562 gnd.n6488 gnd.n352 240.244
R5563 gnd.n6494 gnd.n352 240.244
R5564 gnd.n6494 gnd.n350 240.244
R5565 gnd.n6498 gnd.n350 240.244
R5566 gnd.n6498 gnd.n346 240.244
R5567 gnd.n6504 gnd.n346 240.244
R5568 gnd.n6504 gnd.n344 240.244
R5569 gnd.n6508 gnd.n344 240.244
R5570 gnd.n6508 gnd.n340 240.244
R5571 gnd.n6514 gnd.n340 240.244
R5572 gnd.n6514 gnd.n338 240.244
R5573 gnd.n6518 gnd.n338 240.244
R5574 gnd.n6518 gnd.n334 240.244
R5575 gnd.n6524 gnd.n334 240.244
R5576 gnd.n6524 gnd.n332 240.244
R5577 gnd.n6528 gnd.n332 240.244
R5578 gnd.n6528 gnd.n328 240.244
R5579 gnd.n6534 gnd.n328 240.244
R5580 gnd.n6534 gnd.n326 240.244
R5581 gnd.n6538 gnd.n326 240.244
R5582 gnd.n6538 gnd.n322 240.244
R5583 gnd.n6544 gnd.n322 240.244
R5584 gnd.n6544 gnd.n320 240.244
R5585 gnd.n6548 gnd.n320 240.244
R5586 gnd.n6548 gnd.n316 240.244
R5587 gnd.n6555 gnd.n316 240.244
R5588 gnd.n6555 gnd.n314 240.244
R5589 gnd.n6559 gnd.n314 240.244
R5590 gnd.n6559 gnd.n311 240.244
R5591 gnd.n6565 gnd.n309 240.244
R5592 gnd.n6569 gnd.n309 240.244
R5593 gnd.n6569 gnd.n305 240.244
R5594 gnd.n6575 gnd.n305 240.244
R5595 gnd.n6575 gnd.n303 240.244
R5596 gnd.n6579 gnd.n303 240.244
R5597 gnd.n6579 gnd.n299 240.244
R5598 gnd.n6585 gnd.n299 240.244
R5599 gnd.n6585 gnd.n297 240.244
R5600 gnd.n6589 gnd.n297 240.244
R5601 gnd.n6589 gnd.n293 240.244
R5602 gnd.n6595 gnd.n293 240.244
R5603 gnd.n6595 gnd.n291 240.244
R5604 gnd.n6599 gnd.n291 240.244
R5605 gnd.n6599 gnd.n287 240.244
R5606 gnd.n6605 gnd.n287 240.244
R5607 gnd.n6605 gnd.n285 240.244
R5608 gnd.n6609 gnd.n285 240.244
R5609 gnd.n6609 gnd.n281 240.244
R5610 gnd.n6615 gnd.n281 240.244
R5611 gnd.n6615 gnd.n279 240.244
R5612 gnd.n6619 gnd.n279 240.244
R5613 gnd.n6619 gnd.n275 240.244
R5614 gnd.n6625 gnd.n275 240.244
R5615 gnd.n6625 gnd.n273 240.244
R5616 gnd.n6629 gnd.n273 240.244
R5617 gnd.n6629 gnd.n269 240.244
R5618 gnd.n6635 gnd.n269 240.244
R5619 gnd.n6635 gnd.n267 240.244
R5620 gnd.n6639 gnd.n267 240.244
R5621 gnd.n6639 gnd.n263 240.244
R5622 gnd.n6645 gnd.n263 240.244
R5623 gnd.n6645 gnd.n261 240.244
R5624 gnd.n6649 gnd.n261 240.244
R5625 gnd.n6649 gnd.n257 240.244
R5626 gnd.n6655 gnd.n257 240.244
R5627 gnd.n6655 gnd.n255 240.244
R5628 gnd.n6659 gnd.n255 240.244
R5629 gnd.n6659 gnd.n251 240.244
R5630 gnd.n6665 gnd.n251 240.244
R5631 gnd.n6665 gnd.n249 240.244
R5632 gnd.n6669 gnd.n249 240.244
R5633 gnd.n6669 gnd.n245 240.244
R5634 gnd.n6675 gnd.n245 240.244
R5635 gnd.n6675 gnd.n243 240.244
R5636 gnd.n6679 gnd.n243 240.244
R5637 gnd.n6679 gnd.n239 240.244
R5638 gnd.n6685 gnd.n239 240.244
R5639 gnd.n6685 gnd.n237 240.244
R5640 gnd.n6689 gnd.n237 240.244
R5641 gnd.n6689 gnd.n233 240.244
R5642 gnd.n6695 gnd.n233 240.244
R5643 gnd.n6695 gnd.n231 240.244
R5644 gnd.n6699 gnd.n231 240.244
R5645 gnd.n6699 gnd.n227 240.244
R5646 gnd.n6705 gnd.n227 240.244
R5647 gnd.n6705 gnd.n225 240.244
R5648 gnd.n6709 gnd.n225 240.244
R5649 gnd.n6709 gnd.n221 240.244
R5650 gnd.n6715 gnd.n221 240.244
R5651 gnd.n6715 gnd.n219 240.244
R5652 gnd.n6719 gnd.n219 240.244
R5653 gnd.n6719 gnd.n215 240.244
R5654 gnd.n6725 gnd.n215 240.244
R5655 gnd.n6725 gnd.n213 240.244
R5656 gnd.n6729 gnd.n213 240.244
R5657 gnd.n6729 gnd.n209 240.244
R5658 gnd.n6735 gnd.n209 240.244
R5659 gnd.n6735 gnd.n207 240.244
R5660 gnd.n6739 gnd.n207 240.244
R5661 gnd.n6739 gnd.n203 240.244
R5662 gnd.n6745 gnd.n203 240.244
R5663 gnd.n6745 gnd.n201 240.244
R5664 gnd.n6749 gnd.n201 240.244
R5665 gnd.n6749 gnd.n197 240.244
R5666 gnd.n6755 gnd.n197 240.244
R5667 gnd.n6755 gnd.n195 240.244
R5668 gnd.n6759 gnd.n195 240.244
R5669 gnd.n6759 gnd.n191 240.244
R5670 gnd.n6765 gnd.n191 240.244
R5671 gnd.n6765 gnd.n189 240.244
R5672 gnd.n6770 gnd.n189 240.244
R5673 gnd.n6770 gnd.n185 240.244
R5674 gnd.n6776 gnd.n185 240.244
R5675 gnd.n5968 gnd.n732 240.244
R5676 gnd.n4081 gnd.n732 240.244
R5677 gnd.n4081 gnd.n4078 240.244
R5678 gnd.n4088 gnd.n4078 240.244
R5679 gnd.n4088 gnd.n4079 240.244
R5680 gnd.n4079 gnd.n2118 240.244
R5681 gnd.n4119 gnd.n2118 240.244
R5682 gnd.n4119 gnd.n2116 240.244
R5683 gnd.n4124 gnd.n2116 240.244
R5684 gnd.n4125 gnd.n4124 240.244
R5685 gnd.n4125 gnd.n2113 240.244
R5686 gnd.n4151 gnd.n2113 240.244
R5687 gnd.n4151 gnd.n2114 240.244
R5688 gnd.n4147 gnd.n2114 240.244
R5689 gnd.n4147 gnd.n4146 240.244
R5690 gnd.n4146 gnd.n4145 240.244
R5691 gnd.n4145 gnd.n4133 240.244
R5692 gnd.n4141 gnd.n4133 240.244
R5693 gnd.n4141 gnd.n2093 240.244
R5694 gnd.n4201 gnd.n2093 240.244
R5695 gnd.n4202 gnd.n4201 240.244
R5696 gnd.n4203 gnd.n4202 240.244
R5697 gnd.n4203 gnd.n2089 240.244
R5698 gnd.n4209 gnd.n2089 240.244
R5699 gnd.n4210 gnd.n4209 240.244
R5700 gnd.n4211 gnd.n4210 240.244
R5701 gnd.n4211 gnd.n2085 240.244
R5702 gnd.n4217 gnd.n2085 240.244
R5703 gnd.n4218 gnd.n4217 240.244
R5704 gnd.n4220 gnd.n4218 240.244
R5705 gnd.n4220 gnd.n2081 240.244
R5706 gnd.n4226 gnd.n2081 240.244
R5707 gnd.n4227 gnd.n4226 240.244
R5708 gnd.n4305 gnd.n4227 240.244
R5709 gnd.n4305 gnd.n2077 240.244
R5710 gnd.n4311 gnd.n2077 240.244
R5711 gnd.n4311 gnd.n2066 240.244
R5712 gnd.n4321 gnd.n2066 240.244
R5713 gnd.n4321 gnd.n2062 240.244
R5714 gnd.n4327 gnd.n2062 240.244
R5715 gnd.n4327 gnd.n2053 240.244
R5716 gnd.n4337 gnd.n2053 240.244
R5717 gnd.n4337 gnd.n2049 240.244
R5718 gnd.n4343 gnd.n2049 240.244
R5719 gnd.n4343 gnd.n2039 240.244
R5720 gnd.n4353 gnd.n2039 240.244
R5721 gnd.n4353 gnd.n2035 240.244
R5722 gnd.n4359 gnd.n2035 240.244
R5723 gnd.n4359 gnd.n2025 240.244
R5724 gnd.n4369 gnd.n2025 240.244
R5725 gnd.n4369 gnd.n2021 240.244
R5726 gnd.n4375 gnd.n2021 240.244
R5727 gnd.n4375 gnd.n2011 240.244
R5728 gnd.n4385 gnd.n2011 240.244
R5729 gnd.n4385 gnd.n2007 240.244
R5730 gnd.n4391 gnd.n2007 240.244
R5731 gnd.n4391 gnd.n1996 240.244
R5732 gnd.n4402 gnd.n1996 240.244
R5733 gnd.n4402 gnd.n1991 240.244
R5734 gnd.n4414 gnd.n1991 240.244
R5735 gnd.n4414 gnd.n1992 240.244
R5736 gnd.n4410 gnd.n1992 240.244
R5737 gnd.n4410 gnd.n1205 240.244
R5738 gnd.n5676 gnd.n1205 240.244
R5739 gnd.n5676 gnd.n1206 240.244
R5740 gnd.n5672 gnd.n1206 240.244
R5741 gnd.n5672 gnd.n1212 240.244
R5742 gnd.n1967 gnd.n1212 240.244
R5743 gnd.n4560 gnd.n1967 240.244
R5744 gnd.n4560 gnd.n1962 240.244
R5745 gnd.n4566 gnd.n1962 240.244
R5746 gnd.n4566 gnd.n1939 240.244
R5747 gnd.n4603 gnd.n1939 240.244
R5748 gnd.n4603 gnd.n1934 240.244
R5749 gnd.n4611 gnd.n1934 240.244
R5750 gnd.n4611 gnd.n1935 240.244
R5751 gnd.n1935 gnd.n1918 240.244
R5752 gnd.n4663 gnd.n1918 240.244
R5753 gnd.n4663 gnd.n1913 240.244
R5754 gnd.n4680 gnd.n1913 240.244
R5755 gnd.n4680 gnd.n1914 240.244
R5756 gnd.n4676 gnd.n1914 240.244
R5757 gnd.n4676 gnd.n4675 240.244
R5758 gnd.n4675 gnd.n4674 240.244
R5759 gnd.n4674 gnd.n1881 240.244
R5760 gnd.n4724 gnd.n1881 240.244
R5761 gnd.n4724 gnd.n1877 240.244
R5762 gnd.n4730 gnd.n1877 240.244
R5763 gnd.n4730 gnd.n1858 240.244
R5764 gnd.n4770 gnd.n1858 240.244
R5765 gnd.n4770 gnd.n1853 240.244
R5766 gnd.n4778 gnd.n1853 240.244
R5767 gnd.n4778 gnd.n1854 240.244
R5768 gnd.n1854 gnd.n1837 240.244
R5769 gnd.n4822 gnd.n1837 240.244
R5770 gnd.n4822 gnd.n1832 240.244
R5771 gnd.n4830 gnd.n1832 240.244
R5772 gnd.n4830 gnd.n1833 240.244
R5773 gnd.n1833 gnd.n1810 240.244
R5774 gnd.n4858 gnd.n1810 240.244
R5775 gnd.n4858 gnd.n1806 240.244
R5776 gnd.n4864 gnd.n1806 240.244
R5777 gnd.n4864 gnd.n1754 240.244
R5778 gnd.n5033 gnd.n1754 240.244
R5779 gnd.n5033 gnd.n1750 240.244
R5780 gnd.n5039 gnd.n1750 240.244
R5781 gnd.n5039 gnd.n1742 240.244
R5782 gnd.n5049 gnd.n1742 240.244
R5783 gnd.n5049 gnd.n1738 240.244
R5784 gnd.n5055 gnd.n1738 240.244
R5785 gnd.n5055 gnd.n1729 240.244
R5786 gnd.n5066 gnd.n1729 240.244
R5787 gnd.n5066 gnd.n1725 240.244
R5788 gnd.n5072 gnd.n1725 240.244
R5789 gnd.n5072 gnd.n1717 240.244
R5790 gnd.n5082 gnd.n1717 240.244
R5791 gnd.n5082 gnd.n1713 240.244
R5792 gnd.n5088 gnd.n1713 240.244
R5793 gnd.n5088 gnd.n1704 240.244
R5794 gnd.n5098 gnd.n1704 240.244
R5795 gnd.n5098 gnd.n1700 240.244
R5796 gnd.n5104 gnd.n1700 240.244
R5797 gnd.n5104 gnd.n1691 240.244
R5798 gnd.n5114 gnd.n1691 240.244
R5799 gnd.n5114 gnd.n1687 240.244
R5800 gnd.n5120 gnd.n1687 240.244
R5801 gnd.n5120 gnd.n1678 240.244
R5802 gnd.n5130 gnd.n1678 240.244
R5803 gnd.n5130 gnd.n1674 240.244
R5804 gnd.n5139 gnd.n1674 240.244
R5805 gnd.n5139 gnd.n1665 240.244
R5806 gnd.n5149 gnd.n1665 240.244
R5807 gnd.n5150 gnd.n5149 240.244
R5808 gnd.n5150 gnd.n1306 240.244
R5809 gnd.n1660 gnd.n1306 240.244
R5810 gnd.n5168 gnd.n1660 240.244
R5811 gnd.n5168 gnd.n1661 240.244
R5812 gnd.n5164 gnd.n1661 240.244
R5813 gnd.n5164 gnd.n5163 240.244
R5814 gnd.n5163 gnd.n5162 240.244
R5815 gnd.n5162 gnd.n1629 240.244
R5816 gnd.n5220 gnd.n1629 240.244
R5817 gnd.n5220 gnd.n1625 240.244
R5818 gnd.n5226 gnd.n1625 240.244
R5819 gnd.n5227 gnd.n5226 240.244
R5820 gnd.n5228 gnd.n5227 240.244
R5821 gnd.n5228 gnd.n1621 240.244
R5822 gnd.n5234 gnd.n1621 240.244
R5823 gnd.n5235 gnd.n5234 240.244
R5824 gnd.n5236 gnd.n5235 240.244
R5825 gnd.n5236 gnd.n1616 240.244
R5826 gnd.n5259 gnd.n1616 240.244
R5827 gnd.n5259 gnd.n1617 240.244
R5828 gnd.n5255 gnd.n1617 240.244
R5829 gnd.n5255 gnd.n5254 240.244
R5830 gnd.n5254 gnd.n5253 240.244
R5831 gnd.n5253 gnd.n5244 240.244
R5832 gnd.n5248 gnd.n5244 240.244
R5833 gnd.n5248 gnd.n1587 240.244
R5834 gnd.n5313 gnd.n1587 240.244
R5835 gnd.n5313 gnd.n1588 240.244
R5836 gnd.n5308 gnd.n1588 240.244
R5837 gnd.n5308 gnd.n1592 240.244
R5838 gnd.n1592 gnd.n181 240.244
R5839 gnd.n6782 gnd.n181 240.244
R5840 gnd.n6782 gnd.n182 240.244
R5841 gnd.n6777 gnd.n182 240.244
R5842 gnd.n6138 gnd.n562 240.244
R5843 gnd.n6138 gnd.n565 240.244
R5844 gnd.n6134 gnd.n565 240.244
R5845 gnd.n6134 gnd.n567 240.244
R5846 gnd.n6130 gnd.n567 240.244
R5847 gnd.n6130 gnd.n573 240.244
R5848 gnd.n6126 gnd.n573 240.244
R5849 gnd.n6126 gnd.n575 240.244
R5850 gnd.n6122 gnd.n575 240.244
R5851 gnd.n6122 gnd.n581 240.244
R5852 gnd.n6118 gnd.n581 240.244
R5853 gnd.n6118 gnd.n583 240.244
R5854 gnd.n6114 gnd.n583 240.244
R5855 gnd.n6114 gnd.n589 240.244
R5856 gnd.n6110 gnd.n589 240.244
R5857 gnd.n6110 gnd.n591 240.244
R5858 gnd.n6106 gnd.n591 240.244
R5859 gnd.n6106 gnd.n597 240.244
R5860 gnd.n6102 gnd.n597 240.244
R5861 gnd.n6102 gnd.n599 240.244
R5862 gnd.n6098 gnd.n599 240.244
R5863 gnd.n6098 gnd.n605 240.244
R5864 gnd.n6094 gnd.n605 240.244
R5865 gnd.n6094 gnd.n607 240.244
R5866 gnd.n6090 gnd.n607 240.244
R5867 gnd.n6090 gnd.n613 240.244
R5868 gnd.n6086 gnd.n613 240.244
R5869 gnd.n6086 gnd.n615 240.244
R5870 gnd.n6082 gnd.n615 240.244
R5871 gnd.n6082 gnd.n621 240.244
R5872 gnd.n6078 gnd.n621 240.244
R5873 gnd.n6078 gnd.n623 240.244
R5874 gnd.n6074 gnd.n623 240.244
R5875 gnd.n6074 gnd.n629 240.244
R5876 gnd.n6070 gnd.n629 240.244
R5877 gnd.n6070 gnd.n631 240.244
R5878 gnd.n6066 gnd.n631 240.244
R5879 gnd.n6066 gnd.n637 240.244
R5880 gnd.n6062 gnd.n637 240.244
R5881 gnd.n6062 gnd.n639 240.244
R5882 gnd.n6058 gnd.n639 240.244
R5883 gnd.n6058 gnd.n645 240.244
R5884 gnd.n6054 gnd.n645 240.244
R5885 gnd.n6054 gnd.n647 240.244
R5886 gnd.n6050 gnd.n647 240.244
R5887 gnd.n6050 gnd.n653 240.244
R5888 gnd.n6046 gnd.n653 240.244
R5889 gnd.n6046 gnd.n655 240.244
R5890 gnd.n6042 gnd.n655 240.244
R5891 gnd.n6042 gnd.n661 240.244
R5892 gnd.n6038 gnd.n661 240.244
R5893 gnd.n6038 gnd.n663 240.244
R5894 gnd.n6034 gnd.n663 240.244
R5895 gnd.n6034 gnd.n669 240.244
R5896 gnd.n6030 gnd.n669 240.244
R5897 gnd.n6030 gnd.n671 240.244
R5898 gnd.n6026 gnd.n671 240.244
R5899 gnd.n6026 gnd.n677 240.244
R5900 gnd.n6022 gnd.n677 240.244
R5901 gnd.n6022 gnd.n679 240.244
R5902 gnd.n6018 gnd.n679 240.244
R5903 gnd.n6018 gnd.n685 240.244
R5904 gnd.n6014 gnd.n685 240.244
R5905 gnd.n6014 gnd.n687 240.244
R5906 gnd.n6010 gnd.n687 240.244
R5907 gnd.n6010 gnd.n693 240.244
R5908 gnd.n6006 gnd.n693 240.244
R5909 gnd.n6006 gnd.n695 240.244
R5910 gnd.n6002 gnd.n695 240.244
R5911 gnd.n6002 gnd.n701 240.244
R5912 gnd.n5998 gnd.n701 240.244
R5913 gnd.n5998 gnd.n703 240.244
R5914 gnd.n5994 gnd.n703 240.244
R5915 gnd.n5994 gnd.n709 240.244
R5916 gnd.n5990 gnd.n709 240.244
R5917 gnd.n5990 gnd.n711 240.244
R5918 gnd.n5986 gnd.n711 240.244
R5919 gnd.n5986 gnd.n717 240.244
R5920 gnd.n5982 gnd.n717 240.244
R5921 gnd.n5982 gnd.n719 240.244
R5922 gnd.n5978 gnd.n719 240.244
R5923 gnd.n5978 gnd.n725 240.244
R5924 gnd.n5974 gnd.n725 240.244
R5925 gnd.n5974 gnd.n727 240.244
R5926 gnd.n4298 gnd.n893 240.244
R5927 gnd.n4298 gnd.n4229 240.244
R5928 gnd.n4229 gnd.n2076 240.244
R5929 gnd.n4234 gnd.n2076 240.244
R5930 gnd.n4234 gnd.n2068 240.244
R5931 gnd.n4235 gnd.n2068 240.244
R5932 gnd.n4235 gnd.n2061 240.244
R5933 gnd.n4238 gnd.n2061 240.244
R5934 gnd.n4238 gnd.n2055 240.244
R5935 gnd.n4239 gnd.n2055 240.244
R5936 gnd.n4239 gnd.n2048 240.244
R5937 gnd.n4242 gnd.n2048 240.244
R5938 gnd.n4242 gnd.n2041 240.244
R5939 gnd.n4243 gnd.n2041 240.244
R5940 gnd.n4243 gnd.n2034 240.244
R5941 gnd.n4246 gnd.n2034 240.244
R5942 gnd.n4246 gnd.n2027 240.244
R5943 gnd.n4247 gnd.n2027 240.244
R5944 gnd.n4247 gnd.n2019 240.244
R5945 gnd.n4250 gnd.n2019 240.244
R5946 gnd.n4250 gnd.n2012 240.244
R5947 gnd.n4251 gnd.n2012 240.244
R5948 gnd.n4251 gnd.n2006 240.244
R5949 gnd.n4254 gnd.n2006 240.244
R5950 gnd.n4254 gnd.n1998 240.244
R5951 gnd.n4255 gnd.n1998 240.244
R5952 gnd.n4255 gnd.n1990 240.244
R5953 gnd.n1990 gnd.n1982 240.244
R5954 gnd.n4427 gnd.n1982 240.244
R5955 gnd.n4427 gnd.n4426 240.244
R5956 gnd.n4426 gnd.n1203 240.244
R5957 gnd.n4531 gnd.n1203 240.244
R5958 gnd.n4531 gnd.n1214 240.244
R5959 gnd.n1975 gnd.n1214 240.244
R5960 gnd.n4550 gnd.n1975 240.244
R5961 gnd.n4550 gnd.n1969 240.244
R5962 gnd.n4537 gnd.n1969 240.244
R5963 gnd.n4537 gnd.n1959 240.244
R5964 gnd.n4539 gnd.n1959 240.244
R5965 gnd.n4539 gnd.n1941 240.244
R5966 gnd.n1941 gnd.n1931 240.244
R5967 gnd.n4613 gnd.n1931 240.244
R5968 gnd.n4613 gnd.n1926 240.244
R5969 gnd.n4653 gnd.n1926 240.244
R5970 gnd.n4653 gnd.n1920 240.244
R5971 gnd.n4618 gnd.n1920 240.244
R5972 gnd.n4618 gnd.n1912 240.244
R5973 gnd.n4619 gnd.n1912 240.244
R5974 gnd.n4622 gnd.n4619 240.244
R5975 gnd.n4623 gnd.n4622 240.244
R5976 gnd.n4624 gnd.n4623 240.244
R5977 gnd.n4624 gnd.n1890 240.244
R5978 gnd.n1890 gnd.n1882 240.244
R5979 gnd.n4629 gnd.n1882 240.244
R5980 gnd.n4629 gnd.n1875 240.244
R5981 gnd.n4630 gnd.n1875 240.244
R5982 gnd.n4630 gnd.n1860 240.244
R5983 gnd.n1860 gnd.n1851 240.244
R5984 gnd.n4780 gnd.n1851 240.244
R5985 gnd.n4780 gnd.n1846 240.244
R5986 gnd.n4811 gnd.n1846 240.244
R5987 gnd.n4811 gnd.n1839 240.244
R5988 gnd.n4785 gnd.n1839 240.244
R5989 gnd.n4785 gnd.n1831 240.244
R5990 gnd.n4786 gnd.n1831 240.244
R5991 gnd.n4787 gnd.n4786 240.244
R5992 gnd.n4787 gnd.n1812 240.244
R5993 gnd.n4791 gnd.n1812 240.244
R5994 gnd.n4791 gnd.n1804 240.244
R5995 gnd.n4792 gnd.n1804 240.244
R5996 gnd.n4792 gnd.n1756 240.244
R5997 gnd.n1756 gnd.n1749 240.244
R5998 gnd.n5041 gnd.n1749 240.244
R5999 gnd.n5041 gnd.n1745 240.244
R6000 gnd.n5047 gnd.n1745 240.244
R6001 gnd.n5047 gnd.n1736 240.244
R6002 gnd.n5057 gnd.n1736 240.244
R6003 gnd.n5057 gnd.n1732 240.244
R6004 gnd.n5063 gnd.n1732 240.244
R6005 gnd.n5063 gnd.n1724 240.244
R6006 gnd.n5074 gnd.n1724 240.244
R6007 gnd.n5074 gnd.n1720 240.244
R6008 gnd.n5080 gnd.n1720 240.244
R6009 gnd.n5080 gnd.n1711 240.244
R6010 gnd.n5090 gnd.n1711 240.244
R6011 gnd.n5090 gnd.n1707 240.244
R6012 gnd.n5096 gnd.n1707 240.244
R6013 gnd.n5096 gnd.n1698 240.244
R6014 gnd.n5106 gnd.n1698 240.244
R6015 gnd.n5106 gnd.n1694 240.244
R6016 gnd.n5112 gnd.n1694 240.244
R6017 gnd.n5112 gnd.n1683 240.244
R6018 gnd.n5122 gnd.n1683 240.244
R6019 gnd.n5122 gnd.n1679 240.244
R6020 gnd.n5128 gnd.n1679 240.244
R6021 gnd.n5128 gnd.n1672 240.244
R6022 gnd.n5141 gnd.n1672 240.244
R6023 gnd.n5141 gnd.n1668 240.244
R6024 gnd.n5147 gnd.n1668 240.244
R6025 gnd.n5147 gnd.n1308 240.244
R6026 gnd.n5564 gnd.n1308 240.244
R6027 gnd.n892 gnd.n891 240.244
R6028 gnd.n897 gnd.n891 240.244
R6029 gnd.n899 gnd.n898 240.244
R6030 gnd.n903 gnd.n902 240.244
R6031 gnd.n905 gnd.n904 240.244
R6032 gnd.n915 gnd.n914 240.244
R6033 gnd.n917 gnd.n916 240.244
R6034 gnd.n925 gnd.n924 240.244
R6035 gnd.n933 gnd.n932 240.244
R6036 gnd.n935 gnd.n934 240.244
R6037 gnd.n943 gnd.n942 240.244
R6038 gnd.n951 gnd.n950 240.244
R6039 gnd.n956 gnd.n952 240.244
R6040 gnd.n888 gnd.n874 240.244
R6041 gnd.n4303 gnd.n875 240.244
R6042 gnd.n4303 gnd.n2074 240.244
R6043 gnd.n4313 gnd.n2074 240.244
R6044 gnd.n4313 gnd.n2070 240.244
R6045 gnd.n4319 gnd.n2070 240.244
R6046 gnd.n4319 gnd.n2060 240.244
R6047 gnd.n4329 gnd.n2060 240.244
R6048 gnd.n4329 gnd.n2056 240.244
R6049 gnd.n4335 gnd.n2056 240.244
R6050 gnd.n4335 gnd.n2046 240.244
R6051 gnd.n4345 gnd.n2046 240.244
R6052 gnd.n4345 gnd.n2042 240.244
R6053 gnd.n4351 gnd.n2042 240.244
R6054 gnd.n4351 gnd.n2032 240.244
R6055 gnd.n4361 gnd.n2032 240.244
R6056 gnd.n4361 gnd.n2028 240.244
R6057 gnd.n4367 gnd.n2028 240.244
R6058 gnd.n4367 gnd.n2017 240.244
R6059 gnd.n4377 gnd.n2017 240.244
R6060 gnd.n4377 gnd.n2013 240.244
R6061 gnd.n4383 gnd.n2013 240.244
R6062 gnd.n4383 gnd.n2004 240.244
R6063 gnd.n4393 gnd.n2004 240.244
R6064 gnd.n4393 gnd.n1999 240.244
R6065 gnd.n4400 gnd.n1999 240.244
R6066 gnd.n4400 gnd.n1988 240.244
R6067 gnd.n4416 gnd.n1988 240.244
R6068 gnd.n4417 gnd.n4416 240.244
R6069 gnd.n4417 gnd.n1983 240.244
R6070 gnd.n4424 gnd.n1983 240.244
R6071 gnd.n4424 gnd.n1204 240.244
R6072 gnd.n1215 gnd.n1204 240.244
R6073 gnd.n5670 gnd.n1215 240.244
R6074 gnd.n5670 gnd.n1216 240.244
R6075 gnd.n1221 gnd.n1216 240.244
R6076 gnd.n1222 gnd.n1221 240.244
R6077 gnd.n1223 gnd.n1222 240.244
R6078 gnd.n1961 gnd.n1223 240.244
R6079 gnd.n1961 gnd.n1226 240.244
R6080 gnd.n1227 gnd.n1226 240.244
R6081 gnd.n1228 gnd.n1227 240.244
R6082 gnd.n1933 gnd.n1228 240.244
R6083 gnd.n1933 gnd.n1231 240.244
R6084 gnd.n1232 gnd.n1231 240.244
R6085 gnd.n1233 gnd.n1232 240.244
R6086 gnd.n1909 gnd.n1233 240.244
R6087 gnd.n1909 gnd.n1236 240.244
R6088 gnd.n1237 gnd.n1236 240.244
R6089 gnd.n1238 gnd.n1237 240.244
R6090 gnd.n1893 gnd.n1238 240.244
R6091 gnd.n1893 gnd.n1241 240.244
R6092 gnd.n1242 gnd.n1241 240.244
R6093 gnd.n1243 gnd.n1242 240.244
R6094 gnd.n4627 gnd.n1243 240.244
R6095 gnd.n4627 gnd.n1246 240.244
R6096 gnd.n1247 gnd.n1246 240.244
R6097 gnd.n1248 gnd.n1247 240.244
R6098 gnd.n4743 gnd.n1248 240.244
R6099 gnd.n4743 gnd.n1251 240.244
R6100 gnd.n1252 gnd.n1251 240.244
R6101 gnd.n1253 gnd.n1252 240.244
R6102 gnd.n4820 gnd.n1253 240.244
R6103 gnd.n4820 gnd.n1256 240.244
R6104 gnd.n1257 gnd.n1256 240.244
R6105 gnd.n1258 gnd.n1257 240.244
R6106 gnd.n1817 gnd.n1258 240.244
R6107 gnd.n1817 gnd.n1261 240.244
R6108 gnd.n1262 gnd.n1261 240.244
R6109 gnd.n1263 gnd.n1262 240.244
R6110 gnd.n1796 gnd.n1263 240.244
R6111 gnd.n1796 gnd.n1266 240.244
R6112 gnd.n1267 gnd.n1266 240.244
R6113 gnd.n1268 gnd.n1267 240.244
R6114 gnd.n1743 gnd.n1268 240.244
R6115 gnd.n1743 gnd.n1271 240.244
R6116 gnd.n1272 gnd.n1271 240.244
R6117 gnd.n1273 gnd.n1272 240.244
R6118 gnd.n1730 gnd.n1273 240.244
R6119 gnd.n1730 gnd.n1276 240.244
R6120 gnd.n1277 gnd.n1276 240.244
R6121 gnd.n1278 gnd.n1277 240.244
R6122 gnd.n1718 gnd.n1278 240.244
R6123 gnd.n1718 gnd.n1281 240.244
R6124 gnd.n1282 gnd.n1281 240.244
R6125 gnd.n1283 gnd.n1282 240.244
R6126 gnd.n1705 gnd.n1283 240.244
R6127 gnd.n1705 gnd.n1286 240.244
R6128 gnd.n1287 gnd.n1286 240.244
R6129 gnd.n1288 gnd.n1287 240.244
R6130 gnd.n1692 gnd.n1288 240.244
R6131 gnd.n1692 gnd.n1291 240.244
R6132 gnd.n1292 gnd.n1291 240.244
R6133 gnd.n1293 gnd.n1292 240.244
R6134 gnd.n1685 gnd.n1293 240.244
R6135 gnd.n1685 gnd.n1296 240.244
R6136 gnd.n1297 gnd.n1296 240.244
R6137 gnd.n1298 gnd.n1297 240.244
R6138 gnd.n1666 gnd.n1298 240.244
R6139 gnd.n1666 gnd.n1301 240.244
R6140 gnd.n1302 gnd.n1301 240.244
R6141 gnd.n5566 gnd.n1302 240.244
R6142 gnd.n1314 gnd.n1313 240.244
R6143 gnd.n1638 gnd.n1317 240.244
R6144 gnd.n1319 gnd.n1318 240.244
R6145 gnd.n1641 gnd.n1323 240.244
R6146 gnd.n1644 gnd.n1324 240.244
R6147 gnd.n1333 gnd.n1332 240.244
R6148 gnd.n1646 gnd.n1340 240.244
R6149 gnd.n1649 gnd.n1341 240.244
R6150 gnd.n1349 gnd.n1348 240.244
R6151 gnd.n1651 gnd.n1356 240.244
R6152 gnd.n1654 gnd.n1357 240.244
R6153 gnd.n1365 gnd.n1364 240.244
R6154 gnd.n1657 gnd.n1365 240.244
R6155 gnd.n5172 gnd.n1636 240.244
R6156 gnd.n1185 gnd.n1184 240.132
R6157 gnd.n4881 gnd.n4880 240.132
R6158 gnd.n6146 gnd.n6145 225.874
R6159 gnd.n6147 gnd.n6146 225.874
R6160 gnd.n6147 gnd.n555 225.874
R6161 gnd.n6155 gnd.n555 225.874
R6162 gnd.n6156 gnd.n6155 225.874
R6163 gnd.n6157 gnd.n6156 225.874
R6164 gnd.n6157 gnd.n549 225.874
R6165 gnd.n6165 gnd.n549 225.874
R6166 gnd.n6166 gnd.n6165 225.874
R6167 gnd.n6167 gnd.n6166 225.874
R6168 gnd.n6167 gnd.n543 225.874
R6169 gnd.n6175 gnd.n543 225.874
R6170 gnd.n6176 gnd.n6175 225.874
R6171 gnd.n6177 gnd.n6176 225.874
R6172 gnd.n6177 gnd.n537 225.874
R6173 gnd.n6185 gnd.n537 225.874
R6174 gnd.n6186 gnd.n6185 225.874
R6175 gnd.n6187 gnd.n6186 225.874
R6176 gnd.n6187 gnd.n531 225.874
R6177 gnd.n6195 gnd.n531 225.874
R6178 gnd.n6196 gnd.n6195 225.874
R6179 gnd.n6197 gnd.n6196 225.874
R6180 gnd.n6197 gnd.n525 225.874
R6181 gnd.n6205 gnd.n525 225.874
R6182 gnd.n6206 gnd.n6205 225.874
R6183 gnd.n6207 gnd.n6206 225.874
R6184 gnd.n6207 gnd.n519 225.874
R6185 gnd.n6215 gnd.n519 225.874
R6186 gnd.n6216 gnd.n6215 225.874
R6187 gnd.n6217 gnd.n6216 225.874
R6188 gnd.n6217 gnd.n513 225.874
R6189 gnd.n6225 gnd.n513 225.874
R6190 gnd.n6226 gnd.n6225 225.874
R6191 gnd.n6227 gnd.n6226 225.874
R6192 gnd.n6227 gnd.n507 225.874
R6193 gnd.n6235 gnd.n507 225.874
R6194 gnd.n6236 gnd.n6235 225.874
R6195 gnd.n6237 gnd.n6236 225.874
R6196 gnd.n6237 gnd.n501 225.874
R6197 gnd.n6245 gnd.n501 225.874
R6198 gnd.n6246 gnd.n6245 225.874
R6199 gnd.n6247 gnd.n6246 225.874
R6200 gnd.n6247 gnd.n495 225.874
R6201 gnd.n6255 gnd.n495 225.874
R6202 gnd.n6256 gnd.n6255 225.874
R6203 gnd.n6257 gnd.n6256 225.874
R6204 gnd.n6257 gnd.n489 225.874
R6205 gnd.n6265 gnd.n489 225.874
R6206 gnd.n6266 gnd.n6265 225.874
R6207 gnd.n6267 gnd.n6266 225.874
R6208 gnd.n6267 gnd.n483 225.874
R6209 gnd.n6275 gnd.n483 225.874
R6210 gnd.n6276 gnd.n6275 225.874
R6211 gnd.n6277 gnd.n6276 225.874
R6212 gnd.n6277 gnd.n477 225.874
R6213 gnd.n6285 gnd.n477 225.874
R6214 gnd.n6286 gnd.n6285 225.874
R6215 gnd.n6287 gnd.n6286 225.874
R6216 gnd.n6287 gnd.n471 225.874
R6217 gnd.n6295 gnd.n471 225.874
R6218 gnd.n6296 gnd.n6295 225.874
R6219 gnd.n6297 gnd.n6296 225.874
R6220 gnd.n6297 gnd.n465 225.874
R6221 gnd.n6305 gnd.n465 225.874
R6222 gnd.n6306 gnd.n6305 225.874
R6223 gnd.n6307 gnd.n6306 225.874
R6224 gnd.n6307 gnd.n459 225.874
R6225 gnd.n6315 gnd.n459 225.874
R6226 gnd.n6316 gnd.n6315 225.874
R6227 gnd.n6317 gnd.n6316 225.874
R6228 gnd.n6317 gnd.n453 225.874
R6229 gnd.n6325 gnd.n453 225.874
R6230 gnd.n6326 gnd.n6325 225.874
R6231 gnd.n6327 gnd.n6326 225.874
R6232 gnd.n6327 gnd.n447 225.874
R6233 gnd.n6335 gnd.n447 225.874
R6234 gnd.n6336 gnd.n6335 225.874
R6235 gnd.n6337 gnd.n6336 225.874
R6236 gnd.n6337 gnd.n441 225.874
R6237 gnd.n6345 gnd.n441 225.874
R6238 gnd.n6346 gnd.n6345 225.874
R6239 gnd.n6347 gnd.n6346 225.874
R6240 gnd.n6347 gnd.n435 225.874
R6241 gnd.n6355 gnd.n435 225.874
R6242 gnd.n6356 gnd.n6355 225.874
R6243 gnd.n6357 gnd.n6356 225.874
R6244 gnd.n6357 gnd.n429 225.874
R6245 gnd.n6365 gnd.n429 225.874
R6246 gnd.n6366 gnd.n6365 225.874
R6247 gnd.n6367 gnd.n6366 225.874
R6248 gnd.n6367 gnd.n423 225.874
R6249 gnd.n6375 gnd.n423 225.874
R6250 gnd.n6376 gnd.n6375 225.874
R6251 gnd.n6377 gnd.n6376 225.874
R6252 gnd.n6377 gnd.n417 225.874
R6253 gnd.n6385 gnd.n417 225.874
R6254 gnd.n6386 gnd.n6385 225.874
R6255 gnd.n6387 gnd.n6386 225.874
R6256 gnd.n6387 gnd.n411 225.874
R6257 gnd.n6395 gnd.n411 225.874
R6258 gnd.n6396 gnd.n6395 225.874
R6259 gnd.n6397 gnd.n6396 225.874
R6260 gnd.n6397 gnd.n405 225.874
R6261 gnd.n6405 gnd.n405 225.874
R6262 gnd.n6406 gnd.n6405 225.874
R6263 gnd.n6407 gnd.n6406 225.874
R6264 gnd.n6407 gnd.n399 225.874
R6265 gnd.n6415 gnd.n399 225.874
R6266 gnd.n6416 gnd.n6415 225.874
R6267 gnd.n6417 gnd.n6416 225.874
R6268 gnd.n6417 gnd.n393 225.874
R6269 gnd.n6425 gnd.n393 225.874
R6270 gnd.n6426 gnd.n6425 225.874
R6271 gnd.n6427 gnd.n6426 225.874
R6272 gnd.n6427 gnd.n387 225.874
R6273 gnd.n6435 gnd.n387 225.874
R6274 gnd.n6436 gnd.n6435 225.874
R6275 gnd.n6437 gnd.n6436 225.874
R6276 gnd.n6437 gnd.n381 225.874
R6277 gnd.n6445 gnd.n381 225.874
R6278 gnd.n6446 gnd.n6445 225.874
R6279 gnd.n6447 gnd.n6446 225.874
R6280 gnd.n6447 gnd.n375 225.874
R6281 gnd.n6455 gnd.n375 225.874
R6282 gnd.n6456 gnd.n6455 225.874
R6283 gnd.n6457 gnd.n6456 225.874
R6284 gnd.n6457 gnd.n369 225.874
R6285 gnd.n6465 gnd.n369 225.874
R6286 gnd.n6466 gnd.n6465 225.874
R6287 gnd.n6467 gnd.n6466 225.874
R6288 gnd.n6467 gnd.n363 225.874
R6289 gnd.n6475 gnd.n363 225.874
R6290 gnd.n6476 gnd.n6475 225.874
R6291 gnd.n6477 gnd.n6476 225.874
R6292 gnd.n6477 gnd.n357 225.874
R6293 gnd.n6485 gnd.n357 225.874
R6294 gnd.n6486 gnd.n6485 225.874
R6295 gnd.n6487 gnd.n6486 225.874
R6296 gnd.n6487 gnd.n351 225.874
R6297 gnd.n6495 gnd.n351 225.874
R6298 gnd.n6496 gnd.n6495 225.874
R6299 gnd.n6497 gnd.n6496 225.874
R6300 gnd.n6497 gnd.n345 225.874
R6301 gnd.n6505 gnd.n345 225.874
R6302 gnd.n6506 gnd.n6505 225.874
R6303 gnd.n6507 gnd.n6506 225.874
R6304 gnd.n6507 gnd.n339 225.874
R6305 gnd.n6515 gnd.n339 225.874
R6306 gnd.n6516 gnd.n6515 225.874
R6307 gnd.n6517 gnd.n6516 225.874
R6308 gnd.n6517 gnd.n333 225.874
R6309 gnd.n6525 gnd.n333 225.874
R6310 gnd.n6526 gnd.n6525 225.874
R6311 gnd.n6527 gnd.n6526 225.874
R6312 gnd.n6527 gnd.n327 225.874
R6313 gnd.n6535 gnd.n327 225.874
R6314 gnd.n6536 gnd.n6535 225.874
R6315 gnd.n6537 gnd.n6536 225.874
R6316 gnd.n6537 gnd.n321 225.874
R6317 gnd.n6545 gnd.n321 225.874
R6318 gnd.n6546 gnd.n6545 225.874
R6319 gnd.n6547 gnd.n6546 225.874
R6320 gnd.n6547 gnd.n315 225.874
R6321 gnd.n6556 gnd.n315 225.874
R6322 gnd.n6557 gnd.n6556 225.874
R6323 gnd.n6558 gnd.n6557 225.874
R6324 gnd.n6558 gnd.n310 225.874
R6325 gnd.n2760 gnd.t117 224.174
R6326 gnd.n2270 gnd.t28 224.174
R6327 gnd.n5444 gnd.n1448 213.952
R6328 gnd.n5752 gnd.n5751 213.952
R6329 gnd.n1449 gnd.n1386 199.319
R6330 gnd.n1449 gnd.n1387 199.319
R6331 gnd.n1041 gnd.n996 199.319
R6332 gnd.n1041 gnd.n995 199.319
R6333 gnd.n1186 gnd.n1183 186.49
R6334 gnd.n4882 gnd.n4879 186.49
R6335 gnd.n3535 gnd.n3534 185
R6336 gnd.n3533 gnd.n3532 185
R6337 gnd.n3512 gnd.n3511 185
R6338 gnd.n3527 gnd.n3526 185
R6339 gnd.n3525 gnd.n3524 185
R6340 gnd.n3516 gnd.n3515 185
R6341 gnd.n3519 gnd.n3518 185
R6342 gnd.n3503 gnd.n3502 185
R6343 gnd.n3501 gnd.n3500 185
R6344 gnd.n3480 gnd.n3479 185
R6345 gnd.n3495 gnd.n3494 185
R6346 gnd.n3493 gnd.n3492 185
R6347 gnd.n3484 gnd.n3483 185
R6348 gnd.n3487 gnd.n3486 185
R6349 gnd.n3471 gnd.n3470 185
R6350 gnd.n3469 gnd.n3468 185
R6351 gnd.n3448 gnd.n3447 185
R6352 gnd.n3463 gnd.n3462 185
R6353 gnd.n3461 gnd.n3460 185
R6354 gnd.n3452 gnd.n3451 185
R6355 gnd.n3455 gnd.n3454 185
R6356 gnd.n3440 gnd.n3439 185
R6357 gnd.n3438 gnd.n3437 185
R6358 gnd.n3417 gnd.n3416 185
R6359 gnd.n3432 gnd.n3431 185
R6360 gnd.n3430 gnd.n3429 185
R6361 gnd.n3421 gnd.n3420 185
R6362 gnd.n3424 gnd.n3423 185
R6363 gnd.n3408 gnd.n3407 185
R6364 gnd.n3406 gnd.n3405 185
R6365 gnd.n3385 gnd.n3384 185
R6366 gnd.n3400 gnd.n3399 185
R6367 gnd.n3398 gnd.n3397 185
R6368 gnd.n3389 gnd.n3388 185
R6369 gnd.n3392 gnd.n3391 185
R6370 gnd.n3376 gnd.n3375 185
R6371 gnd.n3374 gnd.n3373 185
R6372 gnd.n3353 gnd.n3352 185
R6373 gnd.n3368 gnd.n3367 185
R6374 gnd.n3366 gnd.n3365 185
R6375 gnd.n3357 gnd.n3356 185
R6376 gnd.n3360 gnd.n3359 185
R6377 gnd.n3344 gnd.n3343 185
R6378 gnd.n3342 gnd.n3341 185
R6379 gnd.n3321 gnd.n3320 185
R6380 gnd.n3336 gnd.n3335 185
R6381 gnd.n3334 gnd.n3333 185
R6382 gnd.n3325 gnd.n3324 185
R6383 gnd.n3328 gnd.n3327 185
R6384 gnd.n3313 gnd.n3312 185
R6385 gnd.n3311 gnd.n3310 185
R6386 gnd.n3290 gnd.n3289 185
R6387 gnd.n3305 gnd.n3304 185
R6388 gnd.n3303 gnd.n3302 185
R6389 gnd.n3294 gnd.n3293 185
R6390 gnd.n3297 gnd.n3296 185
R6391 gnd.n2761 gnd.t116 178.987
R6392 gnd.n2271 gnd.t29 178.987
R6393 gnd.n1 gnd.t172 170.774
R6394 gnd.n9 gnd.t193 170.103
R6395 gnd.n8 gnd.t191 170.103
R6396 gnd.n7 gnd.t152 170.103
R6397 gnd.n6 gnd.t184 170.103
R6398 gnd.n5 gnd.t127 170.103
R6399 gnd.n4 gnd.t137 170.103
R6400 gnd.n3 gnd.t317 170.103
R6401 gnd.n2 gnd.t1 170.103
R6402 gnd.n1 gnd.t165 170.103
R6403 gnd.n4953 gnd.n4952 163.367
R6404 gnd.n4949 gnd.n4948 163.367
R6405 gnd.n4945 gnd.n4944 163.367
R6406 gnd.n4941 gnd.n4940 163.367
R6407 gnd.n4937 gnd.n4936 163.367
R6408 gnd.n4933 gnd.n4932 163.367
R6409 gnd.n4929 gnd.n4928 163.367
R6410 gnd.n4925 gnd.n4924 163.367
R6411 gnd.n4921 gnd.n4920 163.367
R6412 gnd.n4917 gnd.n4916 163.367
R6413 gnd.n4913 gnd.n4912 163.367
R6414 gnd.n4909 gnd.n4908 163.367
R6415 gnd.n4905 gnd.n4904 163.367
R6416 gnd.n4901 gnd.n4900 163.367
R6417 gnd.n4896 gnd.n4895 163.367
R6418 gnd.n4892 gnd.n4891 163.367
R6419 gnd.n5029 gnd.n5028 163.367
R6420 gnd.n5025 gnd.n5024 163.367
R6421 gnd.n5020 gnd.n5019 163.367
R6422 gnd.n5016 gnd.n5015 163.367
R6423 gnd.n5012 gnd.n5011 163.367
R6424 gnd.n5008 gnd.n5007 163.367
R6425 gnd.n5004 gnd.n5003 163.367
R6426 gnd.n5000 gnd.n4999 163.367
R6427 gnd.n4996 gnd.n4995 163.367
R6428 gnd.n4992 gnd.n4991 163.367
R6429 gnd.n4988 gnd.n4987 163.367
R6430 gnd.n4984 gnd.n4983 163.367
R6431 gnd.n4980 gnd.n4979 163.367
R6432 gnd.n4976 gnd.n4975 163.367
R6433 gnd.n4972 gnd.n4971 163.367
R6434 gnd.n4968 gnd.n4967 163.367
R6435 gnd.n4501 gnd.n1202 163.367
R6436 gnd.n4504 gnd.n1202 163.367
R6437 gnd.n4504 gnd.n4433 163.367
R6438 gnd.n4507 gnd.n4433 163.367
R6439 gnd.n4507 gnd.n4435 163.367
R6440 gnd.n4520 gnd.n4435 163.367
R6441 gnd.n4520 gnd.n1974 163.367
R6442 gnd.n4516 gnd.n1974 163.367
R6443 gnd.n4516 gnd.n1970 163.367
R6444 gnd.n4513 gnd.n1970 163.367
R6445 gnd.n4513 gnd.n1958 163.367
R6446 gnd.n1958 gnd.n1953 163.367
R6447 gnd.n4575 gnd.n1953 163.367
R6448 gnd.n4576 gnd.n4575 163.367
R6449 gnd.n4576 gnd.n1942 163.367
R6450 gnd.n1950 gnd.n1942 163.367
R6451 gnd.n4594 gnd.n1950 163.367
R6452 gnd.n4594 gnd.n1951 163.367
R6453 gnd.n4590 gnd.n1951 163.367
R6454 gnd.n4590 gnd.n1925 163.367
R6455 gnd.n4585 gnd.n1925 163.367
R6456 gnd.n4585 gnd.n1921 163.367
R6457 gnd.n4582 gnd.n1921 163.367
R6458 gnd.n4582 gnd.n1911 163.367
R6459 gnd.n1911 gnd.n1902 163.367
R6460 gnd.n4689 gnd.n1902 163.367
R6461 gnd.n4689 gnd.n1900 163.367
R6462 gnd.n4694 gnd.n1900 163.367
R6463 gnd.n4694 gnd.n1892 163.367
R6464 gnd.n4703 gnd.n1892 163.367
R6465 gnd.n4704 gnd.n4703 163.367
R6466 gnd.n4704 gnd.n1889 163.367
R6467 gnd.n4713 gnd.n1889 163.367
R6468 gnd.n4713 gnd.n1883 163.367
R6469 gnd.n4709 gnd.n1883 163.367
R6470 gnd.n4709 gnd.n1874 163.367
R6471 gnd.n1874 gnd.n1869 163.367
R6472 gnd.n4739 gnd.n1869 163.367
R6473 gnd.n4740 gnd.n4739 163.367
R6474 gnd.n4740 gnd.n1861 163.367
R6475 gnd.n4746 gnd.n1861 163.367
R6476 gnd.n4746 gnd.n1866 163.367
R6477 gnd.n4759 gnd.n1866 163.367
R6478 gnd.n4759 gnd.n1867 163.367
R6479 gnd.n1867 gnd.n1845 163.367
R6480 gnd.n4754 gnd.n1845 163.367
R6481 gnd.n4754 gnd.n1840 163.367
R6482 gnd.n4751 gnd.n1840 163.367
R6483 gnd.n4751 gnd.n1830 163.367
R6484 gnd.n1830 gnd.n1822 163.367
R6485 gnd.n4839 gnd.n1822 163.367
R6486 gnd.n4839 gnd.n1819 163.367
R6487 gnd.n4849 gnd.n1819 163.367
R6488 gnd.n4849 gnd.n1820 163.367
R6489 gnd.n1820 gnd.n1813 163.367
R6490 gnd.n4844 gnd.n1813 163.367
R6491 gnd.n4844 gnd.n1803 163.367
R6492 gnd.n1803 gnd.n1794 163.367
R6493 gnd.n4962 gnd.n1794 163.367
R6494 gnd.n4963 gnd.n4962 163.367
R6495 gnd.n1177 gnd.n1176 163.367
R6496 gnd.n5741 gnd.n1176 163.367
R6497 gnd.n5739 gnd.n5738 163.367
R6498 gnd.n5735 gnd.n5734 163.367
R6499 gnd.n5731 gnd.n5730 163.367
R6500 gnd.n5727 gnd.n5726 163.367
R6501 gnd.n5723 gnd.n5722 163.367
R6502 gnd.n5719 gnd.n5718 163.367
R6503 gnd.n5715 gnd.n5714 163.367
R6504 gnd.n5711 gnd.n5710 163.367
R6505 gnd.n5707 gnd.n5706 163.367
R6506 gnd.n5703 gnd.n5702 163.367
R6507 gnd.n5699 gnd.n5698 163.367
R6508 gnd.n5695 gnd.n5694 163.367
R6509 gnd.n5691 gnd.n5690 163.367
R6510 gnd.n5687 gnd.n5686 163.367
R6511 gnd.n5750 gnd.n1142 163.367
R6512 gnd.n4440 gnd.n4439 163.367
R6513 gnd.n4445 gnd.n4444 163.367
R6514 gnd.n4449 gnd.n4448 163.367
R6515 gnd.n4453 gnd.n4452 163.367
R6516 gnd.n4457 gnd.n4456 163.367
R6517 gnd.n4461 gnd.n4460 163.367
R6518 gnd.n4465 gnd.n4464 163.367
R6519 gnd.n4469 gnd.n4468 163.367
R6520 gnd.n4473 gnd.n4472 163.367
R6521 gnd.n4477 gnd.n4476 163.367
R6522 gnd.n4481 gnd.n4480 163.367
R6523 gnd.n4485 gnd.n4484 163.367
R6524 gnd.n4489 gnd.n4488 163.367
R6525 gnd.n4493 gnd.n4492 163.367
R6526 gnd.n4497 gnd.n4496 163.367
R6527 gnd.n5679 gnd.n1178 163.367
R6528 gnd.n5679 gnd.n1200 163.367
R6529 gnd.n4528 gnd.n1200 163.367
R6530 gnd.n4528 gnd.n4434 163.367
R6531 gnd.n4524 gnd.n4434 163.367
R6532 gnd.n4524 gnd.n1973 163.367
R6533 gnd.n4553 gnd.n1973 163.367
R6534 gnd.n4553 gnd.n1971 163.367
R6535 gnd.n4557 gnd.n1971 163.367
R6536 gnd.n4557 gnd.n1956 163.367
R6537 gnd.n4569 gnd.n1956 163.367
R6538 gnd.n4569 gnd.n1954 163.367
R6539 gnd.n4573 gnd.n1954 163.367
R6540 gnd.n4573 gnd.n1944 163.367
R6541 gnd.n4600 gnd.n1944 163.367
R6542 gnd.n4600 gnd.n1945 163.367
R6543 gnd.n4596 gnd.n1945 163.367
R6544 gnd.n4596 gnd.n1948 163.367
R6545 gnd.n1948 gnd.n1924 163.367
R6546 gnd.n4656 gnd.n1924 163.367
R6547 gnd.n4656 gnd.n1922 163.367
R6548 gnd.n4660 gnd.n1922 163.367
R6549 gnd.n4660 gnd.n1908 163.367
R6550 gnd.n4683 gnd.n1908 163.367
R6551 gnd.n4683 gnd.n1906 163.367
R6552 gnd.n4687 gnd.n1906 163.367
R6553 gnd.n4687 gnd.n1898 163.367
R6554 gnd.n4697 gnd.n1898 163.367
R6555 gnd.n4697 gnd.n1896 163.367
R6556 gnd.n4701 gnd.n1896 163.367
R6557 gnd.n4701 gnd.n1887 163.367
R6558 gnd.n4717 gnd.n1887 163.367
R6559 gnd.n4717 gnd.n1885 163.367
R6560 gnd.n4721 gnd.n1885 163.367
R6561 gnd.n4721 gnd.n1873 163.367
R6562 gnd.n4733 gnd.n1873 163.367
R6563 gnd.n4733 gnd.n1871 163.367
R6564 gnd.n4737 gnd.n1871 163.367
R6565 gnd.n4737 gnd.n1862 163.367
R6566 gnd.n4767 gnd.n1862 163.367
R6567 gnd.n4767 gnd.n1863 163.367
R6568 gnd.n4763 gnd.n1863 163.367
R6569 gnd.n4763 gnd.n4762 163.367
R6570 gnd.n4762 gnd.n1843 163.367
R6571 gnd.n4814 gnd.n1843 163.367
R6572 gnd.n4814 gnd.n1841 163.367
R6573 gnd.n4818 gnd.n1841 163.367
R6574 gnd.n4818 gnd.n1828 163.367
R6575 gnd.n4833 gnd.n1828 163.367
R6576 gnd.n4833 gnd.n1826 163.367
R6577 gnd.n4837 gnd.n1826 163.367
R6578 gnd.n4837 gnd.n1816 163.367
R6579 gnd.n4851 gnd.n1816 163.367
R6580 gnd.n4851 gnd.n1814 163.367
R6581 gnd.n4855 gnd.n1814 163.367
R6582 gnd.n4855 gnd.n1801 163.367
R6583 gnd.n4867 gnd.n1801 163.367
R6584 gnd.n4867 gnd.n1798 163.367
R6585 gnd.n4960 gnd.n1798 163.367
R6586 gnd.n4960 gnd.n1799 163.367
R6587 gnd.n4888 gnd.n4887 156.462
R6588 gnd.n3475 gnd.n3443 153.042
R6589 gnd.n3539 gnd.n3538 152.079
R6590 gnd.n3507 gnd.n3506 152.079
R6591 gnd.n3475 gnd.n3474 152.079
R6592 gnd.n1191 gnd.n1190 152
R6593 gnd.n1192 gnd.n1181 152
R6594 gnd.n1194 gnd.n1193 152
R6595 gnd.n1196 gnd.n1179 152
R6596 gnd.n1198 gnd.n1197 152
R6597 gnd.n4886 gnd.n4870 152
R6598 gnd.n4878 gnd.n4871 152
R6599 gnd.n4877 gnd.n4876 152
R6600 gnd.n4875 gnd.n4872 152
R6601 gnd.n4873 gnd.t59 150.546
R6602 gnd.t154 gnd.n3517 147.661
R6603 gnd.t182 gnd.n3485 147.661
R6604 gnd.t170 gnd.n3453 147.661
R6605 gnd.t134 gnd.n3422 147.661
R6606 gnd.t167 gnd.n3390 147.661
R6607 gnd.t178 gnd.n3358 147.661
R6608 gnd.t149 gnd.n3326 147.661
R6609 gnd.t159 gnd.n3295 147.661
R6610 gnd.n6567 gnd.n6566 143.933
R6611 gnd.n6568 gnd.n6567 143.933
R6612 gnd.n6568 gnd.n304 143.933
R6613 gnd.n6576 gnd.n304 143.933
R6614 gnd.n6577 gnd.n6576 143.933
R6615 gnd.n6578 gnd.n6577 143.933
R6616 gnd.n6578 gnd.n298 143.933
R6617 gnd.n6586 gnd.n298 143.933
R6618 gnd.n6587 gnd.n6586 143.933
R6619 gnd.n6588 gnd.n6587 143.933
R6620 gnd.n6588 gnd.n292 143.933
R6621 gnd.n6596 gnd.n292 143.933
R6622 gnd.n6597 gnd.n6596 143.933
R6623 gnd.n6598 gnd.n6597 143.933
R6624 gnd.n6598 gnd.n286 143.933
R6625 gnd.n6606 gnd.n286 143.933
R6626 gnd.n6607 gnd.n6606 143.933
R6627 gnd.n6608 gnd.n6607 143.933
R6628 gnd.n6608 gnd.n280 143.933
R6629 gnd.n6616 gnd.n280 143.933
R6630 gnd.n6617 gnd.n6616 143.933
R6631 gnd.n6618 gnd.n6617 143.933
R6632 gnd.n6618 gnd.n274 143.933
R6633 gnd.n6626 gnd.n274 143.933
R6634 gnd.n6627 gnd.n6626 143.933
R6635 gnd.n6628 gnd.n6627 143.933
R6636 gnd.n6628 gnd.n268 143.933
R6637 gnd.n6636 gnd.n268 143.933
R6638 gnd.n6637 gnd.n6636 143.933
R6639 gnd.n6638 gnd.n6637 143.933
R6640 gnd.n6638 gnd.n262 143.933
R6641 gnd.n6646 gnd.n262 143.933
R6642 gnd.n6647 gnd.n6646 143.933
R6643 gnd.n6648 gnd.n6647 143.933
R6644 gnd.n6648 gnd.n256 143.933
R6645 gnd.n6656 gnd.n256 143.933
R6646 gnd.n6657 gnd.n6656 143.933
R6647 gnd.n6658 gnd.n6657 143.933
R6648 gnd.n6658 gnd.n250 143.933
R6649 gnd.n6666 gnd.n250 143.933
R6650 gnd.n6667 gnd.n6666 143.933
R6651 gnd.n6668 gnd.n6667 143.933
R6652 gnd.n6668 gnd.n244 143.933
R6653 gnd.n6676 gnd.n244 143.933
R6654 gnd.n6677 gnd.n6676 143.933
R6655 gnd.n6678 gnd.n6677 143.933
R6656 gnd.n6678 gnd.n238 143.933
R6657 gnd.n6686 gnd.n238 143.933
R6658 gnd.n6687 gnd.n6686 143.933
R6659 gnd.n6688 gnd.n6687 143.933
R6660 gnd.n6688 gnd.n232 143.933
R6661 gnd.n6696 gnd.n232 143.933
R6662 gnd.n6697 gnd.n6696 143.933
R6663 gnd.n6698 gnd.n6697 143.933
R6664 gnd.n6698 gnd.n226 143.933
R6665 gnd.n6706 gnd.n226 143.933
R6666 gnd.n6707 gnd.n6706 143.933
R6667 gnd.n6708 gnd.n6707 143.933
R6668 gnd.n6708 gnd.n220 143.933
R6669 gnd.n6716 gnd.n220 143.933
R6670 gnd.n6717 gnd.n6716 143.933
R6671 gnd.n6718 gnd.n6717 143.933
R6672 gnd.n6718 gnd.n214 143.933
R6673 gnd.n6726 gnd.n214 143.933
R6674 gnd.n6727 gnd.n6726 143.933
R6675 gnd.n6728 gnd.n6727 143.933
R6676 gnd.n6728 gnd.n208 143.933
R6677 gnd.n6736 gnd.n208 143.933
R6678 gnd.n6737 gnd.n6736 143.933
R6679 gnd.n6738 gnd.n6737 143.933
R6680 gnd.n6738 gnd.n202 143.933
R6681 gnd.n6746 gnd.n202 143.933
R6682 gnd.n6747 gnd.n6746 143.933
R6683 gnd.n6748 gnd.n6747 143.933
R6684 gnd.n6748 gnd.n196 143.933
R6685 gnd.n6756 gnd.n196 143.933
R6686 gnd.n6757 gnd.n6756 143.933
R6687 gnd.n6758 gnd.n6757 143.933
R6688 gnd.n6758 gnd.n190 143.933
R6689 gnd.n6766 gnd.n190 143.933
R6690 gnd.n6767 gnd.n6766 143.933
R6691 gnd.n6769 gnd.n6767 143.933
R6692 gnd.n6769 gnd.n6768 143.933
R6693 gnd.n1790 gnd.n1773 143.351
R6694 gnd.n1158 gnd.n1141 143.351
R6695 gnd.n5749 gnd.n1141 143.351
R6696 gnd.n1188 gnd.t107 130.484
R6697 gnd.n1197 gnd.t101 126.766
R6698 gnd.n1195 gnd.t86 126.766
R6699 gnd.n1181 gnd.t13 126.766
R6700 gnd.n1189 gnd.t62 126.766
R6701 gnd.n4874 gnd.t2 126.766
R6702 gnd.n4876 gnd.t80 126.766
R6703 gnd.n4885 gnd.t98 126.766
R6704 gnd.n4887 gnd.t42 126.766
R6705 gnd.n3534 gnd.n3533 104.615
R6706 gnd.n3533 gnd.n3511 104.615
R6707 gnd.n3526 gnd.n3511 104.615
R6708 gnd.n3526 gnd.n3525 104.615
R6709 gnd.n3525 gnd.n3515 104.615
R6710 gnd.n3518 gnd.n3515 104.615
R6711 gnd.n3502 gnd.n3501 104.615
R6712 gnd.n3501 gnd.n3479 104.615
R6713 gnd.n3494 gnd.n3479 104.615
R6714 gnd.n3494 gnd.n3493 104.615
R6715 gnd.n3493 gnd.n3483 104.615
R6716 gnd.n3486 gnd.n3483 104.615
R6717 gnd.n3470 gnd.n3469 104.615
R6718 gnd.n3469 gnd.n3447 104.615
R6719 gnd.n3462 gnd.n3447 104.615
R6720 gnd.n3462 gnd.n3461 104.615
R6721 gnd.n3461 gnd.n3451 104.615
R6722 gnd.n3454 gnd.n3451 104.615
R6723 gnd.n3439 gnd.n3438 104.615
R6724 gnd.n3438 gnd.n3416 104.615
R6725 gnd.n3431 gnd.n3416 104.615
R6726 gnd.n3431 gnd.n3430 104.615
R6727 gnd.n3430 gnd.n3420 104.615
R6728 gnd.n3423 gnd.n3420 104.615
R6729 gnd.n3407 gnd.n3406 104.615
R6730 gnd.n3406 gnd.n3384 104.615
R6731 gnd.n3399 gnd.n3384 104.615
R6732 gnd.n3399 gnd.n3398 104.615
R6733 gnd.n3398 gnd.n3388 104.615
R6734 gnd.n3391 gnd.n3388 104.615
R6735 gnd.n3375 gnd.n3374 104.615
R6736 gnd.n3374 gnd.n3352 104.615
R6737 gnd.n3367 gnd.n3352 104.615
R6738 gnd.n3367 gnd.n3366 104.615
R6739 gnd.n3366 gnd.n3356 104.615
R6740 gnd.n3359 gnd.n3356 104.615
R6741 gnd.n3343 gnd.n3342 104.615
R6742 gnd.n3342 gnd.n3320 104.615
R6743 gnd.n3335 gnd.n3320 104.615
R6744 gnd.n3335 gnd.n3334 104.615
R6745 gnd.n3334 gnd.n3324 104.615
R6746 gnd.n3327 gnd.n3324 104.615
R6747 gnd.n3312 gnd.n3311 104.615
R6748 gnd.n3311 gnd.n3289 104.615
R6749 gnd.n3304 gnd.n3289 104.615
R6750 gnd.n3304 gnd.n3303 104.615
R6751 gnd.n3303 gnd.n3293 104.615
R6752 gnd.n3296 gnd.n3293 104.615
R6753 gnd.n2686 gnd.t55 100.632
R6754 gnd.n2244 gnd.t112 100.632
R6755 gnd.n7085 gnd.n7084 99.6594
R6756 gnd.n7080 gnd.n6901 99.6594
R6757 gnd.n7076 gnd.n6900 99.6594
R6758 gnd.n7072 gnd.n6899 99.6594
R6759 gnd.n7068 gnd.n6898 99.6594
R6760 gnd.n7064 gnd.n6897 99.6594
R6761 gnd.n7060 gnd.n6896 99.6594
R6762 gnd.n7056 gnd.n6895 99.6594
R6763 gnd.n7049 gnd.n6894 99.6594
R6764 gnd.n7045 gnd.n6893 99.6594
R6765 gnd.n7041 gnd.n6892 99.6594
R6766 gnd.n7037 gnd.n6891 99.6594
R6767 gnd.n7033 gnd.n6890 99.6594
R6768 gnd.n7029 gnd.n6889 99.6594
R6769 gnd.n7025 gnd.n6888 99.6594
R6770 gnd.n7021 gnd.n6887 99.6594
R6771 gnd.n7017 gnd.n6886 99.6594
R6772 gnd.n7013 gnd.n6885 99.6594
R6773 gnd.n7005 gnd.n6884 99.6594
R6774 gnd.n7003 gnd.n6883 99.6594
R6775 gnd.n6999 gnd.n6882 99.6594
R6776 gnd.n6995 gnd.n6881 99.6594
R6777 gnd.n6991 gnd.n6880 99.6594
R6778 gnd.n6987 gnd.n6879 99.6594
R6779 gnd.n6983 gnd.n6878 99.6594
R6780 gnd.n6979 gnd.n6877 99.6594
R6781 gnd.n6975 gnd.n6876 99.6594
R6782 gnd.n6971 gnd.n6875 99.6594
R6783 gnd.n6963 gnd.n6874 99.6594
R6784 gnd.n5496 gnd.n5495 99.6594
R6785 gnd.n5490 gnd.n1375 99.6594
R6786 gnd.n5487 gnd.n1376 99.6594
R6787 gnd.n5483 gnd.n1377 99.6594
R6788 gnd.n5479 gnd.n1378 99.6594
R6789 gnd.n5475 gnd.n1379 99.6594
R6790 gnd.n5471 gnd.n1380 99.6594
R6791 gnd.n5467 gnd.n1381 99.6594
R6792 gnd.n5463 gnd.n1382 99.6594
R6793 gnd.n5458 gnd.n1383 99.6594
R6794 gnd.n5454 gnd.n1384 99.6594
R6795 gnd.n5450 gnd.n1385 99.6594
R6796 gnd.n5446 gnd.n1386 99.6594
R6797 gnd.n5441 gnd.n1388 99.6594
R6798 gnd.n5437 gnd.n1389 99.6594
R6799 gnd.n5433 gnd.n1390 99.6594
R6800 gnd.n5429 gnd.n1391 99.6594
R6801 gnd.n5425 gnd.n1392 99.6594
R6802 gnd.n5421 gnd.n1393 99.6594
R6803 gnd.n5417 gnd.n1394 99.6594
R6804 gnd.n5413 gnd.n1395 99.6594
R6805 gnd.n5409 gnd.n1396 99.6594
R6806 gnd.n5405 gnd.n1397 99.6594
R6807 gnd.n5401 gnd.n1398 99.6594
R6808 gnd.n5397 gnd.n1399 99.6594
R6809 gnd.n5393 gnd.n1400 99.6594
R6810 gnd.n5389 gnd.n1401 99.6594
R6811 gnd.n5385 gnd.n1402 99.6594
R6812 gnd.n5801 gnd.n5800 99.6594
R6813 gnd.n5796 gnd.n1007 99.6594
R6814 gnd.n5792 gnd.n1006 99.6594
R6815 gnd.n5788 gnd.n1005 99.6594
R6816 gnd.n5784 gnd.n1004 99.6594
R6817 gnd.n5780 gnd.n1003 99.6594
R6818 gnd.n5776 gnd.n1002 99.6594
R6819 gnd.n5772 gnd.n1001 99.6594
R6820 gnd.n5767 gnd.n1000 99.6594
R6821 gnd.n5763 gnd.n999 99.6594
R6822 gnd.n5759 gnd.n998 99.6594
R6823 gnd.n5755 gnd.n997 99.6594
R6824 gnd.n1133 gnd.n995 99.6594
R6825 gnd.n1131 gnd.n994 99.6594
R6826 gnd.n1127 gnd.n993 99.6594
R6827 gnd.n1123 gnd.n992 99.6594
R6828 gnd.n1119 gnd.n991 99.6594
R6829 gnd.n1111 gnd.n990 99.6594
R6830 gnd.n1109 gnd.n989 99.6594
R6831 gnd.n1105 gnd.n988 99.6594
R6832 gnd.n1101 gnd.n987 99.6594
R6833 gnd.n1097 gnd.n986 99.6594
R6834 gnd.n1093 gnd.n985 99.6594
R6835 gnd.n1089 gnd.n984 99.6594
R6836 gnd.n1085 gnd.n983 99.6594
R6837 gnd.n1081 gnd.n982 99.6594
R6838 gnd.n1077 gnd.n981 99.6594
R6839 gnd.n1069 gnd.n980 99.6594
R6840 gnd.n3953 gnd.n3745 99.6594
R6841 gnd.n3951 gnd.n3748 99.6594
R6842 gnd.n3947 gnd.n3946 99.6594
R6843 gnd.n3940 gnd.n3753 99.6594
R6844 gnd.n3939 gnd.n3938 99.6594
R6845 gnd.n3932 gnd.n3759 99.6594
R6846 gnd.n3931 gnd.n3930 99.6594
R6847 gnd.n3924 gnd.n3765 99.6594
R6848 gnd.n3923 gnd.n3922 99.6594
R6849 gnd.n3916 gnd.n3771 99.6594
R6850 gnd.n3915 gnd.n3914 99.6594
R6851 gnd.n3908 gnd.n3780 99.6594
R6852 gnd.n3907 gnd.n3906 99.6594
R6853 gnd.n3900 gnd.n3786 99.6594
R6854 gnd.n3899 gnd.n3898 99.6594
R6855 gnd.n3892 gnd.n3792 99.6594
R6856 gnd.n3891 gnd.n3890 99.6594
R6857 gnd.n3884 gnd.n3798 99.6594
R6858 gnd.n3883 gnd.n3882 99.6594
R6859 gnd.n3876 gnd.n3806 99.6594
R6860 gnd.n3875 gnd.n3874 99.6594
R6861 gnd.n3868 gnd.n3812 99.6594
R6862 gnd.n3867 gnd.n3866 99.6594
R6863 gnd.n3860 gnd.n3818 99.6594
R6864 gnd.n3859 gnd.n3858 99.6594
R6865 gnd.n3852 gnd.n3824 99.6594
R6866 gnd.n3851 gnd.n3850 99.6594
R6867 gnd.n3844 gnd.n3830 99.6594
R6868 gnd.n3843 gnd.n3842 99.6594
R6869 gnd.n3657 gnd.n2227 99.6594
R6870 gnd.n3655 gnd.n2226 99.6594
R6871 gnd.n3651 gnd.n2225 99.6594
R6872 gnd.n3647 gnd.n2224 99.6594
R6873 gnd.n3643 gnd.n2223 99.6594
R6874 gnd.n3639 gnd.n2222 99.6594
R6875 gnd.n3635 gnd.n2221 99.6594
R6876 gnd.n3567 gnd.n2220 99.6594
R6877 gnd.n2898 gnd.n2629 99.6594
R6878 gnd.n2655 gnd.n2636 99.6594
R6879 gnd.n2657 gnd.n2637 99.6594
R6880 gnd.n2665 gnd.n2638 99.6594
R6881 gnd.n2667 gnd.n2639 99.6594
R6882 gnd.n2675 gnd.n2640 99.6594
R6883 gnd.n2677 gnd.n2641 99.6594
R6884 gnd.n2685 gnd.n2642 99.6594
R6885 gnd.n6837 gnd.n6816 99.6594
R6886 gnd.n6843 gnd.n6817 99.6594
R6887 gnd.n6847 gnd.n6818 99.6594
R6888 gnd.n6853 gnd.n6819 99.6594
R6889 gnd.n6857 gnd.n6820 99.6594
R6890 gnd.n6863 gnd.n6821 99.6594
R6891 gnd.n6866 gnd.n6822 99.6594
R6892 gnd.n6873 gnd.n6872 99.6594
R6893 gnd.n7088 gnd.n7087 99.6594
R6894 gnd.n1487 gnd.n1403 99.6594
R6895 gnd.n1405 gnd.n1329 99.6594
R6896 gnd.n1406 gnd.n1336 99.6594
R6897 gnd.n1408 gnd.n1407 99.6594
R6898 gnd.n1410 gnd.n1345 99.6594
R6899 gnd.n1411 gnd.n1352 99.6594
R6900 gnd.n1413 gnd.n1412 99.6594
R6901 gnd.n1415 gnd.n1361 99.6594
R6902 gnd.n5498 gnd.n1370 99.6594
R6903 gnd.n3625 gnd.n2207 99.6594
R6904 gnd.n3621 gnd.n2208 99.6594
R6905 gnd.n3617 gnd.n2209 99.6594
R6906 gnd.n3613 gnd.n2210 99.6594
R6907 gnd.n3609 gnd.n2211 99.6594
R6908 gnd.n3605 gnd.n2212 99.6594
R6909 gnd.n3601 gnd.n2213 99.6594
R6910 gnd.n3597 gnd.n2214 99.6594
R6911 gnd.n3593 gnd.n2215 99.6594
R6912 gnd.n3589 gnd.n2216 99.6594
R6913 gnd.n3585 gnd.n2217 99.6594
R6914 gnd.n3581 gnd.n2218 99.6594
R6915 gnd.n3577 gnd.n2219 99.6594
R6916 gnd.n2813 gnd.n2812 99.6594
R6917 gnd.n2807 gnd.n2724 99.6594
R6918 gnd.n2804 gnd.n2725 99.6594
R6919 gnd.n2800 gnd.n2726 99.6594
R6920 gnd.n2796 gnd.n2727 99.6594
R6921 gnd.n2792 gnd.n2728 99.6594
R6922 gnd.n2788 gnd.n2729 99.6594
R6923 gnd.n2784 gnd.n2730 99.6594
R6924 gnd.n2780 gnd.n2731 99.6594
R6925 gnd.n2776 gnd.n2732 99.6594
R6926 gnd.n2772 gnd.n2733 99.6594
R6927 gnd.n2768 gnd.n2734 99.6594
R6928 gnd.n2815 gnd.n2723 99.6594
R6929 gnd.n966 gnd.n911 99.6594
R6930 gnd.n968 gnd.n920 99.6594
R6931 gnd.n970 gnd.n969 99.6594
R6932 gnd.n971 gnd.n929 99.6594
R6933 gnd.n973 gnd.n938 99.6594
R6934 gnd.n975 gnd.n974 99.6594
R6935 gnd.n976 gnd.n947 99.6594
R6936 gnd.n978 gnd.n959 99.6594
R6937 gnd.n5804 gnd.n5803 99.6594
R6938 gnd.n3693 gnd.n2204 99.6594
R6939 gnd.n3696 gnd.n3695 99.6594
R6940 gnd.n3703 gnd.n3702 99.6594
R6941 gnd.n3706 gnd.n3705 99.6594
R6942 gnd.n3713 gnd.n3712 99.6594
R6943 gnd.n3716 gnd.n3715 99.6594
R6944 gnd.n3723 gnd.n3722 99.6594
R6945 gnd.n3726 gnd.n3725 99.6594
R6946 gnd.n3733 gnd.n3732 99.6594
R6947 gnd.n3694 gnd.n3693 99.6594
R6948 gnd.n3695 gnd.n3687 99.6594
R6949 gnd.n3704 gnd.n3703 99.6594
R6950 gnd.n3705 gnd.n3683 99.6594
R6951 gnd.n3714 gnd.n3713 99.6594
R6952 gnd.n3715 gnd.n3679 99.6594
R6953 gnd.n3724 gnd.n3723 99.6594
R6954 gnd.n3725 gnd.n3675 99.6594
R6955 gnd.n3734 gnd.n3733 99.6594
R6956 gnd.n5803 gnd.n964 99.6594
R6957 gnd.n978 gnd.n977 99.6594
R6958 gnd.n976 gnd.n946 99.6594
R6959 gnd.n975 gnd.n939 99.6594
R6960 gnd.n973 gnd.n972 99.6594
R6961 gnd.n971 gnd.n928 99.6594
R6962 gnd.n970 gnd.n921 99.6594
R6963 gnd.n968 gnd.n967 99.6594
R6964 gnd.n966 gnd.n910 99.6594
R6965 gnd.n2813 gnd.n2736 99.6594
R6966 gnd.n2805 gnd.n2724 99.6594
R6967 gnd.n2801 gnd.n2725 99.6594
R6968 gnd.n2797 gnd.n2726 99.6594
R6969 gnd.n2793 gnd.n2727 99.6594
R6970 gnd.n2789 gnd.n2728 99.6594
R6971 gnd.n2785 gnd.n2729 99.6594
R6972 gnd.n2781 gnd.n2730 99.6594
R6973 gnd.n2777 gnd.n2731 99.6594
R6974 gnd.n2773 gnd.n2732 99.6594
R6975 gnd.n2769 gnd.n2733 99.6594
R6976 gnd.n2765 gnd.n2734 99.6594
R6977 gnd.n2816 gnd.n2815 99.6594
R6978 gnd.n3580 gnd.n2219 99.6594
R6979 gnd.n3584 gnd.n2218 99.6594
R6980 gnd.n3588 gnd.n2217 99.6594
R6981 gnd.n3592 gnd.n2216 99.6594
R6982 gnd.n3596 gnd.n2215 99.6594
R6983 gnd.n3600 gnd.n2214 99.6594
R6984 gnd.n3604 gnd.n2213 99.6594
R6985 gnd.n3608 gnd.n2212 99.6594
R6986 gnd.n3612 gnd.n2211 99.6594
R6987 gnd.n3616 gnd.n2210 99.6594
R6988 gnd.n3620 gnd.n2209 99.6594
R6989 gnd.n3624 gnd.n2208 99.6594
R6990 gnd.n2248 gnd.n2207 99.6594
R6991 gnd.n1403 gnd.n1328 99.6594
R6992 gnd.n1405 gnd.n1404 99.6594
R6993 gnd.n1406 gnd.n1337 99.6594
R6994 gnd.n1408 gnd.n1344 99.6594
R6995 gnd.n1410 gnd.n1409 99.6594
R6996 gnd.n1411 gnd.n1353 99.6594
R6997 gnd.n1413 gnd.n1360 99.6594
R6998 gnd.n1415 gnd.n1414 99.6594
R6999 gnd.n5499 gnd.n5498 99.6594
R7000 gnd.n7087 gnd.n6815 99.6594
R7001 gnd.n6873 gnd.n6823 99.6594
R7002 gnd.n6864 gnd.n6822 99.6594
R7003 gnd.n6856 gnd.n6821 99.6594
R7004 gnd.n6854 gnd.n6820 99.6594
R7005 gnd.n6846 gnd.n6819 99.6594
R7006 gnd.n6844 gnd.n6818 99.6594
R7007 gnd.n6836 gnd.n6817 99.6594
R7008 gnd.n6834 gnd.n6816 99.6594
R7009 gnd.n2899 gnd.n2898 99.6594
R7010 gnd.n2658 gnd.n2636 99.6594
R7011 gnd.n2664 gnd.n2637 99.6594
R7012 gnd.n2668 gnd.n2638 99.6594
R7013 gnd.n2674 gnd.n2639 99.6594
R7014 gnd.n2678 gnd.n2640 99.6594
R7015 gnd.n2684 gnd.n2641 99.6594
R7016 gnd.n2642 gnd.n2626 99.6594
R7017 gnd.n3634 gnd.n2220 99.6594
R7018 gnd.n3638 gnd.n2221 99.6594
R7019 gnd.n3642 gnd.n2222 99.6594
R7020 gnd.n3646 gnd.n2223 99.6594
R7021 gnd.n3650 gnd.n2224 99.6594
R7022 gnd.n3654 gnd.n2225 99.6594
R7023 gnd.n3658 gnd.n2226 99.6594
R7024 gnd.n2229 gnd.n2227 99.6594
R7025 gnd.n3954 gnd.n3953 99.6594
R7026 gnd.n3948 gnd.n3748 99.6594
R7027 gnd.n3946 gnd.n3945 99.6594
R7028 gnd.n3941 gnd.n3940 99.6594
R7029 gnd.n3938 gnd.n3937 99.6594
R7030 gnd.n3933 gnd.n3932 99.6594
R7031 gnd.n3930 gnd.n3929 99.6594
R7032 gnd.n3925 gnd.n3924 99.6594
R7033 gnd.n3922 gnd.n3921 99.6594
R7034 gnd.n3917 gnd.n3916 99.6594
R7035 gnd.n3914 gnd.n3913 99.6594
R7036 gnd.n3909 gnd.n3908 99.6594
R7037 gnd.n3906 gnd.n3905 99.6594
R7038 gnd.n3901 gnd.n3900 99.6594
R7039 gnd.n3898 gnd.n3897 99.6594
R7040 gnd.n3893 gnd.n3892 99.6594
R7041 gnd.n3890 gnd.n3889 99.6594
R7042 gnd.n3885 gnd.n3884 99.6594
R7043 gnd.n3882 gnd.n3881 99.6594
R7044 gnd.n3877 gnd.n3876 99.6594
R7045 gnd.n3874 gnd.n3873 99.6594
R7046 gnd.n3869 gnd.n3868 99.6594
R7047 gnd.n3866 gnd.n3865 99.6594
R7048 gnd.n3861 gnd.n3860 99.6594
R7049 gnd.n3858 gnd.n3857 99.6594
R7050 gnd.n3853 gnd.n3852 99.6594
R7051 gnd.n3850 gnd.n3849 99.6594
R7052 gnd.n3845 gnd.n3844 99.6594
R7053 gnd.n3842 gnd.n3841 99.6594
R7054 gnd.n1076 gnd.n980 99.6594
R7055 gnd.n1080 gnd.n981 99.6594
R7056 gnd.n1084 gnd.n982 99.6594
R7057 gnd.n1088 gnd.n983 99.6594
R7058 gnd.n1092 gnd.n984 99.6594
R7059 gnd.n1096 gnd.n985 99.6594
R7060 gnd.n1100 gnd.n986 99.6594
R7061 gnd.n1104 gnd.n987 99.6594
R7062 gnd.n1108 gnd.n988 99.6594
R7063 gnd.n1112 gnd.n989 99.6594
R7064 gnd.n1118 gnd.n990 99.6594
R7065 gnd.n1122 gnd.n991 99.6594
R7066 gnd.n1126 gnd.n992 99.6594
R7067 gnd.n1130 gnd.n993 99.6594
R7068 gnd.n1134 gnd.n994 99.6594
R7069 gnd.n5754 gnd.n996 99.6594
R7070 gnd.n5758 gnd.n997 99.6594
R7071 gnd.n5762 gnd.n998 99.6594
R7072 gnd.n5766 gnd.n999 99.6594
R7073 gnd.n5771 gnd.n1000 99.6594
R7074 gnd.n5775 gnd.n1001 99.6594
R7075 gnd.n5779 gnd.n1002 99.6594
R7076 gnd.n5783 gnd.n1003 99.6594
R7077 gnd.n5787 gnd.n1004 99.6594
R7078 gnd.n5791 gnd.n1005 99.6594
R7079 gnd.n5795 gnd.n1006 99.6594
R7080 gnd.n1009 gnd.n1007 99.6594
R7081 gnd.n5801 gnd.n1008 99.6594
R7082 gnd.n5496 gnd.n1418 99.6594
R7083 gnd.n5488 gnd.n1375 99.6594
R7084 gnd.n5484 gnd.n1376 99.6594
R7085 gnd.n5480 gnd.n1377 99.6594
R7086 gnd.n5476 gnd.n1378 99.6594
R7087 gnd.n5472 gnd.n1379 99.6594
R7088 gnd.n5468 gnd.n1380 99.6594
R7089 gnd.n5464 gnd.n1381 99.6594
R7090 gnd.n5459 gnd.n1382 99.6594
R7091 gnd.n5455 gnd.n1383 99.6594
R7092 gnd.n5451 gnd.n1384 99.6594
R7093 gnd.n5447 gnd.n1385 99.6594
R7094 gnd.n5442 gnd.n1387 99.6594
R7095 gnd.n5438 gnd.n1388 99.6594
R7096 gnd.n5434 gnd.n1389 99.6594
R7097 gnd.n5430 gnd.n1390 99.6594
R7098 gnd.n5426 gnd.n1391 99.6594
R7099 gnd.n5422 gnd.n1392 99.6594
R7100 gnd.n5418 gnd.n1393 99.6594
R7101 gnd.n5414 gnd.n1394 99.6594
R7102 gnd.n5410 gnd.n1395 99.6594
R7103 gnd.n5406 gnd.n1396 99.6594
R7104 gnd.n5402 gnd.n1397 99.6594
R7105 gnd.n5398 gnd.n1398 99.6594
R7106 gnd.n5394 gnd.n1399 99.6594
R7107 gnd.n5390 gnd.n1400 99.6594
R7108 gnd.n5386 gnd.n1401 99.6594
R7109 gnd.n5378 gnd.n1402 99.6594
R7110 gnd.n6970 gnd.n6874 99.6594
R7111 gnd.n6974 gnd.n6875 99.6594
R7112 gnd.n6978 gnd.n6876 99.6594
R7113 gnd.n6982 gnd.n6877 99.6594
R7114 gnd.n6986 gnd.n6878 99.6594
R7115 gnd.n6990 gnd.n6879 99.6594
R7116 gnd.n6994 gnd.n6880 99.6594
R7117 gnd.n6998 gnd.n6881 99.6594
R7118 gnd.n7002 gnd.n6882 99.6594
R7119 gnd.n7006 gnd.n6883 99.6594
R7120 gnd.n7012 gnd.n6884 99.6594
R7121 gnd.n7016 gnd.n6885 99.6594
R7122 gnd.n7020 gnd.n6886 99.6594
R7123 gnd.n7024 gnd.n6887 99.6594
R7124 gnd.n7028 gnd.n6888 99.6594
R7125 gnd.n7032 gnd.n6889 99.6594
R7126 gnd.n7036 gnd.n6890 99.6594
R7127 gnd.n7040 gnd.n6891 99.6594
R7128 gnd.n7044 gnd.n6892 99.6594
R7129 gnd.n7048 gnd.n6893 99.6594
R7130 gnd.n7055 gnd.n6894 99.6594
R7131 gnd.n7059 gnd.n6895 99.6594
R7132 gnd.n7063 gnd.n6896 99.6594
R7133 gnd.n7067 gnd.n6897 99.6594
R7134 gnd.n7071 gnd.n6898 99.6594
R7135 gnd.n7075 gnd.n6899 99.6594
R7136 gnd.n7079 gnd.n6900 99.6594
R7137 gnd.n6903 gnd.n6901 99.6594
R7138 gnd.n7085 gnd.n6902 99.6594
R7139 gnd.n5866 gnd.n5865 99.6594
R7140 gnd.n897 gnd.n877 99.6594
R7141 gnd.n899 gnd.n878 99.6594
R7142 gnd.n903 gnd.n879 99.6594
R7143 gnd.n905 gnd.n880 99.6594
R7144 gnd.n915 gnd.n881 99.6594
R7145 gnd.n917 gnd.n882 99.6594
R7146 gnd.n925 gnd.n883 99.6594
R7147 gnd.n933 gnd.n884 99.6594
R7148 gnd.n935 gnd.n885 99.6594
R7149 gnd.n943 gnd.n886 99.6594
R7150 gnd.n951 gnd.n887 99.6594
R7151 gnd.n956 gnd.n889 99.6594
R7152 gnd.n5868 gnd.n874 99.6594
R7153 gnd.n5866 gnd.n892 99.6594
R7154 gnd.n898 gnd.n877 99.6594
R7155 gnd.n902 gnd.n878 99.6594
R7156 gnd.n904 gnd.n879 99.6594
R7157 gnd.n914 gnd.n880 99.6594
R7158 gnd.n916 gnd.n881 99.6594
R7159 gnd.n924 gnd.n882 99.6594
R7160 gnd.n932 gnd.n883 99.6594
R7161 gnd.n934 gnd.n884 99.6594
R7162 gnd.n942 gnd.n885 99.6594
R7163 gnd.n950 gnd.n886 99.6594
R7164 gnd.n952 gnd.n887 99.6594
R7165 gnd.n889 gnd.n888 99.6594
R7166 gnd.n5869 gnd.n5868 99.6594
R7167 gnd.n1637 gnd.n1313 99.6594
R7168 gnd.n1639 gnd.n1638 99.6594
R7169 gnd.n1640 gnd.n1318 99.6594
R7170 gnd.n1642 gnd.n1641 99.6594
R7171 gnd.n1643 gnd.n1324 99.6594
R7172 gnd.n1645 gnd.n1332 99.6594
R7173 gnd.n1647 gnd.n1646 99.6594
R7174 gnd.n1648 gnd.n1341 99.6594
R7175 gnd.n1650 gnd.n1348 99.6594
R7176 gnd.n1652 gnd.n1651 99.6594
R7177 gnd.n1653 gnd.n1357 99.6594
R7178 gnd.n1655 gnd.n1364 99.6594
R7179 gnd.n1658 gnd.n1657 99.6594
R7180 gnd.n5172 gnd.n5171 99.6594
R7181 gnd.n1655 gnd.n1654 99.6594
R7182 gnd.n1653 gnd.n1356 99.6594
R7183 gnd.n1652 gnd.n1349 99.6594
R7184 gnd.n1650 gnd.n1649 99.6594
R7185 gnd.n1648 gnd.n1340 99.6594
R7186 gnd.n1647 gnd.n1333 99.6594
R7187 gnd.n1645 gnd.n1644 99.6594
R7188 gnd.n1643 gnd.n1323 99.6594
R7189 gnd.n1642 gnd.n1319 99.6594
R7190 gnd.n1640 gnd.n1317 99.6594
R7191 gnd.n1639 gnd.n1314 99.6594
R7192 gnd.n1637 gnd.n1309 99.6594
R7193 gnd.n5171 gnd.n1304 99.6594
R7194 gnd.n1658 gnd.n1636 99.6594
R7195 gnd.n953 gnd.t48 98.63
R7196 gnd.n5500 gnd.t25 98.63
R7197 gnd.n960 gnd.t40 98.63
R7198 gnd.n1438 gnd.t97 98.63
R7199 gnd.n1461 gnd.t106 98.63
R7200 gnd.n5380 gnd.t70 98.63
R7201 gnd.n6965 gnd.t57 98.63
R7202 gnd.n6944 gnd.t75 98.63
R7203 gnd.n7051 gnd.t84 98.63
R7204 gnd.n6812 gnd.t20 98.63
R7205 gnd.n3772 gnd.t51 98.63
R7206 gnd.n3803 gnd.t91 98.63
R7207 gnd.n3835 gnd.t73 98.63
R7208 gnd.n3672 gnd.t37 98.63
R7209 gnd.n1030 gnd.t78 98.63
R7210 gnd.n1071 gnd.t93 98.63
R7211 gnd.n1050 gnd.t119 98.63
R7212 gnd.n1366 gnd.t32 98.63
R7213 gnd.n4436 gnd.t8 88.9408
R7214 gnd.n1791 gnd.t16 88.9408
R7215 gnd.n5683 gnd.t67 88.933
R7216 gnd.n4889 gnd.t11 88.933
R7217 gnd.n6768 gnd.n170 86.3597
R7218 gnd.n1188 gnd.n1187 81.8399
R7219 gnd.n2687 gnd.t54 74.8376
R7220 gnd.n2245 gnd.t113 74.8376
R7221 gnd.n4437 gnd.t7 72.8438
R7222 gnd.n1792 gnd.t17 72.8438
R7223 gnd.n1189 gnd.n1182 72.8411
R7224 gnd.n1195 gnd.n1180 72.8411
R7225 gnd.n4885 gnd.n4884 72.8411
R7226 gnd.n954 gnd.t47 72.836
R7227 gnd.n5684 gnd.t66 72.836
R7228 gnd.n4890 gnd.t12 72.836
R7229 gnd.n5501 gnd.t24 72.836
R7230 gnd.n961 gnd.t41 72.836
R7231 gnd.n1439 gnd.t96 72.836
R7232 gnd.n1462 gnd.t105 72.836
R7233 gnd.n5381 gnd.t69 72.836
R7234 gnd.n6966 gnd.t58 72.836
R7235 gnd.n6945 gnd.t76 72.836
R7236 gnd.n7052 gnd.t85 72.836
R7237 gnd.n6813 gnd.t21 72.836
R7238 gnd.n3773 gnd.t50 72.836
R7239 gnd.n3804 gnd.t90 72.836
R7240 gnd.n3836 gnd.t72 72.836
R7241 gnd.n3673 gnd.t36 72.836
R7242 gnd.n1031 gnd.t79 72.836
R7243 gnd.n1072 gnd.t94 72.836
R7244 gnd.n1051 gnd.t120 72.836
R7245 gnd.n1367 gnd.t33 72.836
R7246 gnd.n4953 gnd.n1757 71.676
R7247 gnd.n4949 gnd.n1758 71.676
R7248 gnd.n4945 gnd.n1759 71.676
R7249 gnd.n4941 gnd.n1760 71.676
R7250 gnd.n4937 gnd.n1761 71.676
R7251 gnd.n4933 gnd.n1762 71.676
R7252 gnd.n4929 gnd.n1763 71.676
R7253 gnd.n4925 gnd.n1764 71.676
R7254 gnd.n4921 gnd.n1765 71.676
R7255 gnd.n4917 gnd.n1766 71.676
R7256 gnd.n4913 gnd.n1767 71.676
R7257 gnd.n4909 gnd.n1768 71.676
R7258 gnd.n4905 gnd.n1769 71.676
R7259 gnd.n4901 gnd.n1770 71.676
R7260 gnd.n4896 gnd.n1771 71.676
R7261 gnd.n4892 gnd.n1772 71.676
R7262 gnd.n5029 gnd.n1790 71.676
R7263 gnd.n5025 gnd.n1789 71.676
R7264 gnd.n5020 gnd.n1788 71.676
R7265 gnd.n5016 gnd.n1787 71.676
R7266 gnd.n5012 gnd.n1786 71.676
R7267 gnd.n5008 gnd.n1785 71.676
R7268 gnd.n5004 gnd.n1784 71.676
R7269 gnd.n5000 gnd.n1783 71.676
R7270 gnd.n4996 gnd.n1782 71.676
R7271 gnd.n4992 gnd.n1781 71.676
R7272 gnd.n4988 gnd.n1780 71.676
R7273 gnd.n4984 gnd.n1779 71.676
R7274 gnd.n4980 gnd.n1778 71.676
R7275 gnd.n4976 gnd.n1777 71.676
R7276 gnd.n4972 gnd.n1776 71.676
R7277 gnd.n4968 gnd.n1775 71.676
R7278 gnd.n4964 gnd.n1774 71.676
R7279 gnd.n5747 gnd.n5746 71.676
R7280 gnd.n5741 gnd.n1144 71.676
R7281 gnd.n5738 gnd.n1145 71.676
R7282 gnd.n5734 gnd.n1146 71.676
R7283 gnd.n5730 gnd.n1147 71.676
R7284 gnd.n5726 gnd.n1148 71.676
R7285 gnd.n5722 gnd.n1149 71.676
R7286 gnd.n5718 gnd.n1150 71.676
R7287 gnd.n5714 gnd.n1151 71.676
R7288 gnd.n5710 gnd.n1152 71.676
R7289 gnd.n5706 gnd.n1153 71.676
R7290 gnd.n5702 gnd.n1154 71.676
R7291 gnd.n5698 gnd.n1155 71.676
R7292 gnd.n5694 gnd.n1156 71.676
R7293 gnd.n5690 gnd.n1157 71.676
R7294 gnd.n5686 gnd.n1158 71.676
R7295 gnd.n1159 gnd.n1142 71.676
R7296 gnd.n4440 gnd.n1160 71.676
R7297 gnd.n4445 gnd.n1161 71.676
R7298 gnd.n4449 gnd.n1162 71.676
R7299 gnd.n4453 gnd.n1163 71.676
R7300 gnd.n4457 gnd.n1164 71.676
R7301 gnd.n4461 gnd.n1165 71.676
R7302 gnd.n4465 gnd.n1166 71.676
R7303 gnd.n4469 gnd.n1167 71.676
R7304 gnd.n4473 gnd.n1168 71.676
R7305 gnd.n4477 gnd.n1169 71.676
R7306 gnd.n4481 gnd.n1170 71.676
R7307 gnd.n4485 gnd.n1171 71.676
R7308 gnd.n4489 gnd.n1172 71.676
R7309 gnd.n4493 gnd.n1173 71.676
R7310 gnd.n4497 gnd.n1174 71.676
R7311 gnd.n5747 gnd.n1177 71.676
R7312 gnd.n5739 gnd.n1144 71.676
R7313 gnd.n5735 gnd.n1145 71.676
R7314 gnd.n5731 gnd.n1146 71.676
R7315 gnd.n5727 gnd.n1147 71.676
R7316 gnd.n5723 gnd.n1148 71.676
R7317 gnd.n5719 gnd.n1149 71.676
R7318 gnd.n5715 gnd.n1150 71.676
R7319 gnd.n5711 gnd.n1151 71.676
R7320 gnd.n5707 gnd.n1152 71.676
R7321 gnd.n5703 gnd.n1153 71.676
R7322 gnd.n5699 gnd.n1154 71.676
R7323 gnd.n5695 gnd.n1155 71.676
R7324 gnd.n5691 gnd.n1156 71.676
R7325 gnd.n5687 gnd.n1157 71.676
R7326 gnd.n5750 gnd.n5749 71.676
R7327 gnd.n4439 gnd.n1159 71.676
R7328 gnd.n4444 gnd.n1160 71.676
R7329 gnd.n4448 gnd.n1161 71.676
R7330 gnd.n4452 gnd.n1162 71.676
R7331 gnd.n4456 gnd.n1163 71.676
R7332 gnd.n4460 gnd.n1164 71.676
R7333 gnd.n4464 gnd.n1165 71.676
R7334 gnd.n4468 gnd.n1166 71.676
R7335 gnd.n4472 gnd.n1167 71.676
R7336 gnd.n4476 gnd.n1168 71.676
R7337 gnd.n4480 gnd.n1169 71.676
R7338 gnd.n4484 gnd.n1170 71.676
R7339 gnd.n4488 gnd.n1171 71.676
R7340 gnd.n4492 gnd.n1172 71.676
R7341 gnd.n4496 gnd.n1173 71.676
R7342 gnd.n4500 gnd.n1174 71.676
R7343 gnd.n4967 gnd.n1774 71.676
R7344 gnd.n4971 gnd.n1775 71.676
R7345 gnd.n4975 gnd.n1776 71.676
R7346 gnd.n4979 gnd.n1777 71.676
R7347 gnd.n4983 gnd.n1778 71.676
R7348 gnd.n4987 gnd.n1779 71.676
R7349 gnd.n4991 gnd.n1780 71.676
R7350 gnd.n4995 gnd.n1781 71.676
R7351 gnd.n4999 gnd.n1782 71.676
R7352 gnd.n5003 gnd.n1783 71.676
R7353 gnd.n5007 gnd.n1784 71.676
R7354 gnd.n5011 gnd.n1785 71.676
R7355 gnd.n5015 gnd.n1786 71.676
R7356 gnd.n5019 gnd.n1787 71.676
R7357 gnd.n5024 gnd.n1788 71.676
R7358 gnd.n5028 gnd.n1789 71.676
R7359 gnd.n4891 gnd.n1773 71.676
R7360 gnd.n4895 gnd.n1772 71.676
R7361 gnd.n4900 gnd.n1771 71.676
R7362 gnd.n4904 gnd.n1770 71.676
R7363 gnd.n4908 gnd.n1769 71.676
R7364 gnd.n4912 gnd.n1768 71.676
R7365 gnd.n4916 gnd.n1767 71.676
R7366 gnd.n4920 gnd.n1766 71.676
R7367 gnd.n4924 gnd.n1765 71.676
R7368 gnd.n4928 gnd.n1764 71.676
R7369 gnd.n4932 gnd.n1763 71.676
R7370 gnd.n4936 gnd.n1762 71.676
R7371 gnd.n4940 gnd.n1761 71.676
R7372 gnd.n4944 gnd.n1760 71.676
R7373 gnd.n4948 gnd.n1759 71.676
R7374 gnd.n4952 gnd.n1758 71.676
R7375 gnd.n4955 gnd.n1757 71.676
R7376 gnd.n10 gnd.t322 69.1507
R7377 gnd.n18 gnd.t195 68.4792
R7378 gnd.n17 gnd.t326 68.4792
R7379 gnd.n16 gnd.t180 68.4792
R7380 gnd.n15 gnd.t189 68.4792
R7381 gnd.n14 gnd.t142 68.4792
R7382 gnd.n13 gnd.t324 68.4792
R7383 gnd.n12 gnd.t174 68.4792
R7384 gnd.n11 gnd.t161 68.4792
R7385 gnd.n10 gnd.t320 68.4792
R7386 gnd.n2814 gnd.n2718 64.369
R7387 gnd.n3961 gnd.n3667 63.0944
R7388 gnd.n4442 gnd.n4437 59.5399
R7389 gnd.n5022 gnd.n1792 59.5399
R7390 gnd.n5685 gnd.n5684 59.5399
R7391 gnd.n4898 gnd.n4890 59.5399
R7392 gnd.n5682 gnd.n1198 59.1804
R7393 gnd.n3666 gnd.n2205 57.3586
R7394 gnd.n2473 gnd.t290 56.407
R7395 gnd.n2438 gnd.t304 56.407
R7396 gnd.n2449 gnd.t276 56.407
R7397 gnd.n2461 gnd.t212 56.407
R7398 gnd.n56 gnd.t270 56.407
R7399 gnd.n21 gnd.t218 56.407
R7400 gnd.n32 gnd.t257 56.407
R7401 gnd.n44 gnd.t298 56.407
R7402 gnd.n2482 gnd.t230 55.8337
R7403 gnd.n2447 gnd.t300 55.8337
R7404 gnd.n2458 gnd.t268 55.8337
R7405 gnd.n2470 gnd.t281 55.8337
R7406 gnd.n65 gnd.t306 55.8337
R7407 gnd.n30 gnd.t204 55.8337
R7408 gnd.n41 gnd.t203 55.8337
R7409 gnd.n53 gnd.t248 55.8337
R7410 gnd.n7086 gnd.n170 55.7653
R7411 gnd.n1186 gnd.n1185 54.358
R7412 gnd.n4882 gnd.n4881 54.358
R7413 gnd.n2473 gnd.n2472 53.0052
R7414 gnd.n2475 gnd.n2474 53.0052
R7415 gnd.n2477 gnd.n2476 53.0052
R7416 gnd.n2479 gnd.n2478 53.0052
R7417 gnd.n2481 gnd.n2480 53.0052
R7418 gnd.n2438 gnd.n2437 53.0052
R7419 gnd.n2440 gnd.n2439 53.0052
R7420 gnd.n2442 gnd.n2441 53.0052
R7421 gnd.n2444 gnd.n2443 53.0052
R7422 gnd.n2446 gnd.n2445 53.0052
R7423 gnd.n2449 gnd.n2448 53.0052
R7424 gnd.n2451 gnd.n2450 53.0052
R7425 gnd.n2453 gnd.n2452 53.0052
R7426 gnd.n2455 gnd.n2454 53.0052
R7427 gnd.n2457 gnd.n2456 53.0052
R7428 gnd.n2461 gnd.n2460 53.0052
R7429 gnd.n2463 gnd.n2462 53.0052
R7430 gnd.n2465 gnd.n2464 53.0052
R7431 gnd.n2467 gnd.n2466 53.0052
R7432 gnd.n2469 gnd.n2468 53.0052
R7433 gnd.n64 gnd.n63 53.0052
R7434 gnd.n62 gnd.n61 53.0052
R7435 gnd.n60 gnd.n59 53.0052
R7436 gnd.n58 gnd.n57 53.0052
R7437 gnd.n56 gnd.n55 53.0052
R7438 gnd.n29 gnd.n28 53.0052
R7439 gnd.n27 gnd.n26 53.0052
R7440 gnd.n25 gnd.n24 53.0052
R7441 gnd.n23 gnd.n22 53.0052
R7442 gnd.n21 gnd.n20 53.0052
R7443 gnd.n40 gnd.n39 53.0052
R7444 gnd.n38 gnd.n37 53.0052
R7445 gnd.n36 gnd.n35 53.0052
R7446 gnd.n34 gnd.n33 53.0052
R7447 gnd.n32 gnd.n31 53.0052
R7448 gnd.n52 gnd.n51 53.0052
R7449 gnd.n50 gnd.n49 53.0052
R7450 gnd.n48 gnd.n47 53.0052
R7451 gnd.n46 gnd.n45 53.0052
R7452 gnd.n44 gnd.n43 53.0052
R7453 gnd.n4873 gnd.n4872 52.4801
R7454 gnd.n3518 gnd.t154 52.3082
R7455 gnd.n3486 gnd.t182 52.3082
R7456 gnd.n3454 gnd.t170 52.3082
R7457 gnd.n3423 gnd.t134 52.3082
R7458 gnd.n3391 gnd.t167 52.3082
R7459 gnd.n3359 gnd.t178 52.3082
R7460 gnd.n3327 gnd.t149 52.3082
R7461 gnd.n3296 gnd.t159 52.3082
R7462 gnd.n3348 gnd.n3316 51.4173
R7463 gnd.n3412 gnd.n3411 50.455
R7464 gnd.n3380 gnd.n3379 50.455
R7465 gnd.n3348 gnd.n3347 50.455
R7466 gnd.n2761 gnd.n2760 45.1884
R7467 gnd.n2271 gnd.n2270 45.1884
R7468 gnd.n4957 gnd.n4888 44.3322
R7469 gnd.n1189 gnd.n1188 44.3189
R7470 gnd.n955 gnd.n954 42.4732
R7471 gnd.n1368 gnd.n1367 42.4732
R7472 gnd.n5502 gnd.n5501 42.2793
R7473 gnd.n2762 gnd.n2761 42.2793
R7474 gnd.n2272 gnd.n2271 42.2793
R7475 gnd.n2688 gnd.n2687 42.2793
R7476 gnd.n3633 gnd.n2245 42.2793
R7477 gnd.n5806 gnd.n961 42.2793
R7478 gnd.n5461 gnd.n1439 42.2793
R7479 gnd.n5424 gnd.n1462 42.2793
R7480 gnd.n5384 gnd.n5381 42.2793
R7481 gnd.n6969 gnd.n6966 42.2793
R7482 gnd.n7011 gnd.n6945 42.2793
R7483 gnd.n7053 gnd.n7052 42.2793
R7484 gnd.n6814 gnd.n6813 42.2793
R7485 gnd.n3774 gnd.n3773 42.2793
R7486 gnd.n3805 gnd.n3804 42.2793
R7487 gnd.n3837 gnd.n3836 42.2793
R7488 gnd.n3674 gnd.n3673 42.2793
R7489 gnd.n5769 gnd.n1031 42.2793
R7490 gnd.n1075 gnd.n1072 42.2793
R7491 gnd.n1117 gnd.n1051 42.2793
R7492 gnd.n1187 gnd.n1186 41.6274
R7493 gnd.n4883 gnd.n4882 41.6274
R7494 gnd.n1196 gnd.n1195 40.8975
R7495 gnd.n4886 gnd.n4885 40.8975
R7496 gnd.n6137 gnd.n561 37.8532
R7497 gnd.n6137 gnd.n6136 37.8532
R7498 gnd.n6136 gnd.n6135 37.8532
R7499 gnd.n6135 gnd.n566 37.8532
R7500 gnd.n6129 gnd.n566 37.8532
R7501 gnd.n6129 gnd.n6128 37.8532
R7502 gnd.n6128 gnd.n6127 37.8532
R7503 gnd.n6127 gnd.n574 37.8532
R7504 gnd.n6121 gnd.n574 37.8532
R7505 gnd.n6121 gnd.n6120 37.8532
R7506 gnd.n6120 gnd.n6119 37.8532
R7507 gnd.n6119 gnd.n582 37.8532
R7508 gnd.n6113 gnd.n582 37.8532
R7509 gnd.n6113 gnd.n6112 37.8532
R7510 gnd.n6112 gnd.n6111 37.8532
R7511 gnd.n6111 gnd.n590 37.8532
R7512 gnd.n6105 gnd.n590 37.8532
R7513 gnd.n6105 gnd.n6104 37.8532
R7514 gnd.n6104 gnd.n6103 37.8532
R7515 gnd.n6103 gnd.n598 37.8532
R7516 gnd.n6097 gnd.n598 37.8532
R7517 gnd.n6097 gnd.n6096 37.8532
R7518 gnd.n6096 gnd.n6095 37.8532
R7519 gnd.n6095 gnd.n606 37.8532
R7520 gnd.n6089 gnd.n606 37.8532
R7521 gnd.n6089 gnd.n6088 37.8532
R7522 gnd.n6088 gnd.n6087 37.8532
R7523 gnd.n6087 gnd.n614 37.8532
R7524 gnd.n6081 gnd.n614 37.8532
R7525 gnd.n6081 gnd.n6080 37.8532
R7526 gnd.n6080 gnd.n6079 37.8532
R7527 gnd.n6079 gnd.n622 37.8532
R7528 gnd.n6073 gnd.n622 37.8532
R7529 gnd.n6073 gnd.n6072 37.8532
R7530 gnd.n6072 gnd.n6071 37.8532
R7531 gnd.n6071 gnd.n630 37.8532
R7532 gnd.n6065 gnd.n630 37.8532
R7533 gnd.n6065 gnd.n6064 37.8532
R7534 gnd.n6064 gnd.n6063 37.8532
R7535 gnd.n6063 gnd.n638 37.8532
R7536 gnd.n6057 gnd.n638 37.8532
R7537 gnd.n6057 gnd.n6056 37.8532
R7538 gnd.n6056 gnd.n6055 37.8532
R7539 gnd.n6055 gnd.n646 37.8532
R7540 gnd.n6049 gnd.n646 37.8532
R7541 gnd.n6049 gnd.n6048 37.8532
R7542 gnd.n6048 gnd.n6047 37.8532
R7543 gnd.n6047 gnd.n654 37.8532
R7544 gnd.n6041 gnd.n654 37.8532
R7545 gnd.n6041 gnd.n6040 37.8532
R7546 gnd.n6040 gnd.n6039 37.8532
R7547 gnd.n6039 gnd.n662 37.8532
R7548 gnd.n6033 gnd.n662 37.8532
R7549 gnd.n6033 gnd.n6032 37.8532
R7550 gnd.n6032 gnd.n6031 37.8532
R7551 gnd.n6031 gnd.n670 37.8532
R7552 gnd.n6025 gnd.n670 37.8532
R7553 gnd.n6025 gnd.n6024 37.8532
R7554 gnd.n6024 gnd.n6023 37.8532
R7555 gnd.n6023 gnd.n678 37.8532
R7556 gnd.n6017 gnd.n678 37.8532
R7557 gnd.n6017 gnd.n6016 37.8532
R7558 gnd.n6016 gnd.n6015 37.8532
R7559 gnd.n6015 gnd.n686 37.8532
R7560 gnd.n6009 gnd.n686 37.8532
R7561 gnd.n6009 gnd.n6008 37.8532
R7562 gnd.n6008 gnd.n6007 37.8532
R7563 gnd.n6007 gnd.n694 37.8532
R7564 gnd.n6001 gnd.n694 37.8532
R7565 gnd.n6001 gnd.n6000 37.8532
R7566 gnd.n6000 gnd.n5999 37.8532
R7567 gnd.n5999 gnd.n702 37.8532
R7568 gnd.n5993 gnd.n702 37.8532
R7569 gnd.n5993 gnd.n5992 37.8532
R7570 gnd.n5992 gnd.n5991 37.8532
R7571 gnd.n5991 gnd.n710 37.8532
R7572 gnd.n5985 gnd.n710 37.8532
R7573 gnd.n5985 gnd.n5984 37.8532
R7574 gnd.n5984 gnd.n5983 37.8532
R7575 gnd.n5983 gnd.n718 37.8532
R7576 gnd.n5977 gnd.n718 37.8532
R7577 gnd.n5977 gnd.n5976 37.8532
R7578 gnd.n5976 gnd.n5975 37.8532
R7579 gnd.n1195 gnd.n1194 35.055
R7580 gnd.n1190 gnd.n1189 35.055
R7581 gnd.n4875 gnd.n4874 35.055
R7582 gnd.n4885 gnd.n4871 35.055
R7583 gnd.n4965 gnd.n1793 32.3127
R7584 gnd.n4502 gnd.n4499 32.3127
R7585 gnd.n2824 gnd.n2718 31.8661
R7586 gnd.n2824 gnd.n2823 31.8661
R7587 gnd.n2832 gnd.n2707 31.8661
R7588 gnd.n2840 gnd.n2707 31.8661
R7589 gnd.n2840 gnd.n2701 31.8661
R7590 gnd.n2848 gnd.n2701 31.8661
R7591 gnd.n2848 gnd.n2694 31.8661
R7592 gnd.n2886 gnd.n2694 31.8661
R7593 gnd.n2896 gnd.n2627 31.8661
R7594 gnd.n3961 gnd.n3744 31.8661
R7595 gnd.n3979 gnd.n2185 31.8661
R7596 gnd.n3989 gnd.n2185 31.8661
R7597 gnd.n3989 gnd.n2179 31.8661
R7598 gnd.n3999 gnd.n2179 31.8661
R7599 gnd.n4014 gnd.n2160 31.8661
R7600 gnd.n4024 gnd.n2160 31.8661
R7601 gnd.n4036 gnd.n2154 31.8661
R7602 gnd.n4054 gnd.n2144 31.8661
R7603 gnd.n965 gnd.n862 31.8661
R7604 gnd.n4219 gnd.n979 31.8661
R7605 gnd.n4219 gnd.n876 31.8661
R7606 gnd.n4228 gnd.n890 31.8661
R7607 gnd.n4304 gnd.n4228 31.8661
R7608 gnd.n4312 gnd.n2075 31.8661
R7609 gnd.n4312 gnd.n2067 31.8661
R7610 gnd.n4320 gnd.n2067 31.8661
R7611 gnd.n4320 gnd.n2069 31.8661
R7612 gnd.n4328 gnd.n2054 31.8661
R7613 gnd.n4336 gnd.n2054 31.8661
R7614 gnd.n4336 gnd.n2047 31.8661
R7615 gnd.n4344 gnd.n2047 31.8661
R7616 gnd.n4352 gnd.n2040 31.8661
R7617 gnd.n4352 gnd.n2033 31.8661
R7618 gnd.n4360 gnd.n2033 31.8661
R7619 gnd.n4368 gnd.n2026 31.8661
R7620 gnd.n4368 gnd.n2018 31.8661
R7621 gnd.n4376 gnd.n2018 31.8661
R7622 gnd.n4376 gnd.n2020 31.8661
R7623 gnd.n4384 gnd.n2005 31.8661
R7624 gnd.n4392 gnd.n2005 31.8661
R7625 gnd.n4392 gnd.n1997 31.8661
R7626 gnd.n4401 gnd.n1997 31.8661
R7627 gnd.n4415 gnd.n1989 31.8661
R7628 gnd.n4415 gnd.n1143 31.8661
R7629 gnd.n5040 gnd.n1744 31.8661
R7630 gnd.n5048 gnd.n1744 31.8661
R7631 gnd.n5056 gnd.n1737 31.8661
R7632 gnd.n5056 gnd.n1731 31.8661
R7633 gnd.n5065 gnd.n1731 31.8661
R7634 gnd.n5065 gnd.n5064 31.8661
R7635 gnd.n5073 gnd.n1719 31.8661
R7636 gnd.n5081 gnd.n1719 31.8661
R7637 gnd.n5081 gnd.n1712 31.8661
R7638 gnd.n5089 gnd.n1712 31.8661
R7639 gnd.n5097 gnd.n1706 31.8661
R7640 gnd.n5097 gnd.n1699 31.8661
R7641 gnd.n5105 gnd.n1699 31.8661
R7642 gnd.n5113 gnd.n1693 31.8661
R7643 gnd.n5113 gnd.n1684 31.8661
R7644 gnd.n5121 gnd.n1684 31.8661
R7645 gnd.n5121 gnd.n1686 31.8661
R7646 gnd.n5129 gnd.n1673 31.8661
R7647 gnd.n5140 gnd.n1673 31.8661
R7648 gnd.n5140 gnd.n1667 31.8661
R7649 gnd.n5148 gnd.n1667 31.8661
R7650 gnd.n5565 gnd.n1305 31.8661
R7651 gnd.n5565 gnd.n1307 31.8661
R7652 gnd.n5169 gnd.n1659 31.8661
R7653 gnd.n1659 gnd.n1374 31.8661
R7654 gnd.n1484 gnd.n1416 31.8661
R7655 gnd.n7183 gnd.n111 31.8661
R7656 gnd.n7177 gnd.n120 31.8661
R7657 gnd.n7171 gnd.n130 31.8661
R7658 gnd.n7171 gnd.n133 31.8661
R7659 gnd.n7165 gnd.n142 31.8661
R7660 gnd.n7159 gnd.n142 31.8661
R7661 gnd.n7159 gnd.n152 31.8661
R7662 gnd.n7153 gnd.n152 31.8661
R7663 gnd.n7147 gnd.n167 31.8661
R7664 gnd.t198 gnd.n2154 30.9101
R7665 gnd.n7177 gnd.t223 30.9101
R7666 gnd.t0 gnd.n1989 28.9982
R7667 gnd.n5048 gnd.t179 28.9982
R7668 gnd.n4360 gnd.t164 27.0862
R7669 gnd.t325 gnd.n1706 27.0862
R7670 gnd.n5748 gnd.n1143 25.8116
R7671 gnd.n954 gnd.n953 25.7944
R7672 gnd.n5501 gnd.n5500 25.7944
R7673 gnd.n2687 gnd.n2686 25.7944
R7674 gnd.n2245 gnd.n2244 25.7944
R7675 gnd.n961 gnd.n960 25.7944
R7676 gnd.n1439 gnd.n1438 25.7944
R7677 gnd.n1462 gnd.n1461 25.7944
R7678 gnd.n5381 gnd.n5380 25.7944
R7679 gnd.n6966 gnd.n6965 25.7944
R7680 gnd.n6945 gnd.n6944 25.7944
R7681 gnd.n7052 gnd.n7051 25.7944
R7682 gnd.n6813 gnd.n6812 25.7944
R7683 gnd.n3773 gnd.n3772 25.7944
R7684 gnd.n3804 gnd.n3803 25.7944
R7685 gnd.n3836 gnd.n3835 25.7944
R7686 gnd.n3673 gnd.n3672 25.7944
R7687 gnd.n1031 gnd.n1030 25.7944
R7688 gnd.n1072 gnd.n1071 25.7944
R7689 gnd.n1051 gnd.n1050 25.7944
R7690 gnd.n1367 gnd.n1366 25.7944
R7691 gnd.n2908 gnd.n2628 24.8557
R7692 gnd.n2918 gnd.n2611 24.8557
R7693 gnd.n2614 gnd.n2602 24.8557
R7694 gnd.n2939 gnd.n2603 24.8557
R7695 gnd.n2949 gnd.n2583 24.8557
R7696 gnd.n2959 gnd.n2958 24.8557
R7697 gnd.n2569 gnd.n2567 24.8557
R7698 gnd.n2990 gnd.n2989 24.8557
R7699 gnd.n3005 gnd.n2552 24.8557
R7700 gnd.n3059 gnd.n2491 24.8557
R7701 gnd.n3015 gnd.n2492 24.8557
R7702 gnd.n3052 gnd.n2503 24.8557
R7703 gnd.n2541 gnd.n2540 24.8557
R7704 gnd.n3046 gnd.n3045 24.8557
R7705 gnd.n2527 gnd.n2514 24.8557
R7706 gnd.n3085 gnd.n3084 24.8557
R7707 gnd.n3095 gnd.n2423 24.8557
R7708 gnd.n3107 gnd.n2415 24.8557
R7709 gnd.n3106 gnd.n2403 24.8557
R7710 gnd.n3125 gnd.n3124 24.8557
R7711 gnd.n3135 gnd.n2396 24.8557
R7712 gnd.n3146 gnd.n2384 24.8557
R7713 gnd.n3170 gnd.n3169 24.8557
R7714 gnd.n3181 gnd.n2367 24.8557
R7715 gnd.n3180 gnd.n2369 24.8557
R7716 gnd.n3192 gnd.n2360 24.8557
R7717 gnd.n3210 gnd.n3209 24.8557
R7718 gnd.n2351 gnd.n2340 24.8557
R7719 gnd.n3231 gnd.n2328 24.8557
R7720 gnd.n3259 gnd.n3258 24.8557
R7721 gnd.n3270 gnd.n2313 24.8557
R7722 gnd.n3281 gnd.n2306 24.8557
R7723 gnd.n3280 gnd.n2294 24.8557
R7724 gnd.n3553 gnd.n3552 24.8557
R7725 gnd.n3575 gnd.n2279 24.8557
R7726 gnd.n4304 gnd.t46 24.537
R7727 gnd.t321 gnd.n2040 24.537
R7728 gnd.n5105 gnd.t192 24.537
R7729 gnd.t31 gnd.n1305 24.537
R7730 gnd.n5867 gnd.n890 23.8997
R7731 gnd.n5170 gnd.n1307 23.8997
R7732 gnd.n2929 gnd.t158 23.2624
R7733 gnd.n5975 gnd.n726 22.7121
R7734 gnd.n2630 gnd.t53 22.6251
R7735 gnd.t160 gnd.n1175 22.6251
R7736 gnd.t151 gnd.n5031 22.6251
R7737 gnd.n4036 gnd.t236 21.9878
R7738 gnd.n120 gnd.t215 21.9878
R7739 gnd.n5678 gnd.n1201 21.6691
R7740 gnd.n4529 gnd.n1213 21.6691
R7741 gnd.n4601 gnd.n1943 21.6691
R7742 gnd.n4688 gnd.n1903 21.6691
R7743 gnd.n4696 gnd.n4695 21.6691
R7744 gnd.n4716 gnd.n1888 21.6691
R7745 gnd.n4722 gnd.n1884 21.6691
R7746 gnd.n4813 gnd.n1844 21.6691
R7747 gnd.n4838 gnd.n1823 21.6691
R7748 gnd.n4866 gnd.n1802 21.6691
R7749 gnd.t133 gnd.n2635 21.3504
R7750 gnd.n4595 gnd.n1949 21.0318
R7751 gnd.n4588 gnd.n1932 21.0318
R7752 gnd.n4744 gnd.n1852 21.0318
R7753 gnd.n4761 gnd.n4760 21.0318
R7754 gnd.n5040 gnd.t43 21.0318
R7755 gnd.t121 gnd.n2341 20.7131
R7756 gnd.n2144 gnd.n2134 20.7131
R7757 gnd.t251 gnd.n733 20.7131
R7758 gnd.n7116 gnd.t209 20.7131
R7759 gnd.n111 gnd.n104 20.7131
R7760 gnd.n5682 gnd.n5681 20.1371
R7761 gnd.n4958 gnd.n4957 20.1371
R7762 gnd.t131 gnd.n2376 20.0758
R7763 gnd.n4014 gnd.t229 20.0758
R7764 gnd.t202 gnd.n133 20.0758
R7765 gnd.n1184 gnd.t88 19.8005
R7766 gnd.n1184 gnd.t14 19.8005
R7767 gnd.n1183 gnd.t64 19.8005
R7768 gnd.n1183 gnd.t109 19.8005
R7769 gnd.n4880 gnd.t4 19.8005
R7770 gnd.n4880 gnd.t82 19.8005
R7771 gnd.n4879 gnd.t100 19.8005
R7772 gnd.n4879 gnd.t44 19.8005
R7773 gnd.n5802 gnd.n979 19.7572
R7774 gnd.n4538 gnd.n1940 19.7572
R7775 gnd.n4662 gnd.n1919 19.7572
R7776 gnd.n1870 gnd.n1859 19.7572
R7777 gnd.n4821 gnd.n1838 19.7572
R7778 gnd.n5497 gnd.n1374 19.7572
R7779 gnd.n1180 gnd.n1179 19.5087
R7780 gnd.n1193 gnd.n1180 19.5087
R7781 gnd.n1191 gnd.n1182 19.5087
R7782 gnd.n4884 gnd.n4878 19.5087
R7783 gnd.n3096 gnd.t168 19.4385
R7784 gnd.n2069 gnd.t171 19.4385
R7785 gnd.n5129 gnd.t194 19.4385
R7786 gnd.n4302 gnd.n4299 19.3944
R7787 gnd.n4302 gnd.n2073 19.3944
R7788 gnd.n4314 gnd.n2073 19.3944
R7789 gnd.n4314 gnd.n2071 19.3944
R7790 gnd.n4318 gnd.n2071 19.3944
R7791 gnd.n4318 gnd.n2059 19.3944
R7792 gnd.n4330 gnd.n2059 19.3944
R7793 gnd.n4330 gnd.n2057 19.3944
R7794 gnd.n4334 gnd.n2057 19.3944
R7795 gnd.n4334 gnd.n2045 19.3944
R7796 gnd.n4346 gnd.n2045 19.3944
R7797 gnd.n4346 gnd.n2043 19.3944
R7798 gnd.n4350 gnd.n2043 19.3944
R7799 gnd.n4350 gnd.n2031 19.3944
R7800 gnd.n4362 gnd.n2031 19.3944
R7801 gnd.n4362 gnd.n2029 19.3944
R7802 gnd.n4366 gnd.n2029 19.3944
R7803 gnd.n4366 gnd.n2016 19.3944
R7804 gnd.n4378 gnd.n2016 19.3944
R7805 gnd.n4378 gnd.n2014 19.3944
R7806 gnd.n4382 gnd.n2014 19.3944
R7807 gnd.n4382 gnd.n2003 19.3944
R7808 gnd.n4394 gnd.n2003 19.3944
R7809 gnd.n4394 gnd.n2000 19.3944
R7810 gnd.n4399 gnd.n2000 19.3944
R7811 gnd.n4399 gnd.n2001 19.3944
R7812 gnd.n2001 gnd.n1987 19.3944
R7813 gnd.n4418 gnd.n1987 19.3944
R7814 gnd.n4418 gnd.n1984 19.3944
R7815 gnd.n4423 gnd.n1984 19.3944
R7816 gnd.n4423 gnd.n1985 19.3944
R7817 gnd.n1985 gnd.n1217 19.3944
R7818 gnd.n5669 gnd.n1217 19.3944
R7819 gnd.n5669 gnd.n1218 19.3944
R7820 gnd.n5665 gnd.n1218 19.3944
R7821 gnd.n5665 gnd.n5664 19.3944
R7822 gnd.n5664 gnd.n5663 19.3944
R7823 gnd.n5663 gnd.n1224 19.3944
R7824 gnd.n5659 gnd.n1224 19.3944
R7825 gnd.n5659 gnd.n5658 19.3944
R7826 gnd.n5658 gnd.n5657 19.3944
R7827 gnd.n5657 gnd.n1229 19.3944
R7828 gnd.n5653 gnd.n1229 19.3944
R7829 gnd.n5653 gnd.n5652 19.3944
R7830 gnd.n5652 gnd.n5651 19.3944
R7831 gnd.n5651 gnd.n1234 19.3944
R7832 gnd.n5647 gnd.n1234 19.3944
R7833 gnd.n5647 gnd.n5646 19.3944
R7834 gnd.n5646 gnd.n5645 19.3944
R7835 gnd.n5645 gnd.n1239 19.3944
R7836 gnd.n5641 gnd.n1239 19.3944
R7837 gnd.n5641 gnd.n5640 19.3944
R7838 gnd.n5640 gnd.n5639 19.3944
R7839 gnd.n5639 gnd.n1244 19.3944
R7840 gnd.n5635 gnd.n1244 19.3944
R7841 gnd.n5635 gnd.n5634 19.3944
R7842 gnd.n5634 gnd.n5633 19.3944
R7843 gnd.n5633 gnd.n1249 19.3944
R7844 gnd.n5629 gnd.n1249 19.3944
R7845 gnd.n5629 gnd.n5628 19.3944
R7846 gnd.n5628 gnd.n5627 19.3944
R7847 gnd.n5627 gnd.n1254 19.3944
R7848 gnd.n5623 gnd.n1254 19.3944
R7849 gnd.n5623 gnd.n5622 19.3944
R7850 gnd.n5622 gnd.n5621 19.3944
R7851 gnd.n5621 gnd.n1259 19.3944
R7852 gnd.n5617 gnd.n1259 19.3944
R7853 gnd.n5617 gnd.n5616 19.3944
R7854 gnd.n5616 gnd.n5615 19.3944
R7855 gnd.n5615 gnd.n1264 19.3944
R7856 gnd.n5611 gnd.n1264 19.3944
R7857 gnd.n5611 gnd.n5610 19.3944
R7858 gnd.n5610 gnd.n5609 19.3944
R7859 gnd.n5609 gnd.n1269 19.3944
R7860 gnd.n5605 gnd.n1269 19.3944
R7861 gnd.n5605 gnd.n5604 19.3944
R7862 gnd.n5604 gnd.n5603 19.3944
R7863 gnd.n5603 gnd.n1274 19.3944
R7864 gnd.n5599 gnd.n1274 19.3944
R7865 gnd.n5599 gnd.n5598 19.3944
R7866 gnd.n5598 gnd.n5597 19.3944
R7867 gnd.n5597 gnd.n1279 19.3944
R7868 gnd.n5593 gnd.n1279 19.3944
R7869 gnd.n5593 gnd.n5592 19.3944
R7870 gnd.n5592 gnd.n5591 19.3944
R7871 gnd.n5591 gnd.n1284 19.3944
R7872 gnd.n5587 gnd.n1284 19.3944
R7873 gnd.n5587 gnd.n5586 19.3944
R7874 gnd.n5586 gnd.n5585 19.3944
R7875 gnd.n5585 gnd.n1289 19.3944
R7876 gnd.n5581 gnd.n1289 19.3944
R7877 gnd.n5581 gnd.n5580 19.3944
R7878 gnd.n5580 gnd.n5579 19.3944
R7879 gnd.n5579 gnd.n1294 19.3944
R7880 gnd.n5575 gnd.n1294 19.3944
R7881 gnd.n5575 gnd.n5574 19.3944
R7882 gnd.n5574 gnd.n5573 19.3944
R7883 gnd.n5573 gnd.n1299 19.3944
R7884 gnd.n5569 gnd.n1299 19.3944
R7885 gnd.n5569 gnd.n5568 19.3944
R7886 gnd.n5568 gnd.n5567 19.3944
R7887 gnd.n957 gnd.n873 19.3944
R7888 gnd.n5871 gnd.n873 19.3944
R7889 gnd.n5871 gnd.n5870 19.3944
R7890 gnd.n5864 gnd.n5863 19.3944
R7891 gnd.n5863 gnd.n895 19.3944
R7892 gnd.n5859 gnd.n895 19.3944
R7893 gnd.n5859 gnd.n5858 19.3944
R7894 gnd.n5858 gnd.n5857 19.3944
R7895 gnd.n5857 gnd.n900 19.3944
R7896 gnd.n5852 gnd.n900 19.3944
R7897 gnd.n5852 gnd.n5851 19.3944
R7898 gnd.n5851 gnd.n5850 19.3944
R7899 gnd.n5850 gnd.n906 19.3944
R7900 gnd.n5843 gnd.n906 19.3944
R7901 gnd.n5843 gnd.n5842 19.3944
R7902 gnd.n5842 gnd.n918 19.3944
R7903 gnd.n5835 gnd.n918 19.3944
R7904 gnd.n5835 gnd.n5834 19.3944
R7905 gnd.n5834 gnd.n926 19.3944
R7906 gnd.n5827 gnd.n926 19.3944
R7907 gnd.n5827 gnd.n5826 19.3944
R7908 gnd.n5826 gnd.n936 19.3944
R7909 gnd.n5819 gnd.n936 19.3944
R7910 gnd.n5819 gnd.n5818 19.3944
R7911 gnd.n5818 gnd.n944 19.3944
R7912 gnd.n5811 gnd.n944 19.3944
R7913 gnd.n5811 gnd.n5810 19.3944
R7914 gnd.n5543 gnd.n1327 19.3944
R7915 gnd.n5543 gnd.n5542 19.3944
R7916 gnd.n5542 gnd.n1330 19.3944
R7917 gnd.n5535 gnd.n1330 19.3944
R7918 gnd.n5535 gnd.n5534 19.3944
R7919 gnd.n5534 gnd.n1338 19.3944
R7920 gnd.n5527 gnd.n1338 19.3944
R7921 gnd.n5527 gnd.n5526 19.3944
R7922 gnd.n5526 gnd.n1346 19.3944
R7923 gnd.n5519 gnd.n1346 19.3944
R7924 gnd.n5519 gnd.n5518 19.3944
R7925 gnd.n5518 gnd.n1354 19.3944
R7926 gnd.n5511 gnd.n1354 19.3944
R7927 gnd.n5511 gnd.n5510 19.3944
R7928 gnd.n5510 gnd.n1362 19.3944
R7929 gnd.n5503 gnd.n1362 19.3944
R7930 gnd.n2811 gnd.n2810 19.3944
R7931 gnd.n2810 gnd.n2809 19.3944
R7932 gnd.n2809 gnd.n2808 19.3944
R7933 gnd.n2808 gnd.n2806 19.3944
R7934 gnd.n2806 gnd.n2803 19.3944
R7935 gnd.n2803 gnd.n2802 19.3944
R7936 gnd.n2802 gnd.n2799 19.3944
R7937 gnd.n2799 gnd.n2798 19.3944
R7938 gnd.n2798 gnd.n2795 19.3944
R7939 gnd.n2795 gnd.n2794 19.3944
R7940 gnd.n2794 gnd.n2791 19.3944
R7941 gnd.n2791 gnd.n2790 19.3944
R7942 gnd.n2790 gnd.n2787 19.3944
R7943 gnd.n2787 gnd.n2786 19.3944
R7944 gnd.n2786 gnd.n2783 19.3944
R7945 gnd.n2783 gnd.n2782 19.3944
R7946 gnd.n2782 gnd.n2779 19.3944
R7947 gnd.n2779 gnd.n2778 19.3944
R7948 gnd.n2778 gnd.n2775 19.3944
R7949 gnd.n2775 gnd.n2774 19.3944
R7950 gnd.n2774 gnd.n2771 19.3944
R7951 gnd.n2771 gnd.n2770 19.3944
R7952 gnd.n2767 gnd.n2766 19.3944
R7953 gnd.n2766 gnd.n2722 19.3944
R7954 gnd.n2817 gnd.n2722 19.3944
R7955 gnd.n3583 gnd.n3582 19.3944
R7956 gnd.n3582 gnd.n3579 19.3944
R7957 gnd.n3579 gnd.n3578 19.3944
R7958 gnd.n3628 gnd.n3627 19.3944
R7959 gnd.n3627 gnd.n3626 19.3944
R7960 gnd.n3626 gnd.n3623 19.3944
R7961 gnd.n3623 gnd.n3622 19.3944
R7962 gnd.n3622 gnd.n3619 19.3944
R7963 gnd.n3619 gnd.n3618 19.3944
R7964 gnd.n3618 gnd.n3615 19.3944
R7965 gnd.n3615 gnd.n3614 19.3944
R7966 gnd.n3614 gnd.n3611 19.3944
R7967 gnd.n3611 gnd.n3610 19.3944
R7968 gnd.n3610 gnd.n3607 19.3944
R7969 gnd.n3607 gnd.n3606 19.3944
R7970 gnd.n3606 gnd.n3603 19.3944
R7971 gnd.n3603 gnd.n3602 19.3944
R7972 gnd.n3602 gnd.n3599 19.3944
R7973 gnd.n3599 gnd.n3598 19.3944
R7974 gnd.n3598 gnd.n3595 19.3944
R7975 gnd.n3595 gnd.n3594 19.3944
R7976 gnd.n3594 gnd.n3591 19.3944
R7977 gnd.n3591 gnd.n3590 19.3944
R7978 gnd.n3590 gnd.n3587 19.3944
R7979 gnd.n3587 gnd.n3586 19.3944
R7980 gnd.n2910 gnd.n2619 19.3944
R7981 gnd.n2920 gnd.n2619 19.3944
R7982 gnd.n2921 gnd.n2920 19.3944
R7983 gnd.n2921 gnd.n2600 19.3944
R7984 gnd.n2941 gnd.n2600 19.3944
R7985 gnd.n2941 gnd.n2592 19.3944
R7986 gnd.n2951 gnd.n2592 19.3944
R7987 gnd.n2952 gnd.n2951 19.3944
R7988 gnd.n2953 gnd.n2952 19.3944
R7989 gnd.n2953 gnd.n2575 19.3944
R7990 gnd.n2970 gnd.n2575 19.3944
R7991 gnd.n2973 gnd.n2970 19.3944
R7992 gnd.n2973 gnd.n2972 19.3944
R7993 gnd.n2972 gnd.n2548 19.3944
R7994 gnd.n3012 gnd.n2548 19.3944
R7995 gnd.n3012 gnd.n2545 19.3944
R7996 gnd.n3018 gnd.n2545 19.3944
R7997 gnd.n3019 gnd.n3018 19.3944
R7998 gnd.n3019 gnd.n2543 19.3944
R7999 gnd.n3025 gnd.n2543 19.3944
R8000 gnd.n3028 gnd.n3025 19.3944
R8001 gnd.n3030 gnd.n3028 19.3944
R8002 gnd.n3036 gnd.n3030 19.3944
R8003 gnd.n3036 gnd.n3035 19.3944
R8004 gnd.n3035 gnd.n2418 19.3944
R8005 gnd.n3102 gnd.n2418 19.3944
R8006 gnd.n3103 gnd.n3102 19.3944
R8007 gnd.n3103 gnd.n2411 19.3944
R8008 gnd.n3114 gnd.n2411 19.3944
R8009 gnd.n3115 gnd.n3114 19.3944
R8010 gnd.n3115 gnd.n2394 19.3944
R8011 gnd.n2394 gnd.n2392 19.3944
R8012 gnd.n3139 gnd.n2392 19.3944
R8013 gnd.n3140 gnd.n3139 19.3944
R8014 gnd.n3140 gnd.n2363 19.3944
R8015 gnd.n3187 gnd.n2363 19.3944
R8016 gnd.n3188 gnd.n3187 19.3944
R8017 gnd.n3188 gnd.n2356 19.3944
R8018 gnd.n3199 gnd.n2356 19.3944
R8019 gnd.n3200 gnd.n3199 19.3944
R8020 gnd.n3200 gnd.n2339 19.3944
R8021 gnd.n2339 gnd.n2337 19.3944
R8022 gnd.n3224 gnd.n2337 19.3944
R8023 gnd.n3225 gnd.n3224 19.3944
R8024 gnd.n3225 gnd.n2309 19.3944
R8025 gnd.n3276 gnd.n2309 19.3944
R8026 gnd.n3277 gnd.n3276 19.3944
R8027 gnd.n3277 gnd.n2302 19.3944
R8028 gnd.n3544 gnd.n2302 19.3944
R8029 gnd.n3545 gnd.n3544 19.3944
R8030 gnd.n3545 gnd.n2283 19.3944
R8031 gnd.n3570 gnd.n2283 19.3944
R8032 gnd.n3570 gnd.n2284 19.3944
R8033 gnd.n2901 gnd.n2900 19.3944
R8034 gnd.n2900 gnd.n2633 19.3944
R8035 gnd.n2656 gnd.n2633 19.3944
R8036 gnd.n2659 gnd.n2656 19.3944
R8037 gnd.n2659 gnd.n2652 19.3944
R8038 gnd.n2663 gnd.n2652 19.3944
R8039 gnd.n2666 gnd.n2663 19.3944
R8040 gnd.n2669 gnd.n2666 19.3944
R8041 gnd.n2669 gnd.n2650 19.3944
R8042 gnd.n2673 gnd.n2650 19.3944
R8043 gnd.n2676 gnd.n2673 19.3944
R8044 gnd.n2679 gnd.n2676 19.3944
R8045 gnd.n2679 gnd.n2648 19.3944
R8046 gnd.n2683 gnd.n2648 19.3944
R8047 gnd.n2906 gnd.n2905 19.3944
R8048 gnd.n2905 gnd.n2609 19.3944
R8049 gnd.n2931 gnd.n2609 19.3944
R8050 gnd.n2931 gnd.n2607 19.3944
R8051 gnd.n2937 gnd.n2607 19.3944
R8052 gnd.n2937 gnd.n2936 19.3944
R8053 gnd.n2936 gnd.n2581 19.3944
R8054 gnd.n2961 gnd.n2581 19.3944
R8055 gnd.n2961 gnd.n2579 19.3944
R8056 gnd.n2965 gnd.n2579 19.3944
R8057 gnd.n2965 gnd.n2559 19.3944
R8058 gnd.n2992 gnd.n2559 19.3944
R8059 gnd.n2992 gnd.n2557 19.3944
R8060 gnd.n3002 gnd.n2557 19.3944
R8061 gnd.n3002 gnd.n3001 19.3944
R8062 gnd.n3001 gnd.n3000 19.3944
R8063 gnd.n3000 gnd.n2506 19.3944
R8064 gnd.n3050 gnd.n2506 19.3944
R8065 gnd.n3050 gnd.n3049 19.3944
R8066 gnd.n3049 gnd.n3048 19.3944
R8067 gnd.n3048 gnd.n2510 19.3944
R8068 gnd.n2530 gnd.n2510 19.3944
R8069 gnd.n2530 gnd.n2428 19.3944
R8070 gnd.n3087 gnd.n2428 19.3944
R8071 gnd.n3087 gnd.n2426 19.3944
R8072 gnd.n3093 gnd.n2426 19.3944
R8073 gnd.n3093 gnd.n3092 19.3944
R8074 gnd.n3092 gnd.n2401 19.3944
R8075 gnd.n3127 gnd.n2401 19.3944
R8076 gnd.n3127 gnd.n2399 19.3944
R8077 gnd.n3133 gnd.n2399 19.3944
R8078 gnd.n3133 gnd.n3132 19.3944
R8079 gnd.n3132 gnd.n2374 19.3944
R8080 gnd.n3172 gnd.n2374 19.3944
R8081 gnd.n3172 gnd.n2372 19.3944
R8082 gnd.n3178 gnd.n2372 19.3944
R8083 gnd.n3178 gnd.n3177 19.3944
R8084 gnd.n3177 gnd.n2346 19.3944
R8085 gnd.n3212 gnd.n2346 19.3944
R8086 gnd.n3212 gnd.n2344 19.3944
R8087 gnd.n3218 gnd.n2344 19.3944
R8088 gnd.n3218 gnd.n3217 19.3944
R8089 gnd.n3217 gnd.n2319 19.3944
R8090 gnd.n3261 gnd.n2319 19.3944
R8091 gnd.n3261 gnd.n2317 19.3944
R8092 gnd.n3267 gnd.n2317 19.3944
R8093 gnd.n3267 gnd.n3266 19.3944
R8094 gnd.n3266 gnd.n2292 19.3944
R8095 gnd.n3555 gnd.n2292 19.3944
R8096 gnd.n3555 gnd.n2290 19.3944
R8097 gnd.n3563 gnd.n2290 19.3944
R8098 gnd.n3563 gnd.n3562 19.3944
R8099 gnd.n3562 gnd.n3561 19.3944
R8100 gnd.n3664 gnd.n3663 19.3944
R8101 gnd.n3663 gnd.n2231 19.3944
R8102 gnd.n3659 gnd.n2231 19.3944
R8103 gnd.n3659 gnd.n3656 19.3944
R8104 gnd.n3656 gnd.n3653 19.3944
R8105 gnd.n3653 gnd.n3652 19.3944
R8106 gnd.n3652 gnd.n3649 19.3944
R8107 gnd.n3649 gnd.n3648 19.3944
R8108 gnd.n3648 gnd.n3645 19.3944
R8109 gnd.n3645 gnd.n3644 19.3944
R8110 gnd.n3644 gnd.n3641 19.3944
R8111 gnd.n3641 gnd.n3640 19.3944
R8112 gnd.n3640 gnd.n3637 19.3944
R8113 gnd.n3637 gnd.n3636 19.3944
R8114 gnd.n2821 gnd.n2720 19.3944
R8115 gnd.n2821 gnd.n2711 19.3944
R8116 gnd.n2834 gnd.n2711 19.3944
R8117 gnd.n2834 gnd.n2709 19.3944
R8118 gnd.n2838 gnd.n2709 19.3944
R8119 gnd.n2838 gnd.n2699 19.3944
R8120 gnd.n2850 gnd.n2699 19.3944
R8121 gnd.n2850 gnd.n2697 19.3944
R8122 gnd.n2884 gnd.n2697 19.3944
R8123 gnd.n2884 gnd.n2883 19.3944
R8124 gnd.n2883 gnd.n2882 19.3944
R8125 gnd.n2882 gnd.n2881 19.3944
R8126 gnd.n2881 gnd.n2878 19.3944
R8127 gnd.n2878 gnd.n2877 19.3944
R8128 gnd.n2877 gnd.n2876 19.3944
R8129 gnd.n2876 gnd.n2874 19.3944
R8130 gnd.n2874 gnd.n2873 19.3944
R8131 gnd.n2873 gnd.n2870 19.3944
R8132 gnd.n2870 gnd.n2869 19.3944
R8133 gnd.n2869 gnd.n2868 19.3944
R8134 gnd.n2868 gnd.n2866 19.3944
R8135 gnd.n2866 gnd.n2565 19.3944
R8136 gnd.n2981 gnd.n2565 19.3944
R8137 gnd.n2981 gnd.n2563 19.3944
R8138 gnd.n2987 gnd.n2563 19.3944
R8139 gnd.n2987 gnd.n2986 19.3944
R8140 gnd.n2986 gnd.n2487 19.3944
R8141 gnd.n3061 gnd.n2487 19.3944
R8142 gnd.n3061 gnd.n2488 19.3944
R8143 gnd.n2535 gnd.n2534 19.3944
R8144 gnd.n2538 gnd.n2537 19.3944
R8145 gnd.n2525 gnd.n2524 19.3944
R8146 gnd.n3080 gnd.n2433 19.3944
R8147 gnd.n3080 gnd.n3079 19.3944
R8148 gnd.n3079 gnd.n3078 19.3944
R8149 gnd.n3078 gnd.n3076 19.3944
R8150 gnd.n3076 gnd.n3075 19.3944
R8151 gnd.n3075 gnd.n3073 19.3944
R8152 gnd.n3073 gnd.n3072 19.3944
R8153 gnd.n3072 gnd.n2382 19.3944
R8154 gnd.n3148 gnd.n2382 19.3944
R8155 gnd.n3148 gnd.n2380 19.3944
R8156 gnd.n3167 gnd.n2380 19.3944
R8157 gnd.n3167 gnd.n3166 19.3944
R8158 gnd.n3166 gnd.n3165 19.3944
R8159 gnd.n3165 gnd.n3163 19.3944
R8160 gnd.n3163 gnd.n3162 19.3944
R8161 gnd.n3162 gnd.n3160 19.3944
R8162 gnd.n3160 gnd.n3159 19.3944
R8163 gnd.n3159 gnd.n2326 19.3944
R8164 gnd.n3233 gnd.n2326 19.3944
R8165 gnd.n3233 gnd.n2324 19.3944
R8166 gnd.n3256 gnd.n2324 19.3944
R8167 gnd.n3256 gnd.n3255 19.3944
R8168 gnd.n3255 gnd.n3254 19.3944
R8169 gnd.n3254 gnd.n3251 19.3944
R8170 gnd.n3251 gnd.n3250 19.3944
R8171 gnd.n3250 gnd.n3248 19.3944
R8172 gnd.n3248 gnd.n3247 19.3944
R8173 gnd.n3247 gnd.n3245 19.3944
R8174 gnd.n3245 gnd.n2278 19.3944
R8175 gnd.n2826 gnd.n2716 19.3944
R8176 gnd.n2826 gnd.n2714 19.3944
R8177 gnd.n2830 gnd.n2714 19.3944
R8178 gnd.n2830 gnd.n2705 19.3944
R8179 gnd.n2842 gnd.n2705 19.3944
R8180 gnd.n2842 gnd.n2703 19.3944
R8181 gnd.n2846 gnd.n2703 19.3944
R8182 gnd.n2846 gnd.n2692 19.3944
R8183 gnd.n2888 gnd.n2692 19.3944
R8184 gnd.n2888 gnd.n2646 19.3944
R8185 gnd.n2894 gnd.n2646 19.3944
R8186 gnd.n2894 gnd.n2893 19.3944
R8187 gnd.n2893 gnd.n2624 19.3944
R8188 gnd.n2915 gnd.n2624 19.3944
R8189 gnd.n2915 gnd.n2617 19.3944
R8190 gnd.n2926 gnd.n2617 19.3944
R8191 gnd.n2926 gnd.n2925 19.3944
R8192 gnd.n2925 gnd.n2598 19.3944
R8193 gnd.n2946 gnd.n2598 19.3944
R8194 gnd.n2946 gnd.n2588 19.3944
R8195 gnd.n2956 gnd.n2588 19.3944
R8196 gnd.n2956 gnd.n2571 19.3944
R8197 gnd.n2977 gnd.n2571 19.3944
R8198 gnd.n2977 gnd.n2976 19.3944
R8199 gnd.n2976 gnd.n2550 19.3944
R8200 gnd.n3007 gnd.n2550 19.3944
R8201 gnd.n3007 gnd.n2495 19.3944
R8202 gnd.n3057 gnd.n2495 19.3944
R8203 gnd.n3057 gnd.n3056 19.3944
R8204 gnd.n3056 gnd.n3055 19.3944
R8205 gnd.n3055 gnd.n2499 19.3944
R8206 gnd.n2517 gnd.n2499 19.3944
R8207 gnd.n3043 gnd.n2517 19.3944
R8208 gnd.n3043 gnd.n3042 19.3944
R8209 gnd.n3042 gnd.n3041 19.3944
R8210 gnd.n3041 gnd.n2521 19.3944
R8211 gnd.n2521 gnd.n2420 19.3944
R8212 gnd.n3098 gnd.n2420 19.3944
R8213 gnd.n3098 gnd.n2413 19.3944
R8214 gnd.n3109 gnd.n2413 19.3944
R8215 gnd.n3109 gnd.n2409 19.3944
R8216 gnd.n3122 gnd.n2409 19.3944
R8217 gnd.n3122 gnd.n3121 19.3944
R8218 gnd.n3121 gnd.n2388 19.3944
R8219 gnd.n3144 gnd.n2388 19.3944
R8220 gnd.n3144 gnd.n3143 19.3944
R8221 gnd.n3143 gnd.n2365 19.3944
R8222 gnd.n3183 gnd.n2365 19.3944
R8223 gnd.n3183 gnd.n2358 19.3944
R8224 gnd.n3194 gnd.n2358 19.3944
R8225 gnd.n3194 gnd.n2354 19.3944
R8226 gnd.n3207 gnd.n2354 19.3944
R8227 gnd.n3207 gnd.n3206 19.3944
R8228 gnd.n3206 gnd.n2333 19.3944
R8229 gnd.n3229 gnd.n2333 19.3944
R8230 gnd.n3229 gnd.n3228 19.3944
R8231 gnd.n3228 gnd.n2311 19.3944
R8232 gnd.n3272 gnd.n2311 19.3944
R8233 gnd.n3272 gnd.n2304 19.3944
R8234 gnd.n3283 gnd.n2304 19.3944
R8235 gnd.n3283 gnd.n2300 19.3944
R8236 gnd.n3550 gnd.n2300 19.3944
R8237 gnd.n3550 gnd.n3549 19.3944
R8238 gnd.n3549 gnd.n2281 19.3944
R8239 gnd.n3573 gnd.n2281 19.3944
R8240 gnd.n5847 gnd.n909 19.3944
R8241 gnd.n5847 gnd.n5846 19.3944
R8242 gnd.n5846 gnd.n912 19.3944
R8243 gnd.n5839 gnd.n912 19.3944
R8244 gnd.n5839 gnd.n5838 19.3944
R8245 gnd.n5838 gnd.n922 19.3944
R8246 gnd.n5831 gnd.n922 19.3944
R8247 gnd.n5831 gnd.n5830 19.3944
R8248 gnd.n5830 gnd.n930 19.3944
R8249 gnd.n5823 gnd.n930 19.3944
R8250 gnd.n5823 gnd.n5822 19.3944
R8251 gnd.n5822 gnd.n940 19.3944
R8252 gnd.n5815 gnd.n940 19.3944
R8253 gnd.n5815 gnd.n5814 19.3944
R8254 gnd.n5814 gnd.n948 19.3944
R8255 gnd.n5807 gnd.n948 19.3944
R8256 gnd.n6564 gnd.n308 19.3944
R8257 gnd.n6570 gnd.n308 19.3944
R8258 gnd.n6570 gnd.n306 19.3944
R8259 gnd.n6574 gnd.n306 19.3944
R8260 gnd.n6574 gnd.n302 19.3944
R8261 gnd.n6580 gnd.n302 19.3944
R8262 gnd.n6580 gnd.n300 19.3944
R8263 gnd.n6584 gnd.n300 19.3944
R8264 gnd.n6584 gnd.n296 19.3944
R8265 gnd.n6590 gnd.n296 19.3944
R8266 gnd.n6590 gnd.n294 19.3944
R8267 gnd.n6594 gnd.n294 19.3944
R8268 gnd.n6594 gnd.n290 19.3944
R8269 gnd.n6600 gnd.n290 19.3944
R8270 gnd.n6600 gnd.n288 19.3944
R8271 gnd.n6604 gnd.n288 19.3944
R8272 gnd.n6604 gnd.n284 19.3944
R8273 gnd.n6610 gnd.n284 19.3944
R8274 gnd.n6610 gnd.n282 19.3944
R8275 gnd.n6614 gnd.n282 19.3944
R8276 gnd.n6614 gnd.n278 19.3944
R8277 gnd.n6620 gnd.n278 19.3944
R8278 gnd.n6620 gnd.n276 19.3944
R8279 gnd.n6624 gnd.n276 19.3944
R8280 gnd.n6624 gnd.n272 19.3944
R8281 gnd.n6630 gnd.n272 19.3944
R8282 gnd.n6630 gnd.n270 19.3944
R8283 gnd.n6634 gnd.n270 19.3944
R8284 gnd.n6634 gnd.n266 19.3944
R8285 gnd.n6640 gnd.n266 19.3944
R8286 gnd.n6640 gnd.n264 19.3944
R8287 gnd.n6644 gnd.n264 19.3944
R8288 gnd.n6644 gnd.n260 19.3944
R8289 gnd.n6650 gnd.n260 19.3944
R8290 gnd.n6650 gnd.n258 19.3944
R8291 gnd.n6654 gnd.n258 19.3944
R8292 gnd.n6654 gnd.n254 19.3944
R8293 gnd.n6660 gnd.n254 19.3944
R8294 gnd.n6660 gnd.n252 19.3944
R8295 gnd.n6664 gnd.n252 19.3944
R8296 gnd.n6664 gnd.n248 19.3944
R8297 gnd.n6670 gnd.n248 19.3944
R8298 gnd.n6670 gnd.n246 19.3944
R8299 gnd.n6674 gnd.n246 19.3944
R8300 gnd.n6674 gnd.n242 19.3944
R8301 gnd.n6680 gnd.n242 19.3944
R8302 gnd.n6680 gnd.n240 19.3944
R8303 gnd.n6684 gnd.n240 19.3944
R8304 gnd.n6684 gnd.n236 19.3944
R8305 gnd.n6690 gnd.n236 19.3944
R8306 gnd.n6690 gnd.n234 19.3944
R8307 gnd.n6694 gnd.n234 19.3944
R8308 gnd.n6694 gnd.n230 19.3944
R8309 gnd.n6700 gnd.n230 19.3944
R8310 gnd.n6700 gnd.n228 19.3944
R8311 gnd.n6704 gnd.n228 19.3944
R8312 gnd.n6704 gnd.n224 19.3944
R8313 gnd.n6710 gnd.n224 19.3944
R8314 gnd.n6710 gnd.n222 19.3944
R8315 gnd.n6714 gnd.n222 19.3944
R8316 gnd.n6714 gnd.n218 19.3944
R8317 gnd.n6720 gnd.n218 19.3944
R8318 gnd.n6720 gnd.n216 19.3944
R8319 gnd.n6724 gnd.n216 19.3944
R8320 gnd.n6724 gnd.n212 19.3944
R8321 gnd.n6730 gnd.n212 19.3944
R8322 gnd.n6730 gnd.n210 19.3944
R8323 gnd.n6734 gnd.n210 19.3944
R8324 gnd.n6734 gnd.n206 19.3944
R8325 gnd.n6740 gnd.n206 19.3944
R8326 gnd.n6740 gnd.n204 19.3944
R8327 gnd.n6744 gnd.n204 19.3944
R8328 gnd.n6744 gnd.n200 19.3944
R8329 gnd.n6750 gnd.n200 19.3944
R8330 gnd.n6750 gnd.n198 19.3944
R8331 gnd.n6754 gnd.n198 19.3944
R8332 gnd.n6754 gnd.n194 19.3944
R8333 gnd.n6760 gnd.n194 19.3944
R8334 gnd.n6760 gnd.n192 19.3944
R8335 gnd.n6764 gnd.n192 19.3944
R8336 gnd.n6764 gnd.n188 19.3944
R8337 gnd.n6771 gnd.n188 19.3944
R8338 gnd.n6771 gnd.n186 19.3944
R8339 gnd.n6775 gnd.n186 19.3944
R8340 gnd.n6143 gnd.n559 19.3944
R8341 gnd.n6149 gnd.n559 19.3944
R8342 gnd.n6149 gnd.n557 19.3944
R8343 gnd.n6153 gnd.n557 19.3944
R8344 gnd.n6153 gnd.n553 19.3944
R8345 gnd.n6159 gnd.n553 19.3944
R8346 gnd.n6159 gnd.n551 19.3944
R8347 gnd.n6163 gnd.n551 19.3944
R8348 gnd.n6163 gnd.n547 19.3944
R8349 gnd.n6169 gnd.n547 19.3944
R8350 gnd.n6169 gnd.n545 19.3944
R8351 gnd.n6173 gnd.n545 19.3944
R8352 gnd.n6173 gnd.n541 19.3944
R8353 gnd.n6179 gnd.n541 19.3944
R8354 gnd.n6179 gnd.n539 19.3944
R8355 gnd.n6183 gnd.n539 19.3944
R8356 gnd.n6183 gnd.n535 19.3944
R8357 gnd.n6189 gnd.n535 19.3944
R8358 gnd.n6189 gnd.n533 19.3944
R8359 gnd.n6193 gnd.n533 19.3944
R8360 gnd.n6193 gnd.n529 19.3944
R8361 gnd.n6199 gnd.n529 19.3944
R8362 gnd.n6199 gnd.n527 19.3944
R8363 gnd.n6203 gnd.n527 19.3944
R8364 gnd.n6203 gnd.n523 19.3944
R8365 gnd.n6209 gnd.n523 19.3944
R8366 gnd.n6209 gnd.n521 19.3944
R8367 gnd.n6213 gnd.n521 19.3944
R8368 gnd.n6213 gnd.n517 19.3944
R8369 gnd.n6219 gnd.n517 19.3944
R8370 gnd.n6219 gnd.n515 19.3944
R8371 gnd.n6223 gnd.n515 19.3944
R8372 gnd.n6223 gnd.n511 19.3944
R8373 gnd.n6229 gnd.n511 19.3944
R8374 gnd.n6229 gnd.n509 19.3944
R8375 gnd.n6233 gnd.n509 19.3944
R8376 gnd.n6233 gnd.n505 19.3944
R8377 gnd.n6239 gnd.n505 19.3944
R8378 gnd.n6239 gnd.n503 19.3944
R8379 gnd.n6243 gnd.n503 19.3944
R8380 gnd.n6243 gnd.n499 19.3944
R8381 gnd.n6249 gnd.n499 19.3944
R8382 gnd.n6249 gnd.n497 19.3944
R8383 gnd.n6253 gnd.n497 19.3944
R8384 gnd.n6253 gnd.n493 19.3944
R8385 gnd.n6259 gnd.n493 19.3944
R8386 gnd.n6259 gnd.n491 19.3944
R8387 gnd.n6263 gnd.n491 19.3944
R8388 gnd.n6263 gnd.n487 19.3944
R8389 gnd.n6269 gnd.n487 19.3944
R8390 gnd.n6269 gnd.n485 19.3944
R8391 gnd.n6273 gnd.n485 19.3944
R8392 gnd.n6273 gnd.n481 19.3944
R8393 gnd.n6279 gnd.n481 19.3944
R8394 gnd.n6279 gnd.n479 19.3944
R8395 gnd.n6283 gnd.n479 19.3944
R8396 gnd.n6283 gnd.n475 19.3944
R8397 gnd.n6289 gnd.n475 19.3944
R8398 gnd.n6289 gnd.n473 19.3944
R8399 gnd.n6293 gnd.n473 19.3944
R8400 gnd.n6293 gnd.n469 19.3944
R8401 gnd.n6299 gnd.n469 19.3944
R8402 gnd.n6299 gnd.n467 19.3944
R8403 gnd.n6303 gnd.n467 19.3944
R8404 gnd.n6303 gnd.n463 19.3944
R8405 gnd.n6309 gnd.n463 19.3944
R8406 gnd.n6309 gnd.n461 19.3944
R8407 gnd.n6313 gnd.n461 19.3944
R8408 gnd.n6313 gnd.n457 19.3944
R8409 gnd.n6319 gnd.n457 19.3944
R8410 gnd.n6319 gnd.n455 19.3944
R8411 gnd.n6323 gnd.n455 19.3944
R8412 gnd.n6323 gnd.n451 19.3944
R8413 gnd.n6329 gnd.n451 19.3944
R8414 gnd.n6329 gnd.n449 19.3944
R8415 gnd.n6333 gnd.n449 19.3944
R8416 gnd.n6333 gnd.n445 19.3944
R8417 gnd.n6339 gnd.n445 19.3944
R8418 gnd.n6339 gnd.n443 19.3944
R8419 gnd.n6343 gnd.n443 19.3944
R8420 gnd.n6343 gnd.n439 19.3944
R8421 gnd.n6349 gnd.n439 19.3944
R8422 gnd.n6349 gnd.n437 19.3944
R8423 gnd.n6353 gnd.n437 19.3944
R8424 gnd.n6353 gnd.n433 19.3944
R8425 gnd.n6359 gnd.n433 19.3944
R8426 gnd.n6359 gnd.n431 19.3944
R8427 gnd.n6363 gnd.n431 19.3944
R8428 gnd.n6363 gnd.n427 19.3944
R8429 gnd.n6369 gnd.n427 19.3944
R8430 gnd.n6369 gnd.n425 19.3944
R8431 gnd.n6373 gnd.n425 19.3944
R8432 gnd.n6373 gnd.n421 19.3944
R8433 gnd.n6379 gnd.n421 19.3944
R8434 gnd.n6379 gnd.n419 19.3944
R8435 gnd.n6383 gnd.n419 19.3944
R8436 gnd.n6383 gnd.n415 19.3944
R8437 gnd.n6389 gnd.n415 19.3944
R8438 gnd.n6389 gnd.n413 19.3944
R8439 gnd.n6393 gnd.n413 19.3944
R8440 gnd.n6393 gnd.n409 19.3944
R8441 gnd.n6399 gnd.n409 19.3944
R8442 gnd.n6399 gnd.n407 19.3944
R8443 gnd.n6403 gnd.n407 19.3944
R8444 gnd.n6403 gnd.n403 19.3944
R8445 gnd.n6409 gnd.n403 19.3944
R8446 gnd.n6409 gnd.n401 19.3944
R8447 gnd.n6413 gnd.n401 19.3944
R8448 gnd.n6413 gnd.n397 19.3944
R8449 gnd.n6419 gnd.n397 19.3944
R8450 gnd.n6419 gnd.n395 19.3944
R8451 gnd.n6423 gnd.n395 19.3944
R8452 gnd.n6423 gnd.n391 19.3944
R8453 gnd.n6429 gnd.n391 19.3944
R8454 gnd.n6429 gnd.n389 19.3944
R8455 gnd.n6433 gnd.n389 19.3944
R8456 gnd.n6433 gnd.n385 19.3944
R8457 gnd.n6439 gnd.n385 19.3944
R8458 gnd.n6439 gnd.n383 19.3944
R8459 gnd.n6443 gnd.n383 19.3944
R8460 gnd.n6443 gnd.n379 19.3944
R8461 gnd.n6449 gnd.n379 19.3944
R8462 gnd.n6449 gnd.n377 19.3944
R8463 gnd.n6453 gnd.n377 19.3944
R8464 gnd.n6453 gnd.n373 19.3944
R8465 gnd.n6459 gnd.n373 19.3944
R8466 gnd.n6459 gnd.n371 19.3944
R8467 gnd.n6463 gnd.n371 19.3944
R8468 gnd.n6463 gnd.n367 19.3944
R8469 gnd.n6469 gnd.n367 19.3944
R8470 gnd.n6469 gnd.n365 19.3944
R8471 gnd.n6473 gnd.n365 19.3944
R8472 gnd.n6473 gnd.n361 19.3944
R8473 gnd.n6479 gnd.n361 19.3944
R8474 gnd.n6479 gnd.n359 19.3944
R8475 gnd.n6483 gnd.n359 19.3944
R8476 gnd.n6483 gnd.n355 19.3944
R8477 gnd.n6489 gnd.n355 19.3944
R8478 gnd.n6489 gnd.n353 19.3944
R8479 gnd.n6493 gnd.n353 19.3944
R8480 gnd.n6493 gnd.n349 19.3944
R8481 gnd.n6499 gnd.n349 19.3944
R8482 gnd.n6499 gnd.n347 19.3944
R8483 gnd.n6503 gnd.n347 19.3944
R8484 gnd.n6503 gnd.n343 19.3944
R8485 gnd.n6509 gnd.n343 19.3944
R8486 gnd.n6509 gnd.n341 19.3944
R8487 gnd.n6513 gnd.n341 19.3944
R8488 gnd.n6513 gnd.n337 19.3944
R8489 gnd.n6519 gnd.n337 19.3944
R8490 gnd.n6519 gnd.n335 19.3944
R8491 gnd.n6523 gnd.n335 19.3944
R8492 gnd.n6523 gnd.n331 19.3944
R8493 gnd.n6529 gnd.n331 19.3944
R8494 gnd.n6529 gnd.n329 19.3944
R8495 gnd.n6533 gnd.n329 19.3944
R8496 gnd.n6533 gnd.n325 19.3944
R8497 gnd.n6539 gnd.n325 19.3944
R8498 gnd.n6539 gnd.n323 19.3944
R8499 gnd.n6543 gnd.n323 19.3944
R8500 gnd.n6543 gnd.n319 19.3944
R8501 gnd.n6549 gnd.n319 19.3944
R8502 gnd.n6549 gnd.n317 19.3944
R8503 gnd.n6554 gnd.n317 19.3944
R8504 gnd.n6554 gnd.n313 19.3944
R8505 gnd.n6560 gnd.n313 19.3944
R8506 gnd.n6561 gnd.n6560 19.3944
R8507 gnd.n5494 gnd.n5493 19.3944
R8508 gnd.n5493 gnd.n5492 19.3944
R8509 gnd.n5492 gnd.n5491 19.3944
R8510 gnd.n5491 gnd.n5489 19.3944
R8511 gnd.n5489 gnd.n5486 19.3944
R8512 gnd.n5486 gnd.n5485 19.3944
R8513 gnd.n5485 gnd.n5482 19.3944
R8514 gnd.n5482 gnd.n5481 19.3944
R8515 gnd.n5481 gnd.n5478 19.3944
R8516 gnd.n5478 gnd.n5477 19.3944
R8517 gnd.n5477 gnd.n5474 19.3944
R8518 gnd.n5474 gnd.n5473 19.3944
R8519 gnd.n5473 gnd.n5470 19.3944
R8520 gnd.n5470 gnd.n5469 19.3944
R8521 gnd.n5469 gnd.n5466 19.3944
R8522 gnd.n5466 gnd.n5465 19.3944
R8523 gnd.n5465 gnd.n5462 19.3944
R8524 gnd.n5460 gnd.n5457 19.3944
R8525 gnd.n5457 gnd.n5456 19.3944
R8526 gnd.n5456 gnd.n5453 19.3944
R8527 gnd.n5453 gnd.n5452 19.3944
R8528 gnd.n5452 gnd.n5449 19.3944
R8529 gnd.n5449 gnd.n5448 19.3944
R8530 gnd.n5448 gnd.n5445 19.3944
R8531 gnd.n5443 gnd.n5440 19.3944
R8532 gnd.n5440 gnd.n5439 19.3944
R8533 gnd.n5439 gnd.n5436 19.3944
R8534 gnd.n5436 gnd.n5435 19.3944
R8535 gnd.n5435 gnd.n5432 19.3944
R8536 gnd.n5432 gnd.n5431 19.3944
R8537 gnd.n5431 gnd.n5428 19.3944
R8538 gnd.n5428 gnd.n5427 19.3944
R8539 gnd.n5423 gnd.n5420 19.3944
R8540 gnd.n5420 gnd.n5419 19.3944
R8541 gnd.n5419 gnd.n5416 19.3944
R8542 gnd.n5416 gnd.n5415 19.3944
R8543 gnd.n5415 gnd.n5412 19.3944
R8544 gnd.n5412 gnd.n5411 19.3944
R8545 gnd.n5411 gnd.n5408 19.3944
R8546 gnd.n5408 gnd.n5407 19.3944
R8547 gnd.n5407 gnd.n5404 19.3944
R8548 gnd.n5404 gnd.n5403 19.3944
R8549 gnd.n5403 gnd.n5400 19.3944
R8550 gnd.n5400 gnd.n5399 19.3944
R8551 gnd.n5399 gnd.n5396 19.3944
R8552 gnd.n5396 gnd.n5395 19.3944
R8553 gnd.n5395 gnd.n5392 19.3944
R8554 gnd.n5392 gnd.n5391 19.3944
R8555 gnd.n5391 gnd.n5388 19.3944
R8556 gnd.n5388 gnd.n5387 19.3944
R8557 gnd.n5371 gnd.n1483 19.3944
R8558 gnd.n5371 gnd.n5370 19.3944
R8559 gnd.n5370 gnd.n1492 19.3944
R8560 gnd.n5185 gnd.n1492 19.3944
R8561 gnd.n5188 gnd.n5185 19.3944
R8562 gnd.n5189 gnd.n5188 19.3944
R8563 gnd.n5194 gnd.n5189 19.3944
R8564 gnd.n5195 gnd.n5194 19.3944
R8565 gnd.n5199 gnd.n5195 19.3944
R8566 gnd.n5199 gnd.n5198 19.3944
R8567 gnd.n5198 gnd.n5197 19.3944
R8568 gnd.n5197 gnd.n1611 19.3944
R8569 gnd.n5271 gnd.n1611 19.3944
R8570 gnd.n5272 gnd.n5271 19.3944
R8571 gnd.n5274 gnd.n5272 19.3944
R8572 gnd.n5274 gnd.n1605 19.3944
R8573 gnd.n5290 gnd.n1605 19.3944
R8574 gnd.n5291 gnd.n5290 19.3944
R8575 gnd.n5292 gnd.n5291 19.3944
R8576 gnd.n5292 gnd.n1601 19.3944
R8577 gnd.n5300 gnd.n1601 19.3944
R8578 gnd.n5302 gnd.n5300 19.3944
R8579 gnd.n5302 gnd.n5301 19.3944
R8580 gnd.n5301 gnd.n178 19.3944
R8581 gnd.n6789 gnd.n178 19.3944
R8582 gnd.n6789 gnd.n174 19.3944
R8583 gnd.n7118 gnd.n174 19.3944
R8584 gnd.n7119 gnd.n7118 19.3944
R8585 gnd.n7122 gnd.n7119 19.3944
R8586 gnd.n7123 gnd.n7122 19.3944
R8587 gnd.n7125 gnd.n7123 19.3944
R8588 gnd.n7126 gnd.n7125 19.3944
R8589 gnd.n7129 gnd.n7126 19.3944
R8590 gnd.n7130 gnd.n7129 19.3944
R8591 gnd.n7132 gnd.n7130 19.3944
R8592 gnd.n7133 gnd.n7132 19.3944
R8593 gnd.n7136 gnd.n7133 19.3944
R8594 gnd.n7137 gnd.n7136 19.3944
R8595 gnd.n7139 gnd.n7137 19.3944
R8596 gnd.n7140 gnd.n7139 19.3944
R8597 gnd.n7142 gnd.n7140 19.3944
R8598 gnd.n7143 gnd.n7142 19.3944
R8599 gnd.n5374 gnd.n5373 19.3944
R8600 gnd.n5373 gnd.n1490 19.3944
R8601 gnd.n1514 gnd.n1490 19.3944
R8602 gnd.n5360 gnd.n1514 19.3944
R8603 gnd.n5360 gnd.n5359 19.3944
R8604 gnd.n5359 gnd.n5358 19.3944
R8605 gnd.n5358 gnd.n1519 19.3944
R8606 gnd.n5348 gnd.n1519 19.3944
R8607 gnd.n5348 gnd.n5347 19.3944
R8608 gnd.n5347 gnd.n5346 19.3944
R8609 gnd.n5346 gnd.n1539 19.3944
R8610 gnd.n5336 gnd.n1539 19.3944
R8611 gnd.n5336 gnd.n5335 19.3944
R8612 gnd.n5335 gnd.n5334 19.3944
R8613 gnd.n5334 gnd.n1559 19.3944
R8614 gnd.n5324 gnd.n1559 19.3944
R8615 gnd.n5324 gnd.n5323 19.3944
R8616 gnd.n5323 gnd.n5322 19.3944
R8617 gnd.n5322 gnd.n1576 19.3944
R8618 gnd.n5295 gnd.n1576 19.3944
R8619 gnd.n5295 gnd.n1599 19.3944
R8620 gnd.n5304 gnd.n1599 19.3944
R8621 gnd.n5304 gnd.n180 19.3944
R8622 gnd.n6786 gnd.n180 19.3944
R8623 gnd.n6786 gnd.n96 19.3944
R8624 gnd.n7193 gnd.n96 19.3944
R8625 gnd.n7193 gnd.n7192 19.3944
R8626 gnd.n7192 gnd.n7191 19.3944
R8627 gnd.n7191 gnd.n100 19.3944
R8628 gnd.n7181 gnd.n100 19.3944
R8629 gnd.n7181 gnd.n7180 19.3944
R8630 gnd.n7180 gnd.n7179 19.3944
R8631 gnd.n7179 gnd.n118 19.3944
R8632 gnd.n7169 gnd.n118 19.3944
R8633 gnd.n7169 gnd.n7168 19.3944
R8634 gnd.n7168 gnd.n7167 19.3944
R8635 gnd.n7167 gnd.n138 19.3944
R8636 gnd.n7157 gnd.n138 19.3944
R8637 gnd.n7157 gnd.n7156 19.3944
R8638 gnd.n7156 gnd.n7155 19.3944
R8639 gnd.n7155 gnd.n157 19.3944
R8640 gnd.n7145 gnd.n157 19.3944
R8641 gnd.n7007 gnd.n6943 19.3944
R8642 gnd.n7007 gnd.n7004 19.3944
R8643 gnd.n7004 gnd.n7001 19.3944
R8644 gnd.n7001 gnd.n7000 19.3944
R8645 gnd.n7000 gnd.n6997 19.3944
R8646 gnd.n6997 gnd.n6996 19.3944
R8647 gnd.n6996 gnd.n6993 19.3944
R8648 gnd.n6993 gnd.n6992 19.3944
R8649 gnd.n6992 gnd.n6989 19.3944
R8650 gnd.n6989 gnd.n6988 19.3944
R8651 gnd.n6988 gnd.n6985 19.3944
R8652 gnd.n6985 gnd.n6984 19.3944
R8653 gnd.n6984 gnd.n6981 19.3944
R8654 gnd.n6981 gnd.n6980 19.3944
R8655 gnd.n6980 gnd.n6977 19.3944
R8656 gnd.n6977 gnd.n6976 19.3944
R8657 gnd.n6976 gnd.n6973 19.3944
R8658 gnd.n6973 gnd.n6972 19.3944
R8659 gnd.n7050 gnd.n7047 19.3944
R8660 gnd.n7047 gnd.n7046 19.3944
R8661 gnd.n7046 gnd.n7043 19.3944
R8662 gnd.n7043 gnd.n7042 19.3944
R8663 gnd.n7042 gnd.n7039 19.3944
R8664 gnd.n7039 gnd.n7038 19.3944
R8665 gnd.n7038 gnd.n7035 19.3944
R8666 gnd.n7035 gnd.n7034 19.3944
R8667 gnd.n7034 gnd.n7031 19.3944
R8668 gnd.n7031 gnd.n7030 19.3944
R8669 gnd.n7030 gnd.n7027 19.3944
R8670 gnd.n7027 gnd.n7026 19.3944
R8671 gnd.n7026 gnd.n7023 19.3944
R8672 gnd.n7023 gnd.n7022 19.3944
R8673 gnd.n7022 gnd.n7019 19.3944
R8674 gnd.n7019 gnd.n7018 19.3944
R8675 gnd.n7018 gnd.n7015 19.3944
R8676 gnd.n7015 gnd.n7014 19.3944
R8677 gnd.n6905 gnd.n6904 19.3944
R8678 gnd.n7083 gnd.n6904 19.3944
R8679 gnd.n7083 gnd.n7082 19.3944
R8680 gnd.n7082 gnd.n7081 19.3944
R8681 gnd.n7081 gnd.n7078 19.3944
R8682 gnd.n7078 gnd.n7077 19.3944
R8683 gnd.n7077 gnd.n7074 19.3944
R8684 gnd.n7074 gnd.n7073 19.3944
R8685 gnd.n7073 gnd.n7070 19.3944
R8686 gnd.n7070 gnd.n7069 19.3944
R8687 gnd.n7069 gnd.n7066 19.3944
R8688 gnd.n7066 gnd.n7065 19.3944
R8689 gnd.n7065 gnd.n7062 19.3944
R8690 gnd.n7062 gnd.n7061 19.3944
R8691 gnd.n7061 gnd.n7058 19.3944
R8692 gnd.n7058 gnd.n7057 19.3944
R8693 gnd.n7057 gnd.n7054 19.3944
R8694 gnd.n6835 gnd.n6833 19.3944
R8695 gnd.n6838 gnd.n6835 19.3944
R8696 gnd.n6838 gnd.n6830 19.3944
R8697 gnd.n6842 gnd.n6830 19.3944
R8698 gnd.n6845 gnd.n6842 19.3944
R8699 gnd.n6848 gnd.n6845 19.3944
R8700 gnd.n6848 gnd.n6828 19.3944
R8701 gnd.n6852 gnd.n6828 19.3944
R8702 gnd.n6855 gnd.n6852 19.3944
R8703 gnd.n6858 gnd.n6855 19.3944
R8704 gnd.n6858 gnd.n6826 19.3944
R8705 gnd.n6862 gnd.n6826 19.3944
R8706 gnd.n6865 gnd.n6862 19.3944
R8707 gnd.n6867 gnd.n6865 19.3944
R8708 gnd.n6867 gnd.n6824 19.3944
R8709 gnd.n6871 gnd.n6824 19.3944
R8710 gnd.n5216 gnd.n1630 19.3944
R8711 gnd.n5216 gnd.n1631 19.3944
R8712 gnd.n5212 gnd.n1631 19.3944
R8713 gnd.n5212 gnd.n5211 19.3944
R8714 gnd.n5211 gnd.n5210 19.3944
R8715 gnd.n5210 gnd.n5182 19.3944
R8716 gnd.n5206 gnd.n5182 19.3944
R8717 gnd.n5206 gnd.n5205 19.3944
R8718 gnd.n5205 gnd.n5204 19.3944
R8719 gnd.n5204 gnd.n1614 19.3944
R8720 gnd.n5263 gnd.n1614 19.3944
R8721 gnd.n5263 gnd.n1612 19.3944
R8722 gnd.n5267 gnd.n1612 19.3944
R8723 gnd.n5267 gnd.n1609 19.3944
R8724 gnd.n5278 gnd.n1609 19.3944
R8725 gnd.n5278 gnd.n1606 19.3944
R8726 gnd.n5286 gnd.n1606 19.3944
R8727 gnd.n5286 gnd.n1607 19.3944
R8728 gnd.n5282 gnd.n1607 19.3944
R8729 gnd.n5282 gnd.n5281 19.3944
R8730 gnd.n5281 gnd.n68 19.3944
R8731 gnd.n7206 gnd.n68 19.3944
R8732 gnd.n7206 gnd.n7205 19.3944
R8733 gnd.n7205 gnd.n71 19.3944
R8734 gnd.n6793 gnd.n71 19.3944
R8735 gnd.n6793 gnd.n175 19.3944
R8736 gnd.n7114 gnd.n175 19.3944
R8737 gnd.n7114 gnd.n7113 19.3944
R8738 gnd.n7113 gnd.n7112 19.3944
R8739 gnd.n7112 gnd.n7110 19.3944
R8740 gnd.n7110 gnd.n7109 19.3944
R8741 gnd.n7109 gnd.n7107 19.3944
R8742 gnd.n7107 gnd.n7106 19.3944
R8743 gnd.n7106 gnd.n7104 19.3944
R8744 gnd.n7104 gnd.n7103 19.3944
R8745 gnd.n7103 gnd.n7101 19.3944
R8746 gnd.n7101 gnd.n7100 19.3944
R8747 gnd.n7100 gnd.n7098 19.3944
R8748 gnd.n7098 gnd.n7097 19.3944
R8749 gnd.n7097 gnd.n7095 19.3944
R8750 gnd.n7095 gnd.n7094 19.3944
R8751 gnd.n7094 gnd.n7092 19.3944
R8752 gnd.n1500 gnd.n1499 19.3944
R8753 gnd.n5366 gnd.n1499 19.3944
R8754 gnd.n5366 gnd.n5365 19.3944
R8755 gnd.n5365 gnd.n5364 19.3944
R8756 gnd.n5364 gnd.n1506 19.3944
R8757 gnd.n5354 gnd.n1506 19.3944
R8758 gnd.n5354 gnd.n5353 19.3944
R8759 gnd.n5353 gnd.n5352 19.3944
R8760 gnd.n5352 gnd.n1529 19.3944
R8761 gnd.n5342 gnd.n1529 19.3944
R8762 gnd.n5342 gnd.n5341 19.3944
R8763 gnd.n5341 gnd.n5340 19.3944
R8764 gnd.n5340 gnd.n1550 19.3944
R8765 gnd.n5330 gnd.n1550 19.3944
R8766 gnd.n5330 gnd.n5329 19.3944
R8767 gnd.n5329 gnd.n5328 19.3944
R8768 gnd.n5318 gnd.n5317 19.3944
R8769 gnd.n1584 gnd.n1583 19.3944
R8770 gnd.n1594 gnd.n1593 19.3944
R8771 gnd.n7201 gnd.n7200 19.3944
R8772 gnd.n7197 gnd.n80 19.3944
R8773 gnd.n7197 gnd.n87 19.3944
R8774 gnd.n7187 gnd.n87 19.3944
R8775 gnd.n7187 gnd.n7186 19.3944
R8776 gnd.n7186 gnd.n7185 19.3944
R8777 gnd.n7185 gnd.n109 19.3944
R8778 gnd.n7175 gnd.n109 19.3944
R8779 gnd.n7175 gnd.n7174 19.3944
R8780 gnd.n7174 gnd.n7173 19.3944
R8781 gnd.n7173 gnd.n128 19.3944
R8782 gnd.n7163 gnd.n128 19.3944
R8783 gnd.n7163 gnd.n7162 19.3944
R8784 gnd.n7162 gnd.n7161 19.3944
R8785 gnd.n7161 gnd.n148 19.3944
R8786 gnd.n7151 gnd.n148 19.3944
R8787 gnd.n7151 gnd.n7150 19.3944
R8788 gnd.n7150 gnd.n7149 19.3944
R8789 gnd.n5969 gnd.n731 19.3944
R8790 gnd.n4083 gnd.n4082 19.3944
R8791 gnd.n4087 gnd.n4086 19.3944
R8792 gnd.n4120 gnd.n2117 19.3944
R8793 gnd.n4123 gnd.n4122 19.3944
R8794 gnd.n4127 gnd.n4126 19.3944
R8795 gnd.n4150 gnd.n4127 19.3944
R8796 gnd.n4150 gnd.n4149 19.3944
R8797 gnd.n4149 gnd.n4148 19.3944
R8798 gnd.n4148 gnd.n4132 19.3944
R8799 gnd.n4144 gnd.n4132 19.3944
R8800 gnd.n4144 gnd.n4143 19.3944
R8801 gnd.n4143 gnd.n4142 19.3944
R8802 gnd.n4142 gnd.n4140 19.3944
R8803 gnd.n4140 gnd.n2094 19.3944
R8804 gnd.n2094 gnd.n2092 19.3944
R8805 gnd.n4204 gnd.n2092 19.3944
R8806 gnd.n4204 gnd.n2090 19.3944
R8807 gnd.n4208 gnd.n2090 19.3944
R8808 gnd.n4208 gnd.n2088 19.3944
R8809 gnd.n4212 gnd.n2088 19.3944
R8810 gnd.n4212 gnd.n2086 19.3944
R8811 gnd.n4216 gnd.n2086 19.3944
R8812 gnd.n4216 gnd.n2084 19.3944
R8813 gnd.n4221 gnd.n2084 19.3944
R8814 gnd.n4221 gnd.n2082 19.3944
R8815 gnd.n4225 gnd.n2082 19.3944
R8816 gnd.n4225 gnd.n2080 19.3944
R8817 gnd.n4306 gnd.n2080 19.3944
R8818 gnd.n4306 gnd.n2078 19.3944
R8819 gnd.n4310 gnd.n2078 19.3944
R8820 gnd.n4310 gnd.n2065 19.3944
R8821 gnd.n4322 gnd.n2065 19.3944
R8822 gnd.n4322 gnd.n2063 19.3944
R8823 gnd.n4326 gnd.n2063 19.3944
R8824 gnd.n4326 gnd.n2052 19.3944
R8825 gnd.n4338 gnd.n2052 19.3944
R8826 gnd.n4338 gnd.n2050 19.3944
R8827 gnd.n4342 gnd.n2050 19.3944
R8828 gnd.n4342 gnd.n2038 19.3944
R8829 gnd.n4354 gnd.n2038 19.3944
R8830 gnd.n4354 gnd.n2036 19.3944
R8831 gnd.n4358 gnd.n2036 19.3944
R8832 gnd.n4358 gnd.n2024 19.3944
R8833 gnd.n4370 gnd.n2024 19.3944
R8834 gnd.n4370 gnd.n2022 19.3944
R8835 gnd.n4374 gnd.n2022 19.3944
R8836 gnd.n4374 gnd.n2010 19.3944
R8837 gnd.n4386 gnd.n2010 19.3944
R8838 gnd.n4386 gnd.n2008 19.3944
R8839 gnd.n4390 gnd.n2008 19.3944
R8840 gnd.n4390 gnd.n1995 19.3944
R8841 gnd.n4403 gnd.n1995 19.3944
R8842 gnd.n4403 gnd.n1993 19.3944
R8843 gnd.n4413 gnd.n1993 19.3944
R8844 gnd.n4413 gnd.n4412 19.3944
R8845 gnd.n4412 gnd.n4411 19.3944
R8846 gnd.n4411 gnd.n1207 19.3944
R8847 gnd.n5675 gnd.n1207 19.3944
R8848 gnd.n5675 gnd.n5674 19.3944
R8849 gnd.n5674 gnd.n5673 19.3944
R8850 gnd.n5673 gnd.n1211 19.3944
R8851 gnd.n1966 gnd.n1211 19.3944
R8852 gnd.n4561 gnd.n1966 19.3944
R8853 gnd.n4561 gnd.n1963 19.3944
R8854 gnd.n4565 gnd.n1963 19.3944
R8855 gnd.n4565 gnd.n1938 19.3944
R8856 gnd.n4604 gnd.n1938 19.3944
R8857 gnd.n4604 gnd.n1936 19.3944
R8858 gnd.n4610 gnd.n1936 19.3944
R8859 gnd.n4610 gnd.n4609 19.3944
R8860 gnd.n4609 gnd.n1917 19.3944
R8861 gnd.n4664 gnd.n1917 19.3944
R8862 gnd.n4664 gnd.n1915 19.3944
R8863 gnd.n4679 gnd.n1915 19.3944
R8864 gnd.n4679 gnd.n4678 19.3944
R8865 gnd.n4678 gnd.n4677 19.3944
R8866 gnd.n4677 gnd.n4670 19.3944
R8867 gnd.n4673 gnd.n4670 19.3944
R8868 gnd.n4673 gnd.n1880 19.3944
R8869 gnd.n4725 gnd.n1880 19.3944
R8870 gnd.n4725 gnd.n1878 19.3944
R8871 gnd.n4729 gnd.n1878 19.3944
R8872 gnd.n4729 gnd.n1857 19.3944
R8873 gnd.n4771 gnd.n1857 19.3944
R8874 gnd.n4771 gnd.n1855 19.3944
R8875 gnd.n4777 gnd.n1855 19.3944
R8876 gnd.n4777 gnd.n4776 19.3944
R8877 gnd.n4776 gnd.n1836 19.3944
R8878 gnd.n4823 gnd.n1836 19.3944
R8879 gnd.n4823 gnd.n1834 19.3944
R8880 gnd.n4829 gnd.n1834 19.3944
R8881 gnd.n4829 gnd.n4828 19.3944
R8882 gnd.n4828 gnd.n1809 19.3944
R8883 gnd.n4859 gnd.n1809 19.3944
R8884 gnd.n4859 gnd.n1807 19.3944
R8885 gnd.n4863 gnd.n1807 19.3944
R8886 gnd.n4863 gnd.n1753 19.3944
R8887 gnd.n5034 gnd.n1753 19.3944
R8888 gnd.n5034 gnd.n1751 19.3944
R8889 gnd.n5038 gnd.n1751 19.3944
R8890 gnd.n5038 gnd.n1741 19.3944
R8891 gnd.n5050 gnd.n1741 19.3944
R8892 gnd.n5050 gnd.n1739 19.3944
R8893 gnd.n5054 gnd.n1739 19.3944
R8894 gnd.n5054 gnd.n1728 19.3944
R8895 gnd.n5067 gnd.n1728 19.3944
R8896 gnd.n5067 gnd.n1726 19.3944
R8897 gnd.n5071 gnd.n1726 19.3944
R8898 gnd.n5071 gnd.n1716 19.3944
R8899 gnd.n5083 gnd.n1716 19.3944
R8900 gnd.n5083 gnd.n1714 19.3944
R8901 gnd.n5087 gnd.n1714 19.3944
R8902 gnd.n5087 gnd.n1703 19.3944
R8903 gnd.n5099 gnd.n1703 19.3944
R8904 gnd.n5099 gnd.n1701 19.3944
R8905 gnd.n5103 gnd.n1701 19.3944
R8906 gnd.n5103 gnd.n1690 19.3944
R8907 gnd.n5115 gnd.n1690 19.3944
R8908 gnd.n5115 gnd.n1688 19.3944
R8909 gnd.n5119 gnd.n1688 19.3944
R8910 gnd.n5119 gnd.n1677 19.3944
R8911 gnd.n5131 gnd.n1677 19.3944
R8912 gnd.n5131 gnd.n1675 19.3944
R8913 gnd.n5138 gnd.n1675 19.3944
R8914 gnd.n5138 gnd.n5137 19.3944
R8915 gnd.n5137 gnd.n1664 19.3944
R8916 gnd.n5151 gnd.n1664 19.3944
R8917 gnd.n5152 gnd.n5151 19.3944
R8918 gnd.n5152 gnd.n1662 19.3944
R8919 gnd.n5167 gnd.n1662 19.3944
R8920 gnd.n5167 gnd.n5166 19.3944
R8921 gnd.n5166 gnd.n5165 19.3944
R8922 gnd.n5165 gnd.n5158 19.3944
R8923 gnd.n5161 gnd.n5158 19.3944
R8924 gnd.n5161 gnd.n1628 19.3944
R8925 gnd.n5221 gnd.n1628 19.3944
R8926 gnd.n5221 gnd.n1626 19.3944
R8927 gnd.n5225 gnd.n1626 19.3944
R8928 gnd.n5225 gnd.n1624 19.3944
R8929 gnd.n5229 gnd.n1624 19.3944
R8930 gnd.n5229 gnd.n1622 19.3944
R8931 gnd.n5233 gnd.n1622 19.3944
R8932 gnd.n5233 gnd.n1620 19.3944
R8933 gnd.n5237 gnd.n1620 19.3944
R8934 gnd.n5237 gnd.n1618 19.3944
R8935 gnd.n5258 gnd.n1618 19.3944
R8936 gnd.n5258 gnd.n5257 19.3944
R8937 gnd.n5257 gnd.n5256 19.3944
R8938 gnd.n5256 gnd.n5243 19.3944
R8939 gnd.n5252 gnd.n5243 19.3944
R8940 gnd.n5252 gnd.n5251 19.3944
R8941 gnd.n5249 gnd.n5247 19.3944
R8942 gnd.n5312 gnd.n5311 19.3944
R8943 gnd.n5309 gnd.n1591 19.3944
R8944 gnd.n6781 gnd.n183 19.3944
R8945 gnd.n6779 gnd.n6778 19.3944
R8946 gnd.n3956 gnd.n3955 19.3944
R8947 gnd.n3955 gnd.n3747 19.3944
R8948 gnd.n3950 gnd.n3747 19.3944
R8949 gnd.n3950 gnd.n3949 19.3944
R8950 gnd.n3949 gnd.n3752 19.3944
R8951 gnd.n3944 gnd.n3752 19.3944
R8952 gnd.n3944 gnd.n3943 19.3944
R8953 gnd.n3943 gnd.n3942 19.3944
R8954 gnd.n3942 gnd.n3758 19.3944
R8955 gnd.n3936 gnd.n3758 19.3944
R8956 gnd.n3936 gnd.n3935 19.3944
R8957 gnd.n3935 gnd.n3934 19.3944
R8958 gnd.n3934 gnd.n3764 19.3944
R8959 gnd.n3928 gnd.n3764 19.3944
R8960 gnd.n3928 gnd.n3927 19.3944
R8961 gnd.n3927 gnd.n3926 19.3944
R8962 gnd.n3926 gnd.n3770 19.3944
R8963 gnd.n3920 gnd.n3919 19.3944
R8964 gnd.n3919 gnd.n3918 19.3944
R8965 gnd.n3918 gnd.n3779 19.3944
R8966 gnd.n3912 gnd.n3779 19.3944
R8967 gnd.n3912 gnd.n3911 19.3944
R8968 gnd.n3911 gnd.n3910 19.3944
R8969 gnd.n3910 gnd.n3785 19.3944
R8970 gnd.n3904 gnd.n3785 19.3944
R8971 gnd.n3904 gnd.n3903 19.3944
R8972 gnd.n3903 gnd.n3902 19.3944
R8973 gnd.n3902 gnd.n3791 19.3944
R8974 gnd.n3896 gnd.n3791 19.3944
R8975 gnd.n3896 gnd.n3895 19.3944
R8976 gnd.n3895 gnd.n3894 19.3944
R8977 gnd.n3894 gnd.n3797 19.3944
R8978 gnd.n3888 gnd.n3797 19.3944
R8979 gnd.n3888 gnd.n3887 19.3944
R8980 gnd.n3887 gnd.n3886 19.3944
R8981 gnd.n3880 gnd.n3879 19.3944
R8982 gnd.n3879 gnd.n3878 19.3944
R8983 gnd.n3878 gnd.n3811 19.3944
R8984 gnd.n3872 gnd.n3811 19.3944
R8985 gnd.n3872 gnd.n3871 19.3944
R8986 gnd.n3871 gnd.n3870 19.3944
R8987 gnd.n3870 gnd.n3817 19.3944
R8988 gnd.n3864 gnd.n3817 19.3944
R8989 gnd.n3864 gnd.n3863 19.3944
R8990 gnd.n3863 gnd.n3862 19.3944
R8991 gnd.n3862 gnd.n3823 19.3944
R8992 gnd.n3856 gnd.n3823 19.3944
R8993 gnd.n3856 gnd.n3855 19.3944
R8994 gnd.n3855 gnd.n3854 19.3944
R8995 gnd.n3854 gnd.n3829 19.3944
R8996 gnd.n3848 gnd.n3829 19.3944
R8997 gnd.n3848 gnd.n3847 19.3944
R8998 gnd.n3847 gnd.n3846 19.3944
R8999 gnd.n3692 gnd.n3691 19.3944
R9000 gnd.n3697 gnd.n3692 19.3944
R9001 gnd.n3697 gnd.n3688 19.3944
R9002 gnd.n3701 gnd.n3688 19.3944
R9003 gnd.n3701 gnd.n3686 19.3944
R9004 gnd.n3707 gnd.n3686 19.3944
R9005 gnd.n3707 gnd.n3684 19.3944
R9006 gnd.n3711 gnd.n3684 19.3944
R9007 gnd.n3711 gnd.n3682 19.3944
R9008 gnd.n3717 gnd.n3682 19.3944
R9009 gnd.n3717 gnd.n3680 19.3944
R9010 gnd.n3721 gnd.n3680 19.3944
R9011 gnd.n3721 gnd.n3678 19.3944
R9012 gnd.n3727 gnd.n3678 19.3944
R9013 gnd.n3727 gnd.n3676 19.3944
R9014 gnd.n3731 gnd.n3676 19.3944
R9015 gnd.n3742 gnd.n3670 19.3944
R9016 gnd.n3742 gnd.n3741 19.3944
R9017 gnd.n3741 gnd.n2183 19.3944
R9018 gnd.n3991 gnd.n2183 19.3944
R9019 gnd.n3991 gnd.n2181 19.3944
R9020 gnd.n3997 gnd.n2181 19.3944
R9021 gnd.n3997 gnd.n3996 19.3944
R9022 gnd.n3996 gnd.n2158 19.3944
R9023 gnd.n4026 gnd.n2158 19.3944
R9024 gnd.n4026 gnd.n2156 19.3944
R9025 gnd.n4034 gnd.n2156 19.3944
R9026 gnd.n4034 gnd.n4033 19.3944
R9027 gnd.n4033 gnd.n4032 19.3944
R9028 gnd.n4032 gnd.n2132 19.3944
R9029 gnd.n4066 gnd.n2132 19.3944
R9030 gnd.n4066 gnd.n2130 19.3944
R9031 gnd.n4070 gnd.n2130 19.3944
R9032 gnd.n4070 gnd.n2127 19.3944
R9033 gnd.n4092 gnd.n2127 19.3944
R9034 gnd.n4092 gnd.n2125 19.3944
R9035 gnd.n4096 gnd.n2125 19.3944
R9036 gnd.n4096 gnd.n2120 19.3944
R9037 gnd.n4115 gnd.n2120 19.3944
R9038 gnd.n4115 gnd.n2121 19.3944
R9039 gnd.n4111 gnd.n2121 19.3944
R9040 gnd.n4111 gnd.n2111 19.3944
R9041 gnd.n4155 gnd.n2111 19.3944
R9042 gnd.n4155 gnd.n2109 19.3944
R9043 gnd.n4159 gnd.n2109 19.3944
R9044 gnd.n4159 gnd.n2105 19.3944
R9045 gnd.n4169 gnd.n2105 19.3944
R9046 gnd.n4169 gnd.n2103 19.3944
R9047 gnd.n4173 gnd.n2103 19.3944
R9048 gnd.n4173 gnd.n2096 19.3944
R9049 gnd.n4197 gnd.n2096 19.3944
R9050 gnd.n4197 gnd.n2097 19.3944
R9051 gnd.n4193 gnd.n2097 19.3944
R9052 gnd.n4193 gnd.n4192 19.3944
R9053 gnd.n4192 gnd.n4191 19.3944
R9054 gnd.n4191 gnd.n868 19.3944
R9055 gnd.n5876 gnd.n868 19.3944
R9056 gnd.n5876 gnd.n869 19.3944
R9057 gnd.n3966 gnd.n2201 19.3944
R9058 gnd.n3967 gnd.n3966 19.3944
R9059 gnd.n3969 gnd.n3967 19.3944
R9060 gnd.n3970 gnd.n3969 19.3944
R9061 gnd.n3970 gnd.n2176 19.3944
R9062 gnd.n4001 gnd.n2176 19.3944
R9063 gnd.n4002 gnd.n4001 19.3944
R9064 gnd.n4004 gnd.n4002 19.3944
R9065 gnd.n4005 gnd.n4004 19.3944
R9066 gnd.n4005 gnd.n2151 19.3944
R9067 gnd.n4038 gnd.n2151 19.3944
R9068 gnd.n4039 gnd.n4038 19.3944
R9069 gnd.n4041 gnd.n4039 19.3944
R9070 gnd.n4042 gnd.n4041 19.3944
R9071 gnd.n4044 gnd.n4042 19.3944
R9072 gnd.n4044 gnd.n2128 19.3944
R9073 gnd.n4074 gnd.n2128 19.3944
R9074 gnd.n4075 gnd.n4074 19.3944
R9075 gnd.n4076 gnd.n4075 19.3944
R9076 gnd.n4076 gnd.n2123 19.3944
R9077 gnd.n4100 gnd.n2123 19.3944
R9078 gnd.n4101 gnd.n4100 19.3944
R9079 gnd.n4102 gnd.n4101 19.3944
R9080 gnd.n4103 gnd.n4102 19.3944
R9081 gnd.n4107 gnd.n4103 19.3944
R9082 gnd.n4107 gnd.n4106 19.3944
R9083 gnd.n4106 gnd.n4105 19.3944
R9084 gnd.n4105 gnd.n2107 19.3944
R9085 gnd.n4163 gnd.n2107 19.3944
R9086 gnd.n4164 gnd.n4163 19.3944
R9087 gnd.n4165 gnd.n4164 19.3944
R9088 gnd.n4165 gnd.n2101 19.3944
R9089 gnd.n4177 gnd.n2101 19.3944
R9090 gnd.n4178 gnd.n4177 19.3944
R9091 gnd.n4179 gnd.n4178 19.3944
R9092 gnd.n4180 gnd.n4179 19.3944
R9093 gnd.n4184 gnd.n4180 19.3944
R9094 gnd.n4185 gnd.n4184 19.3944
R9095 gnd.n4186 gnd.n4185 19.3944
R9096 gnd.n4186 gnd.n866 19.3944
R9097 gnd.n5880 gnd.n866 19.3944
R9098 gnd.n5881 gnd.n5880 19.3944
R9099 gnd.n3963 gnd.n2198 19.3944
R9100 gnd.n3977 gnd.n2198 19.3944
R9101 gnd.n3977 gnd.n3976 19.3944
R9102 gnd.n3976 gnd.n3975 19.3944
R9103 gnd.n3975 gnd.n3974 19.3944
R9104 gnd.n3974 gnd.n2173 19.3944
R9105 gnd.n4012 gnd.n2173 19.3944
R9106 gnd.n4012 gnd.n4011 19.3944
R9107 gnd.n4011 gnd.n4010 19.3944
R9108 gnd.n4010 gnd.n4009 19.3944
R9109 gnd.n4009 gnd.n2147 19.3944
R9110 gnd.n4052 gnd.n2147 19.3944
R9111 gnd.n4052 gnd.n4051 19.3944
R9112 gnd.n4051 gnd.n4050 19.3944
R9113 gnd.n4050 gnd.n4049 19.3944
R9114 gnd.n4049 gnd.n4047 19.3944
R9115 gnd.n4047 gnd.n750 19.3944
R9116 gnd.n5957 gnd.n750 19.3944
R9117 gnd.n5957 gnd.n5956 19.3944
R9118 gnd.n5956 gnd.n5955 19.3944
R9119 gnd.n5955 gnd.n754 19.3944
R9120 gnd.n5944 gnd.n754 19.3944
R9121 gnd.n5944 gnd.n5943 19.3944
R9122 gnd.n5943 gnd.n5942 19.3944
R9123 gnd.n5942 gnd.n770 19.3944
R9124 gnd.n5931 gnd.n770 19.3944
R9125 gnd.n5931 gnd.n5930 19.3944
R9126 gnd.n5930 gnd.n5929 19.3944
R9127 gnd.n5929 gnd.n788 19.3944
R9128 gnd.n5919 gnd.n788 19.3944
R9129 gnd.n5919 gnd.n5918 19.3944
R9130 gnd.n5918 gnd.n5917 19.3944
R9131 gnd.n5917 gnd.n807 19.3944
R9132 gnd.n5907 gnd.n807 19.3944
R9133 gnd.n5907 gnd.n5906 19.3944
R9134 gnd.n5906 gnd.n5905 19.3944
R9135 gnd.n5905 gnd.n828 19.3944
R9136 gnd.n5895 gnd.n828 19.3944
R9137 gnd.n5895 gnd.n5894 19.3944
R9138 gnd.n5894 gnd.n5893 19.3944
R9139 gnd.n5893 gnd.n848 19.3944
R9140 gnd.n5883 gnd.n848 19.3944
R9141 gnd.n1011 gnd.n1010 19.3944
R9142 gnd.n5799 gnd.n1010 19.3944
R9143 gnd.n5799 gnd.n5798 19.3944
R9144 gnd.n5798 gnd.n5797 19.3944
R9145 gnd.n5797 gnd.n5794 19.3944
R9146 gnd.n5794 gnd.n5793 19.3944
R9147 gnd.n5793 gnd.n5790 19.3944
R9148 gnd.n5790 gnd.n5789 19.3944
R9149 gnd.n5789 gnd.n5786 19.3944
R9150 gnd.n5786 gnd.n5785 19.3944
R9151 gnd.n5785 gnd.n5782 19.3944
R9152 gnd.n5782 gnd.n5781 19.3944
R9153 gnd.n5781 gnd.n5778 19.3944
R9154 gnd.n5778 gnd.n5777 19.3944
R9155 gnd.n5777 gnd.n5774 19.3944
R9156 gnd.n5774 gnd.n5773 19.3944
R9157 gnd.n5773 gnd.n5770 19.3944
R9158 gnd.n1113 gnd.n1049 19.3944
R9159 gnd.n1113 gnd.n1110 19.3944
R9160 gnd.n1110 gnd.n1107 19.3944
R9161 gnd.n1107 gnd.n1106 19.3944
R9162 gnd.n1106 gnd.n1103 19.3944
R9163 gnd.n1103 gnd.n1102 19.3944
R9164 gnd.n1102 gnd.n1099 19.3944
R9165 gnd.n1099 gnd.n1098 19.3944
R9166 gnd.n1098 gnd.n1095 19.3944
R9167 gnd.n1095 gnd.n1094 19.3944
R9168 gnd.n1094 gnd.n1091 19.3944
R9169 gnd.n1091 gnd.n1090 19.3944
R9170 gnd.n1090 gnd.n1087 19.3944
R9171 gnd.n1087 gnd.n1086 19.3944
R9172 gnd.n1086 gnd.n1083 19.3944
R9173 gnd.n1083 gnd.n1082 19.3944
R9174 gnd.n1082 gnd.n1079 19.3944
R9175 gnd.n1079 gnd.n1078 19.3944
R9176 gnd.n1135 gnd.n1040 19.3944
R9177 gnd.n1135 gnd.n1132 19.3944
R9178 gnd.n1132 gnd.n1129 19.3944
R9179 gnd.n1129 gnd.n1128 19.3944
R9180 gnd.n1128 gnd.n1125 19.3944
R9181 gnd.n1125 gnd.n1124 19.3944
R9182 gnd.n1124 gnd.n1121 19.3944
R9183 gnd.n1121 gnd.n1120 19.3944
R9184 gnd.n5768 gnd.n5765 19.3944
R9185 gnd.n5765 gnd.n5764 19.3944
R9186 gnd.n5764 gnd.n5761 19.3944
R9187 gnd.n5761 gnd.n5760 19.3944
R9188 gnd.n5760 gnd.n5757 19.3944
R9189 gnd.n5757 gnd.n5756 19.3944
R9190 gnd.n5756 gnd.n5753 19.3944
R9191 gnd.n3959 gnd.n2192 19.3944
R9192 gnd.n3981 gnd.n2192 19.3944
R9193 gnd.n3981 gnd.n2190 19.3944
R9194 gnd.n3987 gnd.n2190 19.3944
R9195 gnd.n3987 gnd.n3986 19.3944
R9196 gnd.n3986 gnd.n2167 19.3944
R9197 gnd.n4016 gnd.n2167 19.3944
R9198 gnd.n4016 gnd.n2165 19.3944
R9199 gnd.n4022 gnd.n2165 19.3944
R9200 gnd.n4022 gnd.n4021 19.3944
R9201 gnd.n4021 gnd.n2140 19.3944
R9202 gnd.n4056 gnd.n2140 19.3944
R9203 gnd.n4056 gnd.n2138 19.3944
R9204 gnd.n4061 gnd.n2138 19.3944
R9205 gnd.n4061 gnd.n740 19.3944
R9206 gnd.n5964 gnd.n740 19.3944
R9207 gnd.n5962 gnd.n5961 19.3944
R9208 gnd.n5951 gnd.n760 19.3944
R9209 gnd.n5949 gnd.n5948 19.3944
R9210 gnd.n5938 gnd.n777 19.3944
R9211 gnd.n5936 gnd.n5935 19.3944
R9212 gnd.n5935 gnd.n778 19.3944
R9213 gnd.n5925 gnd.n778 19.3944
R9214 gnd.n5925 gnd.n5924 19.3944
R9215 gnd.n5924 gnd.n5923 19.3944
R9216 gnd.n5923 gnd.n798 19.3944
R9217 gnd.n5913 gnd.n798 19.3944
R9218 gnd.n5913 gnd.n5912 19.3944
R9219 gnd.n5912 gnd.n5911 19.3944
R9220 gnd.n5911 gnd.n818 19.3944
R9221 gnd.n5901 gnd.n818 19.3944
R9222 gnd.n5901 gnd.n5900 19.3944
R9223 gnd.n5900 gnd.n5899 19.3944
R9224 gnd.n5899 gnd.n838 19.3944
R9225 gnd.n5889 gnd.n838 19.3944
R9226 gnd.n5889 gnd.n5888 19.3944
R9227 gnd.n5888 gnd.n5887 19.3944
R9228 gnd.n6140 gnd.n6139 19.3944
R9229 gnd.n6139 gnd.n564 19.3944
R9230 gnd.n6133 gnd.n564 19.3944
R9231 gnd.n6133 gnd.n6132 19.3944
R9232 gnd.n6132 gnd.n6131 19.3944
R9233 gnd.n6131 gnd.n572 19.3944
R9234 gnd.n6125 gnd.n572 19.3944
R9235 gnd.n6125 gnd.n6124 19.3944
R9236 gnd.n6124 gnd.n6123 19.3944
R9237 gnd.n6123 gnd.n580 19.3944
R9238 gnd.n6117 gnd.n580 19.3944
R9239 gnd.n6117 gnd.n6116 19.3944
R9240 gnd.n6116 gnd.n6115 19.3944
R9241 gnd.n6115 gnd.n588 19.3944
R9242 gnd.n6109 gnd.n588 19.3944
R9243 gnd.n6109 gnd.n6108 19.3944
R9244 gnd.n6108 gnd.n6107 19.3944
R9245 gnd.n6107 gnd.n596 19.3944
R9246 gnd.n6101 gnd.n596 19.3944
R9247 gnd.n6101 gnd.n6100 19.3944
R9248 gnd.n6100 gnd.n6099 19.3944
R9249 gnd.n6099 gnd.n604 19.3944
R9250 gnd.n6093 gnd.n604 19.3944
R9251 gnd.n6093 gnd.n6092 19.3944
R9252 gnd.n6092 gnd.n6091 19.3944
R9253 gnd.n6091 gnd.n612 19.3944
R9254 gnd.n6085 gnd.n612 19.3944
R9255 gnd.n6085 gnd.n6084 19.3944
R9256 gnd.n6084 gnd.n6083 19.3944
R9257 gnd.n6083 gnd.n620 19.3944
R9258 gnd.n6077 gnd.n620 19.3944
R9259 gnd.n6077 gnd.n6076 19.3944
R9260 gnd.n6076 gnd.n6075 19.3944
R9261 gnd.n6075 gnd.n628 19.3944
R9262 gnd.n6069 gnd.n628 19.3944
R9263 gnd.n6069 gnd.n6068 19.3944
R9264 gnd.n6068 gnd.n6067 19.3944
R9265 gnd.n6067 gnd.n636 19.3944
R9266 gnd.n6061 gnd.n636 19.3944
R9267 gnd.n6061 gnd.n6060 19.3944
R9268 gnd.n6060 gnd.n6059 19.3944
R9269 gnd.n6059 gnd.n644 19.3944
R9270 gnd.n6053 gnd.n644 19.3944
R9271 gnd.n6053 gnd.n6052 19.3944
R9272 gnd.n6052 gnd.n6051 19.3944
R9273 gnd.n6051 gnd.n652 19.3944
R9274 gnd.n6045 gnd.n652 19.3944
R9275 gnd.n6045 gnd.n6044 19.3944
R9276 gnd.n6044 gnd.n6043 19.3944
R9277 gnd.n6043 gnd.n660 19.3944
R9278 gnd.n6037 gnd.n660 19.3944
R9279 gnd.n6037 gnd.n6036 19.3944
R9280 gnd.n6036 gnd.n6035 19.3944
R9281 gnd.n6035 gnd.n668 19.3944
R9282 gnd.n6029 gnd.n668 19.3944
R9283 gnd.n6029 gnd.n6028 19.3944
R9284 gnd.n6028 gnd.n6027 19.3944
R9285 gnd.n6027 gnd.n676 19.3944
R9286 gnd.n6021 gnd.n676 19.3944
R9287 gnd.n6021 gnd.n6020 19.3944
R9288 gnd.n6020 gnd.n6019 19.3944
R9289 gnd.n6019 gnd.n684 19.3944
R9290 gnd.n6013 gnd.n684 19.3944
R9291 gnd.n6013 gnd.n6012 19.3944
R9292 gnd.n6012 gnd.n6011 19.3944
R9293 gnd.n6011 gnd.n692 19.3944
R9294 gnd.n6005 gnd.n692 19.3944
R9295 gnd.n6005 gnd.n6004 19.3944
R9296 gnd.n6004 gnd.n6003 19.3944
R9297 gnd.n6003 gnd.n700 19.3944
R9298 gnd.n5997 gnd.n700 19.3944
R9299 gnd.n5997 gnd.n5996 19.3944
R9300 gnd.n5996 gnd.n5995 19.3944
R9301 gnd.n5995 gnd.n708 19.3944
R9302 gnd.n5989 gnd.n708 19.3944
R9303 gnd.n5989 gnd.n5988 19.3944
R9304 gnd.n5988 gnd.n5987 19.3944
R9305 gnd.n5987 gnd.n716 19.3944
R9306 gnd.n5981 gnd.n716 19.3944
R9307 gnd.n5981 gnd.n5980 19.3944
R9308 gnd.n5980 gnd.n5979 19.3944
R9309 gnd.n5979 gnd.n724 19.3944
R9310 gnd.n5973 gnd.n724 19.3944
R9311 gnd.n5973 gnd.n5972 19.3944
R9312 gnd.n4297 gnd.n4230 19.3944
R9313 gnd.n4297 gnd.n4231 19.3944
R9314 gnd.n4293 gnd.n4231 19.3944
R9315 gnd.n4293 gnd.n4292 19.3944
R9316 gnd.n4292 gnd.n4291 19.3944
R9317 gnd.n4291 gnd.n4236 19.3944
R9318 gnd.n4287 gnd.n4236 19.3944
R9319 gnd.n4287 gnd.n4286 19.3944
R9320 gnd.n4286 gnd.n4285 19.3944
R9321 gnd.n4285 gnd.n4240 19.3944
R9322 gnd.n4281 gnd.n4240 19.3944
R9323 gnd.n4281 gnd.n4280 19.3944
R9324 gnd.n4280 gnd.n4279 19.3944
R9325 gnd.n4279 gnd.n4244 19.3944
R9326 gnd.n4275 gnd.n4244 19.3944
R9327 gnd.n4275 gnd.n4274 19.3944
R9328 gnd.n4274 gnd.n4273 19.3944
R9329 gnd.n4273 gnd.n4248 19.3944
R9330 gnd.n4269 gnd.n4248 19.3944
R9331 gnd.n4269 gnd.n4268 19.3944
R9332 gnd.n4268 gnd.n4267 19.3944
R9333 gnd.n4267 gnd.n4252 19.3944
R9334 gnd.n4263 gnd.n4252 19.3944
R9335 gnd.n4263 gnd.n4262 19.3944
R9336 gnd.n4262 gnd.n4261 19.3944
R9337 gnd.n4261 gnd.n4256 19.3944
R9338 gnd.n4257 gnd.n4256 19.3944
R9339 gnd.n4257 gnd.n1981 19.3944
R9340 gnd.n4428 gnd.n1981 19.3944
R9341 gnd.n4428 gnd.n1979 19.3944
R9342 gnd.n4432 gnd.n1979 19.3944
R9343 gnd.n4532 gnd.n4432 19.3944
R9344 gnd.n4533 gnd.n4532 19.3944
R9345 gnd.n4533 gnd.n1976 19.3944
R9346 gnd.n4549 gnd.n1976 19.3944
R9347 gnd.n4549 gnd.n1977 19.3944
R9348 gnd.n4545 gnd.n1977 19.3944
R9349 gnd.n4545 gnd.n4544 19.3944
R9350 gnd.n4544 gnd.n4543 19.3944
R9351 gnd.n4543 gnd.n4540 19.3944
R9352 gnd.n4540 gnd.n1930 19.3944
R9353 gnd.n4614 gnd.n1930 19.3944
R9354 gnd.n4614 gnd.n1927 19.3944
R9355 gnd.n4652 gnd.n1927 19.3944
R9356 gnd.n4652 gnd.n1928 19.3944
R9357 gnd.n4648 gnd.n1928 19.3944
R9358 gnd.n4648 gnd.n4647 19.3944
R9359 gnd.n4647 gnd.n4646 19.3944
R9360 gnd.n4646 gnd.n4620 19.3944
R9361 gnd.n4642 gnd.n4620 19.3944
R9362 gnd.n4642 gnd.n4641 19.3944
R9363 gnd.n4641 gnd.n4640 19.3944
R9364 gnd.n4640 gnd.n4625 19.3944
R9365 gnd.n4636 gnd.n4625 19.3944
R9366 gnd.n4636 gnd.n4635 19.3944
R9367 gnd.n4635 gnd.n4634 19.3944
R9368 gnd.n4634 gnd.n4631 19.3944
R9369 gnd.n4631 gnd.n1850 19.3944
R9370 gnd.n4781 gnd.n1850 19.3944
R9371 gnd.n4781 gnd.n1847 19.3944
R9372 gnd.n4810 gnd.n1847 19.3944
R9373 gnd.n4810 gnd.n1848 19.3944
R9374 gnd.n4806 gnd.n1848 19.3944
R9375 gnd.n4806 gnd.n4805 19.3944
R9376 gnd.n4805 gnd.n4804 19.3944
R9377 gnd.n4804 gnd.n4788 19.3944
R9378 gnd.n4800 gnd.n4788 19.3944
R9379 gnd.n4800 gnd.n4799 19.3944
R9380 gnd.n4799 gnd.n4798 19.3944
R9381 gnd.n4798 gnd.n4793 19.3944
R9382 gnd.n4794 gnd.n4793 19.3944
R9383 gnd.n4794 gnd.n1748 19.3944
R9384 gnd.n5042 gnd.n1748 19.3944
R9385 gnd.n5042 gnd.n1746 19.3944
R9386 gnd.n5046 gnd.n1746 19.3944
R9387 gnd.n5046 gnd.n1735 19.3944
R9388 gnd.n5058 gnd.n1735 19.3944
R9389 gnd.n5058 gnd.n1733 19.3944
R9390 gnd.n5062 gnd.n1733 19.3944
R9391 gnd.n5062 gnd.n1723 19.3944
R9392 gnd.n5075 gnd.n1723 19.3944
R9393 gnd.n5075 gnd.n1721 19.3944
R9394 gnd.n5079 gnd.n1721 19.3944
R9395 gnd.n5079 gnd.n1710 19.3944
R9396 gnd.n5091 gnd.n1710 19.3944
R9397 gnd.n5091 gnd.n1708 19.3944
R9398 gnd.n5095 gnd.n1708 19.3944
R9399 gnd.n5095 gnd.n1697 19.3944
R9400 gnd.n5107 gnd.n1697 19.3944
R9401 gnd.n5107 gnd.n1695 19.3944
R9402 gnd.n5111 gnd.n1695 19.3944
R9403 gnd.n5111 gnd.n1682 19.3944
R9404 gnd.n5123 gnd.n1682 19.3944
R9405 gnd.n5123 gnd.n1680 19.3944
R9406 gnd.n5127 gnd.n1680 19.3944
R9407 gnd.n5127 gnd.n1671 19.3944
R9408 gnd.n5142 gnd.n1671 19.3944
R9409 gnd.n5142 gnd.n1669 19.3944
R9410 gnd.n5146 gnd.n1669 19.3944
R9411 gnd.n5146 gnd.n1310 19.3944
R9412 gnd.n5563 gnd.n1310 19.3944
R9413 gnd.n5560 gnd.n5559 19.3944
R9414 gnd.n5559 gnd.n5558 19.3944
R9415 gnd.n5558 gnd.n1315 19.3944
R9416 gnd.n5554 gnd.n1315 19.3944
R9417 gnd.n5554 gnd.n5553 19.3944
R9418 gnd.n5553 gnd.n5552 19.3944
R9419 gnd.n5552 gnd.n1320 19.3944
R9420 gnd.n5547 gnd.n1320 19.3944
R9421 gnd.n5547 gnd.n5546 19.3944
R9422 gnd.n5546 gnd.n1325 19.3944
R9423 gnd.n5539 gnd.n1325 19.3944
R9424 gnd.n5539 gnd.n5538 19.3944
R9425 gnd.n5538 gnd.n1334 19.3944
R9426 gnd.n5531 gnd.n1334 19.3944
R9427 gnd.n5531 gnd.n5530 19.3944
R9428 gnd.n5530 gnd.n1342 19.3944
R9429 gnd.n5523 gnd.n1342 19.3944
R9430 gnd.n5523 gnd.n5522 19.3944
R9431 gnd.n5522 gnd.n1350 19.3944
R9432 gnd.n5515 gnd.n1350 19.3944
R9433 gnd.n5515 gnd.n5514 19.3944
R9434 gnd.n5514 gnd.n1358 19.3944
R9435 gnd.n5507 gnd.n1358 19.3944
R9436 gnd.n5507 gnd.n5506 19.3944
R9437 gnd.n1656 gnd.n1635 19.3944
R9438 gnd.n5174 gnd.n1635 19.3944
R9439 gnd.n5174 gnd.n5173 19.3944
R9440 gnd.n5967 gnd.n733 19.1199
R9441 gnd.n5966 gnd.n736 19.1199
R9442 gnd.n5959 gnd.n747 19.1199
R9443 gnd.n4090 gnd.n4089 19.1199
R9444 gnd.n5953 gnd.n758 19.1199
R9445 gnd.n4098 gnd.n763 19.1199
R9446 gnd.n4117 gnd.n772 19.1199
R9447 gnd.n5940 gnd.n775 19.1199
R9448 gnd.n4109 gnd.n780 19.1199
R9449 gnd.n5933 gnd.n783 19.1199
R9450 gnd.n4153 gnd.n4152 19.1199
R9451 gnd.n5927 gnd.n792 19.1199
R9452 gnd.n4161 gnd.n800 19.1199
R9453 gnd.n4167 gnd.n809 19.1199
R9454 gnd.n5915 gnd.n812 19.1199
R9455 gnd.n4175 gnd.n820 19.1199
R9456 gnd.n5909 gnd.n823 19.1199
R9457 gnd.n4200 gnd.n4199 19.1199
R9458 gnd.n5903 gnd.n832 19.1199
R9459 gnd.n4182 gnd.n840 19.1199
R9460 gnd.n5897 gnd.n843 19.1199
R9461 gnd.n4188 gnd.n850 19.1199
R9462 gnd.n5878 gnd.n859 19.1199
R9463 gnd.n5885 gnd.n862 19.1199
R9464 gnd.n5376 gnd.n1484 19.1199
R9465 gnd.n5218 gnd.n1486 19.1199
R9466 gnd.n5179 gnd.n1495 19.1199
R9467 gnd.n5362 gnd.n1508 19.1199
R9468 gnd.n5186 gnd.n1511 19.1199
R9469 gnd.n5356 gnd.n1521 19.1199
R9470 gnd.n5192 gnd.n5191 19.1199
R9471 gnd.n5350 gnd.n1531 19.1199
R9472 gnd.n5201 gnd.n1534 19.1199
R9473 gnd.n5344 gnd.n1541 19.1199
R9474 gnd.n5261 gnd.n1544 19.1199
R9475 gnd.n5269 gnd.n1554 19.1199
R9476 gnd.n5332 gnd.n1561 19.1199
R9477 gnd.n5276 gnd.n1610 19.1199
R9478 gnd.n5326 gnd.n1568 19.1199
R9479 gnd.n5288 gnd.n1571 19.1199
R9480 gnd.n5320 gnd.n1578 19.1199
R9481 gnd.n5315 gnd.n1581 19.1199
R9482 gnd.n1604 gnd.n1596 19.1199
R9483 gnd.n5307 gnd.n5306 19.1199
R9484 gnd.n7203 gnd.n73 19.1199
R9485 gnd.n6784 gnd.n75 19.1199
R9486 gnd.n7195 gnd.n90 19.1199
R9487 gnd.n7116 gnd.n93 19.1199
R9488 gnd.n3053 gnd.t140 18.8012
R9489 gnd.n3038 gnd.t181 18.8012
R9490 gnd.t221 gnd.n744 18.8012
R9491 gnd.n6783 gnd.t225 18.8012
R9492 gnd.n2897 gnd.n2896 18.4825
R9493 gnd.n4568 gnd.n1957 18.4825
R9494 gnd.n4832 gnd.n4831 18.4825
R9495 gnd.n5445 gnd.n5444 18.4247
R9496 gnd.n5753 gnd.n5752 18.4247
R9497 gnd.n5503 gnd.n5502 18.2308
R9498 gnd.n5807 gnd.n5806 18.2308
R9499 gnd.n6871 gnd.n6814 18.2308
R9500 gnd.n3731 gnd.n3674 18.2308
R9501 gnd.t122 gnd.n2577 18.1639
R9502 gnd.n2605 gnd.t187 17.5266
R9503 gnd.n4589 gnd.t136 17.5266
R9504 gnd.n4745 gnd.t141 17.5266
R9505 gnd.n4530 gnd.t87 17.2079
R9506 gnd.n4551 gnd.n1968 17.2079
R9507 gnd.n3004 gnd.t156 16.8893
R9508 gnd.n3744 gnd.t35 16.8893
R9509 gnd.n4384 gnd.t319 16.8893
R9510 gnd.n4850 gnd.t188 16.8893
R9511 gnd.n5064 gnd.t190 16.8893
R9512 gnd.n167 gnd.t19 16.8893
R9513 gnd.n5427 gnd.n5424 16.6793
R9514 gnd.n7014 gnd.n7011 16.6793
R9515 gnd.n3886 gnd.n3805 16.6793
R9516 gnd.n1120 gnd.n1117 16.6793
R9517 gnd.t81 gnd.n1805 16.5706
R9518 gnd.n2832 gnd.t115 16.2519
R9519 gnd.n2532 gnd.t132 16.2519
R9520 gnd.n4437 gnd.n4436 16.0975
R9521 gnd.n1792 gnd.n1791 16.0975
R9522 gnd.n5684 gnd.n5683 16.0975
R9523 gnd.n4890 gnd.n4889 16.0975
R9524 gnd.n4523 gnd.n4522 15.9333
R9525 gnd.n4682 gnd.t135 15.9333
R9526 gnd.n4702 gnd.n1894 15.9333
R9527 gnd.n4702 gnd.n1895 15.9333
R9528 gnd.n4732 gnd.t128 15.9333
R9529 gnd.n3519 gnd.n3517 15.6674
R9530 gnd.n3487 gnd.n3485 15.6674
R9531 gnd.n3455 gnd.n3453 15.6674
R9532 gnd.n3424 gnd.n3422 15.6674
R9533 gnd.n3392 gnd.n3390 15.6674
R9534 gnd.n3360 gnd.n3358 15.6674
R9535 gnd.n3328 gnd.n3326 15.6674
R9536 gnd.n3297 gnd.n3295 15.6674
R9537 gnd.n2823 gnd.t115 15.6146
R9538 gnd.t27 gnd.n2286 15.6146
R9539 gnd.t111 gnd.n2287 15.6146
R9540 gnd.n5384 gnd.n5379 15.3217
R9541 gnd.n6969 gnd.n6964 15.3217
R9542 gnd.n3840 gnd.n3837 15.3217
R9543 gnd.n1075 gnd.n1070 15.3217
R9544 gnd.n4581 gnd.t147 15.296
R9545 gnd.n1876 gnd.t130 15.296
R9546 gnd.n4874 gnd.n4873 15.0827
R9547 gnd.n1187 gnd.n1182 15.0481
R9548 gnd.n4884 gnd.n4883 15.0481
R9549 gnd.n3191 gnd.t186 14.9773
R9550 gnd.n3979 gnd.t35 14.9773
R9551 gnd.n5891 gnd.t39 14.9773
R9552 gnd.n2020 gnd.t319 14.9773
R9553 gnd.n5073 gnd.t190 14.9773
R9554 gnd.n5368 gnd.t23 14.9773
R9555 gnd.n7153 gnd.t19 14.9773
R9556 gnd.n5677 gnd.t87 14.6587
R9557 gnd.n4559 gnd.n1968 14.6587
R9558 gnd.n4512 gnd.t108 14.6587
R9559 gnd.n1825 gnd.n1824 14.6587
R9560 gnd.n1805 gnd.n1797 14.6587
R9561 gnd.n4961 gnd.t99 14.6587
R9562 gnd.n3269 gnd.t155 14.34
R9563 gnd.t316 gnd.t63 14.34
R9564 gnd.n2979 gnd.t169 13.7027
R9565 gnd.n2689 gnd.n2688 13.5763
R9566 gnd.n3633 gnd.n2243 13.5763
R9567 gnd.n2897 gnd.n2635 13.384
R9568 gnd.n4568 gnd.n4567 13.384
R9569 gnd.n4682 gnd.n1910 13.384
R9570 gnd.t124 gnd.n1899 13.384
R9571 gnd.n4715 gnd.t129 13.384
R9572 gnd.n4732 gnd.n4731 13.384
R9573 gnd.n4832 gnd.n1829 13.384
R9574 gnd.n1198 gnd.n1179 13.1884
R9575 gnd.n1193 gnd.n1192 13.1884
R9576 gnd.n1192 gnd.n1191 13.1884
R9577 gnd.n4877 gnd.n4872 13.1884
R9578 gnd.n4878 gnd.n4877 13.1884
R9579 gnd.n1194 gnd.n1181 13.146
R9580 gnd.n1190 gnd.n1181 13.146
R9581 gnd.n4876 gnd.n4875 13.146
R9582 gnd.n4876 gnd.n4871 13.146
R9583 gnd.n3520 gnd.n3516 12.8005
R9584 gnd.n3488 gnd.n3484 12.8005
R9585 gnd.n3456 gnd.n3452 12.8005
R9586 gnd.n3425 gnd.n3421 12.8005
R9587 gnd.n3393 gnd.n3389 12.8005
R9588 gnd.n3361 gnd.n3357 12.8005
R9589 gnd.n3329 gnd.n3325 12.8005
R9590 gnd.n3298 gnd.n3294 12.8005
R9591 gnd.n5967 gnd.n5966 12.7467
R9592 gnd.n4072 gnd.n736 12.7467
R9593 gnd.n5959 gnd.n744 12.7467
R9594 gnd.n4090 gnd.n747 12.7467
R9595 gnd.n4098 gnd.n758 12.7467
R9596 gnd.n5946 gnd.n763 12.7467
R9597 gnd.n4118 gnd.n4117 12.7467
R9598 gnd.n5940 gnd.n772 12.7467
R9599 gnd.n5933 gnd.n780 12.7467
R9600 gnd.n4153 gnd.n783 12.7467
R9601 gnd.n4161 gnd.n792 12.7467
R9602 gnd.n5921 gnd.n800 12.7467
R9603 gnd.n4167 gnd.n2106 12.7467
R9604 gnd.n5915 gnd.n809 12.7467
R9605 gnd.n5909 gnd.n820 12.7467
R9606 gnd.n4199 gnd.n823 12.7467
R9607 gnd.n4182 gnd.n832 12.7467
R9608 gnd.n5897 gnd.n840 12.7467
R9609 gnd.n4188 gnd.n843 12.7467
R9610 gnd.n5891 gnd.n850 12.7467
R9611 gnd.n5878 gnd.n867 12.7467
R9612 gnd.n5885 gnd.n859 12.7467
R9613 gnd.n5376 gnd.n1486 12.7467
R9614 gnd.n5219 gnd.n5218 12.7467
R9615 gnd.n5368 gnd.n1495 12.7467
R9616 gnd.n5179 gnd.n1508 12.7467
R9617 gnd.n5362 gnd.n1511 12.7467
R9618 gnd.n5186 gnd.n1521 12.7467
R9619 gnd.n5192 gnd.n1531 12.7467
R9620 gnd.n5350 gnd.n1534 12.7467
R9621 gnd.n5344 gnd.n1544 12.7467
R9622 gnd.n5261 gnd.n5260 12.7467
R9623 gnd.n5338 gnd.n1554 12.7467
R9624 gnd.n5269 gnd.n1561 12.7467
R9625 gnd.n5276 gnd.n1568 12.7467
R9626 gnd.n5326 gnd.n1571 12.7467
R9627 gnd.n5320 gnd.n1581 12.7467
R9628 gnd.n5315 gnd.n5314 12.7467
R9629 gnd.n5297 gnd.n1604 12.7467
R9630 gnd.n5307 gnd.n1596 12.7467
R9631 gnd.n7203 gnd.n75 12.7467
R9632 gnd.n6784 gnd.n6783 12.7467
R9633 gnd.n6791 gnd.n90 12.7467
R9634 gnd.n7195 gnd.n93 12.7467
R9635 gnd.t240 gnd.n775 12.4281
R9636 gnd.n4328 gnd.t171 12.4281
R9637 gnd.n1686 gnd.t194 12.4281
R9638 gnd.t196 gnd.n1578 12.4281
R9639 gnd.n2688 gnd.n2683 12.4126
R9640 gnd.n3636 gnd.n3633 12.4126
R9641 gnd.n5745 gnd.n5682 12.1761
R9642 gnd.n4957 gnd.n4956 12.1761
R9643 gnd.n5802 gnd.n965 12.1094
R9644 gnd.n4523 gnd.t6 12.1094
R9645 gnd.n4602 gnd.n1940 12.1094
R9646 gnd.n4654 gnd.n1919 12.1094
R9647 gnd.n4769 gnd.n1859 12.1094
R9648 gnd.n4812 gnd.n1838 12.1094
R9649 gnd.n4856 gnd.t10 12.1094
R9650 gnd.n5497 gnd.n1416 12.1094
R9651 gnd.n3524 gnd.n3523 12.0247
R9652 gnd.n3492 gnd.n3491 12.0247
R9653 gnd.n3460 gnd.n3459 12.0247
R9654 gnd.n3429 gnd.n3428 12.0247
R9655 gnd.n3397 gnd.n3396 12.0247
R9656 gnd.n3365 gnd.n3364 12.0247
R9657 gnd.n3333 gnd.n3332 12.0247
R9658 gnd.n3302 gnd.n3301 12.0247
R9659 gnd.n3999 gnd.t229 11.7908
R9660 gnd.t253 gnd.n812 11.7908
R9661 gnd.n5903 gnd.t211 11.7908
R9662 gnd.n5356 gnd.t217 11.7908
R9663 gnd.t219 gnd.n1541 11.7908
R9664 gnd.n7165 gnd.t202 11.7908
R9665 gnd.n1960 gnd.t125 11.4721
R9666 gnd.n4750 gnd.t144 11.4721
R9667 gnd.n4857 gnd.t3 11.4721
R9668 gnd.n3527 gnd.n3514 11.249
R9669 gnd.n3495 gnd.n3482 11.249
R9670 gnd.n3463 gnd.n3450 11.249
R9671 gnd.n3432 gnd.n3419 11.249
R9672 gnd.n3400 gnd.n3387 11.249
R9673 gnd.n3368 gnd.n3355 11.249
R9674 gnd.n3336 gnd.n3323 11.249
R9675 gnd.n3305 gnd.n3292 11.249
R9676 gnd.n2967 gnd.t169 11.1535
R9677 gnd.n4063 gnd.n2134 11.1535
R9678 gnd.n4063 gnd.t251 11.1535
R9679 gnd.n5927 gnd.t200 11.1535
R9680 gnd.n5332 gnd.t205 11.1535
R9681 gnd.n7189 gnd.t209 11.1535
R9682 gnd.n7189 gnd.n104 11.1535
R9683 gnd.n4612 gnd.n1932 10.8348
R9684 gnd.n4779 gnd.n1852 10.8348
R9685 gnd.n5387 gnd.n5384 10.6672
R9686 gnd.n6972 gnd.n6969 10.6672
R9687 gnd.n3846 gnd.n3837 10.6672
R9688 gnd.n1078 gnd.n1075 10.6672
R9689 gnd.n5027 gnd.n5026 10.6151
R9690 gnd.n5026 gnd.n5023 10.6151
R9691 gnd.n5021 gnd.n5018 10.6151
R9692 gnd.n5018 gnd.n5017 10.6151
R9693 gnd.n5017 gnd.n5014 10.6151
R9694 gnd.n5014 gnd.n5013 10.6151
R9695 gnd.n5013 gnd.n5010 10.6151
R9696 gnd.n5010 gnd.n5009 10.6151
R9697 gnd.n5009 gnd.n5006 10.6151
R9698 gnd.n5006 gnd.n5005 10.6151
R9699 gnd.n5005 gnd.n5002 10.6151
R9700 gnd.n5002 gnd.n5001 10.6151
R9701 gnd.n5001 gnd.n4998 10.6151
R9702 gnd.n4998 gnd.n4997 10.6151
R9703 gnd.n4997 gnd.n4994 10.6151
R9704 gnd.n4994 gnd.n4993 10.6151
R9705 gnd.n4993 gnd.n4990 10.6151
R9706 gnd.n4990 gnd.n4989 10.6151
R9707 gnd.n4989 gnd.n4986 10.6151
R9708 gnd.n4986 gnd.n4985 10.6151
R9709 gnd.n4985 gnd.n4982 10.6151
R9710 gnd.n4982 gnd.n4981 10.6151
R9711 gnd.n4981 gnd.n4978 10.6151
R9712 gnd.n4978 gnd.n4977 10.6151
R9713 gnd.n4977 gnd.n4974 10.6151
R9714 gnd.n4974 gnd.n4973 10.6151
R9715 gnd.n4973 gnd.n4970 10.6151
R9716 gnd.n4970 gnd.n4969 10.6151
R9717 gnd.n4969 gnd.n4966 10.6151
R9718 gnd.n4966 gnd.n4965 10.6151
R9719 gnd.n4503 gnd.n4502 10.6151
R9720 gnd.n4505 gnd.n4503 10.6151
R9721 gnd.n4506 gnd.n4505 10.6151
R9722 gnd.n4508 gnd.n4506 10.6151
R9723 gnd.n4509 gnd.n4508 10.6151
R9724 gnd.n4519 gnd.n4509 10.6151
R9725 gnd.n4519 gnd.n4518 10.6151
R9726 gnd.n4518 gnd.n4517 10.6151
R9727 gnd.n4517 gnd.n4515 10.6151
R9728 gnd.n4515 gnd.n4514 10.6151
R9729 gnd.n4514 gnd.n4511 10.6151
R9730 gnd.n4511 gnd.n4510 10.6151
R9731 gnd.n4510 gnd.n1952 10.6151
R9732 gnd.n4577 gnd.n1952 10.6151
R9733 gnd.n4578 gnd.n4577 10.6151
R9734 gnd.n4579 gnd.n4578 10.6151
R9735 gnd.n4593 gnd.n4579 10.6151
R9736 gnd.n4593 gnd.n4592 10.6151
R9737 gnd.n4592 gnd.n4591 10.6151
R9738 gnd.n4591 gnd.n4587 10.6151
R9739 gnd.n4587 gnd.n4586 10.6151
R9740 gnd.n4586 gnd.n4584 10.6151
R9741 gnd.n4584 gnd.n4583 10.6151
R9742 gnd.n4583 gnd.n4580 10.6151
R9743 gnd.n4580 gnd.n1901 10.6151
R9744 gnd.n4690 gnd.n1901 10.6151
R9745 gnd.n4691 gnd.n4690 10.6151
R9746 gnd.n4693 gnd.n4691 10.6151
R9747 gnd.n4693 gnd.n4692 10.6151
R9748 gnd.n4692 gnd.n1891 10.6151
R9749 gnd.n4705 gnd.n1891 10.6151
R9750 gnd.n4706 gnd.n4705 10.6151
R9751 gnd.n4712 gnd.n4706 10.6151
R9752 gnd.n4712 gnd.n4711 10.6151
R9753 gnd.n4711 gnd.n4710 10.6151
R9754 gnd.n4710 gnd.n4708 10.6151
R9755 gnd.n4708 gnd.n4707 10.6151
R9756 gnd.n4707 gnd.n1868 10.6151
R9757 gnd.n4741 gnd.n1868 10.6151
R9758 gnd.n4742 gnd.n4741 10.6151
R9759 gnd.n4747 gnd.n4742 10.6151
R9760 gnd.n4748 gnd.n4747 10.6151
R9761 gnd.n4758 gnd.n4748 10.6151
R9762 gnd.n4758 gnd.n4757 10.6151
R9763 gnd.n4757 gnd.n4756 10.6151
R9764 gnd.n4756 gnd.n4755 10.6151
R9765 gnd.n4755 gnd.n4753 10.6151
R9766 gnd.n4753 gnd.n4752 10.6151
R9767 gnd.n4752 gnd.n4749 10.6151
R9768 gnd.n4749 gnd.n1821 10.6151
R9769 gnd.n4840 gnd.n1821 10.6151
R9770 gnd.n4841 gnd.n4840 10.6151
R9771 gnd.n4848 gnd.n4841 10.6151
R9772 gnd.n4848 gnd.n4847 10.6151
R9773 gnd.n4847 gnd.n4846 10.6151
R9774 gnd.n4846 gnd.n4845 10.6151
R9775 gnd.n4845 gnd.n4843 10.6151
R9776 gnd.n4843 gnd.n4842 10.6151
R9777 gnd.n4842 gnd.n1795 10.6151
R9778 gnd.n1795 gnd.n1793 10.6151
R9779 gnd.n4438 gnd.n1139 10.6151
R9780 gnd.n4441 gnd.n4438 10.6151
R9781 gnd.n4446 gnd.n4443 10.6151
R9782 gnd.n4447 gnd.n4446 10.6151
R9783 gnd.n4450 gnd.n4447 10.6151
R9784 gnd.n4451 gnd.n4450 10.6151
R9785 gnd.n4454 gnd.n4451 10.6151
R9786 gnd.n4455 gnd.n4454 10.6151
R9787 gnd.n4458 gnd.n4455 10.6151
R9788 gnd.n4459 gnd.n4458 10.6151
R9789 gnd.n4462 gnd.n4459 10.6151
R9790 gnd.n4463 gnd.n4462 10.6151
R9791 gnd.n4466 gnd.n4463 10.6151
R9792 gnd.n4467 gnd.n4466 10.6151
R9793 gnd.n4470 gnd.n4467 10.6151
R9794 gnd.n4471 gnd.n4470 10.6151
R9795 gnd.n4474 gnd.n4471 10.6151
R9796 gnd.n4475 gnd.n4474 10.6151
R9797 gnd.n4478 gnd.n4475 10.6151
R9798 gnd.n4479 gnd.n4478 10.6151
R9799 gnd.n4482 gnd.n4479 10.6151
R9800 gnd.n4483 gnd.n4482 10.6151
R9801 gnd.n4486 gnd.n4483 10.6151
R9802 gnd.n4487 gnd.n4486 10.6151
R9803 gnd.n4490 gnd.n4487 10.6151
R9804 gnd.n4491 gnd.n4490 10.6151
R9805 gnd.n4494 gnd.n4491 10.6151
R9806 gnd.n4495 gnd.n4494 10.6151
R9807 gnd.n4498 gnd.n4495 10.6151
R9808 gnd.n4499 gnd.n4498 10.6151
R9809 gnd.n5745 gnd.n5744 10.6151
R9810 gnd.n5744 gnd.n5743 10.6151
R9811 gnd.n5743 gnd.n5742 10.6151
R9812 gnd.n5742 gnd.n5740 10.6151
R9813 gnd.n5740 gnd.n5737 10.6151
R9814 gnd.n5737 gnd.n5736 10.6151
R9815 gnd.n5736 gnd.n5733 10.6151
R9816 gnd.n5733 gnd.n5732 10.6151
R9817 gnd.n5732 gnd.n5729 10.6151
R9818 gnd.n5729 gnd.n5728 10.6151
R9819 gnd.n5728 gnd.n5725 10.6151
R9820 gnd.n5725 gnd.n5724 10.6151
R9821 gnd.n5724 gnd.n5721 10.6151
R9822 gnd.n5721 gnd.n5720 10.6151
R9823 gnd.n5720 gnd.n5717 10.6151
R9824 gnd.n5717 gnd.n5716 10.6151
R9825 gnd.n5716 gnd.n5713 10.6151
R9826 gnd.n5713 gnd.n5712 10.6151
R9827 gnd.n5712 gnd.n5709 10.6151
R9828 gnd.n5709 gnd.n5708 10.6151
R9829 gnd.n5708 gnd.n5705 10.6151
R9830 gnd.n5705 gnd.n5704 10.6151
R9831 gnd.n5704 gnd.n5701 10.6151
R9832 gnd.n5701 gnd.n5700 10.6151
R9833 gnd.n5700 gnd.n5697 10.6151
R9834 gnd.n5697 gnd.n5696 10.6151
R9835 gnd.n5696 gnd.n5693 10.6151
R9836 gnd.n5693 gnd.n5692 10.6151
R9837 gnd.n5689 gnd.n5688 10.6151
R9838 gnd.n5688 gnd.n1140 10.6151
R9839 gnd.n4956 gnd.n4954 10.6151
R9840 gnd.n4954 gnd.n4951 10.6151
R9841 gnd.n4951 gnd.n4950 10.6151
R9842 gnd.n4950 gnd.n4947 10.6151
R9843 gnd.n4947 gnd.n4946 10.6151
R9844 gnd.n4946 gnd.n4943 10.6151
R9845 gnd.n4943 gnd.n4942 10.6151
R9846 gnd.n4942 gnd.n4939 10.6151
R9847 gnd.n4939 gnd.n4938 10.6151
R9848 gnd.n4938 gnd.n4935 10.6151
R9849 gnd.n4935 gnd.n4934 10.6151
R9850 gnd.n4934 gnd.n4931 10.6151
R9851 gnd.n4931 gnd.n4930 10.6151
R9852 gnd.n4930 gnd.n4927 10.6151
R9853 gnd.n4927 gnd.n4926 10.6151
R9854 gnd.n4926 gnd.n4923 10.6151
R9855 gnd.n4923 gnd.n4922 10.6151
R9856 gnd.n4922 gnd.n4919 10.6151
R9857 gnd.n4919 gnd.n4918 10.6151
R9858 gnd.n4918 gnd.n4915 10.6151
R9859 gnd.n4915 gnd.n4914 10.6151
R9860 gnd.n4914 gnd.n4911 10.6151
R9861 gnd.n4911 gnd.n4910 10.6151
R9862 gnd.n4910 gnd.n4907 10.6151
R9863 gnd.n4907 gnd.n4906 10.6151
R9864 gnd.n4906 gnd.n4903 10.6151
R9865 gnd.n4903 gnd.n4902 10.6151
R9866 gnd.n4902 gnd.n4899 10.6151
R9867 gnd.n4897 gnd.n4894 10.6151
R9868 gnd.n4894 gnd.n4893 10.6151
R9869 gnd.n5681 gnd.n5680 10.6151
R9870 gnd.n5680 gnd.n1199 10.6151
R9871 gnd.n4527 gnd.n1199 10.6151
R9872 gnd.n4527 gnd.n4526 10.6151
R9873 gnd.n4526 gnd.n4525 10.6151
R9874 gnd.n4525 gnd.n1972 10.6151
R9875 gnd.n4554 gnd.n1972 10.6151
R9876 gnd.n4555 gnd.n4554 10.6151
R9877 gnd.n4556 gnd.n4555 10.6151
R9878 gnd.n4556 gnd.n1955 10.6151
R9879 gnd.n4570 gnd.n1955 10.6151
R9880 gnd.n4571 gnd.n4570 10.6151
R9881 gnd.n4572 gnd.n4571 10.6151
R9882 gnd.n4572 gnd.n1946 10.6151
R9883 gnd.n4599 gnd.n1946 10.6151
R9884 gnd.n4599 gnd.n4598 10.6151
R9885 gnd.n4598 gnd.n4597 10.6151
R9886 gnd.n4597 gnd.n1947 10.6151
R9887 gnd.n1947 gnd.n1923 10.6151
R9888 gnd.n4657 gnd.n1923 10.6151
R9889 gnd.n4658 gnd.n4657 10.6151
R9890 gnd.n4659 gnd.n4658 10.6151
R9891 gnd.n4659 gnd.n1907 10.6151
R9892 gnd.n4684 gnd.n1907 10.6151
R9893 gnd.n4685 gnd.n4684 10.6151
R9894 gnd.n4686 gnd.n4685 10.6151
R9895 gnd.n4686 gnd.n1897 10.6151
R9896 gnd.n4698 gnd.n1897 10.6151
R9897 gnd.n4699 gnd.n4698 10.6151
R9898 gnd.n4700 gnd.n4699 10.6151
R9899 gnd.n4700 gnd.n1886 10.6151
R9900 gnd.n4718 gnd.n1886 10.6151
R9901 gnd.n4719 gnd.n4718 10.6151
R9902 gnd.n4720 gnd.n4719 10.6151
R9903 gnd.n4720 gnd.n1872 10.6151
R9904 gnd.n4734 gnd.n1872 10.6151
R9905 gnd.n4735 gnd.n4734 10.6151
R9906 gnd.n4736 gnd.n4735 10.6151
R9907 gnd.n4736 gnd.n1864 10.6151
R9908 gnd.n4766 gnd.n1864 10.6151
R9909 gnd.n4766 gnd.n4765 10.6151
R9910 gnd.n4765 gnd.n4764 10.6151
R9911 gnd.n4764 gnd.n1865 10.6151
R9912 gnd.n1865 gnd.n1842 10.6151
R9913 gnd.n4815 gnd.n1842 10.6151
R9914 gnd.n4816 gnd.n4815 10.6151
R9915 gnd.n4817 gnd.n4816 10.6151
R9916 gnd.n4817 gnd.n1827 10.6151
R9917 gnd.n4834 gnd.n1827 10.6151
R9918 gnd.n4835 gnd.n4834 10.6151
R9919 gnd.n4836 gnd.n4835 10.6151
R9920 gnd.n4836 gnd.n1815 10.6151
R9921 gnd.n4852 gnd.n1815 10.6151
R9922 gnd.n4853 gnd.n4852 10.6151
R9923 gnd.n4854 gnd.n4853 10.6151
R9924 gnd.n4854 gnd.n1800 10.6151
R9925 gnd.n4868 gnd.n1800 10.6151
R9926 gnd.n4869 gnd.n4868 10.6151
R9927 gnd.n4959 gnd.n4869 10.6151
R9928 gnd.n4959 gnd.n4958 10.6151
R9929 gnd.n2886 gnd.t133 10.5161
R9930 gnd.n2331 gnd.t166 10.5161
R9931 gnd.n3252 gnd.t155 10.5161
R9932 gnd.n5953 gnd.t207 10.5161
R9933 gnd.n5946 gnd.t213 10.5161
R9934 gnd.n5297 gnd.t243 10.5161
R9935 gnd.n5306 gnd.t245 10.5161
R9936 gnd.n3528 gnd.n3512 10.4732
R9937 gnd.n3496 gnd.n3480 10.4732
R9938 gnd.n3464 gnd.n3448 10.4732
R9939 gnd.n3433 gnd.n3417 10.4732
R9940 gnd.n3401 gnd.n3385 10.4732
R9941 gnd.n3369 gnd.n3353 10.4732
R9942 gnd.n3337 gnd.n3321 10.4732
R9943 gnd.n3306 gnd.n3290 10.4732
R9944 gnd.n4574 gnd.t125 10.1975
R9945 gnd.n4819 gnd.t144 10.1975
R9946 gnd.t186 gnd.n2348 9.87883
R9947 gnd.n4054 gnd.t236 9.87883
R9948 gnd.n5921 gnd.t264 9.87883
R9949 gnd.n5338 gnd.t227 9.87883
R9950 gnd.n7183 gnd.t215 9.87883
R9951 gnd.n3532 gnd.n3531 9.69747
R9952 gnd.n3500 gnd.n3499 9.69747
R9953 gnd.n3468 gnd.n3467 9.69747
R9954 gnd.n3437 gnd.n3436 9.69747
R9955 gnd.n3405 gnd.n3404 9.69747
R9956 gnd.n3373 gnd.n3372 9.69747
R9957 gnd.n3341 gnd.n3340 9.69747
R9958 gnd.n3310 gnd.n3309 9.69747
R9959 gnd.n4655 gnd.n4654 9.56018
R9960 gnd.n4769 gnd.n4768 9.56018
R9961 gnd.t60 gnd.n1818 9.56018
R9962 gnd.n3538 gnd.n3537 9.45567
R9963 gnd.n3506 gnd.n3505 9.45567
R9964 gnd.n3474 gnd.n3473 9.45567
R9965 gnd.n3443 gnd.n3442 9.45567
R9966 gnd.n3411 gnd.n3410 9.45567
R9967 gnd.n3379 gnd.n3378 9.45567
R9968 gnd.n3347 gnd.n3346 9.45567
R9969 gnd.n3316 gnd.n3315 9.45567
R9970 gnd.n5424 gnd.n5423 9.30959
R9971 gnd.n7011 gnd.n6943 9.30959
R9972 gnd.n3880 gnd.n3805 9.30959
R9973 gnd.n1117 gnd.n1049 9.30959
R9974 gnd.n3537 gnd.n3536 9.3005
R9975 gnd.n3510 gnd.n3509 9.3005
R9976 gnd.n3531 gnd.n3530 9.3005
R9977 gnd.n3529 gnd.n3528 9.3005
R9978 gnd.n3514 gnd.n3513 9.3005
R9979 gnd.n3523 gnd.n3522 9.3005
R9980 gnd.n3521 gnd.n3520 9.3005
R9981 gnd.n3505 gnd.n3504 9.3005
R9982 gnd.n3478 gnd.n3477 9.3005
R9983 gnd.n3499 gnd.n3498 9.3005
R9984 gnd.n3497 gnd.n3496 9.3005
R9985 gnd.n3482 gnd.n3481 9.3005
R9986 gnd.n3491 gnd.n3490 9.3005
R9987 gnd.n3489 gnd.n3488 9.3005
R9988 gnd.n3473 gnd.n3472 9.3005
R9989 gnd.n3446 gnd.n3445 9.3005
R9990 gnd.n3467 gnd.n3466 9.3005
R9991 gnd.n3465 gnd.n3464 9.3005
R9992 gnd.n3450 gnd.n3449 9.3005
R9993 gnd.n3459 gnd.n3458 9.3005
R9994 gnd.n3457 gnd.n3456 9.3005
R9995 gnd.n3442 gnd.n3441 9.3005
R9996 gnd.n3415 gnd.n3414 9.3005
R9997 gnd.n3436 gnd.n3435 9.3005
R9998 gnd.n3434 gnd.n3433 9.3005
R9999 gnd.n3419 gnd.n3418 9.3005
R10000 gnd.n3428 gnd.n3427 9.3005
R10001 gnd.n3426 gnd.n3425 9.3005
R10002 gnd.n3410 gnd.n3409 9.3005
R10003 gnd.n3383 gnd.n3382 9.3005
R10004 gnd.n3404 gnd.n3403 9.3005
R10005 gnd.n3402 gnd.n3401 9.3005
R10006 gnd.n3387 gnd.n3386 9.3005
R10007 gnd.n3396 gnd.n3395 9.3005
R10008 gnd.n3394 gnd.n3393 9.3005
R10009 gnd.n3378 gnd.n3377 9.3005
R10010 gnd.n3351 gnd.n3350 9.3005
R10011 gnd.n3372 gnd.n3371 9.3005
R10012 gnd.n3370 gnd.n3369 9.3005
R10013 gnd.n3355 gnd.n3354 9.3005
R10014 gnd.n3364 gnd.n3363 9.3005
R10015 gnd.n3362 gnd.n3361 9.3005
R10016 gnd.n3346 gnd.n3345 9.3005
R10017 gnd.n3319 gnd.n3318 9.3005
R10018 gnd.n3340 gnd.n3339 9.3005
R10019 gnd.n3338 gnd.n3337 9.3005
R10020 gnd.n3323 gnd.n3322 9.3005
R10021 gnd.n3332 gnd.n3331 9.3005
R10022 gnd.n3330 gnd.n3329 9.3005
R10023 gnd.n3315 gnd.n3314 9.3005
R10024 gnd.n3288 gnd.n3287 9.3005
R10025 gnd.n3309 gnd.n3308 9.3005
R10026 gnd.n3307 gnd.n3306 9.3005
R10027 gnd.n3292 gnd.n3291 9.3005
R10028 gnd.n3301 gnd.n3300 9.3005
R10029 gnd.n3299 gnd.n3298 9.3005
R10030 gnd.n3663 gnd.n3662 9.3005
R10031 gnd.n3661 gnd.n2231 9.3005
R10032 gnd.n3660 gnd.n3659 9.3005
R10033 gnd.n3656 gnd.n2232 9.3005
R10034 gnd.n3653 gnd.n2233 9.3005
R10035 gnd.n3652 gnd.n2234 9.3005
R10036 gnd.n3649 gnd.n2235 9.3005
R10037 gnd.n3648 gnd.n2236 9.3005
R10038 gnd.n3645 gnd.n2237 9.3005
R10039 gnd.n3644 gnd.n2238 9.3005
R10040 gnd.n3641 gnd.n2239 9.3005
R10041 gnd.n3640 gnd.n2240 9.3005
R10042 gnd.n3637 gnd.n2241 9.3005
R10043 gnd.n3636 gnd.n2242 9.3005
R10044 gnd.n3633 gnd.n3632 9.3005
R10045 gnd.n3631 gnd.n2243 9.3005
R10046 gnd.n3664 gnd.n2230 9.3005
R10047 gnd.n2905 gnd.n2904 9.3005
R10048 gnd.n2609 gnd.n2608 9.3005
R10049 gnd.n2932 gnd.n2931 9.3005
R10050 gnd.n2933 gnd.n2607 9.3005
R10051 gnd.n2937 gnd.n2934 9.3005
R10052 gnd.n2936 gnd.n2935 9.3005
R10053 gnd.n2581 gnd.n2580 9.3005
R10054 gnd.n2962 gnd.n2961 9.3005
R10055 gnd.n2963 gnd.n2579 9.3005
R10056 gnd.n2965 gnd.n2964 9.3005
R10057 gnd.n2559 gnd.n2558 9.3005
R10058 gnd.n2993 gnd.n2992 9.3005
R10059 gnd.n2994 gnd.n2557 9.3005
R10060 gnd.n3002 gnd.n2995 9.3005
R10061 gnd.n3001 gnd.n2996 9.3005
R10062 gnd.n3000 gnd.n2998 9.3005
R10063 gnd.n2997 gnd.n2506 9.3005
R10064 gnd.n3050 gnd.n2507 9.3005
R10065 gnd.n3049 gnd.n2508 9.3005
R10066 gnd.n3048 gnd.n2509 9.3005
R10067 gnd.n2528 gnd.n2510 9.3005
R10068 gnd.n2530 gnd.n2529 9.3005
R10069 gnd.n2428 gnd.n2427 9.3005
R10070 gnd.n3088 gnd.n3087 9.3005
R10071 gnd.n3089 gnd.n2426 9.3005
R10072 gnd.n3093 gnd.n3090 9.3005
R10073 gnd.n3092 gnd.n3091 9.3005
R10074 gnd.n2401 gnd.n2400 9.3005
R10075 gnd.n3128 gnd.n3127 9.3005
R10076 gnd.n3129 gnd.n2399 9.3005
R10077 gnd.n3133 gnd.n3130 9.3005
R10078 gnd.n3132 gnd.n3131 9.3005
R10079 gnd.n2374 gnd.n2373 9.3005
R10080 gnd.n3173 gnd.n3172 9.3005
R10081 gnd.n3174 gnd.n2372 9.3005
R10082 gnd.n3178 gnd.n3175 9.3005
R10083 gnd.n3177 gnd.n3176 9.3005
R10084 gnd.n2346 gnd.n2345 9.3005
R10085 gnd.n3213 gnd.n3212 9.3005
R10086 gnd.n3214 gnd.n2344 9.3005
R10087 gnd.n3218 gnd.n3215 9.3005
R10088 gnd.n3217 gnd.n3216 9.3005
R10089 gnd.n2319 gnd.n2318 9.3005
R10090 gnd.n3262 gnd.n3261 9.3005
R10091 gnd.n3263 gnd.n2317 9.3005
R10092 gnd.n3267 gnd.n3264 9.3005
R10093 gnd.n3266 gnd.n3265 9.3005
R10094 gnd.n2292 gnd.n2291 9.3005
R10095 gnd.n3556 gnd.n3555 9.3005
R10096 gnd.n3557 gnd.n2290 9.3005
R10097 gnd.n3563 gnd.n3558 9.3005
R10098 gnd.n3562 gnd.n3559 9.3005
R10099 gnd.n3561 gnd.n3560 9.3005
R10100 gnd.n2906 gnd.n2903 9.3005
R10101 gnd.n2688 gnd.n2647 9.3005
R10102 gnd.n2683 gnd.n2682 9.3005
R10103 gnd.n2681 gnd.n2648 9.3005
R10104 gnd.n2680 gnd.n2679 9.3005
R10105 gnd.n2676 gnd.n2649 9.3005
R10106 gnd.n2673 gnd.n2672 9.3005
R10107 gnd.n2671 gnd.n2650 9.3005
R10108 gnd.n2670 gnd.n2669 9.3005
R10109 gnd.n2666 gnd.n2651 9.3005
R10110 gnd.n2663 gnd.n2662 9.3005
R10111 gnd.n2661 gnd.n2652 9.3005
R10112 gnd.n2660 gnd.n2659 9.3005
R10113 gnd.n2656 gnd.n2654 9.3005
R10114 gnd.n2653 gnd.n2633 9.3005
R10115 gnd.n2900 gnd.n2632 9.3005
R10116 gnd.n2902 gnd.n2901 9.3005
R10117 gnd.n2690 gnd.n2689 9.3005
R10118 gnd.n2913 gnd.n2619 9.3005
R10119 gnd.n2920 gnd.n2620 9.3005
R10120 gnd.n2922 gnd.n2921 9.3005
R10121 gnd.n2923 gnd.n2600 9.3005
R10122 gnd.n2942 gnd.n2941 9.3005
R10123 gnd.n2944 gnd.n2592 9.3005
R10124 gnd.n2951 gnd.n2594 9.3005
R10125 gnd.n2952 gnd.n2589 9.3005
R10126 gnd.n2954 gnd.n2953 9.3005
R10127 gnd.n2590 gnd.n2575 9.3005
R10128 gnd.n2970 gnd.n2573 9.3005
R10129 gnd.n2974 gnd.n2973 9.3005
R10130 gnd.n2972 gnd.n2549 9.3005
R10131 gnd.n3009 gnd.n2548 9.3005
R10132 gnd.n3012 gnd.n3011 9.3005
R10133 gnd.n2545 gnd.n2544 9.3005
R10134 gnd.n3018 gnd.n2546 9.3005
R10135 gnd.n3020 gnd.n3019 9.3005
R10136 gnd.n3022 gnd.n2543 9.3005
R10137 gnd.n3025 gnd.n3024 9.3005
R10138 gnd.n3028 gnd.n3026 9.3005
R10139 gnd.n3030 gnd.n3029 9.3005
R10140 gnd.n3036 gnd.n3031 9.3005
R10141 gnd.n3035 gnd.n3034 9.3005
R10142 gnd.n2419 gnd.n2418 9.3005
R10143 gnd.n3102 gnd.n3101 9.3005
R10144 gnd.n3103 gnd.n2412 9.3005
R10145 gnd.n3111 gnd.n2411 9.3005
R10146 gnd.n3114 gnd.n3113 9.3005
R10147 gnd.n3116 gnd.n3115 9.3005
R10148 gnd.n3119 gnd.n2394 9.3005
R10149 gnd.n3117 gnd.n2392 9.3005
R10150 gnd.n3139 gnd.n2390 9.3005
R10151 gnd.n3141 gnd.n3140 9.3005
R10152 gnd.n2364 gnd.n2363 9.3005
R10153 gnd.n3187 gnd.n3186 9.3005
R10154 gnd.n3188 gnd.n2357 9.3005
R10155 gnd.n3196 gnd.n2356 9.3005
R10156 gnd.n3199 gnd.n3198 9.3005
R10157 gnd.n3201 gnd.n3200 9.3005
R10158 gnd.n3204 gnd.n2339 9.3005
R10159 gnd.n3202 gnd.n2337 9.3005
R10160 gnd.n3224 gnd.n2335 9.3005
R10161 gnd.n3226 gnd.n3225 9.3005
R10162 gnd.n2310 gnd.n2309 9.3005
R10163 gnd.n3276 gnd.n3275 9.3005
R10164 gnd.n3277 gnd.n2303 9.3005
R10165 gnd.n3285 gnd.n2302 9.3005
R10166 gnd.n3544 gnd.n3543 9.3005
R10167 gnd.n3546 gnd.n3545 9.3005
R10168 gnd.n3547 gnd.n2283 9.3005
R10169 gnd.n3571 gnd.n3570 9.3005
R10170 gnd.n2284 gnd.n2246 9.3005
R10171 gnd.n2911 gnd.n2910 9.3005
R10172 gnd.n3627 gnd.n2247 9.3005
R10173 gnd.n3626 gnd.n2249 9.3005
R10174 gnd.n3623 gnd.n2250 9.3005
R10175 gnd.n3622 gnd.n2251 9.3005
R10176 gnd.n3619 gnd.n2252 9.3005
R10177 gnd.n3618 gnd.n2253 9.3005
R10178 gnd.n3615 gnd.n2254 9.3005
R10179 gnd.n3614 gnd.n2255 9.3005
R10180 gnd.n3611 gnd.n2256 9.3005
R10181 gnd.n3610 gnd.n2257 9.3005
R10182 gnd.n3607 gnd.n2258 9.3005
R10183 gnd.n3606 gnd.n2259 9.3005
R10184 gnd.n3603 gnd.n2260 9.3005
R10185 gnd.n3602 gnd.n2261 9.3005
R10186 gnd.n3599 gnd.n2262 9.3005
R10187 gnd.n3598 gnd.n2263 9.3005
R10188 gnd.n3595 gnd.n2264 9.3005
R10189 gnd.n3594 gnd.n2265 9.3005
R10190 gnd.n3591 gnd.n2266 9.3005
R10191 gnd.n3590 gnd.n2267 9.3005
R10192 gnd.n3587 gnd.n2268 9.3005
R10193 gnd.n3586 gnd.n2269 9.3005
R10194 gnd.n3583 gnd.n2273 9.3005
R10195 gnd.n3582 gnd.n2274 9.3005
R10196 gnd.n3579 gnd.n2275 9.3005
R10197 gnd.n3578 gnd.n2276 9.3005
R10198 gnd.n3629 gnd.n3628 9.3005
R10199 gnd.n3080 gnd.n3064 9.3005
R10200 gnd.n3079 gnd.n3065 9.3005
R10201 gnd.n3078 gnd.n3066 9.3005
R10202 gnd.n3076 gnd.n3067 9.3005
R10203 gnd.n3075 gnd.n3068 9.3005
R10204 gnd.n3073 gnd.n3069 9.3005
R10205 gnd.n3072 gnd.n3070 9.3005
R10206 gnd.n2382 gnd.n2381 9.3005
R10207 gnd.n3149 gnd.n3148 9.3005
R10208 gnd.n3150 gnd.n2380 9.3005
R10209 gnd.n3167 gnd.n3151 9.3005
R10210 gnd.n3166 gnd.n3152 9.3005
R10211 gnd.n3165 gnd.n3153 9.3005
R10212 gnd.n3163 gnd.n3154 9.3005
R10213 gnd.n3162 gnd.n3155 9.3005
R10214 gnd.n3160 gnd.n3156 9.3005
R10215 gnd.n3159 gnd.n3157 9.3005
R10216 gnd.n2326 gnd.n2325 9.3005
R10217 gnd.n3234 gnd.n3233 9.3005
R10218 gnd.n3235 gnd.n2324 9.3005
R10219 gnd.n3256 gnd.n3236 9.3005
R10220 gnd.n3255 gnd.n3237 9.3005
R10221 gnd.n3254 gnd.n3238 9.3005
R10222 gnd.n3251 gnd.n3239 9.3005
R10223 gnd.n3250 gnd.n3240 9.3005
R10224 gnd.n3248 gnd.n3241 9.3005
R10225 gnd.n3247 gnd.n3242 9.3005
R10226 gnd.n3245 gnd.n3244 9.3005
R10227 gnd.n3243 gnd.n2278 9.3005
R10228 gnd.n2821 gnd.n2820 9.3005
R10229 gnd.n2711 gnd.n2710 9.3005
R10230 gnd.n2835 gnd.n2834 9.3005
R10231 gnd.n2836 gnd.n2709 9.3005
R10232 gnd.n2838 gnd.n2837 9.3005
R10233 gnd.n2699 gnd.n2698 9.3005
R10234 gnd.n2851 gnd.n2850 9.3005
R10235 gnd.n2852 gnd.n2697 9.3005
R10236 gnd.n2884 gnd.n2853 9.3005
R10237 gnd.n2883 gnd.n2854 9.3005
R10238 gnd.n2882 gnd.n2855 9.3005
R10239 gnd.n2881 gnd.n2856 9.3005
R10240 gnd.n2878 gnd.n2857 9.3005
R10241 gnd.n2877 gnd.n2858 9.3005
R10242 gnd.n2876 gnd.n2859 9.3005
R10243 gnd.n2874 gnd.n2860 9.3005
R10244 gnd.n2873 gnd.n2861 9.3005
R10245 gnd.n2870 gnd.n2862 9.3005
R10246 gnd.n2869 gnd.n2863 9.3005
R10247 gnd.n2868 gnd.n2864 9.3005
R10248 gnd.n2866 gnd.n2865 9.3005
R10249 gnd.n2565 gnd.n2564 9.3005
R10250 gnd.n2982 gnd.n2981 9.3005
R10251 gnd.n2983 gnd.n2563 9.3005
R10252 gnd.n2987 gnd.n2984 9.3005
R10253 gnd.n2986 gnd.n2985 9.3005
R10254 gnd.n2487 gnd.n2486 9.3005
R10255 gnd.n3062 gnd.n3061 9.3005
R10256 gnd.n2819 gnd.n2720 9.3005
R10257 gnd.n2722 gnd.n2721 9.3005
R10258 gnd.n2766 gnd.n2764 9.3005
R10259 gnd.n2767 gnd.n2763 9.3005
R10260 gnd.n2770 gnd.n2759 9.3005
R10261 gnd.n2771 gnd.n2758 9.3005
R10262 gnd.n2774 gnd.n2757 9.3005
R10263 gnd.n2775 gnd.n2756 9.3005
R10264 gnd.n2778 gnd.n2755 9.3005
R10265 gnd.n2779 gnd.n2754 9.3005
R10266 gnd.n2782 gnd.n2753 9.3005
R10267 gnd.n2783 gnd.n2752 9.3005
R10268 gnd.n2786 gnd.n2751 9.3005
R10269 gnd.n2787 gnd.n2750 9.3005
R10270 gnd.n2790 gnd.n2749 9.3005
R10271 gnd.n2791 gnd.n2748 9.3005
R10272 gnd.n2794 gnd.n2747 9.3005
R10273 gnd.n2795 gnd.n2746 9.3005
R10274 gnd.n2798 gnd.n2745 9.3005
R10275 gnd.n2799 gnd.n2744 9.3005
R10276 gnd.n2802 gnd.n2743 9.3005
R10277 gnd.n2803 gnd.n2742 9.3005
R10278 gnd.n2806 gnd.n2741 9.3005
R10279 gnd.n2808 gnd.n2740 9.3005
R10280 gnd.n2809 gnd.n2739 9.3005
R10281 gnd.n2810 gnd.n2738 9.3005
R10282 gnd.n2811 gnd.n2737 9.3005
R10283 gnd.n2818 gnd.n2817 9.3005
R10284 gnd.n2827 gnd.n2826 9.3005
R10285 gnd.n2828 gnd.n2714 9.3005
R10286 gnd.n2830 gnd.n2829 9.3005
R10287 gnd.n2705 gnd.n2704 9.3005
R10288 gnd.n2843 gnd.n2842 9.3005
R10289 gnd.n2844 gnd.n2703 9.3005
R10290 gnd.n2846 gnd.n2845 9.3005
R10291 gnd.n2692 gnd.n2691 9.3005
R10292 gnd.n2889 gnd.n2888 9.3005
R10293 gnd.n2890 gnd.n2646 9.3005
R10294 gnd.n2894 gnd.n2892 9.3005
R10295 gnd.n2893 gnd.n2625 9.3005
R10296 gnd.n2912 gnd.n2624 9.3005
R10297 gnd.n2915 gnd.n2914 9.3005
R10298 gnd.n2618 gnd.n2617 9.3005
R10299 gnd.n2926 gnd.n2924 9.3005
R10300 gnd.n2925 gnd.n2599 9.3005
R10301 gnd.n2943 gnd.n2598 9.3005
R10302 gnd.n2946 gnd.n2945 9.3005
R10303 gnd.n2593 gnd.n2588 9.3005
R10304 gnd.n2956 gnd.n2955 9.3005
R10305 gnd.n2591 gnd.n2571 9.3005
R10306 gnd.n2977 gnd.n2572 9.3005
R10307 gnd.n2976 gnd.n2975 9.3005
R10308 gnd.n2574 gnd.n2550 9.3005
R10309 gnd.n3008 gnd.n3007 9.3005
R10310 gnd.n3010 gnd.n2495 9.3005
R10311 gnd.n3057 gnd.n2496 9.3005
R10312 gnd.n3056 gnd.n2497 9.3005
R10313 gnd.n3055 gnd.n2498 9.3005
R10314 gnd.n3021 gnd.n2499 9.3005
R10315 gnd.n3023 gnd.n2517 9.3005
R10316 gnd.n3043 gnd.n2518 9.3005
R10317 gnd.n3042 gnd.n2519 9.3005
R10318 gnd.n3041 gnd.n2520 9.3005
R10319 gnd.n3032 gnd.n2521 9.3005
R10320 gnd.n3033 gnd.n2420 9.3005
R10321 gnd.n3099 gnd.n3098 9.3005
R10322 gnd.n3100 gnd.n2413 9.3005
R10323 gnd.n3110 gnd.n3109 9.3005
R10324 gnd.n3112 gnd.n2409 9.3005
R10325 gnd.n3122 gnd.n2410 9.3005
R10326 gnd.n3121 gnd.n3120 9.3005
R10327 gnd.n3118 gnd.n2388 9.3005
R10328 gnd.n3144 gnd.n2389 9.3005
R10329 gnd.n3143 gnd.n3142 9.3005
R10330 gnd.n2391 gnd.n2365 9.3005
R10331 gnd.n3184 gnd.n3183 9.3005
R10332 gnd.n3185 gnd.n2358 9.3005
R10333 gnd.n3195 gnd.n3194 9.3005
R10334 gnd.n3197 gnd.n2354 9.3005
R10335 gnd.n3207 gnd.n2355 9.3005
R10336 gnd.n3206 gnd.n3205 9.3005
R10337 gnd.n3203 gnd.n2333 9.3005
R10338 gnd.n3229 gnd.n2334 9.3005
R10339 gnd.n3228 gnd.n3227 9.3005
R10340 gnd.n2336 gnd.n2311 9.3005
R10341 gnd.n3273 gnd.n3272 9.3005
R10342 gnd.n3274 gnd.n2304 9.3005
R10343 gnd.n3284 gnd.n3283 9.3005
R10344 gnd.n3542 gnd.n2300 9.3005
R10345 gnd.n3550 gnd.n2301 9.3005
R10346 gnd.n3549 gnd.n3548 9.3005
R10347 gnd.n2282 gnd.n2281 9.3005
R10348 gnd.n3573 gnd.n3572 9.3005
R10349 gnd.n2716 gnd.n2715 9.3005
R10350 gnd.n6143 gnd.n6142 9.3005
R10351 gnd.n559 gnd.n558 9.3005
R10352 gnd.n6150 gnd.n6149 9.3005
R10353 gnd.n6151 gnd.n557 9.3005
R10354 gnd.n6153 gnd.n6152 9.3005
R10355 gnd.n553 gnd.n552 9.3005
R10356 gnd.n6160 gnd.n6159 9.3005
R10357 gnd.n6161 gnd.n551 9.3005
R10358 gnd.n6163 gnd.n6162 9.3005
R10359 gnd.n547 gnd.n546 9.3005
R10360 gnd.n6170 gnd.n6169 9.3005
R10361 gnd.n6171 gnd.n545 9.3005
R10362 gnd.n6173 gnd.n6172 9.3005
R10363 gnd.n541 gnd.n540 9.3005
R10364 gnd.n6180 gnd.n6179 9.3005
R10365 gnd.n6181 gnd.n539 9.3005
R10366 gnd.n6183 gnd.n6182 9.3005
R10367 gnd.n535 gnd.n534 9.3005
R10368 gnd.n6190 gnd.n6189 9.3005
R10369 gnd.n6191 gnd.n533 9.3005
R10370 gnd.n6193 gnd.n6192 9.3005
R10371 gnd.n529 gnd.n528 9.3005
R10372 gnd.n6200 gnd.n6199 9.3005
R10373 gnd.n6201 gnd.n527 9.3005
R10374 gnd.n6203 gnd.n6202 9.3005
R10375 gnd.n523 gnd.n522 9.3005
R10376 gnd.n6210 gnd.n6209 9.3005
R10377 gnd.n6211 gnd.n521 9.3005
R10378 gnd.n6213 gnd.n6212 9.3005
R10379 gnd.n517 gnd.n516 9.3005
R10380 gnd.n6220 gnd.n6219 9.3005
R10381 gnd.n6221 gnd.n515 9.3005
R10382 gnd.n6223 gnd.n6222 9.3005
R10383 gnd.n511 gnd.n510 9.3005
R10384 gnd.n6230 gnd.n6229 9.3005
R10385 gnd.n6231 gnd.n509 9.3005
R10386 gnd.n6233 gnd.n6232 9.3005
R10387 gnd.n505 gnd.n504 9.3005
R10388 gnd.n6240 gnd.n6239 9.3005
R10389 gnd.n6241 gnd.n503 9.3005
R10390 gnd.n6243 gnd.n6242 9.3005
R10391 gnd.n499 gnd.n498 9.3005
R10392 gnd.n6250 gnd.n6249 9.3005
R10393 gnd.n6251 gnd.n497 9.3005
R10394 gnd.n6253 gnd.n6252 9.3005
R10395 gnd.n493 gnd.n492 9.3005
R10396 gnd.n6260 gnd.n6259 9.3005
R10397 gnd.n6261 gnd.n491 9.3005
R10398 gnd.n6263 gnd.n6262 9.3005
R10399 gnd.n487 gnd.n486 9.3005
R10400 gnd.n6270 gnd.n6269 9.3005
R10401 gnd.n6271 gnd.n485 9.3005
R10402 gnd.n6273 gnd.n6272 9.3005
R10403 gnd.n481 gnd.n480 9.3005
R10404 gnd.n6280 gnd.n6279 9.3005
R10405 gnd.n6281 gnd.n479 9.3005
R10406 gnd.n6283 gnd.n6282 9.3005
R10407 gnd.n475 gnd.n474 9.3005
R10408 gnd.n6290 gnd.n6289 9.3005
R10409 gnd.n6291 gnd.n473 9.3005
R10410 gnd.n6293 gnd.n6292 9.3005
R10411 gnd.n469 gnd.n468 9.3005
R10412 gnd.n6300 gnd.n6299 9.3005
R10413 gnd.n6301 gnd.n467 9.3005
R10414 gnd.n6303 gnd.n6302 9.3005
R10415 gnd.n463 gnd.n462 9.3005
R10416 gnd.n6310 gnd.n6309 9.3005
R10417 gnd.n6311 gnd.n461 9.3005
R10418 gnd.n6313 gnd.n6312 9.3005
R10419 gnd.n457 gnd.n456 9.3005
R10420 gnd.n6320 gnd.n6319 9.3005
R10421 gnd.n6321 gnd.n455 9.3005
R10422 gnd.n6323 gnd.n6322 9.3005
R10423 gnd.n451 gnd.n450 9.3005
R10424 gnd.n6330 gnd.n6329 9.3005
R10425 gnd.n6331 gnd.n449 9.3005
R10426 gnd.n6333 gnd.n6332 9.3005
R10427 gnd.n445 gnd.n444 9.3005
R10428 gnd.n6340 gnd.n6339 9.3005
R10429 gnd.n6341 gnd.n443 9.3005
R10430 gnd.n6343 gnd.n6342 9.3005
R10431 gnd.n439 gnd.n438 9.3005
R10432 gnd.n6350 gnd.n6349 9.3005
R10433 gnd.n6351 gnd.n437 9.3005
R10434 gnd.n6353 gnd.n6352 9.3005
R10435 gnd.n433 gnd.n432 9.3005
R10436 gnd.n6360 gnd.n6359 9.3005
R10437 gnd.n6361 gnd.n431 9.3005
R10438 gnd.n6363 gnd.n6362 9.3005
R10439 gnd.n427 gnd.n426 9.3005
R10440 gnd.n6370 gnd.n6369 9.3005
R10441 gnd.n6371 gnd.n425 9.3005
R10442 gnd.n6373 gnd.n6372 9.3005
R10443 gnd.n421 gnd.n420 9.3005
R10444 gnd.n6380 gnd.n6379 9.3005
R10445 gnd.n6381 gnd.n419 9.3005
R10446 gnd.n6383 gnd.n6382 9.3005
R10447 gnd.n415 gnd.n414 9.3005
R10448 gnd.n6390 gnd.n6389 9.3005
R10449 gnd.n6391 gnd.n413 9.3005
R10450 gnd.n6393 gnd.n6392 9.3005
R10451 gnd.n409 gnd.n408 9.3005
R10452 gnd.n6400 gnd.n6399 9.3005
R10453 gnd.n6401 gnd.n407 9.3005
R10454 gnd.n6403 gnd.n6402 9.3005
R10455 gnd.n403 gnd.n402 9.3005
R10456 gnd.n6410 gnd.n6409 9.3005
R10457 gnd.n6411 gnd.n401 9.3005
R10458 gnd.n6413 gnd.n6412 9.3005
R10459 gnd.n397 gnd.n396 9.3005
R10460 gnd.n6420 gnd.n6419 9.3005
R10461 gnd.n6421 gnd.n395 9.3005
R10462 gnd.n6423 gnd.n6422 9.3005
R10463 gnd.n391 gnd.n390 9.3005
R10464 gnd.n6430 gnd.n6429 9.3005
R10465 gnd.n6431 gnd.n389 9.3005
R10466 gnd.n6433 gnd.n6432 9.3005
R10467 gnd.n385 gnd.n384 9.3005
R10468 gnd.n6440 gnd.n6439 9.3005
R10469 gnd.n6441 gnd.n383 9.3005
R10470 gnd.n6443 gnd.n6442 9.3005
R10471 gnd.n379 gnd.n378 9.3005
R10472 gnd.n6450 gnd.n6449 9.3005
R10473 gnd.n6451 gnd.n377 9.3005
R10474 gnd.n6453 gnd.n6452 9.3005
R10475 gnd.n373 gnd.n372 9.3005
R10476 gnd.n6460 gnd.n6459 9.3005
R10477 gnd.n6461 gnd.n371 9.3005
R10478 gnd.n6463 gnd.n6462 9.3005
R10479 gnd.n367 gnd.n366 9.3005
R10480 gnd.n6470 gnd.n6469 9.3005
R10481 gnd.n6471 gnd.n365 9.3005
R10482 gnd.n6473 gnd.n6472 9.3005
R10483 gnd.n361 gnd.n360 9.3005
R10484 gnd.n6480 gnd.n6479 9.3005
R10485 gnd.n6481 gnd.n359 9.3005
R10486 gnd.n6483 gnd.n6482 9.3005
R10487 gnd.n355 gnd.n354 9.3005
R10488 gnd.n6490 gnd.n6489 9.3005
R10489 gnd.n6491 gnd.n353 9.3005
R10490 gnd.n6493 gnd.n6492 9.3005
R10491 gnd.n349 gnd.n348 9.3005
R10492 gnd.n6500 gnd.n6499 9.3005
R10493 gnd.n6501 gnd.n347 9.3005
R10494 gnd.n6503 gnd.n6502 9.3005
R10495 gnd.n343 gnd.n342 9.3005
R10496 gnd.n6510 gnd.n6509 9.3005
R10497 gnd.n6511 gnd.n341 9.3005
R10498 gnd.n6513 gnd.n6512 9.3005
R10499 gnd.n337 gnd.n336 9.3005
R10500 gnd.n6520 gnd.n6519 9.3005
R10501 gnd.n6521 gnd.n335 9.3005
R10502 gnd.n6523 gnd.n6522 9.3005
R10503 gnd.n331 gnd.n330 9.3005
R10504 gnd.n6530 gnd.n6529 9.3005
R10505 gnd.n6531 gnd.n329 9.3005
R10506 gnd.n6533 gnd.n6532 9.3005
R10507 gnd.n325 gnd.n324 9.3005
R10508 gnd.n6540 gnd.n6539 9.3005
R10509 gnd.n6541 gnd.n323 9.3005
R10510 gnd.n6543 gnd.n6542 9.3005
R10511 gnd.n319 gnd.n318 9.3005
R10512 gnd.n6550 gnd.n6549 9.3005
R10513 gnd.n6551 gnd.n317 9.3005
R10514 gnd.n6554 gnd.n6553 9.3005
R10515 gnd.n6552 gnd.n313 9.3005
R10516 gnd.n6560 gnd.n312 9.3005
R10517 gnd.n6562 gnd.n6561 9.3005
R10518 gnd.n308 gnd.n307 9.3005
R10519 gnd.n6571 gnd.n6570 9.3005
R10520 gnd.n6572 gnd.n306 9.3005
R10521 gnd.n6574 gnd.n6573 9.3005
R10522 gnd.n302 gnd.n301 9.3005
R10523 gnd.n6581 gnd.n6580 9.3005
R10524 gnd.n6582 gnd.n300 9.3005
R10525 gnd.n6584 gnd.n6583 9.3005
R10526 gnd.n296 gnd.n295 9.3005
R10527 gnd.n6591 gnd.n6590 9.3005
R10528 gnd.n6592 gnd.n294 9.3005
R10529 gnd.n6594 gnd.n6593 9.3005
R10530 gnd.n290 gnd.n289 9.3005
R10531 gnd.n6601 gnd.n6600 9.3005
R10532 gnd.n6602 gnd.n288 9.3005
R10533 gnd.n6604 gnd.n6603 9.3005
R10534 gnd.n284 gnd.n283 9.3005
R10535 gnd.n6611 gnd.n6610 9.3005
R10536 gnd.n6612 gnd.n282 9.3005
R10537 gnd.n6614 gnd.n6613 9.3005
R10538 gnd.n278 gnd.n277 9.3005
R10539 gnd.n6621 gnd.n6620 9.3005
R10540 gnd.n6622 gnd.n276 9.3005
R10541 gnd.n6624 gnd.n6623 9.3005
R10542 gnd.n272 gnd.n271 9.3005
R10543 gnd.n6631 gnd.n6630 9.3005
R10544 gnd.n6632 gnd.n270 9.3005
R10545 gnd.n6634 gnd.n6633 9.3005
R10546 gnd.n266 gnd.n265 9.3005
R10547 gnd.n6641 gnd.n6640 9.3005
R10548 gnd.n6642 gnd.n264 9.3005
R10549 gnd.n6644 gnd.n6643 9.3005
R10550 gnd.n260 gnd.n259 9.3005
R10551 gnd.n6651 gnd.n6650 9.3005
R10552 gnd.n6652 gnd.n258 9.3005
R10553 gnd.n6654 gnd.n6653 9.3005
R10554 gnd.n254 gnd.n253 9.3005
R10555 gnd.n6661 gnd.n6660 9.3005
R10556 gnd.n6662 gnd.n252 9.3005
R10557 gnd.n6664 gnd.n6663 9.3005
R10558 gnd.n248 gnd.n247 9.3005
R10559 gnd.n6671 gnd.n6670 9.3005
R10560 gnd.n6672 gnd.n246 9.3005
R10561 gnd.n6674 gnd.n6673 9.3005
R10562 gnd.n242 gnd.n241 9.3005
R10563 gnd.n6681 gnd.n6680 9.3005
R10564 gnd.n6682 gnd.n240 9.3005
R10565 gnd.n6684 gnd.n6683 9.3005
R10566 gnd.n236 gnd.n235 9.3005
R10567 gnd.n6691 gnd.n6690 9.3005
R10568 gnd.n6692 gnd.n234 9.3005
R10569 gnd.n6694 gnd.n6693 9.3005
R10570 gnd.n230 gnd.n229 9.3005
R10571 gnd.n6701 gnd.n6700 9.3005
R10572 gnd.n6702 gnd.n228 9.3005
R10573 gnd.n6704 gnd.n6703 9.3005
R10574 gnd.n224 gnd.n223 9.3005
R10575 gnd.n6711 gnd.n6710 9.3005
R10576 gnd.n6712 gnd.n222 9.3005
R10577 gnd.n6714 gnd.n6713 9.3005
R10578 gnd.n218 gnd.n217 9.3005
R10579 gnd.n6721 gnd.n6720 9.3005
R10580 gnd.n6722 gnd.n216 9.3005
R10581 gnd.n6724 gnd.n6723 9.3005
R10582 gnd.n212 gnd.n211 9.3005
R10583 gnd.n6731 gnd.n6730 9.3005
R10584 gnd.n6732 gnd.n210 9.3005
R10585 gnd.n6734 gnd.n6733 9.3005
R10586 gnd.n206 gnd.n205 9.3005
R10587 gnd.n6741 gnd.n6740 9.3005
R10588 gnd.n6742 gnd.n204 9.3005
R10589 gnd.n6744 gnd.n6743 9.3005
R10590 gnd.n200 gnd.n199 9.3005
R10591 gnd.n6751 gnd.n6750 9.3005
R10592 gnd.n6752 gnd.n198 9.3005
R10593 gnd.n6754 gnd.n6753 9.3005
R10594 gnd.n194 gnd.n193 9.3005
R10595 gnd.n6761 gnd.n6760 9.3005
R10596 gnd.n6762 gnd.n192 9.3005
R10597 gnd.n6764 gnd.n6763 9.3005
R10598 gnd.n188 gnd.n187 9.3005
R10599 gnd.n6772 gnd.n6771 9.3005
R10600 gnd.n6773 gnd.n186 9.3005
R10601 gnd.n6775 gnd.n6774 9.3005
R10602 gnd.n6564 gnd.n6563 9.3005
R10603 gnd.n7207 gnd.n7206 9.3005
R10604 gnd.n7205 gnd.n69 9.3005
R10605 gnd.n176 gnd.n71 9.3005
R10606 gnd.n6794 gnd.n6793 9.3005
R10607 gnd.n6795 gnd.n175 9.3005
R10608 gnd.n7114 gnd.n6796 9.3005
R10609 gnd.n7113 gnd.n6797 9.3005
R10610 gnd.n7112 gnd.n6798 9.3005
R10611 gnd.n7110 gnd.n6799 9.3005
R10612 gnd.n7109 gnd.n6800 9.3005
R10613 gnd.n7107 gnd.n6801 9.3005
R10614 gnd.n7106 gnd.n6802 9.3005
R10615 gnd.n7104 gnd.n6803 9.3005
R10616 gnd.n7103 gnd.n6804 9.3005
R10617 gnd.n7101 gnd.n6805 9.3005
R10618 gnd.n7100 gnd.n6806 9.3005
R10619 gnd.n7098 gnd.n6807 9.3005
R10620 gnd.n7097 gnd.n6808 9.3005
R10621 gnd.n7095 gnd.n6809 9.3005
R10622 gnd.n7094 gnd.n6810 9.3005
R10623 gnd.n7092 gnd.n7091 9.3005
R10624 gnd.n6835 gnd.n6831 9.3005
R10625 gnd.n6839 gnd.n6838 9.3005
R10626 gnd.n6840 gnd.n6830 9.3005
R10627 gnd.n6842 gnd.n6841 9.3005
R10628 gnd.n6845 gnd.n6829 9.3005
R10629 gnd.n6849 gnd.n6848 9.3005
R10630 gnd.n6850 gnd.n6828 9.3005
R10631 gnd.n6852 gnd.n6851 9.3005
R10632 gnd.n6855 gnd.n6827 9.3005
R10633 gnd.n6859 gnd.n6858 9.3005
R10634 gnd.n6860 gnd.n6826 9.3005
R10635 gnd.n6862 gnd.n6861 9.3005
R10636 gnd.n6865 gnd.n6825 9.3005
R10637 gnd.n6868 gnd.n6867 9.3005
R10638 gnd.n6869 gnd.n6824 9.3005
R10639 gnd.n6871 gnd.n6870 9.3005
R10640 gnd.n6814 gnd.n6811 9.3005
R10641 gnd.n7090 gnd.n7089 9.3005
R10642 gnd.n6833 gnd.n6832 9.3005
R10643 gnd.n6907 gnd.n6904 9.3005
R10644 gnd.n7083 gnd.n6908 9.3005
R10645 gnd.n7082 gnd.n6909 9.3005
R10646 gnd.n7081 gnd.n6910 9.3005
R10647 gnd.n7078 gnd.n6911 9.3005
R10648 gnd.n7077 gnd.n6912 9.3005
R10649 gnd.n7074 gnd.n6913 9.3005
R10650 gnd.n7073 gnd.n6914 9.3005
R10651 gnd.n7070 gnd.n6915 9.3005
R10652 gnd.n7069 gnd.n6916 9.3005
R10653 gnd.n7066 gnd.n6917 9.3005
R10654 gnd.n7065 gnd.n6918 9.3005
R10655 gnd.n7062 gnd.n6919 9.3005
R10656 gnd.n7061 gnd.n6920 9.3005
R10657 gnd.n7058 gnd.n6921 9.3005
R10658 gnd.n7057 gnd.n6922 9.3005
R10659 gnd.n7054 gnd.n6923 9.3005
R10660 gnd.n7050 gnd.n6924 9.3005
R10661 gnd.n7047 gnd.n6925 9.3005
R10662 gnd.n7046 gnd.n6926 9.3005
R10663 gnd.n7043 gnd.n6927 9.3005
R10664 gnd.n7042 gnd.n6928 9.3005
R10665 gnd.n7039 gnd.n6929 9.3005
R10666 gnd.n7038 gnd.n6930 9.3005
R10667 gnd.n7035 gnd.n6931 9.3005
R10668 gnd.n7034 gnd.n6932 9.3005
R10669 gnd.n7031 gnd.n6933 9.3005
R10670 gnd.n7030 gnd.n6934 9.3005
R10671 gnd.n7027 gnd.n6935 9.3005
R10672 gnd.n7026 gnd.n6936 9.3005
R10673 gnd.n7023 gnd.n6937 9.3005
R10674 gnd.n7022 gnd.n6938 9.3005
R10675 gnd.n7019 gnd.n6939 9.3005
R10676 gnd.n7018 gnd.n6940 9.3005
R10677 gnd.n7015 gnd.n6941 9.3005
R10678 gnd.n7014 gnd.n6942 9.3005
R10679 gnd.n7011 gnd.n7010 9.3005
R10680 gnd.n7009 gnd.n6943 9.3005
R10681 gnd.n7008 gnd.n7007 9.3005
R10682 gnd.n7004 gnd.n6946 9.3005
R10683 gnd.n7001 gnd.n6947 9.3005
R10684 gnd.n7000 gnd.n6948 9.3005
R10685 gnd.n6997 gnd.n6949 9.3005
R10686 gnd.n6996 gnd.n6950 9.3005
R10687 gnd.n6993 gnd.n6951 9.3005
R10688 gnd.n6992 gnd.n6952 9.3005
R10689 gnd.n6989 gnd.n6953 9.3005
R10690 gnd.n6988 gnd.n6954 9.3005
R10691 gnd.n6985 gnd.n6955 9.3005
R10692 gnd.n6984 gnd.n6956 9.3005
R10693 gnd.n6981 gnd.n6957 9.3005
R10694 gnd.n6980 gnd.n6958 9.3005
R10695 gnd.n6977 gnd.n6959 9.3005
R10696 gnd.n6976 gnd.n6960 9.3005
R10697 gnd.n6973 gnd.n6961 9.3005
R10698 gnd.n6972 gnd.n6962 9.3005
R10699 gnd.n6969 gnd.n6968 9.3005
R10700 gnd.n6967 gnd.n6964 9.3005
R10701 gnd.n6906 gnd.n6905 9.3005
R10702 gnd.n5373 gnd.n5372 9.3005
R10703 gnd.n1491 gnd.n1490 9.3005
R10704 gnd.n1515 gnd.n1514 9.3005
R10705 gnd.n5360 gnd.n1516 9.3005
R10706 gnd.n5359 gnd.n1517 9.3005
R10707 gnd.n5358 gnd.n1518 9.3005
R10708 gnd.n5190 gnd.n1519 9.3005
R10709 gnd.n5348 gnd.n1536 9.3005
R10710 gnd.n5347 gnd.n1537 9.3005
R10711 gnd.n5346 gnd.n1538 9.3005
R10712 gnd.n5196 gnd.n1539 9.3005
R10713 gnd.n5336 gnd.n1556 9.3005
R10714 gnd.n5335 gnd.n1557 9.3005
R10715 gnd.n5334 gnd.n1558 9.3005
R10716 gnd.n5273 gnd.n1559 9.3005
R10717 gnd.n5324 gnd.n1573 9.3005
R10718 gnd.n5323 gnd.n1574 9.3005
R10719 gnd.n5322 gnd.n1575 9.3005
R10720 gnd.n5293 gnd.n1576 9.3005
R10721 gnd.n5295 gnd.n5294 9.3005
R10722 gnd.n1600 gnd.n1599 9.3005
R10723 gnd.n5304 gnd.n5303 9.3005
R10724 gnd.n180 gnd.n179 9.3005
R10725 gnd.n6787 gnd.n6786 9.3005
R10726 gnd.n6788 gnd.n96 9.3005
R10727 gnd.n7193 gnd.n97 9.3005
R10728 gnd.n7192 gnd.n98 9.3005
R10729 gnd.n7191 gnd.n99 9.3005
R10730 gnd.n7120 gnd.n100 9.3005
R10731 gnd.n7181 gnd.n115 9.3005
R10732 gnd.n7180 gnd.n116 9.3005
R10733 gnd.n7179 gnd.n117 9.3005
R10734 gnd.n7127 gnd.n118 9.3005
R10735 gnd.n7169 gnd.n135 9.3005
R10736 gnd.n7168 gnd.n136 9.3005
R10737 gnd.n7167 gnd.n137 9.3005
R10738 gnd.n7134 gnd.n138 9.3005
R10739 gnd.n7157 gnd.n154 9.3005
R10740 gnd.n7156 gnd.n155 9.3005
R10741 gnd.n7155 gnd.n156 9.3005
R10742 gnd.n172 gnd.n157 9.3005
R10743 gnd.n7145 gnd.n7144 9.3005
R10744 gnd.n5374 gnd.n1489 9.3005
R10745 gnd.n5372 gnd.n5371 9.3005
R10746 gnd.n5370 gnd.n1491 9.3005
R10747 gnd.n1515 gnd.n1492 9.3005
R10748 gnd.n5185 gnd.n1516 9.3005
R10749 gnd.n5188 gnd.n1517 9.3005
R10750 gnd.n5189 gnd.n1518 9.3005
R10751 gnd.n5194 gnd.n5190 9.3005
R10752 gnd.n5195 gnd.n1536 9.3005
R10753 gnd.n5199 gnd.n1537 9.3005
R10754 gnd.n5198 gnd.n1538 9.3005
R10755 gnd.n5197 gnd.n5196 9.3005
R10756 gnd.n1611 gnd.n1556 9.3005
R10757 gnd.n5271 gnd.n1557 9.3005
R10758 gnd.n5272 gnd.n1558 9.3005
R10759 gnd.n5274 gnd.n5273 9.3005
R10760 gnd.n1605 gnd.n1573 9.3005
R10761 gnd.n5290 gnd.n1574 9.3005
R10762 gnd.n5291 gnd.n1575 9.3005
R10763 gnd.n5293 gnd.n5292 9.3005
R10764 gnd.n5294 gnd.n1601 9.3005
R10765 gnd.n5300 gnd.n1600 9.3005
R10766 gnd.n5303 gnd.n5302 9.3005
R10767 gnd.n5301 gnd.n179 9.3005
R10768 gnd.n6787 gnd.n178 9.3005
R10769 gnd.n6789 gnd.n6788 9.3005
R10770 gnd.n174 gnd.n97 9.3005
R10771 gnd.n7118 gnd.n98 9.3005
R10772 gnd.n7119 gnd.n99 9.3005
R10773 gnd.n7122 gnd.n7120 9.3005
R10774 gnd.n7123 gnd.n115 9.3005
R10775 gnd.n7125 gnd.n116 9.3005
R10776 gnd.n7126 gnd.n117 9.3005
R10777 gnd.n7129 gnd.n7127 9.3005
R10778 gnd.n7130 gnd.n135 9.3005
R10779 gnd.n7132 gnd.n136 9.3005
R10780 gnd.n7133 gnd.n137 9.3005
R10781 gnd.n7136 gnd.n7134 9.3005
R10782 gnd.n7137 gnd.n154 9.3005
R10783 gnd.n7139 gnd.n155 9.3005
R10784 gnd.n7140 gnd.n156 9.3005
R10785 gnd.n7142 gnd.n172 9.3005
R10786 gnd.n7144 gnd.n7143 9.3005
R10787 gnd.n1489 gnd.n1483 9.3005
R10788 gnd.n5384 gnd.n5383 9.3005
R10789 gnd.n5387 gnd.n1481 9.3005
R10790 gnd.n5388 gnd.n1480 9.3005
R10791 gnd.n5391 gnd.n1479 9.3005
R10792 gnd.n5392 gnd.n1478 9.3005
R10793 gnd.n5395 gnd.n1477 9.3005
R10794 gnd.n5396 gnd.n1476 9.3005
R10795 gnd.n5399 gnd.n1475 9.3005
R10796 gnd.n5400 gnd.n1474 9.3005
R10797 gnd.n5403 gnd.n1473 9.3005
R10798 gnd.n5404 gnd.n1472 9.3005
R10799 gnd.n5407 gnd.n1471 9.3005
R10800 gnd.n5408 gnd.n1470 9.3005
R10801 gnd.n5411 gnd.n1469 9.3005
R10802 gnd.n5412 gnd.n1468 9.3005
R10803 gnd.n5415 gnd.n1467 9.3005
R10804 gnd.n5416 gnd.n1466 9.3005
R10805 gnd.n5419 gnd.n1465 9.3005
R10806 gnd.n5420 gnd.n1464 9.3005
R10807 gnd.n5423 gnd.n1463 9.3005
R10808 gnd.n5427 gnd.n1459 9.3005
R10809 gnd.n5428 gnd.n1458 9.3005
R10810 gnd.n5431 gnd.n1457 9.3005
R10811 gnd.n5432 gnd.n1456 9.3005
R10812 gnd.n5435 gnd.n1455 9.3005
R10813 gnd.n5436 gnd.n1454 9.3005
R10814 gnd.n5439 gnd.n1453 9.3005
R10815 gnd.n5440 gnd.n1452 9.3005
R10816 gnd.n5443 gnd.n1451 9.3005
R10817 gnd.n5445 gnd.n1447 9.3005
R10818 gnd.n5448 gnd.n1446 9.3005
R10819 gnd.n5449 gnd.n1445 9.3005
R10820 gnd.n5452 gnd.n1444 9.3005
R10821 gnd.n5453 gnd.n1443 9.3005
R10822 gnd.n5456 gnd.n1442 9.3005
R10823 gnd.n5457 gnd.n1441 9.3005
R10824 gnd.n5460 gnd.n1440 9.3005
R10825 gnd.n5462 gnd.n1437 9.3005
R10826 gnd.n5465 gnd.n1436 9.3005
R10827 gnd.n5466 gnd.n1435 9.3005
R10828 gnd.n5469 gnd.n1434 9.3005
R10829 gnd.n5470 gnd.n1433 9.3005
R10830 gnd.n5473 gnd.n1432 9.3005
R10831 gnd.n5474 gnd.n1431 9.3005
R10832 gnd.n5477 gnd.n1430 9.3005
R10833 gnd.n5478 gnd.n1429 9.3005
R10834 gnd.n5481 gnd.n1428 9.3005
R10835 gnd.n5482 gnd.n1427 9.3005
R10836 gnd.n5485 gnd.n1426 9.3005
R10837 gnd.n5486 gnd.n1425 9.3005
R10838 gnd.n5489 gnd.n1424 9.3005
R10839 gnd.n5491 gnd.n1423 9.3005
R10840 gnd.n5492 gnd.n1422 9.3005
R10841 gnd.n5493 gnd.n1421 9.3005
R10842 gnd.n5494 gnd.n1420 9.3005
R10843 gnd.n5424 gnd.n1460 9.3005
R10844 gnd.n5382 gnd.n5379 9.3005
R10845 gnd.n1502 gnd.n1499 9.3005
R10846 gnd.n5366 gnd.n1503 9.3005
R10847 gnd.n5365 gnd.n1504 9.3005
R10848 gnd.n5364 gnd.n1505 9.3005
R10849 gnd.n1525 gnd.n1506 9.3005
R10850 gnd.n5354 gnd.n1526 9.3005
R10851 gnd.n5353 gnd.n1527 9.3005
R10852 gnd.n5352 gnd.n1528 9.3005
R10853 gnd.n1546 gnd.n1529 9.3005
R10854 gnd.n5342 gnd.n1547 9.3005
R10855 gnd.n5341 gnd.n1548 9.3005
R10856 gnd.n5340 gnd.n1549 9.3005
R10857 gnd.n1565 gnd.n1550 9.3005
R10858 gnd.n5330 gnd.n1566 9.3005
R10859 gnd.n5329 gnd.n82 9.3005
R10860 gnd.n87 gnd.n81 9.3005
R10861 gnd.n7187 gnd.n106 9.3005
R10862 gnd.n7186 gnd.n107 9.3005
R10863 gnd.n7185 gnd.n108 9.3005
R10864 gnd.n124 gnd.n109 9.3005
R10865 gnd.n7175 gnd.n125 9.3005
R10866 gnd.n7174 gnd.n126 9.3005
R10867 gnd.n7173 gnd.n127 9.3005
R10868 gnd.n144 gnd.n128 9.3005
R10869 gnd.n7163 gnd.n145 9.3005
R10870 gnd.n7162 gnd.n146 9.3005
R10871 gnd.n7161 gnd.n147 9.3005
R10872 gnd.n162 gnd.n148 9.3005
R10873 gnd.n7151 gnd.n163 9.3005
R10874 gnd.n7150 gnd.n164 9.3005
R10875 gnd.n7149 gnd.n165 9.3005
R10876 gnd.n1501 gnd.n1500 9.3005
R10877 gnd.n7198 gnd.n7197 9.3005
R10878 gnd.n4128 gnd.n4127 9.3005
R10879 gnd.n4150 gnd.n4129 9.3005
R10880 gnd.n4149 gnd.n4130 9.3005
R10881 gnd.n4148 gnd.n4131 9.3005
R10882 gnd.n4134 gnd.n4132 9.3005
R10883 gnd.n4144 gnd.n4135 9.3005
R10884 gnd.n4143 gnd.n4136 9.3005
R10885 gnd.n4142 gnd.n4137 9.3005
R10886 gnd.n4140 gnd.n4139 9.3005
R10887 gnd.n4138 gnd.n2094 9.3005
R10888 gnd.n2092 gnd.n2091 9.3005
R10889 gnd.n4205 gnd.n4204 9.3005
R10890 gnd.n4206 gnd.n2090 9.3005
R10891 gnd.n4208 gnd.n4207 9.3005
R10892 gnd.n2088 gnd.n2087 9.3005
R10893 gnd.n4213 gnd.n4212 9.3005
R10894 gnd.n4214 gnd.n2086 9.3005
R10895 gnd.n4216 gnd.n4215 9.3005
R10896 gnd.n2084 gnd.n2083 9.3005
R10897 gnd.n4222 gnd.n4221 9.3005
R10898 gnd.n4223 gnd.n2082 9.3005
R10899 gnd.n4225 gnd.n4224 9.3005
R10900 gnd.n2080 gnd.n2079 9.3005
R10901 gnd.n4307 gnd.n4306 9.3005
R10902 gnd.n4308 gnd.n2078 9.3005
R10903 gnd.n4310 gnd.n4309 9.3005
R10904 gnd.n2065 gnd.n2064 9.3005
R10905 gnd.n4323 gnd.n4322 9.3005
R10906 gnd.n4324 gnd.n2063 9.3005
R10907 gnd.n4326 gnd.n4325 9.3005
R10908 gnd.n2052 gnd.n2051 9.3005
R10909 gnd.n4339 gnd.n4338 9.3005
R10910 gnd.n4340 gnd.n2050 9.3005
R10911 gnd.n4342 gnd.n4341 9.3005
R10912 gnd.n2038 gnd.n2037 9.3005
R10913 gnd.n4355 gnd.n4354 9.3005
R10914 gnd.n4356 gnd.n2036 9.3005
R10915 gnd.n4358 gnd.n4357 9.3005
R10916 gnd.n2024 gnd.n2023 9.3005
R10917 gnd.n4371 gnd.n4370 9.3005
R10918 gnd.n4372 gnd.n2022 9.3005
R10919 gnd.n4374 gnd.n4373 9.3005
R10920 gnd.n2010 gnd.n2009 9.3005
R10921 gnd.n4387 gnd.n4386 9.3005
R10922 gnd.n4388 gnd.n2008 9.3005
R10923 gnd.n4390 gnd.n4389 9.3005
R10924 gnd.n1995 gnd.n1994 9.3005
R10925 gnd.n4404 gnd.n4403 9.3005
R10926 gnd.n4405 gnd.n1993 9.3005
R10927 gnd.n4413 gnd.n4406 9.3005
R10928 gnd.n4412 gnd.n4407 9.3005
R10929 gnd.n4411 gnd.n4409 9.3005
R10930 gnd.n4408 gnd.n1207 9.3005
R10931 gnd.n5675 gnd.n1208 9.3005
R10932 gnd.n5674 gnd.n1209 9.3005
R10933 gnd.n5673 gnd.n1210 9.3005
R10934 gnd.n1964 gnd.n1211 9.3005
R10935 gnd.n1966 gnd.n1965 9.3005
R10936 gnd.n4562 gnd.n4561 9.3005
R10937 gnd.n4563 gnd.n1963 9.3005
R10938 gnd.n4565 gnd.n4564 9.3005
R10939 gnd.n1938 gnd.n1937 9.3005
R10940 gnd.n4605 gnd.n4604 9.3005
R10941 gnd.n4606 gnd.n1936 9.3005
R10942 gnd.n4610 gnd.n4607 9.3005
R10943 gnd.n4609 gnd.n4608 9.3005
R10944 gnd.n1917 gnd.n1916 9.3005
R10945 gnd.n4665 gnd.n4664 9.3005
R10946 gnd.n4666 gnd.n1915 9.3005
R10947 gnd.n4679 gnd.n4667 9.3005
R10948 gnd.n4678 gnd.n4668 9.3005
R10949 gnd.n4677 gnd.n4669 9.3005
R10950 gnd.n4671 gnd.n4670 9.3005
R10951 gnd.n4673 gnd.n4672 9.3005
R10952 gnd.n1880 gnd.n1879 9.3005
R10953 gnd.n4726 gnd.n4725 9.3005
R10954 gnd.n4727 gnd.n1878 9.3005
R10955 gnd.n4729 gnd.n4728 9.3005
R10956 gnd.n1857 gnd.n1856 9.3005
R10957 gnd.n4772 gnd.n4771 9.3005
R10958 gnd.n4773 gnd.n1855 9.3005
R10959 gnd.n4777 gnd.n4774 9.3005
R10960 gnd.n4776 gnd.n4775 9.3005
R10961 gnd.n1836 gnd.n1835 9.3005
R10962 gnd.n4824 gnd.n4823 9.3005
R10963 gnd.n4825 gnd.n1834 9.3005
R10964 gnd.n4829 gnd.n4826 9.3005
R10965 gnd.n4828 gnd.n4827 9.3005
R10966 gnd.n1809 gnd.n1808 9.3005
R10967 gnd.n4860 gnd.n4859 9.3005
R10968 gnd.n4861 gnd.n1807 9.3005
R10969 gnd.n4863 gnd.n4862 9.3005
R10970 gnd.n1753 gnd.n1752 9.3005
R10971 gnd.n5035 gnd.n5034 9.3005
R10972 gnd.n5036 gnd.n1751 9.3005
R10973 gnd.n5038 gnd.n5037 9.3005
R10974 gnd.n1741 gnd.n1740 9.3005
R10975 gnd.n5051 gnd.n5050 9.3005
R10976 gnd.n5052 gnd.n1739 9.3005
R10977 gnd.n5054 gnd.n5053 9.3005
R10978 gnd.n1728 gnd.n1727 9.3005
R10979 gnd.n5068 gnd.n5067 9.3005
R10980 gnd.n5069 gnd.n1726 9.3005
R10981 gnd.n5071 gnd.n5070 9.3005
R10982 gnd.n1716 gnd.n1715 9.3005
R10983 gnd.n5084 gnd.n5083 9.3005
R10984 gnd.n5085 gnd.n1714 9.3005
R10985 gnd.n5087 gnd.n5086 9.3005
R10986 gnd.n1703 gnd.n1702 9.3005
R10987 gnd.n5100 gnd.n5099 9.3005
R10988 gnd.n5101 gnd.n1701 9.3005
R10989 gnd.n5103 gnd.n5102 9.3005
R10990 gnd.n1690 gnd.n1689 9.3005
R10991 gnd.n5116 gnd.n5115 9.3005
R10992 gnd.n5117 gnd.n1688 9.3005
R10993 gnd.n5119 gnd.n5118 9.3005
R10994 gnd.n1677 gnd.n1676 9.3005
R10995 gnd.n5132 gnd.n5131 9.3005
R10996 gnd.n5133 gnd.n1675 9.3005
R10997 gnd.n5138 gnd.n5134 9.3005
R10998 gnd.n5137 gnd.n5136 9.3005
R10999 gnd.n5135 gnd.n1664 9.3005
R11000 gnd.n5151 gnd.n1663 9.3005
R11001 gnd.n5153 gnd.n5152 9.3005
R11002 gnd.n5154 gnd.n1662 9.3005
R11003 gnd.n5167 gnd.n5155 9.3005
R11004 gnd.n5166 gnd.n5156 9.3005
R11005 gnd.n5165 gnd.n5157 9.3005
R11006 gnd.n5159 gnd.n5158 9.3005
R11007 gnd.n5161 gnd.n5160 9.3005
R11008 gnd.n1628 gnd.n1627 9.3005
R11009 gnd.n5222 gnd.n5221 9.3005
R11010 gnd.n5223 gnd.n1626 9.3005
R11011 gnd.n5225 gnd.n5224 9.3005
R11012 gnd.n1624 gnd.n1623 9.3005
R11013 gnd.n5230 gnd.n5229 9.3005
R11014 gnd.n5231 gnd.n1622 9.3005
R11015 gnd.n5233 gnd.n5232 9.3005
R11016 gnd.n1620 gnd.n1619 9.3005
R11017 gnd.n5238 gnd.n5237 9.3005
R11018 gnd.n5239 gnd.n1618 9.3005
R11019 gnd.n5258 gnd.n5240 9.3005
R11020 gnd.n5257 gnd.n5241 9.3005
R11021 gnd.n5256 gnd.n5242 9.3005
R11022 gnd.n5245 gnd.n5243 9.3005
R11023 gnd.n5252 gnd.n5246 9.3005
R11024 gnd.n6778 gnd.n184 9.3005
R11025 gnd.n4096 gnd.n4095 9.3005
R11026 gnd.n3742 gnd.n3739 9.3005
R11027 gnd.n3741 gnd.n3740 9.3005
R11028 gnd.n2183 gnd.n2182 9.3005
R11029 gnd.n3992 gnd.n3991 9.3005
R11030 gnd.n3993 gnd.n2181 9.3005
R11031 gnd.n3997 gnd.n3994 9.3005
R11032 gnd.n3996 gnd.n3995 9.3005
R11033 gnd.n2158 gnd.n2157 9.3005
R11034 gnd.n4027 gnd.n4026 9.3005
R11035 gnd.n4028 gnd.n2156 9.3005
R11036 gnd.n4034 gnd.n4029 9.3005
R11037 gnd.n4033 gnd.n4030 9.3005
R11038 gnd.n4032 gnd.n4031 9.3005
R11039 gnd.n2132 gnd.n2131 9.3005
R11040 gnd.n4067 gnd.n4066 9.3005
R11041 gnd.n4068 gnd.n2130 9.3005
R11042 gnd.n4070 gnd.n4069 9.3005
R11043 gnd.n2127 gnd.n2126 9.3005
R11044 gnd.n4093 gnd.n4092 9.3005
R11045 gnd.n4094 gnd.n2125 9.3005
R11046 gnd.n3738 gnd.n3670 9.3005
R11047 gnd.n3731 gnd.n3730 9.3005
R11048 gnd.n3729 gnd.n3676 9.3005
R11049 gnd.n3728 gnd.n3727 9.3005
R11050 gnd.n3678 gnd.n3677 9.3005
R11051 gnd.n3721 gnd.n3720 9.3005
R11052 gnd.n3719 gnd.n3680 9.3005
R11053 gnd.n3718 gnd.n3717 9.3005
R11054 gnd.n3682 gnd.n3681 9.3005
R11055 gnd.n3711 gnd.n3710 9.3005
R11056 gnd.n3709 gnd.n3684 9.3005
R11057 gnd.n3708 gnd.n3707 9.3005
R11058 gnd.n3686 gnd.n3685 9.3005
R11059 gnd.n3701 gnd.n3700 9.3005
R11060 gnd.n3699 gnd.n3688 9.3005
R11061 gnd.n3698 gnd.n3697 9.3005
R11062 gnd.n3692 gnd.n3689 9.3005
R11063 gnd.n3691 gnd.n3690 9.3005
R11064 gnd.n3674 gnd.n3671 9.3005
R11065 gnd.n3737 gnd.n3736 9.3005
R11066 gnd.n5753 gnd.n1039 9.3005
R11067 gnd.n5756 gnd.n1038 9.3005
R11068 gnd.n5757 gnd.n1037 9.3005
R11069 gnd.n5760 gnd.n1036 9.3005
R11070 gnd.n5761 gnd.n1035 9.3005
R11071 gnd.n5764 gnd.n1034 9.3005
R11072 gnd.n5765 gnd.n1033 9.3005
R11073 gnd.n5768 gnd.n1032 9.3005
R11074 gnd.n5770 gnd.n1029 9.3005
R11075 gnd.n5773 gnd.n1028 9.3005
R11076 gnd.n5774 gnd.n1027 9.3005
R11077 gnd.n5777 gnd.n1026 9.3005
R11078 gnd.n5778 gnd.n1025 9.3005
R11079 gnd.n5781 gnd.n1024 9.3005
R11080 gnd.n5782 gnd.n1023 9.3005
R11081 gnd.n5785 gnd.n1022 9.3005
R11082 gnd.n5786 gnd.n1021 9.3005
R11083 gnd.n5789 gnd.n1020 9.3005
R11084 gnd.n5790 gnd.n1019 9.3005
R11085 gnd.n5793 gnd.n1018 9.3005
R11086 gnd.n5794 gnd.n1017 9.3005
R11087 gnd.n5797 gnd.n1016 9.3005
R11088 gnd.n5798 gnd.n1015 9.3005
R11089 gnd.n5799 gnd.n1014 9.3005
R11090 gnd.n1013 gnd.n1010 9.3005
R11091 gnd.n1012 gnd.n1011 9.3005
R11092 gnd.n1136 gnd.n1135 9.3005
R11093 gnd.n1132 gnd.n1042 9.3005
R11094 gnd.n1129 gnd.n1043 9.3005
R11095 gnd.n1128 gnd.n1044 9.3005
R11096 gnd.n1125 gnd.n1045 9.3005
R11097 gnd.n1124 gnd.n1046 9.3005
R11098 gnd.n1121 gnd.n1047 9.3005
R11099 gnd.n1120 gnd.n1048 9.3005
R11100 gnd.n1117 gnd.n1116 9.3005
R11101 gnd.n1115 gnd.n1049 9.3005
R11102 gnd.n1114 gnd.n1113 9.3005
R11103 gnd.n1110 gnd.n1052 9.3005
R11104 gnd.n1107 gnd.n1053 9.3005
R11105 gnd.n1106 gnd.n1054 9.3005
R11106 gnd.n1103 gnd.n1055 9.3005
R11107 gnd.n1102 gnd.n1056 9.3005
R11108 gnd.n1099 gnd.n1057 9.3005
R11109 gnd.n1098 gnd.n1058 9.3005
R11110 gnd.n1095 gnd.n1059 9.3005
R11111 gnd.n1094 gnd.n1060 9.3005
R11112 gnd.n1091 gnd.n1061 9.3005
R11113 gnd.n1090 gnd.n1062 9.3005
R11114 gnd.n1087 gnd.n1063 9.3005
R11115 gnd.n1086 gnd.n1064 9.3005
R11116 gnd.n1083 gnd.n1065 9.3005
R11117 gnd.n1082 gnd.n1066 9.3005
R11118 gnd.n1079 gnd.n1067 9.3005
R11119 gnd.n1078 gnd.n1068 9.3005
R11120 gnd.n1075 gnd.n1074 9.3005
R11121 gnd.n1073 gnd.n1070 9.3005
R11122 gnd.n1137 gnd.n1040 9.3005
R11123 gnd.n3965 gnd.n2198 9.3005
R11124 gnd.n3977 gnd.n2199 9.3005
R11125 gnd.n3976 gnd.n2200 9.3005
R11126 gnd.n3975 gnd.n3971 9.3005
R11127 gnd.n3974 gnd.n3972 9.3005
R11128 gnd.n2177 gnd.n2173 9.3005
R11129 gnd.n4012 gnd.n2174 9.3005
R11130 gnd.n4011 gnd.n2175 9.3005
R11131 gnd.n4010 gnd.n4006 9.3005
R11132 gnd.n4009 gnd.n4007 9.3005
R11133 gnd.n2152 gnd.n2147 9.3005
R11134 gnd.n4052 gnd.n2148 9.3005
R11135 gnd.n4051 gnd.n2149 9.3005
R11136 gnd.n4050 gnd.n2150 9.3005
R11137 gnd.n4049 gnd.n4045 9.3005
R11138 gnd.n4047 gnd.n4046 9.3005
R11139 gnd.n2129 gnd.n750 9.3005
R11140 gnd.n5957 gnd.n751 9.3005
R11141 gnd.n5956 gnd.n752 9.3005
R11142 gnd.n5955 gnd.n753 9.3005
R11143 gnd.n2124 gnd.n754 9.3005
R11144 gnd.n5944 gnd.n767 9.3005
R11145 gnd.n5943 gnd.n768 9.3005
R11146 gnd.n5942 gnd.n769 9.3005
R11147 gnd.n4104 gnd.n770 9.3005
R11148 gnd.n5931 gnd.n785 9.3005
R11149 gnd.n5930 gnd.n786 9.3005
R11150 gnd.n5929 gnd.n787 9.3005
R11151 gnd.n2108 gnd.n788 9.3005
R11152 gnd.n5919 gnd.n804 9.3005
R11153 gnd.n5918 gnd.n805 9.3005
R11154 gnd.n5917 gnd.n806 9.3005
R11155 gnd.n2102 gnd.n807 9.3005
R11156 gnd.n5907 gnd.n825 9.3005
R11157 gnd.n5906 gnd.n826 9.3005
R11158 gnd.n5905 gnd.n827 9.3005
R11159 gnd.n4181 gnd.n828 9.3005
R11160 gnd.n5895 gnd.n845 9.3005
R11161 gnd.n5894 gnd.n846 9.3005
R11162 gnd.n5893 gnd.n847 9.3005
R11163 gnd.n864 gnd.n848 9.3005
R11164 gnd.n5883 gnd.n5882 9.3005
R11165 gnd.n3964 gnd.n3963 9.3005
R11166 gnd.n3966 gnd.n3965 9.3005
R11167 gnd.n3967 gnd.n2199 9.3005
R11168 gnd.n3969 gnd.n2200 9.3005
R11169 gnd.n3971 gnd.n3970 9.3005
R11170 gnd.n3972 gnd.n2176 9.3005
R11171 gnd.n4001 gnd.n2177 9.3005
R11172 gnd.n4002 gnd.n2174 9.3005
R11173 gnd.n4004 gnd.n2175 9.3005
R11174 gnd.n4006 gnd.n4005 9.3005
R11175 gnd.n4007 gnd.n2151 9.3005
R11176 gnd.n4038 gnd.n2152 9.3005
R11177 gnd.n4039 gnd.n2148 9.3005
R11178 gnd.n4041 gnd.n2149 9.3005
R11179 gnd.n4042 gnd.n2150 9.3005
R11180 gnd.n4045 gnd.n4044 9.3005
R11181 gnd.n4046 gnd.n2128 9.3005
R11182 gnd.n4074 gnd.n2129 9.3005
R11183 gnd.n4075 gnd.n751 9.3005
R11184 gnd.n4076 gnd.n752 9.3005
R11185 gnd.n2123 gnd.n753 9.3005
R11186 gnd.n4100 gnd.n2124 9.3005
R11187 gnd.n4101 gnd.n767 9.3005
R11188 gnd.n4102 gnd.n768 9.3005
R11189 gnd.n4103 gnd.n769 9.3005
R11190 gnd.n4107 gnd.n4104 9.3005
R11191 gnd.n4106 gnd.n785 9.3005
R11192 gnd.n4105 gnd.n786 9.3005
R11193 gnd.n2107 gnd.n787 9.3005
R11194 gnd.n4163 gnd.n2108 9.3005
R11195 gnd.n4164 gnd.n804 9.3005
R11196 gnd.n4165 gnd.n805 9.3005
R11197 gnd.n2101 gnd.n806 9.3005
R11198 gnd.n4177 gnd.n2102 9.3005
R11199 gnd.n4178 gnd.n825 9.3005
R11200 gnd.n4179 gnd.n826 9.3005
R11201 gnd.n4180 gnd.n827 9.3005
R11202 gnd.n4184 gnd.n4181 9.3005
R11203 gnd.n4185 gnd.n845 9.3005
R11204 gnd.n4186 gnd.n846 9.3005
R11205 gnd.n866 gnd.n847 9.3005
R11206 gnd.n5880 gnd.n864 9.3005
R11207 gnd.n5882 gnd.n5881 9.3005
R11208 gnd.n3964 gnd.n2201 9.3005
R11209 gnd.n3838 gnd.n3837 9.3005
R11210 gnd.n3846 gnd.n3834 9.3005
R11211 gnd.n3847 gnd.n3833 9.3005
R11212 gnd.n3848 gnd.n3832 9.3005
R11213 gnd.n3831 gnd.n3829 9.3005
R11214 gnd.n3854 gnd.n3828 9.3005
R11215 gnd.n3855 gnd.n3827 9.3005
R11216 gnd.n3856 gnd.n3826 9.3005
R11217 gnd.n3825 gnd.n3823 9.3005
R11218 gnd.n3862 gnd.n3822 9.3005
R11219 gnd.n3863 gnd.n3821 9.3005
R11220 gnd.n3864 gnd.n3820 9.3005
R11221 gnd.n3819 gnd.n3817 9.3005
R11222 gnd.n3870 gnd.n3816 9.3005
R11223 gnd.n3871 gnd.n3815 9.3005
R11224 gnd.n3872 gnd.n3814 9.3005
R11225 gnd.n3813 gnd.n3811 9.3005
R11226 gnd.n3878 gnd.n3810 9.3005
R11227 gnd.n3879 gnd.n3809 9.3005
R11228 gnd.n3880 gnd.n3808 9.3005
R11229 gnd.n3886 gnd.n3802 9.3005
R11230 gnd.n3887 gnd.n3801 9.3005
R11231 gnd.n3888 gnd.n3800 9.3005
R11232 gnd.n3799 gnd.n3797 9.3005
R11233 gnd.n3894 gnd.n3796 9.3005
R11234 gnd.n3895 gnd.n3795 9.3005
R11235 gnd.n3896 gnd.n3794 9.3005
R11236 gnd.n3793 gnd.n3791 9.3005
R11237 gnd.n3902 gnd.n3790 9.3005
R11238 gnd.n3903 gnd.n3789 9.3005
R11239 gnd.n3904 gnd.n3788 9.3005
R11240 gnd.n3787 gnd.n3785 9.3005
R11241 gnd.n3910 gnd.n3784 9.3005
R11242 gnd.n3911 gnd.n3783 9.3005
R11243 gnd.n3912 gnd.n3782 9.3005
R11244 gnd.n3781 gnd.n3779 9.3005
R11245 gnd.n3918 gnd.n3778 9.3005
R11246 gnd.n3919 gnd.n3777 9.3005
R11247 gnd.n3920 gnd.n3776 9.3005
R11248 gnd.n3775 gnd.n3770 9.3005
R11249 gnd.n3926 gnd.n3769 9.3005
R11250 gnd.n3927 gnd.n3768 9.3005
R11251 gnd.n3928 gnd.n3767 9.3005
R11252 gnd.n3766 gnd.n3764 9.3005
R11253 gnd.n3934 gnd.n3763 9.3005
R11254 gnd.n3935 gnd.n3762 9.3005
R11255 gnd.n3936 gnd.n3761 9.3005
R11256 gnd.n3760 gnd.n3758 9.3005
R11257 gnd.n3942 gnd.n3757 9.3005
R11258 gnd.n3943 gnd.n3756 9.3005
R11259 gnd.n3944 gnd.n3755 9.3005
R11260 gnd.n3754 gnd.n3752 9.3005
R11261 gnd.n3949 gnd.n3751 9.3005
R11262 gnd.n3950 gnd.n3750 9.3005
R11263 gnd.n3749 gnd.n3747 9.3005
R11264 gnd.n3955 gnd.n3746 9.3005
R11265 gnd.n3957 gnd.n3956 9.3005
R11266 gnd.n3807 gnd.n3805 9.3005
R11267 gnd.n3840 gnd.n3839 9.3005
R11268 gnd.n2192 gnd.n2191 9.3005
R11269 gnd.n3982 gnd.n3981 9.3005
R11270 gnd.n3983 gnd.n2190 9.3005
R11271 gnd.n3987 gnd.n3984 9.3005
R11272 gnd.n3986 gnd.n3985 9.3005
R11273 gnd.n2167 gnd.n2166 9.3005
R11274 gnd.n4017 gnd.n4016 9.3005
R11275 gnd.n4018 gnd.n2165 9.3005
R11276 gnd.n4022 gnd.n4019 9.3005
R11277 gnd.n4021 gnd.n4020 9.3005
R11278 gnd.n2140 gnd.n2139 9.3005
R11279 gnd.n4057 gnd.n4056 9.3005
R11280 gnd.n4058 gnd.n2138 9.3005
R11281 gnd.n4061 gnd.n4060 9.3005
R11282 gnd.n4059 gnd.n740 9.3005
R11283 gnd.n794 gnd.n778 9.3005
R11284 gnd.n5925 gnd.n795 9.3005
R11285 gnd.n5924 gnd.n796 9.3005
R11286 gnd.n5923 gnd.n797 9.3005
R11287 gnd.n814 gnd.n798 9.3005
R11288 gnd.n5913 gnd.n815 9.3005
R11289 gnd.n5912 gnd.n816 9.3005
R11290 gnd.n5911 gnd.n817 9.3005
R11291 gnd.n834 gnd.n818 9.3005
R11292 gnd.n5901 gnd.n835 9.3005
R11293 gnd.n5900 gnd.n836 9.3005
R11294 gnd.n5899 gnd.n837 9.3005
R11295 gnd.n854 gnd.n838 9.3005
R11296 gnd.n5889 gnd.n855 9.3005
R11297 gnd.n5888 gnd.n856 9.3005
R11298 gnd.n5887 gnd.n857 9.3005
R11299 gnd.n3959 gnd.n3958 9.3005
R11300 gnd.n5935 gnd.n741 9.3005
R11301 gnd.n5970 gnd.n5969 9.3005
R11302 gnd.n5973 gnd.n729 9.3005
R11303 gnd.n728 gnd.n724 9.3005
R11304 gnd.n5979 gnd.n723 9.3005
R11305 gnd.n5980 gnd.n722 9.3005
R11306 gnd.n5981 gnd.n721 9.3005
R11307 gnd.n720 gnd.n716 9.3005
R11308 gnd.n5987 gnd.n715 9.3005
R11309 gnd.n5988 gnd.n714 9.3005
R11310 gnd.n5989 gnd.n713 9.3005
R11311 gnd.n712 gnd.n708 9.3005
R11312 gnd.n5995 gnd.n707 9.3005
R11313 gnd.n5996 gnd.n706 9.3005
R11314 gnd.n5997 gnd.n705 9.3005
R11315 gnd.n704 gnd.n700 9.3005
R11316 gnd.n6003 gnd.n699 9.3005
R11317 gnd.n6004 gnd.n698 9.3005
R11318 gnd.n6005 gnd.n697 9.3005
R11319 gnd.n696 gnd.n692 9.3005
R11320 gnd.n6011 gnd.n691 9.3005
R11321 gnd.n6012 gnd.n690 9.3005
R11322 gnd.n6013 gnd.n689 9.3005
R11323 gnd.n688 gnd.n684 9.3005
R11324 gnd.n6019 gnd.n683 9.3005
R11325 gnd.n6020 gnd.n682 9.3005
R11326 gnd.n6021 gnd.n681 9.3005
R11327 gnd.n680 gnd.n676 9.3005
R11328 gnd.n6027 gnd.n675 9.3005
R11329 gnd.n6028 gnd.n674 9.3005
R11330 gnd.n6029 gnd.n673 9.3005
R11331 gnd.n672 gnd.n668 9.3005
R11332 gnd.n6035 gnd.n667 9.3005
R11333 gnd.n6036 gnd.n666 9.3005
R11334 gnd.n6037 gnd.n665 9.3005
R11335 gnd.n664 gnd.n660 9.3005
R11336 gnd.n6043 gnd.n659 9.3005
R11337 gnd.n6044 gnd.n658 9.3005
R11338 gnd.n6045 gnd.n657 9.3005
R11339 gnd.n656 gnd.n652 9.3005
R11340 gnd.n6051 gnd.n651 9.3005
R11341 gnd.n6052 gnd.n650 9.3005
R11342 gnd.n6053 gnd.n649 9.3005
R11343 gnd.n648 gnd.n644 9.3005
R11344 gnd.n6059 gnd.n643 9.3005
R11345 gnd.n6060 gnd.n642 9.3005
R11346 gnd.n6061 gnd.n641 9.3005
R11347 gnd.n640 gnd.n636 9.3005
R11348 gnd.n6067 gnd.n635 9.3005
R11349 gnd.n6068 gnd.n634 9.3005
R11350 gnd.n6069 gnd.n633 9.3005
R11351 gnd.n632 gnd.n628 9.3005
R11352 gnd.n6075 gnd.n627 9.3005
R11353 gnd.n6076 gnd.n626 9.3005
R11354 gnd.n6077 gnd.n625 9.3005
R11355 gnd.n624 gnd.n620 9.3005
R11356 gnd.n6083 gnd.n619 9.3005
R11357 gnd.n6084 gnd.n618 9.3005
R11358 gnd.n6085 gnd.n617 9.3005
R11359 gnd.n616 gnd.n612 9.3005
R11360 gnd.n6091 gnd.n611 9.3005
R11361 gnd.n6092 gnd.n610 9.3005
R11362 gnd.n6093 gnd.n609 9.3005
R11363 gnd.n608 gnd.n604 9.3005
R11364 gnd.n6099 gnd.n603 9.3005
R11365 gnd.n6100 gnd.n602 9.3005
R11366 gnd.n6101 gnd.n601 9.3005
R11367 gnd.n600 gnd.n596 9.3005
R11368 gnd.n6107 gnd.n595 9.3005
R11369 gnd.n6108 gnd.n594 9.3005
R11370 gnd.n6109 gnd.n593 9.3005
R11371 gnd.n592 gnd.n588 9.3005
R11372 gnd.n6115 gnd.n587 9.3005
R11373 gnd.n6116 gnd.n586 9.3005
R11374 gnd.n6117 gnd.n585 9.3005
R11375 gnd.n584 gnd.n580 9.3005
R11376 gnd.n6123 gnd.n579 9.3005
R11377 gnd.n6124 gnd.n578 9.3005
R11378 gnd.n6125 gnd.n577 9.3005
R11379 gnd.n576 gnd.n572 9.3005
R11380 gnd.n6131 gnd.n571 9.3005
R11381 gnd.n6132 gnd.n570 9.3005
R11382 gnd.n6133 gnd.n569 9.3005
R11383 gnd.n568 gnd.n564 9.3005
R11384 gnd.n6139 gnd.n563 9.3005
R11385 gnd.n6141 gnd.n6140 9.3005
R11386 gnd.n5972 gnd.n5971 9.3005
R11387 gnd.n5173 gnd.n1632 9.3005
R11388 gnd.n4302 gnd.n4301 9.3005
R11389 gnd.n2073 gnd.n2072 9.3005
R11390 gnd.n4315 gnd.n4314 9.3005
R11391 gnd.n4316 gnd.n2071 9.3005
R11392 gnd.n4318 gnd.n4317 9.3005
R11393 gnd.n2059 gnd.n2058 9.3005
R11394 gnd.n4331 gnd.n4330 9.3005
R11395 gnd.n4332 gnd.n2057 9.3005
R11396 gnd.n4334 gnd.n4333 9.3005
R11397 gnd.n2045 gnd.n2044 9.3005
R11398 gnd.n4347 gnd.n4346 9.3005
R11399 gnd.n4348 gnd.n2043 9.3005
R11400 gnd.n4350 gnd.n4349 9.3005
R11401 gnd.n2031 gnd.n2030 9.3005
R11402 gnd.n4363 gnd.n4362 9.3005
R11403 gnd.n4364 gnd.n2029 9.3005
R11404 gnd.n4366 gnd.n4365 9.3005
R11405 gnd.n2016 gnd.n2015 9.3005
R11406 gnd.n4379 gnd.n4378 9.3005
R11407 gnd.n4380 gnd.n2014 9.3005
R11408 gnd.n4382 gnd.n4381 9.3005
R11409 gnd.n2003 gnd.n2002 9.3005
R11410 gnd.n4395 gnd.n4394 9.3005
R11411 gnd.n4396 gnd.n2000 9.3005
R11412 gnd.n4399 gnd.n4398 9.3005
R11413 gnd.n4397 gnd.n2001 9.3005
R11414 gnd.n1987 gnd.n1986 9.3005
R11415 gnd.n4419 gnd.n4418 9.3005
R11416 gnd.n4420 gnd.n1984 9.3005
R11417 gnd.n4423 gnd.n4422 9.3005
R11418 gnd.n4421 gnd.n1985 9.3005
R11419 gnd.n1219 gnd.n1217 9.3005
R11420 gnd.n5669 gnd.n5668 9.3005
R11421 gnd.n5667 gnd.n1218 9.3005
R11422 gnd.n5666 gnd.n5665 9.3005
R11423 gnd.n5664 gnd.n1220 9.3005
R11424 gnd.n5663 gnd.n5662 9.3005
R11425 gnd.n5661 gnd.n1224 9.3005
R11426 gnd.n5660 gnd.n5659 9.3005
R11427 gnd.n5658 gnd.n1225 9.3005
R11428 gnd.n5657 gnd.n5656 9.3005
R11429 gnd.n5655 gnd.n1229 9.3005
R11430 gnd.n5654 gnd.n5653 9.3005
R11431 gnd.n5652 gnd.n1230 9.3005
R11432 gnd.n5651 gnd.n5650 9.3005
R11433 gnd.n5649 gnd.n1234 9.3005
R11434 gnd.n5648 gnd.n5647 9.3005
R11435 gnd.n5646 gnd.n1235 9.3005
R11436 gnd.n5645 gnd.n5644 9.3005
R11437 gnd.n5643 gnd.n1239 9.3005
R11438 gnd.n5642 gnd.n5641 9.3005
R11439 gnd.n5640 gnd.n1240 9.3005
R11440 gnd.n5639 gnd.n5638 9.3005
R11441 gnd.n5637 gnd.n1244 9.3005
R11442 gnd.n5636 gnd.n5635 9.3005
R11443 gnd.n5634 gnd.n1245 9.3005
R11444 gnd.n5633 gnd.n5632 9.3005
R11445 gnd.n5631 gnd.n1249 9.3005
R11446 gnd.n5630 gnd.n5629 9.3005
R11447 gnd.n5628 gnd.n1250 9.3005
R11448 gnd.n5627 gnd.n5626 9.3005
R11449 gnd.n5625 gnd.n1254 9.3005
R11450 gnd.n5624 gnd.n5623 9.3005
R11451 gnd.n5622 gnd.n1255 9.3005
R11452 gnd.n5621 gnd.n5620 9.3005
R11453 gnd.n5619 gnd.n1259 9.3005
R11454 gnd.n5618 gnd.n5617 9.3005
R11455 gnd.n5616 gnd.n1260 9.3005
R11456 gnd.n5615 gnd.n5614 9.3005
R11457 gnd.n5613 gnd.n1264 9.3005
R11458 gnd.n5612 gnd.n5611 9.3005
R11459 gnd.n5610 gnd.n1265 9.3005
R11460 gnd.n5609 gnd.n5608 9.3005
R11461 gnd.n5607 gnd.n1269 9.3005
R11462 gnd.n5606 gnd.n5605 9.3005
R11463 gnd.n5604 gnd.n1270 9.3005
R11464 gnd.n5603 gnd.n5602 9.3005
R11465 gnd.n5601 gnd.n1274 9.3005
R11466 gnd.n5600 gnd.n5599 9.3005
R11467 gnd.n5598 gnd.n1275 9.3005
R11468 gnd.n5597 gnd.n5596 9.3005
R11469 gnd.n5595 gnd.n1279 9.3005
R11470 gnd.n5594 gnd.n5593 9.3005
R11471 gnd.n5592 gnd.n1280 9.3005
R11472 gnd.n5591 gnd.n5590 9.3005
R11473 gnd.n5589 gnd.n1284 9.3005
R11474 gnd.n5588 gnd.n5587 9.3005
R11475 gnd.n5586 gnd.n1285 9.3005
R11476 gnd.n5585 gnd.n5584 9.3005
R11477 gnd.n5583 gnd.n1289 9.3005
R11478 gnd.n5582 gnd.n5581 9.3005
R11479 gnd.n5580 gnd.n1290 9.3005
R11480 gnd.n5579 gnd.n5578 9.3005
R11481 gnd.n5577 gnd.n1294 9.3005
R11482 gnd.n5576 gnd.n5575 9.3005
R11483 gnd.n5574 gnd.n1295 9.3005
R11484 gnd.n5573 gnd.n5572 9.3005
R11485 gnd.n5571 gnd.n1299 9.3005
R11486 gnd.n5570 gnd.n5569 9.3005
R11487 gnd.n5568 gnd.n1300 9.3005
R11488 gnd.n5567 gnd.n1303 9.3005
R11489 gnd.n4300 gnd.n4299 9.3005
R11490 gnd.n5870 gnd.n871 9.3005
R11491 gnd.n2122 gnd.n2120 9.3005
R11492 gnd.n4115 gnd.n4114 9.3005
R11493 gnd.n4113 gnd.n2121 9.3005
R11494 gnd.n4112 gnd.n4111 9.3005
R11495 gnd.n2111 gnd.n2110 9.3005
R11496 gnd.n4156 gnd.n4155 9.3005
R11497 gnd.n4157 gnd.n2109 9.3005
R11498 gnd.n4159 gnd.n4158 9.3005
R11499 gnd.n2105 gnd.n2104 9.3005
R11500 gnd.n4170 gnd.n4169 9.3005
R11501 gnd.n4171 gnd.n2103 9.3005
R11502 gnd.n4173 gnd.n4172 9.3005
R11503 gnd.n2098 gnd.n2096 9.3005
R11504 gnd.n4197 gnd.n4196 9.3005
R11505 gnd.n4195 gnd.n2097 9.3005
R11506 gnd.n4194 gnd.n4193 9.3005
R11507 gnd.n4192 gnd.n2099 9.3005
R11508 gnd.n4191 gnd.n4190 9.3005
R11509 gnd.n870 gnd.n868 9.3005
R11510 gnd.n5876 gnd.n5875 9.3005
R11511 gnd.n5874 gnd.n869 9.3005
R11512 gnd.n5848 gnd.n5847 9.3005
R11513 gnd.n5846 gnd.n5845 9.3005
R11514 gnd.n913 gnd.n912 9.3005
R11515 gnd.n5840 gnd.n5839 9.3005
R11516 gnd.n5838 gnd.n5837 9.3005
R11517 gnd.n923 gnd.n922 9.3005
R11518 gnd.n5832 gnd.n5831 9.3005
R11519 gnd.n5830 gnd.n5829 9.3005
R11520 gnd.n931 gnd.n930 9.3005
R11521 gnd.n5824 gnd.n5823 9.3005
R11522 gnd.n5822 gnd.n5821 9.3005
R11523 gnd.n941 gnd.n940 9.3005
R11524 gnd.n5816 gnd.n5815 9.3005
R11525 gnd.n5814 gnd.n5813 9.3005
R11526 gnd.n949 gnd.n948 9.3005
R11527 gnd.n5808 gnd.n5807 9.3005
R11528 gnd.n5806 gnd.n963 9.3005
R11529 gnd.n5805 gnd.n872 9.3005
R11530 gnd.n909 gnd.n907 9.3005
R11531 gnd.n5872 gnd.n5871 9.3005
R11532 gnd.n962 gnd.n873 9.3005
R11533 gnd.n958 gnd.n957 9.3005
R11534 gnd.n5810 gnd.n5809 9.3005
R11535 gnd.n5812 gnd.n5811 9.3005
R11536 gnd.n945 gnd.n944 9.3005
R11537 gnd.n5818 gnd.n5817 9.3005
R11538 gnd.n5820 gnd.n5819 9.3005
R11539 gnd.n937 gnd.n936 9.3005
R11540 gnd.n5826 gnd.n5825 9.3005
R11541 gnd.n5828 gnd.n5827 9.3005
R11542 gnd.n927 gnd.n926 9.3005
R11543 gnd.n5834 gnd.n5833 9.3005
R11544 gnd.n5836 gnd.n5835 9.3005
R11545 gnd.n919 gnd.n918 9.3005
R11546 gnd.n5842 gnd.n5841 9.3005
R11547 gnd.n5844 gnd.n5843 9.3005
R11548 gnd.n908 gnd.n906 9.3005
R11549 gnd.n5850 gnd.n5849 9.3005
R11550 gnd.n5851 gnd.n901 9.3005
R11551 gnd.n5853 gnd.n5852 9.3005
R11552 gnd.n5855 gnd.n900 9.3005
R11553 gnd.n5857 gnd.n5856 9.3005
R11554 gnd.n5858 gnd.n896 9.3005
R11555 gnd.n5860 gnd.n5859 9.3005
R11556 gnd.n5861 gnd.n895 9.3005
R11557 gnd.n5863 gnd.n5862 9.3005
R11558 gnd.n5864 gnd.n894 9.3005
R11559 gnd.n4297 gnd.n4296 9.3005
R11560 gnd.n4295 gnd.n4231 9.3005
R11561 gnd.n4294 gnd.n4293 9.3005
R11562 gnd.n4292 gnd.n4233 9.3005
R11563 gnd.n4291 gnd.n4290 9.3005
R11564 gnd.n4289 gnd.n4236 9.3005
R11565 gnd.n4288 gnd.n4287 9.3005
R11566 gnd.n4286 gnd.n4237 9.3005
R11567 gnd.n4285 gnd.n4284 9.3005
R11568 gnd.n4283 gnd.n4240 9.3005
R11569 gnd.n4282 gnd.n4281 9.3005
R11570 gnd.n4280 gnd.n4241 9.3005
R11571 gnd.n4279 gnd.n4278 9.3005
R11572 gnd.n4277 gnd.n4244 9.3005
R11573 gnd.n4276 gnd.n4275 9.3005
R11574 gnd.n4274 gnd.n4245 9.3005
R11575 gnd.n4273 gnd.n4272 9.3005
R11576 gnd.n4271 gnd.n4248 9.3005
R11577 gnd.n4270 gnd.n4269 9.3005
R11578 gnd.n4268 gnd.n4249 9.3005
R11579 gnd.n4267 gnd.n4266 9.3005
R11580 gnd.n4265 gnd.n4252 9.3005
R11581 gnd.n4264 gnd.n4263 9.3005
R11582 gnd.n4262 gnd.n4253 9.3005
R11583 gnd.n4261 gnd.n4260 9.3005
R11584 gnd.n4259 gnd.n4256 9.3005
R11585 gnd.n4258 gnd.n4257 9.3005
R11586 gnd.n1981 gnd.n1980 9.3005
R11587 gnd.n4429 gnd.n4428 9.3005
R11588 gnd.n4430 gnd.n1979 9.3005
R11589 gnd.n4432 gnd.n4431 9.3005
R11590 gnd.n4532 gnd.n1978 9.3005
R11591 gnd.n4534 gnd.n4533 9.3005
R11592 gnd.n4535 gnd.n1976 9.3005
R11593 gnd.n4549 gnd.n4548 9.3005
R11594 gnd.n4547 gnd.n1977 9.3005
R11595 gnd.n4546 gnd.n4545 9.3005
R11596 gnd.n4544 gnd.n4536 9.3005
R11597 gnd.n4543 gnd.n4542 9.3005
R11598 gnd.n4541 gnd.n4540 9.3005
R11599 gnd.n1930 gnd.n1929 9.3005
R11600 gnd.n4615 gnd.n4614 9.3005
R11601 gnd.n4616 gnd.n1927 9.3005
R11602 gnd.n4652 gnd.n4651 9.3005
R11603 gnd.n4650 gnd.n1928 9.3005
R11604 gnd.n4649 gnd.n4648 9.3005
R11605 gnd.n4647 gnd.n4617 9.3005
R11606 gnd.n4646 gnd.n4645 9.3005
R11607 gnd.n4644 gnd.n4620 9.3005
R11608 gnd.n4643 gnd.n4642 9.3005
R11609 gnd.n4641 gnd.n4621 9.3005
R11610 gnd.n4640 gnd.n4639 9.3005
R11611 gnd.n4638 gnd.n4625 9.3005
R11612 gnd.n4637 gnd.n4636 9.3005
R11613 gnd.n4635 gnd.n4626 9.3005
R11614 gnd.n4634 gnd.n4633 9.3005
R11615 gnd.n4632 gnd.n4631 9.3005
R11616 gnd.n1850 gnd.n1849 9.3005
R11617 gnd.n4782 gnd.n4781 9.3005
R11618 gnd.n4783 gnd.n1847 9.3005
R11619 gnd.n4810 gnd.n4809 9.3005
R11620 gnd.n4808 gnd.n1848 9.3005
R11621 gnd.n4807 gnd.n4806 9.3005
R11622 gnd.n4805 gnd.n4784 9.3005
R11623 gnd.n4804 gnd.n4803 9.3005
R11624 gnd.n4802 gnd.n4788 9.3005
R11625 gnd.n4801 gnd.n4800 9.3005
R11626 gnd.n4799 gnd.n4789 9.3005
R11627 gnd.n4798 gnd.n4797 9.3005
R11628 gnd.n4796 gnd.n4793 9.3005
R11629 gnd.n4795 gnd.n4794 9.3005
R11630 gnd.n1748 gnd.n1747 9.3005
R11631 gnd.n5043 gnd.n5042 9.3005
R11632 gnd.n5044 gnd.n1746 9.3005
R11633 gnd.n5046 gnd.n5045 9.3005
R11634 gnd.n1735 gnd.n1734 9.3005
R11635 gnd.n5059 gnd.n5058 9.3005
R11636 gnd.n5060 gnd.n1733 9.3005
R11637 gnd.n5062 gnd.n5061 9.3005
R11638 gnd.n1723 gnd.n1722 9.3005
R11639 gnd.n5076 gnd.n5075 9.3005
R11640 gnd.n5077 gnd.n1721 9.3005
R11641 gnd.n5079 gnd.n5078 9.3005
R11642 gnd.n1710 gnd.n1709 9.3005
R11643 gnd.n5092 gnd.n5091 9.3005
R11644 gnd.n5093 gnd.n1708 9.3005
R11645 gnd.n5095 gnd.n5094 9.3005
R11646 gnd.n1697 gnd.n1696 9.3005
R11647 gnd.n5108 gnd.n5107 9.3005
R11648 gnd.n5109 gnd.n1695 9.3005
R11649 gnd.n5111 gnd.n5110 9.3005
R11650 gnd.n1682 gnd.n1681 9.3005
R11651 gnd.n5124 gnd.n5123 9.3005
R11652 gnd.n5125 gnd.n1680 9.3005
R11653 gnd.n5127 gnd.n5126 9.3005
R11654 gnd.n1671 gnd.n1670 9.3005
R11655 gnd.n5143 gnd.n5142 9.3005
R11656 gnd.n5144 gnd.n1669 9.3005
R11657 gnd.n5146 gnd.n5145 9.3005
R11658 gnd.n1311 gnd.n1310 9.3005
R11659 gnd.n5563 gnd.n5562 9.3005
R11660 gnd.n4232 gnd.n4230 9.3005
R11661 gnd.n5559 gnd.n1312 9.3005
R11662 gnd.n5558 gnd.n5557 9.3005
R11663 gnd.n5556 gnd.n1315 9.3005
R11664 gnd.n5555 gnd.n5554 9.3005
R11665 gnd.n5553 gnd.n1316 9.3005
R11666 gnd.n5552 gnd.n5551 9.3005
R11667 gnd.n5561 gnd.n5560 9.3005
R11668 gnd.n5504 gnd.n5503 9.3005
R11669 gnd.n1363 gnd.n1362 9.3005
R11670 gnd.n5510 gnd.n5509 9.3005
R11671 gnd.n5512 gnd.n5511 9.3005
R11672 gnd.n1355 gnd.n1354 9.3005
R11673 gnd.n5518 gnd.n5517 9.3005
R11674 gnd.n5520 gnd.n5519 9.3005
R11675 gnd.n1347 gnd.n1346 9.3005
R11676 gnd.n5526 gnd.n5525 9.3005
R11677 gnd.n5528 gnd.n5527 9.3005
R11678 gnd.n1339 gnd.n1338 9.3005
R11679 gnd.n5534 gnd.n5533 9.3005
R11680 gnd.n5536 gnd.n5535 9.3005
R11681 gnd.n1331 gnd.n1330 9.3005
R11682 gnd.n5542 gnd.n5541 9.3005
R11683 gnd.n5544 gnd.n5543 9.3005
R11684 gnd.n1327 gnd.n1322 9.3005
R11685 gnd.n5502 gnd.n1372 9.3005
R11686 gnd.n1633 gnd.n1371 9.3005
R11687 gnd.n5549 gnd.n1320 9.3005
R11688 gnd.n5548 gnd.n5547 9.3005
R11689 gnd.n5546 gnd.n5545 9.3005
R11690 gnd.n1326 gnd.n1325 9.3005
R11691 gnd.n5540 gnd.n5539 9.3005
R11692 gnd.n5538 gnd.n5537 9.3005
R11693 gnd.n1335 gnd.n1334 9.3005
R11694 gnd.n5532 gnd.n5531 9.3005
R11695 gnd.n5530 gnd.n5529 9.3005
R11696 gnd.n1343 gnd.n1342 9.3005
R11697 gnd.n5524 gnd.n5523 9.3005
R11698 gnd.n5522 gnd.n5521 9.3005
R11699 gnd.n1351 gnd.n1350 9.3005
R11700 gnd.n5516 gnd.n5515 9.3005
R11701 gnd.n5514 gnd.n5513 9.3005
R11702 gnd.n1359 gnd.n1358 9.3005
R11703 gnd.n5508 gnd.n5507 9.3005
R11704 gnd.n5506 gnd.n5505 9.3005
R11705 gnd.n1656 gnd.n1369 9.3005
R11706 gnd.n1635 gnd.n1634 9.3005
R11707 gnd.n5175 gnd.n5174 9.3005
R11708 gnd.n5216 gnd.n5215 9.3005
R11709 gnd.n5214 gnd.n1631 9.3005
R11710 gnd.n5213 gnd.n5212 9.3005
R11711 gnd.n5211 gnd.n5178 9.3005
R11712 gnd.n5210 gnd.n5209 9.3005
R11713 gnd.n5208 gnd.n5182 9.3005
R11714 gnd.n5207 gnd.n5206 9.3005
R11715 gnd.n5205 gnd.n5183 9.3005
R11716 gnd.n5204 gnd.n5203 9.3005
R11717 gnd.n1614 gnd.n1613 9.3005
R11718 gnd.n5264 gnd.n5263 9.3005
R11719 gnd.n5265 gnd.n1612 9.3005
R11720 gnd.n5267 gnd.n5266 9.3005
R11721 gnd.n1609 gnd.n1608 9.3005
R11722 gnd.n5279 gnd.n5278 9.3005
R11723 gnd.n5280 gnd.n1606 9.3005
R11724 gnd.n5286 gnd.n5285 9.3005
R11725 gnd.n5284 gnd.n1607 9.3005
R11726 gnd.n5283 gnd.n5282 9.3005
R11727 gnd.n5281 gnd.n67 9.3005
R11728 gnd.n5177 gnd.n1630 9.3005
R11729 gnd.n7208 gnd.n68 9.3005
R11730 gnd.t123 gnd.n2395 9.24152
R11731 gnd.n2297 gnd.t27 9.24152
R11732 gnd.n3565 gnd.t111 9.24152
R11733 gnd.n2106 gnd.t264 9.24152
R11734 gnd.n5032 gnd.t151 9.24152
R11735 gnd.n5260 gnd.t227 9.24152
R11736 gnd.t177 gnd.t123 8.92286
R11737 gnd.n4602 gnd.t146 8.92286
R11738 gnd.n4595 gnd.t162 8.92286
R11739 gnd.n4761 gnd.t150 8.92286
R11740 gnd.t163 gnd.n4812 8.92286
R11741 gnd.n3535 gnd.n3510 8.92171
R11742 gnd.n3503 gnd.n3478 8.92171
R11743 gnd.n3471 gnd.n3446 8.92171
R11744 gnd.n3440 gnd.n3415 8.92171
R11745 gnd.n3408 gnd.n3383 8.92171
R11746 gnd.n3376 gnd.n3351 8.92171
R11747 gnd.n3344 gnd.n3319 8.92171
R11748 gnd.n3313 gnd.n3288 8.92171
R11749 gnd.n4888 gnd.n4870 8.72777
R11750 gnd.n3039 gnd.t132 8.60421
R11751 gnd.n4118 gnd.t213 8.60421
R11752 gnd.t323 gnd.n1904 8.60421
R11753 gnd.n4714 gnd.t126 8.60421
R11754 gnd.n5314 gnd.t243 8.60421
R11755 gnd.n2459 gnd.n2447 8.43656
R11756 gnd.n42 gnd.n30 8.43656
R11757 gnd.n4567 gnd.n1960 8.28555
R11758 gnd.n4581 gnd.n1910 8.28555
R11759 gnd.n4731 gnd.n1876 8.28555
R11760 gnd.n4750 gnd.n1829 8.28555
R11761 gnd.n3536 gnd.n3508 8.14595
R11762 gnd.n3504 gnd.n3476 8.14595
R11763 gnd.n3472 gnd.n3444 8.14595
R11764 gnd.n3441 gnd.n3413 8.14595
R11765 gnd.n3409 gnd.n3381 8.14595
R11766 gnd.n3377 gnd.n3349 8.14595
R11767 gnd.n3345 gnd.n3317 8.14595
R11768 gnd.n3314 gnd.n3286 8.14595
R11769 gnd.n4095 gnd.n0 8.10675
R11770 gnd.n7209 gnd.n7208 8.10675
R11771 gnd.n3541 gnd.n3540 7.97301
R11772 gnd.t156 gnd.n2554 7.9669
R11773 gnd.n5867 gnd.n876 7.9669
R11774 gnd.n5170 gnd.n5169 7.9669
R11775 gnd.n7209 gnd.n66 7.78567
R11776 gnd.n5502 gnd.n1371 7.75808
R11777 gnd.n5806 gnd.n5805 7.75808
R11778 gnd.n7089 gnd.n6814 7.75808
R11779 gnd.n3736 gnd.n3674 7.75808
R11780 gnd.t166 gnd.n726 7.64824
R11781 gnd.n1824 gnd.t60 7.64824
R11782 gnd.n2484 gnd.n2483 7.53171
R11783 gnd.n2948 gnd.t187 7.32958
R11784 gnd.t46 gnd.n2075 7.32958
R11785 gnd.n4344 gnd.t321 7.32958
R11786 gnd.t192 gnd.n1693 7.32958
R11787 gnd.n5148 gnd.t31 7.32958
R11788 gnd.n7147 gnd.n170 7.32958
R11789 gnd.n1197 gnd.n1196 7.30353
R11790 gnd.n4887 gnd.n4886 7.30353
R11791 gnd.n2908 gnd.n2627 7.01093
R11792 gnd.n2630 gnd.n2628 7.01093
R11793 gnd.n2918 gnd.n2917 7.01093
R11794 gnd.n2929 gnd.n2611 7.01093
R11795 gnd.n2928 gnd.n2614 7.01093
R11796 gnd.n2939 gnd.n2602 7.01093
R11797 gnd.n2605 gnd.n2603 7.01093
R11798 gnd.n2949 gnd.n2948 7.01093
R11799 gnd.n2959 gnd.n2583 7.01093
R11800 gnd.n2958 gnd.n2586 7.01093
R11801 gnd.n2967 gnd.n2577 7.01093
R11802 gnd.n2979 gnd.n2567 7.01093
R11803 gnd.n2989 gnd.n2552 7.01093
R11804 gnd.n3005 gnd.n3004 7.01093
R11805 gnd.n2554 gnd.n2491 7.01093
R11806 gnd.n3059 gnd.n2492 7.01093
R11807 gnd.n3053 gnd.n3052 7.01093
R11808 gnd.n2541 gnd.n2503 7.01093
R11809 gnd.n3045 gnd.n2514 7.01093
R11810 gnd.n2532 gnd.n2527 7.01093
R11811 gnd.n3039 gnd.n3038 7.01093
R11812 gnd.n3085 gnd.n2430 7.01093
R11813 gnd.n3084 gnd.n3083 7.01093
R11814 gnd.n3096 gnd.n3095 7.01093
R11815 gnd.n2423 gnd.n2415 7.01093
R11816 gnd.n3125 gnd.n2403 7.01093
R11817 gnd.n3124 gnd.n2406 7.01093
R11818 gnd.n3135 gnd.n2395 7.01093
R11819 gnd.n2396 gnd.n2384 7.01093
R11820 gnd.n3146 gnd.n2385 7.01093
R11821 gnd.n3170 gnd.n2376 7.01093
R11822 gnd.n3169 gnd.n2367 7.01093
R11823 gnd.n3192 gnd.n3191 7.01093
R11824 gnd.n3210 gnd.n2348 7.01093
R11825 gnd.n3209 gnd.n2351 7.01093
R11826 gnd.n3220 gnd.n2340 7.01093
R11827 gnd.n2341 gnd.n2328 7.01093
R11828 gnd.n3231 gnd.n2329 7.01093
R11829 gnd.n3258 gnd.n2313 7.01093
R11830 gnd.n3270 gnd.n3269 7.01093
R11831 gnd.n3252 gnd.n2306 7.01093
R11832 gnd.n3281 gnd.n3280 7.01093
R11833 gnd.n3553 gnd.n2294 7.01093
R11834 gnd.n3552 gnd.n2297 7.01093
R11835 gnd.n3565 gnd.n2286 7.01093
R11836 gnd.n2287 gnd.n2279 7.01093
R11837 gnd.n3575 gnd.n2205 7.01093
R11838 gnd.n5678 gnd.n5677 7.01093
R11839 gnd.n4559 gnd.n4558 7.01093
R11840 gnd.n4558 gnd.t108 7.01093
R11841 gnd.n4688 gnd.n1905 7.01093
R11842 gnd.n4723 gnd.n4722 7.01093
R11843 gnd.n4838 gnd.n1825 7.01093
R11844 gnd.n4961 gnd.n1797 7.01093
R11845 gnd.t99 gnd.n1755 7.01093
R11846 gnd.n2586 gnd.t122 6.69227
R11847 gnd.n2406 gnd.t177 6.69227
R11848 gnd.n2329 gnd.n726 6.69227
R11849 gnd.n3259 gnd.t318 6.69227
R11850 gnd.n5023 gnd.n5022 6.5566
R11851 gnd.n4442 gnd.n4441 6.5566
R11852 gnd.n5689 gnd.n5685 6.5566
R11853 gnd.n4898 gnd.n4897 6.5566
R11854 gnd.n4425 gnd.t102 6.37362
R11855 gnd.n4661 gnd.t147 6.37362
R11856 gnd.n4738 gnd.t130 6.37362
R11857 gnd.n957 gnd.n955 6.20656
R11858 gnd.n1656 gnd.n1368 6.20656
R11859 gnd.t148 gnd.n3015 6.05496
R11860 gnd.n3016 gnd.t140 6.05496
R11861 gnd.t181 gnd.n2430 6.05496
R11862 gnd.t185 gnd.n3180 6.05496
R11863 gnd.n5748 gnd.n1175 6.05496
R11864 gnd.n1905 gnd.t323 6.05496
R11865 gnd.n4723 gnd.t126 6.05496
R11866 gnd.n5031 gnd.n5030 6.05496
R11867 gnd.n3538 gnd.n3508 5.81868
R11868 gnd.n3506 gnd.n3476 5.81868
R11869 gnd.n3474 gnd.n3444 5.81868
R11870 gnd.n3443 gnd.n3413 5.81868
R11871 gnd.n3411 gnd.n3381 5.81868
R11872 gnd.n3379 gnd.n3349 5.81868
R11873 gnd.n3347 gnd.n3317 5.81868
R11874 gnd.n3316 gnd.n3286 5.81868
R11875 gnd.n5671 gnd.n1213 5.73631
R11876 gnd.n4522 gnd.n4521 5.73631
R11877 gnd.n4695 gnd.n1894 5.73631
R11878 gnd.n1895 gnd.n1888 5.73631
R11879 gnd.n4857 gnd.n1811 5.73631
R11880 gnd.n4790 gnd.n1802 5.73631
R11881 gnd.n5027 gnd.n1448 5.62001
R11882 gnd.n5751 gnd.n1139 5.62001
R11883 gnd.n5751 gnd.n1140 5.62001
R11884 gnd.n4893 gnd.n1448 5.62001
R11885 gnd.n2767 gnd.n2762 5.4308
R11886 gnd.n3583 gnd.n2272 5.4308
R11887 gnd.n3083 gnd.t168 5.41765
R11888 gnd.t176 gnd.n3106 5.41765
R11889 gnd.t153 gnd.n2360 5.41765
R11890 gnd.n3536 gnd.n3535 5.04292
R11891 gnd.n3504 gnd.n3503 5.04292
R11892 gnd.n3472 gnd.n3471 5.04292
R11893 gnd.n3441 gnd.n3440 5.04292
R11894 gnd.n3409 gnd.n3408 5.04292
R11895 gnd.n3377 gnd.n3376 5.04292
R11896 gnd.n3345 gnd.n3344 5.04292
R11897 gnd.n3314 gnd.n3313 5.04292
R11898 gnd.n3046 gnd.t175 4.78034
R11899 gnd.n2385 gnd.t131 4.78034
R11900 gnd.t164 gnd.n2026 4.78034
R11901 gnd.n4521 gnd.t316 4.78034
R11902 gnd.t188 gnd.n1811 4.78034
R11903 gnd.n5030 gnd.t43 4.78034
R11904 gnd.n5089 gnd.t325 4.78034
R11905 gnd.n2488 gnd.n2485 4.74817
R11906 gnd.n2538 gnd.n2436 4.74817
R11907 gnd.n2525 gnd.n2435 4.74817
R11908 gnd.n2434 gnd.n2433 4.74817
R11909 gnd.n2534 gnd.n2485 4.74817
R11910 gnd.n2535 gnd.n2436 4.74817
R11911 gnd.n2537 gnd.n2435 4.74817
R11912 gnd.n2524 gnd.n2434 4.74817
R11913 gnd.n5317 gnd.n86 4.74817
R11914 gnd.n1584 gnd.n85 4.74817
R11915 gnd.n1594 gnd.n84 4.74817
R11916 gnd.n7201 gnd.n79 4.74817
R11917 gnd.n7199 gnd.n80 4.74817
R11918 gnd.n5328 gnd.n86 4.74817
R11919 gnd.n5318 gnd.n85 4.74817
R11920 gnd.n1583 gnd.n84 4.74817
R11921 gnd.n1593 gnd.n79 4.74817
R11922 gnd.n7200 gnd.n7199 4.74817
R11923 gnd.n4080 gnd.n731 4.74817
R11924 gnd.n4087 gnd.n4084 4.74817
R11925 gnd.n4085 gnd.n2117 4.74817
R11926 gnd.n4122 gnd.n4121 4.74817
R11927 gnd.n4126 gnd.n2115 4.74817
R11928 gnd.n5250 gnd.n5249 4.74817
R11929 gnd.n5312 gnd.n1589 4.74817
R11930 gnd.n5310 gnd.n5309 4.74817
R11931 gnd.n1590 gnd.n183 4.74817
R11932 gnd.n6780 gnd.n6779 4.74817
R11933 gnd.n5251 gnd.n5250 4.74817
R11934 gnd.n5247 gnd.n1589 4.74817
R11935 gnd.n5311 gnd.n5310 4.74817
R11936 gnd.n1591 gnd.n1590 4.74817
R11937 gnd.n6781 gnd.n6780 4.74817
R11938 gnd.n5963 gnd.n5962 4.74817
R11939 gnd.n760 gnd.n742 4.74817
R11940 gnd.n5950 gnd.n5949 4.74817
R11941 gnd.n777 gnd.n761 4.74817
R11942 gnd.n5937 gnd.n5936 4.74817
R11943 gnd.n5964 gnd.n5963 4.74817
R11944 gnd.n5961 gnd.n742 4.74817
R11945 gnd.n5951 gnd.n5950 4.74817
R11946 gnd.n5948 gnd.n761 4.74817
R11947 gnd.n5938 gnd.n5937 4.74817
R11948 gnd.n4082 gnd.n4080 4.74817
R11949 gnd.n4084 gnd.n4083 4.74817
R11950 gnd.n4086 gnd.n4085 4.74817
R11951 gnd.n4121 gnd.n4120 4.74817
R11952 gnd.n4123 gnd.n2115 4.74817
R11953 gnd.n2483 gnd.n2482 4.74296
R11954 gnd.n66 gnd.n65 4.74296
R11955 gnd.n2459 gnd.n2458 4.7074
R11956 gnd.n2471 gnd.n2470 4.7074
R11957 gnd.n42 gnd.n41 4.7074
R11958 gnd.n54 gnd.n53 4.7074
R11959 gnd.n2483 gnd.n2471 4.65959
R11960 gnd.n66 gnd.n54 4.65959
R11961 gnd.n5444 gnd.n1450 4.6132
R11962 gnd.n5752 gnd.n1138 4.6132
R11963 gnd.n4530 gnd.n4529 4.46168
R11964 gnd.n4552 gnd.n4551 4.46168
R11965 gnd.n4696 gnd.n1899 4.46168
R11966 gnd.n4716 gnd.n4715 4.46168
R11967 gnd.n4850 gnd.n1818 4.46168
R11968 gnd.t3 gnd.n4856 4.46168
R11969 gnd.n4866 gnd.n4865 4.46168
R11970 gnd.n4883 gnd.n4870 4.46111
R11971 gnd.n3521 gnd.n3517 4.38594
R11972 gnd.n3489 gnd.n3485 4.38594
R11973 gnd.n3457 gnd.n3453 4.38594
R11974 gnd.n3426 gnd.n3422 4.38594
R11975 gnd.n3394 gnd.n3390 4.38594
R11976 gnd.n3362 gnd.n3358 4.38594
R11977 gnd.n3330 gnd.n3326 4.38594
R11978 gnd.n3299 gnd.n3295 4.38594
R11979 gnd.n3532 gnd.n3510 4.26717
R11980 gnd.n3500 gnd.n3478 4.26717
R11981 gnd.n3468 gnd.n3446 4.26717
R11982 gnd.n3437 gnd.n3415 4.26717
R11983 gnd.n3405 gnd.n3383 4.26717
R11984 gnd.n3373 gnd.n3351 4.26717
R11985 gnd.n3341 gnd.n3319 4.26717
R11986 gnd.n3310 gnd.n3288 4.26717
R11987 gnd.n2990 gnd.t139 4.14303
R11988 gnd.n3220 gnd.t121 4.14303
R11989 gnd.n867 gnd.t39 4.14303
R11990 gnd.n5219 gnd.t23 4.14303
R11991 gnd.n3540 gnd.n3539 4.08274
R11992 gnd.n5022 gnd.n5021 4.05904
R11993 gnd.n4443 gnd.n4442 4.05904
R11994 gnd.n5692 gnd.n5685 4.05904
R11995 gnd.n4899 gnd.n4898 4.05904
R11996 gnd.n19 gnd.n9 3.99943
R11997 gnd.n5671 gnd.t6 3.82437
R11998 gnd.n1904 gnd.t124 3.82437
R11999 gnd.t129 gnd.n4714 3.82437
R12000 gnd.n4790 gnd.t10 3.82437
R12001 gnd.n3063 gnd.n2484 3.81325
R12002 gnd.n2471 gnd.n2459 3.72967
R12003 gnd.n54 gnd.n42 3.72967
R12004 gnd.n3540 gnd.n3412 3.70378
R12005 gnd.n19 gnd.n18 3.60163
R12006 gnd.n3531 gnd.n3512 3.49141
R12007 gnd.n3499 gnd.n3480 3.49141
R12008 gnd.n3467 gnd.n3448 3.49141
R12009 gnd.n3436 gnd.n3417 3.49141
R12010 gnd.n3404 gnd.n3385 3.49141
R12011 gnd.n3372 gnd.n3353 3.49141
R12012 gnd.n3340 gnd.n3321 3.49141
R12013 gnd.n3309 gnd.n3290 3.49141
R12014 gnd.n5462 gnd.n5461 3.29747
R12015 gnd.n5461 gnd.n5460 3.29747
R12016 gnd.n7053 gnd.n7050 3.29747
R12017 gnd.n7054 gnd.n7053 3.29747
R12018 gnd.n3774 gnd.n3770 3.29747
R12019 gnd.n3920 gnd.n3774 3.29747
R12020 gnd.n5770 gnd.n5769 3.29747
R12021 gnd.n5769 gnd.n5768 3.29747
R12022 gnd.n4425 gnd.n1201 3.18706
R12023 gnd.n4655 gnd.t157 3.18706
R12024 gnd.n4681 gnd.n1903 3.18706
R12025 gnd.n4628 gnd.n1884 3.18706
R12026 gnd.n4768 gnd.t138 3.18706
R12027 gnd.n5032 gnd.n1755 3.18706
R12028 gnd.n2569 gnd.t139 2.8684
R12029 gnd.n4401 gnd.t0 2.8684
R12030 gnd.t102 gnd.t160 2.8684
R12031 gnd.t179 gnd.n1737 2.8684
R12032 gnd.n2472 gnd.t274 2.82907
R12033 gnd.n2472 gnd.t315 2.82907
R12034 gnd.n2474 gnd.t241 2.82907
R12035 gnd.n2474 gnd.t307 2.82907
R12036 gnd.n2476 gnd.t208 2.82907
R12037 gnd.n2476 gnd.t293 2.82907
R12038 gnd.n2478 gnd.t310 2.82907
R12039 gnd.n2478 gnd.t238 2.82907
R12040 gnd.n2480 gnd.t262 2.82907
R12041 gnd.n2480 gnd.t247 2.82907
R12042 gnd.n2437 gnd.t279 2.82907
R12043 gnd.n2437 gnd.t291 2.82907
R12044 gnd.n2439 gnd.t299 2.82907
R12045 gnd.n2439 gnd.t311 2.82907
R12046 gnd.n2441 gnd.t271 2.82907
R12047 gnd.n2441 gnd.t283 2.82907
R12048 gnd.n2443 gnd.t292 2.82907
R12049 gnd.n2443 gnd.t222 2.82907
R12050 gnd.n2445 gnd.t282 2.82907
R12051 gnd.n2445 gnd.t278 2.82907
R12052 gnd.n2448 gnd.t265 2.82907
R12053 gnd.n2448 gnd.t254 2.82907
R12054 gnd.n2450 gnd.t255 2.82907
R12055 gnd.n2450 gnd.t277 2.82907
R12056 gnd.n2452 gnd.t235 2.82907
R12057 gnd.n2452 gnd.t263 2.82907
R12058 gnd.n2454 gnd.t266 2.82907
R12059 gnd.n2454 gnd.t249 2.82907
R12060 gnd.n2456 gnd.t199 2.82907
R12061 gnd.n2456 gnd.t237 2.82907
R12062 gnd.n2460 gnd.t303 2.82907
R12063 gnd.n2460 gnd.t269 2.82907
R12064 gnd.n2462 gnd.t287 2.82907
R12065 gnd.n2462 gnd.t201 2.82907
R12066 gnd.n2464 gnd.t273 2.82907
R12067 gnd.n2464 gnd.t214 2.82907
R12068 gnd.n2466 gnd.t252 2.82907
R12069 gnd.n2466 gnd.t285 2.82907
R12070 gnd.n2468 gnd.t297 2.82907
R12071 gnd.n2468 gnd.t289 2.82907
R12072 gnd.n63 gnd.t314 2.82907
R12073 gnd.n63 gnd.t234 2.82907
R12074 gnd.n61 gnd.t312 2.82907
R12075 gnd.n61 gnd.t288 2.82907
R12076 gnd.n59 gnd.t272 2.82907
R12077 gnd.n59 gnd.t305 2.82907
R12078 gnd.n57 gnd.t286 2.82907
R12079 gnd.n57 gnd.t313 2.82907
R12080 gnd.n55 gnd.t296 2.82907
R12081 gnd.n55 gnd.t228 2.82907
R12082 gnd.n28 gnd.t294 2.82907
R12083 gnd.n28 gnd.t275 2.82907
R12084 gnd.n26 gnd.t259 2.82907
R12085 gnd.n26 gnd.t309 2.82907
R12086 gnd.n24 gnd.t302 2.82907
R12087 gnd.n24 gnd.t250 2.82907
R12088 gnd.n22 gnd.t233 2.82907
R12089 gnd.n22 gnd.t197 2.82907
R12090 gnd.n20 gnd.t308 2.82907
R12091 gnd.n20 gnd.t295 2.82907
R12092 gnd.n39 gnd.t216 2.82907
R12093 gnd.n39 gnd.t224 2.82907
R12094 gnd.n37 gnd.t226 2.82907
R12095 gnd.n37 gnd.t242 2.82907
R12096 gnd.n35 gnd.t244 2.82907
R12097 gnd.n35 gnd.t258 2.82907
R12098 gnd.n33 gnd.t256 2.82907
R12099 gnd.n33 gnd.t231 2.82907
R12100 gnd.n31 gnd.t232 2.82907
R12101 gnd.n31 gnd.t239 2.82907
R12102 gnd.n51 gnd.t267 2.82907
R12103 gnd.n51 gnd.t284 2.82907
R12104 gnd.n49 gnd.t260 2.82907
R12105 gnd.n49 gnd.t210 2.82907
R12106 gnd.n47 gnd.t301 2.82907
R12107 gnd.n47 gnd.t246 2.82907
R12108 gnd.n45 gnd.t206 2.82907
R12109 gnd.n45 gnd.t261 2.82907
R12110 gnd.n43 gnd.t220 2.82907
R12111 gnd.n43 gnd.t280 2.82907
R12112 gnd.n3528 gnd.n3527 2.71565
R12113 gnd.n3496 gnd.n3495 2.71565
R12114 gnd.n3464 gnd.n3463 2.71565
R12115 gnd.n3433 gnd.n3432 2.71565
R12116 gnd.n3401 gnd.n3400 2.71565
R12117 gnd.n3369 gnd.n3368 2.71565
R12118 gnd.n3337 gnd.n3336 2.71565
R12119 gnd.n3306 gnd.n3305 2.71565
R12120 gnd.n4552 gnd.t63 2.54975
R12121 gnd.t135 gnd.n4681 2.54975
R12122 gnd.n4628 gnd.t128 2.54975
R12123 gnd.n3063 gnd.n2485 2.27742
R12124 gnd.n3063 gnd.n2436 2.27742
R12125 gnd.n3063 gnd.n2435 2.27742
R12126 gnd.n3063 gnd.n2434 2.27742
R12127 gnd.n7198 gnd.n86 2.27742
R12128 gnd.n7198 gnd.n85 2.27742
R12129 gnd.n7198 gnd.n84 2.27742
R12130 gnd.n7198 gnd.n79 2.27742
R12131 gnd.n7199 gnd.n7198 2.27742
R12132 gnd.n5250 gnd.n83 2.27742
R12133 gnd.n1589 gnd.n83 2.27742
R12134 gnd.n5310 gnd.n83 2.27742
R12135 gnd.n1590 gnd.n83 2.27742
R12136 gnd.n6780 gnd.n83 2.27742
R12137 gnd.n5963 gnd.n741 2.27742
R12138 gnd.n742 gnd.n741 2.27742
R12139 gnd.n5950 gnd.n741 2.27742
R12140 gnd.n761 gnd.n741 2.27742
R12141 gnd.n5937 gnd.n741 2.27742
R12142 gnd.n4080 gnd.n730 2.27742
R12143 gnd.n4084 gnd.n730 2.27742
R12144 gnd.n4085 gnd.n730 2.27742
R12145 gnd.n4121 gnd.n730 2.27742
R12146 gnd.n2115 gnd.n730 2.27742
R12147 gnd.n2917 gnd.t53 2.23109
R12148 gnd.n2540 gnd.t175 2.23109
R12149 gnd.n4089 gnd.t207 2.23109
R12150 gnd.t245 gnd.n73 2.23109
R12151 gnd.n3524 gnd.n3514 1.93989
R12152 gnd.n3492 gnd.n3482 1.93989
R12153 gnd.n3460 gnd.n3450 1.93989
R12154 gnd.n3429 gnd.n3419 1.93989
R12155 gnd.n3397 gnd.n3387 1.93989
R12156 gnd.n3365 gnd.n3355 1.93989
R12157 gnd.n3333 gnd.n3323 1.93989
R12158 gnd.n3302 gnd.n3292 1.93989
R12159 gnd.n4512 gnd.t143 1.91244
R12160 gnd.n4612 gnd.t162 1.91244
R12161 gnd.n4662 gnd.n4661 1.91244
R12162 gnd.n4738 gnd.n1870 1.91244
R12163 gnd.n4779 gnd.t150 1.91244
R12164 gnd.t145 gnd.n1823 1.91244
R12165 gnd.t158 gnd.n2928 1.59378
R12166 gnd.n3107 gnd.t176 1.59378
R12167 gnd.n2369 gnd.t153 1.59378
R12168 gnd.n4152 gnd.t200 1.59378
R12169 gnd.n4538 gnd.t173 1.59378
R12170 gnd.n4821 gnd.t183 1.59378
R12171 gnd.n1610 gnd.t205 1.59378
R12172 gnd.t143 gnd.n1957 1.27512
R12173 gnd.n4831 gnd.t145 1.27512
R12174 gnd.n2770 gnd.n2762 1.16414
R12175 gnd.n3586 gnd.n2272 1.16414
R12176 gnd.n3523 gnd.n3516 1.16414
R12177 gnd.n3491 gnd.n3484 1.16414
R12178 gnd.n3459 gnd.n3452 1.16414
R12179 gnd.n3428 gnd.n3421 1.16414
R12180 gnd.n3396 gnd.n3389 1.16414
R12181 gnd.n3364 gnd.n3357 1.16414
R12182 gnd.n3332 gnd.n3325 1.16414
R12183 gnd.n3301 gnd.n3294 1.16414
R12184 gnd.n5444 gnd.n5443 0.970197
R12185 gnd.n5752 gnd.n1040 0.970197
R12186 gnd.n3507 gnd.n3475 0.962709
R12187 gnd.n3539 gnd.n3507 0.962709
R12188 gnd.n3380 gnd.n3348 0.962709
R12189 gnd.n3412 gnd.n3380 0.962709
R12190 gnd.n3016 gnd.t148 0.956468
R12191 gnd.n3181 gnd.t185 0.956468
R12192 gnd.n4024 gnd.t198 0.956468
R12193 gnd.n4175 gnd.t253 0.956468
R12194 gnd.n4200 gnd.t211 0.956468
R12195 gnd.t136 gnd.t157 0.956468
R12196 gnd.t141 gnd.t138 0.956468
R12197 gnd.n5191 gnd.t217 0.956468
R12198 gnd.n5201 gnd.t219 0.956468
R12199 gnd.n130 gnd.t223 0.956468
R12200 gnd.n2 gnd.n1 0.672012
R12201 gnd.n3 gnd.n2 0.672012
R12202 gnd.n4 gnd.n3 0.672012
R12203 gnd.n5 gnd.n4 0.672012
R12204 gnd.n6 gnd.n5 0.672012
R12205 gnd.n7 gnd.n6 0.672012
R12206 gnd.n8 gnd.n7 0.672012
R12207 gnd.n9 gnd.n8 0.672012
R12208 gnd.n11 gnd.n10 0.672012
R12209 gnd.n12 gnd.n11 0.672012
R12210 gnd.n13 gnd.n12 0.672012
R12211 gnd.n14 gnd.n13 0.672012
R12212 gnd.n15 gnd.n14 0.672012
R12213 gnd.n16 gnd.n15 0.672012
R12214 gnd.n17 gnd.n16 0.672012
R12215 gnd.n18 gnd.n17 0.672012
R12216 gnd.t146 gnd.n4601 0.637812
R12217 gnd.n1949 gnd.n1943 0.637812
R12218 gnd.n4589 gnd.n4588 0.637812
R12219 gnd.n4745 gnd.n4744 0.637812
R12220 gnd.n4760 gnd.n1844 0.637812
R12221 gnd.n4813 gnd.t163 0.637812
R12222 gnd.n4865 gnd.t81 0.637812
R12223 gnd gnd.n0 0.624033
R12224 gnd.n2482 gnd.n2481 0.573776
R12225 gnd.n2481 gnd.n2479 0.573776
R12226 gnd.n2479 gnd.n2477 0.573776
R12227 gnd.n2477 gnd.n2475 0.573776
R12228 gnd.n2475 gnd.n2473 0.573776
R12229 gnd.n2447 gnd.n2446 0.573776
R12230 gnd.n2446 gnd.n2444 0.573776
R12231 gnd.n2444 gnd.n2442 0.573776
R12232 gnd.n2442 gnd.n2440 0.573776
R12233 gnd.n2440 gnd.n2438 0.573776
R12234 gnd.n2458 gnd.n2457 0.573776
R12235 gnd.n2457 gnd.n2455 0.573776
R12236 gnd.n2455 gnd.n2453 0.573776
R12237 gnd.n2453 gnd.n2451 0.573776
R12238 gnd.n2451 gnd.n2449 0.573776
R12239 gnd.n2470 gnd.n2469 0.573776
R12240 gnd.n2469 gnd.n2467 0.573776
R12241 gnd.n2467 gnd.n2465 0.573776
R12242 gnd.n2465 gnd.n2463 0.573776
R12243 gnd.n2463 gnd.n2461 0.573776
R12244 gnd.n58 gnd.n56 0.573776
R12245 gnd.n60 gnd.n58 0.573776
R12246 gnd.n62 gnd.n60 0.573776
R12247 gnd.n64 gnd.n62 0.573776
R12248 gnd.n65 gnd.n64 0.573776
R12249 gnd.n23 gnd.n21 0.573776
R12250 gnd.n25 gnd.n23 0.573776
R12251 gnd.n27 gnd.n25 0.573776
R12252 gnd.n29 gnd.n27 0.573776
R12253 gnd.n30 gnd.n29 0.573776
R12254 gnd.n34 gnd.n32 0.573776
R12255 gnd.n36 gnd.n34 0.573776
R12256 gnd.n38 gnd.n36 0.573776
R12257 gnd.n40 gnd.n38 0.573776
R12258 gnd.n41 gnd.n40 0.573776
R12259 gnd.n46 gnd.n44 0.573776
R12260 gnd.n48 gnd.n46 0.573776
R12261 gnd.n50 gnd.n48 0.573776
R12262 gnd.n52 gnd.n50 0.573776
R12263 gnd.n53 gnd.n52 0.573776
R12264 gnd.n7091 gnd.n7090 0.532512
R12265 gnd.n3738 gnd.n3737 0.532512
R12266 gnd.n6906 gnd.n165 0.497451
R12267 gnd.n1012 gnd.n857 0.497451
R12268 gnd.n1501 gnd.n1420 0.497451
R12269 gnd.n3958 gnd.n3957 0.497451
R12270 gnd.n3243 gnd.n2276 0.486781
R12271 gnd.n2819 gnd.n2818 0.48678
R12272 gnd.n3560 gnd.n2230 0.480683
R12273 gnd.n2903 gnd.n2902 0.480683
R12274 gnd.n6142 gnd.n6141 0.480683
R12275 gnd.n6563 gnd.n6562 0.480683
R12276 gnd.n6774 gnd.n184 0.480683
R12277 gnd.n5971 gnd.n5970 0.480683
R12278 gnd.n7210 gnd.n7209 0.4705
R12279 gnd.n1632 gnd.n1303 0.451719
R12280 gnd.n4300 gnd.n871 0.451719
R12281 gnd.n4232 gnd.n894 0.451719
R12282 gnd.n5562 gnd.n5561 0.451719
R12283 gnd.n7198 gnd.n83 0.4255
R12284 gnd.n741 gnd.n730 0.4255
R12285 gnd.n5810 gnd.n955 0.388379
R12286 gnd.n3520 gnd.n3519 0.388379
R12287 gnd.n3488 gnd.n3487 0.388379
R12288 gnd.n3456 gnd.n3455 0.388379
R12289 gnd.n3425 gnd.n3424 0.388379
R12290 gnd.n3393 gnd.n3392 0.388379
R12291 gnd.n3361 gnd.n3360 0.388379
R12292 gnd.n3329 gnd.n3328 0.388379
R12293 gnd.n3298 gnd.n3297 0.388379
R12294 gnd.n5506 gnd.n1368 0.388379
R12295 gnd.n7210 gnd.n19 0.374463
R12296 gnd gnd.n7210 0.367492
R12297 gnd.n2331 gnd.t318 0.319156
R12298 gnd.n4072 gnd.t221 0.319156
R12299 gnd.n4109 gnd.t240 0.319156
R12300 gnd.n4574 gnd.t173 0.319156
R12301 gnd.t183 gnd.n4819 0.319156
R12302 gnd.n5288 gnd.t196 0.319156
R12303 gnd.n6791 gnd.t225 0.319156
R12304 gnd.n2737 gnd.n2715 0.311721
R12305 gnd.n5874 gnd.n5873 0.302329
R12306 gnd.n5177 gnd.n5176 0.302329
R12307 gnd.n6832 gnd.n173 0.293183
R12308 gnd.n3690 gnd.n2203 0.293183
R12309 gnd.n3631 gnd.n3630 0.268793
R12310 gnd.n6967 gnd.n173 0.258122
R12311 gnd.n5382 gnd.n1321 0.258122
R12312 gnd.n1073 gnd.n865 0.258122
R12313 gnd.n3839 gnd.n2203 0.258122
R12314 gnd.n3630 gnd.n3629 0.241354
R12315 gnd.n1450 gnd.n1447 0.229039
R12316 gnd.n1451 gnd.n1450 0.229039
R12317 gnd.n1138 gnd.n1039 0.229039
R12318 gnd.n1138 gnd.n1137 0.229039
R12319 gnd.n2891 gnd.n2690 0.206293
R12320 gnd.n3537 gnd.n3509 0.155672
R12321 gnd.n3530 gnd.n3509 0.155672
R12322 gnd.n3530 gnd.n3529 0.155672
R12323 gnd.n3529 gnd.n3513 0.155672
R12324 gnd.n3522 gnd.n3513 0.155672
R12325 gnd.n3522 gnd.n3521 0.155672
R12326 gnd.n3505 gnd.n3477 0.155672
R12327 gnd.n3498 gnd.n3477 0.155672
R12328 gnd.n3498 gnd.n3497 0.155672
R12329 gnd.n3497 gnd.n3481 0.155672
R12330 gnd.n3490 gnd.n3481 0.155672
R12331 gnd.n3490 gnd.n3489 0.155672
R12332 gnd.n3473 gnd.n3445 0.155672
R12333 gnd.n3466 gnd.n3445 0.155672
R12334 gnd.n3466 gnd.n3465 0.155672
R12335 gnd.n3465 gnd.n3449 0.155672
R12336 gnd.n3458 gnd.n3449 0.155672
R12337 gnd.n3458 gnd.n3457 0.155672
R12338 gnd.n3442 gnd.n3414 0.155672
R12339 gnd.n3435 gnd.n3414 0.155672
R12340 gnd.n3435 gnd.n3434 0.155672
R12341 gnd.n3434 gnd.n3418 0.155672
R12342 gnd.n3427 gnd.n3418 0.155672
R12343 gnd.n3427 gnd.n3426 0.155672
R12344 gnd.n3410 gnd.n3382 0.155672
R12345 gnd.n3403 gnd.n3382 0.155672
R12346 gnd.n3403 gnd.n3402 0.155672
R12347 gnd.n3402 gnd.n3386 0.155672
R12348 gnd.n3395 gnd.n3386 0.155672
R12349 gnd.n3395 gnd.n3394 0.155672
R12350 gnd.n3378 gnd.n3350 0.155672
R12351 gnd.n3371 gnd.n3350 0.155672
R12352 gnd.n3371 gnd.n3370 0.155672
R12353 gnd.n3370 gnd.n3354 0.155672
R12354 gnd.n3363 gnd.n3354 0.155672
R12355 gnd.n3363 gnd.n3362 0.155672
R12356 gnd.n3346 gnd.n3318 0.155672
R12357 gnd.n3339 gnd.n3318 0.155672
R12358 gnd.n3339 gnd.n3338 0.155672
R12359 gnd.n3338 gnd.n3322 0.155672
R12360 gnd.n3331 gnd.n3322 0.155672
R12361 gnd.n3331 gnd.n3330 0.155672
R12362 gnd.n3315 gnd.n3287 0.155672
R12363 gnd.n3308 gnd.n3287 0.155672
R12364 gnd.n3308 gnd.n3307 0.155672
R12365 gnd.n3307 gnd.n3291 0.155672
R12366 gnd.n3300 gnd.n3291 0.155672
R12367 gnd.n3300 gnd.n3299 0.155672
R12368 gnd.n3662 gnd.n2230 0.152939
R12369 gnd.n3662 gnd.n3661 0.152939
R12370 gnd.n3661 gnd.n3660 0.152939
R12371 gnd.n3660 gnd.n2232 0.152939
R12372 gnd.n2233 gnd.n2232 0.152939
R12373 gnd.n2234 gnd.n2233 0.152939
R12374 gnd.n2235 gnd.n2234 0.152939
R12375 gnd.n2236 gnd.n2235 0.152939
R12376 gnd.n2237 gnd.n2236 0.152939
R12377 gnd.n2238 gnd.n2237 0.152939
R12378 gnd.n2239 gnd.n2238 0.152939
R12379 gnd.n2240 gnd.n2239 0.152939
R12380 gnd.n2241 gnd.n2240 0.152939
R12381 gnd.n2242 gnd.n2241 0.152939
R12382 gnd.n3632 gnd.n2242 0.152939
R12383 gnd.n3632 gnd.n3631 0.152939
R12384 gnd.n2904 gnd.n2903 0.152939
R12385 gnd.n2904 gnd.n2608 0.152939
R12386 gnd.n2932 gnd.n2608 0.152939
R12387 gnd.n2933 gnd.n2932 0.152939
R12388 gnd.n2934 gnd.n2933 0.152939
R12389 gnd.n2935 gnd.n2934 0.152939
R12390 gnd.n2935 gnd.n2580 0.152939
R12391 gnd.n2962 gnd.n2580 0.152939
R12392 gnd.n2963 gnd.n2962 0.152939
R12393 gnd.n2964 gnd.n2963 0.152939
R12394 gnd.n2964 gnd.n2558 0.152939
R12395 gnd.n2993 gnd.n2558 0.152939
R12396 gnd.n2994 gnd.n2993 0.152939
R12397 gnd.n2995 gnd.n2994 0.152939
R12398 gnd.n2996 gnd.n2995 0.152939
R12399 gnd.n2998 gnd.n2996 0.152939
R12400 gnd.n2998 gnd.n2997 0.152939
R12401 gnd.n2997 gnd.n2507 0.152939
R12402 gnd.n2508 gnd.n2507 0.152939
R12403 gnd.n2509 gnd.n2508 0.152939
R12404 gnd.n2528 gnd.n2509 0.152939
R12405 gnd.n2529 gnd.n2528 0.152939
R12406 gnd.n2529 gnd.n2427 0.152939
R12407 gnd.n3088 gnd.n2427 0.152939
R12408 gnd.n3089 gnd.n3088 0.152939
R12409 gnd.n3090 gnd.n3089 0.152939
R12410 gnd.n3091 gnd.n3090 0.152939
R12411 gnd.n3091 gnd.n2400 0.152939
R12412 gnd.n3128 gnd.n2400 0.152939
R12413 gnd.n3129 gnd.n3128 0.152939
R12414 gnd.n3130 gnd.n3129 0.152939
R12415 gnd.n3131 gnd.n3130 0.152939
R12416 gnd.n3131 gnd.n2373 0.152939
R12417 gnd.n3173 gnd.n2373 0.152939
R12418 gnd.n3174 gnd.n3173 0.152939
R12419 gnd.n3175 gnd.n3174 0.152939
R12420 gnd.n3176 gnd.n3175 0.152939
R12421 gnd.n3176 gnd.n2345 0.152939
R12422 gnd.n3213 gnd.n2345 0.152939
R12423 gnd.n3214 gnd.n3213 0.152939
R12424 gnd.n3215 gnd.n3214 0.152939
R12425 gnd.n3216 gnd.n3215 0.152939
R12426 gnd.n3216 gnd.n2318 0.152939
R12427 gnd.n3262 gnd.n2318 0.152939
R12428 gnd.n3263 gnd.n3262 0.152939
R12429 gnd.n3264 gnd.n3263 0.152939
R12430 gnd.n3265 gnd.n3264 0.152939
R12431 gnd.n3265 gnd.n2291 0.152939
R12432 gnd.n3556 gnd.n2291 0.152939
R12433 gnd.n3557 gnd.n3556 0.152939
R12434 gnd.n3558 gnd.n3557 0.152939
R12435 gnd.n3559 gnd.n3558 0.152939
R12436 gnd.n3560 gnd.n3559 0.152939
R12437 gnd.n2902 gnd.n2632 0.152939
R12438 gnd.n2653 gnd.n2632 0.152939
R12439 gnd.n2654 gnd.n2653 0.152939
R12440 gnd.n2660 gnd.n2654 0.152939
R12441 gnd.n2661 gnd.n2660 0.152939
R12442 gnd.n2662 gnd.n2661 0.152939
R12443 gnd.n2662 gnd.n2651 0.152939
R12444 gnd.n2670 gnd.n2651 0.152939
R12445 gnd.n2671 gnd.n2670 0.152939
R12446 gnd.n2672 gnd.n2671 0.152939
R12447 gnd.n2672 gnd.n2649 0.152939
R12448 gnd.n2680 gnd.n2649 0.152939
R12449 gnd.n2681 gnd.n2680 0.152939
R12450 gnd.n2682 gnd.n2681 0.152939
R12451 gnd.n2682 gnd.n2647 0.152939
R12452 gnd.n2690 gnd.n2647 0.152939
R12453 gnd.n3629 gnd.n2247 0.152939
R12454 gnd.n2249 gnd.n2247 0.152939
R12455 gnd.n2250 gnd.n2249 0.152939
R12456 gnd.n2251 gnd.n2250 0.152939
R12457 gnd.n2252 gnd.n2251 0.152939
R12458 gnd.n2253 gnd.n2252 0.152939
R12459 gnd.n2254 gnd.n2253 0.152939
R12460 gnd.n2255 gnd.n2254 0.152939
R12461 gnd.n2256 gnd.n2255 0.152939
R12462 gnd.n2257 gnd.n2256 0.152939
R12463 gnd.n2258 gnd.n2257 0.152939
R12464 gnd.n2259 gnd.n2258 0.152939
R12465 gnd.n2260 gnd.n2259 0.152939
R12466 gnd.n2261 gnd.n2260 0.152939
R12467 gnd.n2262 gnd.n2261 0.152939
R12468 gnd.n2263 gnd.n2262 0.152939
R12469 gnd.n2264 gnd.n2263 0.152939
R12470 gnd.n2265 gnd.n2264 0.152939
R12471 gnd.n2266 gnd.n2265 0.152939
R12472 gnd.n2267 gnd.n2266 0.152939
R12473 gnd.n2268 gnd.n2267 0.152939
R12474 gnd.n2269 gnd.n2268 0.152939
R12475 gnd.n2273 gnd.n2269 0.152939
R12476 gnd.n2274 gnd.n2273 0.152939
R12477 gnd.n2275 gnd.n2274 0.152939
R12478 gnd.n2276 gnd.n2275 0.152939
R12479 gnd.n3065 gnd.n3064 0.152939
R12480 gnd.n3066 gnd.n3065 0.152939
R12481 gnd.n3067 gnd.n3066 0.152939
R12482 gnd.n3068 gnd.n3067 0.152939
R12483 gnd.n3069 gnd.n3068 0.152939
R12484 gnd.n3070 gnd.n3069 0.152939
R12485 gnd.n3070 gnd.n2381 0.152939
R12486 gnd.n3149 gnd.n2381 0.152939
R12487 gnd.n3150 gnd.n3149 0.152939
R12488 gnd.n3151 gnd.n3150 0.152939
R12489 gnd.n3152 gnd.n3151 0.152939
R12490 gnd.n3153 gnd.n3152 0.152939
R12491 gnd.n3154 gnd.n3153 0.152939
R12492 gnd.n3155 gnd.n3154 0.152939
R12493 gnd.n3156 gnd.n3155 0.152939
R12494 gnd.n3157 gnd.n3156 0.152939
R12495 gnd.n3157 gnd.n2325 0.152939
R12496 gnd.n3234 gnd.n2325 0.152939
R12497 gnd.n3235 gnd.n3234 0.152939
R12498 gnd.n3236 gnd.n3235 0.152939
R12499 gnd.n3237 gnd.n3236 0.152939
R12500 gnd.n3238 gnd.n3237 0.152939
R12501 gnd.n3239 gnd.n3238 0.152939
R12502 gnd.n3240 gnd.n3239 0.152939
R12503 gnd.n3241 gnd.n3240 0.152939
R12504 gnd.n3242 gnd.n3241 0.152939
R12505 gnd.n3244 gnd.n3242 0.152939
R12506 gnd.n3244 gnd.n3243 0.152939
R12507 gnd.n2820 gnd.n2819 0.152939
R12508 gnd.n2820 gnd.n2710 0.152939
R12509 gnd.n2835 gnd.n2710 0.152939
R12510 gnd.n2836 gnd.n2835 0.152939
R12511 gnd.n2837 gnd.n2836 0.152939
R12512 gnd.n2837 gnd.n2698 0.152939
R12513 gnd.n2851 gnd.n2698 0.152939
R12514 gnd.n2852 gnd.n2851 0.152939
R12515 gnd.n2853 gnd.n2852 0.152939
R12516 gnd.n2854 gnd.n2853 0.152939
R12517 gnd.n2855 gnd.n2854 0.152939
R12518 gnd.n2856 gnd.n2855 0.152939
R12519 gnd.n2857 gnd.n2856 0.152939
R12520 gnd.n2858 gnd.n2857 0.152939
R12521 gnd.n2859 gnd.n2858 0.152939
R12522 gnd.n2860 gnd.n2859 0.152939
R12523 gnd.n2861 gnd.n2860 0.152939
R12524 gnd.n2862 gnd.n2861 0.152939
R12525 gnd.n2863 gnd.n2862 0.152939
R12526 gnd.n2864 gnd.n2863 0.152939
R12527 gnd.n2865 gnd.n2864 0.152939
R12528 gnd.n2865 gnd.n2564 0.152939
R12529 gnd.n2982 gnd.n2564 0.152939
R12530 gnd.n2983 gnd.n2982 0.152939
R12531 gnd.n2984 gnd.n2983 0.152939
R12532 gnd.n2985 gnd.n2984 0.152939
R12533 gnd.n2985 gnd.n2486 0.152939
R12534 gnd.n3062 gnd.n2486 0.152939
R12535 gnd.n2738 gnd.n2737 0.152939
R12536 gnd.n2739 gnd.n2738 0.152939
R12537 gnd.n2740 gnd.n2739 0.152939
R12538 gnd.n2741 gnd.n2740 0.152939
R12539 gnd.n2742 gnd.n2741 0.152939
R12540 gnd.n2743 gnd.n2742 0.152939
R12541 gnd.n2744 gnd.n2743 0.152939
R12542 gnd.n2745 gnd.n2744 0.152939
R12543 gnd.n2746 gnd.n2745 0.152939
R12544 gnd.n2747 gnd.n2746 0.152939
R12545 gnd.n2748 gnd.n2747 0.152939
R12546 gnd.n2749 gnd.n2748 0.152939
R12547 gnd.n2750 gnd.n2749 0.152939
R12548 gnd.n2751 gnd.n2750 0.152939
R12549 gnd.n2752 gnd.n2751 0.152939
R12550 gnd.n2753 gnd.n2752 0.152939
R12551 gnd.n2754 gnd.n2753 0.152939
R12552 gnd.n2755 gnd.n2754 0.152939
R12553 gnd.n2756 gnd.n2755 0.152939
R12554 gnd.n2757 gnd.n2756 0.152939
R12555 gnd.n2758 gnd.n2757 0.152939
R12556 gnd.n2759 gnd.n2758 0.152939
R12557 gnd.n2763 gnd.n2759 0.152939
R12558 gnd.n2764 gnd.n2763 0.152939
R12559 gnd.n2764 gnd.n2721 0.152939
R12560 gnd.n2818 gnd.n2721 0.152939
R12561 gnd.n6142 gnd.n558 0.152939
R12562 gnd.n6150 gnd.n558 0.152939
R12563 gnd.n6151 gnd.n6150 0.152939
R12564 gnd.n6152 gnd.n6151 0.152939
R12565 gnd.n6152 gnd.n552 0.152939
R12566 gnd.n6160 gnd.n552 0.152939
R12567 gnd.n6161 gnd.n6160 0.152939
R12568 gnd.n6162 gnd.n6161 0.152939
R12569 gnd.n6162 gnd.n546 0.152939
R12570 gnd.n6170 gnd.n546 0.152939
R12571 gnd.n6171 gnd.n6170 0.152939
R12572 gnd.n6172 gnd.n6171 0.152939
R12573 gnd.n6172 gnd.n540 0.152939
R12574 gnd.n6180 gnd.n540 0.152939
R12575 gnd.n6181 gnd.n6180 0.152939
R12576 gnd.n6182 gnd.n6181 0.152939
R12577 gnd.n6182 gnd.n534 0.152939
R12578 gnd.n6190 gnd.n534 0.152939
R12579 gnd.n6191 gnd.n6190 0.152939
R12580 gnd.n6192 gnd.n6191 0.152939
R12581 gnd.n6192 gnd.n528 0.152939
R12582 gnd.n6200 gnd.n528 0.152939
R12583 gnd.n6201 gnd.n6200 0.152939
R12584 gnd.n6202 gnd.n6201 0.152939
R12585 gnd.n6202 gnd.n522 0.152939
R12586 gnd.n6210 gnd.n522 0.152939
R12587 gnd.n6211 gnd.n6210 0.152939
R12588 gnd.n6212 gnd.n6211 0.152939
R12589 gnd.n6212 gnd.n516 0.152939
R12590 gnd.n6220 gnd.n516 0.152939
R12591 gnd.n6221 gnd.n6220 0.152939
R12592 gnd.n6222 gnd.n6221 0.152939
R12593 gnd.n6222 gnd.n510 0.152939
R12594 gnd.n6230 gnd.n510 0.152939
R12595 gnd.n6231 gnd.n6230 0.152939
R12596 gnd.n6232 gnd.n6231 0.152939
R12597 gnd.n6232 gnd.n504 0.152939
R12598 gnd.n6240 gnd.n504 0.152939
R12599 gnd.n6241 gnd.n6240 0.152939
R12600 gnd.n6242 gnd.n6241 0.152939
R12601 gnd.n6242 gnd.n498 0.152939
R12602 gnd.n6250 gnd.n498 0.152939
R12603 gnd.n6251 gnd.n6250 0.152939
R12604 gnd.n6252 gnd.n6251 0.152939
R12605 gnd.n6252 gnd.n492 0.152939
R12606 gnd.n6260 gnd.n492 0.152939
R12607 gnd.n6261 gnd.n6260 0.152939
R12608 gnd.n6262 gnd.n6261 0.152939
R12609 gnd.n6262 gnd.n486 0.152939
R12610 gnd.n6270 gnd.n486 0.152939
R12611 gnd.n6271 gnd.n6270 0.152939
R12612 gnd.n6272 gnd.n6271 0.152939
R12613 gnd.n6272 gnd.n480 0.152939
R12614 gnd.n6280 gnd.n480 0.152939
R12615 gnd.n6281 gnd.n6280 0.152939
R12616 gnd.n6282 gnd.n6281 0.152939
R12617 gnd.n6282 gnd.n474 0.152939
R12618 gnd.n6290 gnd.n474 0.152939
R12619 gnd.n6291 gnd.n6290 0.152939
R12620 gnd.n6292 gnd.n6291 0.152939
R12621 gnd.n6292 gnd.n468 0.152939
R12622 gnd.n6300 gnd.n468 0.152939
R12623 gnd.n6301 gnd.n6300 0.152939
R12624 gnd.n6302 gnd.n6301 0.152939
R12625 gnd.n6302 gnd.n462 0.152939
R12626 gnd.n6310 gnd.n462 0.152939
R12627 gnd.n6311 gnd.n6310 0.152939
R12628 gnd.n6312 gnd.n6311 0.152939
R12629 gnd.n6312 gnd.n456 0.152939
R12630 gnd.n6320 gnd.n456 0.152939
R12631 gnd.n6321 gnd.n6320 0.152939
R12632 gnd.n6322 gnd.n6321 0.152939
R12633 gnd.n6322 gnd.n450 0.152939
R12634 gnd.n6330 gnd.n450 0.152939
R12635 gnd.n6331 gnd.n6330 0.152939
R12636 gnd.n6332 gnd.n6331 0.152939
R12637 gnd.n6332 gnd.n444 0.152939
R12638 gnd.n6340 gnd.n444 0.152939
R12639 gnd.n6341 gnd.n6340 0.152939
R12640 gnd.n6342 gnd.n6341 0.152939
R12641 gnd.n6342 gnd.n438 0.152939
R12642 gnd.n6350 gnd.n438 0.152939
R12643 gnd.n6351 gnd.n6350 0.152939
R12644 gnd.n6352 gnd.n6351 0.152939
R12645 gnd.n6352 gnd.n432 0.152939
R12646 gnd.n6360 gnd.n432 0.152939
R12647 gnd.n6361 gnd.n6360 0.152939
R12648 gnd.n6362 gnd.n6361 0.152939
R12649 gnd.n6362 gnd.n426 0.152939
R12650 gnd.n6370 gnd.n426 0.152939
R12651 gnd.n6371 gnd.n6370 0.152939
R12652 gnd.n6372 gnd.n6371 0.152939
R12653 gnd.n6372 gnd.n420 0.152939
R12654 gnd.n6380 gnd.n420 0.152939
R12655 gnd.n6381 gnd.n6380 0.152939
R12656 gnd.n6382 gnd.n6381 0.152939
R12657 gnd.n6382 gnd.n414 0.152939
R12658 gnd.n6390 gnd.n414 0.152939
R12659 gnd.n6391 gnd.n6390 0.152939
R12660 gnd.n6392 gnd.n6391 0.152939
R12661 gnd.n6392 gnd.n408 0.152939
R12662 gnd.n6400 gnd.n408 0.152939
R12663 gnd.n6401 gnd.n6400 0.152939
R12664 gnd.n6402 gnd.n6401 0.152939
R12665 gnd.n6402 gnd.n402 0.152939
R12666 gnd.n6410 gnd.n402 0.152939
R12667 gnd.n6411 gnd.n6410 0.152939
R12668 gnd.n6412 gnd.n6411 0.152939
R12669 gnd.n6412 gnd.n396 0.152939
R12670 gnd.n6420 gnd.n396 0.152939
R12671 gnd.n6421 gnd.n6420 0.152939
R12672 gnd.n6422 gnd.n6421 0.152939
R12673 gnd.n6422 gnd.n390 0.152939
R12674 gnd.n6430 gnd.n390 0.152939
R12675 gnd.n6431 gnd.n6430 0.152939
R12676 gnd.n6432 gnd.n6431 0.152939
R12677 gnd.n6432 gnd.n384 0.152939
R12678 gnd.n6440 gnd.n384 0.152939
R12679 gnd.n6441 gnd.n6440 0.152939
R12680 gnd.n6442 gnd.n6441 0.152939
R12681 gnd.n6442 gnd.n378 0.152939
R12682 gnd.n6450 gnd.n378 0.152939
R12683 gnd.n6451 gnd.n6450 0.152939
R12684 gnd.n6452 gnd.n6451 0.152939
R12685 gnd.n6452 gnd.n372 0.152939
R12686 gnd.n6460 gnd.n372 0.152939
R12687 gnd.n6461 gnd.n6460 0.152939
R12688 gnd.n6462 gnd.n6461 0.152939
R12689 gnd.n6462 gnd.n366 0.152939
R12690 gnd.n6470 gnd.n366 0.152939
R12691 gnd.n6471 gnd.n6470 0.152939
R12692 gnd.n6472 gnd.n6471 0.152939
R12693 gnd.n6472 gnd.n360 0.152939
R12694 gnd.n6480 gnd.n360 0.152939
R12695 gnd.n6481 gnd.n6480 0.152939
R12696 gnd.n6482 gnd.n6481 0.152939
R12697 gnd.n6482 gnd.n354 0.152939
R12698 gnd.n6490 gnd.n354 0.152939
R12699 gnd.n6491 gnd.n6490 0.152939
R12700 gnd.n6492 gnd.n6491 0.152939
R12701 gnd.n6492 gnd.n348 0.152939
R12702 gnd.n6500 gnd.n348 0.152939
R12703 gnd.n6501 gnd.n6500 0.152939
R12704 gnd.n6502 gnd.n6501 0.152939
R12705 gnd.n6502 gnd.n342 0.152939
R12706 gnd.n6510 gnd.n342 0.152939
R12707 gnd.n6511 gnd.n6510 0.152939
R12708 gnd.n6512 gnd.n6511 0.152939
R12709 gnd.n6512 gnd.n336 0.152939
R12710 gnd.n6520 gnd.n336 0.152939
R12711 gnd.n6521 gnd.n6520 0.152939
R12712 gnd.n6522 gnd.n6521 0.152939
R12713 gnd.n6522 gnd.n330 0.152939
R12714 gnd.n6530 gnd.n330 0.152939
R12715 gnd.n6531 gnd.n6530 0.152939
R12716 gnd.n6532 gnd.n6531 0.152939
R12717 gnd.n6532 gnd.n324 0.152939
R12718 gnd.n6540 gnd.n324 0.152939
R12719 gnd.n6541 gnd.n6540 0.152939
R12720 gnd.n6542 gnd.n6541 0.152939
R12721 gnd.n6542 gnd.n318 0.152939
R12722 gnd.n6550 gnd.n318 0.152939
R12723 gnd.n6551 gnd.n6550 0.152939
R12724 gnd.n6553 gnd.n6551 0.152939
R12725 gnd.n6553 gnd.n6552 0.152939
R12726 gnd.n6552 gnd.n312 0.152939
R12727 gnd.n6562 gnd.n312 0.152939
R12728 gnd.n6563 gnd.n307 0.152939
R12729 gnd.n6571 gnd.n307 0.152939
R12730 gnd.n6572 gnd.n6571 0.152939
R12731 gnd.n6573 gnd.n6572 0.152939
R12732 gnd.n6573 gnd.n301 0.152939
R12733 gnd.n6581 gnd.n301 0.152939
R12734 gnd.n6582 gnd.n6581 0.152939
R12735 gnd.n6583 gnd.n6582 0.152939
R12736 gnd.n6583 gnd.n295 0.152939
R12737 gnd.n6591 gnd.n295 0.152939
R12738 gnd.n6592 gnd.n6591 0.152939
R12739 gnd.n6593 gnd.n6592 0.152939
R12740 gnd.n6593 gnd.n289 0.152939
R12741 gnd.n6601 gnd.n289 0.152939
R12742 gnd.n6602 gnd.n6601 0.152939
R12743 gnd.n6603 gnd.n6602 0.152939
R12744 gnd.n6603 gnd.n283 0.152939
R12745 gnd.n6611 gnd.n283 0.152939
R12746 gnd.n6612 gnd.n6611 0.152939
R12747 gnd.n6613 gnd.n6612 0.152939
R12748 gnd.n6613 gnd.n277 0.152939
R12749 gnd.n6621 gnd.n277 0.152939
R12750 gnd.n6622 gnd.n6621 0.152939
R12751 gnd.n6623 gnd.n6622 0.152939
R12752 gnd.n6623 gnd.n271 0.152939
R12753 gnd.n6631 gnd.n271 0.152939
R12754 gnd.n6632 gnd.n6631 0.152939
R12755 gnd.n6633 gnd.n6632 0.152939
R12756 gnd.n6633 gnd.n265 0.152939
R12757 gnd.n6641 gnd.n265 0.152939
R12758 gnd.n6642 gnd.n6641 0.152939
R12759 gnd.n6643 gnd.n6642 0.152939
R12760 gnd.n6643 gnd.n259 0.152939
R12761 gnd.n6651 gnd.n259 0.152939
R12762 gnd.n6652 gnd.n6651 0.152939
R12763 gnd.n6653 gnd.n6652 0.152939
R12764 gnd.n6653 gnd.n253 0.152939
R12765 gnd.n6661 gnd.n253 0.152939
R12766 gnd.n6662 gnd.n6661 0.152939
R12767 gnd.n6663 gnd.n6662 0.152939
R12768 gnd.n6663 gnd.n247 0.152939
R12769 gnd.n6671 gnd.n247 0.152939
R12770 gnd.n6672 gnd.n6671 0.152939
R12771 gnd.n6673 gnd.n6672 0.152939
R12772 gnd.n6673 gnd.n241 0.152939
R12773 gnd.n6681 gnd.n241 0.152939
R12774 gnd.n6682 gnd.n6681 0.152939
R12775 gnd.n6683 gnd.n6682 0.152939
R12776 gnd.n6683 gnd.n235 0.152939
R12777 gnd.n6691 gnd.n235 0.152939
R12778 gnd.n6692 gnd.n6691 0.152939
R12779 gnd.n6693 gnd.n6692 0.152939
R12780 gnd.n6693 gnd.n229 0.152939
R12781 gnd.n6701 gnd.n229 0.152939
R12782 gnd.n6702 gnd.n6701 0.152939
R12783 gnd.n6703 gnd.n6702 0.152939
R12784 gnd.n6703 gnd.n223 0.152939
R12785 gnd.n6711 gnd.n223 0.152939
R12786 gnd.n6712 gnd.n6711 0.152939
R12787 gnd.n6713 gnd.n6712 0.152939
R12788 gnd.n6713 gnd.n217 0.152939
R12789 gnd.n6721 gnd.n217 0.152939
R12790 gnd.n6722 gnd.n6721 0.152939
R12791 gnd.n6723 gnd.n6722 0.152939
R12792 gnd.n6723 gnd.n211 0.152939
R12793 gnd.n6731 gnd.n211 0.152939
R12794 gnd.n6732 gnd.n6731 0.152939
R12795 gnd.n6733 gnd.n6732 0.152939
R12796 gnd.n6733 gnd.n205 0.152939
R12797 gnd.n6741 gnd.n205 0.152939
R12798 gnd.n6742 gnd.n6741 0.152939
R12799 gnd.n6743 gnd.n6742 0.152939
R12800 gnd.n6743 gnd.n199 0.152939
R12801 gnd.n6751 gnd.n199 0.152939
R12802 gnd.n6752 gnd.n6751 0.152939
R12803 gnd.n6753 gnd.n6752 0.152939
R12804 gnd.n6753 gnd.n193 0.152939
R12805 gnd.n6761 gnd.n193 0.152939
R12806 gnd.n6762 gnd.n6761 0.152939
R12807 gnd.n6763 gnd.n6762 0.152939
R12808 gnd.n6763 gnd.n187 0.152939
R12809 gnd.n6772 gnd.n187 0.152939
R12810 gnd.n6773 gnd.n6772 0.152939
R12811 gnd.n6774 gnd.n6773 0.152939
R12812 gnd.n7198 gnd.n81 0.152939
R12813 gnd.n106 gnd.n81 0.152939
R12814 gnd.n107 gnd.n106 0.152939
R12815 gnd.n108 gnd.n107 0.152939
R12816 gnd.n124 gnd.n108 0.152939
R12817 gnd.n125 gnd.n124 0.152939
R12818 gnd.n126 gnd.n125 0.152939
R12819 gnd.n127 gnd.n126 0.152939
R12820 gnd.n144 gnd.n127 0.152939
R12821 gnd.n145 gnd.n144 0.152939
R12822 gnd.n146 gnd.n145 0.152939
R12823 gnd.n147 gnd.n146 0.152939
R12824 gnd.n162 gnd.n147 0.152939
R12825 gnd.n163 gnd.n162 0.152939
R12826 gnd.n164 gnd.n163 0.152939
R12827 gnd.n165 gnd.n164 0.152939
R12828 gnd.n7207 gnd.n69 0.152939
R12829 gnd.n176 gnd.n69 0.152939
R12830 gnd.n6794 gnd.n176 0.152939
R12831 gnd.n6795 gnd.n6794 0.152939
R12832 gnd.n6796 gnd.n6795 0.152939
R12833 gnd.n6797 gnd.n6796 0.152939
R12834 gnd.n6798 gnd.n6797 0.152939
R12835 gnd.n6799 gnd.n6798 0.152939
R12836 gnd.n6800 gnd.n6799 0.152939
R12837 gnd.n6801 gnd.n6800 0.152939
R12838 gnd.n6802 gnd.n6801 0.152939
R12839 gnd.n6803 gnd.n6802 0.152939
R12840 gnd.n6804 gnd.n6803 0.152939
R12841 gnd.n6805 gnd.n6804 0.152939
R12842 gnd.n6806 gnd.n6805 0.152939
R12843 gnd.n6807 gnd.n6806 0.152939
R12844 gnd.n6808 gnd.n6807 0.152939
R12845 gnd.n6809 gnd.n6808 0.152939
R12846 gnd.n6810 gnd.n6809 0.152939
R12847 gnd.n7091 gnd.n6810 0.152939
R12848 gnd.n6832 gnd.n6831 0.152939
R12849 gnd.n6839 gnd.n6831 0.152939
R12850 gnd.n6840 gnd.n6839 0.152939
R12851 gnd.n6841 gnd.n6840 0.152939
R12852 gnd.n6841 gnd.n6829 0.152939
R12853 gnd.n6849 gnd.n6829 0.152939
R12854 gnd.n6850 gnd.n6849 0.152939
R12855 gnd.n6851 gnd.n6850 0.152939
R12856 gnd.n6851 gnd.n6827 0.152939
R12857 gnd.n6859 gnd.n6827 0.152939
R12858 gnd.n6860 gnd.n6859 0.152939
R12859 gnd.n6861 gnd.n6860 0.152939
R12860 gnd.n6861 gnd.n6825 0.152939
R12861 gnd.n6868 gnd.n6825 0.152939
R12862 gnd.n6869 gnd.n6868 0.152939
R12863 gnd.n6870 gnd.n6869 0.152939
R12864 gnd.n6870 gnd.n6811 0.152939
R12865 gnd.n7090 gnd.n6811 0.152939
R12866 gnd.n6907 gnd.n6906 0.152939
R12867 gnd.n6908 gnd.n6907 0.152939
R12868 gnd.n6909 gnd.n6908 0.152939
R12869 gnd.n6910 gnd.n6909 0.152939
R12870 gnd.n6911 gnd.n6910 0.152939
R12871 gnd.n6912 gnd.n6911 0.152939
R12872 gnd.n6913 gnd.n6912 0.152939
R12873 gnd.n6914 gnd.n6913 0.152939
R12874 gnd.n6915 gnd.n6914 0.152939
R12875 gnd.n6916 gnd.n6915 0.152939
R12876 gnd.n6917 gnd.n6916 0.152939
R12877 gnd.n6918 gnd.n6917 0.152939
R12878 gnd.n6919 gnd.n6918 0.152939
R12879 gnd.n6920 gnd.n6919 0.152939
R12880 gnd.n6921 gnd.n6920 0.152939
R12881 gnd.n6922 gnd.n6921 0.152939
R12882 gnd.n6923 gnd.n6922 0.152939
R12883 gnd.n6924 gnd.n6923 0.152939
R12884 gnd.n6925 gnd.n6924 0.152939
R12885 gnd.n6926 gnd.n6925 0.152939
R12886 gnd.n6927 gnd.n6926 0.152939
R12887 gnd.n6928 gnd.n6927 0.152939
R12888 gnd.n6929 gnd.n6928 0.152939
R12889 gnd.n6930 gnd.n6929 0.152939
R12890 gnd.n6931 gnd.n6930 0.152939
R12891 gnd.n6932 gnd.n6931 0.152939
R12892 gnd.n6933 gnd.n6932 0.152939
R12893 gnd.n6934 gnd.n6933 0.152939
R12894 gnd.n6935 gnd.n6934 0.152939
R12895 gnd.n6936 gnd.n6935 0.152939
R12896 gnd.n6937 gnd.n6936 0.152939
R12897 gnd.n6938 gnd.n6937 0.152939
R12898 gnd.n6939 gnd.n6938 0.152939
R12899 gnd.n6940 gnd.n6939 0.152939
R12900 gnd.n6941 gnd.n6940 0.152939
R12901 gnd.n6942 gnd.n6941 0.152939
R12902 gnd.n7010 gnd.n6942 0.152939
R12903 gnd.n7010 gnd.n7009 0.152939
R12904 gnd.n7009 gnd.n7008 0.152939
R12905 gnd.n7008 gnd.n6946 0.152939
R12906 gnd.n6947 gnd.n6946 0.152939
R12907 gnd.n6948 gnd.n6947 0.152939
R12908 gnd.n6949 gnd.n6948 0.152939
R12909 gnd.n6950 gnd.n6949 0.152939
R12910 gnd.n6951 gnd.n6950 0.152939
R12911 gnd.n6952 gnd.n6951 0.152939
R12912 gnd.n6953 gnd.n6952 0.152939
R12913 gnd.n6954 gnd.n6953 0.152939
R12914 gnd.n6955 gnd.n6954 0.152939
R12915 gnd.n6956 gnd.n6955 0.152939
R12916 gnd.n6957 gnd.n6956 0.152939
R12917 gnd.n6958 gnd.n6957 0.152939
R12918 gnd.n6959 gnd.n6958 0.152939
R12919 gnd.n6960 gnd.n6959 0.152939
R12920 gnd.n6961 gnd.n6960 0.152939
R12921 gnd.n6962 gnd.n6961 0.152939
R12922 gnd.n6968 gnd.n6962 0.152939
R12923 gnd.n6968 gnd.n6967 0.152939
R12924 gnd.n1421 gnd.n1420 0.152939
R12925 gnd.n1422 gnd.n1421 0.152939
R12926 gnd.n1423 gnd.n1422 0.152939
R12927 gnd.n1424 gnd.n1423 0.152939
R12928 gnd.n1425 gnd.n1424 0.152939
R12929 gnd.n1426 gnd.n1425 0.152939
R12930 gnd.n1427 gnd.n1426 0.152939
R12931 gnd.n1428 gnd.n1427 0.152939
R12932 gnd.n1429 gnd.n1428 0.152939
R12933 gnd.n1430 gnd.n1429 0.152939
R12934 gnd.n1431 gnd.n1430 0.152939
R12935 gnd.n1432 gnd.n1431 0.152939
R12936 gnd.n1433 gnd.n1432 0.152939
R12937 gnd.n1434 gnd.n1433 0.152939
R12938 gnd.n1435 gnd.n1434 0.152939
R12939 gnd.n1436 gnd.n1435 0.152939
R12940 gnd.n1437 gnd.n1436 0.152939
R12941 gnd.n1440 gnd.n1437 0.152939
R12942 gnd.n1441 gnd.n1440 0.152939
R12943 gnd.n1442 gnd.n1441 0.152939
R12944 gnd.n1443 gnd.n1442 0.152939
R12945 gnd.n1444 gnd.n1443 0.152939
R12946 gnd.n1445 gnd.n1444 0.152939
R12947 gnd.n1446 gnd.n1445 0.152939
R12948 gnd.n1447 gnd.n1446 0.152939
R12949 gnd.n1452 gnd.n1451 0.152939
R12950 gnd.n1453 gnd.n1452 0.152939
R12951 gnd.n1454 gnd.n1453 0.152939
R12952 gnd.n1455 gnd.n1454 0.152939
R12953 gnd.n1456 gnd.n1455 0.152939
R12954 gnd.n1457 gnd.n1456 0.152939
R12955 gnd.n1458 gnd.n1457 0.152939
R12956 gnd.n1459 gnd.n1458 0.152939
R12957 gnd.n1460 gnd.n1459 0.152939
R12958 gnd.n1463 gnd.n1460 0.152939
R12959 gnd.n1464 gnd.n1463 0.152939
R12960 gnd.n1465 gnd.n1464 0.152939
R12961 gnd.n1466 gnd.n1465 0.152939
R12962 gnd.n1467 gnd.n1466 0.152939
R12963 gnd.n1468 gnd.n1467 0.152939
R12964 gnd.n1469 gnd.n1468 0.152939
R12965 gnd.n1470 gnd.n1469 0.152939
R12966 gnd.n1471 gnd.n1470 0.152939
R12967 gnd.n1472 gnd.n1471 0.152939
R12968 gnd.n1473 gnd.n1472 0.152939
R12969 gnd.n1474 gnd.n1473 0.152939
R12970 gnd.n1475 gnd.n1474 0.152939
R12971 gnd.n1476 gnd.n1475 0.152939
R12972 gnd.n1477 gnd.n1476 0.152939
R12973 gnd.n1478 gnd.n1477 0.152939
R12974 gnd.n1479 gnd.n1478 0.152939
R12975 gnd.n1480 gnd.n1479 0.152939
R12976 gnd.n1481 gnd.n1480 0.152939
R12977 gnd.n5383 gnd.n1481 0.152939
R12978 gnd.n5383 gnd.n5382 0.152939
R12979 gnd.n1502 gnd.n1501 0.152939
R12980 gnd.n1503 gnd.n1502 0.152939
R12981 gnd.n1504 gnd.n1503 0.152939
R12982 gnd.n1505 gnd.n1504 0.152939
R12983 gnd.n1525 gnd.n1505 0.152939
R12984 gnd.n1526 gnd.n1525 0.152939
R12985 gnd.n1527 gnd.n1526 0.152939
R12986 gnd.n1528 gnd.n1527 0.152939
R12987 gnd.n1546 gnd.n1528 0.152939
R12988 gnd.n1547 gnd.n1546 0.152939
R12989 gnd.n1548 gnd.n1547 0.152939
R12990 gnd.n1549 gnd.n1548 0.152939
R12991 gnd.n1565 gnd.n1549 0.152939
R12992 gnd.n1566 gnd.n1565 0.152939
R12993 gnd.n1566 gnd.n82 0.152939
R12994 gnd.n7198 gnd.n82 0.152939
R12995 gnd.n4129 gnd.n4128 0.152939
R12996 gnd.n4130 gnd.n4129 0.152939
R12997 gnd.n4131 gnd.n4130 0.152939
R12998 gnd.n4134 gnd.n4131 0.152939
R12999 gnd.n4135 gnd.n4134 0.152939
R13000 gnd.n4136 gnd.n4135 0.152939
R13001 gnd.n4137 gnd.n4136 0.152939
R13002 gnd.n4139 gnd.n4137 0.152939
R13003 gnd.n4139 gnd.n4138 0.152939
R13004 gnd.n4138 gnd.n2091 0.152939
R13005 gnd.n4205 gnd.n2091 0.152939
R13006 gnd.n4206 gnd.n4205 0.152939
R13007 gnd.n4207 gnd.n4206 0.152939
R13008 gnd.n4207 gnd.n2087 0.152939
R13009 gnd.n4213 gnd.n2087 0.152939
R13010 gnd.n4214 gnd.n4213 0.152939
R13011 gnd.n4215 gnd.n4214 0.152939
R13012 gnd.n4215 gnd.n2083 0.152939
R13013 gnd.n4222 gnd.n2083 0.152939
R13014 gnd.n4223 gnd.n4222 0.152939
R13015 gnd.n4224 gnd.n4223 0.152939
R13016 gnd.n4224 gnd.n2079 0.152939
R13017 gnd.n4307 gnd.n2079 0.152939
R13018 gnd.n4308 gnd.n4307 0.152939
R13019 gnd.n4309 gnd.n4308 0.152939
R13020 gnd.n4309 gnd.n2064 0.152939
R13021 gnd.n4323 gnd.n2064 0.152939
R13022 gnd.n4324 gnd.n4323 0.152939
R13023 gnd.n4325 gnd.n4324 0.152939
R13024 gnd.n4325 gnd.n2051 0.152939
R13025 gnd.n4339 gnd.n2051 0.152939
R13026 gnd.n4340 gnd.n4339 0.152939
R13027 gnd.n4341 gnd.n4340 0.152939
R13028 gnd.n4341 gnd.n2037 0.152939
R13029 gnd.n4355 gnd.n2037 0.152939
R13030 gnd.n4356 gnd.n4355 0.152939
R13031 gnd.n4357 gnd.n4356 0.152939
R13032 gnd.n4357 gnd.n2023 0.152939
R13033 gnd.n4371 gnd.n2023 0.152939
R13034 gnd.n4372 gnd.n4371 0.152939
R13035 gnd.n4373 gnd.n4372 0.152939
R13036 gnd.n4373 gnd.n2009 0.152939
R13037 gnd.n4387 gnd.n2009 0.152939
R13038 gnd.n4388 gnd.n4387 0.152939
R13039 gnd.n4389 gnd.n4388 0.152939
R13040 gnd.n4389 gnd.n1994 0.152939
R13041 gnd.n4404 gnd.n1994 0.152939
R13042 gnd.n4405 gnd.n4404 0.152939
R13043 gnd.n4406 gnd.n4405 0.152939
R13044 gnd.n4407 gnd.n4406 0.152939
R13045 gnd.n4409 gnd.n4407 0.152939
R13046 gnd.n4409 gnd.n4408 0.152939
R13047 gnd.n4408 gnd.n1208 0.152939
R13048 gnd.n1209 gnd.n1208 0.152939
R13049 gnd.n1210 gnd.n1209 0.152939
R13050 gnd.n1964 gnd.n1210 0.152939
R13051 gnd.n1965 gnd.n1964 0.152939
R13052 gnd.n4562 gnd.n1965 0.152939
R13053 gnd.n4563 gnd.n4562 0.152939
R13054 gnd.n4564 gnd.n4563 0.152939
R13055 gnd.n4564 gnd.n1937 0.152939
R13056 gnd.n4605 gnd.n1937 0.152939
R13057 gnd.n4606 gnd.n4605 0.152939
R13058 gnd.n4607 gnd.n4606 0.152939
R13059 gnd.n4608 gnd.n4607 0.152939
R13060 gnd.n4608 gnd.n1916 0.152939
R13061 gnd.n4665 gnd.n1916 0.152939
R13062 gnd.n4666 gnd.n4665 0.152939
R13063 gnd.n4667 gnd.n4666 0.152939
R13064 gnd.n4668 gnd.n4667 0.152939
R13065 gnd.n4669 gnd.n4668 0.152939
R13066 gnd.n4671 gnd.n4669 0.152939
R13067 gnd.n4672 gnd.n4671 0.152939
R13068 gnd.n4672 gnd.n1879 0.152939
R13069 gnd.n4726 gnd.n1879 0.152939
R13070 gnd.n4727 gnd.n4726 0.152939
R13071 gnd.n4728 gnd.n4727 0.152939
R13072 gnd.n4728 gnd.n1856 0.152939
R13073 gnd.n4772 gnd.n1856 0.152939
R13074 gnd.n4773 gnd.n4772 0.152939
R13075 gnd.n4774 gnd.n4773 0.152939
R13076 gnd.n4775 gnd.n4774 0.152939
R13077 gnd.n4775 gnd.n1835 0.152939
R13078 gnd.n4824 gnd.n1835 0.152939
R13079 gnd.n4825 gnd.n4824 0.152939
R13080 gnd.n4826 gnd.n4825 0.152939
R13081 gnd.n4827 gnd.n4826 0.152939
R13082 gnd.n4827 gnd.n1808 0.152939
R13083 gnd.n4860 gnd.n1808 0.152939
R13084 gnd.n4861 gnd.n4860 0.152939
R13085 gnd.n4862 gnd.n4861 0.152939
R13086 gnd.n4862 gnd.n1752 0.152939
R13087 gnd.n5035 gnd.n1752 0.152939
R13088 gnd.n5036 gnd.n5035 0.152939
R13089 gnd.n5037 gnd.n5036 0.152939
R13090 gnd.n5037 gnd.n1740 0.152939
R13091 gnd.n5051 gnd.n1740 0.152939
R13092 gnd.n5052 gnd.n5051 0.152939
R13093 gnd.n5053 gnd.n5052 0.152939
R13094 gnd.n5053 gnd.n1727 0.152939
R13095 gnd.n5068 gnd.n1727 0.152939
R13096 gnd.n5069 gnd.n5068 0.152939
R13097 gnd.n5070 gnd.n5069 0.152939
R13098 gnd.n5070 gnd.n1715 0.152939
R13099 gnd.n5084 gnd.n1715 0.152939
R13100 gnd.n5085 gnd.n5084 0.152939
R13101 gnd.n5086 gnd.n5085 0.152939
R13102 gnd.n5086 gnd.n1702 0.152939
R13103 gnd.n5100 gnd.n1702 0.152939
R13104 gnd.n5101 gnd.n5100 0.152939
R13105 gnd.n5102 gnd.n5101 0.152939
R13106 gnd.n5102 gnd.n1689 0.152939
R13107 gnd.n5116 gnd.n1689 0.152939
R13108 gnd.n5117 gnd.n5116 0.152939
R13109 gnd.n5118 gnd.n5117 0.152939
R13110 gnd.n5118 gnd.n1676 0.152939
R13111 gnd.n5132 gnd.n1676 0.152939
R13112 gnd.n5133 gnd.n5132 0.152939
R13113 gnd.n5134 gnd.n5133 0.152939
R13114 gnd.n5136 gnd.n5134 0.152939
R13115 gnd.n5136 gnd.n5135 0.152939
R13116 gnd.n5135 gnd.n1663 0.152939
R13117 gnd.n5153 gnd.n1663 0.152939
R13118 gnd.n5154 gnd.n5153 0.152939
R13119 gnd.n5155 gnd.n5154 0.152939
R13120 gnd.n5156 gnd.n5155 0.152939
R13121 gnd.n5157 gnd.n5156 0.152939
R13122 gnd.n5159 gnd.n5157 0.152939
R13123 gnd.n5160 gnd.n5159 0.152939
R13124 gnd.n5160 gnd.n1627 0.152939
R13125 gnd.n5222 gnd.n1627 0.152939
R13126 gnd.n5223 gnd.n5222 0.152939
R13127 gnd.n5224 gnd.n5223 0.152939
R13128 gnd.n5224 gnd.n1623 0.152939
R13129 gnd.n5230 gnd.n1623 0.152939
R13130 gnd.n5231 gnd.n5230 0.152939
R13131 gnd.n5232 gnd.n5231 0.152939
R13132 gnd.n5232 gnd.n1619 0.152939
R13133 gnd.n5238 gnd.n1619 0.152939
R13134 gnd.n5239 gnd.n5238 0.152939
R13135 gnd.n5240 gnd.n5239 0.152939
R13136 gnd.n5241 gnd.n5240 0.152939
R13137 gnd.n5242 gnd.n5241 0.152939
R13138 gnd.n5245 gnd.n5242 0.152939
R13139 gnd.n5246 gnd.n5245 0.152939
R13140 gnd.n3739 gnd.n3738 0.152939
R13141 gnd.n3740 gnd.n3739 0.152939
R13142 gnd.n3740 gnd.n2182 0.152939
R13143 gnd.n3992 gnd.n2182 0.152939
R13144 gnd.n3993 gnd.n3992 0.152939
R13145 gnd.n3994 gnd.n3993 0.152939
R13146 gnd.n3995 gnd.n3994 0.152939
R13147 gnd.n3995 gnd.n2157 0.152939
R13148 gnd.n4027 gnd.n2157 0.152939
R13149 gnd.n4028 gnd.n4027 0.152939
R13150 gnd.n4029 gnd.n4028 0.152939
R13151 gnd.n4030 gnd.n4029 0.152939
R13152 gnd.n4031 gnd.n4030 0.152939
R13153 gnd.n4031 gnd.n2131 0.152939
R13154 gnd.n4067 gnd.n2131 0.152939
R13155 gnd.n4068 gnd.n4067 0.152939
R13156 gnd.n4069 gnd.n4068 0.152939
R13157 gnd.n4069 gnd.n2126 0.152939
R13158 gnd.n4093 gnd.n2126 0.152939
R13159 gnd.n4094 gnd.n4093 0.152939
R13160 gnd.n3690 gnd.n3689 0.152939
R13161 gnd.n3698 gnd.n3689 0.152939
R13162 gnd.n3699 gnd.n3698 0.152939
R13163 gnd.n3700 gnd.n3699 0.152939
R13164 gnd.n3700 gnd.n3685 0.152939
R13165 gnd.n3708 gnd.n3685 0.152939
R13166 gnd.n3709 gnd.n3708 0.152939
R13167 gnd.n3710 gnd.n3709 0.152939
R13168 gnd.n3710 gnd.n3681 0.152939
R13169 gnd.n3718 gnd.n3681 0.152939
R13170 gnd.n3719 gnd.n3718 0.152939
R13171 gnd.n3720 gnd.n3719 0.152939
R13172 gnd.n3720 gnd.n3677 0.152939
R13173 gnd.n3728 gnd.n3677 0.152939
R13174 gnd.n3729 gnd.n3728 0.152939
R13175 gnd.n3730 gnd.n3729 0.152939
R13176 gnd.n3730 gnd.n3671 0.152939
R13177 gnd.n3737 gnd.n3671 0.152939
R13178 gnd.n794 gnd.n741 0.152939
R13179 gnd.n795 gnd.n794 0.152939
R13180 gnd.n796 gnd.n795 0.152939
R13181 gnd.n797 gnd.n796 0.152939
R13182 gnd.n814 gnd.n797 0.152939
R13183 gnd.n815 gnd.n814 0.152939
R13184 gnd.n816 gnd.n815 0.152939
R13185 gnd.n817 gnd.n816 0.152939
R13186 gnd.n834 gnd.n817 0.152939
R13187 gnd.n835 gnd.n834 0.152939
R13188 gnd.n836 gnd.n835 0.152939
R13189 gnd.n837 gnd.n836 0.152939
R13190 gnd.n854 gnd.n837 0.152939
R13191 gnd.n855 gnd.n854 0.152939
R13192 gnd.n856 gnd.n855 0.152939
R13193 gnd.n857 gnd.n856 0.152939
R13194 gnd.n1013 gnd.n1012 0.152939
R13195 gnd.n1014 gnd.n1013 0.152939
R13196 gnd.n1015 gnd.n1014 0.152939
R13197 gnd.n1016 gnd.n1015 0.152939
R13198 gnd.n1017 gnd.n1016 0.152939
R13199 gnd.n1018 gnd.n1017 0.152939
R13200 gnd.n1019 gnd.n1018 0.152939
R13201 gnd.n1020 gnd.n1019 0.152939
R13202 gnd.n1021 gnd.n1020 0.152939
R13203 gnd.n1022 gnd.n1021 0.152939
R13204 gnd.n1023 gnd.n1022 0.152939
R13205 gnd.n1024 gnd.n1023 0.152939
R13206 gnd.n1025 gnd.n1024 0.152939
R13207 gnd.n1026 gnd.n1025 0.152939
R13208 gnd.n1027 gnd.n1026 0.152939
R13209 gnd.n1028 gnd.n1027 0.152939
R13210 gnd.n1029 gnd.n1028 0.152939
R13211 gnd.n1032 gnd.n1029 0.152939
R13212 gnd.n1033 gnd.n1032 0.152939
R13213 gnd.n1034 gnd.n1033 0.152939
R13214 gnd.n1035 gnd.n1034 0.152939
R13215 gnd.n1036 gnd.n1035 0.152939
R13216 gnd.n1037 gnd.n1036 0.152939
R13217 gnd.n1038 gnd.n1037 0.152939
R13218 gnd.n1039 gnd.n1038 0.152939
R13219 gnd.n1137 gnd.n1136 0.152939
R13220 gnd.n1136 gnd.n1042 0.152939
R13221 gnd.n1043 gnd.n1042 0.152939
R13222 gnd.n1044 gnd.n1043 0.152939
R13223 gnd.n1045 gnd.n1044 0.152939
R13224 gnd.n1046 gnd.n1045 0.152939
R13225 gnd.n1047 gnd.n1046 0.152939
R13226 gnd.n1048 gnd.n1047 0.152939
R13227 gnd.n1116 gnd.n1048 0.152939
R13228 gnd.n1116 gnd.n1115 0.152939
R13229 gnd.n1115 gnd.n1114 0.152939
R13230 gnd.n1114 gnd.n1052 0.152939
R13231 gnd.n1053 gnd.n1052 0.152939
R13232 gnd.n1054 gnd.n1053 0.152939
R13233 gnd.n1055 gnd.n1054 0.152939
R13234 gnd.n1056 gnd.n1055 0.152939
R13235 gnd.n1057 gnd.n1056 0.152939
R13236 gnd.n1058 gnd.n1057 0.152939
R13237 gnd.n1059 gnd.n1058 0.152939
R13238 gnd.n1060 gnd.n1059 0.152939
R13239 gnd.n1061 gnd.n1060 0.152939
R13240 gnd.n1062 gnd.n1061 0.152939
R13241 gnd.n1063 gnd.n1062 0.152939
R13242 gnd.n1064 gnd.n1063 0.152939
R13243 gnd.n1065 gnd.n1064 0.152939
R13244 gnd.n1066 gnd.n1065 0.152939
R13245 gnd.n1067 gnd.n1066 0.152939
R13246 gnd.n1068 gnd.n1067 0.152939
R13247 gnd.n1074 gnd.n1068 0.152939
R13248 gnd.n1074 gnd.n1073 0.152939
R13249 gnd.n3957 gnd.n3746 0.152939
R13250 gnd.n3749 gnd.n3746 0.152939
R13251 gnd.n3750 gnd.n3749 0.152939
R13252 gnd.n3751 gnd.n3750 0.152939
R13253 gnd.n3754 gnd.n3751 0.152939
R13254 gnd.n3755 gnd.n3754 0.152939
R13255 gnd.n3756 gnd.n3755 0.152939
R13256 gnd.n3757 gnd.n3756 0.152939
R13257 gnd.n3760 gnd.n3757 0.152939
R13258 gnd.n3761 gnd.n3760 0.152939
R13259 gnd.n3762 gnd.n3761 0.152939
R13260 gnd.n3763 gnd.n3762 0.152939
R13261 gnd.n3766 gnd.n3763 0.152939
R13262 gnd.n3767 gnd.n3766 0.152939
R13263 gnd.n3768 gnd.n3767 0.152939
R13264 gnd.n3769 gnd.n3768 0.152939
R13265 gnd.n3775 gnd.n3769 0.152939
R13266 gnd.n3776 gnd.n3775 0.152939
R13267 gnd.n3777 gnd.n3776 0.152939
R13268 gnd.n3778 gnd.n3777 0.152939
R13269 gnd.n3781 gnd.n3778 0.152939
R13270 gnd.n3782 gnd.n3781 0.152939
R13271 gnd.n3783 gnd.n3782 0.152939
R13272 gnd.n3784 gnd.n3783 0.152939
R13273 gnd.n3787 gnd.n3784 0.152939
R13274 gnd.n3788 gnd.n3787 0.152939
R13275 gnd.n3789 gnd.n3788 0.152939
R13276 gnd.n3790 gnd.n3789 0.152939
R13277 gnd.n3793 gnd.n3790 0.152939
R13278 gnd.n3794 gnd.n3793 0.152939
R13279 gnd.n3795 gnd.n3794 0.152939
R13280 gnd.n3796 gnd.n3795 0.152939
R13281 gnd.n3799 gnd.n3796 0.152939
R13282 gnd.n3800 gnd.n3799 0.152939
R13283 gnd.n3801 gnd.n3800 0.152939
R13284 gnd.n3802 gnd.n3801 0.152939
R13285 gnd.n3807 gnd.n3802 0.152939
R13286 gnd.n3808 gnd.n3807 0.152939
R13287 gnd.n3809 gnd.n3808 0.152939
R13288 gnd.n3810 gnd.n3809 0.152939
R13289 gnd.n3813 gnd.n3810 0.152939
R13290 gnd.n3814 gnd.n3813 0.152939
R13291 gnd.n3815 gnd.n3814 0.152939
R13292 gnd.n3816 gnd.n3815 0.152939
R13293 gnd.n3819 gnd.n3816 0.152939
R13294 gnd.n3820 gnd.n3819 0.152939
R13295 gnd.n3821 gnd.n3820 0.152939
R13296 gnd.n3822 gnd.n3821 0.152939
R13297 gnd.n3825 gnd.n3822 0.152939
R13298 gnd.n3826 gnd.n3825 0.152939
R13299 gnd.n3827 gnd.n3826 0.152939
R13300 gnd.n3828 gnd.n3827 0.152939
R13301 gnd.n3831 gnd.n3828 0.152939
R13302 gnd.n3832 gnd.n3831 0.152939
R13303 gnd.n3833 gnd.n3832 0.152939
R13304 gnd.n3834 gnd.n3833 0.152939
R13305 gnd.n3838 gnd.n3834 0.152939
R13306 gnd.n3839 gnd.n3838 0.152939
R13307 gnd.n3958 gnd.n2191 0.152939
R13308 gnd.n3982 gnd.n2191 0.152939
R13309 gnd.n3983 gnd.n3982 0.152939
R13310 gnd.n3984 gnd.n3983 0.152939
R13311 gnd.n3985 gnd.n3984 0.152939
R13312 gnd.n3985 gnd.n2166 0.152939
R13313 gnd.n4017 gnd.n2166 0.152939
R13314 gnd.n4018 gnd.n4017 0.152939
R13315 gnd.n4019 gnd.n4018 0.152939
R13316 gnd.n4020 gnd.n4019 0.152939
R13317 gnd.n4020 gnd.n2139 0.152939
R13318 gnd.n4057 gnd.n2139 0.152939
R13319 gnd.n4058 gnd.n4057 0.152939
R13320 gnd.n4060 gnd.n4058 0.152939
R13321 gnd.n4060 gnd.n4059 0.152939
R13322 gnd.n4059 gnd.n741 0.152939
R13323 gnd.n6141 gnd.n563 0.152939
R13324 gnd.n568 gnd.n563 0.152939
R13325 gnd.n569 gnd.n568 0.152939
R13326 gnd.n570 gnd.n569 0.152939
R13327 gnd.n571 gnd.n570 0.152939
R13328 gnd.n576 gnd.n571 0.152939
R13329 gnd.n577 gnd.n576 0.152939
R13330 gnd.n578 gnd.n577 0.152939
R13331 gnd.n579 gnd.n578 0.152939
R13332 gnd.n584 gnd.n579 0.152939
R13333 gnd.n585 gnd.n584 0.152939
R13334 gnd.n586 gnd.n585 0.152939
R13335 gnd.n587 gnd.n586 0.152939
R13336 gnd.n592 gnd.n587 0.152939
R13337 gnd.n593 gnd.n592 0.152939
R13338 gnd.n594 gnd.n593 0.152939
R13339 gnd.n595 gnd.n594 0.152939
R13340 gnd.n600 gnd.n595 0.152939
R13341 gnd.n601 gnd.n600 0.152939
R13342 gnd.n602 gnd.n601 0.152939
R13343 gnd.n603 gnd.n602 0.152939
R13344 gnd.n608 gnd.n603 0.152939
R13345 gnd.n609 gnd.n608 0.152939
R13346 gnd.n610 gnd.n609 0.152939
R13347 gnd.n611 gnd.n610 0.152939
R13348 gnd.n616 gnd.n611 0.152939
R13349 gnd.n617 gnd.n616 0.152939
R13350 gnd.n618 gnd.n617 0.152939
R13351 gnd.n619 gnd.n618 0.152939
R13352 gnd.n624 gnd.n619 0.152939
R13353 gnd.n625 gnd.n624 0.152939
R13354 gnd.n626 gnd.n625 0.152939
R13355 gnd.n627 gnd.n626 0.152939
R13356 gnd.n632 gnd.n627 0.152939
R13357 gnd.n633 gnd.n632 0.152939
R13358 gnd.n634 gnd.n633 0.152939
R13359 gnd.n635 gnd.n634 0.152939
R13360 gnd.n640 gnd.n635 0.152939
R13361 gnd.n641 gnd.n640 0.152939
R13362 gnd.n642 gnd.n641 0.152939
R13363 gnd.n643 gnd.n642 0.152939
R13364 gnd.n648 gnd.n643 0.152939
R13365 gnd.n649 gnd.n648 0.152939
R13366 gnd.n650 gnd.n649 0.152939
R13367 gnd.n651 gnd.n650 0.152939
R13368 gnd.n656 gnd.n651 0.152939
R13369 gnd.n657 gnd.n656 0.152939
R13370 gnd.n658 gnd.n657 0.152939
R13371 gnd.n659 gnd.n658 0.152939
R13372 gnd.n664 gnd.n659 0.152939
R13373 gnd.n665 gnd.n664 0.152939
R13374 gnd.n666 gnd.n665 0.152939
R13375 gnd.n667 gnd.n666 0.152939
R13376 gnd.n672 gnd.n667 0.152939
R13377 gnd.n673 gnd.n672 0.152939
R13378 gnd.n674 gnd.n673 0.152939
R13379 gnd.n675 gnd.n674 0.152939
R13380 gnd.n680 gnd.n675 0.152939
R13381 gnd.n681 gnd.n680 0.152939
R13382 gnd.n682 gnd.n681 0.152939
R13383 gnd.n683 gnd.n682 0.152939
R13384 gnd.n688 gnd.n683 0.152939
R13385 gnd.n689 gnd.n688 0.152939
R13386 gnd.n690 gnd.n689 0.152939
R13387 gnd.n691 gnd.n690 0.152939
R13388 gnd.n696 gnd.n691 0.152939
R13389 gnd.n697 gnd.n696 0.152939
R13390 gnd.n698 gnd.n697 0.152939
R13391 gnd.n699 gnd.n698 0.152939
R13392 gnd.n704 gnd.n699 0.152939
R13393 gnd.n705 gnd.n704 0.152939
R13394 gnd.n706 gnd.n705 0.152939
R13395 gnd.n707 gnd.n706 0.152939
R13396 gnd.n712 gnd.n707 0.152939
R13397 gnd.n713 gnd.n712 0.152939
R13398 gnd.n714 gnd.n713 0.152939
R13399 gnd.n715 gnd.n714 0.152939
R13400 gnd.n720 gnd.n715 0.152939
R13401 gnd.n721 gnd.n720 0.152939
R13402 gnd.n722 gnd.n721 0.152939
R13403 gnd.n723 gnd.n722 0.152939
R13404 gnd.n728 gnd.n723 0.152939
R13405 gnd.n729 gnd.n728 0.152939
R13406 gnd.n5971 gnd.n729 0.152939
R13407 gnd.n4301 gnd.n4300 0.152939
R13408 gnd.n4301 gnd.n2072 0.152939
R13409 gnd.n4315 gnd.n2072 0.152939
R13410 gnd.n4316 gnd.n4315 0.152939
R13411 gnd.n4317 gnd.n4316 0.152939
R13412 gnd.n4317 gnd.n2058 0.152939
R13413 gnd.n4331 gnd.n2058 0.152939
R13414 gnd.n4332 gnd.n4331 0.152939
R13415 gnd.n4333 gnd.n4332 0.152939
R13416 gnd.n4333 gnd.n2044 0.152939
R13417 gnd.n4347 gnd.n2044 0.152939
R13418 gnd.n4348 gnd.n4347 0.152939
R13419 gnd.n4349 gnd.n4348 0.152939
R13420 gnd.n4349 gnd.n2030 0.152939
R13421 gnd.n4363 gnd.n2030 0.152939
R13422 gnd.n4364 gnd.n4363 0.152939
R13423 gnd.n4365 gnd.n4364 0.152939
R13424 gnd.n4365 gnd.n2015 0.152939
R13425 gnd.n4379 gnd.n2015 0.152939
R13426 gnd.n4380 gnd.n4379 0.152939
R13427 gnd.n4381 gnd.n4380 0.152939
R13428 gnd.n4381 gnd.n2002 0.152939
R13429 gnd.n4395 gnd.n2002 0.152939
R13430 gnd.n4396 gnd.n4395 0.152939
R13431 gnd.n4398 gnd.n4396 0.152939
R13432 gnd.n4398 gnd.n4397 0.152939
R13433 gnd.n4397 gnd.n1986 0.152939
R13434 gnd.n4419 gnd.n1986 0.152939
R13435 gnd.n4420 gnd.n4419 0.152939
R13436 gnd.n4422 gnd.n4420 0.152939
R13437 gnd.n4422 gnd.n4421 0.152939
R13438 gnd.n4421 gnd.n1219 0.152939
R13439 gnd.n5668 gnd.n1219 0.152939
R13440 gnd.n5668 gnd.n5667 0.152939
R13441 gnd.n5667 gnd.n5666 0.152939
R13442 gnd.n5666 gnd.n1220 0.152939
R13443 gnd.n5662 gnd.n1220 0.152939
R13444 gnd.n5662 gnd.n5661 0.152939
R13445 gnd.n5661 gnd.n5660 0.152939
R13446 gnd.n5660 gnd.n1225 0.152939
R13447 gnd.n5656 gnd.n1225 0.152939
R13448 gnd.n5656 gnd.n5655 0.152939
R13449 gnd.n5655 gnd.n5654 0.152939
R13450 gnd.n5654 gnd.n1230 0.152939
R13451 gnd.n5650 gnd.n1230 0.152939
R13452 gnd.n5650 gnd.n5649 0.152939
R13453 gnd.n5649 gnd.n5648 0.152939
R13454 gnd.n5648 gnd.n1235 0.152939
R13455 gnd.n5644 gnd.n1235 0.152939
R13456 gnd.n5644 gnd.n5643 0.152939
R13457 gnd.n5643 gnd.n5642 0.152939
R13458 gnd.n5642 gnd.n1240 0.152939
R13459 gnd.n5638 gnd.n1240 0.152939
R13460 gnd.n5638 gnd.n5637 0.152939
R13461 gnd.n5637 gnd.n5636 0.152939
R13462 gnd.n5636 gnd.n1245 0.152939
R13463 gnd.n5632 gnd.n1245 0.152939
R13464 gnd.n5632 gnd.n5631 0.152939
R13465 gnd.n5631 gnd.n5630 0.152939
R13466 gnd.n5630 gnd.n1250 0.152939
R13467 gnd.n5626 gnd.n1250 0.152939
R13468 gnd.n5626 gnd.n5625 0.152939
R13469 gnd.n5625 gnd.n5624 0.152939
R13470 gnd.n5624 gnd.n1255 0.152939
R13471 gnd.n5620 gnd.n1255 0.152939
R13472 gnd.n5620 gnd.n5619 0.152939
R13473 gnd.n5619 gnd.n5618 0.152939
R13474 gnd.n5618 gnd.n1260 0.152939
R13475 gnd.n5614 gnd.n1260 0.152939
R13476 gnd.n5614 gnd.n5613 0.152939
R13477 gnd.n5613 gnd.n5612 0.152939
R13478 gnd.n5612 gnd.n1265 0.152939
R13479 gnd.n5608 gnd.n1265 0.152939
R13480 gnd.n5608 gnd.n5607 0.152939
R13481 gnd.n5607 gnd.n5606 0.152939
R13482 gnd.n5606 gnd.n1270 0.152939
R13483 gnd.n5602 gnd.n1270 0.152939
R13484 gnd.n5602 gnd.n5601 0.152939
R13485 gnd.n5601 gnd.n5600 0.152939
R13486 gnd.n5600 gnd.n1275 0.152939
R13487 gnd.n5596 gnd.n1275 0.152939
R13488 gnd.n5596 gnd.n5595 0.152939
R13489 gnd.n5595 gnd.n5594 0.152939
R13490 gnd.n5594 gnd.n1280 0.152939
R13491 gnd.n5590 gnd.n1280 0.152939
R13492 gnd.n5590 gnd.n5589 0.152939
R13493 gnd.n5589 gnd.n5588 0.152939
R13494 gnd.n5588 gnd.n1285 0.152939
R13495 gnd.n5584 gnd.n1285 0.152939
R13496 gnd.n5584 gnd.n5583 0.152939
R13497 gnd.n5583 gnd.n5582 0.152939
R13498 gnd.n5582 gnd.n1290 0.152939
R13499 gnd.n5578 gnd.n1290 0.152939
R13500 gnd.n5578 gnd.n5577 0.152939
R13501 gnd.n5577 gnd.n5576 0.152939
R13502 gnd.n5576 gnd.n1295 0.152939
R13503 gnd.n5572 gnd.n1295 0.152939
R13504 gnd.n5572 gnd.n5571 0.152939
R13505 gnd.n5571 gnd.n5570 0.152939
R13506 gnd.n5570 gnd.n1300 0.152939
R13507 gnd.n1303 gnd.n1300 0.152939
R13508 gnd.n4114 gnd.n2122 0.152939
R13509 gnd.n4114 gnd.n4113 0.152939
R13510 gnd.n4113 gnd.n4112 0.152939
R13511 gnd.n4112 gnd.n2110 0.152939
R13512 gnd.n4156 gnd.n2110 0.152939
R13513 gnd.n4157 gnd.n4156 0.152939
R13514 gnd.n4158 gnd.n4157 0.152939
R13515 gnd.n4158 gnd.n2104 0.152939
R13516 gnd.n4170 gnd.n2104 0.152939
R13517 gnd.n4171 gnd.n4170 0.152939
R13518 gnd.n4172 gnd.n4171 0.152939
R13519 gnd.n4172 gnd.n2098 0.152939
R13520 gnd.n4196 gnd.n2098 0.152939
R13521 gnd.n4196 gnd.n4195 0.152939
R13522 gnd.n4195 gnd.n4194 0.152939
R13523 gnd.n4194 gnd.n2099 0.152939
R13524 gnd.n4190 gnd.n2099 0.152939
R13525 gnd.n4190 gnd.n870 0.152939
R13526 gnd.n5875 gnd.n870 0.152939
R13527 gnd.n5875 gnd.n5874 0.152939
R13528 gnd.n5862 gnd.n894 0.152939
R13529 gnd.n5862 gnd.n5861 0.152939
R13530 gnd.n5861 gnd.n5860 0.152939
R13531 gnd.n5860 gnd.n896 0.152939
R13532 gnd.n5856 gnd.n896 0.152939
R13533 gnd.n5856 gnd.n5855 0.152939
R13534 gnd.n4296 gnd.n4232 0.152939
R13535 gnd.n4296 gnd.n4295 0.152939
R13536 gnd.n4295 gnd.n4294 0.152939
R13537 gnd.n4294 gnd.n4233 0.152939
R13538 gnd.n4290 gnd.n4233 0.152939
R13539 gnd.n4290 gnd.n4289 0.152939
R13540 gnd.n4289 gnd.n4288 0.152939
R13541 gnd.n4288 gnd.n4237 0.152939
R13542 gnd.n4284 gnd.n4237 0.152939
R13543 gnd.n4284 gnd.n4283 0.152939
R13544 gnd.n4283 gnd.n4282 0.152939
R13545 gnd.n4282 gnd.n4241 0.152939
R13546 gnd.n4278 gnd.n4241 0.152939
R13547 gnd.n4278 gnd.n4277 0.152939
R13548 gnd.n4277 gnd.n4276 0.152939
R13549 gnd.n4276 gnd.n4245 0.152939
R13550 gnd.n4272 gnd.n4245 0.152939
R13551 gnd.n4272 gnd.n4271 0.152939
R13552 gnd.n4271 gnd.n4270 0.152939
R13553 gnd.n4270 gnd.n4249 0.152939
R13554 gnd.n4266 gnd.n4249 0.152939
R13555 gnd.n4266 gnd.n4265 0.152939
R13556 gnd.n4265 gnd.n4264 0.152939
R13557 gnd.n4264 gnd.n4253 0.152939
R13558 gnd.n4260 gnd.n4253 0.152939
R13559 gnd.n4260 gnd.n4259 0.152939
R13560 gnd.n4259 gnd.n4258 0.152939
R13561 gnd.n4258 gnd.n1980 0.152939
R13562 gnd.n4429 gnd.n1980 0.152939
R13563 gnd.n4430 gnd.n4429 0.152939
R13564 gnd.n4431 gnd.n4430 0.152939
R13565 gnd.n4431 gnd.n1978 0.152939
R13566 gnd.n4534 gnd.n1978 0.152939
R13567 gnd.n4535 gnd.n4534 0.152939
R13568 gnd.n4548 gnd.n4535 0.152939
R13569 gnd.n4548 gnd.n4547 0.152939
R13570 gnd.n4547 gnd.n4546 0.152939
R13571 gnd.n4546 gnd.n4536 0.152939
R13572 gnd.n4542 gnd.n4536 0.152939
R13573 gnd.n4542 gnd.n4541 0.152939
R13574 gnd.n4541 gnd.n1929 0.152939
R13575 gnd.n4615 gnd.n1929 0.152939
R13576 gnd.n4616 gnd.n4615 0.152939
R13577 gnd.n4651 gnd.n4616 0.152939
R13578 gnd.n4651 gnd.n4650 0.152939
R13579 gnd.n4650 gnd.n4649 0.152939
R13580 gnd.n4649 gnd.n4617 0.152939
R13581 gnd.n4645 gnd.n4617 0.152939
R13582 gnd.n4645 gnd.n4644 0.152939
R13583 gnd.n4644 gnd.n4643 0.152939
R13584 gnd.n4643 gnd.n4621 0.152939
R13585 gnd.n4639 gnd.n4621 0.152939
R13586 gnd.n4639 gnd.n4638 0.152939
R13587 gnd.n4638 gnd.n4637 0.152939
R13588 gnd.n4637 gnd.n4626 0.152939
R13589 gnd.n4633 gnd.n4626 0.152939
R13590 gnd.n4633 gnd.n4632 0.152939
R13591 gnd.n4632 gnd.n1849 0.152939
R13592 gnd.n4782 gnd.n1849 0.152939
R13593 gnd.n4783 gnd.n4782 0.152939
R13594 gnd.n4809 gnd.n4783 0.152939
R13595 gnd.n4809 gnd.n4808 0.152939
R13596 gnd.n4808 gnd.n4807 0.152939
R13597 gnd.n4807 gnd.n4784 0.152939
R13598 gnd.n4803 gnd.n4784 0.152939
R13599 gnd.n4803 gnd.n4802 0.152939
R13600 gnd.n4802 gnd.n4801 0.152939
R13601 gnd.n4801 gnd.n4789 0.152939
R13602 gnd.n4797 gnd.n4789 0.152939
R13603 gnd.n4797 gnd.n4796 0.152939
R13604 gnd.n4796 gnd.n4795 0.152939
R13605 gnd.n4795 gnd.n1747 0.152939
R13606 gnd.n5043 gnd.n1747 0.152939
R13607 gnd.n5044 gnd.n5043 0.152939
R13608 gnd.n5045 gnd.n5044 0.152939
R13609 gnd.n5045 gnd.n1734 0.152939
R13610 gnd.n5059 gnd.n1734 0.152939
R13611 gnd.n5060 gnd.n5059 0.152939
R13612 gnd.n5061 gnd.n5060 0.152939
R13613 gnd.n5061 gnd.n1722 0.152939
R13614 gnd.n5076 gnd.n1722 0.152939
R13615 gnd.n5077 gnd.n5076 0.152939
R13616 gnd.n5078 gnd.n5077 0.152939
R13617 gnd.n5078 gnd.n1709 0.152939
R13618 gnd.n5092 gnd.n1709 0.152939
R13619 gnd.n5093 gnd.n5092 0.152939
R13620 gnd.n5094 gnd.n5093 0.152939
R13621 gnd.n5094 gnd.n1696 0.152939
R13622 gnd.n5108 gnd.n1696 0.152939
R13623 gnd.n5109 gnd.n5108 0.152939
R13624 gnd.n5110 gnd.n5109 0.152939
R13625 gnd.n5110 gnd.n1681 0.152939
R13626 gnd.n5124 gnd.n1681 0.152939
R13627 gnd.n5125 gnd.n5124 0.152939
R13628 gnd.n5126 gnd.n5125 0.152939
R13629 gnd.n5126 gnd.n1670 0.152939
R13630 gnd.n5143 gnd.n1670 0.152939
R13631 gnd.n5144 gnd.n5143 0.152939
R13632 gnd.n5145 gnd.n5144 0.152939
R13633 gnd.n5145 gnd.n1311 0.152939
R13634 gnd.n5562 gnd.n1311 0.152939
R13635 gnd.n5561 gnd.n1312 0.152939
R13636 gnd.n5557 gnd.n1312 0.152939
R13637 gnd.n5557 gnd.n5556 0.152939
R13638 gnd.n5556 gnd.n5555 0.152939
R13639 gnd.n5555 gnd.n1316 0.152939
R13640 gnd.n5551 gnd.n1316 0.152939
R13641 gnd.n5215 gnd.n5177 0.152939
R13642 gnd.n5215 gnd.n5214 0.152939
R13643 gnd.n5214 gnd.n5213 0.152939
R13644 gnd.n5213 gnd.n5178 0.152939
R13645 gnd.n5209 gnd.n5178 0.152939
R13646 gnd.n5209 gnd.n5208 0.152939
R13647 gnd.n5208 gnd.n5207 0.152939
R13648 gnd.n5207 gnd.n5183 0.152939
R13649 gnd.n5203 gnd.n5183 0.152939
R13650 gnd.n5203 gnd.n1613 0.152939
R13651 gnd.n5264 gnd.n1613 0.152939
R13652 gnd.n5265 gnd.n5264 0.152939
R13653 gnd.n5266 gnd.n5265 0.152939
R13654 gnd.n5266 gnd.n1608 0.152939
R13655 gnd.n5279 gnd.n1608 0.152939
R13656 gnd.n5280 gnd.n5279 0.152939
R13657 gnd.n5285 gnd.n5280 0.152939
R13658 gnd.n5285 gnd.n5284 0.152939
R13659 gnd.n5284 gnd.n5283 0.152939
R13660 gnd.n5283 gnd.n67 0.152939
R13661 gnd.n7208 gnd.n7207 0.145814
R13662 gnd.n4095 gnd.n4094 0.145814
R13663 gnd.n4095 gnd.n2122 0.145814
R13664 gnd.n7208 gnd.n67 0.145814
R13665 gnd.n5855 gnd.n5854 0.128549
R13666 gnd.n5551 gnd.n5550 0.128549
R13667 gnd.n2484 gnd.n0 0.127478
R13668 gnd.n4128 gnd.n730 0.0919634
R13669 gnd.n5246 gnd.n83 0.0919634
R13670 gnd.n3064 gnd.n3063 0.0767195
R13671 gnd.n3063 gnd.n3062 0.0767195
R13672 gnd.n5854 gnd.n865 0.063
R13673 gnd.n5550 gnd.n1321 0.063
R13674 gnd.n184 gnd.n83 0.0614756
R13675 gnd.n5970 gnd.n730 0.0614756
R13676 gnd.n1489 gnd.n1321 0.0538288
R13677 gnd.n7144 gnd.n173 0.0538288
R13678 gnd.n3964 gnd.n2203 0.0538288
R13679 gnd.n5882 gnd.n865 0.0538288
R13680 gnd.n3630 gnd.n2246 0.0477147
R13681 gnd.n2827 gnd.n2715 0.0442063
R13682 gnd.n2828 gnd.n2827 0.0442063
R13683 gnd.n2829 gnd.n2828 0.0442063
R13684 gnd.n2829 gnd.n2704 0.0442063
R13685 gnd.n2843 gnd.n2704 0.0442063
R13686 gnd.n2844 gnd.n2843 0.0442063
R13687 gnd.n2845 gnd.n2844 0.0442063
R13688 gnd.n2845 gnd.n2691 0.0442063
R13689 gnd.n2889 gnd.n2691 0.0442063
R13690 gnd.n2890 gnd.n2889 0.0442063
R13691 gnd.n2892 gnd.n2625 0.0344674
R13692 gnd.n5372 gnd.n1489 0.0344674
R13693 gnd.n5372 gnd.n1491 0.0344674
R13694 gnd.n1515 gnd.n1491 0.0344674
R13695 gnd.n1516 gnd.n1515 0.0344674
R13696 gnd.n1517 gnd.n1516 0.0344674
R13697 gnd.n1518 gnd.n1517 0.0344674
R13698 gnd.n5190 gnd.n1518 0.0344674
R13699 gnd.n5190 gnd.n1536 0.0344674
R13700 gnd.n1537 gnd.n1536 0.0344674
R13701 gnd.n1538 gnd.n1537 0.0344674
R13702 gnd.n5196 gnd.n1538 0.0344674
R13703 gnd.n5196 gnd.n1556 0.0344674
R13704 gnd.n1557 gnd.n1556 0.0344674
R13705 gnd.n1558 gnd.n1557 0.0344674
R13706 gnd.n5273 gnd.n1558 0.0344674
R13707 gnd.n5273 gnd.n1573 0.0344674
R13708 gnd.n1574 gnd.n1573 0.0344674
R13709 gnd.n1575 gnd.n1574 0.0344674
R13710 gnd.n5293 gnd.n1575 0.0344674
R13711 gnd.n5294 gnd.n5293 0.0344674
R13712 gnd.n5294 gnd.n1600 0.0344674
R13713 gnd.n5303 gnd.n1600 0.0344674
R13714 gnd.n5303 gnd.n179 0.0344674
R13715 gnd.n6787 gnd.n179 0.0344674
R13716 gnd.n6788 gnd.n6787 0.0344674
R13717 gnd.n6788 gnd.n97 0.0344674
R13718 gnd.n98 gnd.n97 0.0344674
R13719 gnd.n99 gnd.n98 0.0344674
R13720 gnd.n7120 gnd.n99 0.0344674
R13721 gnd.n7120 gnd.n115 0.0344674
R13722 gnd.n116 gnd.n115 0.0344674
R13723 gnd.n117 gnd.n116 0.0344674
R13724 gnd.n7127 gnd.n117 0.0344674
R13725 gnd.n7127 gnd.n135 0.0344674
R13726 gnd.n136 gnd.n135 0.0344674
R13727 gnd.n137 gnd.n136 0.0344674
R13728 gnd.n7134 gnd.n137 0.0344674
R13729 gnd.n7134 gnd.n154 0.0344674
R13730 gnd.n155 gnd.n154 0.0344674
R13731 gnd.n156 gnd.n155 0.0344674
R13732 gnd.n172 gnd.n156 0.0344674
R13733 gnd.n7144 gnd.n172 0.0344674
R13734 gnd.n3965 gnd.n3964 0.0344674
R13735 gnd.n3965 gnd.n2199 0.0344674
R13736 gnd.n2200 gnd.n2199 0.0344674
R13737 gnd.n3971 gnd.n2200 0.0344674
R13738 gnd.n3972 gnd.n3971 0.0344674
R13739 gnd.n3972 gnd.n2177 0.0344674
R13740 gnd.n2177 gnd.n2174 0.0344674
R13741 gnd.n2175 gnd.n2174 0.0344674
R13742 gnd.n4006 gnd.n2175 0.0344674
R13743 gnd.n4007 gnd.n4006 0.0344674
R13744 gnd.n4007 gnd.n2152 0.0344674
R13745 gnd.n2152 gnd.n2148 0.0344674
R13746 gnd.n2149 gnd.n2148 0.0344674
R13747 gnd.n2150 gnd.n2149 0.0344674
R13748 gnd.n4045 gnd.n2150 0.0344674
R13749 gnd.n4046 gnd.n4045 0.0344674
R13750 gnd.n4046 gnd.n2129 0.0344674
R13751 gnd.n2129 gnd.n751 0.0344674
R13752 gnd.n752 gnd.n751 0.0344674
R13753 gnd.n753 gnd.n752 0.0344674
R13754 gnd.n2124 gnd.n753 0.0344674
R13755 gnd.n2124 gnd.n767 0.0344674
R13756 gnd.n768 gnd.n767 0.0344674
R13757 gnd.n769 gnd.n768 0.0344674
R13758 gnd.n4104 gnd.n769 0.0344674
R13759 gnd.n4104 gnd.n785 0.0344674
R13760 gnd.n786 gnd.n785 0.0344674
R13761 gnd.n787 gnd.n786 0.0344674
R13762 gnd.n2108 gnd.n787 0.0344674
R13763 gnd.n2108 gnd.n804 0.0344674
R13764 gnd.n805 gnd.n804 0.0344674
R13765 gnd.n806 gnd.n805 0.0344674
R13766 gnd.n2102 gnd.n806 0.0344674
R13767 gnd.n2102 gnd.n825 0.0344674
R13768 gnd.n826 gnd.n825 0.0344674
R13769 gnd.n827 gnd.n826 0.0344674
R13770 gnd.n4181 gnd.n827 0.0344674
R13771 gnd.n4181 gnd.n845 0.0344674
R13772 gnd.n846 gnd.n845 0.0344674
R13773 gnd.n847 gnd.n846 0.0344674
R13774 gnd.n864 gnd.n847 0.0344674
R13775 gnd.n5882 gnd.n864 0.0344674
R13776 gnd.n5853 gnd.n901 0.0343753
R13777 gnd.n5549 gnd.n5548 0.0343753
R13778 gnd.n5873 gnd.n5872 0.0296328
R13779 gnd.n5176 gnd.n5175 0.0296328
R13780 gnd.n2912 gnd.n2911 0.0269946
R13781 gnd.n2914 gnd.n2913 0.0269946
R13782 gnd.n2620 gnd.n2618 0.0269946
R13783 gnd.n2924 gnd.n2922 0.0269946
R13784 gnd.n2923 gnd.n2599 0.0269946
R13785 gnd.n2943 gnd.n2942 0.0269946
R13786 gnd.n2945 gnd.n2944 0.0269946
R13787 gnd.n2594 gnd.n2593 0.0269946
R13788 gnd.n2955 gnd.n2589 0.0269946
R13789 gnd.n2954 gnd.n2591 0.0269946
R13790 gnd.n2590 gnd.n2572 0.0269946
R13791 gnd.n2975 gnd.n2573 0.0269946
R13792 gnd.n2974 gnd.n2574 0.0269946
R13793 gnd.n3008 gnd.n2549 0.0269946
R13794 gnd.n3010 gnd.n3009 0.0269946
R13795 gnd.n3011 gnd.n2496 0.0269946
R13796 gnd.n2544 gnd.n2497 0.0269946
R13797 gnd.n2546 gnd.n2498 0.0269946
R13798 gnd.n3021 gnd.n3020 0.0269946
R13799 gnd.n3023 gnd.n3022 0.0269946
R13800 gnd.n3024 gnd.n2518 0.0269946
R13801 gnd.n3026 gnd.n2519 0.0269946
R13802 gnd.n3029 gnd.n2520 0.0269946
R13803 gnd.n3032 gnd.n3031 0.0269946
R13804 gnd.n3034 gnd.n3033 0.0269946
R13805 gnd.n3099 gnd.n2419 0.0269946
R13806 gnd.n3101 gnd.n3100 0.0269946
R13807 gnd.n3110 gnd.n2412 0.0269946
R13808 gnd.n3112 gnd.n3111 0.0269946
R13809 gnd.n3113 gnd.n2410 0.0269946
R13810 gnd.n3120 gnd.n3116 0.0269946
R13811 gnd.n3119 gnd.n3118 0.0269946
R13812 gnd.n3117 gnd.n2389 0.0269946
R13813 gnd.n3142 gnd.n2390 0.0269946
R13814 gnd.n3141 gnd.n2391 0.0269946
R13815 gnd.n3184 gnd.n2364 0.0269946
R13816 gnd.n3186 gnd.n3185 0.0269946
R13817 gnd.n3195 gnd.n2357 0.0269946
R13818 gnd.n3197 gnd.n3196 0.0269946
R13819 gnd.n3198 gnd.n2355 0.0269946
R13820 gnd.n3205 gnd.n3201 0.0269946
R13821 gnd.n3204 gnd.n3203 0.0269946
R13822 gnd.n3202 gnd.n2334 0.0269946
R13823 gnd.n3227 gnd.n2335 0.0269946
R13824 gnd.n3226 gnd.n2336 0.0269946
R13825 gnd.n3273 gnd.n2310 0.0269946
R13826 gnd.n3275 gnd.n3274 0.0269946
R13827 gnd.n3284 gnd.n2303 0.0269946
R13828 gnd.n3543 gnd.n2301 0.0269946
R13829 gnd.n3548 gnd.n3546 0.0269946
R13830 gnd.n3547 gnd.n2282 0.0269946
R13831 gnd.n3572 gnd.n3571 0.0269946
R13832 gnd.n5849 gnd.n907 0.022519
R13833 gnd.n5848 gnd.n908 0.022519
R13834 gnd.n5845 gnd.n5844 0.022519
R13835 gnd.n5841 gnd.n913 0.022519
R13836 gnd.n5840 gnd.n919 0.022519
R13837 gnd.n5837 gnd.n5836 0.022519
R13838 gnd.n5833 gnd.n923 0.022519
R13839 gnd.n5832 gnd.n927 0.022519
R13840 gnd.n5829 gnd.n5828 0.022519
R13841 gnd.n5825 gnd.n931 0.022519
R13842 gnd.n5824 gnd.n937 0.022519
R13843 gnd.n5821 gnd.n5820 0.022519
R13844 gnd.n5817 gnd.n941 0.022519
R13845 gnd.n5816 gnd.n945 0.022519
R13846 gnd.n5813 gnd.n5812 0.022519
R13847 gnd.n5809 gnd.n949 0.022519
R13848 gnd.n5808 gnd.n958 0.022519
R13849 gnd.n963 gnd.n962 0.022519
R13850 gnd.n5872 gnd.n872 0.022519
R13851 gnd.n5545 gnd.n1322 0.022519
R13852 gnd.n5544 gnd.n1326 0.022519
R13853 gnd.n5541 gnd.n5540 0.022519
R13854 gnd.n5537 gnd.n1331 0.022519
R13855 gnd.n5536 gnd.n1335 0.022519
R13856 gnd.n5533 gnd.n5532 0.022519
R13857 gnd.n5529 gnd.n1339 0.022519
R13858 gnd.n5528 gnd.n1343 0.022519
R13859 gnd.n5525 gnd.n5524 0.022519
R13860 gnd.n5521 gnd.n1347 0.022519
R13861 gnd.n5520 gnd.n1351 0.022519
R13862 gnd.n5517 gnd.n5516 0.022519
R13863 gnd.n5513 gnd.n1355 0.022519
R13864 gnd.n5512 gnd.n1359 0.022519
R13865 gnd.n5509 gnd.n5508 0.022519
R13866 gnd.n5505 gnd.n1363 0.022519
R13867 gnd.n5504 gnd.n1369 0.022519
R13868 gnd.n1634 gnd.n1372 0.022519
R13869 gnd.n5175 gnd.n1633 0.022519
R13870 gnd.n5176 gnd.n1632 0.0218415
R13871 gnd.n5873 gnd.n871 0.0218415
R13872 gnd.n2892 gnd.n2891 0.0202011
R13873 gnd.n2891 gnd.n2890 0.0148637
R13874 gnd.n3541 gnd.n3285 0.0144266
R13875 gnd.n3542 gnd.n3541 0.0130679
R13876 gnd.n907 gnd.n901 0.0123564
R13877 gnd.n5849 gnd.n5848 0.0123564
R13878 gnd.n5845 gnd.n908 0.0123564
R13879 gnd.n5844 gnd.n913 0.0123564
R13880 gnd.n5841 gnd.n5840 0.0123564
R13881 gnd.n5837 gnd.n919 0.0123564
R13882 gnd.n5836 gnd.n923 0.0123564
R13883 gnd.n5833 gnd.n5832 0.0123564
R13884 gnd.n5829 gnd.n927 0.0123564
R13885 gnd.n5828 gnd.n931 0.0123564
R13886 gnd.n5825 gnd.n5824 0.0123564
R13887 gnd.n5821 gnd.n937 0.0123564
R13888 gnd.n5820 gnd.n941 0.0123564
R13889 gnd.n5817 gnd.n5816 0.0123564
R13890 gnd.n5813 gnd.n945 0.0123564
R13891 gnd.n5812 gnd.n949 0.0123564
R13892 gnd.n5809 gnd.n5808 0.0123564
R13893 gnd.n963 gnd.n958 0.0123564
R13894 gnd.n962 gnd.n872 0.0123564
R13895 gnd.n5548 gnd.n1322 0.0123564
R13896 gnd.n5545 gnd.n5544 0.0123564
R13897 gnd.n5541 gnd.n1326 0.0123564
R13898 gnd.n5540 gnd.n1331 0.0123564
R13899 gnd.n5537 gnd.n5536 0.0123564
R13900 gnd.n5533 gnd.n1335 0.0123564
R13901 gnd.n5532 gnd.n1339 0.0123564
R13902 gnd.n5529 gnd.n5528 0.0123564
R13903 gnd.n5525 gnd.n1343 0.0123564
R13904 gnd.n5524 gnd.n1347 0.0123564
R13905 gnd.n5521 gnd.n5520 0.0123564
R13906 gnd.n5517 gnd.n1351 0.0123564
R13907 gnd.n5516 gnd.n1355 0.0123564
R13908 gnd.n5513 gnd.n5512 0.0123564
R13909 gnd.n5509 gnd.n1359 0.0123564
R13910 gnd.n5508 gnd.n1363 0.0123564
R13911 gnd.n5505 gnd.n5504 0.0123564
R13912 gnd.n1372 gnd.n1369 0.0123564
R13913 gnd.n1634 gnd.n1633 0.0123564
R13914 gnd.n2911 gnd.n2625 0.00797283
R13915 gnd.n2913 gnd.n2912 0.00797283
R13916 gnd.n2914 gnd.n2620 0.00797283
R13917 gnd.n2922 gnd.n2618 0.00797283
R13918 gnd.n2924 gnd.n2923 0.00797283
R13919 gnd.n2942 gnd.n2599 0.00797283
R13920 gnd.n2944 gnd.n2943 0.00797283
R13921 gnd.n2945 gnd.n2594 0.00797283
R13922 gnd.n2593 gnd.n2589 0.00797283
R13923 gnd.n2955 gnd.n2954 0.00797283
R13924 gnd.n2591 gnd.n2590 0.00797283
R13925 gnd.n2573 gnd.n2572 0.00797283
R13926 gnd.n2975 gnd.n2974 0.00797283
R13927 gnd.n2574 gnd.n2549 0.00797283
R13928 gnd.n3009 gnd.n3008 0.00797283
R13929 gnd.n3011 gnd.n3010 0.00797283
R13930 gnd.n2544 gnd.n2496 0.00797283
R13931 gnd.n2546 gnd.n2497 0.00797283
R13932 gnd.n3020 gnd.n2498 0.00797283
R13933 gnd.n3022 gnd.n3021 0.00797283
R13934 gnd.n3024 gnd.n3023 0.00797283
R13935 gnd.n3026 gnd.n2518 0.00797283
R13936 gnd.n3029 gnd.n2519 0.00797283
R13937 gnd.n3031 gnd.n2520 0.00797283
R13938 gnd.n3034 gnd.n3032 0.00797283
R13939 gnd.n3033 gnd.n2419 0.00797283
R13940 gnd.n3101 gnd.n3099 0.00797283
R13941 gnd.n3100 gnd.n2412 0.00797283
R13942 gnd.n3111 gnd.n3110 0.00797283
R13943 gnd.n3113 gnd.n3112 0.00797283
R13944 gnd.n3116 gnd.n2410 0.00797283
R13945 gnd.n3120 gnd.n3119 0.00797283
R13946 gnd.n3118 gnd.n3117 0.00797283
R13947 gnd.n2390 gnd.n2389 0.00797283
R13948 gnd.n3142 gnd.n3141 0.00797283
R13949 gnd.n2391 gnd.n2364 0.00797283
R13950 gnd.n3186 gnd.n3184 0.00797283
R13951 gnd.n3185 gnd.n2357 0.00797283
R13952 gnd.n3196 gnd.n3195 0.00797283
R13953 gnd.n3198 gnd.n3197 0.00797283
R13954 gnd.n3201 gnd.n2355 0.00797283
R13955 gnd.n3205 gnd.n3204 0.00797283
R13956 gnd.n3203 gnd.n3202 0.00797283
R13957 gnd.n2335 gnd.n2334 0.00797283
R13958 gnd.n3227 gnd.n3226 0.00797283
R13959 gnd.n2336 gnd.n2310 0.00797283
R13960 gnd.n3275 gnd.n3273 0.00797283
R13961 gnd.n3274 gnd.n2303 0.00797283
R13962 gnd.n3285 gnd.n3284 0.00797283
R13963 gnd.n3543 gnd.n3542 0.00797283
R13964 gnd.n3546 gnd.n2301 0.00797283
R13965 gnd.n3548 gnd.n3547 0.00797283
R13966 gnd.n3571 gnd.n2282 0.00797283
R13967 gnd.n3572 gnd.n2246 0.00797283
R13968 gnd.n5854 gnd.n5853 0.00592005
R13969 gnd.n5550 gnd.n5549 0.00592005
R13970 a_n7636_8799.n219 a_n7636_8799.t56 485.149
R13971 a_n7636_8799.n238 a_n7636_8799.t68 485.149
R13972 a_n7636_8799.n258 a_n7636_8799.t105 485.149
R13973 a_n7636_8799.n158 a_n7636_8799.t127 485.149
R13974 a_n7636_8799.n177 a_n7636_8799.t142 485.149
R13975 a_n7636_8799.n197 a_n7636_8799.t104 485.149
R13976 a_n7636_8799.n53 a_n7636_8799.t78 485.135
R13977 a_n7636_8799.n231 a_n7636_8799.t77 464.166
R13978 a_n7636_8799.n213 a_n7636_8799.t50 464.166
R13979 a_n7636_8799.n230 a_n7636_8799.t126 464.166
R13980 a_n7636_8799.n229 a_n7636_8799.t81 464.166
R13981 a_n7636_8799.n214 a_n7636_8799.t57 464.166
R13982 a_n7636_8799.n228 a_n7636_8799.t132 464.166
R13983 a_n7636_8799.n227 a_n7636_8799.t98 464.166
R13984 a_n7636_8799.n215 a_n7636_8799.t96 464.166
R13985 a_n7636_8799.n226 a_n7636_8799.t31 464.166
R13986 a_n7636_8799.n225 a_n7636_8799.t102 464.166
R13987 a_n7636_8799.n216 a_n7636_8799.t101 464.166
R13988 a_n7636_8799.n224 a_n7636_8799.t33 464.166
R13989 a_n7636_8799.n223 a_n7636_8799.t32 464.166
R13990 a_n7636_8799.n217 a_n7636_8799.t118 464.166
R13991 a_n7636_8799.n222 a_n7636_8799.t52 464.166
R13992 a_n7636_8799.n221 a_n7636_8799.t36 464.166
R13993 a_n7636_8799.n218 a_n7636_8799.t122 464.166
R13994 a_n7636_8799.n220 a_n7636_8799.t80 464.166
R13995 a_n7636_8799.n68 a_n7636_8799.t88 485.135
R13996 a_n7636_8799.n250 a_n7636_8799.t87 464.166
R13997 a_n7636_8799.n232 a_n7636_8799.t65 464.166
R13998 a_n7636_8799.n249 a_n7636_8799.t141 464.166
R13999 a_n7636_8799.n248 a_n7636_8799.t94 464.166
R14000 a_n7636_8799.n233 a_n7636_8799.t67 464.166
R14001 a_n7636_8799.n247 a_n7636_8799.t147 464.166
R14002 a_n7636_8799.n246 a_n7636_8799.t111 464.166
R14003 a_n7636_8799.n234 a_n7636_8799.t110 464.166
R14004 a_n7636_8799.n245 a_n7636_8799.t41 464.166
R14005 a_n7636_8799.n244 a_n7636_8799.t114 464.166
R14006 a_n7636_8799.n235 a_n7636_8799.t113 464.166
R14007 a_n7636_8799.n243 a_n7636_8799.t45 464.166
R14008 a_n7636_8799.n242 a_n7636_8799.t44 464.166
R14009 a_n7636_8799.n236 a_n7636_8799.t135 464.166
R14010 a_n7636_8799.n241 a_n7636_8799.t66 464.166
R14011 a_n7636_8799.n240 a_n7636_8799.t48 464.166
R14012 a_n7636_8799.n237 a_n7636_8799.t136 464.166
R14013 a_n7636_8799.n239 a_n7636_8799.t95 464.166
R14014 a_n7636_8799.n83 a_n7636_8799.t146 485.135
R14015 a_n7636_8799.n270 a_n7636_8799.t43 464.166
R14016 a_n7636_8799.n252 a_n7636_8799.t93 464.166
R14017 a_n7636_8799.n269 a_n7636_8799.t30 464.166
R14018 a_n7636_8799.n268 a_n7636_8799.t117 464.166
R14019 a_n7636_8799.n253 a_n7636_8799.t54 464.166
R14020 a_n7636_8799.n267 a_n7636_8799.t100 464.166
R14021 a_n7636_8799.n266 a_n7636_8799.t35 464.166
R14022 a_n7636_8799.n254 a_n7636_8799.t60 464.166
R14023 a_n7636_8799.n265 a_n7636_8799.t140 464.166
R14024 a_n7636_8799.n264 a_n7636_8799.t109 464.166
R14025 a_n7636_8799.n255 a_n7636_8799.t134 464.166
R14026 a_n7636_8799.n263 a_n7636_8799.t91 464.166
R14027 a_n7636_8799.n262 a_n7636_8799.t112 464.166
R14028 a_n7636_8799.n256 a_n7636_8799.t47 464.166
R14029 a_n7636_8799.n261 a_n7636_8799.t131 464.166
R14030 a_n7636_8799.n260 a_n7636_8799.t72 464.166
R14031 a_n7636_8799.n257 a_n7636_8799.t123 464.166
R14032 a_n7636_8799.n259 a_n7636_8799.t59 464.166
R14033 a_n7636_8799.n159 a_n7636_8799.t129 464.166
R14034 a_n7636_8799.n160 a_n7636_8799.t79 464.166
R14035 a_n7636_8799.n161 a_n7636_8799.t108 464.166
R14036 a_n7636_8799.n162 a_n7636_8799.t125 464.166
R14037 a_n7636_8799.n157 a_n7636_8799.t75 464.166
R14038 a_n7636_8799.n163 a_n7636_8799.t76 464.166
R14039 a_n7636_8799.n164 a_n7636_8799.t106 464.166
R14040 a_n7636_8799.n165 a_n7636_8799.t63 464.166
R14041 a_n7636_8799.n166 a_n7636_8799.t64 464.166
R14042 a_n7636_8799.n156 a_n7636_8799.t103 464.166
R14043 a_n7636_8799.n167 a_n7636_8799.t28 464.166
R14044 a_n7636_8799.n155 a_n7636_8799.t61 464.166
R14045 a_n7636_8799.n168 a_n7636_8799.t84 464.166
R14046 a_n7636_8799.n169 a_n7636_8799.t128 464.166
R14047 a_n7636_8799.n170 a_n7636_8799.t40 464.166
R14048 a_n7636_8799.n171 a_n7636_8799.t58 464.166
R14049 a_n7636_8799.n154 a_n7636_8799.t124 464.166
R14050 a_n7636_8799.n172 a_n7636_8799.t37 464.166
R14051 a_n7636_8799.n178 a_n7636_8799.t145 464.166
R14052 a_n7636_8799.n179 a_n7636_8799.t89 464.166
R14053 a_n7636_8799.n180 a_n7636_8799.t121 464.166
R14054 a_n7636_8799.n181 a_n7636_8799.t139 464.166
R14055 a_n7636_8799.n176 a_n7636_8799.t85 464.166
R14056 a_n7636_8799.n182 a_n7636_8799.t86 464.166
R14057 a_n7636_8799.n183 a_n7636_8799.t119 464.166
R14058 a_n7636_8799.n184 a_n7636_8799.t73 464.166
R14059 a_n7636_8799.n185 a_n7636_8799.t74 464.166
R14060 a_n7636_8799.n175 a_n7636_8799.t115 464.166
R14061 a_n7636_8799.n186 a_n7636_8799.t39 464.166
R14062 a_n7636_8799.n174 a_n7636_8799.t70 464.166
R14063 a_n7636_8799.n187 a_n7636_8799.t97 464.166
R14064 a_n7636_8799.n188 a_n7636_8799.t143 464.166
R14065 a_n7636_8799.n189 a_n7636_8799.t55 464.166
R14066 a_n7636_8799.n190 a_n7636_8799.t69 464.166
R14067 a_n7636_8799.n173 a_n7636_8799.t137 464.166
R14068 a_n7636_8799.n191 a_n7636_8799.t49 464.166
R14069 a_n7636_8799.n198 a_n7636_8799.t82 464.166
R14070 a_n7636_8799.n199 a_n7636_8799.t120 464.166
R14071 a_n7636_8799.n200 a_n7636_8799.t71 464.166
R14072 a_n7636_8799.n201 a_n7636_8799.t130 464.166
R14073 a_n7636_8799.n196 a_n7636_8799.t46 464.166
R14074 a_n7636_8799.n202 a_n7636_8799.t29 464.166
R14075 a_n7636_8799.n203 a_n7636_8799.t90 464.166
R14076 a_n7636_8799.n204 a_n7636_8799.t133 464.166
R14077 a_n7636_8799.n205 a_n7636_8799.t107 464.166
R14078 a_n7636_8799.n195 a_n7636_8799.t138 464.166
R14079 a_n7636_8799.n206 a_n7636_8799.t83 464.166
R14080 a_n7636_8799.n194 a_n7636_8799.t34 464.166
R14081 a_n7636_8799.n207 a_n7636_8799.t99 464.166
R14082 a_n7636_8799.n208 a_n7636_8799.t53 464.166
R14083 a_n7636_8799.n209 a_n7636_8799.t116 464.166
R14084 a_n7636_8799.n210 a_n7636_8799.t62 464.166
R14085 a_n7636_8799.n193 a_n7636_8799.t92 464.166
R14086 a_n7636_8799.n211 a_n7636_8799.t42 464.166
R14087 a_n7636_8799.n41 a_n7636_8799.n67 71.7212
R14088 a_n7636_8799.n67 a_n7636_8799.n218 17.8606
R14089 a_n7636_8799.n66 a_n7636_8799.n41 76.9909
R14090 a_n7636_8799.n221 a_n7636_8799.n66 7.32118
R14091 a_n7636_8799.n65 a_n7636_8799.n40 78.3454
R14092 a_n7636_8799.n40 a_n7636_8799.n64 72.8951
R14093 a_n7636_8799.n63 a_n7636_8799.n42 70.1674
R14094 a_n7636_8799.n224 a_n7636_8799.n63 20.9683
R14095 a_n7636_8799.n42 a_n7636_8799.n62 72.3034
R14096 a_n7636_8799.n62 a_n7636_8799.n216 16.6962
R14097 a_n7636_8799.n61 a_n7636_8799.n43 77.6622
R14098 a_n7636_8799.n225 a_n7636_8799.n61 5.97853
R14099 a_n7636_8799.n60 a_n7636_8799.n43 77.6622
R14100 a_n7636_8799.n44 a_n7636_8799.n59 72.3034
R14101 a_n7636_8799.n58 a_n7636_8799.n44 70.1674
R14102 a_n7636_8799.n228 a_n7636_8799.n58 20.9683
R14103 a_n7636_8799.n46 a_n7636_8799.n57 72.8951
R14104 a_n7636_8799.n57 a_n7636_8799.n214 15.5127
R14105 a_n7636_8799.n56 a_n7636_8799.n46 78.3454
R14106 a_n7636_8799.n229 a_n7636_8799.n56 4.61226
R14107 a_n7636_8799.n55 a_n7636_8799.n45 76.9909
R14108 a_n7636_8799.n45 a_n7636_8799.n54 71.7212
R14109 a_n7636_8799.n231 a_n7636_8799.n53 20.9683
R14110 a_n7636_8799.n47 a_n7636_8799.n53 70.1674
R14111 a_n7636_8799.n33 a_n7636_8799.n82 71.7212
R14112 a_n7636_8799.n82 a_n7636_8799.n237 17.8606
R14113 a_n7636_8799.n81 a_n7636_8799.n33 76.9909
R14114 a_n7636_8799.n240 a_n7636_8799.n81 7.32118
R14115 a_n7636_8799.n80 a_n7636_8799.n32 78.3454
R14116 a_n7636_8799.n32 a_n7636_8799.n79 72.8951
R14117 a_n7636_8799.n78 a_n7636_8799.n34 70.1674
R14118 a_n7636_8799.n243 a_n7636_8799.n78 20.9683
R14119 a_n7636_8799.n34 a_n7636_8799.n77 72.3034
R14120 a_n7636_8799.n77 a_n7636_8799.n235 16.6962
R14121 a_n7636_8799.n76 a_n7636_8799.n35 77.6622
R14122 a_n7636_8799.n244 a_n7636_8799.n76 5.97853
R14123 a_n7636_8799.n75 a_n7636_8799.n35 77.6622
R14124 a_n7636_8799.n36 a_n7636_8799.n74 72.3034
R14125 a_n7636_8799.n73 a_n7636_8799.n36 70.1674
R14126 a_n7636_8799.n247 a_n7636_8799.n73 20.9683
R14127 a_n7636_8799.n38 a_n7636_8799.n72 72.8951
R14128 a_n7636_8799.n72 a_n7636_8799.n233 15.5127
R14129 a_n7636_8799.n71 a_n7636_8799.n38 78.3454
R14130 a_n7636_8799.n248 a_n7636_8799.n71 4.61226
R14131 a_n7636_8799.n70 a_n7636_8799.n37 76.9909
R14132 a_n7636_8799.n37 a_n7636_8799.n69 71.7212
R14133 a_n7636_8799.n250 a_n7636_8799.n68 20.9683
R14134 a_n7636_8799.n39 a_n7636_8799.n68 70.1674
R14135 a_n7636_8799.n25 a_n7636_8799.n97 71.7212
R14136 a_n7636_8799.n97 a_n7636_8799.n257 17.8606
R14137 a_n7636_8799.n96 a_n7636_8799.n25 76.9909
R14138 a_n7636_8799.n260 a_n7636_8799.n96 7.32118
R14139 a_n7636_8799.n95 a_n7636_8799.n24 78.3454
R14140 a_n7636_8799.n24 a_n7636_8799.n94 72.8951
R14141 a_n7636_8799.n93 a_n7636_8799.n26 70.1674
R14142 a_n7636_8799.n263 a_n7636_8799.n93 20.9683
R14143 a_n7636_8799.n26 a_n7636_8799.n92 72.3034
R14144 a_n7636_8799.n92 a_n7636_8799.n255 16.6962
R14145 a_n7636_8799.n91 a_n7636_8799.n27 77.6622
R14146 a_n7636_8799.n264 a_n7636_8799.n91 5.97853
R14147 a_n7636_8799.n90 a_n7636_8799.n27 77.6622
R14148 a_n7636_8799.n28 a_n7636_8799.n89 72.3034
R14149 a_n7636_8799.n88 a_n7636_8799.n28 70.1674
R14150 a_n7636_8799.n267 a_n7636_8799.n88 20.9683
R14151 a_n7636_8799.n30 a_n7636_8799.n87 72.8951
R14152 a_n7636_8799.n87 a_n7636_8799.n253 15.5127
R14153 a_n7636_8799.n86 a_n7636_8799.n30 78.3454
R14154 a_n7636_8799.n268 a_n7636_8799.n86 4.61226
R14155 a_n7636_8799.n85 a_n7636_8799.n29 76.9909
R14156 a_n7636_8799.n29 a_n7636_8799.n84 71.7212
R14157 a_n7636_8799.n270 a_n7636_8799.n83 20.9683
R14158 a_n7636_8799.n31 a_n7636_8799.n83 70.1674
R14159 a_n7636_8799.n17 a_n7636_8799.n112 70.1674
R14160 a_n7636_8799.n172 a_n7636_8799.n112 20.9683
R14161 a_n7636_8799.n111 a_n7636_8799.n17 71.7212
R14162 a_n7636_8799.n111 a_n7636_8799.n154 17.8606
R14163 a_n7636_8799.n16 a_n7636_8799.n110 76.9909
R14164 a_n7636_8799.n171 a_n7636_8799.n110 7.32118
R14165 a_n7636_8799.n109 a_n7636_8799.n16 78.3454
R14166 a_n7636_8799.n18 a_n7636_8799.n108 72.8951
R14167 a_n7636_8799.n107 a_n7636_8799.n18 70.1674
R14168 a_n7636_8799.n107 a_n7636_8799.n155 20.9683
R14169 a_n7636_8799.n19 a_n7636_8799.n106 72.3034
R14170 a_n7636_8799.n167 a_n7636_8799.n106 16.6962
R14171 a_n7636_8799.n105 a_n7636_8799.n19 77.6622
R14172 a_n7636_8799.n105 a_n7636_8799.n156 5.97853
R14173 a_n7636_8799.n20 a_n7636_8799.n104 77.6622
R14174 a_n7636_8799.n103 a_n7636_8799.n20 72.3034
R14175 a_n7636_8799.n21 a_n7636_8799.n102 70.1674
R14176 a_n7636_8799.n163 a_n7636_8799.n102 20.9683
R14177 a_n7636_8799.n101 a_n7636_8799.n21 72.8951
R14178 a_n7636_8799.n101 a_n7636_8799.n157 15.5127
R14179 a_n7636_8799.n22 a_n7636_8799.n100 78.3454
R14180 a_n7636_8799.n162 a_n7636_8799.n100 4.61226
R14181 a_n7636_8799.n99 a_n7636_8799.n22 76.9909
R14182 a_n7636_8799.n98 a_n7636_8799.n160 17.8606
R14183 a_n7636_8799.n98 a_n7636_8799.n23 71.7212
R14184 a_n7636_8799.n9 a_n7636_8799.n127 70.1674
R14185 a_n7636_8799.n191 a_n7636_8799.n127 20.9683
R14186 a_n7636_8799.n126 a_n7636_8799.n9 71.7212
R14187 a_n7636_8799.n126 a_n7636_8799.n173 17.8606
R14188 a_n7636_8799.n8 a_n7636_8799.n125 76.9909
R14189 a_n7636_8799.n190 a_n7636_8799.n125 7.32118
R14190 a_n7636_8799.n124 a_n7636_8799.n8 78.3454
R14191 a_n7636_8799.n10 a_n7636_8799.n123 72.8951
R14192 a_n7636_8799.n122 a_n7636_8799.n10 70.1674
R14193 a_n7636_8799.n122 a_n7636_8799.n174 20.9683
R14194 a_n7636_8799.n11 a_n7636_8799.n121 72.3034
R14195 a_n7636_8799.n186 a_n7636_8799.n121 16.6962
R14196 a_n7636_8799.n120 a_n7636_8799.n11 77.6622
R14197 a_n7636_8799.n120 a_n7636_8799.n175 5.97853
R14198 a_n7636_8799.n12 a_n7636_8799.n119 77.6622
R14199 a_n7636_8799.n118 a_n7636_8799.n12 72.3034
R14200 a_n7636_8799.n13 a_n7636_8799.n117 70.1674
R14201 a_n7636_8799.n182 a_n7636_8799.n117 20.9683
R14202 a_n7636_8799.n116 a_n7636_8799.n13 72.8951
R14203 a_n7636_8799.n116 a_n7636_8799.n176 15.5127
R14204 a_n7636_8799.n14 a_n7636_8799.n115 78.3454
R14205 a_n7636_8799.n181 a_n7636_8799.n115 4.61226
R14206 a_n7636_8799.n114 a_n7636_8799.n14 76.9909
R14207 a_n7636_8799.n113 a_n7636_8799.n179 17.8606
R14208 a_n7636_8799.n113 a_n7636_8799.n15 71.7212
R14209 a_n7636_8799.n1 a_n7636_8799.n142 70.1674
R14210 a_n7636_8799.n211 a_n7636_8799.n142 20.9683
R14211 a_n7636_8799.n141 a_n7636_8799.n1 71.7212
R14212 a_n7636_8799.n141 a_n7636_8799.n193 17.8606
R14213 a_n7636_8799.n0 a_n7636_8799.n140 76.9909
R14214 a_n7636_8799.n210 a_n7636_8799.n140 7.32118
R14215 a_n7636_8799.n139 a_n7636_8799.n0 78.3454
R14216 a_n7636_8799.n2 a_n7636_8799.n138 72.8951
R14217 a_n7636_8799.n137 a_n7636_8799.n2 70.1674
R14218 a_n7636_8799.n137 a_n7636_8799.n194 20.9683
R14219 a_n7636_8799.n3 a_n7636_8799.n136 72.3034
R14220 a_n7636_8799.n206 a_n7636_8799.n136 16.6962
R14221 a_n7636_8799.n135 a_n7636_8799.n3 77.6622
R14222 a_n7636_8799.n135 a_n7636_8799.n195 5.97853
R14223 a_n7636_8799.n4 a_n7636_8799.n134 77.6622
R14224 a_n7636_8799.n133 a_n7636_8799.n4 72.3034
R14225 a_n7636_8799.n5 a_n7636_8799.n132 70.1674
R14226 a_n7636_8799.n202 a_n7636_8799.n132 20.9683
R14227 a_n7636_8799.n131 a_n7636_8799.n5 72.8951
R14228 a_n7636_8799.n131 a_n7636_8799.n196 15.5127
R14229 a_n7636_8799.n6 a_n7636_8799.n130 78.3454
R14230 a_n7636_8799.n201 a_n7636_8799.n130 4.61226
R14231 a_n7636_8799.n129 a_n7636_8799.n6 76.9909
R14232 a_n7636_8799.n128 a_n7636_8799.n199 17.8606
R14233 a_n7636_8799.n128 a_n7636_8799.n7 71.7212
R14234 a_n7636_8799.n48 a_n7636_8799.n143 98.9633
R14235 a_n7636_8799.n49 a_n7636_8799.n276 98.9631
R14236 a_n7636_8799.n49 a_n7636_8799.n275 98.6055
R14237 a_n7636_8799.n48 a_n7636_8799.n145 98.6055
R14238 a_n7636_8799.n48 a_n7636_8799.n144 98.6055
R14239 a_n7636_8799.n277 a_n7636_8799.n49 98.6054
R14240 a_n7636_8799.n51 a_n7636_8799.n146 81.2902
R14241 a_n7636_8799.n52 a_n7636_8799.n150 81.2902
R14242 a_n7636_8799.n52 a_n7636_8799.n148 81.2902
R14243 a_n7636_8799.n50 a_n7636_8799.n152 80.9324
R14244 a_n7636_8799.n51 a_n7636_8799.n153 80.9324
R14245 a_n7636_8799.n51 a_n7636_8799.n147 80.9324
R14246 a_n7636_8799.n52 a_n7636_8799.n151 80.9324
R14247 a_n7636_8799.n52 a_n7636_8799.n149 80.9324
R14248 a_n7636_8799.n41 a_n7636_8799.n219 70.4033
R14249 a_n7636_8799.n33 a_n7636_8799.n238 70.4033
R14250 a_n7636_8799.n25 a_n7636_8799.n258 70.4033
R14251 a_n7636_8799.n158 a_n7636_8799.n23 70.4033
R14252 a_n7636_8799.n177 a_n7636_8799.n15 70.4033
R14253 a_n7636_8799.n197 a_n7636_8799.n7 70.4033
R14254 a_n7636_8799.n230 a_n7636_8799.n229 48.2005
R14255 a_n7636_8799.n58 a_n7636_8799.n227 20.9683
R14256 a_n7636_8799.n226 a_n7636_8799.n225 48.2005
R14257 a_n7636_8799.n63 a_n7636_8799.n223 20.9683
R14258 a_n7636_8799.n222 a_n7636_8799.n221 48.2005
R14259 a_n7636_8799.n249 a_n7636_8799.n248 48.2005
R14260 a_n7636_8799.n73 a_n7636_8799.n246 20.9683
R14261 a_n7636_8799.n245 a_n7636_8799.n244 48.2005
R14262 a_n7636_8799.n78 a_n7636_8799.n242 20.9683
R14263 a_n7636_8799.n241 a_n7636_8799.n240 48.2005
R14264 a_n7636_8799.n269 a_n7636_8799.n268 48.2005
R14265 a_n7636_8799.n88 a_n7636_8799.n266 20.9683
R14266 a_n7636_8799.n265 a_n7636_8799.n264 48.2005
R14267 a_n7636_8799.n93 a_n7636_8799.n262 20.9683
R14268 a_n7636_8799.n261 a_n7636_8799.n260 48.2005
R14269 a_n7636_8799.n162 a_n7636_8799.n161 48.2005
R14270 a_n7636_8799.n164 a_n7636_8799.n102 20.9683
R14271 a_n7636_8799.n166 a_n7636_8799.n156 48.2005
R14272 a_n7636_8799.n168 a_n7636_8799.n107 20.9683
R14273 a_n7636_8799.n171 a_n7636_8799.n170 48.2005
R14274 a_n7636_8799.t38 a_n7636_8799.n112 485.135
R14275 a_n7636_8799.n181 a_n7636_8799.n180 48.2005
R14276 a_n7636_8799.n183 a_n7636_8799.n117 20.9683
R14277 a_n7636_8799.n185 a_n7636_8799.n175 48.2005
R14278 a_n7636_8799.n187 a_n7636_8799.n122 20.9683
R14279 a_n7636_8799.n190 a_n7636_8799.n189 48.2005
R14280 a_n7636_8799.t51 a_n7636_8799.n127 485.135
R14281 a_n7636_8799.n201 a_n7636_8799.n200 48.2005
R14282 a_n7636_8799.n203 a_n7636_8799.n132 20.9683
R14283 a_n7636_8799.n205 a_n7636_8799.n195 48.2005
R14284 a_n7636_8799.n207 a_n7636_8799.n137 20.9683
R14285 a_n7636_8799.n210 a_n7636_8799.n209 48.2005
R14286 a_n7636_8799.t144 a_n7636_8799.n142 485.135
R14287 a_n7636_8799.n54 a_n7636_8799.n213 17.8606
R14288 a_n7636_8799.n220 a_n7636_8799.n67 25.894
R14289 a_n7636_8799.n69 a_n7636_8799.n232 17.8606
R14290 a_n7636_8799.n239 a_n7636_8799.n82 25.894
R14291 a_n7636_8799.n84 a_n7636_8799.n252 17.8606
R14292 a_n7636_8799.n259 a_n7636_8799.n97 25.894
R14293 a_n7636_8799.n172 a_n7636_8799.n111 25.894
R14294 a_n7636_8799.n191 a_n7636_8799.n126 25.894
R14295 a_n7636_8799.n211 a_n7636_8799.n141 25.894
R14296 a_n7636_8799.n65 a_n7636_8799.n217 43.3183
R14297 a_n7636_8799.n80 a_n7636_8799.n236 43.3183
R14298 a_n7636_8799.n95 a_n7636_8799.n256 43.3183
R14299 a_n7636_8799.n169 a_n7636_8799.n109 43.3183
R14300 a_n7636_8799.n188 a_n7636_8799.n124 43.3183
R14301 a_n7636_8799.n208 a_n7636_8799.n139 43.3183
R14302 a_n7636_8799.n59 a_n7636_8799.n215 16.6962
R14303 a_n7636_8799.n224 a_n7636_8799.n62 27.6507
R14304 a_n7636_8799.n74 a_n7636_8799.n234 16.6962
R14305 a_n7636_8799.n243 a_n7636_8799.n77 27.6507
R14306 a_n7636_8799.n89 a_n7636_8799.n254 16.6962
R14307 a_n7636_8799.n263 a_n7636_8799.n92 27.6507
R14308 a_n7636_8799.n165 a_n7636_8799.n103 16.6962
R14309 a_n7636_8799.n155 a_n7636_8799.n106 27.6507
R14310 a_n7636_8799.n184 a_n7636_8799.n118 16.6962
R14311 a_n7636_8799.n174 a_n7636_8799.n121 27.6507
R14312 a_n7636_8799.n204 a_n7636_8799.n133 16.6962
R14313 a_n7636_8799.n194 a_n7636_8799.n136 27.6507
R14314 a_n7636_8799.n60 a_n7636_8799.n215 41.7634
R14315 a_n7636_8799.n75 a_n7636_8799.n234 41.7634
R14316 a_n7636_8799.n90 a_n7636_8799.n254 41.7634
R14317 a_n7636_8799.n104 a_n7636_8799.n165 41.7634
R14318 a_n7636_8799.n119 a_n7636_8799.n184 41.7634
R14319 a_n7636_8799.n134 a_n7636_8799.n204 41.7634
R14320 a_n7636_8799.n228 a_n7636_8799.n57 29.3885
R14321 a_n7636_8799.n64 a_n7636_8799.n217 15.5127
R14322 a_n7636_8799.n247 a_n7636_8799.n72 29.3885
R14323 a_n7636_8799.n79 a_n7636_8799.n236 15.5127
R14324 a_n7636_8799.n267 a_n7636_8799.n87 29.3885
R14325 a_n7636_8799.n94 a_n7636_8799.n256 15.5127
R14326 a_n7636_8799.n163 a_n7636_8799.n101 29.3885
R14327 a_n7636_8799.n169 a_n7636_8799.n108 15.5127
R14328 a_n7636_8799.n182 a_n7636_8799.n116 29.3885
R14329 a_n7636_8799.n188 a_n7636_8799.n123 15.5127
R14330 a_n7636_8799.n202 a_n7636_8799.n131 29.3885
R14331 a_n7636_8799.n208 a_n7636_8799.n138 15.5127
R14332 a_n7636_8799.n55 a_n7636_8799.n213 40.1848
R14333 a_n7636_8799.n70 a_n7636_8799.n232 40.1848
R14334 a_n7636_8799.n85 a_n7636_8799.n252 40.1848
R14335 a_n7636_8799.n160 a_n7636_8799.n99 40.1848
R14336 a_n7636_8799.n179 a_n7636_8799.n114 40.1848
R14337 a_n7636_8799.n199 a_n7636_8799.n129 40.1848
R14338 a_n7636_8799.n220 a_n7636_8799.n219 20.9576
R14339 a_n7636_8799.n239 a_n7636_8799.n238 20.9576
R14340 a_n7636_8799.n259 a_n7636_8799.n258 20.9576
R14341 a_n7636_8799.n159 a_n7636_8799.n158 20.9576
R14342 a_n7636_8799.n178 a_n7636_8799.n177 20.9576
R14343 a_n7636_8799.n198 a_n7636_8799.n197 20.9576
R14344 a_n7636_8799.n55 a_n7636_8799.n230 7.32118
R14345 a_n7636_8799.n66 a_n7636_8799.n218 40.1848
R14346 a_n7636_8799.n70 a_n7636_8799.n249 7.32118
R14347 a_n7636_8799.n81 a_n7636_8799.n237 40.1848
R14348 a_n7636_8799.n85 a_n7636_8799.n269 7.32118
R14349 a_n7636_8799.n96 a_n7636_8799.n257 40.1848
R14350 a_n7636_8799.n161 a_n7636_8799.n99 7.32118
R14351 a_n7636_8799.n154 a_n7636_8799.n110 40.1848
R14352 a_n7636_8799.n180 a_n7636_8799.n114 7.32118
R14353 a_n7636_8799.n173 a_n7636_8799.n125 40.1848
R14354 a_n7636_8799.n200 a_n7636_8799.n129 7.32118
R14355 a_n7636_8799.n193 a_n7636_8799.n140 40.1848
R14356 a_n7636_8799.n223 a_n7636_8799.n64 29.3885
R14357 a_n7636_8799.n242 a_n7636_8799.n79 29.3885
R14358 a_n7636_8799.n262 a_n7636_8799.n94 29.3885
R14359 a_n7636_8799.n108 a_n7636_8799.n168 29.3885
R14360 a_n7636_8799.n123 a_n7636_8799.n187 29.3885
R14361 a_n7636_8799.n138 a_n7636_8799.n207 29.3885
R14362 a_n7636_8799.n60 a_n7636_8799.n226 5.97853
R14363 a_n7636_8799.n61 a_n7636_8799.n216 41.7634
R14364 a_n7636_8799.n75 a_n7636_8799.n245 5.97853
R14365 a_n7636_8799.n76 a_n7636_8799.n235 41.7634
R14366 a_n7636_8799.n90 a_n7636_8799.n265 5.97853
R14367 a_n7636_8799.n91 a_n7636_8799.n255 41.7634
R14368 a_n7636_8799.n166 a_n7636_8799.n104 5.97853
R14369 a_n7636_8799.n167 a_n7636_8799.n105 41.7634
R14370 a_n7636_8799.n185 a_n7636_8799.n119 5.97853
R14371 a_n7636_8799.n186 a_n7636_8799.n120 41.7634
R14372 a_n7636_8799.n205 a_n7636_8799.n134 5.97853
R14373 a_n7636_8799.n206 a_n7636_8799.n135 41.7634
R14374 a_n7636_8799.n273 a_n7636_8799.n51 12.3339
R14375 a_n7636_8799.n274 a_n7636_8799.n273 11.4887
R14376 a_n7636_8799.n227 a_n7636_8799.n59 27.6507
R14377 a_n7636_8799.n246 a_n7636_8799.n74 27.6507
R14378 a_n7636_8799.n266 a_n7636_8799.n89 27.6507
R14379 a_n7636_8799.n164 a_n7636_8799.n103 27.6507
R14380 a_n7636_8799.n183 a_n7636_8799.n118 27.6507
R14381 a_n7636_8799.n203 a_n7636_8799.n133 27.6507
R14382 a_n7636_8799.n56 a_n7636_8799.n214 43.3183
R14383 a_n7636_8799.n65 a_n7636_8799.n222 4.61226
R14384 a_n7636_8799.n71 a_n7636_8799.n233 43.3183
R14385 a_n7636_8799.n80 a_n7636_8799.n241 4.61226
R14386 a_n7636_8799.n86 a_n7636_8799.n253 43.3183
R14387 a_n7636_8799.n95 a_n7636_8799.n261 4.61226
R14388 a_n7636_8799.n157 a_n7636_8799.n100 43.3183
R14389 a_n7636_8799.n170 a_n7636_8799.n109 4.61226
R14390 a_n7636_8799.n176 a_n7636_8799.n115 43.3183
R14391 a_n7636_8799.n189 a_n7636_8799.n124 4.61226
R14392 a_n7636_8799.n196 a_n7636_8799.n130 43.3183
R14393 a_n7636_8799.n50 a_n7636_8799.n52 31.7978
R14394 a_n7636_8799.n49 a_n7636_8799.n274 30.6769
R14395 a_n7636_8799.n209 a_n7636_8799.n139 4.61226
R14396 a_n7636_8799.n251 a_n7636_8799.n47 9.04406
R14397 a_n7636_8799.n192 a_n7636_8799.n17 9.04406
R14398 a_n7636_8799.n231 a_n7636_8799.n54 25.894
R14399 a_n7636_8799.n250 a_n7636_8799.n69 25.894
R14400 a_n7636_8799.n270 a_n7636_8799.n84 25.894
R14401 a_n7636_8799.n98 a_n7636_8799.n159 25.894
R14402 a_n7636_8799.n113 a_n7636_8799.n178 25.894
R14403 a_n7636_8799.n128 a_n7636_8799.n198 25.894
R14404 a_n7636_8799.n274 a_n7636_8799.n48 18.4882
R14405 a_n7636_8799.n272 a_n7636_8799.n212 6.81251
R14406 a_n7636_8799.n272 a_n7636_8799.n271 6.5703
R14407 a_n7636_8799.n251 a_n7636_8799.n39 4.93611
R14408 a_n7636_8799.n271 a_n7636_8799.n31 4.93611
R14409 a_n7636_8799.n192 a_n7636_8799.n9 4.93611
R14410 a_n7636_8799.n212 a_n7636_8799.n1 4.93611
R14411 a_n7636_8799.n271 a_n7636_8799.n251 4.10845
R14412 a_n7636_8799.n212 a_n7636_8799.n192 4.10845
R14413 a_n7636_8799.n276 a_n7636_8799.t26 3.61217
R14414 a_n7636_8799.n276 a_n7636_8799.t4 3.61217
R14415 a_n7636_8799.n275 a_n7636_8799.t19 3.61217
R14416 a_n7636_8799.n275 a_n7636_8799.t10 3.61217
R14417 a_n7636_8799.n145 a_n7636_8799.t15 3.61217
R14418 a_n7636_8799.n145 a_n7636_8799.t2 3.61217
R14419 a_n7636_8799.n144 a_n7636_8799.t22 3.61217
R14420 a_n7636_8799.n144 a_n7636_8799.t1 3.61217
R14421 a_n7636_8799.n143 a_n7636_8799.t3 3.61217
R14422 a_n7636_8799.n143 a_n7636_8799.t5 3.61217
R14423 a_n7636_8799.t0 a_n7636_8799.n277 3.61217
R14424 a_n7636_8799.n277 a_n7636_8799.t25 3.61217
R14425 a_n7636_8799.n273 a_n7636_8799.n272 3.4105
R14426 a_n7636_8799.n152 a_n7636_8799.t20 2.82907
R14427 a_n7636_8799.n152 a_n7636_8799.t6 2.82907
R14428 a_n7636_8799.n153 a_n7636_8799.t24 2.82907
R14429 a_n7636_8799.n153 a_n7636_8799.t18 2.82907
R14430 a_n7636_8799.n147 a_n7636_8799.t14 2.82907
R14431 a_n7636_8799.n147 a_n7636_8799.t16 2.82907
R14432 a_n7636_8799.n146 a_n7636_8799.t11 2.82907
R14433 a_n7636_8799.n146 a_n7636_8799.t23 2.82907
R14434 a_n7636_8799.n150 a_n7636_8799.t21 2.82907
R14435 a_n7636_8799.n150 a_n7636_8799.t9 2.82907
R14436 a_n7636_8799.n151 a_n7636_8799.t13 2.82907
R14437 a_n7636_8799.n151 a_n7636_8799.t27 2.82907
R14438 a_n7636_8799.n149 a_n7636_8799.t7 2.82907
R14439 a_n7636_8799.n149 a_n7636_8799.t17 2.82907
R14440 a_n7636_8799.n148 a_n7636_8799.t12 2.82907
R14441 a_n7636_8799.n148 a_n7636_8799.t8 2.82907
R14442 a_n7636_8799.n41 a_n7636_8799.n40 1.13686
R14443 a_n7636_8799.n33 a_n7636_8799.n32 1.13686
R14444 a_n7636_8799.n25 a_n7636_8799.n24 1.13686
R14445 a_n7636_8799.n17 a_n7636_8799.n16 1.13686
R14446 a_n7636_8799.n9 a_n7636_8799.n8 1.13686
R14447 a_n7636_8799.n1 a_n7636_8799.n0 1.13686
R14448 a_n7636_8799.n46 a_n7636_8799.n45 0.758076
R14449 a_n7636_8799.n46 a_n7636_8799.n44 0.758076
R14450 a_n7636_8799.n44 a_n7636_8799.n43 0.758076
R14451 a_n7636_8799.n43 a_n7636_8799.n42 0.758076
R14452 a_n7636_8799.n40 a_n7636_8799.n42 0.758076
R14453 a_n7636_8799.n38 a_n7636_8799.n37 0.758076
R14454 a_n7636_8799.n38 a_n7636_8799.n36 0.758076
R14455 a_n7636_8799.n36 a_n7636_8799.n35 0.758076
R14456 a_n7636_8799.n35 a_n7636_8799.n34 0.758076
R14457 a_n7636_8799.n32 a_n7636_8799.n34 0.758076
R14458 a_n7636_8799.n30 a_n7636_8799.n29 0.758076
R14459 a_n7636_8799.n30 a_n7636_8799.n28 0.758076
R14460 a_n7636_8799.n28 a_n7636_8799.n27 0.758076
R14461 a_n7636_8799.n27 a_n7636_8799.n26 0.758076
R14462 a_n7636_8799.n24 a_n7636_8799.n26 0.758076
R14463 a_n7636_8799.n21 a_n7636_8799.n22 0.758076
R14464 a_n7636_8799.n20 a_n7636_8799.n21 0.758076
R14465 a_n7636_8799.n19 a_n7636_8799.n20 0.758076
R14466 a_n7636_8799.n18 a_n7636_8799.n19 0.758076
R14467 a_n7636_8799.n16 a_n7636_8799.n18 0.758076
R14468 a_n7636_8799.n13 a_n7636_8799.n14 0.758076
R14469 a_n7636_8799.n12 a_n7636_8799.n13 0.758076
R14470 a_n7636_8799.n11 a_n7636_8799.n12 0.758076
R14471 a_n7636_8799.n10 a_n7636_8799.n11 0.758076
R14472 a_n7636_8799.n8 a_n7636_8799.n10 0.758076
R14473 a_n7636_8799.n5 a_n7636_8799.n6 0.758076
R14474 a_n7636_8799.n4 a_n7636_8799.n5 0.758076
R14475 a_n7636_8799.n3 a_n7636_8799.n4 0.758076
R14476 a_n7636_8799.n2 a_n7636_8799.n3 0.758076
R14477 a_n7636_8799.n0 a_n7636_8799.n2 0.758076
R14478 a_n7636_8799.n51 a_n7636_8799.n50 0.716017
R14479 a_n7636_8799.n6 a_n7636_8799.n7 0.568682
R14480 a_n7636_8799.n14 a_n7636_8799.n15 0.568682
R14481 a_n7636_8799.n22 a_n7636_8799.n23 0.568682
R14482 a_n7636_8799.n29 a_n7636_8799.n31 0.568682
R14483 a_n7636_8799.n37 a_n7636_8799.n39 0.568682
R14484 a_n7636_8799.n45 a_n7636_8799.n47 0.568682
R14485 vdd.n327 vdd.n291 756.745
R14486 vdd.n268 vdd.n232 756.745
R14487 vdd.n225 vdd.n189 756.745
R14488 vdd.n166 vdd.n130 756.745
R14489 vdd.n124 vdd.n88 756.745
R14490 vdd.n65 vdd.n29 756.745
R14491 vdd.n1746 vdd.n1710 756.745
R14492 vdd.n1805 vdd.n1769 756.745
R14493 vdd.n1644 vdd.n1608 756.745
R14494 vdd.n1703 vdd.n1667 756.745
R14495 vdd.n1543 vdd.n1507 756.745
R14496 vdd.n1602 vdd.n1566 756.745
R14497 vdd.n2177 vdd.t265 640.208
R14498 vdd.n965 vdd.t250 640.208
R14499 vdd.n2151 vdd.t211 640.208
R14500 vdd.n957 vdd.t275 640.208
R14501 vdd.n2922 vdd.t226 640.208
R14502 vdd.n2642 vdd.t272 640.208
R14503 vdd.n832 vdd.t254 640.208
R14504 vdd.n2639 vdd.t258 640.208
R14505 vdd.n799 vdd.t262 640.208
R14506 vdd.n1027 vdd.t268 640.208
R14507 vdd.n1317 vdd.t241 592.009
R14508 vdd.n1355 vdd.t230 592.009
R14509 vdd.n1251 vdd.t244 592.009
R14510 vdd.n2333 vdd.t222 592.009
R14511 vdd.n1970 vdd.t234 592.009
R14512 vdd.n1930 vdd.t247 592.009
R14513 vdd.n426 vdd.t237 592.009
R14514 vdd.n440 vdd.t278 592.009
R14515 vdd.n452 vdd.t284 592.009
R14516 vdd.n768 vdd.t215 592.009
R14517 vdd.n3184 vdd.t219 592.009
R14518 vdd.n688 vdd.t281 592.009
R14519 vdd.n328 vdd.n327 585
R14520 vdd.n326 vdd.n293 585
R14521 vdd.n325 vdd.n324 585
R14522 vdd.n296 vdd.n294 585
R14523 vdd.n319 vdd.n318 585
R14524 vdd.n317 vdd.n316 585
R14525 vdd.n300 vdd.n299 585
R14526 vdd.n311 vdd.n310 585
R14527 vdd.n309 vdd.n308 585
R14528 vdd.n304 vdd.n303 585
R14529 vdd.n269 vdd.n268 585
R14530 vdd.n267 vdd.n234 585
R14531 vdd.n266 vdd.n265 585
R14532 vdd.n237 vdd.n235 585
R14533 vdd.n260 vdd.n259 585
R14534 vdd.n258 vdd.n257 585
R14535 vdd.n241 vdd.n240 585
R14536 vdd.n252 vdd.n251 585
R14537 vdd.n250 vdd.n249 585
R14538 vdd.n245 vdd.n244 585
R14539 vdd.n226 vdd.n225 585
R14540 vdd.n224 vdd.n191 585
R14541 vdd.n223 vdd.n222 585
R14542 vdd.n194 vdd.n192 585
R14543 vdd.n217 vdd.n216 585
R14544 vdd.n215 vdd.n214 585
R14545 vdd.n198 vdd.n197 585
R14546 vdd.n209 vdd.n208 585
R14547 vdd.n207 vdd.n206 585
R14548 vdd.n202 vdd.n201 585
R14549 vdd.n167 vdd.n166 585
R14550 vdd.n165 vdd.n132 585
R14551 vdd.n164 vdd.n163 585
R14552 vdd.n135 vdd.n133 585
R14553 vdd.n158 vdd.n157 585
R14554 vdd.n156 vdd.n155 585
R14555 vdd.n139 vdd.n138 585
R14556 vdd.n150 vdd.n149 585
R14557 vdd.n148 vdd.n147 585
R14558 vdd.n143 vdd.n142 585
R14559 vdd.n125 vdd.n124 585
R14560 vdd.n123 vdd.n90 585
R14561 vdd.n122 vdd.n121 585
R14562 vdd.n93 vdd.n91 585
R14563 vdd.n116 vdd.n115 585
R14564 vdd.n114 vdd.n113 585
R14565 vdd.n97 vdd.n96 585
R14566 vdd.n108 vdd.n107 585
R14567 vdd.n106 vdd.n105 585
R14568 vdd.n101 vdd.n100 585
R14569 vdd.n66 vdd.n65 585
R14570 vdd.n64 vdd.n31 585
R14571 vdd.n63 vdd.n62 585
R14572 vdd.n34 vdd.n32 585
R14573 vdd.n57 vdd.n56 585
R14574 vdd.n55 vdd.n54 585
R14575 vdd.n38 vdd.n37 585
R14576 vdd.n49 vdd.n48 585
R14577 vdd.n47 vdd.n46 585
R14578 vdd.n42 vdd.n41 585
R14579 vdd.n1747 vdd.n1746 585
R14580 vdd.n1745 vdd.n1712 585
R14581 vdd.n1744 vdd.n1743 585
R14582 vdd.n1715 vdd.n1713 585
R14583 vdd.n1738 vdd.n1737 585
R14584 vdd.n1736 vdd.n1735 585
R14585 vdd.n1719 vdd.n1718 585
R14586 vdd.n1730 vdd.n1729 585
R14587 vdd.n1728 vdd.n1727 585
R14588 vdd.n1723 vdd.n1722 585
R14589 vdd.n1806 vdd.n1805 585
R14590 vdd.n1804 vdd.n1771 585
R14591 vdd.n1803 vdd.n1802 585
R14592 vdd.n1774 vdd.n1772 585
R14593 vdd.n1797 vdd.n1796 585
R14594 vdd.n1795 vdd.n1794 585
R14595 vdd.n1778 vdd.n1777 585
R14596 vdd.n1789 vdd.n1788 585
R14597 vdd.n1787 vdd.n1786 585
R14598 vdd.n1782 vdd.n1781 585
R14599 vdd.n1645 vdd.n1644 585
R14600 vdd.n1643 vdd.n1610 585
R14601 vdd.n1642 vdd.n1641 585
R14602 vdd.n1613 vdd.n1611 585
R14603 vdd.n1636 vdd.n1635 585
R14604 vdd.n1634 vdd.n1633 585
R14605 vdd.n1617 vdd.n1616 585
R14606 vdd.n1628 vdd.n1627 585
R14607 vdd.n1626 vdd.n1625 585
R14608 vdd.n1621 vdd.n1620 585
R14609 vdd.n1704 vdd.n1703 585
R14610 vdd.n1702 vdd.n1669 585
R14611 vdd.n1701 vdd.n1700 585
R14612 vdd.n1672 vdd.n1670 585
R14613 vdd.n1695 vdd.n1694 585
R14614 vdd.n1693 vdd.n1692 585
R14615 vdd.n1676 vdd.n1675 585
R14616 vdd.n1687 vdd.n1686 585
R14617 vdd.n1685 vdd.n1684 585
R14618 vdd.n1680 vdd.n1679 585
R14619 vdd.n1544 vdd.n1543 585
R14620 vdd.n1542 vdd.n1509 585
R14621 vdd.n1541 vdd.n1540 585
R14622 vdd.n1512 vdd.n1510 585
R14623 vdd.n1535 vdd.n1534 585
R14624 vdd.n1533 vdd.n1532 585
R14625 vdd.n1516 vdd.n1515 585
R14626 vdd.n1527 vdd.n1526 585
R14627 vdd.n1525 vdd.n1524 585
R14628 vdd.n1520 vdd.n1519 585
R14629 vdd.n1603 vdd.n1602 585
R14630 vdd.n1601 vdd.n1568 585
R14631 vdd.n1600 vdd.n1599 585
R14632 vdd.n1571 vdd.n1569 585
R14633 vdd.n1594 vdd.n1593 585
R14634 vdd.n1592 vdd.n1591 585
R14635 vdd.n1575 vdd.n1574 585
R14636 vdd.n1586 vdd.n1585 585
R14637 vdd.n1584 vdd.n1583 585
R14638 vdd.n1579 vdd.n1578 585
R14639 vdd.n3356 vdd.n392 509.269
R14640 vdd.n3352 vdd.n393 509.269
R14641 vdd.n3224 vdd.n685 509.269
R14642 vdd.n3221 vdd.n684 509.269
R14643 vdd.n2328 vdd.n1075 509.269
R14644 vdd.n2331 vdd.n2330 509.269
R14645 vdd.n1224 vdd.n1188 509.269
R14646 vdd.n1420 vdd.n1189 509.269
R14647 vdd.n305 vdd.t144 329.043
R14648 vdd.n246 vdd.t119 329.043
R14649 vdd.n203 vdd.t134 329.043
R14650 vdd.n144 vdd.t104 329.043
R14651 vdd.n102 vdd.t83 329.043
R14652 vdd.n43 vdd.t18 329.043
R14653 vdd.n1724 vdd.t164 329.043
R14654 vdd.n1783 vdd.t50 329.043
R14655 vdd.n1622 vdd.t149 329.043
R14656 vdd.n1681 vdd.t26 329.043
R14657 vdd.n1521 vdd.t22 329.043
R14658 vdd.n1580 vdd.t84 329.043
R14659 vdd.n1317 vdd.t243 319.788
R14660 vdd.n1355 vdd.t233 319.788
R14661 vdd.n1251 vdd.t246 319.788
R14662 vdd.n2333 vdd.t224 319.788
R14663 vdd.n1970 vdd.t235 319.788
R14664 vdd.n1930 vdd.t248 319.788
R14665 vdd.n426 vdd.t239 319.788
R14666 vdd.n440 vdd.t279 319.788
R14667 vdd.n452 vdd.t285 319.788
R14668 vdd.n768 vdd.t218 319.788
R14669 vdd.n3184 vdd.t221 319.788
R14670 vdd.n688 vdd.t283 319.788
R14671 vdd.n1318 vdd.t242 303.69
R14672 vdd.n1356 vdd.t232 303.69
R14673 vdd.n1252 vdd.t245 303.69
R14674 vdd.n2334 vdd.t225 303.69
R14675 vdd.n1971 vdd.t236 303.69
R14676 vdd.n1931 vdd.t249 303.69
R14677 vdd.n427 vdd.t240 303.69
R14678 vdd.n441 vdd.t280 303.69
R14679 vdd.n453 vdd.t286 303.69
R14680 vdd.n769 vdd.t217 303.69
R14681 vdd.n3185 vdd.t220 303.69
R14682 vdd.n689 vdd.t282 303.69
R14683 vdd.n2865 vdd.n913 297.074
R14684 vdd.n3058 vdd.n809 297.074
R14685 vdd.n2995 vdd.n806 297.074
R14686 vdd.n2788 vdd.n914 297.074
R14687 vdd.n2603 vdd.n954 297.074
R14688 vdd.n2534 vdd.n2533 297.074
R14689 vdd.n2280 vdd.n1050 297.074
R14690 vdd.n2376 vdd.n1048 297.074
R14691 vdd.n2974 vdd.n807 297.074
R14692 vdd.n3061 vdd.n3060 297.074
R14693 vdd.n2637 vdd.n915 297.074
R14694 vdd.n2863 vdd.n916 297.074
R14695 vdd.n2531 vdd.n963 297.074
R14696 vdd.n961 vdd.n936 297.074
R14697 vdd.n2217 vdd.n1051 297.074
R14698 vdd.n2374 vdd.n1052 297.074
R14699 vdd.n2976 vdd.n807 185
R14700 vdd.n3059 vdd.n807 185
R14701 vdd.n2978 vdd.n2977 185
R14702 vdd.n2977 vdd.n805 185
R14703 vdd.n2979 vdd.n839 185
R14704 vdd.n2989 vdd.n839 185
R14705 vdd.n2980 vdd.n848 185
R14706 vdd.n848 vdd.n846 185
R14707 vdd.n2982 vdd.n2981 185
R14708 vdd.n2983 vdd.n2982 185
R14709 vdd.n2935 vdd.n847 185
R14710 vdd.n847 vdd.n843 185
R14711 vdd.n2934 vdd.n2933 185
R14712 vdd.n2933 vdd.n2932 185
R14713 vdd.n850 vdd.n849 185
R14714 vdd.n851 vdd.n850 185
R14715 vdd.n2925 vdd.n2924 185
R14716 vdd.n2926 vdd.n2925 185
R14717 vdd.n2921 vdd.n860 185
R14718 vdd.n860 vdd.n857 185
R14719 vdd.n2920 vdd.n2919 185
R14720 vdd.n2919 vdd.n2918 185
R14721 vdd.n862 vdd.n861 185
R14722 vdd.n870 vdd.n862 185
R14723 vdd.n2911 vdd.n2910 185
R14724 vdd.n2912 vdd.n2911 185
R14725 vdd.n2909 vdd.n871 185
R14726 vdd.n2760 vdd.n871 185
R14727 vdd.n2908 vdd.n2907 185
R14728 vdd.n2907 vdd.n2906 185
R14729 vdd.n873 vdd.n872 185
R14730 vdd.n874 vdd.n873 185
R14731 vdd.n2899 vdd.n2898 185
R14732 vdd.n2900 vdd.n2899 185
R14733 vdd.n2897 vdd.n883 185
R14734 vdd.n883 vdd.n880 185
R14735 vdd.n2896 vdd.n2895 185
R14736 vdd.n2895 vdd.n2894 185
R14737 vdd.n885 vdd.n884 185
R14738 vdd.n893 vdd.n885 185
R14739 vdd.n2887 vdd.n2886 185
R14740 vdd.n2888 vdd.n2887 185
R14741 vdd.n2885 vdd.n894 185
R14742 vdd.n900 vdd.n894 185
R14743 vdd.n2884 vdd.n2883 185
R14744 vdd.n2883 vdd.n2882 185
R14745 vdd.n896 vdd.n895 185
R14746 vdd.n897 vdd.n896 185
R14747 vdd.n2875 vdd.n2874 185
R14748 vdd.n2876 vdd.n2875 185
R14749 vdd.n2873 vdd.n906 185
R14750 vdd.n2781 vdd.n906 185
R14751 vdd.n2872 vdd.n2871 185
R14752 vdd.n2871 vdd.n2870 185
R14753 vdd.n908 vdd.n907 185
R14754 vdd.t200 vdd.n908 185
R14755 vdd.n2863 vdd.n2862 185
R14756 vdd.n2864 vdd.n2863 185
R14757 vdd.n2861 vdd.n916 185
R14758 vdd.n2860 vdd.n2859 185
R14759 vdd.n918 vdd.n917 185
R14760 vdd.n2646 vdd.n2645 185
R14761 vdd.n2648 vdd.n2647 185
R14762 vdd.n2650 vdd.n2649 185
R14763 vdd.n2652 vdd.n2651 185
R14764 vdd.n2654 vdd.n2653 185
R14765 vdd.n2656 vdd.n2655 185
R14766 vdd.n2658 vdd.n2657 185
R14767 vdd.n2660 vdd.n2659 185
R14768 vdd.n2662 vdd.n2661 185
R14769 vdd.n2664 vdd.n2663 185
R14770 vdd.n2666 vdd.n2665 185
R14771 vdd.n2668 vdd.n2667 185
R14772 vdd.n2670 vdd.n2669 185
R14773 vdd.n2672 vdd.n2671 185
R14774 vdd.n2674 vdd.n2673 185
R14775 vdd.n2676 vdd.n2675 185
R14776 vdd.n2678 vdd.n2677 185
R14777 vdd.n2680 vdd.n2679 185
R14778 vdd.n2682 vdd.n2681 185
R14779 vdd.n2684 vdd.n2683 185
R14780 vdd.n2686 vdd.n2685 185
R14781 vdd.n2688 vdd.n2687 185
R14782 vdd.n2690 vdd.n2689 185
R14783 vdd.n2692 vdd.n2691 185
R14784 vdd.n2694 vdd.n2693 185
R14785 vdd.n2696 vdd.n2695 185
R14786 vdd.n2698 vdd.n2697 185
R14787 vdd.n2700 vdd.n2699 185
R14788 vdd.n2702 vdd.n2701 185
R14789 vdd.n2704 vdd.n2703 185
R14790 vdd.n2706 vdd.n2705 185
R14791 vdd.n2707 vdd.n2637 185
R14792 vdd.n2857 vdd.n2637 185
R14793 vdd.n3062 vdd.n3061 185
R14794 vdd.n3063 vdd.n798 185
R14795 vdd.n3065 vdd.n3064 185
R14796 vdd.n3067 vdd.n796 185
R14797 vdd.n3069 vdd.n3068 185
R14798 vdd.n3070 vdd.n795 185
R14799 vdd.n3072 vdd.n3071 185
R14800 vdd.n3074 vdd.n793 185
R14801 vdd.n3076 vdd.n3075 185
R14802 vdd.n3077 vdd.n792 185
R14803 vdd.n3079 vdd.n3078 185
R14804 vdd.n3081 vdd.n790 185
R14805 vdd.n3083 vdd.n3082 185
R14806 vdd.n3084 vdd.n789 185
R14807 vdd.n3086 vdd.n3085 185
R14808 vdd.n3088 vdd.n788 185
R14809 vdd.n3089 vdd.n786 185
R14810 vdd.n3092 vdd.n3091 185
R14811 vdd.n787 vdd.n785 185
R14812 vdd.n2948 vdd.n2947 185
R14813 vdd.n2950 vdd.n2949 185
R14814 vdd.n2952 vdd.n2944 185
R14815 vdd.n2954 vdd.n2953 185
R14816 vdd.n2955 vdd.n2943 185
R14817 vdd.n2957 vdd.n2956 185
R14818 vdd.n2959 vdd.n2941 185
R14819 vdd.n2961 vdd.n2960 185
R14820 vdd.n2962 vdd.n2940 185
R14821 vdd.n2964 vdd.n2963 185
R14822 vdd.n2966 vdd.n2938 185
R14823 vdd.n2968 vdd.n2967 185
R14824 vdd.n2969 vdd.n2937 185
R14825 vdd.n2971 vdd.n2970 185
R14826 vdd.n2973 vdd.n2936 185
R14827 vdd.n2975 vdd.n2974 185
R14828 vdd.n2974 vdd.n692 185
R14829 vdd.n3060 vdd.n802 185
R14830 vdd.n3060 vdd.n3059 185
R14831 vdd.n2712 vdd.n804 185
R14832 vdd.n805 vdd.n804 185
R14833 vdd.n2713 vdd.n838 185
R14834 vdd.n2989 vdd.n838 185
R14835 vdd.n2715 vdd.n2714 185
R14836 vdd.n2714 vdd.n846 185
R14837 vdd.n2716 vdd.n845 185
R14838 vdd.n2983 vdd.n845 185
R14839 vdd.n2718 vdd.n2717 185
R14840 vdd.n2717 vdd.n843 185
R14841 vdd.n2719 vdd.n853 185
R14842 vdd.n2932 vdd.n853 185
R14843 vdd.n2721 vdd.n2720 185
R14844 vdd.n2720 vdd.n851 185
R14845 vdd.n2722 vdd.n859 185
R14846 vdd.n2926 vdd.n859 185
R14847 vdd.n2724 vdd.n2723 185
R14848 vdd.n2723 vdd.n857 185
R14849 vdd.n2725 vdd.n864 185
R14850 vdd.n2918 vdd.n864 185
R14851 vdd.n2727 vdd.n2726 185
R14852 vdd.n2726 vdd.n870 185
R14853 vdd.n2728 vdd.n869 185
R14854 vdd.n2912 vdd.n869 185
R14855 vdd.n2762 vdd.n2761 185
R14856 vdd.n2761 vdd.n2760 185
R14857 vdd.n2763 vdd.n876 185
R14858 vdd.n2906 vdd.n876 185
R14859 vdd.n2765 vdd.n2764 185
R14860 vdd.n2764 vdd.n874 185
R14861 vdd.n2766 vdd.n882 185
R14862 vdd.n2900 vdd.n882 185
R14863 vdd.n2768 vdd.n2767 185
R14864 vdd.n2767 vdd.n880 185
R14865 vdd.n2769 vdd.n887 185
R14866 vdd.n2894 vdd.n887 185
R14867 vdd.n2771 vdd.n2770 185
R14868 vdd.n2770 vdd.n893 185
R14869 vdd.n2772 vdd.n892 185
R14870 vdd.n2888 vdd.n892 185
R14871 vdd.n2774 vdd.n2773 185
R14872 vdd.n2773 vdd.n900 185
R14873 vdd.n2775 vdd.n899 185
R14874 vdd.n2882 vdd.n899 185
R14875 vdd.n2777 vdd.n2776 185
R14876 vdd.n2776 vdd.n897 185
R14877 vdd.n2778 vdd.n905 185
R14878 vdd.n2876 vdd.n905 185
R14879 vdd.n2780 vdd.n2779 185
R14880 vdd.n2781 vdd.n2780 185
R14881 vdd.n2711 vdd.n910 185
R14882 vdd.n2870 vdd.n910 185
R14883 vdd.n2710 vdd.n2709 185
R14884 vdd.n2709 vdd.t200 185
R14885 vdd.n2708 vdd.n915 185
R14886 vdd.n2864 vdd.n915 185
R14887 vdd.n2328 vdd.n2327 185
R14888 vdd.n2329 vdd.n2328 185
R14889 vdd.n1076 vdd.n1074 185
R14890 vdd.n1894 vdd.n1074 185
R14891 vdd.n1897 vdd.n1896 185
R14892 vdd.n1896 vdd.n1895 185
R14893 vdd.n1079 vdd.n1078 185
R14894 vdd.n1080 vdd.n1079 185
R14895 vdd.n1883 vdd.n1882 185
R14896 vdd.n1884 vdd.n1883 185
R14897 vdd.n1088 vdd.n1087 185
R14898 vdd.n1875 vdd.n1087 185
R14899 vdd.n1878 vdd.n1877 185
R14900 vdd.n1877 vdd.n1876 185
R14901 vdd.n1091 vdd.n1090 185
R14902 vdd.n1098 vdd.n1091 185
R14903 vdd.n1866 vdd.n1865 185
R14904 vdd.n1867 vdd.n1866 185
R14905 vdd.n1100 vdd.n1099 185
R14906 vdd.n1099 vdd.n1097 185
R14907 vdd.n1861 vdd.n1860 185
R14908 vdd.n1860 vdd.n1859 185
R14909 vdd.n1103 vdd.n1102 185
R14910 vdd.n1104 vdd.n1103 185
R14911 vdd.n1850 vdd.n1849 185
R14912 vdd.n1851 vdd.n1850 185
R14913 vdd.n1111 vdd.n1110 185
R14914 vdd.n1842 vdd.n1110 185
R14915 vdd.n1845 vdd.n1844 185
R14916 vdd.n1844 vdd.n1843 185
R14917 vdd.n1114 vdd.n1113 185
R14918 vdd.n1120 vdd.n1114 185
R14919 vdd.n1833 vdd.n1832 185
R14920 vdd.n1834 vdd.n1833 185
R14921 vdd.n1122 vdd.n1121 185
R14922 vdd.n1825 vdd.n1121 185
R14923 vdd.n1828 vdd.n1827 185
R14924 vdd.n1827 vdd.n1826 185
R14925 vdd.n1125 vdd.n1124 185
R14926 vdd.n1126 vdd.n1125 185
R14927 vdd.n1816 vdd.n1815 185
R14928 vdd.n1817 vdd.n1816 185
R14929 vdd.n1134 vdd.n1133 185
R14930 vdd.n1133 vdd.n1132 185
R14931 vdd.n1504 vdd.n1503 185
R14932 vdd.n1503 vdd.n1502 185
R14933 vdd.n1137 vdd.n1136 185
R14934 vdd.n1143 vdd.n1137 185
R14935 vdd.n1493 vdd.n1492 185
R14936 vdd.n1494 vdd.n1493 185
R14937 vdd.n1145 vdd.n1144 185
R14938 vdd.n1485 vdd.n1144 185
R14939 vdd.n1488 vdd.n1487 185
R14940 vdd.n1487 vdd.n1486 185
R14941 vdd.n1148 vdd.n1147 185
R14942 vdd.n1155 vdd.n1148 185
R14943 vdd.n1476 vdd.n1475 185
R14944 vdd.n1477 vdd.n1476 185
R14945 vdd.n1157 vdd.n1156 185
R14946 vdd.n1156 vdd.n1154 185
R14947 vdd.n1471 vdd.n1470 185
R14948 vdd.n1470 vdd.n1469 185
R14949 vdd.n1160 vdd.n1159 185
R14950 vdd.n1161 vdd.n1160 185
R14951 vdd.n1460 vdd.n1459 185
R14952 vdd.n1461 vdd.n1460 185
R14953 vdd.n1168 vdd.n1167 185
R14954 vdd.n1452 vdd.n1167 185
R14955 vdd.n1455 vdd.n1454 185
R14956 vdd.n1454 vdd.n1453 185
R14957 vdd.n1171 vdd.n1170 185
R14958 vdd.n1177 vdd.n1171 185
R14959 vdd.n1443 vdd.n1442 185
R14960 vdd.n1444 vdd.n1443 185
R14961 vdd.n1179 vdd.n1178 185
R14962 vdd.n1435 vdd.n1178 185
R14963 vdd.n1438 vdd.n1437 185
R14964 vdd.n1437 vdd.n1436 185
R14965 vdd.n1182 vdd.n1181 185
R14966 vdd.n1183 vdd.n1182 185
R14967 vdd.n1426 vdd.n1425 185
R14968 vdd.n1427 vdd.n1426 185
R14969 vdd.n1190 vdd.n1189 185
R14970 vdd.n1225 vdd.n1189 185
R14971 vdd.n1421 vdd.n1420 185
R14972 vdd.n1193 vdd.n1192 185
R14973 vdd.n1417 vdd.n1416 185
R14974 vdd.n1418 vdd.n1417 185
R14975 vdd.n1227 vdd.n1226 185
R14976 vdd.n1412 vdd.n1229 185
R14977 vdd.n1411 vdd.n1230 185
R14978 vdd.n1410 vdd.n1231 185
R14979 vdd.n1233 vdd.n1232 185
R14980 vdd.n1406 vdd.n1235 185
R14981 vdd.n1405 vdd.n1236 185
R14982 vdd.n1404 vdd.n1237 185
R14983 vdd.n1239 vdd.n1238 185
R14984 vdd.n1400 vdd.n1241 185
R14985 vdd.n1399 vdd.n1242 185
R14986 vdd.n1398 vdd.n1243 185
R14987 vdd.n1245 vdd.n1244 185
R14988 vdd.n1394 vdd.n1247 185
R14989 vdd.n1393 vdd.n1248 185
R14990 vdd.n1392 vdd.n1249 185
R14991 vdd.n1253 vdd.n1250 185
R14992 vdd.n1388 vdd.n1255 185
R14993 vdd.n1387 vdd.n1256 185
R14994 vdd.n1386 vdd.n1257 185
R14995 vdd.n1259 vdd.n1258 185
R14996 vdd.n1382 vdd.n1261 185
R14997 vdd.n1381 vdd.n1262 185
R14998 vdd.n1380 vdd.n1263 185
R14999 vdd.n1265 vdd.n1264 185
R15000 vdd.n1376 vdd.n1267 185
R15001 vdd.n1375 vdd.n1268 185
R15002 vdd.n1374 vdd.n1269 185
R15003 vdd.n1271 vdd.n1270 185
R15004 vdd.n1370 vdd.n1273 185
R15005 vdd.n1369 vdd.n1274 185
R15006 vdd.n1368 vdd.n1275 185
R15007 vdd.n1277 vdd.n1276 185
R15008 vdd.n1364 vdd.n1279 185
R15009 vdd.n1363 vdd.n1280 185
R15010 vdd.n1362 vdd.n1281 185
R15011 vdd.n1283 vdd.n1282 185
R15012 vdd.n1358 vdd.n1285 185
R15013 vdd.n1357 vdd.n1354 185
R15014 vdd.n1353 vdd.n1286 185
R15015 vdd.n1288 vdd.n1287 185
R15016 vdd.n1349 vdd.n1290 185
R15017 vdd.n1348 vdd.n1291 185
R15018 vdd.n1347 vdd.n1292 185
R15019 vdd.n1294 vdd.n1293 185
R15020 vdd.n1343 vdd.n1296 185
R15021 vdd.n1342 vdd.n1297 185
R15022 vdd.n1341 vdd.n1298 185
R15023 vdd.n1300 vdd.n1299 185
R15024 vdd.n1337 vdd.n1302 185
R15025 vdd.n1336 vdd.n1303 185
R15026 vdd.n1335 vdd.n1304 185
R15027 vdd.n1306 vdd.n1305 185
R15028 vdd.n1331 vdd.n1308 185
R15029 vdd.n1330 vdd.n1309 185
R15030 vdd.n1329 vdd.n1310 185
R15031 vdd.n1312 vdd.n1311 185
R15032 vdd.n1325 vdd.n1314 185
R15033 vdd.n1324 vdd.n1315 185
R15034 vdd.n1323 vdd.n1316 185
R15035 vdd.n1320 vdd.n1224 185
R15036 vdd.n1418 vdd.n1224 185
R15037 vdd.n2332 vdd.n2331 185
R15038 vdd.n2336 vdd.n1069 185
R15039 vdd.n1999 vdd.n1068 185
R15040 vdd.n2002 vdd.n2001 185
R15041 vdd.n2004 vdd.n2003 185
R15042 vdd.n2007 vdd.n2006 185
R15043 vdd.n2009 vdd.n2008 185
R15044 vdd.n2011 vdd.n1997 185
R15045 vdd.n2013 vdd.n2012 185
R15046 vdd.n2014 vdd.n1991 185
R15047 vdd.n2016 vdd.n2015 185
R15048 vdd.n2018 vdd.n1989 185
R15049 vdd.n2020 vdd.n2019 185
R15050 vdd.n2021 vdd.n1984 185
R15051 vdd.n2023 vdd.n2022 185
R15052 vdd.n2025 vdd.n1982 185
R15053 vdd.n2027 vdd.n2026 185
R15054 vdd.n2028 vdd.n1978 185
R15055 vdd.n2030 vdd.n2029 185
R15056 vdd.n2032 vdd.n1975 185
R15057 vdd.n2034 vdd.n2033 185
R15058 vdd.n1976 vdd.n1969 185
R15059 vdd.n2038 vdd.n1973 185
R15060 vdd.n2039 vdd.n1965 185
R15061 vdd.n2041 vdd.n2040 185
R15062 vdd.n2043 vdd.n1963 185
R15063 vdd.n2045 vdd.n2044 185
R15064 vdd.n2046 vdd.n1958 185
R15065 vdd.n2048 vdd.n2047 185
R15066 vdd.n2050 vdd.n1956 185
R15067 vdd.n2052 vdd.n2051 185
R15068 vdd.n2053 vdd.n1951 185
R15069 vdd.n2055 vdd.n2054 185
R15070 vdd.n2057 vdd.n1949 185
R15071 vdd.n2059 vdd.n2058 185
R15072 vdd.n2060 vdd.n1944 185
R15073 vdd.n2062 vdd.n2061 185
R15074 vdd.n2064 vdd.n1942 185
R15075 vdd.n2066 vdd.n2065 185
R15076 vdd.n2067 vdd.n1938 185
R15077 vdd.n2069 vdd.n2068 185
R15078 vdd.n2071 vdd.n1935 185
R15079 vdd.n2073 vdd.n2072 185
R15080 vdd.n1936 vdd.n1929 185
R15081 vdd.n2077 vdd.n1933 185
R15082 vdd.n2078 vdd.n1925 185
R15083 vdd.n2080 vdd.n2079 185
R15084 vdd.n2082 vdd.n1923 185
R15085 vdd.n2084 vdd.n2083 185
R15086 vdd.n2085 vdd.n1918 185
R15087 vdd.n2087 vdd.n2086 185
R15088 vdd.n2089 vdd.n1916 185
R15089 vdd.n2091 vdd.n2090 185
R15090 vdd.n2092 vdd.n1911 185
R15091 vdd.n2094 vdd.n2093 185
R15092 vdd.n2096 vdd.n1910 185
R15093 vdd.n2097 vdd.n1907 185
R15094 vdd.n2100 vdd.n2099 185
R15095 vdd.n1909 vdd.n1905 185
R15096 vdd.n2317 vdd.n1903 185
R15097 vdd.n2319 vdd.n2318 185
R15098 vdd.n2321 vdd.n1901 185
R15099 vdd.n2323 vdd.n2322 185
R15100 vdd.n2324 vdd.n1075 185
R15101 vdd.n2330 vdd.n1072 185
R15102 vdd.n2330 vdd.n2329 185
R15103 vdd.n1083 vdd.n1071 185
R15104 vdd.n1894 vdd.n1071 185
R15105 vdd.n1893 vdd.n1892 185
R15106 vdd.n1895 vdd.n1893 185
R15107 vdd.n1082 vdd.n1081 185
R15108 vdd.n1081 vdd.n1080 185
R15109 vdd.n1886 vdd.n1885 185
R15110 vdd.n1885 vdd.n1884 185
R15111 vdd.n1086 vdd.n1085 185
R15112 vdd.n1875 vdd.n1086 185
R15113 vdd.n1874 vdd.n1873 185
R15114 vdd.n1876 vdd.n1874 185
R15115 vdd.n1093 vdd.n1092 185
R15116 vdd.n1098 vdd.n1092 185
R15117 vdd.n1869 vdd.n1868 185
R15118 vdd.n1868 vdd.n1867 185
R15119 vdd.n1096 vdd.n1095 185
R15120 vdd.n1097 vdd.n1096 185
R15121 vdd.n1858 vdd.n1857 185
R15122 vdd.n1859 vdd.n1858 185
R15123 vdd.n1106 vdd.n1105 185
R15124 vdd.n1105 vdd.n1104 185
R15125 vdd.n1853 vdd.n1852 185
R15126 vdd.n1852 vdd.n1851 185
R15127 vdd.n1109 vdd.n1108 185
R15128 vdd.n1842 vdd.n1109 185
R15129 vdd.n1841 vdd.n1840 185
R15130 vdd.n1843 vdd.n1841 185
R15131 vdd.n1116 vdd.n1115 185
R15132 vdd.n1120 vdd.n1115 185
R15133 vdd.n1836 vdd.n1835 185
R15134 vdd.n1835 vdd.n1834 185
R15135 vdd.n1119 vdd.n1118 185
R15136 vdd.n1825 vdd.n1119 185
R15137 vdd.n1824 vdd.n1823 185
R15138 vdd.n1826 vdd.n1824 185
R15139 vdd.n1128 vdd.n1127 185
R15140 vdd.n1127 vdd.n1126 185
R15141 vdd.n1819 vdd.n1818 185
R15142 vdd.n1818 vdd.n1817 185
R15143 vdd.n1131 vdd.n1130 185
R15144 vdd.n1132 vdd.n1131 185
R15145 vdd.n1501 vdd.n1500 185
R15146 vdd.n1502 vdd.n1501 185
R15147 vdd.n1139 vdd.n1138 185
R15148 vdd.n1143 vdd.n1138 185
R15149 vdd.n1496 vdd.n1495 185
R15150 vdd.n1495 vdd.n1494 185
R15151 vdd.n1142 vdd.n1141 185
R15152 vdd.n1485 vdd.n1142 185
R15153 vdd.n1484 vdd.n1483 185
R15154 vdd.n1486 vdd.n1484 185
R15155 vdd.n1150 vdd.n1149 185
R15156 vdd.n1155 vdd.n1149 185
R15157 vdd.n1479 vdd.n1478 185
R15158 vdd.n1478 vdd.n1477 185
R15159 vdd.n1153 vdd.n1152 185
R15160 vdd.n1154 vdd.n1153 185
R15161 vdd.n1468 vdd.n1467 185
R15162 vdd.n1469 vdd.n1468 185
R15163 vdd.n1163 vdd.n1162 185
R15164 vdd.n1162 vdd.n1161 185
R15165 vdd.n1463 vdd.n1462 185
R15166 vdd.n1462 vdd.n1461 185
R15167 vdd.n1166 vdd.n1165 185
R15168 vdd.n1452 vdd.n1166 185
R15169 vdd.n1451 vdd.n1450 185
R15170 vdd.n1453 vdd.n1451 185
R15171 vdd.n1173 vdd.n1172 185
R15172 vdd.n1177 vdd.n1172 185
R15173 vdd.n1446 vdd.n1445 185
R15174 vdd.n1445 vdd.n1444 185
R15175 vdd.n1176 vdd.n1175 185
R15176 vdd.n1435 vdd.n1176 185
R15177 vdd.n1434 vdd.n1433 185
R15178 vdd.n1436 vdd.n1434 185
R15179 vdd.n1185 vdd.n1184 185
R15180 vdd.n1184 vdd.n1183 185
R15181 vdd.n1429 vdd.n1428 185
R15182 vdd.n1428 vdd.n1427 185
R15183 vdd.n1188 vdd.n1187 185
R15184 vdd.n1225 vdd.n1188 185
R15185 vdd.n956 vdd.n954 185
R15186 vdd.n2532 vdd.n954 185
R15187 vdd.n2454 vdd.n973 185
R15188 vdd.n973 vdd.t292 185
R15189 vdd.n2456 vdd.n2455 185
R15190 vdd.n2457 vdd.n2456 185
R15191 vdd.n2453 vdd.n972 185
R15192 vdd.n2156 vdd.n972 185
R15193 vdd.n2452 vdd.n2451 185
R15194 vdd.n2451 vdd.n2450 185
R15195 vdd.n975 vdd.n974 185
R15196 vdd.n976 vdd.n975 185
R15197 vdd.n2441 vdd.n2440 185
R15198 vdd.n2442 vdd.n2441 185
R15199 vdd.n2439 vdd.n986 185
R15200 vdd.n986 vdd.n983 185
R15201 vdd.n2438 vdd.n2437 185
R15202 vdd.n2437 vdd.n2436 185
R15203 vdd.n988 vdd.n987 185
R15204 vdd.n989 vdd.n988 185
R15205 vdd.n2429 vdd.n2428 185
R15206 vdd.n2430 vdd.n2429 185
R15207 vdd.n2427 vdd.n997 185
R15208 vdd.n1002 vdd.n997 185
R15209 vdd.n2426 vdd.n2425 185
R15210 vdd.n2425 vdd.n2424 185
R15211 vdd.n999 vdd.n998 185
R15212 vdd.n1008 vdd.n999 185
R15213 vdd.n2417 vdd.n2416 185
R15214 vdd.n2418 vdd.n2417 185
R15215 vdd.n2415 vdd.n1009 185
R15216 vdd.n2257 vdd.n1009 185
R15217 vdd.n2414 vdd.n2413 185
R15218 vdd.n2413 vdd.n2412 185
R15219 vdd.n1011 vdd.n1010 185
R15220 vdd.n1012 vdd.n1011 185
R15221 vdd.n2405 vdd.n2404 185
R15222 vdd.n2406 vdd.n2405 185
R15223 vdd.n2403 vdd.n1021 185
R15224 vdd.n1021 vdd.n1018 185
R15225 vdd.n2402 vdd.n2401 185
R15226 vdd.n2401 vdd.n2400 185
R15227 vdd.n1023 vdd.n1022 185
R15228 vdd.n1033 vdd.n1023 185
R15229 vdd.n2392 vdd.n2391 185
R15230 vdd.n2393 vdd.n2392 185
R15231 vdd.n2390 vdd.n1034 185
R15232 vdd.n1034 vdd.n1030 185
R15233 vdd.n2389 vdd.n2388 185
R15234 vdd.n2388 vdd.n2387 185
R15235 vdd.n1036 vdd.n1035 185
R15236 vdd.n1037 vdd.n1036 185
R15237 vdd.n2380 vdd.n2379 185
R15238 vdd.n2381 vdd.n2380 185
R15239 vdd.n2378 vdd.n1046 185
R15240 vdd.n1046 vdd.n1043 185
R15241 vdd.n2377 vdd.n2376 185
R15242 vdd.n2376 vdd.n2375 185
R15243 vdd.n1048 vdd.n1047 185
R15244 vdd.n2112 vdd.n2111 185
R15245 vdd.n2113 vdd.n2109 185
R15246 vdd.n2109 vdd.n1049 185
R15247 vdd.n2115 vdd.n2114 185
R15248 vdd.n2117 vdd.n2108 185
R15249 vdd.n2120 vdd.n2119 185
R15250 vdd.n2121 vdd.n2107 185
R15251 vdd.n2123 vdd.n2122 185
R15252 vdd.n2125 vdd.n2106 185
R15253 vdd.n2128 vdd.n2127 185
R15254 vdd.n2129 vdd.n2105 185
R15255 vdd.n2131 vdd.n2130 185
R15256 vdd.n2133 vdd.n2104 185
R15257 vdd.n2136 vdd.n2135 185
R15258 vdd.n2137 vdd.n2103 185
R15259 vdd.n2139 vdd.n2138 185
R15260 vdd.n2141 vdd.n2102 185
R15261 vdd.n2314 vdd.n2142 185
R15262 vdd.n2313 vdd.n2312 185
R15263 vdd.n2310 vdd.n2143 185
R15264 vdd.n2308 vdd.n2307 185
R15265 vdd.n2306 vdd.n2144 185
R15266 vdd.n2305 vdd.n2304 185
R15267 vdd.n2302 vdd.n2145 185
R15268 vdd.n2300 vdd.n2299 185
R15269 vdd.n2298 vdd.n2146 185
R15270 vdd.n2297 vdd.n2296 185
R15271 vdd.n2294 vdd.n2147 185
R15272 vdd.n2292 vdd.n2291 185
R15273 vdd.n2290 vdd.n2148 185
R15274 vdd.n2289 vdd.n2288 185
R15275 vdd.n2286 vdd.n2149 185
R15276 vdd.n2284 vdd.n2283 185
R15277 vdd.n2282 vdd.n2150 185
R15278 vdd.n2281 vdd.n2280 185
R15279 vdd.n2535 vdd.n2534 185
R15280 vdd.n2537 vdd.n2536 185
R15281 vdd.n2539 vdd.n2538 185
R15282 vdd.n2542 vdd.n2541 185
R15283 vdd.n2544 vdd.n2543 185
R15284 vdd.n2546 vdd.n2545 185
R15285 vdd.n2548 vdd.n2547 185
R15286 vdd.n2550 vdd.n2549 185
R15287 vdd.n2552 vdd.n2551 185
R15288 vdd.n2554 vdd.n2553 185
R15289 vdd.n2556 vdd.n2555 185
R15290 vdd.n2558 vdd.n2557 185
R15291 vdd.n2560 vdd.n2559 185
R15292 vdd.n2562 vdd.n2561 185
R15293 vdd.n2564 vdd.n2563 185
R15294 vdd.n2566 vdd.n2565 185
R15295 vdd.n2568 vdd.n2567 185
R15296 vdd.n2570 vdd.n2569 185
R15297 vdd.n2572 vdd.n2571 185
R15298 vdd.n2574 vdd.n2573 185
R15299 vdd.n2576 vdd.n2575 185
R15300 vdd.n2578 vdd.n2577 185
R15301 vdd.n2580 vdd.n2579 185
R15302 vdd.n2582 vdd.n2581 185
R15303 vdd.n2584 vdd.n2583 185
R15304 vdd.n2586 vdd.n2585 185
R15305 vdd.n2588 vdd.n2587 185
R15306 vdd.n2590 vdd.n2589 185
R15307 vdd.n2592 vdd.n2591 185
R15308 vdd.n2594 vdd.n2593 185
R15309 vdd.n2596 vdd.n2595 185
R15310 vdd.n2598 vdd.n2597 185
R15311 vdd.n2600 vdd.n2599 185
R15312 vdd.n2601 vdd.n955 185
R15313 vdd.n2603 vdd.n2602 185
R15314 vdd.n2604 vdd.n2603 185
R15315 vdd.n2533 vdd.n959 185
R15316 vdd.n2533 vdd.n2532 185
R15317 vdd.n2154 vdd.n960 185
R15318 vdd.t292 vdd.n960 185
R15319 vdd.n2155 vdd.n970 185
R15320 vdd.n2457 vdd.n970 185
R15321 vdd.n2158 vdd.n2157 185
R15322 vdd.n2157 vdd.n2156 185
R15323 vdd.n2159 vdd.n977 185
R15324 vdd.n2450 vdd.n977 185
R15325 vdd.n2161 vdd.n2160 185
R15326 vdd.n2160 vdd.n976 185
R15327 vdd.n2162 vdd.n984 185
R15328 vdd.n2442 vdd.n984 185
R15329 vdd.n2164 vdd.n2163 185
R15330 vdd.n2163 vdd.n983 185
R15331 vdd.n2165 vdd.n990 185
R15332 vdd.n2436 vdd.n990 185
R15333 vdd.n2167 vdd.n2166 185
R15334 vdd.n2166 vdd.n989 185
R15335 vdd.n2168 vdd.n995 185
R15336 vdd.n2430 vdd.n995 185
R15337 vdd.n2170 vdd.n2169 185
R15338 vdd.n2169 vdd.n1002 185
R15339 vdd.n2171 vdd.n1000 185
R15340 vdd.n2424 vdd.n1000 185
R15341 vdd.n2173 vdd.n2172 185
R15342 vdd.n2172 vdd.n1008 185
R15343 vdd.n2174 vdd.n1006 185
R15344 vdd.n2418 vdd.n1006 185
R15345 vdd.n2259 vdd.n2258 185
R15346 vdd.n2258 vdd.n2257 185
R15347 vdd.n2260 vdd.n1013 185
R15348 vdd.n2412 vdd.n1013 185
R15349 vdd.n2262 vdd.n2261 185
R15350 vdd.n2261 vdd.n1012 185
R15351 vdd.n2263 vdd.n1019 185
R15352 vdd.n2406 vdd.n1019 185
R15353 vdd.n2265 vdd.n2264 185
R15354 vdd.n2264 vdd.n1018 185
R15355 vdd.n2266 vdd.n1024 185
R15356 vdd.n2400 vdd.n1024 185
R15357 vdd.n2268 vdd.n2267 185
R15358 vdd.n2267 vdd.n1033 185
R15359 vdd.n2269 vdd.n1031 185
R15360 vdd.n2393 vdd.n1031 185
R15361 vdd.n2271 vdd.n2270 185
R15362 vdd.n2270 vdd.n1030 185
R15363 vdd.n2272 vdd.n1038 185
R15364 vdd.n2387 vdd.n1038 185
R15365 vdd.n2274 vdd.n2273 185
R15366 vdd.n2273 vdd.n1037 185
R15367 vdd.n2275 vdd.n1044 185
R15368 vdd.n2381 vdd.n1044 185
R15369 vdd.n2277 vdd.n2276 185
R15370 vdd.n2276 vdd.n1043 185
R15371 vdd.n2278 vdd.n1050 185
R15372 vdd.n2375 vdd.n1050 185
R15373 vdd.n3357 vdd.n3356 185
R15374 vdd.n3356 vdd.n3355 185
R15375 vdd.n3358 vdd.n387 185
R15376 vdd.n387 vdd.n386 185
R15377 vdd.n3360 vdd.n3359 185
R15378 vdd.n3361 vdd.n3360 185
R15379 vdd.n382 vdd.n381 185
R15380 vdd.n3362 vdd.n382 185
R15381 vdd.n3365 vdd.n3364 185
R15382 vdd.n3364 vdd.n3363 185
R15383 vdd.n3366 vdd.n376 185
R15384 vdd.n376 vdd.n375 185
R15385 vdd.n3368 vdd.n3367 185
R15386 vdd.n3369 vdd.n3368 185
R15387 vdd.n371 vdd.n370 185
R15388 vdd.n3370 vdd.n371 185
R15389 vdd.n3373 vdd.n3372 185
R15390 vdd.n3372 vdd.n3371 185
R15391 vdd.n3374 vdd.n365 185
R15392 vdd.n3331 vdd.n365 185
R15393 vdd.n3376 vdd.n3375 185
R15394 vdd.n3377 vdd.n3376 185
R15395 vdd.n360 vdd.n359 185
R15396 vdd.n3378 vdd.n360 185
R15397 vdd.n3381 vdd.n3380 185
R15398 vdd.n3380 vdd.n3379 185
R15399 vdd.n3382 vdd.n354 185
R15400 vdd.n361 vdd.n354 185
R15401 vdd.n3384 vdd.n3383 185
R15402 vdd.n3385 vdd.n3384 185
R15403 vdd.n350 vdd.n349 185
R15404 vdd.n3386 vdd.n350 185
R15405 vdd.n3389 vdd.n3388 185
R15406 vdd.n3388 vdd.n3387 185
R15407 vdd.n3390 vdd.n345 185
R15408 vdd.n345 vdd.n344 185
R15409 vdd.n3392 vdd.n3391 185
R15410 vdd.n3393 vdd.n3392 185
R15411 vdd.n339 vdd.n337 185
R15412 vdd.n3394 vdd.n339 185
R15413 vdd.n3397 vdd.n3396 185
R15414 vdd.n3396 vdd.n3395 185
R15415 vdd.n338 vdd.n336 185
R15416 vdd.n340 vdd.n338 185
R15417 vdd.n3307 vdd.n3306 185
R15418 vdd.n3308 vdd.n3307 185
R15419 vdd.n635 vdd.n634 185
R15420 vdd.n634 vdd.n633 185
R15421 vdd.n3302 vdd.n3301 185
R15422 vdd.n3301 vdd.n3300 185
R15423 vdd.n638 vdd.n637 185
R15424 vdd.n644 vdd.n638 185
R15425 vdd.n3288 vdd.n3287 185
R15426 vdd.n3289 vdd.n3288 185
R15427 vdd.n646 vdd.n645 185
R15428 vdd.n3280 vdd.n645 185
R15429 vdd.n3283 vdd.n3282 185
R15430 vdd.n3282 vdd.n3281 185
R15431 vdd.n649 vdd.n648 185
R15432 vdd.n656 vdd.n649 185
R15433 vdd.n3271 vdd.n3270 185
R15434 vdd.n3272 vdd.n3271 185
R15435 vdd.n658 vdd.n657 185
R15436 vdd.n657 vdd.n655 185
R15437 vdd.n3266 vdd.n3265 185
R15438 vdd.n3265 vdd.n3264 185
R15439 vdd.n661 vdd.n660 185
R15440 vdd.n662 vdd.n661 185
R15441 vdd.n3255 vdd.n3254 185
R15442 vdd.n3256 vdd.n3255 185
R15443 vdd.n669 vdd.n668 185
R15444 vdd.n3247 vdd.n668 185
R15445 vdd.n3250 vdd.n3249 185
R15446 vdd.n3249 vdd.n3248 185
R15447 vdd.n672 vdd.n671 185
R15448 vdd.n679 vdd.n672 185
R15449 vdd.n3238 vdd.n3237 185
R15450 vdd.n3239 vdd.n3238 185
R15451 vdd.n681 vdd.n680 185
R15452 vdd.n680 vdd.n678 185
R15453 vdd.n3233 vdd.n3232 185
R15454 vdd.n3232 vdd.n3231 185
R15455 vdd.n684 vdd.n683 185
R15456 vdd.n723 vdd.n684 185
R15457 vdd.n3221 vdd.n3220 185
R15458 vdd.n3219 vdd.n725 185
R15459 vdd.n3218 vdd.n724 185
R15460 vdd.n3223 vdd.n724 185
R15461 vdd.n729 vdd.n728 185
R15462 vdd.n733 vdd.n732 185
R15463 vdd.n3214 vdd.n734 185
R15464 vdd.n3213 vdd.n3212 185
R15465 vdd.n3211 vdd.n3210 185
R15466 vdd.n3209 vdd.n3208 185
R15467 vdd.n3207 vdd.n3206 185
R15468 vdd.n3205 vdd.n3204 185
R15469 vdd.n3203 vdd.n3202 185
R15470 vdd.n3201 vdd.n3200 185
R15471 vdd.n3199 vdd.n3198 185
R15472 vdd.n3197 vdd.n3196 185
R15473 vdd.n3195 vdd.n3194 185
R15474 vdd.n3193 vdd.n3192 185
R15475 vdd.n3191 vdd.n3190 185
R15476 vdd.n3189 vdd.n3188 185
R15477 vdd.n3187 vdd.n3186 185
R15478 vdd.n3178 vdd.n747 185
R15479 vdd.n3180 vdd.n3179 185
R15480 vdd.n3177 vdd.n3176 185
R15481 vdd.n3175 vdd.n3174 185
R15482 vdd.n3173 vdd.n3172 185
R15483 vdd.n3171 vdd.n3170 185
R15484 vdd.n3169 vdd.n3168 185
R15485 vdd.n3167 vdd.n3166 185
R15486 vdd.n3165 vdd.n3164 185
R15487 vdd.n3163 vdd.n3162 185
R15488 vdd.n3161 vdd.n3160 185
R15489 vdd.n3159 vdd.n3158 185
R15490 vdd.n3157 vdd.n3156 185
R15491 vdd.n3155 vdd.n3154 185
R15492 vdd.n3153 vdd.n3152 185
R15493 vdd.n3151 vdd.n3150 185
R15494 vdd.n3149 vdd.n3148 185
R15495 vdd.n3147 vdd.n3146 185
R15496 vdd.n3145 vdd.n3144 185
R15497 vdd.n3143 vdd.n3142 185
R15498 vdd.n3141 vdd.n3140 185
R15499 vdd.n3139 vdd.n3138 185
R15500 vdd.n3132 vdd.n767 185
R15501 vdd.n3134 vdd.n3133 185
R15502 vdd.n3131 vdd.n3130 185
R15503 vdd.n3129 vdd.n3128 185
R15504 vdd.n3127 vdd.n3126 185
R15505 vdd.n3125 vdd.n3124 185
R15506 vdd.n3123 vdd.n3122 185
R15507 vdd.n3121 vdd.n3120 185
R15508 vdd.n3119 vdd.n3118 185
R15509 vdd.n3117 vdd.n3116 185
R15510 vdd.n3115 vdd.n3114 185
R15511 vdd.n3113 vdd.n3112 185
R15512 vdd.n3111 vdd.n3110 185
R15513 vdd.n3109 vdd.n3108 185
R15514 vdd.n3107 vdd.n3106 185
R15515 vdd.n3105 vdd.n3104 185
R15516 vdd.n3103 vdd.n3102 185
R15517 vdd.n3101 vdd.n3100 185
R15518 vdd.n3099 vdd.n3098 185
R15519 vdd.n3097 vdd.n3096 185
R15520 vdd.n3095 vdd.n691 185
R15521 vdd.n3225 vdd.n3224 185
R15522 vdd.n3224 vdd.n3223 185
R15523 vdd.n3352 vdd.n3351 185
R15524 vdd.n618 vdd.n425 185
R15525 vdd.n617 vdd.n616 185
R15526 vdd.n615 vdd.n614 185
R15527 vdd.n613 vdd.n430 185
R15528 vdd.n609 vdd.n608 185
R15529 vdd.n607 vdd.n606 185
R15530 vdd.n605 vdd.n604 185
R15531 vdd.n603 vdd.n432 185
R15532 vdd.n599 vdd.n598 185
R15533 vdd.n597 vdd.n596 185
R15534 vdd.n595 vdd.n594 185
R15535 vdd.n593 vdd.n434 185
R15536 vdd.n589 vdd.n588 185
R15537 vdd.n587 vdd.n586 185
R15538 vdd.n585 vdd.n584 185
R15539 vdd.n583 vdd.n436 185
R15540 vdd.n579 vdd.n578 185
R15541 vdd.n577 vdd.n576 185
R15542 vdd.n575 vdd.n574 185
R15543 vdd.n573 vdd.n438 185
R15544 vdd.n569 vdd.n568 185
R15545 vdd.n567 vdd.n566 185
R15546 vdd.n565 vdd.n564 185
R15547 vdd.n563 vdd.n442 185
R15548 vdd.n559 vdd.n558 185
R15549 vdd.n557 vdd.n556 185
R15550 vdd.n555 vdd.n554 185
R15551 vdd.n553 vdd.n444 185
R15552 vdd.n549 vdd.n548 185
R15553 vdd.n547 vdd.n546 185
R15554 vdd.n545 vdd.n544 185
R15555 vdd.n543 vdd.n446 185
R15556 vdd.n539 vdd.n538 185
R15557 vdd.n537 vdd.n536 185
R15558 vdd.n535 vdd.n534 185
R15559 vdd.n533 vdd.n448 185
R15560 vdd.n529 vdd.n528 185
R15561 vdd.n527 vdd.n526 185
R15562 vdd.n525 vdd.n524 185
R15563 vdd.n523 vdd.n450 185
R15564 vdd.n519 vdd.n518 185
R15565 vdd.n517 vdd.n516 185
R15566 vdd.n515 vdd.n514 185
R15567 vdd.n513 vdd.n454 185
R15568 vdd.n509 vdd.n508 185
R15569 vdd.n507 vdd.n506 185
R15570 vdd.n505 vdd.n504 185
R15571 vdd.n503 vdd.n456 185
R15572 vdd.n499 vdd.n498 185
R15573 vdd.n497 vdd.n496 185
R15574 vdd.n495 vdd.n494 185
R15575 vdd.n493 vdd.n458 185
R15576 vdd.n489 vdd.n488 185
R15577 vdd.n487 vdd.n486 185
R15578 vdd.n485 vdd.n484 185
R15579 vdd.n483 vdd.n460 185
R15580 vdd.n479 vdd.n478 185
R15581 vdd.n477 vdd.n476 185
R15582 vdd.n475 vdd.n474 185
R15583 vdd.n473 vdd.n462 185
R15584 vdd.n469 vdd.n468 185
R15585 vdd.n467 vdd.n466 185
R15586 vdd.n465 vdd.n392 185
R15587 vdd.n3348 vdd.n393 185
R15588 vdd.n3355 vdd.n393 185
R15589 vdd.n3347 vdd.n3346 185
R15590 vdd.n3346 vdd.n386 185
R15591 vdd.n3345 vdd.n385 185
R15592 vdd.n3361 vdd.n385 185
R15593 vdd.n621 vdd.n384 185
R15594 vdd.n3362 vdd.n384 185
R15595 vdd.n3341 vdd.n383 185
R15596 vdd.n3363 vdd.n383 185
R15597 vdd.n3340 vdd.n3339 185
R15598 vdd.n3339 vdd.n375 185
R15599 vdd.n3338 vdd.n374 185
R15600 vdd.n3369 vdd.n374 185
R15601 vdd.n623 vdd.n373 185
R15602 vdd.n3370 vdd.n373 185
R15603 vdd.n3334 vdd.n372 185
R15604 vdd.n3371 vdd.n372 185
R15605 vdd.n3333 vdd.n3332 185
R15606 vdd.n3332 vdd.n3331 185
R15607 vdd.n3330 vdd.n364 185
R15608 vdd.n3377 vdd.n364 185
R15609 vdd.n625 vdd.n363 185
R15610 vdd.n3378 vdd.n363 185
R15611 vdd.n3326 vdd.n362 185
R15612 vdd.n3379 vdd.n362 185
R15613 vdd.n3325 vdd.n3324 185
R15614 vdd.n3324 vdd.n361 185
R15615 vdd.n3323 vdd.n353 185
R15616 vdd.n3385 vdd.n353 185
R15617 vdd.n627 vdd.n352 185
R15618 vdd.n3386 vdd.n352 185
R15619 vdd.n3319 vdd.n351 185
R15620 vdd.n3387 vdd.n351 185
R15621 vdd.n3318 vdd.n3317 185
R15622 vdd.n3317 vdd.n344 185
R15623 vdd.n3316 vdd.n343 185
R15624 vdd.n3393 vdd.n343 185
R15625 vdd.n629 vdd.n342 185
R15626 vdd.n3394 vdd.n342 185
R15627 vdd.n3312 vdd.n341 185
R15628 vdd.n3395 vdd.n341 185
R15629 vdd.n3311 vdd.n3310 185
R15630 vdd.n3310 vdd.n340 185
R15631 vdd.n3309 vdd.n631 185
R15632 vdd.n3309 vdd.n3308 185
R15633 vdd.n3297 vdd.n632 185
R15634 vdd.n633 vdd.n632 185
R15635 vdd.n3299 vdd.n3298 185
R15636 vdd.n3300 vdd.n3299 185
R15637 vdd.n640 vdd.n639 185
R15638 vdd.n644 vdd.n639 185
R15639 vdd.n3291 vdd.n3290 185
R15640 vdd.n3290 vdd.n3289 185
R15641 vdd.n643 vdd.n642 185
R15642 vdd.n3280 vdd.n643 185
R15643 vdd.n3279 vdd.n3278 185
R15644 vdd.n3281 vdd.n3279 185
R15645 vdd.n651 vdd.n650 185
R15646 vdd.n656 vdd.n650 185
R15647 vdd.n3274 vdd.n3273 185
R15648 vdd.n3273 vdd.n3272 185
R15649 vdd.n654 vdd.n653 185
R15650 vdd.n655 vdd.n654 185
R15651 vdd.n3263 vdd.n3262 185
R15652 vdd.n3264 vdd.n3263 185
R15653 vdd.n664 vdd.n663 185
R15654 vdd.n663 vdd.n662 185
R15655 vdd.n3258 vdd.n3257 185
R15656 vdd.n3257 vdd.n3256 185
R15657 vdd.n667 vdd.n666 185
R15658 vdd.n3247 vdd.n667 185
R15659 vdd.n3246 vdd.n3245 185
R15660 vdd.n3248 vdd.n3246 185
R15661 vdd.n674 vdd.n673 185
R15662 vdd.n679 vdd.n673 185
R15663 vdd.n3241 vdd.n3240 185
R15664 vdd.n3240 vdd.n3239 185
R15665 vdd.n677 vdd.n676 185
R15666 vdd.n678 vdd.n677 185
R15667 vdd.n3230 vdd.n3229 185
R15668 vdd.n3231 vdd.n3230 185
R15669 vdd.n686 vdd.n685 185
R15670 vdd.n723 vdd.n685 185
R15671 vdd.n913 vdd.n912 185
R15672 vdd.n2855 vdd.n2854 185
R15673 vdd.n2853 vdd.n2638 185
R15674 vdd.n2857 vdd.n2638 185
R15675 vdd.n2852 vdd.n2851 185
R15676 vdd.n2850 vdd.n2849 185
R15677 vdd.n2848 vdd.n2847 185
R15678 vdd.n2846 vdd.n2845 185
R15679 vdd.n2844 vdd.n2843 185
R15680 vdd.n2842 vdd.n2841 185
R15681 vdd.n2840 vdd.n2839 185
R15682 vdd.n2838 vdd.n2837 185
R15683 vdd.n2836 vdd.n2835 185
R15684 vdd.n2834 vdd.n2833 185
R15685 vdd.n2832 vdd.n2831 185
R15686 vdd.n2830 vdd.n2829 185
R15687 vdd.n2828 vdd.n2827 185
R15688 vdd.n2826 vdd.n2825 185
R15689 vdd.n2824 vdd.n2823 185
R15690 vdd.n2822 vdd.n2821 185
R15691 vdd.n2820 vdd.n2819 185
R15692 vdd.n2818 vdd.n2817 185
R15693 vdd.n2816 vdd.n2815 185
R15694 vdd.n2814 vdd.n2813 185
R15695 vdd.n2812 vdd.n2811 185
R15696 vdd.n2810 vdd.n2809 185
R15697 vdd.n2808 vdd.n2807 185
R15698 vdd.n2806 vdd.n2805 185
R15699 vdd.n2804 vdd.n2803 185
R15700 vdd.n2802 vdd.n2801 185
R15701 vdd.n2800 vdd.n2799 185
R15702 vdd.n2798 vdd.n2797 185
R15703 vdd.n2796 vdd.n2795 185
R15704 vdd.n2793 vdd.n2792 185
R15705 vdd.n2791 vdd.n2790 185
R15706 vdd.n2789 vdd.n2788 185
R15707 vdd.n2995 vdd.n2994 185
R15708 vdd.n2997 vdd.n834 185
R15709 vdd.n2999 vdd.n2998 185
R15710 vdd.n3001 vdd.n831 185
R15711 vdd.n3003 vdd.n3002 185
R15712 vdd.n3005 vdd.n829 185
R15713 vdd.n3007 vdd.n3006 185
R15714 vdd.n3008 vdd.n828 185
R15715 vdd.n3010 vdd.n3009 185
R15716 vdd.n3012 vdd.n826 185
R15717 vdd.n3014 vdd.n3013 185
R15718 vdd.n3015 vdd.n825 185
R15719 vdd.n3017 vdd.n3016 185
R15720 vdd.n3019 vdd.n823 185
R15721 vdd.n3021 vdd.n3020 185
R15722 vdd.n3022 vdd.n822 185
R15723 vdd.n3024 vdd.n3023 185
R15724 vdd.n3026 vdd.n731 185
R15725 vdd.n3028 vdd.n3027 185
R15726 vdd.n3030 vdd.n820 185
R15727 vdd.n3032 vdd.n3031 185
R15728 vdd.n3033 vdd.n819 185
R15729 vdd.n3035 vdd.n3034 185
R15730 vdd.n3037 vdd.n817 185
R15731 vdd.n3039 vdd.n3038 185
R15732 vdd.n3040 vdd.n816 185
R15733 vdd.n3042 vdd.n3041 185
R15734 vdd.n3044 vdd.n814 185
R15735 vdd.n3046 vdd.n3045 185
R15736 vdd.n3047 vdd.n813 185
R15737 vdd.n3049 vdd.n3048 185
R15738 vdd.n3051 vdd.n812 185
R15739 vdd.n3052 vdd.n811 185
R15740 vdd.n3055 vdd.n3054 185
R15741 vdd.n3056 vdd.n809 185
R15742 vdd.n809 vdd.n692 185
R15743 vdd.n2993 vdd.n806 185
R15744 vdd.n3059 vdd.n806 185
R15745 vdd.n2992 vdd.n2991 185
R15746 vdd.n2991 vdd.n805 185
R15747 vdd.n2990 vdd.n836 185
R15748 vdd.n2990 vdd.n2989 185
R15749 vdd.n2744 vdd.n837 185
R15750 vdd.n846 vdd.n837 185
R15751 vdd.n2745 vdd.n844 185
R15752 vdd.n2983 vdd.n844 185
R15753 vdd.n2747 vdd.n2746 185
R15754 vdd.n2746 vdd.n843 185
R15755 vdd.n2748 vdd.n852 185
R15756 vdd.n2932 vdd.n852 185
R15757 vdd.n2750 vdd.n2749 185
R15758 vdd.n2749 vdd.n851 185
R15759 vdd.n2751 vdd.n858 185
R15760 vdd.n2926 vdd.n858 185
R15761 vdd.n2753 vdd.n2752 185
R15762 vdd.n2752 vdd.n857 185
R15763 vdd.n2754 vdd.n863 185
R15764 vdd.n2918 vdd.n863 185
R15765 vdd.n2756 vdd.n2755 185
R15766 vdd.n2755 vdd.n870 185
R15767 vdd.n2757 vdd.n868 185
R15768 vdd.n2912 vdd.n868 185
R15769 vdd.n2759 vdd.n2758 185
R15770 vdd.n2760 vdd.n2759 185
R15771 vdd.n2743 vdd.n875 185
R15772 vdd.n2906 vdd.n875 185
R15773 vdd.n2742 vdd.n2741 185
R15774 vdd.n2741 vdd.n874 185
R15775 vdd.n2740 vdd.n881 185
R15776 vdd.n2900 vdd.n881 185
R15777 vdd.n2739 vdd.n2738 185
R15778 vdd.n2738 vdd.n880 185
R15779 vdd.n2737 vdd.n886 185
R15780 vdd.n2894 vdd.n886 185
R15781 vdd.n2736 vdd.n2735 185
R15782 vdd.n2735 vdd.n893 185
R15783 vdd.n2734 vdd.n891 185
R15784 vdd.n2888 vdd.n891 185
R15785 vdd.n2733 vdd.n2732 185
R15786 vdd.n2732 vdd.n900 185
R15787 vdd.n2731 vdd.n898 185
R15788 vdd.n2882 vdd.n898 185
R15789 vdd.n2730 vdd.n2729 185
R15790 vdd.n2729 vdd.n897 185
R15791 vdd.n2641 vdd.n904 185
R15792 vdd.n2876 vdd.n904 185
R15793 vdd.n2783 vdd.n2782 185
R15794 vdd.n2782 vdd.n2781 185
R15795 vdd.n2784 vdd.n909 185
R15796 vdd.n2870 vdd.n909 185
R15797 vdd.n2786 vdd.n2785 185
R15798 vdd.n2785 vdd.t200 185
R15799 vdd.n2787 vdd.n914 185
R15800 vdd.n2864 vdd.n914 185
R15801 vdd.n2866 vdd.n2865 185
R15802 vdd.n2865 vdd.n2864 185
R15803 vdd.n2867 vdd.n911 185
R15804 vdd.n911 vdd.t200 185
R15805 vdd.n2869 vdd.n2868 185
R15806 vdd.n2870 vdd.n2869 185
R15807 vdd.n903 vdd.n902 185
R15808 vdd.n2781 vdd.n903 185
R15809 vdd.n2878 vdd.n2877 185
R15810 vdd.n2877 vdd.n2876 185
R15811 vdd.n2879 vdd.n901 185
R15812 vdd.n901 vdd.n897 185
R15813 vdd.n2881 vdd.n2880 185
R15814 vdd.n2882 vdd.n2881 185
R15815 vdd.n890 vdd.n889 185
R15816 vdd.n900 vdd.n890 185
R15817 vdd.n2890 vdd.n2889 185
R15818 vdd.n2889 vdd.n2888 185
R15819 vdd.n2891 vdd.n888 185
R15820 vdd.n893 vdd.n888 185
R15821 vdd.n2893 vdd.n2892 185
R15822 vdd.n2894 vdd.n2893 185
R15823 vdd.n879 vdd.n878 185
R15824 vdd.n880 vdd.n879 185
R15825 vdd.n2902 vdd.n2901 185
R15826 vdd.n2901 vdd.n2900 185
R15827 vdd.n2903 vdd.n877 185
R15828 vdd.n877 vdd.n874 185
R15829 vdd.n2905 vdd.n2904 185
R15830 vdd.n2906 vdd.n2905 185
R15831 vdd.n867 vdd.n866 185
R15832 vdd.n2760 vdd.n867 185
R15833 vdd.n2914 vdd.n2913 185
R15834 vdd.n2913 vdd.n2912 185
R15835 vdd.n2915 vdd.n865 185
R15836 vdd.n870 vdd.n865 185
R15837 vdd.n2917 vdd.n2916 185
R15838 vdd.n2918 vdd.n2917 185
R15839 vdd.n856 vdd.n855 185
R15840 vdd.n857 vdd.n856 185
R15841 vdd.n2928 vdd.n2927 185
R15842 vdd.n2927 vdd.n2926 185
R15843 vdd.n2929 vdd.n854 185
R15844 vdd.n854 vdd.n851 185
R15845 vdd.n2931 vdd.n2930 185
R15846 vdd.n2932 vdd.n2931 185
R15847 vdd.n842 vdd.n841 185
R15848 vdd.n843 vdd.n842 185
R15849 vdd.n2985 vdd.n2984 185
R15850 vdd.n2984 vdd.n2983 185
R15851 vdd.n2986 vdd.n840 185
R15852 vdd.n846 vdd.n840 185
R15853 vdd.n2988 vdd.n2987 185
R15854 vdd.n2989 vdd.n2988 185
R15855 vdd.n810 vdd.n808 185
R15856 vdd.n808 vdd.n805 185
R15857 vdd.n3058 vdd.n3057 185
R15858 vdd.n3059 vdd.n3058 185
R15859 vdd.n2531 vdd.n2530 185
R15860 vdd.n2532 vdd.n2531 185
R15861 vdd.n964 vdd.n962 185
R15862 vdd.n962 vdd.t292 185
R15863 vdd.n2446 vdd.n971 185
R15864 vdd.n2457 vdd.n971 185
R15865 vdd.n2447 vdd.n980 185
R15866 vdd.n2156 vdd.n980 185
R15867 vdd.n2449 vdd.n2448 185
R15868 vdd.n2450 vdd.n2449 185
R15869 vdd.n2445 vdd.n979 185
R15870 vdd.n979 vdd.n976 185
R15871 vdd.n2444 vdd.n2443 185
R15872 vdd.n2443 vdd.n2442 185
R15873 vdd.n982 vdd.n981 185
R15874 vdd.n983 vdd.n982 185
R15875 vdd.n2435 vdd.n2434 185
R15876 vdd.n2436 vdd.n2435 185
R15877 vdd.n2433 vdd.n992 185
R15878 vdd.n992 vdd.n989 185
R15879 vdd.n2432 vdd.n2431 185
R15880 vdd.n2431 vdd.n2430 185
R15881 vdd.n994 vdd.n993 185
R15882 vdd.n1002 vdd.n994 185
R15883 vdd.n2423 vdd.n2422 185
R15884 vdd.n2424 vdd.n2423 185
R15885 vdd.n2421 vdd.n1003 185
R15886 vdd.n1008 vdd.n1003 185
R15887 vdd.n2420 vdd.n2419 185
R15888 vdd.n2419 vdd.n2418 185
R15889 vdd.n1005 vdd.n1004 185
R15890 vdd.n2257 vdd.n1005 185
R15891 vdd.n2411 vdd.n2410 185
R15892 vdd.n2412 vdd.n2411 185
R15893 vdd.n2409 vdd.n1015 185
R15894 vdd.n1015 vdd.n1012 185
R15895 vdd.n2408 vdd.n2407 185
R15896 vdd.n2407 vdd.n2406 185
R15897 vdd.n1017 vdd.n1016 185
R15898 vdd.n1018 vdd.n1017 185
R15899 vdd.n2399 vdd.n2398 185
R15900 vdd.n2400 vdd.n2399 185
R15901 vdd.n2396 vdd.n1026 185
R15902 vdd.n1033 vdd.n1026 185
R15903 vdd.n2395 vdd.n2394 185
R15904 vdd.n2394 vdd.n2393 185
R15905 vdd.n1029 vdd.n1028 185
R15906 vdd.n1030 vdd.n1029 185
R15907 vdd.n2386 vdd.n2385 185
R15908 vdd.n2387 vdd.n2386 185
R15909 vdd.n2384 vdd.n1040 185
R15910 vdd.n1040 vdd.n1037 185
R15911 vdd.n2383 vdd.n2382 185
R15912 vdd.n2382 vdd.n2381 185
R15913 vdd.n1042 vdd.n1041 185
R15914 vdd.n1043 vdd.n1042 185
R15915 vdd.n2374 vdd.n2373 185
R15916 vdd.n2375 vdd.n2374 185
R15917 vdd.n2462 vdd.n936 185
R15918 vdd.n2604 vdd.n936 185
R15919 vdd.n2464 vdd.n2463 185
R15920 vdd.n2466 vdd.n2465 185
R15921 vdd.n2468 vdd.n2467 185
R15922 vdd.n2470 vdd.n2469 185
R15923 vdd.n2472 vdd.n2471 185
R15924 vdd.n2474 vdd.n2473 185
R15925 vdd.n2476 vdd.n2475 185
R15926 vdd.n2478 vdd.n2477 185
R15927 vdd.n2480 vdd.n2479 185
R15928 vdd.n2482 vdd.n2481 185
R15929 vdd.n2484 vdd.n2483 185
R15930 vdd.n2486 vdd.n2485 185
R15931 vdd.n2488 vdd.n2487 185
R15932 vdd.n2490 vdd.n2489 185
R15933 vdd.n2492 vdd.n2491 185
R15934 vdd.n2494 vdd.n2493 185
R15935 vdd.n2496 vdd.n2495 185
R15936 vdd.n2498 vdd.n2497 185
R15937 vdd.n2500 vdd.n2499 185
R15938 vdd.n2502 vdd.n2501 185
R15939 vdd.n2504 vdd.n2503 185
R15940 vdd.n2506 vdd.n2505 185
R15941 vdd.n2508 vdd.n2507 185
R15942 vdd.n2510 vdd.n2509 185
R15943 vdd.n2512 vdd.n2511 185
R15944 vdd.n2514 vdd.n2513 185
R15945 vdd.n2516 vdd.n2515 185
R15946 vdd.n2518 vdd.n2517 185
R15947 vdd.n2520 vdd.n2519 185
R15948 vdd.n2522 vdd.n2521 185
R15949 vdd.n2524 vdd.n2523 185
R15950 vdd.n2526 vdd.n2525 185
R15951 vdd.n2528 vdd.n2527 185
R15952 vdd.n2529 vdd.n963 185
R15953 vdd.n2461 vdd.n961 185
R15954 vdd.n2532 vdd.n961 185
R15955 vdd.n2460 vdd.n2459 185
R15956 vdd.n2459 vdd.t292 185
R15957 vdd.n2458 vdd.n968 185
R15958 vdd.n2458 vdd.n2457 185
R15959 vdd.n2238 vdd.n969 185
R15960 vdd.n2156 vdd.n969 185
R15961 vdd.n2239 vdd.n978 185
R15962 vdd.n2450 vdd.n978 185
R15963 vdd.n2241 vdd.n2240 185
R15964 vdd.n2240 vdd.n976 185
R15965 vdd.n2242 vdd.n985 185
R15966 vdd.n2442 vdd.n985 185
R15967 vdd.n2244 vdd.n2243 185
R15968 vdd.n2243 vdd.n983 185
R15969 vdd.n2245 vdd.n991 185
R15970 vdd.n2436 vdd.n991 185
R15971 vdd.n2247 vdd.n2246 185
R15972 vdd.n2246 vdd.n989 185
R15973 vdd.n2248 vdd.n996 185
R15974 vdd.n2430 vdd.n996 185
R15975 vdd.n2250 vdd.n2249 185
R15976 vdd.n2249 vdd.n1002 185
R15977 vdd.n2251 vdd.n1001 185
R15978 vdd.n2424 vdd.n1001 185
R15979 vdd.n2253 vdd.n2252 185
R15980 vdd.n2252 vdd.n1008 185
R15981 vdd.n2254 vdd.n1007 185
R15982 vdd.n2418 vdd.n1007 185
R15983 vdd.n2256 vdd.n2255 185
R15984 vdd.n2257 vdd.n2256 185
R15985 vdd.n2237 vdd.n1014 185
R15986 vdd.n2412 vdd.n1014 185
R15987 vdd.n2236 vdd.n2235 185
R15988 vdd.n2235 vdd.n1012 185
R15989 vdd.n2234 vdd.n1020 185
R15990 vdd.n2406 vdd.n1020 185
R15991 vdd.n2233 vdd.n2232 185
R15992 vdd.n2232 vdd.n1018 185
R15993 vdd.n2231 vdd.n1025 185
R15994 vdd.n2400 vdd.n1025 185
R15995 vdd.n2230 vdd.n2229 185
R15996 vdd.n2229 vdd.n1033 185
R15997 vdd.n2228 vdd.n1032 185
R15998 vdd.n2393 vdd.n1032 185
R15999 vdd.n2227 vdd.n2226 185
R16000 vdd.n2226 vdd.n1030 185
R16001 vdd.n2225 vdd.n1039 185
R16002 vdd.n2387 vdd.n1039 185
R16003 vdd.n2224 vdd.n2223 185
R16004 vdd.n2223 vdd.n1037 185
R16005 vdd.n2222 vdd.n1045 185
R16006 vdd.n2381 vdd.n1045 185
R16007 vdd.n2221 vdd.n2220 185
R16008 vdd.n2220 vdd.n1043 185
R16009 vdd.n2219 vdd.n1051 185
R16010 vdd.n2375 vdd.n1051 185
R16011 vdd.n2372 vdd.n1052 185
R16012 vdd.n2371 vdd.n2370 185
R16013 vdd.n2368 vdd.n1053 185
R16014 vdd.n2366 vdd.n2365 185
R16015 vdd.n2364 vdd.n1054 185
R16016 vdd.n2363 vdd.n2362 185
R16017 vdd.n2360 vdd.n1055 185
R16018 vdd.n2358 vdd.n2357 185
R16019 vdd.n2356 vdd.n1056 185
R16020 vdd.n2355 vdd.n2354 185
R16021 vdd.n2352 vdd.n1057 185
R16022 vdd.n2350 vdd.n2349 185
R16023 vdd.n2348 vdd.n1058 185
R16024 vdd.n2347 vdd.n2346 185
R16025 vdd.n2344 vdd.n1059 185
R16026 vdd.n2342 vdd.n2341 185
R16027 vdd.n2340 vdd.n1060 185
R16028 vdd.n2339 vdd.n1062 185
R16029 vdd.n2184 vdd.n1063 185
R16030 vdd.n2187 vdd.n2186 185
R16031 vdd.n2189 vdd.n2188 185
R16032 vdd.n2191 vdd.n2183 185
R16033 vdd.n2194 vdd.n2193 185
R16034 vdd.n2195 vdd.n2182 185
R16035 vdd.n2197 vdd.n2196 185
R16036 vdd.n2199 vdd.n2181 185
R16037 vdd.n2202 vdd.n2201 185
R16038 vdd.n2203 vdd.n2180 185
R16039 vdd.n2205 vdd.n2204 185
R16040 vdd.n2207 vdd.n2179 185
R16041 vdd.n2210 vdd.n2209 185
R16042 vdd.n2211 vdd.n2176 185
R16043 vdd.n2214 vdd.n2213 185
R16044 vdd.n2216 vdd.n2175 185
R16045 vdd.n2218 vdd.n2217 185
R16046 vdd.n2217 vdd.n1049 185
R16047 vdd.n327 vdd.n326 171.744
R16048 vdd.n326 vdd.n325 171.744
R16049 vdd.n325 vdd.n294 171.744
R16050 vdd.n318 vdd.n294 171.744
R16051 vdd.n318 vdd.n317 171.744
R16052 vdd.n317 vdd.n299 171.744
R16053 vdd.n310 vdd.n299 171.744
R16054 vdd.n310 vdd.n309 171.744
R16055 vdd.n309 vdd.n303 171.744
R16056 vdd.n268 vdd.n267 171.744
R16057 vdd.n267 vdd.n266 171.744
R16058 vdd.n266 vdd.n235 171.744
R16059 vdd.n259 vdd.n235 171.744
R16060 vdd.n259 vdd.n258 171.744
R16061 vdd.n258 vdd.n240 171.744
R16062 vdd.n251 vdd.n240 171.744
R16063 vdd.n251 vdd.n250 171.744
R16064 vdd.n250 vdd.n244 171.744
R16065 vdd.n225 vdd.n224 171.744
R16066 vdd.n224 vdd.n223 171.744
R16067 vdd.n223 vdd.n192 171.744
R16068 vdd.n216 vdd.n192 171.744
R16069 vdd.n216 vdd.n215 171.744
R16070 vdd.n215 vdd.n197 171.744
R16071 vdd.n208 vdd.n197 171.744
R16072 vdd.n208 vdd.n207 171.744
R16073 vdd.n207 vdd.n201 171.744
R16074 vdd.n166 vdd.n165 171.744
R16075 vdd.n165 vdd.n164 171.744
R16076 vdd.n164 vdd.n133 171.744
R16077 vdd.n157 vdd.n133 171.744
R16078 vdd.n157 vdd.n156 171.744
R16079 vdd.n156 vdd.n138 171.744
R16080 vdd.n149 vdd.n138 171.744
R16081 vdd.n149 vdd.n148 171.744
R16082 vdd.n148 vdd.n142 171.744
R16083 vdd.n124 vdd.n123 171.744
R16084 vdd.n123 vdd.n122 171.744
R16085 vdd.n122 vdd.n91 171.744
R16086 vdd.n115 vdd.n91 171.744
R16087 vdd.n115 vdd.n114 171.744
R16088 vdd.n114 vdd.n96 171.744
R16089 vdd.n107 vdd.n96 171.744
R16090 vdd.n107 vdd.n106 171.744
R16091 vdd.n106 vdd.n100 171.744
R16092 vdd.n65 vdd.n64 171.744
R16093 vdd.n64 vdd.n63 171.744
R16094 vdd.n63 vdd.n32 171.744
R16095 vdd.n56 vdd.n32 171.744
R16096 vdd.n56 vdd.n55 171.744
R16097 vdd.n55 vdd.n37 171.744
R16098 vdd.n48 vdd.n37 171.744
R16099 vdd.n48 vdd.n47 171.744
R16100 vdd.n47 vdd.n41 171.744
R16101 vdd.n1746 vdd.n1745 171.744
R16102 vdd.n1745 vdd.n1744 171.744
R16103 vdd.n1744 vdd.n1713 171.744
R16104 vdd.n1737 vdd.n1713 171.744
R16105 vdd.n1737 vdd.n1736 171.744
R16106 vdd.n1736 vdd.n1718 171.744
R16107 vdd.n1729 vdd.n1718 171.744
R16108 vdd.n1729 vdd.n1728 171.744
R16109 vdd.n1728 vdd.n1722 171.744
R16110 vdd.n1805 vdd.n1804 171.744
R16111 vdd.n1804 vdd.n1803 171.744
R16112 vdd.n1803 vdd.n1772 171.744
R16113 vdd.n1796 vdd.n1772 171.744
R16114 vdd.n1796 vdd.n1795 171.744
R16115 vdd.n1795 vdd.n1777 171.744
R16116 vdd.n1788 vdd.n1777 171.744
R16117 vdd.n1788 vdd.n1787 171.744
R16118 vdd.n1787 vdd.n1781 171.744
R16119 vdd.n1644 vdd.n1643 171.744
R16120 vdd.n1643 vdd.n1642 171.744
R16121 vdd.n1642 vdd.n1611 171.744
R16122 vdd.n1635 vdd.n1611 171.744
R16123 vdd.n1635 vdd.n1634 171.744
R16124 vdd.n1634 vdd.n1616 171.744
R16125 vdd.n1627 vdd.n1616 171.744
R16126 vdd.n1627 vdd.n1626 171.744
R16127 vdd.n1626 vdd.n1620 171.744
R16128 vdd.n1703 vdd.n1702 171.744
R16129 vdd.n1702 vdd.n1701 171.744
R16130 vdd.n1701 vdd.n1670 171.744
R16131 vdd.n1694 vdd.n1670 171.744
R16132 vdd.n1694 vdd.n1693 171.744
R16133 vdd.n1693 vdd.n1675 171.744
R16134 vdd.n1686 vdd.n1675 171.744
R16135 vdd.n1686 vdd.n1685 171.744
R16136 vdd.n1685 vdd.n1679 171.744
R16137 vdd.n1543 vdd.n1542 171.744
R16138 vdd.n1542 vdd.n1541 171.744
R16139 vdd.n1541 vdd.n1510 171.744
R16140 vdd.n1534 vdd.n1510 171.744
R16141 vdd.n1534 vdd.n1533 171.744
R16142 vdd.n1533 vdd.n1515 171.744
R16143 vdd.n1526 vdd.n1515 171.744
R16144 vdd.n1526 vdd.n1525 171.744
R16145 vdd.n1525 vdd.n1519 171.744
R16146 vdd.n1602 vdd.n1601 171.744
R16147 vdd.n1601 vdd.n1600 171.744
R16148 vdd.n1600 vdd.n1569 171.744
R16149 vdd.n1593 vdd.n1569 171.744
R16150 vdd.n1593 vdd.n1592 171.744
R16151 vdd.n1592 vdd.n1574 171.744
R16152 vdd.n1585 vdd.n1574 171.744
R16153 vdd.n1585 vdd.n1584 171.744
R16154 vdd.n1584 vdd.n1578 171.744
R16155 vdd.n468 vdd.n467 146.341
R16156 vdd.n474 vdd.n473 146.341
R16157 vdd.n478 vdd.n477 146.341
R16158 vdd.n484 vdd.n483 146.341
R16159 vdd.n488 vdd.n487 146.341
R16160 vdd.n494 vdd.n493 146.341
R16161 vdd.n498 vdd.n497 146.341
R16162 vdd.n504 vdd.n503 146.341
R16163 vdd.n508 vdd.n507 146.341
R16164 vdd.n514 vdd.n513 146.341
R16165 vdd.n518 vdd.n517 146.341
R16166 vdd.n524 vdd.n523 146.341
R16167 vdd.n528 vdd.n527 146.341
R16168 vdd.n534 vdd.n533 146.341
R16169 vdd.n538 vdd.n537 146.341
R16170 vdd.n544 vdd.n543 146.341
R16171 vdd.n548 vdd.n547 146.341
R16172 vdd.n554 vdd.n553 146.341
R16173 vdd.n558 vdd.n557 146.341
R16174 vdd.n564 vdd.n563 146.341
R16175 vdd.n568 vdd.n567 146.341
R16176 vdd.n574 vdd.n573 146.341
R16177 vdd.n578 vdd.n577 146.341
R16178 vdd.n584 vdd.n583 146.341
R16179 vdd.n588 vdd.n587 146.341
R16180 vdd.n594 vdd.n593 146.341
R16181 vdd.n598 vdd.n597 146.341
R16182 vdd.n604 vdd.n603 146.341
R16183 vdd.n608 vdd.n607 146.341
R16184 vdd.n614 vdd.n613 146.341
R16185 vdd.n616 vdd.n425 146.341
R16186 vdd.n3230 vdd.n685 146.341
R16187 vdd.n3230 vdd.n677 146.341
R16188 vdd.n3240 vdd.n677 146.341
R16189 vdd.n3240 vdd.n673 146.341
R16190 vdd.n3246 vdd.n673 146.341
R16191 vdd.n3246 vdd.n667 146.341
R16192 vdd.n3257 vdd.n667 146.341
R16193 vdd.n3257 vdd.n663 146.341
R16194 vdd.n3263 vdd.n663 146.341
R16195 vdd.n3263 vdd.n654 146.341
R16196 vdd.n3273 vdd.n654 146.341
R16197 vdd.n3273 vdd.n650 146.341
R16198 vdd.n3279 vdd.n650 146.341
R16199 vdd.n3279 vdd.n643 146.341
R16200 vdd.n3290 vdd.n643 146.341
R16201 vdd.n3290 vdd.n639 146.341
R16202 vdd.n3299 vdd.n639 146.341
R16203 vdd.n3299 vdd.n632 146.341
R16204 vdd.n3309 vdd.n632 146.341
R16205 vdd.n3310 vdd.n3309 146.341
R16206 vdd.n3310 vdd.n341 146.341
R16207 vdd.n342 vdd.n341 146.341
R16208 vdd.n343 vdd.n342 146.341
R16209 vdd.n3317 vdd.n343 146.341
R16210 vdd.n3317 vdd.n351 146.341
R16211 vdd.n352 vdd.n351 146.341
R16212 vdd.n353 vdd.n352 146.341
R16213 vdd.n3324 vdd.n353 146.341
R16214 vdd.n3324 vdd.n362 146.341
R16215 vdd.n363 vdd.n362 146.341
R16216 vdd.n364 vdd.n363 146.341
R16217 vdd.n3332 vdd.n364 146.341
R16218 vdd.n3332 vdd.n372 146.341
R16219 vdd.n373 vdd.n372 146.341
R16220 vdd.n374 vdd.n373 146.341
R16221 vdd.n3339 vdd.n374 146.341
R16222 vdd.n3339 vdd.n383 146.341
R16223 vdd.n384 vdd.n383 146.341
R16224 vdd.n385 vdd.n384 146.341
R16225 vdd.n3346 vdd.n385 146.341
R16226 vdd.n3346 vdd.n393 146.341
R16227 vdd.n725 vdd.n724 146.341
R16228 vdd.n728 vdd.n724 146.341
R16229 vdd.n734 vdd.n733 146.341
R16230 vdd.n3212 vdd.n3211 146.341
R16231 vdd.n3208 vdd.n3207 146.341
R16232 vdd.n3204 vdd.n3203 146.341
R16233 vdd.n3200 vdd.n3199 146.341
R16234 vdd.n3196 vdd.n3195 146.341
R16235 vdd.n3192 vdd.n3191 146.341
R16236 vdd.n3188 vdd.n3187 146.341
R16237 vdd.n3179 vdd.n3178 146.341
R16238 vdd.n3176 vdd.n3175 146.341
R16239 vdd.n3172 vdd.n3171 146.341
R16240 vdd.n3168 vdd.n3167 146.341
R16241 vdd.n3164 vdd.n3163 146.341
R16242 vdd.n3160 vdd.n3159 146.341
R16243 vdd.n3156 vdd.n3155 146.341
R16244 vdd.n3152 vdd.n3151 146.341
R16245 vdd.n3148 vdd.n3147 146.341
R16246 vdd.n3144 vdd.n3143 146.341
R16247 vdd.n3140 vdd.n3139 146.341
R16248 vdd.n3133 vdd.n3132 146.341
R16249 vdd.n3130 vdd.n3129 146.341
R16250 vdd.n3126 vdd.n3125 146.341
R16251 vdd.n3122 vdd.n3121 146.341
R16252 vdd.n3118 vdd.n3117 146.341
R16253 vdd.n3114 vdd.n3113 146.341
R16254 vdd.n3110 vdd.n3109 146.341
R16255 vdd.n3106 vdd.n3105 146.341
R16256 vdd.n3102 vdd.n3101 146.341
R16257 vdd.n3098 vdd.n3097 146.341
R16258 vdd.n3224 vdd.n691 146.341
R16259 vdd.n3232 vdd.n684 146.341
R16260 vdd.n3232 vdd.n680 146.341
R16261 vdd.n3238 vdd.n680 146.341
R16262 vdd.n3238 vdd.n672 146.341
R16263 vdd.n3249 vdd.n672 146.341
R16264 vdd.n3249 vdd.n668 146.341
R16265 vdd.n3255 vdd.n668 146.341
R16266 vdd.n3255 vdd.n661 146.341
R16267 vdd.n3265 vdd.n661 146.341
R16268 vdd.n3265 vdd.n657 146.341
R16269 vdd.n3271 vdd.n657 146.341
R16270 vdd.n3271 vdd.n649 146.341
R16271 vdd.n3282 vdd.n649 146.341
R16272 vdd.n3282 vdd.n645 146.341
R16273 vdd.n3288 vdd.n645 146.341
R16274 vdd.n3288 vdd.n638 146.341
R16275 vdd.n3301 vdd.n638 146.341
R16276 vdd.n3301 vdd.n634 146.341
R16277 vdd.n3307 vdd.n634 146.341
R16278 vdd.n3307 vdd.n338 146.341
R16279 vdd.n3396 vdd.n338 146.341
R16280 vdd.n3396 vdd.n339 146.341
R16281 vdd.n3392 vdd.n339 146.341
R16282 vdd.n3392 vdd.n345 146.341
R16283 vdd.n3388 vdd.n345 146.341
R16284 vdd.n3388 vdd.n350 146.341
R16285 vdd.n3384 vdd.n350 146.341
R16286 vdd.n3384 vdd.n354 146.341
R16287 vdd.n3380 vdd.n354 146.341
R16288 vdd.n3380 vdd.n360 146.341
R16289 vdd.n3376 vdd.n360 146.341
R16290 vdd.n3376 vdd.n365 146.341
R16291 vdd.n3372 vdd.n365 146.341
R16292 vdd.n3372 vdd.n371 146.341
R16293 vdd.n3368 vdd.n371 146.341
R16294 vdd.n3368 vdd.n376 146.341
R16295 vdd.n3364 vdd.n376 146.341
R16296 vdd.n3364 vdd.n382 146.341
R16297 vdd.n3360 vdd.n382 146.341
R16298 vdd.n3360 vdd.n387 146.341
R16299 vdd.n3356 vdd.n387 146.341
R16300 vdd.n2322 vdd.n2321 146.341
R16301 vdd.n2319 vdd.n1903 146.341
R16302 vdd.n2099 vdd.n1909 146.341
R16303 vdd.n2097 vdd.n2096 146.341
R16304 vdd.n2094 vdd.n1911 146.341
R16305 vdd.n2090 vdd.n2089 146.341
R16306 vdd.n2087 vdd.n1918 146.341
R16307 vdd.n2083 vdd.n2082 146.341
R16308 vdd.n2080 vdd.n1925 146.341
R16309 vdd.n1936 vdd.n1933 146.341
R16310 vdd.n2072 vdd.n2071 146.341
R16311 vdd.n2069 vdd.n1938 146.341
R16312 vdd.n2065 vdd.n2064 146.341
R16313 vdd.n2062 vdd.n1944 146.341
R16314 vdd.n2058 vdd.n2057 146.341
R16315 vdd.n2055 vdd.n1951 146.341
R16316 vdd.n2051 vdd.n2050 146.341
R16317 vdd.n2048 vdd.n1958 146.341
R16318 vdd.n2044 vdd.n2043 146.341
R16319 vdd.n2041 vdd.n1965 146.341
R16320 vdd.n1976 vdd.n1973 146.341
R16321 vdd.n2033 vdd.n2032 146.341
R16322 vdd.n2030 vdd.n1978 146.341
R16323 vdd.n2026 vdd.n2025 146.341
R16324 vdd.n2023 vdd.n1984 146.341
R16325 vdd.n2019 vdd.n2018 146.341
R16326 vdd.n2016 vdd.n1991 146.341
R16327 vdd.n2012 vdd.n2011 146.341
R16328 vdd.n2009 vdd.n2006 146.341
R16329 vdd.n2004 vdd.n2001 146.341
R16330 vdd.n1999 vdd.n1069 146.341
R16331 vdd.n1428 vdd.n1188 146.341
R16332 vdd.n1428 vdd.n1184 146.341
R16333 vdd.n1434 vdd.n1184 146.341
R16334 vdd.n1434 vdd.n1176 146.341
R16335 vdd.n1445 vdd.n1176 146.341
R16336 vdd.n1445 vdd.n1172 146.341
R16337 vdd.n1451 vdd.n1172 146.341
R16338 vdd.n1451 vdd.n1166 146.341
R16339 vdd.n1462 vdd.n1166 146.341
R16340 vdd.n1462 vdd.n1162 146.341
R16341 vdd.n1468 vdd.n1162 146.341
R16342 vdd.n1468 vdd.n1153 146.341
R16343 vdd.n1478 vdd.n1153 146.341
R16344 vdd.n1478 vdd.n1149 146.341
R16345 vdd.n1484 vdd.n1149 146.341
R16346 vdd.n1484 vdd.n1142 146.341
R16347 vdd.n1495 vdd.n1142 146.341
R16348 vdd.n1495 vdd.n1138 146.341
R16349 vdd.n1501 vdd.n1138 146.341
R16350 vdd.n1501 vdd.n1131 146.341
R16351 vdd.n1818 vdd.n1131 146.341
R16352 vdd.n1818 vdd.n1127 146.341
R16353 vdd.n1824 vdd.n1127 146.341
R16354 vdd.n1824 vdd.n1119 146.341
R16355 vdd.n1835 vdd.n1119 146.341
R16356 vdd.n1835 vdd.n1115 146.341
R16357 vdd.n1841 vdd.n1115 146.341
R16358 vdd.n1841 vdd.n1109 146.341
R16359 vdd.n1852 vdd.n1109 146.341
R16360 vdd.n1852 vdd.n1105 146.341
R16361 vdd.n1858 vdd.n1105 146.341
R16362 vdd.n1858 vdd.n1096 146.341
R16363 vdd.n1868 vdd.n1096 146.341
R16364 vdd.n1868 vdd.n1092 146.341
R16365 vdd.n1874 vdd.n1092 146.341
R16366 vdd.n1874 vdd.n1086 146.341
R16367 vdd.n1885 vdd.n1086 146.341
R16368 vdd.n1885 vdd.n1081 146.341
R16369 vdd.n1893 vdd.n1081 146.341
R16370 vdd.n1893 vdd.n1071 146.341
R16371 vdd.n2330 vdd.n1071 146.341
R16372 vdd.n1417 vdd.n1193 146.341
R16373 vdd.n1417 vdd.n1226 146.341
R16374 vdd.n1230 vdd.n1229 146.341
R16375 vdd.n1232 vdd.n1231 146.341
R16376 vdd.n1236 vdd.n1235 146.341
R16377 vdd.n1238 vdd.n1237 146.341
R16378 vdd.n1242 vdd.n1241 146.341
R16379 vdd.n1244 vdd.n1243 146.341
R16380 vdd.n1248 vdd.n1247 146.341
R16381 vdd.n1250 vdd.n1249 146.341
R16382 vdd.n1256 vdd.n1255 146.341
R16383 vdd.n1258 vdd.n1257 146.341
R16384 vdd.n1262 vdd.n1261 146.341
R16385 vdd.n1264 vdd.n1263 146.341
R16386 vdd.n1268 vdd.n1267 146.341
R16387 vdd.n1270 vdd.n1269 146.341
R16388 vdd.n1274 vdd.n1273 146.341
R16389 vdd.n1276 vdd.n1275 146.341
R16390 vdd.n1280 vdd.n1279 146.341
R16391 vdd.n1282 vdd.n1281 146.341
R16392 vdd.n1354 vdd.n1285 146.341
R16393 vdd.n1287 vdd.n1286 146.341
R16394 vdd.n1291 vdd.n1290 146.341
R16395 vdd.n1293 vdd.n1292 146.341
R16396 vdd.n1297 vdd.n1296 146.341
R16397 vdd.n1299 vdd.n1298 146.341
R16398 vdd.n1303 vdd.n1302 146.341
R16399 vdd.n1305 vdd.n1304 146.341
R16400 vdd.n1309 vdd.n1308 146.341
R16401 vdd.n1311 vdd.n1310 146.341
R16402 vdd.n1315 vdd.n1314 146.341
R16403 vdd.n1316 vdd.n1224 146.341
R16404 vdd.n1426 vdd.n1189 146.341
R16405 vdd.n1426 vdd.n1182 146.341
R16406 vdd.n1437 vdd.n1182 146.341
R16407 vdd.n1437 vdd.n1178 146.341
R16408 vdd.n1443 vdd.n1178 146.341
R16409 vdd.n1443 vdd.n1171 146.341
R16410 vdd.n1454 vdd.n1171 146.341
R16411 vdd.n1454 vdd.n1167 146.341
R16412 vdd.n1460 vdd.n1167 146.341
R16413 vdd.n1460 vdd.n1160 146.341
R16414 vdd.n1470 vdd.n1160 146.341
R16415 vdd.n1470 vdd.n1156 146.341
R16416 vdd.n1476 vdd.n1156 146.341
R16417 vdd.n1476 vdd.n1148 146.341
R16418 vdd.n1487 vdd.n1148 146.341
R16419 vdd.n1487 vdd.n1144 146.341
R16420 vdd.n1493 vdd.n1144 146.341
R16421 vdd.n1493 vdd.n1137 146.341
R16422 vdd.n1503 vdd.n1137 146.341
R16423 vdd.n1503 vdd.n1133 146.341
R16424 vdd.n1816 vdd.n1133 146.341
R16425 vdd.n1816 vdd.n1125 146.341
R16426 vdd.n1827 vdd.n1125 146.341
R16427 vdd.n1827 vdd.n1121 146.341
R16428 vdd.n1833 vdd.n1121 146.341
R16429 vdd.n1833 vdd.n1114 146.341
R16430 vdd.n1844 vdd.n1114 146.341
R16431 vdd.n1844 vdd.n1110 146.341
R16432 vdd.n1850 vdd.n1110 146.341
R16433 vdd.n1850 vdd.n1103 146.341
R16434 vdd.n1860 vdd.n1103 146.341
R16435 vdd.n1860 vdd.n1099 146.341
R16436 vdd.n1866 vdd.n1099 146.341
R16437 vdd.n1866 vdd.n1091 146.341
R16438 vdd.n1877 vdd.n1091 146.341
R16439 vdd.n1877 vdd.n1087 146.341
R16440 vdd.n1883 vdd.n1087 146.341
R16441 vdd.n1883 vdd.n1079 146.341
R16442 vdd.n1896 vdd.n1079 146.341
R16443 vdd.n1896 vdd.n1074 146.341
R16444 vdd.n2328 vdd.n1074 146.341
R16445 vdd.n1073 vdd.n1049 141.707
R16446 vdd.n3223 vdd.n692 141.707
R16447 vdd.n2177 vdd.t267 127.284
R16448 vdd.n965 vdd.t252 127.284
R16449 vdd.n2151 vdd.t214 127.284
R16450 vdd.n957 vdd.t276 127.284
R16451 vdd.n2922 vdd.t228 127.284
R16452 vdd.n2922 vdd.t229 127.284
R16453 vdd.n2642 vdd.t274 127.284
R16454 vdd.n832 vdd.t256 127.284
R16455 vdd.n2639 vdd.t261 127.284
R16456 vdd.n799 vdd.t263 127.284
R16457 vdd.n1027 vdd.t270 127.284
R16458 vdd.n1027 vdd.t271 127.284
R16459 vdd.n22 vdd.n20 117.314
R16460 vdd.n17 vdd.n15 117.314
R16461 vdd.n27 vdd.n26 116.927
R16462 vdd.n24 vdd.n23 116.927
R16463 vdd.n22 vdd.n21 116.927
R16464 vdd.n17 vdd.n16 116.927
R16465 vdd.n19 vdd.n18 116.927
R16466 vdd.n27 vdd.n25 116.927
R16467 vdd.n2178 vdd.t266 111.188
R16468 vdd.n966 vdd.t253 111.188
R16469 vdd.n2152 vdd.t213 111.188
R16470 vdd.n958 vdd.t277 111.188
R16471 vdd.n2643 vdd.t273 111.188
R16472 vdd.n833 vdd.t257 111.188
R16473 vdd.n2640 vdd.t260 111.188
R16474 vdd.n800 vdd.t264 111.188
R16475 vdd.n2865 vdd.n911 99.5127
R16476 vdd.n2869 vdd.n911 99.5127
R16477 vdd.n2869 vdd.n903 99.5127
R16478 vdd.n2877 vdd.n903 99.5127
R16479 vdd.n2877 vdd.n901 99.5127
R16480 vdd.n2881 vdd.n901 99.5127
R16481 vdd.n2881 vdd.n890 99.5127
R16482 vdd.n2889 vdd.n890 99.5127
R16483 vdd.n2889 vdd.n888 99.5127
R16484 vdd.n2893 vdd.n888 99.5127
R16485 vdd.n2893 vdd.n879 99.5127
R16486 vdd.n2901 vdd.n879 99.5127
R16487 vdd.n2901 vdd.n877 99.5127
R16488 vdd.n2905 vdd.n877 99.5127
R16489 vdd.n2905 vdd.n867 99.5127
R16490 vdd.n2913 vdd.n867 99.5127
R16491 vdd.n2913 vdd.n865 99.5127
R16492 vdd.n2917 vdd.n865 99.5127
R16493 vdd.n2917 vdd.n856 99.5127
R16494 vdd.n2927 vdd.n856 99.5127
R16495 vdd.n2927 vdd.n854 99.5127
R16496 vdd.n2931 vdd.n854 99.5127
R16497 vdd.n2931 vdd.n842 99.5127
R16498 vdd.n2984 vdd.n842 99.5127
R16499 vdd.n2984 vdd.n840 99.5127
R16500 vdd.n2988 vdd.n840 99.5127
R16501 vdd.n2988 vdd.n808 99.5127
R16502 vdd.n3058 vdd.n808 99.5127
R16503 vdd.n3054 vdd.n809 99.5127
R16504 vdd.n3052 vdd.n3051 99.5127
R16505 vdd.n3049 vdd.n813 99.5127
R16506 vdd.n3045 vdd.n3044 99.5127
R16507 vdd.n3042 vdd.n816 99.5127
R16508 vdd.n3038 vdd.n3037 99.5127
R16509 vdd.n3035 vdd.n819 99.5127
R16510 vdd.n3031 vdd.n3030 99.5127
R16511 vdd.n3028 vdd.n3026 99.5127
R16512 vdd.n3024 vdd.n822 99.5127
R16513 vdd.n3020 vdd.n3019 99.5127
R16514 vdd.n3017 vdd.n825 99.5127
R16515 vdd.n3013 vdd.n3012 99.5127
R16516 vdd.n3010 vdd.n828 99.5127
R16517 vdd.n3006 vdd.n3005 99.5127
R16518 vdd.n3003 vdd.n831 99.5127
R16519 vdd.n2998 vdd.n2997 99.5127
R16520 vdd.n2785 vdd.n914 99.5127
R16521 vdd.n2785 vdd.n909 99.5127
R16522 vdd.n2782 vdd.n909 99.5127
R16523 vdd.n2782 vdd.n904 99.5127
R16524 vdd.n2729 vdd.n904 99.5127
R16525 vdd.n2729 vdd.n898 99.5127
R16526 vdd.n2732 vdd.n898 99.5127
R16527 vdd.n2732 vdd.n891 99.5127
R16528 vdd.n2735 vdd.n891 99.5127
R16529 vdd.n2735 vdd.n886 99.5127
R16530 vdd.n2738 vdd.n886 99.5127
R16531 vdd.n2738 vdd.n881 99.5127
R16532 vdd.n2741 vdd.n881 99.5127
R16533 vdd.n2741 vdd.n875 99.5127
R16534 vdd.n2759 vdd.n875 99.5127
R16535 vdd.n2759 vdd.n868 99.5127
R16536 vdd.n2755 vdd.n868 99.5127
R16537 vdd.n2755 vdd.n863 99.5127
R16538 vdd.n2752 vdd.n863 99.5127
R16539 vdd.n2752 vdd.n858 99.5127
R16540 vdd.n2749 vdd.n858 99.5127
R16541 vdd.n2749 vdd.n852 99.5127
R16542 vdd.n2746 vdd.n852 99.5127
R16543 vdd.n2746 vdd.n844 99.5127
R16544 vdd.n844 vdd.n837 99.5127
R16545 vdd.n2990 vdd.n837 99.5127
R16546 vdd.n2991 vdd.n2990 99.5127
R16547 vdd.n2991 vdd.n806 99.5127
R16548 vdd.n2855 vdd.n2638 99.5127
R16549 vdd.n2851 vdd.n2638 99.5127
R16550 vdd.n2849 vdd.n2848 99.5127
R16551 vdd.n2845 vdd.n2844 99.5127
R16552 vdd.n2841 vdd.n2840 99.5127
R16553 vdd.n2837 vdd.n2836 99.5127
R16554 vdd.n2833 vdd.n2832 99.5127
R16555 vdd.n2829 vdd.n2828 99.5127
R16556 vdd.n2825 vdd.n2824 99.5127
R16557 vdd.n2821 vdd.n2820 99.5127
R16558 vdd.n2817 vdd.n2816 99.5127
R16559 vdd.n2813 vdd.n2812 99.5127
R16560 vdd.n2809 vdd.n2808 99.5127
R16561 vdd.n2805 vdd.n2804 99.5127
R16562 vdd.n2801 vdd.n2800 99.5127
R16563 vdd.n2797 vdd.n2796 99.5127
R16564 vdd.n2792 vdd.n2791 99.5127
R16565 vdd.n2603 vdd.n955 99.5127
R16566 vdd.n2599 vdd.n2598 99.5127
R16567 vdd.n2595 vdd.n2594 99.5127
R16568 vdd.n2591 vdd.n2590 99.5127
R16569 vdd.n2587 vdd.n2586 99.5127
R16570 vdd.n2583 vdd.n2582 99.5127
R16571 vdd.n2579 vdd.n2578 99.5127
R16572 vdd.n2575 vdd.n2574 99.5127
R16573 vdd.n2571 vdd.n2570 99.5127
R16574 vdd.n2567 vdd.n2566 99.5127
R16575 vdd.n2563 vdd.n2562 99.5127
R16576 vdd.n2559 vdd.n2558 99.5127
R16577 vdd.n2555 vdd.n2554 99.5127
R16578 vdd.n2551 vdd.n2550 99.5127
R16579 vdd.n2547 vdd.n2546 99.5127
R16580 vdd.n2543 vdd.n2542 99.5127
R16581 vdd.n2538 vdd.n2537 99.5127
R16582 vdd.n2276 vdd.n1050 99.5127
R16583 vdd.n2276 vdd.n1044 99.5127
R16584 vdd.n2273 vdd.n1044 99.5127
R16585 vdd.n2273 vdd.n1038 99.5127
R16586 vdd.n2270 vdd.n1038 99.5127
R16587 vdd.n2270 vdd.n1031 99.5127
R16588 vdd.n2267 vdd.n1031 99.5127
R16589 vdd.n2267 vdd.n1024 99.5127
R16590 vdd.n2264 vdd.n1024 99.5127
R16591 vdd.n2264 vdd.n1019 99.5127
R16592 vdd.n2261 vdd.n1019 99.5127
R16593 vdd.n2261 vdd.n1013 99.5127
R16594 vdd.n2258 vdd.n1013 99.5127
R16595 vdd.n2258 vdd.n1006 99.5127
R16596 vdd.n2172 vdd.n1006 99.5127
R16597 vdd.n2172 vdd.n1000 99.5127
R16598 vdd.n2169 vdd.n1000 99.5127
R16599 vdd.n2169 vdd.n995 99.5127
R16600 vdd.n2166 vdd.n995 99.5127
R16601 vdd.n2166 vdd.n990 99.5127
R16602 vdd.n2163 vdd.n990 99.5127
R16603 vdd.n2163 vdd.n984 99.5127
R16604 vdd.n2160 vdd.n984 99.5127
R16605 vdd.n2160 vdd.n977 99.5127
R16606 vdd.n2157 vdd.n977 99.5127
R16607 vdd.n2157 vdd.n970 99.5127
R16608 vdd.n970 vdd.n960 99.5127
R16609 vdd.n2533 vdd.n960 99.5127
R16610 vdd.n2111 vdd.n2109 99.5127
R16611 vdd.n2115 vdd.n2109 99.5127
R16612 vdd.n2119 vdd.n2117 99.5127
R16613 vdd.n2123 vdd.n2107 99.5127
R16614 vdd.n2127 vdd.n2125 99.5127
R16615 vdd.n2131 vdd.n2105 99.5127
R16616 vdd.n2135 vdd.n2133 99.5127
R16617 vdd.n2139 vdd.n2103 99.5127
R16618 vdd.n2142 vdd.n2141 99.5127
R16619 vdd.n2312 vdd.n2310 99.5127
R16620 vdd.n2308 vdd.n2144 99.5127
R16621 vdd.n2304 vdd.n2302 99.5127
R16622 vdd.n2300 vdd.n2146 99.5127
R16623 vdd.n2296 vdd.n2294 99.5127
R16624 vdd.n2292 vdd.n2148 99.5127
R16625 vdd.n2288 vdd.n2286 99.5127
R16626 vdd.n2284 vdd.n2150 99.5127
R16627 vdd.n2376 vdd.n1046 99.5127
R16628 vdd.n2380 vdd.n1046 99.5127
R16629 vdd.n2380 vdd.n1036 99.5127
R16630 vdd.n2388 vdd.n1036 99.5127
R16631 vdd.n2388 vdd.n1034 99.5127
R16632 vdd.n2392 vdd.n1034 99.5127
R16633 vdd.n2392 vdd.n1023 99.5127
R16634 vdd.n2401 vdd.n1023 99.5127
R16635 vdd.n2401 vdd.n1021 99.5127
R16636 vdd.n2405 vdd.n1021 99.5127
R16637 vdd.n2405 vdd.n1011 99.5127
R16638 vdd.n2413 vdd.n1011 99.5127
R16639 vdd.n2413 vdd.n1009 99.5127
R16640 vdd.n2417 vdd.n1009 99.5127
R16641 vdd.n2417 vdd.n999 99.5127
R16642 vdd.n2425 vdd.n999 99.5127
R16643 vdd.n2425 vdd.n997 99.5127
R16644 vdd.n2429 vdd.n997 99.5127
R16645 vdd.n2429 vdd.n988 99.5127
R16646 vdd.n2437 vdd.n988 99.5127
R16647 vdd.n2437 vdd.n986 99.5127
R16648 vdd.n2441 vdd.n986 99.5127
R16649 vdd.n2441 vdd.n975 99.5127
R16650 vdd.n2451 vdd.n975 99.5127
R16651 vdd.n2451 vdd.n972 99.5127
R16652 vdd.n2456 vdd.n972 99.5127
R16653 vdd.n2456 vdd.n973 99.5127
R16654 vdd.n973 vdd.n954 99.5127
R16655 vdd.n2974 vdd.n2973 99.5127
R16656 vdd.n2971 vdd.n2937 99.5127
R16657 vdd.n2967 vdd.n2966 99.5127
R16658 vdd.n2964 vdd.n2940 99.5127
R16659 vdd.n2960 vdd.n2959 99.5127
R16660 vdd.n2957 vdd.n2943 99.5127
R16661 vdd.n2953 vdd.n2952 99.5127
R16662 vdd.n2950 vdd.n2947 99.5127
R16663 vdd.n3091 vdd.n787 99.5127
R16664 vdd.n3089 vdd.n3088 99.5127
R16665 vdd.n3086 vdd.n789 99.5127
R16666 vdd.n3082 vdd.n3081 99.5127
R16667 vdd.n3079 vdd.n792 99.5127
R16668 vdd.n3075 vdd.n3074 99.5127
R16669 vdd.n3072 vdd.n795 99.5127
R16670 vdd.n3068 vdd.n3067 99.5127
R16671 vdd.n3065 vdd.n798 99.5127
R16672 vdd.n2709 vdd.n915 99.5127
R16673 vdd.n2709 vdd.n910 99.5127
R16674 vdd.n2780 vdd.n910 99.5127
R16675 vdd.n2780 vdd.n905 99.5127
R16676 vdd.n2776 vdd.n905 99.5127
R16677 vdd.n2776 vdd.n899 99.5127
R16678 vdd.n2773 vdd.n899 99.5127
R16679 vdd.n2773 vdd.n892 99.5127
R16680 vdd.n2770 vdd.n892 99.5127
R16681 vdd.n2770 vdd.n887 99.5127
R16682 vdd.n2767 vdd.n887 99.5127
R16683 vdd.n2767 vdd.n882 99.5127
R16684 vdd.n2764 vdd.n882 99.5127
R16685 vdd.n2764 vdd.n876 99.5127
R16686 vdd.n2761 vdd.n876 99.5127
R16687 vdd.n2761 vdd.n869 99.5127
R16688 vdd.n2726 vdd.n869 99.5127
R16689 vdd.n2726 vdd.n864 99.5127
R16690 vdd.n2723 vdd.n864 99.5127
R16691 vdd.n2723 vdd.n859 99.5127
R16692 vdd.n2720 vdd.n859 99.5127
R16693 vdd.n2720 vdd.n853 99.5127
R16694 vdd.n2717 vdd.n853 99.5127
R16695 vdd.n2717 vdd.n845 99.5127
R16696 vdd.n2714 vdd.n845 99.5127
R16697 vdd.n2714 vdd.n838 99.5127
R16698 vdd.n838 vdd.n804 99.5127
R16699 vdd.n3060 vdd.n804 99.5127
R16700 vdd.n2859 vdd.n918 99.5127
R16701 vdd.n2647 vdd.n2646 99.5127
R16702 vdd.n2651 vdd.n2650 99.5127
R16703 vdd.n2655 vdd.n2654 99.5127
R16704 vdd.n2659 vdd.n2658 99.5127
R16705 vdd.n2663 vdd.n2662 99.5127
R16706 vdd.n2667 vdd.n2666 99.5127
R16707 vdd.n2671 vdd.n2670 99.5127
R16708 vdd.n2675 vdd.n2674 99.5127
R16709 vdd.n2679 vdd.n2678 99.5127
R16710 vdd.n2683 vdd.n2682 99.5127
R16711 vdd.n2687 vdd.n2686 99.5127
R16712 vdd.n2691 vdd.n2690 99.5127
R16713 vdd.n2695 vdd.n2694 99.5127
R16714 vdd.n2699 vdd.n2698 99.5127
R16715 vdd.n2703 vdd.n2702 99.5127
R16716 vdd.n2705 vdd.n2637 99.5127
R16717 vdd.n2863 vdd.n908 99.5127
R16718 vdd.n2871 vdd.n908 99.5127
R16719 vdd.n2871 vdd.n906 99.5127
R16720 vdd.n2875 vdd.n906 99.5127
R16721 vdd.n2875 vdd.n896 99.5127
R16722 vdd.n2883 vdd.n896 99.5127
R16723 vdd.n2883 vdd.n894 99.5127
R16724 vdd.n2887 vdd.n894 99.5127
R16725 vdd.n2887 vdd.n885 99.5127
R16726 vdd.n2895 vdd.n885 99.5127
R16727 vdd.n2895 vdd.n883 99.5127
R16728 vdd.n2899 vdd.n883 99.5127
R16729 vdd.n2899 vdd.n873 99.5127
R16730 vdd.n2907 vdd.n873 99.5127
R16731 vdd.n2907 vdd.n871 99.5127
R16732 vdd.n2911 vdd.n871 99.5127
R16733 vdd.n2911 vdd.n862 99.5127
R16734 vdd.n2919 vdd.n862 99.5127
R16735 vdd.n2919 vdd.n860 99.5127
R16736 vdd.n2925 vdd.n860 99.5127
R16737 vdd.n2925 vdd.n850 99.5127
R16738 vdd.n2933 vdd.n850 99.5127
R16739 vdd.n2933 vdd.n847 99.5127
R16740 vdd.n2982 vdd.n847 99.5127
R16741 vdd.n2982 vdd.n848 99.5127
R16742 vdd.n848 vdd.n839 99.5127
R16743 vdd.n2977 vdd.n839 99.5127
R16744 vdd.n2977 vdd.n807 99.5127
R16745 vdd.n2527 vdd.n2526 99.5127
R16746 vdd.n2523 vdd.n2522 99.5127
R16747 vdd.n2519 vdd.n2518 99.5127
R16748 vdd.n2515 vdd.n2514 99.5127
R16749 vdd.n2511 vdd.n2510 99.5127
R16750 vdd.n2507 vdd.n2506 99.5127
R16751 vdd.n2503 vdd.n2502 99.5127
R16752 vdd.n2499 vdd.n2498 99.5127
R16753 vdd.n2495 vdd.n2494 99.5127
R16754 vdd.n2491 vdd.n2490 99.5127
R16755 vdd.n2487 vdd.n2486 99.5127
R16756 vdd.n2483 vdd.n2482 99.5127
R16757 vdd.n2479 vdd.n2478 99.5127
R16758 vdd.n2475 vdd.n2474 99.5127
R16759 vdd.n2471 vdd.n2470 99.5127
R16760 vdd.n2467 vdd.n2466 99.5127
R16761 vdd.n2463 vdd.n936 99.5127
R16762 vdd.n2220 vdd.n1051 99.5127
R16763 vdd.n2220 vdd.n1045 99.5127
R16764 vdd.n2223 vdd.n1045 99.5127
R16765 vdd.n2223 vdd.n1039 99.5127
R16766 vdd.n2226 vdd.n1039 99.5127
R16767 vdd.n2226 vdd.n1032 99.5127
R16768 vdd.n2229 vdd.n1032 99.5127
R16769 vdd.n2229 vdd.n1025 99.5127
R16770 vdd.n2232 vdd.n1025 99.5127
R16771 vdd.n2232 vdd.n1020 99.5127
R16772 vdd.n2235 vdd.n1020 99.5127
R16773 vdd.n2235 vdd.n1014 99.5127
R16774 vdd.n2256 vdd.n1014 99.5127
R16775 vdd.n2256 vdd.n1007 99.5127
R16776 vdd.n2252 vdd.n1007 99.5127
R16777 vdd.n2252 vdd.n1001 99.5127
R16778 vdd.n2249 vdd.n1001 99.5127
R16779 vdd.n2249 vdd.n996 99.5127
R16780 vdd.n2246 vdd.n996 99.5127
R16781 vdd.n2246 vdd.n991 99.5127
R16782 vdd.n2243 vdd.n991 99.5127
R16783 vdd.n2243 vdd.n985 99.5127
R16784 vdd.n2240 vdd.n985 99.5127
R16785 vdd.n2240 vdd.n978 99.5127
R16786 vdd.n978 vdd.n969 99.5127
R16787 vdd.n2458 vdd.n969 99.5127
R16788 vdd.n2459 vdd.n2458 99.5127
R16789 vdd.n2459 vdd.n961 99.5127
R16790 vdd.n2370 vdd.n2368 99.5127
R16791 vdd.n2366 vdd.n1054 99.5127
R16792 vdd.n2362 vdd.n2360 99.5127
R16793 vdd.n2358 vdd.n1056 99.5127
R16794 vdd.n2354 vdd.n2352 99.5127
R16795 vdd.n2350 vdd.n1058 99.5127
R16796 vdd.n2346 vdd.n2344 99.5127
R16797 vdd.n2342 vdd.n1060 99.5127
R16798 vdd.n2184 vdd.n1062 99.5127
R16799 vdd.n2189 vdd.n2186 99.5127
R16800 vdd.n2193 vdd.n2191 99.5127
R16801 vdd.n2197 vdd.n2182 99.5127
R16802 vdd.n2201 vdd.n2199 99.5127
R16803 vdd.n2205 vdd.n2180 99.5127
R16804 vdd.n2209 vdd.n2207 99.5127
R16805 vdd.n2214 vdd.n2176 99.5127
R16806 vdd.n2217 vdd.n2216 99.5127
R16807 vdd.n2374 vdd.n1042 99.5127
R16808 vdd.n2382 vdd.n1042 99.5127
R16809 vdd.n2382 vdd.n1040 99.5127
R16810 vdd.n2386 vdd.n1040 99.5127
R16811 vdd.n2386 vdd.n1029 99.5127
R16812 vdd.n2394 vdd.n1029 99.5127
R16813 vdd.n2394 vdd.n1026 99.5127
R16814 vdd.n2399 vdd.n1026 99.5127
R16815 vdd.n2399 vdd.n1017 99.5127
R16816 vdd.n2407 vdd.n1017 99.5127
R16817 vdd.n2407 vdd.n1015 99.5127
R16818 vdd.n2411 vdd.n1015 99.5127
R16819 vdd.n2411 vdd.n1005 99.5127
R16820 vdd.n2419 vdd.n1005 99.5127
R16821 vdd.n2419 vdd.n1003 99.5127
R16822 vdd.n2423 vdd.n1003 99.5127
R16823 vdd.n2423 vdd.n994 99.5127
R16824 vdd.n2431 vdd.n994 99.5127
R16825 vdd.n2431 vdd.n992 99.5127
R16826 vdd.n2435 vdd.n992 99.5127
R16827 vdd.n2435 vdd.n982 99.5127
R16828 vdd.n2443 vdd.n982 99.5127
R16829 vdd.n2443 vdd.n979 99.5127
R16830 vdd.n2449 vdd.n979 99.5127
R16831 vdd.n2449 vdd.n980 99.5127
R16832 vdd.n980 vdd.n971 99.5127
R16833 vdd.n971 vdd.n962 99.5127
R16834 vdd.n2531 vdd.n962 99.5127
R16835 vdd.n9 vdd.n7 98.9633
R16836 vdd.n2 vdd.n0 98.9633
R16837 vdd.n9 vdd.n8 98.6055
R16838 vdd.n11 vdd.n10 98.6055
R16839 vdd.n13 vdd.n12 98.6055
R16840 vdd.n6 vdd.n5 98.6055
R16841 vdd.n4 vdd.n3 98.6055
R16842 vdd.n2 vdd.n1 98.6055
R16843 vdd.t144 vdd.n303 85.8723
R16844 vdd.t119 vdd.n244 85.8723
R16845 vdd.t134 vdd.n201 85.8723
R16846 vdd.t104 vdd.n142 85.8723
R16847 vdd.t83 vdd.n100 85.8723
R16848 vdd.t18 vdd.n41 85.8723
R16849 vdd.t164 vdd.n1722 85.8723
R16850 vdd.t50 vdd.n1781 85.8723
R16851 vdd.t149 vdd.n1620 85.8723
R16852 vdd.t26 vdd.n1679 85.8723
R16853 vdd.t22 vdd.n1519 85.8723
R16854 vdd.t84 vdd.n1578 85.8723
R16855 vdd.n2923 vdd.n2922 78.546
R16856 vdd.n2397 vdd.n1027 78.546
R16857 vdd.n290 vdd.n289 75.1835
R16858 vdd.n288 vdd.n287 75.1835
R16859 vdd.n286 vdd.n285 75.1835
R16860 vdd.n284 vdd.n283 75.1835
R16861 vdd.n282 vdd.n281 75.1835
R16862 vdd.n280 vdd.n279 75.1835
R16863 vdd.n278 vdd.n277 75.1835
R16864 vdd.n276 vdd.n275 75.1835
R16865 vdd.n274 vdd.n273 75.1835
R16866 vdd.n188 vdd.n187 75.1835
R16867 vdd.n186 vdd.n185 75.1835
R16868 vdd.n184 vdd.n183 75.1835
R16869 vdd.n182 vdd.n181 75.1835
R16870 vdd.n180 vdd.n179 75.1835
R16871 vdd.n178 vdd.n177 75.1835
R16872 vdd.n176 vdd.n175 75.1835
R16873 vdd.n174 vdd.n173 75.1835
R16874 vdd.n172 vdd.n171 75.1835
R16875 vdd.n87 vdd.n86 75.1835
R16876 vdd.n85 vdd.n84 75.1835
R16877 vdd.n83 vdd.n82 75.1835
R16878 vdd.n81 vdd.n80 75.1835
R16879 vdd.n79 vdd.n78 75.1835
R16880 vdd.n77 vdd.n76 75.1835
R16881 vdd.n75 vdd.n74 75.1835
R16882 vdd.n73 vdd.n72 75.1835
R16883 vdd.n71 vdd.n70 75.1835
R16884 vdd.n1752 vdd.n1751 75.1835
R16885 vdd.n1754 vdd.n1753 75.1835
R16886 vdd.n1756 vdd.n1755 75.1835
R16887 vdd.n1758 vdd.n1757 75.1835
R16888 vdd.n1760 vdd.n1759 75.1835
R16889 vdd.n1762 vdd.n1761 75.1835
R16890 vdd.n1764 vdd.n1763 75.1835
R16891 vdd.n1766 vdd.n1765 75.1835
R16892 vdd.n1768 vdd.n1767 75.1835
R16893 vdd.n1650 vdd.n1649 75.1835
R16894 vdd.n1652 vdd.n1651 75.1835
R16895 vdd.n1654 vdd.n1653 75.1835
R16896 vdd.n1656 vdd.n1655 75.1835
R16897 vdd.n1658 vdd.n1657 75.1835
R16898 vdd.n1660 vdd.n1659 75.1835
R16899 vdd.n1662 vdd.n1661 75.1835
R16900 vdd.n1664 vdd.n1663 75.1835
R16901 vdd.n1666 vdd.n1665 75.1835
R16902 vdd.n1549 vdd.n1548 75.1835
R16903 vdd.n1551 vdd.n1550 75.1835
R16904 vdd.n1553 vdd.n1552 75.1835
R16905 vdd.n1555 vdd.n1554 75.1835
R16906 vdd.n1557 vdd.n1556 75.1835
R16907 vdd.n1559 vdd.n1558 75.1835
R16908 vdd.n1561 vdd.n1560 75.1835
R16909 vdd.n1563 vdd.n1562 75.1835
R16910 vdd.n1565 vdd.n1564 75.1835
R16911 vdd.n2858 vdd.n2857 72.8958
R16912 vdd.n2857 vdd.n2621 72.8958
R16913 vdd.n2857 vdd.n2622 72.8958
R16914 vdd.n2857 vdd.n2623 72.8958
R16915 vdd.n2857 vdd.n2624 72.8958
R16916 vdd.n2857 vdd.n2625 72.8958
R16917 vdd.n2857 vdd.n2626 72.8958
R16918 vdd.n2857 vdd.n2627 72.8958
R16919 vdd.n2857 vdd.n2628 72.8958
R16920 vdd.n2857 vdd.n2629 72.8958
R16921 vdd.n2857 vdd.n2630 72.8958
R16922 vdd.n2857 vdd.n2631 72.8958
R16923 vdd.n2857 vdd.n2632 72.8958
R16924 vdd.n2857 vdd.n2633 72.8958
R16925 vdd.n2857 vdd.n2634 72.8958
R16926 vdd.n2857 vdd.n2635 72.8958
R16927 vdd.n2857 vdd.n2636 72.8958
R16928 vdd.n803 vdd.n692 72.8958
R16929 vdd.n3066 vdd.n692 72.8958
R16930 vdd.n797 vdd.n692 72.8958
R16931 vdd.n3073 vdd.n692 72.8958
R16932 vdd.n794 vdd.n692 72.8958
R16933 vdd.n3080 vdd.n692 72.8958
R16934 vdd.n791 vdd.n692 72.8958
R16935 vdd.n3087 vdd.n692 72.8958
R16936 vdd.n3090 vdd.n692 72.8958
R16937 vdd.n2946 vdd.n692 72.8958
R16938 vdd.n2951 vdd.n692 72.8958
R16939 vdd.n2945 vdd.n692 72.8958
R16940 vdd.n2958 vdd.n692 72.8958
R16941 vdd.n2942 vdd.n692 72.8958
R16942 vdd.n2965 vdd.n692 72.8958
R16943 vdd.n2939 vdd.n692 72.8958
R16944 vdd.n2972 vdd.n692 72.8958
R16945 vdd.n2110 vdd.n1049 72.8958
R16946 vdd.n2116 vdd.n1049 72.8958
R16947 vdd.n2118 vdd.n1049 72.8958
R16948 vdd.n2124 vdd.n1049 72.8958
R16949 vdd.n2126 vdd.n1049 72.8958
R16950 vdd.n2132 vdd.n1049 72.8958
R16951 vdd.n2134 vdd.n1049 72.8958
R16952 vdd.n2140 vdd.n1049 72.8958
R16953 vdd.n2311 vdd.n1049 72.8958
R16954 vdd.n2309 vdd.n1049 72.8958
R16955 vdd.n2303 vdd.n1049 72.8958
R16956 vdd.n2301 vdd.n1049 72.8958
R16957 vdd.n2295 vdd.n1049 72.8958
R16958 vdd.n2293 vdd.n1049 72.8958
R16959 vdd.n2287 vdd.n1049 72.8958
R16960 vdd.n2285 vdd.n1049 72.8958
R16961 vdd.n2279 vdd.n1049 72.8958
R16962 vdd.n2604 vdd.n937 72.8958
R16963 vdd.n2604 vdd.n938 72.8958
R16964 vdd.n2604 vdd.n939 72.8958
R16965 vdd.n2604 vdd.n940 72.8958
R16966 vdd.n2604 vdd.n941 72.8958
R16967 vdd.n2604 vdd.n942 72.8958
R16968 vdd.n2604 vdd.n943 72.8958
R16969 vdd.n2604 vdd.n944 72.8958
R16970 vdd.n2604 vdd.n945 72.8958
R16971 vdd.n2604 vdd.n946 72.8958
R16972 vdd.n2604 vdd.n947 72.8958
R16973 vdd.n2604 vdd.n948 72.8958
R16974 vdd.n2604 vdd.n949 72.8958
R16975 vdd.n2604 vdd.n950 72.8958
R16976 vdd.n2604 vdd.n951 72.8958
R16977 vdd.n2604 vdd.n952 72.8958
R16978 vdd.n2604 vdd.n953 72.8958
R16979 vdd.n2857 vdd.n2856 72.8958
R16980 vdd.n2857 vdd.n2605 72.8958
R16981 vdd.n2857 vdd.n2606 72.8958
R16982 vdd.n2857 vdd.n2607 72.8958
R16983 vdd.n2857 vdd.n2608 72.8958
R16984 vdd.n2857 vdd.n2609 72.8958
R16985 vdd.n2857 vdd.n2610 72.8958
R16986 vdd.n2857 vdd.n2611 72.8958
R16987 vdd.n2857 vdd.n2612 72.8958
R16988 vdd.n2857 vdd.n2613 72.8958
R16989 vdd.n2857 vdd.n2614 72.8958
R16990 vdd.n2857 vdd.n2615 72.8958
R16991 vdd.n2857 vdd.n2616 72.8958
R16992 vdd.n2857 vdd.n2617 72.8958
R16993 vdd.n2857 vdd.n2618 72.8958
R16994 vdd.n2857 vdd.n2619 72.8958
R16995 vdd.n2857 vdd.n2620 72.8958
R16996 vdd.n2996 vdd.n692 72.8958
R16997 vdd.n835 vdd.n692 72.8958
R16998 vdd.n3004 vdd.n692 72.8958
R16999 vdd.n830 vdd.n692 72.8958
R17000 vdd.n3011 vdd.n692 72.8958
R17001 vdd.n827 vdd.n692 72.8958
R17002 vdd.n3018 vdd.n692 72.8958
R17003 vdd.n824 vdd.n692 72.8958
R17004 vdd.n3025 vdd.n692 72.8958
R17005 vdd.n3029 vdd.n692 72.8958
R17006 vdd.n821 vdd.n692 72.8958
R17007 vdd.n3036 vdd.n692 72.8958
R17008 vdd.n818 vdd.n692 72.8958
R17009 vdd.n3043 vdd.n692 72.8958
R17010 vdd.n815 vdd.n692 72.8958
R17011 vdd.n3050 vdd.n692 72.8958
R17012 vdd.n3053 vdd.n692 72.8958
R17013 vdd.n2604 vdd.n935 72.8958
R17014 vdd.n2604 vdd.n934 72.8958
R17015 vdd.n2604 vdd.n933 72.8958
R17016 vdd.n2604 vdd.n932 72.8958
R17017 vdd.n2604 vdd.n931 72.8958
R17018 vdd.n2604 vdd.n930 72.8958
R17019 vdd.n2604 vdd.n929 72.8958
R17020 vdd.n2604 vdd.n928 72.8958
R17021 vdd.n2604 vdd.n927 72.8958
R17022 vdd.n2604 vdd.n926 72.8958
R17023 vdd.n2604 vdd.n925 72.8958
R17024 vdd.n2604 vdd.n924 72.8958
R17025 vdd.n2604 vdd.n923 72.8958
R17026 vdd.n2604 vdd.n922 72.8958
R17027 vdd.n2604 vdd.n921 72.8958
R17028 vdd.n2604 vdd.n920 72.8958
R17029 vdd.n2604 vdd.n919 72.8958
R17030 vdd.n2369 vdd.n1049 72.8958
R17031 vdd.n2367 vdd.n1049 72.8958
R17032 vdd.n2361 vdd.n1049 72.8958
R17033 vdd.n2359 vdd.n1049 72.8958
R17034 vdd.n2353 vdd.n1049 72.8958
R17035 vdd.n2351 vdd.n1049 72.8958
R17036 vdd.n2345 vdd.n1049 72.8958
R17037 vdd.n2343 vdd.n1049 72.8958
R17038 vdd.n1061 vdd.n1049 72.8958
R17039 vdd.n2185 vdd.n1049 72.8958
R17040 vdd.n2190 vdd.n1049 72.8958
R17041 vdd.n2192 vdd.n1049 72.8958
R17042 vdd.n2198 vdd.n1049 72.8958
R17043 vdd.n2200 vdd.n1049 72.8958
R17044 vdd.n2206 vdd.n1049 72.8958
R17045 vdd.n2208 vdd.n1049 72.8958
R17046 vdd.n2215 vdd.n1049 72.8958
R17047 vdd.n1419 vdd.n1418 66.2847
R17048 vdd.n1418 vdd.n1194 66.2847
R17049 vdd.n1418 vdd.n1195 66.2847
R17050 vdd.n1418 vdd.n1196 66.2847
R17051 vdd.n1418 vdd.n1197 66.2847
R17052 vdd.n1418 vdd.n1198 66.2847
R17053 vdd.n1418 vdd.n1199 66.2847
R17054 vdd.n1418 vdd.n1200 66.2847
R17055 vdd.n1418 vdd.n1201 66.2847
R17056 vdd.n1418 vdd.n1202 66.2847
R17057 vdd.n1418 vdd.n1203 66.2847
R17058 vdd.n1418 vdd.n1204 66.2847
R17059 vdd.n1418 vdd.n1205 66.2847
R17060 vdd.n1418 vdd.n1206 66.2847
R17061 vdd.n1418 vdd.n1207 66.2847
R17062 vdd.n1418 vdd.n1208 66.2847
R17063 vdd.n1418 vdd.n1209 66.2847
R17064 vdd.n1418 vdd.n1210 66.2847
R17065 vdd.n1418 vdd.n1211 66.2847
R17066 vdd.n1418 vdd.n1212 66.2847
R17067 vdd.n1418 vdd.n1213 66.2847
R17068 vdd.n1418 vdd.n1214 66.2847
R17069 vdd.n1418 vdd.n1215 66.2847
R17070 vdd.n1418 vdd.n1216 66.2847
R17071 vdd.n1418 vdd.n1217 66.2847
R17072 vdd.n1418 vdd.n1218 66.2847
R17073 vdd.n1418 vdd.n1219 66.2847
R17074 vdd.n1418 vdd.n1220 66.2847
R17075 vdd.n1418 vdd.n1221 66.2847
R17076 vdd.n1418 vdd.n1222 66.2847
R17077 vdd.n1418 vdd.n1223 66.2847
R17078 vdd.n1073 vdd.n1070 66.2847
R17079 vdd.n2000 vdd.n1073 66.2847
R17080 vdd.n2005 vdd.n1073 66.2847
R17081 vdd.n2010 vdd.n1073 66.2847
R17082 vdd.n1998 vdd.n1073 66.2847
R17083 vdd.n2017 vdd.n1073 66.2847
R17084 vdd.n1990 vdd.n1073 66.2847
R17085 vdd.n2024 vdd.n1073 66.2847
R17086 vdd.n1983 vdd.n1073 66.2847
R17087 vdd.n2031 vdd.n1073 66.2847
R17088 vdd.n1977 vdd.n1073 66.2847
R17089 vdd.n1972 vdd.n1073 66.2847
R17090 vdd.n2042 vdd.n1073 66.2847
R17091 vdd.n1964 vdd.n1073 66.2847
R17092 vdd.n2049 vdd.n1073 66.2847
R17093 vdd.n1957 vdd.n1073 66.2847
R17094 vdd.n2056 vdd.n1073 66.2847
R17095 vdd.n1950 vdd.n1073 66.2847
R17096 vdd.n2063 vdd.n1073 66.2847
R17097 vdd.n1943 vdd.n1073 66.2847
R17098 vdd.n2070 vdd.n1073 66.2847
R17099 vdd.n1937 vdd.n1073 66.2847
R17100 vdd.n1932 vdd.n1073 66.2847
R17101 vdd.n2081 vdd.n1073 66.2847
R17102 vdd.n1924 vdd.n1073 66.2847
R17103 vdd.n2088 vdd.n1073 66.2847
R17104 vdd.n1917 vdd.n1073 66.2847
R17105 vdd.n2095 vdd.n1073 66.2847
R17106 vdd.n2098 vdd.n1073 66.2847
R17107 vdd.n1908 vdd.n1073 66.2847
R17108 vdd.n2320 vdd.n1073 66.2847
R17109 vdd.n1902 vdd.n1073 66.2847
R17110 vdd.n3223 vdd.n3222 66.2847
R17111 vdd.n3223 vdd.n693 66.2847
R17112 vdd.n3223 vdd.n694 66.2847
R17113 vdd.n3223 vdd.n695 66.2847
R17114 vdd.n3223 vdd.n696 66.2847
R17115 vdd.n3223 vdd.n697 66.2847
R17116 vdd.n3223 vdd.n698 66.2847
R17117 vdd.n3223 vdd.n699 66.2847
R17118 vdd.n3223 vdd.n700 66.2847
R17119 vdd.n3223 vdd.n701 66.2847
R17120 vdd.n3223 vdd.n702 66.2847
R17121 vdd.n3223 vdd.n703 66.2847
R17122 vdd.n3223 vdd.n704 66.2847
R17123 vdd.n3223 vdd.n705 66.2847
R17124 vdd.n3223 vdd.n706 66.2847
R17125 vdd.n3223 vdd.n707 66.2847
R17126 vdd.n3223 vdd.n708 66.2847
R17127 vdd.n3223 vdd.n709 66.2847
R17128 vdd.n3223 vdd.n710 66.2847
R17129 vdd.n3223 vdd.n711 66.2847
R17130 vdd.n3223 vdd.n712 66.2847
R17131 vdd.n3223 vdd.n713 66.2847
R17132 vdd.n3223 vdd.n714 66.2847
R17133 vdd.n3223 vdd.n715 66.2847
R17134 vdd.n3223 vdd.n716 66.2847
R17135 vdd.n3223 vdd.n717 66.2847
R17136 vdd.n3223 vdd.n718 66.2847
R17137 vdd.n3223 vdd.n719 66.2847
R17138 vdd.n3223 vdd.n720 66.2847
R17139 vdd.n3223 vdd.n721 66.2847
R17140 vdd.n3223 vdd.n722 66.2847
R17141 vdd.n3354 vdd.n3353 66.2847
R17142 vdd.n3354 vdd.n424 66.2847
R17143 vdd.n3354 vdd.n423 66.2847
R17144 vdd.n3354 vdd.n422 66.2847
R17145 vdd.n3354 vdd.n421 66.2847
R17146 vdd.n3354 vdd.n420 66.2847
R17147 vdd.n3354 vdd.n419 66.2847
R17148 vdd.n3354 vdd.n418 66.2847
R17149 vdd.n3354 vdd.n417 66.2847
R17150 vdd.n3354 vdd.n416 66.2847
R17151 vdd.n3354 vdd.n415 66.2847
R17152 vdd.n3354 vdd.n414 66.2847
R17153 vdd.n3354 vdd.n413 66.2847
R17154 vdd.n3354 vdd.n412 66.2847
R17155 vdd.n3354 vdd.n411 66.2847
R17156 vdd.n3354 vdd.n410 66.2847
R17157 vdd.n3354 vdd.n409 66.2847
R17158 vdd.n3354 vdd.n408 66.2847
R17159 vdd.n3354 vdd.n407 66.2847
R17160 vdd.n3354 vdd.n406 66.2847
R17161 vdd.n3354 vdd.n405 66.2847
R17162 vdd.n3354 vdd.n404 66.2847
R17163 vdd.n3354 vdd.n403 66.2847
R17164 vdd.n3354 vdd.n402 66.2847
R17165 vdd.n3354 vdd.n401 66.2847
R17166 vdd.n3354 vdd.n400 66.2847
R17167 vdd.n3354 vdd.n399 66.2847
R17168 vdd.n3354 vdd.n398 66.2847
R17169 vdd.n3354 vdd.n397 66.2847
R17170 vdd.n3354 vdd.n396 66.2847
R17171 vdd.n3354 vdd.n395 66.2847
R17172 vdd.n3354 vdd.n394 66.2847
R17173 vdd.n467 vdd.n394 52.4337
R17174 vdd.n473 vdd.n395 52.4337
R17175 vdd.n477 vdd.n396 52.4337
R17176 vdd.n483 vdd.n397 52.4337
R17177 vdd.n487 vdd.n398 52.4337
R17178 vdd.n493 vdd.n399 52.4337
R17179 vdd.n497 vdd.n400 52.4337
R17180 vdd.n503 vdd.n401 52.4337
R17181 vdd.n507 vdd.n402 52.4337
R17182 vdd.n513 vdd.n403 52.4337
R17183 vdd.n517 vdd.n404 52.4337
R17184 vdd.n523 vdd.n405 52.4337
R17185 vdd.n527 vdd.n406 52.4337
R17186 vdd.n533 vdd.n407 52.4337
R17187 vdd.n537 vdd.n408 52.4337
R17188 vdd.n543 vdd.n409 52.4337
R17189 vdd.n547 vdd.n410 52.4337
R17190 vdd.n553 vdd.n411 52.4337
R17191 vdd.n557 vdd.n412 52.4337
R17192 vdd.n563 vdd.n413 52.4337
R17193 vdd.n567 vdd.n414 52.4337
R17194 vdd.n573 vdd.n415 52.4337
R17195 vdd.n577 vdd.n416 52.4337
R17196 vdd.n583 vdd.n417 52.4337
R17197 vdd.n587 vdd.n418 52.4337
R17198 vdd.n593 vdd.n419 52.4337
R17199 vdd.n597 vdd.n420 52.4337
R17200 vdd.n603 vdd.n421 52.4337
R17201 vdd.n607 vdd.n422 52.4337
R17202 vdd.n613 vdd.n423 52.4337
R17203 vdd.n616 vdd.n424 52.4337
R17204 vdd.n3353 vdd.n3352 52.4337
R17205 vdd.n3222 vdd.n3221 52.4337
R17206 vdd.n728 vdd.n693 52.4337
R17207 vdd.n734 vdd.n694 52.4337
R17208 vdd.n3211 vdd.n695 52.4337
R17209 vdd.n3207 vdd.n696 52.4337
R17210 vdd.n3203 vdd.n697 52.4337
R17211 vdd.n3199 vdd.n698 52.4337
R17212 vdd.n3195 vdd.n699 52.4337
R17213 vdd.n3191 vdd.n700 52.4337
R17214 vdd.n3187 vdd.n701 52.4337
R17215 vdd.n3179 vdd.n702 52.4337
R17216 vdd.n3175 vdd.n703 52.4337
R17217 vdd.n3171 vdd.n704 52.4337
R17218 vdd.n3167 vdd.n705 52.4337
R17219 vdd.n3163 vdd.n706 52.4337
R17220 vdd.n3159 vdd.n707 52.4337
R17221 vdd.n3155 vdd.n708 52.4337
R17222 vdd.n3151 vdd.n709 52.4337
R17223 vdd.n3147 vdd.n710 52.4337
R17224 vdd.n3143 vdd.n711 52.4337
R17225 vdd.n3139 vdd.n712 52.4337
R17226 vdd.n3133 vdd.n713 52.4337
R17227 vdd.n3129 vdd.n714 52.4337
R17228 vdd.n3125 vdd.n715 52.4337
R17229 vdd.n3121 vdd.n716 52.4337
R17230 vdd.n3117 vdd.n717 52.4337
R17231 vdd.n3113 vdd.n718 52.4337
R17232 vdd.n3109 vdd.n719 52.4337
R17233 vdd.n3105 vdd.n720 52.4337
R17234 vdd.n3101 vdd.n721 52.4337
R17235 vdd.n3097 vdd.n722 52.4337
R17236 vdd.n2322 vdd.n1902 52.4337
R17237 vdd.n2320 vdd.n2319 52.4337
R17238 vdd.n1909 vdd.n1908 52.4337
R17239 vdd.n2098 vdd.n2097 52.4337
R17240 vdd.n2095 vdd.n2094 52.4337
R17241 vdd.n2090 vdd.n1917 52.4337
R17242 vdd.n2088 vdd.n2087 52.4337
R17243 vdd.n2083 vdd.n1924 52.4337
R17244 vdd.n2081 vdd.n2080 52.4337
R17245 vdd.n1933 vdd.n1932 52.4337
R17246 vdd.n2072 vdd.n1937 52.4337
R17247 vdd.n2070 vdd.n2069 52.4337
R17248 vdd.n2065 vdd.n1943 52.4337
R17249 vdd.n2063 vdd.n2062 52.4337
R17250 vdd.n2058 vdd.n1950 52.4337
R17251 vdd.n2056 vdd.n2055 52.4337
R17252 vdd.n2051 vdd.n1957 52.4337
R17253 vdd.n2049 vdd.n2048 52.4337
R17254 vdd.n2044 vdd.n1964 52.4337
R17255 vdd.n2042 vdd.n2041 52.4337
R17256 vdd.n1973 vdd.n1972 52.4337
R17257 vdd.n2033 vdd.n1977 52.4337
R17258 vdd.n2031 vdd.n2030 52.4337
R17259 vdd.n2026 vdd.n1983 52.4337
R17260 vdd.n2024 vdd.n2023 52.4337
R17261 vdd.n2019 vdd.n1990 52.4337
R17262 vdd.n2017 vdd.n2016 52.4337
R17263 vdd.n2012 vdd.n1998 52.4337
R17264 vdd.n2010 vdd.n2009 52.4337
R17265 vdd.n2005 vdd.n2004 52.4337
R17266 vdd.n2000 vdd.n1999 52.4337
R17267 vdd.n2331 vdd.n1070 52.4337
R17268 vdd.n1420 vdd.n1419 52.4337
R17269 vdd.n1226 vdd.n1194 52.4337
R17270 vdd.n1230 vdd.n1195 52.4337
R17271 vdd.n1232 vdd.n1196 52.4337
R17272 vdd.n1236 vdd.n1197 52.4337
R17273 vdd.n1238 vdd.n1198 52.4337
R17274 vdd.n1242 vdd.n1199 52.4337
R17275 vdd.n1244 vdd.n1200 52.4337
R17276 vdd.n1248 vdd.n1201 52.4337
R17277 vdd.n1250 vdd.n1202 52.4337
R17278 vdd.n1256 vdd.n1203 52.4337
R17279 vdd.n1258 vdd.n1204 52.4337
R17280 vdd.n1262 vdd.n1205 52.4337
R17281 vdd.n1264 vdd.n1206 52.4337
R17282 vdd.n1268 vdd.n1207 52.4337
R17283 vdd.n1270 vdd.n1208 52.4337
R17284 vdd.n1274 vdd.n1209 52.4337
R17285 vdd.n1276 vdd.n1210 52.4337
R17286 vdd.n1280 vdd.n1211 52.4337
R17287 vdd.n1282 vdd.n1212 52.4337
R17288 vdd.n1354 vdd.n1213 52.4337
R17289 vdd.n1287 vdd.n1214 52.4337
R17290 vdd.n1291 vdd.n1215 52.4337
R17291 vdd.n1293 vdd.n1216 52.4337
R17292 vdd.n1297 vdd.n1217 52.4337
R17293 vdd.n1299 vdd.n1218 52.4337
R17294 vdd.n1303 vdd.n1219 52.4337
R17295 vdd.n1305 vdd.n1220 52.4337
R17296 vdd.n1309 vdd.n1221 52.4337
R17297 vdd.n1311 vdd.n1222 52.4337
R17298 vdd.n1315 vdd.n1223 52.4337
R17299 vdd.n1419 vdd.n1193 52.4337
R17300 vdd.n1229 vdd.n1194 52.4337
R17301 vdd.n1231 vdd.n1195 52.4337
R17302 vdd.n1235 vdd.n1196 52.4337
R17303 vdd.n1237 vdd.n1197 52.4337
R17304 vdd.n1241 vdd.n1198 52.4337
R17305 vdd.n1243 vdd.n1199 52.4337
R17306 vdd.n1247 vdd.n1200 52.4337
R17307 vdd.n1249 vdd.n1201 52.4337
R17308 vdd.n1255 vdd.n1202 52.4337
R17309 vdd.n1257 vdd.n1203 52.4337
R17310 vdd.n1261 vdd.n1204 52.4337
R17311 vdd.n1263 vdd.n1205 52.4337
R17312 vdd.n1267 vdd.n1206 52.4337
R17313 vdd.n1269 vdd.n1207 52.4337
R17314 vdd.n1273 vdd.n1208 52.4337
R17315 vdd.n1275 vdd.n1209 52.4337
R17316 vdd.n1279 vdd.n1210 52.4337
R17317 vdd.n1281 vdd.n1211 52.4337
R17318 vdd.n1285 vdd.n1212 52.4337
R17319 vdd.n1286 vdd.n1213 52.4337
R17320 vdd.n1290 vdd.n1214 52.4337
R17321 vdd.n1292 vdd.n1215 52.4337
R17322 vdd.n1296 vdd.n1216 52.4337
R17323 vdd.n1298 vdd.n1217 52.4337
R17324 vdd.n1302 vdd.n1218 52.4337
R17325 vdd.n1304 vdd.n1219 52.4337
R17326 vdd.n1308 vdd.n1220 52.4337
R17327 vdd.n1310 vdd.n1221 52.4337
R17328 vdd.n1314 vdd.n1222 52.4337
R17329 vdd.n1316 vdd.n1223 52.4337
R17330 vdd.n1070 vdd.n1069 52.4337
R17331 vdd.n2001 vdd.n2000 52.4337
R17332 vdd.n2006 vdd.n2005 52.4337
R17333 vdd.n2011 vdd.n2010 52.4337
R17334 vdd.n1998 vdd.n1991 52.4337
R17335 vdd.n2018 vdd.n2017 52.4337
R17336 vdd.n1990 vdd.n1984 52.4337
R17337 vdd.n2025 vdd.n2024 52.4337
R17338 vdd.n1983 vdd.n1978 52.4337
R17339 vdd.n2032 vdd.n2031 52.4337
R17340 vdd.n1977 vdd.n1976 52.4337
R17341 vdd.n1972 vdd.n1965 52.4337
R17342 vdd.n2043 vdd.n2042 52.4337
R17343 vdd.n1964 vdd.n1958 52.4337
R17344 vdd.n2050 vdd.n2049 52.4337
R17345 vdd.n1957 vdd.n1951 52.4337
R17346 vdd.n2057 vdd.n2056 52.4337
R17347 vdd.n1950 vdd.n1944 52.4337
R17348 vdd.n2064 vdd.n2063 52.4337
R17349 vdd.n1943 vdd.n1938 52.4337
R17350 vdd.n2071 vdd.n2070 52.4337
R17351 vdd.n1937 vdd.n1936 52.4337
R17352 vdd.n1932 vdd.n1925 52.4337
R17353 vdd.n2082 vdd.n2081 52.4337
R17354 vdd.n1924 vdd.n1918 52.4337
R17355 vdd.n2089 vdd.n2088 52.4337
R17356 vdd.n1917 vdd.n1911 52.4337
R17357 vdd.n2096 vdd.n2095 52.4337
R17358 vdd.n2099 vdd.n2098 52.4337
R17359 vdd.n1908 vdd.n1903 52.4337
R17360 vdd.n2321 vdd.n2320 52.4337
R17361 vdd.n1902 vdd.n1075 52.4337
R17362 vdd.n3222 vdd.n725 52.4337
R17363 vdd.n733 vdd.n693 52.4337
R17364 vdd.n3212 vdd.n694 52.4337
R17365 vdd.n3208 vdd.n695 52.4337
R17366 vdd.n3204 vdd.n696 52.4337
R17367 vdd.n3200 vdd.n697 52.4337
R17368 vdd.n3196 vdd.n698 52.4337
R17369 vdd.n3192 vdd.n699 52.4337
R17370 vdd.n3188 vdd.n700 52.4337
R17371 vdd.n3178 vdd.n701 52.4337
R17372 vdd.n3176 vdd.n702 52.4337
R17373 vdd.n3172 vdd.n703 52.4337
R17374 vdd.n3168 vdd.n704 52.4337
R17375 vdd.n3164 vdd.n705 52.4337
R17376 vdd.n3160 vdd.n706 52.4337
R17377 vdd.n3156 vdd.n707 52.4337
R17378 vdd.n3152 vdd.n708 52.4337
R17379 vdd.n3148 vdd.n709 52.4337
R17380 vdd.n3144 vdd.n710 52.4337
R17381 vdd.n3140 vdd.n711 52.4337
R17382 vdd.n3132 vdd.n712 52.4337
R17383 vdd.n3130 vdd.n713 52.4337
R17384 vdd.n3126 vdd.n714 52.4337
R17385 vdd.n3122 vdd.n715 52.4337
R17386 vdd.n3118 vdd.n716 52.4337
R17387 vdd.n3114 vdd.n717 52.4337
R17388 vdd.n3110 vdd.n718 52.4337
R17389 vdd.n3106 vdd.n719 52.4337
R17390 vdd.n3102 vdd.n720 52.4337
R17391 vdd.n3098 vdd.n721 52.4337
R17392 vdd.n722 vdd.n691 52.4337
R17393 vdd.n3353 vdd.n425 52.4337
R17394 vdd.n614 vdd.n424 52.4337
R17395 vdd.n608 vdd.n423 52.4337
R17396 vdd.n604 vdd.n422 52.4337
R17397 vdd.n598 vdd.n421 52.4337
R17398 vdd.n594 vdd.n420 52.4337
R17399 vdd.n588 vdd.n419 52.4337
R17400 vdd.n584 vdd.n418 52.4337
R17401 vdd.n578 vdd.n417 52.4337
R17402 vdd.n574 vdd.n416 52.4337
R17403 vdd.n568 vdd.n415 52.4337
R17404 vdd.n564 vdd.n414 52.4337
R17405 vdd.n558 vdd.n413 52.4337
R17406 vdd.n554 vdd.n412 52.4337
R17407 vdd.n548 vdd.n411 52.4337
R17408 vdd.n544 vdd.n410 52.4337
R17409 vdd.n538 vdd.n409 52.4337
R17410 vdd.n534 vdd.n408 52.4337
R17411 vdd.n528 vdd.n407 52.4337
R17412 vdd.n524 vdd.n406 52.4337
R17413 vdd.n518 vdd.n405 52.4337
R17414 vdd.n514 vdd.n404 52.4337
R17415 vdd.n508 vdd.n403 52.4337
R17416 vdd.n504 vdd.n402 52.4337
R17417 vdd.n498 vdd.n401 52.4337
R17418 vdd.n494 vdd.n400 52.4337
R17419 vdd.n488 vdd.n399 52.4337
R17420 vdd.n484 vdd.n398 52.4337
R17421 vdd.n478 vdd.n397 52.4337
R17422 vdd.n474 vdd.n396 52.4337
R17423 vdd.n468 vdd.n395 52.4337
R17424 vdd.n394 vdd.n392 52.4337
R17425 vdd.t294 vdd.t196 51.4683
R17426 vdd.n274 vdd.n272 42.0461
R17427 vdd.n172 vdd.n170 42.0461
R17428 vdd.n71 vdd.n69 42.0461
R17429 vdd.n1752 vdd.n1750 42.0461
R17430 vdd.n1650 vdd.n1648 42.0461
R17431 vdd.n1549 vdd.n1547 42.0461
R17432 vdd.n332 vdd.n331 41.6884
R17433 vdd.n230 vdd.n229 41.6884
R17434 vdd.n129 vdd.n128 41.6884
R17435 vdd.n1810 vdd.n1809 41.6884
R17436 vdd.n1708 vdd.n1707 41.6884
R17437 vdd.n1607 vdd.n1606 41.6884
R17438 vdd.n1319 vdd.n1318 41.1157
R17439 vdd.n1357 vdd.n1356 41.1157
R17440 vdd.n1253 vdd.n1252 41.1157
R17441 vdd.n428 vdd.n427 41.1157
R17442 vdd.n566 vdd.n441 41.1157
R17443 vdd.n454 vdd.n453 41.1157
R17444 vdd.n3053 vdd.n3052 39.2114
R17445 vdd.n3050 vdd.n3049 39.2114
R17446 vdd.n3045 vdd.n815 39.2114
R17447 vdd.n3043 vdd.n3042 39.2114
R17448 vdd.n3038 vdd.n818 39.2114
R17449 vdd.n3036 vdd.n3035 39.2114
R17450 vdd.n3031 vdd.n821 39.2114
R17451 vdd.n3029 vdd.n3028 39.2114
R17452 vdd.n3025 vdd.n3024 39.2114
R17453 vdd.n3020 vdd.n824 39.2114
R17454 vdd.n3018 vdd.n3017 39.2114
R17455 vdd.n3013 vdd.n827 39.2114
R17456 vdd.n3011 vdd.n3010 39.2114
R17457 vdd.n3006 vdd.n830 39.2114
R17458 vdd.n3004 vdd.n3003 39.2114
R17459 vdd.n2998 vdd.n835 39.2114
R17460 vdd.n2996 vdd.n2995 39.2114
R17461 vdd.n2856 vdd.n913 39.2114
R17462 vdd.n2851 vdd.n2605 39.2114
R17463 vdd.n2848 vdd.n2606 39.2114
R17464 vdd.n2844 vdd.n2607 39.2114
R17465 vdd.n2840 vdd.n2608 39.2114
R17466 vdd.n2836 vdd.n2609 39.2114
R17467 vdd.n2832 vdd.n2610 39.2114
R17468 vdd.n2828 vdd.n2611 39.2114
R17469 vdd.n2824 vdd.n2612 39.2114
R17470 vdd.n2820 vdd.n2613 39.2114
R17471 vdd.n2816 vdd.n2614 39.2114
R17472 vdd.n2812 vdd.n2615 39.2114
R17473 vdd.n2808 vdd.n2616 39.2114
R17474 vdd.n2804 vdd.n2617 39.2114
R17475 vdd.n2800 vdd.n2618 39.2114
R17476 vdd.n2796 vdd.n2619 39.2114
R17477 vdd.n2791 vdd.n2620 39.2114
R17478 vdd.n2599 vdd.n953 39.2114
R17479 vdd.n2595 vdd.n952 39.2114
R17480 vdd.n2591 vdd.n951 39.2114
R17481 vdd.n2587 vdd.n950 39.2114
R17482 vdd.n2583 vdd.n949 39.2114
R17483 vdd.n2579 vdd.n948 39.2114
R17484 vdd.n2575 vdd.n947 39.2114
R17485 vdd.n2571 vdd.n946 39.2114
R17486 vdd.n2567 vdd.n945 39.2114
R17487 vdd.n2563 vdd.n944 39.2114
R17488 vdd.n2559 vdd.n943 39.2114
R17489 vdd.n2555 vdd.n942 39.2114
R17490 vdd.n2551 vdd.n941 39.2114
R17491 vdd.n2547 vdd.n940 39.2114
R17492 vdd.n2543 vdd.n939 39.2114
R17493 vdd.n2538 vdd.n938 39.2114
R17494 vdd.n2534 vdd.n937 39.2114
R17495 vdd.n2110 vdd.n1048 39.2114
R17496 vdd.n2116 vdd.n2115 39.2114
R17497 vdd.n2119 vdd.n2118 39.2114
R17498 vdd.n2124 vdd.n2123 39.2114
R17499 vdd.n2127 vdd.n2126 39.2114
R17500 vdd.n2132 vdd.n2131 39.2114
R17501 vdd.n2135 vdd.n2134 39.2114
R17502 vdd.n2140 vdd.n2139 39.2114
R17503 vdd.n2311 vdd.n2142 39.2114
R17504 vdd.n2310 vdd.n2309 39.2114
R17505 vdd.n2303 vdd.n2144 39.2114
R17506 vdd.n2302 vdd.n2301 39.2114
R17507 vdd.n2295 vdd.n2146 39.2114
R17508 vdd.n2294 vdd.n2293 39.2114
R17509 vdd.n2287 vdd.n2148 39.2114
R17510 vdd.n2286 vdd.n2285 39.2114
R17511 vdd.n2279 vdd.n2150 39.2114
R17512 vdd.n2972 vdd.n2971 39.2114
R17513 vdd.n2967 vdd.n2939 39.2114
R17514 vdd.n2965 vdd.n2964 39.2114
R17515 vdd.n2960 vdd.n2942 39.2114
R17516 vdd.n2958 vdd.n2957 39.2114
R17517 vdd.n2953 vdd.n2945 39.2114
R17518 vdd.n2951 vdd.n2950 39.2114
R17519 vdd.n2946 vdd.n787 39.2114
R17520 vdd.n3090 vdd.n3089 39.2114
R17521 vdd.n3087 vdd.n3086 39.2114
R17522 vdd.n3082 vdd.n791 39.2114
R17523 vdd.n3080 vdd.n3079 39.2114
R17524 vdd.n3075 vdd.n794 39.2114
R17525 vdd.n3073 vdd.n3072 39.2114
R17526 vdd.n3068 vdd.n797 39.2114
R17527 vdd.n3066 vdd.n3065 39.2114
R17528 vdd.n3061 vdd.n803 39.2114
R17529 vdd.n2858 vdd.n916 39.2114
R17530 vdd.n2621 vdd.n918 39.2114
R17531 vdd.n2647 vdd.n2622 39.2114
R17532 vdd.n2651 vdd.n2623 39.2114
R17533 vdd.n2655 vdd.n2624 39.2114
R17534 vdd.n2659 vdd.n2625 39.2114
R17535 vdd.n2663 vdd.n2626 39.2114
R17536 vdd.n2667 vdd.n2627 39.2114
R17537 vdd.n2671 vdd.n2628 39.2114
R17538 vdd.n2675 vdd.n2629 39.2114
R17539 vdd.n2679 vdd.n2630 39.2114
R17540 vdd.n2683 vdd.n2631 39.2114
R17541 vdd.n2687 vdd.n2632 39.2114
R17542 vdd.n2691 vdd.n2633 39.2114
R17543 vdd.n2695 vdd.n2634 39.2114
R17544 vdd.n2699 vdd.n2635 39.2114
R17545 vdd.n2703 vdd.n2636 39.2114
R17546 vdd.n2859 vdd.n2858 39.2114
R17547 vdd.n2646 vdd.n2621 39.2114
R17548 vdd.n2650 vdd.n2622 39.2114
R17549 vdd.n2654 vdd.n2623 39.2114
R17550 vdd.n2658 vdd.n2624 39.2114
R17551 vdd.n2662 vdd.n2625 39.2114
R17552 vdd.n2666 vdd.n2626 39.2114
R17553 vdd.n2670 vdd.n2627 39.2114
R17554 vdd.n2674 vdd.n2628 39.2114
R17555 vdd.n2678 vdd.n2629 39.2114
R17556 vdd.n2682 vdd.n2630 39.2114
R17557 vdd.n2686 vdd.n2631 39.2114
R17558 vdd.n2690 vdd.n2632 39.2114
R17559 vdd.n2694 vdd.n2633 39.2114
R17560 vdd.n2698 vdd.n2634 39.2114
R17561 vdd.n2702 vdd.n2635 39.2114
R17562 vdd.n2705 vdd.n2636 39.2114
R17563 vdd.n803 vdd.n798 39.2114
R17564 vdd.n3067 vdd.n3066 39.2114
R17565 vdd.n797 vdd.n795 39.2114
R17566 vdd.n3074 vdd.n3073 39.2114
R17567 vdd.n794 vdd.n792 39.2114
R17568 vdd.n3081 vdd.n3080 39.2114
R17569 vdd.n791 vdd.n789 39.2114
R17570 vdd.n3088 vdd.n3087 39.2114
R17571 vdd.n3091 vdd.n3090 39.2114
R17572 vdd.n2947 vdd.n2946 39.2114
R17573 vdd.n2952 vdd.n2951 39.2114
R17574 vdd.n2945 vdd.n2943 39.2114
R17575 vdd.n2959 vdd.n2958 39.2114
R17576 vdd.n2942 vdd.n2940 39.2114
R17577 vdd.n2966 vdd.n2965 39.2114
R17578 vdd.n2939 vdd.n2937 39.2114
R17579 vdd.n2973 vdd.n2972 39.2114
R17580 vdd.n2111 vdd.n2110 39.2114
R17581 vdd.n2117 vdd.n2116 39.2114
R17582 vdd.n2118 vdd.n2107 39.2114
R17583 vdd.n2125 vdd.n2124 39.2114
R17584 vdd.n2126 vdd.n2105 39.2114
R17585 vdd.n2133 vdd.n2132 39.2114
R17586 vdd.n2134 vdd.n2103 39.2114
R17587 vdd.n2141 vdd.n2140 39.2114
R17588 vdd.n2312 vdd.n2311 39.2114
R17589 vdd.n2309 vdd.n2308 39.2114
R17590 vdd.n2304 vdd.n2303 39.2114
R17591 vdd.n2301 vdd.n2300 39.2114
R17592 vdd.n2296 vdd.n2295 39.2114
R17593 vdd.n2293 vdd.n2292 39.2114
R17594 vdd.n2288 vdd.n2287 39.2114
R17595 vdd.n2285 vdd.n2284 39.2114
R17596 vdd.n2280 vdd.n2279 39.2114
R17597 vdd.n2537 vdd.n937 39.2114
R17598 vdd.n2542 vdd.n938 39.2114
R17599 vdd.n2546 vdd.n939 39.2114
R17600 vdd.n2550 vdd.n940 39.2114
R17601 vdd.n2554 vdd.n941 39.2114
R17602 vdd.n2558 vdd.n942 39.2114
R17603 vdd.n2562 vdd.n943 39.2114
R17604 vdd.n2566 vdd.n944 39.2114
R17605 vdd.n2570 vdd.n945 39.2114
R17606 vdd.n2574 vdd.n946 39.2114
R17607 vdd.n2578 vdd.n947 39.2114
R17608 vdd.n2582 vdd.n948 39.2114
R17609 vdd.n2586 vdd.n949 39.2114
R17610 vdd.n2590 vdd.n950 39.2114
R17611 vdd.n2594 vdd.n951 39.2114
R17612 vdd.n2598 vdd.n952 39.2114
R17613 vdd.n955 vdd.n953 39.2114
R17614 vdd.n2856 vdd.n2855 39.2114
R17615 vdd.n2849 vdd.n2605 39.2114
R17616 vdd.n2845 vdd.n2606 39.2114
R17617 vdd.n2841 vdd.n2607 39.2114
R17618 vdd.n2837 vdd.n2608 39.2114
R17619 vdd.n2833 vdd.n2609 39.2114
R17620 vdd.n2829 vdd.n2610 39.2114
R17621 vdd.n2825 vdd.n2611 39.2114
R17622 vdd.n2821 vdd.n2612 39.2114
R17623 vdd.n2817 vdd.n2613 39.2114
R17624 vdd.n2813 vdd.n2614 39.2114
R17625 vdd.n2809 vdd.n2615 39.2114
R17626 vdd.n2805 vdd.n2616 39.2114
R17627 vdd.n2801 vdd.n2617 39.2114
R17628 vdd.n2797 vdd.n2618 39.2114
R17629 vdd.n2792 vdd.n2619 39.2114
R17630 vdd.n2788 vdd.n2620 39.2114
R17631 vdd.n2997 vdd.n2996 39.2114
R17632 vdd.n835 vdd.n831 39.2114
R17633 vdd.n3005 vdd.n3004 39.2114
R17634 vdd.n830 vdd.n828 39.2114
R17635 vdd.n3012 vdd.n3011 39.2114
R17636 vdd.n827 vdd.n825 39.2114
R17637 vdd.n3019 vdd.n3018 39.2114
R17638 vdd.n824 vdd.n822 39.2114
R17639 vdd.n3026 vdd.n3025 39.2114
R17640 vdd.n3030 vdd.n3029 39.2114
R17641 vdd.n821 vdd.n819 39.2114
R17642 vdd.n3037 vdd.n3036 39.2114
R17643 vdd.n818 vdd.n816 39.2114
R17644 vdd.n3044 vdd.n3043 39.2114
R17645 vdd.n815 vdd.n813 39.2114
R17646 vdd.n3051 vdd.n3050 39.2114
R17647 vdd.n3054 vdd.n3053 39.2114
R17648 vdd.n963 vdd.n919 39.2114
R17649 vdd.n2526 vdd.n920 39.2114
R17650 vdd.n2522 vdd.n921 39.2114
R17651 vdd.n2518 vdd.n922 39.2114
R17652 vdd.n2514 vdd.n923 39.2114
R17653 vdd.n2510 vdd.n924 39.2114
R17654 vdd.n2506 vdd.n925 39.2114
R17655 vdd.n2502 vdd.n926 39.2114
R17656 vdd.n2498 vdd.n927 39.2114
R17657 vdd.n2494 vdd.n928 39.2114
R17658 vdd.n2490 vdd.n929 39.2114
R17659 vdd.n2486 vdd.n930 39.2114
R17660 vdd.n2482 vdd.n931 39.2114
R17661 vdd.n2478 vdd.n932 39.2114
R17662 vdd.n2474 vdd.n933 39.2114
R17663 vdd.n2470 vdd.n934 39.2114
R17664 vdd.n2466 vdd.n935 39.2114
R17665 vdd.n2369 vdd.n1052 39.2114
R17666 vdd.n2368 vdd.n2367 39.2114
R17667 vdd.n2361 vdd.n1054 39.2114
R17668 vdd.n2360 vdd.n2359 39.2114
R17669 vdd.n2353 vdd.n1056 39.2114
R17670 vdd.n2352 vdd.n2351 39.2114
R17671 vdd.n2345 vdd.n1058 39.2114
R17672 vdd.n2344 vdd.n2343 39.2114
R17673 vdd.n1061 vdd.n1060 39.2114
R17674 vdd.n2185 vdd.n2184 39.2114
R17675 vdd.n2190 vdd.n2189 39.2114
R17676 vdd.n2193 vdd.n2192 39.2114
R17677 vdd.n2198 vdd.n2197 39.2114
R17678 vdd.n2201 vdd.n2200 39.2114
R17679 vdd.n2206 vdd.n2205 39.2114
R17680 vdd.n2209 vdd.n2208 39.2114
R17681 vdd.n2215 vdd.n2214 39.2114
R17682 vdd.n2463 vdd.n935 39.2114
R17683 vdd.n2467 vdd.n934 39.2114
R17684 vdd.n2471 vdd.n933 39.2114
R17685 vdd.n2475 vdd.n932 39.2114
R17686 vdd.n2479 vdd.n931 39.2114
R17687 vdd.n2483 vdd.n930 39.2114
R17688 vdd.n2487 vdd.n929 39.2114
R17689 vdd.n2491 vdd.n928 39.2114
R17690 vdd.n2495 vdd.n927 39.2114
R17691 vdd.n2499 vdd.n926 39.2114
R17692 vdd.n2503 vdd.n925 39.2114
R17693 vdd.n2507 vdd.n924 39.2114
R17694 vdd.n2511 vdd.n923 39.2114
R17695 vdd.n2515 vdd.n922 39.2114
R17696 vdd.n2519 vdd.n921 39.2114
R17697 vdd.n2523 vdd.n920 39.2114
R17698 vdd.n2527 vdd.n919 39.2114
R17699 vdd.n2370 vdd.n2369 39.2114
R17700 vdd.n2367 vdd.n2366 39.2114
R17701 vdd.n2362 vdd.n2361 39.2114
R17702 vdd.n2359 vdd.n2358 39.2114
R17703 vdd.n2354 vdd.n2353 39.2114
R17704 vdd.n2351 vdd.n2350 39.2114
R17705 vdd.n2346 vdd.n2345 39.2114
R17706 vdd.n2343 vdd.n2342 39.2114
R17707 vdd.n1062 vdd.n1061 39.2114
R17708 vdd.n2186 vdd.n2185 39.2114
R17709 vdd.n2191 vdd.n2190 39.2114
R17710 vdd.n2192 vdd.n2182 39.2114
R17711 vdd.n2199 vdd.n2198 39.2114
R17712 vdd.n2200 vdd.n2180 39.2114
R17713 vdd.n2207 vdd.n2206 39.2114
R17714 vdd.n2208 vdd.n2176 39.2114
R17715 vdd.n2216 vdd.n2215 39.2114
R17716 vdd.n2335 vdd.n2334 37.2369
R17717 vdd.n2038 vdd.n1971 37.2369
R17718 vdd.n2077 vdd.n1931 37.2369
R17719 vdd.n3138 vdd.n769 37.2369
R17720 vdd.n3186 vdd.n3185 37.2369
R17721 vdd.n690 vdd.n689 37.2369
R17722 vdd.n2377 vdd.n1047 31.6883
R17723 vdd.n2602 vdd.n956 31.6883
R17724 vdd.n2535 vdd.n959 31.6883
R17725 vdd.n2281 vdd.n2278 31.6883
R17726 vdd.n2789 vdd.n2787 31.6883
R17727 vdd.n2994 vdd.n2993 31.6883
R17728 vdd.n2866 vdd.n912 31.6883
R17729 vdd.n3057 vdd.n3056 31.6883
R17730 vdd.n2976 vdd.n2975 31.6883
R17731 vdd.n3062 vdd.n802 31.6883
R17732 vdd.n2708 vdd.n2707 31.6883
R17733 vdd.n2862 vdd.n2861 31.6883
R17734 vdd.n2373 vdd.n2372 31.6883
R17735 vdd.n2530 vdd.n2529 31.6883
R17736 vdd.n2462 vdd.n2461 31.6883
R17737 vdd.n2219 vdd.n2218 31.6883
R17738 vdd.n2212 vdd.n2178 30.449
R17739 vdd.n967 vdd.n966 30.449
R17740 vdd.n2153 vdd.n2152 30.449
R17741 vdd.n2540 vdd.n958 30.449
R17742 vdd.n2644 vdd.n2643 30.449
R17743 vdd.n3000 vdd.n833 30.449
R17744 vdd.n2794 vdd.n2640 30.449
R17745 vdd.n801 vdd.n800 30.449
R17746 vdd.n1418 vdd.n1225 22.2201
R17747 vdd.n2329 vdd.n1073 22.2201
R17748 vdd.n3223 vdd.n723 22.2201
R17749 vdd.n3355 vdd.n3354 22.2201
R17750 vdd.n1429 vdd.n1187 19.3944
R17751 vdd.n1429 vdd.n1185 19.3944
R17752 vdd.n1433 vdd.n1185 19.3944
R17753 vdd.n1433 vdd.n1175 19.3944
R17754 vdd.n1446 vdd.n1175 19.3944
R17755 vdd.n1446 vdd.n1173 19.3944
R17756 vdd.n1450 vdd.n1173 19.3944
R17757 vdd.n1450 vdd.n1165 19.3944
R17758 vdd.n1463 vdd.n1165 19.3944
R17759 vdd.n1463 vdd.n1163 19.3944
R17760 vdd.n1467 vdd.n1163 19.3944
R17761 vdd.n1467 vdd.n1152 19.3944
R17762 vdd.n1479 vdd.n1152 19.3944
R17763 vdd.n1479 vdd.n1150 19.3944
R17764 vdd.n1483 vdd.n1150 19.3944
R17765 vdd.n1483 vdd.n1141 19.3944
R17766 vdd.n1496 vdd.n1141 19.3944
R17767 vdd.n1496 vdd.n1139 19.3944
R17768 vdd.n1500 vdd.n1139 19.3944
R17769 vdd.n1500 vdd.n1130 19.3944
R17770 vdd.n1819 vdd.n1130 19.3944
R17771 vdd.n1819 vdd.n1128 19.3944
R17772 vdd.n1823 vdd.n1128 19.3944
R17773 vdd.n1823 vdd.n1118 19.3944
R17774 vdd.n1836 vdd.n1118 19.3944
R17775 vdd.n1836 vdd.n1116 19.3944
R17776 vdd.n1840 vdd.n1116 19.3944
R17777 vdd.n1840 vdd.n1108 19.3944
R17778 vdd.n1853 vdd.n1108 19.3944
R17779 vdd.n1853 vdd.n1106 19.3944
R17780 vdd.n1857 vdd.n1106 19.3944
R17781 vdd.n1857 vdd.n1095 19.3944
R17782 vdd.n1869 vdd.n1095 19.3944
R17783 vdd.n1869 vdd.n1093 19.3944
R17784 vdd.n1873 vdd.n1093 19.3944
R17785 vdd.n1873 vdd.n1085 19.3944
R17786 vdd.n1886 vdd.n1085 19.3944
R17787 vdd.n1886 vdd.n1082 19.3944
R17788 vdd.n1892 vdd.n1082 19.3944
R17789 vdd.n1892 vdd.n1083 19.3944
R17790 vdd.n1083 vdd.n1072 19.3944
R17791 vdd.n1353 vdd.n1288 19.3944
R17792 vdd.n1349 vdd.n1288 19.3944
R17793 vdd.n1349 vdd.n1348 19.3944
R17794 vdd.n1348 vdd.n1347 19.3944
R17795 vdd.n1347 vdd.n1294 19.3944
R17796 vdd.n1343 vdd.n1294 19.3944
R17797 vdd.n1343 vdd.n1342 19.3944
R17798 vdd.n1342 vdd.n1341 19.3944
R17799 vdd.n1341 vdd.n1300 19.3944
R17800 vdd.n1337 vdd.n1300 19.3944
R17801 vdd.n1337 vdd.n1336 19.3944
R17802 vdd.n1336 vdd.n1335 19.3944
R17803 vdd.n1335 vdd.n1306 19.3944
R17804 vdd.n1331 vdd.n1306 19.3944
R17805 vdd.n1331 vdd.n1330 19.3944
R17806 vdd.n1330 vdd.n1329 19.3944
R17807 vdd.n1329 vdd.n1312 19.3944
R17808 vdd.n1325 vdd.n1312 19.3944
R17809 vdd.n1325 vdd.n1324 19.3944
R17810 vdd.n1324 vdd.n1323 19.3944
R17811 vdd.n1388 vdd.n1387 19.3944
R17812 vdd.n1387 vdd.n1386 19.3944
R17813 vdd.n1386 vdd.n1259 19.3944
R17814 vdd.n1382 vdd.n1259 19.3944
R17815 vdd.n1382 vdd.n1381 19.3944
R17816 vdd.n1381 vdd.n1380 19.3944
R17817 vdd.n1380 vdd.n1265 19.3944
R17818 vdd.n1376 vdd.n1265 19.3944
R17819 vdd.n1376 vdd.n1375 19.3944
R17820 vdd.n1375 vdd.n1374 19.3944
R17821 vdd.n1374 vdd.n1271 19.3944
R17822 vdd.n1370 vdd.n1271 19.3944
R17823 vdd.n1370 vdd.n1369 19.3944
R17824 vdd.n1369 vdd.n1368 19.3944
R17825 vdd.n1368 vdd.n1277 19.3944
R17826 vdd.n1364 vdd.n1277 19.3944
R17827 vdd.n1364 vdd.n1363 19.3944
R17828 vdd.n1363 vdd.n1362 19.3944
R17829 vdd.n1362 vdd.n1283 19.3944
R17830 vdd.n1358 vdd.n1283 19.3944
R17831 vdd.n1421 vdd.n1192 19.3944
R17832 vdd.n1416 vdd.n1192 19.3944
R17833 vdd.n1416 vdd.n1227 19.3944
R17834 vdd.n1412 vdd.n1227 19.3944
R17835 vdd.n1412 vdd.n1411 19.3944
R17836 vdd.n1411 vdd.n1410 19.3944
R17837 vdd.n1410 vdd.n1233 19.3944
R17838 vdd.n1406 vdd.n1233 19.3944
R17839 vdd.n1406 vdd.n1405 19.3944
R17840 vdd.n1405 vdd.n1404 19.3944
R17841 vdd.n1404 vdd.n1239 19.3944
R17842 vdd.n1400 vdd.n1239 19.3944
R17843 vdd.n1400 vdd.n1399 19.3944
R17844 vdd.n1399 vdd.n1398 19.3944
R17845 vdd.n1398 vdd.n1245 19.3944
R17846 vdd.n1394 vdd.n1245 19.3944
R17847 vdd.n1394 vdd.n1393 19.3944
R17848 vdd.n1393 vdd.n1392 19.3944
R17849 vdd.n2034 vdd.n1969 19.3944
R17850 vdd.n2034 vdd.n1975 19.3944
R17851 vdd.n2029 vdd.n1975 19.3944
R17852 vdd.n2029 vdd.n2028 19.3944
R17853 vdd.n2028 vdd.n2027 19.3944
R17854 vdd.n2027 vdd.n1982 19.3944
R17855 vdd.n2022 vdd.n1982 19.3944
R17856 vdd.n2022 vdd.n2021 19.3944
R17857 vdd.n2021 vdd.n2020 19.3944
R17858 vdd.n2020 vdd.n1989 19.3944
R17859 vdd.n2015 vdd.n1989 19.3944
R17860 vdd.n2015 vdd.n2014 19.3944
R17861 vdd.n2014 vdd.n2013 19.3944
R17862 vdd.n2013 vdd.n1997 19.3944
R17863 vdd.n2008 vdd.n1997 19.3944
R17864 vdd.n2008 vdd.n2007 19.3944
R17865 vdd.n2003 vdd.n2002 19.3944
R17866 vdd.n2336 vdd.n1068 19.3944
R17867 vdd.n2073 vdd.n1929 19.3944
R17868 vdd.n2073 vdd.n1935 19.3944
R17869 vdd.n2068 vdd.n1935 19.3944
R17870 vdd.n2068 vdd.n2067 19.3944
R17871 vdd.n2067 vdd.n2066 19.3944
R17872 vdd.n2066 vdd.n1942 19.3944
R17873 vdd.n2061 vdd.n1942 19.3944
R17874 vdd.n2061 vdd.n2060 19.3944
R17875 vdd.n2060 vdd.n2059 19.3944
R17876 vdd.n2059 vdd.n1949 19.3944
R17877 vdd.n2054 vdd.n1949 19.3944
R17878 vdd.n2054 vdd.n2053 19.3944
R17879 vdd.n2053 vdd.n2052 19.3944
R17880 vdd.n2052 vdd.n1956 19.3944
R17881 vdd.n2047 vdd.n1956 19.3944
R17882 vdd.n2047 vdd.n2046 19.3944
R17883 vdd.n2046 vdd.n2045 19.3944
R17884 vdd.n2045 vdd.n1963 19.3944
R17885 vdd.n2040 vdd.n1963 19.3944
R17886 vdd.n2040 vdd.n2039 19.3944
R17887 vdd.n2324 vdd.n2323 19.3944
R17888 vdd.n2323 vdd.n1901 19.3944
R17889 vdd.n2318 vdd.n2317 19.3944
R17890 vdd.n2100 vdd.n1905 19.3944
R17891 vdd.n2100 vdd.n1907 19.3944
R17892 vdd.n1910 vdd.n1907 19.3944
R17893 vdd.n2093 vdd.n1910 19.3944
R17894 vdd.n2093 vdd.n2092 19.3944
R17895 vdd.n2092 vdd.n2091 19.3944
R17896 vdd.n2091 vdd.n1916 19.3944
R17897 vdd.n2086 vdd.n1916 19.3944
R17898 vdd.n2086 vdd.n2085 19.3944
R17899 vdd.n2085 vdd.n2084 19.3944
R17900 vdd.n2084 vdd.n1923 19.3944
R17901 vdd.n2079 vdd.n1923 19.3944
R17902 vdd.n2079 vdd.n2078 19.3944
R17903 vdd.n1425 vdd.n1190 19.3944
R17904 vdd.n1425 vdd.n1181 19.3944
R17905 vdd.n1438 vdd.n1181 19.3944
R17906 vdd.n1438 vdd.n1179 19.3944
R17907 vdd.n1442 vdd.n1179 19.3944
R17908 vdd.n1442 vdd.n1170 19.3944
R17909 vdd.n1455 vdd.n1170 19.3944
R17910 vdd.n1455 vdd.n1168 19.3944
R17911 vdd.n1459 vdd.n1168 19.3944
R17912 vdd.n1459 vdd.n1159 19.3944
R17913 vdd.n1471 vdd.n1159 19.3944
R17914 vdd.n1471 vdd.n1157 19.3944
R17915 vdd.n1475 vdd.n1157 19.3944
R17916 vdd.n1475 vdd.n1147 19.3944
R17917 vdd.n1488 vdd.n1147 19.3944
R17918 vdd.n1488 vdd.n1145 19.3944
R17919 vdd.n1492 vdd.n1145 19.3944
R17920 vdd.n1492 vdd.n1136 19.3944
R17921 vdd.n1504 vdd.n1136 19.3944
R17922 vdd.n1504 vdd.n1134 19.3944
R17923 vdd.n1815 vdd.n1134 19.3944
R17924 vdd.n1815 vdd.n1124 19.3944
R17925 vdd.n1828 vdd.n1124 19.3944
R17926 vdd.n1828 vdd.n1122 19.3944
R17927 vdd.n1832 vdd.n1122 19.3944
R17928 vdd.n1832 vdd.n1113 19.3944
R17929 vdd.n1845 vdd.n1113 19.3944
R17930 vdd.n1845 vdd.n1111 19.3944
R17931 vdd.n1849 vdd.n1111 19.3944
R17932 vdd.n1849 vdd.n1102 19.3944
R17933 vdd.n1861 vdd.n1102 19.3944
R17934 vdd.n1861 vdd.n1100 19.3944
R17935 vdd.n1865 vdd.n1100 19.3944
R17936 vdd.n1865 vdd.n1090 19.3944
R17937 vdd.n1878 vdd.n1090 19.3944
R17938 vdd.n1878 vdd.n1088 19.3944
R17939 vdd.n1882 vdd.n1088 19.3944
R17940 vdd.n1882 vdd.n1078 19.3944
R17941 vdd.n1897 vdd.n1078 19.3944
R17942 vdd.n1897 vdd.n1076 19.3944
R17943 vdd.n2327 vdd.n1076 19.3944
R17944 vdd.n3229 vdd.n686 19.3944
R17945 vdd.n3229 vdd.n676 19.3944
R17946 vdd.n3241 vdd.n676 19.3944
R17947 vdd.n3241 vdd.n674 19.3944
R17948 vdd.n3245 vdd.n674 19.3944
R17949 vdd.n3245 vdd.n666 19.3944
R17950 vdd.n3258 vdd.n666 19.3944
R17951 vdd.n3258 vdd.n664 19.3944
R17952 vdd.n3262 vdd.n664 19.3944
R17953 vdd.n3262 vdd.n653 19.3944
R17954 vdd.n3274 vdd.n653 19.3944
R17955 vdd.n3274 vdd.n651 19.3944
R17956 vdd.n3278 vdd.n651 19.3944
R17957 vdd.n3278 vdd.n642 19.3944
R17958 vdd.n3291 vdd.n642 19.3944
R17959 vdd.n3291 vdd.n640 19.3944
R17960 vdd.n3298 vdd.n640 19.3944
R17961 vdd.n3298 vdd.n3297 19.3944
R17962 vdd.n3297 vdd.n631 19.3944
R17963 vdd.n3311 vdd.n631 19.3944
R17964 vdd.n3312 vdd.n3311 19.3944
R17965 vdd.n3312 vdd.n629 19.3944
R17966 vdd.n3316 vdd.n629 19.3944
R17967 vdd.n3318 vdd.n3316 19.3944
R17968 vdd.n3319 vdd.n3318 19.3944
R17969 vdd.n3319 vdd.n627 19.3944
R17970 vdd.n3323 vdd.n627 19.3944
R17971 vdd.n3325 vdd.n3323 19.3944
R17972 vdd.n3326 vdd.n3325 19.3944
R17973 vdd.n3326 vdd.n625 19.3944
R17974 vdd.n3330 vdd.n625 19.3944
R17975 vdd.n3333 vdd.n3330 19.3944
R17976 vdd.n3334 vdd.n3333 19.3944
R17977 vdd.n3334 vdd.n623 19.3944
R17978 vdd.n3338 vdd.n623 19.3944
R17979 vdd.n3340 vdd.n3338 19.3944
R17980 vdd.n3341 vdd.n3340 19.3944
R17981 vdd.n3341 vdd.n621 19.3944
R17982 vdd.n3345 vdd.n621 19.3944
R17983 vdd.n3347 vdd.n3345 19.3944
R17984 vdd.n3348 vdd.n3347 19.3944
R17985 vdd.n569 vdd.n438 19.3944
R17986 vdd.n575 vdd.n438 19.3944
R17987 vdd.n576 vdd.n575 19.3944
R17988 vdd.n579 vdd.n576 19.3944
R17989 vdd.n579 vdd.n436 19.3944
R17990 vdd.n585 vdd.n436 19.3944
R17991 vdd.n586 vdd.n585 19.3944
R17992 vdd.n589 vdd.n586 19.3944
R17993 vdd.n589 vdd.n434 19.3944
R17994 vdd.n595 vdd.n434 19.3944
R17995 vdd.n596 vdd.n595 19.3944
R17996 vdd.n599 vdd.n596 19.3944
R17997 vdd.n599 vdd.n432 19.3944
R17998 vdd.n605 vdd.n432 19.3944
R17999 vdd.n606 vdd.n605 19.3944
R18000 vdd.n609 vdd.n606 19.3944
R18001 vdd.n609 vdd.n430 19.3944
R18002 vdd.n615 vdd.n430 19.3944
R18003 vdd.n617 vdd.n615 19.3944
R18004 vdd.n618 vdd.n617 19.3944
R18005 vdd.n516 vdd.n515 19.3944
R18006 vdd.n519 vdd.n516 19.3944
R18007 vdd.n519 vdd.n450 19.3944
R18008 vdd.n525 vdd.n450 19.3944
R18009 vdd.n526 vdd.n525 19.3944
R18010 vdd.n529 vdd.n526 19.3944
R18011 vdd.n529 vdd.n448 19.3944
R18012 vdd.n535 vdd.n448 19.3944
R18013 vdd.n536 vdd.n535 19.3944
R18014 vdd.n539 vdd.n536 19.3944
R18015 vdd.n539 vdd.n446 19.3944
R18016 vdd.n545 vdd.n446 19.3944
R18017 vdd.n546 vdd.n545 19.3944
R18018 vdd.n549 vdd.n546 19.3944
R18019 vdd.n549 vdd.n444 19.3944
R18020 vdd.n555 vdd.n444 19.3944
R18021 vdd.n556 vdd.n555 19.3944
R18022 vdd.n559 vdd.n556 19.3944
R18023 vdd.n559 vdd.n442 19.3944
R18024 vdd.n565 vdd.n442 19.3944
R18025 vdd.n466 vdd.n465 19.3944
R18026 vdd.n469 vdd.n466 19.3944
R18027 vdd.n469 vdd.n462 19.3944
R18028 vdd.n475 vdd.n462 19.3944
R18029 vdd.n476 vdd.n475 19.3944
R18030 vdd.n479 vdd.n476 19.3944
R18031 vdd.n479 vdd.n460 19.3944
R18032 vdd.n485 vdd.n460 19.3944
R18033 vdd.n486 vdd.n485 19.3944
R18034 vdd.n489 vdd.n486 19.3944
R18035 vdd.n489 vdd.n458 19.3944
R18036 vdd.n495 vdd.n458 19.3944
R18037 vdd.n496 vdd.n495 19.3944
R18038 vdd.n499 vdd.n496 19.3944
R18039 vdd.n499 vdd.n456 19.3944
R18040 vdd.n505 vdd.n456 19.3944
R18041 vdd.n506 vdd.n505 19.3944
R18042 vdd.n509 vdd.n506 19.3944
R18043 vdd.n3233 vdd.n683 19.3944
R18044 vdd.n3233 vdd.n681 19.3944
R18045 vdd.n3237 vdd.n681 19.3944
R18046 vdd.n3237 vdd.n671 19.3944
R18047 vdd.n3250 vdd.n671 19.3944
R18048 vdd.n3250 vdd.n669 19.3944
R18049 vdd.n3254 vdd.n669 19.3944
R18050 vdd.n3254 vdd.n660 19.3944
R18051 vdd.n3266 vdd.n660 19.3944
R18052 vdd.n3266 vdd.n658 19.3944
R18053 vdd.n3270 vdd.n658 19.3944
R18054 vdd.n3270 vdd.n648 19.3944
R18055 vdd.n3283 vdd.n648 19.3944
R18056 vdd.n3283 vdd.n646 19.3944
R18057 vdd.n3287 vdd.n646 19.3944
R18058 vdd.n3287 vdd.n637 19.3944
R18059 vdd.n3302 vdd.n637 19.3944
R18060 vdd.n3302 vdd.n635 19.3944
R18061 vdd.n3306 vdd.n635 19.3944
R18062 vdd.n3306 vdd.n336 19.3944
R18063 vdd.n3397 vdd.n336 19.3944
R18064 vdd.n3397 vdd.n337 19.3944
R18065 vdd.n3391 vdd.n337 19.3944
R18066 vdd.n3391 vdd.n3390 19.3944
R18067 vdd.n3390 vdd.n3389 19.3944
R18068 vdd.n3389 vdd.n349 19.3944
R18069 vdd.n3383 vdd.n349 19.3944
R18070 vdd.n3383 vdd.n3382 19.3944
R18071 vdd.n3382 vdd.n3381 19.3944
R18072 vdd.n3381 vdd.n359 19.3944
R18073 vdd.n3375 vdd.n359 19.3944
R18074 vdd.n3375 vdd.n3374 19.3944
R18075 vdd.n3374 vdd.n3373 19.3944
R18076 vdd.n3373 vdd.n370 19.3944
R18077 vdd.n3367 vdd.n370 19.3944
R18078 vdd.n3367 vdd.n3366 19.3944
R18079 vdd.n3366 vdd.n3365 19.3944
R18080 vdd.n3365 vdd.n381 19.3944
R18081 vdd.n3359 vdd.n381 19.3944
R18082 vdd.n3359 vdd.n3358 19.3944
R18083 vdd.n3358 vdd.n3357 19.3944
R18084 vdd.n3180 vdd.n747 19.3944
R18085 vdd.n3180 vdd.n3177 19.3944
R18086 vdd.n3177 vdd.n3174 19.3944
R18087 vdd.n3174 vdd.n3173 19.3944
R18088 vdd.n3173 vdd.n3170 19.3944
R18089 vdd.n3170 vdd.n3169 19.3944
R18090 vdd.n3169 vdd.n3166 19.3944
R18091 vdd.n3166 vdd.n3165 19.3944
R18092 vdd.n3165 vdd.n3162 19.3944
R18093 vdd.n3162 vdd.n3161 19.3944
R18094 vdd.n3161 vdd.n3158 19.3944
R18095 vdd.n3158 vdd.n3157 19.3944
R18096 vdd.n3157 vdd.n3154 19.3944
R18097 vdd.n3154 vdd.n3153 19.3944
R18098 vdd.n3153 vdd.n3150 19.3944
R18099 vdd.n3150 vdd.n3149 19.3944
R18100 vdd.n3149 vdd.n3146 19.3944
R18101 vdd.n3146 vdd.n3145 19.3944
R18102 vdd.n3145 vdd.n3142 19.3944
R18103 vdd.n3142 vdd.n3141 19.3944
R18104 vdd.n3220 vdd.n3219 19.3944
R18105 vdd.n3219 vdd.n3218 19.3944
R18106 vdd.n732 vdd.n729 19.3944
R18107 vdd.n3214 vdd.n3213 19.3944
R18108 vdd.n3213 vdd.n3210 19.3944
R18109 vdd.n3210 vdd.n3209 19.3944
R18110 vdd.n3209 vdd.n3206 19.3944
R18111 vdd.n3206 vdd.n3205 19.3944
R18112 vdd.n3205 vdd.n3202 19.3944
R18113 vdd.n3202 vdd.n3201 19.3944
R18114 vdd.n3201 vdd.n3198 19.3944
R18115 vdd.n3198 vdd.n3197 19.3944
R18116 vdd.n3197 vdd.n3194 19.3944
R18117 vdd.n3194 vdd.n3193 19.3944
R18118 vdd.n3193 vdd.n3190 19.3944
R18119 vdd.n3190 vdd.n3189 19.3944
R18120 vdd.n3134 vdd.n767 19.3944
R18121 vdd.n3134 vdd.n3131 19.3944
R18122 vdd.n3131 vdd.n3128 19.3944
R18123 vdd.n3128 vdd.n3127 19.3944
R18124 vdd.n3127 vdd.n3124 19.3944
R18125 vdd.n3124 vdd.n3123 19.3944
R18126 vdd.n3123 vdd.n3120 19.3944
R18127 vdd.n3120 vdd.n3119 19.3944
R18128 vdd.n3119 vdd.n3116 19.3944
R18129 vdd.n3116 vdd.n3115 19.3944
R18130 vdd.n3115 vdd.n3112 19.3944
R18131 vdd.n3112 vdd.n3111 19.3944
R18132 vdd.n3111 vdd.n3108 19.3944
R18133 vdd.n3108 vdd.n3107 19.3944
R18134 vdd.n3107 vdd.n3104 19.3944
R18135 vdd.n3104 vdd.n3103 19.3944
R18136 vdd.n3100 vdd.n3099 19.3944
R18137 vdd.n3096 vdd.n3095 19.3944
R18138 vdd.n1357 vdd.n1353 19.0066
R18139 vdd.n2038 vdd.n1969 19.0066
R18140 vdd.n569 vdd.n566 19.0066
R18141 vdd.n3138 vdd.n767 19.0066
R18142 vdd.n2178 vdd.n2177 16.0975
R18143 vdd.n966 vdd.n965 16.0975
R18144 vdd.n1318 vdd.n1317 16.0975
R18145 vdd.n1356 vdd.n1355 16.0975
R18146 vdd.n1252 vdd.n1251 16.0975
R18147 vdd.n2334 vdd.n2333 16.0975
R18148 vdd.n1971 vdd.n1970 16.0975
R18149 vdd.n1931 vdd.n1930 16.0975
R18150 vdd.n2152 vdd.n2151 16.0975
R18151 vdd.n958 vdd.n957 16.0975
R18152 vdd.n2643 vdd.n2642 16.0975
R18153 vdd.n427 vdd.n426 16.0975
R18154 vdd.n441 vdd.n440 16.0975
R18155 vdd.n453 vdd.n452 16.0975
R18156 vdd.n769 vdd.n768 16.0975
R18157 vdd.n3185 vdd.n3184 16.0975
R18158 vdd.n833 vdd.n832 16.0975
R18159 vdd.n2640 vdd.n2639 16.0975
R18160 vdd.n689 vdd.n688 16.0975
R18161 vdd.n800 vdd.n799 16.0975
R18162 vdd.t196 vdd.n2604 15.4182
R18163 vdd.n2857 vdd.t294 15.4182
R18164 vdd.n28 vdd.n27 14.5458
R18165 vdd.n2375 vdd.n1049 14.5112
R18166 vdd.n3059 vdd.n692 14.5112
R18167 vdd.n328 vdd.n293 13.1884
R18168 vdd.n269 vdd.n234 13.1884
R18169 vdd.n226 vdd.n191 13.1884
R18170 vdd.n167 vdd.n132 13.1884
R18171 vdd.n125 vdd.n90 13.1884
R18172 vdd.n66 vdd.n31 13.1884
R18173 vdd.n1747 vdd.n1712 13.1884
R18174 vdd.n1806 vdd.n1771 13.1884
R18175 vdd.n1645 vdd.n1610 13.1884
R18176 vdd.n1704 vdd.n1669 13.1884
R18177 vdd.n1544 vdd.n1509 13.1884
R18178 vdd.n1603 vdd.n1568 13.1884
R18179 vdd.n1388 vdd.n1253 12.9944
R18180 vdd.n1392 vdd.n1253 12.9944
R18181 vdd.n2077 vdd.n1929 12.9944
R18182 vdd.n2078 vdd.n2077 12.9944
R18183 vdd.n515 vdd.n454 12.9944
R18184 vdd.n509 vdd.n454 12.9944
R18185 vdd.n3186 vdd.n747 12.9944
R18186 vdd.n3189 vdd.n3186 12.9944
R18187 vdd.n329 vdd.n291 12.8005
R18188 vdd.n324 vdd.n295 12.8005
R18189 vdd.n270 vdd.n232 12.8005
R18190 vdd.n265 vdd.n236 12.8005
R18191 vdd.n227 vdd.n189 12.8005
R18192 vdd.n222 vdd.n193 12.8005
R18193 vdd.n168 vdd.n130 12.8005
R18194 vdd.n163 vdd.n134 12.8005
R18195 vdd.n126 vdd.n88 12.8005
R18196 vdd.n121 vdd.n92 12.8005
R18197 vdd.n67 vdd.n29 12.8005
R18198 vdd.n62 vdd.n33 12.8005
R18199 vdd.n1748 vdd.n1710 12.8005
R18200 vdd.n1743 vdd.n1714 12.8005
R18201 vdd.n1807 vdd.n1769 12.8005
R18202 vdd.n1802 vdd.n1773 12.8005
R18203 vdd.n1646 vdd.n1608 12.8005
R18204 vdd.n1641 vdd.n1612 12.8005
R18205 vdd.n1705 vdd.n1667 12.8005
R18206 vdd.n1700 vdd.n1671 12.8005
R18207 vdd.n1545 vdd.n1507 12.8005
R18208 vdd.n1540 vdd.n1511 12.8005
R18209 vdd.n1604 vdd.n1566 12.8005
R18210 vdd.n1599 vdd.n1570 12.8005
R18211 vdd.n323 vdd.n296 12.0247
R18212 vdd.n264 vdd.n237 12.0247
R18213 vdd.n221 vdd.n194 12.0247
R18214 vdd.n162 vdd.n135 12.0247
R18215 vdd.n120 vdd.n93 12.0247
R18216 vdd.n61 vdd.n34 12.0247
R18217 vdd.n1742 vdd.n1715 12.0247
R18218 vdd.n1801 vdd.n1774 12.0247
R18219 vdd.n1640 vdd.n1613 12.0247
R18220 vdd.n1699 vdd.n1672 12.0247
R18221 vdd.n1539 vdd.n1512 12.0247
R18222 vdd.n1598 vdd.n1571 12.0247
R18223 vdd.n1427 vdd.n1183 11.337
R18224 vdd.n1436 vdd.n1183 11.337
R18225 vdd.n1436 vdd.n1435 11.337
R18226 vdd.n1444 vdd.n1177 11.337
R18227 vdd.n1453 vdd.n1452 11.337
R18228 vdd.n1469 vdd.n1161 11.337
R18229 vdd.n1477 vdd.n1154 11.337
R18230 vdd.n1486 vdd.n1485 11.337
R18231 vdd.n1494 vdd.n1143 11.337
R18232 vdd.n1817 vdd.n1132 11.337
R18233 vdd.n1826 vdd.n1126 11.337
R18234 vdd.n1834 vdd.n1120 11.337
R18235 vdd.n1843 vdd.n1842 11.337
R18236 vdd.n1859 vdd.n1104 11.337
R18237 vdd.n1867 vdd.n1097 11.337
R18238 vdd.n1876 vdd.n1875 11.337
R18239 vdd.n1884 vdd.n1080 11.337
R18240 vdd.n1895 vdd.n1080 11.337
R18241 vdd.n1895 vdd.n1894 11.337
R18242 vdd.n3231 vdd.n678 11.337
R18243 vdd.n3239 vdd.n678 11.337
R18244 vdd.n3239 vdd.n679 11.337
R18245 vdd.n3248 vdd.n3247 11.337
R18246 vdd.n3264 vdd.n662 11.337
R18247 vdd.n3272 vdd.n655 11.337
R18248 vdd.n3281 vdd.n3280 11.337
R18249 vdd.n3289 vdd.n644 11.337
R18250 vdd.n3308 vdd.n633 11.337
R18251 vdd.n3395 vdd.n340 11.337
R18252 vdd.n3393 vdd.n344 11.337
R18253 vdd.n3387 vdd.n3386 11.337
R18254 vdd.n3379 vdd.n361 11.337
R18255 vdd.n3378 vdd.n3377 11.337
R18256 vdd.n3371 vdd.n3370 11.337
R18257 vdd.n3369 vdd.n375 11.337
R18258 vdd.n3363 vdd.n3362 11.337
R18259 vdd.n3362 vdd.n3361 11.337
R18260 vdd.n3361 vdd.n386 11.337
R18261 vdd.n320 vdd.n319 11.249
R18262 vdd.n261 vdd.n260 11.249
R18263 vdd.n218 vdd.n217 11.249
R18264 vdd.n159 vdd.n158 11.249
R18265 vdd.n117 vdd.n116 11.249
R18266 vdd.n58 vdd.n57 11.249
R18267 vdd.n1739 vdd.n1738 11.249
R18268 vdd.n1798 vdd.n1797 11.249
R18269 vdd.n1637 vdd.n1636 11.249
R18270 vdd.n1696 vdd.n1695 11.249
R18271 vdd.n1536 vdd.n1535 11.249
R18272 vdd.n1595 vdd.n1594 11.249
R18273 vdd.n1225 vdd.t231 11.2237
R18274 vdd.n3355 vdd.t238 11.2237
R18275 vdd.n2532 vdd.t204 11.1103
R18276 vdd.n2864 vdd.t193 11.1103
R18277 vdd.t35 vdd.n1098 10.7702
R18278 vdd.n3256 vdd.t97 10.7702
R18279 vdd.n305 vdd.n304 10.7238
R18280 vdd.n246 vdd.n245 10.7238
R18281 vdd.n203 vdd.n202 10.7238
R18282 vdd.n144 vdd.n143 10.7238
R18283 vdd.n102 vdd.n101 10.7238
R18284 vdd.n43 vdd.n42 10.7238
R18285 vdd.n1724 vdd.n1723 10.7238
R18286 vdd.n1783 vdd.n1782 10.7238
R18287 vdd.n1622 vdd.n1621 10.7238
R18288 vdd.n1681 vdd.n1680 10.7238
R18289 vdd.n1521 vdd.n1520 10.7238
R18290 vdd.n1580 vdd.n1579 10.7238
R18291 vdd.n2378 vdd.n2377 10.6151
R18292 vdd.n2379 vdd.n2378 10.6151
R18293 vdd.n2379 vdd.n1035 10.6151
R18294 vdd.n2389 vdd.n1035 10.6151
R18295 vdd.n2390 vdd.n2389 10.6151
R18296 vdd.n2391 vdd.n2390 10.6151
R18297 vdd.n2391 vdd.n1022 10.6151
R18298 vdd.n2402 vdd.n1022 10.6151
R18299 vdd.n2403 vdd.n2402 10.6151
R18300 vdd.n2404 vdd.n2403 10.6151
R18301 vdd.n2404 vdd.n1010 10.6151
R18302 vdd.n2414 vdd.n1010 10.6151
R18303 vdd.n2415 vdd.n2414 10.6151
R18304 vdd.n2416 vdd.n2415 10.6151
R18305 vdd.n2416 vdd.n998 10.6151
R18306 vdd.n2426 vdd.n998 10.6151
R18307 vdd.n2427 vdd.n2426 10.6151
R18308 vdd.n2428 vdd.n2427 10.6151
R18309 vdd.n2428 vdd.n987 10.6151
R18310 vdd.n2438 vdd.n987 10.6151
R18311 vdd.n2439 vdd.n2438 10.6151
R18312 vdd.n2440 vdd.n2439 10.6151
R18313 vdd.n2440 vdd.n974 10.6151
R18314 vdd.n2452 vdd.n974 10.6151
R18315 vdd.n2453 vdd.n2452 10.6151
R18316 vdd.n2455 vdd.n2453 10.6151
R18317 vdd.n2455 vdd.n2454 10.6151
R18318 vdd.n2454 vdd.n956 10.6151
R18319 vdd.n2602 vdd.n2601 10.6151
R18320 vdd.n2601 vdd.n2600 10.6151
R18321 vdd.n2600 vdd.n2597 10.6151
R18322 vdd.n2597 vdd.n2596 10.6151
R18323 vdd.n2596 vdd.n2593 10.6151
R18324 vdd.n2593 vdd.n2592 10.6151
R18325 vdd.n2592 vdd.n2589 10.6151
R18326 vdd.n2589 vdd.n2588 10.6151
R18327 vdd.n2588 vdd.n2585 10.6151
R18328 vdd.n2585 vdd.n2584 10.6151
R18329 vdd.n2584 vdd.n2581 10.6151
R18330 vdd.n2581 vdd.n2580 10.6151
R18331 vdd.n2580 vdd.n2577 10.6151
R18332 vdd.n2577 vdd.n2576 10.6151
R18333 vdd.n2576 vdd.n2573 10.6151
R18334 vdd.n2573 vdd.n2572 10.6151
R18335 vdd.n2572 vdd.n2569 10.6151
R18336 vdd.n2569 vdd.n2568 10.6151
R18337 vdd.n2568 vdd.n2565 10.6151
R18338 vdd.n2565 vdd.n2564 10.6151
R18339 vdd.n2564 vdd.n2561 10.6151
R18340 vdd.n2561 vdd.n2560 10.6151
R18341 vdd.n2560 vdd.n2557 10.6151
R18342 vdd.n2557 vdd.n2556 10.6151
R18343 vdd.n2556 vdd.n2553 10.6151
R18344 vdd.n2553 vdd.n2552 10.6151
R18345 vdd.n2552 vdd.n2549 10.6151
R18346 vdd.n2549 vdd.n2548 10.6151
R18347 vdd.n2548 vdd.n2545 10.6151
R18348 vdd.n2545 vdd.n2544 10.6151
R18349 vdd.n2544 vdd.n2541 10.6151
R18350 vdd.n2539 vdd.n2536 10.6151
R18351 vdd.n2536 vdd.n2535 10.6151
R18352 vdd.n2278 vdd.n2277 10.6151
R18353 vdd.n2277 vdd.n2275 10.6151
R18354 vdd.n2275 vdd.n2274 10.6151
R18355 vdd.n2274 vdd.n2272 10.6151
R18356 vdd.n2272 vdd.n2271 10.6151
R18357 vdd.n2271 vdd.n2269 10.6151
R18358 vdd.n2269 vdd.n2268 10.6151
R18359 vdd.n2268 vdd.n2266 10.6151
R18360 vdd.n2266 vdd.n2265 10.6151
R18361 vdd.n2265 vdd.n2263 10.6151
R18362 vdd.n2263 vdd.n2262 10.6151
R18363 vdd.n2262 vdd.n2260 10.6151
R18364 vdd.n2260 vdd.n2259 10.6151
R18365 vdd.n2259 vdd.n2174 10.6151
R18366 vdd.n2174 vdd.n2173 10.6151
R18367 vdd.n2173 vdd.n2171 10.6151
R18368 vdd.n2171 vdd.n2170 10.6151
R18369 vdd.n2170 vdd.n2168 10.6151
R18370 vdd.n2168 vdd.n2167 10.6151
R18371 vdd.n2167 vdd.n2165 10.6151
R18372 vdd.n2165 vdd.n2164 10.6151
R18373 vdd.n2164 vdd.n2162 10.6151
R18374 vdd.n2162 vdd.n2161 10.6151
R18375 vdd.n2161 vdd.n2159 10.6151
R18376 vdd.n2159 vdd.n2158 10.6151
R18377 vdd.n2158 vdd.n2155 10.6151
R18378 vdd.n2155 vdd.n2154 10.6151
R18379 vdd.n2154 vdd.n959 10.6151
R18380 vdd.n2112 vdd.n1047 10.6151
R18381 vdd.n2113 vdd.n2112 10.6151
R18382 vdd.n2114 vdd.n2113 10.6151
R18383 vdd.n2114 vdd.n2108 10.6151
R18384 vdd.n2120 vdd.n2108 10.6151
R18385 vdd.n2121 vdd.n2120 10.6151
R18386 vdd.n2122 vdd.n2121 10.6151
R18387 vdd.n2122 vdd.n2106 10.6151
R18388 vdd.n2128 vdd.n2106 10.6151
R18389 vdd.n2129 vdd.n2128 10.6151
R18390 vdd.n2130 vdd.n2129 10.6151
R18391 vdd.n2130 vdd.n2104 10.6151
R18392 vdd.n2136 vdd.n2104 10.6151
R18393 vdd.n2137 vdd.n2136 10.6151
R18394 vdd.n2138 vdd.n2137 10.6151
R18395 vdd.n2138 vdd.n2102 10.6151
R18396 vdd.n2314 vdd.n2102 10.6151
R18397 vdd.n2314 vdd.n2313 10.6151
R18398 vdd.n2313 vdd.n2143 10.6151
R18399 vdd.n2307 vdd.n2143 10.6151
R18400 vdd.n2307 vdd.n2306 10.6151
R18401 vdd.n2306 vdd.n2305 10.6151
R18402 vdd.n2305 vdd.n2145 10.6151
R18403 vdd.n2299 vdd.n2145 10.6151
R18404 vdd.n2299 vdd.n2298 10.6151
R18405 vdd.n2298 vdd.n2297 10.6151
R18406 vdd.n2297 vdd.n2147 10.6151
R18407 vdd.n2291 vdd.n2147 10.6151
R18408 vdd.n2291 vdd.n2290 10.6151
R18409 vdd.n2290 vdd.n2289 10.6151
R18410 vdd.n2289 vdd.n2149 10.6151
R18411 vdd.n2283 vdd.n2282 10.6151
R18412 vdd.n2282 vdd.n2281 10.6151
R18413 vdd.n2787 vdd.n2786 10.6151
R18414 vdd.n2786 vdd.n2784 10.6151
R18415 vdd.n2784 vdd.n2783 10.6151
R18416 vdd.n2783 vdd.n2641 10.6151
R18417 vdd.n2730 vdd.n2641 10.6151
R18418 vdd.n2731 vdd.n2730 10.6151
R18419 vdd.n2733 vdd.n2731 10.6151
R18420 vdd.n2734 vdd.n2733 10.6151
R18421 vdd.n2736 vdd.n2734 10.6151
R18422 vdd.n2737 vdd.n2736 10.6151
R18423 vdd.n2739 vdd.n2737 10.6151
R18424 vdd.n2740 vdd.n2739 10.6151
R18425 vdd.n2742 vdd.n2740 10.6151
R18426 vdd.n2743 vdd.n2742 10.6151
R18427 vdd.n2758 vdd.n2743 10.6151
R18428 vdd.n2758 vdd.n2757 10.6151
R18429 vdd.n2757 vdd.n2756 10.6151
R18430 vdd.n2756 vdd.n2754 10.6151
R18431 vdd.n2754 vdd.n2753 10.6151
R18432 vdd.n2753 vdd.n2751 10.6151
R18433 vdd.n2751 vdd.n2750 10.6151
R18434 vdd.n2750 vdd.n2748 10.6151
R18435 vdd.n2748 vdd.n2747 10.6151
R18436 vdd.n2747 vdd.n2745 10.6151
R18437 vdd.n2745 vdd.n2744 10.6151
R18438 vdd.n2744 vdd.n836 10.6151
R18439 vdd.n2992 vdd.n836 10.6151
R18440 vdd.n2993 vdd.n2992 10.6151
R18441 vdd.n2854 vdd.n912 10.6151
R18442 vdd.n2854 vdd.n2853 10.6151
R18443 vdd.n2853 vdd.n2852 10.6151
R18444 vdd.n2852 vdd.n2850 10.6151
R18445 vdd.n2850 vdd.n2847 10.6151
R18446 vdd.n2847 vdd.n2846 10.6151
R18447 vdd.n2846 vdd.n2843 10.6151
R18448 vdd.n2843 vdd.n2842 10.6151
R18449 vdd.n2842 vdd.n2839 10.6151
R18450 vdd.n2839 vdd.n2838 10.6151
R18451 vdd.n2838 vdd.n2835 10.6151
R18452 vdd.n2835 vdd.n2834 10.6151
R18453 vdd.n2834 vdd.n2831 10.6151
R18454 vdd.n2831 vdd.n2830 10.6151
R18455 vdd.n2830 vdd.n2827 10.6151
R18456 vdd.n2827 vdd.n2826 10.6151
R18457 vdd.n2826 vdd.n2823 10.6151
R18458 vdd.n2823 vdd.n2822 10.6151
R18459 vdd.n2822 vdd.n2819 10.6151
R18460 vdd.n2819 vdd.n2818 10.6151
R18461 vdd.n2818 vdd.n2815 10.6151
R18462 vdd.n2815 vdd.n2814 10.6151
R18463 vdd.n2814 vdd.n2811 10.6151
R18464 vdd.n2811 vdd.n2810 10.6151
R18465 vdd.n2810 vdd.n2807 10.6151
R18466 vdd.n2807 vdd.n2806 10.6151
R18467 vdd.n2806 vdd.n2803 10.6151
R18468 vdd.n2803 vdd.n2802 10.6151
R18469 vdd.n2802 vdd.n2799 10.6151
R18470 vdd.n2799 vdd.n2798 10.6151
R18471 vdd.n2798 vdd.n2795 10.6151
R18472 vdd.n2793 vdd.n2790 10.6151
R18473 vdd.n2790 vdd.n2789 10.6151
R18474 vdd.n2867 vdd.n2866 10.6151
R18475 vdd.n2868 vdd.n2867 10.6151
R18476 vdd.n2868 vdd.n902 10.6151
R18477 vdd.n2878 vdd.n902 10.6151
R18478 vdd.n2879 vdd.n2878 10.6151
R18479 vdd.n2880 vdd.n2879 10.6151
R18480 vdd.n2880 vdd.n889 10.6151
R18481 vdd.n2890 vdd.n889 10.6151
R18482 vdd.n2891 vdd.n2890 10.6151
R18483 vdd.n2892 vdd.n2891 10.6151
R18484 vdd.n2892 vdd.n878 10.6151
R18485 vdd.n2902 vdd.n878 10.6151
R18486 vdd.n2903 vdd.n2902 10.6151
R18487 vdd.n2904 vdd.n2903 10.6151
R18488 vdd.n2904 vdd.n866 10.6151
R18489 vdd.n2914 vdd.n866 10.6151
R18490 vdd.n2915 vdd.n2914 10.6151
R18491 vdd.n2916 vdd.n2915 10.6151
R18492 vdd.n2916 vdd.n855 10.6151
R18493 vdd.n2928 vdd.n855 10.6151
R18494 vdd.n2929 vdd.n2928 10.6151
R18495 vdd.n2930 vdd.n2929 10.6151
R18496 vdd.n2930 vdd.n841 10.6151
R18497 vdd.n2985 vdd.n841 10.6151
R18498 vdd.n2986 vdd.n2985 10.6151
R18499 vdd.n2987 vdd.n2986 10.6151
R18500 vdd.n2987 vdd.n810 10.6151
R18501 vdd.n3057 vdd.n810 10.6151
R18502 vdd.n3056 vdd.n3055 10.6151
R18503 vdd.n3055 vdd.n811 10.6151
R18504 vdd.n812 vdd.n811 10.6151
R18505 vdd.n3048 vdd.n812 10.6151
R18506 vdd.n3048 vdd.n3047 10.6151
R18507 vdd.n3047 vdd.n3046 10.6151
R18508 vdd.n3046 vdd.n814 10.6151
R18509 vdd.n3041 vdd.n814 10.6151
R18510 vdd.n3041 vdd.n3040 10.6151
R18511 vdd.n3040 vdd.n3039 10.6151
R18512 vdd.n3039 vdd.n817 10.6151
R18513 vdd.n3034 vdd.n817 10.6151
R18514 vdd.n3034 vdd.n3033 10.6151
R18515 vdd.n3033 vdd.n3032 10.6151
R18516 vdd.n3032 vdd.n820 10.6151
R18517 vdd.n3027 vdd.n820 10.6151
R18518 vdd.n3027 vdd.n731 10.6151
R18519 vdd.n3023 vdd.n731 10.6151
R18520 vdd.n3023 vdd.n3022 10.6151
R18521 vdd.n3022 vdd.n3021 10.6151
R18522 vdd.n3021 vdd.n823 10.6151
R18523 vdd.n3016 vdd.n823 10.6151
R18524 vdd.n3016 vdd.n3015 10.6151
R18525 vdd.n3015 vdd.n3014 10.6151
R18526 vdd.n3014 vdd.n826 10.6151
R18527 vdd.n3009 vdd.n826 10.6151
R18528 vdd.n3009 vdd.n3008 10.6151
R18529 vdd.n3008 vdd.n3007 10.6151
R18530 vdd.n3007 vdd.n829 10.6151
R18531 vdd.n3002 vdd.n829 10.6151
R18532 vdd.n3002 vdd.n3001 10.6151
R18533 vdd.n2999 vdd.n834 10.6151
R18534 vdd.n2994 vdd.n834 10.6151
R18535 vdd.n2975 vdd.n2936 10.6151
R18536 vdd.n2970 vdd.n2936 10.6151
R18537 vdd.n2970 vdd.n2969 10.6151
R18538 vdd.n2969 vdd.n2968 10.6151
R18539 vdd.n2968 vdd.n2938 10.6151
R18540 vdd.n2963 vdd.n2938 10.6151
R18541 vdd.n2963 vdd.n2962 10.6151
R18542 vdd.n2962 vdd.n2961 10.6151
R18543 vdd.n2961 vdd.n2941 10.6151
R18544 vdd.n2956 vdd.n2941 10.6151
R18545 vdd.n2956 vdd.n2955 10.6151
R18546 vdd.n2955 vdd.n2954 10.6151
R18547 vdd.n2954 vdd.n2944 10.6151
R18548 vdd.n2949 vdd.n2944 10.6151
R18549 vdd.n2949 vdd.n2948 10.6151
R18550 vdd.n2948 vdd.n785 10.6151
R18551 vdd.n3092 vdd.n785 10.6151
R18552 vdd.n3092 vdd.n786 10.6151
R18553 vdd.n788 vdd.n786 10.6151
R18554 vdd.n3085 vdd.n788 10.6151
R18555 vdd.n3085 vdd.n3084 10.6151
R18556 vdd.n3084 vdd.n3083 10.6151
R18557 vdd.n3083 vdd.n790 10.6151
R18558 vdd.n3078 vdd.n790 10.6151
R18559 vdd.n3078 vdd.n3077 10.6151
R18560 vdd.n3077 vdd.n3076 10.6151
R18561 vdd.n3076 vdd.n793 10.6151
R18562 vdd.n3071 vdd.n793 10.6151
R18563 vdd.n3071 vdd.n3070 10.6151
R18564 vdd.n3070 vdd.n3069 10.6151
R18565 vdd.n3069 vdd.n796 10.6151
R18566 vdd.n3064 vdd.n3063 10.6151
R18567 vdd.n3063 vdd.n3062 10.6151
R18568 vdd.n2710 vdd.n2708 10.6151
R18569 vdd.n2711 vdd.n2710 10.6151
R18570 vdd.n2779 vdd.n2711 10.6151
R18571 vdd.n2779 vdd.n2778 10.6151
R18572 vdd.n2778 vdd.n2777 10.6151
R18573 vdd.n2777 vdd.n2775 10.6151
R18574 vdd.n2775 vdd.n2774 10.6151
R18575 vdd.n2774 vdd.n2772 10.6151
R18576 vdd.n2772 vdd.n2771 10.6151
R18577 vdd.n2771 vdd.n2769 10.6151
R18578 vdd.n2769 vdd.n2768 10.6151
R18579 vdd.n2768 vdd.n2766 10.6151
R18580 vdd.n2766 vdd.n2765 10.6151
R18581 vdd.n2765 vdd.n2763 10.6151
R18582 vdd.n2763 vdd.n2762 10.6151
R18583 vdd.n2762 vdd.n2728 10.6151
R18584 vdd.n2728 vdd.n2727 10.6151
R18585 vdd.n2727 vdd.n2725 10.6151
R18586 vdd.n2725 vdd.n2724 10.6151
R18587 vdd.n2724 vdd.n2722 10.6151
R18588 vdd.n2722 vdd.n2721 10.6151
R18589 vdd.n2721 vdd.n2719 10.6151
R18590 vdd.n2719 vdd.n2718 10.6151
R18591 vdd.n2718 vdd.n2716 10.6151
R18592 vdd.n2716 vdd.n2715 10.6151
R18593 vdd.n2715 vdd.n2713 10.6151
R18594 vdd.n2713 vdd.n2712 10.6151
R18595 vdd.n2712 vdd.n802 10.6151
R18596 vdd.n2861 vdd.n2860 10.6151
R18597 vdd.n2860 vdd.n917 10.6151
R18598 vdd.n2645 vdd.n917 10.6151
R18599 vdd.n2648 vdd.n2645 10.6151
R18600 vdd.n2649 vdd.n2648 10.6151
R18601 vdd.n2652 vdd.n2649 10.6151
R18602 vdd.n2653 vdd.n2652 10.6151
R18603 vdd.n2656 vdd.n2653 10.6151
R18604 vdd.n2657 vdd.n2656 10.6151
R18605 vdd.n2660 vdd.n2657 10.6151
R18606 vdd.n2661 vdd.n2660 10.6151
R18607 vdd.n2664 vdd.n2661 10.6151
R18608 vdd.n2665 vdd.n2664 10.6151
R18609 vdd.n2668 vdd.n2665 10.6151
R18610 vdd.n2669 vdd.n2668 10.6151
R18611 vdd.n2672 vdd.n2669 10.6151
R18612 vdd.n2673 vdd.n2672 10.6151
R18613 vdd.n2676 vdd.n2673 10.6151
R18614 vdd.n2677 vdd.n2676 10.6151
R18615 vdd.n2680 vdd.n2677 10.6151
R18616 vdd.n2681 vdd.n2680 10.6151
R18617 vdd.n2684 vdd.n2681 10.6151
R18618 vdd.n2685 vdd.n2684 10.6151
R18619 vdd.n2688 vdd.n2685 10.6151
R18620 vdd.n2689 vdd.n2688 10.6151
R18621 vdd.n2692 vdd.n2689 10.6151
R18622 vdd.n2693 vdd.n2692 10.6151
R18623 vdd.n2696 vdd.n2693 10.6151
R18624 vdd.n2697 vdd.n2696 10.6151
R18625 vdd.n2700 vdd.n2697 10.6151
R18626 vdd.n2701 vdd.n2700 10.6151
R18627 vdd.n2706 vdd.n2704 10.6151
R18628 vdd.n2707 vdd.n2706 10.6151
R18629 vdd.n2862 vdd.n907 10.6151
R18630 vdd.n2872 vdd.n907 10.6151
R18631 vdd.n2873 vdd.n2872 10.6151
R18632 vdd.n2874 vdd.n2873 10.6151
R18633 vdd.n2874 vdd.n895 10.6151
R18634 vdd.n2884 vdd.n895 10.6151
R18635 vdd.n2885 vdd.n2884 10.6151
R18636 vdd.n2886 vdd.n2885 10.6151
R18637 vdd.n2886 vdd.n884 10.6151
R18638 vdd.n2896 vdd.n884 10.6151
R18639 vdd.n2897 vdd.n2896 10.6151
R18640 vdd.n2898 vdd.n2897 10.6151
R18641 vdd.n2898 vdd.n872 10.6151
R18642 vdd.n2908 vdd.n872 10.6151
R18643 vdd.n2909 vdd.n2908 10.6151
R18644 vdd.n2910 vdd.n2909 10.6151
R18645 vdd.n2910 vdd.n861 10.6151
R18646 vdd.n2920 vdd.n861 10.6151
R18647 vdd.n2921 vdd.n2920 10.6151
R18648 vdd.n2924 vdd.n2921 10.6151
R18649 vdd.n2934 vdd.n849 10.6151
R18650 vdd.n2935 vdd.n2934 10.6151
R18651 vdd.n2981 vdd.n2935 10.6151
R18652 vdd.n2981 vdd.n2980 10.6151
R18653 vdd.n2980 vdd.n2979 10.6151
R18654 vdd.n2979 vdd.n2978 10.6151
R18655 vdd.n2978 vdd.n2976 10.6151
R18656 vdd.n2373 vdd.n1041 10.6151
R18657 vdd.n2383 vdd.n1041 10.6151
R18658 vdd.n2384 vdd.n2383 10.6151
R18659 vdd.n2385 vdd.n2384 10.6151
R18660 vdd.n2385 vdd.n1028 10.6151
R18661 vdd.n2395 vdd.n1028 10.6151
R18662 vdd.n2396 vdd.n2395 10.6151
R18663 vdd.n2398 vdd.n1016 10.6151
R18664 vdd.n2408 vdd.n1016 10.6151
R18665 vdd.n2409 vdd.n2408 10.6151
R18666 vdd.n2410 vdd.n2409 10.6151
R18667 vdd.n2410 vdd.n1004 10.6151
R18668 vdd.n2420 vdd.n1004 10.6151
R18669 vdd.n2421 vdd.n2420 10.6151
R18670 vdd.n2422 vdd.n2421 10.6151
R18671 vdd.n2422 vdd.n993 10.6151
R18672 vdd.n2432 vdd.n993 10.6151
R18673 vdd.n2433 vdd.n2432 10.6151
R18674 vdd.n2434 vdd.n2433 10.6151
R18675 vdd.n2434 vdd.n981 10.6151
R18676 vdd.n2444 vdd.n981 10.6151
R18677 vdd.n2445 vdd.n2444 10.6151
R18678 vdd.n2448 vdd.n2445 10.6151
R18679 vdd.n2448 vdd.n2447 10.6151
R18680 vdd.n2447 vdd.n2446 10.6151
R18681 vdd.n2446 vdd.n964 10.6151
R18682 vdd.n2530 vdd.n964 10.6151
R18683 vdd.n2529 vdd.n2528 10.6151
R18684 vdd.n2528 vdd.n2525 10.6151
R18685 vdd.n2525 vdd.n2524 10.6151
R18686 vdd.n2524 vdd.n2521 10.6151
R18687 vdd.n2521 vdd.n2520 10.6151
R18688 vdd.n2520 vdd.n2517 10.6151
R18689 vdd.n2517 vdd.n2516 10.6151
R18690 vdd.n2516 vdd.n2513 10.6151
R18691 vdd.n2513 vdd.n2512 10.6151
R18692 vdd.n2512 vdd.n2509 10.6151
R18693 vdd.n2509 vdd.n2508 10.6151
R18694 vdd.n2508 vdd.n2505 10.6151
R18695 vdd.n2505 vdd.n2504 10.6151
R18696 vdd.n2504 vdd.n2501 10.6151
R18697 vdd.n2501 vdd.n2500 10.6151
R18698 vdd.n2500 vdd.n2497 10.6151
R18699 vdd.n2497 vdd.n2496 10.6151
R18700 vdd.n2496 vdd.n2493 10.6151
R18701 vdd.n2493 vdd.n2492 10.6151
R18702 vdd.n2492 vdd.n2489 10.6151
R18703 vdd.n2489 vdd.n2488 10.6151
R18704 vdd.n2488 vdd.n2485 10.6151
R18705 vdd.n2485 vdd.n2484 10.6151
R18706 vdd.n2484 vdd.n2481 10.6151
R18707 vdd.n2481 vdd.n2480 10.6151
R18708 vdd.n2480 vdd.n2477 10.6151
R18709 vdd.n2477 vdd.n2476 10.6151
R18710 vdd.n2476 vdd.n2473 10.6151
R18711 vdd.n2473 vdd.n2472 10.6151
R18712 vdd.n2472 vdd.n2469 10.6151
R18713 vdd.n2469 vdd.n2468 10.6151
R18714 vdd.n2465 vdd.n2464 10.6151
R18715 vdd.n2464 vdd.n2462 10.6151
R18716 vdd.n2221 vdd.n2219 10.6151
R18717 vdd.n2222 vdd.n2221 10.6151
R18718 vdd.n2224 vdd.n2222 10.6151
R18719 vdd.n2225 vdd.n2224 10.6151
R18720 vdd.n2227 vdd.n2225 10.6151
R18721 vdd.n2228 vdd.n2227 10.6151
R18722 vdd.n2230 vdd.n2228 10.6151
R18723 vdd.n2231 vdd.n2230 10.6151
R18724 vdd.n2233 vdd.n2231 10.6151
R18725 vdd.n2234 vdd.n2233 10.6151
R18726 vdd.n2236 vdd.n2234 10.6151
R18727 vdd.n2237 vdd.n2236 10.6151
R18728 vdd.n2255 vdd.n2237 10.6151
R18729 vdd.n2255 vdd.n2254 10.6151
R18730 vdd.n2254 vdd.n2253 10.6151
R18731 vdd.n2253 vdd.n2251 10.6151
R18732 vdd.n2251 vdd.n2250 10.6151
R18733 vdd.n2250 vdd.n2248 10.6151
R18734 vdd.n2248 vdd.n2247 10.6151
R18735 vdd.n2247 vdd.n2245 10.6151
R18736 vdd.n2245 vdd.n2244 10.6151
R18737 vdd.n2244 vdd.n2242 10.6151
R18738 vdd.n2242 vdd.n2241 10.6151
R18739 vdd.n2241 vdd.n2239 10.6151
R18740 vdd.n2239 vdd.n2238 10.6151
R18741 vdd.n2238 vdd.n968 10.6151
R18742 vdd.n2460 vdd.n968 10.6151
R18743 vdd.n2461 vdd.n2460 10.6151
R18744 vdd.n2372 vdd.n2371 10.6151
R18745 vdd.n2371 vdd.n1053 10.6151
R18746 vdd.n2365 vdd.n1053 10.6151
R18747 vdd.n2365 vdd.n2364 10.6151
R18748 vdd.n2364 vdd.n2363 10.6151
R18749 vdd.n2363 vdd.n1055 10.6151
R18750 vdd.n2357 vdd.n1055 10.6151
R18751 vdd.n2357 vdd.n2356 10.6151
R18752 vdd.n2356 vdd.n2355 10.6151
R18753 vdd.n2355 vdd.n1057 10.6151
R18754 vdd.n2349 vdd.n1057 10.6151
R18755 vdd.n2349 vdd.n2348 10.6151
R18756 vdd.n2348 vdd.n2347 10.6151
R18757 vdd.n2347 vdd.n1059 10.6151
R18758 vdd.n2341 vdd.n1059 10.6151
R18759 vdd.n2341 vdd.n2340 10.6151
R18760 vdd.n2340 vdd.n2339 10.6151
R18761 vdd.n2339 vdd.n1063 10.6151
R18762 vdd.n2187 vdd.n1063 10.6151
R18763 vdd.n2188 vdd.n2187 10.6151
R18764 vdd.n2188 vdd.n2183 10.6151
R18765 vdd.n2194 vdd.n2183 10.6151
R18766 vdd.n2195 vdd.n2194 10.6151
R18767 vdd.n2196 vdd.n2195 10.6151
R18768 vdd.n2196 vdd.n2181 10.6151
R18769 vdd.n2202 vdd.n2181 10.6151
R18770 vdd.n2203 vdd.n2202 10.6151
R18771 vdd.n2204 vdd.n2203 10.6151
R18772 vdd.n2204 vdd.n2179 10.6151
R18773 vdd.n2210 vdd.n2179 10.6151
R18774 vdd.n2211 vdd.n2210 10.6151
R18775 vdd.n2213 vdd.n2175 10.6151
R18776 vdd.n2218 vdd.n2175 10.6151
R18777 vdd.n1851 vdd.t23 10.5435
R18778 vdd.n656 vdd.t132 10.5435
R18779 vdd.n316 vdd.n298 10.4732
R18780 vdd.n257 vdd.n239 10.4732
R18781 vdd.n214 vdd.n196 10.4732
R18782 vdd.n155 vdd.n137 10.4732
R18783 vdd.n113 vdd.n95 10.4732
R18784 vdd.n54 vdd.n36 10.4732
R18785 vdd.n1735 vdd.n1717 10.4732
R18786 vdd.n1794 vdd.n1776 10.4732
R18787 vdd.n1633 vdd.n1615 10.4732
R18788 vdd.n1692 vdd.n1674 10.4732
R18789 vdd.n1532 vdd.n1514 10.4732
R18790 vdd.n1591 vdd.n1573 10.4732
R18791 vdd.t112 vdd.n1825 10.3167
R18792 vdd.n3300 vdd.t75 10.3167
R18793 vdd.n1502 vdd.t43 10.09
R18794 vdd.n3394 vdd.t41 10.09
R18795 vdd.t109 vdd.n1155 9.86327
R18796 vdd.n3385 vdd.t39 9.86327
R18797 vdd.n315 vdd.n300 9.69747
R18798 vdd.n256 vdd.n241 9.69747
R18799 vdd.n213 vdd.n198 9.69747
R18800 vdd.n154 vdd.n139 9.69747
R18801 vdd.n112 vdd.n97 9.69747
R18802 vdd.n53 vdd.n38 9.69747
R18803 vdd.n1734 vdd.n1719 9.69747
R18804 vdd.n1793 vdd.n1778 9.69747
R18805 vdd.n1632 vdd.n1617 9.69747
R18806 vdd.n1691 vdd.n1676 9.69747
R18807 vdd.n1531 vdd.n1516 9.69747
R18808 vdd.n1590 vdd.n1575 9.69747
R18809 vdd.n2315 vdd.n2314 9.67831
R18810 vdd.n3216 vdd.n731 9.67831
R18811 vdd.n3093 vdd.n3092 9.67831
R18812 vdd.n2339 vdd.n2338 9.67831
R18813 vdd.n1461 vdd.t60 9.63654
R18814 vdd.n3331 vdd.t37 9.63654
R18815 vdd.n331 vdd.n330 9.45567
R18816 vdd.n272 vdd.n271 9.45567
R18817 vdd.n229 vdd.n228 9.45567
R18818 vdd.n170 vdd.n169 9.45567
R18819 vdd.n128 vdd.n127 9.45567
R18820 vdd.n69 vdd.n68 9.45567
R18821 vdd.n1750 vdd.n1749 9.45567
R18822 vdd.n1809 vdd.n1808 9.45567
R18823 vdd.n1648 vdd.n1647 9.45567
R18824 vdd.n1707 vdd.n1706 9.45567
R18825 vdd.n1547 vdd.n1546 9.45567
R18826 vdd.n1606 vdd.n1605 9.45567
R18827 vdd.n1435 vdd.t25 9.40981
R18828 vdd.n3363 vdd.t82 9.40981
R18829 vdd.n2075 vdd.n1929 9.3005
R18830 vdd.n2074 vdd.n2073 9.3005
R18831 vdd.n1935 vdd.n1934 9.3005
R18832 vdd.n2068 vdd.n1939 9.3005
R18833 vdd.n2067 vdd.n1940 9.3005
R18834 vdd.n2066 vdd.n1941 9.3005
R18835 vdd.n1945 vdd.n1942 9.3005
R18836 vdd.n2061 vdd.n1946 9.3005
R18837 vdd.n2060 vdd.n1947 9.3005
R18838 vdd.n2059 vdd.n1948 9.3005
R18839 vdd.n1952 vdd.n1949 9.3005
R18840 vdd.n2054 vdd.n1953 9.3005
R18841 vdd.n2053 vdd.n1954 9.3005
R18842 vdd.n2052 vdd.n1955 9.3005
R18843 vdd.n1959 vdd.n1956 9.3005
R18844 vdd.n2047 vdd.n1960 9.3005
R18845 vdd.n2046 vdd.n1961 9.3005
R18846 vdd.n2045 vdd.n1962 9.3005
R18847 vdd.n1966 vdd.n1963 9.3005
R18848 vdd.n2040 vdd.n1967 9.3005
R18849 vdd.n2039 vdd.n1968 9.3005
R18850 vdd.n2038 vdd.n2037 9.3005
R18851 vdd.n2036 vdd.n1969 9.3005
R18852 vdd.n2035 vdd.n2034 9.3005
R18853 vdd.n1975 vdd.n1974 9.3005
R18854 vdd.n2029 vdd.n1979 9.3005
R18855 vdd.n2028 vdd.n1980 9.3005
R18856 vdd.n2027 vdd.n1981 9.3005
R18857 vdd.n1985 vdd.n1982 9.3005
R18858 vdd.n2022 vdd.n1986 9.3005
R18859 vdd.n2021 vdd.n1987 9.3005
R18860 vdd.n2020 vdd.n1988 9.3005
R18861 vdd.n1992 vdd.n1989 9.3005
R18862 vdd.n2015 vdd.n1993 9.3005
R18863 vdd.n2014 vdd.n1994 9.3005
R18864 vdd.n2013 vdd.n1995 9.3005
R18865 vdd.n1997 vdd.n1996 9.3005
R18866 vdd.n2008 vdd.n1064 9.3005
R18867 vdd.n2077 vdd.n2076 9.3005
R18868 vdd.n2101 vdd.n2100 9.3005
R18869 vdd.n1907 vdd.n1906 9.3005
R18870 vdd.n1912 vdd.n1910 9.3005
R18871 vdd.n2093 vdd.n1913 9.3005
R18872 vdd.n2092 vdd.n1914 9.3005
R18873 vdd.n2091 vdd.n1915 9.3005
R18874 vdd.n1919 vdd.n1916 9.3005
R18875 vdd.n2086 vdd.n1920 9.3005
R18876 vdd.n2085 vdd.n1921 9.3005
R18877 vdd.n2084 vdd.n1922 9.3005
R18878 vdd.n1926 vdd.n1923 9.3005
R18879 vdd.n2079 vdd.n1927 9.3005
R18880 vdd.n2078 vdd.n1928 9.3005
R18881 vdd.n2323 vdd.n1900 9.3005
R18882 vdd.n2325 vdd.n2324 9.3005
R18883 vdd.n1815 vdd.n1814 9.3005
R18884 vdd.n1124 vdd.n1123 9.3005
R18885 vdd.n1829 vdd.n1828 9.3005
R18886 vdd.n1830 vdd.n1122 9.3005
R18887 vdd.n1832 vdd.n1831 9.3005
R18888 vdd.n1113 vdd.n1112 9.3005
R18889 vdd.n1846 vdd.n1845 9.3005
R18890 vdd.n1847 vdd.n1111 9.3005
R18891 vdd.n1849 vdd.n1848 9.3005
R18892 vdd.n1102 vdd.n1101 9.3005
R18893 vdd.n1862 vdd.n1861 9.3005
R18894 vdd.n1863 vdd.n1100 9.3005
R18895 vdd.n1865 vdd.n1864 9.3005
R18896 vdd.n1090 vdd.n1089 9.3005
R18897 vdd.n1879 vdd.n1878 9.3005
R18898 vdd.n1880 vdd.n1088 9.3005
R18899 vdd.n1882 vdd.n1881 9.3005
R18900 vdd.n1078 vdd.n1077 9.3005
R18901 vdd.n1898 vdd.n1897 9.3005
R18902 vdd.n1899 vdd.n1076 9.3005
R18903 vdd.n2327 vdd.n2326 9.3005
R18904 vdd.n307 vdd.n306 9.3005
R18905 vdd.n302 vdd.n301 9.3005
R18906 vdd.n313 vdd.n312 9.3005
R18907 vdd.n315 vdd.n314 9.3005
R18908 vdd.n298 vdd.n297 9.3005
R18909 vdd.n321 vdd.n320 9.3005
R18910 vdd.n323 vdd.n322 9.3005
R18911 vdd.n295 vdd.n292 9.3005
R18912 vdd.n330 vdd.n329 9.3005
R18913 vdd.n248 vdd.n247 9.3005
R18914 vdd.n243 vdd.n242 9.3005
R18915 vdd.n254 vdd.n253 9.3005
R18916 vdd.n256 vdd.n255 9.3005
R18917 vdd.n239 vdd.n238 9.3005
R18918 vdd.n262 vdd.n261 9.3005
R18919 vdd.n264 vdd.n263 9.3005
R18920 vdd.n236 vdd.n233 9.3005
R18921 vdd.n271 vdd.n270 9.3005
R18922 vdd.n205 vdd.n204 9.3005
R18923 vdd.n200 vdd.n199 9.3005
R18924 vdd.n211 vdd.n210 9.3005
R18925 vdd.n213 vdd.n212 9.3005
R18926 vdd.n196 vdd.n195 9.3005
R18927 vdd.n219 vdd.n218 9.3005
R18928 vdd.n221 vdd.n220 9.3005
R18929 vdd.n193 vdd.n190 9.3005
R18930 vdd.n228 vdd.n227 9.3005
R18931 vdd.n146 vdd.n145 9.3005
R18932 vdd.n141 vdd.n140 9.3005
R18933 vdd.n152 vdd.n151 9.3005
R18934 vdd.n154 vdd.n153 9.3005
R18935 vdd.n137 vdd.n136 9.3005
R18936 vdd.n160 vdd.n159 9.3005
R18937 vdd.n162 vdd.n161 9.3005
R18938 vdd.n134 vdd.n131 9.3005
R18939 vdd.n169 vdd.n168 9.3005
R18940 vdd.n104 vdd.n103 9.3005
R18941 vdd.n99 vdd.n98 9.3005
R18942 vdd.n110 vdd.n109 9.3005
R18943 vdd.n112 vdd.n111 9.3005
R18944 vdd.n95 vdd.n94 9.3005
R18945 vdd.n118 vdd.n117 9.3005
R18946 vdd.n120 vdd.n119 9.3005
R18947 vdd.n92 vdd.n89 9.3005
R18948 vdd.n127 vdd.n126 9.3005
R18949 vdd.n45 vdd.n44 9.3005
R18950 vdd.n40 vdd.n39 9.3005
R18951 vdd.n51 vdd.n50 9.3005
R18952 vdd.n53 vdd.n52 9.3005
R18953 vdd.n36 vdd.n35 9.3005
R18954 vdd.n59 vdd.n58 9.3005
R18955 vdd.n61 vdd.n60 9.3005
R18956 vdd.n33 vdd.n30 9.3005
R18957 vdd.n68 vdd.n67 9.3005
R18958 vdd.n3138 vdd.n3137 9.3005
R18959 vdd.n3141 vdd.n766 9.3005
R18960 vdd.n3142 vdd.n765 9.3005
R18961 vdd.n3145 vdd.n764 9.3005
R18962 vdd.n3146 vdd.n763 9.3005
R18963 vdd.n3149 vdd.n762 9.3005
R18964 vdd.n3150 vdd.n761 9.3005
R18965 vdd.n3153 vdd.n760 9.3005
R18966 vdd.n3154 vdd.n759 9.3005
R18967 vdd.n3157 vdd.n758 9.3005
R18968 vdd.n3158 vdd.n757 9.3005
R18969 vdd.n3161 vdd.n756 9.3005
R18970 vdd.n3162 vdd.n755 9.3005
R18971 vdd.n3165 vdd.n754 9.3005
R18972 vdd.n3166 vdd.n753 9.3005
R18973 vdd.n3169 vdd.n752 9.3005
R18974 vdd.n3170 vdd.n751 9.3005
R18975 vdd.n3173 vdd.n750 9.3005
R18976 vdd.n3174 vdd.n749 9.3005
R18977 vdd.n3177 vdd.n748 9.3005
R18978 vdd.n3181 vdd.n3180 9.3005
R18979 vdd.n3182 vdd.n747 9.3005
R18980 vdd.n3186 vdd.n3183 9.3005
R18981 vdd.n3189 vdd.n746 9.3005
R18982 vdd.n3190 vdd.n745 9.3005
R18983 vdd.n3193 vdd.n744 9.3005
R18984 vdd.n3194 vdd.n743 9.3005
R18985 vdd.n3197 vdd.n742 9.3005
R18986 vdd.n3198 vdd.n741 9.3005
R18987 vdd.n3201 vdd.n740 9.3005
R18988 vdd.n3202 vdd.n739 9.3005
R18989 vdd.n3205 vdd.n738 9.3005
R18990 vdd.n3206 vdd.n737 9.3005
R18991 vdd.n3209 vdd.n736 9.3005
R18992 vdd.n3210 vdd.n735 9.3005
R18993 vdd.n3213 vdd.n730 9.3005
R18994 vdd.n3219 vdd.n727 9.3005
R18995 vdd.n3220 vdd.n726 9.3005
R18996 vdd.n3234 vdd.n3233 9.3005
R18997 vdd.n3235 vdd.n681 9.3005
R18998 vdd.n3237 vdd.n3236 9.3005
R18999 vdd.n671 vdd.n670 9.3005
R19000 vdd.n3251 vdd.n3250 9.3005
R19001 vdd.n3252 vdd.n669 9.3005
R19002 vdd.n3254 vdd.n3253 9.3005
R19003 vdd.n660 vdd.n659 9.3005
R19004 vdd.n3267 vdd.n3266 9.3005
R19005 vdd.n3268 vdd.n658 9.3005
R19006 vdd.n3270 vdd.n3269 9.3005
R19007 vdd.n648 vdd.n647 9.3005
R19008 vdd.n3284 vdd.n3283 9.3005
R19009 vdd.n3285 vdd.n646 9.3005
R19010 vdd.n3287 vdd.n3286 9.3005
R19011 vdd.n637 vdd.n636 9.3005
R19012 vdd.n3303 vdd.n3302 9.3005
R19013 vdd.n3304 vdd.n635 9.3005
R19014 vdd.n3306 vdd.n3305 9.3005
R19015 vdd.n336 vdd.n334 9.3005
R19016 vdd.n683 vdd.n682 9.3005
R19017 vdd.n3398 vdd.n3397 9.3005
R19018 vdd.n337 vdd.n335 9.3005
R19019 vdd.n3391 vdd.n346 9.3005
R19020 vdd.n3390 vdd.n347 9.3005
R19021 vdd.n3389 vdd.n348 9.3005
R19022 vdd.n355 vdd.n349 9.3005
R19023 vdd.n3383 vdd.n356 9.3005
R19024 vdd.n3382 vdd.n357 9.3005
R19025 vdd.n3381 vdd.n358 9.3005
R19026 vdd.n366 vdd.n359 9.3005
R19027 vdd.n3375 vdd.n367 9.3005
R19028 vdd.n3374 vdd.n368 9.3005
R19029 vdd.n3373 vdd.n369 9.3005
R19030 vdd.n377 vdd.n370 9.3005
R19031 vdd.n3367 vdd.n378 9.3005
R19032 vdd.n3366 vdd.n379 9.3005
R19033 vdd.n3365 vdd.n380 9.3005
R19034 vdd.n388 vdd.n381 9.3005
R19035 vdd.n3359 vdd.n389 9.3005
R19036 vdd.n3358 vdd.n390 9.3005
R19037 vdd.n3357 vdd.n391 9.3005
R19038 vdd.n466 vdd.n463 9.3005
R19039 vdd.n470 vdd.n469 9.3005
R19040 vdd.n471 vdd.n462 9.3005
R19041 vdd.n475 vdd.n472 9.3005
R19042 vdd.n476 vdd.n461 9.3005
R19043 vdd.n480 vdd.n479 9.3005
R19044 vdd.n481 vdd.n460 9.3005
R19045 vdd.n485 vdd.n482 9.3005
R19046 vdd.n486 vdd.n459 9.3005
R19047 vdd.n490 vdd.n489 9.3005
R19048 vdd.n491 vdd.n458 9.3005
R19049 vdd.n495 vdd.n492 9.3005
R19050 vdd.n496 vdd.n457 9.3005
R19051 vdd.n500 vdd.n499 9.3005
R19052 vdd.n501 vdd.n456 9.3005
R19053 vdd.n505 vdd.n502 9.3005
R19054 vdd.n506 vdd.n455 9.3005
R19055 vdd.n510 vdd.n509 9.3005
R19056 vdd.n511 vdd.n454 9.3005
R19057 vdd.n515 vdd.n512 9.3005
R19058 vdd.n516 vdd.n451 9.3005
R19059 vdd.n520 vdd.n519 9.3005
R19060 vdd.n521 vdd.n450 9.3005
R19061 vdd.n525 vdd.n522 9.3005
R19062 vdd.n526 vdd.n449 9.3005
R19063 vdd.n530 vdd.n529 9.3005
R19064 vdd.n531 vdd.n448 9.3005
R19065 vdd.n535 vdd.n532 9.3005
R19066 vdd.n536 vdd.n447 9.3005
R19067 vdd.n540 vdd.n539 9.3005
R19068 vdd.n541 vdd.n446 9.3005
R19069 vdd.n545 vdd.n542 9.3005
R19070 vdd.n546 vdd.n445 9.3005
R19071 vdd.n550 vdd.n549 9.3005
R19072 vdd.n551 vdd.n444 9.3005
R19073 vdd.n555 vdd.n552 9.3005
R19074 vdd.n556 vdd.n443 9.3005
R19075 vdd.n560 vdd.n559 9.3005
R19076 vdd.n561 vdd.n442 9.3005
R19077 vdd.n565 vdd.n562 9.3005
R19078 vdd.n566 vdd.n439 9.3005
R19079 vdd.n570 vdd.n569 9.3005
R19080 vdd.n571 vdd.n438 9.3005
R19081 vdd.n575 vdd.n572 9.3005
R19082 vdd.n576 vdd.n437 9.3005
R19083 vdd.n580 vdd.n579 9.3005
R19084 vdd.n581 vdd.n436 9.3005
R19085 vdd.n585 vdd.n582 9.3005
R19086 vdd.n586 vdd.n435 9.3005
R19087 vdd.n590 vdd.n589 9.3005
R19088 vdd.n591 vdd.n434 9.3005
R19089 vdd.n595 vdd.n592 9.3005
R19090 vdd.n596 vdd.n433 9.3005
R19091 vdd.n600 vdd.n599 9.3005
R19092 vdd.n601 vdd.n432 9.3005
R19093 vdd.n605 vdd.n602 9.3005
R19094 vdd.n606 vdd.n431 9.3005
R19095 vdd.n610 vdd.n609 9.3005
R19096 vdd.n611 vdd.n430 9.3005
R19097 vdd.n615 vdd.n612 9.3005
R19098 vdd.n617 vdd.n429 9.3005
R19099 vdd.n619 vdd.n618 9.3005
R19100 vdd.n3351 vdd.n3350 9.3005
R19101 vdd.n465 vdd.n464 9.3005
R19102 vdd.n3229 vdd.n3228 9.3005
R19103 vdd.n676 vdd.n675 9.3005
R19104 vdd.n3242 vdd.n3241 9.3005
R19105 vdd.n3243 vdd.n674 9.3005
R19106 vdd.n3245 vdd.n3244 9.3005
R19107 vdd.n666 vdd.n665 9.3005
R19108 vdd.n3259 vdd.n3258 9.3005
R19109 vdd.n3260 vdd.n664 9.3005
R19110 vdd.n3262 vdd.n3261 9.3005
R19111 vdd.n653 vdd.n652 9.3005
R19112 vdd.n3275 vdd.n3274 9.3005
R19113 vdd.n3276 vdd.n651 9.3005
R19114 vdd.n3278 vdd.n3277 9.3005
R19115 vdd.n642 vdd.n641 9.3005
R19116 vdd.n3292 vdd.n3291 9.3005
R19117 vdd.n3293 vdd.n640 9.3005
R19118 vdd.n3298 vdd.n3294 9.3005
R19119 vdd.n3297 vdd.n3296 9.3005
R19120 vdd.n3295 vdd.n631 9.3005
R19121 vdd.n3311 vdd.n630 9.3005
R19122 vdd.n3313 vdd.n3312 9.3005
R19123 vdd.n3314 vdd.n629 9.3005
R19124 vdd.n3316 vdd.n3315 9.3005
R19125 vdd.n3318 vdd.n628 9.3005
R19126 vdd.n3320 vdd.n3319 9.3005
R19127 vdd.n3321 vdd.n627 9.3005
R19128 vdd.n3323 vdd.n3322 9.3005
R19129 vdd.n3325 vdd.n626 9.3005
R19130 vdd.n3327 vdd.n3326 9.3005
R19131 vdd.n3328 vdd.n625 9.3005
R19132 vdd.n3330 vdd.n3329 9.3005
R19133 vdd.n3333 vdd.n624 9.3005
R19134 vdd.n3335 vdd.n3334 9.3005
R19135 vdd.n3336 vdd.n623 9.3005
R19136 vdd.n3338 vdd.n3337 9.3005
R19137 vdd.n3340 vdd.n622 9.3005
R19138 vdd.n3342 vdd.n3341 9.3005
R19139 vdd.n3343 vdd.n621 9.3005
R19140 vdd.n3345 vdd.n3344 9.3005
R19141 vdd.n3347 vdd.n620 9.3005
R19142 vdd.n3349 vdd.n3348 9.3005
R19143 vdd.n3227 vdd.n686 9.3005
R19144 vdd.n3226 vdd.n3225 9.3005
R19145 vdd.n3095 vdd.n687 9.3005
R19146 vdd.n3104 vdd.n783 9.3005
R19147 vdd.n3107 vdd.n782 9.3005
R19148 vdd.n3108 vdd.n781 9.3005
R19149 vdd.n3111 vdd.n780 9.3005
R19150 vdd.n3112 vdd.n779 9.3005
R19151 vdd.n3115 vdd.n778 9.3005
R19152 vdd.n3116 vdd.n777 9.3005
R19153 vdd.n3119 vdd.n776 9.3005
R19154 vdd.n3120 vdd.n775 9.3005
R19155 vdd.n3123 vdd.n774 9.3005
R19156 vdd.n3124 vdd.n773 9.3005
R19157 vdd.n3127 vdd.n772 9.3005
R19158 vdd.n3128 vdd.n771 9.3005
R19159 vdd.n3131 vdd.n770 9.3005
R19160 vdd.n3135 vdd.n3134 9.3005
R19161 vdd.n3136 vdd.n767 9.3005
R19162 vdd.n2337 vdd.n2336 9.3005
R19163 vdd.n2332 vdd.n1067 9.3005
R19164 vdd.n1430 vdd.n1429 9.3005
R19165 vdd.n1431 vdd.n1185 9.3005
R19166 vdd.n1433 vdd.n1432 9.3005
R19167 vdd.n1175 vdd.n1174 9.3005
R19168 vdd.n1447 vdd.n1446 9.3005
R19169 vdd.n1448 vdd.n1173 9.3005
R19170 vdd.n1450 vdd.n1449 9.3005
R19171 vdd.n1165 vdd.n1164 9.3005
R19172 vdd.n1464 vdd.n1463 9.3005
R19173 vdd.n1465 vdd.n1163 9.3005
R19174 vdd.n1467 vdd.n1466 9.3005
R19175 vdd.n1152 vdd.n1151 9.3005
R19176 vdd.n1480 vdd.n1479 9.3005
R19177 vdd.n1481 vdd.n1150 9.3005
R19178 vdd.n1483 vdd.n1482 9.3005
R19179 vdd.n1141 vdd.n1140 9.3005
R19180 vdd.n1497 vdd.n1496 9.3005
R19181 vdd.n1498 vdd.n1139 9.3005
R19182 vdd.n1500 vdd.n1499 9.3005
R19183 vdd.n1130 vdd.n1129 9.3005
R19184 vdd.n1820 vdd.n1819 9.3005
R19185 vdd.n1821 vdd.n1128 9.3005
R19186 vdd.n1823 vdd.n1822 9.3005
R19187 vdd.n1118 vdd.n1117 9.3005
R19188 vdd.n1837 vdd.n1836 9.3005
R19189 vdd.n1838 vdd.n1116 9.3005
R19190 vdd.n1840 vdd.n1839 9.3005
R19191 vdd.n1108 vdd.n1107 9.3005
R19192 vdd.n1854 vdd.n1853 9.3005
R19193 vdd.n1855 vdd.n1106 9.3005
R19194 vdd.n1857 vdd.n1856 9.3005
R19195 vdd.n1095 vdd.n1094 9.3005
R19196 vdd.n1870 vdd.n1869 9.3005
R19197 vdd.n1871 vdd.n1093 9.3005
R19198 vdd.n1873 vdd.n1872 9.3005
R19199 vdd.n1085 vdd.n1084 9.3005
R19200 vdd.n1887 vdd.n1886 9.3005
R19201 vdd.n1888 vdd.n1082 9.3005
R19202 vdd.n1892 vdd.n1891 9.3005
R19203 vdd.n1890 vdd.n1083 9.3005
R19204 vdd.n1889 vdd.n1072 9.3005
R19205 vdd.n1187 vdd.n1186 9.3005
R19206 vdd.n1323 vdd.n1322 9.3005
R19207 vdd.n1324 vdd.n1313 9.3005
R19208 vdd.n1326 vdd.n1325 9.3005
R19209 vdd.n1327 vdd.n1312 9.3005
R19210 vdd.n1329 vdd.n1328 9.3005
R19211 vdd.n1330 vdd.n1307 9.3005
R19212 vdd.n1332 vdd.n1331 9.3005
R19213 vdd.n1333 vdd.n1306 9.3005
R19214 vdd.n1335 vdd.n1334 9.3005
R19215 vdd.n1336 vdd.n1301 9.3005
R19216 vdd.n1338 vdd.n1337 9.3005
R19217 vdd.n1339 vdd.n1300 9.3005
R19218 vdd.n1341 vdd.n1340 9.3005
R19219 vdd.n1342 vdd.n1295 9.3005
R19220 vdd.n1344 vdd.n1343 9.3005
R19221 vdd.n1345 vdd.n1294 9.3005
R19222 vdd.n1347 vdd.n1346 9.3005
R19223 vdd.n1348 vdd.n1289 9.3005
R19224 vdd.n1350 vdd.n1349 9.3005
R19225 vdd.n1351 vdd.n1288 9.3005
R19226 vdd.n1353 vdd.n1352 9.3005
R19227 vdd.n1357 vdd.n1284 9.3005
R19228 vdd.n1359 vdd.n1358 9.3005
R19229 vdd.n1360 vdd.n1283 9.3005
R19230 vdd.n1362 vdd.n1361 9.3005
R19231 vdd.n1363 vdd.n1278 9.3005
R19232 vdd.n1365 vdd.n1364 9.3005
R19233 vdd.n1366 vdd.n1277 9.3005
R19234 vdd.n1368 vdd.n1367 9.3005
R19235 vdd.n1369 vdd.n1272 9.3005
R19236 vdd.n1371 vdd.n1370 9.3005
R19237 vdd.n1372 vdd.n1271 9.3005
R19238 vdd.n1374 vdd.n1373 9.3005
R19239 vdd.n1375 vdd.n1266 9.3005
R19240 vdd.n1377 vdd.n1376 9.3005
R19241 vdd.n1378 vdd.n1265 9.3005
R19242 vdd.n1380 vdd.n1379 9.3005
R19243 vdd.n1381 vdd.n1260 9.3005
R19244 vdd.n1383 vdd.n1382 9.3005
R19245 vdd.n1384 vdd.n1259 9.3005
R19246 vdd.n1386 vdd.n1385 9.3005
R19247 vdd.n1387 vdd.n1254 9.3005
R19248 vdd.n1389 vdd.n1388 9.3005
R19249 vdd.n1390 vdd.n1253 9.3005
R19250 vdd.n1392 vdd.n1391 9.3005
R19251 vdd.n1393 vdd.n1246 9.3005
R19252 vdd.n1395 vdd.n1394 9.3005
R19253 vdd.n1396 vdd.n1245 9.3005
R19254 vdd.n1398 vdd.n1397 9.3005
R19255 vdd.n1399 vdd.n1240 9.3005
R19256 vdd.n1401 vdd.n1400 9.3005
R19257 vdd.n1402 vdd.n1239 9.3005
R19258 vdd.n1404 vdd.n1403 9.3005
R19259 vdd.n1405 vdd.n1234 9.3005
R19260 vdd.n1407 vdd.n1406 9.3005
R19261 vdd.n1408 vdd.n1233 9.3005
R19262 vdd.n1410 vdd.n1409 9.3005
R19263 vdd.n1411 vdd.n1228 9.3005
R19264 vdd.n1413 vdd.n1412 9.3005
R19265 vdd.n1414 vdd.n1227 9.3005
R19266 vdd.n1416 vdd.n1415 9.3005
R19267 vdd.n1192 vdd.n1191 9.3005
R19268 vdd.n1422 vdd.n1421 9.3005
R19269 vdd.n1321 vdd.n1320 9.3005
R19270 vdd.n1425 vdd.n1424 9.3005
R19271 vdd.n1181 vdd.n1180 9.3005
R19272 vdd.n1439 vdd.n1438 9.3005
R19273 vdd.n1440 vdd.n1179 9.3005
R19274 vdd.n1442 vdd.n1441 9.3005
R19275 vdd.n1170 vdd.n1169 9.3005
R19276 vdd.n1456 vdd.n1455 9.3005
R19277 vdd.n1457 vdd.n1168 9.3005
R19278 vdd.n1459 vdd.n1458 9.3005
R19279 vdd.n1159 vdd.n1158 9.3005
R19280 vdd.n1472 vdd.n1471 9.3005
R19281 vdd.n1473 vdd.n1157 9.3005
R19282 vdd.n1475 vdd.n1474 9.3005
R19283 vdd.n1147 vdd.n1146 9.3005
R19284 vdd.n1489 vdd.n1488 9.3005
R19285 vdd.n1490 vdd.n1145 9.3005
R19286 vdd.n1492 vdd.n1491 9.3005
R19287 vdd.n1136 vdd.n1135 9.3005
R19288 vdd.n1505 vdd.n1504 9.3005
R19289 vdd.n1506 vdd.n1134 9.3005
R19290 vdd.n1423 vdd.n1190 9.3005
R19291 vdd.n1726 vdd.n1725 9.3005
R19292 vdd.n1721 vdd.n1720 9.3005
R19293 vdd.n1732 vdd.n1731 9.3005
R19294 vdd.n1734 vdd.n1733 9.3005
R19295 vdd.n1717 vdd.n1716 9.3005
R19296 vdd.n1740 vdd.n1739 9.3005
R19297 vdd.n1742 vdd.n1741 9.3005
R19298 vdd.n1714 vdd.n1711 9.3005
R19299 vdd.n1749 vdd.n1748 9.3005
R19300 vdd.n1785 vdd.n1784 9.3005
R19301 vdd.n1780 vdd.n1779 9.3005
R19302 vdd.n1791 vdd.n1790 9.3005
R19303 vdd.n1793 vdd.n1792 9.3005
R19304 vdd.n1776 vdd.n1775 9.3005
R19305 vdd.n1799 vdd.n1798 9.3005
R19306 vdd.n1801 vdd.n1800 9.3005
R19307 vdd.n1773 vdd.n1770 9.3005
R19308 vdd.n1808 vdd.n1807 9.3005
R19309 vdd.n1624 vdd.n1623 9.3005
R19310 vdd.n1619 vdd.n1618 9.3005
R19311 vdd.n1630 vdd.n1629 9.3005
R19312 vdd.n1632 vdd.n1631 9.3005
R19313 vdd.n1615 vdd.n1614 9.3005
R19314 vdd.n1638 vdd.n1637 9.3005
R19315 vdd.n1640 vdd.n1639 9.3005
R19316 vdd.n1612 vdd.n1609 9.3005
R19317 vdd.n1647 vdd.n1646 9.3005
R19318 vdd.n1683 vdd.n1682 9.3005
R19319 vdd.n1678 vdd.n1677 9.3005
R19320 vdd.n1689 vdd.n1688 9.3005
R19321 vdd.n1691 vdd.n1690 9.3005
R19322 vdd.n1674 vdd.n1673 9.3005
R19323 vdd.n1697 vdd.n1696 9.3005
R19324 vdd.n1699 vdd.n1698 9.3005
R19325 vdd.n1671 vdd.n1668 9.3005
R19326 vdd.n1706 vdd.n1705 9.3005
R19327 vdd.n1523 vdd.n1522 9.3005
R19328 vdd.n1518 vdd.n1517 9.3005
R19329 vdd.n1529 vdd.n1528 9.3005
R19330 vdd.n1531 vdd.n1530 9.3005
R19331 vdd.n1514 vdd.n1513 9.3005
R19332 vdd.n1537 vdd.n1536 9.3005
R19333 vdd.n1539 vdd.n1538 9.3005
R19334 vdd.n1511 vdd.n1508 9.3005
R19335 vdd.n1546 vdd.n1545 9.3005
R19336 vdd.n1582 vdd.n1581 9.3005
R19337 vdd.n1577 vdd.n1576 9.3005
R19338 vdd.n1588 vdd.n1587 9.3005
R19339 vdd.n1590 vdd.n1589 9.3005
R19340 vdd.n1573 vdd.n1572 9.3005
R19341 vdd.n1596 vdd.n1595 9.3005
R19342 vdd.n1598 vdd.n1597 9.3005
R19343 vdd.n1570 vdd.n1567 9.3005
R19344 vdd.n1605 vdd.n1604 9.3005
R19345 vdd.n1461 vdd.t56 9.18308
R19346 vdd.n3331 vdd.t125 9.18308
R19347 vdd.n1155 vdd.t107 8.95635
R19348 vdd.n2329 vdd.t223 8.95635
R19349 vdd.n723 vdd.t216 8.95635
R19350 vdd.t71 vdd.n3385 8.95635
R19351 vdd.n312 vdd.n311 8.92171
R19352 vdd.n253 vdd.n252 8.92171
R19353 vdd.n210 vdd.n209 8.92171
R19354 vdd.n151 vdd.n150 8.92171
R19355 vdd.n109 vdd.n108 8.92171
R19356 vdd.n50 vdd.n49 8.92171
R19357 vdd.n1731 vdd.n1730 8.92171
R19358 vdd.n1790 vdd.n1789 8.92171
R19359 vdd.n1629 vdd.n1628 8.92171
R19360 vdd.n1688 vdd.n1687 8.92171
R19361 vdd.n1528 vdd.n1527 8.92171
R19362 vdd.n1587 vdd.n1586 8.92171
R19363 vdd.n231 vdd.n129 8.81535
R19364 vdd.n1709 vdd.n1607 8.81535
R19365 vdd.n1502 vdd.t79 8.72962
R19366 vdd.t68 vdd.n3394 8.72962
R19367 vdd.n1825 vdd.t128 8.50289
R19368 vdd.n3300 vdd.t73 8.50289
R19369 vdd.n28 vdd.n14 8.42249
R19370 vdd.n1851 vdd.t65 8.27616
R19371 vdd.t58 vdd.n656 8.27616
R19372 vdd.n3400 vdd.n3399 8.16225
R19373 vdd.n1813 vdd.n1812 8.16225
R19374 vdd.n308 vdd.n302 8.14595
R19375 vdd.n249 vdd.n243 8.14595
R19376 vdd.n206 vdd.n200 8.14595
R19377 vdd.n147 vdd.n141 8.14595
R19378 vdd.n105 vdd.n99 8.14595
R19379 vdd.n46 vdd.n40 8.14595
R19380 vdd.n1727 vdd.n1721 8.14595
R19381 vdd.n1786 vdd.n1780 8.14595
R19382 vdd.n1625 vdd.n1619 8.14595
R19383 vdd.n1684 vdd.n1678 8.14595
R19384 vdd.n1524 vdd.n1518 8.14595
R19385 vdd.n1583 vdd.n1577 8.14595
R19386 vdd.n2923 vdd.n849 8.11757
R19387 vdd.n2397 vdd.n2396 8.11757
R19388 vdd.n1098 vdd.t151 8.04943
R19389 vdd.n3256 vdd.t105 8.04943
R19390 vdd.n2375 vdd.n1043 7.70933
R19391 vdd.n2381 vdd.n1043 7.70933
R19392 vdd.n2387 vdd.n1037 7.70933
R19393 vdd.n2387 vdd.n1030 7.70933
R19394 vdd.n2393 vdd.n1030 7.70933
R19395 vdd.n2393 vdd.n1033 7.70933
R19396 vdd.n2400 vdd.n1018 7.70933
R19397 vdd.n2406 vdd.n1018 7.70933
R19398 vdd.n2412 vdd.n1012 7.70933
R19399 vdd.n2418 vdd.n1008 7.70933
R19400 vdd.n2424 vdd.n1002 7.70933
R19401 vdd.n2436 vdd.n989 7.70933
R19402 vdd.n2442 vdd.n983 7.70933
R19403 vdd.n2442 vdd.n976 7.70933
R19404 vdd.n2450 vdd.n976 7.70933
R19405 vdd.n2457 vdd.t292 7.70933
R19406 vdd.n2532 vdd.t292 7.70933
R19407 vdd.n2864 vdd.t200 7.70933
R19408 vdd.n2870 vdd.t200 7.70933
R19409 vdd.n2876 vdd.n897 7.70933
R19410 vdd.n2882 vdd.n897 7.70933
R19411 vdd.n2882 vdd.n900 7.70933
R19412 vdd.n2888 vdd.n893 7.70933
R19413 vdd.n2900 vdd.n880 7.70933
R19414 vdd.n2906 vdd.n874 7.70933
R19415 vdd.n2912 vdd.n870 7.70933
R19416 vdd.n2918 vdd.n857 7.70933
R19417 vdd.n2926 vdd.n857 7.70933
R19418 vdd.n2932 vdd.n851 7.70933
R19419 vdd.n2932 vdd.n843 7.70933
R19420 vdd.n2983 vdd.n843 7.70933
R19421 vdd.n2983 vdd.n846 7.70933
R19422 vdd.n2989 vdd.n805 7.70933
R19423 vdd.n3059 vdd.n805 7.70933
R19424 vdd.n307 vdd.n304 7.3702
R19425 vdd.n248 vdd.n245 7.3702
R19426 vdd.n205 vdd.n202 7.3702
R19427 vdd.n146 vdd.n143 7.3702
R19428 vdd.n104 vdd.n101 7.3702
R19429 vdd.n45 vdd.n42 7.3702
R19430 vdd.n1726 vdd.n1723 7.3702
R19431 vdd.n1785 vdd.n1782 7.3702
R19432 vdd.n1624 vdd.n1621 7.3702
R19433 vdd.n1683 vdd.n1680 7.3702
R19434 vdd.n1523 vdd.n1520 7.3702
R19435 vdd.n1582 vdd.n1579 7.3702
R19436 vdd.n1884 vdd.t21 7.1425
R19437 vdd.n679 vdd.t17 7.1425
R19438 vdd.n1358 vdd.n1357 6.98232
R19439 vdd.n2039 vdd.n2038 6.98232
R19440 vdd.n566 vdd.n565 6.98232
R19441 vdd.n3141 vdd.n3138 6.98232
R19442 vdd.t130 vdd.n1097 6.91577
R19443 vdd.n3264 vdd.t27 6.91577
R19444 vdd.n1843 vdd.t89 6.68904
R19445 vdd.n3280 vdd.t14 6.68904
R19446 vdd.t33 vdd.n1126 6.46231
R19447 vdd.n3308 vdd.t29 6.46231
R19448 vdd.n3400 vdd.n333 6.38151
R19449 vdd.n1812 vdd.n1811 6.38151
R19450 vdd.n1494 vdd.t62 6.23558
R19451 vdd.t100 vdd.n344 6.23558
R19452 vdd.t31 vdd.n1154 6.00885
R19453 vdd.n2412 vdd.t5 6.00885
R19454 vdd.n2912 vdd.t11 6.00885
R19455 vdd.n3379 vdd.t45 6.00885
R19456 vdd.n1033 vdd.t269 5.89549
R19457 vdd.t227 vdd.n851 5.89549
R19458 vdd.n308 vdd.n307 5.81868
R19459 vdd.n249 vdd.n248 5.81868
R19460 vdd.n206 vdd.n205 5.81868
R19461 vdd.n147 vdd.n146 5.81868
R19462 vdd.n105 vdd.n104 5.81868
R19463 vdd.n46 vdd.n45 5.81868
R19464 vdd.n1727 vdd.n1726 5.81868
R19465 vdd.n1786 vdd.n1785 5.81868
R19466 vdd.n1625 vdd.n1624 5.81868
R19467 vdd.n1684 vdd.n1683 5.81868
R19468 vdd.n1524 vdd.n1523 5.81868
R19469 vdd.n1583 vdd.n1582 5.81868
R19470 vdd.n1453 vdd.t19 5.78212
R19471 vdd.t212 vdd.n1037 5.78212
R19472 vdd.n2156 vdd.t251 5.78212
R19473 vdd.n2781 vdd.t259 5.78212
R19474 vdd.n846 vdd.t255 5.78212
R19475 vdd.n3370 vdd.t94 5.78212
R19476 vdd.n2540 vdd.n2539 5.77611
R19477 vdd.n2283 vdd.n2153 5.77611
R19478 vdd.n2794 vdd.n2793 5.77611
R19479 vdd.n3000 vdd.n2999 5.77611
R19480 vdd.n3064 vdd.n801 5.77611
R19481 vdd.n2704 vdd.n2644 5.77611
R19482 vdd.n2465 vdd.n967 5.77611
R19483 vdd.n2213 vdd.n2212 5.77611
R19484 vdd.n1320 vdd.n1319 5.62474
R19485 vdd.n2335 vdd.n2332 5.62474
R19486 vdd.n3351 vdd.n428 5.62474
R19487 vdd.n3225 vdd.n690 5.62474
R19488 vdd.n1177 vdd.t19 5.55539
R19489 vdd.t94 vdd.n3369 5.55539
R19490 vdd.t2 vdd.n989 5.44203
R19491 vdd.n893 vdd.t12 5.44203
R19492 vdd.n1469 vdd.t31 5.32866
R19493 vdd.t45 vdd.n3378 5.32866
R19494 vdd.n1485 vdd.t62 5.10193
R19495 vdd.t184 vdd.n1012 5.10193
R19496 vdd.n1002 vdd.t198 5.10193
R19497 vdd.t183 vdd.n880 5.10193
R19498 vdd.n870 vdd.t192 5.10193
R19499 vdd.n3387 vdd.t100 5.10193
R19500 vdd.n311 vdd.n302 5.04292
R19501 vdd.n252 vdd.n243 5.04292
R19502 vdd.n209 vdd.n200 5.04292
R19503 vdd.n150 vdd.n141 5.04292
R19504 vdd.n108 vdd.n99 5.04292
R19505 vdd.n49 vdd.n40 5.04292
R19506 vdd.n1730 vdd.n1721 5.04292
R19507 vdd.n1789 vdd.n1780 5.04292
R19508 vdd.n1628 vdd.n1619 5.04292
R19509 vdd.n1687 vdd.n1678 5.04292
R19510 vdd.n1527 vdd.n1518 5.04292
R19511 vdd.n1586 vdd.n1577 5.04292
R19512 vdd.n1817 vdd.t33 4.8752
R19513 vdd.t195 vdd.t206 4.8752
R19514 vdd.t182 vdd.t289 4.8752
R19515 vdd.t0 vdd.t179 4.8752
R19516 vdd.t185 vdd.t187 4.8752
R19517 vdd.t29 vdd.n340 4.8752
R19518 vdd.n2541 vdd.n2540 4.83952
R19519 vdd.n2153 vdd.n2149 4.83952
R19520 vdd.n2795 vdd.n2794 4.83952
R19521 vdd.n3001 vdd.n3000 4.83952
R19522 vdd.n801 vdd.n796 4.83952
R19523 vdd.n2701 vdd.n2644 4.83952
R19524 vdd.n2468 vdd.n967 4.83952
R19525 vdd.n2212 vdd.n2211 4.83952
R19526 vdd.n2007 vdd.n1065 4.74817
R19527 vdd.n2002 vdd.n1066 4.74817
R19528 vdd.n1904 vdd.n1901 4.74817
R19529 vdd.n2316 vdd.n1905 4.74817
R19530 vdd.n2318 vdd.n1904 4.74817
R19531 vdd.n2317 vdd.n2316 4.74817
R19532 vdd.n3218 vdd.n3217 4.74817
R19533 vdd.n3215 vdd.n3214 4.74817
R19534 vdd.n3215 vdd.n732 4.74817
R19535 vdd.n3217 vdd.n729 4.74817
R19536 vdd.n3100 vdd.n784 4.74817
R19537 vdd.n3096 vdd.n3094 4.74817
R19538 vdd.n3099 vdd.n3094 4.74817
R19539 vdd.n3103 vdd.n784 4.74817
R19540 vdd.n2003 vdd.n1065 4.74817
R19541 vdd.n1068 vdd.n1066 4.74817
R19542 vdd.n333 vdd.n332 4.7074
R19543 vdd.n231 vdd.n230 4.7074
R19544 vdd.n1811 vdd.n1810 4.7074
R19545 vdd.n1709 vdd.n1708 4.7074
R19546 vdd.n1120 vdd.t89 4.64847
R19547 vdd.n3289 vdd.t14 4.64847
R19548 vdd.n2418 vdd.t287 4.53511
R19549 vdd.n2906 vdd.t190 4.53511
R19550 vdd.n1859 vdd.t130 4.42174
R19551 vdd.t27 vdd.n655 4.42174
R19552 vdd.n2450 vdd.t6 4.30838
R19553 vdd.n2876 vdd.t176 4.30838
R19554 vdd.n312 vdd.n300 4.26717
R19555 vdd.n253 vdd.n241 4.26717
R19556 vdd.n210 vdd.n198 4.26717
R19557 vdd.n151 vdd.n139 4.26717
R19558 vdd.n109 vdd.n97 4.26717
R19559 vdd.n50 vdd.n38 4.26717
R19560 vdd.n1731 vdd.n1719 4.26717
R19561 vdd.n1790 vdd.n1778 4.26717
R19562 vdd.n1629 vdd.n1617 4.26717
R19563 vdd.n1688 vdd.n1676 4.26717
R19564 vdd.n1528 vdd.n1516 4.26717
R19565 vdd.n1587 vdd.n1575 4.26717
R19566 vdd.n1875 vdd.t21 4.19501
R19567 vdd.n3248 vdd.t17 4.19501
R19568 vdd.n333 vdd.n231 4.10845
R19569 vdd.n1811 vdd.n1709 4.10845
R19570 vdd.n289 vdd.t55 4.06363
R19571 vdd.n289 vdd.t117 4.06363
R19572 vdd.n287 vdd.t148 4.06363
R19573 vdd.n287 vdd.t166 4.06363
R19574 vdd.n285 vdd.t169 4.06363
R19575 vdd.n285 vdd.t64 4.06363
R19576 vdd.n283 vdd.t87 4.06363
R19577 vdd.n283 vdd.t160 4.06363
R19578 vdd.n281 vdd.t170 4.06363
R19579 vdd.n281 vdd.t86 4.06363
R19580 vdd.n279 vdd.t91 4.06363
R19581 vdd.n279 vdd.t93 4.06363
R19582 vdd.n277 vdd.t143 4.06363
R19583 vdd.n277 vdd.t16 4.06363
R19584 vdd.n275 vdd.t51 4.06363
R19585 vdd.n275 vdd.t116 4.06363
R19586 vdd.n273 vdd.t121 4.06363
R19587 vdd.n273 vdd.t150 4.06363
R19588 vdd.n187 vdd.t38 4.06363
R19589 vdd.n187 vdd.t95 4.06363
R19590 vdd.n185 vdd.t135 4.06363
R19591 vdd.n185 vdd.t153 4.06363
R19592 vdd.n183 vdd.t157 4.06363
R19593 vdd.n183 vdd.t40 4.06363
R19594 vdd.n181 vdd.t70 4.06363
R19595 vdd.n181 vdd.t156 4.06363
R19596 vdd.n179 vdd.t162 4.06363
R19597 vdd.n179 vdd.t69 4.06363
R19598 vdd.n177 vdd.t74 4.06363
R19599 vdd.n177 vdd.t76 4.06363
R19600 vdd.n175 vdd.t133 4.06363
R19601 vdd.n175 vdd.t15 4.06363
R19602 vdd.n173 vdd.t28 4.06363
R19603 vdd.n173 vdd.t96 4.06363
R19604 vdd.n171 vdd.t106 4.06363
R19605 vdd.n171 vdd.t136 4.06363
R19606 vdd.n86 vdd.t54 4.06363
R19607 vdd.n86 vdd.t141 4.06363
R19608 vdd.n84 vdd.t46 4.06363
R19609 vdd.n84 vdd.t126 4.06363
R19610 vdd.n82 vdd.t72 4.06363
R19611 vdd.n82 vdd.t154 4.06363
R19612 vdd.n80 vdd.t42 4.06363
R19613 vdd.n80 vdd.t101 4.06363
R19614 vdd.n78 vdd.t30 4.06363
R19615 vdd.n78 vdd.t77 4.06363
R19616 vdd.n76 vdd.t167 4.06363
R19617 vdd.n76 vdd.t140 4.06363
R19618 vdd.n74 vdd.t146 4.06363
R19619 vdd.n74 vdd.t88 4.06363
R19620 vdd.n72 vdd.t171 4.06363
R19621 vdd.n72 vdd.t59 4.06363
R19622 vdd.n70 vdd.t158 4.06363
R19623 vdd.n70 vdd.t98 4.06363
R19624 vdd.n1751 vdd.t53 4.06363
R19625 vdd.n1751 vdd.t165 4.06363
R19626 vdd.n1753 vdd.t159 4.06363
R19627 vdd.n1753 vdd.t142 4.06363
R19628 vdd.n1755 vdd.t111 4.06363
R19629 vdd.n1755 vdd.t49 4.06363
R19630 vdd.n1757 vdd.t173 4.06363
R19631 vdd.n1757 vdd.t139 4.06363
R19632 vdd.n1759 vdd.t115 4.06363
R19633 vdd.n1759 vdd.t85 4.06363
R19634 vdd.n1761 vdd.t81 4.06363
R19635 vdd.n1761 vdd.t137 4.06363
R19636 vdd.n1763 vdd.t122 4.06363
R19637 vdd.n1763 vdd.t120 4.06363
R19638 vdd.n1765 vdd.t78 4.06363
R19639 vdd.n1765 vdd.t52 4.06363
R19640 vdd.n1767 vdd.t48 4.06363
R19641 vdd.n1767 vdd.t118 4.06363
R19642 vdd.n1649 vdd.t36 4.06363
R19643 vdd.n1649 vdd.t152 4.06363
R19644 vdd.n1651 vdd.t145 4.06363
R19645 vdd.n1651 vdd.t131 4.06363
R19646 vdd.n1653 vdd.t92 4.06363
R19647 vdd.n1653 vdd.t24 4.06363
R19648 vdd.n1655 vdd.t163 4.06363
R19649 vdd.n1655 vdd.t129 4.06363
R19650 vdd.n1657 vdd.t123 4.06363
R19651 vdd.n1657 vdd.t67 4.06363
R19652 vdd.n1659 vdd.t63 4.06363
R19653 vdd.n1659 vdd.t124 4.06363
R19654 vdd.n1661 vdd.t110 4.06363
R19655 vdd.n1661 vdd.t108 4.06363
R19656 vdd.n1663 vdd.t57 4.06363
R19657 vdd.n1663 vdd.t32 4.06363
R19658 vdd.n1665 vdd.t20 4.06363
R19659 vdd.n1665 vdd.t103 4.06363
R19660 vdd.n1548 vdd.t99 4.06363
R19661 vdd.n1548 vdd.t161 4.06363
R19662 vdd.n1550 vdd.t66 4.06363
R19663 vdd.n1550 vdd.t138 4.06363
R19664 vdd.n1552 vdd.t90 4.06363
R19665 vdd.n1552 vdd.t147 4.06363
R19666 vdd.n1554 vdd.t113 4.06363
R19667 vdd.n1554 vdd.t168 4.06363
R19668 vdd.n1556 vdd.t80 4.06363
R19669 vdd.n1556 vdd.t34 4.06363
R19670 vdd.n1558 vdd.t102 4.06363
R19671 vdd.n1558 vdd.t44 4.06363
R19672 vdd.n1560 vdd.t155 4.06363
R19673 vdd.n1560 vdd.t172 4.06363
R19674 vdd.n1562 vdd.t127 4.06363
R19675 vdd.n1562 vdd.t47 4.06363
R19676 vdd.n1564 vdd.t114 4.06363
R19677 vdd.n1564 vdd.t61 4.06363
R19678 vdd.n26 vdd.t203 3.9605
R19679 vdd.n26 vdd.t10 3.9605
R19680 vdd.n23 vdd.t181 3.9605
R19681 vdd.n23 vdd.t202 3.9605
R19682 vdd.n21 vdd.t180 3.9605
R19683 vdd.n21 vdd.t189 3.9605
R19684 vdd.n20 vdd.t210 3.9605
R19685 vdd.n20 vdd.t9 3.9605
R19686 vdd.n15 vdd.t291 3.9605
R19687 vdd.n15 vdd.t188 3.9605
R19688 vdd.n16 vdd.t209 3.9605
R19689 vdd.n16 vdd.t8 3.9605
R19690 vdd.n18 vdd.t174 3.9605
R19691 vdd.n18 vdd.t208 3.9605
R19692 vdd.n25 vdd.t175 3.9605
R19693 vdd.n25 vdd.t199 3.9605
R19694 vdd.n7 vdd.t186 3.61217
R19695 vdd.n7 vdd.t191 3.61217
R19696 vdd.n8 vdd.t1 3.61217
R19697 vdd.n8 vdd.t13 3.61217
R19698 vdd.n10 vdd.t201 3.61217
R19699 vdd.n10 vdd.t177 3.61217
R19700 vdd.n12 vdd.t295 3.61217
R19701 vdd.n12 vdd.t194 3.61217
R19702 vdd.n5 vdd.t205 3.61217
R19703 vdd.n5 vdd.t197 3.61217
R19704 vdd.n3 vdd.t7 3.61217
R19705 vdd.n3 vdd.t293 3.61217
R19706 vdd.n1 vdd.t3 3.61217
R19707 vdd.n1 vdd.t290 3.61217
R19708 vdd.n0 vdd.t288 3.61217
R19709 vdd.n0 vdd.t207 3.61217
R19710 vdd.n316 vdd.n315 3.49141
R19711 vdd.n257 vdd.n256 3.49141
R19712 vdd.n214 vdd.n213 3.49141
R19713 vdd.n155 vdd.n154 3.49141
R19714 vdd.n113 vdd.n112 3.49141
R19715 vdd.n54 vdd.n53 3.49141
R19716 vdd.n1735 vdd.n1734 3.49141
R19717 vdd.n1794 vdd.n1793 3.49141
R19718 vdd.n1633 vdd.n1632 3.49141
R19719 vdd.n1692 vdd.n1691 3.49141
R19720 vdd.n1532 vdd.n1531 3.49141
R19721 vdd.n1591 vdd.n1590 3.49141
R19722 vdd.n2156 vdd.t6 3.40145
R19723 vdd.n2604 vdd.t204 3.40145
R19724 vdd.n2857 vdd.t193 3.40145
R19725 vdd.n2781 vdd.t176 3.40145
R19726 vdd.n1876 vdd.t151 3.28809
R19727 vdd.n3247 vdd.t105 3.28809
R19728 vdd.n2257 vdd.t287 3.17472
R19729 vdd.n2760 vdd.t190 3.17472
R19730 vdd.t65 vdd.n1104 3.06136
R19731 vdd.n3272 vdd.t58 3.06136
R19732 vdd.n1834 vdd.t128 2.83463
R19733 vdd.n644 vdd.t73 2.83463
R19734 vdd.n319 vdd.n298 2.71565
R19735 vdd.n260 vdd.n239 2.71565
R19736 vdd.n217 vdd.n196 2.71565
R19737 vdd.n158 vdd.n137 2.71565
R19738 vdd.n116 vdd.n95 2.71565
R19739 vdd.n57 vdd.n36 2.71565
R19740 vdd.n1738 vdd.n1717 2.71565
R19741 vdd.n1797 vdd.n1776 2.71565
R19742 vdd.n1636 vdd.n1615 2.71565
R19743 vdd.n1695 vdd.n1674 2.71565
R19744 vdd.n1535 vdd.n1514 2.71565
R19745 vdd.n1594 vdd.n1573 2.71565
R19746 vdd.t79 vdd.n1132 2.6079
R19747 vdd.n2406 vdd.t184 2.6079
R19748 vdd.n2430 vdd.t198 2.6079
R19749 vdd.n2894 vdd.t183 2.6079
R19750 vdd.n2918 vdd.t192 2.6079
R19751 vdd.n3395 vdd.t68 2.6079
R19752 vdd.n2924 vdd.n2923 2.49806
R19753 vdd.n2398 vdd.n2397 2.49806
R19754 vdd.n306 vdd.n305 2.4129
R19755 vdd.n247 vdd.n246 2.4129
R19756 vdd.n204 vdd.n203 2.4129
R19757 vdd.n145 vdd.n144 2.4129
R19758 vdd.n103 vdd.n102 2.4129
R19759 vdd.n44 vdd.n43 2.4129
R19760 vdd.n1725 vdd.n1724 2.4129
R19761 vdd.n1784 vdd.n1783 2.4129
R19762 vdd.n1623 vdd.n1622 2.4129
R19763 vdd.n1682 vdd.n1681 2.4129
R19764 vdd.n1522 vdd.n1521 2.4129
R19765 vdd.n1581 vdd.n1580 2.4129
R19766 vdd.n1486 vdd.t107 2.38117
R19767 vdd.n1894 vdd.t223 2.38117
R19768 vdd.n3231 vdd.t216 2.38117
R19769 vdd.n3386 vdd.t71 2.38117
R19770 vdd.n2315 vdd.n1904 2.27742
R19771 vdd.n2316 vdd.n2315 2.27742
R19772 vdd.n3216 vdd.n3215 2.27742
R19773 vdd.n3217 vdd.n3216 2.27742
R19774 vdd.n3094 vdd.n3093 2.27742
R19775 vdd.n3093 vdd.n784 2.27742
R19776 vdd.n2338 vdd.n1065 2.27742
R19777 vdd.n2338 vdd.n1066 2.27742
R19778 vdd.n2430 vdd.t2 2.2678
R19779 vdd.n2894 vdd.t12 2.2678
R19780 vdd.t56 vdd.n1161 2.15444
R19781 vdd.n3377 vdd.t125 2.15444
R19782 vdd.t289 vdd.n983 2.04107
R19783 vdd.n900 vdd.t0 2.04107
R19784 vdd.n320 vdd.n296 1.93989
R19785 vdd.n261 vdd.n237 1.93989
R19786 vdd.n218 vdd.n194 1.93989
R19787 vdd.n159 vdd.n135 1.93989
R19788 vdd.n117 vdd.n93 1.93989
R19789 vdd.n58 vdd.n34 1.93989
R19790 vdd.n1739 vdd.n1715 1.93989
R19791 vdd.n1798 vdd.n1774 1.93989
R19792 vdd.n1637 vdd.n1613 1.93989
R19793 vdd.n1696 vdd.n1672 1.93989
R19794 vdd.n1536 vdd.n1512 1.93989
R19795 vdd.n1595 vdd.n1571 1.93989
R19796 vdd.n1444 vdd.t25 1.92771
R19797 vdd.n2381 vdd.t212 1.92771
R19798 vdd.n2457 vdd.t251 1.92771
R19799 vdd.n2870 vdd.t259 1.92771
R19800 vdd.n2989 vdd.t255 1.92771
R19801 vdd.t82 vdd.n375 1.92771
R19802 vdd.n1452 vdd.t60 1.70098
R19803 vdd.n2257 vdd.t5 1.70098
R19804 vdd.n1008 vdd.t195 1.70098
R19805 vdd.t187 vdd.n874 1.70098
R19806 vdd.n2760 vdd.t11 1.70098
R19807 vdd.n3371 vdd.t37 1.70098
R19808 vdd.n1477 vdd.t109 1.47425
R19809 vdd.n361 vdd.t39 1.47425
R19810 vdd.n1143 vdd.t43 1.24752
R19811 vdd.t41 vdd.n3393 1.24752
R19812 vdd.n331 vdd.n291 1.16414
R19813 vdd.n324 vdd.n323 1.16414
R19814 vdd.n272 vdd.n232 1.16414
R19815 vdd.n265 vdd.n264 1.16414
R19816 vdd.n229 vdd.n189 1.16414
R19817 vdd.n222 vdd.n221 1.16414
R19818 vdd.n170 vdd.n130 1.16414
R19819 vdd.n163 vdd.n162 1.16414
R19820 vdd.n128 vdd.n88 1.16414
R19821 vdd.n121 vdd.n120 1.16414
R19822 vdd.n69 vdd.n29 1.16414
R19823 vdd.n62 vdd.n61 1.16414
R19824 vdd.n1750 vdd.n1710 1.16414
R19825 vdd.n1743 vdd.n1742 1.16414
R19826 vdd.n1809 vdd.n1769 1.16414
R19827 vdd.n1802 vdd.n1801 1.16414
R19828 vdd.n1648 vdd.n1608 1.16414
R19829 vdd.n1641 vdd.n1640 1.16414
R19830 vdd.n1707 vdd.n1667 1.16414
R19831 vdd.n1700 vdd.n1699 1.16414
R19832 vdd.n1547 vdd.n1507 1.16414
R19833 vdd.n1540 vdd.n1539 1.16414
R19834 vdd.n1606 vdd.n1566 1.16414
R19835 vdd.n1599 vdd.n1598 1.16414
R19836 vdd.n2424 vdd.t206 1.13415
R19837 vdd.n2900 vdd.t185 1.13415
R19838 vdd.n1826 vdd.t112 1.02079
R19839 vdd.t269 vdd.t4 1.02079
R19840 vdd.t178 vdd.t227 1.02079
R19841 vdd.t75 vdd.n633 1.02079
R19842 vdd.n1323 vdd.n1319 0.970197
R19843 vdd.n2336 vdd.n2335 0.970197
R19844 vdd.n618 vdd.n428 0.970197
R19845 vdd.n3095 vdd.n690 0.970197
R19846 vdd.n1812 vdd.n28 0.90431
R19847 vdd vdd.n3400 0.896477
R19848 vdd.n1842 vdd.t23 0.794056
R19849 vdd.n2400 vdd.t4 0.794056
R19850 vdd.n2436 vdd.t182 0.794056
R19851 vdd.n2888 vdd.t179 0.794056
R19852 vdd.n2926 vdd.t178 0.794056
R19853 vdd.n3281 vdd.t132 0.794056
R19854 vdd.n1867 vdd.t35 0.567326
R19855 vdd.t97 vdd.n662 0.567326
R19856 vdd.n2326 vdd.n2325 0.530988
R19857 vdd.n726 vdd.n682 0.530988
R19858 vdd.n464 vdd.n391 0.530988
R19859 vdd.n3350 vdd.n3349 0.530988
R19860 vdd.n3227 vdd.n3226 0.530988
R19861 vdd.n1889 vdd.n1067 0.530988
R19862 vdd.n1321 vdd.n1186 0.530988
R19863 vdd.n1423 vdd.n1422 0.530988
R19864 vdd.n4 vdd.n2 0.459552
R19865 vdd.n11 vdd.n9 0.459552
R19866 vdd.n329 vdd.n328 0.388379
R19867 vdd.n295 vdd.n293 0.388379
R19868 vdd.n270 vdd.n269 0.388379
R19869 vdd.n236 vdd.n234 0.388379
R19870 vdd.n227 vdd.n226 0.388379
R19871 vdd.n193 vdd.n191 0.388379
R19872 vdd.n168 vdd.n167 0.388379
R19873 vdd.n134 vdd.n132 0.388379
R19874 vdd.n126 vdd.n125 0.388379
R19875 vdd.n92 vdd.n90 0.388379
R19876 vdd.n67 vdd.n66 0.388379
R19877 vdd.n33 vdd.n31 0.388379
R19878 vdd.n1748 vdd.n1747 0.388379
R19879 vdd.n1714 vdd.n1712 0.388379
R19880 vdd.n1807 vdd.n1806 0.388379
R19881 vdd.n1773 vdd.n1771 0.388379
R19882 vdd.n1646 vdd.n1645 0.388379
R19883 vdd.n1612 vdd.n1610 0.388379
R19884 vdd.n1705 vdd.n1704 0.388379
R19885 vdd.n1671 vdd.n1669 0.388379
R19886 vdd.n1545 vdd.n1544 0.388379
R19887 vdd.n1511 vdd.n1509 0.388379
R19888 vdd.n1604 vdd.n1603 0.388379
R19889 vdd.n1570 vdd.n1568 0.388379
R19890 vdd.n19 vdd.n17 0.387128
R19891 vdd.n24 vdd.n22 0.387128
R19892 vdd.n6 vdd.n4 0.358259
R19893 vdd.n13 vdd.n11 0.358259
R19894 vdd.n276 vdd.n274 0.358259
R19895 vdd.n278 vdd.n276 0.358259
R19896 vdd.n280 vdd.n278 0.358259
R19897 vdd.n282 vdd.n280 0.358259
R19898 vdd.n284 vdd.n282 0.358259
R19899 vdd.n286 vdd.n284 0.358259
R19900 vdd.n288 vdd.n286 0.358259
R19901 vdd.n290 vdd.n288 0.358259
R19902 vdd.n332 vdd.n290 0.358259
R19903 vdd.n174 vdd.n172 0.358259
R19904 vdd.n176 vdd.n174 0.358259
R19905 vdd.n178 vdd.n176 0.358259
R19906 vdd.n180 vdd.n178 0.358259
R19907 vdd.n182 vdd.n180 0.358259
R19908 vdd.n184 vdd.n182 0.358259
R19909 vdd.n186 vdd.n184 0.358259
R19910 vdd.n188 vdd.n186 0.358259
R19911 vdd.n230 vdd.n188 0.358259
R19912 vdd.n73 vdd.n71 0.358259
R19913 vdd.n75 vdd.n73 0.358259
R19914 vdd.n77 vdd.n75 0.358259
R19915 vdd.n79 vdd.n77 0.358259
R19916 vdd.n81 vdd.n79 0.358259
R19917 vdd.n83 vdd.n81 0.358259
R19918 vdd.n85 vdd.n83 0.358259
R19919 vdd.n87 vdd.n85 0.358259
R19920 vdd.n129 vdd.n87 0.358259
R19921 vdd.n1810 vdd.n1768 0.358259
R19922 vdd.n1768 vdd.n1766 0.358259
R19923 vdd.n1766 vdd.n1764 0.358259
R19924 vdd.n1764 vdd.n1762 0.358259
R19925 vdd.n1762 vdd.n1760 0.358259
R19926 vdd.n1760 vdd.n1758 0.358259
R19927 vdd.n1758 vdd.n1756 0.358259
R19928 vdd.n1756 vdd.n1754 0.358259
R19929 vdd.n1754 vdd.n1752 0.358259
R19930 vdd.n1708 vdd.n1666 0.358259
R19931 vdd.n1666 vdd.n1664 0.358259
R19932 vdd.n1664 vdd.n1662 0.358259
R19933 vdd.n1662 vdd.n1660 0.358259
R19934 vdd.n1660 vdd.n1658 0.358259
R19935 vdd.n1658 vdd.n1656 0.358259
R19936 vdd.n1656 vdd.n1654 0.358259
R19937 vdd.n1654 vdd.n1652 0.358259
R19938 vdd.n1652 vdd.n1650 0.358259
R19939 vdd.n1607 vdd.n1565 0.358259
R19940 vdd.n1565 vdd.n1563 0.358259
R19941 vdd.n1563 vdd.n1561 0.358259
R19942 vdd.n1561 vdd.n1559 0.358259
R19943 vdd.n1559 vdd.n1557 0.358259
R19944 vdd.n1557 vdd.n1555 0.358259
R19945 vdd.n1555 vdd.n1553 0.358259
R19946 vdd.n1553 vdd.n1551 0.358259
R19947 vdd.n1551 vdd.n1549 0.358259
R19948 vdd.n14 vdd.n6 0.334552
R19949 vdd.n14 vdd.n13 0.334552
R19950 vdd.n27 vdd.n19 0.21707
R19951 vdd.n27 vdd.n24 0.21707
R19952 vdd.n330 vdd.n292 0.155672
R19953 vdd.n322 vdd.n292 0.155672
R19954 vdd.n322 vdd.n321 0.155672
R19955 vdd.n321 vdd.n297 0.155672
R19956 vdd.n314 vdd.n297 0.155672
R19957 vdd.n314 vdd.n313 0.155672
R19958 vdd.n313 vdd.n301 0.155672
R19959 vdd.n306 vdd.n301 0.155672
R19960 vdd.n271 vdd.n233 0.155672
R19961 vdd.n263 vdd.n233 0.155672
R19962 vdd.n263 vdd.n262 0.155672
R19963 vdd.n262 vdd.n238 0.155672
R19964 vdd.n255 vdd.n238 0.155672
R19965 vdd.n255 vdd.n254 0.155672
R19966 vdd.n254 vdd.n242 0.155672
R19967 vdd.n247 vdd.n242 0.155672
R19968 vdd.n228 vdd.n190 0.155672
R19969 vdd.n220 vdd.n190 0.155672
R19970 vdd.n220 vdd.n219 0.155672
R19971 vdd.n219 vdd.n195 0.155672
R19972 vdd.n212 vdd.n195 0.155672
R19973 vdd.n212 vdd.n211 0.155672
R19974 vdd.n211 vdd.n199 0.155672
R19975 vdd.n204 vdd.n199 0.155672
R19976 vdd.n169 vdd.n131 0.155672
R19977 vdd.n161 vdd.n131 0.155672
R19978 vdd.n161 vdd.n160 0.155672
R19979 vdd.n160 vdd.n136 0.155672
R19980 vdd.n153 vdd.n136 0.155672
R19981 vdd.n153 vdd.n152 0.155672
R19982 vdd.n152 vdd.n140 0.155672
R19983 vdd.n145 vdd.n140 0.155672
R19984 vdd.n127 vdd.n89 0.155672
R19985 vdd.n119 vdd.n89 0.155672
R19986 vdd.n119 vdd.n118 0.155672
R19987 vdd.n118 vdd.n94 0.155672
R19988 vdd.n111 vdd.n94 0.155672
R19989 vdd.n111 vdd.n110 0.155672
R19990 vdd.n110 vdd.n98 0.155672
R19991 vdd.n103 vdd.n98 0.155672
R19992 vdd.n68 vdd.n30 0.155672
R19993 vdd.n60 vdd.n30 0.155672
R19994 vdd.n60 vdd.n59 0.155672
R19995 vdd.n59 vdd.n35 0.155672
R19996 vdd.n52 vdd.n35 0.155672
R19997 vdd.n52 vdd.n51 0.155672
R19998 vdd.n51 vdd.n39 0.155672
R19999 vdd.n44 vdd.n39 0.155672
R20000 vdd.n1749 vdd.n1711 0.155672
R20001 vdd.n1741 vdd.n1711 0.155672
R20002 vdd.n1741 vdd.n1740 0.155672
R20003 vdd.n1740 vdd.n1716 0.155672
R20004 vdd.n1733 vdd.n1716 0.155672
R20005 vdd.n1733 vdd.n1732 0.155672
R20006 vdd.n1732 vdd.n1720 0.155672
R20007 vdd.n1725 vdd.n1720 0.155672
R20008 vdd.n1808 vdd.n1770 0.155672
R20009 vdd.n1800 vdd.n1770 0.155672
R20010 vdd.n1800 vdd.n1799 0.155672
R20011 vdd.n1799 vdd.n1775 0.155672
R20012 vdd.n1792 vdd.n1775 0.155672
R20013 vdd.n1792 vdd.n1791 0.155672
R20014 vdd.n1791 vdd.n1779 0.155672
R20015 vdd.n1784 vdd.n1779 0.155672
R20016 vdd.n1647 vdd.n1609 0.155672
R20017 vdd.n1639 vdd.n1609 0.155672
R20018 vdd.n1639 vdd.n1638 0.155672
R20019 vdd.n1638 vdd.n1614 0.155672
R20020 vdd.n1631 vdd.n1614 0.155672
R20021 vdd.n1631 vdd.n1630 0.155672
R20022 vdd.n1630 vdd.n1618 0.155672
R20023 vdd.n1623 vdd.n1618 0.155672
R20024 vdd.n1706 vdd.n1668 0.155672
R20025 vdd.n1698 vdd.n1668 0.155672
R20026 vdd.n1698 vdd.n1697 0.155672
R20027 vdd.n1697 vdd.n1673 0.155672
R20028 vdd.n1690 vdd.n1673 0.155672
R20029 vdd.n1690 vdd.n1689 0.155672
R20030 vdd.n1689 vdd.n1677 0.155672
R20031 vdd.n1682 vdd.n1677 0.155672
R20032 vdd.n1546 vdd.n1508 0.155672
R20033 vdd.n1538 vdd.n1508 0.155672
R20034 vdd.n1538 vdd.n1537 0.155672
R20035 vdd.n1537 vdd.n1513 0.155672
R20036 vdd.n1530 vdd.n1513 0.155672
R20037 vdd.n1530 vdd.n1529 0.155672
R20038 vdd.n1529 vdd.n1517 0.155672
R20039 vdd.n1522 vdd.n1517 0.155672
R20040 vdd.n1605 vdd.n1567 0.155672
R20041 vdd.n1597 vdd.n1567 0.155672
R20042 vdd.n1597 vdd.n1596 0.155672
R20043 vdd.n1596 vdd.n1572 0.155672
R20044 vdd.n1589 vdd.n1572 0.155672
R20045 vdd.n1589 vdd.n1588 0.155672
R20046 vdd.n1588 vdd.n1576 0.155672
R20047 vdd.n1581 vdd.n1576 0.155672
R20048 vdd.n2101 vdd.n1906 0.152939
R20049 vdd.n1912 vdd.n1906 0.152939
R20050 vdd.n1913 vdd.n1912 0.152939
R20051 vdd.n1914 vdd.n1913 0.152939
R20052 vdd.n1915 vdd.n1914 0.152939
R20053 vdd.n1919 vdd.n1915 0.152939
R20054 vdd.n1920 vdd.n1919 0.152939
R20055 vdd.n1921 vdd.n1920 0.152939
R20056 vdd.n1922 vdd.n1921 0.152939
R20057 vdd.n1926 vdd.n1922 0.152939
R20058 vdd.n1927 vdd.n1926 0.152939
R20059 vdd.n1928 vdd.n1927 0.152939
R20060 vdd.n2076 vdd.n1928 0.152939
R20061 vdd.n2076 vdd.n2075 0.152939
R20062 vdd.n2075 vdd.n2074 0.152939
R20063 vdd.n2074 vdd.n1934 0.152939
R20064 vdd.n1939 vdd.n1934 0.152939
R20065 vdd.n1940 vdd.n1939 0.152939
R20066 vdd.n1941 vdd.n1940 0.152939
R20067 vdd.n1945 vdd.n1941 0.152939
R20068 vdd.n1946 vdd.n1945 0.152939
R20069 vdd.n1947 vdd.n1946 0.152939
R20070 vdd.n1948 vdd.n1947 0.152939
R20071 vdd.n1952 vdd.n1948 0.152939
R20072 vdd.n1953 vdd.n1952 0.152939
R20073 vdd.n1954 vdd.n1953 0.152939
R20074 vdd.n1955 vdd.n1954 0.152939
R20075 vdd.n1959 vdd.n1955 0.152939
R20076 vdd.n1960 vdd.n1959 0.152939
R20077 vdd.n1961 vdd.n1960 0.152939
R20078 vdd.n1962 vdd.n1961 0.152939
R20079 vdd.n1966 vdd.n1962 0.152939
R20080 vdd.n1967 vdd.n1966 0.152939
R20081 vdd.n1968 vdd.n1967 0.152939
R20082 vdd.n2037 vdd.n1968 0.152939
R20083 vdd.n2037 vdd.n2036 0.152939
R20084 vdd.n2036 vdd.n2035 0.152939
R20085 vdd.n2035 vdd.n1974 0.152939
R20086 vdd.n1979 vdd.n1974 0.152939
R20087 vdd.n1980 vdd.n1979 0.152939
R20088 vdd.n1981 vdd.n1980 0.152939
R20089 vdd.n1985 vdd.n1981 0.152939
R20090 vdd.n1986 vdd.n1985 0.152939
R20091 vdd.n1987 vdd.n1986 0.152939
R20092 vdd.n1988 vdd.n1987 0.152939
R20093 vdd.n1992 vdd.n1988 0.152939
R20094 vdd.n1993 vdd.n1992 0.152939
R20095 vdd.n1994 vdd.n1993 0.152939
R20096 vdd.n1995 vdd.n1994 0.152939
R20097 vdd.n1996 vdd.n1995 0.152939
R20098 vdd.n1996 vdd.n1064 0.152939
R20099 vdd.n2325 vdd.n1900 0.152939
R20100 vdd.n1814 vdd.n1123 0.152939
R20101 vdd.n1829 vdd.n1123 0.152939
R20102 vdd.n1830 vdd.n1829 0.152939
R20103 vdd.n1831 vdd.n1830 0.152939
R20104 vdd.n1831 vdd.n1112 0.152939
R20105 vdd.n1846 vdd.n1112 0.152939
R20106 vdd.n1847 vdd.n1846 0.152939
R20107 vdd.n1848 vdd.n1847 0.152939
R20108 vdd.n1848 vdd.n1101 0.152939
R20109 vdd.n1862 vdd.n1101 0.152939
R20110 vdd.n1863 vdd.n1862 0.152939
R20111 vdd.n1864 vdd.n1863 0.152939
R20112 vdd.n1864 vdd.n1089 0.152939
R20113 vdd.n1879 vdd.n1089 0.152939
R20114 vdd.n1880 vdd.n1879 0.152939
R20115 vdd.n1881 vdd.n1880 0.152939
R20116 vdd.n1881 vdd.n1077 0.152939
R20117 vdd.n1898 vdd.n1077 0.152939
R20118 vdd.n1899 vdd.n1898 0.152939
R20119 vdd.n2326 vdd.n1899 0.152939
R20120 vdd.n735 vdd.n730 0.152939
R20121 vdd.n736 vdd.n735 0.152939
R20122 vdd.n737 vdd.n736 0.152939
R20123 vdd.n738 vdd.n737 0.152939
R20124 vdd.n739 vdd.n738 0.152939
R20125 vdd.n740 vdd.n739 0.152939
R20126 vdd.n741 vdd.n740 0.152939
R20127 vdd.n742 vdd.n741 0.152939
R20128 vdd.n743 vdd.n742 0.152939
R20129 vdd.n744 vdd.n743 0.152939
R20130 vdd.n745 vdd.n744 0.152939
R20131 vdd.n746 vdd.n745 0.152939
R20132 vdd.n3183 vdd.n746 0.152939
R20133 vdd.n3183 vdd.n3182 0.152939
R20134 vdd.n3182 vdd.n3181 0.152939
R20135 vdd.n3181 vdd.n748 0.152939
R20136 vdd.n749 vdd.n748 0.152939
R20137 vdd.n750 vdd.n749 0.152939
R20138 vdd.n751 vdd.n750 0.152939
R20139 vdd.n752 vdd.n751 0.152939
R20140 vdd.n753 vdd.n752 0.152939
R20141 vdd.n754 vdd.n753 0.152939
R20142 vdd.n755 vdd.n754 0.152939
R20143 vdd.n756 vdd.n755 0.152939
R20144 vdd.n757 vdd.n756 0.152939
R20145 vdd.n758 vdd.n757 0.152939
R20146 vdd.n759 vdd.n758 0.152939
R20147 vdd.n760 vdd.n759 0.152939
R20148 vdd.n761 vdd.n760 0.152939
R20149 vdd.n762 vdd.n761 0.152939
R20150 vdd.n763 vdd.n762 0.152939
R20151 vdd.n764 vdd.n763 0.152939
R20152 vdd.n765 vdd.n764 0.152939
R20153 vdd.n766 vdd.n765 0.152939
R20154 vdd.n3137 vdd.n766 0.152939
R20155 vdd.n3137 vdd.n3136 0.152939
R20156 vdd.n3136 vdd.n3135 0.152939
R20157 vdd.n3135 vdd.n770 0.152939
R20158 vdd.n771 vdd.n770 0.152939
R20159 vdd.n772 vdd.n771 0.152939
R20160 vdd.n773 vdd.n772 0.152939
R20161 vdd.n774 vdd.n773 0.152939
R20162 vdd.n775 vdd.n774 0.152939
R20163 vdd.n776 vdd.n775 0.152939
R20164 vdd.n777 vdd.n776 0.152939
R20165 vdd.n778 vdd.n777 0.152939
R20166 vdd.n779 vdd.n778 0.152939
R20167 vdd.n780 vdd.n779 0.152939
R20168 vdd.n781 vdd.n780 0.152939
R20169 vdd.n782 vdd.n781 0.152939
R20170 vdd.n783 vdd.n782 0.152939
R20171 vdd.n727 vdd.n726 0.152939
R20172 vdd.n3234 vdd.n682 0.152939
R20173 vdd.n3235 vdd.n3234 0.152939
R20174 vdd.n3236 vdd.n3235 0.152939
R20175 vdd.n3236 vdd.n670 0.152939
R20176 vdd.n3251 vdd.n670 0.152939
R20177 vdd.n3252 vdd.n3251 0.152939
R20178 vdd.n3253 vdd.n3252 0.152939
R20179 vdd.n3253 vdd.n659 0.152939
R20180 vdd.n3267 vdd.n659 0.152939
R20181 vdd.n3268 vdd.n3267 0.152939
R20182 vdd.n3269 vdd.n3268 0.152939
R20183 vdd.n3269 vdd.n647 0.152939
R20184 vdd.n3284 vdd.n647 0.152939
R20185 vdd.n3285 vdd.n3284 0.152939
R20186 vdd.n3286 vdd.n3285 0.152939
R20187 vdd.n3286 vdd.n636 0.152939
R20188 vdd.n3303 vdd.n636 0.152939
R20189 vdd.n3304 vdd.n3303 0.152939
R20190 vdd.n3305 vdd.n3304 0.152939
R20191 vdd.n3305 vdd.n334 0.152939
R20192 vdd.n3398 vdd.n335 0.152939
R20193 vdd.n346 vdd.n335 0.152939
R20194 vdd.n347 vdd.n346 0.152939
R20195 vdd.n348 vdd.n347 0.152939
R20196 vdd.n355 vdd.n348 0.152939
R20197 vdd.n356 vdd.n355 0.152939
R20198 vdd.n357 vdd.n356 0.152939
R20199 vdd.n358 vdd.n357 0.152939
R20200 vdd.n366 vdd.n358 0.152939
R20201 vdd.n367 vdd.n366 0.152939
R20202 vdd.n368 vdd.n367 0.152939
R20203 vdd.n369 vdd.n368 0.152939
R20204 vdd.n377 vdd.n369 0.152939
R20205 vdd.n378 vdd.n377 0.152939
R20206 vdd.n379 vdd.n378 0.152939
R20207 vdd.n380 vdd.n379 0.152939
R20208 vdd.n388 vdd.n380 0.152939
R20209 vdd.n389 vdd.n388 0.152939
R20210 vdd.n390 vdd.n389 0.152939
R20211 vdd.n391 vdd.n390 0.152939
R20212 vdd.n464 vdd.n463 0.152939
R20213 vdd.n470 vdd.n463 0.152939
R20214 vdd.n471 vdd.n470 0.152939
R20215 vdd.n472 vdd.n471 0.152939
R20216 vdd.n472 vdd.n461 0.152939
R20217 vdd.n480 vdd.n461 0.152939
R20218 vdd.n481 vdd.n480 0.152939
R20219 vdd.n482 vdd.n481 0.152939
R20220 vdd.n482 vdd.n459 0.152939
R20221 vdd.n490 vdd.n459 0.152939
R20222 vdd.n491 vdd.n490 0.152939
R20223 vdd.n492 vdd.n491 0.152939
R20224 vdd.n492 vdd.n457 0.152939
R20225 vdd.n500 vdd.n457 0.152939
R20226 vdd.n501 vdd.n500 0.152939
R20227 vdd.n502 vdd.n501 0.152939
R20228 vdd.n502 vdd.n455 0.152939
R20229 vdd.n510 vdd.n455 0.152939
R20230 vdd.n511 vdd.n510 0.152939
R20231 vdd.n512 vdd.n511 0.152939
R20232 vdd.n512 vdd.n451 0.152939
R20233 vdd.n520 vdd.n451 0.152939
R20234 vdd.n521 vdd.n520 0.152939
R20235 vdd.n522 vdd.n521 0.152939
R20236 vdd.n522 vdd.n449 0.152939
R20237 vdd.n530 vdd.n449 0.152939
R20238 vdd.n531 vdd.n530 0.152939
R20239 vdd.n532 vdd.n531 0.152939
R20240 vdd.n532 vdd.n447 0.152939
R20241 vdd.n540 vdd.n447 0.152939
R20242 vdd.n541 vdd.n540 0.152939
R20243 vdd.n542 vdd.n541 0.152939
R20244 vdd.n542 vdd.n445 0.152939
R20245 vdd.n550 vdd.n445 0.152939
R20246 vdd.n551 vdd.n550 0.152939
R20247 vdd.n552 vdd.n551 0.152939
R20248 vdd.n552 vdd.n443 0.152939
R20249 vdd.n560 vdd.n443 0.152939
R20250 vdd.n561 vdd.n560 0.152939
R20251 vdd.n562 vdd.n561 0.152939
R20252 vdd.n562 vdd.n439 0.152939
R20253 vdd.n570 vdd.n439 0.152939
R20254 vdd.n571 vdd.n570 0.152939
R20255 vdd.n572 vdd.n571 0.152939
R20256 vdd.n572 vdd.n437 0.152939
R20257 vdd.n580 vdd.n437 0.152939
R20258 vdd.n581 vdd.n580 0.152939
R20259 vdd.n582 vdd.n581 0.152939
R20260 vdd.n582 vdd.n435 0.152939
R20261 vdd.n590 vdd.n435 0.152939
R20262 vdd.n591 vdd.n590 0.152939
R20263 vdd.n592 vdd.n591 0.152939
R20264 vdd.n592 vdd.n433 0.152939
R20265 vdd.n600 vdd.n433 0.152939
R20266 vdd.n601 vdd.n600 0.152939
R20267 vdd.n602 vdd.n601 0.152939
R20268 vdd.n602 vdd.n431 0.152939
R20269 vdd.n610 vdd.n431 0.152939
R20270 vdd.n611 vdd.n610 0.152939
R20271 vdd.n612 vdd.n611 0.152939
R20272 vdd.n612 vdd.n429 0.152939
R20273 vdd.n619 vdd.n429 0.152939
R20274 vdd.n3350 vdd.n619 0.152939
R20275 vdd.n3228 vdd.n3227 0.152939
R20276 vdd.n3228 vdd.n675 0.152939
R20277 vdd.n3242 vdd.n675 0.152939
R20278 vdd.n3243 vdd.n3242 0.152939
R20279 vdd.n3244 vdd.n3243 0.152939
R20280 vdd.n3244 vdd.n665 0.152939
R20281 vdd.n3259 vdd.n665 0.152939
R20282 vdd.n3260 vdd.n3259 0.152939
R20283 vdd.n3261 vdd.n3260 0.152939
R20284 vdd.n3261 vdd.n652 0.152939
R20285 vdd.n3275 vdd.n652 0.152939
R20286 vdd.n3276 vdd.n3275 0.152939
R20287 vdd.n3277 vdd.n3276 0.152939
R20288 vdd.n3277 vdd.n641 0.152939
R20289 vdd.n3292 vdd.n641 0.152939
R20290 vdd.n3293 vdd.n3292 0.152939
R20291 vdd.n3294 vdd.n3293 0.152939
R20292 vdd.n3296 vdd.n3294 0.152939
R20293 vdd.n3296 vdd.n3295 0.152939
R20294 vdd.n3295 vdd.n630 0.152939
R20295 vdd.n3313 vdd.n630 0.152939
R20296 vdd.n3314 vdd.n3313 0.152939
R20297 vdd.n3315 vdd.n3314 0.152939
R20298 vdd.n3315 vdd.n628 0.152939
R20299 vdd.n3320 vdd.n628 0.152939
R20300 vdd.n3321 vdd.n3320 0.152939
R20301 vdd.n3322 vdd.n3321 0.152939
R20302 vdd.n3322 vdd.n626 0.152939
R20303 vdd.n3327 vdd.n626 0.152939
R20304 vdd.n3328 vdd.n3327 0.152939
R20305 vdd.n3329 vdd.n3328 0.152939
R20306 vdd.n3329 vdd.n624 0.152939
R20307 vdd.n3335 vdd.n624 0.152939
R20308 vdd.n3336 vdd.n3335 0.152939
R20309 vdd.n3337 vdd.n3336 0.152939
R20310 vdd.n3337 vdd.n622 0.152939
R20311 vdd.n3342 vdd.n622 0.152939
R20312 vdd.n3343 vdd.n3342 0.152939
R20313 vdd.n3344 vdd.n3343 0.152939
R20314 vdd.n3344 vdd.n620 0.152939
R20315 vdd.n3349 vdd.n620 0.152939
R20316 vdd.n3226 vdd.n687 0.152939
R20317 vdd.n2337 vdd.n1067 0.152939
R20318 vdd.n1430 vdd.n1186 0.152939
R20319 vdd.n1431 vdd.n1430 0.152939
R20320 vdd.n1432 vdd.n1431 0.152939
R20321 vdd.n1432 vdd.n1174 0.152939
R20322 vdd.n1447 vdd.n1174 0.152939
R20323 vdd.n1448 vdd.n1447 0.152939
R20324 vdd.n1449 vdd.n1448 0.152939
R20325 vdd.n1449 vdd.n1164 0.152939
R20326 vdd.n1464 vdd.n1164 0.152939
R20327 vdd.n1465 vdd.n1464 0.152939
R20328 vdd.n1466 vdd.n1465 0.152939
R20329 vdd.n1466 vdd.n1151 0.152939
R20330 vdd.n1480 vdd.n1151 0.152939
R20331 vdd.n1481 vdd.n1480 0.152939
R20332 vdd.n1482 vdd.n1481 0.152939
R20333 vdd.n1482 vdd.n1140 0.152939
R20334 vdd.n1497 vdd.n1140 0.152939
R20335 vdd.n1498 vdd.n1497 0.152939
R20336 vdd.n1499 vdd.n1498 0.152939
R20337 vdd.n1499 vdd.n1129 0.152939
R20338 vdd.n1820 vdd.n1129 0.152939
R20339 vdd.n1821 vdd.n1820 0.152939
R20340 vdd.n1822 vdd.n1821 0.152939
R20341 vdd.n1822 vdd.n1117 0.152939
R20342 vdd.n1837 vdd.n1117 0.152939
R20343 vdd.n1838 vdd.n1837 0.152939
R20344 vdd.n1839 vdd.n1838 0.152939
R20345 vdd.n1839 vdd.n1107 0.152939
R20346 vdd.n1854 vdd.n1107 0.152939
R20347 vdd.n1855 vdd.n1854 0.152939
R20348 vdd.n1856 vdd.n1855 0.152939
R20349 vdd.n1856 vdd.n1094 0.152939
R20350 vdd.n1870 vdd.n1094 0.152939
R20351 vdd.n1871 vdd.n1870 0.152939
R20352 vdd.n1872 vdd.n1871 0.152939
R20353 vdd.n1872 vdd.n1084 0.152939
R20354 vdd.n1887 vdd.n1084 0.152939
R20355 vdd.n1888 vdd.n1887 0.152939
R20356 vdd.n1891 vdd.n1888 0.152939
R20357 vdd.n1891 vdd.n1890 0.152939
R20358 vdd.n1890 vdd.n1889 0.152939
R20359 vdd.n1422 vdd.n1191 0.152939
R20360 vdd.n1415 vdd.n1191 0.152939
R20361 vdd.n1415 vdd.n1414 0.152939
R20362 vdd.n1414 vdd.n1413 0.152939
R20363 vdd.n1413 vdd.n1228 0.152939
R20364 vdd.n1409 vdd.n1228 0.152939
R20365 vdd.n1409 vdd.n1408 0.152939
R20366 vdd.n1408 vdd.n1407 0.152939
R20367 vdd.n1407 vdd.n1234 0.152939
R20368 vdd.n1403 vdd.n1234 0.152939
R20369 vdd.n1403 vdd.n1402 0.152939
R20370 vdd.n1402 vdd.n1401 0.152939
R20371 vdd.n1401 vdd.n1240 0.152939
R20372 vdd.n1397 vdd.n1240 0.152939
R20373 vdd.n1397 vdd.n1396 0.152939
R20374 vdd.n1396 vdd.n1395 0.152939
R20375 vdd.n1395 vdd.n1246 0.152939
R20376 vdd.n1391 vdd.n1246 0.152939
R20377 vdd.n1391 vdd.n1390 0.152939
R20378 vdd.n1390 vdd.n1389 0.152939
R20379 vdd.n1389 vdd.n1254 0.152939
R20380 vdd.n1385 vdd.n1254 0.152939
R20381 vdd.n1385 vdd.n1384 0.152939
R20382 vdd.n1384 vdd.n1383 0.152939
R20383 vdd.n1383 vdd.n1260 0.152939
R20384 vdd.n1379 vdd.n1260 0.152939
R20385 vdd.n1379 vdd.n1378 0.152939
R20386 vdd.n1378 vdd.n1377 0.152939
R20387 vdd.n1377 vdd.n1266 0.152939
R20388 vdd.n1373 vdd.n1266 0.152939
R20389 vdd.n1373 vdd.n1372 0.152939
R20390 vdd.n1372 vdd.n1371 0.152939
R20391 vdd.n1371 vdd.n1272 0.152939
R20392 vdd.n1367 vdd.n1272 0.152939
R20393 vdd.n1367 vdd.n1366 0.152939
R20394 vdd.n1366 vdd.n1365 0.152939
R20395 vdd.n1365 vdd.n1278 0.152939
R20396 vdd.n1361 vdd.n1278 0.152939
R20397 vdd.n1361 vdd.n1360 0.152939
R20398 vdd.n1360 vdd.n1359 0.152939
R20399 vdd.n1359 vdd.n1284 0.152939
R20400 vdd.n1352 vdd.n1284 0.152939
R20401 vdd.n1352 vdd.n1351 0.152939
R20402 vdd.n1351 vdd.n1350 0.152939
R20403 vdd.n1350 vdd.n1289 0.152939
R20404 vdd.n1346 vdd.n1289 0.152939
R20405 vdd.n1346 vdd.n1345 0.152939
R20406 vdd.n1345 vdd.n1344 0.152939
R20407 vdd.n1344 vdd.n1295 0.152939
R20408 vdd.n1340 vdd.n1295 0.152939
R20409 vdd.n1340 vdd.n1339 0.152939
R20410 vdd.n1339 vdd.n1338 0.152939
R20411 vdd.n1338 vdd.n1301 0.152939
R20412 vdd.n1334 vdd.n1301 0.152939
R20413 vdd.n1334 vdd.n1333 0.152939
R20414 vdd.n1333 vdd.n1332 0.152939
R20415 vdd.n1332 vdd.n1307 0.152939
R20416 vdd.n1328 vdd.n1307 0.152939
R20417 vdd.n1328 vdd.n1327 0.152939
R20418 vdd.n1327 vdd.n1326 0.152939
R20419 vdd.n1326 vdd.n1313 0.152939
R20420 vdd.n1322 vdd.n1313 0.152939
R20421 vdd.n1322 vdd.n1321 0.152939
R20422 vdd.n1424 vdd.n1423 0.152939
R20423 vdd.n1424 vdd.n1180 0.152939
R20424 vdd.n1439 vdd.n1180 0.152939
R20425 vdd.n1440 vdd.n1439 0.152939
R20426 vdd.n1441 vdd.n1440 0.152939
R20427 vdd.n1441 vdd.n1169 0.152939
R20428 vdd.n1456 vdd.n1169 0.152939
R20429 vdd.n1457 vdd.n1456 0.152939
R20430 vdd.n1458 vdd.n1457 0.152939
R20431 vdd.n1458 vdd.n1158 0.152939
R20432 vdd.n1472 vdd.n1158 0.152939
R20433 vdd.n1473 vdd.n1472 0.152939
R20434 vdd.n1474 vdd.n1473 0.152939
R20435 vdd.n1474 vdd.n1146 0.152939
R20436 vdd.n1489 vdd.n1146 0.152939
R20437 vdd.n1490 vdd.n1489 0.152939
R20438 vdd.n1491 vdd.n1490 0.152939
R20439 vdd.n1491 vdd.n1135 0.152939
R20440 vdd.n1505 vdd.n1135 0.152939
R20441 vdd.n1506 vdd.n1505 0.152939
R20442 vdd.n1427 vdd.t231 0.113865
R20443 vdd.t238 vdd.n386 0.113865
R20444 vdd.n2315 vdd.n1900 0.110256
R20445 vdd.n3216 vdd.n727 0.110256
R20446 vdd.n3093 vdd.n687 0.110256
R20447 vdd.n2338 vdd.n2337 0.110256
R20448 vdd.n1814 vdd.n1813 0.0695946
R20449 vdd.n3399 vdd.n334 0.0695946
R20450 vdd.n3399 vdd.n3398 0.0695946
R20451 vdd.n1813 vdd.n1506 0.0695946
R20452 vdd.n2315 vdd.n2101 0.0431829
R20453 vdd.n2338 vdd.n1064 0.0431829
R20454 vdd.n3216 vdd.n730 0.0431829
R20455 vdd.n3093 vdd.n783 0.0431829
R20456 vdd vdd.n28 0.00833333
R20457 CSoutput.n19 CSoutput.t208 184.661
R20458 CSoutput.n78 CSoutput.n77 165.8
R20459 CSoutput.n76 CSoutput.n0 165.8
R20460 CSoutput.n75 CSoutput.n74 165.8
R20461 CSoutput.n73 CSoutput.n72 165.8
R20462 CSoutput.n71 CSoutput.n2 165.8
R20463 CSoutput.n69 CSoutput.n68 165.8
R20464 CSoutput.n67 CSoutput.n3 165.8
R20465 CSoutput.n66 CSoutput.n65 165.8
R20466 CSoutput.n63 CSoutput.n4 165.8
R20467 CSoutput.n61 CSoutput.n60 165.8
R20468 CSoutput.n59 CSoutput.n5 165.8
R20469 CSoutput.n58 CSoutput.n57 165.8
R20470 CSoutput.n55 CSoutput.n6 165.8
R20471 CSoutput.n54 CSoutput.n53 165.8
R20472 CSoutput.n52 CSoutput.n51 165.8
R20473 CSoutput.n50 CSoutput.n8 165.8
R20474 CSoutput.n48 CSoutput.n47 165.8
R20475 CSoutput.n46 CSoutput.n9 165.8
R20476 CSoutput.n45 CSoutput.n44 165.8
R20477 CSoutput.n42 CSoutput.n10 165.8
R20478 CSoutput.n41 CSoutput.n40 165.8
R20479 CSoutput.n39 CSoutput.n38 165.8
R20480 CSoutput.n37 CSoutput.n12 165.8
R20481 CSoutput.n35 CSoutput.n34 165.8
R20482 CSoutput.n33 CSoutput.n13 165.8
R20483 CSoutput.n32 CSoutput.n31 165.8
R20484 CSoutput.n29 CSoutput.n14 165.8
R20485 CSoutput.n28 CSoutput.n27 165.8
R20486 CSoutput.n26 CSoutput.n25 165.8
R20487 CSoutput.n24 CSoutput.n16 165.8
R20488 CSoutput.n22 CSoutput.n21 165.8
R20489 CSoutput.n20 CSoutput.n17 165.8
R20490 CSoutput.n77 CSoutput.t212 162.194
R20491 CSoutput.n18 CSoutput.t198 120.501
R20492 CSoutput.n23 CSoutput.t200 120.501
R20493 CSoutput.n15 CSoutput.t213 120.501
R20494 CSoutput.n30 CSoutput.t201 120.501
R20495 CSoutput.n36 CSoutput.t204 120.501
R20496 CSoutput.n11 CSoutput.t196 120.501
R20497 CSoutput.n43 CSoutput.t209 120.501
R20498 CSoutput.n49 CSoutput.t205 120.501
R20499 CSoutput.n7 CSoutput.t199 120.501
R20500 CSoutput.n56 CSoutput.t195 120.501
R20501 CSoutput.n62 CSoutput.t206 120.501
R20502 CSoutput.n64 CSoutput.t207 120.501
R20503 CSoutput.n70 CSoutput.t197 120.501
R20504 CSoutput.n1 CSoutput.t193 120.501
R20505 CSoutput.n330 CSoutput.n328 103.469
R20506 CSoutput.n310 CSoutput.n308 103.469
R20507 CSoutput.n291 CSoutput.n289 103.469
R20508 CSoutput.n120 CSoutput.n118 103.469
R20509 CSoutput.n100 CSoutput.n98 103.469
R20510 CSoutput.n81 CSoutput.n79 103.469
R20511 CSoutput.n344 CSoutput.n343 103.111
R20512 CSoutput.n342 CSoutput.n341 103.111
R20513 CSoutput.n340 CSoutput.n339 103.111
R20514 CSoutput.n338 CSoutput.n337 103.111
R20515 CSoutput.n336 CSoutput.n335 103.111
R20516 CSoutput.n334 CSoutput.n333 103.111
R20517 CSoutput.n332 CSoutput.n331 103.111
R20518 CSoutput.n330 CSoutput.n329 103.111
R20519 CSoutput.n326 CSoutput.n325 103.111
R20520 CSoutput.n324 CSoutput.n323 103.111
R20521 CSoutput.n322 CSoutput.n321 103.111
R20522 CSoutput.n320 CSoutput.n319 103.111
R20523 CSoutput.n318 CSoutput.n317 103.111
R20524 CSoutput.n316 CSoutput.n315 103.111
R20525 CSoutput.n314 CSoutput.n313 103.111
R20526 CSoutput.n312 CSoutput.n311 103.111
R20527 CSoutput.n310 CSoutput.n309 103.111
R20528 CSoutput.n307 CSoutput.n306 103.111
R20529 CSoutput.n305 CSoutput.n304 103.111
R20530 CSoutput.n303 CSoutput.n302 103.111
R20531 CSoutput.n301 CSoutput.n300 103.111
R20532 CSoutput.n299 CSoutput.n298 103.111
R20533 CSoutput.n297 CSoutput.n296 103.111
R20534 CSoutput.n295 CSoutput.n294 103.111
R20535 CSoutput.n293 CSoutput.n292 103.111
R20536 CSoutput.n291 CSoutput.n290 103.111
R20537 CSoutput.n120 CSoutput.n119 103.111
R20538 CSoutput.n122 CSoutput.n121 103.111
R20539 CSoutput.n124 CSoutput.n123 103.111
R20540 CSoutput.n126 CSoutput.n125 103.111
R20541 CSoutput.n128 CSoutput.n127 103.111
R20542 CSoutput.n130 CSoutput.n129 103.111
R20543 CSoutput.n132 CSoutput.n131 103.111
R20544 CSoutput.n134 CSoutput.n133 103.111
R20545 CSoutput.n136 CSoutput.n135 103.111
R20546 CSoutput.n100 CSoutput.n99 103.111
R20547 CSoutput.n102 CSoutput.n101 103.111
R20548 CSoutput.n104 CSoutput.n103 103.111
R20549 CSoutput.n106 CSoutput.n105 103.111
R20550 CSoutput.n108 CSoutput.n107 103.111
R20551 CSoutput.n110 CSoutput.n109 103.111
R20552 CSoutput.n112 CSoutput.n111 103.111
R20553 CSoutput.n114 CSoutput.n113 103.111
R20554 CSoutput.n116 CSoutput.n115 103.111
R20555 CSoutput.n81 CSoutput.n80 103.111
R20556 CSoutput.n83 CSoutput.n82 103.111
R20557 CSoutput.n85 CSoutput.n84 103.111
R20558 CSoutput.n87 CSoutput.n86 103.111
R20559 CSoutput.n89 CSoutput.n88 103.111
R20560 CSoutput.n91 CSoutput.n90 103.111
R20561 CSoutput.n93 CSoutput.n92 103.111
R20562 CSoutput.n95 CSoutput.n94 103.111
R20563 CSoutput.n97 CSoutput.n96 103.111
R20564 CSoutput.n346 CSoutput.n345 103.111
R20565 CSoutput.n374 CSoutput.n372 81.5057
R20566 CSoutput.n362 CSoutput.n360 81.5057
R20567 CSoutput.n351 CSoutput.n349 81.5057
R20568 CSoutput.n410 CSoutput.n408 81.5057
R20569 CSoutput.n398 CSoutput.n396 81.5057
R20570 CSoutput.n387 CSoutput.n385 81.5057
R20571 CSoutput.n382 CSoutput.n381 80.9324
R20572 CSoutput.n380 CSoutput.n379 80.9324
R20573 CSoutput.n378 CSoutput.n377 80.9324
R20574 CSoutput.n376 CSoutput.n375 80.9324
R20575 CSoutput.n374 CSoutput.n373 80.9324
R20576 CSoutput.n370 CSoutput.n369 80.9324
R20577 CSoutput.n368 CSoutput.n367 80.9324
R20578 CSoutput.n366 CSoutput.n365 80.9324
R20579 CSoutput.n364 CSoutput.n363 80.9324
R20580 CSoutput.n362 CSoutput.n361 80.9324
R20581 CSoutput.n359 CSoutput.n358 80.9324
R20582 CSoutput.n357 CSoutput.n356 80.9324
R20583 CSoutput.n355 CSoutput.n354 80.9324
R20584 CSoutput.n353 CSoutput.n352 80.9324
R20585 CSoutput.n351 CSoutput.n350 80.9324
R20586 CSoutput.n410 CSoutput.n409 80.9324
R20587 CSoutput.n412 CSoutput.n411 80.9324
R20588 CSoutput.n414 CSoutput.n413 80.9324
R20589 CSoutput.n416 CSoutput.n415 80.9324
R20590 CSoutput.n418 CSoutput.n417 80.9324
R20591 CSoutput.n398 CSoutput.n397 80.9324
R20592 CSoutput.n400 CSoutput.n399 80.9324
R20593 CSoutput.n402 CSoutput.n401 80.9324
R20594 CSoutput.n404 CSoutput.n403 80.9324
R20595 CSoutput.n406 CSoutput.n405 80.9324
R20596 CSoutput.n387 CSoutput.n386 80.9324
R20597 CSoutput.n389 CSoutput.n388 80.9324
R20598 CSoutput.n391 CSoutput.n390 80.9324
R20599 CSoutput.n393 CSoutput.n392 80.9324
R20600 CSoutput.n395 CSoutput.n394 80.9324
R20601 CSoutput.n25 CSoutput.n24 48.1486
R20602 CSoutput.n69 CSoutput.n3 48.1486
R20603 CSoutput.n38 CSoutput.n37 48.1486
R20604 CSoutput.n42 CSoutput.n41 48.1486
R20605 CSoutput.n51 CSoutput.n50 48.1486
R20606 CSoutput.n55 CSoutput.n54 48.1486
R20607 CSoutput.n22 CSoutput.n17 46.462
R20608 CSoutput.n72 CSoutput.n71 46.462
R20609 CSoutput.n20 CSoutput.n19 44.9055
R20610 CSoutput.n29 CSoutput.n28 43.7635
R20611 CSoutput.n65 CSoutput.n63 43.7635
R20612 CSoutput.n35 CSoutput.n13 41.7396
R20613 CSoutput.n57 CSoutput.n5 41.7396
R20614 CSoutput.n44 CSoutput.n9 37.0171
R20615 CSoutput.n48 CSoutput.n9 37.0171
R20616 CSoutput.n76 CSoutput.n75 34.9932
R20617 CSoutput.n31 CSoutput.n13 32.2947
R20618 CSoutput.n61 CSoutput.n5 32.2947
R20619 CSoutput.n30 CSoutput.n29 29.6014
R20620 CSoutput.n63 CSoutput.n62 29.6014
R20621 CSoutput.n19 CSoutput.n18 28.4085
R20622 CSoutput.n18 CSoutput.n17 25.1176
R20623 CSoutput.n72 CSoutput.n1 25.1176
R20624 CSoutput.n43 CSoutput.n42 22.0922
R20625 CSoutput.n50 CSoutput.n49 22.0922
R20626 CSoutput.n77 CSoutput.n76 21.8586
R20627 CSoutput.n37 CSoutput.n36 18.9681
R20628 CSoutput.n56 CSoutput.n55 18.9681
R20629 CSoutput.n25 CSoutput.n15 17.6292
R20630 CSoutput.n64 CSoutput.n3 17.6292
R20631 CSoutput.n24 CSoutput.n23 15.844
R20632 CSoutput.n70 CSoutput.n69 15.844
R20633 CSoutput.n38 CSoutput.n11 14.5051
R20634 CSoutput.n54 CSoutput.n7 14.5051
R20635 CSoutput.n421 CSoutput.n78 11.4982
R20636 CSoutput.n41 CSoutput.n11 11.3811
R20637 CSoutput.n51 CSoutput.n7 11.3811
R20638 CSoutput.n23 CSoutput.n22 10.0422
R20639 CSoutput.n71 CSoutput.n70 10.0422
R20640 CSoutput.n327 CSoutput.n307 9.25285
R20641 CSoutput.n117 CSoutput.n97 9.25285
R20642 CSoutput.n371 CSoutput.n359 8.98182
R20643 CSoutput.n407 CSoutput.n395 8.98182
R20644 CSoutput.n384 CSoutput.n348 8.76129
R20645 CSoutput.n28 CSoutput.n15 8.25698
R20646 CSoutput.n65 CSoutput.n64 8.25698
R20647 CSoutput.n348 CSoutput.n347 7.12641
R20648 CSoutput.n138 CSoutput.n137 7.12641
R20649 CSoutput.n36 CSoutput.n35 6.91809
R20650 CSoutput.n57 CSoutput.n56 6.91809
R20651 CSoutput.n384 CSoutput.n383 6.02792
R20652 CSoutput.n420 CSoutput.n419 6.02792
R20653 CSoutput.n383 CSoutput.n382 5.25266
R20654 CSoutput.n371 CSoutput.n370 5.25266
R20655 CSoutput.n419 CSoutput.n418 5.25266
R20656 CSoutput.n407 CSoutput.n406 5.25266
R20657 CSoutput.n421 CSoutput.n138 5.16885
R20658 CSoutput.n347 CSoutput.n346 5.1449
R20659 CSoutput.n327 CSoutput.n326 5.1449
R20660 CSoutput.n137 CSoutput.n136 5.1449
R20661 CSoutput.n117 CSoutput.n116 5.1449
R20662 CSoutput.n229 CSoutput.n182 4.5005
R20663 CSoutput.n198 CSoutput.n182 4.5005
R20664 CSoutput.n193 CSoutput.n177 4.5005
R20665 CSoutput.n193 CSoutput.n179 4.5005
R20666 CSoutput.n193 CSoutput.n176 4.5005
R20667 CSoutput.n193 CSoutput.n180 4.5005
R20668 CSoutput.n193 CSoutput.n175 4.5005
R20669 CSoutput.n193 CSoutput.t210 4.5005
R20670 CSoutput.n193 CSoutput.n174 4.5005
R20671 CSoutput.n193 CSoutput.n181 4.5005
R20672 CSoutput.n193 CSoutput.n182 4.5005
R20673 CSoutput.n191 CSoutput.n177 4.5005
R20674 CSoutput.n191 CSoutput.n179 4.5005
R20675 CSoutput.n191 CSoutput.n176 4.5005
R20676 CSoutput.n191 CSoutput.n180 4.5005
R20677 CSoutput.n191 CSoutput.n175 4.5005
R20678 CSoutput.n191 CSoutput.t210 4.5005
R20679 CSoutput.n191 CSoutput.n174 4.5005
R20680 CSoutput.n191 CSoutput.n181 4.5005
R20681 CSoutput.n191 CSoutput.n182 4.5005
R20682 CSoutput.n190 CSoutput.n177 4.5005
R20683 CSoutput.n190 CSoutput.n179 4.5005
R20684 CSoutput.n190 CSoutput.n176 4.5005
R20685 CSoutput.n190 CSoutput.n180 4.5005
R20686 CSoutput.n190 CSoutput.n175 4.5005
R20687 CSoutput.n190 CSoutput.t210 4.5005
R20688 CSoutput.n190 CSoutput.n174 4.5005
R20689 CSoutput.n190 CSoutput.n181 4.5005
R20690 CSoutput.n190 CSoutput.n182 4.5005
R20691 CSoutput.n275 CSoutput.n177 4.5005
R20692 CSoutput.n275 CSoutput.n179 4.5005
R20693 CSoutput.n275 CSoutput.n176 4.5005
R20694 CSoutput.n275 CSoutput.n180 4.5005
R20695 CSoutput.n275 CSoutput.n175 4.5005
R20696 CSoutput.n275 CSoutput.t210 4.5005
R20697 CSoutput.n275 CSoutput.n174 4.5005
R20698 CSoutput.n275 CSoutput.n181 4.5005
R20699 CSoutput.n275 CSoutput.n182 4.5005
R20700 CSoutput.n273 CSoutput.n177 4.5005
R20701 CSoutput.n273 CSoutput.n179 4.5005
R20702 CSoutput.n273 CSoutput.n176 4.5005
R20703 CSoutput.n273 CSoutput.n180 4.5005
R20704 CSoutput.n273 CSoutput.n175 4.5005
R20705 CSoutput.n273 CSoutput.t210 4.5005
R20706 CSoutput.n273 CSoutput.n174 4.5005
R20707 CSoutput.n273 CSoutput.n181 4.5005
R20708 CSoutput.n271 CSoutput.n177 4.5005
R20709 CSoutput.n271 CSoutput.n179 4.5005
R20710 CSoutput.n271 CSoutput.n176 4.5005
R20711 CSoutput.n271 CSoutput.n180 4.5005
R20712 CSoutput.n271 CSoutput.n175 4.5005
R20713 CSoutput.n271 CSoutput.t210 4.5005
R20714 CSoutput.n271 CSoutput.n174 4.5005
R20715 CSoutput.n271 CSoutput.n181 4.5005
R20716 CSoutput.n201 CSoutput.n177 4.5005
R20717 CSoutput.n201 CSoutput.n179 4.5005
R20718 CSoutput.n201 CSoutput.n176 4.5005
R20719 CSoutput.n201 CSoutput.n180 4.5005
R20720 CSoutput.n201 CSoutput.n175 4.5005
R20721 CSoutput.n201 CSoutput.t210 4.5005
R20722 CSoutput.n201 CSoutput.n174 4.5005
R20723 CSoutput.n201 CSoutput.n181 4.5005
R20724 CSoutput.n201 CSoutput.n182 4.5005
R20725 CSoutput.n200 CSoutput.n177 4.5005
R20726 CSoutput.n200 CSoutput.n179 4.5005
R20727 CSoutput.n200 CSoutput.n176 4.5005
R20728 CSoutput.n200 CSoutput.n180 4.5005
R20729 CSoutput.n200 CSoutput.n175 4.5005
R20730 CSoutput.n200 CSoutput.t210 4.5005
R20731 CSoutput.n200 CSoutput.n174 4.5005
R20732 CSoutput.n200 CSoutput.n181 4.5005
R20733 CSoutput.n200 CSoutput.n182 4.5005
R20734 CSoutput.n204 CSoutput.n177 4.5005
R20735 CSoutput.n204 CSoutput.n179 4.5005
R20736 CSoutput.n204 CSoutput.n176 4.5005
R20737 CSoutput.n204 CSoutput.n180 4.5005
R20738 CSoutput.n204 CSoutput.n175 4.5005
R20739 CSoutput.n204 CSoutput.t210 4.5005
R20740 CSoutput.n204 CSoutput.n174 4.5005
R20741 CSoutput.n204 CSoutput.n181 4.5005
R20742 CSoutput.n204 CSoutput.n182 4.5005
R20743 CSoutput.n203 CSoutput.n177 4.5005
R20744 CSoutput.n203 CSoutput.n179 4.5005
R20745 CSoutput.n203 CSoutput.n176 4.5005
R20746 CSoutput.n203 CSoutput.n180 4.5005
R20747 CSoutput.n203 CSoutput.n175 4.5005
R20748 CSoutput.n203 CSoutput.t210 4.5005
R20749 CSoutput.n203 CSoutput.n174 4.5005
R20750 CSoutput.n203 CSoutput.n181 4.5005
R20751 CSoutput.n203 CSoutput.n182 4.5005
R20752 CSoutput.n186 CSoutput.n177 4.5005
R20753 CSoutput.n186 CSoutput.n179 4.5005
R20754 CSoutput.n186 CSoutput.n176 4.5005
R20755 CSoutput.n186 CSoutput.n180 4.5005
R20756 CSoutput.n186 CSoutput.n175 4.5005
R20757 CSoutput.n186 CSoutput.t210 4.5005
R20758 CSoutput.n186 CSoutput.n174 4.5005
R20759 CSoutput.n186 CSoutput.n181 4.5005
R20760 CSoutput.n186 CSoutput.n182 4.5005
R20761 CSoutput.n278 CSoutput.n177 4.5005
R20762 CSoutput.n278 CSoutput.n179 4.5005
R20763 CSoutput.n278 CSoutput.n176 4.5005
R20764 CSoutput.n278 CSoutput.n180 4.5005
R20765 CSoutput.n278 CSoutput.n175 4.5005
R20766 CSoutput.n278 CSoutput.t210 4.5005
R20767 CSoutput.n278 CSoutput.n174 4.5005
R20768 CSoutput.n278 CSoutput.n181 4.5005
R20769 CSoutput.n278 CSoutput.n182 4.5005
R20770 CSoutput.n265 CSoutput.n236 4.5005
R20771 CSoutput.n265 CSoutput.n242 4.5005
R20772 CSoutput.n223 CSoutput.n212 4.5005
R20773 CSoutput.n223 CSoutput.n214 4.5005
R20774 CSoutput.n223 CSoutput.n211 4.5005
R20775 CSoutput.n223 CSoutput.n215 4.5005
R20776 CSoutput.n223 CSoutput.n210 4.5005
R20777 CSoutput.n223 CSoutput.t203 4.5005
R20778 CSoutput.n223 CSoutput.n209 4.5005
R20779 CSoutput.n223 CSoutput.n216 4.5005
R20780 CSoutput.n265 CSoutput.n223 4.5005
R20781 CSoutput.n244 CSoutput.n212 4.5005
R20782 CSoutput.n244 CSoutput.n214 4.5005
R20783 CSoutput.n244 CSoutput.n211 4.5005
R20784 CSoutput.n244 CSoutput.n215 4.5005
R20785 CSoutput.n244 CSoutput.n210 4.5005
R20786 CSoutput.n244 CSoutput.t203 4.5005
R20787 CSoutput.n244 CSoutput.n209 4.5005
R20788 CSoutput.n244 CSoutput.n216 4.5005
R20789 CSoutput.n265 CSoutput.n244 4.5005
R20790 CSoutput.n222 CSoutput.n212 4.5005
R20791 CSoutput.n222 CSoutput.n214 4.5005
R20792 CSoutput.n222 CSoutput.n211 4.5005
R20793 CSoutput.n222 CSoutput.n215 4.5005
R20794 CSoutput.n222 CSoutput.n210 4.5005
R20795 CSoutput.n222 CSoutput.t203 4.5005
R20796 CSoutput.n222 CSoutput.n209 4.5005
R20797 CSoutput.n222 CSoutput.n216 4.5005
R20798 CSoutput.n265 CSoutput.n222 4.5005
R20799 CSoutput.n246 CSoutput.n212 4.5005
R20800 CSoutput.n246 CSoutput.n214 4.5005
R20801 CSoutput.n246 CSoutput.n211 4.5005
R20802 CSoutput.n246 CSoutput.n215 4.5005
R20803 CSoutput.n246 CSoutput.n210 4.5005
R20804 CSoutput.n246 CSoutput.t203 4.5005
R20805 CSoutput.n246 CSoutput.n209 4.5005
R20806 CSoutput.n246 CSoutput.n216 4.5005
R20807 CSoutput.n265 CSoutput.n246 4.5005
R20808 CSoutput.n212 CSoutput.n207 4.5005
R20809 CSoutput.n214 CSoutput.n207 4.5005
R20810 CSoutput.n211 CSoutput.n207 4.5005
R20811 CSoutput.n215 CSoutput.n207 4.5005
R20812 CSoutput.n210 CSoutput.n207 4.5005
R20813 CSoutput.t203 CSoutput.n207 4.5005
R20814 CSoutput.n209 CSoutput.n207 4.5005
R20815 CSoutput.n216 CSoutput.n207 4.5005
R20816 CSoutput.n268 CSoutput.n212 4.5005
R20817 CSoutput.n268 CSoutput.n214 4.5005
R20818 CSoutput.n268 CSoutput.n211 4.5005
R20819 CSoutput.n268 CSoutput.n215 4.5005
R20820 CSoutput.n268 CSoutput.n210 4.5005
R20821 CSoutput.n268 CSoutput.t203 4.5005
R20822 CSoutput.n268 CSoutput.n209 4.5005
R20823 CSoutput.n268 CSoutput.n216 4.5005
R20824 CSoutput.n266 CSoutput.n212 4.5005
R20825 CSoutput.n266 CSoutput.n214 4.5005
R20826 CSoutput.n266 CSoutput.n211 4.5005
R20827 CSoutput.n266 CSoutput.n215 4.5005
R20828 CSoutput.n266 CSoutput.n210 4.5005
R20829 CSoutput.n266 CSoutput.t203 4.5005
R20830 CSoutput.n266 CSoutput.n209 4.5005
R20831 CSoutput.n266 CSoutput.n216 4.5005
R20832 CSoutput.n266 CSoutput.n265 4.5005
R20833 CSoutput.n248 CSoutput.n212 4.5005
R20834 CSoutput.n248 CSoutput.n214 4.5005
R20835 CSoutput.n248 CSoutput.n211 4.5005
R20836 CSoutput.n248 CSoutput.n215 4.5005
R20837 CSoutput.n248 CSoutput.n210 4.5005
R20838 CSoutput.n248 CSoutput.t203 4.5005
R20839 CSoutput.n248 CSoutput.n209 4.5005
R20840 CSoutput.n248 CSoutput.n216 4.5005
R20841 CSoutput.n265 CSoutput.n248 4.5005
R20842 CSoutput.n220 CSoutput.n212 4.5005
R20843 CSoutput.n220 CSoutput.n214 4.5005
R20844 CSoutput.n220 CSoutput.n211 4.5005
R20845 CSoutput.n220 CSoutput.n215 4.5005
R20846 CSoutput.n220 CSoutput.n210 4.5005
R20847 CSoutput.n220 CSoutput.t203 4.5005
R20848 CSoutput.n220 CSoutput.n209 4.5005
R20849 CSoutput.n220 CSoutput.n216 4.5005
R20850 CSoutput.n265 CSoutput.n220 4.5005
R20851 CSoutput.n250 CSoutput.n212 4.5005
R20852 CSoutput.n250 CSoutput.n214 4.5005
R20853 CSoutput.n250 CSoutput.n211 4.5005
R20854 CSoutput.n250 CSoutput.n215 4.5005
R20855 CSoutput.n250 CSoutput.n210 4.5005
R20856 CSoutput.n250 CSoutput.t203 4.5005
R20857 CSoutput.n250 CSoutput.n209 4.5005
R20858 CSoutput.n250 CSoutput.n216 4.5005
R20859 CSoutput.n265 CSoutput.n250 4.5005
R20860 CSoutput.n219 CSoutput.n212 4.5005
R20861 CSoutput.n219 CSoutput.n214 4.5005
R20862 CSoutput.n219 CSoutput.n211 4.5005
R20863 CSoutput.n219 CSoutput.n215 4.5005
R20864 CSoutput.n219 CSoutput.n210 4.5005
R20865 CSoutput.n219 CSoutput.t203 4.5005
R20866 CSoutput.n219 CSoutput.n209 4.5005
R20867 CSoutput.n219 CSoutput.n216 4.5005
R20868 CSoutput.n265 CSoutput.n219 4.5005
R20869 CSoutput.n264 CSoutput.n212 4.5005
R20870 CSoutput.n264 CSoutput.n214 4.5005
R20871 CSoutput.n264 CSoutput.n211 4.5005
R20872 CSoutput.n264 CSoutput.n215 4.5005
R20873 CSoutput.n264 CSoutput.n210 4.5005
R20874 CSoutput.n264 CSoutput.t203 4.5005
R20875 CSoutput.n264 CSoutput.n209 4.5005
R20876 CSoutput.n264 CSoutput.n216 4.5005
R20877 CSoutput.n265 CSoutput.n264 4.5005
R20878 CSoutput.n263 CSoutput.n148 4.5005
R20879 CSoutput.n164 CSoutput.n148 4.5005
R20880 CSoutput.n159 CSoutput.n143 4.5005
R20881 CSoutput.n159 CSoutput.n145 4.5005
R20882 CSoutput.n159 CSoutput.n142 4.5005
R20883 CSoutput.n159 CSoutput.n146 4.5005
R20884 CSoutput.n159 CSoutput.n141 4.5005
R20885 CSoutput.n159 CSoutput.t202 4.5005
R20886 CSoutput.n159 CSoutput.n140 4.5005
R20887 CSoutput.n159 CSoutput.n147 4.5005
R20888 CSoutput.n159 CSoutput.n148 4.5005
R20889 CSoutput.n157 CSoutput.n143 4.5005
R20890 CSoutput.n157 CSoutput.n145 4.5005
R20891 CSoutput.n157 CSoutput.n142 4.5005
R20892 CSoutput.n157 CSoutput.n146 4.5005
R20893 CSoutput.n157 CSoutput.n141 4.5005
R20894 CSoutput.n157 CSoutput.t202 4.5005
R20895 CSoutput.n157 CSoutput.n140 4.5005
R20896 CSoutput.n157 CSoutput.n147 4.5005
R20897 CSoutput.n157 CSoutput.n148 4.5005
R20898 CSoutput.n156 CSoutput.n143 4.5005
R20899 CSoutput.n156 CSoutput.n145 4.5005
R20900 CSoutput.n156 CSoutput.n142 4.5005
R20901 CSoutput.n156 CSoutput.n146 4.5005
R20902 CSoutput.n156 CSoutput.n141 4.5005
R20903 CSoutput.n156 CSoutput.t202 4.5005
R20904 CSoutput.n156 CSoutput.n140 4.5005
R20905 CSoutput.n156 CSoutput.n147 4.5005
R20906 CSoutput.n156 CSoutput.n148 4.5005
R20907 CSoutput.n285 CSoutput.n143 4.5005
R20908 CSoutput.n285 CSoutput.n145 4.5005
R20909 CSoutput.n285 CSoutput.n142 4.5005
R20910 CSoutput.n285 CSoutput.n146 4.5005
R20911 CSoutput.n285 CSoutput.n141 4.5005
R20912 CSoutput.n285 CSoutput.t202 4.5005
R20913 CSoutput.n285 CSoutput.n140 4.5005
R20914 CSoutput.n285 CSoutput.n147 4.5005
R20915 CSoutput.n285 CSoutput.n148 4.5005
R20916 CSoutput.n283 CSoutput.n143 4.5005
R20917 CSoutput.n283 CSoutput.n145 4.5005
R20918 CSoutput.n283 CSoutput.n142 4.5005
R20919 CSoutput.n283 CSoutput.n146 4.5005
R20920 CSoutput.n283 CSoutput.n141 4.5005
R20921 CSoutput.n283 CSoutput.t202 4.5005
R20922 CSoutput.n283 CSoutput.n140 4.5005
R20923 CSoutput.n283 CSoutput.n147 4.5005
R20924 CSoutput.n281 CSoutput.n143 4.5005
R20925 CSoutput.n281 CSoutput.n145 4.5005
R20926 CSoutput.n281 CSoutput.n142 4.5005
R20927 CSoutput.n281 CSoutput.n146 4.5005
R20928 CSoutput.n281 CSoutput.n141 4.5005
R20929 CSoutput.n281 CSoutput.t202 4.5005
R20930 CSoutput.n281 CSoutput.n140 4.5005
R20931 CSoutput.n281 CSoutput.n147 4.5005
R20932 CSoutput.n167 CSoutput.n143 4.5005
R20933 CSoutput.n167 CSoutput.n145 4.5005
R20934 CSoutput.n167 CSoutput.n142 4.5005
R20935 CSoutput.n167 CSoutput.n146 4.5005
R20936 CSoutput.n167 CSoutput.n141 4.5005
R20937 CSoutput.n167 CSoutput.t202 4.5005
R20938 CSoutput.n167 CSoutput.n140 4.5005
R20939 CSoutput.n167 CSoutput.n147 4.5005
R20940 CSoutput.n167 CSoutput.n148 4.5005
R20941 CSoutput.n166 CSoutput.n143 4.5005
R20942 CSoutput.n166 CSoutput.n145 4.5005
R20943 CSoutput.n166 CSoutput.n142 4.5005
R20944 CSoutput.n166 CSoutput.n146 4.5005
R20945 CSoutput.n166 CSoutput.n141 4.5005
R20946 CSoutput.n166 CSoutput.t202 4.5005
R20947 CSoutput.n166 CSoutput.n140 4.5005
R20948 CSoutput.n166 CSoutput.n147 4.5005
R20949 CSoutput.n166 CSoutput.n148 4.5005
R20950 CSoutput.n170 CSoutput.n143 4.5005
R20951 CSoutput.n170 CSoutput.n145 4.5005
R20952 CSoutput.n170 CSoutput.n142 4.5005
R20953 CSoutput.n170 CSoutput.n146 4.5005
R20954 CSoutput.n170 CSoutput.n141 4.5005
R20955 CSoutput.n170 CSoutput.t202 4.5005
R20956 CSoutput.n170 CSoutput.n140 4.5005
R20957 CSoutput.n170 CSoutput.n147 4.5005
R20958 CSoutput.n170 CSoutput.n148 4.5005
R20959 CSoutput.n169 CSoutput.n143 4.5005
R20960 CSoutput.n169 CSoutput.n145 4.5005
R20961 CSoutput.n169 CSoutput.n142 4.5005
R20962 CSoutput.n169 CSoutput.n146 4.5005
R20963 CSoutput.n169 CSoutput.n141 4.5005
R20964 CSoutput.n169 CSoutput.t202 4.5005
R20965 CSoutput.n169 CSoutput.n140 4.5005
R20966 CSoutput.n169 CSoutput.n147 4.5005
R20967 CSoutput.n169 CSoutput.n148 4.5005
R20968 CSoutput.n152 CSoutput.n143 4.5005
R20969 CSoutput.n152 CSoutput.n145 4.5005
R20970 CSoutput.n152 CSoutput.n142 4.5005
R20971 CSoutput.n152 CSoutput.n146 4.5005
R20972 CSoutput.n152 CSoutput.n141 4.5005
R20973 CSoutput.n152 CSoutput.t202 4.5005
R20974 CSoutput.n152 CSoutput.n140 4.5005
R20975 CSoutput.n152 CSoutput.n147 4.5005
R20976 CSoutput.n152 CSoutput.n148 4.5005
R20977 CSoutput.n288 CSoutput.n143 4.5005
R20978 CSoutput.n288 CSoutput.n145 4.5005
R20979 CSoutput.n288 CSoutput.n142 4.5005
R20980 CSoutput.n288 CSoutput.n146 4.5005
R20981 CSoutput.n288 CSoutput.n141 4.5005
R20982 CSoutput.n288 CSoutput.t202 4.5005
R20983 CSoutput.n288 CSoutput.n140 4.5005
R20984 CSoutput.n288 CSoutput.n147 4.5005
R20985 CSoutput.n288 CSoutput.n148 4.5005
R20986 CSoutput.n347 CSoutput.n327 4.10845
R20987 CSoutput.n137 CSoutput.n117 4.10845
R20988 CSoutput.n345 CSoutput.t67 4.06363
R20989 CSoutput.n345 CSoutput.t91 4.06363
R20990 CSoutput.n343 CSoutput.t111 4.06363
R20991 CSoutput.n343 CSoutput.t25 4.06363
R20992 CSoutput.n341 CSoutput.t29 4.06363
R20993 CSoutput.n341 CSoutput.t95 4.06363
R20994 CSoutput.n339 CSoutput.t114 4.06363
R20995 CSoutput.n339 CSoutput.t115 4.06363
R20996 CSoutput.n337 CSoutput.t45 4.06363
R20997 CSoutput.n337 CSoutput.t46 4.06363
R20998 CSoutput.n335 CSoutput.t51 4.06363
R20999 CSoutput.n335 CSoutput.t116 4.06363
R21000 CSoutput.n333 CSoutput.t15 4.06363
R21001 CSoutput.n333 CSoutput.t49 4.06363
R21002 CSoutput.n331 CSoutput.t66 4.06363
R21003 CSoutput.n331 CSoutput.t90 4.06363
R21004 CSoutput.n329 CSoutput.t97 4.06363
R21005 CSoutput.n329 CSoutput.t21 4.06363
R21006 CSoutput.n328 CSoutput.t69 4.06363
R21007 CSoutput.n328 CSoutput.t70 4.06363
R21008 CSoutput.n325 CSoutput.t52 4.06363
R21009 CSoutput.n325 CSoutput.t79 4.06363
R21010 CSoutput.n323 CSoutput.t99 4.06363
R21011 CSoutput.n323 CSoutput.t11 4.06363
R21012 CSoutput.n321 CSoutput.t12 4.06363
R21013 CSoutput.n321 CSoutput.t81 4.06363
R21014 CSoutput.n319 CSoutput.t102 4.06363
R21015 CSoutput.n319 CSoutput.t103 4.06363
R21016 CSoutput.n317 CSoutput.t33 4.06363
R21017 CSoutput.n317 CSoutput.t34 4.06363
R21018 CSoutput.n315 CSoutput.t37 4.06363
R21019 CSoutput.n315 CSoutput.t106 4.06363
R21020 CSoutput.n313 CSoutput.t0 4.06363
R21021 CSoutput.n313 CSoutput.t36 4.06363
R21022 CSoutput.n311 CSoutput.t53 4.06363
R21023 CSoutput.n311 CSoutput.t80 4.06363
R21024 CSoutput.n309 CSoutput.t82 4.06363
R21025 CSoutput.n309 CSoutput.t6 4.06363
R21026 CSoutput.n308 CSoutput.t59 4.06363
R21027 CSoutput.n308 CSoutput.t60 4.06363
R21028 CSoutput.n306 CSoutput.t88 4.06363
R21029 CSoutput.n306 CSoutput.t42 4.06363
R21030 CSoutput.n304 CSoutput.t75 4.06363
R21031 CSoutput.n304 CSoutput.t24 4.06363
R21032 CSoutput.n302 CSoutput.t100 4.06363
R21033 CSoutput.n302 CSoutput.t16 4.06363
R21034 CSoutput.n300 CSoutput.t56 4.06363
R21035 CSoutput.n300 CSoutput.t35 4.06363
R21036 CSoutput.n298 CSoutput.t38 4.06363
R21037 CSoutput.n298 CSoutput.t13 4.06363
R21038 CSoutput.n296 CSoutput.t87 4.06363
R21039 CSoutput.n296 CSoutput.t7 4.06363
R21040 CSoutput.n294 CSoutput.t47 4.06363
R21041 CSoutput.n294 CSoutput.t112 4.06363
R21042 CSoutput.n292 CSoutput.t30 4.06363
R21043 CSoutput.n292 CSoutput.t93 4.06363
R21044 CSoutput.n290 CSoutput.t54 4.06363
R21045 CSoutput.n290 CSoutput.t117 4.06363
R21046 CSoutput.n289 CSoutput.t1 4.06363
R21047 CSoutput.n289 CSoutput.t104 4.06363
R21048 CSoutput.n118 CSoutput.t110 4.06363
R21049 CSoutput.n118 CSoutput.t109 4.06363
R21050 CSoutput.n119 CSoutput.t89 4.06363
R21051 CSoutput.n119 CSoutput.t23 4.06363
R21052 CSoutput.n121 CSoutput.t19 4.06363
R21053 CSoutput.n121 CSoutput.t107 4.06363
R21054 CSoutput.n123 CSoutput.t86 4.06363
R21055 CSoutput.n123 CSoutput.t63 4.06363
R21056 CSoutput.n125 CSoutput.t44 4.06363
R21057 CSoutput.n125 CSoutput.t119 4.06363
R21058 CSoutput.n127 CSoutput.t84 4.06363
R21059 CSoutput.n127 CSoutput.t83 4.06363
R21060 CSoutput.n129 CSoutput.t71 4.06363
R21061 CSoutput.n129 CSoutput.t41 4.06363
R21062 CSoutput.n131 CSoutput.t22 4.06363
R21063 CSoutput.n131 CSoutput.t72 4.06363
R21064 CSoutput.n133 CSoutput.t68 4.06363
R21065 CSoutput.n133 CSoutput.t39 4.06363
R21066 CSoutput.n135 CSoutput.t20 4.06363
R21067 CSoutput.n135 CSoutput.t18 4.06363
R21068 CSoutput.n98 CSoutput.t98 4.06363
R21069 CSoutput.n98 CSoutput.t96 4.06363
R21070 CSoutput.n99 CSoutput.t78 4.06363
R21071 CSoutput.n99 CSoutput.t10 4.06363
R21072 CSoutput.n101 CSoutput.t4 4.06363
R21073 CSoutput.n101 CSoutput.t92 4.06363
R21074 CSoutput.n103 CSoutput.t77 4.06363
R21075 CSoutput.n103 CSoutput.t50 4.06363
R21076 CSoutput.n105 CSoutput.t32 4.06363
R21077 CSoutput.n105 CSoutput.t108 4.06363
R21078 CSoutput.n107 CSoutput.t74 4.06363
R21079 CSoutput.n107 CSoutput.t73 4.06363
R21080 CSoutput.n109 CSoutput.t61 4.06363
R21081 CSoutput.n109 CSoutput.t28 4.06363
R21082 CSoutput.n111 CSoutput.t8 4.06363
R21083 CSoutput.n111 CSoutput.t62 4.06363
R21084 CSoutput.n113 CSoutput.t58 4.06363
R21085 CSoutput.n113 CSoutput.t26 4.06363
R21086 CSoutput.n115 CSoutput.t5 4.06363
R21087 CSoutput.n115 CSoutput.t2 4.06363
R21088 CSoutput.n79 CSoutput.t105 4.06363
R21089 CSoutput.n79 CSoutput.t3 4.06363
R21090 CSoutput.n80 CSoutput.t85 4.06363
R21091 CSoutput.n80 CSoutput.t55 4.06363
R21092 CSoutput.n82 CSoutput.t94 4.06363
R21093 CSoutput.n82 CSoutput.t31 4.06363
R21094 CSoutput.n84 CSoutput.t113 4.06363
R21095 CSoutput.n84 CSoutput.t48 4.06363
R21096 CSoutput.n86 CSoutput.t9 4.06363
R21097 CSoutput.n86 CSoutput.t64 4.06363
R21098 CSoutput.n88 CSoutput.t14 4.06363
R21099 CSoutput.n88 CSoutput.t40 4.06363
R21100 CSoutput.n90 CSoutput.t118 4.06363
R21101 CSoutput.n90 CSoutput.t57 4.06363
R21102 CSoutput.n92 CSoutput.t17 4.06363
R21103 CSoutput.n92 CSoutput.t101 4.06363
R21104 CSoutput.n94 CSoutput.t27 4.06363
R21105 CSoutput.n94 CSoutput.t76 4.06363
R21106 CSoutput.n96 CSoutput.t43 4.06363
R21107 CSoutput.n96 CSoutput.t65 4.06363
R21108 CSoutput.n44 CSoutput.n43 3.79402
R21109 CSoutput.n49 CSoutput.n48 3.79402
R21110 CSoutput.n383 CSoutput.n371 3.72967
R21111 CSoutput.n419 CSoutput.n407 3.72967
R21112 CSoutput.n421 CSoutput.n420 3.57343
R21113 CSoutput.n420 CSoutput.n384 3.04641
R21114 CSoutput.n381 CSoutput.t164 2.82907
R21115 CSoutput.n381 CSoutput.t121 2.82907
R21116 CSoutput.n379 CSoutput.t190 2.82907
R21117 CSoutput.n379 CSoutput.t179 2.82907
R21118 CSoutput.n377 CSoutput.t146 2.82907
R21119 CSoutput.n377 CSoutput.t155 2.82907
R21120 CSoutput.n375 CSoutput.t120 2.82907
R21121 CSoutput.n375 CSoutput.t186 2.82907
R21122 CSoutput.n373 CSoutput.t180 2.82907
R21123 CSoutput.n373 CSoutput.t135 2.82907
R21124 CSoutput.n372 CSoutput.t128 2.82907
R21125 CSoutput.n372 CSoutput.t189 2.82907
R21126 CSoutput.n369 CSoutput.t131 2.82907
R21127 CSoutput.n369 CSoutput.t141 2.82907
R21128 CSoutput.n367 CSoutput.t139 2.82907
R21129 CSoutput.n367 CSoutput.t127 2.82907
R21130 CSoutput.n365 CSoutput.t152 2.82907
R21131 CSoutput.n365 CSoutput.t132 2.82907
R21132 CSoutput.n363 CSoutput.t133 2.82907
R21133 CSoutput.n363 CSoutput.t140 2.82907
R21134 CSoutput.n361 CSoutput.t138 2.82907
R21135 CSoutput.n361 CSoutput.t150 2.82907
R21136 CSoutput.n360 CSoutput.t151 2.82907
R21137 CSoutput.n360 CSoutput.t134 2.82907
R21138 CSoutput.n358 CSoutput.t173 2.82907
R21139 CSoutput.n358 CSoutput.t143 2.82907
R21140 CSoutput.n356 CSoutput.t124 2.82907
R21141 CSoutput.n356 CSoutput.t159 2.82907
R21142 CSoutput.n354 CSoutput.t142 2.82907
R21143 CSoutput.n354 CSoutput.t153 2.82907
R21144 CSoutput.n352 CSoutput.t154 2.82907
R21145 CSoutput.n352 CSoutput.t185 2.82907
R21146 CSoutput.n350 CSoutput.t169 2.82907
R21147 CSoutput.n350 CSoutput.t122 2.82907
R21148 CSoutput.n349 CSoutput.t182 2.82907
R21149 CSoutput.n349 CSoutput.t129 2.82907
R21150 CSoutput.n408 CSoutput.t177 2.82907
R21151 CSoutput.n408 CSoutput.t188 2.82907
R21152 CSoutput.n409 CSoutput.t191 2.82907
R21153 CSoutput.n409 CSoutput.t168 2.82907
R21154 CSoutput.n411 CSoutput.t172 2.82907
R21155 CSoutput.n411 CSoutput.t183 2.82907
R21156 CSoutput.n413 CSoutput.t130 2.82907
R21157 CSoutput.n413 CSoutput.t162 2.82907
R21158 CSoutput.n415 CSoutput.t167 2.82907
R21159 CSoutput.n415 CSoutput.t178 2.82907
R21160 CSoutput.n417 CSoutput.t184 2.82907
R21161 CSoutput.n417 CSoutput.t171 2.82907
R21162 CSoutput.n396 CSoutput.t148 2.82907
R21163 CSoutput.n396 CSoutput.t165 2.82907
R21164 CSoutput.n397 CSoutput.t166 2.82907
R21165 CSoutput.n397 CSoutput.t157 2.82907
R21166 CSoutput.n399 CSoutput.t156 2.82907
R21167 CSoutput.n399 CSoutput.t149 2.82907
R21168 CSoutput.n401 CSoutput.t144 2.82907
R21169 CSoutput.n401 CSoutput.t136 2.82907
R21170 CSoutput.n403 CSoutput.t137 2.82907
R21171 CSoutput.n403 CSoutput.t158 2.82907
R21172 CSoutput.n405 CSoutput.t160 2.82907
R21173 CSoutput.n405 CSoutput.t123 2.82907
R21174 CSoutput.n385 CSoutput.t161 2.82907
R21175 CSoutput.n385 CSoutput.t125 2.82907
R21176 CSoutput.n386 CSoutput.t145 2.82907
R21177 CSoutput.n386 CSoutput.t187 2.82907
R21178 CSoutput.n388 CSoutput.t126 2.82907
R21179 CSoutput.n388 CSoutput.t175 2.82907
R21180 CSoutput.n390 CSoutput.t174 2.82907
R21181 CSoutput.n390 CSoutput.t163 2.82907
R21182 CSoutput.n392 CSoutput.t176 2.82907
R21183 CSoutput.n392 CSoutput.t147 2.82907
R21184 CSoutput.n394 CSoutput.t170 2.82907
R21185 CSoutput.n394 CSoutput.t181 2.82907
R21186 CSoutput.n348 CSoutput.n138 2.57547
R21187 CSoutput.n75 CSoutput.n1 2.45513
R21188 CSoutput.n229 CSoutput.n227 2.251
R21189 CSoutput.n229 CSoutput.n226 2.251
R21190 CSoutput.n229 CSoutput.n225 2.251
R21191 CSoutput.n229 CSoutput.n224 2.251
R21192 CSoutput.n198 CSoutput.n197 2.251
R21193 CSoutput.n198 CSoutput.n196 2.251
R21194 CSoutput.n198 CSoutput.n195 2.251
R21195 CSoutput.n198 CSoutput.n194 2.251
R21196 CSoutput.n271 CSoutput.n270 2.251
R21197 CSoutput.n236 CSoutput.n234 2.251
R21198 CSoutput.n236 CSoutput.n233 2.251
R21199 CSoutput.n236 CSoutput.n232 2.251
R21200 CSoutput.n254 CSoutput.n236 2.251
R21201 CSoutput.n242 CSoutput.n241 2.251
R21202 CSoutput.n242 CSoutput.n240 2.251
R21203 CSoutput.n242 CSoutput.n239 2.251
R21204 CSoutput.n242 CSoutput.n238 2.251
R21205 CSoutput.n268 CSoutput.n208 2.251
R21206 CSoutput.n263 CSoutput.n261 2.251
R21207 CSoutput.n263 CSoutput.n260 2.251
R21208 CSoutput.n263 CSoutput.n259 2.251
R21209 CSoutput.n263 CSoutput.n258 2.251
R21210 CSoutput.n164 CSoutput.n163 2.251
R21211 CSoutput.n164 CSoutput.n162 2.251
R21212 CSoutput.n164 CSoutput.n161 2.251
R21213 CSoutput.n164 CSoutput.n160 2.251
R21214 CSoutput.n281 CSoutput.n280 2.251
R21215 CSoutput.n198 CSoutput.n178 2.2505
R21216 CSoutput.n193 CSoutput.n178 2.2505
R21217 CSoutput.n191 CSoutput.n178 2.2505
R21218 CSoutput.n190 CSoutput.n178 2.2505
R21219 CSoutput.n275 CSoutput.n178 2.2505
R21220 CSoutput.n273 CSoutput.n178 2.2505
R21221 CSoutput.n271 CSoutput.n178 2.2505
R21222 CSoutput.n201 CSoutput.n178 2.2505
R21223 CSoutput.n200 CSoutput.n178 2.2505
R21224 CSoutput.n204 CSoutput.n178 2.2505
R21225 CSoutput.n203 CSoutput.n178 2.2505
R21226 CSoutput.n186 CSoutput.n178 2.2505
R21227 CSoutput.n278 CSoutput.n178 2.2505
R21228 CSoutput.n278 CSoutput.n277 2.2505
R21229 CSoutput.n242 CSoutput.n213 2.2505
R21230 CSoutput.n223 CSoutput.n213 2.2505
R21231 CSoutput.n244 CSoutput.n213 2.2505
R21232 CSoutput.n222 CSoutput.n213 2.2505
R21233 CSoutput.n246 CSoutput.n213 2.2505
R21234 CSoutput.n213 CSoutput.n207 2.2505
R21235 CSoutput.n268 CSoutput.n213 2.2505
R21236 CSoutput.n266 CSoutput.n213 2.2505
R21237 CSoutput.n248 CSoutput.n213 2.2505
R21238 CSoutput.n220 CSoutput.n213 2.2505
R21239 CSoutput.n250 CSoutput.n213 2.2505
R21240 CSoutput.n219 CSoutput.n213 2.2505
R21241 CSoutput.n264 CSoutput.n213 2.2505
R21242 CSoutput.n264 CSoutput.n217 2.2505
R21243 CSoutput.n164 CSoutput.n144 2.2505
R21244 CSoutput.n159 CSoutput.n144 2.2505
R21245 CSoutput.n157 CSoutput.n144 2.2505
R21246 CSoutput.n156 CSoutput.n144 2.2505
R21247 CSoutput.n285 CSoutput.n144 2.2505
R21248 CSoutput.n283 CSoutput.n144 2.2505
R21249 CSoutput.n281 CSoutput.n144 2.2505
R21250 CSoutput.n167 CSoutput.n144 2.2505
R21251 CSoutput.n166 CSoutput.n144 2.2505
R21252 CSoutput.n170 CSoutput.n144 2.2505
R21253 CSoutput.n169 CSoutput.n144 2.2505
R21254 CSoutput.n152 CSoutput.n144 2.2505
R21255 CSoutput.n288 CSoutput.n144 2.2505
R21256 CSoutput.n288 CSoutput.n287 2.2505
R21257 CSoutput.n206 CSoutput.n199 2.25024
R21258 CSoutput.n206 CSoutput.n192 2.25024
R21259 CSoutput.n274 CSoutput.n206 2.25024
R21260 CSoutput.n206 CSoutput.n202 2.25024
R21261 CSoutput.n206 CSoutput.n205 2.25024
R21262 CSoutput.n206 CSoutput.n173 2.25024
R21263 CSoutput.n256 CSoutput.n253 2.25024
R21264 CSoutput.n256 CSoutput.n252 2.25024
R21265 CSoutput.n256 CSoutput.n251 2.25024
R21266 CSoutput.n256 CSoutput.n218 2.25024
R21267 CSoutput.n256 CSoutput.n255 2.25024
R21268 CSoutput.n257 CSoutput.n256 2.25024
R21269 CSoutput.n172 CSoutput.n165 2.25024
R21270 CSoutput.n172 CSoutput.n158 2.25024
R21271 CSoutput.n284 CSoutput.n172 2.25024
R21272 CSoutput.n172 CSoutput.n168 2.25024
R21273 CSoutput.n172 CSoutput.n171 2.25024
R21274 CSoutput.n172 CSoutput.n139 2.25024
R21275 CSoutput.n273 CSoutput.n183 1.50111
R21276 CSoutput.n221 CSoutput.n207 1.50111
R21277 CSoutput.n283 CSoutput.n149 1.50111
R21278 CSoutput.n229 CSoutput.n228 1.501
R21279 CSoutput.n236 CSoutput.n235 1.501
R21280 CSoutput.n263 CSoutput.n262 1.501
R21281 CSoutput.n277 CSoutput.n188 1.12536
R21282 CSoutput.n277 CSoutput.n189 1.12536
R21283 CSoutput.n277 CSoutput.n276 1.12536
R21284 CSoutput.n237 CSoutput.n217 1.12536
R21285 CSoutput.n243 CSoutput.n217 1.12536
R21286 CSoutput.n245 CSoutput.n217 1.12536
R21287 CSoutput.n287 CSoutput.n154 1.12536
R21288 CSoutput.n287 CSoutput.n155 1.12536
R21289 CSoutput.n287 CSoutput.n286 1.12536
R21290 CSoutput.n277 CSoutput.n184 1.12536
R21291 CSoutput.n277 CSoutput.n185 1.12536
R21292 CSoutput.n277 CSoutput.n187 1.12536
R21293 CSoutput.n267 CSoutput.n217 1.12536
R21294 CSoutput.n247 CSoutput.n217 1.12536
R21295 CSoutput.n249 CSoutput.n217 1.12536
R21296 CSoutput.n287 CSoutput.n150 1.12536
R21297 CSoutput.n287 CSoutput.n151 1.12536
R21298 CSoutput.n287 CSoutput.n153 1.12536
R21299 CSoutput.n31 CSoutput.n30 0.669944
R21300 CSoutput.n62 CSoutput.n61 0.669944
R21301 CSoutput.n376 CSoutput.n374 0.573776
R21302 CSoutput.n378 CSoutput.n376 0.573776
R21303 CSoutput.n380 CSoutput.n378 0.573776
R21304 CSoutput.n382 CSoutput.n380 0.573776
R21305 CSoutput.n364 CSoutput.n362 0.573776
R21306 CSoutput.n366 CSoutput.n364 0.573776
R21307 CSoutput.n368 CSoutput.n366 0.573776
R21308 CSoutput.n370 CSoutput.n368 0.573776
R21309 CSoutput.n353 CSoutput.n351 0.573776
R21310 CSoutput.n355 CSoutput.n353 0.573776
R21311 CSoutput.n357 CSoutput.n355 0.573776
R21312 CSoutput.n359 CSoutput.n357 0.573776
R21313 CSoutput.n418 CSoutput.n416 0.573776
R21314 CSoutput.n416 CSoutput.n414 0.573776
R21315 CSoutput.n414 CSoutput.n412 0.573776
R21316 CSoutput.n412 CSoutput.n410 0.573776
R21317 CSoutput.n406 CSoutput.n404 0.573776
R21318 CSoutput.n404 CSoutput.n402 0.573776
R21319 CSoutput.n402 CSoutput.n400 0.573776
R21320 CSoutput.n400 CSoutput.n398 0.573776
R21321 CSoutput.n395 CSoutput.n393 0.573776
R21322 CSoutput.n393 CSoutput.n391 0.573776
R21323 CSoutput.n391 CSoutput.n389 0.573776
R21324 CSoutput.n389 CSoutput.n387 0.573776
R21325 CSoutput.n421 CSoutput.n288 0.53442
R21326 CSoutput.n332 CSoutput.n330 0.358259
R21327 CSoutput.n334 CSoutput.n332 0.358259
R21328 CSoutput.n336 CSoutput.n334 0.358259
R21329 CSoutput.n338 CSoutput.n336 0.358259
R21330 CSoutput.n340 CSoutput.n338 0.358259
R21331 CSoutput.n342 CSoutput.n340 0.358259
R21332 CSoutput.n344 CSoutput.n342 0.358259
R21333 CSoutput.n346 CSoutput.n344 0.358259
R21334 CSoutput.n312 CSoutput.n310 0.358259
R21335 CSoutput.n314 CSoutput.n312 0.358259
R21336 CSoutput.n316 CSoutput.n314 0.358259
R21337 CSoutput.n318 CSoutput.n316 0.358259
R21338 CSoutput.n320 CSoutput.n318 0.358259
R21339 CSoutput.n322 CSoutput.n320 0.358259
R21340 CSoutput.n324 CSoutput.n322 0.358259
R21341 CSoutput.n326 CSoutput.n324 0.358259
R21342 CSoutput.n293 CSoutput.n291 0.358259
R21343 CSoutput.n295 CSoutput.n293 0.358259
R21344 CSoutput.n297 CSoutput.n295 0.358259
R21345 CSoutput.n299 CSoutput.n297 0.358259
R21346 CSoutput.n301 CSoutput.n299 0.358259
R21347 CSoutput.n303 CSoutput.n301 0.358259
R21348 CSoutput.n305 CSoutput.n303 0.358259
R21349 CSoutput.n307 CSoutput.n305 0.358259
R21350 CSoutput.n136 CSoutput.n134 0.358259
R21351 CSoutput.n134 CSoutput.n132 0.358259
R21352 CSoutput.n132 CSoutput.n130 0.358259
R21353 CSoutput.n130 CSoutput.n128 0.358259
R21354 CSoutput.n128 CSoutput.n126 0.358259
R21355 CSoutput.n126 CSoutput.n124 0.358259
R21356 CSoutput.n124 CSoutput.n122 0.358259
R21357 CSoutput.n122 CSoutput.n120 0.358259
R21358 CSoutput.n116 CSoutput.n114 0.358259
R21359 CSoutput.n114 CSoutput.n112 0.358259
R21360 CSoutput.n112 CSoutput.n110 0.358259
R21361 CSoutput.n110 CSoutput.n108 0.358259
R21362 CSoutput.n108 CSoutput.n106 0.358259
R21363 CSoutput.n106 CSoutput.n104 0.358259
R21364 CSoutput.n104 CSoutput.n102 0.358259
R21365 CSoutput.n102 CSoutput.n100 0.358259
R21366 CSoutput.n97 CSoutput.n95 0.358259
R21367 CSoutput.n95 CSoutput.n93 0.358259
R21368 CSoutput.n93 CSoutput.n91 0.358259
R21369 CSoutput.n91 CSoutput.n89 0.358259
R21370 CSoutput.n89 CSoutput.n87 0.358259
R21371 CSoutput.n87 CSoutput.n85 0.358259
R21372 CSoutput.n85 CSoutput.n83 0.358259
R21373 CSoutput.n83 CSoutput.n81 0.358259
R21374 CSoutput.n21 CSoutput.n20 0.169105
R21375 CSoutput.n21 CSoutput.n16 0.169105
R21376 CSoutput.n26 CSoutput.n16 0.169105
R21377 CSoutput.n27 CSoutput.n26 0.169105
R21378 CSoutput.n27 CSoutput.n14 0.169105
R21379 CSoutput.n32 CSoutput.n14 0.169105
R21380 CSoutput.n33 CSoutput.n32 0.169105
R21381 CSoutput.n34 CSoutput.n33 0.169105
R21382 CSoutput.n34 CSoutput.n12 0.169105
R21383 CSoutput.n39 CSoutput.n12 0.169105
R21384 CSoutput.n40 CSoutput.n39 0.169105
R21385 CSoutput.n40 CSoutput.n10 0.169105
R21386 CSoutput.n45 CSoutput.n10 0.169105
R21387 CSoutput.n46 CSoutput.n45 0.169105
R21388 CSoutput.n47 CSoutput.n46 0.169105
R21389 CSoutput.n47 CSoutput.n8 0.169105
R21390 CSoutput.n52 CSoutput.n8 0.169105
R21391 CSoutput.n53 CSoutput.n52 0.169105
R21392 CSoutput.n53 CSoutput.n6 0.169105
R21393 CSoutput.n58 CSoutput.n6 0.169105
R21394 CSoutput.n59 CSoutput.n58 0.169105
R21395 CSoutput.n60 CSoutput.n59 0.169105
R21396 CSoutput.n60 CSoutput.n4 0.169105
R21397 CSoutput.n66 CSoutput.n4 0.169105
R21398 CSoutput.n67 CSoutput.n66 0.169105
R21399 CSoutput.n68 CSoutput.n67 0.169105
R21400 CSoutput.n68 CSoutput.n2 0.169105
R21401 CSoutput.n73 CSoutput.n2 0.169105
R21402 CSoutput.n74 CSoutput.n73 0.169105
R21403 CSoutput.n74 CSoutput.n0 0.169105
R21404 CSoutput.n78 CSoutput.n0 0.169105
R21405 CSoutput.n231 CSoutput.n230 0.0910737
R21406 CSoutput.n282 CSoutput.n279 0.0723685
R21407 CSoutput.n236 CSoutput.n231 0.0522944
R21408 CSoutput.n279 CSoutput.n278 0.0499135
R21409 CSoutput.n230 CSoutput.n229 0.0499135
R21410 CSoutput.n264 CSoutput.n263 0.0464294
R21411 CSoutput.n272 CSoutput.n269 0.0391444
R21412 CSoutput.n231 CSoutput.t211 0.023435
R21413 CSoutput.n279 CSoutput.t192 0.02262
R21414 CSoutput.n230 CSoutput.t194 0.02262
R21415 CSoutput CSoutput.n421 0.0052
R21416 CSoutput.n201 CSoutput.n184 0.00365111
R21417 CSoutput.n204 CSoutput.n185 0.00365111
R21418 CSoutput.n187 CSoutput.n186 0.00365111
R21419 CSoutput.n229 CSoutput.n188 0.00365111
R21420 CSoutput.n193 CSoutput.n189 0.00365111
R21421 CSoutput.n276 CSoutput.n190 0.00365111
R21422 CSoutput.n267 CSoutput.n266 0.00365111
R21423 CSoutput.n247 CSoutput.n220 0.00365111
R21424 CSoutput.n249 CSoutput.n219 0.00365111
R21425 CSoutput.n237 CSoutput.n236 0.00365111
R21426 CSoutput.n243 CSoutput.n223 0.00365111
R21427 CSoutput.n245 CSoutput.n222 0.00365111
R21428 CSoutput.n167 CSoutput.n150 0.00365111
R21429 CSoutput.n170 CSoutput.n151 0.00365111
R21430 CSoutput.n153 CSoutput.n152 0.00365111
R21431 CSoutput.n263 CSoutput.n154 0.00365111
R21432 CSoutput.n159 CSoutput.n155 0.00365111
R21433 CSoutput.n286 CSoutput.n156 0.00365111
R21434 CSoutput.n198 CSoutput.n188 0.00340054
R21435 CSoutput.n191 CSoutput.n189 0.00340054
R21436 CSoutput.n276 CSoutput.n275 0.00340054
R21437 CSoutput.n271 CSoutput.n184 0.00340054
R21438 CSoutput.n200 CSoutput.n185 0.00340054
R21439 CSoutput.n203 CSoutput.n187 0.00340054
R21440 CSoutput.n242 CSoutput.n237 0.00340054
R21441 CSoutput.n244 CSoutput.n243 0.00340054
R21442 CSoutput.n246 CSoutput.n245 0.00340054
R21443 CSoutput.n268 CSoutput.n267 0.00340054
R21444 CSoutput.n248 CSoutput.n247 0.00340054
R21445 CSoutput.n250 CSoutput.n249 0.00340054
R21446 CSoutput.n164 CSoutput.n154 0.00340054
R21447 CSoutput.n157 CSoutput.n155 0.00340054
R21448 CSoutput.n286 CSoutput.n285 0.00340054
R21449 CSoutput.n281 CSoutput.n150 0.00340054
R21450 CSoutput.n166 CSoutput.n151 0.00340054
R21451 CSoutput.n169 CSoutput.n153 0.00340054
R21452 CSoutput.n199 CSoutput.n193 0.00252698
R21453 CSoutput.n192 CSoutput.n190 0.00252698
R21454 CSoutput.n274 CSoutput.n273 0.00252698
R21455 CSoutput.n202 CSoutput.n200 0.00252698
R21456 CSoutput.n205 CSoutput.n203 0.00252698
R21457 CSoutput.n278 CSoutput.n173 0.00252698
R21458 CSoutput.n199 CSoutput.n198 0.00252698
R21459 CSoutput.n192 CSoutput.n191 0.00252698
R21460 CSoutput.n275 CSoutput.n274 0.00252698
R21461 CSoutput.n202 CSoutput.n201 0.00252698
R21462 CSoutput.n205 CSoutput.n204 0.00252698
R21463 CSoutput.n186 CSoutput.n173 0.00252698
R21464 CSoutput.n253 CSoutput.n223 0.00252698
R21465 CSoutput.n252 CSoutput.n222 0.00252698
R21466 CSoutput.n251 CSoutput.n207 0.00252698
R21467 CSoutput.n248 CSoutput.n218 0.00252698
R21468 CSoutput.n255 CSoutput.n250 0.00252698
R21469 CSoutput.n264 CSoutput.n257 0.00252698
R21470 CSoutput.n253 CSoutput.n242 0.00252698
R21471 CSoutput.n252 CSoutput.n244 0.00252698
R21472 CSoutput.n251 CSoutput.n246 0.00252698
R21473 CSoutput.n266 CSoutput.n218 0.00252698
R21474 CSoutput.n255 CSoutput.n220 0.00252698
R21475 CSoutput.n257 CSoutput.n219 0.00252698
R21476 CSoutput.n165 CSoutput.n159 0.00252698
R21477 CSoutput.n158 CSoutput.n156 0.00252698
R21478 CSoutput.n284 CSoutput.n283 0.00252698
R21479 CSoutput.n168 CSoutput.n166 0.00252698
R21480 CSoutput.n171 CSoutput.n169 0.00252698
R21481 CSoutput.n288 CSoutput.n139 0.00252698
R21482 CSoutput.n165 CSoutput.n164 0.00252698
R21483 CSoutput.n158 CSoutput.n157 0.00252698
R21484 CSoutput.n285 CSoutput.n284 0.00252698
R21485 CSoutput.n168 CSoutput.n167 0.00252698
R21486 CSoutput.n171 CSoutput.n170 0.00252698
R21487 CSoutput.n152 CSoutput.n139 0.00252698
R21488 CSoutput.n273 CSoutput.n272 0.0020275
R21489 CSoutput.n272 CSoutput.n271 0.0020275
R21490 CSoutput.n269 CSoutput.n207 0.0020275
R21491 CSoutput.n269 CSoutput.n268 0.0020275
R21492 CSoutput.n283 CSoutput.n282 0.0020275
R21493 CSoutput.n282 CSoutput.n281 0.0020275
R21494 CSoutput.n183 CSoutput.n182 0.00166668
R21495 CSoutput.n265 CSoutput.n221 0.00166668
R21496 CSoutput.n149 CSoutput.n148 0.00166668
R21497 CSoutput.n287 CSoutput.n149 0.00133328
R21498 CSoutput.n221 CSoutput.n217 0.00133328
R21499 CSoutput.n277 CSoutput.n183 0.00133328
R21500 CSoutput.n280 CSoutput.n172 0.001
R21501 CSoutput.n258 CSoutput.n172 0.001
R21502 CSoutput.n160 CSoutput.n140 0.001
R21503 CSoutput.n259 CSoutput.n140 0.001
R21504 CSoutput.n161 CSoutput.n141 0.001
R21505 CSoutput.n260 CSoutput.n141 0.001
R21506 CSoutput.n162 CSoutput.n142 0.001
R21507 CSoutput.n261 CSoutput.n142 0.001
R21508 CSoutput.n163 CSoutput.n143 0.001
R21509 CSoutput.n262 CSoutput.n143 0.001
R21510 CSoutput.n256 CSoutput.n208 0.001
R21511 CSoutput.n256 CSoutput.n254 0.001
R21512 CSoutput.n238 CSoutput.n209 0.001
R21513 CSoutput.n232 CSoutput.n209 0.001
R21514 CSoutput.n239 CSoutput.n210 0.001
R21515 CSoutput.n233 CSoutput.n210 0.001
R21516 CSoutput.n240 CSoutput.n211 0.001
R21517 CSoutput.n234 CSoutput.n211 0.001
R21518 CSoutput.n241 CSoutput.n212 0.001
R21519 CSoutput.n235 CSoutput.n212 0.001
R21520 CSoutput.n270 CSoutput.n206 0.001
R21521 CSoutput.n224 CSoutput.n206 0.001
R21522 CSoutput.n194 CSoutput.n174 0.001
R21523 CSoutput.n225 CSoutput.n174 0.001
R21524 CSoutput.n195 CSoutput.n175 0.001
R21525 CSoutput.n226 CSoutput.n175 0.001
R21526 CSoutput.n196 CSoutput.n176 0.001
R21527 CSoutput.n227 CSoutput.n176 0.001
R21528 CSoutput.n197 CSoutput.n177 0.001
R21529 CSoutput.n228 CSoutput.n177 0.001
R21530 CSoutput.n228 CSoutput.n178 0.001
R21531 CSoutput.n227 CSoutput.n179 0.001
R21532 CSoutput.n226 CSoutput.n180 0.001
R21533 CSoutput.n225 CSoutput.t210 0.001
R21534 CSoutput.n224 CSoutput.n181 0.001
R21535 CSoutput.n197 CSoutput.n179 0.001
R21536 CSoutput.n196 CSoutput.n180 0.001
R21537 CSoutput.n195 CSoutput.t210 0.001
R21538 CSoutput.n194 CSoutput.n181 0.001
R21539 CSoutput.n270 CSoutput.n182 0.001
R21540 CSoutput.n235 CSoutput.n213 0.001
R21541 CSoutput.n234 CSoutput.n214 0.001
R21542 CSoutput.n233 CSoutput.n215 0.001
R21543 CSoutput.n232 CSoutput.t203 0.001
R21544 CSoutput.n254 CSoutput.n216 0.001
R21545 CSoutput.n241 CSoutput.n214 0.001
R21546 CSoutput.n240 CSoutput.n215 0.001
R21547 CSoutput.n239 CSoutput.t203 0.001
R21548 CSoutput.n238 CSoutput.n216 0.001
R21549 CSoutput.n265 CSoutput.n208 0.001
R21550 CSoutput.n262 CSoutput.n144 0.001
R21551 CSoutput.n261 CSoutput.n145 0.001
R21552 CSoutput.n260 CSoutput.n146 0.001
R21553 CSoutput.n259 CSoutput.t202 0.001
R21554 CSoutput.n258 CSoutput.n147 0.001
R21555 CSoutput.n163 CSoutput.n145 0.001
R21556 CSoutput.n162 CSoutput.n146 0.001
R21557 CSoutput.n161 CSoutput.t202 0.001
R21558 CSoutput.n160 CSoutput.n147 0.001
R21559 CSoutput.n280 CSoutput.n148 0.001
R21560 a_n1986_13878.n3 a_n1986_13878.t30 539.01
R21561 a_n1986_13878.n91 a_n1986_13878.t22 512.366
R21562 a_n1986_13878.n90 a_n1986_13878.t10 512.366
R21563 a_n1986_13878.n52 a_n1986_13878.t12 512.366
R21564 a_n1986_13878.n89 a_n1986_13878.t26 512.366
R21565 a_n1986_13878.n7 a_n1986_13878.t66 539.01
R21566 a_n1986_13878.n80 a_n1986_13878.t49 512.366
R21567 a_n1986_13878.n79 a_n1986_13878.t53 512.366
R21568 a_n1986_13878.n53 a_n1986_13878.t43 512.366
R21569 a_n1986_13878.n78 a_n1986_13878.t58 512.366
R21570 a_n1986_13878.n20 a_n1986_13878.t18 539.01
R21571 a_n1986_13878.n61 a_n1986_13878.t20 512.366
R21572 a_n1986_13878.n62 a_n1986_13878.t24 512.366
R21573 a_n1986_13878.n56 a_n1986_13878.t16 512.366
R21574 a_n1986_13878.n63 a_n1986_13878.t32 512.366
R21575 a_n1986_13878.n24 a_n1986_13878.t61 539.01
R21576 a_n1986_13878.n58 a_n1986_13878.t62 512.366
R21577 a_n1986_13878.n59 a_n1986_13878.t41 512.366
R21578 a_n1986_13878.n57 a_n1986_13878.t48 512.366
R21579 a_n1986_13878.n60 a_n1986_13878.t57 512.366
R21580 a_n1986_13878.n75 a_n1986_13878.t55 512.366
R21581 a_n1986_13878.n65 a_n1986_13878.t46 512.366
R21582 a_n1986_13878.n76 a_n1986_13878.t40 512.366
R21583 a_n1986_13878.n73 a_n1986_13878.t63 512.366
R21584 a_n1986_13878.n66 a_n1986_13878.t52 512.366
R21585 a_n1986_13878.n74 a_n1986_13878.t51 512.366
R21586 a_n1986_13878.n71 a_n1986_13878.t59 512.366
R21587 a_n1986_13878.n67 a_n1986_13878.t44 512.366
R21588 a_n1986_13878.n72 a_n1986_13878.t45 512.366
R21589 a_n1986_13878.n69 a_n1986_13878.t47 512.366
R21590 a_n1986_13878.n68 a_n1986_13878.t56 512.366
R21591 a_n1986_13878.n70 a_n1986_13878.t67 512.366
R21592 a_n1986_13878.n51 a_n1986_13878.n0 70.3058
R21593 a_n1986_13878.n48 a_n1986_13878.n5 70.3058
R21594 a_n1986_13878.n17 a_n1986_13878.n37 70.3058
R21595 a_n1986_13878.n21 a_n1986_13878.n34 70.3058
R21596 a_n1986_13878.n33 a_n1986_13878.n22 70.1674
R21597 a_n1986_13878.n33 a_n1986_13878.n57 20.9683
R21598 a_n1986_13878.n22 a_n1986_13878.n32 75.0448
R21599 a_n1986_13878.n59 a_n1986_13878.n32 11.2134
R21600 a_n1986_13878.n23 a_n1986_13878.n24 44.8194
R21601 a_n1986_13878.n36 a_n1986_13878.n18 70.1674
R21602 a_n1986_13878.n36 a_n1986_13878.n56 20.9683
R21603 a_n1986_13878.n18 a_n1986_13878.n35 75.0448
R21604 a_n1986_13878.n62 a_n1986_13878.n35 11.2134
R21605 a_n1986_13878.n19 a_n1986_13878.n20 44.8194
R21606 a_n1986_13878.n8 a_n1986_13878.n45 70.1674
R21607 a_n1986_13878.n10 a_n1986_13878.n43 70.1674
R21608 a_n1986_13878.n12 a_n1986_13878.n41 70.1674
R21609 a_n1986_13878.n15 a_n1986_13878.n39 70.1674
R21610 a_n1986_13878.n70 a_n1986_13878.n39 20.9683
R21611 a_n1986_13878.n38 a_n1986_13878.n16 75.0448
R21612 a_n1986_13878.n38 a_n1986_13878.n68 11.2134
R21613 a_n1986_13878.n16 a_n1986_13878.n69 161.3
R21614 a_n1986_13878.n72 a_n1986_13878.n41 20.9683
R21615 a_n1986_13878.n40 a_n1986_13878.n13 75.0448
R21616 a_n1986_13878.n40 a_n1986_13878.n67 11.2134
R21617 a_n1986_13878.n13 a_n1986_13878.n71 161.3
R21618 a_n1986_13878.n74 a_n1986_13878.n43 20.9683
R21619 a_n1986_13878.n42 a_n1986_13878.n11 75.0448
R21620 a_n1986_13878.n42 a_n1986_13878.n66 11.2134
R21621 a_n1986_13878.n11 a_n1986_13878.n73 161.3
R21622 a_n1986_13878.n76 a_n1986_13878.n45 20.9683
R21623 a_n1986_13878.n44 a_n1986_13878.n9 75.0448
R21624 a_n1986_13878.n44 a_n1986_13878.n65 11.2134
R21625 a_n1986_13878.n9 a_n1986_13878.n75 161.3
R21626 a_n1986_13878.n6 a_n1986_13878.n47 70.1674
R21627 a_n1986_13878.n47 a_n1986_13878.n53 20.9683
R21628 a_n1986_13878.n46 a_n1986_13878.n6 75.0448
R21629 a_n1986_13878.n79 a_n1986_13878.n46 11.2134
R21630 a_n1986_13878.n4 a_n1986_13878.n7 44.8194
R21631 a_n1986_13878.n2 a_n1986_13878.n50 70.1674
R21632 a_n1986_13878.n50 a_n1986_13878.n52 20.9683
R21633 a_n1986_13878.n49 a_n1986_13878.n2 75.0448
R21634 a_n1986_13878.n90 a_n1986_13878.n49 11.2134
R21635 a_n1986_13878.n1 a_n1986_13878.n3 44.8194
R21636 a_n1986_13878.n30 a_n1986_13878.n87 81.2902
R21637 a_n1986_13878.n31 a_n1986_13878.n83 81.2902
R21638 a_n1986_13878.n31 a_n1986_13878.n81 81.2902
R21639 a_n1986_13878.n30 a_n1986_13878.n88 80.9324
R21640 a_n1986_13878.n30 a_n1986_13878.n86 80.9324
R21641 a_n1986_13878.n29 a_n1986_13878.n85 80.9324
R21642 a_n1986_13878.n31 a_n1986_13878.n84 80.9324
R21643 a_n1986_13878.n31 a_n1986_13878.n82 80.9324
R21644 a_n1986_13878.n28 a_n1986_13878.t15 74.6477
R21645 a_n1986_13878.n25 a_n1986_13878.t19 74.6477
R21646 a_n1986_13878.n27 a_n1986_13878.t31 74.2899
R21647 a_n1986_13878.n26 a_n1986_13878.t29 74.2897
R21648 a_n1986_13878.n28 a_n1986_13878.n93 70.6783
R21649 a_n1986_13878.n26 a_n1986_13878.n55 70.6783
R21650 a_n1986_13878.n25 a_n1986_13878.n54 70.6783
R21651 a_n1986_13878.n94 a_n1986_13878.n28 70.6782
R21652 a_n1986_13878.n91 a_n1986_13878.n90 48.2005
R21653 a_n1986_13878.n89 a_n1986_13878.n50 20.9683
R21654 a_n1986_13878.n80 a_n1986_13878.n79 48.2005
R21655 a_n1986_13878.n78 a_n1986_13878.n47 20.9683
R21656 a_n1986_13878.n62 a_n1986_13878.n61 48.2005
R21657 a_n1986_13878.n63 a_n1986_13878.n36 20.9683
R21658 a_n1986_13878.n59 a_n1986_13878.n58 48.2005
R21659 a_n1986_13878.n60 a_n1986_13878.n33 20.9683
R21660 a_n1986_13878.n75 a_n1986_13878.n65 48.2005
R21661 a_n1986_13878.t60 a_n1986_13878.n45 533.335
R21662 a_n1986_13878.n73 a_n1986_13878.n66 48.2005
R21663 a_n1986_13878.t65 a_n1986_13878.n43 533.335
R21664 a_n1986_13878.n71 a_n1986_13878.n67 48.2005
R21665 a_n1986_13878.t54 a_n1986_13878.n41 533.335
R21666 a_n1986_13878.n69 a_n1986_13878.n68 48.2005
R21667 a_n1986_13878.t50 a_n1986_13878.n39 533.335
R21668 a_n1986_13878.n51 a_n1986_13878.t14 533.058
R21669 a_n1986_13878.n48 a_n1986_13878.t64 533.058
R21670 a_n1986_13878.t28 a_n1986_13878.n37 533.058
R21671 a_n1986_13878.t42 a_n1986_13878.n34 533.058
R21672 a_n1986_13878.n49 a_n1986_13878.n52 35.3134
R21673 a_n1986_13878.n46 a_n1986_13878.n53 35.3134
R21674 a_n1986_13878.n56 a_n1986_13878.n35 35.3134
R21675 a_n1986_13878.n57 a_n1986_13878.n32 35.3134
R21676 a_n1986_13878.n76 a_n1986_13878.n44 35.3134
R21677 a_n1986_13878.n74 a_n1986_13878.n42 35.3134
R21678 a_n1986_13878.n72 a_n1986_13878.n40 35.3134
R21679 a_n1986_13878.n70 a_n1986_13878.n38 35.3134
R21680 a_n1986_13878.n29 a_n1986_13878.n31 31.0592
R21681 a_n1986_13878.n0 a_n1986_13878.n30 23.891
R21682 a_n1986_13878.n23 a_n1986_13878.n14 12.046
R21683 a_n1986_13878.n5 a_n1986_13878.n77 11.8414
R21684 a_n1986_13878.n92 a_n1986_13878.n1 10.5365
R21685 a_n1986_13878.n64 a_n1986_13878.n26 9.50122
R21686 a_n1986_13878.n16 a_n1986_13878.n14 7.47588
R21687 a_n1986_13878.n77 a_n1986_13878.n8 7.47588
R21688 a_n1986_13878.n64 a_n1986_13878.n17 6.70126
R21689 a_n1986_13878.n27 a_n1986_13878.n92 5.65783
R21690 a_n1986_13878.n77 a_n1986_13878.n64 5.3452
R21691 a_n1986_13878.n19 a_n1986_13878.n21 3.95126
R21692 a_n1986_13878.n93 a_n1986_13878.t13 3.61217
R21693 a_n1986_13878.n93 a_n1986_13878.t27 3.61217
R21694 a_n1986_13878.n55 a_n1986_13878.t17 3.61217
R21695 a_n1986_13878.n55 a_n1986_13878.t33 3.61217
R21696 a_n1986_13878.n54 a_n1986_13878.t21 3.61217
R21697 a_n1986_13878.n54 a_n1986_13878.t25 3.61217
R21698 a_n1986_13878.n94 a_n1986_13878.t23 3.61217
R21699 a_n1986_13878.t11 a_n1986_13878.n94 3.61217
R21700 a_n1986_13878.n0 a_n1986_13878.n4 3.42095
R21701 a_n1986_13878.n87 a_n1986_13878.t5 2.82907
R21702 a_n1986_13878.n87 a_n1986_13878.t0 2.82907
R21703 a_n1986_13878.n88 a_n1986_13878.t35 2.82907
R21704 a_n1986_13878.n88 a_n1986_13878.t9 2.82907
R21705 a_n1986_13878.n86 a_n1986_13878.t38 2.82907
R21706 a_n1986_13878.n86 a_n1986_13878.t37 2.82907
R21707 a_n1986_13878.n85 a_n1986_13878.t7 2.82907
R21708 a_n1986_13878.n85 a_n1986_13878.t1 2.82907
R21709 a_n1986_13878.n83 a_n1986_13878.t8 2.82907
R21710 a_n1986_13878.n83 a_n1986_13878.t39 2.82907
R21711 a_n1986_13878.n84 a_n1986_13878.t34 2.82907
R21712 a_n1986_13878.n84 a_n1986_13878.t36 2.82907
R21713 a_n1986_13878.n82 a_n1986_13878.t4 2.82907
R21714 a_n1986_13878.n82 a_n1986_13878.t6 2.82907
R21715 a_n1986_13878.n81 a_n1986_13878.t3 2.82907
R21716 a_n1986_13878.n81 a_n1986_13878.t2 2.82907
R21717 a_n1986_13878.n92 a_n1986_13878.n14 1.30542
R21718 a_n1986_13878.n11 a_n1986_13878.n12 1.04595
R21719 a_n1986_13878.n3 a_n1986_13878.n91 13.657
R21720 a_n1986_13878.n89 a_n1986_13878.n51 21.4216
R21721 a_n1986_13878.n7 a_n1986_13878.n80 13.657
R21722 a_n1986_13878.n78 a_n1986_13878.n48 21.4216
R21723 a_n1986_13878.n61 a_n1986_13878.n20 13.657
R21724 a_n1986_13878.n37 a_n1986_13878.n63 21.4216
R21725 a_n1986_13878.n58 a_n1986_13878.n24 13.657
R21726 a_n1986_13878.n34 a_n1986_13878.n60 21.4216
R21727 a_n1986_13878.n2 a_n1986_13878.n0 1.2505
R21728 a_n1986_13878.n23 a_n1986_13878.n22 0.758076
R21729 a_n1986_13878.n22 a_n1986_13878.n21 0.758076
R21730 a_n1986_13878.n19 a_n1986_13878.n18 0.758076
R21731 a_n1986_13878.n18 a_n1986_13878.n17 0.758076
R21732 a_n1986_13878.n16 a_n1986_13878.n15 0.758076
R21733 a_n1986_13878.n13 a_n1986_13878.n12 0.758076
R21734 a_n1986_13878.n11 a_n1986_13878.n10 0.758076
R21735 a_n1986_13878.n9 a_n1986_13878.n8 0.758076
R21736 a_n1986_13878.n6 a_n1986_13878.n4 0.758076
R21737 a_n1986_13878.n6 a_n1986_13878.n5 0.758076
R21738 a_n1986_13878.n2 a_n1986_13878.n1 0.758076
R21739 a_n1986_13878.n30 a_n1986_13878.n29 0.716017
R21740 a_n1986_13878.n28 a_n1986_13878.n27 0.716017
R21741 a_n1986_13878.n26 a_n1986_13878.n25 0.716017
R21742 a_n1986_13878.n13 a_n1986_13878.n15 0.67853
R21743 a_n1986_13878.n9 a_n1986_13878.n10 0.67853
R21744 a_n1808_13878.n17 a_n1808_13878.n16 98.9632
R21745 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R21746 a_n1808_13878.n16 a_n1808_13878.n15 98.6055
R21747 a_n1808_13878.n4 a_n1808_13878.n3 98.6055
R21748 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R21749 a_n1808_13878.n14 a_n1808_13878.n13 98.6054
R21750 a_n1808_13878.n6 a_n1808_13878.t13 74.6477
R21751 a_n1808_13878.n11 a_n1808_13878.t14 74.2899
R21752 a_n1808_13878.n8 a_n1808_13878.t15 74.2899
R21753 a_n1808_13878.n7 a_n1808_13878.t12 74.2899
R21754 a_n1808_13878.n10 a_n1808_13878.n9 70.6783
R21755 a_n1808_13878.n6 a_n1808_13878.n5 70.6783
R21756 a_n1808_13878.n12 a_n1808_13878.n4 13.5694
R21757 a_n1808_13878.n14 a_n1808_13878.n12 11.5762
R21758 a_n1808_13878.n12 a_n1808_13878.n11 6.2408
R21759 a_n1808_13878.n13 a_n1808_13878.t9 3.61217
R21760 a_n1808_13878.n13 a_n1808_13878.t10 3.61217
R21761 a_n1808_13878.n15 a_n1808_13878.t0 3.61217
R21762 a_n1808_13878.n15 a_n1808_13878.t5 3.61217
R21763 a_n1808_13878.n9 a_n1808_13878.t18 3.61217
R21764 a_n1808_13878.n9 a_n1808_13878.t19 3.61217
R21765 a_n1808_13878.n5 a_n1808_13878.t16 3.61217
R21766 a_n1808_13878.n5 a_n1808_13878.t17 3.61217
R21767 a_n1808_13878.n3 a_n1808_13878.t6 3.61217
R21768 a_n1808_13878.n3 a_n1808_13878.t1 3.61217
R21769 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R21770 a_n1808_13878.n1 a_n1808_13878.t3 3.61217
R21771 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R21772 a_n1808_13878.n0 a_n1808_13878.t4 3.61217
R21773 a_n1808_13878.n17 a_n1808_13878.t7 3.61217
R21774 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R21775 a_n1808_13878.n7 a_n1808_13878.n6 0.358259
R21776 a_n1808_13878.n10 a_n1808_13878.n8 0.358259
R21777 a_n1808_13878.n11 a_n1808_13878.n10 0.358259
R21778 a_n1808_13878.n16 a_n1808_13878.n14 0.358259
R21779 a_n1808_13878.n4 a_n1808_13878.n2 0.146627
R21780 a_n1808_13878.n8 a_n1808_13878.n7 0.101793
R21781 diffpairibias.n0 diffpairibias.t27 436.822
R21782 diffpairibias.n27 diffpairibias.t24 435.479
R21783 diffpairibias.n26 diffpairibias.t21 435.479
R21784 diffpairibias.n25 diffpairibias.t22 435.479
R21785 diffpairibias.n24 diffpairibias.t26 435.479
R21786 diffpairibias.n23 diffpairibias.t20 435.479
R21787 diffpairibias.n0 diffpairibias.t23 435.479
R21788 diffpairibias.n1 diffpairibias.t28 435.479
R21789 diffpairibias.n2 diffpairibias.t25 435.479
R21790 diffpairibias.n3 diffpairibias.t29 435.479
R21791 diffpairibias.n13 diffpairibias.t14 377.536
R21792 diffpairibias.n13 diffpairibias.t0 376.193
R21793 diffpairibias.n14 diffpairibias.t10 376.193
R21794 diffpairibias.n15 diffpairibias.t12 376.193
R21795 diffpairibias.n16 diffpairibias.t6 376.193
R21796 diffpairibias.n17 diffpairibias.t2 376.193
R21797 diffpairibias.n18 diffpairibias.t16 376.193
R21798 diffpairibias.n19 diffpairibias.t4 376.193
R21799 diffpairibias.n20 diffpairibias.t18 376.193
R21800 diffpairibias.n21 diffpairibias.t8 376.193
R21801 diffpairibias.n4 diffpairibias.t15 113.368
R21802 diffpairibias.n4 diffpairibias.t1 112.698
R21803 diffpairibias.n5 diffpairibias.t11 112.698
R21804 diffpairibias.n6 diffpairibias.t13 112.698
R21805 diffpairibias.n7 diffpairibias.t7 112.698
R21806 diffpairibias.n8 diffpairibias.t3 112.698
R21807 diffpairibias.n9 diffpairibias.t17 112.698
R21808 diffpairibias.n10 diffpairibias.t5 112.698
R21809 diffpairibias.n11 diffpairibias.t19 112.698
R21810 diffpairibias.n12 diffpairibias.t9 112.698
R21811 diffpairibias.n22 diffpairibias.n21 4.77242
R21812 diffpairibias.n22 diffpairibias.n12 4.30807
R21813 diffpairibias.n23 diffpairibias.n22 4.13945
R21814 diffpairibias.n21 diffpairibias.n20 1.34352
R21815 diffpairibias.n20 diffpairibias.n19 1.34352
R21816 diffpairibias.n19 diffpairibias.n18 1.34352
R21817 diffpairibias.n18 diffpairibias.n17 1.34352
R21818 diffpairibias.n17 diffpairibias.n16 1.34352
R21819 diffpairibias.n16 diffpairibias.n15 1.34352
R21820 diffpairibias.n15 diffpairibias.n14 1.34352
R21821 diffpairibias.n14 diffpairibias.n13 1.34352
R21822 diffpairibias.n3 diffpairibias.n2 1.34352
R21823 diffpairibias.n2 diffpairibias.n1 1.34352
R21824 diffpairibias.n1 diffpairibias.n0 1.34352
R21825 diffpairibias.n24 diffpairibias.n23 1.34352
R21826 diffpairibias.n25 diffpairibias.n24 1.34352
R21827 diffpairibias.n26 diffpairibias.n25 1.34352
R21828 diffpairibias.n27 diffpairibias.n26 1.34352
R21829 diffpairibias.n28 diffpairibias.n27 0.862419
R21830 diffpairibias diffpairibias.n28 0.684875
R21831 diffpairibias.n12 diffpairibias.n11 0.672012
R21832 diffpairibias.n11 diffpairibias.n10 0.672012
R21833 diffpairibias.n10 diffpairibias.n9 0.672012
R21834 diffpairibias.n9 diffpairibias.n8 0.672012
R21835 diffpairibias.n8 diffpairibias.n7 0.672012
R21836 diffpairibias.n7 diffpairibias.n6 0.672012
R21837 diffpairibias.n6 diffpairibias.n5 0.672012
R21838 diffpairibias.n5 diffpairibias.n4 0.672012
R21839 diffpairibias.n28 diffpairibias.n3 0.190907
R21840 a_n3827_n3924.n35 a_n3827_n3924.t31 214.994
R21841 a_n3827_n3924.t38 a_n3827_n3924.n42 214.994
R21842 a_n3827_n3924.n35 a_n3827_n3924.t35 214.321
R21843 a_n3827_n3924.n0 a_n3827_n3924.t30 214.321
R21844 a_n3827_n3924.n36 a_n3827_n3924.t33 214.321
R21845 a_n3827_n3924.n37 a_n3827_n3924.t29 214.321
R21846 a_n3827_n3924.n38 a_n3827_n3924.t34 214.321
R21847 a_n3827_n3924.n39 a_n3827_n3924.t37 214.321
R21848 a_n3827_n3924.n41 a_n3827_n3924.t36 214.321
R21849 a_n3827_n3924.n42 a_n3827_n3924.t32 214.321
R21850 a_n3827_n3924.n10 a_n3827_n3924.t15 55.8337
R21851 a_n3827_n3924.n9 a_n3827_n3924.t0 55.8337
R21852 a_n3827_n3924.n2 a_n3827_n3924.t7 55.8337
R21853 a_n3827_n3924.n17 a_n3827_n3924.t9 55.8335
R21854 a_n3827_n3924.n33 a_n3827_n3924.t40 55.8335
R21855 a_n3827_n3924.n26 a_n3827_n3924.t3 55.8335
R21856 a_n3827_n3924.n25 a_n3827_n3924.t13 55.8335
R21857 a_n3827_n3924.n18 a_n3827_n3924.t16 55.8335
R21858 a_n3827_n3924.n16 a_n3827_n3924.n15 53.0052
R21859 a_n3827_n3924.n14 a_n3827_n3924.n13 53.0052
R21860 a_n3827_n3924.n12 a_n3827_n3924.n11 53.0052
R21861 a_n3827_n3924.n8 a_n3827_n3924.n7 53.0052
R21862 a_n3827_n3924.n6 a_n3827_n3924.n5 53.0052
R21863 a_n3827_n3924.n4 a_n3827_n3924.n3 53.0052
R21864 a_n3827_n3924.n32 a_n3827_n3924.n31 53.0051
R21865 a_n3827_n3924.n30 a_n3827_n3924.n29 53.0051
R21866 a_n3827_n3924.n28 a_n3827_n3924.n27 53.0051
R21867 a_n3827_n3924.n24 a_n3827_n3924.n23 53.0051
R21868 a_n3827_n3924.n22 a_n3827_n3924.n21 53.0051
R21869 a_n3827_n3924.n20 a_n3827_n3924.n19 53.0051
R21870 a_n3827_n3924.n2 a_n3827_n3924.n1 12.1555
R21871 a_n3827_n3924.n34 a_n3827_n3924.n17 12.1555
R21872 a_n3827_n3924.n18 a_n3827_n3924.n1 5.07593
R21873 a_n3827_n3924.n34 a_n3827_n3924.n33 5.07593
R21874 a_n3827_n3924.n31 a_n3827_n3924.t25 2.82907
R21875 a_n3827_n3924.n31 a_n3827_n3924.t8 2.82907
R21876 a_n3827_n3924.n29 a_n3827_n3924.t6 2.82907
R21877 a_n3827_n3924.n29 a_n3827_n3924.t14 2.82907
R21878 a_n3827_n3924.n27 a_n3827_n3924.t2 2.82907
R21879 a_n3827_n3924.n27 a_n3827_n3924.t4 2.82907
R21880 a_n3827_n3924.n23 a_n3827_n3924.t41 2.82907
R21881 a_n3827_n3924.n23 a_n3827_n3924.t24 2.82907
R21882 a_n3827_n3924.n21 a_n3827_n3924.t21 2.82907
R21883 a_n3827_n3924.n21 a_n3827_n3924.t17 2.82907
R21884 a_n3827_n3924.n19 a_n3827_n3924.t12 2.82907
R21885 a_n3827_n3924.n19 a_n3827_n3924.t10 2.82907
R21886 a_n3827_n3924.n15 a_n3827_n3924.t22 2.82907
R21887 a_n3827_n3924.n15 a_n3827_n3924.t23 2.82907
R21888 a_n3827_n3924.n13 a_n3827_n3924.t20 2.82907
R21889 a_n3827_n3924.n13 a_n3827_n3924.t28 2.82907
R21890 a_n3827_n3924.n11 a_n3827_n3924.t27 2.82907
R21891 a_n3827_n3924.n11 a_n3827_n3924.t18 2.82907
R21892 a_n3827_n3924.n7 a_n3827_n3924.t11 2.82907
R21893 a_n3827_n3924.n7 a_n3827_n3924.t5 2.82907
R21894 a_n3827_n3924.n5 a_n3827_n3924.t26 2.82907
R21895 a_n3827_n3924.n5 a_n3827_n3924.t19 2.82907
R21896 a_n3827_n3924.n3 a_n3827_n3924.t1 2.82907
R21897 a_n3827_n3924.n3 a_n3827_n3924.t39 2.82907
R21898 a_n3827_n3924.n40 a_n3827_n3924.n1 1.95694
R21899 a_n3827_n3924.n0 a_n3827_n3924.n34 1.95694
R21900 a_n3827_n3924.n42 a_n3827_n3924.n41 0.672012
R21901 a_n3827_n3924.n39 a_n3827_n3924.n38 0.672012
R21902 a_n3827_n3924.n38 a_n3827_n3924.n37 0.672012
R21903 a_n3827_n3924.n37 a_n3827_n3924.n36 0.672012
R21904 a_n3827_n3924.n36 a_n3827_n3924.n0 0.672012
R21905 a_n3827_n3924.n0 a_n3827_n3924.n35 0.672012
R21906 a_n3827_n3924.n41 a_n3827_n3924.n40 0.511401
R21907 a_n3827_n3924.n4 a_n3827_n3924.n2 0.358259
R21908 a_n3827_n3924.n6 a_n3827_n3924.n4 0.358259
R21909 a_n3827_n3924.n8 a_n3827_n3924.n6 0.358259
R21910 a_n3827_n3924.n9 a_n3827_n3924.n8 0.358259
R21911 a_n3827_n3924.n12 a_n3827_n3924.n10 0.358259
R21912 a_n3827_n3924.n14 a_n3827_n3924.n12 0.358259
R21913 a_n3827_n3924.n16 a_n3827_n3924.n14 0.358259
R21914 a_n3827_n3924.n17 a_n3827_n3924.n16 0.358259
R21915 a_n3827_n3924.n20 a_n3827_n3924.n18 0.358259
R21916 a_n3827_n3924.n22 a_n3827_n3924.n20 0.358259
R21917 a_n3827_n3924.n24 a_n3827_n3924.n22 0.358259
R21918 a_n3827_n3924.n25 a_n3827_n3924.n24 0.358259
R21919 a_n3827_n3924.n28 a_n3827_n3924.n26 0.358259
R21920 a_n3827_n3924.n30 a_n3827_n3924.n28 0.358259
R21921 a_n3827_n3924.n32 a_n3827_n3924.n30 0.358259
R21922 a_n3827_n3924.n33 a_n3827_n3924.n32 0.358259
R21923 a_n3827_n3924.n10 a_n3827_n3924.n9 0.235414
R21924 a_n3827_n3924.n26 a_n3827_n3924.n25 0.235414
R21925 a_n3827_n3924.n40 a_n3827_n3924.n39 0.16111
R21926 a_n1986_8322.n6 a_n1986_8322.t17 74.6477
R21927 a_n1986_8322.n1 a_n1986_8322.t3 74.6477
R21928 a_n1986_8322.n16 a_n1986_8322.t12 74.6474
R21929 a_n1986_8322.n14 a_n1986_8322.t5 74.2899
R21930 a_n1986_8322.n7 a_n1986_8322.t15 74.2899
R21931 a_n1986_8322.n8 a_n1986_8322.t18 74.2899
R21932 a_n1986_8322.n11 a_n1986_8322.t19 74.2899
R21933 a_n1986_8322.n4 a_n1986_8322.t2 74.2899
R21934 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R21935 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R21936 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R21937 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R21938 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R21939 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R21940 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R21941 a_n1986_8322.n13 a_n1986_8322.t0 9.94227
R21942 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R21943 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R21944 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R21945 a_n1986_8322.n15 a_n1986_8322.t10 3.61217
R21946 a_n1986_8322.n15 a_n1986_8322.t7 3.61217
R21947 a_n1986_8322.n5 a_n1986_8322.t21 3.61217
R21948 a_n1986_8322.n5 a_n1986_8322.t20 3.61217
R21949 a_n1986_8322.n9 a_n1986_8322.t16 3.61217
R21950 a_n1986_8322.n9 a_n1986_8322.t14 3.61217
R21951 a_n1986_8322.n0 a_n1986_8322.t11 3.61217
R21952 a_n1986_8322.n0 a_n1986_8322.t6 3.61217
R21953 a_n1986_8322.n2 a_n1986_8322.t9 3.61217
R21954 a_n1986_8322.n2 a_n1986_8322.t8 3.61217
R21955 a_n1986_8322.n18 a_n1986_8322.t4 3.61217
R21956 a_n1986_8322.t13 a_n1986_8322.n18 3.61217
R21957 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R21958 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R21959 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R21960 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R21961 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R21962 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R21963 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R21964 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R21965 a_n1986_8322.t0 a_n1986_8322.t1 0.057021
R21966 plus.n27 plus.t19 436.949
R21967 plus.n5 plus.t11 436.949
R21968 plus.n28 plus.t5 415.966
R21969 plus.n30 plus.t17 415.966
R21970 plus.n34 plus.t20 415.966
R21971 plus.n35 plus.t10 415.966
R21972 plus.n23 plus.t6 415.966
R21973 plus.n41 plus.t9 415.966
R21974 plus.n42 plus.t16 415.966
R21975 plus.n20 plus.t7 415.966
R21976 plus.n19 plus.t15 415.966
R21977 plus.n1 plus.t12 415.966
R21978 plus.n13 plus.t18 415.966
R21979 plus.n12 plus.t14 415.966
R21980 plus.n4 plus.t8 415.966
R21981 plus.n6 plus.t13 415.966
R21982 plus.n46 plus.t4 243.97
R21983 plus.n46 plus.n45 223.454
R21984 plus.n48 plus.n47 223.454
R21985 plus.n43 plus.n42 161.3
R21986 plus.n41 plus.n22 161.3
R21987 plus.n40 plus.n39 161.3
R21988 plus.n38 plus.n23 161.3
R21989 plus.n37 plus.n36 161.3
R21990 plus.n35 plus.n24 161.3
R21991 plus.n34 plus.n33 161.3
R21992 plus.n32 plus.n25 161.3
R21993 plus.n31 plus.n30 161.3
R21994 plus.n29 plus.n26 161.3
R21995 plus.n8 plus.n7 161.3
R21996 plus.n9 plus.n4 161.3
R21997 plus.n11 plus.n10 161.3
R21998 plus.n12 plus.n3 161.3
R21999 plus.n13 plus.n2 161.3
R22000 plus.n15 plus.n14 161.3
R22001 plus.n16 plus.n1 161.3
R22002 plus.n18 plus.n17 161.3
R22003 plus.n19 plus.n0 161.3
R22004 plus.n21 plus.n20 161.3
R22005 plus.n27 plus.n26 70.4033
R22006 plus.n8 plus.n5 70.4033
R22007 plus.n35 plus.n34 48.2005
R22008 plus.n42 plus.n41 48.2005
R22009 plus.n20 plus.n19 48.2005
R22010 plus.n13 plus.n12 48.2005
R22011 plus.n30 plus.n29 37.246
R22012 plus.n40 plus.n23 37.246
R22013 plus.n18 plus.n1 37.246
R22014 plus.n7 plus.n4 37.246
R22015 plus.n30 plus.n25 35.7853
R22016 plus.n36 plus.n23 35.7853
R22017 plus.n14 plus.n1 35.7853
R22018 plus.n11 plus.n4 35.7853
R22019 plus.n44 plus.n43 28.5744
R22020 plus.n28 plus.n27 20.9576
R22021 plus.n6 plus.n5 20.9576
R22022 plus.n45 plus.t0 19.8005
R22023 plus.n45 plus.t1 19.8005
R22024 plus.n47 plus.t3 19.8005
R22025 plus.n47 plus.t2 19.8005
R22026 plus plus.n49 14.1603
R22027 plus.n34 plus.n25 12.4157
R22028 plus.n36 plus.n35 12.4157
R22029 plus.n14 plus.n13 12.4157
R22030 plus.n12 plus.n11 12.4157
R22031 plus.n44 plus.n21 11.76
R22032 plus.n29 plus.n28 10.955
R22033 plus.n41 plus.n40 10.955
R22034 plus.n19 plus.n18 10.955
R22035 plus.n7 plus.n6 10.955
R22036 plus.n49 plus.n48 5.40567
R22037 plus.n49 plus.n44 1.188
R22038 plus.n48 plus.n46 0.716017
R22039 plus.n31 plus.n26 0.189894
R22040 plus.n32 plus.n31 0.189894
R22041 plus.n33 plus.n32 0.189894
R22042 plus.n33 plus.n24 0.189894
R22043 plus.n37 plus.n24 0.189894
R22044 plus.n38 plus.n37 0.189894
R22045 plus.n39 plus.n38 0.189894
R22046 plus.n39 plus.n22 0.189894
R22047 plus.n43 plus.n22 0.189894
R22048 plus.n21 plus.n0 0.189894
R22049 plus.n17 plus.n0 0.189894
R22050 plus.n17 plus.n16 0.189894
R22051 plus.n16 plus.n15 0.189894
R22052 plus.n15 plus.n2 0.189894
R22053 plus.n3 plus.n2 0.189894
R22054 plus.n10 plus.n3 0.189894
R22055 plus.n10 plus.n9 0.189894
R22056 plus.n9 plus.n8 0.189894
R22057 outputibias.n27 outputibias.n1 289.615
R22058 outputibias.n58 outputibias.n32 289.615
R22059 outputibias.n90 outputibias.n64 289.615
R22060 outputibias.n122 outputibias.n96 289.615
R22061 outputibias.n28 outputibias.n27 185
R22062 outputibias.n26 outputibias.n25 185
R22063 outputibias.n5 outputibias.n4 185
R22064 outputibias.n20 outputibias.n19 185
R22065 outputibias.n18 outputibias.n17 185
R22066 outputibias.n9 outputibias.n8 185
R22067 outputibias.n12 outputibias.n11 185
R22068 outputibias.n59 outputibias.n58 185
R22069 outputibias.n57 outputibias.n56 185
R22070 outputibias.n36 outputibias.n35 185
R22071 outputibias.n51 outputibias.n50 185
R22072 outputibias.n49 outputibias.n48 185
R22073 outputibias.n40 outputibias.n39 185
R22074 outputibias.n43 outputibias.n42 185
R22075 outputibias.n91 outputibias.n90 185
R22076 outputibias.n89 outputibias.n88 185
R22077 outputibias.n68 outputibias.n67 185
R22078 outputibias.n83 outputibias.n82 185
R22079 outputibias.n81 outputibias.n80 185
R22080 outputibias.n72 outputibias.n71 185
R22081 outputibias.n75 outputibias.n74 185
R22082 outputibias.n123 outputibias.n122 185
R22083 outputibias.n121 outputibias.n120 185
R22084 outputibias.n100 outputibias.n99 185
R22085 outputibias.n115 outputibias.n114 185
R22086 outputibias.n113 outputibias.n112 185
R22087 outputibias.n104 outputibias.n103 185
R22088 outputibias.n107 outputibias.n106 185
R22089 outputibias.n0 outputibias.t10 178.945
R22090 outputibias.n133 outputibias.t8 177.018
R22091 outputibias.n132 outputibias.t11 177.018
R22092 outputibias.n0 outputibias.t9 177.018
R22093 outputibias.t7 outputibias.n10 147.661
R22094 outputibias.t1 outputibias.n41 147.661
R22095 outputibias.t3 outputibias.n73 147.661
R22096 outputibias.t5 outputibias.n105 147.661
R22097 outputibias.n128 outputibias.t6 132.363
R22098 outputibias.n128 outputibias.t0 130.436
R22099 outputibias.n129 outputibias.t2 130.436
R22100 outputibias.n130 outputibias.t4 130.436
R22101 outputibias.n27 outputibias.n26 104.615
R22102 outputibias.n26 outputibias.n4 104.615
R22103 outputibias.n19 outputibias.n4 104.615
R22104 outputibias.n19 outputibias.n18 104.615
R22105 outputibias.n18 outputibias.n8 104.615
R22106 outputibias.n11 outputibias.n8 104.615
R22107 outputibias.n58 outputibias.n57 104.615
R22108 outputibias.n57 outputibias.n35 104.615
R22109 outputibias.n50 outputibias.n35 104.615
R22110 outputibias.n50 outputibias.n49 104.615
R22111 outputibias.n49 outputibias.n39 104.615
R22112 outputibias.n42 outputibias.n39 104.615
R22113 outputibias.n90 outputibias.n89 104.615
R22114 outputibias.n89 outputibias.n67 104.615
R22115 outputibias.n82 outputibias.n67 104.615
R22116 outputibias.n82 outputibias.n81 104.615
R22117 outputibias.n81 outputibias.n71 104.615
R22118 outputibias.n74 outputibias.n71 104.615
R22119 outputibias.n122 outputibias.n121 104.615
R22120 outputibias.n121 outputibias.n99 104.615
R22121 outputibias.n114 outputibias.n99 104.615
R22122 outputibias.n114 outputibias.n113 104.615
R22123 outputibias.n113 outputibias.n103 104.615
R22124 outputibias.n106 outputibias.n103 104.615
R22125 outputibias.n63 outputibias.n31 95.6354
R22126 outputibias.n63 outputibias.n62 94.6732
R22127 outputibias.n95 outputibias.n94 94.6732
R22128 outputibias.n127 outputibias.n126 94.6732
R22129 outputibias.n11 outputibias.t7 52.3082
R22130 outputibias.n42 outputibias.t1 52.3082
R22131 outputibias.n74 outputibias.t3 52.3082
R22132 outputibias.n106 outputibias.t5 52.3082
R22133 outputibias.n12 outputibias.n10 15.6674
R22134 outputibias.n43 outputibias.n41 15.6674
R22135 outputibias.n75 outputibias.n73 15.6674
R22136 outputibias.n107 outputibias.n105 15.6674
R22137 outputibias.n13 outputibias.n9 12.8005
R22138 outputibias.n44 outputibias.n40 12.8005
R22139 outputibias.n76 outputibias.n72 12.8005
R22140 outputibias.n108 outputibias.n104 12.8005
R22141 outputibias.n17 outputibias.n16 12.0247
R22142 outputibias.n48 outputibias.n47 12.0247
R22143 outputibias.n80 outputibias.n79 12.0247
R22144 outputibias.n112 outputibias.n111 12.0247
R22145 outputibias.n20 outputibias.n7 11.249
R22146 outputibias.n51 outputibias.n38 11.249
R22147 outputibias.n83 outputibias.n70 11.249
R22148 outputibias.n115 outputibias.n102 11.249
R22149 outputibias.n21 outputibias.n5 10.4732
R22150 outputibias.n52 outputibias.n36 10.4732
R22151 outputibias.n84 outputibias.n68 10.4732
R22152 outputibias.n116 outputibias.n100 10.4732
R22153 outputibias.n25 outputibias.n24 9.69747
R22154 outputibias.n56 outputibias.n55 9.69747
R22155 outputibias.n88 outputibias.n87 9.69747
R22156 outputibias.n120 outputibias.n119 9.69747
R22157 outputibias.n31 outputibias.n30 9.45567
R22158 outputibias.n62 outputibias.n61 9.45567
R22159 outputibias.n94 outputibias.n93 9.45567
R22160 outputibias.n126 outputibias.n125 9.45567
R22161 outputibias.n30 outputibias.n29 9.3005
R22162 outputibias.n3 outputibias.n2 9.3005
R22163 outputibias.n24 outputibias.n23 9.3005
R22164 outputibias.n22 outputibias.n21 9.3005
R22165 outputibias.n7 outputibias.n6 9.3005
R22166 outputibias.n16 outputibias.n15 9.3005
R22167 outputibias.n14 outputibias.n13 9.3005
R22168 outputibias.n61 outputibias.n60 9.3005
R22169 outputibias.n34 outputibias.n33 9.3005
R22170 outputibias.n55 outputibias.n54 9.3005
R22171 outputibias.n53 outputibias.n52 9.3005
R22172 outputibias.n38 outputibias.n37 9.3005
R22173 outputibias.n47 outputibias.n46 9.3005
R22174 outputibias.n45 outputibias.n44 9.3005
R22175 outputibias.n93 outputibias.n92 9.3005
R22176 outputibias.n66 outputibias.n65 9.3005
R22177 outputibias.n87 outputibias.n86 9.3005
R22178 outputibias.n85 outputibias.n84 9.3005
R22179 outputibias.n70 outputibias.n69 9.3005
R22180 outputibias.n79 outputibias.n78 9.3005
R22181 outputibias.n77 outputibias.n76 9.3005
R22182 outputibias.n125 outputibias.n124 9.3005
R22183 outputibias.n98 outputibias.n97 9.3005
R22184 outputibias.n119 outputibias.n118 9.3005
R22185 outputibias.n117 outputibias.n116 9.3005
R22186 outputibias.n102 outputibias.n101 9.3005
R22187 outputibias.n111 outputibias.n110 9.3005
R22188 outputibias.n109 outputibias.n108 9.3005
R22189 outputibias.n28 outputibias.n3 8.92171
R22190 outputibias.n59 outputibias.n34 8.92171
R22191 outputibias.n91 outputibias.n66 8.92171
R22192 outputibias.n123 outputibias.n98 8.92171
R22193 outputibias.n29 outputibias.n1 8.14595
R22194 outputibias.n60 outputibias.n32 8.14595
R22195 outputibias.n92 outputibias.n64 8.14595
R22196 outputibias.n124 outputibias.n96 8.14595
R22197 outputibias.n31 outputibias.n1 5.81868
R22198 outputibias.n62 outputibias.n32 5.81868
R22199 outputibias.n94 outputibias.n64 5.81868
R22200 outputibias.n126 outputibias.n96 5.81868
R22201 outputibias.n131 outputibias.n130 5.20947
R22202 outputibias.n29 outputibias.n28 5.04292
R22203 outputibias.n60 outputibias.n59 5.04292
R22204 outputibias.n92 outputibias.n91 5.04292
R22205 outputibias.n124 outputibias.n123 5.04292
R22206 outputibias.n131 outputibias.n127 4.42209
R22207 outputibias.n14 outputibias.n10 4.38594
R22208 outputibias.n45 outputibias.n41 4.38594
R22209 outputibias.n77 outputibias.n73 4.38594
R22210 outputibias.n109 outputibias.n105 4.38594
R22211 outputibias.n132 outputibias.n131 4.28454
R22212 outputibias.n25 outputibias.n3 4.26717
R22213 outputibias.n56 outputibias.n34 4.26717
R22214 outputibias.n88 outputibias.n66 4.26717
R22215 outputibias.n120 outputibias.n98 4.26717
R22216 outputibias.n24 outputibias.n5 3.49141
R22217 outputibias.n55 outputibias.n36 3.49141
R22218 outputibias.n87 outputibias.n68 3.49141
R22219 outputibias.n119 outputibias.n100 3.49141
R22220 outputibias.n21 outputibias.n20 2.71565
R22221 outputibias.n52 outputibias.n51 2.71565
R22222 outputibias.n84 outputibias.n83 2.71565
R22223 outputibias.n116 outputibias.n115 2.71565
R22224 outputibias.n17 outputibias.n7 1.93989
R22225 outputibias.n48 outputibias.n38 1.93989
R22226 outputibias.n80 outputibias.n70 1.93989
R22227 outputibias.n112 outputibias.n102 1.93989
R22228 outputibias.n130 outputibias.n129 1.9266
R22229 outputibias.n129 outputibias.n128 1.9266
R22230 outputibias.n133 outputibias.n132 1.92658
R22231 outputibias.n134 outputibias.n133 1.29913
R22232 outputibias.n16 outputibias.n9 1.16414
R22233 outputibias.n47 outputibias.n40 1.16414
R22234 outputibias.n79 outputibias.n72 1.16414
R22235 outputibias.n111 outputibias.n104 1.16414
R22236 outputibias.n127 outputibias.n95 0.962709
R22237 outputibias.n95 outputibias.n63 0.962709
R22238 outputibias.n13 outputibias.n12 0.388379
R22239 outputibias.n44 outputibias.n43 0.388379
R22240 outputibias.n76 outputibias.n75 0.388379
R22241 outputibias.n108 outputibias.n107 0.388379
R22242 outputibias.n134 outputibias.n0 0.337251
R22243 outputibias outputibias.n134 0.302375
R22244 outputibias.n30 outputibias.n2 0.155672
R22245 outputibias.n23 outputibias.n2 0.155672
R22246 outputibias.n23 outputibias.n22 0.155672
R22247 outputibias.n22 outputibias.n6 0.155672
R22248 outputibias.n15 outputibias.n6 0.155672
R22249 outputibias.n15 outputibias.n14 0.155672
R22250 outputibias.n61 outputibias.n33 0.155672
R22251 outputibias.n54 outputibias.n33 0.155672
R22252 outputibias.n54 outputibias.n53 0.155672
R22253 outputibias.n53 outputibias.n37 0.155672
R22254 outputibias.n46 outputibias.n37 0.155672
R22255 outputibias.n46 outputibias.n45 0.155672
R22256 outputibias.n93 outputibias.n65 0.155672
R22257 outputibias.n86 outputibias.n65 0.155672
R22258 outputibias.n86 outputibias.n85 0.155672
R22259 outputibias.n85 outputibias.n69 0.155672
R22260 outputibias.n78 outputibias.n69 0.155672
R22261 outputibias.n78 outputibias.n77 0.155672
R22262 outputibias.n125 outputibias.n97 0.155672
R22263 outputibias.n118 outputibias.n97 0.155672
R22264 outputibias.n118 outputibias.n117 0.155672
R22265 outputibias.n117 outputibias.n101 0.155672
R22266 outputibias.n110 outputibias.n101 0.155672
R22267 outputibias.n110 outputibias.n109 0.155672
R22268 output.n41 output.n15 289.615
R22269 output.n72 output.n46 289.615
R22270 output.n104 output.n78 289.615
R22271 output.n136 output.n110 289.615
R22272 output.n77 output.n45 197.26
R22273 output.n77 output.n76 196.298
R22274 output.n109 output.n108 196.298
R22275 output.n141 output.n140 196.298
R22276 output.n42 output.n41 185
R22277 output.n40 output.n39 185
R22278 output.n19 output.n18 185
R22279 output.n34 output.n33 185
R22280 output.n32 output.n31 185
R22281 output.n23 output.n22 185
R22282 output.n26 output.n25 185
R22283 output.n73 output.n72 185
R22284 output.n71 output.n70 185
R22285 output.n50 output.n49 185
R22286 output.n65 output.n64 185
R22287 output.n63 output.n62 185
R22288 output.n54 output.n53 185
R22289 output.n57 output.n56 185
R22290 output.n105 output.n104 185
R22291 output.n103 output.n102 185
R22292 output.n82 output.n81 185
R22293 output.n97 output.n96 185
R22294 output.n95 output.n94 185
R22295 output.n86 output.n85 185
R22296 output.n89 output.n88 185
R22297 output.n137 output.n136 185
R22298 output.n135 output.n134 185
R22299 output.n114 output.n113 185
R22300 output.n129 output.n128 185
R22301 output.n127 output.n126 185
R22302 output.n118 output.n117 185
R22303 output.n121 output.n120 185
R22304 output.t1 output.n24 147.661
R22305 output.t2 output.n55 147.661
R22306 output.t3 output.n87 147.661
R22307 output.t0 output.n119 147.661
R22308 output.n41 output.n40 104.615
R22309 output.n40 output.n18 104.615
R22310 output.n33 output.n18 104.615
R22311 output.n33 output.n32 104.615
R22312 output.n32 output.n22 104.615
R22313 output.n25 output.n22 104.615
R22314 output.n72 output.n71 104.615
R22315 output.n71 output.n49 104.615
R22316 output.n64 output.n49 104.615
R22317 output.n64 output.n63 104.615
R22318 output.n63 output.n53 104.615
R22319 output.n56 output.n53 104.615
R22320 output.n104 output.n103 104.615
R22321 output.n103 output.n81 104.615
R22322 output.n96 output.n81 104.615
R22323 output.n96 output.n95 104.615
R22324 output.n95 output.n85 104.615
R22325 output.n88 output.n85 104.615
R22326 output.n136 output.n135 104.615
R22327 output.n135 output.n113 104.615
R22328 output.n128 output.n113 104.615
R22329 output.n128 output.n127 104.615
R22330 output.n127 output.n117 104.615
R22331 output.n120 output.n117 104.615
R22332 output.n1 output.t5 77.056
R22333 output.n14 output.t7 76.6694
R22334 output.n1 output.n0 72.7095
R22335 output.n3 output.n2 72.7095
R22336 output.n5 output.n4 72.7095
R22337 output.n7 output.n6 72.7095
R22338 output.n9 output.n8 72.7095
R22339 output.n11 output.n10 72.7095
R22340 output.n13 output.n12 72.7095
R22341 output.n25 output.t1 52.3082
R22342 output.n56 output.t2 52.3082
R22343 output.n88 output.t3 52.3082
R22344 output.n120 output.t0 52.3082
R22345 output.n26 output.n24 15.6674
R22346 output.n57 output.n55 15.6674
R22347 output.n89 output.n87 15.6674
R22348 output.n121 output.n119 15.6674
R22349 output.n27 output.n23 12.8005
R22350 output.n58 output.n54 12.8005
R22351 output.n90 output.n86 12.8005
R22352 output.n122 output.n118 12.8005
R22353 output.n31 output.n30 12.0247
R22354 output.n62 output.n61 12.0247
R22355 output.n94 output.n93 12.0247
R22356 output.n126 output.n125 12.0247
R22357 output.n34 output.n21 11.249
R22358 output.n65 output.n52 11.249
R22359 output.n97 output.n84 11.249
R22360 output.n129 output.n116 11.249
R22361 output.n35 output.n19 10.4732
R22362 output.n66 output.n50 10.4732
R22363 output.n98 output.n82 10.4732
R22364 output.n130 output.n114 10.4732
R22365 output.n39 output.n38 9.69747
R22366 output.n70 output.n69 9.69747
R22367 output.n102 output.n101 9.69747
R22368 output.n134 output.n133 9.69747
R22369 output.n45 output.n44 9.45567
R22370 output.n76 output.n75 9.45567
R22371 output.n108 output.n107 9.45567
R22372 output.n140 output.n139 9.45567
R22373 output.n44 output.n43 9.3005
R22374 output.n17 output.n16 9.3005
R22375 output.n38 output.n37 9.3005
R22376 output.n36 output.n35 9.3005
R22377 output.n21 output.n20 9.3005
R22378 output.n30 output.n29 9.3005
R22379 output.n28 output.n27 9.3005
R22380 output.n75 output.n74 9.3005
R22381 output.n48 output.n47 9.3005
R22382 output.n69 output.n68 9.3005
R22383 output.n67 output.n66 9.3005
R22384 output.n52 output.n51 9.3005
R22385 output.n61 output.n60 9.3005
R22386 output.n59 output.n58 9.3005
R22387 output.n107 output.n106 9.3005
R22388 output.n80 output.n79 9.3005
R22389 output.n101 output.n100 9.3005
R22390 output.n99 output.n98 9.3005
R22391 output.n84 output.n83 9.3005
R22392 output.n93 output.n92 9.3005
R22393 output.n91 output.n90 9.3005
R22394 output.n139 output.n138 9.3005
R22395 output.n112 output.n111 9.3005
R22396 output.n133 output.n132 9.3005
R22397 output.n131 output.n130 9.3005
R22398 output.n116 output.n115 9.3005
R22399 output.n125 output.n124 9.3005
R22400 output.n123 output.n122 9.3005
R22401 output.n42 output.n17 8.92171
R22402 output.n73 output.n48 8.92171
R22403 output.n105 output.n80 8.92171
R22404 output.n137 output.n112 8.92171
R22405 output output.n141 8.15037
R22406 output.n43 output.n15 8.14595
R22407 output.n74 output.n46 8.14595
R22408 output.n106 output.n78 8.14595
R22409 output.n138 output.n110 8.14595
R22410 output.n45 output.n15 5.81868
R22411 output.n76 output.n46 5.81868
R22412 output.n108 output.n78 5.81868
R22413 output.n140 output.n110 5.81868
R22414 output.n43 output.n42 5.04292
R22415 output.n74 output.n73 5.04292
R22416 output.n106 output.n105 5.04292
R22417 output.n138 output.n137 5.04292
R22418 output.n28 output.n24 4.38594
R22419 output.n59 output.n55 4.38594
R22420 output.n91 output.n87 4.38594
R22421 output.n123 output.n119 4.38594
R22422 output.n39 output.n17 4.26717
R22423 output.n70 output.n48 4.26717
R22424 output.n102 output.n80 4.26717
R22425 output.n134 output.n112 4.26717
R22426 output.n0 output.t16 3.9605
R22427 output.n0 output.t19 3.9605
R22428 output.n2 output.t9 3.9605
R22429 output.n2 output.t8 3.9605
R22430 output.n4 output.t14 3.9605
R22431 output.n4 output.t18 3.9605
R22432 output.n6 output.t6 3.9605
R22433 output.n6 output.t10 3.9605
R22434 output.n8 output.t11 3.9605
R22435 output.n8 output.t17 3.9605
R22436 output.n10 output.t4 3.9605
R22437 output.n10 output.t12 3.9605
R22438 output.n12 output.t15 3.9605
R22439 output.n12 output.t13 3.9605
R22440 output.n38 output.n19 3.49141
R22441 output.n69 output.n50 3.49141
R22442 output.n101 output.n82 3.49141
R22443 output.n133 output.n114 3.49141
R22444 output.n35 output.n34 2.71565
R22445 output.n66 output.n65 2.71565
R22446 output.n98 output.n97 2.71565
R22447 output.n130 output.n129 2.71565
R22448 output.n31 output.n21 1.93989
R22449 output.n62 output.n52 1.93989
R22450 output.n94 output.n84 1.93989
R22451 output.n126 output.n116 1.93989
R22452 output.n30 output.n23 1.16414
R22453 output.n61 output.n54 1.16414
R22454 output.n93 output.n86 1.16414
R22455 output.n125 output.n118 1.16414
R22456 output.n141 output.n109 0.962709
R22457 output.n109 output.n77 0.962709
R22458 output.n27 output.n26 0.388379
R22459 output.n58 output.n57 0.388379
R22460 output.n90 output.n89 0.388379
R22461 output.n122 output.n121 0.388379
R22462 output.n14 output.n13 0.387128
R22463 output.n13 output.n11 0.387128
R22464 output.n11 output.n9 0.387128
R22465 output.n9 output.n7 0.387128
R22466 output.n7 output.n5 0.387128
R22467 output.n5 output.n3 0.387128
R22468 output.n3 output.n1 0.387128
R22469 output.n44 output.n16 0.155672
R22470 output.n37 output.n16 0.155672
R22471 output.n37 output.n36 0.155672
R22472 output.n36 output.n20 0.155672
R22473 output.n29 output.n20 0.155672
R22474 output.n29 output.n28 0.155672
R22475 output.n75 output.n47 0.155672
R22476 output.n68 output.n47 0.155672
R22477 output.n68 output.n67 0.155672
R22478 output.n67 output.n51 0.155672
R22479 output.n60 output.n51 0.155672
R22480 output.n60 output.n59 0.155672
R22481 output.n107 output.n79 0.155672
R22482 output.n100 output.n79 0.155672
R22483 output.n100 output.n99 0.155672
R22484 output.n99 output.n83 0.155672
R22485 output.n92 output.n83 0.155672
R22486 output.n92 output.n91 0.155672
R22487 output.n139 output.n111 0.155672
R22488 output.n132 output.n111 0.155672
R22489 output.n132 output.n131 0.155672
R22490 output.n131 output.n115 0.155672
R22491 output.n124 output.n115 0.155672
R22492 output.n124 output.n123 0.155672
R22493 output output.n14 0.126227
R22494 minus.n27 minus.t20 436.949
R22495 minus.n5 minus.t11 436.949
R22496 minus.n42 minus.t17 415.966
R22497 minus.n41 minus.t10 415.966
R22498 minus.n23 minus.t5 415.966
R22499 minus.n35 minus.t13 415.966
R22500 minus.n34 minus.t9 415.966
R22501 minus.n26 minus.t19 415.966
R22502 minus.n28 minus.t7 415.966
R22503 minus.n6 minus.t14 415.966
R22504 minus.n8 minus.t8 415.966
R22505 minus.n12 minus.t12 415.966
R22506 minus.n13 minus.t18 415.966
R22507 minus.n1 minus.t15 415.966
R22508 minus.n19 minus.t16 415.966
R22509 minus.n20 minus.t6 415.966
R22510 minus.n48 minus.t1 243.255
R22511 minus.n47 minus.n45 224.169
R22512 minus.n47 minus.n46 223.454
R22513 minus.n30 minus.n29 161.3
R22514 minus.n31 minus.n26 161.3
R22515 minus.n33 minus.n32 161.3
R22516 minus.n34 minus.n25 161.3
R22517 minus.n35 minus.n24 161.3
R22518 minus.n37 minus.n36 161.3
R22519 minus.n38 minus.n23 161.3
R22520 minus.n40 minus.n39 161.3
R22521 minus.n41 minus.n22 161.3
R22522 minus.n43 minus.n42 161.3
R22523 minus.n21 minus.n20 161.3
R22524 minus.n19 minus.n0 161.3
R22525 minus.n18 minus.n17 161.3
R22526 minus.n16 minus.n1 161.3
R22527 minus.n15 minus.n14 161.3
R22528 minus.n13 minus.n2 161.3
R22529 minus.n12 minus.n11 161.3
R22530 minus.n10 minus.n3 161.3
R22531 minus.n9 minus.n8 161.3
R22532 minus.n7 minus.n4 161.3
R22533 minus.n30 minus.n27 70.4033
R22534 minus.n5 minus.n4 70.4033
R22535 minus.n42 minus.n41 48.2005
R22536 minus.n35 minus.n34 48.2005
R22537 minus.n13 minus.n12 48.2005
R22538 minus.n20 minus.n19 48.2005
R22539 minus.n40 minus.n23 37.246
R22540 minus.n29 minus.n26 37.246
R22541 minus.n8 minus.n7 37.246
R22542 minus.n18 minus.n1 37.246
R22543 minus.n36 minus.n23 35.7853
R22544 minus.n33 minus.n26 35.7853
R22545 minus.n8 minus.n3 35.7853
R22546 minus.n14 minus.n1 35.7853
R22547 minus.n44 minus.n43 28.7903
R22548 minus.n28 minus.n27 20.9576
R22549 minus.n6 minus.n5 20.9576
R22550 minus.n46 minus.t3 19.8005
R22551 minus.n46 minus.t4 19.8005
R22552 minus.n45 minus.t2 19.8005
R22553 minus.n45 minus.t0 19.8005
R22554 minus.n36 minus.n35 12.4157
R22555 minus.n34 minus.n33 12.4157
R22556 minus.n12 minus.n3 12.4157
R22557 minus.n14 minus.n13 12.4157
R22558 minus.n44 minus.n21 11.9759
R22559 minus minus.n49 11.7381
R22560 minus.n41 minus.n40 10.955
R22561 minus.n29 minus.n28 10.955
R22562 minus.n7 minus.n6 10.955
R22563 minus.n19 minus.n18 10.955
R22564 minus.n49 minus.n48 4.80222
R22565 minus.n49 minus.n44 0.972091
R22566 minus.n48 minus.n47 0.716017
R22567 minus.n43 minus.n22 0.189894
R22568 minus.n39 minus.n22 0.189894
R22569 minus.n39 minus.n38 0.189894
R22570 minus.n38 minus.n37 0.189894
R22571 minus.n37 minus.n24 0.189894
R22572 minus.n25 minus.n24 0.189894
R22573 minus.n32 minus.n25 0.189894
R22574 minus.n32 minus.n31 0.189894
R22575 minus.n31 minus.n30 0.189894
R22576 minus.n9 minus.n4 0.189894
R22577 minus.n10 minus.n9 0.189894
R22578 minus.n11 minus.n10 0.189894
R22579 minus.n11 minus.n2 0.189894
R22580 minus.n15 minus.n2 0.189894
R22581 minus.n16 minus.n15 0.189894
R22582 minus.n17 minus.n16 0.189894
R22583 minus.n17 minus.n0 0.189894
R22584 minus.n21 minus.n0 0.189894
C0 plus commonsourceibias 0.268404f
C1 output outputibias 2.34152f
C2 vdd output 7.23429f
C3 CSoutput output 6.13881f
C4 CSoutput outputibias 0.032386f
C5 vdd CSoutput 0.140616p
C6 commonsourceibias output 0.006808f
C7 minus diffpairibias 1.62e-19
C8 CSoutput minus 2.92106f
C9 vdd plus 0.0849f
C10 plus diffpairibias 2.39e-19
C11 commonsourceibias outputibias 0.003832f
C12 vdd commonsourceibias 0.004218f
C13 CSoutput plus 0.826585f
C14 commonsourceibias diffpairibias 0.064336f
C15 CSoutput commonsourceibias 42.3358f
C16 minus plus 8.493211f
C17 minus commonsourceibias 0.323331f
C18 diffpairibias gnd 60.002533f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.145046p
C22 plus gnd 28.75359f
C23 minus gnd 25.09441f
C24 CSoutput gnd 0.107728p
C25 vdd gnd 0.438684p
C26 minus.n0 gnd 0.031169f
C27 minus.t15 gnd 0.314894f
C28 minus.n1 gnd 0.145585f
C29 minus.n2 gnd 0.031169f
C30 minus.n3 gnd 0.007073f
C31 minus.n4 gnd 0.099236f
C32 minus.t11 gnd 0.32173f
C33 minus.n5 gnd 0.13571f
C34 minus.t14 gnd 0.314894f
C35 minus.n6 gnd 0.14376f
C36 minus.n7 gnd 0.007073f
C37 minus.t8 gnd 0.314894f
C38 minus.n8 gnd 0.145585f
C39 minus.n9 gnd 0.031169f
C40 minus.n10 gnd 0.031169f
C41 minus.n11 gnd 0.031169f
C42 minus.t12 gnd 0.314894f
C43 minus.n12 gnd 0.143952f
C44 minus.t18 gnd 0.314894f
C45 minus.n13 gnd 0.143952f
C46 minus.n14 gnd 0.007073f
C47 minus.n15 gnd 0.031169f
C48 minus.n16 gnd 0.031169f
C49 minus.n17 gnd 0.031169f
C50 minus.n18 gnd 0.007073f
C51 minus.t16 gnd 0.314894f
C52 minus.n19 gnd 0.14376f
C53 minus.t6 gnd 0.314894f
C54 minus.n20 gnd 0.142318f
C55 minus.n21 gnd 0.352319f
C56 minus.n22 gnd 0.031169f
C57 minus.t17 gnd 0.314894f
C58 minus.t10 gnd 0.314894f
C59 minus.t5 gnd 0.314894f
C60 minus.n23 gnd 0.145585f
C61 minus.n24 gnd 0.031169f
C62 minus.t13 gnd 0.314894f
C63 minus.t9 gnd 0.314894f
C64 minus.n25 gnd 0.031169f
C65 minus.t19 gnd 0.314894f
C66 minus.n26 gnd 0.145585f
C67 minus.t20 gnd 0.32173f
C68 minus.n27 gnd 0.13571f
C69 minus.t7 gnd 0.314894f
C70 minus.n28 gnd 0.14376f
C71 minus.n29 gnd 0.007073f
C72 minus.n30 gnd 0.099236f
C73 minus.n31 gnd 0.031169f
C74 minus.n32 gnd 0.031169f
C75 minus.n33 gnd 0.007073f
C76 minus.n34 gnd 0.143952f
C77 minus.n35 gnd 0.143952f
C78 minus.n36 gnd 0.007073f
C79 minus.n37 gnd 0.031169f
C80 minus.n38 gnd 0.031169f
C81 minus.n39 gnd 0.031169f
C82 minus.n40 gnd 0.007073f
C83 minus.n41 gnd 0.14376f
C84 minus.n42 gnd 0.142318f
C85 minus.n43 gnd 0.838903f
C86 minus.n44 gnd 1.29085f
C87 minus.t2 gnd 0.009608f
C88 minus.t0 gnd 0.009608f
C89 minus.n45 gnd 0.031595f
C90 minus.t3 gnd 0.009608f
C91 minus.t4 gnd 0.009608f
C92 minus.n46 gnd 0.031162f
C93 minus.n47 gnd 0.265951f
C94 minus.t1 gnd 0.053479f
C95 minus.n48 gnd 0.145127f
C96 minus.n49 gnd 2.094f
C97 output.t5 gnd 0.464308f
C98 output.t16 gnd 0.044422f
C99 output.t19 gnd 0.044422f
C100 output.n0 gnd 0.364624f
C101 output.n1 gnd 0.614102f
C102 output.t9 gnd 0.044422f
C103 output.t8 gnd 0.044422f
C104 output.n2 gnd 0.364624f
C105 output.n3 gnd 0.350265f
C106 output.t14 gnd 0.044422f
C107 output.t18 gnd 0.044422f
C108 output.n4 gnd 0.364624f
C109 output.n5 gnd 0.350265f
C110 output.t6 gnd 0.044422f
C111 output.t10 gnd 0.044422f
C112 output.n6 gnd 0.364624f
C113 output.n7 gnd 0.350265f
C114 output.t11 gnd 0.044422f
C115 output.t17 gnd 0.044422f
C116 output.n8 gnd 0.364624f
C117 output.n9 gnd 0.350265f
C118 output.t4 gnd 0.044422f
C119 output.t12 gnd 0.044422f
C120 output.n10 gnd 0.364624f
C121 output.n11 gnd 0.350265f
C122 output.t15 gnd 0.044422f
C123 output.t13 gnd 0.044422f
C124 output.n12 gnd 0.364624f
C125 output.n13 gnd 0.350265f
C126 output.t7 gnd 0.462979f
C127 output.n14 gnd 0.28994f
C128 output.n15 gnd 0.015803f
C129 output.n16 gnd 0.011243f
C130 output.n17 gnd 0.006041f
C131 output.n18 gnd 0.01428f
C132 output.n19 gnd 0.006397f
C133 output.n20 gnd 0.011243f
C134 output.n21 gnd 0.006041f
C135 output.n22 gnd 0.01428f
C136 output.n23 gnd 0.006397f
C137 output.n24 gnd 0.048111f
C138 output.t1 gnd 0.023274f
C139 output.n25 gnd 0.01071f
C140 output.n26 gnd 0.008435f
C141 output.n27 gnd 0.006041f
C142 output.n28 gnd 0.267512f
C143 output.n29 gnd 0.011243f
C144 output.n30 gnd 0.006041f
C145 output.n31 gnd 0.006397f
C146 output.n32 gnd 0.01428f
C147 output.n33 gnd 0.01428f
C148 output.n34 gnd 0.006397f
C149 output.n35 gnd 0.006041f
C150 output.n36 gnd 0.011243f
C151 output.n37 gnd 0.011243f
C152 output.n38 gnd 0.006041f
C153 output.n39 gnd 0.006397f
C154 output.n40 gnd 0.01428f
C155 output.n41 gnd 0.030913f
C156 output.n42 gnd 0.006397f
C157 output.n43 gnd 0.006041f
C158 output.n44 gnd 0.025987f
C159 output.n45 gnd 0.097665f
C160 output.n46 gnd 0.015803f
C161 output.n47 gnd 0.011243f
C162 output.n48 gnd 0.006041f
C163 output.n49 gnd 0.01428f
C164 output.n50 gnd 0.006397f
C165 output.n51 gnd 0.011243f
C166 output.n52 gnd 0.006041f
C167 output.n53 gnd 0.01428f
C168 output.n54 gnd 0.006397f
C169 output.n55 gnd 0.048111f
C170 output.t2 gnd 0.023274f
C171 output.n56 gnd 0.01071f
C172 output.n57 gnd 0.008435f
C173 output.n58 gnd 0.006041f
C174 output.n59 gnd 0.267512f
C175 output.n60 gnd 0.011243f
C176 output.n61 gnd 0.006041f
C177 output.n62 gnd 0.006397f
C178 output.n63 gnd 0.01428f
C179 output.n64 gnd 0.01428f
C180 output.n65 gnd 0.006397f
C181 output.n66 gnd 0.006041f
C182 output.n67 gnd 0.011243f
C183 output.n68 gnd 0.011243f
C184 output.n69 gnd 0.006041f
C185 output.n70 gnd 0.006397f
C186 output.n71 gnd 0.01428f
C187 output.n72 gnd 0.030913f
C188 output.n73 gnd 0.006397f
C189 output.n74 gnd 0.006041f
C190 output.n75 gnd 0.025987f
C191 output.n76 gnd 0.09306f
C192 output.n77 gnd 1.65264f
C193 output.n78 gnd 0.015803f
C194 output.n79 gnd 0.011243f
C195 output.n80 gnd 0.006041f
C196 output.n81 gnd 0.01428f
C197 output.n82 gnd 0.006397f
C198 output.n83 gnd 0.011243f
C199 output.n84 gnd 0.006041f
C200 output.n85 gnd 0.01428f
C201 output.n86 gnd 0.006397f
C202 output.n87 gnd 0.048111f
C203 output.t3 gnd 0.023274f
C204 output.n88 gnd 0.01071f
C205 output.n89 gnd 0.008435f
C206 output.n90 gnd 0.006041f
C207 output.n91 gnd 0.267512f
C208 output.n92 gnd 0.011243f
C209 output.n93 gnd 0.006041f
C210 output.n94 gnd 0.006397f
C211 output.n95 gnd 0.01428f
C212 output.n96 gnd 0.01428f
C213 output.n97 gnd 0.006397f
C214 output.n98 gnd 0.006041f
C215 output.n99 gnd 0.011243f
C216 output.n100 gnd 0.011243f
C217 output.n101 gnd 0.006041f
C218 output.n102 gnd 0.006397f
C219 output.n103 gnd 0.01428f
C220 output.n104 gnd 0.030913f
C221 output.n105 gnd 0.006397f
C222 output.n106 gnd 0.006041f
C223 output.n107 gnd 0.025987f
C224 output.n108 gnd 0.09306f
C225 output.n109 gnd 0.713089f
C226 output.n110 gnd 0.015803f
C227 output.n111 gnd 0.011243f
C228 output.n112 gnd 0.006041f
C229 output.n113 gnd 0.01428f
C230 output.n114 gnd 0.006397f
C231 output.n115 gnd 0.011243f
C232 output.n116 gnd 0.006041f
C233 output.n117 gnd 0.01428f
C234 output.n118 gnd 0.006397f
C235 output.n119 gnd 0.048111f
C236 output.t0 gnd 0.023274f
C237 output.n120 gnd 0.01071f
C238 output.n121 gnd 0.008435f
C239 output.n122 gnd 0.006041f
C240 output.n123 gnd 0.267512f
C241 output.n124 gnd 0.011243f
C242 output.n125 gnd 0.006041f
C243 output.n126 gnd 0.006397f
C244 output.n127 gnd 0.01428f
C245 output.n128 gnd 0.01428f
C246 output.n129 gnd 0.006397f
C247 output.n130 gnd 0.006041f
C248 output.n131 gnd 0.011243f
C249 output.n132 gnd 0.011243f
C250 output.n133 gnd 0.006041f
C251 output.n134 gnd 0.006397f
C252 output.n135 gnd 0.01428f
C253 output.n136 gnd 0.030913f
C254 output.n137 gnd 0.006397f
C255 output.n138 gnd 0.006041f
C256 output.n139 gnd 0.025987f
C257 output.n140 gnd 0.09306f
C258 output.n141 gnd 1.67353f
C259 outputibias.t9 gnd 0.11477f
C260 outputibias.t10 gnd 0.115567f
C261 outputibias.n0 gnd 0.130108f
C262 outputibias.n1 gnd 0.001372f
C263 outputibias.n2 gnd 9.76e-19
C264 outputibias.n3 gnd 5.24e-19
C265 outputibias.n4 gnd 0.001239f
C266 outputibias.n5 gnd 5.55e-19
C267 outputibias.n6 gnd 9.76e-19
C268 outputibias.n7 gnd 5.24e-19
C269 outputibias.n8 gnd 0.001239f
C270 outputibias.n9 gnd 5.55e-19
C271 outputibias.n10 gnd 0.004176f
C272 outputibias.t7 gnd 0.00202f
C273 outputibias.n11 gnd 9.3e-19
C274 outputibias.n12 gnd 7.32e-19
C275 outputibias.n13 gnd 5.24e-19
C276 outputibias.n14 gnd 0.02322f
C277 outputibias.n15 gnd 9.76e-19
C278 outputibias.n16 gnd 5.24e-19
C279 outputibias.n17 gnd 5.55e-19
C280 outputibias.n18 gnd 0.001239f
C281 outputibias.n19 gnd 0.001239f
C282 outputibias.n20 gnd 5.55e-19
C283 outputibias.n21 gnd 5.24e-19
C284 outputibias.n22 gnd 9.76e-19
C285 outputibias.n23 gnd 9.76e-19
C286 outputibias.n24 gnd 5.24e-19
C287 outputibias.n25 gnd 5.55e-19
C288 outputibias.n26 gnd 0.001239f
C289 outputibias.n27 gnd 0.002683f
C290 outputibias.n28 gnd 5.55e-19
C291 outputibias.n29 gnd 5.24e-19
C292 outputibias.n30 gnd 0.002256f
C293 outputibias.n31 gnd 0.005781f
C294 outputibias.n32 gnd 0.001372f
C295 outputibias.n33 gnd 9.76e-19
C296 outputibias.n34 gnd 5.24e-19
C297 outputibias.n35 gnd 0.001239f
C298 outputibias.n36 gnd 5.55e-19
C299 outputibias.n37 gnd 9.76e-19
C300 outputibias.n38 gnd 5.24e-19
C301 outputibias.n39 gnd 0.001239f
C302 outputibias.n40 gnd 5.55e-19
C303 outputibias.n41 gnd 0.004176f
C304 outputibias.t1 gnd 0.00202f
C305 outputibias.n42 gnd 9.3e-19
C306 outputibias.n43 gnd 7.32e-19
C307 outputibias.n44 gnd 5.24e-19
C308 outputibias.n45 gnd 0.02322f
C309 outputibias.n46 gnd 9.76e-19
C310 outputibias.n47 gnd 5.24e-19
C311 outputibias.n48 gnd 5.55e-19
C312 outputibias.n49 gnd 0.001239f
C313 outputibias.n50 gnd 0.001239f
C314 outputibias.n51 gnd 5.55e-19
C315 outputibias.n52 gnd 5.24e-19
C316 outputibias.n53 gnd 9.76e-19
C317 outputibias.n54 gnd 9.76e-19
C318 outputibias.n55 gnd 5.24e-19
C319 outputibias.n56 gnd 5.55e-19
C320 outputibias.n57 gnd 0.001239f
C321 outputibias.n58 gnd 0.002683f
C322 outputibias.n59 gnd 5.55e-19
C323 outputibias.n60 gnd 5.24e-19
C324 outputibias.n61 gnd 0.002256f
C325 outputibias.n62 gnd 0.005197f
C326 outputibias.n63 gnd 0.121892f
C327 outputibias.n64 gnd 0.001372f
C328 outputibias.n65 gnd 9.76e-19
C329 outputibias.n66 gnd 5.24e-19
C330 outputibias.n67 gnd 0.001239f
C331 outputibias.n68 gnd 5.55e-19
C332 outputibias.n69 gnd 9.76e-19
C333 outputibias.n70 gnd 5.24e-19
C334 outputibias.n71 gnd 0.001239f
C335 outputibias.n72 gnd 5.55e-19
C336 outputibias.n73 gnd 0.004176f
C337 outputibias.t3 gnd 0.00202f
C338 outputibias.n74 gnd 9.3e-19
C339 outputibias.n75 gnd 7.32e-19
C340 outputibias.n76 gnd 5.24e-19
C341 outputibias.n77 gnd 0.02322f
C342 outputibias.n78 gnd 9.76e-19
C343 outputibias.n79 gnd 5.24e-19
C344 outputibias.n80 gnd 5.55e-19
C345 outputibias.n81 gnd 0.001239f
C346 outputibias.n82 gnd 0.001239f
C347 outputibias.n83 gnd 5.55e-19
C348 outputibias.n84 gnd 5.24e-19
C349 outputibias.n85 gnd 9.76e-19
C350 outputibias.n86 gnd 9.76e-19
C351 outputibias.n87 gnd 5.24e-19
C352 outputibias.n88 gnd 5.55e-19
C353 outputibias.n89 gnd 0.001239f
C354 outputibias.n90 gnd 0.002683f
C355 outputibias.n91 gnd 5.55e-19
C356 outputibias.n92 gnd 5.24e-19
C357 outputibias.n93 gnd 0.002256f
C358 outputibias.n94 gnd 0.005197f
C359 outputibias.n95 gnd 0.064513f
C360 outputibias.n96 gnd 0.001372f
C361 outputibias.n97 gnd 9.76e-19
C362 outputibias.n98 gnd 5.24e-19
C363 outputibias.n99 gnd 0.001239f
C364 outputibias.n100 gnd 5.55e-19
C365 outputibias.n101 gnd 9.76e-19
C366 outputibias.n102 gnd 5.24e-19
C367 outputibias.n103 gnd 0.001239f
C368 outputibias.n104 gnd 5.55e-19
C369 outputibias.n105 gnd 0.004176f
C370 outputibias.t5 gnd 0.00202f
C371 outputibias.n106 gnd 9.3e-19
C372 outputibias.n107 gnd 7.32e-19
C373 outputibias.n108 gnd 5.24e-19
C374 outputibias.n109 gnd 0.02322f
C375 outputibias.n110 gnd 9.76e-19
C376 outputibias.n111 gnd 5.24e-19
C377 outputibias.n112 gnd 5.55e-19
C378 outputibias.n113 gnd 0.001239f
C379 outputibias.n114 gnd 0.001239f
C380 outputibias.n115 gnd 5.55e-19
C381 outputibias.n116 gnd 5.24e-19
C382 outputibias.n117 gnd 9.76e-19
C383 outputibias.n118 gnd 9.76e-19
C384 outputibias.n119 gnd 5.24e-19
C385 outputibias.n120 gnd 5.55e-19
C386 outputibias.n121 gnd 0.001239f
C387 outputibias.n122 gnd 0.002683f
C388 outputibias.n123 gnd 5.55e-19
C389 outputibias.n124 gnd 5.24e-19
C390 outputibias.n125 gnd 0.002256f
C391 outputibias.n126 gnd 0.005197f
C392 outputibias.n127 gnd 0.084814f
C393 outputibias.t4 gnd 0.108319f
C394 outputibias.t2 gnd 0.108319f
C395 outputibias.t0 gnd 0.108319f
C396 outputibias.t6 gnd 0.109238f
C397 outputibias.n128 gnd 0.134674f
C398 outputibias.n129 gnd 0.07244f
C399 outputibias.n130 gnd 0.079818f
C400 outputibias.n131 gnd 0.164901f
C401 outputibias.t11 gnd 0.11477f
C402 outputibias.n132 gnd 0.067481f
C403 outputibias.t8 gnd 0.11477f
C404 outputibias.n133 gnd 0.065115f
C405 outputibias.n134 gnd 0.029159f
C406 plus.n0 gnd 0.022256f
C407 plus.t7 gnd 0.224852f
C408 plus.t15 gnd 0.224852f
C409 plus.t12 gnd 0.224852f
C410 plus.n1 gnd 0.103956f
C411 plus.n2 gnd 0.022256f
C412 plus.t18 gnd 0.224852f
C413 plus.n3 gnd 0.022256f
C414 plus.t14 gnd 0.224852f
C415 plus.t8 gnd 0.224852f
C416 plus.n4 gnd 0.103956f
C417 plus.t11 gnd 0.229734f
C418 plus.n5 gnd 0.096905f
C419 plus.t13 gnd 0.224852f
C420 plus.n6 gnd 0.102653f
C421 plus.n7 gnd 0.00505f
C422 plus.n8 gnd 0.07086f
C423 plus.n9 gnd 0.022256f
C424 plus.n10 gnd 0.022256f
C425 plus.n11 gnd 0.00505f
C426 plus.n12 gnd 0.10279f
C427 plus.n13 gnd 0.10279f
C428 plus.n14 gnd 0.00505f
C429 plus.n15 gnd 0.022256f
C430 plus.n16 gnd 0.022256f
C431 plus.n17 gnd 0.022256f
C432 plus.n18 gnd 0.00505f
C433 plus.n19 gnd 0.102653f
C434 plus.n20 gnd 0.101624f
C435 plus.n21 gnd 0.24583f
C436 plus.n22 gnd 0.022256f
C437 plus.t6 gnd 0.224852f
C438 plus.n23 gnd 0.103956f
C439 plus.n24 gnd 0.022256f
C440 plus.n25 gnd 0.00505f
C441 plus.t20 gnd 0.224852f
C442 plus.n26 gnd 0.07086f
C443 plus.t5 gnd 0.224852f
C444 plus.t19 gnd 0.229734f
C445 plus.n27 gnd 0.096905f
C446 plus.n28 gnd 0.102653f
C447 plus.n29 gnd 0.00505f
C448 plus.t17 gnd 0.224852f
C449 plus.n30 gnd 0.103956f
C450 plus.n31 gnd 0.022256f
C451 plus.n32 gnd 0.022256f
C452 plus.n33 gnd 0.022256f
C453 plus.n34 gnd 0.10279f
C454 plus.t10 gnd 0.224852f
C455 plus.n35 gnd 0.10279f
C456 plus.n36 gnd 0.00505f
C457 plus.n37 gnd 0.022256f
C458 plus.n38 gnd 0.022256f
C459 plus.n39 gnd 0.022256f
C460 plus.n40 gnd 0.00505f
C461 plus.t9 gnd 0.224852f
C462 plus.n41 gnd 0.102653f
C463 plus.t16 gnd 0.224852f
C464 plus.n42 gnd 0.101624f
C465 plus.n43 gnd 0.590081f
C466 plus.n44 gnd 0.912967f
C467 plus.t4 gnd 0.038421f
C468 plus.t0 gnd 0.006861f
C469 plus.t1 gnd 0.006861f
C470 plus.n45 gnd 0.022251f
C471 plus.n46 gnd 0.172738f
C472 plus.t3 gnd 0.006861f
C473 plus.t2 gnd 0.006861f
C474 plus.n47 gnd 0.022251f
C475 plus.n48 gnd 0.129661f
C476 plus.n49 gnd 2.32639f
C477 a_n1986_8322.t1 gnd 49.333103f
C478 a_n1986_8322.t0 gnd 75.3563f
C479 a_n1986_8322.t4 gnd 0.093486f
C480 a_n1986_8322.t3 gnd 0.875352f
C481 a_n1986_8322.t11 gnd 0.093486f
C482 a_n1986_8322.t6 gnd 0.093486f
C483 a_n1986_8322.n0 gnd 0.658513f
C484 a_n1986_8322.n1 gnd 0.735791f
C485 a_n1986_8322.t9 gnd 0.093486f
C486 a_n1986_8322.t8 gnd 0.093486f
C487 a_n1986_8322.n2 gnd 0.658513f
C488 a_n1986_8322.n3 gnd 0.373846f
C489 a_n1986_8322.t2 gnd 0.873609f
C490 a_n1986_8322.n4 gnd 1.39826f
C491 a_n1986_8322.t17 gnd 0.875352f
C492 a_n1986_8322.t21 gnd 0.093486f
C493 a_n1986_8322.t20 gnd 0.093486f
C494 a_n1986_8322.n5 gnd 0.658513f
C495 a_n1986_8322.n6 gnd 0.735791f
C496 a_n1986_8322.t15 gnd 0.873609f
C497 a_n1986_8322.n7 gnd 0.37026f
C498 a_n1986_8322.t18 gnd 0.873609f
C499 a_n1986_8322.n8 gnd 0.37026f
C500 a_n1986_8322.t16 gnd 0.093486f
C501 a_n1986_8322.t14 gnd 0.093486f
C502 a_n1986_8322.n9 gnd 0.658513f
C503 a_n1986_8322.n10 gnd 0.373846f
C504 a_n1986_8322.t19 gnd 0.873609f
C505 a_n1986_8322.n11 gnd 0.871879f
C506 a_n1986_8322.n12 gnd 1.58991f
C507 a_n1986_8322.n13 gnd 3.44798f
C508 a_n1986_8322.t5 gnd 0.873609f
C509 a_n1986_8322.n14 gnd 0.766135f
C510 a_n1986_8322.t12 gnd 0.875349f
C511 a_n1986_8322.t10 gnd 0.093486f
C512 a_n1986_8322.t7 gnd 0.093486f
C513 a_n1986_8322.n15 gnd 0.658513f
C514 a_n1986_8322.n16 gnd 0.735793f
C515 a_n1986_8322.n17 gnd 0.373844f
C516 a_n1986_8322.n18 gnd 0.658514f
C517 a_n1986_8322.t13 gnd 0.093486f
C518 a_n3827_n3924.n0 gnd 0.947295f
C519 a_n3827_n3924.n1 gnd 0.829256f
C520 a_n3827_n3924.t7 gnd 0.923252f
C521 a_n3827_n3924.n2 gnd 0.796733f
C522 a_n3827_n3924.t1 gnd 0.088833f
C523 a_n3827_n3924.t39 gnd 0.088833f
C524 a_n3827_n3924.n3 gnd 0.72551f
C525 a_n3827_n3924.n4 gnd 0.294242f
C526 a_n3827_n3924.t26 gnd 0.088833f
C527 a_n3827_n3924.t19 gnd 0.088833f
C528 a_n3827_n3924.n5 gnd 0.72551f
C529 a_n3827_n3924.n6 gnd 0.294242f
C530 a_n3827_n3924.t11 gnd 0.088833f
C531 a_n3827_n3924.t5 gnd 0.088833f
C532 a_n3827_n3924.n7 gnd 0.72551f
C533 a_n3827_n3924.n8 gnd 0.294242f
C534 a_n3827_n3924.t0 gnd 0.923252f
C535 a_n3827_n3924.n9 gnd 0.313344f
C536 a_n3827_n3924.t15 gnd 0.923252f
C537 a_n3827_n3924.n10 gnd 0.313344f
C538 a_n3827_n3924.t27 gnd 0.088833f
C539 a_n3827_n3924.t18 gnd 0.088833f
C540 a_n3827_n3924.n11 gnd 0.72551f
C541 a_n3827_n3924.n12 gnd 0.294242f
C542 a_n3827_n3924.t20 gnd 0.088833f
C543 a_n3827_n3924.t28 gnd 0.088833f
C544 a_n3827_n3924.n13 gnd 0.72551f
C545 a_n3827_n3924.n14 gnd 0.294242f
C546 a_n3827_n3924.t22 gnd 0.088833f
C547 a_n3827_n3924.t23 gnd 0.088833f
C548 a_n3827_n3924.n15 gnd 0.72551f
C549 a_n3827_n3924.n16 gnd 0.294242f
C550 a_n3827_n3924.t9 gnd 0.923249f
C551 a_n3827_n3924.n17 gnd 0.796737f
C552 a_n3827_n3924.t16 gnd 0.923249f
C553 a_n3827_n3924.n18 gnd 0.506437f
C554 a_n3827_n3924.t12 gnd 0.088833f
C555 a_n3827_n3924.t10 gnd 0.088833f
C556 a_n3827_n3924.n19 gnd 0.725509f
C557 a_n3827_n3924.n20 gnd 0.294243f
C558 a_n3827_n3924.t21 gnd 0.088833f
C559 a_n3827_n3924.t17 gnd 0.088833f
C560 a_n3827_n3924.n21 gnd 0.725509f
C561 a_n3827_n3924.n22 gnd 0.294243f
C562 a_n3827_n3924.t41 gnd 0.088833f
C563 a_n3827_n3924.t24 gnd 0.088833f
C564 a_n3827_n3924.n23 gnd 0.725509f
C565 a_n3827_n3924.n24 gnd 0.294243f
C566 a_n3827_n3924.t13 gnd 0.923249f
C567 a_n3827_n3924.n25 gnd 0.313347f
C568 a_n3827_n3924.t3 gnd 0.923249f
C569 a_n3827_n3924.n26 gnd 0.313347f
C570 a_n3827_n3924.t2 gnd 0.088833f
C571 a_n3827_n3924.t4 gnd 0.088833f
C572 a_n3827_n3924.n27 gnd 0.725509f
C573 a_n3827_n3924.n28 gnd 0.294243f
C574 a_n3827_n3924.t6 gnd 0.088833f
C575 a_n3827_n3924.t14 gnd 0.088833f
C576 a_n3827_n3924.n29 gnd 0.725509f
C577 a_n3827_n3924.n30 gnd 0.294243f
C578 a_n3827_n3924.t25 gnd 0.088833f
C579 a_n3827_n3924.t8 gnd 0.088833f
C580 a_n3827_n3924.n31 gnd 0.725509f
C581 a_n3827_n3924.n32 gnd 0.294243f
C582 a_n3827_n3924.t40 gnd 0.923249f
C583 a_n3827_n3924.n33 gnd 0.506437f
C584 a_n3827_n3924.n34 gnd 0.829256f
C585 a_n3827_n3924.t31 gnd 1.15026f
C586 a_n3827_n3924.t35 gnd 1.14712f
C587 a_n3827_n3924.n35 gnd 1.80223f
C588 a_n3827_n3924.t30 gnd 1.14712f
C589 a_n3827_n3924.t33 gnd 1.14712f
C590 a_n3827_n3924.n36 gnd 0.807936f
C591 a_n3827_n3924.t29 gnd 1.14712f
C592 a_n3827_n3924.n37 gnd 0.807936f
C593 a_n3827_n3924.t34 gnd 1.14712f
C594 a_n3827_n3924.n38 gnd 0.807936f
C595 a_n3827_n3924.t37 gnd 1.14712f
C596 a_n3827_n3924.n39 gnd 0.57544f
C597 a_n3827_n3924.n40 gnd 0.436676f
C598 a_n3827_n3924.t36 gnd 1.14712f
C599 a_n3827_n3924.n41 gnd 0.734847f
C600 a_n3827_n3924.t32 gnd 1.14712f
C601 a_n3827_n3924.n42 gnd 1.33048f
C602 a_n3827_n3924.t38 gnd 1.14876f
C603 diffpairibias.t27 gnd 0.090128f
C604 diffpairibias.t23 gnd 0.08996f
C605 diffpairibias.n0 gnd 0.105991f
C606 diffpairibias.t28 gnd 0.08996f
C607 diffpairibias.n1 gnd 0.051736f
C608 diffpairibias.t25 gnd 0.08996f
C609 diffpairibias.n2 gnd 0.051736f
C610 diffpairibias.t29 gnd 0.08996f
C611 diffpairibias.n3 gnd 0.041084f
C612 diffpairibias.t15 gnd 0.086371f
C613 diffpairibias.t1 gnd 0.085993f
C614 diffpairibias.n4 gnd 0.13579f
C615 diffpairibias.t11 gnd 0.085993f
C616 diffpairibias.n5 gnd 0.072463f
C617 diffpairibias.t13 gnd 0.085993f
C618 diffpairibias.n6 gnd 0.072463f
C619 diffpairibias.t7 gnd 0.085993f
C620 diffpairibias.n7 gnd 0.072463f
C621 diffpairibias.t3 gnd 0.085993f
C622 diffpairibias.n8 gnd 0.072463f
C623 diffpairibias.t17 gnd 0.085993f
C624 diffpairibias.n9 gnd 0.072463f
C625 diffpairibias.t5 gnd 0.085993f
C626 diffpairibias.n10 gnd 0.072463f
C627 diffpairibias.t19 gnd 0.085993f
C628 diffpairibias.n11 gnd 0.072463f
C629 diffpairibias.t9 gnd 0.085993f
C630 diffpairibias.n12 gnd 0.102883f
C631 diffpairibias.t14 gnd 0.086899f
C632 diffpairibias.t0 gnd 0.086748f
C633 diffpairibias.n13 gnd 0.094648f
C634 diffpairibias.t10 gnd 0.086748f
C635 diffpairibias.n14 gnd 0.052262f
C636 diffpairibias.t12 gnd 0.086748f
C637 diffpairibias.n15 gnd 0.052262f
C638 diffpairibias.t6 gnd 0.086748f
C639 diffpairibias.n16 gnd 0.052262f
C640 diffpairibias.t2 gnd 0.086748f
C641 diffpairibias.n17 gnd 0.052262f
C642 diffpairibias.t16 gnd 0.086748f
C643 diffpairibias.n18 gnd 0.052262f
C644 diffpairibias.t4 gnd 0.086748f
C645 diffpairibias.n19 gnd 0.052262f
C646 diffpairibias.t18 gnd 0.086748f
C647 diffpairibias.n20 gnd 0.052262f
C648 diffpairibias.t8 gnd 0.086748f
C649 diffpairibias.n21 gnd 0.061849f
C650 diffpairibias.n22 gnd 0.233513f
C651 diffpairibias.t20 gnd 0.08996f
C652 diffpairibias.n23 gnd 0.051747f
C653 diffpairibias.t26 gnd 0.08996f
C654 diffpairibias.n24 gnd 0.051736f
C655 diffpairibias.t22 gnd 0.08996f
C656 diffpairibias.n25 gnd 0.051736f
C657 diffpairibias.t21 gnd 0.08996f
C658 diffpairibias.n26 gnd 0.051736f
C659 diffpairibias.t24 gnd 0.08996f
C660 diffpairibias.n27 gnd 0.04729f
C661 diffpairibias.n28 gnd 0.047711f
C662 a_n1808_13878.t7 gnd 0.185195f
C663 a_n1808_13878.t2 gnd 0.185195f
C664 a_n1808_13878.t4 gnd 0.185195f
C665 a_n1808_13878.n0 gnd 1.4598f
C666 a_n1808_13878.t8 gnd 0.185195f
C667 a_n1808_13878.t3 gnd 0.185195f
C668 a_n1808_13878.n1 gnd 1.45825f
C669 a_n1808_13878.n2 gnd 2.03762f
C670 a_n1808_13878.t6 gnd 0.185195f
C671 a_n1808_13878.t1 gnd 0.185195f
C672 a_n1808_13878.n3 gnd 1.45825f
C673 a_n1808_13878.n4 gnd 3.69301f
C674 a_n1808_13878.t13 gnd 1.73408f
C675 a_n1808_13878.t16 gnd 0.185195f
C676 a_n1808_13878.t17 gnd 0.185195f
C677 a_n1808_13878.n5 gnd 1.30452f
C678 a_n1808_13878.n6 gnd 1.4576f
C679 a_n1808_13878.t12 gnd 1.73062f
C680 a_n1808_13878.n7 gnd 0.733487f
C681 a_n1808_13878.t15 gnd 1.73062f
C682 a_n1808_13878.n8 gnd 0.733487f
C683 a_n1808_13878.t18 gnd 0.185195f
C684 a_n1808_13878.t19 gnd 0.185195f
C685 a_n1808_13878.n9 gnd 1.30452f
C686 a_n1808_13878.n10 gnd 0.74059f
C687 a_n1808_13878.t14 gnd 1.73062f
C688 a_n1808_13878.n11 gnd 1.7272f
C689 a_n1808_13878.n12 gnd 2.51438f
C690 a_n1808_13878.t9 gnd 0.185195f
C691 a_n1808_13878.t10 gnd 0.185195f
C692 a_n1808_13878.n13 gnd 1.45825f
C693 a_n1808_13878.n14 gnd 1.80025f
C694 a_n1808_13878.t0 gnd 0.185195f
C695 a_n1808_13878.t5 gnd 0.185195f
C696 a_n1808_13878.n15 gnd 1.45825f
C697 a_n1808_13878.n16 gnd 1.31079f
C698 a_n1808_13878.n17 gnd 1.46067f
C699 a_n1808_13878.t11 gnd 0.185195f
C700 a_n1986_13878.n0 gnd 3.20192f
C701 a_n1986_13878.n1 gnd 0.64915f
C702 a_n1986_13878.n2 gnd 0.219304f
C703 a_n1986_13878.n3 gnd 0.286909f
C704 a_n1986_13878.n4 gnd 0.452885f
C705 a_n1986_13878.n5 gnd 0.674778f
C706 a_n1986_13878.n6 gnd 0.219304f
C707 a_n1986_13878.n7 gnd 0.286909f
C708 a_n1986_13878.n8 gnd 0.534226f
C709 a_n1986_13878.n9 gnd 0.208083f
C710 a_n1986_13878.n10 gnd 0.153257f
C711 a_n1986_13878.n11 gnd 0.240872f
C712 a_n1986_13878.n12 gnd 0.186046f
C713 a_n1986_13878.n13 gnd 0.208083f
C714 a_n1986_13878.n14 gnd 1.02197f
C715 a_n1986_13878.n15 gnd 0.153257f
C716 a_n1986_13878.n16 gnd 0.589052f
C717 a_n1986_13878.n17 gnd 0.439018f
C718 a_n1986_13878.n18 gnd 0.219304f
C719 a_n1986_13878.n19 gnd 0.500138f
C720 a_n1986_13878.n20 gnd 0.286909f
C721 a_n1986_13878.n21 gnd 0.445312f
C722 a_n1986_13878.n22 gnd 0.219304f
C723 a_n1986_13878.n23 gnd 0.742922f
C724 a_n1986_13878.n24 gnd 0.286909f
C725 a_n1986_13878.n25 gnd 1.19721f
C726 a_n1986_13878.n26 gnd 1.9455f
C727 a_n1986_13878.n27 gnd 1.1624f
C728 a_n1986_13878.n28 gnd 1.8055f
C729 a_n1986_13878.n29 gnd 2.46475f
C730 a_n1986_13878.n30 gnd 3.82161f
C731 a_n1986_13878.n31 gnd 3.20861f
C732 a_n1986_13878.n32 gnd 0.008491f
C733 a_n1986_13878.n34 gnd 0.290112f
C734 a_n1986_13878.n35 gnd 0.008491f
C735 a_n1986_13878.n37 gnd 0.290112f
C736 a_n1986_13878.n38 gnd 0.008491f
C737 a_n1986_13878.n39 gnd 0.2897f
C738 a_n1986_13878.n40 gnd 0.008491f
C739 a_n1986_13878.n41 gnd 0.2897f
C740 a_n1986_13878.n42 gnd 0.008491f
C741 a_n1986_13878.n43 gnd 0.2897f
C742 a_n1986_13878.n44 gnd 0.008491f
C743 a_n1986_13878.n45 gnd 0.2897f
C744 a_n1986_13878.n46 gnd 0.008491f
C745 a_n1986_13878.n48 gnd 0.290112f
C746 a_n1986_13878.n49 gnd 0.008491f
C747 a_n1986_13878.n51 gnd 0.290112f
C748 a_n1986_13878.t23 gnd 0.152112f
C749 a_n1986_13878.t30 gnd 0.722451f
C750 a_n1986_13878.t22 gnd 0.707549f
C751 a_n1986_13878.t10 gnd 0.707549f
C752 a_n1986_13878.t12 gnd 0.707549f
C753 a_n1986_13878.n52 gnd 0.311083f
C754 a_n1986_13878.t26 gnd 0.707549f
C755 a_n1986_13878.t14 gnd 0.719248f
C756 a_n1986_13878.t66 gnd 0.722451f
C757 a_n1986_13878.t49 gnd 0.707549f
C758 a_n1986_13878.t53 gnd 0.707549f
C759 a_n1986_13878.t43 gnd 0.707549f
C760 a_n1986_13878.n53 gnd 0.311083f
C761 a_n1986_13878.t58 gnd 0.707549f
C762 a_n1986_13878.t64 gnd 0.719248f
C763 a_n1986_13878.t19 gnd 1.4243f
C764 a_n1986_13878.t21 gnd 0.152112f
C765 a_n1986_13878.t25 gnd 0.152112f
C766 a_n1986_13878.n54 gnd 1.07147f
C767 a_n1986_13878.t17 gnd 0.152112f
C768 a_n1986_13878.t33 gnd 0.152112f
C769 a_n1986_13878.n55 gnd 1.07147f
C770 a_n1986_13878.t29 gnd 1.42146f
C771 a_n1986_13878.t16 gnd 0.707549f
C772 a_n1986_13878.n56 gnd 0.311083f
C773 a_n1986_13878.t32 gnd 0.707549f
C774 a_n1986_13878.t20 gnd 0.707549f
C775 a_n1986_13878.t48 gnd 0.707549f
C776 a_n1986_13878.n57 gnd 0.311083f
C777 a_n1986_13878.t57 gnd 0.707549f
C778 a_n1986_13878.t62 gnd 0.707549f
C779 a_n1986_13878.t61 gnd 0.722451f
C780 a_n1986_13878.n58 gnd 0.313741f
C781 a_n1986_13878.t41 gnd 0.707549f
C782 a_n1986_13878.n59 gnd 0.307133f
C783 a_n1986_13878.n60 gnd 0.313742f
C784 a_n1986_13878.t42 gnd 0.719248f
C785 a_n1986_13878.t18 gnd 0.722451f
C786 a_n1986_13878.n61 gnd 0.313741f
C787 a_n1986_13878.t24 gnd 0.707549f
C788 a_n1986_13878.n62 gnd 0.307133f
C789 a_n1986_13878.n63 gnd 0.313742f
C790 a_n1986_13878.t28 gnd 0.719248f
C791 a_n1986_13878.n64 gnd 1.14966f
C792 a_n1986_13878.t46 gnd 0.707549f
C793 a_n1986_13878.n65 gnd 0.307133f
C794 a_n1986_13878.t52 gnd 0.707549f
C795 a_n1986_13878.n66 gnd 0.307133f
C796 a_n1986_13878.t44 gnd 0.707549f
C797 a_n1986_13878.n67 gnd 0.307133f
C798 a_n1986_13878.t56 gnd 0.707549f
C799 a_n1986_13878.n68 gnd 0.307133f
C800 a_n1986_13878.t47 gnd 0.707549f
C801 a_n1986_13878.n69 gnd 0.301556f
C802 a_n1986_13878.t67 gnd 0.707549f
C803 a_n1986_13878.n70 gnd 0.311083f
C804 a_n1986_13878.t50 gnd 0.719405f
C805 a_n1986_13878.t59 gnd 0.707549f
C806 a_n1986_13878.n71 gnd 0.301556f
C807 a_n1986_13878.t45 gnd 0.707549f
C808 a_n1986_13878.n72 gnd 0.311083f
C809 a_n1986_13878.t54 gnd 0.719405f
C810 a_n1986_13878.t63 gnd 0.707549f
C811 a_n1986_13878.n73 gnd 0.301556f
C812 a_n1986_13878.t51 gnd 0.707549f
C813 a_n1986_13878.n74 gnd 0.311083f
C814 a_n1986_13878.t65 gnd 0.719405f
C815 a_n1986_13878.t55 gnd 0.707549f
C816 a_n1986_13878.n75 gnd 0.301556f
C817 a_n1986_13878.t40 gnd 0.707549f
C818 a_n1986_13878.n76 gnd 0.311083f
C819 a_n1986_13878.t60 gnd 0.719405f
C820 a_n1986_13878.n77 gnd 1.35928f
C821 a_n1986_13878.n78 gnd 0.313742f
C822 a_n1986_13878.n79 gnd 0.307133f
C823 a_n1986_13878.n80 gnd 0.313741f
C824 a_n1986_13878.t3 gnd 0.118309f
C825 a_n1986_13878.t2 gnd 0.118309f
C826 a_n1986_13878.n81 gnd 1.04709f
C827 a_n1986_13878.t4 gnd 0.118309f
C828 a_n1986_13878.t6 gnd 0.118309f
C829 a_n1986_13878.n82 gnd 1.04542f
C830 a_n1986_13878.t8 gnd 0.118309f
C831 a_n1986_13878.t39 gnd 0.118309f
C832 a_n1986_13878.n83 gnd 1.04709f
C833 a_n1986_13878.t34 gnd 0.118309f
C834 a_n1986_13878.t36 gnd 0.118309f
C835 a_n1986_13878.n84 gnd 1.04542f
C836 a_n1986_13878.t7 gnd 0.118309f
C837 a_n1986_13878.t1 gnd 0.118309f
C838 a_n1986_13878.n85 gnd 1.04542f
C839 a_n1986_13878.t38 gnd 0.118309f
C840 a_n1986_13878.t37 gnd 0.118309f
C841 a_n1986_13878.n86 gnd 1.04542f
C842 a_n1986_13878.t5 gnd 0.118309f
C843 a_n1986_13878.t0 gnd 0.118309f
C844 a_n1986_13878.n87 gnd 1.04709f
C845 a_n1986_13878.t35 gnd 0.118309f
C846 a_n1986_13878.t9 gnd 0.118309f
C847 a_n1986_13878.n88 gnd 1.04542f
C848 a_n1986_13878.n89 gnd 0.313742f
C849 a_n1986_13878.n90 gnd 0.307133f
C850 a_n1986_13878.n91 gnd 0.313741f
C851 a_n1986_13878.n92 gnd 0.799185f
C852 a_n1986_13878.t31 gnd 1.42146f
C853 a_n1986_13878.t15 gnd 1.4243f
C854 a_n1986_13878.t13 gnd 0.152112f
C855 a_n1986_13878.t27 gnd 0.152112f
C856 a_n1986_13878.n93 gnd 1.07147f
C857 a_n1986_13878.n94 gnd 1.07148f
C858 a_n1986_13878.t11 gnd 0.152112f
C859 CSoutput.n0 gnd 0.048923f
C860 CSoutput.t193 gnd 0.323618f
C861 CSoutput.n1 gnd 0.14613f
C862 CSoutput.n2 gnd 0.048923f
C863 CSoutput.t197 gnd 0.323618f
C864 CSoutput.n3 gnd 0.038776f
C865 CSoutput.n4 gnd 0.048923f
C866 CSoutput.t206 gnd 0.323618f
C867 CSoutput.n5 gnd 0.033437f
C868 CSoutput.n6 gnd 0.048923f
C869 CSoutput.t195 gnd 0.323618f
C870 CSoutput.t199 gnd 0.323618f
C871 CSoutput.n7 gnd 0.144537f
C872 CSoutput.n8 gnd 0.048923f
C873 CSoutput.t205 gnd 0.323618f
C874 CSoutput.n9 gnd 0.03188f
C875 CSoutput.n10 gnd 0.048923f
C876 CSoutput.t209 gnd 0.323618f
C877 CSoutput.t196 gnd 0.323618f
C878 CSoutput.n11 gnd 0.144537f
C879 CSoutput.n12 gnd 0.048923f
C880 CSoutput.t204 gnd 0.323618f
C881 CSoutput.n13 gnd 0.033437f
C882 CSoutput.n14 gnd 0.048923f
C883 CSoutput.t201 gnd 0.323618f
C884 CSoutput.t213 gnd 0.323618f
C885 CSoutput.n15 gnd 0.144537f
C886 CSoutput.n16 gnd 0.048923f
C887 CSoutput.t200 gnd 0.323618f
C888 CSoutput.n17 gnd 0.035712f
C889 CSoutput.t208 gnd 0.386732f
C890 CSoutput.t198 gnd 0.323618f
C891 CSoutput.n18 gnd 0.184518f
C892 CSoutput.n19 gnd 0.179046f
C893 CSoutput.n20 gnd 0.207715f
C894 CSoutput.n21 gnd 0.048923f
C895 CSoutput.n22 gnd 0.040832f
C896 CSoutput.n23 gnd 0.144537f
C897 CSoutput.n24 gnd 0.039361f
C898 CSoutput.n25 gnd 0.038776f
C899 CSoutput.n26 gnd 0.048923f
C900 CSoutput.n27 gnd 0.048923f
C901 CSoutput.n28 gnd 0.040518f
C902 CSoutput.n29 gnd 0.034401f
C903 CSoutput.n30 gnd 0.147755f
C904 CSoutput.n31 gnd 0.034875f
C905 CSoutput.n32 gnd 0.048923f
C906 CSoutput.n33 gnd 0.048923f
C907 CSoutput.n34 gnd 0.048923f
C908 CSoutput.n35 gnd 0.040087f
C909 CSoutput.n36 gnd 0.144537f
C910 CSoutput.n37 gnd 0.038337f
C911 CSoutput.n38 gnd 0.0398f
C912 CSoutput.n39 gnd 0.048923f
C913 CSoutput.n40 gnd 0.048923f
C914 CSoutput.n41 gnd 0.040824f
C915 CSoutput.n42 gnd 0.037313f
C916 CSoutput.n43 gnd 0.144537f
C917 CSoutput.n44 gnd 0.038259f
C918 CSoutput.n45 gnd 0.048923f
C919 CSoutput.n46 gnd 0.048923f
C920 CSoutput.n47 gnd 0.048923f
C921 CSoutput.n48 gnd 0.038259f
C922 CSoutput.n49 gnd 0.144537f
C923 CSoutput.n50 gnd 0.037313f
C924 CSoutput.n51 gnd 0.040824f
C925 CSoutput.n52 gnd 0.048923f
C926 CSoutput.n53 gnd 0.048923f
C927 CSoutput.n54 gnd 0.0398f
C928 CSoutput.n55 gnd 0.038337f
C929 CSoutput.n56 gnd 0.144537f
C930 CSoutput.n57 gnd 0.040087f
C931 CSoutput.n58 gnd 0.048923f
C932 CSoutput.n59 gnd 0.048923f
C933 CSoutput.n60 gnd 0.048923f
C934 CSoutput.n61 gnd 0.034875f
C935 CSoutput.n62 gnd 0.147755f
C936 CSoutput.n63 gnd 0.034401f
C937 CSoutput.t207 gnd 0.323618f
C938 CSoutput.n64 gnd 0.144537f
C939 CSoutput.n65 gnd 0.040518f
C940 CSoutput.n66 gnd 0.048923f
C941 CSoutput.n67 gnd 0.048923f
C942 CSoutput.n68 gnd 0.048923f
C943 CSoutput.n69 gnd 0.039361f
C944 CSoutput.n70 gnd 0.144537f
C945 CSoutput.n71 gnd 0.040832f
C946 CSoutput.n72 gnd 0.035712f
C947 CSoutput.n73 gnd 0.048923f
C948 CSoutput.n74 gnd 0.048923f
C949 CSoutput.n75 gnd 0.037036f
C950 CSoutput.n76 gnd 0.021996f
C951 CSoutput.t212 gnd 0.363608f
C952 CSoutput.n77 gnd 0.180626f
C953 CSoutput.n78 gnd 0.738931f
C954 CSoutput.t105 gnd 0.061025f
C955 CSoutput.t3 gnd 0.061025f
C956 CSoutput.n79 gnd 0.472477f
C957 CSoutput.t85 gnd 0.061025f
C958 CSoutput.t55 gnd 0.061025f
C959 CSoutput.n80 gnd 0.471634f
C960 CSoutput.n81 gnd 0.478708f
C961 CSoutput.t94 gnd 0.061025f
C962 CSoutput.t31 gnd 0.061025f
C963 CSoutput.n82 gnd 0.471634f
C964 CSoutput.n83 gnd 0.235887f
C965 CSoutput.t113 gnd 0.061025f
C966 CSoutput.t48 gnd 0.061025f
C967 CSoutput.n84 gnd 0.471634f
C968 CSoutput.n85 gnd 0.235887f
C969 CSoutput.t9 gnd 0.061025f
C970 CSoutput.t64 gnd 0.061025f
C971 CSoutput.n86 gnd 0.471634f
C972 CSoutput.n87 gnd 0.235887f
C973 CSoutput.t14 gnd 0.061025f
C974 CSoutput.t40 gnd 0.061025f
C975 CSoutput.n88 gnd 0.471634f
C976 CSoutput.n89 gnd 0.235887f
C977 CSoutput.t118 gnd 0.061025f
C978 CSoutput.t57 gnd 0.061025f
C979 CSoutput.n90 gnd 0.471634f
C980 CSoutput.n91 gnd 0.235887f
C981 CSoutput.t17 gnd 0.061025f
C982 CSoutput.t101 gnd 0.061025f
C983 CSoutput.n92 gnd 0.471634f
C984 CSoutput.n93 gnd 0.235887f
C985 CSoutput.t27 gnd 0.061025f
C986 CSoutput.t76 gnd 0.061025f
C987 CSoutput.n94 gnd 0.471634f
C988 CSoutput.n95 gnd 0.235887f
C989 CSoutput.t43 gnd 0.061025f
C990 CSoutput.t65 gnd 0.061025f
C991 CSoutput.n96 gnd 0.471634f
C992 CSoutput.n97 gnd 0.432562f
C993 CSoutput.t98 gnd 0.061025f
C994 CSoutput.t96 gnd 0.061025f
C995 CSoutput.n98 gnd 0.472477f
C996 CSoutput.t78 gnd 0.061025f
C997 CSoutput.t10 gnd 0.061025f
C998 CSoutput.n99 gnd 0.471634f
C999 CSoutput.n100 gnd 0.478708f
C1000 CSoutput.t4 gnd 0.061025f
C1001 CSoutput.t92 gnd 0.061025f
C1002 CSoutput.n101 gnd 0.471634f
C1003 CSoutput.n102 gnd 0.235887f
C1004 CSoutput.t77 gnd 0.061025f
C1005 CSoutput.t50 gnd 0.061025f
C1006 CSoutput.n103 gnd 0.471634f
C1007 CSoutput.n104 gnd 0.235887f
C1008 CSoutput.t32 gnd 0.061025f
C1009 CSoutput.t108 gnd 0.061025f
C1010 CSoutput.n105 gnd 0.471634f
C1011 CSoutput.n106 gnd 0.235887f
C1012 CSoutput.t74 gnd 0.061025f
C1013 CSoutput.t73 gnd 0.061025f
C1014 CSoutput.n107 gnd 0.471634f
C1015 CSoutput.n108 gnd 0.235887f
C1016 CSoutput.t61 gnd 0.061025f
C1017 CSoutput.t28 gnd 0.061025f
C1018 CSoutput.n109 gnd 0.471634f
C1019 CSoutput.n110 gnd 0.235887f
C1020 CSoutput.t8 gnd 0.061025f
C1021 CSoutput.t62 gnd 0.061025f
C1022 CSoutput.n111 gnd 0.471634f
C1023 CSoutput.n112 gnd 0.235887f
C1024 CSoutput.t58 gnd 0.061025f
C1025 CSoutput.t26 gnd 0.061025f
C1026 CSoutput.n113 gnd 0.471634f
C1027 CSoutput.n114 gnd 0.235887f
C1028 CSoutput.t5 gnd 0.061025f
C1029 CSoutput.t2 gnd 0.061025f
C1030 CSoutput.n115 gnd 0.471634f
C1031 CSoutput.n116 gnd 0.351767f
C1032 CSoutput.n117 gnd 0.443576f
C1033 CSoutput.t110 gnd 0.061025f
C1034 CSoutput.t109 gnd 0.061025f
C1035 CSoutput.n118 gnd 0.472477f
C1036 CSoutput.t89 gnd 0.061025f
C1037 CSoutput.t23 gnd 0.061025f
C1038 CSoutput.n119 gnd 0.471634f
C1039 CSoutput.n120 gnd 0.478708f
C1040 CSoutput.t19 gnd 0.061025f
C1041 CSoutput.t107 gnd 0.061025f
C1042 CSoutput.n121 gnd 0.471634f
C1043 CSoutput.n122 gnd 0.235887f
C1044 CSoutput.t86 gnd 0.061025f
C1045 CSoutput.t63 gnd 0.061025f
C1046 CSoutput.n123 gnd 0.471634f
C1047 CSoutput.n124 gnd 0.235887f
C1048 CSoutput.t44 gnd 0.061025f
C1049 CSoutput.t119 gnd 0.061025f
C1050 CSoutput.n125 gnd 0.471634f
C1051 CSoutput.n126 gnd 0.235887f
C1052 CSoutput.t84 gnd 0.061025f
C1053 CSoutput.t83 gnd 0.061025f
C1054 CSoutput.n127 gnd 0.471634f
C1055 CSoutput.n128 gnd 0.235887f
C1056 CSoutput.t71 gnd 0.061025f
C1057 CSoutput.t41 gnd 0.061025f
C1058 CSoutput.n129 gnd 0.471634f
C1059 CSoutput.n130 gnd 0.235887f
C1060 CSoutput.t22 gnd 0.061025f
C1061 CSoutput.t72 gnd 0.061025f
C1062 CSoutput.n131 gnd 0.471634f
C1063 CSoutput.n132 gnd 0.235887f
C1064 CSoutput.t68 gnd 0.061025f
C1065 CSoutput.t39 gnd 0.061025f
C1066 CSoutput.n133 gnd 0.471634f
C1067 CSoutput.n134 gnd 0.235887f
C1068 CSoutput.t20 gnd 0.061025f
C1069 CSoutput.t18 gnd 0.061025f
C1070 CSoutput.n135 gnd 0.471634f
C1071 CSoutput.n136 gnd 0.351767f
C1072 CSoutput.n137 gnd 0.495804f
C1073 CSoutput.n138 gnd 9.09012f
C1074 CSoutput.n140 gnd 0.865447f
C1075 CSoutput.n141 gnd 0.649085f
C1076 CSoutput.n142 gnd 0.865447f
C1077 CSoutput.n143 gnd 0.865447f
C1078 CSoutput.n144 gnd 2.33005f
C1079 CSoutput.n145 gnd 0.865447f
C1080 CSoutput.n146 gnd 0.865447f
C1081 CSoutput.t202 gnd 1.08181f
C1082 CSoutput.n147 gnd 0.865447f
C1083 CSoutput.n148 gnd 0.865447f
C1084 CSoutput.n152 gnd 0.865447f
C1085 CSoutput.n156 gnd 0.865447f
C1086 CSoutput.n157 gnd 0.865447f
C1087 CSoutput.n159 gnd 0.865447f
C1088 CSoutput.n164 gnd 0.865447f
C1089 CSoutput.n166 gnd 0.865447f
C1090 CSoutput.n167 gnd 0.865447f
C1091 CSoutput.n169 gnd 0.865447f
C1092 CSoutput.n170 gnd 0.865447f
C1093 CSoutput.n172 gnd 0.865447f
C1094 CSoutput.t192 gnd 14.4615f
C1095 CSoutput.n174 gnd 0.865447f
C1096 CSoutput.n175 gnd 0.649085f
C1097 CSoutput.n176 gnd 0.865447f
C1098 CSoutput.n177 gnd 0.865447f
C1099 CSoutput.n178 gnd 2.33005f
C1100 CSoutput.n179 gnd 0.865447f
C1101 CSoutput.n180 gnd 0.865447f
C1102 CSoutput.t210 gnd 1.08181f
C1103 CSoutput.n181 gnd 0.865447f
C1104 CSoutput.n182 gnd 0.865447f
C1105 CSoutput.n186 gnd 0.865447f
C1106 CSoutput.n190 gnd 0.865447f
C1107 CSoutput.n191 gnd 0.865447f
C1108 CSoutput.n193 gnd 0.865447f
C1109 CSoutput.n198 gnd 0.865447f
C1110 CSoutput.n200 gnd 0.865447f
C1111 CSoutput.n201 gnd 0.865447f
C1112 CSoutput.n203 gnd 0.865447f
C1113 CSoutput.n204 gnd 0.865447f
C1114 CSoutput.n206 gnd 0.865447f
C1115 CSoutput.n207 gnd 0.649085f
C1116 CSoutput.n209 gnd 0.865447f
C1117 CSoutput.n210 gnd 0.649085f
C1118 CSoutput.n211 gnd 0.865447f
C1119 CSoutput.n212 gnd 0.865447f
C1120 CSoutput.n213 gnd 2.33005f
C1121 CSoutput.n214 gnd 0.865447f
C1122 CSoutput.n215 gnd 0.865447f
C1123 CSoutput.t203 gnd 1.08181f
C1124 CSoutput.n216 gnd 0.865447f
C1125 CSoutput.n217 gnd 2.33005f
C1126 CSoutput.n219 gnd 0.865447f
C1127 CSoutput.n220 gnd 0.865447f
C1128 CSoutput.n222 gnd 0.865447f
C1129 CSoutput.n223 gnd 0.865447f
C1130 CSoutput.t211 gnd 14.2258f
C1131 CSoutput.t194 gnd 14.4615f
C1132 CSoutput.n229 gnd 2.71503f
C1133 CSoutput.n230 gnd 11.0601f
C1134 CSoutput.n231 gnd 11.522901f
C1135 CSoutput.n236 gnd 2.94111f
C1136 CSoutput.n242 gnd 0.865447f
C1137 CSoutput.n244 gnd 0.865447f
C1138 CSoutput.n246 gnd 0.865447f
C1139 CSoutput.n248 gnd 0.865447f
C1140 CSoutput.n250 gnd 0.865447f
C1141 CSoutput.n256 gnd 0.865447f
C1142 CSoutput.n263 gnd 1.58776f
C1143 CSoutput.n264 gnd 1.58776f
C1144 CSoutput.n265 gnd 0.865447f
C1145 CSoutput.n266 gnd 0.865447f
C1146 CSoutput.n268 gnd 0.649085f
C1147 CSoutput.n269 gnd 0.555883f
C1148 CSoutput.n271 gnd 0.649085f
C1149 CSoutput.n272 gnd 0.555883f
C1150 CSoutput.n273 gnd 0.649085f
C1151 CSoutput.n275 gnd 0.865447f
C1152 CSoutput.n277 gnd 2.33005f
C1153 CSoutput.n278 gnd 2.71503f
C1154 CSoutput.n279 gnd 10.1724f
C1155 CSoutput.n281 gnd 0.649085f
C1156 CSoutput.n282 gnd 1.67014f
C1157 CSoutput.n283 gnd 0.649085f
C1158 CSoutput.n285 gnd 0.865447f
C1159 CSoutput.n287 gnd 2.33005f
C1160 CSoutput.n288 gnd 5.07522f
C1161 CSoutput.t1 gnd 0.061025f
C1162 CSoutput.t104 gnd 0.061025f
C1163 CSoutput.n289 gnd 0.472477f
C1164 CSoutput.t54 gnd 0.061025f
C1165 CSoutput.t117 gnd 0.061025f
C1166 CSoutput.n290 gnd 0.471634f
C1167 CSoutput.n291 gnd 0.478708f
C1168 CSoutput.t30 gnd 0.061025f
C1169 CSoutput.t93 gnd 0.061025f
C1170 CSoutput.n292 gnd 0.471634f
C1171 CSoutput.n293 gnd 0.235887f
C1172 CSoutput.t47 gnd 0.061025f
C1173 CSoutput.t112 gnd 0.061025f
C1174 CSoutput.n294 gnd 0.471634f
C1175 CSoutput.n295 gnd 0.235887f
C1176 CSoutput.t87 gnd 0.061025f
C1177 CSoutput.t7 gnd 0.061025f
C1178 CSoutput.n296 gnd 0.471634f
C1179 CSoutput.n297 gnd 0.235887f
C1180 CSoutput.t38 gnd 0.061025f
C1181 CSoutput.t13 gnd 0.061025f
C1182 CSoutput.n298 gnd 0.471634f
C1183 CSoutput.n299 gnd 0.235887f
C1184 CSoutput.t56 gnd 0.061025f
C1185 CSoutput.t35 gnd 0.061025f
C1186 CSoutput.n300 gnd 0.471634f
C1187 CSoutput.n301 gnd 0.235887f
C1188 CSoutput.t100 gnd 0.061025f
C1189 CSoutput.t16 gnd 0.061025f
C1190 CSoutput.n302 gnd 0.471634f
C1191 CSoutput.n303 gnd 0.235887f
C1192 CSoutput.t75 gnd 0.061025f
C1193 CSoutput.t24 gnd 0.061025f
C1194 CSoutput.n304 gnd 0.471634f
C1195 CSoutput.n305 gnd 0.235887f
C1196 CSoutput.t88 gnd 0.061025f
C1197 CSoutput.t42 gnd 0.061025f
C1198 CSoutput.n306 gnd 0.471634f
C1199 CSoutput.n307 gnd 0.432562f
C1200 CSoutput.t59 gnd 0.061025f
C1201 CSoutput.t60 gnd 0.061025f
C1202 CSoutput.n308 gnd 0.472477f
C1203 CSoutput.t82 gnd 0.061025f
C1204 CSoutput.t6 gnd 0.061025f
C1205 CSoutput.n309 gnd 0.471634f
C1206 CSoutput.n310 gnd 0.478708f
C1207 CSoutput.t53 gnd 0.061025f
C1208 CSoutput.t80 gnd 0.061025f
C1209 CSoutput.n311 gnd 0.471634f
C1210 CSoutput.n312 gnd 0.235887f
C1211 CSoutput.t0 gnd 0.061025f
C1212 CSoutput.t36 gnd 0.061025f
C1213 CSoutput.n313 gnd 0.471634f
C1214 CSoutput.n314 gnd 0.235887f
C1215 CSoutput.t37 gnd 0.061025f
C1216 CSoutput.t106 gnd 0.061025f
C1217 CSoutput.n315 gnd 0.471634f
C1218 CSoutput.n316 gnd 0.235887f
C1219 CSoutput.t33 gnd 0.061025f
C1220 CSoutput.t34 gnd 0.061025f
C1221 CSoutput.n317 gnd 0.471634f
C1222 CSoutput.n318 gnd 0.235887f
C1223 CSoutput.t102 gnd 0.061025f
C1224 CSoutput.t103 gnd 0.061025f
C1225 CSoutput.n319 gnd 0.471634f
C1226 CSoutput.n320 gnd 0.235887f
C1227 CSoutput.t12 gnd 0.061025f
C1228 CSoutput.t81 gnd 0.061025f
C1229 CSoutput.n321 gnd 0.471634f
C1230 CSoutput.n322 gnd 0.235887f
C1231 CSoutput.t99 gnd 0.061025f
C1232 CSoutput.t11 gnd 0.061025f
C1233 CSoutput.n323 gnd 0.471634f
C1234 CSoutput.n324 gnd 0.235887f
C1235 CSoutput.t52 gnd 0.061025f
C1236 CSoutput.t79 gnd 0.061025f
C1237 CSoutput.n325 gnd 0.471634f
C1238 CSoutput.n326 gnd 0.351767f
C1239 CSoutput.n327 gnd 0.443576f
C1240 CSoutput.t69 gnd 0.061025f
C1241 CSoutput.t70 gnd 0.061025f
C1242 CSoutput.n328 gnd 0.472477f
C1243 CSoutput.t97 gnd 0.061025f
C1244 CSoutput.t21 gnd 0.061025f
C1245 CSoutput.n329 gnd 0.471634f
C1246 CSoutput.n330 gnd 0.478708f
C1247 CSoutput.t66 gnd 0.061025f
C1248 CSoutput.t90 gnd 0.061025f
C1249 CSoutput.n331 gnd 0.471634f
C1250 CSoutput.n332 gnd 0.235887f
C1251 CSoutput.t15 gnd 0.061025f
C1252 CSoutput.t49 gnd 0.061025f
C1253 CSoutput.n333 gnd 0.471634f
C1254 CSoutput.n334 gnd 0.235887f
C1255 CSoutput.t51 gnd 0.061025f
C1256 CSoutput.t116 gnd 0.061025f
C1257 CSoutput.n335 gnd 0.471634f
C1258 CSoutput.n336 gnd 0.235887f
C1259 CSoutput.t45 gnd 0.061025f
C1260 CSoutput.t46 gnd 0.061025f
C1261 CSoutput.n337 gnd 0.471634f
C1262 CSoutput.n338 gnd 0.235887f
C1263 CSoutput.t114 gnd 0.061025f
C1264 CSoutput.t115 gnd 0.061025f
C1265 CSoutput.n339 gnd 0.471634f
C1266 CSoutput.n340 gnd 0.235887f
C1267 CSoutput.t29 gnd 0.061025f
C1268 CSoutput.t95 gnd 0.061025f
C1269 CSoutput.n341 gnd 0.471634f
C1270 CSoutput.n342 gnd 0.235887f
C1271 CSoutput.t111 gnd 0.061025f
C1272 CSoutput.t25 gnd 0.061025f
C1273 CSoutput.n343 gnd 0.471634f
C1274 CSoutput.n344 gnd 0.235887f
C1275 CSoutput.t67 gnd 0.061025f
C1276 CSoutput.t91 gnd 0.061025f
C1277 CSoutput.n345 gnd 0.471632f
C1278 CSoutput.n346 gnd 0.351769f
C1279 CSoutput.n347 gnd 0.495804f
C1280 CSoutput.n348 gnd 13.025901f
C1281 CSoutput.t182 gnd 0.053397f
C1282 CSoutput.t129 gnd 0.053397f
C1283 CSoutput.n349 gnd 0.473413f
C1284 CSoutput.t169 gnd 0.053397f
C1285 CSoutput.t122 gnd 0.053397f
C1286 CSoutput.n350 gnd 0.471834f
C1287 CSoutput.n351 gnd 0.439661f
C1288 CSoutput.t154 gnd 0.053397f
C1289 CSoutput.t185 gnd 0.053397f
C1290 CSoutput.n352 gnd 0.471834f
C1291 CSoutput.n353 gnd 0.216732f
C1292 CSoutput.t142 gnd 0.053397f
C1293 CSoutput.t153 gnd 0.053397f
C1294 CSoutput.n354 gnd 0.471834f
C1295 CSoutput.n355 gnd 0.216732f
C1296 CSoutput.t124 gnd 0.053397f
C1297 CSoutput.t159 gnd 0.053397f
C1298 CSoutput.n356 gnd 0.471834f
C1299 CSoutput.n357 gnd 0.216732f
C1300 CSoutput.t173 gnd 0.053397f
C1301 CSoutput.t143 gnd 0.053397f
C1302 CSoutput.n358 gnd 0.471834f
C1303 CSoutput.n359 gnd 0.399751f
C1304 CSoutput.t151 gnd 0.053397f
C1305 CSoutput.t134 gnd 0.053397f
C1306 CSoutput.n360 gnd 0.473413f
C1307 CSoutput.t138 gnd 0.053397f
C1308 CSoutput.t150 gnd 0.053397f
C1309 CSoutput.n361 gnd 0.471834f
C1310 CSoutput.n362 gnd 0.439661f
C1311 CSoutput.t133 gnd 0.053397f
C1312 CSoutput.t140 gnd 0.053397f
C1313 CSoutput.n363 gnd 0.471834f
C1314 CSoutput.n364 gnd 0.216732f
C1315 CSoutput.t152 gnd 0.053397f
C1316 CSoutput.t132 gnd 0.053397f
C1317 CSoutput.n365 gnd 0.471834f
C1318 CSoutput.n366 gnd 0.216732f
C1319 CSoutput.t139 gnd 0.053397f
C1320 CSoutput.t127 gnd 0.053397f
C1321 CSoutput.n367 gnd 0.471834f
C1322 CSoutput.n368 gnd 0.216732f
C1323 CSoutput.t131 gnd 0.053397f
C1324 CSoutput.t141 gnd 0.053397f
C1325 CSoutput.n369 gnd 0.471834f
C1326 CSoutput.n370 gnd 0.329046f
C1327 CSoutput.n371 gnd 0.415029f
C1328 CSoutput.t128 gnd 0.053397f
C1329 CSoutput.t189 gnd 0.053397f
C1330 CSoutput.n372 gnd 0.473413f
C1331 CSoutput.t180 gnd 0.053397f
C1332 CSoutput.t135 gnd 0.053397f
C1333 CSoutput.n373 gnd 0.471834f
C1334 CSoutput.n374 gnd 0.439661f
C1335 CSoutput.t120 gnd 0.053397f
C1336 CSoutput.t186 gnd 0.053397f
C1337 CSoutput.n375 gnd 0.471834f
C1338 CSoutput.n376 gnd 0.216732f
C1339 CSoutput.t146 gnd 0.053397f
C1340 CSoutput.t155 gnd 0.053397f
C1341 CSoutput.n377 gnd 0.471834f
C1342 CSoutput.n378 gnd 0.216732f
C1343 CSoutput.t190 gnd 0.053397f
C1344 CSoutput.t179 gnd 0.053397f
C1345 CSoutput.n379 gnd 0.471834f
C1346 CSoutput.n380 gnd 0.216732f
C1347 CSoutput.t164 gnd 0.053397f
C1348 CSoutput.t121 gnd 0.053397f
C1349 CSoutput.n381 gnd 0.471834f
C1350 CSoutput.n382 gnd 0.329046f
C1351 CSoutput.n383 gnd 0.445676f
C1352 CSoutput.n384 gnd 13.3417f
C1353 CSoutput.t161 gnd 0.053397f
C1354 CSoutput.t125 gnd 0.053397f
C1355 CSoutput.n385 gnd 0.473413f
C1356 CSoutput.t145 gnd 0.053397f
C1357 CSoutput.t187 gnd 0.053397f
C1358 CSoutput.n386 gnd 0.471834f
C1359 CSoutput.n387 gnd 0.439661f
C1360 CSoutput.t126 gnd 0.053397f
C1361 CSoutput.t175 gnd 0.053397f
C1362 CSoutput.n388 gnd 0.471834f
C1363 CSoutput.n389 gnd 0.216732f
C1364 CSoutput.t174 gnd 0.053397f
C1365 CSoutput.t163 gnd 0.053397f
C1366 CSoutput.n390 gnd 0.471834f
C1367 CSoutput.n391 gnd 0.216732f
C1368 CSoutput.t176 gnd 0.053397f
C1369 CSoutput.t147 gnd 0.053397f
C1370 CSoutput.n392 gnd 0.471834f
C1371 CSoutput.n393 gnd 0.216732f
C1372 CSoutput.t170 gnd 0.053397f
C1373 CSoutput.t181 gnd 0.053397f
C1374 CSoutput.n394 gnd 0.471834f
C1375 CSoutput.n395 gnd 0.399751f
C1376 CSoutput.t148 gnd 0.053397f
C1377 CSoutput.t165 gnd 0.053397f
C1378 CSoutput.n396 gnd 0.473413f
C1379 CSoutput.t166 gnd 0.053397f
C1380 CSoutput.t157 gnd 0.053397f
C1381 CSoutput.n397 gnd 0.471834f
C1382 CSoutput.n398 gnd 0.439661f
C1383 CSoutput.t156 gnd 0.053397f
C1384 CSoutput.t149 gnd 0.053397f
C1385 CSoutput.n399 gnd 0.471834f
C1386 CSoutput.n400 gnd 0.216732f
C1387 CSoutput.t144 gnd 0.053397f
C1388 CSoutput.t136 gnd 0.053397f
C1389 CSoutput.n401 gnd 0.471834f
C1390 CSoutput.n402 gnd 0.216732f
C1391 CSoutput.t137 gnd 0.053397f
C1392 CSoutput.t158 gnd 0.053397f
C1393 CSoutput.n403 gnd 0.471834f
C1394 CSoutput.n404 gnd 0.216732f
C1395 CSoutput.t160 gnd 0.053397f
C1396 CSoutput.t123 gnd 0.053397f
C1397 CSoutput.n405 gnd 0.471834f
C1398 CSoutput.n406 gnd 0.329046f
C1399 CSoutput.n407 gnd 0.415029f
C1400 CSoutput.t177 gnd 0.053397f
C1401 CSoutput.t188 gnd 0.053397f
C1402 CSoutput.n408 gnd 0.473413f
C1403 CSoutput.t191 gnd 0.053397f
C1404 CSoutput.t168 gnd 0.053397f
C1405 CSoutput.n409 gnd 0.471834f
C1406 CSoutput.n410 gnd 0.439661f
C1407 CSoutput.t172 gnd 0.053397f
C1408 CSoutput.t183 gnd 0.053397f
C1409 CSoutput.n411 gnd 0.471834f
C1410 CSoutput.n412 gnd 0.216732f
C1411 CSoutput.t130 gnd 0.053397f
C1412 CSoutput.t162 gnd 0.053397f
C1413 CSoutput.n413 gnd 0.471834f
C1414 CSoutput.n414 gnd 0.216732f
C1415 CSoutput.t167 gnd 0.053397f
C1416 CSoutput.t178 gnd 0.053397f
C1417 CSoutput.n415 gnd 0.471834f
C1418 CSoutput.n416 gnd 0.216732f
C1419 CSoutput.t184 gnd 0.053397f
C1420 CSoutput.t171 gnd 0.053397f
C1421 CSoutput.n417 gnd 0.471834f
C1422 CSoutput.n418 gnd 0.329046f
C1423 CSoutput.n419 gnd 0.445676f
C1424 CSoutput.n420 gnd 7.67865f
C1425 CSoutput.n421 gnd 14.832201f
C1426 vdd.t288 gnd 0.040769f
C1427 vdd.t207 gnd 0.040769f
C1428 vdd.n0 gnd 0.321549f
C1429 vdd.t3 gnd 0.040769f
C1430 vdd.t290 gnd 0.040769f
C1431 vdd.n1 gnd 0.321019f
C1432 vdd.n2 gnd 0.29604f
C1433 vdd.t7 gnd 0.040769f
C1434 vdd.t293 gnd 0.040769f
C1435 vdd.n3 gnd 0.321019f
C1436 vdd.n4 gnd 0.149719f
C1437 vdd.t205 gnd 0.040769f
C1438 vdd.t197 gnd 0.040769f
C1439 vdd.n5 gnd 0.321019f
C1440 vdd.n6 gnd 0.140483f
C1441 vdd.t186 gnd 0.040769f
C1442 vdd.t191 gnd 0.040769f
C1443 vdd.n7 gnd 0.321549f
C1444 vdd.t1 gnd 0.040769f
C1445 vdd.t13 gnd 0.040769f
C1446 vdd.n8 gnd 0.321019f
C1447 vdd.n9 gnd 0.29604f
C1448 vdd.t201 gnd 0.040769f
C1449 vdd.t177 gnd 0.040769f
C1450 vdd.n10 gnd 0.321019f
C1451 vdd.n11 gnd 0.149719f
C1452 vdd.t295 gnd 0.040769f
C1453 vdd.t194 gnd 0.040769f
C1454 vdd.n12 gnd 0.321019f
C1455 vdd.n13 gnd 0.140483f
C1456 vdd.n14 gnd 0.099319f
C1457 vdd.t291 gnd 0.022649f
C1458 vdd.t188 gnd 0.022649f
C1459 vdd.n15 gnd 0.208477f
C1460 vdd.t209 gnd 0.022649f
C1461 vdd.t8 gnd 0.022649f
C1462 vdd.n16 gnd 0.207867f
C1463 vdd.n17 gnd 0.361754f
C1464 vdd.t174 gnd 0.022649f
C1465 vdd.t208 gnd 0.022649f
C1466 vdd.n18 gnd 0.207867f
C1467 vdd.n19 gnd 0.149662f
C1468 vdd.t210 gnd 0.022649f
C1469 vdd.t9 gnd 0.022649f
C1470 vdd.n20 gnd 0.208477f
C1471 vdd.t180 gnd 0.022649f
C1472 vdd.t189 gnd 0.022649f
C1473 vdd.n21 gnd 0.207867f
C1474 vdd.n22 gnd 0.361754f
C1475 vdd.t181 gnd 0.022649f
C1476 vdd.t202 gnd 0.022649f
C1477 vdd.n23 gnd 0.207867f
C1478 vdd.n24 gnd 0.149662f
C1479 vdd.t175 gnd 0.022649f
C1480 vdd.t199 gnd 0.022649f
C1481 vdd.n25 gnd 0.207867f
C1482 vdd.t203 gnd 0.022649f
C1483 vdd.t10 gnd 0.022649f
C1484 vdd.n26 gnd 0.207867f
C1485 vdd.n27 gnd 22.7579f
C1486 vdd.n28 gnd 8.6933f
C1487 vdd.n29 gnd 0.006177f
C1488 vdd.n30 gnd 0.005732f
C1489 vdd.n31 gnd 0.003171f
C1490 vdd.n32 gnd 0.007281f
C1491 vdd.n33 gnd 0.00308f
C1492 vdd.n34 gnd 0.003262f
C1493 vdd.n35 gnd 0.005732f
C1494 vdd.n36 gnd 0.00308f
C1495 vdd.n37 gnd 0.007281f
C1496 vdd.n38 gnd 0.003262f
C1497 vdd.n39 gnd 0.005732f
C1498 vdd.n40 gnd 0.00308f
C1499 vdd.n41 gnd 0.005461f
C1500 vdd.n42 gnd 0.005477f
C1501 vdd.t18 gnd 0.015642f
C1502 vdd.n43 gnd 0.034803f
C1503 vdd.n44 gnd 0.181124f
C1504 vdd.n45 gnd 0.00308f
C1505 vdd.n46 gnd 0.003262f
C1506 vdd.n47 gnd 0.007281f
C1507 vdd.n48 gnd 0.007281f
C1508 vdd.n49 gnd 0.003262f
C1509 vdd.n50 gnd 0.00308f
C1510 vdd.n51 gnd 0.005732f
C1511 vdd.n52 gnd 0.005732f
C1512 vdd.n53 gnd 0.00308f
C1513 vdd.n54 gnd 0.003262f
C1514 vdd.n55 gnd 0.007281f
C1515 vdd.n56 gnd 0.007281f
C1516 vdd.n57 gnd 0.003262f
C1517 vdd.n58 gnd 0.00308f
C1518 vdd.n59 gnd 0.005732f
C1519 vdd.n60 gnd 0.005732f
C1520 vdd.n61 gnd 0.00308f
C1521 vdd.n62 gnd 0.003262f
C1522 vdd.n63 gnd 0.007281f
C1523 vdd.n64 gnd 0.007281f
C1524 vdd.n65 gnd 0.017213f
C1525 vdd.n66 gnd 0.003171f
C1526 vdd.n67 gnd 0.00308f
C1527 vdd.n68 gnd 0.014816f
C1528 vdd.n69 gnd 0.010344f
C1529 vdd.t158 gnd 0.036239f
C1530 vdd.t98 gnd 0.036239f
C1531 vdd.n70 gnd 0.249058f
C1532 vdd.n71 gnd 0.195846f
C1533 vdd.t171 gnd 0.036239f
C1534 vdd.t59 gnd 0.036239f
C1535 vdd.n72 gnd 0.249058f
C1536 vdd.n73 gnd 0.158047f
C1537 vdd.t146 gnd 0.036239f
C1538 vdd.t88 gnd 0.036239f
C1539 vdd.n74 gnd 0.249058f
C1540 vdd.n75 gnd 0.158047f
C1541 vdd.t167 gnd 0.036239f
C1542 vdd.t140 gnd 0.036239f
C1543 vdd.n76 gnd 0.249058f
C1544 vdd.n77 gnd 0.158047f
C1545 vdd.t30 gnd 0.036239f
C1546 vdd.t77 gnd 0.036239f
C1547 vdd.n78 gnd 0.249058f
C1548 vdd.n79 gnd 0.158047f
C1549 vdd.t42 gnd 0.036239f
C1550 vdd.t101 gnd 0.036239f
C1551 vdd.n80 gnd 0.249058f
C1552 vdd.n81 gnd 0.158047f
C1553 vdd.t72 gnd 0.036239f
C1554 vdd.t154 gnd 0.036239f
C1555 vdd.n82 gnd 0.249058f
C1556 vdd.n83 gnd 0.158047f
C1557 vdd.t46 gnd 0.036239f
C1558 vdd.t126 gnd 0.036239f
C1559 vdd.n84 gnd 0.249058f
C1560 vdd.n85 gnd 0.158047f
C1561 vdd.t54 gnd 0.036239f
C1562 vdd.t141 gnd 0.036239f
C1563 vdd.n86 gnd 0.249058f
C1564 vdd.n87 gnd 0.158047f
C1565 vdd.n88 gnd 0.006177f
C1566 vdd.n89 gnd 0.005732f
C1567 vdd.n90 gnd 0.003171f
C1568 vdd.n91 gnd 0.007281f
C1569 vdd.n92 gnd 0.00308f
C1570 vdd.n93 gnd 0.003262f
C1571 vdd.n94 gnd 0.005732f
C1572 vdd.n95 gnd 0.00308f
C1573 vdd.n96 gnd 0.007281f
C1574 vdd.n97 gnd 0.003262f
C1575 vdd.n98 gnd 0.005732f
C1576 vdd.n99 gnd 0.00308f
C1577 vdd.n100 gnd 0.005461f
C1578 vdd.n101 gnd 0.005477f
C1579 vdd.t83 gnd 0.015642f
C1580 vdd.n102 gnd 0.034803f
C1581 vdd.n103 gnd 0.181124f
C1582 vdd.n104 gnd 0.00308f
C1583 vdd.n105 gnd 0.003262f
C1584 vdd.n106 gnd 0.007281f
C1585 vdd.n107 gnd 0.007281f
C1586 vdd.n108 gnd 0.003262f
C1587 vdd.n109 gnd 0.00308f
C1588 vdd.n110 gnd 0.005732f
C1589 vdd.n111 gnd 0.005732f
C1590 vdd.n112 gnd 0.00308f
C1591 vdd.n113 gnd 0.003262f
C1592 vdd.n114 gnd 0.007281f
C1593 vdd.n115 gnd 0.007281f
C1594 vdd.n116 gnd 0.003262f
C1595 vdd.n117 gnd 0.00308f
C1596 vdd.n118 gnd 0.005732f
C1597 vdd.n119 gnd 0.005732f
C1598 vdd.n120 gnd 0.00308f
C1599 vdd.n121 gnd 0.003262f
C1600 vdd.n122 gnd 0.007281f
C1601 vdd.n123 gnd 0.007281f
C1602 vdd.n124 gnd 0.017213f
C1603 vdd.n125 gnd 0.003171f
C1604 vdd.n126 gnd 0.00308f
C1605 vdd.n127 gnd 0.014816f
C1606 vdd.n128 gnd 0.010019f
C1607 vdd.n129 gnd 0.117588f
C1608 vdd.n130 gnd 0.006177f
C1609 vdd.n131 gnd 0.005732f
C1610 vdd.n132 gnd 0.003171f
C1611 vdd.n133 gnd 0.007281f
C1612 vdd.n134 gnd 0.00308f
C1613 vdd.n135 gnd 0.003262f
C1614 vdd.n136 gnd 0.005732f
C1615 vdd.n137 gnd 0.00308f
C1616 vdd.n138 gnd 0.007281f
C1617 vdd.n139 gnd 0.003262f
C1618 vdd.n140 gnd 0.005732f
C1619 vdd.n141 gnd 0.00308f
C1620 vdd.n142 gnd 0.005461f
C1621 vdd.n143 gnd 0.005477f
C1622 vdd.t104 gnd 0.015642f
C1623 vdd.n144 gnd 0.034803f
C1624 vdd.n145 gnd 0.181124f
C1625 vdd.n146 gnd 0.00308f
C1626 vdd.n147 gnd 0.003262f
C1627 vdd.n148 gnd 0.007281f
C1628 vdd.n149 gnd 0.007281f
C1629 vdd.n150 gnd 0.003262f
C1630 vdd.n151 gnd 0.00308f
C1631 vdd.n152 gnd 0.005732f
C1632 vdd.n153 gnd 0.005732f
C1633 vdd.n154 gnd 0.00308f
C1634 vdd.n155 gnd 0.003262f
C1635 vdd.n156 gnd 0.007281f
C1636 vdd.n157 gnd 0.007281f
C1637 vdd.n158 gnd 0.003262f
C1638 vdd.n159 gnd 0.00308f
C1639 vdd.n160 gnd 0.005732f
C1640 vdd.n161 gnd 0.005732f
C1641 vdd.n162 gnd 0.00308f
C1642 vdd.n163 gnd 0.003262f
C1643 vdd.n164 gnd 0.007281f
C1644 vdd.n165 gnd 0.007281f
C1645 vdd.n166 gnd 0.017213f
C1646 vdd.n167 gnd 0.003171f
C1647 vdd.n168 gnd 0.00308f
C1648 vdd.n169 gnd 0.014816f
C1649 vdd.n170 gnd 0.010344f
C1650 vdd.t106 gnd 0.036239f
C1651 vdd.t136 gnd 0.036239f
C1652 vdd.n171 gnd 0.249058f
C1653 vdd.n172 gnd 0.195846f
C1654 vdd.t28 gnd 0.036239f
C1655 vdd.t96 gnd 0.036239f
C1656 vdd.n173 gnd 0.249058f
C1657 vdd.n174 gnd 0.158047f
C1658 vdd.t133 gnd 0.036239f
C1659 vdd.t15 gnd 0.036239f
C1660 vdd.n175 gnd 0.249058f
C1661 vdd.n176 gnd 0.158047f
C1662 vdd.t74 gnd 0.036239f
C1663 vdd.t76 gnd 0.036239f
C1664 vdd.n177 gnd 0.249058f
C1665 vdd.n178 gnd 0.158047f
C1666 vdd.t162 gnd 0.036239f
C1667 vdd.t69 gnd 0.036239f
C1668 vdd.n179 gnd 0.249058f
C1669 vdd.n180 gnd 0.158047f
C1670 vdd.t70 gnd 0.036239f
C1671 vdd.t156 gnd 0.036239f
C1672 vdd.n181 gnd 0.249058f
C1673 vdd.n182 gnd 0.158047f
C1674 vdd.t157 gnd 0.036239f
C1675 vdd.t40 gnd 0.036239f
C1676 vdd.n183 gnd 0.249058f
C1677 vdd.n184 gnd 0.158047f
C1678 vdd.t135 gnd 0.036239f
C1679 vdd.t153 gnd 0.036239f
C1680 vdd.n185 gnd 0.249058f
C1681 vdd.n186 gnd 0.158047f
C1682 vdd.t38 gnd 0.036239f
C1683 vdd.t95 gnd 0.036239f
C1684 vdd.n187 gnd 0.249058f
C1685 vdd.n188 gnd 0.158047f
C1686 vdd.n189 gnd 0.006177f
C1687 vdd.n190 gnd 0.005732f
C1688 vdd.n191 gnd 0.003171f
C1689 vdd.n192 gnd 0.007281f
C1690 vdd.n193 gnd 0.00308f
C1691 vdd.n194 gnd 0.003262f
C1692 vdd.n195 gnd 0.005732f
C1693 vdd.n196 gnd 0.00308f
C1694 vdd.n197 gnd 0.007281f
C1695 vdd.n198 gnd 0.003262f
C1696 vdd.n199 gnd 0.005732f
C1697 vdd.n200 gnd 0.00308f
C1698 vdd.n201 gnd 0.005461f
C1699 vdd.n202 gnd 0.005477f
C1700 vdd.t134 gnd 0.015642f
C1701 vdd.n203 gnd 0.034803f
C1702 vdd.n204 gnd 0.181124f
C1703 vdd.n205 gnd 0.00308f
C1704 vdd.n206 gnd 0.003262f
C1705 vdd.n207 gnd 0.007281f
C1706 vdd.n208 gnd 0.007281f
C1707 vdd.n209 gnd 0.003262f
C1708 vdd.n210 gnd 0.00308f
C1709 vdd.n211 gnd 0.005732f
C1710 vdd.n212 gnd 0.005732f
C1711 vdd.n213 gnd 0.00308f
C1712 vdd.n214 gnd 0.003262f
C1713 vdd.n215 gnd 0.007281f
C1714 vdd.n216 gnd 0.007281f
C1715 vdd.n217 gnd 0.003262f
C1716 vdd.n218 gnd 0.00308f
C1717 vdd.n219 gnd 0.005732f
C1718 vdd.n220 gnd 0.005732f
C1719 vdd.n221 gnd 0.00308f
C1720 vdd.n222 gnd 0.003262f
C1721 vdd.n223 gnd 0.007281f
C1722 vdd.n224 gnd 0.007281f
C1723 vdd.n225 gnd 0.017213f
C1724 vdd.n226 gnd 0.003171f
C1725 vdd.n227 gnd 0.00308f
C1726 vdd.n228 gnd 0.014816f
C1727 vdd.n229 gnd 0.010019f
C1728 vdd.n230 gnd 0.069953f
C1729 vdd.n231 gnd 0.252058f
C1730 vdd.n232 gnd 0.006177f
C1731 vdd.n233 gnd 0.005732f
C1732 vdd.n234 gnd 0.003171f
C1733 vdd.n235 gnd 0.007281f
C1734 vdd.n236 gnd 0.00308f
C1735 vdd.n237 gnd 0.003262f
C1736 vdd.n238 gnd 0.005732f
C1737 vdd.n239 gnd 0.00308f
C1738 vdd.n240 gnd 0.007281f
C1739 vdd.n241 gnd 0.003262f
C1740 vdd.n242 gnd 0.005732f
C1741 vdd.n243 gnd 0.00308f
C1742 vdd.n244 gnd 0.005461f
C1743 vdd.n245 gnd 0.005477f
C1744 vdd.t119 gnd 0.015642f
C1745 vdd.n246 gnd 0.034803f
C1746 vdd.n247 gnd 0.181124f
C1747 vdd.n248 gnd 0.00308f
C1748 vdd.n249 gnd 0.003262f
C1749 vdd.n250 gnd 0.007281f
C1750 vdd.n251 gnd 0.007281f
C1751 vdd.n252 gnd 0.003262f
C1752 vdd.n253 gnd 0.00308f
C1753 vdd.n254 gnd 0.005732f
C1754 vdd.n255 gnd 0.005732f
C1755 vdd.n256 gnd 0.00308f
C1756 vdd.n257 gnd 0.003262f
C1757 vdd.n258 gnd 0.007281f
C1758 vdd.n259 gnd 0.007281f
C1759 vdd.n260 gnd 0.003262f
C1760 vdd.n261 gnd 0.00308f
C1761 vdd.n262 gnd 0.005732f
C1762 vdd.n263 gnd 0.005732f
C1763 vdd.n264 gnd 0.00308f
C1764 vdd.n265 gnd 0.003262f
C1765 vdd.n266 gnd 0.007281f
C1766 vdd.n267 gnd 0.007281f
C1767 vdd.n268 gnd 0.017213f
C1768 vdd.n269 gnd 0.003171f
C1769 vdd.n270 gnd 0.00308f
C1770 vdd.n271 gnd 0.014816f
C1771 vdd.n272 gnd 0.010344f
C1772 vdd.t121 gnd 0.036239f
C1773 vdd.t150 gnd 0.036239f
C1774 vdd.n273 gnd 0.249058f
C1775 vdd.n274 gnd 0.195846f
C1776 vdd.t51 gnd 0.036239f
C1777 vdd.t116 gnd 0.036239f
C1778 vdd.n275 gnd 0.249058f
C1779 vdd.n276 gnd 0.158047f
C1780 vdd.t143 gnd 0.036239f
C1781 vdd.t16 gnd 0.036239f
C1782 vdd.n277 gnd 0.249058f
C1783 vdd.n278 gnd 0.158047f
C1784 vdd.t91 gnd 0.036239f
C1785 vdd.t93 gnd 0.036239f
C1786 vdd.n279 gnd 0.249058f
C1787 vdd.n280 gnd 0.158047f
C1788 vdd.t170 gnd 0.036239f
C1789 vdd.t86 gnd 0.036239f
C1790 vdd.n281 gnd 0.249058f
C1791 vdd.n282 gnd 0.158047f
C1792 vdd.t87 gnd 0.036239f
C1793 vdd.t160 gnd 0.036239f
C1794 vdd.n283 gnd 0.249058f
C1795 vdd.n284 gnd 0.158047f
C1796 vdd.t169 gnd 0.036239f
C1797 vdd.t64 gnd 0.036239f
C1798 vdd.n285 gnd 0.249058f
C1799 vdd.n286 gnd 0.158047f
C1800 vdd.t148 gnd 0.036239f
C1801 vdd.t166 gnd 0.036239f
C1802 vdd.n287 gnd 0.249058f
C1803 vdd.n288 gnd 0.158047f
C1804 vdd.t55 gnd 0.036239f
C1805 vdd.t117 gnd 0.036239f
C1806 vdd.n289 gnd 0.249058f
C1807 vdd.n290 gnd 0.158047f
C1808 vdd.n291 gnd 0.006177f
C1809 vdd.n292 gnd 0.005732f
C1810 vdd.n293 gnd 0.003171f
C1811 vdd.n294 gnd 0.007281f
C1812 vdd.n295 gnd 0.00308f
C1813 vdd.n296 gnd 0.003262f
C1814 vdd.n297 gnd 0.005732f
C1815 vdd.n298 gnd 0.00308f
C1816 vdd.n299 gnd 0.007281f
C1817 vdd.n300 gnd 0.003262f
C1818 vdd.n301 gnd 0.005732f
C1819 vdd.n302 gnd 0.00308f
C1820 vdd.n303 gnd 0.005461f
C1821 vdd.n304 gnd 0.005477f
C1822 vdd.t144 gnd 0.015642f
C1823 vdd.n305 gnd 0.034803f
C1824 vdd.n306 gnd 0.181124f
C1825 vdd.n307 gnd 0.00308f
C1826 vdd.n308 gnd 0.003262f
C1827 vdd.n309 gnd 0.007281f
C1828 vdd.n310 gnd 0.007281f
C1829 vdd.n311 gnd 0.003262f
C1830 vdd.n312 gnd 0.00308f
C1831 vdd.n313 gnd 0.005732f
C1832 vdd.n314 gnd 0.005732f
C1833 vdd.n315 gnd 0.00308f
C1834 vdd.n316 gnd 0.003262f
C1835 vdd.n317 gnd 0.007281f
C1836 vdd.n318 gnd 0.007281f
C1837 vdd.n319 gnd 0.003262f
C1838 vdd.n320 gnd 0.00308f
C1839 vdd.n321 gnd 0.005732f
C1840 vdd.n322 gnd 0.005732f
C1841 vdd.n323 gnd 0.00308f
C1842 vdd.n324 gnd 0.003262f
C1843 vdd.n325 gnd 0.007281f
C1844 vdd.n326 gnd 0.007281f
C1845 vdd.n327 gnd 0.017213f
C1846 vdd.n328 gnd 0.003171f
C1847 vdd.n329 gnd 0.00308f
C1848 vdd.n330 gnd 0.014816f
C1849 vdd.n331 gnd 0.010019f
C1850 vdd.n332 gnd 0.069953f
C1851 vdd.n333 gnd 0.288552f
C1852 vdd.n334 gnd 0.008651f
C1853 vdd.n335 gnd 0.011256f
C1854 vdd.n336 gnd 0.00906f
C1855 vdd.n337 gnd 0.00906f
C1856 vdd.n338 gnd 0.011256f
C1857 vdd.n339 gnd 0.011256f
C1858 vdd.n340 gnd 0.822471f
C1859 vdd.n341 gnd 0.011256f
C1860 vdd.n342 gnd 0.011256f
C1861 vdd.n343 gnd 0.011256f
C1862 vdd.n344 gnd 0.89149f
C1863 vdd.n345 gnd 0.011256f
C1864 vdd.n346 gnd 0.011256f
C1865 vdd.n347 gnd 0.011256f
C1866 vdd.n348 gnd 0.011256f
C1867 vdd.n349 gnd 0.00906f
C1868 vdd.n350 gnd 0.011256f
C1869 vdd.t100 gnd 0.575155f
C1870 vdd.n351 gnd 0.011256f
C1871 vdd.n352 gnd 0.011256f
C1872 vdd.n353 gnd 0.011256f
C1873 vdd.t39 gnd 0.575155f
C1874 vdd.n354 gnd 0.011256f
C1875 vdd.n355 gnd 0.011256f
C1876 vdd.n356 gnd 0.011256f
C1877 vdd.n357 gnd 0.011256f
C1878 vdd.n358 gnd 0.011256f
C1879 vdd.n359 gnd 0.00906f
C1880 vdd.n360 gnd 0.011256f
C1881 vdd.n361 gnd 0.649925f
C1882 vdd.n362 gnd 0.011256f
C1883 vdd.n363 gnd 0.011256f
C1884 vdd.n364 gnd 0.011256f
C1885 vdd.t125 gnd 0.575155f
C1886 vdd.n365 gnd 0.011256f
C1887 vdd.n366 gnd 0.011256f
C1888 vdd.n367 gnd 0.011256f
C1889 vdd.n368 gnd 0.011256f
C1890 vdd.n369 gnd 0.011256f
C1891 vdd.n370 gnd 0.00906f
C1892 vdd.n371 gnd 0.011256f
C1893 vdd.t37 gnd 0.575155f
C1894 vdd.n372 gnd 0.011256f
C1895 vdd.n373 gnd 0.011256f
C1896 vdd.n374 gnd 0.011256f
C1897 vdd.n375 gnd 0.672931f
C1898 vdd.n376 gnd 0.011256f
C1899 vdd.n377 gnd 0.011256f
C1900 vdd.n378 gnd 0.011256f
C1901 vdd.n379 gnd 0.011256f
C1902 vdd.n380 gnd 0.011256f
C1903 vdd.n381 gnd 0.00906f
C1904 vdd.n382 gnd 0.011256f
C1905 vdd.t82 gnd 0.575155f
C1906 vdd.n383 gnd 0.011256f
C1907 vdd.n384 gnd 0.011256f
C1908 vdd.n385 gnd 0.011256f
C1909 vdd.n386 gnd 0.580906f
C1910 vdd.n387 gnd 0.011256f
C1911 vdd.n388 gnd 0.011256f
C1912 vdd.n389 gnd 0.011256f
C1913 vdd.n390 gnd 0.011256f
C1914 vdd.n391 gnd 0.027229f
C1915 vdd.n392 gnd 0.027813f
C1916 vdd.t238 gnd 0.575155f
C1917 vdd.n393 gnd 0.027229f
C1918 vdd.n425 gnd 0.011256f
C1919 vdd.t240 gnd 0.138478f
C1920 vdd.t239 gnd 0.147995f
C1921 vdd.t237 gnd 0.180851f
C1922 vdd.n426 gnd 0.231825f
C1923 vdd.n427 gnd 0.195681f
C1924 vdd.n428 gnd 0.014858f
C1925 vdd.n429 gnd 0.011256f
C1926 vdd.n430 gnd 0.00906f
C1927 vdd.n431 gnd 0.011256f
C1928 vdd.n432 gnd 0.00906f
C1929 vdd.n433 gnd 0.011256f
C1930 vdd.n434 gnd 0.00906f
C1931 vdd.n435 gnd 0.011256f
C1932 vdd.n436 gnd 0.00906f
C1933 vdd.n437 gnd 0.011256f
C1934 vdd.n438 gnd 0.00906f
C1935 vdd.n439 gnd 0.011256f
C1936 vdd.t280 gnd 0.138478f
C1937 vdd.t279 gnd 0.147995f
C1938 vdd.t278 gnd 0.180851f
C1939 vdd.n440 gnd 0.231825f
C1940 vdd.n441 gnd 0.195681f
C1941 vdd.n442 gnd 0.00906f
C1942 vdd.n443 gnd 0.011256f
C1943 vdd.n444 gnd 0.00906f
C1944 vdd.n445 gnd 0.011256f
C1945 vdd.n446 gnd 0.00906f
C1946 vdd.n447 gnd 0.011256f
C1947 vdd.n448 gnd 0.00906f
C1948 vdd.n449 gnd 0.011256f
C1949 vdd.n450 gnd 0.00906f
C1950 vdd.n451 gnd 0.011256f
C1951 vdd.t286 gnd 0.138478f
C1952 vdd.t285 gnd 0.147995f
C1953 vdd.t284 gnd 0.180851f
C1954 vdd.n452 gnd 0.231825f
C1955 vdd.n453 gnd 0.195681f
C1956 vdd.n454 gnd 0.019388f
C1957 vdd.n455 gnd 0.011256f
C1958 vdd.n456 gnd 0.00906f
C1959 vdd.n457 gnd 0.011256f
C1960 vdd.n458 gnd 0.00906f
C1961 vdd.n459 gnd 0.011256f
C1962 vdd.n460 gnd 0.00906f
C1963 vdd.n461 gnd 0.011256f
C1964 vdd.n462 gnd 0.00906f
C1965 vdd.n463 gnd 0.011256f
C1966 vdd.n464 gnd 0.027813f
C1967 vdd.n465 gnd 0.00752f
C1968 vdd.n466 gnd 0.00906f
C1969 vdd.n467 gnd 0.011256f
C1970 vdd.n468 gnd 0.011256f
C1971 vdd.n469 gnd 0.00906f
C1972 vdd.n470 gnd 0.011256f
C1973 vdd.n471 gnd 0.011256f
C1974 vdd.n472 gnd 0.011256f
C1975 vdd.n473 gnd 0.011256f
C1976 vdd.n474 gnd 0.011256f
C1977 vdd.n475 gnd 0.00906f
C1978 vdd.n476 gnd 0.00906f
C1979 vdd.n477 gnd 0.011256f
C1980 vdd.n478 gnd 0.011256f
C1981 vdd.n479 gnd 0.00906f
C1982 vdd.n480 gnd 0.011256f
C1983 vdd.n481 gnd 0.011256f
C1984 vdd.n482 gnd 0.011256f
C1985 vdd.n483 gnd 0.011256f
C1986 vdd.n484 gnd 0.011256f
C1987 vdd.n485 gnd 0.00906f
C1988 vdd.n486 gnd 0.00906f
C1989 vdd.n487 gnd 0.011256f
C1990 vdd.n488 gnd 0.011256f
C1991 vdd.n489 gnd 0.00906f
C1992 vdd.n490 gnd 0.011256f
C1993 vdd.n491 gnd 0.011256f
C1994 vdd.n492 gnd 0.011256f
C1995 vdd.n493 gnd 0.011256f
C1996 vdd.n494 gnd 0.011256f
C1997 vdd.n495 gnd 0.00906f
C1998 vdd.n496 gnd 0.00906f
C1999 vdd.n497 gnd 0.011256f
C2000 vdd.n498 gnd 0.011256f
C2001 vdd.n499 gnd 0.00906f
C2002 vdd.n500 gnd 0.011256f
C2003 vdd.n501 gnd 0.011256f
C2004 vdd.n502 gnd 0.011256f
C2005 vdd.n503 gnd 0.011256f
C2006 vdd.n504 gnd 0.011256f
C2007 vdd.n505 gnd 0.00906f
C2008 vdd.n506 gnd 0.00906f
C2009 vdd.n507 gnd 0.011256f
C2010 vdd.n508 gnd 0.011256f
C2011 vdd.n509 gnd 0.007565f
C2012 vdd.n510 gnd 0.011256f
C2013 vdd.n511 gnd 0.011256f
C2014 vdd.n512 gnd 0.011256f
C2015 vdd.n513 gnd 0.011256f
C2016 vdd.n514 gnd 0.011256f
C2017 vdd.n515 gnd 0.007565f
C2018 vdd.n516 gnd 0.00906f
C2019 vdd.n517 gnd 0.011256f
C2020 vdd.n518 gnd 0.011256f
C2021 vdd.n519 gnd 0.00906f
C2022 vdd.n520 gnd 0.011256f
C2023 vdd.n521 gnd 0.011256f
C2024 vdd.n522 gnd 0.011256f
C2025 vdd.n523 gnd 0.011256f
C2026 vdd.n524 gnd 0.011256f
C2027 vdd.n525 gnd 0.00906f
C2028 vdd.n526 gnd 0.00906f
C2029 vdd.n527 gnd 0.011256f
C2030 vdd.n528 gnd 0.011256f
C2031 vdd.n529 gnd 0.00906f
C2032 vdd.n530 gnd 0.011256f
C2033 vdd.n531 gnd 0.011256f
C2034 vdd.n532 gnd 0.011256f
C2035 vdd.n533 gnd 0.011256f
C2036 vdd.n534 gnd 0.011256f
C2037 vdd.n535 gnd 0.00906f
C2038 vdd.n536 gnd 0.00906f
C2039 vdd.n537 gnd 0.011256f
C2040 vdd.n538 gnd 0.011256f
C2041 vdd.n539 gnd 0.00906f
C2042 vdd.n540 gnd 0.011256f
C2043 vdd.n541 gnd 0.011256f
C2044 vdd.n542 gnd 0.011256f
C2045 vdd.n543 gnd 0.011256f
C2046 vdd.n544 gnd 0.011256f
C2047 vdd.n545 gnd 0.00906f
C2048 vdd.n546 gnd 0.00906f
C2049 vdd.n547 gnd 0.011256f
C2050 vdd.n548 gnd 0.011256f
C2051 vdd.n549 gnd 0.00906f
C2052 vdd.n550 gnd 0.011256f
C2053 vdd.n551 gnd 0.011256f
C2054 vdd.n552 gnd 0.011256f
C2055 vdd.n553 gnd 0.011256f
C2056 vdd.n554 gnd 0.011256f
C2057 vdd.n555 gnd 0.00906f
C2058 vdd.n556 gnd 0.00906f
C2059 vdd.n557 gnd 0.011256f
C2060 vdd.n558 gnd 0.011256f
C2061 vdd.n559 gnd 0.00906f
C2062 vdd.n560 gnd 0.011256f
C2063 vdd.n561 gnd 0.011256f
C2064 vdd.n562 gnd 0.011256f
C2065 vdd.n563 gnd 0.011256f
C2066 vdd.n564 gnd 0.011256f
C2067 vdd.n565 gnd 0.006161f
C2068 vdd.n566 gnd 0.019388f
C2069 vdd.n567 gnd 0.011256f
C2070 vdd.n568 gnd 0.011256f
C2071 vdd.n569 gnd 0.008969f
C2072 vdd.n570 gnd 0.011256f
C2073 vdd.n571 gnd 0.011256f
C2074 vdd.n572 gnd 0.011256f
C2075 vdd.n573 gnd 0.011256f
C2076 vdd.n574 gnd 0.011256f
C2077 vdd.n575 gnd 0.00906f
C2078 vdd.n576 gnd 0.00906f
C2079 vdd.n577 gnd 0.011256f
C2080 vdd.n578 gnd 0.011256f
C2081 vdd.n579 gnd 0.00906f
C2082 vdd.n580 gnd 0.011256f
C2083 vdd.n581 gnd 0.011256f
C2084 vdd.n582 gnd 0.011256f
C2085 vdd.n583 gnd 0.011256f
C2086 vdd.n584 gnd 0.011256f
C2087 vdd.n585 gnd 0.00906f
C2088 vdd.n586 gnd 0.00906f
C2089 vdd.n587 gnd 0.011256f
C2090 vdd.n588 gnd 0.011256f
C2091 vdd.n589 gnd 0.00906f
C2092 vdd.n590 gnd 0.011256f
C2093 vdd.n591 gnd 0.011256f
C2094 vdd.n592 gnd 0.011256f
C2095 vdd.n593 gnd 0.011256f
C2096 vdd.n594 gnd 0.011256f
C2097 vdd.n595 gnd 0.00906f
C2098 vdd.n596 gnd 0.00906f
C2099 vdd.n597 gnd 0.011256f
C2100 vdd.n598 gnd 0.011256f
C2101 vdd.n599 gnd 0.00906f
C2102 vdd.n600 gnd 0.011256f
C2103 vdd.n601 gnd 0.011256f
C2104 vdd.n602 gnd 0.011256f
C2105 vdd.n603 gnd 0.011256f
C2106 vdd.n604 gnd 0.011256f
C2107 vdd.n605 gnd 0.00906f
C2108 vdd.n606 gnd 0.00906f
C2109 vdd.n607 gnd 0.011256f
C2110 vdd.n608 gnd 0.011256f
C2111 vdd.n609 gnd 0.00906f
C2112 vdd.n610 gnd 0.011256f
C2113 vdd.n611 gnd 0.011256f
C2114 vdd.n612 gnd 0.011256f
C2115 vdd.n613 gnd 0.011256f
C2116 vdd.n614 gnd 0.011256f
C2117 vdd.n615 gnd 0.00906f
C2118 vdd.n616 gnd 0.011256f
C2119 vdd.n617 gnd 0.00906f
C2120 vdd.n618 gnd 0.004756f
C2121 vdd.n619 gnd 0.011256f
C2122 vdd.n620 gnd 0.011256f
C2123 vdd.n621 gnd 0.00906f
C2124 vdd.n622 gnd 0.011256f
C2125 vdd.n623 gnd 0.00906f
C2126 vdd.n624 gnd 0.011256f
C2127 vdd.n625 gnd 0.00906f
C2128 vdd.n626 gnd 0.011256f
C2129 vdd.n627 gnd 0.00906f
C2130 vdd.n628 gnd 0.011256f
C2131 vdd.n629 gnd 0.00906f
C2132 vdd.n630 gnd 0.011256f
C2133 vdd.n631 gnd 0.00906f
C2134 vdd.n632 gnd 0.011256f
C2135 vdd.n633 gnd 0.626919f
C2136 vdd.t29 gnd 0.575155f
C2137 vdd.n634 gnd 0.011256f
C2138 vdd.n635 gnd 0.00906f
C2139 vdd.n636 gnd 0.011256f
C2140 vdd.n637 gnd 0.00906f
C2141 vdd.n638 gnd 0.011256f
C2142 vdd.t73 gnd 0.575155f
C2143 vdd.n639 gnd 0.011256f
C2144 vdd.n640 gnd 0.00906f
C2145 vdd.n641 gnd 0.011256f
C2146 vdd.n642 gnd 0.00906f
C2147 vdd.n643 gnd 0.011256f
C2148 vdd.t14 gnd 0.575155f
C2149 vdd.n644 gnd 0.718943f
C2150 vdd.n645 gnd 0.011256f
C2151 vdd.n646 gnd 0.00906f
C2152 vdd.n647 gnd 0.011256f
C2153 vdd.n648 gnd 0.00906f
C2154 vdd.n649 gnd 0.011256f
C2155 vdd.t132 gnd 0.575155f
C2156 vdd.n650 gnd 0.011256f
C2157 vdd.n651 gnd 0.00906f
C2158 vdd.n652 gnd 0.011256f
C2159 vdd.n653 gnd 0.00906f
C2160 vdd.n654 gnd 0.011256f
C2161 vdd.n655 gnd 0.799465f
C2162 vdd.n656 gnd 0.954757f
C2163 vdd.t58 gnd 0.575155f
C2164 vdd.n657 gnd 0.011256f
C2165 vdd.n658 gnd 0.00906f
C2166 vdd.n659 gnd 0.011256f
C2167 vdd.n660 gnd 0.00906f
C2168 vdd.n661 gnd 0.011256f
C2169 vdd.n662 gnd 0.603912f
C2170 vdd.n663 gnd 0.011256f
C2171 vdd.n664 gnd 0.00906f
C2172 vdd.n665 gnd 0.011256f
C2173 vdd.n666 gnd 0.00906f
C2174 vdd.n667 gnd 0.011256f
C2175 vdd.t105 gnd 0.575155f
C2176 vdd.t97 gnd 0.575155f
C2177 vdd.n668 gnd 0.011256f
C2178 vdd.n669 gnd 0.00906f
C2179 vdd.n670 gnd 0.011256f
C2180 vdd.n671 gnd 0.00906f
C2181 vdd.n672 gnd 0.011256f
C2182 vdd.t17 gnd 0.575155f
C2183 vdd.n673 gnd 0.011256f
C2184 vdd.n674 gnd 0.00906f
C2185 vdd.n675 gnd 0.011256f
C2186 vdd.n676 gnd 0.00906f
C2187 vdd.n677 gnd 0.011256f
C2188 vdd.n678 gnd 1.15031f
C2189 vdd.n679 gnd 0.937502f
C2190 vdd.n680 gnd 0.011256f
C2191 vdd.n681 gnd 0.00906f
C2192 vdd.n682 gnd 0.027229f
C2193 vdd.n683 gnd 0.00752f
C2194 vdd.n684 gnd 0.027229f
C2195 vdd.t216 gnd 0.575155f
C2196 vdd.n685 gnd 0.027229f
C2197 vdd.n686 gnd 0.00752f
C2198 vdd.n687 gnd 0.00968f
C2199 vdd.t282 gnd 0.138478f
C2200 vdd.t283 gnd 0.147995f
C2201 vdd.t281 gnd 0.180851f
C2202 vdd.n688 gnd 0.231825f
C2203 vdd.n689 gnd 0.194775f
C2204 vdd.n690 gnd 0.013952f
C2205 vdd.n691 gnd 0.011256f
C2206 vdd.n692 gnd 7.92563f
C2207 vdd.n723 gnd 1.58168f
C2208 vdd.n724 gnd 0.011256f
C2209 vdd.n725 gnd 0.011256f
C2210 vdd.n726 gnd 0.027813f
C2211 vdd.n727 gnd 0.00968f
C2212 vdd.n728 gnd 0.011256f
C2213 vdd.n729 gnd 0.00906f
C2214 vdd.n730 gnd 0.007204f
C2215 vdd.n731 gnd 0.018393f
C2216 vdd.n732 gnd 0.00906f
C2217 vdd.n733 gnd 0.011256f
C2218 vdd.n734 gnd 0.011256f
C2219 vdd.n735 gnd 0.011256f
C2220 vdd.n736 gnd 0.011256f
C2221 vdd.n737 gnd 0.011256f
C2222 vdd.n738 gnd 0.011256f
C2223 vdd.n739 gnd 0.011256f
C2224 vdd.n740 gnd 0.011256f
C2225 vdd.n741 gnd 0.011256f
C2226 vdd.n742 gnd 0.011256f
C2227 vdd.n743 gnd 0.011256f
C2228 vdd.n744 gnd 0.011256f
C2229 vdd.n745 gnd 0.011256f
C2230 vdd.n746 gnd 0.011256f
C2231 vdd.n747 gnd 0.007565f
C2232 vdd.n748 gnd 0.011256f
C2233 vdd.n749 gnd 0.011256f
C2234 vdd.n750 gnd 0.011256f
C2235 vdd.n751 gnd 0.011256f
C2236 vdd.n752 gnd 0.011256f
C2237 vdd.n753 gnd 0.011256f
C2238 vdd.n754 gnd 0.011256f
C2239 vdd.n755 gnd 0.011256f
C2240 vdd.n756 gnd 0.011256f
C2241 vdd.n757 gnd 0.011256f
C2242 vdd.n758 gnd 0.011256f
C2243 vdd.n759 gnd 0.011256f
C2244 vdd.n760 gnd 0.011256f
C2245 vdd.n761 gnd 0.011256f
C2246 vdd.n762 gnd 0.011256f
C2247 vdd.n763 gnd 0.011256f
C2248 vdd.n764 gnd 0.011256f
C2249 vdd.n765 gnd 0.011256f
C2250 vdd.n766 gnd 0.011256f
C2251 vdd.n767 gnd 0.008969f
C2252 vdd.t217 gnd 0.138478f
C2253 vdd.t218 gnd 0.147995f
C2254 vdd.t215 gnd 0.180851f
C2255 vdd.n768 gnd 0.231825f
C2256 vdd.n769 gnd 0.194775f
C2257 vdd.n770 gnd 0.011256f
C2258 vdd.n771 gnd 0.011256f
C2259 vdd.n772 gnd 0.011256f
C2260 vdd.n773 gnd 0.011256f
C2261 vdd.n774 gnd 0.011256f
C2262 vdd.n775 gnd 0.011256f
C2263 vdd.n776 gnd 0.011256f
C2264 vdd.n777 gnd 0.011256f
C2265 vdd.n778 gnd 0.011256f
C2266 vdd.n779 gnd 0.011256f
C2267 vdd.n780 gnd 0.011256f
C2268 vdd.n781 gnd 0.011256f
C2269 vdd.n782 gnd 0.011256f
C2270 vdd.n783 gnd 0.007204f
C2271 vdd.n785 gnd 0.007654f
C2272 vdd.n786 gnd 0.007654f
C2273 vdd.n787 gnd 0.007654f
C2274 vdd.n788 gnd 0.007654f
C2275 vdd.n789 gnd 0.007654f
C2276 vdd.n790 gnd 0.007654f
C2277 vdd.n792 gnd 0.007654f
C2278 vdd.n793 gnd 0.007654f
C2279 vdd.n795 gnd 0.007654f
C2280 vdd.n796 gnd 0.005572f
C2281 vdd.n798 gnd 0.007654f
C2282 vdd.t264 gnd 0.3093f
C2283 vdd.t263 gnd 0.316607f
C2284 vdd.t262 gnd 0.201923f
C2285 vdd.n799 gnd 0.109128f
C2286 vdd.n800 gnd 0.061901f
C2287 vdd.n801 gnd 0.010939f
C2288 vdd.n802 gnd 0.017889f
C2289 vdd.n804 gnd 0.007654f
C2290 vdd.n805 gnd 0.78221f
C2291 vdd.n806 gnd 0.016957f
C2292 vdd.n807 gnd 0.016957f
C2293 vdd.n808 gnd 0.007654f
C2294 vdd.n809 gnd 0.018162f
C2295 vdd.n810 gnd 0.007654f
C2296 vdd.n811 gnd 0.007654f
C2297 vdd.n812 gnd 0.007654f
C2298 vdd.n813 gnd 0.007654f
C2299 vdd.n814 gnd 0.007654f
C2300 vdd.n816 gnd 0.007654f
C2301 vdd.n817 gnd 0.007654f
C2302 vdd.n819 gnd 0.007654f
C2303 vdd.n820 gnd 0.007654f
C2304 vdd.n822 gnd 0.007654f
C2305 vdd.n823 gnd 0.007654f
C2306 vdd.n825 gnd 0.007654f
C2307 vdd.n826 gnd 0.007654f
C2308 vdd.n828 gnd 0.007654f
C2309 vdd.n829 gnd 0.007654f
C2310 vdd.n831 gnd 0.007654f
C2311 vdd.t257 gnd 0.3093f
C2312 vdd.t256 gnd 0.316607f
C2313 vdd.t254 gnd 0.201923f
C2314 vdd.n832 gnd 0.109128f
C2315 vdd.n833 gnd 0.061901f
C2316 vdd.n834 gnd 0.007654f
C2317 vdd.n836 gnd 0.007654f
C2318 vdd.n837 gnd 0.007654f
C2319 vdd.t255 gnd 0.391105f
C2320 vdd.n838 gnd 0.007654f
C2321 vdd.n839 gnd 0.007654f
C2322 vdd.n840 gnd 0.007654f
C2323 vdd.n841 gnd 0.007654f
C2324 vdd.n842 gnd 0.007654f
C2325 vdd.n843 gnd 0.78221f
C2326 vdd.n844 gnd 0.007654f
C2327 vdd.n845 gnd 0.007654f
C2328 vdd.n846 gnd 0.684434f
C2329 vdd.n847 gnd 0.007654f
C2330 vdd.n848 gnd 0.007654f
C2331 vdd.n849 gnd 0.006754f
C2332 vdd.n850 gnd 0.007654f
C2333 vdd.n851 gnd 0.690186f
C2334 vdd.n852 gnd 0.007654f
C2335 vdd.n853 gnd 0.007654f
C2336 vdd.n854 gnd 0.007654f
C2337 vdd.n855 gnd 0.007654f
C2338 vdd.n856 gnd 0.007654f
C2339 vdd.n857 gnd 0.78221f
C2340 vdd.n858 gnd 0.007654f
C2341 vdd.n859 gnd 0.007654f
C2342 vdd.t227 gnd 0.350844f
C2343 vdd.t178 gnd 0.092025f
C2344 vdd.n860 gnd 0.007654f
C2345 vdd.n861 gnd 0.007654f
C2346 vdd.n862 gnd 0.007654f
C2347 vdd.t192 gnd 0.391105f
C2348 vdd.n863 gnd 0.007654f
C2349 vdd.n864 gnd 0.007654f
C2350 vdd.n865 gnd 0.007654f
C2351 vdd.n866 gnd 0.007654f
C2352 vdd.n867 gnd 0.007654f
C2353 vdd.t11 gnd 0.391105f
C2354 vdd.n868 gnd 0.007654f
C2355 vdd.n869 gnd 0.007654f
C2356 vdd.n870 gnd 0.649925f
C2357 vdd.n871 gnd 0.007654f
C2358 vdd.n872 gnd 0.007654f
C2359 vdd.n873 gnd 0.007654f
C2360 vdd.n874 gnd 0.477378f
C2361 vdd.n875 gnd 0.007654f
C2362 vdd.n876 gnd 0.007654f
C2363 vdd.t190 gnd 0.391105f
C2364 vdd.n877 gnd 0.007654f
C2365 vdd.n878 gnd 0.007654f
C2366 vdd.n879 gnd 0.007654f
C2367 vdd.n880 gnd 0.649925f
C2368 vdd.n881 gnd 0.007654f
C2369 vdd.n882 gnd 0.007654f
C2370 vdd.t187 gnd 0.33359f
C2371 vdd.t185 gnd 0.304832f
C2372 vdd.n883 gnd 0.007654f
C2373 vdd.n884 gnd 0.007654f
C2374 vdd.n885 gnd 0.007654f
C2375 vdd.t12 gnd 0.391105f
C2376 vdd.n886 gnd 0.007654f
C2377 vdd.n887 gnd 0.007654f
C2378 vdd.t183 gnd 0.391105f
C2379 vdd.n888 gnd 0.007654f
C2380 vdd.n889 gnd 0.007654f
C2381 vdd.n890 gnd 0.007654f
C2382 vdd.t179 gnd 0.287577f
C2383 vdd.n891 gnd 0.007654f
C2384 vdd.n892 gnd 0.007654f
C2385 vdd.n893 gnd 0.667179f
C2386 vdd.n894 gnd 0.007654f
C2387 vdd.n895 gnd 0.007654f
C2388 vdd.n896 gnd 0.007654f
C2389 vdd.n897 gnd 0.78221f
C2390 vdd.n898 gnd 0.007654f
C2391 vdd.n899 gnd 0.007654f
C2392 vdd.t0 gnd 0.350844f
C2393 vdd.n900 gnd 0.494633f
C2394 vdd.n901 gnd 0.007654f
C2395 vdd.n902 gnd 0.007654f
C2396 vdd.n903 gnd 0.007654f
C2397 vdd.t176 gnd 0.391105f
C2398 vdd.n904 gnd 0.007654f
C2399 vdd.n905 gnd 0.007654f
C2400 vdd.n906 gnd 0.007654f
C2401 vdd.n907 gnd 0.007654f
C2402 vdd.n908 gnd 0.007654f
C2403 vdd.t200 gnd 0.78221f
C2404 vdd.n909 gnd 0.007654f
C2405 vdd.n910 gnd 0.007654f
C2406 vdd.t259 gnd 0.391105f
C2407 vdd.n911 gnd 0.007654f
C2408 vdd.n912 gnd 0.018162f
C2409 vdd.n913 gnd 0.018162f
C2410 vdd.t193 gnd 0.736198f
C2411 vdd.n914 gnd 0.016957f
C2412 vdd.n915 gnd 0.016957f
C2413 vdd.n916 gnd 0.018162f
C2414 vdd.n917 gnd 0.007654f
C2415 vdd.n918 gnd 0.007654f
C2416 vdd.t204 gnd 0.736198f
C2417 vdd.n936 gnd 0.018162f
C2418 vdd.n954 gnd 0.016957f
C2419 vdd.n955 gnd 0.007654f
C2420 vdd.n956 gnd 0.016957f
C2421 vdd.t277 gnd 0.3093f
C2422 vdd.t276 gnd 0.316607f
C2423 vdd.t275 gnd 0.201923f
C2424 vdd.n957 gnd 0.109128f
C2425 vdd.n958 gnd 0.061901f
C2426 vdd.n959 gnd 0.017889f
C2427 vdd.n960 gnd 0.007654f
C2428 vdd.t292 gnd 0.78221f
C2429 vdd.n961 gnd 0.016957f
C2430 vdd.n962 gnd 0.007654f
C2431 vdd.n963 gnd 0.018162f
C2432 vdd.n964 gnd 0.007654f
C2433 vdd.t253 gnd 0.3093f
C2434 vdd.t252 gnd 0.316607f
C2435 vdd.t250 gnd 0.201923f
C2436 vdd.n965 gnd 0.109128f
C2437 vdd.n966 gnd 0.061901f
C2438 vdd.n967 gnd 0.010939f
C2439 vdd.n968 gnd 0.007654f
C2440 vdd.n969 gnd 0.007654f
C2441 vdd.t251 gnd 0.391105f
C2442 vdd.n970 gnd 0.007654f
C2443 vdd.n971 gnd 0.007654f
C2444 vdd.n972 gnd 0.007654f
C2445 vdd.n973 gnd 0.007654f
C2446 vdd.n974 gnd 0.007654f
C2447 vdd.n975 gnd 0.007654f
C2448 vdd.n976 gnd 0.78221f
C2449 vdd.n977 gnd 0.007654f
C2450 vdd.n978 gnd 0.007654f
C2451 vdd.t6 gnd 0.391105f
C2452 vdd.n979 gnd 0.007654f
C2453 vdd.n980 gnd 0.007654f
C2454 vdd.n981 gnd 0.007654f
C2455 vdd.n982 gnd 0.007654f
C2456 vdd.n983 gnd 0.494633f
C2457 vdd.n984 gnd 0.007654f
C2458 vdd.n985 gnd 0.007654f
C2459 vdd.n986 gnd 0.007654f
C2460 vdd.n987 gnd 0.007654f
C2461 vdd.n988 gnd 0.007654f
C2462 vdd.n989 gnd 0.667179f
C2463 vdd.n990 gnd 0.007654f
C2464 vdd.n991 gnd 0.007654f
C2465 vdd.t289 gnd 0.350844f
C2466 vdd.t182 gnd 0.287577f
C2467 vdd.n992 gnd 0.007654f
C2468 vdd.n993 gnd 0.007654f
C2469 vdd.n994 gnd 0.007654f
C2470 vdd.t198 gnd 0.391105f
C2471 vdd.n995 gnd 0.007654f
C2472 vdd.n996 gnd 0.007654f
C2473 vdd.t2 gnd 0.391105f
C2474 vdd.n997 gnd 0.007654f
C2475 vdd.n998 gnd 0.007654f
C2476 vdd.n999 gnd 0.007654f
C2477 vdd.t206 gnd 0.304832f
C2478 vdd.n1000 gnd 0.007654f
C2479 vdd.n1001 gnd 0.007654f
C2480 vdd.n1002 gnd 0.649925f
C2481 vdd.n1003 gnd 0.007654f
C2482 vdd.n1004 gnd 0.007654f
C2483 vdd.n1005 gnd 0.007654f
C2484 vdd.t287 gnd 0.391105f
C2485 vdd.n1006 gnd 0.007654f
C2486 vdd.n1007 gnd 0.007654f
C2487 vdd.t195 gnd 0.33359f
C2488 vdd.n1008 gnd 0.477378f
C2489 vdd.n1009 gnd 0.007654f
C2490 vdd.n1010 gnd 0.007654f
C2491 vdd.n1011 gnd 0.007654f
C2492 vdd.n1012 gnd 0.649925f
C2493 vdd.n1013 gnd 0.007654f
C2494 vdd.n1014 gnd 0.007654f
C2495 vdd.t5 gnd 0.391105f
C2496 vdd.n1015 gnd 0.007654f
C2497 vdd.n1016 gnd 0.007654f
C2498 vdd.n1017 gnd 0.007654f
C2499 vdd.n1018 gnd 0.78221f
C2500 vdd.n1019 gnd 0.007654f
C2501 vdd.n1020 gnd 0.007654f
C2502 vdd.t184 gnd 0.391105f
C2503 vdd.n1021 gnd 0.007654f
C2504 vdd.n1022 gnd 0.007654f
C2505 vdd.n1023 gnd 0.007654f
C2506 vdd.t4 gnd 0.092025f
C2507 vdd.n1024 gnd 0.007654f
C2508 vdd.n1025 gnd 0.007654f
C2509 vdd.n1026 gnd 0.007654f
C2510 vdd.t270 gnd 0.316607f
C2511 vdd.t268 gnd 0.201923f
C2512 vdd.t271 gnd 0.316607f
C2513 vdd.n1027 gnd 0.177946f
C2514 vdd.n1028 gnd 0.007654f
C2515 vdd.n1029 gnd 0.007654f
C2516 vdd.n1030 gnd 0.78221f
C2517 vdd.n1031 gnd 0.007654f
C2518 vdd.n1032 gnd 0.007654f
C2519 vdd.t269 gnd 0.350844f
C2520 vdd.n1033 gnd 0.690186f
C2521 vdd.n1034 gnd 0.007654f
C2522 vdd.n1035 gnd 0.007654f
C2523 vdd.n1036 gnd 0.007654f
C2524 vdd.n1037 gnd 0.684434f
C2525 vdd.n1038 gnd 0.007654f
C2526 vdd.n1039 gnd 0.007654f
C2527 vdd.n1040 gnd 0.007654f
C2528 vdd.n1041 gnd 0.007654f
C2529 vdd.n1042 gnd 0.007654f
C2530 vdd.n1043 gnd 0.78221f
C2531 vdd.n1044 gnd 0.007654f
C2532 vdd.n1045 gnd 0.007654f
C2533 vdd.t212 gnd 0.391105f
C2534 vdd.n1046 gnd 0.007654f
C2535 vdd.n1047 gnd 0.018162f
C2536 vdd.n1048 gnd 0.018162f
C2537 vdd.n1049 gnd 7.92563f
C2538 vdd.n1050 gnd 0.016957f
C2539 vdd.n1051 gnd 0.016957f
C2540 vdd.n1052 gnd 0.018162f
C2541 vdd.n1053 gnd 0.007654f
C2542 vdd.n1054 gnd 0.007654f
C2543 vdd.n1055 gnd 0.007654f
C2544 vdd.n1056 gnd 0.007654f
C2545 vdd.n1057 gnd 0.007654f
C2546 vdd.n1058 gnd 0.007654f
C2547 vdd.n1059 gnd 0.007654f
C2548 vdd.n1060 gnd 0.007654f
C2549 vdd.n1062 gnd 0.007654f
C2550 vdd.n1063 gnd 0.007654f
C2551 vdd.n1064 gnd 0.007204f
C2552 vdd.n1067 gnd 0.027813f
C2553 vdd.n1068 gnd 0.00906f
C2554 vdd.n1069 gnd 0.011256f
C2555 vdd.n1071 gnd 0.011256f
C2556 vdd.n1072 gnd 0.00752f
C2557 vdd.t223 gnd 0.575155f
C2558 vdd.n1073 gnd 8.31674f
C2559 vdd.n1074 gnd 0.011256f
C2560 vdd.n1075 gnd 0.027813f
C2561 vdd.n1076 gnd 0.00906f
C2562 vdd.n1077 gnd 0.011256f
C2563 vdd.n1078 gnd 0.00906f
C2564 vdd.n1079 gnd 0.011256f
C2565 vdd.n1080 gnd 1.15031f
C2566 vdd.n1081 gnd 0.011256f
C2567 vdd.n1082 gnd 0.00906f
C2568 vdd.n1083 gnd 0.00906f
C2569 vdd.n1084 gnd 0.011256f
C2570 vdd.n1085 gnd 0.00906f
C2571 vdd.n1086 gnd 0.011256f
C2572 vdd.t21 gnd 0.575155f
C2573 vdd.n1087 gnd 0.011256f
C2574 vdd.n1088 gnd 0.00906f
C2575 vdd.n1089 gnd 0.011256f
C2576 vdd.n1090 gnd 0.00906f
C2577 vdd.n1091 gnd 0.011256f
C2578 vdd.t151 gnd 0.575155f
C2579 vdd.n1092 gnd 0.011256f
C2580 vdd.n1093 gnd 0.00906f
C2581 vdd.n1094 gnd 0.011256f
C2582 vdd.n1095 gnd 0.00906f
C2583 vdd.n1096 gnd 0.011256f
C2584 vdd.n1097 gnd 0.925999f
C2585 vdd.n1098 gnd 0.954757f
C2586 vdd.t35 gnd 0.575155f
C2587 vdd.n1099 gnd 0.011256f
C2588 vdd.n1100 gnd 0.00906f
C2589 vdd.n1101 gnd 0.011256f
C2590 vdd.n1102 gnd 0.00906f
C2591 vdd.n1103 gnd 0.011256f
C2592 vdd.n1104 gnd 0.730446f
C2593 vdd.n1105 gnd 0.011256f
C2594 vdd.n1106 gnd 0.00906f
C2595 vdd.n1107 gnd 0.011256f
C2596 vdd.n1108 gnd 0.00906f
C2597 vdd.n1109 gnd 0.011256f
C2598 vdd.t23 gnd 0.575155f
C2599 vdd.t65 gnd 0.575155f
C2600 vdd.n1110 gnd 0.011256f
C2601 vdd.n1111 gnd 0.00906f
C2602 vdd.n1112 gnd 0.011256f
C2603 vdd.n1113 gnd 0.00906f
C2604 vdd.n1114 gnd 0.011256f
C2605 vdd.t89 gnd 0.575155f
C2606 vdd.n1115 gnd 0.011256f
C2607 vdd.n1116 gnd 0.00906f
C2608 vdd.n1117 gnd 0.011256f
C2609 vdd.n1118 gnd 0.00906f
C2610 vdd.n1119 gnd 0.011256f
C2611 vdd.t128 gnd 0.575155f
C2612 vdd.n1120 gnd 0.810968f
C2613 vdd.n1121 gnd 0.011256f
C2614 vdd.n1122 gnd 0.00906f
C2615 vdd.n1123 gnd 0.011256f
C2616 vdd.n1124 gnd 0.00906f
C2617 vdd.n1125 gnd 0.011256f
C2618 vdd.n1126 gnd 0.902993f
C2619 vdd.n1127 gnd 0.011256f
C2620 vdd.n1128 gnd 0.00906f
C2621 vdd.n1129 gnd 0.011256f
C2622 vdd.n1130 gnd 0.00906f
C2623 vdd.n1131 gnd 0.011256f
C2624 vdd.n1132 gnd 0.70744f
C2625 vdd.t33 gnd 0.575155f
C2626 vdd.n1133 gnd 0.011256f
C2627 vdd.n1134 gnd 0.00906f
C2628 vdd.n1135 gnd 0.011256f
C2629 vdd.n1136 gnd 0.00906f
C2630 vdd.n1137 gnd 0.011256f
C2631 vdd.t43 gnd 0.575155f
C2632 vdd.n1138 gnd 0.011256f
C2633 vdd.n1139 gnd 0.00906f
C2634 vdd.n1140 gnd 0.011256f
C2635 vdd.n1141 gnd 0.00906f
C2636 vdd.n1142 gnd 0.011256f
C2637 vdd.t62 gnd 0.575155f
C2638 vdd.n1143 gnd 0.638422f
C2639 vdd.n1144 gnd 0.011256f
C2640 vdd.n1145 gnd 0.00906f
C2641 vdd.n1146 gnd 0.011256f
C2642 vdd.n1147 gnd 0.00906f
C2643 vdd.n1148 gnd 0.011256f
C2644 vdd.t107 gnd 0.575155f
C2645 vdd.n1149 gnd 0.011256f
C2646 vdd.n1150 gnd 0.00906f
C2647 vdd.n1151 gnd 0.011256f
C2648 vdd.n1152 gnd 0.00906f
C2649 vdd.n1153 gnd 0.011256f
C2650 vdd.n1154 gnd 0.879987f
C2651 vdd.n1155 gnd 0.954757f
C2652 vdd.t109 gnd 0.575155f
C2653 vdd.n1156 gnd 0.011256f
C2654 vdd.n1157 gnd 0.00906f
C2655 vdd.n1158 gnd 0.011256f
C2656 vdd.n1159 gnd 0.00906f
C2657 vdd.n1160 gnd 0.011256f
C2658 vdd.n1161 gnd 0.684434f
C2659 vdd.n1162 gnd 0.011256f
C2660 vdd.n1163 gnd 0.00906f
C2661 vdd.n1164 gnd 0.011256f
C2662 vdd.n1165 gnd 0.00906f
C2663 vdd.n1166 gnd 0.011256f
C2664 vdd.t60 gnd 0.575155f
C2665 vdd.t56 gnd 0.575155f
C2666 vdd.n1167 gnd 0.011256f
C2667 vdd.n1168 gnd 0.00906f
C2668 vdd.n1169 gnd 0.011256f
C2669 vdd.n1170 gnd 0.00906f
C2670 vdd.n1171 gnd 0.011256f
C2671 vdd.t19 gnd 0.575155f
C2672 vdd.n1172 gnd 0.011256f
C2673 vdd.n1173 gnd 0.00906f
C2674 vdd.n1174 gnd 0.011256f
C2675 vdd.n1175 gnd 0.00906f
C2676 vdd.n1176 gnd 0.011256f
C2677 vdd.t25 gnd 0.575155f
C2678 vdd.n1177 gnd 0.85698f
C2679 vdd.n1178 gnd 0.011256f
C2680 vdd.n1179 gnd 0.00906f
C2681 vdd.n1180 gnd 0.011256f
C2682 vdd.n1181 gnd 0.00906f
C2683 vdd.n1182 gnd 0.011256f
C2684 vdd.n1183 gnd 1.15031f
C2685 vdd.n1184 gnd 0.011256f
C2686 vdd.n1185 gnd 0.00906f
C2687 vdd.n1186 gnd 0.027229f
C2688 vdd.n1187 gnd 0.00752f
C2689 vdd.n1188 gnd 0.027229f
C2690 vdd.t231 gnd 0.575155f
C2691 vdd.n1189 gnd 0.027229f
C2692 vdd.n1190 gnd 0.00752f
C2693 vdd.n1191 gnd 0.011256f
C2694 vdd.n1192 gnd 0.00906f
C2695 vdd.n1193 gnd 0.011256f
C2696 vdd.n1224 gnd 0.027813f
C2697 vdd.n1225 gnd 1.69671f
C2698 vdd.n1226 gnd 0.011256f
C2699 vdd.n1227 gnd 0.00906f
C2700 vdd.n1228 gnd 0.011256f
C2701 vdd.n1229 gnd 0.011256f
C2702 vdd.n1230 gnd 0.011256f
C2703 vdd.n1231 gnd 0.011256f
C2704 vdd.n1232 gnd 0.011256f
C2705 vdd.n1233 gnd 0.00906f
C2706 vdd.n1234 gnd 0.011256f
C2707 vdd.n1235 gnd 0.011256f
C2708 vdd.n1236 gnd 0.011256f
C2709 vdd.n1237 gnd 0.011256f
C2710 vdd.n1238 gnd 0.011256f
C2711 vdd.n1239 gnd 0.00906f
C2712 vdd.n1240 gnd 0.011256f
C2713 vdd.n1241 gnd 0.011256f
C2714 vdd.n1242 gnd 0.011256f
C2715 vdd.n1243 gnd 0.011256f
C2716 vdd.n1244 gnd 0.011256f
C2717 vdd.n1245 gnd 0.00906f
C2718 vdd.n1246 gnd 0.011256f
C2719 vdd.n1247 gnd 0.011256f
C2720 vdd.n1248 gnd 0.011256f
C2721 vdd.n1249 gnd 0.011256f
C2722 vdd.n1250 gnd 0.011256f
C2723 vdd.t245 gnd 0.138478f
C2724 vdd.t246 gnd 0.147995f
C2725 vdd.t244 gnd 0.180851f
C2726 vdd.n1251 gnd 0.231825f
C2727 vdd.n1252 gnd 0.195681f
C2728 vdd.n1253 gnd 0.019388f
C2729 vdd.n1254 gnd 0.011256f
C2730 vdd.n1255 gnd 0.011256f
C2731 vdd.n1256 gnd 0.011256f
C2732 vdd.n1257 gnd 0.011256f
C2733 vdd.n1258 gnd 0.011256f
C2734 vdd.n1259 gnd 0.00906f
C2735 vdd.n1260 gnd 0.011256f
C2736 vdd.n1261 gnd 0.011256f
C2737 vdd.n1262 gnd 0.011256f
C2738 vdd.n1263 gnd 0.011256f
C2739 vdd.n1264 gnd 0.011256f
C2740 vdd.n1265 gnd 0.00906f
C2741 vdd.n1266 gnd 0.011256f
C2742 vdd.n1267 gnd 0.011256f
C2743 vdd.n1268 gnd 0.011256f
C2744 vdd.n1269 gnd 0.011256f
C2745 vdd.n1270 gnd 0.011256f
C2746 vdd.n1271 gnd 0.00906f
C2747 vdd.n1272 gnd 0.011256f
C2748 vdd.n1273 gnd 0.011256f
C2749 vdd.n1274 gnd 0.011256f
C2750 vdd.n1275 gnd 0.011256f
C2751 vdd.n1276 gnd 0.011256f
C2752 vdd.n1277 gnd 0.00906f
C2753 vdd.n1278 gnd 0.011256f
C2754 vdd.n1279 gnd 0.011256f
C2755 vdd.n1280 gnd 0.011256f
C2756 vdd.n1281 gnd 0.011256f
C2757 vdd.n1282 gnd 0.011256f
C2758 vdd.n1283 gnd 0.00906f
C2759 vdd.n1284 gnd 0.011256f
C2760 vdd.n1285 gnd 0.011256f
C2761 vdd.n1286 gnd 0.011256f
C2762 vdd.n1287 gnd 0.011256f
C2763 vdd.n1288 gnd 0.00906f
C2764 vdd.n1289 gnd 0.011256f
C2765 vdd.n1290 gnd 0.011256f
C2766 vdd.n1291 gnd 0.011256f
C2767 vdd.n1292 gnd 0.011256f
C2768 vdd.n1293 gnd 0.011256f
C2769 vdd.n1294 gnd 0.00906f
C2770 vdd.n1295 gnd 0.011256f
C2771 vdd.n1296 gnd 0.011256f
C2772 vdd.n1297 gnd 0.011256f
C2773 vdd.n1298 gnd 0.011256f
C2774 vdd.n1299 gnd 0.011256f
C2775 vdd.n1300 gnd 0.00906f
C2776 vdd.n1301 gnd 0.011256f
C2777 vdd.n1302 gnd 0.011256f
C2778 vdd.n1303 gnd 0.011256f
C2779 vdd.n1304 gnd 0.011256f
C2780 vdd.n1305 gnd 0.011256f
C2781 vdd.n1306 gnd 0.00906f
C2782 vdd.n1307 gnd 0.011256f
C2783 vdd.n1308 gnd 0.011256f
C2784 vdd.n1309 gnd 0.011256f
C2785 vdd.n1310 gnd 0.011256f
C2786 vdd.n1311 gnd 0.011256f
C2787 vdd.n1312 gnd 0.00906f
C2788 vdd.n1313 gnd 0.011256f
C2789 vdd.n1314 gnd 0.011256f
C2790 vdd.n1315 gnd 0.011256f
C2791 vdd.n1316 gnd 0.011256f
C2792 vdd.t242 gnd 0.138478f
C2793 vdd.t243 gnd 0.147995f
C2794 vdd.t241 gnd 0.180851f
C2795 vdd.n1317 gnd 0.231825f
C2796 vdd.n1318 gnd 0.195681f
C2797 vdd.n1319 gnd 0.014858f
C2798 vdd.n1320 gnd 0.004303f
C2799 vdd.n1321 gnd 0.027813f
C2800 vdd.n1322 gnd 0.011256f
C2801 vdd.n1323 gnd 0.004756f
C2802 vdd.n1324 gnd 0.00906f
C2803 vdd.n1325 gnd 0.00906f
C2804 vdd.n1326 gnd 0.011256f
C2805 vdd.n1327 gnd 0.011256f
C2806 vdd.n1328 gnd 0.011256f
C2807 vdd.n1329 gnd 0.00906f
C2808 vdd.n1330 gnd 0.00906f
C2809 vdd.n1331 gnd 0.00906f
C2810 vdd.n1332 gnd 0.011256f
C2811 vdd.n1333 gnd 0.011256f
C2812 vdd.n1334 gnd 0.011256f
C2813 vdd.n1335 gnd 0.00906f
C2814 vdd.n1336 gnd 0.00906f
C2815 vdd.n1337 gnd 0.00906f
C2816 vdd.n1338 gnd 0.011256f
C2817 vdd.n1339 gnd 0.011256f
C2818 vdd.n1340 gnd 0.011256f
C2819 vdd.n1341 gnd 0.00906f
C2820 vdd.n1342 gnd 0.00906f
C2821 vdd.n1343 gnd 0.00906f
C2822 vdd.n1344 gnd 0.011256f
C2823 vdd.n1345 gnd 0.011256f
C2824 vdd.n1346 gnd 0.011256f
C2825 vdd.n1347 gnd 0.00906f
C2826 vdd.n1348 gnd 0.00906f
C2827 vdd.n1349 gnd 0.00906f
C2828 vdd.n1350 gnd 0.011256f
C2829 vdd.n1351 gnd 0.011256f
C2830 vdd.n1352 gnd 0.011256f
C2831 vdd.n1353 gnd 0.008969f
C2832 vdd.n1354 gnd 0.011256f
C2833 vdd.t232 gnd 0.138478f
C2834 vdd.t233 gnd 0.147995f
C2835 vdd.t230 gnd 0.180851f
C2836 vdd.n1355 gnd 0.231825f
C2837 vdd.n1356 gnd 0.195681f
C2838 vdd.n1357 gnd 0.019388f
C2839 vdd.n1358 gnd 0.006161f
C2840 vdd.n1359 gnd 0.011256f
C2841 vdd.n1360 gnd 0.011256f
C2842 vdd.n1361 gnd 0.011256f
C2843 vdd.n1362 gnd 0.00906f
C2844 vdd.n1363 gnd 0.00906f
C2845 vdd.n1364 gnd 0.00906f
C2846 vdd.n1365 gnd 0.011256f
C2847 vdd.n1366 gnd 0.011256f
C2848 vdd.n1367 gnd 0.011256f
C2849 vdd.n1368 gnd 0.00906f
C2850 vdd.n1369 gnd 0.00906f
C2851 vdd.n1370 gnd 0.00906f
C2852 vdd.n1371 gnd 0.011256f
C2853 vdd.n1372 gnd 0.011256f
C2854 vdd.n1373 gnd 0.011256f
C2855 vdd.n1374 gnd 0.00906f
C2856 vdd.n1375 gnd 0.00906f
C2857 vdd.n1376 gnd 0.00906f
C2858 vdd.n1377 gnd 0.011256f
C2859 vdd.n1378 gnd 0.011256f
C2860 vdd.n1379 gnd 0.011256f
C2861 vdd.n1380 gnd 0.00906f
C2862 vdd.n1381 gnd 0.00906f
C2863 vdd.n1382 gnd 0.00906f
C2864 vdd.n1383 gnd 0.011256f
C2865 vdd.n1384 gnd 0.011256f
C2866 vdd.n1385 gnd 0.011256f
C2867 vdd.n1386 gnd 0.00906f
C2868 vdd.n1387 gnd 0.00906f
C2869 vdd.n1388 gnd 0.007565f
C2870 vdd.n1389 gnd 0.011256f
C2871 vdd.n1390 gnd 0.011256f
C2872 vdd.n1391 gnd 0.011256f
C2873 vdd.n1392 gnd 0.007565f
C2874 vdd.n1393 gnd 0.00906f
C2875 vdd.n1394 gnd 0.00906f
C2876 vdd.n1395 gnd 0.011256f
C2877 vdd.n1396 gnd 0.011256f
C2878 vdd.n1397 gnd 0.011256f
C2879 vdd.n1398 gnd 0.00906f
C2880 vdd.n1399 gnd 0.00906f
C2881 vdd.n1400 gnd 0.00906f
C2882 vdd.n1401 gnd 0.011256f
C2883 vdd.n1402 gnd 0.011256f
C2884 vdd.n1403 gnd 0.011256f
C2885 vdd.n1404 gnd 0.00906f
C2886 vdd.n1405 gnd 0.00906f
C2887 vdd.n1406 gnd 0.00906f
C2888 vdd.n1407 gnd 0.011256f
C2889 vdd.n1408 gnd 0.011256f
C2890 vdd.n1409 gnd 0.011256f
C2891 vdd.n1410 gnd 0.00906f
C2892 vdd.n1411 gnd 0.00906f
C2893 vdd.n1412 gnd 0.00906f
C2894 vdd.n1413 gnd 0.011256f
C2895 vdd.n1414 gnd 0.011256f
C2896 vdd.n1415 gnd 0.011256f
C2897 vdd.n1416 gnd 0.00906f
C2898 vdd.n1417 gnd 0.011256f
C2899 vdd.n1418 gnd 2.72623f
C2900 vdd.n1420 gnd 0.027813f
C2901 vdd.n1421 gnd 0.00752f
C2902 vdd.n1422 gnd 0.027813f
C2903 vdd.n1423 gnd 0.027229f
C2904 vdd.n1424 gnd 0.011256f
C2905 vdd.n1425 gnd 0.00906f
C2906 vdd.n1426 gnd 0.011256f
C2907 vdd.n1427 gnd 0.580906f
C2908 vdd.n1428 gnd 0.011256f
C2909 vdd.n1429 gnd 0.00906f
C2910 vdd.n1430 gnd 0.011256f
C2911 vdd.n1431 gnd 0.011256f
C2912 vdd.n1432 gnd 0.011256f
C2913 vdd.n1433 gnd 0.00906f
C2914 vdd.n1434 gnd 0.011256f
C2915 vdd.n1435 gnd 1.05253f
C2916 vdd.n1436 gnd 1.15031f
C2917 vdd.n1437 gnd 0.011256f
C2918 vdd.n1438 gnd 0.00906f
C2919 vdd.n1439 gnd 0.011256f
C2920 vdd.n1440 gnd 0.011256f
C2921 vdd.n1441 gnd 0.011256f
C2922 vdd.n1442 gnd 0.00906f
C2923 vdd.n1443 gnd 0.011256f
C2924 vdd.n1444 gnd 0.672931f
C2925 vdd.n1445 gnd 0.011256f
C2926 vdd.n1446 gnd 0.00906f
C2927 vdd.n1447 gnd 0.011256f
C2928 vdd.n1448 gnd 0.011256f
C2929 vdd.n1449 gnd 0.011256f
C2930 vdd.n1450 gnd 0.00906f
C2931 vdd.n1451 gnd 0.011256f
C2932 vdd.n1452 gnd 0.661428f
C2933 vdd.n1453 gnd 0.868483f
C2934 vdd.n1454 gnd 0.011256f
C2935 vdd.n1455 gnd 0.00906f
C2936 vdd.n1456 gnd 0.011256f
C2937 vdd.n1457 gnd 0.011256f
C2938 vdd.n1458 gnd 0.011256f
C2939 vdd.n1459 gnd 0.00906f
C2940 vdd.n1460 gnd 0.011256f
C2941 vdd.n1461 gnd 0.954757f
C2942 vdd.n1462 gnd 0.011256f
C2943 vdd.n1463 gnd 0.00906f
C2944 vdd.n1464 gnd 0.011256f
C2945 vdd.n1465 gnd 0.011256f
C2946 vdd.n1466 gnd 0.011256f
C2947 vdd.n1467 gnd 0.00906f
C2948 vdd.n1468 gnd 0.011256f
C2949 vdd.t31 gnd 0.575155f
C2950 vdd.n1469 gnd 0.845477f
C2951 vdd.n1470 gnd 0.011256f
C2952 vdd.n1471 gnd 0.00906f
C2953 vdd.n1472 gnd 0.011256f
C2954 vdd.n1473 gnd 0.011256f
C2955 vdd.n1474 gnd 0.011256f
C2956 vdd.n1475 gnd 0.00906f
C2957 vdd.n1476 gnd 0.011256f
C2958 vdd.n1477 gnd 0.649925f
C2959 vdd.n1478 gnd 0.011256f
C2960 vdd.n1479 gnd 0.00906f
C2961 vdd.n1480 gnd 0.011256f
C2962 vdd.n1481 gnd 0.011256f
C2963 vdd.n1482 gnd 0.011256f
C2964 vdd.n1483 gnd 0.00906f
C2965 vdd.n1484 gnd 0.011256f
C2966 vdd.n1485 gnd 0.833974f
C2967 vdd.n1486 gnd 0.695937f
C2968 vdd.n1487 gnd 0.011256f
C2969 vdd.n1488 gnd 0.00906f
C2970 vdd.n1489 gnd 0.011256f
C2971 vdd.n1490 gnd 0.011256f
C2972 vdd.n1491 gnd 0.011256f
C2973 vdd.n1492 gnd 0.00906f
C2974 vdd.n1493 gnd 0.011256f
C2975 vdd.n1494 gnd 0.89149f
C2976 vdd.n1495 gnd 0.011256f
C2977 vdd.n1496 gnd 0.00906f
C2978 vdd.n1497 gnd 0.011256f
C2979 vdd.n1498 gnd 0.011256f
C2980 vdd.n1499 gnd 0.011256f
C2981 vdd.n1500 gnd 0.00906f
C2982 vdd.n1501 gnd 0.011256f
C2983 vdd.t79 gnd 0.575155f
C2984 vdd.n1502 gnd 0.954757f
C2985 vdd.n1503 gnd 0.011256f
C2986 vdd.n1504 gnd 0.00906f
C2987 vdd.n1505 gnd 0.011256f
C2988 vdd.n1506 gnd 0.008651f
C2989 vdd.n1507 gnd 0.006177f
C2990 vdd.n1508 gnd 0.005732f
C2991 vdd.n1509 gnd 0.003171f
C2992 vdd.n1510 gnd 0.007281f
C2993 vdd.n1511 gnd 0.00308f
C2994 vdd.n1512 gnd 0.003262f
C2995 vdd.n1513 gnd 0.005732f
C2996 vdd.n1514 gnd 0.00308f
C2997 vdd.n1515 gnd 0.007281f
C2998 vdd.n1516 gnd 0.003262f
C2999 vdd.n1517 gnd 0.005732f
C3000 vdd.n1518 gnd 0.00308f
C3001 vdd.n1519 gnd 0.005461f
C3002 vdd.n1520 gnd 0.005477f
C3003 vdd.t22 gnd 0.015642f
C3004 vdd.n1521 gnd 0.034803f
C3005 vdd.n1522 gnd 0.181124f
C3006 vdd.n1523 gnd 0.00308f
C3007 vdd.n1524 gnd 0.003262f
C3008 vdd.n1525 gnd 0.007281f
C3009 vdd.n1526 gnd 0.007281f
C3010 vdd.n1527 gnd 0.003262f
C3011 vdd.n1528 gnd 0.00308f
C3012 vdd.n1529 gnd 0.005732f
C3013 vdd.n1530 gnd 0.005732f
C3014 vdd.n1531 gnd 0.00308f
C3015 vdd.n1532 gnd 0.003262f
C3016 vdd.n1533 gnd 0.007281f
C3017 vdd.n1534 gnd 0.007281f
C3018 vdd.n1535 gnd 0.003262f
C3019 vdd.n1536 gnd 0.00308f
C3020 vdd.n1537 gnd 0.005732f
C3021 vdd.n1538 gnd 0.005732f
C3022 vdd.n1539 gnd 0.00308f
C3023 vdd.n1540 gnd 0.003262f
C3024 vdd.n1541 gnd 0.007281f
C3025 vdd.n1542 gnd 0.007281f
C3026 vdd.n1543 gnd 0.017213f
C3027 vdd.n1544 gnd 0.003171f
C3028 vdd.n1545 gnd 0.00308f
C3029 vdd.n1546 gnd 0.014816f
C3030 vdd.n1547 gnd 0.010344f
C3031 vdd.t99 gnd 0.036239f
C3032 vdd.t161 gnd 0.036239f
C3033 vdd.n1548 gnd 0.249058f
C3034 vdd.n1549 gnd 0.195846f
C3035 vdd.t66 gnd 0.036239f
C3036 vdd.t138 gnd 0.036239f
C3037 vdd.n1550 gnd 0.249058f
C3038 vdd.n1551 gnd 0.158047f
C3039 vdd.t90 gnd 0.036239f
C3040 vdd.t147 gnd 0.036239f
C3041 vdd.n1552 gnd 0.249058f
C3042 vdd.n1553 gnd 0.158047f
C3043 vdd.t113 gnd 0.036239f
C3044 vdd.t168 gnd 0.036239f
C3045 vdd.n1554 gnd 0.249058f
C3046 vdd.n1555 gnd 0.158047f
C3047 vdd.t80 gnd 0.036239f
C3048 vdd.t34 gnd 0.036239f
C3049 vdd.n1556 gnd 0.249058f
C3050 vdd.n1557 gnd 0.158047f
C3051 vdd.t102 gnd 0.036239f
C3052 vdd.t44 gnd 0.036239f
C3053 vdd.n1558 gnd 0.249058f
C3054 vdd.n1559 gnd 0.158047f
C3055 vdd.t155 gnd 0.036239f
C3056 vdd.t172 gnd 0.036239f
C3057 vdd.n1560 gnd 0.249058f
C3058 vdd.n1561 gnd 0.158047f
C3059 vdd.t127 gnd 0.036239f
C3060 vdd.t47 gnd 0.036239f
C3061 vdd.n1562 gnd 0.249058f
C3062 vdd.n1563 gnd 0.158047f
C3063 vdd.t114 gnd 0.036239f
C3064 vdd.t61 gnd 0.036239f
C3065 vdd.n1564 gnd 0.249058f
C3066 vdd.n1565 gnd 0.158047f
C3067 vdd.n1566 gnd 0.006177f
C3068 vdd.n1567 gnd 0.005732f
C3069 vdd.n1568 gnd 0.003171f
C3070 vdd.n1569 gnd 0.007281f
C3071 vdd.n1570 gnd 0.00308f
C3072 vdd.n1571 gnd 0.003262f
C3073 vdd.n1572 gnd 0.005732f
C3074 vdd.n1573 gnd 0.00308f
C3075 vdd.n1574 gnd 0.007281f
C3076 vdd.n1575 gnd 0.003262f
C3077 vdd.n1576 gnd 0.005732f
C3078 vdd.n1577 gnd 0.00308f
C3079 vdd.n1578 gnd 0.005461f
C3080 vdd.n1579 gnd 0.005477f
C3081 vdd.t84 gnd 0.015642f
C3082 vdd.n1580 gnd 0.034803f
C3083 vdd.n1581 gnd 0.181124f
C3084 vdd.n1582 gnd 0.00308f
C3085 vdd.n1583 gnd 0.003262f
C3086 vdd.n1584 gnd 0.007281f
C3087 vdd.n1585 gnd 0.007281f
C3088 vdd.n1586 gnd 0.003262f
C3089 vdd.n1587 gnd 0.00308f
C3090 vdd.n1588 gnd 0.005732f
C3091 vdd.n1589 gnd 0.005732f
C3092 vdd.n1590 gnd 0.00308f
C3093 vdd.n1591 gnd 0.003262f
C3094 vdd.n1592 gnd 0.007281f
C3095 vdd.n1593 gnd 0.007281f
C3096 vdd.n1594 gnd 0.003262f
C3097 vdd.n1595 gnd 0.00308f
C3098 vdd.n1596 gnd 0.005732f
C3099 vdd.n1597 gnd 0.005732f
C3100 vdd.n1598 gnd 0.00308f
C3101 vdd.n1599 gnd 0.003262f
C3102 vdd.n1600 gnd 0.007281f
C3103 vdd.n1601 gnd 0.007281f
C3104 vdd.n1602 gnd 0.017213f
C3105 vdd.n1603 gnd 0.003171f
C3106 vdd.n1604 gnd 0.00308f
C3107 vdd.n1605 gnd 0.014816f
C3108 vdd.n1606 gnd 0.010019f
C3109 vdd.n1607 gnd 0.117588f
C3110 vdd.n1608 gnd 0.006177f
C3111 vdd.n1609 gnd 0.005732f
C3112 vdd.n1610 gnd 0.003171f
C3113 vdd.n1611 gnd 0.007281f
C3114 vdd.n1612 gnd 0.00308f
C3115 vdd.n1613 gnd 0.003262f
C3116 vdd.n1614 gnd 0.005732f
C3117 vdd.n1615 gnd 0.00308f
C3118 vdd.n1616 gnd 0.007281f
C3119 vdd.n1617 gnd 0.003262f
C3120 vdd.n1618 gnd 0.005732f
C3121 vdd.n1619 gnd 0.00308f
C3122 vdd.n1620 gnd 0.005461f
C3123 vdd.n1621 gnd 0.005477f
C3124 vdd.t149 gnd 0.015642f
C3125 vdd.n1622 gnd 0.034803f
C3126 vdd.n1623 gnd 0.181124f
C3127 vdd.n1624 gnd 0.00308f
C3128 vdd.n1625 gnd 0.003262f
C3129 vdd.n1626 gnd 0.007281f
C3130 vdd.n1627 gnd 0.007281f
C3131 vdd.n1628 gnd 0.003262f
C3132 vdd.n1629 gnd 0.00308f
C3133 vdd.n1630 gnd 0.005732f
C3134 vdd.n1631 gnd 0.005732f
C3135 vdd.n1632 gnd 0.00308f
C3136 vdd.n1633 gnd 0.003262f
C3137 vdd.n1634 gnd 0.007281f
C3138 vdd.n1635 gnd 0.007281f
C3139 vdd.n1636 gnd 0.003262f
C3140 vdd.n1637 gnd 0.00308f
C3141 vdd.n1638 gnd 0.005732f
C3142 vdd.n1639 gnd 0.005732f
C3143 vdd.n1640 gnd 0.00308f
C3144 vdd.n1641 gnd 0.003262f
C3145 vdd.n1642 gnd 0.007281f
C3146 vdd.n1643 gnd 0.007281f
C3147 vdd.n1644 gnd 0.017213f
C3148 vdd.n1645 gnd 0.003171f
C3149 vdd.n1646 gnd 0.00308f
C3150 vdd.n1647 gnd 0.014816f
C3151 vdd.n1648 gnd 0.010344f
C3152 vdd.t36 gnd 0.036239f
C3153 vdd.t152 gnd 0.036239f
C3154 vdd.n1649 gnd 0.249058f
C3155 vdd.n1650 gnd 0.195846f
C3156 vdd.t145 gnd 0.036239f
C3157 vdd.t131 gnd 0.036239f
C3158 vdd.n1651 gnd 0.249058f
C3159 vdd.n1652 gnd 0.158047f
C3160 vdd.t92 gnd 0.036239f
C3161 vdd.t24 gnd 0.036239f
C3162 vdd.n1653 gnd 0.249058f
C3163 vdd.n1654 gnd 0.158047f
C3164 vdd.t163 gnd 0.036239f
C3165 vdd.t129 gnd 0.036239f
C3166 vdd.n1655 gnd 0.249058f
C3167 vdd.n1656 gnd 0.158047f
C3168 vdd.t123 gnd 0.036239f
C3169 vdd.t67 gnd 0.036239f
C3170 vdd.n1657 gnd 0.249058f
C3171 vdd.n1658 gnd 0.158047f
C3172 vdd.t63 gnd 0.036239f
C3173 vdd.t124 gnd 0.036239f
C3174 vdd.n1659 gnd 0.249058f
C3175 vdd.n1660 gnd 0.158047f
C3176 vdd.t110 gnd 0.036239f
C3177 vdd.t108 gnd 0.036239f
C3178 vdd.n1661 gnd 0.249058f
C3179 vdd.n1662 gnd 0.158047f
C3180 vdd.t57 gnd 0.036239f
C3181 vdd.t32 gnd 0.036239f
C3182 vdd.n1663 gnd 0.249058f
C3183 vdd.n1664 gnd 0.158047f
C3184 vdd.t20 gnd 0.036239f
C3185 vdd.t103 gnd 0.036239f
C3186 vdd.n1665 gnd 0.249058f
C3187 vdd.n1666 gnd 0.158047f
C3188 vdd.n1667 gnd 0.006177f
C3189 vdd.n1668 gnd 0.005732f
C3190 vdd.n1669 gnd 0.003171f
C3191 vdd.n1670 gnd 0.007281f
C3192 vdd.n1671 gnd 0.00308f
C3193 vdd.n1672 gnd 0.003262f
C3194 vdd.n1673 gnd 0.005732f
C3195 vdd.n1674 gnd 0.00308f
C3196 vdd.n1675 gnd 0.007281f
C3197 vdd.n1676 gnd 0.003262f
C3198 vdd.n1677 gnd 0.005732f
C3199 vdd.n1678 gnd 0.00308f
C3200 vdd.n1679 gnd 0.005461f
C3201 vdd.n1680 gnd 0.005477f
C3202 vdd.t26 gnd 0.015642f
C3203 vdd.n1681 gnd 0.034803f
C3204 vdd.n1682 gnd 0.181124f
C3205 vdd.n1683 gnd 0.00308f
C3206 vdd.n1684 gnd 0.003262f
C3207 vdd.n1685 gnd 0.007281f
C3208 vdd.n1686 gnd 0.007281f
C3209 vdd.n1687 gnd 0.003262f
C3210 vdd.n1688 gnd 0.00308f
C3211 vdd.n1689 gnd 0.005732f
C3212 vdd.n1690 gnd 0.005732f
C3213 vdd.n1691 gnd 0.00308f
C3214 vdd.n1692 gnd 0.003262f
C3215 vdd.n1693 gnd 0.007281f
C3216 vdd.n1694 gnd 0.007281f
C3217 vdd.n1695 gnd 0.003262f
C3218 vdd.n1696 gnd 0.00308f
C3219 vdd.n1697 gnd 0.005732f
C3220 vdd.n1698 gnd 0.005732f
C3221 vdd.n1699 gnd 0.00308f
C3222 vdd.n1700 gnd 0.003262f
C3223 vdd.n1701 gnd 0.007281f
C3224 vdd.n1702 gnd 0.007281f
C3225 vdd.n1703 gnd 0.017213f
C3226 vdd.n1704 gnd 0.003171f
C3227 vdd.n1705 gnd 0.00308f
C3228 vdd.n1706 gnd 0.014816f
C3229 vdd.n1707 gnd 0.010019f
C3230 vdd.n1708 gnd 0.069953f
C3231 vdd.n1709 gnd 0.252058f
C3232 vdd.n1710 gnd 0.006177f
C3233 vdd.n1711 gnd 0.005732f
C3234 vdd.n1712 gnd 0.003171f
C3235 vdd.n1713 gnd 0.007281f
C3236 vdd.n1714 gnd 0.00308f
C3237 vdd.n1715 gnd 0.003262f
C3238 vdd.n1716 gnd 0.005732f
C3239 vdd.n1717 gnd 0.00308f
C3240 vdd.n1718 gnd 0.007281f
C3241 vdd.n1719 gnd 0.003262f
C3242 vdd.n1720 gnd 0.005732f
C3243 vdd.n1721 gnd 0.00308f
C3244 vdd.n1722 gnd 0.005461f
C3245 vdd.n1723 gnd 0.005477f
C3246 vdd.t164 gnd 0.015642f
C3247 vdd.n1724 gnd 0.034803f
C3248 vdd.n1725 gnd 0.181124f
C3249 vdd.n1726 gnd 0.00308f
C3250 vdd.n1727 gnd 0.003262f
C3251 vdd.n1728 gnd 0.007281f
C3252 vdd.n1729 gnd 0.007281f
C3253 vdd.n1730 gnd 0.003262f
C3254 vdd.n1731 gnd 0.00308f
C3255 vdd.n1732 gnd 0.005732f
C3256 vdd.n1733 gnd 0.005732f
C3257 vdd.n1734 gnd 0.00308f
C3258 vdd.n1735 gnd 0.003262f
C3259 vdd.n1736 gnd 0.007281f
C3260 vdd.n1737 gnd 0.007281f
C3261 vdd.n1738 gnd 0.003262f
C3262 vdd.n1739 gnd 0.00308f
C3263 vdd.n1740 gnd 0.005732f
C3264 vdd.n1741 gnd 0.005732f
C3265 vdd.n1742 gnd 0.00308f
C3266 vdd.n1743 gnd 0.003262f
C3267 vdd.n1744 gnd 0.007281f
C3268 vdd.n1745 gnd 0.007281f
C3269 vdd.n1746 gnd 0.017213f
C3270 vdd.n1747 gnd 0.003171f
C3271 vdd.n1748 gnd 0.00308f
C3272 vdd.n1749 gnd 0.014816f
C3273 vdd.n1750 gnd 0.010344f
C3274 vdd.t53 gnd 0.036239f
C3275 vdd.t165 gnd 0.036239f
C3276 vdd.n1751 gnd 0.249058f
C3277 vdd.n1752 gnd 0.195846f
C3278 vdd.t159 gnd 0.036239f
C3279 vdd.t142 gnd 0.036239f
C3280 vdd.n1753 gnd 0.249058f
C3281 vdd.n1754 gnd 0.158047f
C3282 vdd.t111 gnd 0.036239f
C3283 vdd.t49 gnd 0.036239f
C3284 vdd.n1755 gnd 0.249058f
C3285 vdd.n1756 gnd 0.158047f
C3286 vdd.t173 gnd 0.036239f
C3287 vdd.t139 gnd 0.036239f
C3288 vdd.n1757 gnd 0.249058f
C3289 vdd.n1758 gnd 0.158047f
C3290 vdd.t115 gnd 0.036239f
C3291 vdd.t85 gnd 0.036239f
C3292 vdd.n1759 gnd 0.249058f
C3293 vdd.n1760 gnd 0.158047f
C3294 vdd.t81 gnd 0.036239f
C3295 vdd.t137 gnd 0.036239f
C3296 vdd.n1761 gnd 0.249058f
C3297 vdd.n1762 gnd 0.158047f
C3298 vdd.t122 gnd 0.036239f
C3299 vdd.t120 gnd 0.036239f
C3300 vdd.n1763 gnd 0.249058f
C3301 vdd.n1764 gnd 0.158047f
C3302 vdd.t78 gnd 0.036239f
C3303 vdd.t52 gnd 0.036239f
C3304 vdd.n1765 gnd 0.249058f
C3305 vdd.n1766 gnd 0.158047f
C3306 vdd.t48 gnd 0.036239f
C3307 vdd.t118 gnd 0.036239f
C3308 vdd.n1767 gnd 0.249058f
C3309 vdd.n1768 gnd 0.158047f
C3310 vdd.n1769 gnd 0.006177f
C3311 vdd.n1770 gnd 0.005732f
C3312 vdd.n1771 gnd 0.003171f
C3313 vdd.n1772 gnd 0.007281f
C3314 vdd.n1773 gnd 0.00308f
C3315 vdd.n1774 gnd 0.003262f
C3316 vdd.n1775 gnd 0.005732f
C3317 vdd.n1776 gnd 0.00308f
C3318 vdd.n1777 gnd 0.007281f
C3319 vdd.n1778 gnd 0.003262f
C3320 vdd.n1779 gnd 0.005732f
C3321 vdd.n1780 gnd 0.00308f
C3322 vdd.n1781 gnd 0.005461f
C3323 vdd.n1782 gnd 0.005477f
C3324 vdd.t50 gnd 0.015642f
C3325 vdd.n1783 gnd 0.034803f
C3326 vdd.n1784 gnd 0.181124f
C3327 vdd.n1785 gnd 0.00308f
C3328 vdd.n1786 gnd 0.003262f
C3329 vdd.n1787 gnd 0.007281f
C3330 vdd.n1788 gnd 0.007281f
C3331 vdd.n1789 gnd 0.003262f
C3332 vdd.n1790 gnd 0.00308f
C3333 vdd.n1791 gnd 0.005732f
C3334 vdd.n1792 gnd 0.005732f
C3335 vdd.n1793 gnd 0.00308f
C3336 vdd.n1794 gnd 0.003262f
C3337 vdd.n1795 gnd 0.007281f
C3338 vdd.n1796 gnd 0.007281f
C3339 vdd.n1797 gnd 0.003262f
C3340 vdd.n1798 gnd 0.00308f
C3341 vdd.n1799 gnd 0.005732f
C3342 vdd.n1800 gnd 0.005732f
C3343 vdd.n1801 gnd 0.00308f
C3344 vdd.n1802 gnd 0.003262f
C3345 vdd.n1803 gnd 0.007281f
C3346 vdd.n1804 gnd 0.007281f
C3347 vdd.n1805 gnd 0.017213f
C3348 vdd.n1806 gnd 0.003171f
C3349 vdd.n1807 gnd 0.00308f
C3350 vdd.n1808 gnd 0.014816f
C3351 vdd.n1809 gnd 0.010019f
C3352 vdd.n1810 gnd 0.069953f
C3353 vdd.n1811 gnd 0.288552f
C3354 vdd.n1812 gnd 2.89099f
C3355 vdd.n1813 gnd 0.663921f
C3356 vdd.n1814 gnd 0.008651f
C3357 vdd.n1815 gnd 0.00906f
C3358 vdd.n1816 gnd 0.011256f
C3359 vdd.n1817 gnd 0.822471f
C3360 vdd.n1818 gnd 0.011256f
C3361 vdd.n1819 gnd 0.00906f
C3362 vdd.n1820 gnd 0.011256f
C3363 vdd.n1821 gnd 0.011256f
C3364 vdd.n1822 gnd 0.011256f
C3365 vdd.n1823 gnd 0.00906f
C3366 vdd.n1824 gnd 0.011256f
C3367 vdd.n1825 gnd 0.954757f
C3368 vdd.t112 gnd 0.575155f
C3369 vdd.n1826 gnd 0.626919f
C3370 vdd.n1827 gnd 0.011256f
C3371 vdd.n1828 gnd 0.00906f
C3372 vdd.n1829 gnd 0.011256f
C3373 vdd.n1830 gnd 0.011256f
C3374 vdd.n1831 gnd 0.011256f
C3375 vdd.n1832 gnd 0.00906f
C3376 vdd.n1833 gnd 0.011256f
C3377 vdd.n1834 gnd 0.718943f
C3378 vdd.n1835 gnd 0.011256f
C3379 vdd.n1836 gnd 0.00906f
C3380 vdd.n1837 gnd 0.011256f
C3381 vdd.n1838 gnd 0.011256f
C3382 vdd.n1839 gnd 0.011256f
C3383 vdd.n1840 gnd 0.00906f
C3384 vdd.n1841 gnd 0.011256f
C3385 vdd.n1842 gnd 0.615415f
C3386 vdd.n1843 gnd 0.914496f
C3387 vdd.n1844 gnd 0.011256f
C3388 vdd.n1845 gnd 0.00906f
C3389 vdd.n1846 gnd 0.011256f
C3390 vdd.n1847 gnd 0.011256f
C3391 vdd.n1848 gnd 0.011256f
C3392 vdd.n1849 gnd 0.00906f
C3393 vdd.n1850 gnd 0.011256f
C3394 vdd.n1851 gnd 0.954757f
C3395 vdd.n1852 gnd 0.011256f
C3396 vdd.n1853 gnd 0.00906f
C3397 vdd.n1854 gnd 0.011256f
C3398 vdd.n1855 gnd 0.011256f
C3399 vdd.n1856 gnd 0.011256f
C3400 vdd.n1857 gnd 0.00906f
C3401 vdd.n1858 gnd 0.011256f
C3402 vdd.t130 gnd 0.575155f
C3403 vdd.n1859 gnd 0.799465f
C3404 vdd.n1860 gnd 0.011256f
C3405 vdd.n1861 gnd 0.00906f
C3406 vdd.n1862 gnd 0.011256f
C3407 vdd.n1863 gnd 0.011256f
C3408 vdd.n1864 gnd 0.011256f
C3409 vdd.n1865 gnd 0.00906f
C3410 vdd.n1866 gnd 0.011256f
C3411 vdd.n1867 gnd 0.603912f
C3412 vdd.n1868 gnd 0.011256f
C3413 vdd.n1869 gnd 0.00906f
C3414 vdd.n1870 gnd 0.011256f
C3415 vdd.n1871 gnd 0.011256f
C3416 vdd.n1872 gnd 0.011256f
C3417 vdd.n1873 gnd 0.00906f
C3418 vdd.n1874 gnd 0.011256f
C3419 vdd.n1875 gnd 0.787962f
C3420 vdd.n1876 gnd 0.741949f
C3421 vdd.n1877 gnd 0.011256f
C3422 vdd.n1878 gnd 0.00906f
C3423 vdd.n1879 gnd 0.011256f
C3424 vdd.n1880 gnd 0.011256f
C3425 vdd.n1881 gnd 0.011256f
C3426 vdd.n1882 gnd 0.00906f
C3427 vdd.n1883 gnd 0.011256f
C3428 vdd.n1884 gnd 0.937502f
C3429 vdd.n1885 gnd 0.011256f
C3430 vdd.n1886 gnd 0.00906f
C3431 vdd.n1887 gnd 0.011256f
C3432 vdd.n1888 gnd 0.011256f
C3433 vdd.n1889 gnd 0.027229f
C3434 vdd.n1890 gnd 0.011256f
C3435 vdd.n1891 gnd 0.011256f
C3436 vdd.n1892 gnd 0.00906f
C3437 vdd.n1893 gnd 0.011256f
C3438 vdd.n1894 gnd 0.695937f
C3439 vdd.n1895 gnd 1.15031f
C3440 vdd.n1896 gnd 0.011256f
C3441 vdd.n1897 gnd 0.00906f
C3442 vdd.n1898 gnd 0.011256f
C3443 vdd.n1899 gnd 0.011256f
C3444 vdd.n1900 gnd 0.00968f
C3445 vdd.n1901 gnd 0.00906f
C3446 vdd.n1903 gnd 0.011256f
C3447 vdd.n1905 gnd 0.00906f
C3448 vdd.n1906 gnd 0.011256f
C3449 vdd.n1907 gnd 0.00906f
C3450 vdd.n1909 gnd 0.011256f
C3451 vdd.n1910 gnd 0.00906f
C3452 vdd.n1911 gnd 0.011256f
C3453 vdd.n1912 gnd 0.011256f
C3454 vdd.n1913 gnd 0.011256f
C3455 vdd.n1914 gnd 0.011256f
C3456 vdd.n1915 gnd 0.011256f
C3457 vdd.n1916 gnd 0.00906f
C3458 vdd.n1918 gnd 0.011256f
C3459 vdd.n1919 gnd 0.011256f
C3460 vdd.n1920 gnd 0.011256f
C3461 vdd.n1921 gnd 0.011256f
C3462 vdd.n1922 gnd 0.011256f
C3463 vdd.n1923 gnd 0.00906f
C3464 vdd.n1925 gnd 0.011256f
C3465 vdd.n1926 gnd 0.011256f
C3466 vdd.n1927 gnd 0.011256f
C3467 vdd.n1928 gnd 0.011256f
C3468 vdd.n1929 gnd 0.007565f
C3469 vdd.t249 gnd 0.138478f
C3470 vdd.t248 gnd 0.147995f
C3471 vdd.t247 gnd 0.180851f
C3472 vdd.n1930 gnd 0.231825f
C3473 vdd.n1931 gnd 0.194775f
C3474 vdd.n1933 gnd 0.011256f
C3475 vdd.n1934 gnd 0.011256f
C3476 vdd.n1935 gnd 0.00906f
C3477 vdd.n1936 gnd 0.011256f
C3478 vdd.n1938 gnd 0.011256f
C3479 vdd.n1939 gnd 0.011256f
C3480 vdd.n1940 gnd 0.011256f
C3481 vdd.n1941 gnd 0.011256f
C3482 vdd.n1942 gnd 0.00906f
C3483 vdd.n1944 gnd 0.011256f
C3484 vdd.n1945 gnd 0.011256f
C3485 vdd.n1946 gnd 0.011256f
C3486 vdd.n1947 gnd 0.011256f
C3487 vdd.n1948 gnd 0.011256f
C3488 vdd.n1949 gnd 0.00906f
C3489 vdd.n1951 gnd 0.011256f
C3490 vdd.n1952 gnd 0.011256f
C3491 vdd.n1953 gnd 0.011256f
C3492 vdd.n1954 gnd 0.011256f
C3493 vdd.n1955 gnd 0.011256f
C3494 vdd.n1956 gnd 0.00906f
C3495 vdd.n1958 gnd 0.011256f
C3496 vdd.n1959 gnd 0.011256f
C3497 vdd.n1960 gnd 0.011256f
C3498 vdd.n1961 gnd 0.011256f
C3499 vdd.n1962 gnd 0.011256f
C3500 vdd.n1963 gnd 0.00906f
C3501 vdd.n1965 gnd 0.011256f
C3502 vdd.n1966 gnd 0.011256f
C3503 vdd.n1967 gnd 0.011256f
C3504 vdd.n1968 gnd 0.011256f
C3505 vdd.n1969 gnd 0.008969f
C3506 vdd.t236 gnd 0.138478f
C3507 vdd.t235 gnd 0.147995f
C3508 vdd.t234 gnd 0.180851f
C3509 vdd.n1970 gnd 0.231825f
C3510 vdd.n1971 gnd 0.194775f
C3511 vdd.n1973 gnd 0.011256f
C3512 vdd.n1974 gnd 0.011256f
C3513 vdd.n1975 gnd 0.00906f
C3514 vdd.n1976 gnd 0.011256f
C3515 vdd.n1978 gnd 0.011256f
C3516 vdd.n1979 gnd 0.011256f
C3517 vdd.n1980 gnd 0.011256f
C3518 vdd.n1981 gnd 0.011256f
C3519 vdd.n1982 gnd 0.00906f
C3520 vdd.n1984 gnd 0.011256f
C3521 vdd.n1985 gnd 0.011256f
C3522 vdd.n1986 gnd 0.011256f
C3523 vdd.n1987 gnd 0.011256f
C3524 vdd.n1988 gnd 0.011256f
C3525 vdd.n1989 gnd 0.00906f
C3526 vdd.n1991 gnd 0.011256f
C3527 vdd.n1992 gnd 0.011256f
C3528 vdd.n1993 gnd 0.011256f
C3529 vdd.n1994 gnd 0.011256f
C3530 vdd.n1995 gnd 0.011256f
C3531 vdd.n1996 gnd 0.011256f
C3532 vdd.n1997 gnd 0.00906f
C3533 vdd.n1999 gnd 0.011256f
C3534 vdd.n2001 gnd 0.011256f
C3535 vdd.n2002 gnd 0.00906f
C3536 vdd.n2003 gnd 0.00906f
C3537 vdd.n2004 gnd 0.011256f
C3538 vdd.n2006 gnd 0.011256f
C3539 vdd.n2007 gnd 0.00906f
C3540 vdd.n2008 gnd 0.00906f
C3541 vdd.n2009 gnd 0.011256f
C3542 vdd.n2011 gnd 0.011256f
C3543 vdd.n2012 gnd 0.011256f
C3544 vdd.n2013 gnd 0.00906f
C3545 vdd.n2014 gnd 0.00906f
C3546 vdd.n2015 gnd 0.00906f
C3547 vdd.n2016 gnd 0.011256f
C3548 vdd.n2018 gnd 0.011256f
C3549 vdd.n2019 gnd 0.011256f
C3550 vdd.n2020 gnd 0.00906f
C3551 vdd.n2021 gnd 0.00906f
C3552 vdd.n2022 gnd 0.00906f
C3553 vdd.n2023 gnd 0.011256f
C3554 vdd.n2025 gnd 0.011256f
C3555 vdd.n2026 gnd 0.011256f
C3556 vdd.n2027 gnd 0.00906f
C3557 vdd.n2028 gnd 0.00906f
C3558 vdd.n2029 gnd 0.00906f
C3559 vdd.n2030 gnd 0.011256f
C3560 vdd.n2032 gnd 0.011256f
C3561 vdd.n2033 gnd 0.011256f
C3562 vdd.n2034 gnd 0.00906f
C3563 vdd.n2035 gnd 0.011256f
C3564 vdd.n2036 gnd 0.011256f
C3565 vdd.n2037 gnd 0.011256f
C3566 vdd.n2038 gnd 0.018482f
C3567 vdd.n2039 gnd 0.006161f
C3568 vdd.n2040 gnd 0.00906f
C3569 vdd.n2041 gnd 0.011256f
C3570 vdd.n2043 gnd 0.011256f
C3571 vdd.n2044 gnd 0.011256f
C3572 vdd.n2045 gnd 0.00906f
C3573 vdd.n2046 gnd 0.00906f
C3574 vdd.n2047 gnd 0.00906f
C3575 vdd.n2048 gnd 0.011256f
C3576 vdd.n2050 gnd 0.011256f
C3577 vdd.n2051 gnd 0.011256f
C3578 vdd.n2052 gnd 0.00906f
C3579 vdd.n2053 gnd 0.00906f
C3580 vdd.n2054 gnd 0.00906f
C3581 vdd.n2055 gnd 0.011256f
C3582 vdd.n2057 gnd 0.011256f
C3583 vdd.n2058 gnd 0.011256f
C3584 vdd.n2059 gnd 0.00906f
C3585 vdd.n2060 gnd 0.00906f
C3586 vdd.n2061 gnd 0.00906f
C3587 vdd.n2062 gnd 0.011256f
C3588 vdd.n2064 gnd 0.011256f
C3589 vdd.n2065 gnd 0.011256f
C3590 vdd.n2066 gnd 0.00906f
C3591 vdd.n2067 gnd 0.00906f
C3592 vdd.n2068 gnd 0.00906f
C3593 vdd.n2069 gnd 0.011256f
C3594 vdd.n2071 gnd 0.011256f
C3595 vdd.n2072 gnd 0.011256f
C3596 vdd.n2073 gnd 0.00906f
C3597 vdd.n2074 gnd 0.011256f
C3598 vdd.n2075 gnd 0.011256f
C3599 vdd.n2076 gnd 0.011256f
C3600 vdd.n2077 gnd 0.018482f
C3601 vdd.n2078 gnd 0.007565f
C3602 vdd.n2079 gnd 0.00906f
C3603 vdd.n2080 gnd 0.011256f
C3604 vdd.n2082 gnd 0.011256f
C3605 vdd.n2083 gnd 0.011256f
C3606 vdd.n2084 gnd 0.00906f
C3607 vdd.n2085 gnd 0.00906f
C3608 vdd.n2086 gnd 0.00906f
C3609 vdd.n2087 gnd 0.011256f
C3610 vdd.n2089 gnd 0.011256f
C3611 vdd.n2090 gnd 0.011256f
C3612 vdd.n2091 gnd 0.00906f
C3613 vdd.n2092 gnd 0.00906f
C3614 vdd.n2093 gnd 0.00906f
C3615 vdd.n2094 gnd 0.011256f
C3616 vdd.n2096 gnd 0.011256f
C3617 vdd.n2097 gnd 0.011256f
C3618 vdd.n2099 gnd 0.011256f
C3619 vdd.n2100 gnd 0.00906f
C3620 vdd.n2101 gnd 0.007204f
C3621 vdd.n2102 gnd 0.007654f
C3622 vdd.n2103 gnd 0.007654f
C3623 vdd.n2104 gnd 0.007654f
C3624 vdd.n2105 gnd 0.007654f
C3625 vdd.n2106 gnd 0.007654f
C3626 vdd.n2107 gnd 0.007654f
C3627 vdd.n2108 gnd 0.007654f
C3628 vdd.n2109 gnd 0.007654f
C3629 vdd.n2111 gnd 0.007654f
C3630 vdd.n2112 gnd 0.007654f
C3631 vdd.n2113 gnd 0.007654f
C3632 vdd.n2114 gnd 0.007654f
C3633 vdd.n2115 gnd 0.007654f
C3634 vdd.n2117 gnd 0.007654f
C3635 vdd.n2119 gnd 0.007654f
C3636 vdd.n2120 gnd 0.007654f
C3637 vdd.n2121 gnd 0.007654f
C3638 vdd.n2122 gnd 0.007654f
C3639 vdd.n2123 gnd 0.007654f
C3640 vdd.n2125 gnd 0.007654f
C3641 vdd.n2127 gnd 0.007654f
C3642 vdd.n2128 gnd 0.007654f
C3643 vdd.n2129 gnd 0.007654f
C3644 vdd.n2130 gnd 0.007654f
C3645 vdd.n2131 gnd 0.007654f
C3646 vdd.n2133 gnd 0.007654f
C3647 vdd.n2135 gnd 0.007654f
C3648 vdd.n2136 gnd 0.007654f
C3649 vdd.n2137 gnd 0.007654f
C3650 vdd.n2138 gnd 0.007654f
C3651 vdd.n2139 gnd 0.007654f
C3652 vdd.n2141 gnd 0.007654f
C3653 vdd.n2142 gnd 0.007654f
C3654 vdd.n2143 gnd 0.007654f
C3655 vdd.n2144 gnd 0.007654f
C3656 vdd.n2145 gnd 0.007654f
C3657 vdd.n2146 gnd 0.007654f
C3658 vdd.n2147 gnd 0.007654f
C3659 vdd.n2148 gnd 0.007654f
C3660 vdd.n2149 gnd 0.005572f
C3661 vdd.n2150 gnd 0.007654f
C3662 vdd.t213 gnd 0.3093f
C3663 vdd.t214 gnd 0.316607f
C3664 vdd.t211 gnd 0.201923f
C3665 vdd.n2151 gnd 0.109128f
C3666 vdd.n2152 gnd 0.061901f
C3667 vdd.n2153 gnd 0.010939f
C3668 vdd.n2154 gnd 0.007654f
C3669 vdd.n2155 gnd 0.007654f
C3670 vdd.n2156 gnd 0.465875f
C3671 vdd.n2157 gnd 0.007654f
C3672 vdd.n2158 gnd 0.007654f
C3673 vdd.n2159 gnd 0.007654f
C3674 vdd.n2160 gnd 0.007654f
C3675 vdd.n2161 gnd 0.007654f
C3676 vdd.n2162 gnd 0.007654f
C3677 vdd.n2163 gnd 0.007654f
C3678 vdd.n2164 gnd 0.007654f
C3679 vdd.n2165 gnd 0.007654f
C3680 vdd.n2166 gnd 0.007654f
C3681 vdd.n2167 gnd 0.007654f
C3682 vdd.n2168 gnd 0.007654f
C3683 vdd.n2169 gnd 0.007654f
C3684 vdd.n2170 gnd 0.007654f
C3685 vdd.n2171 gnd 0.007654f
C3686 vdd.n2172 gnd 0.007654f
C3687 vdd.n2173 gnd 0.007654f
C3688 vdd.n2174 gnd 0.007654f
C3689 vdd.n2175 gnd 0.007654f
C3690 vdd.n2176 gnd 0.007654f
C3691 vdd.t266 gnd 0.3093f
C3692 vdd.t267 gnd 0.316607f
C3693 vdd.t265 gnd 0.201923f
C3694 vdd.n2177 gnd 0.109128f
C3695 vdd.n2178 gnd 0.061901f
C3696 vdd.n2179 gnd 0.007654f
C3697 vdd.n2180 gnd 0.007654f
C3698 vdd.n2181 gnd 0.007654f
C3699 vdd.n2182 gnd 0.007654f
C3700 vdd.n2183 gnd 0.007654f
C3701 vdd.n2184 gnd 0.007654f
C3702 vdd.n2186 gnd 0.007654f
C3703 vdd.n2187 gnd 0.007654f
C3704 vdd.n2188 gnd 0.007654f
C3705 vdd.n2189 gnd 0.007654f
C3706 vdd.n2191 gnd 0.007654f
C3707 vdd.n2193 gnd 0.007654f
C3708 vdd.n2194 gnd 0.007654f
C3709 vdd.n2195 gnd 0.007654f
C3710 vdd.n2196 gnd 0.007654f
C3711 vdd.n2197 gnd 0.007654f
C3712 vdd.n2199 gnd 0.007654f
C3713 vdd.n2201 gnd 0.007654f
C3714 vdd.n2202 gnd 0.007654f
C3715 vdd.n2203 gnd 0.007654f
C3716 vdd.n2204 gnd 0.007654f
C3717 vdd.n2205 gnd 0.007654f
C3718 vdd.n2207 gnd 0.007654f
C3719 vdd.n2209 gnd 0.007654f
C3720 vdd.n2210 gnd 0.007654f
C3721 vdd.n2211 gnd 0.005572f
C3722 vdd.n2212 gnd 0.010939f
C3723 vdd.n2213 gnd 0.005909f
C3724 vdd.n2214 gnd 0.007654f
C3725 vdd.n2216 gnd 0.007654f
C3726 vdd.n2217 gnd 0.018162f
C3727 vdd.n2218 gnd 0.018162f
C3728 vdd.n2219 gnd 0.016957f
C3729 vdd.n2220 gnd 0.007654f
C3730 vdd.n2221 gnd 0.007654f
C3731 vdd.n2222 gnd 0.007654f
C3732 vdd.n2223 gnd 0.007654f
C3733 vdd.n2224 gnd 0.007654f
C3734 vdd.n2225 gnd 0.007654f
C3735 vdd.n2226 gnd 0.007654f
C3736 vdd.n2227 gnd 0.007654f
C3737 vdd.n2228 gnd 0.007654f
C3738 vdd.n2229 gnd 0.007654f
C3739 vdd.n2230 gnd 0.007654f
C3740 vdd.n2231 gnd 0.007654f
C3741 vdd.n2232 gnd 0.007654f
C3742 vdd.n2233 gnd 0.007654f
C3743 vdd.n2234 gnd 0.007654f
C3744 vdd.n2235 gnd 0.007654f
C3745 vdd.n2236 gnd 0.007654f
C3746 vdd.n2237 gnd 0.007654f
C3747 vdd.n2238 gnd 0.007654f
C3748 vdd.n2239 gnd 0.007654f
C3749 vdd.n2240 gnd 0.007654f
C3750 vdd.n2241 gnd 0.007654f
C3751 vdd.n2242 gnd 0.007654f
C3752 vdd.n2243 gnd 0.007654f
C3753 vdd.n2244 gnd 0.007654f
C3754 vdd.n2245 gnd 0.007654f
C3755 vdd.n2246 gnd 0.007654f
C3756 vdd.n2247 gnd 0.007654f
C3757 vdd.n2248 gnd 0.007654f
C3758 vdd.n2249 gnd 0.007654f
C3759 vdd.n2250 gnd 0.007654f
C3760 vdd.n2251 gnd 0.007654f
C3761 vdd.n2252 gnd 0.007654f
C3762 vdd.n2253 gnd 0.007654f
C3763 vdd.n2254 gnd 0.007654f
C3764 vdd.n2255 gnd 0.007654f
C3765 vdd.n2256 gnd 0.007654f
C3766 vdd.n2257 gnd 0.247316f
C3767 vdd.n2258 gnd 0.007654f
C3768 vdd.n2259 gnd 0.007654f
C3769 vdd.n2260 gnd 0.007654f
C3770 vdd.n2261 gnd 0.007654f
C3771 vdd.n2262 gnd 0.007654f
C3772 vdd.n2263 gnd 0.007654f
C3773 vdd.n2264 gnd 0.007654f
C3774 vdd.n2265 gnd 0.007654f
C3775 vdd.n2266 gnd 0.007654f
C3776 vdd.n2267 gnd 0.007654f
C3777 vdd.n2268 gnd 0.007654f
C3778 vdd.n2269 gnd 0.007654f
C3779 vdd.n2270 gnd 0.007654f
C3780 vdd.n2271 gnd 0.007654f
C3781 vdd.n2272 gnd 0.007654f
C3782 vdd.n2273 gnd 0.007654f
C3783 vdd.n2274 gnd 0.007654f
C3784 vdd.n2275 gnd 0.007654f
C3785 vdd.n2276 gnd 0.007654f
C3786 vdd.n2277 gnd 0.007654f
C3787 vdd.n2278 gnd 0.016957f
C3788 vdd.n2280 gnd 0.018162f
C3789 vdd.n2281 gnd 0.018162f
C3790 vdd.n2282 gnd 0.007654f
C3791 vdd.n2283 gnd 0.005909f
C3792 vdd.n2284 gnd 0.007654f
C3793 vdd.n2286 gnd 0.007654f
C3794 vdd.n2288 gnd 0.007654f
C3795 vdd.n2289 gnd 0.007654f
C3796 vdd.n2290 gnd 0.007654f
C3797 vdd.n2291 gnd 0.007654f
C3798 vdd.n2292 gnd 0.007654f
C3799 vdd.n2294 gnd 0.007654f
C3800 vdd.n2296 gnd 0.007654f
C3801 vdd.n2297 gnd 0.007654f
C3802 vdd.n2298 gnd 0.007654f
C3803 vdd.n2299 gnd 0.007654f
C3804 vdd.n2300 gnd 0.007654f
C3805 vdd.n2302 gnd 0.007654f
C3806 vdd.n2304 gnd 0.007654f
C3807 vdd.n2305 gnd 0.007654f
C3808 vdd.n2306 gnd 0.007654f
C3809 vdd.n2307 gnd 0.007654f
C3810 vdd.n2308 gnd 0.007654f
C3811 vdd.n2310 gnd 0.007654f
C3812 vdd.n2312 gnd 0.007654f
C3813 vdd.n2313 gnd 0.007654f
C3814 vdd.n2314 gnd 0.02283f
C3815 vdd.n2315 gnd 0.676794f
C3816 vdd.n2317 gnd 0.00906f
C3817 vdd.n2318 gnd 0.00906f
C3818 vdd.n2319 gnd 0.011256f
C3819 vdd.n2321 gnd 0.011256f
C3820 vdd.n2322 gnd 0.011256f
C3821 vdd.n2323 gnd 0.00906f
C3822 vdd.n2324 gnd 0.00752f
C3823 vdd.n2325 gnd 0.027813f
C3824 vdd.n2326 gnd 0.027229f
C3825 vdd.n2327 gnd 0.00752f
C3826 vdd.n2328 gnd 0.027229f
C3827 vdd.n2329 gnd 1.58168f
C3828 vdd.n2330 gnd 0.027229f
C3829 vdd.n2331 gnd 0.027813f
C3830 vdd.n2332 gnd 0.004303f
C3831 vdd.t225 gnd 0.138478f
C3832 vdd.t224 gnd 0.147995f
C3833 vdd.t222 gnd 0.180851f
C3834 vdd.n2333 gnd 0.231825f
C3835 vdd.n2334 gnd 0.194775f
C3836 vdd.n2335 gnd 0.013952f
C3837 vdd.n2336 gnd 0.004756f
C3838 vdd.n2337 gnd 0.00968f
C3839 vdd.n2338 gnd 0.676794f
C3840 vdd.n2339 gnd 0.02283f
C3841 vdd.n2340 gnd 0.007654f
C3842 vdd.n2341 gnd 0.007654f
C3843 vdd.n2342 gnd 0.007654f
C3844 vdd.n2344 gnd 0.007654f
C3845 vdd.n2346 gnd 0.007654f
C3846 vdd.n2347 gnd 0.007654f
C3847 vdd.n2348 gnd 0.007654f
C3848 vdd.n2349 gnd 0.007654f
C3849 vdd.n2350 gnd 0.007654f
C3850 vdd.n2352 gnd 0.007654f
C3851 vdd.n2354 gnd 0.007654f
C3852 vdd.n2355 gnd 0.007654f
C3853 vdd.n2356 gnd 0.007654f
C3854 vdd.n2357 gnd 0.007654f
C3855 vdd.n2358 gnd 0.007654f
C3856 vdd.n2360 gnd 0.007654f
C3857 vdd.n2362 gnd 0.007654f
C3858 vdd.n2363 gnd 0.007654f
C3859 vdd.n2364 gnd 0.007654f
C3860 vdd.n2365 gnd 0.007654f
C3861 vdd.n2366 gnd 0.007654f
C3862 vdd.n2368 gnd 0.007654f
C3863 vdd.n2370 gnd 0.007654f
C3864 vdd.n2371 gnd 0.007654f
C3865 vdd.n2372 gnd 0.018162f
C3866 vdd.n2373 gnd 0.016957f
C3867 vdd.n2374 gnd 0.016957f
C3868 vdd.n2375 gnd 1.1273f
C3869 vdd.n2376 gnd 0.016957f
C3870 vdd.n2377 gnd 0.016957f
C3871 vdd.n2378 gnd 0.007654f
C3872 vdd.n2379 gnd 0.007654f
C3873 vdd.n2380 gnd 0.007654f
C3874 vdd.n2381 gnd 0.488881f
C3875 vdd.n2382 gnd 0.007654f
C3876 vdd.n2383 gnd 0.007654f
C3877 vdd.n2384 gnd 0.007654f
C3878 vdd.n2385 gnd 0.007654f
C3879 vdd.n2386 gnd 0.007654f
C3880 vdd.n2387 gnd 0.78221f
C3881 vdd.n2388 gnd 0.007654f
C3882 vdd.n2389 gnd 0.007654f
C3883 vdd.n2390 gnd 0.007654f
C3884 vdd.n2391 gnd 0.007654f
C3885 vdd.n2392 gnd 0.007654f
C3886 vdd.n2393 gnd 0.78221f
C3887 vdd.n2394 gnd 0.007654f
C3888 vdd.n2395 gnd 0.007654f
C3889 vdd.n2396 gnd 0.006754f
C3890 vdd.n2397 gnd 0.022173f
C3891 vdd.n2398 gnd 0.004728f
C3892 vdd.n2399 gnd 0.007654f
C3893 vdd.n2400 gnd 0.431366f
C3894 vdd.n2401 gnd 0.007654f
C3895 vdd.n2402 gnd 0.007654f
C3896 vdd.n2403 gnd 0.007654f
C3897 vdd.n2404 gnd 0.007654f
C3898 vdd.n2405 gnd 0.007654f
C3899 vdd.n2406 gnd 0.523391f
C3900 vdd.n2407 gnd 0.007654f
C3901 vdd.n2408 gnd 0.007654f
C3902 vdd.n2409 gnd 0.007654f
C3903 vdd.n2410 gnd 0.007654f
C3904 vdd.n2411 gnd 0.007654f
C3905 vdd.n2412 gnd 0.695937f
C3906 vdd.n2413 gnd 0.007654f
C3907 vdd.n2414 gnd 0.007654f
C3908 vdd.n2415 gnd 0.007654f
C3909 vdd.n2416 gnd 0.007654f
C3910 vdd.n2417 gnd 0.007654f
C3911 vdd.n2418 gnd 0.621167f
C3912 vdd.n2419 gnd 0.007654f
C3913 vdd.n2420 gnd 0.007654f
C3914 vdd.n2421 gnd 0.007654f
C3915 vdd.n2422 gnd 0.007654f
C3916 vdd.n2423 gnd 0.007654f
C3917 vdd.n2424 gnd 0.448621f
C3918 vdd.n2425 gnd 0.007654f
C3919 vdd.n2426 gnd 0.007654f
C3920 vdd.n2427 gnd 0.007654f
C3921 vdd.n2428 gnd 0.007654f
C3922 vdd.n2429 gnd 0.007654f
C3923 vdd.n2430 gnd 0.247316f
C3924 vdd.n2431 gnd 0.007654f
C3925 vdd.n2432 gnd 0.007654f
C3926 vdd.n2433 gnd 0.007654f
C3927 vdd.n2434 gnd 0.007654f
C3928 vdd.n2435 gnd 0.007654f
C3929 vdd.n2436 gnd 0.431366f
C3930 vdd.n2437 gnd 0.007654f
C3931 vdd.n2438 gnd 0.007654f
C3932 vdd.n2439 gnd 0.007654f
C3933 vdd.n2440 gnd 0.007654f
C3934 vdd.n2441 gnd 0.007654f
C3935 vdd.n2442 gnd 0.78221f
C3936 vdd.n2443 gnd 0.007654f
C3937 vdd.n2444 gnd 0.007654f
C3938 vdd.n2445 gnd 0.007654f
C3939 vdd.n2446 gnd 0.007654f
C3940 vdd.n2447 gnd 0.007654f
C3941 vdd.n2448 gnd 0.007654f
C3942 vdd.n2449 gnd 0.007654f
C3943 vdd.n2450 gnd 0.609664f
C3944 vdd.n2451 gnd 0.007654f
C3945 vdd.n2452 gnd 0.007654f
C3946 vdd.n2453 gnd 0.007654f
C3947 vdd.n2454 gnd 0.007654f
C3948 vdd.n2455 gnd 0.007654f
C3949 vdd.n2456 gnd 0.007654f
C3950 vdd.n2457 gnd 0.488881f
C3951 vdd.n2458 gnd 0.007654f
C3952 vdd.n2459 gnd 0.007654f
C3953 vdd.n2460 gnd 0.007654f
C3954 vdd.n2461 gnd 0.017889f
C3955 vdd.n2462 gnd 0.01723f
C3956 vdd.n2463 gnd 0.007654f
C3957 vdd.n2464 gnd 0.007654f
C3958 vdd.n2465 gnd 0.005909f
C3959 vdd.n2466 gnd 0.007654f
C3960 vdd.n2467 gnd 0.007654f
C3961 vdd.n2468 gnd 0.005572f
C3962 vdd.n2469 gnd 0.007654f
C3963 vdd.n2470 gnd 0.007654f
C3964 vdd.n2471 gnd 0.007654f
C3965 vdd.n2472 gnd 0.007654f
C3966 vdd.n2473 gnd 0.007654f
C3967 vdd.n2474 gnd 0.007654f
C3968 vdd.n2475 gnd 0.007654f
C3969 vdd.n2476 gnd 0.007654f
C3970 vdd.n2477 gnd 0.007654f
C3971 vdd.n2478 gnd 0.007654f
C3972 vdd.n2479 gnd 0.007654f
C3973 vdd.n2480 gnd 0.007654f
C3974 vdd.n2481 gnd 0.007654f
C3975 vdd.n2482 gnd 0.007654f
C3976 vdd.n2483 gnd 0.007654f
C3977 vdd.n2484 gnd 0.007654f
C3978 vdd.n2485 gnd 0.007654f
C3979 vdd.n2486 gnd 0.007654f
C3980 vdd.n2487 gnd 0.007654f
C3981 vdd.n2488 gnd 0.007654f
C3982 vdd.n2489 gnd 0.007654f
C3983 vdd.n2490 gnd 0.007654f
C3984 vdd.n2491 gnd 0.007654f
C3985 vdd.n2492 gnd 0.007654f
C3986 vdd.n2493 gnd 0.007654f
C3987 vdd.n2494 gnd 0.007654f
C3988 vdd.n2495 gnd 0.007654f
C3989 vdd.n2496 gnd 0.007654f
C3990 vdd.n2497 gnd 0.007654f
C3991 vdd.n2498 gnd 0.007654f
C3992 vdd.n2499 gnd 0.007654f
C3993 vdd.n2500 gnd 0.007654f
C3994 vdd.n2501 gnd 0.007654f
C3995 vdd.n2502 gnd 0.007654f
C3996 vdd.n2503 gnd 0.007654f
C3997 vdd.n2504 gnd 0.007654f
C3998 vdd.n2505 gnd 0.007654f
C3999 vdd.n2506 gnd 0.007654f
C4000 vdd.n2507 gnd 0.007654f
C4001 vdd.n2508 gnd 0.007654f
C4002 vdd.n2509 gnd 0.007654f
C4003 vdd.n2510 gnd 0.007654f
C4004 vdd.n2511 gnd 0.007654f
C4005 vdd.n2512 gnd 0.007654f
C4006 vdd.n2513 gnd 0.007654f
C4007 vdd.n2514 gnd 0.007654f
C4008 vdd.n2515 gnd 0.007654f
C4009 vdd.n2516 gnd 0.007654f
C4010 vdd.n2517 gnd 0.007654f
C4011 vdd.n2518 gnd 0.007654f
C4012 vdd.n2519 gnd 0.007654f
C4013 vdd.n2520 gnd 0.007654f
C4014 vdd.n2521 gnd 0.007654f
C4015 vdd.n2522 gnd 0.007654f
C4016 vdd.n2523 gnd 0.007654f
C4017 vdd.n2524 gnd 0.007654f
C4018 vdd.n2525 gnd 0.007654f
C4019 vdd.n2526 gnd 0.007654f
C4020 vdd.n2527 gnd 0.007654f
C4021 vdd.n2528 gnd 0.007654f
C4022 vdd.n2529 gnd 0.018162f
C4023 vdd.n2530 gnd 0.016957f
C4024 vdd.n2531 gnd 0.016957f
C4025 vdd.n2532 gnd 0.954757f
C4026 vdd.n2533 gnd 0.016957f
C4027 vdd.n2534 gnd 0.018162f
C4028 vdd.n2535 gnd 0.01723f
C4029 vdd.n2536 gnd 0.007654f
C4030 vdd.n2537 gnd 0.007654f
C4031 vdd.n2538 gnd 0.007654f
C4032 vdd.n2539 gnd 0.005909f
C4033 vdd.n2540 gnd 0.010939f
C4034 vdd.n2541 gnd 0.005572f
C4035 vdd.n2542 gnd 0.007654f
C4036 vdd.n2543 gnd 0.007654f
C4037 vdd.n2544 gnd 0.007654f
C4038 vdd.n2545 gnd 0.007654f
C4039 vdd.n2546 gnd 0.007654f
C4040 vdd.n2547 gnd 0.007654f
C4041 vdd.n2548 gnd 0.007654f
C4042 vdd.n2549 gnd 0.007654f
C4043 vdd.n2550 gnd 0.007654f
C4044 vdd.n2551 gnd 0.007654f
C4045 vdd.n2552 gnd 0.007654f
C4046 vdd.n2553 gnd 0.007654f
C4047 vdd.n2554 gnd 0.007654f
C4048 vdd.n2555 gnd 0.007654f
C4049 vdd.n2556 gnd 0.007654f
C4050 vdd.n2557 gnd 0.007654f
C4051 vdd.n2558 gnd 0.007654f
C4052 vdd.n2559 gnd 0.007654f
C4053 vdd.n2560 gnd 0.007654f
C4054 vdd.n2561 gnd 0.007654f
C4055 vdd.n2562 gnd 0.007654f
C4056 vdd.n2563 gnd 0.007654f
C4057 vdd.n2564 gnd 0.007654f
C4058 vdd.n2565 gnd 0.007654f
C4059 vdd.n2566 gnd 0.007654f
C4060 vdd.n2567 gnd 0.007654f
C4061 vdd.n2568 gnd 0.007654f
C4062 vdd.n2569 gnd 0.007654f
C4063 vdd.n2570 gnd 0.007654f
C4064 vdd.n2571 gnd 0.007654f
C4065 vdd.n2572 gnd 0.007654f
C4066 vdd.n2573 gnd 0.007654f
C4067 vdd.n2574 gnd 0.007654f
C4068 vdd.n2575 gnd 0.007654f
C4069 vdd.n2576 gnd 0.007654f
C4070 vdd.n2577 gnd 0.007654f
C4071 vdd.n2578 gnd 0.007654f
C4072 vdd.n2579 gnd 0.007654f
C4073 vdd.n2580 gnd 0.007654f
C4074 vdd.n2581 gnd 0.007654f
C4075 vdd.n2582 gnd 0.007654f
C4076 vdd.n2583 gnd 0.007654f
C4077 vdd.n2584 gnd 0.007654f
C4078 vdd.n2585 gnd 0.007654f
C4079 vdd.n2586 gnd 0.007654f
C4080 vdd.n2587 gnd 0.007654f
C4081 vdd.n2588 gnd 0.007654f
C4082 vdd.n2589 gnd 0.007654f
C4083 vdd.n2590 gnd 0.007654f
C4084 vdd.n2591 gnd 0.007654f
C4085 vdd.n2592 gnd 0.007654f
C4086 vdd.n2593 gnd 0.007654f
C4087 vdd.n2594 gnd 0.007654f
C4088 vdd.n2595 gnd 0.007654f
C4089 vdd.n2596 gnd 0.007654f
C4090 vdd.n2597 gnd 0.007654f
C4091 vdd.n2598 gnd 0.007654f
C4092 vdd.n2599 gnd 0.007654f
C4093 vdd.n2600 gnd 0.007654f
C4094 vdd.n2601 gnd 0.007654f
C4095 vdd.n2602 gnd 0.018162f
C4096 vdd.n2603 gnd 0.018162f
C4097 vdd.n2604 gnd 0.954757f
C4098 vdd.t196 gnd 3.39341f
C4099 vdd.t294 gnd 3.39341f
C4100 vdd.n2637 gnd 0.018162f
C4101 vdd.n2638 gnd 0.007654f
C4102 vdd.t260 gnd 0.3093f
C4103 vdd.t261 gnd 0.316607f
C4104 vdd.t258 gnd 0.201923f
C4105 vdd.n2639 gnd 0.109128f
C4106 vdd.n2640 gnd 0.061901f
C4107 vdd.n2641 gnd 0.007654f
C4108 vdd.t273 gnd 0.3093f
C4109 vdd.t274 gnd 0.316607f
C4110 vdd.t272 gnd 0.201923f
C4111 vdd.n2642 gnd 0.109128f
C4112 vdd.n2643 gnd 0.061901f
C4113 vdd.n2644 gnd 0.010939f
C4114 vdd.n2645 gnd 0.007654f
C4115 vdd.n2646 gnd 0.007654f
C4116 vdd.n2647 gnd 0.007654f
C4117 vdd.n2648 gnd 0.007654f
C4118 vdd.n2649 gnd 0.007654f
C4119 vdd.n2650 gnd 0.007654f
C4120 vdd.n2651 gnd 0.007654f
C4121 vdd.n2652 gnd 0.007654f
C4122 vdd.n2653 gnd 0.007654f
C4123 vdd.n2654 gnd 0.007654f
C4124 vdd.n2655 gnd 0.007654f
C4125 vdd.n2656 gnd 0.007654f
C4126 vdd.n2657 gnd 0.007654f
C4127 vdd.n2658 gnd 0.007654f
C4128 vdd.n2659 gnd 0.007654f
C4129 vdd.n2660 gnd 0.007654f
C4130 vdd.n2661 gnd 0.007654f
C4131 vdd.n2662 gnd 0.007654f
C4132 vdd.n2663 gnd 0.007654f
C4133 vdd.n2664 gnd 0.007654f
C4134 vdd.n2665 gnd 0.007654f
C4135 vdd.n2666 gnd 0.007654f
C4136 vdd.n2667 gnd 0.007654f
C4137 vdd.n2668 gnd 0.007654f
C4138 vdd.n2669 gnd 0.007654f
C4139 vdd.n2670 gnd 0.007654f
C4140 vdd.n2671 gnd 0.007654f
C4141 vdd.n2672 gnd 0.007654f
C4142 vdd.n2673 gnd 0.007654f
C4143 vdd.n2674 gnd 0.007654f
C4144 vdd.n2675 gnd 0.007654f
C4145 vdd.n2676 gnd 0.007654f
C4146 vdd.n2677 gnd 0.007654f
C4147 vdd.n2678 gnd 0.007654f
C4148 vdd.n2679 gnd 0.007654f
C4149 vdd.n2680 gnd 0.007654f
C4150 vdd.n2681 gnd 0.007654f
C4151 vdd.n2682 gnd 0.007654f
C4152 vdd.n2683 gnd 0.007654f
C4153 vdd.n2684 gnd 0.007654f
C4154 vdd.n2685 gnd 0.007654f
C4155 vdd.n2686 gnd 0.007654f
C4156 vdd.n2687 gnd 0.007654f
C4157 vdd.n2688 gnd 0.007654f
C4158 vdd.n2689 gnd 0.007654f
C4159 vdd.n2690 gnd 0.007654f
C4160 vdd.n2691 gnd 0.007654f
C4161 vdd.n2692 gnd 0.007654f
C4162 vdd.n2693 gnd 0.007654f
C4163 vdd.n2694 gnd 0.007654f
C4164 vdd.n2695 gnd 0.007654f
C4165 vdd.n2696 gnd 0.007654f
C4166 vdd.n2697 gnd 0.007654f
C4167 vdd.n2698 gnd 0.007654f
C4168 vdd.n2699 gnd 0.007654f
C4169 vdd.n2700 gnd 0.007654f
C4170 vdd.n2701 gnd 0.005572f
C4171 vdd.n2702 gnd 0.007654f
C4172 vdd.n2703 gnd 0.007654f
C4173 vdd.n2704 gnd 0.005909f
C4174 vdd.n2705 gnd 0.007654f
C4175 vdd.n2706 gnd 0.007654f
C4176 vdd.n2707 gnd 0.018162f
C4177 vdd.n2708 gnd 0.016957f
C4178 vdd.n2709 gnd 0.007654f
C4179 vdd.n2710 gnd 0.007654f
C4180 vdd.n2711 gnd 0.007654f
C4181 vdd.n2712 gnd 0.007654f
C4182 vdd.n2713 gnd 0.007654f
C4183 vdd.n2714 gnd 0.007654f
C4184 vdd.n2715 gnd 0.007654f
C4185 vdd.n2716 gnd 0.007654f
C4186 vdd.n2717 gnd 0.007654f
C4187 vdd.n2718 gnd 0.007654f
C4188 vdd.n2719 gnd 0.007654f
C4189 vdd.n2720 gnd 0.007654f
C4190 vdd.n2721 gnd 0.007654f
C4191 vdd.n2722 gnd 0.007654f
C4192 vdd.n2723 gnd 0.007654f
C4193 vdd.n2724 gnd 0.007654f
C4194 vdd.n2725 gnd 0.007654f
C4195 vdd.n2726 gnd 0.007654f
C4196 vdd.n2727 gnd 0.007654f
C4197 vdd.n2728 gnd 0.007654f
C4198 vdd.n2729 gnd 0.007654f
C4199 vdd.n2730 gnd 0.007654f
C4200 vdd.n2731 gnd 0.007654f
C4201 vdd.n2732 gnd 0.007654f
C4202 vdd.n2733 gnd 0.007654f
C4203 vdd.n2734 gnd 0.007654f
C4204 vdd.n2735 gnd 0.007654f
C4205 vdd.n2736 gnd 0.007654f
C4206 vdd.n2737 gnd 0.007654f
C4207 vdd.n2738 gnd 0.007654f
C4208 vdd.n2739 gnd 0.007654f
C4209 vdd.n2740 gnd 0.007654f
C4210 vdd.n2741 gnd 0.007654f
C4211 vdd.n2742 gnd 0.007654f
C4212 vdd.n2743 gnd 0.007654f
C4213 vdd.n2744 gnd 0.007654f
C4214 vdd.n2745 gnd 0.007654f
C4215 vdd.n2746 gnd 0.007654f
C4216 vdd.n2747 gnd 0.007654f
C4217 vdd.n2748 gnd 0.007654f
C4218 vdd.n2749 gnd 0.007654f
C4219 vdd.n2750 gnd 0.007654f
C4220 vdd.n2751 gnd 0.007654f
C4221 vdd.n2752 gnd 0.007654f
C4222 vdd.n2753 gnd 0.007654f
C4223 vdd.n2754 gnd 0.007654f
C4224 vdd.n2755 gnd 0.007654f
C4225 vdd.n2756 gnd 0.007654f
C4226 vdd.n2757 gnd 0.007654f
C4227 vdd.n2758 gnd 0.007654f
C4228 vdd.n2759 gnd 0.007654f
C4229 vdd.n2760 gnd 0.247316f
C4230 vdd.n2761 gnd 0.007654f
C4231 vdd.n2762 gnd 0.007654f
C4232 vdd.n2763 gnd 0.007654f
C4233 vdd.n2764 gnd 0.007654f
C4234 vdd.n2765 gnd 0.007654f
C4235 vdd.n2766 gnd 0.007654f
C4236 vdd.n2767 gnd 0.007654f
C4237 vdd.n2768 gnd 0.007654f
C4238 vdd.n2769 gnd 0.007654f
C4239 vdd.n2770 gnd 0.007654f
C4240 vdd.n2771 gnd 0.007654f
C4241 vdd.n2772 gnd 0.007654f
C4242 vdd.n2773 gnd 0.007654f
C4243 vdd.n2774 gnd 0.007654f
C4244 vdd.n2775 gnd 0.007654f
C4245 vdd.n2776 gnd 0.007654f
C4246 vdd.n2777 gnd 0.007654f
C4247 vdd.n2778 gnd 0.007654f
C4248 vdd.n2779 gnd 0.007654f
C4249 vdd.n2780 gnd 0.007654f
C4250 vdd.n2781 gnd 0.465875f
C4251 vdd.n2782 gnd 0.007654f
C4252 vdd.n2783 gnd 0.007654f
C4253 vdd.n2784 gnd 0.007654f
C4254 vdd.n2785 gnd 0.007654f
C4255 vdd.n2786 gnd 0.007654f
C4256 vdd.n2787 gnd 0.016957f
C4257 vdd.n2788 gnd 0.018162f
C4258 vdd.n2789 gnd 0.018162f
C4259 vdd.n2790 gnd 0.007654f
C4260 vdd.n2791 gnd 0.007654f
C4261 vdd.n2792 gnd 0.007654f
C4262 vdd.n2793 gnd 0.005909f
C4263 vdd.n2794 gnd 0.010939f
C4264 vdd.n2795 gnd 0.005572f
C4265 vdd.n2796 gnd 0.007654f
C4266 vdd.n2797 gnd 0.007654f
C4267 vdd.n2798 gnd 0.007654f
C4268 vdd.n2799 gnd 0.007654f
C4269 vdd.n2800 gnd 0.007654f
C4270 vdd.n2801 gnd 0.007654f
C4271 vdd.n2802 gnd 0.007654f
C4272 vdd.n2803 gnd 0.007654f
C4273 vdd.n2804 gnd 0.007654f
C4274 vdd.n2805 gnd 0.007654f
C4275 vdd.n2806 gnd 0.007654f
C4276 vdd.n2807 gnd 0.007654f
C4277 vdd.n2808 gnd 0.007654f
C4278 vdd.n2809 gnd 0.007654f
C4279 vdd.n2810 gnd 0.007654f
C4280 vdd.n2811 gnd 0.007654f
C4281 vdd.n2812 gnd 0.007654f
C4282 vdd.n2813 gnd 0.007654f
C4283 vdd.n2814 gnd 0.007654f
C4284 vdd.n2815 gnd 0.007654f
C4285 vdd.n2816 gnd 0.007654f
C4286 vdd.n2817 gnd 0.007654f
C4287 vdd.n2818 gnd 0.007654f
C4288 vdd.n2819 gnd 0.007654f
C4289 vdd.n2820 gnd 0.007654f
C4290 vdd.n2821 gnd 0.007654f
C4291 vdd.n2822 gnd 0.007654f
C4292 vdd.n2823 gnd 0.007654f
C4293 vdd.n2824 gnd 0.007654f
C4294 vdd.n2825 gnd 0.007654f
C4295 vdd.n2826 gnd 0.007654f
C4296 vdd.n2827 gnd 0.007654f
C4297 vdd.n2828 gnd 0.007654f
C4298 vdd.n2829 gnd 0.007654f
C4299 vdd.n2830 gnd 0.007654f
C4300 vdd.n2831 gnd 0.007654f
C4301 vdd.n2832 gnd 0.007654f
C4302 vdd.n2833 gnd 0.007654f
C4303 vdd.n2834 gnd 0.007654f
C4304 vdd.n2835 gnd 0.007654f
C4305 vdd.n2836 gnd 0.007654f
C4306 vdd.n2837 gnd 0.007654f
C4307 vdd.n2838 gnd 0.007654f
C4308 vdd.n2839 gnd 0.007654f
C4309 vdd.n2840 gnd 0.007654f
C4310 vdd.n2841 gnd 0.007654f
C4311 vdd.n2842 gnd 0.007654f
C4312 vdd.n2843 gnd 0.007654f
C4313 vdd.n2844 gnd 0.007654f
C4314 vdd.n2845 gnd 0.007654f
C4315 vdd.n2846 gnd 0.007654f
C4316 vdd.n2847 gnd 0.007654f
C4317 vdd.n2848 gnd 0.007654f
C4318 vdd.n2849 gnd 0.007654f
C4319 vdd.n2850 gnd 0.007654f
C4320 vdd.n2851 gnd 0.007654f
C4321 vdd.n2852 gnd 0.007654f
C4322 vdd.n2853 gnd 0.007654f
C4323 vdd.n2854 gnd 0.007654f
C4324 vdd.n2855 gnd 0.007654f
C4325 vdd.n2857 gnd 0.954757f
C4326 vdd.n2859 gnd 0.007654f
C4327 vdd.n2860 gnd 0.007654f
C4328 vdd.n2861 gnd 0.018162f
C4329 vdd.n2862 gnd 0.016957f
C4330 vdd.n2863 gnd 0.016957f
C4331 vdd.n2864 gnd 0.954757f
C4332 vdd.n2865 gnd 0.016957f
C4333 vdd.n2866 gnd 0.016957f
C4334 vdd.n2867 gnd 0.007654f
C4335 vdd.n2868 gnd 0.007654f
C4336 vdd.n2869 gnd 0.007654f
C4337 vdd.n2870 gnd 0.488881f
C4338 vdd.n2871 gnd 0.007654f
C4339 vdd.n2872 gnd 0.007654f
C4340 vdd.n2873 gnd 0.007654f
C4341 vdd.n2874 gnd 0.007654f
C4342 vdd.n2875 gnd 0.007654f
C4343 vdd.n2876 gnd 0.609664f
C4344 vdd.n2877 gnd 0.007654f
C4345 vdd.n2878 gnd 0.007654f
C4346 vdd.n2879 gnd 0.007654f
C4347 vdd.n2880 gnd 0.007654f
C4348 vdd.n2881 gnd 0.007654f
C4349 vdd.n2882 gnd 0.78221f
C4350 vdd.n2883 gnd 0.007654f
C4351 vdd.n2884 gnd 0.007654f
C4352 vdd.n2885 gnd 0.007654f
C4353 vdd.n2886 gnd 0.007654f
C4354 vdd.n2887 gnd 0.007654f
C4355 vdd.n2888 gnd 0.431366f
C4356 vdd.n2889 gnd 0.007654f
C4357 vdd.n2890 gnd 0.007654f
C4358 vdd.n2891 gnd 0.007654f
C4359 vdd.n2892 gnd 0.007654f
C4360 vdd.n2893 gnd 0.007654f
C4361 vdd.n2894 gnd 0.247316f
C4362 vdd.n2895 gnd 0.007654f
C4363 vdd.n2896 gnd 0.007654f
C4364 vdd.n2897 gnd 0.007654f
C4365 vdd.n2898 gnd 0.007654f
C4366 vdd.n2899 gnd 0.007654f
C4367 vdd.n2900 gnd 0.448621f
C4368 vdd.n2901 gnd 0.007654f
C4369 vdd.n2902 gnd 0.007654f
C4370 vdd.n2903 gnd 0.007654f
C4371 vdd.n2904 gnd 0.007654f
C4372 vdd.n2905 gnd 0.007654f
C4373 vdd.n2906 gnd 0.621167f
C4374 vdd.n2907 gnd 0.007654f
C4375 vdd.n2908 gnd 0.007654f
C4376 vdd.n2909 gnd 0.007654f
C4377 vdd.n2910 gnd 0.007654f
C4378 vdd.n2911 gnd 0.007654f
C4379 vdd.n2912 gnd 0.695937f
C4380 vdd.n2913 gnd 0.007654f
C4381 vdd.n2914 gnd 0.007654f
C4382 vdd.n2915 gnd 0.007654f
C4383 vdd.n2916 gnd 0.007654f
C4384 vdd.n2917 gnd 0.007654f
C4385 vdd.n2918 gnd 0.523391f
C4386 vdd.n2919 gnd 0.007654f
C4387 vdd.n2920 gnd 0.007654f
C4388 vdd.n2921 gnd 0.007654f
C4389 vdd.t228 gnd 0.316607f
C4390 vdd.t226 gnd 0.201923f
C4391 vdd.t229 gnd 0.316607f
C4392 vdd.n2922 gnd 0.177946f
C4393 vdd.n2923 gnd 0.022173f
C4394 vdd.n2924 gnd 0.004728f
C4395 vdd.n2925 gnd 0.007654f
C4396 vdd.n2926 gnd 0.431366f
C4397 vdd.n2927 gnd 0.007654f
C4398 vdd.n2928 gnd 0.007654f
C4399 vdd.n2929 gnd 0.007654f
C4400 vdd.n2930 gnd 0.007654f
C4401 vdd.n2931 gnd 0.007654f
C4402 vdd.n2932 gnd 0.78221f
C4403 vdd.n2933 gnd 0.007654f
C4404 vdd.n2934 gnd 0.007654f
C4405 vdd.n2935 gnd 0.007654f
C4406 vdd.n2936 gnd 0.007654f
C4407 vdd.n2937 gnd 0.007654f
C4408 vdd.n2938 gnd 0.007654f
C4409 vdd.n2940 gnd 0.007654f
C4410 vdd.n2941 gnd 0.007654f
C4411 vdd.n2943 gnd 0.007654f
C4412 vdd.n2944 gnd 0.007654f
C4413 vdd.n2947 gnd 0.007654f
C4414 vdd.n2948 gnd 0.007654f
C4415 vdd.n2949 gnd 0.007654f
C4416 vdd.n2950 gnd 0.007654f
C4417 vdd.n2952 gnd 0.007654f
C4418 vdd.n2953 gnd 0.007654f
C4419 vdd.n2954 gnd 0.007654f
C4420 vdd.n2955 gnd 0.007654f
C4421 vdd.n2956 gnd 0.007654f
C4422 vdd.n2957 gnd 0.007654f
C4423 vdd.n2959 gnd 0.007654f
C4424 vdd.n2960 gnd 0.007654f
C4425 vdd.n2961 gnd 0.007654f
C4426 vdd.n2962 gnd 0.007654f
C4427 vdd.n2963 gnd 0.007654f
C4428 vdd.n2964 gnd 0.007654f
C4429 vdd.n2966 gnd 0.007654f
C4430 vdd.n2967 gnd 0.007654f
C4431 vdd.n2968 gnd 0.007654f
C4432 vdd.n2969 gnd 0.007654f
C4433 vdd.n2970 gnd 0.007654f
C4434 vdd.n2971 gnd 0.007654f
C4435 vdd.n2973 gnd 0.007654f
C4436 vdd.n2974 gnd 0.018162f
C4437 vdd.n2975 gnd 0.018162f
C4438 vdd.n2976 gnd 0.016957f
C4439 vdd.n2977 gnd 0.007654f
C4440 vdd.n2978 gnd 0.007654f
C4441 vdd.n2979 gnd 0.007654f
C4442 vdd.n2980 gnd 0.007654f
C4443 vdd.n2981 gnd 0.007654f
C4444 vdd.n2982 gnd 0.007654f
C4445 vdd.n2983 gnd 0.78221f
C4446 vdd.n2984 gnd 0.007654f
C4447 vdd.n2985 gnd 0.007654f
C4448 vdd.n2986 gnd 0.007654f
C4449 vdd.n2987 gnd 0.007654f
C4450 vdd.n2988 gnd 0.007654f
C4451 vdd.n2989 gnd 0.488881f
C4452 vdd.n2990 gnd 0.007654f
C4453 vdd.n2991 gnd 0.007654f
C4454 vdd.n2992 gnd 0.007654f
C4455 vdd.n2993 gnd 0.017889f
C4456 vdd.n2994 gnd 0.01723f
C4457 vdd.n2995 gnd 0.018162f
C4458 vdd.n2997 gnd 0.007654f
C4459 vdd.n2998 gnd 0.007654f
C4460 vdd.n2999 gnd 0.005909f
C4461 vdd.n3000 gnd 0.010939f
C4462 vdd.n3001 gnd 0.005572f
C4463 vdd.n3002 gnd 0.007654f
C4464 vdd.n3003 gnd 0.007654f
C4465 vdd.n3005 gnd 0.007654f
C4466 vdd.n3006 gnd 0.007654f
C4467 vdd.n3007 gnd 0.007654f
C4468 vdd.n3008 gnd 0.007654f
C4469 vdd.n3009 gnd 0.007654f
C4470 vdd.n3010 gnd 0.007654f
C4471 vdd.n3012 gnd 0.007654f
C4472 vdd.n3013 gnd 0.007654f
C4473 vdd.n3014 gnd 0.007654f
C4474 vdd.n3015 gnd 0.007654f
C4475 vdd.n3016 gnd 0.007654f
C4476 vdd.n3017 gnd 0.007654f
C4477 vdd.n3019 gnd 0.007654f
C4478 vdd.n3020 gnd 0.007654f
C4479 vdd.n3021 gnd 0.007654f
C4480 vdd.n3022 gnd 0.007654f
C4481 vdd.n3023 gnd 0.007654f
C4482 vdd.n3024 gnd 0.007654f
C4483 vdd.n3026 gnd 0.007654f
C4484 vdd.n3027 gnd 0.007654f
C4485 vdd.n3028 gnd 0.007654f
C4486 vdd.n3030 gnd 0.007654f
C4487 vdd.n3031 gnd 0.007654f
C4488 vdd.n3032 gnd 0.007654f
C4489 vdd.n3033 gnd 0.007654f
C4490 vdd.n3034 gnd 0.007654f
C4491 vdd.n3035 gnd 0.007654f
C4492 vdd.n3037 gnd 0.007654f
C4493 vdd.n3038 gnd 0.007654f
C4494 vdd.n3039 gnd 0.007654f
C4495 vdd.n3040 gnd 0.007654f
C4496 vdd.n3041 gnd 0.007654f
C4497 vdd.n3042 gnd 0.007654f
C4498 vdd.n3044 gnd 0.007654f
C4499 vdd.n3045 gnd 0.007654f
C4500 vdd.n3046 gnd 0.007654f
C4501 vdd.n3047 gnd 0.007654f
C4502 vdd.n3048 gnd 0.007654f
C4503 vdd.n3049 gnd 0.007654f
C4504 vdd.n3051 gnd 0.007654f
C4505 vdd.n3052 gnd 0.007654f
C4506 vdd.n3054 gnd 0.007654f
C4507 vdd.n3055 gnd 0.007654f
C4508 vdd.n3056 gnd 0.018162f
C4509 vdd.n3057 gnd 0.016957f
C4510 vdd.n3058 gnd 0.016957f
C4511 vdd.n3059 gnd 1.1273f
C4512 vdd.n3060 gnd 0.016957f
C4513 vdd.n3061 gnd 0.018162f
C4514 vdd.n3062 gnd 0.01723f
C4515 vdd.n3063 gnd 0.007654f
C4516 vdd.n3064 gnd 0.005909f
C4517 vdd.n3065 gnd 0.007654f
C4518 vdd.n3067 gnd 0.007654f
C4519 vdd.n3068 gnd 0.007654f
C4520 vdd.n3069 gnd 0.007654f
C4521 vdd.n3070 gnd 0.007654f
C4522 vdd.n3071 gnd 0.007654f
C4523 vdd.n3072 gnd 0.007654f
C4524 vdd.n3074 gnd 0.007654f
C4525 vdd.n3075 gnd 0.007654f
C4526 vdd.n3076 gnd 0.007654f
C4527 vdd.n3077 gnd 0.007654f
C4528 vdd.n3078 gnd 0.007654f
C4529 vdd.n3079 gnd 0.007654f
C4530 vdd.n3081 gnd 0.007654f
C4531 vdd.n3082 gnd 0.007654f
C4532 vdd.n3083 gnd 0.007654f
C4533 vdd.n3084 gnd 0.007654f
C4534 vdd.n3085 gnd 0.007654f
C4535 vdd.n3086 gnd 0.007654f
C4536 vdd.n3088 gnd 0.007654f
C4537 vdd.n3089 gnd 0.007654f
C4538 vdd.n3091 gnd 0.007654f
C4539 vdd.n3092 gnd 0.018393f
C4540 vdd.n3093 gnd 0.681231f
C4541 vdd.n3095 gnd 0.004756f
C4542 vdd.n3096 gnd 0.00906f
C4543 vdd.n3097 gnd 0.011256f
C4544 vdd.n3098 gnd 0.011256f
C4545 vdd.n3099 gnd 0.00906f
C4546 vdd.n3100 gnd 0.00906f
C4547 vdd.n3101 gnd 0.011256f
C4548 vdd.n3102 gnd 0.011256f
C4549 vdd.n3103 gnd 0.00906f
C4550 vdd.n3104 gnd 0.00906f
C4551 vdd.n3105 gnd 0.011256f
C4552 vdd.n3106 gnd 0.011256f
C4553 vdd.n3107 gnd 0.00906f
C4554 vdd.n3108 gnd 0.00906f
C4555 vdd.n3109 gnd 0.011256f
C4556 vdd.n3110 gnd 0.011256f
C4557 vdd.n3111 gnd 0.00906f
C4558 vdd.n3112 gnd 0.00906f
C4559 vdd.n3113 gnd 0.011256f
C4560 vdd.n3114 gnd 0.011256f
C4561 vdd.n3115 gnd 0.00906f
C4562 vdd.n3116 gnd 0.00906f
C4563 vdd.n3117 gnd 0.011256f
C4564 vdd.n3118 gnd 0.011256f
C4565 vdd.n3119 gnd 0.00906f
C4566 vdd.n3120 gnd 0.00906f
C4567 vdd.n3121 gnd 0.011256f
C4568 vdd.n3122 gnd 0.011256f
C4569 vdd.n3123 gnd 0.00906f
C4570 vdd.n3124 gnd 0.00906f
C4571 vdd.n3125 gnd 0.011256f
C4572 vdd.n3126 gnd 0.011256f
C4573 vdd.n3127 gnd 0.00906f
C4574 vdd.n3128 gnd 0.00906f
C4575 vdd.n3129 gnd 0.011256f
C4576 vdd.n3130 gnd 0.011256f
C4577 vdd.n3131 gnd 0.00906f
C4578 vdd.n3132 gnd 0.011256f
C4579 vdd.n3133 gnd 0.011256f
C4580 vdd.n3134 gnd 0.00906f
C4581 vdd.n3135 gnd 0.011256f
C4582 vdd.n3136 gnd 0.011256f
C4583 vdd.n3137 gnd 0.011256f
C4584 vdd.n3138 gnd 0.018482f
C4585 vdd.n3139 gnd 0.011256f
C4586 vdd.n3140 gnd 0.011256f
C4587 vdd.n3141 gnd 0.006161f
C4588 vdd.n3142 gnd 0.00906f
C4589 vdd.n3143 gnd 0.011256f
C4590 vdd.n3144 gnd 0.011256f
C4591 vdd.n3145 gnd 0.00906f
C4592 vdd.n3146 gnd 0.00906f
C4593 vdd.n3147 gnd 0.011256f
C4594 vdd.n3148 gnd 0.011256f
C4595 vdd.n3149 gnd 0.00906f
C4596 vdd.n3150 gnd 0.00906f
C4597 vdd.n3151 gnd 0.011256f
C4598 vdd.n3152 gnd 0.011256f
C4599 vdd.n3153 gnd 0.00906f
C4600 vdd.n3154 gnd 0.00906f
C4601 vdd.n3155 gnd 0.011256f
C4602 vdd.n3156 gnd 0.011256f
C4603 vdd.n3157 gnd 0.00906f
C4604 vdd.n3158 gnd 0.00906f
C4605 vdd.n3159 gnd 0.011256f
C4606 vdd.n3160 gnd 0.011256f
C4607 vdd.n3161 gnd 0.00906f
C4608 vdd.n3162 gnd 0.00906f
C4609 vdd.n3163 gnd 0.011256f
C4610 vdd.n3164 gnd 0.011256f
C4611 vdd.n3165 gnd 0.00906f
C4612 vdd.n3166 gnd 0.00906f
C4613 vdd.n3167 gnd 0.011256f
C4614 vdd.n3168 gnd 0.011256f
C4615 vdd.n3169 gnd 0.00906f
C4616 vdd.n3170 gnd 0.00906f
C4617 vdd.n3171 gnd 0.011256f
C4618 vdd.n3172 gnd 0.011256f
C4619 vdd.n3173 gnd 0.00906f
C4620 vdd.n3174 gnd 0.00906f
C4621 vdd.n3175 gnd 0.011256f
C4622 vdd.n3176 gnd 0.011256f
C4623 vdd.n3177 gnd 0.00906f
C4624 vdd.n3178 gnd 0.011256f
C4625 vdd.n3179 gnd 0.011256f
C4626 vdd.n3180 gnd 0.00906f
C4627 vdd.n3181 gnd 0.011256f
C4628 vdd.n3182 gnd 0.011256f
C4629 vdd.n3183 gnd 0.011256f
C4630 vdd.t220 gnd 0.138478f
C4631 vdd.t221 gnd 0.147995f
C4632 vdd.t219 gnd 0.180851f
C4633 vdd.n3184 gnd 0.231825f
C4634 vdd.n3185 gnd 0.194775f
C4635 vdd.n3186 gnd 0.018482f
C4636 vdd.n3187 gnd 0.011256f
C4637 vdd.n3188 gnd 0.011256f
C4638 vdd.n3189 gnd 0.007565f
C4639 vdd.n3190 gnd 0.00906f
C4640 vdd.n3191 gnd 0.011256f
C4641 vdd.n3192 gnd 0.011256f
C4642 vdd.n3193 gnd 0.00906f
C4643 vdd.n3194 gnd 0.00906f
C4644 vdd.n3195 gnd 0.011256f
C4645 vdd.n3196 gnd 0.011256f
C4646 vdd.n3197 gnd 0.00906f
C4647 vdd.n3198 gnd 0.00906f
C4648 vdd.n3199 gnd 0.011256f
C4649 vdd.n3200 gnd 0.011256f
C4650 vdd.n3201 gnd 0.00906f
C4651 vdd.n3202 gnd 0.00906f
C4652 vdd.n3203 gnd 0.011256f
C4653 vdd.n3204 gnd 0.011256f
C4654 vdd.n3205 gnd 0.00906f
C4655 vdd.n3206 gnd 0.00906f
C4656 vdd.n3207 gnd 0.011256f
C4657 vdd.n3208 gnd 0.011256f
C4658 vdd.n3209 gnd 0.00906f
C4659 vdd.n3210 gnd 0.00906f
C4660 vdd.n3211 gnd 0.011256f
C4661 vdd.n3212 gnd 0.011256f
C4662 vdd.n3213 gnd 0.00906f
C4663 vdd.n3214 gnd 0.00906f
C4664 vdd.n3216 gnd 0.681231f
C4665 vdd.n3218 gnd 0.00906f
C4666 vdd.n3219 gnd 0.00906f
C4667 vdd.n3220 gnd 0.00752f
C4668 vdd.n3221 gnd 0.027813f
C4669 vdd.n3223 gnd 8.31674f
C4670 vdd.n3224 gnd 0.027813f
C4671 vdd.n3225 gnd 0.004303f
C4672 vdd.n3226 gnd 0.027813f
C4673 vdd.n3227 gnd 0.027229f
C4674 vdd.n3228 gnd 0.011256f
C4675 vdd.n3229 gnd 0.00906f
C4676 vdd.n3230 gnd 0.011256f
C4677 vdd.n3231 gnd 0.695937f
C4678 vdd.n3232 gnd 0.011256f
C4679 vdd.n3233 gnd 0.00906f
C4680 vdd.n3234 gnd 0.011256f
C4681 vdd.n3235 gnd 0.011256f
C4682 vdd.n3236 gnd 0.011256f
C4683 vdd.n3237 gnd 0.00906f
C4684 vdd.n3238 gnd 0.011256f
C4685 vdd.n3239 gnd 1.15031f
C4686 vdd.n3240 gnd 0.011256f
C4687 vdd.n3241 gnd 0.00906f
C4688 vdd.n3242 gnd 0.011256f
C4689 vdd.n3243 gnd 0.011256f
C4690 vdd.n3244 gnd 0.011256f
C4691 vdd.n3245 gnd 0.00906f
C4692 vdd.n3246 gnd 0.011256f
C4693 vdd.n3247 gnd 0.741949f
C4694 vdd.n3248 gnd 0.787962f
C4695 vdd.n3249 gnd 0.011256f
C4696 vdd.n3250 gnd 0.00906f
C4697 vdd.n3251 gnd 0.011256f
C4698 vdd.n3252 gnd 0.011256f
C4699 vdd.n3253 gnd 0.011256f
C4700 vdd.n3254 gnd 0.00906f
C4701 vdd.n3255 gnd 0.011256f
C4702 vdd.n3256 gnd 0.954757f
C4703 vdd.n3257 gnd 0.011256f
C4704 vdd.n3258 gnd 0.00906f
C4705 vdd.n3259 gnd 0.011256f
C4706 vdd.n3260 gnd 0.011256f
C4707 vdd.n3261 gnd 0.011256f
C4708 vdd.n3262 gnd 0.00906f
C4709 vdd.n3263 gnd 0.011256f
C4710 vdd.t27 gnd 0.575155f
C4711 vdd.n3264 gnd 0.925999f
C4712 vdd.n3265 gnd 0.011256f
C4713 vdd.n3266 gnd 0.00906f
C4714 vdd.n3267 gnd 0.011256f
C4715 vdd.n3268 gnd 0.011256f
C4716 vdd.n3269 gnd 0.011256f
C4717 vdd.n3270 gnd 0.00906f
C4718 vdd.n3271 gnd 0.011256f
C4719 vdd.n3272 gnd 0.730446f
C4720 vdd.n3273 gnd 0.011256f
C4721 vdd.n3274 gnd 0.00906f
C4722 vdd.n3275 gnd 0.011256f
C4723 vdd.n3276 gnd 0.011256f
C4724 vdd.n3277 gnd 0.011256f
C4725 vdd.n3278 gnd 0.00906f
C4726 vdd.n3279 gnd 0.011256f
C4727 vdd.n3280 gnd 0.914496f
C4728 vdd.n3281 gnd 0.615415f
C4729 vdd.n3282 gnd 0.011256f
C4730 vdd.n3283 gnd 0.00906f
C4731 vdd.n3284 gnd 0.011256f
C4732 vdd.n3285 gnd 0.011256f
C4733 vdd.n3286 gnd 0.011256f
C4734 vdd.n3287 gnd 0.00906f
C4735 vdd.n3288 gnd 0.011256f
C4736 vdd.n3289 gnd 0.810968f
C4737 vdd.n3290 gnd 0.011256f
C4738 vdd.n3291 gnd 0.00906f
C4739 vdd.n3292 gnd 0.011256f
C4740 vdd.n3293 gnd 0.011256f
C4741 vdd.n3294 gnd 0.011256f
C4742 vdd.n3295 gnd 0.011256f
C4743 vdd.n3296 gnd 0.011256f
C4744 vdd.n3297 gnd 0.00906f
C4745 vdd.n3298 gnd 0.00906f
C4746 vdd.n3299 gnd 0.011256f
C4747 vdd.t75 gnd 0.575155f
C4748 vdd.n3300 gnd 0.954757f
C4749 vdd.n3301 gnd 0.011256f
C4750 vdd.n3302 gnd 0.00906f
C4751 vdd.n3303 gnd 0.011256f
C4752 vdd.n3304 gnd 0.011256f
C4753 vdd.n3305 gnd 0.011256f
C4754 vdd.n3306 gnd 0.00906f
C4755 vdd.n3307 gnd 0.011256f
C4756 vdd.n3308 gnd 0.902993f
C4757 vdd.n3309 gnd 0.011256f
C4758 vdd.n3310 gnd 0.011256f
C4759 vdd.n3311 gnd 0.00906f
C4760 vdd.n3312 gnd 0.00906f
C4761 vdd.n3313 gnd 0.011256f
C4762 vdd.n3314 gnd 0.011256f
C4763 vdd.n3315 gnd 0.011256f
C4764 vdd.n3316 gnd 0.00906f
C4765 vdd.n3317 gnd 0.011256f
C4766 vdd.n3318 gnd 0.00906f
C4767 vdd.n3319 gnd 0.00906f
C4768 vdd.n3320 gnd 0.011256f
C4769 vdd.n3321 gnd 0.011256f
C4770 vdd.n3322 gnd 0.011256f
C4771 vdd.n3323 gnd 0.00906f
C4772 vdd.n3324 gnd 0.011256f
C4773 vdd.n3325 gnd 0.00906f
C4774 vdd.n3326 gnd 0.00906f
C4775 vdd.n3327 gnd 0.011256f
C4776 vdd.n3328 gnd 0.011256f
C4777 vdd.n3329 gnd 0.011256f
C4778 vdd.n3330 gnd 0.00906f
C4779 vdd.n3331 gnd 0.954757f
C4780 vdd.n3332 gnd 0.011256f
C4781 vdd.n3333 gnd 0.00906f
C4782 vdd.n3334 gnd 0.00906f
C4783 vdd.n3335 gnd 0.011256f
C4784 vdd.n3336 gnd 0.011256f
C4785 vdd.n3337 gnd 0.011256f
C4786 vdd.n3338 gnd 0.00906f
C4787 vdd.n3339 gnd 0.011256f
C4788 vdd.n3340 gnd 0.00906f
C4789 vdd.n3341 gnd 0.00906f
C4790 vdd.n3342 gnd 0.011256f
C4791 vdd.n3343 gnd 0.011256f
C4792 vdd.n3344 gnd 0.011256f
C4793 vdd.n3345 gnd 0.00906f
C4794 vdd.n3346 gnd 0.011256f
C4795 vdd.n3347 gnd 0.00906f
C4796 vdd.n3348 gnd 0.00752f
C4797 vdd.n3349 gnd 0.027229f
C4798 vdd.n3350 gnd 0.027813f
C4799 vdd.n3351 gnd 0.004303f
C4800 vdd.n3352 gnd 0.027813f
C4801 vdd.n3354 gnd 2.72623f
C4802 vdd.n3355 gnd 1.69671f
C4803 vdd.n3356 gnd 0.027229f
C4804 vdd.n3357 gnd 0.00752f
C4805 vdd.n3358 gnd 0.00906f
C4806 vdd.n3359 gnd 0.00906f
C4807 vdd.n3360 gnd 0.011256f
C4808 vdd.n3361 gnd 1.15031f
C4809 vdd.n3362 gnd 1.15031f
C4810 vdd.n3363 gnd 1.05253f
C4811 vdd.n3364 gnd 0.011256f
C4812 vdd.n3365 gnd 0.00906f
C4813 vdd.n3366 gnd 0.00906f
C4814 vdd.n3367 gnd 0.00906f
C4815 vdd.n3368 gnd 0.011256f
C4816 vdd.n3369 gnd 0.85698f
C4817 vdd.t94 gnd 0.575155f
C4818 vdd.n3370 gnd 0.868483f
C4819 vdd.n3371 gnd 0.661428f
C4820 vdd.n3372 gnd 0.011256f
C4821 vdd.n3373 gnd 0.00906f
C4822 vdd.n3374 gnd 0.00906f
C4823 vdd.n3375 gnd 0.00906f
C4824 vdd.n3376 gnd 0.011256f
C4825 vdd.n3377 gnd 0.684434f
C4826 vdd.n3378 gnd 0.845477f
C4827 vdd.t45 gnd 0.575155f
C4828 vdd.n3379 gnd 0.879987f
C4829 vdd.n3380 gnd 0.011256f
C4830 vdd.n3381 gnd 0.00906f
C4831 vdd.n3382 gnd 0.00906f
C4832 vdd.n3383 gnd 0.00906f
C4833 vdd.n3384 gnd 0.011256f
C4834 vdd.n3385 gnd 0.954757f
C4835 vdd.t71 gnd 0.575155f
C4836 vdd.n3386 gnd 0.695937f
C4837 vdd.n3387 gnd 0.833974f
C4838 vdd.n3388 gnd 0.011256f
C4839 vdd.n3389 gnd 0.00906f
C4840 vdd.n3390 gnd 0.00906f
C4841 vdd.n3391 gnd 0.00906f
C4842 vdd.n3392 gnd 0.011256f
C4843 vdd.n3393 gnd 0.638422f
C4844 vdd.t41 gnd 0.575155f
C4845 vdd.n3394 gnd 0.954757f
C4846 vdd.t68 gnd 0.575155f
C4847 vdd.n3395 gnd 0.70744f
C4848 vdd.n3396 gnd 0.011256f
C4849 vdd.n3397 gnd 0.00906f
C4850 vdd.n3398 gnd 0.008651f
C4851 vdd.n3399 gnd 0.663921f
C4852 vdd.n3400 gnd 2.87832f
C4853 a_n7636_8799.n0 gnd 0.208536f
C4854 a_n7636_8799.n1 gnd 0.286348f
C4855 a_n7636_8799.n2 gnd 0.208536f
C4856 a_n7636_8799.n3 gnd 0.208536f
C4857 a_n7636_8799.n4 gnd 0.208536f
C4858 a_n7636_8799.n5 gnd 0.208536f
C4859 a_n7636_8799.n6 gnd 0.208536f
C4860 a_n7636_8799.n7 gnd 0.21684f
C4861 a_n7636_8799.n8 gnd 0.208536f
C4862 a_n7636_8799.n9 gnd 0.286348f
C4863 a_n7636_8799.n10 gnd 0.208536f
C4864 a_n7636_8799.n11 gnd 0.208536f
C4865 a_n7636_8799.n12 gnd 0.208536f
C4866 a_n7636_8799.n13 gnd 0.208536f
C4867 a_n7636_8799.n14 gnd 0.208536f
C4868 a_n7636_8799.n15 gnd 0.21684f
C4869 a_n7636_8799.n16 gnd 0.208536f
C4870 a_n7636_8799.n17 gnd 0.451989f
C4871 a_n7636_8799.n18 gnd 0.208536f
C4872 a_n7636_8799.n19 gnd 0.208536f
C4873 a_n7636_8799.n20 gnd 0.208536f
C4874 a_n7636_8799.n21 gnd 0.208536f
C4875 a_n7636_8799.n22 gnd 0.208536f
C4876 a_n7636_8799.n23 gnd 0.21684f
C4877 a_n7636_8799.n24 gnd 0.208536f
C4878 a_n7636_8799.n25 gnd 0.321108f
C4879 a_n7636_8799.n26 gnd 0.208536f
C4880 a_n7636_8799.n27 gnd 0.208536f
C4881 a_n7636_8799.n28 gnd 0.208536f
C4882 a_n7636_8799.n29 gnd 0.208536f
C4883 a_n7636_8799.n30 gnd 0.208536f
C4884 a_n7636_8799.n31 gnd 0.182079f
C4885 a_n7636_8799.n32 gnd 0.208536f
C4886 a_n7636_8799.n33 gnd 0.321108f
C4887 a_n7636_8799.n34 gnd 0.208536f
C4888 a_n7636_8799.n35 gnd 0.208536f
C4889 a_n7636_8799.n36 gnd 0.208536f
C4890 a_n7636_8799.n37 gnd 0.208536f
C4891 a_n7636_8799.n38 gnd 0.208536f
C4892 a_n7636_8799.n39 gnd 0.182079f
C4893 a_n7636_8799.n40 gnd 0.208536f
C4894 a_n7636_8799.n41 gnd 0.321108f
C4895 a_n7636_8799.n42 gnd 0.208536f
C4896 a_n7636_8799.n43 gnd 0.208536f
C4897 a_n7636_8799.n44 gnd 0.208536f
C4898 a_n7636_8799.n45 gnd 0.208536f
C4899 a_n7636_8799.n46 gnd 0.208536f
C4900 a_n7636_8799.n47 gnd 0.347721f
C4901 a_n7636_8799.n48 gnd 2.87986f
C4902 a_n7636_8799.n49 gnd 3.94234f
C4903 a_n7636_8799.n50 gnd 2.39774f
C4904 a_n7636_8799.n51 gnd 1.40139f
C4905 a_n7636_8799.n52 gnd 3.10218f
C4906 a_n7636_8799.n53 gnd 0.251058f
C4907 a_n7636_8799.n54 gnd 0.00367f
C4908 a_n7636_8799.n55 gnd 0.009675f
C4909 a_n7636_8799.n56 gnd 0.010571f
C4910 a_n7636_8799.n57 gnd 0.005586f
C4911 a_n7636_8799.n59 gnd 0.004687f
C4912 a_n7636_8799.n60 gnd 0.010137f
C4913 a_n7636_8799.n61 gnd 0.010137f
C4914 a_n7636_8799.n62 gnd 0.004687f
C4915 a_n7636_8799.n64 gnd 0.005586f
C4916 a_n7636_8799.n65 gnd 0.010571f
C4917 a_n7636_8799.n66 gnd 0.009675f
C4918 a_n7636_8799.n67 gnd 0.00367f
C4919 a_n7636_8799.n68 gnd 0.251058f
C4920 a_n7636_8799.n69 gnd 0.00367f
C4921 a_n7636_8799.n70 gnd 0.009675f
C4922 a_n7636_8799.n71 gnd 0.010571f
C4923 a_n7636_8799.n72 gnd 0.005586f
C4924 a_n7636_8799.n74 gnd 0.004687f
C4925 a_n7636_8799.n75 gnd 0.010137f
C4926 a_n7636_8799.n76 gnd 0.010137f
C4927 a_n7636_8799.n77 gnd 0.004687f
C4928 a_n7636_8799.n79 gnd 0.005586f
C4929 a_n7636_8799.n80 gnd 0.010571f
C4930 a_n7636_8799.n81 gnd 0.009675f
C4931 a_n7636_8799.n82 gnd 0.00367f
C4932 a_n7636_8799.n83 gnd 0.251058f
C4933 a_n7636_8799.n84 gnd 0.00367f
C4934 a_n7636_8799.n85 gnd 0.009675f
C4935 a_n7636_8799.n86 gnd 0.010571f
C4936 a_n7636_8799.n87 gnd 0.005586f
C4937 a_n7636_8799.n89 gnd 0.004687f
C4938 a_n7636_8799.n90 gnd 0.010137f
C4939 a_n7636_8799.n91 gnd 0.010137f
C4940 a_n7636_8799.n92 gnd 0.004687f
C4941 a_n7636_8799.n94 gnd 0.005586f
C4942 a_n7636_8799.n95 gnd 0.010571f
C4943 a_n7636_8799.n96 gnd 0.009675f
C4944 a_n7636_8799.n97 gnd 0.00367f
C4945 a_n7636_8799.n98 gnd 0.00367f
C4946 a_n7636_8799.n99 gnd 0.009675f
C4947 a_n7636_8799.n100 gnd 0.010571f
C4948 a_n7636_8799.n101 gnd 0.005586f
C4949 a_n7636_8799.n103 gnd 0.004687f
C4950 a_n7636_8799.n104 gnd 0.010137f
C4951 a_n7636_8799.n105 gnd 0.010137f
C4952 a_n7636_8799.n106 gnd 0.004687f
C4953 a_n7636_8799.n108 gnd 0.005586f
C4954 a_n7636_8799.n109 gnd 0.010571f
C4955 a_n7636_8799.n110 gnd 0.009675f
C4956 a_n7636_8799.n111 gnd 0.00367f
C4957 a_n7636_8799.n112 gnd 0.251058f
C4958 a_n7636_8799.n113 gnd 0.00367f
C4959 a_n7636_8799.n114 gnd 0.009675f
C4960 a_n7636_8799.n115 gnd 0.010571f
C4961 a_n7636_8799.n116 gnd 0.005586f
C4962 a_n7636_8799.n118 gnd 0.004687f
C4963 a_n7636_8799.n119 gnd 0.010137f
C4964 a_n7636_8799.n120 gnd 0.010137f
C4965 a_n7636_8799.n121 gnd 0.004687f
C4966 a_n7636_8799.n123 gnd 0.005586f
C4967 a_n7636_8799.n124 gnd 0.010571f
C4968 a_n7636_8799.n125 gnd 0.009675f
C4969 a_n7636_8799.n126 gnd 0.00367f
C4970 a_n7636_8799.n127 gnd 0.251058f
C4971 a_n7636_8799.n128 gnd 0.00367f
C4972 a_n7636_8799.n129 gnd 0.009675f
C4973 a_n7636_8799.n130 gnd 0.010571f
C4974 a_n7636_8799.n131 gnd 0.005586f
C4975 a_n7636_8799.n133 gnd 0.004687f
C4976 a_n7636_8799.n134 gnd 0.010137f
C4977 a_n7636_8799.n135 gnd 0.010137f
C4978 a_n7636_8799.n136 gnd 0.004687f
C4979 a_n7636_8799.n138 gnd 0.005586f
C4980 a_n7636_8799.n139 gnd 0.010571f
C4981 a_n7636_8799.n140 gnd 0.009675f
C4982 a_n7636_8799.n141 gnd 0.00367f
C4983 a_n7636_8799.n142 gnd 0.251058f
C4984 a_n7636_8799.t25 gnd 0.144643f
C4985 a_n7636_8799.t3 gnd 0.144643f
C4986 a_n7636_8799.t5 gnd 0.144643f
C4987 a_n7636_8799.n143 gnd 1.14082f
C4988 a_n7636_8799.t22 gnd 0.144643f
C4989 a_n7636_8799.t1 gnd 0.144643f
C4990 a_n7636_8799.n144 gnd 1.13894f
C4991 a_n7636_8799.t15 gnd 0.144643f
C4992 a_n7636_8799.t2 gnd 0.144643f
C4993 a_n7636_8799.n145 gnd 1.13894f
C4994 a_n7636_8799.t11 gnd 0.1125f
C4995 a_n7636_8799.t23 gnd 0.1125f
C4996 a_n7636_8799.n146 gnd 0.995675f
C4997 a_n7636_8799.t14 gnd 0.1125f
C4998 a_n7636_8799.t16 gnd 0.1125f
C4999 a_n7636_8799.n147 gnd 0.994091f
C5000 a_n7636_8799.t12 gnd 0.1125f
C5001 a_n7636_8799.t8 gnd 0.1125f
C5002 a_n7636_8799.n148 gnd 0.995674f
C5003 a_n7636_8799.t7 gnd 0.1125f
C5004 a_n7636_8799.t17 gnd 0.1125f
C5005 a_n7636_8799.n149 gnd 0.99409f
C5006 a_n7636_8799.t21 gnd 0.1125f
C5007 a_n7636_8799.t9 gnd 0.1125f
C5008 a_n7636_8799.n150 gnd 0.995674f
C5009 a_n7636_8799.t13 gnd 0.1125f
C5010 a_n7636_8799.t27 gnd 0.1125f
C5011 a_n7636_8799.n151 gnd 0.99409f
C5012 a_n7636_8799.t20 gnd 0.1125f
C5013 a_n7636_8799.t6 gnd 0.1125f
C5014 a_n7636_8799.n152 gnd 0.994091f
C5015 a_n7636_8799.t24 gnd 0.1125f
C5016 a_n7636_8799.t18 gnd 0.1125f
C5017 a_n7636_8799.n153 gnd 0.994091f
C5018 a_n7636_8799.t124 gnd 0.599757f
C5019 a_n7636_8799.n154 gnd 0.270018f
C5020 a_n7636_8799.t40 gnd 0.599757f
C5021 a_n7636_8799.t61 gnd 0.599757f
C5022 a_n7636_8799.n155 gnd 0.271953f
C5023 a_n7636_8799.t84 gnd 0.599757f
C5024 a_n7636_8799.t103 gnd 0.599757f
C5025 a_n7636_8799.n156 gnd 0.265131f
C5026 a_n7636_8799.t63 gnd 0.599757f
C5027 a_n7636_8799.t75 gnd 0.599757f
C5028 a_n7636_8799.n157 gnd 0.269123f
C5029 a_n7636_8799.t108 gnd 0.599757f
C5030 a_n7636_8799.t129 gnd 0.599757f
C5031 a_n7636_8799.t127 gnd 0.611109f
C5032 a_n7636_8799.n158 gnd 0.251423f
C5033 a_n7636_8799.n159 gnd 0.272327f
C5034 a_n7636_8799.t79 gnd 0.599757f
C5035 a_n7636_8799.n160 gnd 0.270018f
C5036 a_n7636_8799.n161 gnd 0.265774f
C5037 a_n7636_8799.t125 gnd 0.599757f
C5038 a_n7636_8799.n162 gnd 0.264488f
C5039 a_n7636_8799.t76 gnd 0.599757f
C5040 a_n7636_8799.n163 gnd 0.271697f
C5041 a_n7636_8799.t106 gnd 0.599757f
C5042 a_n7636_8799.n164 gnd 0.271953f
C5043 a_n7636_8799.n165 gnd 0.269557f
C5044 a_n7636_8799.t64 gnd 0.599757f
C5045 a_n7636_8799.n166 gnd 0.265131f
C5046 a_n7636_8799.t28 gnd 0.599757f
C5047 a_n7636_8799.n167 gnd 0.269557f
C5048 a_n7636_8799.n168 gnd 0.271697f
C5049 a_n7636_8799.t128 gnd 0.599757f
C5050 a_n7636_8799.n169 gnd 0.269123f
C5051 a_n7636_8799.n170 gnd 0.264488f
C5052 a_n7636_8799.t58 gnd 0.599757f
C5053 a_n7636_8799.n171 gnd 0.265774f
C5054 a_n7636_8799.t37 gnd 0.599757f
C5055 a_n7636_8799.n172 gnd 0.272327f
C5056 a_n7636_8799.t38 gnd 0.611098f
C5057 a_n7636_8799.t137 gnd 0.599757f
C5058 a_n7636_8799.n173 gnd 0.270018f
C5059 a_n7636_8799.t55 gnd 0.599757f
C5060 a_n7636_8799.t70 gnd 0.599757f
C5061 a_n7636_8799.n174 gnd 0.271953f
C5062 a_n7636_8799.t97 gnd 0.599757f
C5063 a_n7636_8799.t115 gnd 0.599757f
C5064 a_n7636_8799.n175 gnd 0.265131f
C5065 a_n7636_8799.t73 gnd 0.599757f
C5066 a_n7636_8799.t85 gnd 0.599757f
C5067 a_n7636_8799.n176 gnd 0.269123f
C5068 a_n7636_8799.t121 gnd 0.599757f
C5069 a_n7636_8799.t145 gnd 0.599757f
C5070 a_n7636_8799.t142 gnd 0.611109f
C5071 a_n7636_8799.n177 gnd 0.251423f
C5072 a_n7636_8799.n178 gnd 0.272327f
C5073 a_n7636_8799.t89 gnd 0.599757f
C5074 a_n7636_8799.n179 gnd 0.270018f
C5075 a_n7636_8799.n180 gnd 0.265774f
C5076 a_n7636_8799.t139 gnd 0.599757f
C5077 a_n7636_8799.n181 gnd 0.264488f
C5078 a_n7636_8799.t86 gnd 0.599757f
C5079 a_n7636_8799.n182 gnd 0.271697f
C5080 a_n7636_8799.t119 gnd 0.599757f
C5081 a_n7636_8799.n183 gnd 0.271953f
C5082 a_n7636_8799.n184 gnd 0.269557f
C5083 a_n7636_8799.t74 gnd 0.599757f
C5084 a_n7636_8799.n185 gnd 0.265131f
C5085 a_n7636_8799.t39 gnd 0.599757f
C5086 a_n7636_8799.n186 gnd 0.269557f
C5087 a_n7636_8799.n187 gnd 0.271697f
C5088 a_n7636_8799.t143 gnd 0.599757f
C5089 a_n7636_8799.n188 gnd 0.269123f
C5090 a_n7636_8799.n189 gnd 0.264488f
C5091 a_n7636_8799.t69 gnd 0.599757f
C5092 a_n7636_8799.n190 gnd 0.265774f
C5093 a_n7636_8799.t49 gnd 0.599757f
C5094 a_n7636_8799.n191 gnd 0.272327f
C5095 a_n7636_8799.t51 gnd 0.611098f
C5096 a_n7636_8799.n192 gnd 0.901652f
C5097 a_n7636_8799.t92 gnd 0.599757f
C5098 a_n7636_8799.n193 gnd 0.270018f
C5099 a_n7636_8799.t116 gnd 0.599757f
C5100 a_n7636_8799.t34 gnd 0.599757f
C5101 a_n7636_8799.n194 gnd 0.271953f
C5102 a_n7636_8799.t99 gnd 0.599757f
C5103 a_n7636_8799.t138 gnd 0.599757f
C5104 a_n7636_8799.n195 gnd 0.265131f
C5105 a_n7636_8799.t133 gnd 0.599757f
C5106 a_n7636_8799.t46 gnd 0.599757f
C5107 a_n7636_8799.n196 gnd 0.269123f
C5108 a_n7636_8799.t71 gnd 0.599757f
C5109 a_n7636_8799.t82 gnd 0.599757f
C5110 a_n7636_8799.t104 gnd 0.611109f
C5111 a_n7636_8799.n197 gnd 0.251423f
C5112 a_n7636_8799.n198 gnd 0.272327f
C5113 a_n7636_8799.t120 gnd 0.599757f
C5114 a_n7636_8799.n199 gnd 0.270018f
C5115 a_n7636_8799.n200 gnd 0.265774f
C5116 a_n7636_8799.t130 gnd 0.599757f
C5117 a_n7636_8799.n201 gnd 0.264488f
C5118 a_n7636_8799.t29 gnd 0.599757f
C5119 a_n7636_8799.n202 gnd 0.271697f
C5120 a_n7636_8799.t90 gnd 0.599757f
C5121 a_n7636_8799.n203 gnd 0.271953f
C5122 a_n7636_8799.n204 gnd 0.269557f
C5123 a_n7636_8799.t107 gnd 0.599757f
C5124 a_n7636_8799.n205 gnd 0.265131f
C5125 a_n7636_8799.t83 gnd 0.599757f
C5126 a_n7636_8799.n206 gnd 0.269557f
C5127 a_n7636_8799.n207 gnd 0.271697f
C5128 a_n7636_8799.t53 gnd 0.599757f
C5129 a_n7636_8799.n208 gnd 0.269123f
C5130 a_n7636_8799.n209 gnd 0.264488f
C5131 a_n7636_8799.t62 gnd 0.599757f
C5132 a_n7636_8799.n210 gnd 0.265774f
C5133 a_n7636_8799.t42 gnd 0.599757f
C5134 a_n7636_8799.n211 gnd 0.272327f
C5135 a_n7636_8799.t144 gnd 0.611098f
C5136 a_n7636_8799.n212 gnd 1.40196f
C5137 a_n7636_8799.t78 gnd 0.611098f
C5138 a_n7636_8799.t77 gnd 0.599757f
C5139 a_n7636_8799.t50 gnd 0.599757f
C5140 a_n7636_8799.n213 gnd 0.270018f
C5141 a_n7636_8799.t126 gnd 0.599757f
C5142 a_n7636_8799.t81 gnd 0.599757f
C5143 a_n7636_8799.t57 gnd 0.599757f
C5144 a_n7636_8799.n214 gnd 0.269123f
C5145 a_n7636_8799.t132 gnd 0.599757f
C5146 a_n7636_8799.t98 gnd 0.599757f
C5147 a_n7636_8799.t96 gnd 0.599757f
C5148 a_n7636_8799.n215 gnd 0.269557f
C5149 a_n7636_8799.t31 gnd 0.599757f
C5150 a_n7636_8799.t102 gnd 0.599757f
C5151 a_n7636_8799.t101 gnd 0.599757f
C5152 a_n7636_8799.n216 gnd 0.269557f
C5153 a_n7636_8799.t33 gnd 0.599757f
C5154 a_n7636_8799.t32 gnd 0.599757f
C5155 a_n7636_8799.t118 gnd 0.599757f
C5156 a_n7636_8799.n217 gnd 0.269123f
C5157 a_n7636_8799.t52 gnd 0.599757f
C5158 a_n7636_8799.t36 gnd 0.599757f
C5159 a_n7636_8799.t122 gnd 0.599757f
C5160 a_n7636_8799.n218 gnd 0.270018f
C5161 a_n7636_8799.t56 gnd 0.611109f
C5162 a_n7636_8799.n219 gnd 0.251423f
C5163 a_n7636_8799.t80 gnd 0.599757f
C5164 a_n7636_8799.n220 gnd 0.272327f
C5165 a_n7636_8799.n221 gnd 0.265774f
C5166 a_n7636_8799.n222 gnd 0.264488f
C5167 a_n7636_8799.n223 gnd 0.271697f
C5168 a_n7636_8799.n224 gnd 0.271953f
C5169 a_n7636_8799.n225 gnd 0.265131f
C5170 a_n7636_8799.n226 gnd 0.265131f
C5171 a_n7636_8799.n227 gnd 0.271953f
C5172 a_n7636_8799.n228 gnd 0.271697f
C5173 a_n7636_8799.n229 gnd 0.264488f
C5174 a_n7636_8799.n230 gnd 0.265774f
C5175 a_n7636_8799.n231 gnd 0.272327f
C5176 a_n7636_8799.t88 gnd 0.611098f
C5177 a_n7636_8799.t87 gnd 0.599757f
C5178 a_n7636_8799.t65 gnd 0.599757f
C5179 a_n7636_8799.n232 gnd 0.270018f
C5180 a_n7636_8799.t141 gnd 0.599757f
C5181 a_n7636_8799.t94 gnd 0.599757f
C5182 a_n7636_8799.t67 gnd 0.599757f
C5183 a_n7636_8799.n233 gnd 0.269123f
C5184 a_n7636_8799.t147 gnd 0.599757f
C5185 a_n7636_8799.t111 gnd 0.599757f
C5186 a_n7636_8799.t110 gnd 0.599757f
C5187 a_n7636_8799.n234 gnd 0.269557f
C5188 a_n7636_8799.t41 gnd 0.599757f
C5189 a_n7636_8799.t114 gnd 0.599757f
C5190 a_n7636_8799.t113 gnd 0.599757f
C5191 a_n7636_8799.n235 gnd 0.269557f
C5192 a_n7636_8799.t45 gnd 0.599757f
C5193 a_n7636_8799.t44 gnd 0.599757f
C5194 a_n7636_8799.t135 gnd 0.599757f
C5195 a_n7636_8799.n236 gnd 0.269123f
C5196 a_n7636_8799.t66 gnd 0.599757f
C5197 a_n7636_8799.t48 gnd 0.599757f
C5198 a_n7636_8799.t136 gnd 0.599757f
C5199 a_n7636_8799.n237 gnd 0.270018f
C5200 a_n7636_8799.t68 gnd 0.611109f
C5201 a_n7636_8799.n238 gnd 0.251423f
C5202 a_n7636_8799.t95 gnd 0.599757f
C5203 a_n7636_8799.n239 gnd 0.272327f
C5204 a_n7636_8799.n240 gnd 0.265774f
C5205 a_n7636_8799.n241 gnd 0.264488f
C5206 a_n7636_8799.n242 gnd 0.271697f
C5207 a_n7636_8799.n243 gnd 0.271953f
C5208 a_n7636_8799.n244 gnd 0.265131f
C5209 a_n7636_8799.n245 gnd 0.265131f
C5210 a_n7636_8799.n246 gnd 0.271953f
C5211 a_n7636_8799.n247 gnd 0.271697f
C5212 a_n7636_8799.n248 gnd 0.264488f
C5213 a_n7636_8799.n249 gnd 0.265774f
C5214 a_n7636_8799.n250 gnd 0.272327f
C5215 a_n7636_8799.n251 gnd 0.901652f
C5216 a_n7636_8799.t146 gnd 0.611098f
C5217 a_n7636_8799.t43 gnd 0.599757f
C5218 a_n7636_8799.t93 gnd 0.599757f
C5219 a_n7636_8799.n252 gnd 0.270018f
C5220 a_n7636_8799.t30 gnd 0.599757f
C5221 a_n7636_8799.t117 gnd 0.599757f
C5222 a_n7636_8799.t54 gnd 0.599757f
C5223 a_n7636_8799.n253 gnd 0.269123f
C5224 a_n7636_8799.t100 gnd 0.599757f
C5225 a_n7636_8799.t35 gnd 0.599757f
C5226 a_n7636_8799.t60 gnd 0.599757f
C5227 a_n7636_8799.n254 gnd 0.269557f
C5228 a_n7636_8799.t140 gnd 0.599757f
C5229 a_n7636_8799.t109 gnd 0.599757f
C5230 a_n7636_8799.t134 gnd 0.599757f
C5231 a_n7636_8799.n255 gnd 0.269557f
C5232 a_n7636_8799.t91 gnd 0.599757f
C5233 a_n7636_8799.t112 gnd 0.599757f
C5234 a_n7636_8799.t47 gnd 0.599757f
C5235 a_n7636_8799.n256 gnd 0.269123f
C5236 a_n7636_8799.t131 gnd 0.599757f
C5237 a_n7636_8799.t72 gnd 0.599757f
C5238 a_n7636_8799.t123 gnd 0.599757f
C5239 a_n7636_8799.n257 gnd 0.270018f
C5240 a_n7636_8799.t105 gnd 0.611109f
C5241 a_n7636_8799.n258 gnd 0.251423f
C5242 a_n7636_8799.t59 gnd 0.599757f
C5243 a_n7636_8799.n259 gnd 0.272327f
C5244 a_n7636_8799.n260 gnd 0.265774f
C5245 a_n7636_8799.n261 gnd 0.264488f
C5246 a_n7636_8799.n262 gnd 0.271697f
C5247 a_n7636_8799.n263 gnd 0.271953f
C5248 a_n7636_8799.n264 gnd 0.265131f
C5249 a_n7636_8799.n265 gnd 0.265131f
C5250 a_n7636_8799.n266 gnd 0.271953f
C5251 a_n7636_8799.n267 gnd 0.271697f
C5252 a_n7636_8799.n268 gnd 0.264488f
C5253 a_n7636_8799.n269 gnd 0.265774f
C5254 a_n7636_8799.n270 gnd 0.272327f
C5255 a_n7636_8799.n271 gnd 1.17929f
C5256 a_n7636_8799.n272 gnd 12.302401f
C5257 a_n7636_8799.n273 gnd 4.38935f
C5258 a_n7636_8799.n274 gnd 5.71736f
C5259 a_n7636_8799.t19 gnd 0.144643f
C5260 a_n7636_8799.t10 gnd 0.144643f
C5261 a_n7636_8799.n275 gnd 1.13894f
C5262 a_n7636_8799.t26 gnd 0.144643f
C5263 a_n7636_8799.t4 gnd 0.144643f
C5264 a_n7636_8799.n276 gnd 1.14082f
C5265 a_n7636_8799.n277 gnd 1.13894f
C5266 a_n7636_8799.t0 gnd 0.144643f
C5267 commonsourceibias.n0 gnd 0.012299f
C5268 commonsourceibias.t57 gnd 0.18623f
C5269 commonsourceibias.t110 gnd 0.172196f
C5270 commonsourceibias.n1 gnd 0.068706f
C5271 commonsourceibias.n2 gnd 0.009217f
C5272 commonsourceibias.t70 gnd 0.172196f
C5273 commonsourceibias.n3 gnd 0.007456f
C5274 commonsourceibias.n4 gnd 0.009217f
C5275 commonsourceibias.t117 gnd 0.172196f
C5276 commonsourceibias.n5 gnd 0.008898f
C5277 commonsourceibias.n6 gnd 0.009217f
C5278 commonsourceibias.t85 gnd 0.172196f
C5279 commonsourceibias.n7 gnd 0.068706f
C5280 commonsourceibias.t54 gnd 0.172196f
C5281 commonsourceibias.n8 gnd 0.007444f
C5282 commonsourceibias.n9 gnd 0.012299f
C5283 commonsourceibias.t20 gnd 0.18623f
C5284 commonsourceibias.t28 gnd 0.172196f
C5285 commonsourceibias.n10 gnd 0.068706f
C5286 commonsourceibias.n11 gnd 0.009217f
C5287 commonsourceibias.t0 gnd 0.172196f
C5288 commonsourceibias.n12 gnd 0.007456f
C5289 commonsourceibias.n13 gnd 0.009217f
C5290 commonsourceibias.t36 gnd 0.172196f
C5291 commonsourceibias.n14 gnd 0.008898f
C5292 commonsourceibias.n15 gnd 0.009217f
C5293 commonsourceibias.t14 gnd 0.172196f
C5294 commonsourceibias.n16 gnd 0.068706f
C5295 commonsourceibias.t22 gnd 0.172196f
C5296 commonsourceibias.n17 gnd 0.007444f
C5297 commonsourceibias.n18 gnd 0.009217f
C5298 commonsourceibias.t30 gnd 0.172196f
C5299 commonsourceibias.t12 gnd 0.172196f
C5300 commonsourceibias.n19 gnd 0.068706f
C5301 commonsourceibias.n20 gnd 0.009217f
C5302 commonsourceibias.t38 gnd 0.172196f
C5303 commonsourceibias.n21 gnd 0.068706f
C5304 commonsourceibias.n22 gnd 0.009217f
C5305 commonsourceibias.t16 gnd 0.172196f
C5306 commonsourceibias.n23 gnd 0.068706f
C5307 commonsourceibias.n24 gnd 0.046399f
C5308 commonsourceibias.t4 gnd 0.172196f
C5309 commonsourceibias.t32 gnd 0.194303f
C5310 commonsourceibias.n25 gnd 0.079733f
C5311 commonsourceibias.n26 gnd 0.082545f
C5312 commonsourceibias.n27 gnd 0.01136f
C5313 commonsourceibias.n28 gnd 0.012567f
C5314 commonsourceibias.n29 gnd 0.009217f
C5315 commonsourceibias.n30 gnd 0.009217f
C5316 commonsourceibias.n31 gnd 0.012485f
C5317 commonsourceibias.n32 gnd 0.007456f
C5318 commonsourceibias.n33 gnd 0.01264f
C5319 commonsourceibias.n34 gnd 0.009217f
C5320 commonsourceibias.n35 gnd 0.009217f
C5321 commonsourceibias.n36 gnd 0.012717f
C5322 commonsourceibias.n37 gnd 0.010966f
C5323 commonsourceibias.n38 gnd 0.008898f
C5324 commonsourceibias.n39 gnd 0.009217f
C5325 commonsourceibias.n40 gnd 0.009217f
C5326 commonsourceibias.n41 gnd 0.011274f
C5327 commonsourceibias.n42 gnd 0.012653f
C5328 commonsourceibias.n43 gnd 0.068706f
C5329 commonsourceibias.n44 gnd 0.012568f
C5330 commonsourceibias.n45 gnd 0.009217f
C5331 commonsourceibias.n46 gnd 0.009217f
C5332 commonsourceibias.n47 gnd 0.009217f
C5333 commonsourceibias.n48 gnd 0.012568f
C5334 commonsourceibias.n49 gnd 0.068706f
C5335 commonsourceibias.n50 gnd 0.012653f
C5336 commonsourceibias.n51 gnd 0.011274f
C5337 commonsourceibias.n52 gnd 0.009217f
C5338 commonsourceibias.n53 gnd 0.009217f
C5339 commonsourceibias.n54 gnd 0.009217f
C5340 commonsourceibias.n55 gnd 0.010966f
C5341 commonsourceibias.n56 gnd 0.012717f
C5342 commonsourceibias.n57 gnd 0.068706f
C5343 commonsourceibias.n58 gnd 0.01264f
C5344 commonsourceibias.n59 gnd 0.009217f
C5345 commonsourceibias.n60 gnd 0.009217f
C5346 commonsourceibias.n61 gnd 0.009217f
C5347 commonsourceibias.n62 gnd 0.012485f
C5348 commonsourceibias.n63 gnd 0.068706f
C5349 commonsourceibias.n64 gnd 0.012567f
C5350 commonsourceibias.n65 gnd 0.01136f
C5351 commonsourceibias.n66 gnd 0.009217f
C5352 commonsourceibias.n67 gnd 0.009217f
C5353 commonsourceibias.n68 gnd 0.009349f
C5354 commonsourceibias.n69 gnd 0.009666f
C5355 commonsourceibias.n70 gnd 0.082208f
C5356 commonsourceibias.n71 gnd 0.091197f
C5357 commonsourceibias.t21 gnd 0.019889f
C5358 commonsourceibias.t29 gnd 0.019889f
C5359 commonsourceibias.n72 gnd 0.175743f
C5360 commonsourceibias.n73 gnd 0.151855f
C5361 commonsourceibias.t1 gnd 0.019889f
C5362 commonsourceibias.t37 gnd 0.019889f
C5363 commonsourceibias.n74 gnd 0.175743f
C5364 commonsourceibias.n75 gnd 0.080726f
C5365 commonsourceibias.t15 gnd 0.019889f
C5366 commonsourceibias.t23 gnd 0.019889f
C5367 commonsourceibias.n76 gnd 0.175743f
C5368 commonsourceibias.n77 gnd 0.067443f
C5369 commonsourceibias.t5 gnd 0.019889f
C5370 commonsourceibias.t33 gnd 0.019889f
C5371 commonsourceibias.n78 gnd 0.176331f
C5372 commonsourceibias.t39 gnd 0.019889f
C5373 commonsourceibias.t17 gnd 0.019889f
C5374 commonsourceibias.n79 gnd 0.175743f
C5375 commonsourceibias.n80 gnd 0.16376f
C5376 commonsourceibias.t31 gnd 0.019889f
C5377 commonsourceibias.t13 gnd 0.019889f
C5378 commonsourceibias.n81 gnd 0.175743f
C5379 commonsourceibias.n82 gnd 0.067443f
C5380 commonsourceibias.n83 gnd 0.081666f
C5381 commonsourceibias.n84 gnd 0.009217f
C5382 commonsourceibias.t97 gnd 0.172196f
C5383 commonsourceibias.t86 gnd 0.172196f
C5384 commonsourceibias.n85 gnd 0.068706f
C5385 commonsourceibias.n86 gnd 0.009217f
C5386 commonsourceibias.t115 gnd 0.172196f
C5387 commonsourceibias.n87 gnd 0.068706f
C5388 commonsourceibias.n88 gnd 0.009217f
C5389 commonsourceibias.t80 gnd 0.172196f
C5390 commonsourceibias.n89 gnd 0.068706f
C5391 commonsourceibias.n90 gnd 0.046399f
C5392 commonsourceibias.t66 gnd 0.172196f
C5393 commonsourceibias.t96 gnd 0.194303f
C5394 commonsourceibias.n91 gnd 0.079733f
C5395 commonsourceibias.n92 gnd 0.082545f
C5396 commonsourceibias.n93 gnd 0.01136f
C5397 commonsourceibias.n94 gnd 0.012567f
C5398 commonsourceibias.n95 gnd 0.009217f
C5399 commonsourceibias.n96 gnd 0.009217f
C5400 commonsourceibias.n97 gnd 0.012485f
C5401 commonsourceibias.n98 gnd 0.007456f
C5402 commonsourceibias.n99 gnd 0.01264f
C5403 commonsourceibias.n100 gnd 0.009217f
C5404 commonsourceibias.n101 gnd 0.009217f
C5405 commonsourceibias.n102 gnd 0.012717f
C5406 commonsourceibias.n103 gnd 0.010966f
C5407 commonsourceibias.n104 gnd 0.008898f
C5408 commonsourceibias.n105 gnd 0.009217f
C5409 commonsourceibias.n106 gnd 0.009217f
C5410 commonsourceibias.n107 gnd 0.011274f
C5411 commonsourceibias.n108 gnd 0.012653f
C5412 commonsourceibias.n109 gnd 0.068706f
C5413 commonsourceibias.n110 gnd 0.012568f
C5414 commonsourceibias.n111 gnd 0.009172f
C5415 commonsourceibias.n112 gnd 0.066626f
C5416 commonsourceibias.n113 gnd 0.009172f
C5417 commonsourceibias.n114 gnd 0.012568f
C5418 commonsourceibias.n115 gnd 0.068706f
C5419 commonsourceibias.n116 gnd 0.012653f
C5420 commonsourceibias.n117 gnd 0.011274f
C5421 commonsourceibias.n118 gnd 0.009217f
C5422 commonsourceibias.n119 gnd 0.009217f
C5423 commonsourceibias.n120 gnd 0.009217f
C5424 commonsourceibias.n121 gnd 0.010966f
C5425 commonsourceibias.n122 gnd 0.012717f
C5426 commonsourceibias.n123 gnd 0.068706f
C5427 commonsourceibias.n124 gnd 0.01264f
C5428 commonsourceibias.n125 gnd 0.009217f
C5429 commonsourceibias.n126 gnd 0.009217f
C5430 commonsourceibias.n127 gnd 0.009217f
C5431 commonsourceibias.n128 gnd 0.012485f
C5432 commonsourceibias.n129 gnd 0.068706f
C5433 commonsourceibias.n130 gnd 0.012567f
C5434 commonsourceibias.n131 gnd 0.01136f
C5435 commonsourceibias.n132 gnd 0.009217f
C5436 commonsourceibias.n133 gnd 0.009217f
C5437 commonsourceibias.n134 gnd 0.009349f
C5438 commonsourceibias.n135 gnd 0.009666f
C5439 commonsourceibias.n136 gnd 0.082208f
C5440 commonsourceibias.n137 gnd 0.05322f
C5441 commonsourceibias.n138 gnd 0.012299f
C5442 commonsourceibias.t88 gnd 0.18623f
C5443 commonsourceibias.t105 gnd 0.172196f
C5444 commonsourceibias.n139 gnd 0.068706f
C5445 commonsourceibias.n140 gnd 0.009217f
C5446 commonsourceibias.t101 gnd 0.172196f
C5447 commonsourceibias.n141 gnd 0.007456f
C5448 commonsourceibias.n142 gnd 0.009217f
C5449 commonsourceibias.t89 gnd 0.172196f
C5450 commonsourceibias.n143 gnd 0.008898f
C5451 commonsourceibias.n144 gnd 0.009217f
C5452 commonsourceibias.t106 gnd 0.172196f
C5453 commonsourceibias.n145 gnd 0.068706f
C5454 commonsourceibias.t99 gnd 0.172196f
C5455 commonsourceibias.n146 gnd 0.007444f
C5456 commonsourceibias.n147 gnd 0.009217f
C5457 commonsourceibias.t87 gnd 0.172196f
C5458 commonsourceibias.t107 gnd 0.172196f
C5459 commonsourceibias.n148 gnd 0.068706f
C5460 commonsourceibias.n149 gnd 0.009217f
C5461 commonsourceibias.t100 gnd 0.172196f
C5462 commonsourceibias.n150 gnd 0.068706f
C5463 commonsourceibias.n151 gnd 0.009217f
C5464 commonsourceibias.t112 gnd 0.172196f
C5465 commonsourceibias.n152 gnd 0.068706f
C5466 commonsourceibias.n153 gnd 0.046399f
C5467 commonsourceibias.t108 gnd 0.172196f
C5468 commonsourceibias.t98 gnd 0.194303f
C5469 commonsourceibias.n154 gnd 0.079733f
C5470 commonsourceibias.n155 gnd 0.082545f
C5471 commonsourceibias.n156 gnd 0.01136f
C5472 commonsourceibias.n157 gnd 0.012567f
C5473 commonsourceibias.n158 gnd 0.009217f
C5474 commonsourceibias.n159 gnd 0.009217f
C5475 commonsourceibias.n160 gnd 0.012485f
C5476 commonsourceibias.n161 gnd 0.007456f
C5477 commonsourceibias.n162 gnd 0.01264f
C5478 commonsourceibias.n163 gnd 0.009217f
C5479 commonsourceibias.n164 gnd 0.009217f
C5480 commonsourceibias.n165 gnd 0.012717f
C5481 commonsourceibias.n166 gnd 0.010966f
C5482 commonsourceibias.n167 gnd 0.008898f
C5483 commonsourceibias.n168 gnd 0.009217f
C5484 commonsourceibias.n169 gnd 0.009217f
C5485 commonsourceibias.n170 gnd 0.011274f
C5486 commonsourceibias.n171 gnd 0.012653f
C5487 commonsourceibias.n172 gnd 0.068706f
C5488 commonsourceibias.n173 gnd 0.012568f
C5489 commonsourceibias.n174 gnd 0.009217f
C5490 commonsourceibias.n175 gnd 0.009217f
C5491 commonsourceibias.n176 gnd 0.009217f
C5492 commonsourceibias.n177 gnd 0.012568f
C5493 commonsourceibias.n178 gnd 0.068706f
C5494 commonsourceibias.n179 gnd 0.012653f
C5495 commonsourceibias.n180 gnd 0.011274f
C5496 commonsourceibias.n181 gnd 0.009217f
C5497 commonsourceibias.n182 gnd 0.009217f
C5498 commonsourceibias.n183 gnd 0.009217f
C5499 commonsourceibias.n184 gnd 0.010966f
C5500 commonsourceibias.n185 gnd 0.012717f
C5501 commonsourceibias.n186 gnd 0.068706f
C5502 commonsourceibias.n187 gnd 0.01264f
C5503 commonsourceibias.n188 gnd 0.009217f
C5504 commonsourceibias.n189 gnd 0.009217f
C5505 commonsourceibias.n190 gnd 0.009217f
C5506 commonsourceibias.n191 gnd 0.012485f
C5507 commonsourceibias.n192 gnd 0.068706f
C5508 commonsourceibias.n193 gnd 0.012567f
C5509 commonsourceibias.n194 gnd 0.01136f
C5510 commonsourceibias.n195 gnd 0.009217f
C5511 commonsourceibias.n196 gnd 0.009217f
C5512 commonsourceibias.n197 gnd 0.009349f
C5513 commonsourceibias.n198 gnd 0.009666f
C5514 commonsourceibias.n199 gnd 0.082208f
C5515 commonsourceibias.n200 gnd 0.027976f
C5516 commonsourceibias.n201 gnd 0.147064f
C5517 commonsourceibias.n202 gnd 0.012299f
C5518 commonsourceibias.t50 gnd 0.172196f
C5519 commonsourceibias.n203 gnd 0.068706f
C5520 commonsourceibias.n204 gnd 0.009217f
C5521 commonsourceibias.t59 gnd 0.172196f
C5522 commonsourceibias.n205 gnd 0.007456f
C5523 commonsourceibias.n206 gnd 0.009217f
C5524 commonsourceibias.t104 gnd 0.172196f
C5525 commonsourceibias.n207 gnd 0.008898f
C5526 commonsourceibias.n208 gnd 0.009217f
C5527 commonsourceibias.t119 gnd 0.172196f
C5528 commonsourceibias.n209 gnd 0.068706f
C5529 commonsourceibias.t53 gnd 0.172196f
C5530 commonsourceibias.n210 gnd 0.007444f
C5531 commonsourceibias.n211 gnd 0.009217f
C5532 commonsourceibias.t93 gnd 0.172196f
C5533 commonsourceibias.t84 gnd 0.172196f
C5534 commonsourceibias.n212 gnd 0.068706f
C5535 commonsourceibias.n213 gnd 0.009217f
C5536 commonsourceibias.t49 gnd 0.172196f
C5537 commonsourceibias.n214 gnd 0.068706f
C5538 commonsourceibias.n215 gnd 0.009217f
C5539 commonsourceibias.t60 gnd 0.172196f
C5540 commonsourceibias.n216 gnd 0.068706f
C5541 commonsourceibias.n217 gnd 0.046399f
C5542 commonsourceibias.t75 gnd 0.172196f
C5543 commonsourceibias.t118 gnd 0.194303f
C5544 commonsourceibias.n218 gnd 0.079733f
C5545 commonsourceibias.n219 gnd 0.082545f
C5546 commonsourceibias.n220 gnd 0.01136f
C5547 commonsourceibias.n221 gnd 0.012567f
C5548 commonsourceibias.n222 gnd 0.009217f
C5549 commonsourceibias.n223 gnd 0.009217f
C5550 commonsourceibias.n224 gnd 0.012485f
C5551 commonsourceibias.n225 gnd 0.007456f
C5552 commonsourceibias.n226 gnd 0.01264f
C5553 commonsourceibias.n227 gnd 0.009217f
C5554 commonsourceibias.n228 gnd 0.009217f
C5555 commonsourceibias.n229 gnd 0.012717f
C5556 commonsourceibias.n230 gnd 0.010966f
C5557 commonsourceibias.n231 gnd 0.008898f
C5558 commonsourceibias.n232 gnd 0.009217f
C5559 commonsourceibias.n233 gnd 0.009217f
C5560 commonsourceibias.n234 gnd 0.011274f
C5561 commonsourceibias.n235 gnd 0.012653f
C5562 commonsourceibias.n236 gnd 0.068706f
C5563 commonsourceibias.n237 gnd 0.012568f
C5564 commonsourceibias.n238 gnd 0.009217f
C5565 commonsourceibias.n239 gnd 0.009217f
C5566 commonsourceibias.n240 gnd 0.009217f
C5567 commonsourceibias.n241 gnd 0.012568f
C5568 commonsourceibias.n242 gnd 0.068706f
C5569 commonsourceibias.n243 gnd 0.012653f
C5570 commonsourceibias.n244 gnd 0.011274f
C5571 commonsourceibias.n245 gnd 0.009217f
C5572 commonsourceibias.n246 gnd 0.009217f
C5573 commonsourceibias.n247 gnd 0.009217f
C5574 commonsourceibias.n248 gnd 0.010966f
C5575 commonsourceibias.n249 gnd 0.012717f
C5576 commonsourceibias.n250 gnd 0.068706f
C5577 commonsourceibias.n251 gnd 0.01264f
C5578 commonsourceibias.n252 gnd 0.009217f
C5579 commonsourceibias.n253 gnd 0.009217f
C5580 commonsourceibias.n254 gnd 0.009217f
C5581 commonsourceibias.n255 gnd 0.012485f
C5582 commonsourceibias.n256 gnd 0.068706f
C5583 commonsourceibias.n257 gnd 0.012567f
C5584 commonsourceibias.n258 gnd 0.01136f
C5585 commonsourceibias.n259 gnd 0.009217f
C5586 commonsourceibias.n260 gnd 0.009217f
C5587 commonsourceibias.n261 gnd 0.009349f
C5588 commonsourceibias.n262 gnd 0.009666f
C5589 commonsourceibias.t111 gnd 0.18623f
C5590 commonsourceibias.n263 gnd 0.082208f
C5591 commonsourceibias.n264 gnd 0.027976f
C5592 commonsourceibias.n265 gnd 0.517265f
C5593 commonsourceibias.n266 gnd 0.012299f
C5594 commonsourceibias.t114 gnd 0.18623f
C5595 commonsourceibias.t78 gnd 0.172196f
C5596 commonsourceibias.n267 gnd 0.068706f
C5597 commonsourceibias.n268 gnd 0.009217f
C5598 commonsourceibias.t52 gnd 0.172196f
C5599 commonsourceibias.n269 gnd 0.007456f
C5600 commonsourceibias.n270 gnd 0.009217f
C5601 commonsourceibias.t94 gnd 0.172196f
C5602 commonsourceibias.n271 gnd 0.008898f
C5603 commonsourceibias.n272 gnd 0.009217f
C5604 commonsourceibias.t113 gnd 0.172196f
C5605 commonsourceibias.n273 gnd 0.007444f
C5606 commonsourceibias.n274 gnd 0.009217f
C5607 commonsourceibias.t76 gnd 0.172196f
C5608 commonsourceibias.t65 gnd 0.172196f
C5609 commonsourceibias.n275 gnd 0.068706f
C5610 commonsourceibias.n276 gnd 0.009217f
C5611 commonsourceibias.t92 gnd 0.172196f
C5612 commonsourceibias.n277 gnd 0.068706f
C5613 commonsourceibias.n278 gnd 0.009217f
C5614 commonsourceibias.t63 gnd 0.172196f
C5615 commonsourceibias.n279 gnd 0.068706f
C5616 commonsourceibias.n280 gnd 0.046399f
C5617 commonsourceibias.t58 gnd 0.172196f
C5618 commonsourceibias.t69 gnd 0.194303f
C5619 commonsourceibias.n281 gnd 0.079733f
C5620 commonsourceibias.n282 gnd 0.082545f
C5621 commonsourceibias.n283 gnd 0.01136f
C5622 commonsourceibias.n284 gnd 0.012567f
C5623 commonsourceibias.n285 gnd 0.009217f
C5624 commonsourceibias.n286 gnd 0.009217f
C5625 commonsourceibias.n287 gnd 0.012485f
C5626 commonsourceibias.n288 gnd 0.007456f
C5627 commonsourceibias.n289 gnd 0.01264f
C5628 commonsourceibias.n290 gnd 0.009217f
C5629 commonsourceibias.n291 gnd 0.009217f
C5630 commonsourceibias.n292 gnd 0.012717f
C5631 commonsourceibias.n293 gnd 0.010966f
C5632 commonsourceibias.n294 gnd 0.008898f
C5633 commonsourceibias.n295 gnd 0.009217f
C5634 commonsourceibias.n296 gnd 0.009217f
C5635 commonsourceibias.n297 gnd 0.011274f
C5636 commonsourceibias.n298 gnd 0.012653f
C5637 commonsourceibias.n299 gnd 0.068706f
C5638 commonsourceibias.n300 gnd 0.012568f
C5639 commonsourceibias.n301 gnd 0.009172f
C5640 commonsourceibias.t3 gnd 0.019889f
C5641 commonsourceibias.t45 gnd 0.019889f
C5642 commonsourceibias.n302 gnd 0.176331f
C5643 commonsourceibias.t27 gnd 0.019889f
C5644 commonsourceibias.t11 gnd 0.019889f
C5645 commonsourceibias.n303 gnd 0.175743f
C5646 commonsourceibias.n304 gnd 0.16376f
C5647 commonsourceibias.t7 gnd 0.019889f
C5648 commonsourceibias.t47 gnd 0.019889f
C5649 commonsourceibias.n305 gnd 0.175743f
C5650 commonsourceibias.n306 gnd 0.067443f
C5651 commonsourceibias.n307 gnd 0.012299f
C5652 commonsourceibias.t18 gnd 0.172196f
C5653 commonsourceibias.n308 gnd 0.068706f
C5654 commonsourceibias.n309 gnd 0.009217f
C5655 commonsourceibias.t24 gnd 0.172196f
C5656 commonsourceibias.n310 gnd 0.007456f
C5657 commonsourceibias.n311 gnd 0.009217f
C5658 commonsourceibias.t34 gnd 0.172196f
C5659 commonsourceibias.n312 gnd 0.008898f
C5660 commonsourceibias.n313 gnd 0.009217f
C5661 commonsourceibias.t42 gnd 0.172196f
C5662 commonsourceibias.n314 gnd 0.007444f
C5663 commonsourceibias.n315 gnd 0.009217f
C5664 commonsourceibias.t46 gnd 0.172196f
C5665 commonsourceibias.t6 gnd 0.172196f
C5666 commonsourceibias.n316 gnd 0.068706f
C5667 commonsourceibias.n317 gnd 0.009217f
C5668 commonsourceibias.t10 gnd 0.172196f
C5669 commonsourceibias.n318 gnd 0.068706f
C5670 commonsourceibias.n319 gnd 0.009217f
C5671 commonsourceibias.t26 gnd 0.172196f
C5672 commonsourceibias.n320 gnd 0.068706f
C5673 commonsourceibias.n321 gnd 0.046399f
C5674 commonsourceibias.t44 gnd 0.172196f
C5675 commonsourceibias.t2 gnd 0.194303f
C5676 commonsourceibias.n322 gnd 0.079733f
C5677 commonsourceibias.n323 gnd 0.082545f
C5678 commonsourceibias.n324 gnd 0.01136f
C5679 commonsourceibias.n325 gnd 0.012567f
C5680 commonsourceibias.n326 gnd 0.009217f
C5681 commonsourceibias.n327 gnd 0.009217f
C5682 commonsourceibias.n328 gnd 0.012485f
C5683 commonsourceibias.n329 gnd 0.007456f
C5684 commonsourceibias.n330 gnd 0.01264f
C5685 commonsourceibias.n331 gnd 0.009217f
C5686 commonsourceibias.n332 gnd 0.009217f
C5687 commonsourceibias.n333 gnd 0.012717f
C5688 commonsourceibias.n334 gnd 0.010966f
C5689 commonsourceibias.n335 gnd 0.008898f
C5690 commonsourceibias.n336 gnd 0.009217f
C5691 commonsourceibias.n337 gnd 0.009217f
C5692 commonsourceibias.n338 gnd 0.011274f
C5693 commonsourceibias.n339 gnd 0.012653f
C5694 commonsourceibias.n340 gnd 0.068706f
C5695 commonsourceibias.n341 gnd 0.012568f
C5696 commonsourceibias.n342 gnd 0.009217f
C5697 commonsourceibias.n343 gnd 0.009217f
C5698 commonsourceibias.n344 gnd 0.009217f
C5699 commonsourceibias.n345 gnd 0.012568f
C5700 commonsourceibias.n346 gnd 0.068706f
C5701 commonsourceibias.n347 gnd 0.012653f
C5702 commonsourceibias.t8 gnd 0.172196f
C5703 commonsourceibias.n348 gnd 0.068706f
C5704 commonsourceibias.n349 gnd 0.011274f
C5705 commonsourceibias.n350 gnd 0.009217f
C5706 commonsourceibias.n351 gnd 0.009217f
C5707 commonsourceibias.n352 gnd 0.009217f
C5708 commonsourceibias.n353 gnd 0.010966f
C5709 commonsourceibias.n354 gnd 0.012717f
C5710 commonsourceibias.n355 gnd 0.068706f
C5711 commonsourceibias.n356 gnd 0.01264f
C5712 commonsourceibias.n357 gnd 0.009217f
C5713 commonsourceibias.n358 gnd 0.009217f
C5714 commonsourceibias.n359 gnd 0.009217f
C5715 commonsourceibias.n360 gnd 0.012485f
C5716 commonsourceibias.n361 gnd 0.068706f
C5717 commonsourceibias.n362 gnd 0.012567f
C5718 commonsourceibias.n363 gnd 0.01136f
C5719 commonsourceibias.n364 gnd 0.009217f
C5720 commonsourceibias.n365 gnd 0.009217f
C5721 commonsourceibias.n366 gnd 0.009349f
C5722 commonsourceibias.n367 gnd 0.009666f
C5723 commonsourceibias.t40 gnd 0.18623f
C5724 commonsourceibias.n368 gnd 0.082208f
C5725 commonsourceibias.n369 gnd 0.091197f
C5726 commonsourceibias.t19 gnd 0.019889f
C5727 commonsourceibias.t41 gnd 0.019889f
C5728 commonsourceibias.n370 gnd 0.175743f
C5729 commonsourceibias.n371 gnd 0.151855f
C5730 commonsourceibias.t35 gnd 0.019889f
C5731 commonsourceibias.t25 gnd 0.019889f
C5732 commonsourceibias.n372 gnd 0.175743f
C5733 commonsourceibias.n373 gnd 0.080726f
C5734 commonsourceibias.t43 gnd 0.019889f
C5735 commonsourceibias.t9 gnd 0.019889f
C5736 commonsourceibias.n374 gnd 0.175743f
C5737 commonsourceibias.n375 gnd 0.067443f
C5738 commonsourceibias.n376 gnd 0.081666f
C5739 commonsourceibias.n377 gnd 0.066626f
C5740 commonsourceibias.n378 gnd 0.009172f
C5741 commonsourceibias.n379 gnd 0.012568f
C5742 commonsourceibias.n380 gnd 0.068706f
C5743 commonsourceibias.n381 gnd 0.012653f
C5744 commonsourceibias.t64 gnd 0.172196f
C5745 commonsourceibias.n382 gnd 0.068706f
C5746 commonsourceibias.n383 gnd 0.011274f
C5747 commonsourceibias.n384 gnd 0.009217f
C5748 commonsourceibias.n385 gnd 0.009217f
C5749 commonsourceibias.n386 gnd 0.009217f
C5750 commonsourceibias.n387 gnd 0.010966f
C5751 commonsourceibias.n388 gnd 0.012717f
C5752 commonsourceibias.n389 gnd 0.068706f
C5753 commonsourceibias.n390 gnd 0.01264f
C5754 commonsourceibias.n391 gnd 0.009217f
C5755 commonsourceibias.n392 gnd 0.009217f
C5756 commonsourceibias.n393 gnd 0.009217f
C5757 commonsourceibias.n394 gnd 0.012485f
C5758 commonsourceibias.n395 gnd 0.068706f
C5759 commonsourceibias.n396 gnd 0.012567f
C5760 commonsourceibias.n397 gnd 0.01136f
C5761 commonsourceibias.n398 gnd 0.009217f
C5762 commonsourceibias.n399 gnd 0.009217f
C5763 commonsourceibias.n400 gnd 0.009349f
C5764 commonsourceibias.n401 gnd 0.009666f
C5765 commonsourceibias.n402 gnd 0.082208f
C5766 commonsourceibias.n403 gnd 0.05322f
C5767 commonsourceibias.n404 gnd 0.012299f
C5768 commonsourceibias.t91 gnd 0.172196f
C5769 commonsourceibias.n405 gnd 0.068706f
C5770 commonsourceibias.n406 gnd 0.009217f
C5771 commonsourceibias.t82 gnd 0.172196f
C5772 commonsourceibias.n407 gnd 0.007456f
C5773 commonsourceibias.n408 gnd 0.009217f
C5774 commonsourceibias.t73 gnd 0.172196f
C5775 commonsourceibias.n409 gnd 0.008898f
C5776 commonsourceibias.n410 gnd 0.009217f
C5777 commonsourceibias.t83 gnd 0.172196f
C5778 commonsourceibias.n411 gnd 0.007444f
C5779 commonsourceibias.n412 gnd 0.009217f
C5780 commonsourceibias.t103 gnd 0.172196f
C5781 commonsourceibias.t95 gnd 0.172196f
C5782 commonsourceibias.n413 gnd 0.068706f
C5783 commonsourceibias.n414 gnd 0.009217f
C5784 commonsourceibias.t81 gnd 0.172196f
C5785 commonsourceibias.n415 gnd 0.068706f
C5786 commonsourceibias.n416 gnd 0.009217f
C5787 commonsourceibias.t102 gnd 0.172196f
C5788 commonsourceibias.n417 gnd 0.068706f
C5789 commonsourceibias.n418 gnd 0.046399f
C5790 commonsourceibias.t116 gnd 0.172196f
C5791 commonsourceibias.t79 gnd 0.194303f
C5792 commonsourceibias.n419 gnd 0.079733f
C5793 commonsourceibias.n420 gnd 0.082545f
C5794 commonsourceibias.n421 gnd 0.01136f
C5795 commonsourceibias.n422 gnd 0.012567f
C5796 commonsourceibias.n423 gnd 0.009217f
C5797 commonsourceibias.n424 gnd 0.009217f
C5798 commonsourceibias.n425 gnd 0.012485f
C5799 commonsourceibias.n426 gnd 0.007456f
C5800 commonsourceibias.n427 gnd 0.01264f
C5801 commonsourceibias.n428 gnd 0.009217f
C5802 commonsourceibias.n429 gnd 0.009217f
C5803 commonsourceibias.n430 gnd 0.012717f
C5804 commonsourceibias.n431 gnd 0.010966f
C5805 commonsourceibias.n432 gnd 0.008898f
C5806 commonsourceibias.n433 gnd 0.009217f
C5807 commonsourceibias.n434 gnd 0.009217f
C5808 commonsourceibias.n435 gnd 0.011274f
C5809 commonsourceibias.n436 gnd 0.012653f
C5810 commonsourceibias.n437 gnd 0.068706f
C5811 commonsourceibias.n438 gnd 0.012568f
C5812 commonsourceibias.n439 gnd 0.009217f
C5813 commonsourceibias.n440 gnd 0.009217f
C5814 commonsourceibias.n441 gnd 0.009217f
C5815 commonsourceibias.n442 gnd 0.012568f
C5816 commonsourceibias.n443 gnd 0.068706f
C5817 commonsourceibias.n444 gnd 0.012653f
C5818 commonsourceibias.t90 gnd 0.172196f
C5819 commonsourceibias.n445 gnd 0.068706f
C5820 commonsourceibias.n446 gnd 0.011274f
C5821 commonsourceibias.n447 gnd 0.009217f
C5822 commonsourceibias.n448 gnd 0.009217f
C5823 commonsourceibias.n449 gnd 0.009217f
C5824 commonsourceibias.n450 gnd 0.010966f
C5825 commonsourceibias.n451 gnd 0.012717f
C5826 commonsourceibias.n452 gnd 0.068706f
C5827 commonsourceibias.n453 gnd 0.01264f
C5828 commonsourceibias.n454 gnd 0.009217f
C5829 commonsourceibias.n455 gnd 0.009217f
C5830 commonsourceibias.n456 gnd 0.009217f
C5831 commonsourceibias.n457 gnd 0.012485f
C5832 commonsourceibias.n458 gnd 0.068706f
C5833 commonsourceibias.n459 gnd 0.012567f
C5834 commonsourceibias.n460 gnd 0.01136f
C5835 commonsourceibias.n461 gnd 0.009217f
C5836 commonsourceibias.n462 gnd 0.009217f
C5837 commonsourceibias.n463 gnd 0.009349f
C5838 commonsourceibias.n464 gnd 0.009666f
C5839 commonsourceibias.t74 gnd 0.18623f
C5840 commonsourceibias.n465 gnd 0.082208f
C5841 commonsourceibias.n466 gnd 0.027976f
C5842 commonsourceibias.n467 gnd 0.147064f
C5843 commonsourceibias.n468 gnd 0.012299f
C5844 commonsourceibias.t62 gnd 0.172196f
C5845 commonsourceibias.n469 gnd 0.068706f
C5846 commonsourceibias.n470 gnd 0.009217f
C5847 commonsourceibias.t71 gnd 0.172196f
C5848 commonsourceibias.n471 gnd 0.007456f
C5849 commonsourceibias.n472 gnd 0.009217f
C5850 commonsourceibias.t48 gnd 0.172196f
C5851 commonsourceibias.n473 gnd 0.008898f
C5852 commonsourceibias.n474 gnd 0.009217f
C5853 commonsourceibias.t67 gnd 0.172196f
C5854 commonsourceibias.n475 gnd 0.007444f
C5855 commonsourceibias.n476 gnd 0.009217f
C5856 commonsourceibias.t77 gnd 0.172196f
C5857 commonsourceibias.t109 gnd 0.172196f
C5858 commonsourceibias.n477 gnd 0.068706f
C5859 commonsourceibias.n478 gnd 0.009217f
C5860 commonsourceibias.t61 gnd 0.172196f
C5861 commonsourceibias.n479 gnd 0.068706f
C5862 commonsourceibias.n480 gnd 0.009217f
C5863 commonsourceibias.t72 gnd 0.172196f
C5864 commonsourceibias.n481 gnd 0.068706f
C5865 commonsourceibias.n482 gnd 0.046399f
C5866 commonsourceibias.t68 gnd 0.172196f
C5867 commonsourceibias.t55 gnd 0.194303f
C5868 commonsourceibias.n483 gnd 0.079733f
C5869 commonsourceibias.n484 gnd 0.082545f
C5870 commonsourceibias.n485 gnd 0.01136f
C5871 commonsourceibias.n486 gnd 0.012567f
C5872 commonsourceibias.n487 gnd 0.009217f
C5873 commonsourceibias.n488 gnd 0.009217f
C5874 commonsourceibias.n489 gnd 0.012485f
C5875 commonsourceibias.n490 gnd 0.007456f
C5876 commonsourceibias.n491 gnd 0.01264f
C5877 commonsourceibias.n492 gnd 0.009217f
C5878 commonsourceibias.n493 gnd 0.009217f
C5879 commonsourceibias.n494 gnd 0.012717f
C5880 commonsourceibias.n495 gnd 0.010966f
C5881 commonsourceibias.n496 gnd 0.008898f
C5882 commonsourceibias.n497 gnd 0.009217f
C5883 commonsourceibias.n498 gnd 0.009217f
C5884 commonsourceibias.n499 gnd 0.011274f
C5885 commonsourceibias.n500 gnd 0.012653f
C5886 commonsourceibias.n501 gnd 0.068706f
C5887 commonsourceibias.n502 gnd 0.012568f
C5888 commonsourceibias.n503 gnd 0.009217f
C5889 commonsourceibias.n504 gnd 0.009217f
C5890 commonsourceibias.n505 gnd 0.009217f
C5891 commonsourceibias.n506 gnd 0.012568f
C5892 commonsourceibias.n507 gnd 0.068706f
C5893 commonsourceibias.n508 gnd 0.012653f
C5894 commonsourceibias.t56 gnd 0.172196f
C5895 commonsourceibias.n509 gnd 0.068706f
C5896 commonsourceibias.n510 gnd 0.011274f
C5897 commonsourceibias.n511 gnd 0.009217f
C5898 commonsourceibias.n512 gnd 0.009217f
C5899 commonsourceibias.n513 gnd 0.009217f
C5900 commonsourceibias.n514 gnd 0.010966f
C5901 commonsourceibias.n515 gnd 0.012717f
C5902 commonsourceibias.n516 gnd 0.068706f
C5903 commonsourceibias.n517 gnd 0.01264f
C5904 commonsourceibias.n518 gnd 0.009217f
C5905 commonsourceibias.n519 gnd 0.009217f
C5906 commonsourceibias.n520 gnd 0.009217f
C5907 commonsourceibias.n521 gnd 0.012485f
C5908 commonsourceibias.n522 gnd 0.068706f
C5909 commonsourceibias.n523 gnd 0.012567f
C5910 commonsourceibias.n524 gnd 0.01136f
C5911 commonsourceibias.n525 gnd 0.009217f
C5912 commonsourceibias.n526 gnd 0.009217f
C5913 commonsourceibias.n527 gnd 0.009349f
C5914 commonsourceibias.n528 gnd 0.009666f
C5915 commonsourceibias.t51 gnd 0.18623f
C5916 commonsourceibias.n529 gnd 0.082208f
C5917 commonsourceibias.n530 gnd 0.027976f
C5918 commonsourceibias.n531 gnd 0.194274f
C5919 commonsourceibias.n532 gnd 5.09694f
.ends

