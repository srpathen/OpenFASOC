* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t45 plus.t0 drain_left.t12 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X1 source.t7 minus.t0 drain_right.t23 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X2 drain_right.t22 minus.t1 source.t18 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X3 a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=1
X4 source.t44 plus.t1 drain_left.t15 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X5 drain_left.t6 plus.t2 source.t43 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X6 source.t15 minus.t2 drain_right.t21 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X7 drain_left.t13 plus.t3 source.t42 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X8 drain_left.t10 plus.t4 source.t41 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X9 drain_right.t20 minus.t3 source.t19 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X10 drain_right.t19 minus.t4 source.t20 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X11 source.t16 minus.t5 drain_right.t18 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X12 drain_left.t21 plus.t5 source.t40 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X13 source.t39 plus.t6 drain_left.t5 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X14 drain_left.t14 plus.t7 source.t38 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X15 drain_left.t23 plus.t8 source.t37 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X16 source.t36 plus.t9 drain_left.t8 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X17 drain_right.t17 minus.t6 source.t14 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X18 source.t12 minus.t7 drain_right.t16 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X19 source.t35 plus.t10 drain_left.t1 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X20 drain_left.t11 plus.t11 source.t34 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X21 source.t33 plus.t12 drain_left.t9 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X22 drain_left.t4 plus.t13 source.t32 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X23 drain_right.t15 minus.t8 source.t21 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X24 drain_left.t19 plus.t14 source.t31 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X25 source.t30 plus.t15 drain_left.t18 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X26 source.t0 minus.t9 drain_right.t14 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X27 source.t29 plus.t16 drain_left.t22 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X28 drain_right.t13 minus.t10 source.t10 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X29 source.t28 plus.t17 drain_left.t20 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X30 source.t27 plus.t18 drain_left.t16 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X31 drain_right.t12 minus.t11 source.t8 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X32 drain_right.t11 minus.t12 source.t17 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X33 drain_left.t17 plus.t19 source.t26 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X34 source.t47 minus.t13 drain_right.t10 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X35 drain_right.t9 minus.t14 source.t46 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X36 source.t6 minus.t15 drain_right.t8 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X37 source.t13 minus.t16 drain_right.t7 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X38 drain_right.t6 minus.t17 source.t5 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X39 drain_right.t5 minus.t18 source.t4 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X40 drain_right.t4 minus.t19 source.t3 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X41 drain_left.t7 plus.t20 source.t25 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X42 drain_left.t2 plus.t21 source.t24 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X43 a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X44 a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X45 source.t11 minus.t20 drain_right.t3 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X46 source.t2 minus.t21 drain_right.t2 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X47 source.t23 plus.t22 drain_left.t0 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X48 source.t9 minus.t22 drain_right.t1 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X49 source.t1 minus.t23 drain_right.t0 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X50 a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X51 source.t22 plus.t23 drain_left.t3 a_n4174_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
R0 plus.n15 plus.t23 205.905
R1 plus.n79 plus.t19 205.905
R2 plus.n61 plus.t8 183.883
R3 plus.n124 plus.t6 183.883
R4 plus.n17 plus.n14 161.3
R5 plus.n19 plus.n18 161.3
R6 plus.n21 plus.n20 161.3
R7 plus.n22 plus.n12 161.3
R8 plus.n24 plus.n23 161.3
R9 plus.n26 plus.n25 161.3
R10 plus.n27 plus.n10 161.3
R11 plus.n29 plus.n28 161.3
R12 plus.n31 plus.n30 161.3
R13 plus.n32 plus.n8 161.3
R14 plus.n35 plus.n34 161.3
R15 plus.n36 plus.n7 161.3
R16 plus.n38 plus.n37 161.3
R17 plus.n40 plus.n6 161.3
R18 plus.n43 plus.n42 161.3
R19 plus.n44 plus.n5 161.3
R20 plus.n46 plus.n45 161.3
R21 plus.n47 plus.n4 161.3
R22 plus.n50 plus.n49 161.3
R23 plus.n51 plus.n3 161.3
R24 plus.n53 plus.n52 161.3
R25 plus.n55 plus.n2 161.3
R26 plus.n57 plus.n56 161.3
R27 plus.n59 plus.n58 161.3
R28 plus.n60 plus.n0 161.3
R29 plus.n81 plus.n78 161.3
R30 plus.n83 plus.n82 161.3
R31 plus.n85 plus.n84 161.3
R32 plus.n86 plus.n76 161.3
R33 plus.n88 plus.n87 161.3
R34 plus.n90 plus.n89 161.3
R35 plus.n91 plus.n74 161.3
R36 plus.n93 plus.n92 161.3
R37 plus.n95 plus.n94 161.3
R38 plus.n96 plus.n72 161.3
R39 plus.n99 plus.n98 161.3
R40 plus.n100 plus.n71 161.3
R41 plus.n102 plus.n101 161.3
R42 plus.n104 plus.n69 161.3
R43 plus.n106 plus.n105 161.3
R44 plus.n107 plus.n68 161.3
R45 plus.n109 plus.n108 161.3
R46 plus.n110 plus.n67 161.3
R47 plus.n113 plus.n112 161.3
R48 plus.n114 plus.n66 161.3
R49 plus.n116 plus.n115 161.3
R50 plus.n118 plus.n65 161.3
R51 plus.n120 plus.n119 161.3
R52 plus.n122 plus.n121 161.3
R53 plus.n123 plus.n63 161.3
R54 plus.n1 plus.t10 144.601
R55 plus.n54 plus.t14 144.601
R56 plus.n48 plus.t9 144.601
R57 plus.n41 plus.t11 144.601
R58 plus.n39 plus.t15 144.601
R59 plus.n33 plus.t7 144.601
R60 plus.n9 plus.t12 144.601
R61 plus.n11 plus.t4 144.601
R62 plus.n13 plus.t0 144.601
R63 plus.n16 plus.t2 144.601
R64 plus.n64 plus.t21 144.601
R65 plus.n117 plus.t1 144.601
R66 plus.n111 plus.t5 144.601
R67 plus.n70 plus.t22 144.601
R68 plus.n103 plus.t13 144.601
R69 plus.n97 plus.t18 144.601
R70 plus.n73 plus.t3 144.601
R71 plus.n75 plus.t16 144.601
R72 plus.n77 plus.t20 144.601
R73 plus.n80 plus.t17 144.601
R74 plus.n62 plus.n61 80.6037
R75 plus.n125 plus.n124 80.6037
R76 plus.n56 plus.n55 56.5617
R77 plus.n42 plus.n40 56.5617
R78 plus.n32 plus.n31 56.5617
R79 plus.n18 plus.n17 56.5617
R80 plus.n119 plus.n118 56.5617
R81 plus.n105 plus.n104 56.5617
R82 plus.n96 plus.n95 56.5617
R83 plus.n82 plus.n81 56.5617
R84 plus.n47 plus.n46 56.0773
R85 plus.n27 plus.n26 56.0773
R86 plus.n110 plus.n109 56.0773
R87 plus.n91 plus.n90 56.0773
R88 plus.n61 plus.n60 46.0096
R89 plus.n124 plus.n123 46.0096
R90 plus.n49 plus.n3 41.5458
R91 plus.n23 plus.n22 41.5458
R92 plus.n112 plus.n66 41.5458
R93 plus.n87 plus.n86 41.5458
R94 plus.n38 plus.n7 40.577
R95 plus.n34 plus.n7 40.577
R96 plus.n102 plus.n71 40.577
R97 plus.n98 plus.n71 40.577
R98 plus.n53 plus.n3 39.6083
R99 plus.n22 plus.n21 39.6083
R100 plus.n116 plus.n66 39.6083
R101 plus.n86 plus.n85 39.6083
R102 plus plus.n125 36.8517
R103 plus.n16 plus.n15 33.0515
R104 plus.n80 plus.n79 33.0515
R105 plus.n15 plus.n14 28.5514
R106 plus.n79 plus.n78 28.5514
R107 plus.n60 plus.n59 26.0455
R108 plus.n123 plus.n122 26.0455
R109 plus.n46 plus.n5 25.0767
R110 plus.n28 plus.n27 25.0767
R111 plus.n109 plus.n68 25.0767
R112 plus.n92 plus.n91 25.0767
R113 plus.n42 plus.n41 24.3464
R114 plus.n31 plus.n9 24.3464
R115 plus.n105 plus.n70 24.3464
R116 plus.n95 plus.n73 24.3464
R117 plus.n56 plus.n1 23.8546
R118 plus.n17 plus.n16 23.8546
R119 plus.n119 plus.n64 23.8546
R120 plus.n81 plus.n80 23.8546
R121 plus.n55 plus.n54 16.9689
R122 plus.n18 plus.n13 16.9689
R123 plus.n118 plus.n117 16.9689
R124 plus.n82 plus.n77 16.9689
R125 plus.n40 plus.n39 16.477
R126 plus.n33 plus.n32 16.477
R127 plus.n104 plus.n103 16.477
R128 plus.n97 plus.n96 16.477
R129 plus.n48 plus.n47 15.9852
R130 plus.n26 plus.n11 15.9852
R131 plus.n111 plus.n110 15.9852
R132 plus.n90 plus.n75 15.9852
R133 plus plus.n62 10.1828
R134 plus.n49 plus.n48 8.60764
R135 plus.n23 plus.n11 8.60764
R136 plus.n112 plus.n111 8.60764
R137 plus.n87 plus.n75 8.60764
R138 plus.n39 plus.n38 8.11581
R139 plus.n34 plus.n33 8.11581
R140 plus.n103 plus.n102 8.11581
R141 plus.n98 plus.n97 8.11581
R142 plus.n54 plus.n53 7.62397
R143 plus.n21 plus.n13 7.62397
R144 plus.n117 plus.n116 7.62397
R145 plus.n85 plus.n77 7.62397
R146 plus.n59 plus.n1 0.738255
R147 plus.n122 plus.n64 0.738255
R148 plus.n62 plus.n0 0.285035
R149 plus.n125 plus.n63 0.285035
R150 plus.n41 plus.n5 0.246418
R151 plus.n28 plus.n9 0.246418
R152 plus.n70 plus.n68 0.246418
R153 plus.n92 plus.n73 0.246418
R154 plus.n19 plus.n14 0.189894
R155 plus.n20 plus.n19 0.189894
R156 plus.n20 plus.n12 0.189894
R157 plus.n24 plus.n12 0.189894
R158 plus.n25 plus.n24 0.189894
R159 plus.n25 plus.n10 0.189894
R160 plus.n29 plus.n10 0.189894
R161 plus.n30 plus.n29 0.189894
R162 plus.n30 plus.n8 0.189894
R163 plus.n35 plus.n8 0.189894
R164 plus.n36 plus.n35 0.189894
R165 plus.n37 plus.n36 0.189894
R166 plus.n37 plus.n6 0.189894
R167 plus.n43 plus.n6 0.189894
R168 plus.n44 plus.n43 0.189894
R169 plus.n45 plus.n44 0.189894
R170 plus.n45 plus.n4 0.189894
R171 plus.n50 plus.n4 0.189894
R172 plus.n51 plus.n50 0.189894
R173 plus.n52 plus.n51 0.189894
R174 plus.n52 plus.n2 0.189894
R175 plus.n57 plus.n2 0.189894
R176 plus.n58 plus.n57 0.189894
R177 plus.n58 plus.n0 0.189894
R178 plus.n121 plus.n63 0.189894
R179 plus.n121 plus.n120 0.189894
R180 plus.n120 plus.n65 0.189894
R181 plus.n115 plus.n65 0.189894
R182 plus.n115 plus.n114 0.189894
R183 plus.n114 plus.n113 0.189894
R184 plus.n113 plus.n67 0.189894
R185 plus.n108 plus.n67 0.189894
R186 plus.n108 plus.n107 0.189894
R187 plus.n107 plus.n106 0.189894
R188 plus.n106 plus.n69 0.189894
R189 plus.n101 plus.n69 0.189894
R190 plus.n101 plus.n100 0.189894
R191 plus.n100 plus.n99 0.189894
R192 plus.n99 plus.n72 0.189894
R193 plus.n94 plus.n72 0.189894
R194 plus.n94 plus.n93 0.189894
R195 plus.n93 plus.n74 0.189894
R196 plus.n89 plus.n74 0.189894
R197 plus.n89 plus.n88 0.189894
R198 plus.n88 plus.n76 0.189894
R199 plus.n84 plus.n76 0.189894
R200 plus.n84 plus.n83 0.189894
R201 plus.n83 plus.n78 0.189894
R202 drain_left.n13 drain_left.n11 68.3374
R203 drain_left.n7 drain_left.n5 68.3372
R204 drain_left.n2 drain_left.n0 68.3372
R205 drain_left.n19 drain_left.n18 67.1908
R206 drain_left.n17 drain_left.n16 67.1908
R207 drain_left.n15 drain_left.n14 67.1908
R208 drain_left.n13 drain_left.n12 67.1908
R209 drain_left.n21 drain_left.n20 67.1907
R210 drain_left.n7 drain_left.n6 67.1907
R211 drain_left.n9 drain_left.n8 67.1907
R212 drain_left.n4 drain_left.n3 67.1907
R213 drain_left.n2 drain_left.n1 67.1907
R214 drain_left drain_left.n10 33.7139
R215 drain_left drain_left.n21 6.79977
R216 drain_left.n5 drain_left.t20 3.3005
R217 drain_left.n5 drain_left.t17 3.3005
R218 drain_left.n6 drain_left.t22 3.3005
R219 drain_left.n6 drain_left.t7 3.3005
R220 drain_left.n8 drain_left.t16 3.3005
R221 drain_left.n8 drain_left.t13 3.3005
R222 drain_left.n3 drain_left.t0 3.3005
R223 drain_left.n3 drain_left.t4 3.3005
R224 drain_left.n1 drain_left.t15 3.3005
R225 drain_left.n1 drain_left.t21 3.3005
R226 drain_left.n0 drain_left.t5 3.3005
R227 drain_left.n0 drain_left.t2 3.3005
R228 drain_left.n20 drain_left.t1 3.3005
R229 drain_left.n20 drain_left.t23 3.3005
R230 drain_left.n18 drain_left.t8 3.3005
R231 drain_left.n18 drain_left.t19 3.3005
R232 drain_left.n16 drain_left.t18 3.3005
R233 drain_left.n16 drain_left.t11 3.3005
R234 drain_left.n14 drain_left.t9 3.3005
R235 drain_left.n14 drain_left.t14 3.3005
R236 drain_left.n12 drain_left.t12 3.3005
R237 drain_left.n12 drain_left.t10 3.3005
R238 drain_left.n11 drain_left.t3 3.3005
R239 drain_left.n11 drain_left.t6 3.3005
R240 drain_left.n9 drain_left.n7 1.14705
R241 drain_left.n4 drain_left.n2 1.14705
R242 drain_left.n15 drain_left.n13 1.14705
R243 drain_left.n17 drain_left.n15 1.14705
R244 drain_left.n19 drain_left.n17 1.14705
R245 drain_left.n21 drain_left.n19 1.14705
R246 drain_left.n10 drain_left.n9 0.51843
R247 drain_left.n10 drain_left.n4 0.51843
R248 source.n290 source.n264 289.615
R249 source.n248 source.n222 289.615
R250 source.n216 source.n190 289.615
R251 source.n174 source.n148 289.615
R252 source.n26 source.n0 289.615
R253 source.n68 source.n42 289.615
R254 source.n100 source.n74 289.615
R255 source.n142 source.n116 289.615
R256 source.n275 source.n274 185
R257 source.n272 source.n271 185
R258 source.n281 source.n280 185
R259 source.n283 source.n282 185
R260 source.n268 source.n267 185
R261 source.n289 source.n288 185
R262 source.n291 source.n290 185
R263 source.n233 source.n232 185
R264 source.n230 source.n229 185
R265 source.n239 source.n238 185
R266 source.n241 source.n240 185
R267 source.n226 source.n225 185
R268 source.n247 source.n246 185
R269 source.n249 source.n248 185
R270 source.n201 source.n200 185
R271 source.n198 source.n197 185
R272 source.n207 source.n206 185
R273 source.n209 source.n208 185
R274 source.n194 source.n193 185
R275 source.n215 source.n214 185
R276 source.n217 source.n216 185
R277 source.n159 source.n158 185
R278 source.n156 source.n155 185
R279 source.n165 source.n164 185
R280 source.n167 source.n166 185
R281 source.n152 source.n151 185
R282 source.n173 source.n172 185
R283 source.n175 source.n174 185
R284 source.n27 source.n26 185
R285 source.n25 source.n24 185
R286 source.n4 source.n3 185
R287 source.n19 source.n18 185
R288 source.n17 source.n16 185
R289 source.n8 source.n7 185
R290 source.n11 source.n10 185
R291 source.n69 source.n68 185
R292 source.n67 source.n66 185
R293 source.n46 source.n45 185
R294 source.n61 source.n60 185
R295 source.n59 source.n58 185
R296 source.n50 source.n49 185
R297 source.n53 source.n52 185
R298 source.n101 source.n100 185
R299 source.n99 source.n98 185
R300 source.n78 source.n77 185
R301 source.n93 source.n92 185
R302 source.n91 source.n90 185
R303 source.n82 source.n81 185
R304 source.n85 source.n84 185
R305 source.n143 source.n142 185
R306 source.n141 source.n140 185
R307 source.n120 source.n119 185
R308 source.n135 source.n134 185
R309 source.n133 source.n132 185
R310 source.n124 source.n123 185
R311 source.n127 source.n126 185
R312 source.t8 source.n273 147.661
R313 source.t6 source.n231 147.661
R314 source.t26 source.n199 147.661
R315 source.t39 source.n157 147.661
R316 source.t37 source.n9 147.661
R317 source.t22 source.n51 147.661
R318 source.t46 source.n83 147.661
R319 source.t15 source.n125 147.661
R320 source.n274 source.n271 104.615
R321 source.n281 source.n271 104.615
R322 source.n282 source.n281 104.615
R323 source.n282 source.n267 104.615
R324 source.n289 source.n267 104.615
R325 source.n290 source.n289 104.615
R326 source.n232 source.n229 104.615
R327 source.n239 source.n229 104.615
R328 source.n240 source.n239 104.615
R329 source.n240 source.n225 104.615
R330 source.n247 source.n225 104.615
R331 source.n248 source.n247 104.615
R332 source.n200 source.n197 104.615
R333 source.n207 source.n197 104.615
R334 source.n208 source.n207 104.615
R335 source.n208 source.n193 104.615
R336 source.n215 source.n193 104.615
R337 source.n216 source.n215 104.615
R338 source.n158 source.n155 104.615
R339 source.n165 source.n155 104.615
R340 source.n166 source.n165 104.615
R341 source.n166 source.n151 104.615
R342 source.n173 source.n151 104.615
R343 source.n174 source.n173 104.615
R344 source.n26 source.n25 104.615
R345 source.n25 source.n3 104.615
R346 source.n18 source.n3 104.615
R347 source.n18 source.n17 104.615
R348 source.n17 source.n7 104.615
R349 source.n10 source.n7 104.615
R350 source.n68 source.n67 104.615
R351 source.n67 source.n45 104.615
R352 source.n60 source.n45 104.615
R353 source.n60 source.n59 104.615
R354 source.n59 source.n49 104.615
R355 source.n52 source.n49 104.615
R356 source.n100 source.n99 104.615
R357 source.n99 source.n77 104.615
R358 source.n92 source.n77 104.615
R359 source.n92 source.n91 104.615
R360 source.n91 source.n81 104.615
R361 source.n84 source.n81 104.615
R362 source.n142 source.n141 104.615
R363 source.n141 source.n119 104.615
R364 source.n134 source.n119 104.615
R365 source.n134 source.n133 104.615
R366 source.n133 source.n123 104.615
R367 source.n126 source.n123 104.615
R368 source.n274 source.t8 52.3082
R369 source.n232 source.t6 52.3082
R370 source.n200 source.t26 52.3082
R371 source.n158 source.t39 52.3082
R372 source.n10 source.t37 52.3082
R373 source.n52 source.t22 52.3082
R374 source.n84 source.t46 52.3082
R375 source.n126 source.t15 52.3082
R376 source.n33 source.n32 50.512
R377 source.n35 source.n34 50.512
R378 source.n37 source.n36 50.512
R379 source.n39 source.n38 50.512
R380 source.n41 source.n40 50.512
R381 source.n107 source.n106 50.512
R382 source.n109 source.n108 50.512
R383 source.n111 source.n110 50.512
R384 source.n113 source.n112 50.512
R385 source.n115 source.n114 50.512
R386 source.n263 source.n262 50.5119
R387 source.n261 source.n260 50.5119
R388 source.n259 source.n258 50.5119
R389 source.n257 source.n256 50.5119
R390 source.n255 source.n254 50.5119
R391 source.n189 source.n188 50.5119
R392 source.n187 source.n186 50.5119
R393 source.n185 source.n184 50.5119
R394 source.n183 source.n182 50.5119
R395 source.n181 source.n180 50.5119
R396 source.n295 source.n294 32.1853
R397 source.n253 source.n252 32.1853
R398 source.n221 source.n220 32.1853
R399 source.n179 source.n178 32.1853
R400 source.n31 source.n30 32.1853
R401 source.n73 source.n72 32.1853
R402 source.n105 source.n104 32.1853
R403 source.n147 source.n146 32.1853
R404 source.n179 source.n147 17.8888
R405 source.n275 source.n273 15.6674
R406 source.n233 source.n231 15.6674
R407 source.n201 source.n199 15.6674
R408 source.n159 source.n157 15.6674
R409 source.n11 source.n9 15.6674
R410 source.n53 source.n51 15.6674
R411 source.n85 source.n83 15.6674
R412 source.n127 source.n125 15.6674
R413 source.n276 source.n272 12.8005
R414 source.n234 source.n230 12.8005
R415 source.n202 source.n198 12.8005
R416 source.n160 source.n156 12.8005
R417 source.n12 source.n8 12.8005
R418 source.n54 source.n50 12.8005
R419 source.n86 source.n82 12.8005
R420 source.n128 source.n124 12.8005
R421 source.n296 source.n31 12.0526
R422 source.n280 source.n279 12.0247
R423 source.n238 source.n237 12.0247
R424 source.n206 source.n205 12.0247
R425 source.n164 source.n163 12.0247
R426 source.n16 source.n15 12.0247
R427 source.n58 source.n57 12.0247
R428 source.n90 source.n89 12.0247
R429 source.n132 source.n131 12.0247
R430 source.n283 source.n270 11.249
R431 source.n241 source.n228 11.249
R432 source.n209 source.n196 11.249
R433 source.n167 source.n154 11.249
R434 source.n19 source.n6 11.249
R435 source.n61 source.n48 11.249
R436 source.n93 source.n80 11.249
R437 source.n135 source.n122 11.249
R438 source.n284 source.n268 10.4732
R439 source.n242 source.n226 10.4732
R440 source.n210 source.n194 10.4732
R441 source.n168 source.n152 10.4732
R442 source.n20 source.n4 10.4732
R443 source.n62 source.n46 10.4732
R444 source.n94 source.n78 10.4732
R445 source.n136 source.n120 10.4732
R446 source.n288 source.n287 9.69747
R447 source.n246 source.n245 9.69747
R448 source.n214 source.n213 9.69747
R449 source.n172 source.n171 9.69747
R450 source.n24 source.n23 9.69747
R451 source.n66 source.n65 9.69747
R452 source.n98 source.n97 9.69747
R453 source.n140 source.n139 9.69747
R454 source.n294 source.n293 9.45567
R455 source.n252 source.n251 9.45567
R456 source.n220 source.n219 9.45567
R457 source.n178 source.n177 9.45567
R458 source.n30 source.n29 9.45567
R459 source.n72 source.n71 9.45567
R460 source.n104 source.n103 9.45567
R461 source.n146 source.n145 9.45567
R462 source.n293 source.n292 9.3005
R463 source.n266 source.n265 9.3005
R464 source.n287 source.n286 9.3005
R465 source.n285 source.n284 9.3005
R466 source.n270 source.n269 9.3005
R467 source.n279 source.n278 9.3005
R468 source.n277 source.n276 9.3005
R469 source.n251 source.n250 9.3005
R470 source.n224 source.n223 9.3005
R471 source.n245 source.n244 9.3005
R472 source.n243 source.n242 9.3005
R473 source.n228 source.n227 9.3005
R474 source.n237 source.n236 9.3005
R475 source.n235 source.n234 9.3005
R476 source.n219 source.n218 9.3005
R477 source.n192 source.n191 9.3005
R478 source.n213 source.n212 9.3005
R479 source.n211 source.n210 9.3005
R480 source.n196 source.n195 9.3005
R481 source.n205 source.n204 9.3005
R482 source.n203 source.n202 9.3005
R483 source.n177 source.n176 9.3005
R484 source.n150 source.n149 9.3005
R485 source.n171 source.n170 9.3005
R486 source.n169 source.n168 9.3005
R487 source.n154 source.n153 9.3005
R488 source.n163 source.n162 9.3005
R489 source.n161 source.n160 9.3005
R490 source.n29 source.n28 9.3005
R491 source.n2 source.n1 9.3005
R492 source.n23 source.n22 9.3005
R493 source.n21 source.n20 9.3005
R494 source.n6 source.n5 9.3005
R495 source.n15 source.n14 9.3005
R496 source.n13 source.n12 9.3005
R497 source.n71 source.n70 9.3005
R498 source.n44 source.n43 9.3005
R499 source.n65 source.n64 9.3005
R500 source.n63 source.n62 9.3005
R501 source.n48 source.n47 9.3005
R502 source.n57 source.n56 9.3005
R503 source.n55 source.n54 9.3005
R504 source.n103 source.n102 9.3005
R505 source.n76 source.n75 9.3005
R506 source.n97 source.n96 9.3005
R507 source.n95 source.n94 9.3005
R508 source.n80 source.n79 9.3005
R509 source.n89 source.n88 9.3005
R510 source.n87 source.n86 9.3005
R511 source.n145 source.n144 9.3005
R512 source.n118 source.n117 9.3005
R513 source.n139 source.n138 9.3005
R514 source.n137 source.n136 9.3005
R515 source.n122 source.n121 9.3005
R516 source.n131 source.n130 9.3005
R517 source.n129 source.n128 9.3005
R518 source.n291 source.n266 8.92171
R519 source.n249 source.n224 8.92171
R520 source.n217 source.n192 8.92171
R521 source.n175 source.n150 8.92171
R522 source.n27 source.n2 8.92171
R523 source.n69 source.n44 8.92171
R524 source.n101 source.n76 8.92171
R525 source.n143 source.n118 8.92171
R526 source.n292 source.n264 8.14595
R527 source.n250 source.n222 8.14595
R528 source.n218 source.n190 8.14595
R529 source.n176 source.n148 8.14595
R530 source.n28 source.n0 8.14595
R531 source.n70 source.n42 8.14595
R532 source.n102 source.n74 8.14595
R533 source.n144 source.n116 8.14595
R534 source.n296 source.n295 5.83671
R535 source.n294 source.n264 5.81868
R536 source.n252 source.n222 5.81868
R537 source.n220 source.n190 5.81868
R538 source.n178 source.n148 5.81868
R539 source.n30 source.n0 5.81868
R540 source.n72 source.n42 5.81868
R541 source.n104 source.n74 5.81868
R542 source.n146 source.n116 5.81868
R543 source.n292 source.n291 5.04292
R544 source.n250 source.n249 5.04292
R545 source.n218 source.n217 5.04292
R546 source.n176 source.n175 5.04292
R547 source.n28 source.n27 5.04292
R548 source.n70 source.n69 5.04292
R549 source.n102 source.n101 5.04292
R550 source.n144 source.n143 5.04292
R551 source.n277 source.n273 4.38594
R552 source.n235 source.n231 4.38594
R553 source.n203 source.n199 4.38594
R554 source.n161 source.n157 4.38594
R555 source.n13 source.n9 4.38594
R556 source.n55 source.n51 4.38594
R557 source.n87 source.n83 4.38594
R558 source.n129 source.n125 4.38594
R559 source.n288 source.n266 4.26717
R560 source.n246 source.n224 4.26717
R561 source.n214 source.n192 4.26717
R562 source.n172 source.n150 4.26717
R563 source.n24 source.n2 4.26717
R564 source.n66 source.n44 4.26717
R565 source.n98 source.n76 4.26717
R566 source.n140 source.n118 4.26717
R567 source.n287 source.n268 3.49141
R568 source.n245 source.n226 3.49141
R569 source.n213 source.n194 3.49141
R570 source.n171 source.n152 3.49141
R571 source.n23 source.n4 3.49141
R572 source.n65 source.n46 3.49141
R573 source.n97 source.n78 3.49141
R574 source.n139 source.n120 3.49141
R575 source.n262 source.t21 3.3005
R576 source.n262 source.t1 3.3005
R577 source.n260 source.t19 3.3005
R578 source.n260 source.t13 3.3005
R579 source.n258 source.t5 3.3005
R580 source.n258 source.t47 3.3005
R581 source.n256 source.t3 3.3005
R582 source.n256 source.t0 3.3005
R583 source.n254 source.t17 3.3005
R584 source.n254 source.t2 3.3005
R585 source.n188 source.t25 3.3005
R586 source.n188 source.t28 3.3005
R587 source.n186 source.t42 3.3005
R588 source.n186 source.t29 3.3005
R589 source.n184 source.t32 3.3005
R590 source.n184 source.t27 3.3005
R591 source.n182 source.t40 3.3005
R592 source.n182 source.t23 3.3005
R593 source.n180 source.t24 3.3005
R594 source.n180 source.t44 3.3005
R595 source.n32 source.t31 3.3005
R596 source.n32 source.t35 3.3005
R597 source.n34 source.t34 3.3005
R598 source.n34 source.t36 3.3005
R599 source.n36 source.t38 3.3005
R600 source.n36 source.t30 3.3005
R601 source.n38 source.t41 3.3005
R602 source.n38 source.t33 3.3005
R603 source.n40 source.t43 3.3005
R604 source.n40 source.t45 3.3005
R605 source.n106 source.t4 3.3005
R606 source.n106 source.t11 3.3005
R607 source.n108 source.t20 3.3005
R608 source.n108 source.t9 3.3005
R609 source.n110 source.t14 3.3005
R610 source.n110 source.t7 3.3005
R611 source.n112 source.t18 3.3005
R612 source.n112 source.t16 3.3005
R613 source.n114 source.t10 3.3005
R614 source.n114 source.t12 3.3005
R615 source.n284 source.n283 2.71565
R616 source.n242 source.n241 2.71565
R617 source.n210 source.n209 2.71565
R618 source.n168 source.n167 2.71565
R619 source.n20 source.n19 2.71565
R620 source.n62 source.n61 2.71565
R621 source.n94 source.n93 2.71565
R622 source.n136 source.n135 2.71565
R623 source.n280 source.n270 1.93989
R624 source.n238 source.n228 1.93989
R625 source.n206 source.n196 1.93989
R626 source.n164 source.n154 1.93989
R627 source.n16 source.n6 1.93989
R628 source.n58 source.n48 1.93989
R629 source.n90 source.n80 1.93989
R630 source.n132 source.n122 1.93989
R631 source.n279 source.n272 1.16414
R632 source.n237 source.n230 1.16414
R633 source.n205 source.n198 1.16414
R634 source.n163 source.n156 1.16414
R635 source.n15 source.n8 1.16414
R636 source.n57 source.n50 1.16414
R637 source.n89 source.n82 1.16414
R638 source.n131 source.n124 1.16414
R639 source.n147 source.n115 1.14705
R640 source.n115 source.n113 1.14705
R641 source.n113 source.n111 1.14705
R642 source.n111 source.n109 1.14705
R643 source.n109 source.n107 1.14705
R644 source.n107 source.n105 1.14705
R645 source.n73 source.n41 1.14705
R646 source.n41 source.n39 1.14705
R647 source.n39 source.n37 1.14705
R648 source.n37 source.n35 1.14705
R649 source.n35 source.n33 1.14705
R650 source.n33 source.n31 1.14705
R651 source.n181 source.n179 1.14705
R652 source.n183 source.n181 1.14705
R653 source.n185 source.n183 1.14705
R654 source.n187 source.n185 1.14705
R655 source.n189 source.n187 1.14705
R656 source.n221 source.n189 1.14705
R657 source.n255 source.n253 1.14705
R658 source.n257 source.n255 1.14705
R659 source.n259 source.n257 1.14705
R660 source.n261 source.n259 1.14705
R661 source.n263 source.n261 1.14705
R662 source.n295 source.n263 1.14705
R663 source.n105 source.n73 0.470328
R664 source.n253 source.n221 0.470328
R665 source.n276 source.n275 0.388379
R666 source.n234 source.n233 0.388379
R667 source.n202 source.n201 0.388379
R668 source.n160 source.n159 0.388379
R669 source.n12 source.n11 0.388379
R670 source.n54 source.n53 0.388379
R671 source.n86 source.n85 0.388379
R672 source.n128 source.n127 0.388379
R673 source source.n296 0.188
R674 source.n278 source.n277 0.155672
R675 source.n278 source.n269 0.155672
R676 source.n285 source.n269 0.155672
R677 source.n286 source.n285 0.155672
R678 source.n286 source.n265 0.155672
R679 source.n293 source.n265 0.155672
R680 source.n236 source.n235 0.155672
R681 source.n236 source.n227 0.155672
R682 source.n243 source.n227 0.155672
R683 source.n244 source.n243 0.155672
R684 source.n244 source.n223 0.155672
R685 source.n251 source.n223 0.155672
R686 source.n204 source.n203 0.155672
R687 source.n204 source.n195 0.155672
R688 source.n211 source.n195 0.155672
R689 source.n212 source.n211 0.155672
R690 source.n212 source.n191 0.155672
R691 source.n219 source.n191 0.155672
R692 source.n162 source.n161 0.155672
R693 source.n162 source.n153 0.155672
R694 source.n169 source.n153 0.155672
R695 source.n170 source.n169 0.155672
R696 source.n170 source.n149 0.155672
R697 source.n177 source.n149 0.155672
R698 source.n29 source.n1 0.155672
R699 source.n22 source.n1 0.155672
R700 source.n22 source.n21 0.155672
R701 source.n21 source.n5 0.155672
R702 source.n14 source.n5 0.155672
R703 source.n14 source.n13 0.155672
R704 source.n71 source.n43 0.155672
R705 source.n64 source.n43 0.155672
R706 source.n64 source.n63 0.155672
R707 source.n63 source.n47 0.155672
R708 source.n56 source.n47 0.155672
R709 source.n56 source.n55 0.155672
R710 source.n103 source.n75 0.155672
R711 source.n96 source.n75 0.155672
R712 source.n96 source.n95 0.155672
R713 source.n95 source.n79 0.155672
R714 source.n88 source.n79 0.155672
R715 source.n88 source.n87 0.155672
R716 source.n145 source.n117 0.155672
R717 source.n138 source.n117 0.155672
R718 source.n138 source.n137 0.155672
R719 source.n137 source.n121 0.155672
R720 source.n130 source.n121 0.155672
R721 source.n130 source.n129 0.155672
R722 minus.n16 minus.t14 205.905
R723 minus.n78 minus.t15 205.905
R724 minus.n61 minus.t2 183.883
R725 minus.n124 minus.t11 183.883
R726 minus.n60 minus.n0 161.3
R727 minus.n59 minus.n58 161.3
R728 minus.n57 minus.n56 161.3
R729 minus.n55 minus.n2 161.3
R730 minus.n53 minus.n52 161.3
R731 minus.n51 minus.n3 161.3
R732 minus.n50 minus.n49 161.3
R733 minus.n47 minus.n4 161.3
R734 minus.n46 minus.n45 161.3
R735 minus.n44 minus.n5 161.3
R736 minus.n43 minus.n42 161.3
R737 minus.n41 minus.n6 161.3
R738 minus.n39 minus.n38 161.3
R739 minus.n37 minus.n8 161.3
R740 minus.n36 minus.n35 161.3
R741 minus.n33 minus.n9 161.3
R742 minus.n32 minus.n31 161.3
R743 minus.n30 minus.n29 161.3
R744 minus.n28 minus.n11 161.3
R745 minus.n27 minus.n26 161.3
R746 minus.n25 minus.n24 161.3
R747 minus.n23 minus.n13 161.3
R748 minus.n22 minus.n21 161.3
R749 minus.n20 minus.n19 161.3
R750 minus.n18 minus.n15 161.3
R751 minus.n123 minus.n63 161.3
R752 minus.n122 minus.n121 161.3
R753 minus.n120 minus.n119 161.3
R754 minus.n118 minus.n65 161.3
R755 minus.n116 minus.n115 161.3
R756 minus.n114 minus.n66 161.3
R757 minus.n113 minus.n112 161.3
R758 minus.n110 minus.n67 161.3
R759 minus.n109 minus.n108 161.3
R760 minus.n107 minus.n68 161.3
R761 minus.n106 minus.n105 161.3
R762 minus.n103 minus.n69 161.3
R763 minus.n101 minus.n100 161.3
R764 minus.n99 minus.n70 161.3
R765 minus.n98 minus.n97 161.3
R766 minus.n95 minus.n71 161.3
R767 minus.n94 minus.n93 161.3
R768 minus.n92 minus.n91 161.3
R769 minus.n90 minus.n73 161.3
R770 minus.n89 minus.n88 161.3
R771 minus.n87 minus.n86 161.3
R772 minus.n85 minus.n75 161.3
R773 minus.n84 minus.n83 161.3
R774 minus.n82 minus.n81 161.3
R775 minus.n80 minus.n77 161.3
R776 minus.n17 minus.t20 144.601
R777 minus.n14 minus.t18 144.601
R778 minus.n12 minus.t22 144.601
R779 minus.n10 minus.t4 144.601
R780 minus.n34 minus.t0 144.601
R781 minus.n40 minus.t6 144.601
R782 minus.n7 minus.t5 144.601
R783 minus.n48 minus.t1 144.601
R784 minus.n54 minus.t7 144.601
R785 minus.n1 minus.t10 144.601
R786 minus.n79 minus.t12 144.601
R787 minus.n76 minus.t21 144.601
R788 minus.n74 minus.t19 144.601
R789 minus.n72 minus.t9 144.601
R790 minus.n96 minus.t17 144.601
R791 minus.n102 minus.t13 144.601
R792 minus.n104 minus.t3 144.601
R793 minus.n111 minus.t16 144.601
R794 minus.n117 minus.t8 144.601
R795 minus.n64 minus.t23 144.601
R796 minus.n62 minus.n61 80.6037
R797 minus.n125 minus.n124 80.6037
R798 minus.n19 minus.n18 56.5617
R799 minus.n33 minus.n32 56.5617
R800 minus.n42 minus.n41 56.5617
R801 minus.n56 minus.n55 56.5617
R802 minus.n81 minus.n80 56.5617
R803 minus.n95 minus.n94 56.5617
R804 minus.n105 minus.n103 56.5617
R805 minus.n119 minus.n118 56.5617
R806 minus.n28 minus.n27 56.0773
R807 minus.n47 minus.n46 56.0773
R808 minus.n90 minus.n89 56.0773
R809 minus.n110 minus.n109 56.0773
R810 minus.n61 minus.n60 46.0096
R811 minus.n124 minus.n123 46.0096
R812 minus.n24 minus.n23 41.5458
R813 minus.n49 minus.n3 41.5458
R814 minus.n86 minus.n85 41.5458
R815 minus.n112 minus.n66 41.5458
R816 minus.n126 minus.n62 40.6979
R817 minus.n35 minus.n8 40.577
R818 minus.n39 minus.n8 40.577
R819 minus.n97 minus.n70 40.577
R820 minus.n101 minus.n70 40.577
R821 minus.n23 minus.n22 39.6083
R822 minus.n53 minus.n3 39.6083
R823 minus.n85 minus.n84 39.6083
R824 minus.n116 minus.n66 39.6083
R825 minus.n17 minus.n16 33.0515
R826 minus.n79 minus.n78 33.0515
R827 minus.n16 minus.n15 28.5514
R828 minus.n78 minus.n77 28.5514
R829 minus.n60 minus.n59 26.0455
R830 minus.n123 minus.n122 26.0455
R831 minus.n29 minus.n28 25.0767
R832 minus.n46 minus.n5 25.0767
R833 minus.n91 minus.n90 25.0767
R834 minus.n109 minus.n68 25.0767
R835 minus.n32 minus.n10 24.3464
R836 minus.n42 minus.n7 24.3464
R837 minus.n94 minus.n72 24.3464
R838 minus.n105 minus.n104 24.3464
R839 minus.n18 minus.n17 23.8546
R840 minus.n56 minus.n1 23.8546
R841 minus.n80 minus.n79 23.8546
R842 minus.n119 minus.n64 23.8546
R843 minus.n19 minus.n14 16.9689
R844 minus.n55 minus.n54 16.9689
R845 minus.n81 minus.n76 16.9689
R846 minus.n118 minus.n117 16.9689
R847 minus.n34 minus.n33 16.477
R848 minus.n41 minus.n40 16.477
R849 minus.n96 minus.n95 16.477
R850 minus.n103 minus.n102 16.477
R851 minus.n27 minus.n12 15.9852
R852 minus.n48 minus.n47 15.9852
R853 minus.n89 minus.n74 15.9852
R854 minus.n111 minus.n110 15.9852
R855 minus.n24 minus.n12 8.60764
R856 minus.n49 minus.n48 8.60764
R857 minus.n86 minus.n74 8.60764
R858 minus.n112 minus.n111 8.60764
R859 minus.n35 minus.n34 8.11581
R860 minus.n40 minus.n39 8.11581
R861 minus.n97 minus.n96 8.11581
R862 minus.n102 minus.n101 8.11581
R863 minus.n22 minus.n14 7.62397
R864 minus.n54 minus.n53 7.62397
R865 minus.n84 minus.n76 7.62397
R866 minus.n117 minus.n116 7.62397
R867 minus.n126 minus.n125 6.81155
R868 minus.n59 minus.n1 0.738255
R869 minus.n122 minus.n64 0.738255
R870 minus.n62 minus.n0 0.285035
R871 minus.n125 minus.n63 0.285035
R872 minus.n29 minus.n10 0.246418
R873 minus.n7 minus.n5 0.246418
R874 minus.n91 minus.n72 0.246418
R875 minus.n104 minus.n68 0.246418
R876 minus.n58 minus.n0 0.189894
R877 minus.n58 minus.n57 0.189894
R878 minus.n57 minus.n2 0.189894
R879 minus.n52 minus.n2 0.189894
R880 minus.n52 minus.n51 0.189894
R881 minus.n51 minus.n50 0.189894
R882 minus.n50 minus.n4 0.189894
R883 minus.n45 minus.n4 0.189894
R884 minus.n45 minus.n44 0.189894
R885 minus.n44 minus.n43 0.189894
R886 minus.n43 minus.n6 0.189894
R887 minus.n38 minus.n6 0.189894
R888 minus.n38 minus.n37 0.189894
R889 minus.n37 minus.n36 0.189894
R890 minus.n36 minus.n9 0.189894
R891 minus.n31 minus.n9 0.189894
R892 minus.n31 minus.n30 0.189894
R893 minus.n30 minus.n11 0.189894
R894 minus.n26 minus.n11 0.189894
R895 minus.n26 minus.n25 0.189894
R896 minus.n25 minus.n13 0.189894
R897 minus.n21 minus.n13 0.189894
R898 minus.n21 minus.n20 0.189894
R899 minus.n20 minus.n15 0.189894
R900 minus.n82 minus.n77 0.189894
R901 minus.n83 minus.n82 0.189894
R902 minus.n83 minus.n75 0.189894
R903 minus.n87 minus.n75 0.189894
R904 minus.n88 minus.n87 0.189894
R905 minus.n88 minus.n73 0.189894
R906 minus.n92 minus.n73 0.189894
R907 minus.n93 minus.n92 0.189894
R908 minus.n93 minus.n71 0.189894
R909 minus.n98 minus.n71 0.189894
R910 minus.n99 minus.n98 0.189894
R911 minus.n100 minus.n99 0.189894
R912 minus.n100 minus.n69 0.189894
R913 minus.n106 minus.n69 0.189894
R914 minus.n107 minus.n106 0.189894
R915 minus.n108 minus.n107 0.189894
R916 minus.n108 minus.n67 0.189894
R917 minus.n113 minus.n67 0.189894
R918 minus.n114 minus.n113 0.189894
R919 minus.n115 minus.n114 0.189894
R920 minus.n115 minus.n65 0.189894
R921 minus.n120 minus.n65 0.189894
R922 minus.n121 minus.n120 0.189894
R923 minus.n121 minus.n63 0.189894
R924 minus minus.n126 0.188
R925 drain_right.n7 drain_right.n5 68.3372
R926 drain_right.n2 drain_right.n0 68.3372
R927 drain_right.n13 drain_right.n11 68.3372
R928 drain_right.n13 drain_right.n12 67.1908
R929 drain_right.n15 drain_right.n14 67.1908
R930 drain_right.n17 drain_right.n16 67.1908
R931 drain_right.n19 drain_right.n18 67.1908
R932 drain_right.n21 drain_right.n20 67.1908
R933 drain_right.n7 drain_right.n6 67.1907
R934 drain_right.n9 drain_right.n8 67.1907
R935 drain_right.n4 drain_right.n3 67.1907
R936 drain_right.n2 drain_right.n1 67.1907
R937 drain_right drain_right.n10 33.1606
R938 drain_right drain_right.n21 6.79977
R939 drain_right.n5 drain_right.t0 3.3005
R940 drain_right.n5 drain_right.t12 3.3005
R941 drain_right.n6 drain_right.t7 3.3005
R942 drain_right.n6 drain_right.t15 3.3005
R943 drain_right.n8 drain_right.t10 3.3005
R944 drain_right.n8 drain_right.t20 3.3005
R945 drain_right.n3 drain_right.t14 3.3005
R946 drain_right.n3 drain_right.t6 3.3005
R947 drain_right.n1 drain_right.t2 3.3005
R948 drain_right.n1 drain_right.t4 3.3005
R949 drain_right.n0 drain_right.t8 3.3005
R950 drain_right.n0 drain_right.t11 3.3005
R951 drain_right.n11 drain_right.t3 3.3005
R952 drain_right.n11 drain_right.t9 3.3005
R953 drain_right.n12 drain_right.t1 3.3005
R954 drain_right.n12 drain_right.t5 3.3005
R955 drain_right.n14 drain_right.t23 3.3005
R956 drain_right.n14 drain_right.t19 3.3005
R957 drain_right.n16 drain_right.t18 3.3005
R958 drain_right.n16 drain_right.t17 3.3005
R959 drain_right.n18 drain_right.t16 3.3005
R960 drain_right.n18 drain_right.t22 3.3005
R961 drain_right.n20 drain_right.t21 3.3005
R962 drain_right.n20 drain_right.t13 3.3005
R963 drain_right.n9 drain_right.n7 1.14705
R964 drain_right.n4 drain_right.n2 1.14705
R965 drain_right.n21 drain_right.n19 1.14705
R966 drain_right.n19 drain_right.n17 1.14705
R967 drain_right.n17 drain_right.n15 1.14705
R968 drain_right.n15 drain_right.n13 1.14705
R969 drain_right.n10 drain_right.n9 0.51843
R970 drain_right.n10 drain_right.n4 0.51843
C0 drain_right source 14.663401f
C1 plus drain_left 9.81417f
C2 minus plus 7.245201f
C3 minus drain_left 0.176388f
C4 plus source 10.430599f
C5 source drain_left 14.6592f
C6 minus source 10.416599f
C7 plus drain_right 0.582226f
C8 drain_right drain_left 2.34071f
C9 minus drain_right 9.392559f
C10 drain_right a_n4174_n2088# 7.77518f
C11 drain_left a_n4174_n2088# 8.353439f
C12 source a_n4174_n2088# 6.248529f
C13 minus a_n4174_n2088# 16.520988f
C14 plus a_n4174_n2088# 18.082079f
C15 drain_right.t8 a_n4174_n2088# 0.13356f
C16 drain_right.t11 a_n4174_n2088# 0.13356f
C17 drain_right.n0 a_n4174_n2088# 1.12141f
C18 drain_right.t2 a_n4174_n2088# 0.13356f
C19 drain_right.t4 a_n4174_n2088# 0.13356f
C20 drain_right.n1 a_n4174_n2088# 1.11389f
C21 drain_right.n2 a_n4174_n2088# 0.877362f
C22 drain_right.t14 a_n4174_n2088# 0.13356f
C23 drain_right.t6 a_n4174_n2088# 0.13356f
C24 drain_right.n3 a_n4174_n2088# 1.11389f
C25 drain_right.n4 a_n4174_n2088# 0.38097f
C26 drain_right.t0 a_n4174_n2088# 0.13356f
C27 drain_right.t12 a_n4174_n2088# 0.13356f
C28 drain_right.n5 a_n4174_n2088# 1.12141f
C29 drain_right.t7 a_n4174_n2088# 0.13356f
C30 drain_right.t15 a_n4174_n2088# 0.13356f
C31 drain_right.n6 a_n4174_n2088# 1.11389f
C32 drain_right.n7 a_n4174_n2088# 0.877362f
C33 drain_right.t10 a_n4174_n2088# 0.13356f
C34 drain_right.t20 a_n4174_n2088# 0.13356f
C35 drain_right.n8 a_n4174_n2088# 1.11389f
C36 drain_right.n9 a_n4174_n2088# 0.38097f
C37 drain_right.n10 a_n4174_n2088# 1.67308f
C38 drain_right.t3 a_n4174_n2088# 0.13356f
C39 drain_right.t9 a_n4174_n2088# 0.13356f
C40 drain_right.n11 a_n4174_n2088# 1.12141f
C41 drain_right.t1 a_n4174_n2088# 0.13356f
C42 drain_right.t5 a_n4174_n2088# 0.13356f
C43 drain_right.n12 a_n4174_n2088# 1.1139f
C44 drain_right.n13 a_n4174_n2088# 0.877357f
C45 drain_right.t23 a_n4174_n2088# 0.13356f
C46 drain_right.t19 a_n4174_n2088# 0.13356f
C47 drain_right.n14 a_n4174_n2088# 1.1139f
C48 drain_right.n15 a_n4174_n2088# 0.436762f
C49 drain_right.t18 a_n4174_n2088# 0.13356f
C50 drain_right.t17 a_n4174_n2088# 0.13356f
C51 drain_right.n16 a_n4174_n2088# 1.1139f
C52 drain_right.n17 a_n4174_n2088# 0.436762f
C53 drain_right.t16 a_n4174_n2088# 0.13356f
C54 drain_right.t22 a_n4174_n2088# 0.13356f
C55 drain_right.n18 a_n4174_n2088# 1.1139f
C56 drain_right.n19 a_n4174_n2088# 0.436762f
C57 drain_right.t21 a_n4174_n2088# 0.13356f
C58 drain_right.t13 a_n4174_n2088# 0.13356f
C59 drain_right.n20 a_n4174_n2088# 1.1139f
C60 drain_right.n21 a_n4174_n2088# 0.695958f
C61 minus.n0 a_n4174_n2088# 0.04651f
C62 minus.t10 a_n4174_n2088# 0.553526f
C63 minus.n1 a_n4174_n2088# 0.227271f
C64 minus.n2 a_n4174_n2088# 0.034855f
C65 minus.t7 a_n4174_n2088# 0.553526f
C66 minus.n3 a_n4174_n2088# 0.028196f
C67 minus.n4 a_n4174_n2088# 0.034855f
C68 minus.t1 a_n4174_n2088# 0.553526f
C69 minus.n5 a_n4174_n2088# 0.03365f
C70 minus.n6 a_n4174_n2088# 0.034855f
C71 minus.t5 a_n4174_n2088# 0.553526f
C72 minus.n7 a_n4174_n2088# 0.227271f
C73 minus.t6 a_n4174_n2088# 0.553526f
C74 minus.n8 a_n4174_n2088# 0.028152f
C75 minus.n9 a_n4174_n2088# 0.034855f
C76 minus.t0 a_n4174_n2088# 0.553526f
C77 minus.t4 a_n4174_n2088# 0.553526f
C78 minus.n10 a_n4174_n2088# 0.227271f
C79 minus.n11 a_n4174_n2088# 0.034855f
C80 minus.t22 a_n4174_n2088# 0.553526f
C81 minus.n12 a_n4174_n2088# 0.227271f
C82 minus.n13 a_n4174_n2088# 0.034855f
C83 minus.t18 a_n4174_n2088# 0.553526f
C84 minus.n14 a_n4174_n2088# 0.227271f
C85 minus.n15 a_n4174_n2088# 0.175471f
C86 minus.t20 a_n4174_n2088# 0.553526f
C87 minus.t14 a_n4174_n2088# 0.637223f
C88 minus.n16 a_n4174_n2088# 0.268882f
C89 minus.n17 a_n4174_n2088# 0.279607f
C90 minus.n18 a_n4174_n2088# 0.04296f
C91 minus.n19 a_n4174_n2088# 0.047526f
C92 minus.n20 a_n4174_n2088# 0.034855f
C93 minus.n21 a_n4174_n2088# 0.034855f
C94 minus.n22 a_n4174_n2088# 0.047216f
C95 minus.n23 a_n4174_n2088# 0.028196f
C96 minus.n24 a_n4174_n2088# 0.047801f
C97 minus.n25 a_n4174_n2088# 0.034855f
C98 minus.n26 a_n4174_n2088# 0.034855f
C99 minus.n27 a_n4174_n2088# 0.048093f
C100 minus.n28 a_n4174_n2088# 0.04147f
C101 minus.n29 a_n4174_n2088# 0.03365f
C102 minus.n30 a_n4174_n2088# 0.034855f
C103 minus.n31 a_n4174_n2088# 0.034855f
C104 minus.n32 a_n4174_n2088# 0.042634f
C105 minus.n33 a_n4174_n2088# 0.047853f
C106 minus.n34 a_n4174_n2088# 0.227271f
C107 minus.n35 a_n4174_n2088# 0.047531f
C108 minus.n36 a_n4174_n2088# 0.034855f
C109 minus.n37 a_n4174_n2088# 0.034855f
C110 minus.n38 a_n4174_n2088# 0.034855f
C111 minus.n39 a_n4174_n2088# 0.047531f
C112 minus.n40 a_n4174_n2088# 0.227271f
C113 minus.n41 a_n4174_n2088# 0.047853f
C114 minus.n42 a_n4174_n2088# 0.042634f
C115 minus.n43 a_n4174_n2088# 0.034855f
C116 minus.n44 a_n4174_n2088# 0.034855f
C117 minus.n45 a_n4174_n2088# 0.034855f
C118 minus.n46 a_n4174_n2088# 0.04147f
C119 minus.n47 a_n4174_n2088# 0.048093f
C120 minus.n48 a_n4174_n2088# 0.227271f
C121 minus.n49 a_n4174_n2088# 0.047801f
C122 minus.n50 a_n4174_n2088# 0.034855f
C123 minus.n51 a_n4174_n2088# 0.034855f
C124 minus.n52 a_n4174_n2088# 0.034855f
C125 minus.n53 a_n4174_n2088# 0.047216f
C126 minus.n54 a_n4174_n2088# 0.227271f
C127 minus.n55 a_n4174_n2088# 0.047526f
C128 minus.n56 a_n4174_n2088# 0.04296f
C129 minus.n57 a_n4174_n2088# 0.034855f
C130 minus.n58 a_n4174_n2088# 0.034855f
C131 minus.n59 a_n4174_n2088# 0.035358f
C132 minus.n60 a_n4174_n2088# 0.036553f
C133 minus.t2 a_n4174_n2088# 0.6066f
C134 minus.n61 a_n4174_n2088# 0.27833f
C135 minus.n62 a_n4174_n2088# 1.49307f
C136 minus.n63 a_n4174_n2088# 0.04651f
C137 minus.t23 a_n4174_n2088# 0.553526f
C138 minus.n64 a_n4174_n2088# 0.227271f
C139 minus.n65 a_n4174_n2088# 0.034855f
C140 minus.t8 a_n4174_n2088# 0.553526f
C141 minus.n66 a_n4174_n2088# 0.028196f
C142 minus.n67 a_n4174_n2088# 0.034855f
C143 minus.t16 a_n4174_n2088# 0.553526f
C144 minus.n68 a_n4174_n2088# 0.03365f
C145 minus.n69 a_n4174_n2088# 0.034855f
C146 minus.t13 a_n4174_n2088# 0.553526f
C147 minus.n70 a_n4174_n2088# 0.028152f
C148 minus.n71 a_n4174_n2088# 0.034855f
C149 minus.t17 a_n4174_n2088# 0.553526f
C150 minus.t9 a_n4174_n2088# 0.553526f
C151 minus.n72 a_n4174_n2088# 0.227271f
C152 minus.n73 a_n4174_n2088# 0.034855f
C153 minus.t19 a_n4174_n2088# 0.553526f
C154 minus.n74 a_n4174_n2088# 0.227271f
C155 minus.n75 a_n4174_n2088# 0.034855f
C156 minus.t21 a_n4174_n2088# 0.553526f
C157 minus.n76 a_n4174_n2088# 0.227271f
C158 minus.n77 a_n4174_n2088# 0.175471f
C159 minus.t12 a_n4174_n2088# 0.553526f
C160 minus.t15 a_n4174_n2088# 0.637223f
C161 minus.n78 a_n4174_n2088# 0.268882f
C162 minus.n79 a_n4174_n2088# 0.279607f
C163 minus.n80 a_n4174_n2088# 0.04296f
C164 minus.n81 a_n4174_n2088# 0.047526f
C165 minus.n82 a_n4174_n2088# 0.034855f
C166 minus.n83 a_n4174_n2088# 0.034855f
C167 minus.n84 a_n4174_n2088# 0.047216f
C168 minus.n85 a_n4174_n2088# 0.028196f
C169 minus.n86 a_n4174_n2088# 0.047801f
C170 minus.n87 a_n4174_n2088# 0.034855f
C171 minus.n88 a_n4174_n2088# 0.034855f
C172 minus.n89 a_n4174_n2088# 0.048093f
C173 minus.n90 a_n4174_n2088# 0.04147f
C174 minus.n91 a_n4174_n2088# 0.03365f
C175 minus.n92 a_n4174_n2088# 0.034855f
C176 minus.n93 a_n4174_n2088# 0.034855f
C177 minus.n94 a_n4174_n2088# 0.042634f
C178 minus.n95 a_n4174_n2088# 0.047853f
C179 minus.n96 a_n4174_n2088# 0.227271f
C180 minus.n97 a_n4174_n2088# 0.047531f
C181 minus.n98 a_n4174_n2088# 0.034855f
C182 minus.n99 a_n4174_n2088# 0.034855f
C183 minus.n100 a_n4174_n2088# 0.034855f
C184 minus.n101 a_n4174_n2088# 0.047531f
C185 minus.n102 a_n4174_n2088# 0.227271f
C186 minus.n103 a_n4174_n2088# 0.047853f
C187 minus.t3 a_n4174_n2088# 0.553526f
C188 minus.n104 a_n4174_n2088# 0.227271f
C189 minus.n105 a_n4174_n2088# 0.042634f
C190 minus.n106 a_n4174_n2088# 0.034855f
C191 minus.n107 a_n4174_n2088# 0.034855f
C192 minus.n108 a_n4174_n2088# 0.034855f
C193 minus.n109 a_n4174_n2088# 0.04147f
C194 minus.n110 a_n4174_n2088# 0.048093f
C195 minus.n111 a_n4174_n2088# 0.227271f
C196 minus.n112 a_n4174_n2088# 0.047801f
C197 minus.n113 a_n4174_n2088# 0.034855f
C198 minus.n114 a_n4174_n2088# 0.034855f
C199 minus.n115 a_n4174_n2088# 0.034855f
C200 minus.n116 a_n4174_n2088# 0.047216f
C201 minus.n117 a_n4174_n2088# 0.227271f
C202 minus.n118 a_n4174_n2088# 0.047526f
C203 minus.n119 a_n4174_n2088# 0.04296f
C204 minus.n120 a_n4174_n2088# 0.034855f
C205 minus.n121 a_n4174_n2088# 0.034855f
C206 minus.n122 a_n4174_n2088# 0.035358f
C207 minus.n123 a_n4174_n2088# 0.036553f
C208 minus.t11 a_n4174_n2088# 0.6066f
C209 minus.n124 a_n4174_n2088# 0.27833f
C210 minus.n125 a_n4174_n2088# 0.265241f
C211 minus.n126 a_n4174_n2088# 1.76893f
C212 source.n0 a_n4174_n2088# 0.03673f
C213 source.n1 a_n4174_n2088# 0.026132f
C214 source.n2 a_n4174_n2088# 0.014042f
C215 source.n3 a_n4174_n2088# 0.03319f
C216 source.n4 a_n4174_n2088# 0.014868f
C217 source.n5 a_n4174_n2088# 0.026132f
C218 source.n6 a_n4174_n2088# 0.014042f
C219 source.n7 a_n4174_n2088# 0.03319f
C220 source.n8 a_n4174_n2088# 0.014868f
C221 source.n9 a_n4174_n2088# 0.111825f
C222 source.t37 a_n4174_n2088# 0.054096f
C223 source.n10 a_n4174_n2088# 0.024893f
C224 source.n11 a_n4174_n2088# 0.019605f
C225 source.n12 a_n4174_n2088# 0.014042f
C226 source.n13 a_n4174_n2088# 0.621778f
C227 source.n14 a_n4174_n2088# 0.026132f
C228 source.n15 a_n4174_n2088# 0.014042f
C229 source.n16 a_n4174_n2088# 0.014868f
C230 source.n17 a_n4174_n2088# 0.03319f
C231 source.n18 a_n4174_n2088# 0.03319f
C232 source.n19 a_n4174_n2088# 0.014868f
C233 source.n20 a_n4174_n2088# 0.014042f
C234 source.n21 a_n4174_n2088# 0.026132f
C235 source.n22 a_n4174_n2088# 0.026132f
C236 source.n23 a_n4174_n2088# 0.014042f
C237 source.n24 a_n4174_n2088# 0.014868f
C238 source.n25 a_n4174_n2088# 0.03319f
C239 source.n26 a_n4174_n2088# 0.071851f
C240 source.n27 a_n4174_n2088# 0.014868f
C241 source.n28 a_n4174_n2088# 0.014042f
C242 source.n29 a_n4174_n2088# 0.060402f
C243 source.n30 a_n4174_n2088# 0.040204f
C244 source.n31 a_n4174_n2088# 0.719806f
C245 source.t31 a_n4174_n2088# 0.1239f
C246 source.t35 a_n4174_n2088# 0.1239f
C247 source.n32 a_n4174_n2088# 0.964945f
C248 source.n33 a_n4174_n2088# 0.438043f
C249 source.t34 a_n4174_n2088# 0.1239f
C250 source.t36 a_n4174_n2088# 0.1239f
C251 source.n34 a_n4174_n2088# 0.964945f
C252 source.n35 a_n4174_n2088# 0.438043f
C253 source.t38 a_n4174_n2088# 0.1239f
C254 source.t30 a_n4174_n2088# 0.1239f
C255 source.n36 a_n4174_n2088# 0.964945f
C256 source.n37 a_n4174_n2088# 0.438043f
C257 source.t41 a_n4174_n2088# 0.1239f
C258 source.t33 a_n4174_n2088# 0.1239f
C259 source.n38 a_n4174_n2088# 0.964945f
C260 source.n39 a_n4174_n2088# 0.438043f
C261 source.t43 a_n4174_n2088# 0.1239f
C262 source.t45 a_n4174_n2088# 0.1239f
C263 source.n40 a_n4174_n2088# 0.964945f
C264 source.n41 a_n4174_n2088# 0.438043f
C265 source.n42 a_n4174_n2088# 0.03673f
C266 source.n43 a_n4174_n2088# 0.026132f
C267 source.n44 a_n4174_n2088# 0.014042f
C268 source.n45 a_n4174_n2088# 0.03319f
C269 source.n46 a_n4174_n2088# 0.014868f
C270 source.n47 a_n4174_n2088# 0.026132f
C271 source.n48 a_n4174_n2088# 0.014042f
C272 source.n49 a_n4174_n2088# 0.03319f
C273 source.n50 a_n4174_n2088# 0.014868f
C274 source.n51 a_n4174_n2088# 0.111825f
C275 source.t22 a_n4174_n2088# 0.054096f
C276 source.n52 a_n4174_n2088# 0.024893f
C277 source.n53 a_n4174_n2088# 0.019605f
C278 source.n54 a_n4174_n2088# 0.014042f
C279 source.n55 a_n4174_n2088# 0.621778f
C280 source.n56 a_n4174_n2088# 0.026132f
C281 source.n57 a_n4174_n2088# 0.014042f
C282 source.n58 a_n4174_n2088# 0.014868f
C283 source.n59 a_n4174_n2088# 0.03319f
C284 source.n60 a_n4174_n2088# 0.03319f
C285 source.n61 a_n4174_n2088# 0.014868f
C286 source.n62 a_n4174_n2088# 0.014042f
C287 source.n63 a_n4174_n2088# 0.026132f
C288 source.n64 a_n4174_n2088# 0.026132f
C289 source.n65 a_n4174_n2088# 0.014042f
C290 source.n66 a_n4174_n2088# 0.014868f
C291 source.n67 a_n4174_n2088# 0.03319f
C292 source.n68 a_n4174_n2088# 0.071851f
C293 source.n69 a_n4174_n2088# 0.014868f
C294 source.n70 a_n4174_n2088# 0.014042f
C295 source.n71 a_n4174_n2088# 0.060402f
C296 source.n72 a_n4174_n2088# 0.040204f
C297 source.n73 a_n4174_n2088# 0.158421f
C298 source.n74 a_n4174_n2088# 0.03673f
C299 source.n75 a_n4174_n2088# 0.026132f
C300 source.n76 a_n4174_n2088# 0.014042f
C301 source.n77 a_n4174_n2088# 0.03319f
C302 source.n78 a_n4174_n2088# 0.014868f
C303 source.n79 a_n4174_n2088# 0.026132f
C304 source.n80 a_n4174_n2088# 0.014042f
C305 source.n81 a_n4174_n2088# 0.03319f
C306 source.n82 a_n4174_n2088# 0.014868f
C307 source.n83 a_n4174_n2088# 0.111825f
C308 source.t46 a_n4174_n2088# 0.054096f
C309 source.n84 a_n4174_n2088# 0.024893f
C310 source.n85 a_n4174_n2088# 0.019605f
C311 source.n86 a_n4174_n2088# 0.014042f
C312 source.n87 a_n4174_n2088# 0.621778f
C313 source.n88 a_n4174_n2088# 0.026132f
C314 source.n89 a_n4174_n2088# 0.014042f
C315 source.n90 a_n4174_n2088# 0.014868f
C316 source.n91 a_n4174_n2088# 0.03319f
C317 source.n92 a_n4174_n2088# 0.03319f
C318 source.n93 a_n4174_n2088# 0.014868f
C319 source.n94 a_n4174_n2088# 0.014042f
C320 source.n95 a_n4174_n2088# 0.026132f
C321 source.n96 a_n4174_n2088# 0.026132f
C322 source.n97 a_n4174_n2088# 0.014042f
C323 source.n98 a_n4174_n2088# 0.014868f
C324 source.n99 a_n4174_n2088# 0.03319f
C325 source.n100 a_n4174_n2088# 0.071851f
C326 source.n101 a_n4174_n2088# 0.014868f
C327 source.n102 a_n4174_n2088# 0.014042f
C328 source.n103 a_n4174_n2088# 0.060402f
C329 source.n104 a_n4174_n2088# 0.040204f
C330 source.n105 a_n4174_n2088# 0.158421f
C331 source.t4 a_n4174_n2088# 0.1239f
C332 source.t11 a_n4174_n2088# 0.1239f
C333 source.n106 a_n4174_n2088# 0.964945f
C334 source.n107 a_n4174_n2088# 0.438043f
C335 source.t20 a_n4174_n2088# 0.1239f
C336 source.t9 a_n4174_n2088# 0.1239f
C337 source.n108 a_n4174_n2088# 0.964945f
C338 source.n109 a_n4174_n2088# 0.438043f
C339 source.t14 a_n4174_n2088# 0.1239f
C340 source.t7 a_n4174_n2088# 0.1239f
C341 source.n110 a_n4174_n2088# 0.964945f
C342 source.n111 a_n4174_n2088# 0.438043f
C343 source.t18 a_n4174_n2088# 0.1239f
C344 source.t16 a_n4174_n2088# 0.1239f
C345 source.n112 a_n4174_n2088# 0.964945f
C346 source.n113 a_n4174_n2088# 0.438043f
C347 source.t10 a_n4174_n2088# 0.1239f
C348 source.t12 a_n4174_n2088# 0.1239f
C349 source.n114 a_n4174_n2088# 0.964945f
C350 source.n115 a_n4174_n2088# 0.438043f
C351 source.n116 a_n4174_n2088# 0.03673f
C352 source.n117 a_n4174_n2088# 0.026132f
C353 source.n118 a_n4174_n2088# 0.014042f
C354 source.n119 a_n4174_n2088# 0.03319f
C355 source.n120 a_n4174_n2088# 0.014868f
C356 source.n121 a_n4174_n2088# 0.026132f
C357 source.n122 a_n4174_n2088# 0.014042f
C358 source.n123 a_n4174_n2088# 0.03319f
C359 source.n124 a_n4174_n2088# 0.014868f
C360 source.n125 a_n4174_n2088# 0.111825f
C361 source.t15 a_n4174_n2088# 0.054096f
C362 source.n126 a_n4174_n2088# 0.024893f
C363 source.n127 a_n4174_n2088# 0.019605f
C364 source.n128 a_n4174_n2088# 0.014042f
C365 source.n129 a_n4174_n2088# 0.621778f
C366 source.n130 a_n4174_n2088# 0.026132f
C367 source.n131 a_n4174_n2088# 0.014042f
C368 source.n132 a_n4174_n2088# 0.014868f
C369 source.n133 a_n4174_n2088# 0.03319f
C370 source.n134 a_n4174_n2088# 0.03319f
C371 source.n135 a_n4174_n2088# 0.014868f
C372 source.n136 a_n4174_n2088# 0.014042f
C373 source.n137 a_n4174_n2088# 0.026132f
C374 source.n138 a_n4174_n2088# 0.026132f
C375 source.n139 a_n4174_n2088# 0.014042f
C376 source.n140 a_n4174_n2088# 0.014868f
C377 source.n141 a_n4174_n2088# 0.03319f
C378 source.n142 a_n4174_n2088# 0.071851f
C379 source.n143 a_n4174_n2088# 0.014868f
C380 source.n144 a_n4174_n2088# 0.014042f
C381 source.n145 a_n4174_n2088# 0.060402f
C382 source.n146 a_n4174_n2088# 0.040204f
C383 source.n147 a_n4174_n2088# 1.071f
C384 source.n148 a_n4174_n2088# 0.03673f
C385 source.n149 a_n4174_n2088# 0.026132f
C386 source.n150 a_n4174_n2088# 0.014042f
C387 source.n151 a_n4174_n2088# 0.03319f
C388 source.n152 a_n4174_n2088# 0.014868f
C389 source.n153 a_n4174_n2088# 0.026132f
C390 source.n154 a_n4174_n2088# 0.014042f
C391 source.n155 a_n4174_n2088# 0.03319f
C392 source.n156 a_n4174_n2088# 0.014868f
C393 source.n157 a_n4174_n2088# 0.111825f
C394 source.t39 a_n4174_n2088# 0.054096f
C395 source.n158 a_n4174_n2088# 0.024893f
C396 source.n159 a_n4174_n2088# 0.019605f
C397 source.n160 a_n4174_n2088# 0.014042f
C398 source.n161 a_n4174_n2088# 0.621778f
C399 source.n162 a_n4174_n2088# 0.026132f
C400 source.n163 a_n4174_n2088# 0.014042f
C401 source.n164 a_n4174_n2088# 0.014868f
C402 source.n165 a_n4174_n2088# 0.03319f
C403 source.n166 a_n4174_n2088# 0.03319f
C404 source.n167 a_n4174_n2088# 0.014868f
C405 source.n168 a_n4174_n2088# 0.014042f
C406 source.n169 a_n4174_n2088# 0.026132f
C407 source.n170 a_n4174_n2088# 0.026132f
C408 source.n171 a_n4174_n2088# 0.014042f
C409 source.n172 a_n4174_n2088# 0.014868f
C410 source.n173 a_n4174_n2088# 0.03319f
C411 source.n174 a_n4174_n2088# 0.071851f
C412 source.n175 a_n4174_n2088# 0.014868f
C413 source.n176 a_n4174_n2088# 0.014042f
C414 source.n177 a_n4174_n2088# 0.060402f
C415 source.n178 a_n4174_n2088# 0.040204f
C416 source.n179 a_n4174_n2088# 1.071f
C417 source.t24 a_n4174_n2088# 0.1239f
C418 source.t44 a_n4174_n2088# 0.1239f
C419 source.n180 a_n4174_n2088# 0.964938f
C420 source.n181 a_n4174_n2088# 0.43805f
C421 source.t40 a_n4174_n2088# 0.1239f
C422 source.t23 a_n4174_n2088# 0.1239f
C423 source.n182 a_n4174_n2088# 0.964938f
C424 source.n183 a_n4174_n2088# 0.43805f
C425 source.t32 a_n4174_n2088# 0.1239f
C426 source.t27 a_n4174_n2088# 0.1239f
C427 source.n184 a_n4174_n2088# 0.964938f
C428 source.n185 a_n4174_n2088# 0.43805f
C429 source.t42 a_n4174_n2088# 0.1239f
C430 source.t29 a_n4174_n2088# 0.1239f
C431 source.n186 a_n4174_n2088# 0.964938f
C432 source.n187 a_n4174_n2088# 0.43805f
C433 source.t25 a_n4174_n2088# 0.1239f
C434 source.t28 a_n4174_n2088# 0.1239f
C435 source.n188 a_n4174_n2088# 0.964938f
C436 source.n189 a_n4174_n2088# 0.43805f
C437 source.n190 a_n4174_n2088# 0.03673f
C438 source.n191 a_n4174_n2088# 0.026132f
C439 source.n192 a_n4174_n2088# 0.014042f
C440 source.n193 a_n4174_n2088# 0.03319f
C441 source.n194 a_n4174_n2088# 0.014868f
C442 source.n195 a_n4174_n2088# 0.026132f
C443 source.n196 a_n4174_n2088# 0.014042f
C444 source.n197 a_n4174_n2088# 0.03319f
C445 source.n198 a_n4174_n2088# 0.014868f
C446 source.n199 a_n4174_n2088# 0.111825f
C447 source.t26 a_n4174_n2088# 0.054096f
C448 source.n200 a_n4174_n2088# 0.024893f
C449 source.n201 a_n4174_n2088# 0.019605f
C450 source.n202 a_n4174_n2088# 0.014042f
C451 source.n203 a_n4174_n2088# 0.621778f
C452 source.n204 a_n4174_n2088# 0.026132f
C453 source.n205 a_n4174_n2088# 0.014042f
C454 source.n206 a_n4174_n2088# 0.014868f
C455 source.n207 a_n4174_n2088# 0.03319f
C456 source.n208 a_n4174_n2088# 0.03319f
C457 source.n209 a_n4174_n2088# 0.014868f
C458 source.n210 a_n4174_n2088# 0.014042f
C459 source.n211 a_n4174_n2088# 0.026132f
C460 source.n212 a_n4174_n2088# 0.026132f
C461 source.n213 a_n4174_n2088# 0.014042f
C462 source.n214 a_n4174_n2088# 0.014868f
C463 source.n215 a_n4174_n2088# 0.03319f
C464 source.n216 a_n4174_n2088# 0.071851f
C465 source.n217 a_n4174_n2088# 0.014868f
C466 source.n218 a_n4174_n2088# 0.014042f
C467 source.n219 a_n4174_n2088# 0.060402f
C468 source.n220 a_n4174_n2088# 0.040204f
C469 source.n221 a_n4174_n2088# 0.158421f
C470 source.n222 a_n4174_n2088# 0.03673f
C471 source.n223 a_n4174_n2088# 0.026132f
C472 source.n224 a_n4174_n2088# 0.014042f
C473 source.n225 a_n4174_n2088# 0.03319f
C474 source.n226 a_n4174_n2088# 0.014868f
C475 source.n227 a_n4174_n2088# 0.026132f
C476 source.n228 a_n4174_n2088# 0.014042f
C477 source.n229 a_n4174_n2088# 0.03319f
C478 source.n230 a_n4174_n2088# 0.014868f
C479 source.n231 a_n4174_n2088# 0.111825f
C480 source.t6 a_n4174_n2088# 0.054096f
C481 source.n232 a_n4174_n2088# 0.024893f
C482 source.n233 a_n4174_n2088# 0.019605f
C483 source.n234 a_n4174_n2088# 0.014042f
C484 source.n235 a_n4174_n2088# 0.621778f
C485 source.n236 a_n4174_n2088# 0.026132f
C486 source.n237 a_n4174_n2088# 0.014042f
C487 source.n238 a_n4174_n2088# 0.014868f
C488 source.n239 a_n4174_n2088# 0.03319f
C489 source.n240 a_n4174_n2088# 0.03319f
C490 source.n241 a_n4174_n2088# 0.014868f
C491 source.n242 a_n4174_n2088# 0.014042f
C492 source.n243 a_n4174_n2088# 0.026132f
C493 source.n244 a_n4174_n2088# 0.026132f
C494 source.n245 a_n4174_n2088# 0.014042f
C495 source.n246 a_n4174_n2088# 0.014868f
C496 source.n247 a_n4174_n2088# 0.03319f
C497 source.n248 a_n4174_n2088# 0.071851f
C498 source.n249 a_n4174_n2088# 0.014868f
C499 source.n250 a_n4174_n2088# 0.014042f
C500 source.n251 a_n4174_n2088# 0.060402f
C501 source.n252 a_n4174_n2088# 0.040204f
C502 source.n253 a_n4174_n2088# 0.158421f
C503 source.t17 a_n4174_n2088# 0.1239f
C504 source.t2 a_n4174_n2088# 0.1239f
C505 source.n254 a_n4174_n2088# 0.964938f
C506 source.n255 a_n4174_n2088# 0.43805f
C507 source.t3 a_n4174_n2088# 0.1239f
C508 source.t0 a_n4174_n2088# 0.1239f
C509 source.n256 a_n4174_n2088# 0.964938f
C510 source.n257 a_n4174_n2088# 0.43805f
C511 source.t5 a_n4174_n2088# 0.1239f
C512 source.t47 a_n4174_n2088# 0.1239f
C513 source.n258 a_n4174_n2088# 0.964938f
C514 source.n259 a_n4174_n2088# 0.43805f
C515 source.t19 a_n4174_n2088# 0.1239f
C516 source.t13 a_n4174_n2088# 0.1239f
C517 source.n260 a_n4174_n2088# 0.964938f
C518 source.n261 a_n4174_n2088# 0.43805f
C519 source.t21 a_n4174_n2088# 0.1239f
C520 source.t1 a_n4174_n2088# 0.1239f
C521 source.n262 a_n4174_n2088# 0.964938f
C522 source.n263 a_n4174_n2088# 0.43805f
C523 source.n264 a_n4174_n2088# 0.03673f
C524 source.n265 a_n4174_n2088# 0.026132f
C525 source.n266 a_n4174_n2088# 0.014042f
C526 source.n267 a_n4174_n2088# 0.03319f
C527 source.n268 a_n4174_n2088# 0.014868f
C528 source.n269 a_n4174_n2088# 0.026132f
C529 source.n270 a_n4174_n2088# 0.014042f
C530 source.n271 a_n4174_n2088# 0.03319f
C531 source.n272 a_n4174_n2088# 0.014868f
C532 source.n273 a_n4174_n2088# 0.111825f
C533 source.t8 a_n4174_n2088# 0.054096f
C534 source.n274 a_n4174_n2088# 0.024893f
C535 source.n275 a_n4174_n2088# 0.019605f
C536 source.n276 a_n4174_n2088# 0.014042f
C537 source.n277 a_n4174_n2088# 0.621778f
C538 source.n278 a_n4174_n2088# 0.026132f
C539 source.n279 a_n4174_n2088# 0.014042f
C540 source.n280 a_n4174_n2088# 0.014868f
C541 source.n281 a_n4174_n2088# 0.03319f
C542 source.n282 a_n4174_n2088# 0.03319f
C543 source.n283 a_n4174_n2088# 0.014868f
C544 source.n284 a_n4174_n2088# 0.014042f
C545 source.n285 a_n4174_n2088# 0.026132f
C546 source.n286 a_n4174_n2088# 0.026132f
C547 source.n287 a_n4174_n2088# 0.014042f
C548 source.n288 a_n4174_n2088# 0.014868f
C549 source.n289 a_n4174_n2088# 0.03319f
C550 source.n290 a_n4174_n2088# 0.071851f
C551 source.n291 a_n4174_n2088# 0.014868f
C552 source.n292 a_n4174_n2088# 0.014042f
C553 source.n293 a_n4174_n2088# 0.060402f
C554 source.n294 a_n4174_n2088# 0.040204f
C555 source.n295 a_n4174_n2088# 0.34576f
C556 source.n296 a_n4174_n2088# 1.09502f
C557 drain_left.t5 a_n4174_n2088# 0.13502f
C558 drain_left.t2 a_n4174_n2088# 0.13502f
C559 drain_left.n0 a_n4174_n2088# 1.13367f
C560 drain_left.t15 a_n4174_n2088# 0.13502f
C561 drain_left.t21 a_n4174_n2088# 0.13502f
C562 drain_left.n1 a_n4174_n2088# 1.12607f
C563 drain_left.n2 a_n4174_n2088# 0.886954f
C564 drain_left.t0 a_n4174_n2088# 0.13502f
C565 drain_left.t4 a_n4174_n2088# 0.13502f
C566 drain_left.n3 a_n4174_n2088# 1.12607f
C567 drain_left.n4 a_n4174_n2088# 0.385135f
C568 drain_left.t20 a_n4174_n2088# 0.13502f
C569 drain_left.t17 a_n4174_n2088# 0.13502f
C570 drain_left.n5 a_n4174_n2088# 1.13367f
C571 drain_left.t22 a_n4174_n2088# 0.13502f
C572 drain_left.t7 a_n4174_n2088# 0.13502f
C573 drain_left.n6 a_n4174_n2088# 1.12607f
C574 drain_left.n7 a_n4174_n2088# 0.886954f
C575 drain_left.t16 a_n4174_n2088# 0.13502f
C576 drain_left.t13 a_n4174_n2088# 0.13502f
C577 drain_left.n8 a_n4174_n2088# 1.12607f
C578 drain_left.n9 a_n4174_n2088# 0.385135f
C579 drain_left.n10 a_n4174_n2088# 1.74739f
C580 drain_left.t3 a_n4174_n2088# 0.13502f
C581 drain_left.t6 a_n4174_n2088# 0.13502f
C582 drain_left.n11 a_n4174_n2088# 1.13367f
C583 drain_left.t12 a_n4174_n2088# 0.13502f
C584 drain_left.t10 a_n4174_n2088# 0.13502f
C585 drain_left.n12 a_n4174_n2088# 1.12607f
C586 drain_left.n13 a_n4174_n2088# 0.886943f
C587 drain_left.t9 a_n4174_n2088# 0.13502f
C588 drain_left.t14 a_n4174_n2088# 0.13502f
C589 drain_left.n14 a_n4174_n2088# 1.12607f
C590 drain_left.n15 a_n4174_n2088# 0.441537f
C591 drain_left.t18 a_n4174_n2088# 0.13502f
C592 drain_left.t11 a_n4174_n2088# 0.13502f
C593 drain_left.n16 a_n4174_n2088# 1.12607f
C594 drain_left.n17 a_n4174_n2088# 0.441537f
C595 drain_left.t8 a_n4174_n2088# 0.13502f
C596 drain_left.t19 a_n4174_n2088# 0.13502f
C597 drain_left.n18 a_n4174_n2088# 1.12607f
C598 drain_left.n19 a_n4174_n2088# 0.441537f
C599 drain_left.t1 a_n4174_n2088# 0.13502f
C600 drain_left.t23 a_n4174_n2088# 0.13502f
C601 drain_left.n20 a_n4174_n2088# 1.12607f
C602 drain_left.n21 a_n4174_n2088# 0.703571f
C603 plus.n0 a_n4174_n2088# 0.047323f
C604 plus.t8 a_n4174_n2088# 0.617198f
C605 plus.t10 a_n4174_n2088# 0.563197f
C606 plus.n1 a_n4174_n2088# 0.231242f
C607 plus.n2 a_n4174_n2088# 0.035464f
C608 plus.t14 a_n4174_n2088# 0.563197f
C609 plus.n3 a_n4174_n2088# 0.028689f
C610 plus.n4 a_n4174_n2088# 0.035464f
C611 plus.t9 a_n4174_n2088# 0.563197f
C612 plus.n5 a_n4174_n2088# 0.034238f
C613 plus.n6 a_n4174_n2088# 0.035464f
C614 plus.t15 a_n4174_n2088# 0.563197f
C615 plus.n7 a_n4174_n2088# 0.028643f
C616 plus.n8 a_n4174_n2088# 0.035464f
C617 plus.t7 a_n4174_n2088# 0.563197f
C618 plus.t12 a_n4174_n2088# 0.563197f
C619 plus.n9 a_n4174_n2088# 0.231242f
C620 plus.n10 a_n4174_n2088# 0.035464f
C621 plus.t4 a_n4174_n2088# 0.563197f
C622 plus.n11 a_n4174_n2088# 0.231242f
C623 plus.n12 a_n4174_n2088# 0.035464f
C624 plus.t0 a_n4174_n2088# 0.563197f
C625 plus.n13 a_n4174_n2088# 0.231242f
C626 plus.n14 a_n4174_n2088# 0.178537f
C627 plus.t2 a_n4174_n2088# 0.563197f
C628 plus.t23 a_n4174_n2088# 0.648356f
C629 plus.n15 a_n4174_n2088# 0.273579f
C630 plus.n16 a_n4174_n2088# 0.284492f
C631 plus.n17 a_n4174_n2088# 0.043711f
C632 plus.n18 a_n4174_n2088# 0.048357f
C633 plus.n19 a_n4174_n2088# 0.035464f
C634 plus.n20 a_n4174_n2088# 0.035464f
C635 plus.n21 a_n4174_n2088# 0.048041f
C636 plus.n22 a_n4174_n2088# 0.028689f
C637 plus.n23 a_n4174_n2088# 0.048637f
C638 plus.n24 a_n4174_n2088# 0.035464f
C639 plus.n25 a_n4174_n2088# 0.035464f
C640 plus.n26 a_n4174_n2088# 0.048933f
C641 plus.n27 a_n4174_n2088# 0.042195f
C642 plus.n28 a_n4174_n2088# 0.034238f
C643 plus.n29 a_n4174_n2088# 0.035464f
C644 plus.n30 a_n4174_n2088# 0.035464f
C645 plus.n31 a_n4174_n2088# 0.043379f
C646 plus.n32 a_n4174_n2088# 0.048689f
C647 plus.n33 a_n4174_n2088# 0.231242f
C648 plus.n34 a_n4174_n2088# 0.048361f
C649 plus.n35 a_n4174_n2088# 0.035464f
C650 plus.n36 a_n4174_n2088# 0.035464f
C651 plus.n37 a_n4174_n2088# 0.035464f
C652 plus.n38 a_n4174_n2088# 0.048361f
C653 plus.n39 a_n4174_n2088# 0.231242f
C654 plus.n40 a_n4174_n2088# 0.048689f
C655 plus.t11 a_n4174_n2088# 0.563197f
C656 plus.n41 a_n4174_n2088# 0.231242f
C657 plus.n42 a_n4174_n2088# 0.043379f
C658 plus.n43 a_n4174_n2088# 0.035464f
C659 plus.n44 a_n4174_n2088# 0.035464f
C660 plus.n45 a_n4174_n2088# 0.035464f
C661 plus.n46 a_n4174_n2088# 0.042195f
C662 plus.n47 a_n4174_n2088# 0.048933f
C663 plus.n48 a_n4174_n2088# 0.231242f
C664 plus.n49 a_n4174_n2088# 0.048637f
C665 plus.n50 a_n4174_n2088# 0.035464f
C666 plus.n51 a_n4174_n2088# 0.035464f
C667 plus.n52 a_n4174_n2088# 0.035464f
C668 plus.n53 a_n4174_n2088# 0.048041f
C669 plus.n54 a_n4174_n2088# 0.231242f
C670 plus.n55 a_n4174_n2088# 0.048357f
C671 plus.n56 a_n4174_n2088# 0.043711f
C672 plus.n57 a_n4174_n2088# 0.035464f
C673 plus.n58 a_n4174_n2088# 0.035464f
C674 plus.n59 a_n4174_n2088# 0.035975f
C675 plus.n60 a_n4174_n2088# 0.037192f
C676 plus.n61 a_n4174_n2088# 0.283193f
C677 plus.n62 a_n4174_n2088# 0.343206f
C678 plus.n63 a_n4174_n2088# 0.047323f
C679 plus.t6 a_n4174_n2088# 0.617198f
C680 plus.t21 a_n4174_n2088# 0.563197f
C681 plus.n64 a_n4174_n2088# 0.231242f
C682 plus.n65 a_n4174_n2088# 0.035464f
C683 plus.t1 a_n4174_n2088# 0.563197f
C684 plus.n66 a_n4174_n2088# 0.028689f
C685 plus.n67 a_n4174_n2088# 0.035464f
C686 plus.t5 a_n4174_n2088# 0.563197f
C687 plus.n68 a_n4174_n2088# 0.034238f
C688 plus.n69 a_n4174_n2088# 0.035464f
C689 plus.t22 a_n4174_n2088# 0.563197f
C690 plus.n70 a_n4174_n2088# 0.231242f
C691 plus.t13 a_n4174_n2088# 0.563197f
C692 plus.n71 a_n4174_n2088# 0.028643f
C693 plus.n72 a_n4174_n2088# 0.035464f
C694 plus.t18 a_n4174_n2088# 0.563197f
C695 plus.t3 a_n4174_n2088# 0.563197f
C696 plus.n73 a_n4174_n2088# 0.231242f
C697 plus.n74 a_n4174_n2088# 0.035464f
C698 plus.t16 a_n4174_n2088# 0.563197f
C699 plus.n75 a_n4174_n2088# 0.231242f
C700 plus.n76 a_n4174_n2088# 0.035464f
C701 plus.t20 a_n4174_n2088# 0.563197f
C702 plus.n77 a_n4174_n2088# 0.231242f
C703 plus.n78 a_n4174_n2088# 0.178537f
C704 plus.t17 a_n4174_n2088# 0.563197f
C705 plus.t19 a_n4174_n2088# 0.648356f
C706 plus.n79 a_n4174_n2088# 0.273579f
C707 plus.n80 a_n4174_n2088# 0.284492f
C708 plus.n81 a_n4174_n2088# 0.043711f
C709 plus.n82 a_n4174_n2088# 0.048357f
C710 plus.n83 a_n4174_n2088# 0.035464f
C711 plus.n84 a_n4174_n2088# 0.035464f
C712 plus.n85 a_n4174_n2088# 0.048041f
C713 plus.n86 a_n4174_n2088# 0.028689f
C714 plus.n87 a_n4174_n2088# 0.048637f
C715 plus.n88 a_n4174_n2088# 0.035464f
C716 plus.n89 a_n4174_n2088# 0.035464f
C717 plus.n90 a_n4174_n2088# 0.048933f
C718 plus.n91 a_n4174_n2088# 0.042195f
C719 plus.n92 a_n4174_n2088# 0.034238f
C720 plus.n93 a_n4174_n2088# 0.035464f
C721 plus.n94 a_n4174_n2088# 0.035464f
C722 plus.n95 a_n4174_n2088# 0.043379f
C723 plus.n96 a_n4174_n2088# 0.048689f
C724 plus.n97 a_n4174_n2088# 0.231242f
C725 plus.n98 a_n4174_n2088# 0.048361f
C726 plus.n99 a_n4174_n2088# 0.035464f
C727 plus.n100 a_n4174_n2088# 0.035464f
C728 plus.n101 a_n4174_n2088# 0.035464f
C729 plus.n102 a_n4174_n2088# 0.048361f
C730 plus.n103 a_n4174_n2088# 0.231242f
C731 plus.n104 a_n4174_n2088# 0.048689f
C732 plus.n105 a_n4174_n2088# 0.043379f
C733 plus.n106 a_n4174_n2088# 0.035464f
C734 plus.n107 a_n4174_n2088# 0.035464f
C735 plus.n108 a_n4174_n2088# 0.035464f
C736 plus.n109 a_n4174_n2088# 0.042195f
C737 plus.n110 a_n4174_n2088# 0.048933f
C738 plus.n111 a_n4174_n2088# 0.231242f
C739 plus.n112 a_n4174_n2088# 0.048637f
C740 plus.n113 a_n4174_n2088# 0.035464f
C741 plus.n114 a_n4174_n2088# 0.035464f
C742 plus.n115 a_n4174_n2088# 0.035464f
C743 plus.n116 a_n4174_n2088# 0.048041f
C744 plus.n117 a_n4174_n2088# 0.231242f
C745 plus.n118 a_n4174_n2088# 0.048357f
C746 plus.n119 a_n4174_n2088# 0.043711f
C747 plus.n120 a_n4174_n2088# 0.035464f
C748 plus.n121 a_n4174_n2088# 0.035464f
C749 plus.n122 a_n4174_n2088# 0.035975f
C750 plus.n123 a_n4174_n2088# 0.037192f
C751 plus.n124 a_n4174_n2088# 0.283193f
C752 plus.n125 a_n4174_n2088# 1.38836f
.ends

