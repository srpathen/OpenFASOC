* NGSPICE file created from opamp19.ext - technology: sky130A

.subckt opamp19 gnd CSoutput output vdd plus minus commonsourceibias outputibias diffpairibias
X0 CSoutput.t178 a_n8964_8799.t36 vdd.t298 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X1 CSoutput.t41 commonsourceibias.t48 gnd.t130 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X2 a_n2472_13878.t27 a_n2650_13878.t56 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 a_n2472_13878.t19 a_n2650_13878.t26 a_n2650_13878.t27 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X4 vdd.t297 a_n8964_8799.t37 CSoutput.t177 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 output.t17 CSoutput.t192 vdd.t58 gnd.t306 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X6 gnd.t129 commonsourceibias.t49 CSoutput.t51 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X7 a_n8964_8799.t6 plus.t5 a_n2903_n3924.t19 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X8 CSoutput.t50 commonsourceibias.t50 gnd.t128 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X9 CSoutput.t10 commonsourceibias.t51 gnd.t127 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 CSoutput.t176 a_n8964_8799.t38 vdd.t296 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 CSoutput.t175 a_n8964_8799.t39 vdd.t295 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X12 minus.t4 gnd.t288 gnd.t290 gnd.t289 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X13 vdd.t294 a_n8964_8799.t40 CSoutput.t174 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X14 a_n2650_8322.t27 a_n2650_13878.t57 a_n8964_8799.t27 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X15 CSoutput.t173 a_n8964_8799.t41 vdd.t293 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 vdd.t292 a_n8964_8799.t42 CSoutput.t172 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X17 CSoutput.t171 a_n8964_8799.t43 vdd.t290 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X18 gnd.t126 commonsourceibias.t52 CSoutput.t182 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X19 CSoutput.t18 commonsourceibias.t53 gnd.t125 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X20 gnd.t124 commonsourceibias.t54 CSoutput.t6 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X21 vdd.t291 a_n8964_8799.t44 CSoutput.t170 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 vdd.t289 a_n8964_8799.t45 CSoutput.t169 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X23 CSoutput.t21 commonsourceibias.t55 gnd.t123 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X24 CSoutput.t184 commonsourceibias.t56 gnd.t122 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 a_n2650_13878.t49 minus.t5 a_n2903_n3924.t31 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 CSoutput.t0 commonsourceibias.t57 gnd.t121 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X27 a_n8964_8799.t2 plus.t6 a_n2903_n3924.t18 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 a_n8964_8799.t24 a_n2650_13878.t58 a_n2650_8322.t26 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X29 a_n2650_13878.t52 minus.t6 a_n2903_n3924.t34 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X30 vdd.t288 a_n8964_8799.t46 CSoutput.t168 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 vdd.t287 a_n8964_8799.t47 CSoutput.t167 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X32 gnd.t287 gnd.t284 gnd.t286 gnd.t285 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X33 a_n8964_8799.t25 a_n2650_13878.t59 a_n2650_8322.t25 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X34 CSoutput.t36 commonsourceibias.t58 gnd.t120 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 gnd.t119 commonsourceibias.t59 CSoutput.t183 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 gnd.t283 gnd.t281 gnd.t282 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X37 CSoutput.t29 commonsourceibias.t60 gnd.t118 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 vdd.t59 CSoutput.t193 output.t16 gnd.t305 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X39 CSoutput.t194 a_n2650_8322.t33 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X40 CSoutput.t15 commonsourceibias.t61 gnd.t117 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X41 CSoutput.t166 a_n8964_8799.t48 vdd.t282 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X42 a_n2903_n3924.t17 plus.t7 a_n8964_8799.t21 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X43 a_n2903_n3924.t21 diffpairibias.t16 gnd.t137 gnd.t136 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X44 a_n2903_n3924.t2 minus.t7 a_n2650_13878.t2 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X45 CSoutput.t165 a_n8964_8799.t49 vdd.t286 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X46 gnd.t116 commonsourceibias.t62 CSoutput.t42 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X47 vdd.t285 a_n8964_8799.t50 CSoutput.t164 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X48 CSoutput.t31 commonsourceibias.t63 gnd.t115 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X49 outputibias.t7 outputibias.t6 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X50 gnd.t114 commonsourceibias.t8 commonsourceibias.t9 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 CSoutput.t11 commonsourceibias.t64 gnd.t113 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 CSoutput.t163 a_n8964_8799.t51 vdd.t284 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 vdd.t283 a_n8964_8799.t52 CSoutput.t162 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 vdd.t138 vdd.t136 vdd.t137 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X55 CSoutput.t23 commonsourceibias.t65 gnd.t112 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 a_n2472_13878.t18 a_n2650_13878.t28 a_n2650_13878.t29 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X57 a_n2650_13878.t19 a_n2650_13878.t18 a_n2472_13878.t17 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 gnd.t111 commonsourceibias.t66 CSoutput.t8 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X59 gnd.t280 gnd.t278 plus.t4 gnd.t279 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X60 CSoutput.t161 a_n8964_8799.t53 vdd.t281 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 gnd.t99 commonsourceibias.t10 commonsourceibias.t11 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X62 vdd.t135 vdd.t133 vdd.t134 vdd.t110 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X63 CSoutput.t48 commonsourceibias.t67 gnd.t110 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X64 a_n2903_n3924.t16 plus.t8 a_n8964_8799.t23 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X65 vdd.t280 a_n8964_8799.t54 CSoutput.t160 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 vdd.t279 a_n8964_8799.t55 CSoutput.t159 vdd.t278 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 gnd.t277 gnd.t275 gnd.t276 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X68 gnd.t274 gnd.t272 gnd.t273 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X69 CSoutput.t7 commonsourceibias.t68 gnd.t109 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 diffpairibias.t15 diffpairibias.t14 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X71 a_n2650_13878.t13 a_n2650_13878.t12 a_n2472_13878.t16 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X72 CSoutput.t181 commonsourceibias.t69 gnd.t108 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X73 CSoutput.t158 a_n8964_8799.t56 vdd.t277 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 CSoutput.t2 commonsourceibias.t70 gnd.t107 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X75 gnd.t106 commonsourceibias.t71 CSoutput.t22 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 vdd.t276 a_n8964_8799.t57 CSoutput.t157 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 a_n8964_8799.t17 a_n2650_13878.t60 a_n2650_8322.t24 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X78 CSoutput.t156 a_n8964_8799.t58 vdd.t275 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X79 gnd.t105 commonsourceibias.t72 CSoutput.t191 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 a_n2650_13878.t7 a_n2650_13878.t6 a_n2472_13878.t15 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X81 vdd.t274 a_n8964_8799.t59 CSoutput.t155 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 vdd.t273 a_n8964_8799.t60 CSoutput.t154 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 a_n8964_8799.t18 a_n2650_13878.t61 a_n2650_8322.t23 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X84 CSoutput.t12 commonsourceibias.t73 gnd.t104 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X85 diffpairibias.t13 diffpairibias.t12 gnd.t9 gnd.t8 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X86 CSoutput.t153 a_n8964_8799.t61 vdd.t272 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 gnd.t103 commonsourceibias.t12 commonsourceibias.t13 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 CSoutput.t19 commonsourceibias.t74 gnd.t102 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 gnd.t101 commonsourceibias.t75 CSoutput.t190 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 CSoutput.t13 commonsourceibias.t76 gnd.t100 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 a_n2650_8322.t22 a_n2650_13878.t62 a_n8964_8799.t10 vdd.t17 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X92 gnd.t98 commonsourceibias.t77 CSoutput.t1 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 CSoutput.t152 a_n8964_8799.t62 vdd.t271 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X94 a_n2903_n3924.t0 minus.t8 a_n2650_13878.t0 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X95 a_n2903_n3924.t15 plus.t9 a_n8964_8799.t34 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X96 gnd.t97 commonsourceibias.t78 CSoutput.t16 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X97 vdd.t132 vdd.t130 vdd.t131 vdd.t106 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X98 a_n2903_n3924.t30 diffpairibias.t17 gnd.t161 gnd.t160 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X99 vdd.t270 a_n8964_8799.t63 CSoutput.t151 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X100 gnd.t271 gnd.t269 gnd.t270 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X101 vdd.t27 CSoutput.t195 output.t15 gnd.t304 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X102 vdd.t269 a_n8964_8799.t64 CSoutput.t150 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 a_n2650_13878.t11 a_n2650_13878.t10 a_n2472_13878.t14 vdd.t42 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X104 vdd.t268 a_n8964_8799.t65 CSoutput.t149 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X105 a_n2903_n3924.t14 plus.t10 a_n8964_8799.t1 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X106 vdd.t267 a_n8964_8799.t66 CSoutput.t148 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 gnd.t96 commonsourceibias.t79 CSoutput.t54 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 a_n8964_8799.t11 a_n2650_13878.t63 a_n2650_8322.t21 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X109 a_n2650_13878.t15 a_n2650_13878.t14 a_n2472_13878.t13 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X110 gnd.t268 gnd.t266 gnd.t267 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X111 CSoutput.t196 a_n2650_8322.t32 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X112 vdd.t28 CSoutput.t197 output.t14 gnd.t303 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X113 vdd.t266 a_n8964_8799.t67 CSoutput.t147 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X114 CSoutput.t146 a_n8964_8799.t68 vdd.t265 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 CSoutput.t145 a_n8964_8799.t69 vdd.t264 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 gnd.t95 commonsourceibias.t80 CSoutput.t57 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X117 vdd.t129 vdd.t127 vdd.t128 vdd.t114 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t94 commonsourceibias.t4 commonsourceibias.t5 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X119 gnd.t93 commonsourceibias.t81 CSoutput.t58 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 CSoutput.t144 a_n8964_8799.t70 vdd.t263 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 vdd.t126 vdd.t123 vdd.t125 vdd.t124 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X122 CSoutput.t143 a_n8964_8799.t71 vdd.t262 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X123 vdd.t261 a_n8964_8799.t72 CSoutput.t142 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 vdd.t38 a_n2650_13878.t64 a_n2650_8322.t7 vdd.t37 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 a_n2650_13878.t43 a_n2650_13878.t42 a_n2472_13878.t12 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X126 gnd.t265 gnd.t263 minus.t3 gnd.t264 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X127 vdd.t122 vdd.t120 vdd.t121 vdd.t90 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X128 a_n2650_8322.t6 a_n2650_13878.t65 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 a_n2903_n3924.t24 diffpairibias.t18 gnd.t147 gnd.t146 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X130 CSoutput.t141 a_n8964_8799.t73 vdd.t260 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X131 CSoutput.t55 commonsourceibias.t82 gnd.t92 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X132 CSoutput.t56 commonsourceibias.t83 gnd.t91 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 gnd.t262 gnd.t260 gnd.t261 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X134 gnd.t259 gnd.t257 gnd.t258 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X135 vdd.t34 a_n2650_13878.t66 a_n2472_13878.t26 vdd.t33 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 vdd.t119 vdd.t117 vdd.t118 vdd.t106 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X137 vdd.t116 vdd.t113 vdd.t115 vdd.t114 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X138 gnd.t256 gnd.t254 gnd.t255 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X139 vdd.t259 a_n8964_8799.t74 CSoutput.t140 vdd.t258 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X140 vdd.t257 a_n8964_8799.t75 CSoutput.t139 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 output.t13 CSoutput.t198 vdd.t60 gnd.t302 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X142 a_n8964_8799.t16 plus.t11 a_n2903_n3924.t13 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X143 vdd.t112 vdd.t109 vdd.t111 vdd.t110 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 a_n2650_8322.t5 a_n2650_13878.t67 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X145 a_n8964_8799.t3 a_n2650_13878.t68 a_n2650_8322.t20 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X146 a_n8964_8799.t19 plus.t12 a_n2903_n3924.t12 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X147 CSoutput.t138 a_n8964_8799.t76 vdd.t256 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 diffpairibias.t11 diffpairibias.t10 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X149 vdd.t255 a_n8964_8799.t77 CSoutput.t137 vdd.t254 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 a_n2650_13878.t39 a_n2650_13878.t38 a_n2472_13878.t11 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 vdd.t253 a_n8964_8799.t78 CSoutput.t136 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 CSoutput.t32 commonsourceibias.t84 gnd.t90 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n8964_8799.t4 a_n2650_13878.t69 a_n2650_8322.t19 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X154 CSoutput.t135 a_n8964_8799.t79 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X155 CSoutput.t134 a_n8964_8799.t80 vdd.t252 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 CSoutput.t133 a_n8964_8799.t81 vdd.t251 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 commonsourceibias.t25 commonsourceibias.t24 gnd.t79 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X158 gnd.t89 commonsourceibias.t85 CSoutput.t33 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X159 a_n2472_13878.t10 a_n2650_13878.t36 a_n2650_13878.t37 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 gnd.t253 gnd.t251 gnd.t252 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X161 vdd.t108 vdd.t105 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X162 vdd.t104 vdd.t102 vdd.t103 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X163 output.t1 outputibias.t8 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X164 CSoutput.t132 a_n8964_8799.t82 vdd.t250 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X165 CSoutput.t34 commonsourceibias.t86 gnd.t88 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 vdd.t15 a_n2650_13878.t70 a_n2650_8322.t4 vdd.t14 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X167 a_n2472_13878.t9 a_n2650_13878.t20 a_n2650_13878.t21 vdd.t43 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 vdd.t249 a_n8964_8799.t83 CSoutput.t131 vdd.t234 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X169 vdd.t248 a_n8964_8799.t84 CSoutput.t130 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X170 a_n2650_13878.t54 minus.t9 a_n2903_n3924.t38 gnd.t10 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X171 a_n2903_n3924.t11 plus.t13 a_n8964_8799.t22 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X172 vdd.t101 vdd.t99 vdd.t100 vdd.t90 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X173 gnd.t87 commonsourceibias.t87 CSoutput.t35 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X174 gnd.t86 commonsourceibias.t88 CSoutput.t37 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 a_n2650_13878.t23 a_n2650_13878.t22 a_n2472_13878.t8 vdd.t299 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X176 CSoutput.t199 a_n2650_8322.t31 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X177 commonsourceibias.t45 commonsourceibias.t44 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 vdd.t61 CSoutput.t200 output.t12 gnd.t301 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X179 output.t11 CSoutput.t201 vdd.t62 gnd.t300 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X180 output.t19 outputibias.t9 gnd.t319 gnd.t318 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X181 gnd.t83 commonsourceibias.t89 CSoutput.t38 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X182 plus.t3 gnd.t248 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X183 vdd.t247 a_n8964_8799.t85 CSoutput.t129 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X184 CSoutput.t39 commonsourceibias.t90 gnd.t82 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X185 a_n2903_n3924.t37 diffpairibias.t19 gnd.t314 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X186 gnd.t247 gnd.t245 minus.t2 gnd.t246 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X187 gnd.t244 gnd.t241 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X188 a_n2903_n3924.t25 diffpairibias.t20 gnd.t149 gnd.t148 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X189 output.t10 CSoutput.t202 vdd.t54 gnd.t299 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X190 commonsourceibias.t27 commonsourceibias.t26 gnd.t81 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 a_n8964_8799.t15 plus.t14 a_n2903_n3924.t10 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 vdd.t246 a_n8964_8799.t86 CSoutput.t128 vdd.t234 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X193 vdd.t245 a_n8964_8799.t87 CSoutput.t127 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 CSoutput.t126 a_n8964_8799.t88 vdd.t244 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X195 gnd.t240 gnd.t238 gnd.t239 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X196 CSoutput.t40 commonsourceibias.t91 gnd.t78 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 a_n8964_8799.t30 plus.t15 a_n2903_n3924.t9 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X198 CSoutput.t43 commonsourceibias.t92 gnd.t77 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X199 a_n2472_13878.t7 a_n2650_13878.t30 a_n2650_13878.t31 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X200 gnd.t237 gnd.t235 gnd.t236 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X201 vdd.t98 vdd.t96 vdd.t97 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X202 a_n2650_8322.t18 a_n2650_13878.t71 a_n8964_8799.t9 vdd.t16 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X203 CSoutput.t125 a_n8964_8799.t89 vdd.t243 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X204 CSoutput.t124 a_n8964_8799.t90 vdd.t242 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 CSoutput.t123 a_n8964_8799.t91 vdd.t239 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X206 commonsourceibias.t39 commonsourceibias.t38 gnd.t72 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 diffpairibias.t9 diffpairibias.t8 gnd.t170 gnd.t169 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 a_n2472_13878.t25 a_n2650_13878.t72 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 a_n2650_13878.t51 minus.t10 a_n2903_n3924.t33 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X210 vdd.t32 a_n2650_13878.t73 a_n2472_13878.t24 vdd.t31 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X211 CSoutput.t44 commonsourceibias.t93 gnd.t76 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t52 commonsourceibias.t94 gnd.t75 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 CSoutput.t122 a_n8964_8799.t92 vdd.t237 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 output.t9 CSoutput.t203 vdd.t55 gnd.t298 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X215 gnd.t74 commonsourceibias.t22 commonsourceibias.t23 gnd.t73 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 vdd.t56 CSoutput.t204 output.t8 gnd.t297 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X217 a_n2903_n3924.t8 plus.t16 a_n8964_8799.t12 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X218 vdd.t235 a_n8964_8799.t93 CSoutput.t121 vdd.t234 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X219 vdd.t233 a_n8964_8799.t94 CSoutput.t120 vdd.t232 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X220 vdd.t231 a_n8964_8799.t95 CSoutput.t119 vdd.t230 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X221 commonsourceibias.t37 commonsourceibias.t36 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 CSoutput.t118 a_n8964_8799.t96 vdd.t229 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X223 a_n2472_13878.t6 a_n2650_13878.t4 a_n2650_13878.t5 vdd.t41 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X224 gnd.t69 commonsourceibias.t95 CSoutput.t53 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X225 commonsourceibias.t35 commonsourceibias.t34 gnd.t68 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X226 vdd.t228 a_n8964_8799.t97 CSoutput.t117 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X227 vdd.t57 CSoutput.t205 output.t7 gnd.t296 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X228 outputibias.t5 outputibias.t4 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X229 gnd.t67 commonsourceibias.t32 commonsourceibias.t33 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 a_n2903_n3924.t26 minus.t11 a_n2650_13878.t46 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X231 a_n2650_8322.t17 a_n2650_13878.t74 a_n8964_8799.t5 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 CSoutput.t116 a_n8964_8799.t98 vdd.t227 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 diffpairibias.t7 diffpairibias.t6 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X234 gnd.t234 gnd.t232 gnd.t233 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X235 vdd.t226 a_n8964_8799.t99 CSoutput.t115 vdd.t225 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X236 a_n2472_13878.t5 a_n2650_13878.t34 a_n2650_13878.t35 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X237 commonsourceibias.t31 commonsourceibias.t30 gnd.t66 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X238 CSoutput.t206 a_n2650_8322.t30 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X239 vdd.t11 a_n2650_13878.t75 a_n2650_8322.t3 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X240 vdd.t224 a_n8964_8799.t100 CSoutput.t114 vdd.t223 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 plus.t2 gnd.t229 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X242 gnd.t228 gnd.t226 minus.t1 gnd.t227 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X243 gnd.t65 commonsourceibias.t96 CSoutput.t9 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X244 CSoutput.t113 a_n8964_8799.t101 vdd.t222 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 gnd.t64 commonsourceibias.t28 commonsourceibias.t29 gnd.t63 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 a_n2472_13878.t23 a_n2650_13878.t76 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X247 vdd.t95 vdd.t93 vdd.t94 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X248 CSoutput.t207 a_n2650_8322.t29 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X249 vdd.t221 a_n8964_8799.t102 CSoutput.t112 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 vdd.t219 a_n8964_8799.t103 CSoutput.t111 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X251 CSoutput.t110 a_n8964_8799.t104 vdd.t218 vdd.t217 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 CSoutput.t109 a_n8964_8799.t105 vdd.t216 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X253 vdd.t300 CSoutput.t208 output.t6 gnd.t295 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X254 gnd.t225 gnd.t222 gnd.t224 gnd.t223 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X255 vdd.t215 a_n8964_8799.t106 CSoutput.t108 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 a_n2903_n3924.t27 diffpairibias.t21 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X257 vdd.t23 a_n2650_13878.t77 a_n2650_8322.t2 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X258 a_n2650_8322.t16 a_n2650_13878.t78 a_n8964_8799.t7 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X259 gnd.t62 commonsourceibias.t2 commonsourceibias.t3 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 a_n8964_8799.t35 plus.t17 a_n2903_n3924.t7 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X261 a_n2650_13878.t53 minus.t12 a_n2903_n3924.t35 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X262 CSoutput.t107 a_n8964_8799.t107 vdd.t214 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 vdd.t92 vdd.t89 vdd.t91 vdd.t90 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X264 vdd.t213 a_n8964_8799.t108 CSoutput.t106 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 a_n2903_n3924.t39 minus.t13 a_n2650_13878.t55 gnd.t317 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X266 vdd.t88 vdd.t86 vdd.t87 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X267 vdd.t212 a_n8964_8799.t109 CSoutput.t105 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X268 vdd.t211 a_n8964_8799.t110 CSoutput.t104 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X269 output.t5 CSoutput.t209 vdd.t301 gnd.t294 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X270 gnd.t55 commonsourceibias.t0 commonsourceibias.t1 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 vdd.t85 vdd.t82 vdd.t84 vdd.t83 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X272 a_n2903_n3924.t28 minus.t14 a_n2650_13878.t47 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X273 vdd.t210 a_n8964_8799.t111 CSoutput.t103 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 CSoutput.t102 a_n8964_8799.t112 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 CSoutput.t45 commonsourceibias.t97 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X276 a_n2903_n3924.t29 minus.t15 a_n2650_13878.t48 gnd.t155 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X277 a_n2472_13878.t4 a_n2650_13878.t32 a_n2650_13878.t33 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X278 CSoutput.t101 a_n8964_8799.t113 vdd.t207 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 CSoutput.t100 a_n8964_8799.t114 vdd.t206 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X280 a_n2650_8322.t15 a_n2650_13878.t79 a_n8964_8799.t8 vdd.t13 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X281 vdd.t81 vdd.t79 vdd.t80 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X282 diffpairibias.t5 diffpairibias.t4 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X283 gnd.t221 gnd.t218 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X284 CSoutput.t99 a_n8964_8799.t115 vdd.t205 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t98 a_n8964_8799.t116 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 CSoutput.t97 a_n8964_8799.t117 vdd.t201 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 vdd.t200 a_n8964_8799.t118 CSoutput.t96 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X288 vdd.t78 vdd.t75 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X289 gnd.t217 gnd.t214 gnd.t216 gnd.t215 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X290 CSoutput.t27 commonsourceibias.t98 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X291 output.t4 CSoutput.t210 vdd.t51 gnd.t293 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X292 vdd.t199 a_n8964_8799.t119 CSoutput.t95 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X293 vdd.t52 CSoutput.t211 output.t3 gnd.t292 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X294 a_n2650_8322.t1 a_n2650_13878.t80 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X295 CSoutput.t94 a_n8964_8799.t120 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 output.t0 outputibias.t10 gnd.t142 gnd.t141 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X297 a_n2903_n3924.t1 minus.t16 a_n2650_13878.t1 gnd.t3 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X298 vdd.t195 a_n8964_8799.t121 CSoutput.t93 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X299 gnd.t213 gnd.t211 gnd.t212 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X300 gnd.t57 commonsourceibias.t99 CSoutput.t49 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 CSoutput.t92 a_n8964_8799.t122 vdd.t194 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X302 outputibias.t3 outputibias.t2 gnd.t151 gnd.t150 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X303 vdd.t6 a_n2650_13878.t81 a_n2472_13878.t22 vdd.t5 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X304 vdd.t193 a_n8964_8799.t123 CSoutput.t91 vdd.t192 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 CSoutput.t90 a_n8964_8799.t124 vdd.t191 vdd.t190 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 CSoutput.t89 a_n8964_8799.t125 vdd.t189 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X307 vdd.t188 a_n8964_8799.t126 CSoutput.t88 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X308 vdd.t186 a_n8964_8799.t127 CSoutput.t87 vdd.t185 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 vdd.t184 a_n8964_8799.t128 CSoutput.t86 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 gnd.t210 gnd.t207 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X311 gnd.t56 commonsourceibias.t100 CSoutput.t24 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 gnd.t206 gnd.t204 plus.t1 gnd.t205 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X313 gnd.t54 commonsourceibias.t101 CSoutput.t25 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 gnd.t203 gnd.t201 gnd.t202 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X315 a_n2650_8322.t14 a_n2650_13878.t82 a_n8964_8799.t13 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X316 commonsourceibias.t15 commonsourceibias.t14 gnd.t53 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 a_n8964_8799.t14 a_n2650_13878.t83 a_n2650_8322.t13 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X318 a_n2472_13878.t21 a_n2650_13878.t84 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X319 gnd.t51 commonsourceibias.t102 CSoutput.t28 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t74 vdd.t71 vdd.t73 vdd.t72 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X321 vdd.t183 a_n8964_8799.t129 CSoutput.t85 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 vdd.t70 vdd.t67 vdd.t69 vdd.t68 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X323 CSoutput.t84 a_n8964_8799.t130 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X324 CSoutput.t83 a_n8964_8799.t131 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput.t82 a_n8964_8799.t132 vdd.t142 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X326 vdd.t66 vdd.t63 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X327 a_n2903_n3924.t6 plus.t18 a_n8964_8799.t20 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X328 a_n2650_13878.t3 minus.t17 a_n2903_n3924.t3 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X329 a_n8964_8799.t0 a_n2650_13878.t85 a_n2650_8322.t12 vdd.t2 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X330 gnd.t50 commonsourceibias.t103 CSoutput.t26 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X331 commonsourceibias.t41 commonsourceibias.t40 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 a_n2650_8322.t11 a_n2650_13878.t86 a_n8964_8799.t31 vdd.t45 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X333 gnd.t47 commonsourceibias.t104 CSoutput.t179 gnd.t46 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X334 vdd.t178 a_n8964_8799.t133 CSoutput.t81 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 gnd.t45 commonsourceibias.t16 commonsourceibias.t17 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 output.t2 CSoutput.t212 vdd.t53 gnd.t291 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X337 CSoutput.t80 a_n8964_8799.t134 vdd.t176 vdd.t175 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 CSoutput.t79 a_n8964_8799.t135 vdd.t174 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 CSoutput.t78 a_n8964_8799.t136 vdd.t173 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X340 a_n2472_13878.t3 a_n2650_13878.t8 a_n2650_13878.t9 vdd.t7 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X341 vdd.t172 a_n8964_8799.t137 CSoutput.t77 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X342 gnd.t43 commonsourceibias.t6 commonsourceibias.t7 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X343 commonsourceibias.t43 commonsourceibias.t42 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 outputibias.t1 outputibias.t0 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X345 a_n2903_n3924.t23 minus.t18 a_n2650_13878.t45 gnd.t145 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X346 gnd.t40 commonsourceibias.t105 CSoutput.t180 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 a_n2903_n3924.t36 diffpairibias.t22 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X348 CSoutput.t17 commonsourceibias.t106 gnd.t38 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 vdd.t171 a_n8964_8799.t138 CSoutput.t76 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X350 gnd.t37 commonsourceibias.t107 CSoutput.t20 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 CSoutput.t75 a_n8964_8799.t139 vdd.t170 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 a_n2650_13878.t25 a_n2650_13878.t24 a_n2472_13878.t2 vdd.t26 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X353 gnd.t200 gnd.t197 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X354 a_n8964_8799.t32 a_n2650_13878.t87 a_n2650_8322.t10 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X355 gnd.t196 gnd.t193 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X356 vdd.t144 a_n8964_8799.t140 CSoutput.t74 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 CSoutput.t73 a_n8964_8799.t141 vdd.t169 vdd.t168 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X358 CSoutput.t3 commonsourceibias.t108 gnd.t35 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 gnd.t34 commonsourceibias.t109 CSoutput.t185 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X360 commonsourceibias.t19 commonsourceibias.t18 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X361 diffpairibias.t3 diffpairibias.t2 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X362 gnd.t192 gnd.t189 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X363 vdd.t167 a_n8964_8799.t142 CSoutput.t72 vdd.t166 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 CSoutput.t71 a_n8964_8799.t143 vdd.t165 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 output.t18 outputibias.t11 gnd.t316 gnd.t315 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X366 gnd.t188 gnd.t186 plus.t0 gnd.t187 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X367 minus.t0 gnd.t183 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X368 CSoutput.t70 a_n8964_8799.t144 vdd.t164 vdd.t163 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X369 a_n2650_8322.t9 a_n2650_13878.t88 a_n8964_8799.t33 vdd.t299 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X370 gnd.t30 commonsourceibias.t110 CSoutput.t14 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 a_n2650_13878.t44 minus.t19 a_n2903_n3924.t22 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X372 vdd.t162 a_n8964_8799.t145 CSoutput.t69 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 CSoutput.t68 a_n8964_8799.t146 vdd.t145 vdd.t141 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X374 CSoutput.t67 a_n8964_8799.t147 vdd.t160 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X375 diffpairibias.t1 diffpairibias.t0 gnd.t310 gnd.t309 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X376 commonsourceibias.t47 commonsourceibias.t46 gnd.t29 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X377 gnd.t28 commonsourceibias.t111 CSoutput.t4 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X378 gnd.t182 gnd.t179 gnd.t181 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X379 gnd.t178 gnd.t175 gnd.t177 gnd.t176 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X380 CSoutput.t213 a_n2650_8322.t28 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X381 CSoutput.t186 commonsourceibias.t112 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X382 vdd.t303 a_n2650_13878.t89 a_n2472_13878.t20 vdd.t302 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X383 CSoutput.t66 a_n8964_8799.t148 vdd.t158 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X384 vdd.t156 a_n8964_8799.t149 CSoutput.t65 vdd.t155 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X385 vdd.t154 a_n8964_8799.t150 CSoutput.t64 vdd.t143 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X386 gnd.t25 commonsourceibias.t20 commonsourceibias.t21 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X387 CSoutput.t63 a_n8964_8799.t151 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X388 a_n8964_8799.t29 plus.t19 a_n2903_n3924.t5 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X389 a_n2650_13878.t50 minus.t20 a_n2903_n3924.t32 gnd.t138 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X390 gnd.t23 commonsourceibias.t113 CSoutput.t46 gnd.t22 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X391 gnd.t21 commonsourceibias.t114 CSoutput.t30 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X392 a_n2650_8322.t8 a_n2650_13878.t90 a_n8964_8799.t26 vdd.t46 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X393 vdd.t149 a_n8964_8799.t152 CSoutput.t62 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X394 vdd.t151 a_n8964_8799.t153 CSoutput.t61 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X395 CSoutput.t60 a_n8964_8799.t154 vdd.t147 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 gnd.t19 commonsourceibias.t115 CSoutput.t188 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 a_n2650_8322.t0 a_n2650_13878.t91 vdd.t48 vdd.t47 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X398 gnd.t174 gnd.t171 gnd.t173 gnd.t172 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X399 gnd.t18 commonsourceibias.t116 CSoutput.t189 gnd.t17 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 a_n2472_13878.t1 a_n2650_13878.t16 a_n2650_13878.t17 vdd.t44 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X401 gnd.t16 commonsourceibias.t117 CSoutput.t187 gnd.t15 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 CSoutput.t5 commonsourceibias.t118 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X403 CSoutput.t47 commonsourceibias.t119 gnd.t12 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 a_n2903_n3924.t4 plus.t20 a_n8964_8799.t28 gnd.t152 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X405 a_n2903_n3924.t20 diffpairibias.t23 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X406 CSoutput.t59 a_n8964_8799.t155 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X407 a_n2650_13878.t41 a_n2650_13878.t40 a_n2472_13878.t0 vdd.t9 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 a_n8964_8799.n223 a_n8964_8799.t132 485.149
R1 a_n8964_8799.n242 a_n8964_8799.t146 485.149
R2 a_n8964_8799.n262 a_n8964_8799.t88 485.149
R3 a_n8964_8799.n162 a_n8964_8799.t83 485.149
R4 a_n8964_8799.n181 a_n8964_8799.t93 485.149
R5 a_n8964_8799.n201 a_n8964_8799.t86 485.149
R6 a_n8964_8799.n55 a_n8964_8799.t103 485.135
R7 a_n8964_8799.n235 a_n8964_8799.t39 464.166
R8 a_n8964_8799.n217 a_n8964_8799.t109 464.166
R9 a_n8964_8799.n234 a_n8964_8799.t107 464.166
R10 a_n8964_8799.n233 a_n8964_8799.t45 464.166
R11 a_n8964_8799.n218 a_n8964_8799.t43 464.166
R12 a_n8964_8799.n232 a_n8964_8799.t129 464.166
R13 a_n8964_8799.n231 a_n8964_8799.t61 464.166
R14 a_n8964_8799.n219 a_n8964_8799.t47 464.166
R15 a_n8964_8799.n230 a_n8964_8799.t135 464.166
R16 a_n8964_8799.n229 a_n8964_8799.t87 464.166
R17 a_n8964_8799.n220 a_n8964_8799.t62 464.166
R18 a_n8964_8799.n228 a_n8964_8799.t153 464.166
R19 a_n8964_8799.n227 a_n8964_8799.t105 464.166
R20 a_n8964_8799.n221 a_n8964_8799.t64 464.166
R21 a_n8964_8799.n226 a_n8964_8799.t147 464.166
R22 a_n8964_8799.n225 a_n8964_8799.t108 464.166
R23 a_n8964_8799.n222 a_n8964_8799.t81 464.166
R24 a_n8964_8799.n224 a_n8964_8799.t44 464.166
R25 a_n8964_8799.n70 a_n8964_8799.t119 485.135
R26 a_n8964_8799.n254 a_n8964_8799.t51 464.166
R27 a_n8964_8799.n236 a_n8964_8799.t127 464.166
R28 a_n8964_8799.n253 a_n8964_8799.t125 464.166
R29 a_n8964_8799.n252 a_n8964_8799.t54 464.166
R30 a_n8964_8799.n237 a_n8964_8799.t53 464.166
R31 a_n8964_8799.n251 a_n8964_8799.t145 464.166
R32 a_n8964_8799.n250 a_n8964_8799.t70 464.166
R33 a_n8964_8799.n238 a_n8964_8799.t60 464.166
R34 a_n8964_8799.n249 a_n8964_8799.t148 464.166
R35 a_n8964_8799.n248 a_n8964_8799.t100 464.166
R36 a_n8964_8799.n239 a_n8964_8799.t73 464.166
R37 a_n8964_8799.n247 a_n8964_8799.t46 464.166
R38 a_n8964_8799.n246 a_n8964_8799.t120 464.166
R39 a_n8964_8799.n240 a_n8964_8799.t74 464.166
R40 a_n8964_8799.n245 a_n8964_8799.t38 464.166
R41 a_n8964_8799.n244 a_n8964_8799.t126 464.166
R42 a_n8964_8799.n241 a_n8964_8799.t89 464.166
R43 a_n8964_8799.n243 a_n8964_8799.t55 464.166
R44 a_n8964_8799.n85 a_n8964_8799.t65 485.135
R45 a_n8964_8799.n274 a_n8964_8799.t151 464.166
R46 a_n8964_8799.n256 a_n8964_8799.t118 464.166
R47 a_n8964_8799.n273 a_n8964_8799.t144 464.166
R48 a_n8964_8799.n272 a_n8964_8799.t99 464.166
R49 a_n8964_8799.n257 a_n8964_8799.t124 464.166
R50 a_n8964_8799.n271 a_n8964_8799.t59 464.166
R51 a_n8964_8799.n270 a_n8964_8799.t141 464.166
R52 a_n8964_8799.n258 a_n8964_8799.t77 464.166
R53 a_n8964_8799.n269 a_n8964_8799.t136 464.166
R54 a_n8964_8799.n268 a_n8964_8799.t63 464.166
R55 a_n8964_8799.n259 a_n8964_8799.t112 464.166
R56 a_n8964_8799.n267 a_n8964_8799.t50 464.166
R57 a_n8964_8799.n266 a_n8964_8799.t96 464.166
R58 a_n8964_8799.n260 a_n8964_8799.t72 464.166
R59 a_n8964_8799.n265 a_n8964_8799.t122 464.166
R60 a_n8964_8799.n264 a_n8964_8799.t57 464.166
R61 a_n8964_8799.n261 a_n8964_8799.t104 464.166
R62 a_n8964_8799.n263 a_n8964_8799.t42 464.166
R63 a_n8964_8799.n163 a_n8964_8799.t113 464.166
R64 a_n8964_8799.n164 a_n8964_8799.t40 464.166
R65 a_n8964_8799.n165 a_n8964_8799.t68 464.166
R66 a_n8964_8799.n166 a_n8964_8799.t106 464.166
R67 a_n8964_8799.n161 a_n8964_8799.t143 464.166
R68 a_n8964_8799.n167 a_n8964_8799.t66 464.166
R69 a_n8964_8799.n168 a_n8964_8799.t101 464.166
R70 a_n8964_8799.n169 a_n8964_8799.t138 464.166
R71 a_n8964_8799.n170 a_n8964_8799.t139 464.166
R72 a_n8964_8799.n160 a_n8964_8799.t85 464.166
R73 a_n8964_8799.n171 a_n8964_8799.t117 464.166
R74 a_n8964_8799.n159 a_n8964_8799.t137 464.166
R75 a_n8964_8799.n172 a_n8964_8799.t82 464.166
R76 a_n8964_8799.n173 a_n8964_8799.t84 464.166
R77 a_n8964_8799.n174 a_n8964_8799.t114 464.166
R78 a_n8964_8799.n175 a_n8964_8799.t67 464.166
R79 a_n8964_8799.n158 a_n8964_8799.t69 464.166
R80 a_n8964_8799.n176 a_n8964_8799.t110 464.166
R81 a_n8964_8799.n182 a_n8964_8799.t130 464.166
R82 a_n8964_8799.n183 a_n8964_8799.t52 464.166
R83 a_n8964_8799.n184 a_n8964_8799.t79 464.166
R84 a_n8964_8799.n185 a_n8964_8799.t121 464.166
R85 a_n8964_8799.n180 a_n8964_8799.t155 464.166
R86 a_n8964_8799.n186 a_n8964_8799.t75 464.166
R87 a_n8964_8799.n187 a_n8964_8799.t115 464.166
R88 a_n8964_8799.n188 a_n8964_8799.t152 464.166
R89 a_n8964_8799.n189 a_n8964_8799.t154 464.166
R90 a_n8964_8799.n179 a_n8964_8799.t97 464.166
R91 a_n8964_8799.n190 a_n8964_8799.t134 464.166
R92 a_n8964_8799.n178 a_n8964_8799.t150 464.166
R93 a_n8964_8799.n191 a_n8964_8799.t92 464.166
R94 a_n8964_8799.n192 a_n8964_8799.t94 464.166
R95 a_n8964_8799.n193 a_n8964_8799.t131 464.166
R96 a_n8964_8799.n194 a_n8964_8799.t78 464.166
R97 a_n8964_8799.n177 a_n8964_8799.t80 464.166
R98 a_n8964_8799.n195 a_n8964_8799.t128 464.166
R99 a_n8964_8799.n202 a_n8964_8799.t41 464.166
R100 a_n8964_8799.n203 a_n8964_8799.t102 464.166
R101 a_n8964_8799.n204 a_n8964_8799.t56 464.166
R102 a_n8964_8799.n205 a_n8964_8799.t123 464.166
R103 a_n8964_8799.n200 a_n8964_8799.t71 464.166
R104 a_n8964_8799.n206 a_n8964_8799.t95 464.166
R105 a_n8964_8799.n207 a_n8964_8799.t49 464.166
R106 a_n8964_8799.n208 a_n8964_8799.t111 464.166
R107 a_n8964_8799.n209 a_n8964_8799.t90 464.166
R108 a_n8964_8799.n199 a_n8964_8799.t133 464.166
R109 a_n8964_8799.n210 a_n8964_8799.t76 464.166
R110 a_n8964_8799.n198 a_n8964_8799.t140 464.166
R111 a_n8964_8799.n211 a_n8964_8799.t58 464.166
R112 a_n8964_8799.n212 a_n8964_8799.t37 464.166
R113 a_n8964_8799.n213 a_n8964_8799.t98 464.166
R114 a_n8964_8799.n214 a_n8964_8799.t142 464.166
R115 a_n8964_8799.n197 a_n8964_8799.t116 464.166
R116 a_n8964_8799.n215 a_n8964_8799.t149 464.166
R117 a_n8964_8799.n44 a_n8964_8799.n69 71.7212
R118 a_n8964_8799.n69 a_n8964_8799.n222 17.8606
R119 a_n8964_8799.n68 a_n8964_8799.n44 76.9909
R120 a_n8964_8799.n225 a_n8964_8799.n68 7.32118
R121 a_n8964_8799.n67 a_n8964_8799.n43 78.3454
R122 a_n8964_8799.n43 a_n8964_8799.n66 72.8951
R123 a_n8964_8799.n65 a_n8964_8799.n45 70.1674
R124 a_n8964_8799.n228 a_n8964_8799.n65 20.9683
R125 a_n8964_8799.n45 a_n8964_8799.n64 72.3034
R126 a_n8964_8799.n64 a_n8964_8799.n220 16.6962
R127 a_n8964_8799.n63 a_n8964_8799.n46 77.6622
R128 a_n8964_8799.n229 a_n8964_8799.n63 5.97853
R129 a_n8964_8799.n62 a_n8964_8799.n46 77.6622
R130 a_n8964_8799.n47 a_n8964_8799.n61 72.3034
R131 a_n8964_8799.n60 a_n8964_8799.n47 70.1674
R132 a_n8964_8799.n232 a_n8964_8799.n60 20.9683
R133 a_n8964_8799.n49 a_n8964_8799.n59 72.8951
R134 a_n8964_8799.n59 a_n8964_8799.n218 15.5127
R135 a_n8964_8799.n58 a_n8964_8799.n49 78.3454
R136 a_n8964_8799.n233 a_n8964_8799.n58 4.61226
R137 a_n8964_8799.n57 a_n8964_8799.n48 76.9909
R138 a_n8964_8799.n48 a_n8964_8799.n56 71.7212
R139 a_n8964_8799.n235 a_n8964_8799.n55 20.9683
R140 a_n8964_8799.n50 a_n8964_8799.n55 70.1674
R141 a_n8964_8799.n36 a_n8964_8799.n84 71.7212
R142 a_n8964_8799.n84 a_n8964_8799.n241 17.8606
R143 a_n8964_8799.n83 a_n8964_8799.n36 76.9909
R144 a_n8964_8799.n244 a_n8964_8799.n83 7.32118
R145 a_n8964_8799.n82 a_n8964_8799.n35 78.3454
R146 a_n8964_8799.n35 a_n8964_8799.n81 72.8951
R147 a_n8964_8799.n80 a_n8964_8799.n37 70.1674
R148 a_n8964_8799.n247 a_n8964_8799.n80 20.9683
R149 a_n8964_8799.n37 a_n8964_8799.n79 72.3034
R150 a_n8964_8799.n79 a_n8964_8799.n239 16.6962
R151 a_n8964_8799.n78 a_n8964_8799.n38 77.6622
R152 a_n8964_8799.n248 a_n8964_8799.n78 5.97853
R153 a_n8964_8799.n77 a_n8964_8799.n38 77.6622
R154 a_n8964_8799.n39 a_n8964_8799.n76 72.3034
R155 a_n8964_8799.n75 a_n8964_8799.n39 70.1674
R156 a_n8964_8799.n251 a_n8964_8799.n75 20.9683
R157 a_n8964_8799.n41 a_n8964_8799.n74 72.8951
R158 a_n8964_8799.n74 a_n8964_8799.n237 15.5127
R159 a_n8964_8799.n73 a_n8964_8799.n41 78.3454
R160 a_n8964_8799.n252 a_n8964_8799.n73 4.61226
R161 a_n8964_8799.n72 a_n8964_8799.n40 76.9909
R162 a_n8964_8799.n40 a_n8964_8799.n71 71.7212
R163 a_n8964_8799.n254 a_n8964_8799.n70 20.9683
R164 a_n8964_8799.n42 a_n8964_8799.n70 70.1674
R165 a_n8964_8799.n28 a_n8964_8799.n99 71.7212
R166 a_n8964_8799.n99 a_n8964_8799.n261 17.8606
R167 a_n8964_8799.n98 a_n8964_8799.n28 76.9909
R168 a_n8964_8799.n264 a_n8964_8799.n98 7.32118
R169 a_n8964_8799.n97 a_n8964_8799.n27 78.3454
R170 a_n8964_8799.n27 a_n8964_8799.n96 72.8951
R171 a_n8964_8799.n95 a_n8964_8799.n29 70.1674
R172 a_n8964_8799.n267 a_n8964_8799.n95 20.9683
R173 a_n8964_8799.n29 a_n8964_8799.n94 72.3034
R174 a_n8964_8799.n94 a_n8964_8799.n259 16.6962
R175 a_n8964_8799.n93 a_n8964_8799.n30 77.6622
R176 a_n8964_8799.n268 a_n8964_8799.n93 5.97853
R177 a_n8964_8799.n92 a_n8964_8799.n30 77.6622
R178 a_n8964_8799.n31 a_n8964_8799.n91 72.3034
R179 a_n8964_8799.n90 a_n8964_8799.n31 70.1674
R180 a_n8964_8799.n271 a_n8964_8799.n90 20.9683
R181 a_n8964_8799.n33 a_n8964_8799.n89 72.8951
R182 a_n8964_8799.n89 a_n8964_8799.n257 15.5127
R183 a_n8964_8799.n88 a_n8964_8799.n33 78.3454
R184 a_n8964_8799.n272 a_n8964_8799.n88 4.61226
R185 a_n8964_8799.n87 a_n8964_8799.n32 76.9909
R186 a_n8964_8799.n32 a_n8964_8799.n86 71.7212
R187 a_n8964_8799.n274 a_n8964_8799.n85 20.9683
R188 a_n8964_8799.n34 a_n8964_8799.n85 70.1674
R189 a_n8964_8799.n20 a_n8964_8799.n114 70.1674
R190 a_n8964_8799.n176 a_n8964_8799.n114 20.9683
R191 a_n8964_8799.n113 a_n8964_8799.n20 71.7212
R192 a_n8964_8799.n113 a_n8964_8799.n158 17.8606
R193 a_n8964_8799.n19 a_n8964_8799.n112 76.9909
R194 a_n8964_8799.n175 a_n8964_8799.n112 7.32118
R195 a_n8964_8799.n111 a_n8964_8799.n19 78.3454
R196 a_n8964_8799.n21 a_n8964_8799.n110 72.8951
R197 a_n8964_8799.n109 a_n8964_8799.n21 70.1674
R198 a_n8964_8799.n109 a_n8964_8799.n159 20.9683
R199 a_n8964_8799.n22 a_n8964_8799.n108 72.3034
R200 a_n8964_8799.n171 a_n8964_8799.n108 16.6962
R201 a_n8964_8799.n107 a_n8964_8799.n22 77.6622
R202 a_n8964_8799.n107 a_n8964_8799.n160 5.97853
R203 a_n8964_8799.n23 a_n8964_8799.n106 77.6622
R204 a_n8964_8799.n105 a_n8964_8799.n23 72.3034
R205 a_n8964_8799.n24 a_n8964_8799.n104 70.1674
R206 a_n8964_8799.n167 a_n8964_8799.n104 20.9683
R207 a_n8964_8799.n103 a_n8964_8799.n24 72.8951
R208 a_n8964_8799.n103 a_n8964_8799.n161 15.5127
R209 a_n8964_8799.n25 a_n8964_8799.n102 78.3454
R210 a_n8964_8799.n166 a_n8964_8799.n102 4.61226
R211 a_n8964_8799.n101 a_n8964_8799.n25 76.9909
R212 a_n8964_8799.n100 a_n8964_8799.n164 17.8606
R213 a_n8964_8799.n100 a_n8964_8799.n26 71.7212
R214 a_n8964_8799.n12 a_n8964_8799.n129 70.1674
R215 a_n8964_8799.n195 a_n8964_8799.n129 20.9683
R216 a_n8964_8799.n128 a_n8964_8799.n12 71.7212
R217 a_n8964_8799.n128 a_n8964_8799.n177 17.8606
R218 a_n8964_8799.n11 a_n8964_8799.n127 76.9909
R219 a_n8964_8799.n194 a_n8964_8799.n127 7.32118
R220 a_n8964_8799.n126 a_n8964_8799.n11 78.3454
R221 a_n8964_8799.n13 a_n8964_8799.n125 72.8951
R222 a_n8964_8799.n124 a_n8964_8799.n13 70.1674
R223 a_n8964_8799.n124 a_n8964_8799.n178 20.9683
R224 a_n8964_8799.n14 a_n8964_8799.n123 72.3034
R225 a_n8964_8799.n190 a_n8964_8799.n123 16.6962
R226 a_n8964_8799.n122 a_n8964_8799.n14 77.6622
R227 a_n8964_8799.n122 a_n8964_8799.n179 5.97853
R228 a_n8964_8799.n15 a_n8964_8799.n121 77.6622
R229 a_n8964_8799.n120 a_n8964_8799.n15 72.3034
R230 a_n8964_8799.n16 a_n8964_8799.n119 70.1674
R231 a_n8964_8799.n186 a_n8964_8799.n119 20.9683
R232 a_n8964_8799.n118 a_n8964_8799.n16 72.8951
R233 a_n8964_8799.n118 a_n8964_8799.n180 15.5127
R234 a_n8964_8799.n17 a_n8964_8799.n117 78.3454
R235 a_n8964_8799.n185 a_n8964_8799.n117 4.61226
R236 a_n8964_8799.n116 a_n8964_8799.n17 76.9909
R237 a_n8964_8799.n115 a_n8964_8799.n183 17.8606
R238 a_n8964_8799.n115 a_n8964_8799.n18 71.7212
R239 a_n8964_8799.n4 a_n8964_8799.n144 70.1674
R240 a_n8964_8799.n215 a_n8964_8799.n144 20.9683
R241 a_n8964_8799.n143 a_n8964_8799.n4 71.7212
R242 a_n8964_8799.n143 a_n8964_8799.n197 17.8606
R243 a_n8964_8799.n3 a_n8964_8799.n142 76.9909
R244 a_n8964_8799.n214 a_n8964_8799.n142 7.32118
R245 a_n8964_8799.n141 a_n8964_8799.n3 78.3454
R246 a_n8964_8799.n5 a_n8964_8799.n140 72.8951
R247 a_n8964_8799.n139 a_n8964_8799.n5 70.1674
R248 a_n8964_8799.n139 a_n8964_8799.n198 20.9683
R249 a_n8964_8799.n6 a_n8964_8799.n138 72.3034
R250 a_n8964_8799.n210 a_n8964_8799.n138 16.6962
R251 a_n8964_8799.n137 a_n8964_8799.n6 77.6622
R252 a_n8964_8799.n137 a_n8964_8799.n199 5.97853
R253 a_n8964_8799.n7 a_n8964_8799.n136 77.6622
R254 a_n8964_8799.n135 a_n8964_8799.n7 72.3034
R255 a_n8964_8799.n8 a_n8964_8799.n134 70.1674
R256 a_n8964_8799.n206 a_n8964_8799.n134 20.9683
R257 a_n8964_8799.n133 a_n8964_8799.n8 72.8951
R258 a_n8964_8799.n133 a_n8964_8799.n200 15.5127
R259 a_n8964_8799.n9 a_n8964_8799.n132 78.3454
R260 a_n8964_8799.n205 a_n8964_8799.n132 4.61226
R261 a_n8964_8799.n131 a_n8964_8799.n9 76.9909
R262 a_n8964_8799.n130 a_n8964_8799.n203 17.8606
R263 a_n8964_8799.n130 a_n8964_8799.n10 71.7212
R264 a_n8964_8799.n51 a_n8964_8799.n145 98.9633
R265 a_n8964_8799.n53 a_n8964_8799.n279 98.9631
R266 a_n8964_8799.n53 a_n8964_8799.n280 98.6055
R267 a_n8964_8799.n53 a_n8964_8799.n281 98.6055
R268 a_n8964_8799.n54 a_n8964_8799.n282 98.6055
R269 a_n8964_8799.n52 a_n8964_8799.n149 98.6055
R270 a_n8964_8799.n52 a_n8964_8799.n148 98.6055
R271 a_n8964_8799.n51 a_n8964_8799.n147 98.6055
R272 a_n8964_8799.n51 a_n8964_8799.n146 98.6055
R273 a_n8964_8799.n283 a_n8964_8799.n54 98.6054
R274 a_n8964_8799.n1 a_n8964_8799.n150 81.4626
R275 a_n8964_8799.n2 a_n8964_8799.n154 81.4626
R276 a_n8964_8799.n2 a_n8964_8799.n152 81.4626
R277 a_n8964_8799.n0 a_n8964_8799.n156 80.9324
R278 a_n8964_8799.n1 a_n8964_8799.n157 80.9324
R279 a_n8964_8799.n1 a_n8964_8799.n151 80.9324
R280 a_n8964_8799.n2 a_n8964_8799.n155 80.9324
R281 a_n8964_8799.n2 a_n8964_8799.n153 80.9324
R282 a_n8964_8799.n44 a_n8964_8799.n223 70.4033
R283 a_n8964_8799.n36 a_n8964_8799.n242 70.4033
R284 a_n8964_8799.n28 a_n8964_8799.n262 70.4033
R285 a_n8964_8799.n162 a_n8964_8799.n26 70.4033
R286 a_n8964_8799.n181 a_n8964_8799.n18 70.4033
R287 a_n8964_8799.n201 a_n8964_8799.n10 70.4033
R288 a_n8964_8799.n234 a_n8964_8799.n233 48.2005
R289 a_n8964_8799.n60 a_n8964_8799.n231 20.9683
R290 a_n8964_8799.n230 a_n8964_8799.n229 48.2005
R291 a_n8964_8799.n65 a_n8964_8799.n227 20.9683
R292 a_n8964_8799.n226 a_n8964_8799.n225 48.2005
R293 a_n8964_8799.n253 a_n8964_8799.n252 48.2005
R294 a_n8964_8799.n75 a_n8964_8799.n250 20.9683
R295 a_n8964_8799.n249 a_n8964_8799.n248 48.2005
R296 a_n8964_8799.n80 a_n8964_8799.n246 20.9683
R297 a_n8964_8799.n245 a_n8964_8799.n244 48.2005
R298 a_n8964_8799.n273 a_n8964_8799.n272 48.2005
R299 a_n8964_8799.n90 a_n8964_8799.n270 20.9683
R300 a_n8964_8799.n269 a_n8964_8799.n268 48.2005
R301 a_n8964_8799.n95 a_n8964_8799.n266 20.9683
R302 a_n8964_8799.n265 a_n8964_8799.n264 48.2005
R303 a_n8964_8799.n166 a_n8964_8799.n165 48.2005
R304 a_n8964_8799.n168 a_n8964_8799.n104 20.9683
R305 a_n8964_8799.n170 a_n8964_8799.n160 48.2005
R306 a_n8964_8799.n172 a_n8964_8799.n109 20.9683
R307 a_n8964_8799.n175 a_n8964_8799.n174 48.2005
R308 a_n8964_8799.t36 a_n8964_8799.n114 485.135
R309 a_n8964_8799.n185 a_n8964_8799.n184 48.2005
R310 a_n8964_8799.n187 a_n8964_8799.n119 20.9683
R311 a_n8964_8799.n189 a_n8964_8799.n179 48.2005
R312 a_n8964_8799.n191 a_n8964_8799.n124 20.9683
R313 a_n8964_8799.n194 a_n8964_8799.n193 48.2005
R314 a_n8964_8799.t48 a_n8964_8799.n129 485.135
R315 a_n8964_8799.n205 a_n8964_8799.n204 48.2005
R316 a_n8964_8799.n207 a_n8964_8799.n134 20.9683
R317 a_n8964_8799.n209 a_n8964_8799.n199 48.2005
R318 a_n8964_8799.n211 a_n8964_8799.n139 20.9683
R319 a_n8964_8799.n214 a_n8964_8799.n213 48.2005
R320 a_n8964_8799.t91 a_n8964_8799.n144 485.135
R321 a_n8964_8799.n56 a_n8964_8799.n217 17.8606
R322 a_n8964_8799.n224 a_n8964_8799.n69 25.894
R323 a_n8964_8799.n71 a_n8964_8799.n236 17.8606
R324 a_n8964_8799.n243 a_n8964_8799.n84 25.894
R325 a_n8964_8799.n86 a_n8964_8799.n256 17.8606
R326 a_n8964_8799.n263 a_n8964_8799.n99 25.894
R327 a_n8964_8799.n176 a_n8964_8799.n113 25.894
R328 a_n8964_8799.n195 a_n8964_8799.n128 25.894
R329 a_n8964_8799.n215 a_n8964_8799.n143 25.894
R330 a_n8964_8799.n67 a_n8964_8799.n221 43.3183
R331 a_n8964_8799.n82 a_n8964_8799.n240 43.3183
R332 a_n8964_8799.n97 a_n8964_8799.n260 43.3183
R333 a_n8964_8799.n173 a_n8964_8799.n111 43.3183
R334 a_n8964_8799.n192 a_n8964_8799.n126 43.3183
R335 a_n8964_8799.n212 a_n8964_8799.n141 43.3183
R336 a_n8964_8799.n61 a_n8964_8799.n219 16.6962
R337 a_n8964_8799.n228 a_n8964_8799.n64 27.6507
R338 a_n8964_8799.n76 a_n8964_8799.n238 16.6962
R339 a_n8964_8799.n247 a_n8964_8799.n79 27.6507
R340 a_n8964_8799.n91 a_n8964_8799.n258 16.6962
R341 a_n8964_8799.n267 a_n8964_8799.n94 27.6507
R342 a_n8964_8799.n169 a_n8964_8799.n105 16.6962
R343 a_n8964_8799.n159 a_n8964_8799.n108 27.6507
R344 a_n8964_8799.n188 a_n8964_8799.n120 16.6962
R345 a_n8964_8799.n178 a_n8964_8799.n123 27.6507
R346 a_n8964_8799.n208 a_n8964_8799.n135 16.6962
R347 a_n8964_8799.n198 a_n8964_8799.n138 27.6507
R348 a_n8964_8799.n62 a_n8964_8799.n219 41.7634
R349 a_n8964_8799.n77 a_n8964_8799.n238 41.7634
R350 a_n8964_8799.n92 a_n8964_8799.n258 41.7634
R351 a_n8964_8799.n106 a_n8964_8799.n169 41.7634
R352 a_n8964_8799.n121 a_n8964_8799.n188 41.7634
R353 a_n8964_8799.n136 a_n8964_8799.n208 41.7634
R354 a_n8964_8799.n232 a_n8964_8799.n59 29.3885
R355 a_n8964_8799.n66 a_n8964_8799.n221 15.5127
R356 a_n8964_8799.n251 a_n8964_8799.n74 29.3885
R357 a_n8964_8799.n81 a_n8964_8799.n240 15.5127
R358 a_n8964_8799.n271 a_n8964_8799.n89 29.3885
R359 a_n8964_8799.n96 a_n8964_8799.n260 15.5127
R360 a_n8964_8799.n167 a_n8964_8799.n103 29.3885
R361 a_n8964_8799.n173 a_n8964_8799.n110 15.5127
R362 a_n8964_8799.n186 a_n8964_8799.n118 29.3885
R363 a_n8964_8799.n192 a_n8964_8799.n125 15.5127
R364 a_n8964_8799.n206 a_n8964_8799.n133 29.3885
R365 a_n8964_8799.n212 a_n8964_8799.n140 15.5127
R366 a_n8964_8799.n57 a_n8964_8799.n217 40.1848
R367 a_n8964_8799.n72 a_n8964_8799.n236 40.1848
R368 a_n8964_8799.n87 a_n8964_8799.n256 40.1848
R369 a_n8964_8799.n164 a_n8964_8799.n101 40.1848
R370 a_n8964_8799.n183 a_n8964_8799.n116 40.1848
R371 a_n8964_8799.n203 a_n8964_8799.n131 40.1848
R372 a_n8964_8799.n54 a_n8964_8799.n278 32.8105
R373 a_n8964_8799.n224 a_n8964_8799.n223 20.9576
R374 a_n8964_8799.n243 a_n8964_8799.n242 20.9576
R375 a_n8964_8799.n263 a_n8964_8799.n262 20.9576
R376 a_n8964_8799.n163 a_n8964_8799.n162 20.9576
R377 a_n8964_8799.n182 a_n8964_8799.n181 20.9576
R378 a_n8964_8799.n202 a_n8964_8799.n201 20.9576
R379 a_n8964_8799.n278 a_n8964_8799.n52 19.9322
R380 a_n8964_8799.n57 a_n8964_8799.n234 7.32118
R381 a_n8964_8799.n68 a_n8964_8799.n222 40.1848
R382 a_n8964_8799.n72 a_n8964_8799.n253 7.32118
R383 a_n8964_8799.n83 a_n8964_8799.n241 40.1848
R384 a_n8964_8799.n87 a_n8964_8799.n273 7.32118
R385 a_n8964_8799.n98 a_n8964_8799.n261 40.1848
R386 a_n8964_8799.n165 a_n8964_8799.n101 7.32118
R387 a_n8964_8799.n158 a_n8964_8799.n112 40.1848
R388 a_n8964_8799.n184 a_n8964_8799.n116 7.32118
R389 a_n8964_8799.n177 a_n8964_8799.n127 40.1848
R390 a_n8964_8799.n204 a_n8964_8799.n131 7.32118
R391 a_n8964_8799.n197 a_n8964_8799.n142 40.1848
R392 a_n8964_8799.n227 a_n8964_8799.n66 29.3885
R393 a_n8964_8799.n246 a_n8964_8799.n81 29.3885
R394 a_n8964_8799.n266 a_n8964_8799.n96 29.3885
R395 a_n8964_8799.n110 a_n8964_8799.n172 29.3885
R396 a_n8964_8799.n125 a_n8964_8799.n191 29.3885
R397 a_n8964_8799.n140 a_n8964_8799.n211 29.3885
R398 a_n8964_8799.n62 a_n8964_8799.n230 5.97853
R399 a_n8964_8799.n63 a_n8964_8799.n220 41.7634
R400 a_n8964_8799.n77 a_n8964_8799.n249 5.97853
R401 a_n8964_8799.n78 a_n8964_8799.n239 41.7634
R402 a_n8964_8799.n92 a_n8964_8799.n269 5.97853
R403 a_n8964_8799.n93 a_n8964_8799.n259 41.7634
R404 a_n8964_8799.n170 a_n8964_8799.n106 5.97853
R405 a_n8964_8799.n171 a_n8964_8799.n107 41.7634
R406 a_n8964_8799.n189 a_n8964_8799.n121 5.97853
R407 a_n8964_8799.n190 a_n8964_8799.n122 41.7634
R408 a_n8964_8799.n209 a_n8964_8799.n136 5.97853
R409 a_n8964_8799.n210 a_n8964_8799.n137 41.7634
R410 a_n8964_8799.n277 a_n8964_8799.n1 12.3339
R411 a_n8964_8799.n278 a_n8964_8799.n277 11.4887
R412 a_n8964_8799.n231 a_n8964_8799.n61 27.6507
R413 a_n8964_8799.n250 a_n8964_8799.n76 27.6507
R414 a_n8964_8799.n270 a_n8964_8799.n91 27.6507
R415 a_n8964_8799.n168 a_n8964_8799.n105 27.6507
R416 a_n8964_8799.n187 a_n8964_8799.n120 27.6507
R417 a_n8964_8799.n207 a_n8964_8799.n135 27.6507
R418 a_n8964_8799.n58 a_n8964_8799.n218 43.3183
R419 a_n8964_8799.n67 a_n8964_8799.n226 4.61226
R420 a_n8964_8799.n73 a_n8964_8799.n237 43.3183
R421 a_n8964_8799.n82 a_n8964_8799.n245 4.61226
R422 a_n8964_8799.n88 a_n8964_8799.n257 43.3183
R423 a_n8964_8799.n97 a_n8964_8799.n265 4.61226
R424 a_n8964_8799.n161 a_n8964_8799.n102 43.3183
R425 a_n8964_8799.n174 a_n8964_8799.n111 4.61226
R426 a_n8964_8799.n180 a_n8964_8799.n117 43.3183
R427 a_n8964_8799.n193 a_n8964_8799.n126 4.61226
R428 a_n8964_8799.n200 a_n8964_8799.n132 43.3183
R429 a_n8964_8799.n0 a_n8964_8799.n2 33.2634
R430 a_n8964_8799.n213 a_n8964_8799.n141 4.61226
R431 a_n8964_8799.n255 a_n8964_8799.n50 9.04406
R432 a_n8964_8799.n196 a_n8964_8799.n20 9.04406
R433 a_n8964_8799.n235 a_n8964_8799.n56 25.894
R434 a_n8964_8799.n254 a_n8964_8799.n71 25.894
R435 a_n8964_8799.n274 a_n8964_8799.n86 25.894
R436 a_n8964_8799.n100 a_n8964_8799.n163 25.894
R437 a_n8964_8799.n115 a_n8964_8799.n182 25.894
R438 a_n8964_8799.n130 a_n8964_8799.n202 25.894
R439 a_n8964_8799.n276 a_n8964_8799.n216 7.07069
R440 a_n8964_8799.n276 a_n8964_8799.n275 6.72822
R441 a_n8964_8799.n255 a_n8964_8799.n42 4.93611
R442 a_n8964_8799.n275 a_n8964_8799.n34 4.93611
R443 a_n8964_8799.n196 a_n8964_8799.n12 4.93611
R444 a_n8964_8799.n216 a_n8964_8799.n4 4.93611
R445 a_n8964_8799.n275 a_n8964_8799.n255 4.10845
R446 a_n8964_8799.n216 a_n8964_8799.n196 4.10845
R447 a_n8964_8799.n279 a_n8964_8799.t7 3.61217
R448 a_n8964_8799.n279 a_n8964_8799.t25 3.61217
R449 a_n8964_8799.n280 a_n8964_8799.t27 3.61217
R450 a_n8964_8799.n280 a_n8964_8799.t3 3.61217
R451 a_n8964_8799.n281 a_n8964_8799.t13 3.61217
R452 a_n8964_8799.n281 a_n8964_8799.t14 3.61217
R453 a_n8964_8799.n282 a_n8964_8799.t31 3.61217
R454 a_n8964_8799.n282 a_n8964_8799.t17 3.61217
R455 a_n8964_8799.n149 a_n8964_8799.t9 3.61217
R456 a_n8964_8799.n149 a_n8964_8799.t18 3.61217
R457 a_n8964_8799.n148 a_n8964_8799.t33 3.61217
R458 a_n8964_8799.n148 a_n8964_8799.t24 3.61217
R459 a_n8964_8799.n147 a_n8964_8799.t8 3.61217
R460 a_n8964_8799.n147 a_n8964_8799.t32 3.61217
R461 a_n8964_8799.n146 a_n8964_8799.t5 3.61217
R462 a_n8964_8799.n146 a_n8964_8799.t11 3.61217
R463 a_n8964_8799.n145 a_n8964_8799.t26 3.61217
R464 a_n8964_8799.n145 a_n8964_8799.t4 3.61217
R465 a_n8964_8799.n283 a_n8964_8799.t10 3.61217
R466 a_n8964_8799.t0 a_n8964_8799.n283 3.61217
R467 a_n8964_8799.n277 a_n8964_8799.n276 3.4105
R468 a_n8964_8799.n156 a_n8964_8799.t1 2.82907
R469 a_n8964_8799.n156 a_n8964_8799.t19 2.82907
R470 a_n8964_8799.n157 a_n8964_8799.t22 2.82907
R471 a_n8964_8799.n157 a_n8964_8799.t15 2.82907
R472 a_n8964_8799.n151 a_n8964_8799.t20 2.82907
R473 a_n8964_8799.n151 a_n8964_8799.t35 2.82907
R474 a_n8964_8799.n150 a_n8964_8799.t34 2.82907
R475 a_n8964_8799.n150 a_n8964_8799.t6 2.82907
R476 a_n8964_8799.n154 a_n8964_8799.t23 2.82907
R477 a_n8964_8799.n154 a_n8964_8799.t16 2.82907
R478 a_n8964_8799.n155 a_n8964_8799.t28 2.82907
R479 a_n8964_8799.n155 a_n8964_8799.t29 2.82907
R480 a_n8964_8799.n153 a_n8964_8799.t12 2.82907
R481 a_n8964_8799.n153 a_n8964_8799.t30 2.82907
R482 a_n8964_8799.n152 a_n8964_8799.t21 2.82907
R483 a_n8964_8799.n152 a_n8964_8799.t2 2.82907
R484 a_n8964_8799.n44 a_n8964_8799.n43 1.13686
R485 a_n8964_8799.n36 a_n8964_8799.n35 1.13686
R486 a_n8964_8799.n28 a_n8964_8799.n27 1.13686
R487 a_n8964_8799.n20 a_n8964_8799.n19 1.13686
R488 a_n8964_8799.n12 a_n8964_8799.n11 1.13686
R489 a_n8964_8799.n4 a_n8964_8799.n3 1.13686
R490 a_n8964_8799.n54 a_n8964_8799.n53 1.07378
R491 a_n8964_8799.n52 a_n8964_8799.n51 1.07378
R492 a_n8964_8799.n1 a_n8964_8799.n0 1.06084
R493 a_n8964_8799.n49 a_n8964_8799.n48 0.758076
R494 a_n8964_8799.n49 a_n8964_8799.n47 0.758076
R495 a_n8964_8799.n47 a_n8964_8799.n46 0.758076
R496 a_n8964_8799.n46 a_n8964_8799.n45 0.758076
R497 a_n8964_8799.n43 a_n8964_8799.n45 0.758076
R498 a_n8964_8799.n41 a_n8964_8799.n40 0.758076
R499 a_n8964_8799.n41 a_n8964_8799.n39 0.758076
R500 a_n8964_8799.n39 a_n8964_8799.n38 0.758076
R501 a_n8964_8799.n38 a_n8964_8799.n37 0.758076
R502 a_n8964_8799.n35 a_n8964_8799.n37 0.758076
R503 a_n8964_8799.n33 a_n8964_8799.n32 0.758076
R504 a_n8964_8799.n33 a_n8964_8799.n31 0.758076
R505 a_n8964_8799.n31 a_n8964_8799.n30 0.758076
R506 a_n8964_8799.n30 a_n8964_8799.n29 0.758076
R507 a_n8964_8799.n27 a_n8964_8799.n29 0.758076
R508 a_n8964_8799.n24 a_n8964_8799.n25 0.758076
R509 a_n8964_8799.n23 a_n8964_8799.n24 0.758076
R510 a_n8964_8799.n22 a_n8964_8799.n23 0.758076
R511 a_n8964_8799.n21 a_n8964_8799.n22 0.758076
R512 a_n8964_8799.n19 a_n8964_8799.n21 0.758076
R513 a_n8964_8799.n16 a_n8964_8799.n17 0.758076
R514 a_n8964_8799.n15 a_n8964_8799.n16 0.758076
R515 a_n8964_8799.n14 a_n8964_8799.n15 0.758076
R516 a_n8964_8799.n13 a_n8964_8799.n14 0.758076
R517 a_n8964_8799.n11 a_n8964_8799.n13 0.758076
R518 a_n8964_8799.n8 a_n8964_8799.n9 0.758076
R519 a_n8964_8799.n7 a_n8964_8799.n8 0.758076
R520 a_n8964_8799.n6 a_n8964_8799.n7 0.758076
R521 a_n8964_8799.n5 a_n8964_8799.n6 0.758076
R522 a_n8964_8799.n3 a_n8964_8799.n5 0.758076
R523 a_n8964_8799.n9 a_n8964_8799.n10 0.568682
R524 a_n8964_8799.n17 a_n8964_8799.n18 0.568682
R525 a_n8964_8799.n25 a_n8964_8799.n26 0.568682
R526 a_n8964_8799.n32 a_n8964_8799.n34 0.568682
R527 a_n8964_8799.n40 a_n8964_8799.n42 0.568682
R528 a_n8964_8799.n48 a_n8964_8799.n50 0.568682
R529 vdd.n327 vdd.n291 756.745
R530 vdd.n268 vdd.n232 756.745
R531 vdd.n225 vdd.n189 756.745
R532 vdd.n166 vdd.n130 756.745
R533 vdd.n124 vdd.n88 756.745
R534 vdd.n65 vdd.n29 756.745
R535 vdd.n1826 vdd.n1790 756.745
R536 vdd.n1885 vdd.n1849 756.745
R537 vdd.n1724 vdd.n1688 756.745
R538 vdd.n1783 vdd.n1747 756.745
R539 vdd.n1623 vdd.n1587 756.745
R540 vdd.n1682 vdd.n1646 756.745
R541 vdd.n1136 vdd.t71 640.208
R542 vdd.n997 vdd.t109 640.208
R543 vdd.n1130 vdd.t136 640.208
R544 vdd.n988 vdd.t133 640.208
R545 vdd.n885 vdd.t82 640.208
R546 vdd.n2761 vdd.t127 640.208
R547 vdd.n832 vdd.t96 640.208
R548 vdd.n2830 vdd.t113 640.208
R549 vdd.n799 vdd.t67 640.208
R550 vdd.n1058 vdd.t123 640.208
R551 vdd.n1397 vdd.t105 592.009
R552 vdd.n1435 vdd.t117 592.009
R553 vdd.n1331 vdd.t130 592.009
R554 vdd.n2200 vdd.t89 592.009
R555 vdd.n2050 vdd.t99 592.009
R556 vdd.n2010 vdd.t120 592.009
R557 vdd.n426 vdd.t102 592.009
R558 vdd.n440 vdd.t75 592.009
R559 vdd.n452 vdd.t93 592.009
R560 vdd.n768 vdd.t63 592.009
R561 vdd.n3366 vdd.t79 592.009
R562 vdd.n688 vdd.t86 592.009
R563 vdd.n328 vdd.n327 585
R564 vdd.n326 vdd.n293 585
R565 vdd.n325 vdd.n324 585
R566 vdd.n296 vdd.n294 585
R567 vdd.n319 vdd.n318 585
R568 vdd.n317 vdd.n316 585
R569 vdd.n300 vdd.n299 585
R570 vdd.n311 vdd.n310 585
R571 vdd.n309 vdd.n308 585
R572 vdd.n304 vdd.n303 585
R573 vdd.n269 vdd.n268 585
R574 vdd.n267 vdd.n234 585
R575 vdd.n266 vdd.n265 585
R576 vdd.n237 vdd.n235 585
R577 vdd.n260 vdd.n259 585
R578 vdd.n258 vdd.n257 585
R579 vdd.n241 vdd.n240 585
R580 vdd.n252 vdd.n251 585
R581 vdd.n250 vdd.n249 585
R582 vdd.n245 vdd.n244 585
R583 vdd.n226 vdd.n225 585
R584 vdd.n224 vdd.n191 585
R585 vdd.n223 vdd.n222 585
R586 vdd.n194 vdd.n192 585
R587 vdd.n217 vdd.n216 585
R588 vdd.n215 vdd.n214 585
R589 vdd.n198 vdd.n197 585
R590 vdd.n209 vdd.n208 585
R591 vdd.n207 vdd.n206 585
R592 vdd.n202 vdd.n201 585
R593 vdd.n167 vdd.n166 585
R594 vdd.n165 vdd.n132 585
R595 vdd.n164 vdd.n163 585
R596 vdd.n135 vdd.n133 585
R597 vdd.n158 vdd.n157 585
R598 vdd.n156 vdd.n155 585
R599 vdd.n139 vdd.n138 585
R600 vdd.n150 vdd.n149 585
R601 vdd.n148 vdd.n147 585
R602 vdd.n143 vdd.n142 585
R603 vdd.n125 vdd.n124 585
R604 vdd.n123 vdd.n90 585
R605 vdd.n122 vdd.n121 585
R606 vdd.n93 vdd.n91 585
R607 vdd.n116 vdd.n115 585
R608 vdd.n114 vdd.n113 585
R609 vdd.n97 vdd.n96 585
R610 vdd.n108 vdd.n107 585
R611 vdd.n106 vdd.n105 585
R612 vdd.n101 vdd.n100 585
R613 vdd.n66 vdd.n65 585
R614 vdd.n64 vdd.n31 585
R615 vdd.n63 vdd.n62 585
R616 vdd.n34 vdd.n32 585
R617 vdd.n57 vdd.n56 585
R618 vdd.n55 vdd.n54 585
R619 vdd.n38 vdd.n37 585
R620 vdd.n49 vdd.n48 585
R621 vdd.n47 vdd.n46 585
R622 vdd.n42 vdd.n41 585
R623 vdd.n1827 vdd.n1826 585
R624 vdd.n1825 vdd.n1792 585
R625 vdd.n1824 vdd.n1823 585
R626 vdd.n1795 vdd.n1793 585
R627 vdd.n1818 vdd.n1817 585
R628 vdd.n1816 vdd.n1815 585
R629 vdd.n1799 vdd.n1798 585
R630 vdd.n1810 vdd.n1809 585
R631 vdd.n1808 vdd.n1807 585
R632 vdd.n1803 vdd.n1802 585
R633 vdd.n1886 vdd.n1885 585
R634 vdd.n1884 vdd.n1851 585
R635 vdd.n1883 vdd.n1882 585
R636 vdd.n1854 vdd.n1852 585
R637 vdd.n1877 vdd.n1876 585
R638 vdd.n1875 vdd.n1874 585
R639 vdd.n1858 vdd.n1857 585
R640 vdd.n1869 vdd.n1868 585
R641 vdd.n1867 vdd.n1866 585
R642 vdd.n1862 vdd.n1861 585
R643 vdd.n1725 vdd.n1724 585
R644 vdd.n1723 vdd.n1690 585
R645 vdd.n1722 vdd.n1721 585
R646 vdd.n1693 vdd.n1691 585
R647 vdd.n1716 vdd.n1715 585
R648 vdd.n1714 vdd.n1713 585
R649 vdd.n1697 vdd.n1696 585
R650 vdd.n1708 vdd.n1707 585
R651 vdd.n1706 vdd.n1705 585
R652 vdd.n1701 vdd.n1700 585
R653 vdd.n1784 vdd.n1783 585
R654 vdd.n1782 vdd.n1749 585
R655 vdd.n1781 vdd.n1780 585
R656 vdd.n1752 vdd.n1750 585
R657 vdd.n1775 vdd.n1774 585
R658 vdd.n1773 vdd.n1772 585
R659 vdd.n1756 vdd.n1755 585
R660 vdd.n1767 vdd.n1766 585
R661 vdd.n1765 vdd.n1764 585
R662 vdd.n1760 vdd.n1759 585
R663 vdd.n1624 vdd.n1623 585
R664 vdd.n1622 vdd.n1589 585
R665 vdd.n1621 vdd.n1620 585
R666 vdd.n1592 vdd.n1590 585
R667 vdd.n1615 vdd.n1614 585
R668 vdd.n1613 vdd.n1612 585
R669 vdd.n1596 vdd.n1595 585
R670 vdd.n1607 vdd.n1606 585
R671 vdd.n1605 vdd.n1604 585
R672 vdd.n1600 vdd.n1599 585
R673 vdd.n1683 vdd.n1682 585
R674 vdd.n1681 vdd.n1648 585
R675 vdd.n1680 vdd.n1679 585
R676 vdd.n1651 vdd.n1649 585
R677 vdd.n1674 vdd.n1673 585
R678 vdd.n1672 vdd.n1671 585
R679 vdd.n1655 vdd.n1654 585
R680 vdd.n1666 vdd.n1665 585
R681 vdd.n1664 vdd.n1663 585
R682 vdd.n1659 vdd.n1658 585
R683 vdd.n3538 vdd.n392 509.269
R684 vdd.n3534 vdd.n393 509.269
R685 vdd.n3406 vdd.n685 509.269
R686 vdd.n3403 vdd.n684 509.269
R687 vdd.n2195 vdd.n1155 509.269
R688 vdd.n2198 vdd.n2197 509.269
R689 vdd.n1304 vdd.n1268 509.269
R690 vdd.n1500 vdd.n1269 509.269
R691 vdd.n305 vdd.t142 329.043
R692 vdd.n246 vdd.t219 329.043
R693 vdd.n203 vdd.t145 329.043
R694 vdd.n144 vdd.t199 329.043
R695 vdd.n102 vdd.t244 329.043
R696 vdd.n43 vdd.t268 329.043
R697 vdd.n1804 vdd.t298 329.043
R698 vdd.n1863 vdd.t249 329.043
R699 vdd.n1702 vdd.t282 329.043
R700 vdd.n1761 vdd.t235 329.043
R701 vdd.n1601 vdd.t239 329.043
R702 vdd.n1660 vdd.t246 329.043
R703 vdd.n1397 vdd.t108 319.788
R704 vdd.n1435 vdd.t119 319.788
R705 vdd.n1331 vdd.t132 319.788
R706 vdd.n2200 vdd.t91 319.788
R707 vdd.n2050 vdd.t100 319.788
R708 vdd.n2010 vdd.t121 319.788
R709 vdd.n426 vdd.t103 319.788
R710 vdd.n440 vdd.t77 319.788
R711 vdd.n452 vdd.t94 319.788
R712 vdd.n768 vdd.t66 319.788
R713 vdd.n3366 vdd.t81 319.788
R714 vdd.n688 vdd.t88 319.788
R715 vdd.n1398 vdd.t107 303.69
R716 vdd.n1436 vdd.t118 303.69
R717 vdd.n1332 vdd.t131 303.69
R718 vdd.n2201 vdd.t92 303.69
R719 vdd.n2051 vdd.t101 303.69
R720 vdd.n2011 vdd.t122 303.69
R721 vdd.n427 vdd.t104 303.69
R722 vdd.n441 vdd.t78 303.69
R723 vdd.n453 vdd.t95 303.69
R724 vdd.n769 vdd.t65 303.69
R725 vdd.n3367 vdd.t80 303.69
R726 vdd.n689 vdd.t87 303.69
R727 vdd.n3016 vdd.n947 285.366
R728 vdd.n3240 vdd.n809 285.366
R729 vdd.n3177 vdd.n806 285.366
R730 vdd.n2895 vdd.n944 285.366
R731 vdd.n2725 vdd.n985 285.366
R732 vdd.n2656 vdd.n2655 285.366
R733 vdd.n2396 vdd.n1111 285.366
R734 vdd.n2466 vdd.n1113 285.366
R735 vdd.n3156 vdd.n807 285.366
R736 vdd.n3243 vdd.n3242 285.366
R737 vdd.n3009 vdd.n945 285.366
R738 vdd.n3018 vdd.n943 285.366
R739 vdd.n2653 vdd.n995 285.366
R740 vdd.n993 vdd.n967 285.366
R741 vdd.n2282 vdd.n1112 285.366
R742 vdd.n2468 vdd.n1109 285.366
R743 vdd.n1153 vdd.n1110 216.982
R744 vdd.n3405 vdd.n692 216.982
R745 vdd.n3158 vdd.n807 185
R746 vdd.n3241 vdd.n807 185
R747 vdd.n3160 vdd.n3159 185
R748 vdd.n3159 vdd.n805 185
R749 vdd.n3161 vdd.n839 185
R750 vdd.n3171 vdd.n839 185
R751 vdd.n3162 vdd.n848 185
R752 vdd.n848 vdd.n846 185
R753 vdd.n3164 vdd.n3163 185
R754 vdd.n3165 vdd.n3164 185
R755 vdd.n3117 vdd.n847 185
R756 vdd.n847 vdd.n843 185
R757 vdd.n3116 vdd.n3115 185
R758 vdd.n3115 vdd.n3114 185
R759 vdd.n850 vdd.n849 185
R760 vdd.n851 vdd.n850 185
R761 vdd.n3107 vdd.n3106 185
R762 vdd.n3108 vdd.n3107 185
R763 vdd.n3105 vdd.n859 185
R764 vdd.n864 vdd.n859 185
R765 vdd.n3104 vdd.n3103 185
R766 vdd.n3103 vdd.n3102 185
R767 vdd.n861 vdd.n860 185
R768 vdd.n870 vdd.n861 185
R769 vdd.n3095 vdd.n3094 185
R770 vdd.n3096 vdd.n3095 185
R771 vdd.n3093 vdd.n871 185
R772 vdd.n877 vdd.n871 185
R773 vdd.n3092 vdd.n3091 185
R774 vdd.n3091 vdd.n3090 185
R775 vdd.n873 vdd.n872 185
R776 vdd.n874 vdd.n873 185
R777 vdd.n3083 vdd.n3082 185
R778 vdd.n3084 vdd.n3083 185
R779 vdd.n3081 vdd.n884 185
R780 vdd.n884 vdd.n881 185
R781 vdd.n3079 vdd.n3078 185
R782 vdd.n3078 vdd.n3077 185
R783 vdd.n887 vdd.n886 185
R784 vdd.n888 vdd.n887 185
R785 vdd.n3070 vdd.n3069 185
R786 vdd.n3071 vdd.n3070 185
R787 vdd.n3068 vdd.n896 185
R788 vdd.n901 vdd.n896 185
R789 vdd.n3067 vdd.n3066 185
R790 vdd.n3066 vdd.n3065 185
R791 vdd.n898 vdd.n897 185
R792 vdd.n2977 vdd.n898 185
R793 vdd.n3058 vdd.n3057 185
R794 vdd.n3059 vdd.n3058 185
R795 vdd.n3056 vdd.n908 185
R796 vdd.n908 vdd.n905 185
R797 vdd.n3055 vdd.n3054 185
R798 vdd.n3054 vdd.n3053 185
R799 vdd.n910 vdd.n909 185
R800 vdd.n911 vdd.n910 185
R801 vdd.n3046 vdd.n3045 185
R802 vdd.n3047 vdd.n3046 185
R803 vdd.n3044 vdd.n919 185
R804 vdd.n2989 vdd.n919 185
R805 vdd.n3043 vdd.n3042 185
R806 vdd.n3042 vdd.n3041 185
R807 vdd.n921 vdd.n920 185
R808 vdd.n930 vdd.n921 185
R809 vdd.n3034 vdd.n3033 185
R810 vdd.n3035 vdd.n3034 185
R811 vdd.n3032 vdd.n931 185
R812 vdd.n931 vdd.n927 185
R813 vdd.n3031 vdd.n3030 185
R814 vdd.n3030 vdd.n3029 185
R815 vdd.n933 vdd.n932 185
R816 vdd.n3001 vdd.n933 185
R817 vdd.n3022 vdd.n3021 185
R818 vdd.n3023 vdd.n3022 185
R819 vdd.n3020 vdd.n941 185
R820 vdd.n946 vdd.n941 185
R821 vdd.n3019 vdd.n3018 185
R822 vdd.n3018 vdd.n3017 185
R823 vdd.n943 vdd.n942 185
R824 vdd.n2765 vdd.n2764 185
R825 vdd.n2767 vdd.n2766 185
R826 vdd.n2769 vdd.n2768 185
R827 vdd.n2771 vdd.n2770 185
R828 vdd.n2773 vdd.n2772 185
R829 vdd.n2775 vdd.n2774 185
R830 vdd.n2777 vdd.n2776 185
R831 vdd.n2779 vdd.n2778 185
R832 vdd.n2781 vdd.n2780 185
R833 vdd.n2783 vdd.n2782 185
R834 vdd.n2785 vdd.n2784 185
R835 vdd.n2787 vdd.n2786 185
R836 vdd.n2789 vdd.n2788 185
R837 vdd.n2791 vdd.n2790 185
R838 vdd.n2793 vdd.n2792 185
R839 vdd.n2795 vdd.n2794 185
R840 vdd.n2797 vdd.n2796 185
R841 vdd.n2799 vdd.n2798 185
R842 vdd.n2801 vdd.n2800 185
R843 vdd.n2803 vdd.n2802 185
R844 vdd.n2805 vdd.n2804 185
R845 vdd.n2807 vdd.n2806 185
R846 vdd.n2809 vdd.n2808 185
R847 vdd.n2811 vdd.n2810 185
R848 vdd.n2813 vdd.n2812 185
R849 vdd.n2815 vdd.n2814 185
R850 vdd.n2817 vdd.n2816 185
R851 vdd.n2819 vdd.n2818 185
R852 vdd.n2821 vdd.n2820 185
R853 vdd.n2823 vdd.n2822 185
R854 vdd.n2825 vdd.n2824 185
R855 vdd.n2827 vdd.n2826 185
R856 vdd.n2828 vdd.n2760 185
R857 vdd.n3009 vdd.n3008 185
R858 vdd.n3010 vdd.n3009 185
R859 vdd.n3244 vdd.n3243 185
R860 vdd.n3245 vdd.n798 185
R861 vdd.n3247 vdd.n3246 185
R862 vdd.n3249 vdd.n796 185
R863 vdd.n3251 vdd.n3250 185
R864 vdd.n3252 vdd.n795 185
R865 vdd.n3254 vdd.n3253 185
R866 vdd.n3256 vdd.n793 185
R867 vdd.n3258 vdd.n3257 185
R868 vdd.n3259 vdd.n792 185
R869 vdd.n3261 vdd.n3260 185
R870 vdd.n3263 vdd.n790 185
R871 vdd.n3265 vdd.n3264 185
R872 vdd.n3266 vdd.n789 185
R873 vdd.n3268 vdd.n3267 185
R874 vdd.n3270 vdd.n788 185
R875 vdd.n3271 vdd.n786 185
R876 vdd.n3274 vdd.n3273 185
R877 vdd.n787 vdd.n785 185
R878 vdd.n3130 vdd.n3129 185
R879 vdd.n3132 vdd.n3131 185
R880 vdd.n3134 vdd.n3126 185
R881 vdd.n3136 vdd.n3135 185
R882 vdd.n3137 vdd.n3125 185
R883 vdd.n3139 vdd.n3138 185
R884 vdd.n3141 vdd.n3123 185
R885 vdd.n3143 vdd.n3142 185
R886 vdd.n3144 vdd.n3122 185
R887 vdd.n3146 vdd.n3145 185
R888 vdd.n3148 vdd.n3120 185
R889 vdd.n3150 vdd.n3149 185
R890 vdd.n3151 vdd.n3119 185
R891 vdd.n3153 vdd.n3152 185
R892 vdd.n3155 vdd.n3118 185
R893 vdd.n3157 vdd.n3156 185
R894 vdd.n3156 vdd.n692 185
R895 vdd.n3242 vdd.n802 185
R896 vdd.n3242 vdd.n3241 185
R897 vdd.n2908 vdd.n804 185
R898 vdd.n805 vdd.n804 185
R899 vdd.n2909 vdd.n838 185
R900 vdd.n3171 vdd.n838 185
R901 vdd.n2911 vdd.n2910 185
R902 vdd.n2910 vdd.n846 185
R903 vdd.n2912 vdd.n845 185
R904 vdd.n3165 vdd.n845 185
R905 vdd.n2914 vdd.n2913 185
R906 vdd.n2913 vdd.n843 185
R907 vdd.n2915 vdd.n853 185
R908 vdd.n3114 vdd.n853 185
R909 vdd.n2917 vdd.n2916 185
R910 vdd.n2916 vdd.n851 185
R911 vdd.n2918 vdd.n858 185
R912 vdd.n3108 vdd.n858 185
R913 vdd.n2920 vdd.n2919 185
R914 vdd.n2919 vdd.n864 185
R915 vdd.n2921 vdd.n863 185
R916 vdd.n3102 vdd.n863 185
R917 vdd.n2923 vdd.n2922 185
R918 vdd.n2922 vdd.n870 185
R919 vdd.n2924 vdd.n869 185
R920 vdd.n3096 vdd.n869 185
R921 vdd.n2926 vdd.n2925 185
R922 vdd.n2925 vdd.n877 185
R923 vdd.n2927 vdd.n876 185
R924 vdd.n3090 vdd.n876 185
R925 vdd.n2929 vdd.n2928 185
R926 vdd.n2928 vdd.n874 185
R927 vdd.n2930 vdd.n883 185
R928 vdd.n3084 vdd.n883 185
R929 vdd.n2932 vdd.n2931 185
R930 vdd.n2931 vdd.n881 185
R931 vdd.n2933 vdd.n890 185
R932 vdd.n3077 vdd.n890 185
R933 vdd.n2935 vdd.n2934 185
R934 vdd.n2934 vdd.n888 185
R935 vdd.n2936 vdd.n895 185
R936 vdd.n3071 vdd.n895 185
R937 vdd.n2938 vdd.n2937 185
R938 vdd.n2937 vdd.n901 185
R939 vdd.n2939 vdd.n900 185
R940 vdd.n3065 vdd.n900 185
R941 vdd.n2979 vdd.n2978 185
R942 vdd.n2978 vdd.n2977 185
R943 vdd.n2980 vdd.n907 185
R944 vdd.n3059 vdd.n907 185
R945 vdd.n2982 vdd.n2981 185
R946 vdd.n2981 vdd.n905 185
R947 vdd.n2983 vdd.n913 185
R948 vdd.n3053 vdd.n913 185
R949 vdd.n2985 vdd.n2984 185
R950 vdd.n2984 vdd.n911 185
R951 vdd.n2986 vdd.n918 185
R952 vdd.n3047 vdd.n918 185
R953 vdd.n2988 vdd.n2987 185
R954 vdd.n2989 vdd.n2988 185
R955 vdd.n2907 vdd.n923 185
R956 vdd.n3041 vdd.n923 185
R957 vdd.n2906 vdd.n2905 185
R958 vdd.n2905 vdd.n930 185
R959 vdd.n2904 vdd.n929 185
R960 vdd.n3035 vdd.n929 185
R961 vdd.n2903 vdd.n2902 185
R962 vdd.n2902 vdd.n927 185
R963 vdd.n2829 vdd.n935 185
R964 vdd.n3029 vdd.n935 185
R965 vdd.n3003 vdd.n3002 185
R966 vdd.n3002 vdd.n3001 185
R967 vdd.n3004 vdd.n940 185
R968 vdd.n3023 vdd.n940 185
R969 vdd.n3006 vdd.n3005 185
R970 vdd.n3005 vdd.n946 185
R971 vdd.n3007 vdd.n945 185
R972 vdd.n3017 vdd.n945 185
R973 vdd.n2195 vdd.n2194 185
R974 vdd.n2196 vdd.n2195 185
R975 vdd.n1156 vdd.n1154 185
R976 vdd.n1974 vdd.n1154 185
R977 vdd.n1977 vdd.n1976 185
R978 vdd.n1976 vdd.n1975 185
R979 vdd.n1159 vdd.n1158 185
R980 vdd.n1160 vdd.n1159 185
R981 vdd.n1963 vdd.n1962 185
R982 vdd.n1964 vdd.n1963 185
R983 vdd.n1168 vdd.n1167 185
R984 vdd.n1955 vdd.n1167 185
R985 vdd.n1958 vdd.n1957 185
R986 vdd.n1957 vdd.n1956 185
R987 vdd.n1171 vdd.n1170 185
R988 vdd.n1178 vdd.n1171 185
R989 vdd.n1946 vdd.n1945 185
R990 vdd.n1947 vdd.n1946 185
R991 vdd.n1180 vdd.n1179 185
R992 vdd.n1179 vdd.n1177 185
R993 vdd.n1941 vdd.n1940 185
R994 vdd.n1940 vdd.n1939 185
R995 vdd.n1183 vdd.n1182 185
R996 vdd.n1184 vdd.n1183 185
R997 vdd.n1930 vdd.n1929 185
R998 vdd.n1931 vdd.n1930 185
R999 vdd.n1191 vdd.n1190 185
R1000 vdd.n1922 vdd.n1190 185
R1001 vdd.n1925 vdd.n1924 185
R1002 vdd.n1924 vdd.n1923 185
R1003 vdd.n1194 vdd.n1193 185
R1004 vdd.n1200 vdd.n1194 185
R1005 vdd.n1913 vdd.n1912 185
R1006 vdd.n1914 vdd.n1913 185
R1007 vdd.n1202 vdd.n1201 185
R1008 vdd.n1905 vdd.n1201 185
R1009 vdd.n1908 vdd.n1907 185
R1010 vdd.n1907 vdd.n1906 185
R1011 vdd.n1205 vdd.n1204 185
R1012 vdd.n1206 vdd.n1205 185
R1013 vdd.n1896 vdd.n1895 185
R1014 vdd.n1897 vdd.n1896 185
R1015 vdd.n1214 vdd.n1213 185
R1016 vdd.n1213 vdd.n1212 185
R1017 vdd.n1584 vdd.n1583 185
R1018 vdd.n1583 vdd.n1582 185
R1019 vdd.n1217 vdd.n1216 185
R1020 vdd.n1223 vdd.n1217 185
R1021 vdd.n1573 vdd.n1572 185
R1022 vdd.n1574 vdd.n1573 185
R1023 vdd.n1225 vdd.n1224 185
R1024 vdd.n1565 vdd.n1224 185
R1025 vdd.n1568 vdd.n1567 185
R1026 vdd.n1567 vdd.n1566 185
R1027 vdd.n1228 vdd.n1227 185
R1028 vdd.n1235 vdd.n1228 185
R1029 vdd.n1556 vdd.n1555 185
R1030 vdd.n1557 vdd.n1556 185
R1031 vdd.n1237 vdd.n1236 185
R1032 vdd.n1236 vdd.n1234 185
R1033 vdd.n1551 vdd.n1550 185
R1034 vdd.n1550 vdd.n1549 185
R1035 vdd.n1240 vdd.n1239 185
R1036 vdd.n1241 vdd.n1240 185
R1037 vdd.n1540 vdd.n1539 185
R1038 vdd.n1541 vdd.n1540 185
R1039 vdd.n1248 vdd.n1247 185
R1040 vdd.n1532 vdd.n1247 185
R1041 vdd.n1535 vdd.n1534 185
R1042 vdd.n1534 vdd.n1533 185
R1043 vdd.n1251 vdd.n1250 185
R1044 vdd.n1257 vdd.n1251 185
R1045 vdd.n1523 vdd.n1522 185
R1046 vdd.n1524 vdd.n1523 185
R1047 vdd.n1259 vdd.n1258 185
R1048 vdd.n1515 vdd.n1258 185
R1049 vdd.n1518 vdd.n1517 185
R1050 vdd.n1517 vdd.n1516 185
R1051 vdd.n1262 vdd.n1261 185
R1052 vdd.n1263 vdd.n1262 185
R1053 vdd.n1506 vdd.n1505 185
R1054 vdd.n1507 vdd.n1506 185
R1055 vdd.n1270 vdd.n1269 185
R1056 vdd.n1305 vdd.n1269 185
R1057 vdd.n1501 vdd.n1500 185
R1058 vdd.n1273 vdd.n1272 185
R1059 vdd.n1497 vdd.n1496 185
R1060 vdd.n1498 vdd.n1497 185
R1061 vdd.n1307 vdd.n1306 185
R1062 vdd.n1492 vdd.n1309 185
R1063 vdd.n1491 vdd.n1310 185
R1064 vdd.n1490 vdd.n1311 185
R1065 vdd.n1313 vdd.n1312 185
R1066 vdd.n1486 vdd.n1315 185
R1067 vdd.n1485 vdd.n1316 185
R1068 vdd.n1484 vdd.n1317 185
R1069 vdd.n1319 vdd.n1318 185
R1070 vdd.n1480 vdd.n1321 185
R1071 vdd.n1479 vdd.n1322 185
R1072 vdd.n1478 vdd.n1323 185
R1073 vdd.n1325 vdd.n1324 185
R1074 vdd.n1474 vdd.n1327 185
R1075 vdd.n1473 vdd.n1328 185
R1076 vdd.n1472 vdd.n1329 185
R1077 vdd.n1333 vdd.n1330 185
R1078 vdd.n1468 vdd.n1335 185
R1079 vdd.n1467 vdd.n1336 185
R1080 vdd.n1466 vdd.n1337 185
R1081 vdd.n1339 vdd.n1338 185
R1082 vdd.n1462 vdd.n1341 185
R1083 vdd.n1461 vdd.n1342 185
R1084 vdd.n1460 vdd.n1343 185
R1085 vdd.n1345 vdd.n1344 185
R1086 vdd.n1456 vdd.n1347 185
R1087 vdd.n1455 vdd.n1348 185
R1088 vdd.n1454 vdd.n1349 185
R1089 vdd.n1351 vdd.n1350 185
R1090 vdd.n1450 vdd.n1353 185
R1091 vdd.n1449 vdd.n1354 185
R1092 vdd.n1448 vdd.n1355 185
R1093 vdd.n1357 vdd.n1356 185
R1094 vdd.n1444 vdd.n1359 185
R1095 vdd.n1443 vdd.n1360 185
R1096 vdd.n1442 vdd.n1361 185
R1097 vdd.n1363 vdd.n1362 185
R1098 vdd.n1438 vdd.n1365 185
R1099 vdd.n1437 vdd.n1434 185
R1100 vdd.n1433 vdd.n1366 185
R1101 vdd.n1368 vdd.n1367 185
R1102 vdd.n1429 vdd.n1370 185
R1103 vdd.n1428 vdd.n1371 185
R1104 vdd.n1427 vdd.n1372 185
R1105 vdd.n1374 vdd.n1373 185
R1106 vdd.n1423 vdd.n1376 185
R1107 vdd.n1422 vdd.n1377 185
R1108 vdd.n1421 vdd.n1378 185
R1109 vdd.n1380 vdd.n1379 185
R1110 vdd.n1417 vdd.n1382 185
R1111 vdd.n1416 vdd.n1383 185
R1112 vdd.n1415 vdd.n1384 185
R1113 vdd.n1386 vdd.n1385 185
R1114 vdd.n1411 vdd.n1388 185
R1115 vdd.n1410 vdd.n1389 185
R1116 vdd.n1409 vdd.n1390 185
R1117 vdd.n1392 vdd.n1391 185
R1118 vdd.n1405 vdd.n1394 185
R1119 vdd.n1404 vdd.n1395 185
R1120 vdd.n1403 vdd.n1396 185
R1121 vdd.n1400 vdd.n1304 185
R1122 vdd.n1498 vdd.n1304 185
R1123 vdd.n2199 vdd.n2198 185
R1124 vdd.n2203 vdd.n1149 185
R1125 vdd.n2079 vdd.n1148 185
R1126 vdd.n2082 vdd.n2081 185
R1127 vdd.n2084 vdd.n2083 185
R1128 vdd.n2087 vdd.n2086 185
R1129 vdd.n2089 vdd.n2088 185
R1130 vdd.n2091 vdd.n2077 185
R1131 vdd.n2093 vdd.n2092 185
R1132 vdd.n2094 vdd.n2071 185
R1133 vdd.n2096 vdd.n2095 185
R1134 vdd.n2098 vdd.n2069 185
R1135 vdd.n2100 vdd.n2099 185
R1136 vdd.n2101 vdd.n2064 185
R1137 vdd.n2103 vdd.n2102 185
R1138 vdd.n2105 vdd.n2062 185
R1139 vdd.n2107 vdd.n2106 185
R1140 vdd.n2108 vdd.n2058 185
R1141 vdd.n2110 vdd.n2109 185
R1142 vdd.n2112 vdd.n2055 185
R1143 vdd.n2114 vdd.n2113 185
R1144 vdd.n2056 vdd.n2049 185
R1145 vdd.n2118 vdd.n2053 185
R1146 vdd.n2119 vdd.n2045 185
R1147 vdd.n2121 vdd.n2120 185
R1148 vdd.n2123 vdd.n2043 185
R1149 vdd.n2125 vdd.n2124 185
R1150 vdd.n2126 vdd.n2038 185
R1151 vdd.n2128 vdd.n2127 185
R1152 vdd.n2130 vdd.n2036 185
R1153 vdd.n2132 vdd.n2131 185
R1154 vdd.n2133 vdd.n2031 185
R1155 vdd.n2135 vdd.n2134 185
R1156 vdd.n2137 vdd.n2029 185
R1157 vdd.n2139 vdd.n2138 185
R1158 vdd.n2140 vdd.n2024 185
R1159 vdd.n2142 vdd.n2141 185
R1160 vdd.n2144 vdd.n2022 185
R1161 vdd.n2146 vdd.n2145 185
R1162 vdd.n2147 vdd.n2018 185
R1163 vdd.n2149 vdd.n2148 185
R1164 vdd.n2151 vdd.n2015 185
R1165 vdd.n2153 vdd.n2152 185
R1166 vdd.n2016 vdd.n2009 185
R1167 vdd.n2157 vdd.n2013 185
R1168 vdd.n2158 vdd.n2005 185
R1169 vdd.n2160 vdd.n2159 185
R1170 vdd.n2162 vdd.n2003 185
R1171 vdd.n2164 vdd.n2163 185
R1172 vdd.n2165 vdd.n1998 185
R1173 vdd.n2167 vdd.n2166 185
R1174 vdd.n2169 vdd.n1996 185
R1175 vdd.n2171 vdd.n2170 185
R1176 vdd.n2172 vdd.n1991 185
R1177 vdd.n2174 vdd.n2173 185
R1178 vdd.n2176 vdd.n1990 185
R1179 vdd.n2177 vdd.n1987 185
R1180 vdd.n2180 vdd.n2179 185
R1181 vdd.n1989 vdd.n1985 185
R1182 vdd.n2184 vdd.n1983 185
R1183 vdd.n2186 vdd.n2185 185
R1184 vdd.n2188 vdd.n1981 185
R1185 vdd.n2190 vdd.n2189 185
R1186 vdd.n2191 vdd.n1155 185
R1187 vdd.n2197 vdd.n1152 185
R1188 vdd.n2197 vdd.n2196 185
R1189 vdd.n1163 vdd.n1151 185
R1190 vdd.n1974 vdd.n1151 185
R1191 vdd.n1973 vdd.n1972 185
R1192 vdd.n1975 vdd.n1973 185
R1193 vdd.n1162 vdd.n1161 185
R1194 vdd.n1161 vdd.n1160 185
R1195 vdd.n1966 vdd.n1965 185
R1196 vdd.n1965 vdd.n1964 185
R1197 vdd.n1166 vdd.n1165 185
R1198 vdd.n1955 vdd.n1166 185
R1199 vdd.n1954 vdd.n1953 185
R1200 vdd.n1956 vdd.n1954 185
R1201 vdd.n1173 vdd.n1172 185
R1202 vdd.n1178 vdd.n1172 185
R1203 vdd.n1949 vdd.n1948 185
R1204 vdd.n1948 vdd.n1947 185
R1205 vdd.n1176 vdd.n1175 185
R1206 vdd.n1177 vdd.n1176 185
R1207 vdd.n1938 vdd.n1937 185
R1208 vdd.n1939 vdd.n1938 185
R1209 vdd.n1186 vdd.n1185 185
R1210 vdd.n1185 vdd.n1184 185
R1211 vdd.n1933 vdd.n1932 185
R1212 vdd.n1932 vdd.n1931 185
R1213 vdd.n1189 vdd.n1188 185
R1214 vdd.n1922 vdd.n1189 185
R1215 vdd.n1921 vdd.n1920 185
R1216 vdd.n1923 vdd.n1921 185
R1217 vdd.n1196 vdd.n1195 185
R1218 vdd.n1200 vdd.n1195 185
R1219 vdd.n1916 vdd.n1915 185
R1220 vdd.n1915 vdd.n1914 185
R1221 vdd.n1199 vdd.n1198 185
R1222 vdd.n1905 vdd.n1199 185
R1223 vdd.n1904 vdd.n1903 185
R1224 vdd.n1906 vdd.n1904 185
R1225 vdd.n1208 vdd.n1207 185
R1226 vdd.n1207 vdd.n1206 185
R1227 vdd.n1899 vdd.n1898 185
R1228 vdd.n1898 vdd.n1897 185
R1229 vdd.n1211 vdd.n1210 185
R1230 vdd.n1212 vdd.n1211 185
R1231 vdd.n1581 vdd.n1580 185
R1232 vdd.n1582 vdd.n1581 185
R1233 vdd.n1219 vdd.n1218 185
R1234 vdd.n1223 vdd.n1218 185
R1235 vdd.n1576 vdd.n1575 185
R1236 vdd.n1575 vdd.n1574 185
R1237 vdd.n1222 vdd.n1221 185
R1238 vdd.n1565 vdd.n1222 185
R1239 vdd.n1564 vdd.n1563 185
R1240 vdd.n1566 vdd.n1564 185
R1241 vdd.n1230 vdd.n1229 185
R1242 vdd.n1235 vdd.n1229 185
R1243 vdd.n1559 vdd.n1558 185
R1244 vdd.n1558 vdd.n1557 185
R1245 vdd.n1233 vdd.n1232 185
R1246 vdd.n1234 vdd.n1233 185
R1247 vdd.n1548 vdd.n1547 185
R1248 vdd.n1549 vdd.n1548 185
R1249 vdd.n1243 vdd.n1242 185
R1250 vdd.n1242 vdd.n1241 185
R1251 vdd.n1543 vdd.n1542 185
R1252 vdd.n1542 vdd.n1541 185
R1253 vdd.n1246 vdd.n1245 185
R1254 vdd.n1532 vdd.n1246 185
R1255 vdd.n1531 vdd.n1530 185
R1256 vdd.n1533 vdd.n1531 185
R1257 vdd.n1253 vdd.n1252 185
R1258 vdd.n1257 vdd.n1252 185
R1259 vdd.n1526 vdd.n1525 185
R1260 vdd.n1525 vdd.n1524 185
R1261 vdd.n1256 vdd.n1255 185
R1262 vdd.n1515 vdd.n1256 185
R1263 vdd.n1514 vdd.n1513 185
R1264 vdd.n1516 vdd.n1514 185
R1265 vdd.n1265 vdd.n1264 185
R1266 vdd.n1264 vdd.n1263 185
R1267 vdd.n1509 vdd.n1508 185
R1268 vdd.n1508 vdd.n1507 185
R1269 vdd.n1268 vdd.n1267 185
R1270 vdd.n1305 vdd.n1268 185
R1271 vdd.n987 vdd.n985 185
R1272 vdd.n2654 vdd.n985 185
R1273 vdd.n2576 vdd.n1005 185
R1274 vdd.n1005 vdd.n992 185
R1275 vdd.n2578 vdd.n2577 185
R1276 vdd.n2579 vdd.n2578 185
R1277 vdd.n2575 vdd.n1004 185
R1278 vdd.n2334 vdd.n1004 185
R1279 vdd.n2574 vdd.n2573 185
R1280 vdd.n2573 vdd.n2572 185
R1281 vdd.n1007 vdd.n1006 185
R1282 vdd.n1008 vdd.n1007 185
R1283 vdd.n2563 vdd.n2562 185
R1284 vdd.n2564 vdd.n2563 185
R1285 vdd.n2561 vdd.n1018 185
R1286 vdd.n1018 vdd.n1015 185
R1287 vdd.n2560 vdd.n2559 185
R1288 vdd.n2559 vdd.n2558 185
R1289 vdd.n1020 vdd.n1019 185
R1290 vdd.n2346 vdd.n1020 185
R1291 vdd.n2551 vdd.n2550 185
R1292 vdd.n2552 vdd.n2551 185
R1293 vdd.n2549 vdd.n1028 185
R1294 vdd.n1033 vdd.n1028 185
R1295 vdd.n2548 vdd.n2547 185
R1296 vdd.n2547 vdd.n2546 185
R1297 vdd.n1030 vdd.n1029 185
R1298 vdd.n1039 vdd.n1030 185
R1299 vdd.n2539 vdd.n2538 185
R1300 vdd.n2540 vdd.n2539 185
R1301 vdd.n2537 vdd.n1040 185
R1302 vdd.n2358 vdd.n1040 185
R1303 vdd.n2536 vdd.n2535 185
R1304 vdd.n2535 vdd.n2534 185
R1305 vdd.n1042 vdd.n1041 185
R1306 vdd.n1043 vdd.n1042 185
R1307 vdd.n2527 vdd.n2526 185
R1308 vdd.n2528 vdd.n2527 185
R1309 vdd.n2525 vdd.n1052 185
R1310 vdd.n1052 vdd.n1049 185
R1311 vdd.n2524 vdd.n2523 185
R1312 vdd.n2523 vdd.n2522 185
R1313 vdd.n1054 vdd.n1053 185
R1314 vdd.n1063 vdd.n1054 185
R1315 vdd.n2514 vdd.n2513 185
R1316 vdd.n2515 vdd.n2514 185
R1317 vdd.n2512 vdd.n1064 185
R1318 vdd.n1070 vdd.n1064 185
R1319 vdd.n2511 vdd.n2510 185
R1320 vdd.n2510 vdd.n2509 185
R1321 vdd.n1066 vdd.n1065 185
R1322 vdd.n1067 vdd.n1066 185
R1323 vdd.n2502 vdd.n2501 185
R1324 vdd.n2503 vdd.n2502 185
R1325 vdd.n2500 vdd.n1077 185
R1326 vdd.n1077 vdd.n1074 185
R1327 vdd.n2499 vdd.n2498 185
R1328 vdd.n2498 vdd.n2497 185
R1329 vdd.n1079 vdd.n1078 185
R1330 vdd.n1080 vdd.n1079 185
R1331 vdd.n2490 vdd.n2489 185
R1332 vdd.n2491 vdd.n2490 185
R1333 vdd.n2488 vdd.n1089 185
R1334 vdd.n1089 vdd.n1086 185
R1335 vdd.n2487 vdd.n2486 185
R1336 vdd.n2486 vdd.n2485 185
R1337 vdd.n1091 vdd.n1090 185
R1338 vdd.n1092 vdd.n1091 185
R1339 vdd.n2478 vdd.n2477 185
R1340 vdd.n2479 vdd.n2478 185
R1341 vdd.n2476 vdd.n1101 185
R1342 vdd.n1101 vdd.n1098 185
R1343 vdd.n2475 vdd.n2474 185
R1344 vdd.n2474 vdd.n2473 185
R1345 vdd.n1103 vdd.n1102 185
R1346 vdd.n1104 vdd.n1103 185
R1347 vdd.n2466 vdd.n2465 185
R1348 vdd.n2467 vdd.n2466 185
R1349 vdd.n2464 vdd.n1113 185
R1350 vdd.n2463 vdd.n2462 185
R1351 vdd.n2460 vdd.n1114 185
R1352 vdd.n2460 vdd.n1110 185
R1353 vdd.n2459 vdd.n2458 185
R1354 vdd.n2457 vdd.n2456 185
R1355 vdd.n2455 vdd.n1116 185
R1356 vdd.n2453 vdd.n2452 185
R1357 vdd.n2451 vdd.n1117 185
R1358 vdd.n2450 vdd.n2449 185
R1359 vdd.n2447 vdd.n1118 185
R1360 vdd.n2445 vdd.n2444 185
R1361 vdd.n2443 vdd.n1119 185
R1362 vdd.n2442 vdd.n2441 185
R1363 vdd.n2439 vdd.n1120 185
R1364 vdd.n2437 vdd.n2436 185
R1365 vdd.n2435 vdd.n1121 185
R1366 vdd.n2434 vdd.n2433 185
R1367 vdd.n2431 vdd.n1122 185
R1368 vdd.n2429 vdd.n2428 185
R1369 vdd.n2427 vdd.n1123 185
R1370 vdd.n2426 vdd.n2425 185
R1371 vdd.n2423 vdd.n1124 185
R1372 vdd.n2421 vdd.n2420 185
R1373 vdd.n2419 vdd.n1125 185
R1374 vdd.n2418 vdd.n2417 185
R1375 vdd.n2415 vdd.n1126 185
R1376 vdd.n2413 vdd.n2412 185
R1377 vdd.n2411 vdd.n1127 185
R1378 vdd.n2410 vdd.n2409 185
R1379 vdd.n2407 vdd.n1128 185
R1380 vdd.n2405 vdd.n2404 185
R1381 vdd.n2403 vdd.n1129 185
R1382 vdd.n2401 vdd.n2400 185
R1383 vdd.n2398 vdd.n1132 185
R1384 vdd.n2396 vdd.n2395 185
R1385 vdd.n2657 vdd.n2656 185
R1386 vdd.n2659 vdd.n2658 185
R1387 vdd.n2661 vdd.n2660 185
R1388 vdd.n2664 vdd.n2663 185
R1389 vdd.n2666 vdd.n2665 185
R1390 vdd.n2668 vdd.n2667 185
R1391 vdd.n2670 vdd.n2669 185
R1392 vdd.n2672 vdd.n2671 185
R1393 vdd.n2674 vdd.n2673 185
R1394 vdd.n2676 vdd.n2675 185
R1395 vdd.n2678 vdd.n2677 185
R1396 vdd.n2680 vdd.n2679 185
R1397 vdd.n2682 vdd.n2681 185
R1398 vdd.n2684 vdd.n2683 185
R1399 vdd.n2686 vdd.n2685 185
R1400 vdd.n2688 vdd.n2687 185
R1401 vdd.n2690 vdd.n2689 185
R1402 vdd.n2692 vdd.n2691 185
R1403 vdd.n2694 vdd.n2693 185
R1404 vdd.n2696 vdd.n2695 185
R1405 vdd.n2698 vdd.n2697 185
R1406 vdd.n2700 vdd.n2699 185
R1407 vdd.n2702 vdd.n2701 185
R1408 vdd.n2704 vdd.n2703 185
R1409 vdd.n2706 vdd.n2705 185
R1410 vdd.n2708 vdd.n2707 185
R1411 vdd.n2710 vdd.n2709 185
R1412 vdd.n2712 vdd.n2711 185
R1413 vdd.n2714 vdd.n2713 185
R1414 vdd.n2716 vdd.n2715 185
R1415 vdd.n2718 vdd.n2717 185
R1416 vdd.n2720 vdd.n2719 185
R1417 vdd.n2722 vdd.n2721 185
R1418 vdd.n2723 vdd.n986 185
R1419 vdd.n2725 vdd.n2724 185
R1420 vdd.n2726 vdd.n2725 185
R1421 vdd.n2655 vdd.n990 185
R1422 vdd.n2655 vdd.n2654 185
R1423 vdd.n2332 vdd.n991 185
R1424 vdd.n992 vdd.n991 185
R1425 vdd.n2333 vdd.n1002 185
R1426 vdd.n2579 vdd.n1002 185
R1427 vdd.n2336 vdd.n2335 185
R1428 vdd.n2335 vdd.n2334 185
R1429 vdd.n2337 vdd.n1009 185
R1430 vdd.n2572 vdd.n1009 185
R1431 vdd.n2339 vdd.n2338 185
R1432 vdd.n2338 vdd.n1008 185
R1433 vdd.n2340 vdd.n1016 185
R1434 vdd.n2564 vdd.n1016 185
R1435 vdd.n2342 vdd.n2341 185
R1436 vdd.n2341 vdd.n1015 185
R1437 vdd.n2343 vdd.n1021 185
R1438 vdd.n2558 vdd.n1021 185
R1439 vdd.n2345 vdd.n2344 185
R1440 vdd.n2346 vdd.n2345 185
R1441 vdd.n2331 vdd.n1026 185
R1442 vdd.n2552 vdd.n1026 185
R1443 vdd.n2330 vdd.n2329 185
R1444 vdd.n2329 vdd.n1033 185
R1445 vdd.n2328 vdd.n1031 185
R1446 vdd.n2546 vdd.n1031 185
R1447 vdd.n2327 vdd.n2326 185
R1448 vdd.n2326 vdd.n1039 185
R1449 vdd.n1133 vdd.n1037 185
R1450 vdd.n2540 vdd.n1037 185
R1451 vdd.n2360 vdd.n2359 185
R1452 vdd.n2359 vdd.n2358 185
R1453 vdd.n2361 vdd.n1044 185
R1454 vdd.n2534 vdd.n1044 185
R1455 vdd.n2363 vdd.n2362 185
R1456 vdd.n2362 vdd.n1043 185
R1457 vdd.n2364 vdd.n1050 185
R1458 vdd.n2528 vdd.n1050 185
R1459 vdd.n2366 vdd.n2365 185
R1460 vdd.n2365 vdd.n1049 185
R1461 vdd.n2367 vdd.n1055 185
R1462 vdd.n2522 vdd.n1055 185
R1463 vdd.n2369 vdd.n2368 185
R1464 vdd.n2368 vdd.n1063 185
R1465 vdd.n2370 vdd.n1061 185
R1466 vdd.n2515 vdd.n1061 185
R1467 vdd.n2372 vdd.n2371 185
R1468 vdd.n2371 vdd.n1070 185
R1469 vdd.n2373 vdd.n1068 185
R1470 vdd.n2509 vdd.n1068 185
R1471 vdd.n2375 vdd.n2374 185
R1472 vdd.n2374 vdd.n1067 185
R1473 vdd.n2376 vdd.n1075 185
R1474 vdd.n2503 vdd.n1075 185
R1475 vdd.n2378 vdd.n2377 185
R1476 vdd.n2377 vdd.n1074 185
R1477 vdd.n2379 vdd.n1081 185
R1478 vdd.n2497 vdd.n1081 185
R1479 vdd.n2381 vdd.n2380 185
R1480 vdd.n2380 vdd.n1080 185
R1481 vdd.n2382 vdd.n1087 185
R1482 vdd.n2491 vdd.n1087 185
R1483 vdd.n2384 vdd.n2383 185
R1484 vdd.n2383 vdd.n1086 185
R1485 vdd.n2385 vdd.n1093 185
R1486 vdd.n2485 vdd.n1093 185
R1487 vdd.n2387 vdd.n2386 185
R1488 vdd.n2386 vdd.n1092 185
R1489 vdd.n2388 vdd.n1099 185
R1490 vdd.n2479 vdd.n1099 185
R1491 vdd.n2390 vdd.n2389 185
R1492 vdd.n2389 vdd.n1098 185
R1493 vdd.n2391 vdd.n1105 185
R1494 vdd.n2473 vdd.n1105 185
R1495 vdd.n2393 vdd.n2392 185
R1496 vdd.n2392 vdd.n1104 185
R1497 vdd.n2394 vdd.n1111 185
R1498 vdd.n2467 vdd.n1111 185
R1499 vdd.n3539 vdd.n3538 185
R1500 vdd.n3538 vdd.n3537 185
R1501 vdd.n3540 vdd.n387 185
R1502 vdd.n387 vdd.n386 185
R1503 vdd.n3542 vdd.n3541 185
R1504 vdd.n3543 vdd.n3542 185
R1505 vdd.n382 vdd.n381 185
R1506 vdd.n3544 vdd.n382 185
R1507 vdd.n3547 vdd.n3546 185
R1508 vdd.n3546 vdd.n3545 185
R1509 vdd.n3548 vdd.n376 185
R1510 vdd.n376 vdd.n375 185
R1511 vdd.n3550 vdd.n3549 185
R1512 vdd.n3551 vdd.n3550 185
R1513 vdd.n371 vdd.n370 185
R1514 vdd.n3552 vdd.n371 185
R1515 vdd.n3555 vdd.n3554 185
R1516 vdd.n3554 vdd.n3553 185
R1517 vdd.n3556 vdd.n365 185
R1518 vdd.n3513 vdd.n365 185
R1519 vdd.n3558 vdd.n3557 185
R1520 vdd.n3559 vdd.n3558 185
R1521 vdd.n360 vdd.n359 185
R1522 vdd.n3560 vdd.n360 185
R1523 vdd.n3563 vdd.n3562 185
R1524 vdd.n3562 vdd.n3561 185
R1525 vdd.n3564 vdd.n354 185
R1526 vdd.n361 vdd.n354 185
R1527 vdd.n3566 vdd.n3565 185
R1528 vdd.n3567 vdd.n3566 185
R1529 vdd.n350 vdd.n349 185
R1530 vdd.n3568 vdd.n350 185
R1531 vdd.n3571 vdd.n3570 185
R1532 vdd.n3570 vdd.n3569 185
R1533 vdd.n3572 vdd.n345 185
R1534 vdd.n345 vdd.n344 185
R1535 vdd.n3574 vdd.n3573 185
R1536 vdd.n3575 vdd.n3574 185
R1537 vdd.n339 vdd.n337 185
R1538 vdd.n3576 vdd.n339 185
R1539 vdd.n3579 vdd.n3578 185
R1540 vdd.n3578 vdd.n3577 185
R1541 vdd.n338 vdd.n336 185
R1542 vdd.n340 vdd.n338 185
R1543 vdd.n3489 vdd.n3488 185
R1544 vdd.n3490 vdd.n3489 185
R1545 vdd.n635 vdd.n634 185
R1546 vdd.n634 vdd.n633 185
R1547 vdd.n3484 vdd.n3483 185
R1548 vdd.n3483 vdd.n3482 185
R1549 vdd.n638 vdd.n637 185
R1550 vdd.n644 vdd.n638 185
R1551 vdd.n3470 vdd.n3469 185
R1552 vdd.n3471 vdd.n3470 185
R1553 vdd.n646 vdd.n645 185
R1554 vdd.n3462 vdd.n645 185
R1555 vdd.n3465 vdd.n3464 185
R1556 vdd.n3464 vdd.n3463 185
R1557 vdd.n649 vdd.n648 185
R1558 vdd.n656 vdd.n649 185
R1559 vdd.n3453 vdd.n3452 185
R1560 vdd.n3454 vdd.n3453 185
R1561 vdd.n658 vdd.n657 185
R1562 vdd.n657 vdd.n655 185
R1563 vdd.n3448 vdd.n3447 185
R1564 vdd.n3447 vdd.n3446 185
R1565 vdd.n661 vdd.n660 185
R1566 vdd.n662 vdd.n661 185
R1567 vdd.n3437 vdd.n3436 185
R1568 vdd.n3438 vdd.n3437 185
R1569 vdd.n669 vdd.n668 185
R1570 vdd.n3429 vdd.n668 185
R1571 vdd.n3432 vdd.n3431 185
R1572 vdd.n3431 vdd.n3430 185
R1573 vdd.n672 vdd.n671 185
R1574 vdd.n679 vdd.n672 185
R1575 vdd.n3420 vdd.n3419 185
R1576 vdd.n3421 vdd.n3420 185
R1577 vdd.n681 vdd.n680 185
R1578 vdd.n680 vdd.n678 185
R1579 vdd.n3415 vdd.n3414 185
R1580 vdd.n3414 vdd.n3413 185
R1581 vdd.n684 vdd.n683 185
R1582 vdd.n723 vdd.n684 185
R1583 vdd.n3403 vdd.n3402 185
R1584 vdd.n3401 vdd.n725 185
R1585 vdd.n3400 vdd.n724 185
R1586 vdd.n3405 vdd.n724 185
R1587 vdd.n729 vdd.n728 185
R1588 vdd.n733 vdd.n732 185
R1589 vdd.n3396 vdd.n734 185
R1590 vdd.n3395 vdd.n3394 185
R1591 vdd.n3393 vdd.n3392 185
R1592 vdd.n3391 vdd.n3390 185
R1593 vdd.n3389 vdd.n3388 185
R1594 vdd.n3387 vdd.n3386 185
R1595 vdd.n3385 vdd.n3384 185
R1596 vdd.n3383 vdd.n3382 185
R1597 vdd.n3381 vdd.n3380 185
R1598 vdd.n3379 vdd.n3378 185
R1599 vdd.n3377 vdd.n3376 185
R1600 vdd.n3375 vdd.n3374 185
R1601 vdd.n3373 vdd.n3372 185
R1602 vdd.n3371 vdd.n3370 185
R1603 vdd.n3369 vdd.n3368 185
R1604 vdd.n3360 vdd.n747 185
R1605 vdd.n3362 vdd.n3361 185
R1606 vdd.n3359 vdd.n3358 185
R1607 vdd.n3357 vdd.n3356 185
R1608 vdd.n3355 vdd.n3354 185
R1609 vdd.n3353 vdd.n3352 185
R1610 vdd.n3351 vdd.n3350 185
R1611 vdd.n3349 vdd.n3348 185
R1612 vdd.n3347 vdd.n3346 185
R1613 vdd.n3345 vdd.n3344 185
R1614 vdd.n3343 vdd.n3342 185
R1615 vdd.n3341 vdd.n3340 185
R1616 vdd.n3339 vdd.n3338 185
R1617 vdd.n3337 vdd.n3336 185
R1618 vdd.n3335 vdd.n3334 185
R1619 vdd.n3333 vdd.n3332 185
R1620 vdd.n3331 vdd.n3330 185
R1621 vdd.n3329 vdd.n3328 185
R1622 vdd.n3327 vdd.n3326 185
R1623 vdd.n3325 vdd.n3324 185
R1624 vdd.n3323 vdd.n3322 185
R1625 vdd.n3321 vdd.n3320 185
R1626 vdd.n3314 vdd.n767 185
R1627 vdd.n3316 vdd.n3315 185
R1628 vdd.n3313 vdd.n3312 185
R1629 vdd.n3311 vdd.n3310 185
R1630 vdd.n3309 vdd.n3308 185
R1631 vdd.n3307 vdd.n3306 185
R1632 vdd.n3305 vdd.n3304 185
R1633 vdd.n3303 vdd.n3302 185
R1634 vdd.n3301 vdd.n3300 185
R1635 vdd.n3299 vdd.n3298 185
R1636 vdd.n3297 vdd.n3296 185
R1637 vdd.n3295 vdd.n3294 185
R1638 vdd.n3293 vdd.n3292 185
R1639 vdd.n3291 vdd.n3290 185
R1640 vdd.n3289 vdd.n3288 185
R1641 vdd.n3287 vdd.n3286 185
R1642 vdd.n3285 vdd.n3284 185
R1643 vdd.n3283 vdd.n3282 185
R1644 vdd.n3281 vdd.n3280 185
R1645 vdd.n3279 vdd.n3278 185
R1646 vdd.n3277 vdd.n691 185
R1647 vdd.n3407 vdd.n3406 185
R1648 vdd.n3406 vdd.n3405 185
R1649 vdd.n3534 vdd.n3533 185
R1650 vdd.n618 vdd.n425 185
R1651 vdd.n617 vdd.n616 185
R1652 vdd.n615 vdd.n614 185
R1653 vdd.n613 vdd.n430 185
R1654 vdd.n609 vdd.n608 185
R1655 vdd.n607 vdd.n606 185
R1656 vdd.n605 vdd.n604 185
R1657 vdd.n603 vdd.n432 185
R1658 vdd.n599 vdd.n598 185
R1659 vdd.n597 vdd.n596 185
R1660 vdd.n595 vdd.n594 185
R1661 vdd.n593 vdd.n434 185
R1662 vdd.n589 vdd.n588 185
R1663 vdd.n587 vdd.n586 185
R1664 vdd.n585 vdd.n584 185
R1665 vdd.n583 vdd.n436 185
R1666 vdd.n579 vdd.n578 185
R1667 vdd.n577 vdd.n576 185
R1668 vdd.n575 vdd.n574 185
R1669 vdd.n573 vdd.n438 185
R1670 vdd.n569 vdd.n568 185
R1671 vdd.n567 vdd.n566 185
R1672 vdd.n565 vdd.n564 185
R1673 vdd.n563 vdd.n442 185
R1674 vdd.n559 vdd.n558 185
R1675 vdd.n557 vdd.n556 185
R1676 vdd.n555 vdd.n554 185
R1677 vdd.n553 vdd.n444 185
R1678 vdd.n549 vdd.n548 185
R1679 vdd.n547 vdd.n546 185
R1680 vdd.n545 vdd.n544 185
R1681 vdd.n543 vdd.n446 185
R1682 vdd.n539 vdd.n538 185
R1683 vdd.n537 vdd.n536 185
R1684 vdd.n535 vdd.n534 185
R1685 vdd.n533 vdd.n448 185
R1686 vdd.n529 vdd.n528 185
R1687 vdd.n527 vdd.n526 185
R1688 vdd.n525 vdd.n524 185
R1689 vdd.n523 vdd.n450 185
R1690 vdd.n519 vdd.n518 185
R1691 vdd.n517 vdd.n516 185
R1692 vdd.n515 vdd.n514 185
R1693 vdd.n513 vdd.n454 185
R1694 vdd.n509 vdd.n508 185
R1695 vdd.n507 vdd.n506 185
R1696 vdd.n505 vdd.n504 185
R1697 vdd.n503 vdd.n456 185
R1698 vdd.n499 vdd.n498 185
R1699 vdd.n497 vdd.n496 185
R1700 vdd.n495 vdd.n494 185
R1701 vdd.n493 vdd.n458 185
R1702 vdd.n489 vdd.n488 185
R1703 vdd.n487 vdd.n486 185
R1704 vdd.n485 vdd.n484 185
R1705 vdd.n483 vdd.n460 185
R1706 vdd.n479 vdd.n478 185
R1707 vdd.n477 vdd.n476 185
R1708 vdd.n475 vdd.n474 185
R1709 vdd.n473 vdd.n462 185
R1710 vdd.n469 vdd.n468 185
R1711 vdd.n467 vdd.n466 185
R1712 vdd.n465 vdd.n392 185
R1713 vdd.n3530 vdd.n393 185
R1714 vdd.n3537 vdd.n393 185
R1715 vdd.n3529 vdd.n3528 185
R1716 vdd.n3528 vdd.n386 185
R1717 vdd.n3527 vdd.n385 185
R1718 vdd.n3543 vdd.n385 185
R1719 vdd.n621 vdd.n384 185
R1720 vdd.n3544 vdd.n384 185
R1721 vdd.n3523 vdd.n383 185
R1722 vdd.n3545 vdd.n383 185
R1723 vdd.n3522 vdd.n3521 185
R1724 vdd.n3521 vdd.n375 185
R1725 vdd.n3520 vdd.n374 185
R1726 vdd.n3551 vdd.n374 185
R1727 vdd.n623 vdd.n373 185
R1728 vdd.n3552 vdd.n373 185
R1729 vdd.n3516 vdd.n372 185
R1730 vdd.n3553 vdd.n372 185
R1731 vdd.n3515 vdd.n3514 185
R1732 vdd.n3514 vdd.n3513 185
R1733 vdd.n3512 vdd.n364 185
R1734 vdd.n3559 vdd.n364 185
R1735 vdd.n625 vdd.n363 185
R1736 vdd.n3560 vdd.n363 185
R1737 vdd.n3508 vdd.n362 185
R1738 vdd.n3561 vdd.n362 185
R1739 vdd.n3507 vdd.n3506 185
R1740 vdd.n3506 vdd.n361 185
R1741 vdd.n3505 vdd.n353 185
R1742 vdd.n3567 vdd.n353 185
R1743 vdd.n627 vdd.n352 185
R1744 vdd.n3568 vdd.n352 185
R1745 vdd.n3501 vdd.n351 185
R1746 vdd.n3569 vdd.n351 185
R1747 vdd.n3500 vdd.n3499 185
R1748 vdd.n3499 vdd.n344 185
R1749 vdd.n3498 vdd.n343 185
R1750 vdd.n3575 vdd.n343 185
R1751 vdd.n629 vdd.n342 185
R1752 vdd.n3576 vdd.n342 185
R1753 vdd.n3494 vdd.n341 185
R1754 vdd.n3577 vdd.n341 185
R1755 vdd.n3493 vdd.n3492 185
R1756 vdd.n3492 vdd.n340 185
R1757 vdd.n3491 vdd.n631 185
R1758 vdd.n3491 vdd.n3490 185
R1759 vdd.n3479 vdd.n632 185
R1760 vdd.n633 vdd.n632 185
R1761 vdd.n3481 vdd.n3480 185
R1762 vdd.n3482 vdd.n3481 185
R1763 vdd.n640 vdd.n639 185
R1764 vdd.n644 vdd.n639 185
R1765 vdd.n3473 vdd.n3472 185
R1766 vdd.n3472 vdd.n3471 185
R1767 vdd.n643 vdd.n642 185
R1768 vdd.n3462 vdd.n643 185
R1769 vdd.n3461 vdd.n3460 185
R1770 vdd.n3463 vdd.n3461 185
R1771 vdd.n651 vdd.n650 185
R1772 vdd.n656 vdd.n650 185
R1773 vdd.n3456 vdd.n3455 185
R1774 vdd.n3455 vdd.n3454 185
R1775 vdd.n654 vdd.n653 185
R1776 vdd.n655 vdd.n654 185
R1777 vdd.n3445 vdd.n3444 185
R1778 vdd.n3446 vdd.n3445 185
R1779 vdd.n664 vdd.n663 185
R1780 vdd.n663 vdd.n662 185
R1781 vdd.n3440 vdd.n3439 185
R1782 vdd.n3439 vdd.n3438 185
R1783 vdd.n667 vdd.n666 185
R1784 vdd.n3429 vdd.n667 185
R1785 vdd.n3428 vdd.n3427 185
R1786 vdd.n3430 vdd.n3428 185
R1787 vdd.n674 vdd.n673 185
R1788 vdd.n679 vdd.n673 185
R1789 vdd.n3423 vdd.n3422 185
R1790 vdd.n3422 vdd.n3421 185
R1791 vdd.n677 vdd.n676 185
R1792 vdd.n678 vdd.n677 185
R1793 vdd.n3412 vdd.n3411 185
R1794 vdd.n3413 vdd.n3412 185
R1795 vdd.n686 vdd.n685 185
R1796 vdd.n723 vdd.n685 185
R1797 vdd.n3014 vdd.n947 185
R1798 vdd.n3013 vdd.n3012 185
R1799 vdd.n949 vdd.n948 185
R1800 vdd.n3010 vdd.n949 185
R1801 vdd.n2833 vdd.n2832 185
R1802 vdd.n2835 vdd.n2834 185
R1803 vdd.n2837 vdd.n2836 185
R1804 vdd.n2839 vdd.n2838 185
R1805 vdd.n2841 vdd.n2840 185
R1806 vdd.n2843 vdd.n2842 185
R1807 vdd.n2845 vdd.n2844 185
R1808 vdd.n2847 vdd.n2846 185
R1809 vdd.n2849 vdd.n2848 185
R1810 vdd.n2851 vdd.n2850 185
R1811 vdd.n2853 vdd.n2852 185
R1812 vdd.n2855 vdd.n2854 185
R1813 vdd.n2857 vdd.n2856 185
R1814 vdd.n2859 vdd.n2858 185
R1815 vdd.n2861 vdd.n2860 185
R1816 vdd.n2863 vdd.n2862 185
R1817 vdd.n2865 vdd.n2864 185
R1818 vdd.n2867 vdd.n2866 185
R1819 vdd.n2869 vdd.n2868 185
R1820 vdd.n2871 vdd.n2870 185
R1821 vdd.n2873 vdd.n2872 185
R1822 vdd.n2875 vdd.n2874 185
R1823 vdd.n2877 vdd.n2876 185
R1824 vdd.n2879 vdd.n2878 185
R1825 vdd.n2881 vdd.n2880 185
R1826 vdd.n2883 vdd.n2882 185
R1827 vdd.n2885 vdd.n2884 185
R1828 vdd.n2887 vdd.n2886 185
R1829 vdd.n2889 vdd.n2888 185
R1830 vdd.n2892 vdd.n2891 185
R1831 vdd.n2894 vdd.n2893 185
R1832 vdd.n2896 vdd.n2895 185
R1833 vdd.n3177 vdd.n3176 185
R1834 vdd.n3179 vdd.n834 185
R1835 vdd.n3181 vdd.n3180 185
R1836 vdd.n3183 vdd.n831 185
R1837 vdd.n3185 vdd.n3184 185
R1838 vdd.n3187 vdd.n829 185
R1839 vdd.n3189 vdd.n3188 185
R1840 vdd.n3190 vdd.n828 185
R1841 vdd.n3192 vdd.n3191 185
R1842 vdd.n3194 vdd.n826 185
R1843 vdd.n3196 vdd.n3195 185
R1844 vdd.n3197 vdd.n825 185
R1845 vdd.n3199 vdd.n3198 185
R1846 vdd.n3201 vdd.n823 185
R1847 vdd.n3203 vdd.n3202 185
R1848 vdd.n3204 vdd.n822 185
R1849 vdd.n3206 vdd.n3205 185
R1850 vdd.n3208 vdd.n731 185
R1851 vdd.n3210 vdd.n3209 185
R1852 vdd.n3212 vdd.n820 185
R1853 vdd.n3214 vdd.n3213 185
R1854 vdd.n3215 vdd.n819 185
R1855 vdd.n3217 vdd.n3216 185
R1856 vdd.n3219 vdd.n817 185
R1857 vdd.n3221 vdd.n3220 185
R1858 vdd.n3222 vdd.n816 185
R1859 vdd.n3224 vdd.n3223 185
R1860 vdd.n3226 vdd.n814 185
R1861 vdd.n3228 vdd.n3227 185
R1862 vdd.n3229 vdd.n813 185
R1863 vdd.n3231 vdd.n3230 185
R1864 vdd.n3233 vdd.n812 185
R1865 vdd.n3234 vdd.n811 185
R1866 vdd.n3237 vdd.n3236 185
R1867 vdd.n3238 vdd.n809 185
R1868 vdd.n809 vdd.n692 185
R1869 vdd.n3175 vdd.n806 185
R1870 vdd.n3241 vdd.n806 185
R1871 vdd.n3174 vdd.n3173 185
R1872 vdd.n3173 vdd.n805 185
R1873 vdd.n3172 vdd.n836 185
R1874 vdd.n3172 vdd.n3171 185
R1875 vdd.n2946 vdd.n837 185
R1876 vdd.n846 vdd.n837 185
R1877 vdd.n2947 vdd.n844 185
R1878 vdd.n3165 vdd.n844 185
R1879 vdd.n2949 vdd.n2948 185
R1880 vdd.n2948 vdd.n843 185
R1881 vdd.n2950 vdd.n852 185
R1882 vdd.n3114 vdd.n852 185
R1883 vdd.n2952 vdd.n2951 185
R1884 vdd.n2951 vdd.n851 185
R1885 vdd.n2953 vdd.n857 185
R1886 vdd.n3108 vdd.n857 185
R1887 vdd.n2955 vdd.n2954 185
R1888 vdd.n2954 vdd.n864 185
R1889 vdd.n2956 vdd.n862 185
R1890 vdd.n3102 vdd.n862 185
R1891 vdd.n2958 vdd.n2957 185
R1892 vdd.n2957 vdd.n870 185
R1893 vdd.n2959 vdd.n868 185
R1894 vdd.n3096 vdd.n868 185
R1895 vdd.n2961 vdd.n2960 185
R1896 vdd.n2960 vdd.n877 185
R1897 vdd.n2962 vdd.n875 185
R1898 vdd.n3090 vdd.n875 185
R1899 vdd.n2964 vdd.n2963 185
R1900 vdd.n2963 vdd.n874 185
R1901 vdd.n2965 vdd.n882 185
R1902 vdd.n3084 vdd.n882 185
R1903 vdd.n2967 vdd.n2966 185
R1904 vdd.n2966 vdd.n881 185
R1905 vdd.n2968 vdd.n889 185
R1906 vdd.n3077 vdd.n889 185
R1907 vdd.n2970 vdd.n2969 185
R1908 vdd.n2969 vdd.n888 185
R1909 vdd.n2971 vdd.n894 185
R1910 vdd.n3071 vdd.n894 185
R1911 vdd.n2973 vdd.n2972 185
R1912 vdd.n2972 vdd.n901 185
R1913 vdd.n2974 vdd.n899 185
R1914 vdd.n3065 vdd.n899 185
R1915 vdd.n2976 vdd.n2975 185
R1916 vdd.n2977 vdd.n2976 185
R1917 vdd.n2945 vdd.n906 185
R1918 vdd.n3059 vdd.n906 185
R1919 vdd.n2944 vdd.n2943 185
R1920 vdd.n2943 vdd.n905 185
R1921 vdd.n2942 vdd.n912 185
R1922 vdd.n3053 vdd.n912 185
R1923 vdd.n2941 vdd.n2940 185
R1924 vdd.n2940 vdd.n911 185
R1925 vdd.n2901 vdd.n917 185
R1926 vdd.n3047 vdd.n917 185
R1927 vdd.n2991 vdd.n2990 185
R1928 vdd.n2990 vdd.n2989 185
R1929 vdd.n2992 vdd.n922 185
R1930 vdd.n3041 vdd.n922 185
R1931 vdd.n2994 vdd.n2993 185
R1932 vdd.n2993 vdd.n930 185
R1933 vdd.n2995 vdd.n928 185
R1934 vdd.n3035 vdd.n928 185
R1935 vdd.n2997 vdd.n2996 185
R1936 vdd.n2996 vdd.n927 185
R1937 vdd.n2998 vdd.n934 185
R1938 vdd.n3029 vdd.n934 185
R1939 vdd.n3000 vdd.n2999 185
R1940 vdd.n3001 vdd.n3000 185
R1941 vdd.n2900 vdd.n939 185
R1942 vdd.n3023 vdd.n939 185
R1943 vdd.n2899 vdd.n2898 185
R1944 vdd.n2898 vdd.n946 185
R1945 vdd.n2897 vdd.n944 185
R1946 vdd.n3017 vdd.n944 185
R1947 vdd.n3016 vdd.n3015 185
R1948 vdd.n3017 vdd.n3016 185
R1949 vdd.n938 vdd.n937 185
R1950 vdd.n946 vdd.n938 185
R1951 vdd.n3025 vdd.n3024 185
R1952 vdd.n3024 vdd.n3023 185
R1953 vdd.n3026 vdd.n936 185
R1954 vdd.n3001 vdd.n936 185
R1955 vdd.n3028 vdd.n3027 185
R1956 vdd.n3029 vdd.n3028 185
R1957 vdd.n926 vdd.n925 185
R1958 vdd.n927 vdd.n926 185
R1959 vdd.n3037 vdd.n3036 185
R1960 vdd.n3036 vdd.n3035 185
R1961 vdd.n3038 vdd.n924 185
R1962 vdd.n930 vdd.n924 185
R1963 vdd.n3040 vdd.n3039 185
R1964 vdd.n3041 vdd.n3040 185
R1965 vdd.n916 vdd.n915 185
R1966 vdd.n2989 vdd.n916 185
R1967 vdd.n3049 vdd.n3048 185
R1968 vdd.n3048 vdd.n3047 185
R1969 vdd.n3050 vdd.n914 185
R1970 vdd.n914 vdd.n911 185
R1971 vdd.n3052 vdd.n3051 185
R1972 vdd.n3053 vdd.n3052 185
R1973 vdd.n904 vdd.n903 185
R1974 vdd.n905 vdd.n904 185
R1975 vdd.n3061 vdd.n3060 185
R1976 vdd.n3060 vdd.n3059 185
R1977 vdd.n3062 vdd.n902 185
R1978 vdd.n2977 vdd.n902 185
R1979 vdd.n3064 vdd.n3063 185
R1980 vdd.n3065 vdd.n3064 185
R1981 vdd.n893 vdd.n892 185
R1982 vdd.n901 vdd.n893 185
R1983 vdd.n3073 vdd.n3072 185
R1984 vdd.n3072 vdd.n3071 185
R1985 vdd.n3074 vdd.n891 185
R1986 vdd.n891 vdd.n888 185
R1987 vdd.n3076 vdd.n3075 185
R1988 vdd.n3077 vdd.n3076 185
R1989 vdd.n880 vdd.n879 185
R1990 vdd.n881 vdd.n880 185
R1991 vdd.n3086 vdd.n3085 185
R1992 vdd.n3085 vdd.n3084 185
R1993 vdd.n3087 vdd.n878 185
R1994 vdd.n878 vdd.n874 185
R1995 vdd.n3089 vdd.n3088 185
R1996 vdd.n3090 vdd.n3089 185
R1997 vdd.n867 vdd.n866 185
R1998 vdd.n877 vdd.n867 185
R1999 vdd.n3098 vdd.n3097 185
R2000 vdd.n3097 vdd.n3096 185
R2001 vdd.n3099 vdd.n865 185
R2002 vdd.n870 vdd.n865 185
R2003 vdd.n3101 vdd.n3100 185
R2004 vdd.n3102 vdd.n3101 185
R2005 vdd.n856 vdd.n855 185
R2006 vdd.n864 vdd.n856 185
R2007 vdd.n3110 vdd.n3109 185
R2008 vdd.n3109 vdd.n3108 185
R2009 vdd.n3111 vdd.n854 185
R2010 vdd.n854 vdd.n851 185
R2011 vdd.n3113 vdd.n3112 185
R2012 vdd.n3114 vdd.n3113 185
R2013 vdd.n842 vdd.n841 185
R2014 vdd.n843 vdd.n842 185
R2015 vdd.n3167 vdd.n3166 185
R2016 vdd.n3166 vdd.n3165 185
R2017 vdd.n3168 vdd.n840 185
R2018 vdd.n846 vdd.n840 185
R2019 vdd.n3170 vdd.n3169 185
R2020 vdd.n3171 vdd.n3170 185
R2021 vdd.n810 vdd.n808 185
R2022 vdd.n808 vdd.n805 185
R2023 vdd.n3240 vdd.n3239 185
R2024 vdd.n3241 vdd.n3240 185
R2025 vdd.n2653 vdd.n2652 185
R2026 vdd.n2654 vdd.n2653 185
R2027 vdd.n996 vdd.n994 185
R2028 vdd.n994 vdd.n992 185
R2029 vdd.n2568 vdd.n1003 185
R2030 vdd.n2579 vdd.n1003 185
R2031 vdd.n2569 vdd.n1012 185
R2032 vdd.n2334 vdd.n1012 185
R2033 vdd.n2571 vdd.n2570 185
R2034 vdd.n2572 vdd.n2571 185
R2035 vdd.n2567 vdd.n1011 185
R2036 vdd.n1011 vdd.n1008 185
R2037 vdd.n2566 vdd.n2565 185
R2038 vdd.n2565 vdd.n2564 185
R2039 vdd.n1014 vdd.n1013 185
R2040 vdd.n1015 vdd.n1014 185
R2041 vdd.n2557 vdd.n2556 185
R2042 vdd.n2558 vdd.n2557 185
R2043 vdd.n2555 vdd.n1023 185
R2044 vdd.n2346 vdd.n1023 185
R2045 vdd.n2554 vdd.n2553 185
R2046 vdd.n2553 vdd.n2552 185
R2047 vdd.n1025 vdd.n1024 185
R2048 vdd.n1033 vdd.n1025 185
R2049 vdd.n2545 vdd.n2544 185
R2050 vdd.n2546 vdd.n2545 185
R2051 vdd.n2543 vdd.n1034 185
R2052 vdd.n1039 vdd.n1034 185
R2053 vdd.n2542 vdd.n2541 185
R2054 vdd.n2541 vdd.n2540 185
R2055 vdd.n1036 vdd.n1035 185
R2056 vdd.n2358 vdd.n1036 185
R2057 vdd.n2533 vdd.n2532 185
R2058 vdd.n2534 vdd.n2533 185
R2059 vdd.n2531 vdd.n1046 185
R2060 vdd.n1046 vdd.n1043 185
R2061 vdd.n2530 vdd.n2529 185
R2062 vdd.n2529 vdd.n2528 185
R2063 vdd.n1048 vdd.n1047 185
R2064 vdd.n1049 vdd.n1048 185
R2065 vdd.n2521 vdd.n2520 185
R2066 vdd.n2522 vdd.n2521 185
R2067 vdd.n2518 vdd.n1057 185
R2068 vdd.n1063 vdd.n1057 185
R2069 vdd.n2517 vdd.n2516 185
R2070 vdd.n2516 vdd.n2515 185
R2071 vdd.n1060 vdd.n1059 185
R2072 vdd.n1070 vdd.n1060 185
R2073 vdd.n2508 vdd.n2507 185
R2074 vdd.n2509 vdd.n2508 185
R2075 vdd.n2506 vdd.n1071 185
R2076 vdd.n1071 vdd.n1067 185
R2077 vdd.n2505 vdd.n2504 185
R2078 vdd.n2504 vdd.n2503 185
R2079 vdd.n1073 vdd.n1072 185
R2080 vdd.n1074 vdd.n1073 185
R2081 vdd.n2496 vdd.n2495 185
R2082 vdd.n2497 vdd.n2496 185
R2083 vdd.n2494 vdd.n1083 185
R2084 vdd.n1083 vdd.n1080 185
R2085 vdd.n2493 vdd.n2492 185
R2086 vdd.n2492 vdd.n2491 185
R2087 vdd.n1085 vdd.n1084 185
R2088 vdd.n1086 vdd.n1085 185
R2089 vdd.n2484 vdd.n2483 185
R2090 vdd.n2485 vdd.n2484 185
R2091 vdd.n2482 vdd.n1095 185
R2092 vdd.n1095 vdd.n1092 185
R2093 vdd.n2481 vdd.n2480 185
R2094 vdd.n2480 vdd.n2479 185
R2095 vdd.n1097 vdd.n1096 185
R2096 vdd.n1098 vdd.n1097 185
R2097 vdd.n2472 vdd.n2471 185
R2098 vdd.n2473 vdd.n2472 185
R2099 vdd.n2470 vdd.n1107 185
R2100 vdd.n1107 vdd.n1104 185
R2101 vdd.n2469 vdd.n2468 185
R2102 vdd.n2468 vdd.n2467 185
R2103 vdd.n2584 vdd.n967 185
R2104 vdd.n2726 vdd.n967 185
R2105 vdd.n2586 vdd.n2585 185
R2106 vdd.n2588 vdd.n2587 185
R2107 vdd.n2590 vdd.n2589 185
R2108 vdd.n2592 vdd.n2591 185
R2109 vdd.n2594 vdd.n2593 185
R2110 vdd.n2596 vdd.n2595 185
R2111 vdd.n2598 vdd.n2597 185
R2112 vdd.n2600 vdd.n2599 185
R2113 vdd.n2602 vdd.n2601 185
R2114 vdd.n2604 vdd.n2603 185
R2115 vdd.n2606 vdd.n2605 185
R2116 vdd.n2608 vdd.n2607 185
R2117 vdd.n2610 vdd.n2609 185
R2118 vdd.n2612 vdd.n2611 185
R2119 vdd.n2614 vdd.n2613 185
R2120 vdd.n2616 vdd.n2615 185
R2121 vdd.n2618 vdd.n2617 185
R2122 vdd.n2620 vdd.n2619 185
R2123 vdd.n2622 vdd.n2621 185
R2124 vdd.n2624 vdd.n2623 185
R2125 vdd.n2626 vdd.n2625 185
R2126 vdd.n2628 vdd.n2627 185
R2127 vdd.n2630 vdd.n2629 185
R2128 vdd.n2632 vdd.n2631 185
R2129 vdd.n2634 vdd.n2633 185
R2130 vdd.n2636 vdd.n2635 185
R2131 vdd.n2638 vdd.n2637 185
R2132 vdd.n2640 vdd.n2639 185
R2133 vdd.n2642 vdd.n2641 185
R2134 vdd.n2644 vdd.n2643 185
R2135 vdd.n2646 vdd.n2645 185
R2136 vdd.n2648 vdd.n2647 185
R2137 vdd.n2650 vdd.n2649 185
R2138 vdd.n2651 vdd.n995 185
R2139 vdd.n2583 vdd.n993 185
R2140 vdd.n2654 vdd.n993 185
R2141 vdd.n2582 vdd.n2581 185
R2142 vdd.n2581 vdd.n992 185
R2143 vdd.n2580 vdd.n1000 185
R2144 vdd.n2580 vdd.n2579 185
R2145 vdd.n2318 vdd.n1001 185
R2146 vdd.n2334 vdd.n1001 185
R2147 vdd.n2319 vdd.n1010 185
R2148 vdd.n2572 vdd.n1010 185
R2149 vdd.n2321 vdd.n2320 185
R2150 vdd.n2320 vdd.n1008 185
R2151 vdd.n2322 vdd.n1017 185
R2152 vdd.n2564 vdd.n1017 185
R2153 vdd.n2324 vdd.n2323 185
R2154 vdd.n2323 vdd.n1015 185
R2155 vdd.n2325 vdd.n1022 185
R2156 vdd.n2558 vdd.n1022 185
R2157 vdd.n2348 vdd.n2347 185
R2158 vdd.n2347 vdd.n2346 185
R2159 vdd.n2349 vdd.n1027 185
R2160 vdd.n2552 vdd.n1027 185
R2161 vdd.n2351 vdd.n2350 185
R2162 vdd.n2350 vdd.n1033 185
R2163 vdd.n2352 vdd.n1032 185
R2164 vdd.n2546 vdd.n1032 185
R2165 vdd.n2354 vdd.n2353 185
R2166 vdd.n2353 vdd.n1039 185
R2167 vdd.n2355 vdd.n1038 185
R2168 vdd.n2540 vdd.n1038 185
R2169 vdd.n2357 vdd.n2356 185
R2170 vdd.n2358 vdd.n2357 185
R2171 vdd.n2317 vdd.n1045 185
R2172 vdd.n2534 vdd.n1045 185
R2173 vdd.n2316 vdd.n2315 185
R2174 vdd.n2315 vdd.n1043 185
R2175 vdd.n2314 vdd.n1051 185
R2176 vdd.n2528 vdd.n1051 185
R2177 vdd.n2313 vdd.n2312 185
R2178 vdd.n2312 vdd.n1049 185
R2179 vdd.n2311 vdd.n1056 185
R2180 vdd.n2522 vdd.n1056 185
R2181 vdd.n2310 vdd.n2309 185
R2182 vdd.n2309 vdd.n1063 185
R2183 vdd.n2308 vdd.n1062 185
R2184 vdd.n2515 vdd.n1062 185
R2185 vdd.n2307 vdd.n2306 185
R2186 vdd.n2306 vdd.n1070 185
R2187 vdd.n2305 vdd.n1069 185
R2188 vdd.n2509 vdd.n1069 185
R2189 vdd.n2304 vdd.n2303 185
R2190 vdd.n2303 vdd.n1067 185
R2191 vdd.n2302 vdd.n1076 185
R2192 vdd.n2503 vdd.n1076 185
R2193 vdd.n2301 vdd.n2300 185
R2194 vdd.n2300 vdd.n1074 185
R2195 vdd.n2299 vdd.n1082 185
R2196 vdd.n2497 vdd.n1082 185
R2197 vdd.n2298 vdd.n2297 185
R2198 vdd.n2297 vdd.n1080 185
R2199 vdd.n2296 vdd.n1088 185
R2200 vdd.n2491 vdd.n1088 185
R2201 vdd.n2295 vdd.n2294 185
R2202 vdd.n2294 vdd.n1086 185
R2203 vdd.n2293 vdd.n1094 185
R2204 vdd.n2485 vdd.n1094 185
R2205 vdd.n2292 vdd.n2291 185
R2206 vdd.n2291 vdd.n1092 185
R2207 vdd.n2290 vdd.n1100 185
R2208 vdd.n2479 vdd.n1100 185
R2209 vdd.n2289 vdd.n2288 185
R2210 vdd.n2288 vdd.n1098 185
R2211 vdd.n2287 vdd.n1106 185
R2212 vdd.n2473 vdd.n1106 185
R2213 vdd.n2286 vdd.n2285 185
R2214 vdd.n2285 vdd.n1104 185
R2215 vdd.n2284 vdd.n1112 185
R2216 vdd.n2467 vdd.n1112 185
R2217 vdd.n1109 vdd.n1108 185
R2218 vdd.n2216 vdd.n2214 185
R2219 vdd.n2219 vdd.n2218 185
R2220 vdd.n2220 vdd.n2213 185
R2221 vdd.n2222 vdd.n2221 185
R2222 vdd.n2224 vdd.n2212 185
R2223 vdd.n2227 vdd.n2226 185
R2224 vdd.n2228 vdd.n2211 185
R2225 vdd.n2230 vdd.n2229 185
R2226 vdd.n2232 vdd.n2210 185
R2227 vdd.n2235 vdd.n2234 185
R2228 vdd.n2236 vdd.n2209 185
R2229 vdd.n2238 vdd.n2237 185
R2230 vdd.n2240 vdd.n2208 185
R2231 vdd.n2243 vdd.n2242 185
R2232 vdd.n2244 vdd.n2207 185
R2233 vdd.n2246 vdd.n2245 185
R2234 vdd.n2248 vdd.n2206 185
R2235 vdd.n2251 vdd.n2250 185
R2236 vdd.n2252 vdd.n1143 185
R2237 vdd.n2254 vdd.n2253 185
R2238 vdd.n2256 vdd.n1142 185
R2239 vdd.n2259 vdd.n2258 185
R2240 vdd.n2260 vdd.n1141 185
R2241 vdd.n2262 vdd.n2261 185
R2242 vdd.n2264 vdd.n1140 185
R2243 vdd.n2267 vdd.n2266 185
R2244 vdd.n2268 vdd.n1139 185
R2245 vdd.n2270 vdd.n2269 185
R2246 vdd.n2272 vdd.n1138 185
R2247 vdd.n2275 vdd.n2274 185
R2248 vdd.n2276 vdd.n1135 185
R2249 vdd.n2279 vdd.n2278 185
R2250 vdd.n2281 vdd.n1134 185
R2251 vdd.n2283 vdd.n2282 185
R2252 vdd.n2282 vdd.n1110 185
R2253 vdd.n327 vdd.n326 171.744
R2254 vdd.n326 vdd.n325 171.744
R2255 vdd.n325 vdd.n294 171.744
R2256 vdd.n318 vdd.n294 171.744
R2257 vdd.n318 vdd.n317 171.744
R2258 vdd.n317 vdd.n299 171.744
R2259 vdd.n310 vdd.n299 171.744
R2260 vdd.n310 vdd.n309 171.744
R2261 vdd.n309 vdd.n303 171.744
R2262 vdd.n268 vdd.n267 171.744
R2263 vdd.n267 vdd.n266 171.744
R2264 vdd.n266 vdd.n235 171.744
R2265 vdd.n259 vdd.n235 171.744
R2266 vdd.n259 vdd.n258 171.744
R2267 vdd.n258 vdd.n240 171.744
R2268 vdd.n251 vdd.n240 171.744
R2269 vdd.n251 vdd.n250 171.744
R2270 vdd.n250 vdd.n244 171.744
R2271 vdd.n225 vdd.n224 171.744
R2272 vdd.n224 vdd.n223 171.744
R2273 vdd.n223 vdd.n192 171.744
R2274 vdd.n216 vdd.n192 171.744
R2275 vdd.n216 vdd.n215 171.744
R2276 vdd.n215 vdd.n197 171.744
R2277 vdd.n208 vdd.n197 171.744
R2278 vdd.n208 vdd.n207 171.744
R2279 vdd.n207 vdd.n201 171.744
R2280 vdd.n166 vdd.n165 171.744
R2281 vdd.n165 vdd.n164 171.744
R2282 vdd.n164 vdd.n133 171.744
R2283 vdd.n157 vdd.n133 171.744
R2284 vdd.n157 vdd.n156 171.744
R2285 vdd.n156 vdd.n138 171.744
R2286 vdd.n149 vdd.n138 171.744
R2287 vdd.n149 vdd.n148 171.744
R2288 vdd.n148 vdd.n142 171.744
R2289 vdd.n124 vdd.n123 171.744
R2290 vdd.n123 vdd.n122 171.744
R2291 vdd.n122 vdd.n91 171.744
R2292 vdd.n115 vdd.n91 171.744
R2293 vdd.n115 vdd.n114 171.744
R2294 vdd.n114 vdd.n96 171.744
R2295 vdd.n107 vdd.n96 171.744
R2296 vdd.n107 vdd.n106 171.744
R2297 vdd.n106 vdd.n100 171.744
R2298 vdd.n65 vdd.n64 171.744
R2299 vdd.n64 vdd.n63 171.744
R2300 vdd.n63 vdd.n32 171.744
R2301 vdd.n56 vdd.n32 171.744
R2302 vdd.n56 vdd.n55 171.744
R2303 vdd.n55 vdd.n37 171.744
R2304 vdd.n48 vdd.n37 171.744
R2305 vdd.n48 vdd.n47 171.744
R2306 vdd.n47 vdd.n41 171.744
R2307 vdd.n1826 vdd.n1825 171.744
R2308 vdd.n1825 vdd.n1824 171.744
R2309 vdd.n1824 vdd.n1793 171.744
R2310 vdd.n1817 vdd.n1793 171.744
R2311 vdd.n1817 vdd.n1816 171.744
R2312 vdd.n1816 vdd.n1798 171.744
R2313 vdd.n1809 vdd.n1798 171.744
R2314 vdd.n1809 vdd.n1808 171.744
R2315 vdd.n1808 vdd.n1802 171.744
R2316 vdd.n1885 vdd.n1884 171.744
R2317 vdd.n1884 vdd.n1883 171.744
R2318 vdd.n1883 vdd.n1852 171.744
R2319 vdd.n1876 vdd.n1852 171.744
R2320 vdd.n1876 vdd.n1875 171.744
R2321 vdd.n1875 vdd.n1857 171.744
R2322 vdd.n1868 vdd.n1857 171.744
R2323 vdd.n1868 vdd.n1867 171.744
R2324 vdd.n1867 vdd.n1861 171.744
R2325 vdd.n1724 vdd.n1723 171.744
R2326 vdd.n1723 vdd.n1722 171.744
R2327 vdd.n1722 vdd.n1691 171.744
R2328 vdd.n1715 vdd.n1691 171.744
R2329 vdd.n1715 vdd.n1714 171.744
R2330 vdd.n1714 vdd.n1696 171.744
R2331 vdd.n1707 vdd.n1696 171.744
R2332 vdd.n1707 vdd.n1706 171.744
R2333 vdd.n1706 vdd.n1700 171.744
R2334 vdd.n1783 vdd.n1782 171.744
R2335 vdd.n1782 vdd.n1781 171.744
R2336 vdd.n1781 vdd.n1750 171.744
R2337 vdd.n1774 vdd.n1750 171.744
R2338 vdd.n1774 vdd.n1773 171.744
R2339 vdd.n1773 vdd.n1755 171.744
R2340 vdd.n1766 vdd.n1755 171.744
R2341 vdd.n1766 vdd.n1765 171.744
R2342 vdd.n1765 vdd.n1759 171.744
R2343 vdd.n1623 vdd.n1622 171.744
R2344 vdd.n1622 vdd.n1621 171.744
R2345 vdd.n1621 vdd.n1590 171.744
R2346 vdd.n1614 vdd.n1590 171.744
R2347 vdd.n1614 vdd.n1613 171.744
R2348 vdd.n1613 vdd.n1595 171.744
R2349 vdd.n1606 vdd.n1595 171.744
R2350 vdd.n1606 vdd.n1605 171.744
R2351 vdd.n1605 vdd.n1599 171.744
R2352 vdd.n1682 vdd.n1681 171.744
R2353 vdd.n1681 vdd.n1680 171.744
R2354 vdd.n1680 vdd.n1649 171.744
R2355 vdd.n1673 vdd.n1649 171.744
R2356 vdd.n1673 vdd.n1672 171.744
R2357 vdd.n1672 vdd.n1654 171.744
R2358 vdd.n1665 vdd.n1654 171.744
R2359 vdd.n1665 vdd.n1664 171.744
R2360 vdd.n1664 vdd.n1658 171.744
R2361 vdd.n468 vdd.n467 146.341
R2362 vdd.n474 vdd.n473 146.341
R2363 vdd.n478 vdd.n477 146.341
R2364 vdd.n484 vdd.n483 146.341
R2365 vdd.n488 vdd.n487 146.341
R2366 vdd.n494 vdd.n493 146.341
R2367 vdd.n498 vdd.n497 146.341
R2368 vdd.n504 vdd.n503 146.341
R2369 vdd.n508 vdd.n507 146.341
R2370 vdd.n514 vdd.n513 146.341
R2371 vdd.n518 vdd.n517 146.341
R2372 vdd.n524 vdd.n523 146.341
R2373 vdd.n528 vdd.n527 146.341
R2374 vdd.n534 vdd.n533 146.341
R2375 vdd.n538 vdd.n537 146.341
R2376 vdd.n544 vdd.n543 146.341
R2377 vdd.n548 vdd.n547 146.341
R2378 vdd.n554 vdd.n553 146.341
R2379 vdd.n558 vdd.n557 146.341
R2380 vdd.n564 vdd.n563 146.341
R2381 vdd.n568 vdd.n567 146.341
R2382 vdd.n574 vdd.n573 146.341
R2383 vdd.n578 vdd.n577 146.341
R2384 vdd.n584 vdd.n583 146.341
R2385 vdd.n588 vdd.n587 146.341
R2386 vdd.n594 vdd.n593 146.341
R2387 vdd.n598 vdd.n597 146.341
R2388 vdd.n604 vdd.n603 146.341
R2389 vdd.n608 vdd.n607 146.341
R2390 vdd.n614 vdd.n613 146.341
R2391 vdd.n616 vdd.n425 146.341
R2392 vdd.n3412 vdd.n685 146.341
R2393 vdd.n3412 vdd.n677 146.341
R2394 vdd.n3422 vdd.n677 146.341
R2395 vdd.n3422 vdd.n673 146.341
R2396 vdd.n3428 vdd.n673 146.341
R2397 vdd.n3428 vdd.n667 146.341
R2398 vdd.n3439 vdd.n667 146.341
R2399 vdd.n3439 vdd.n663 146.341
R2400 vdd.n3445 vdd.n663 146.341
R2401 vdd.n3445 vdd.n654 146.341
R2402 vdd.n3455 vdd.n654 146.341
R2403 vdd.n3455 vdd.n650 146.341
R2404 vdd.n3461 vdd.n650 146.341
R2405 vdd.n3461 vdd.n643 146.341
R2406 vdd.n3472 vdd.n643 146.341
R2407 vdd.n3472 vdd.n639 146.341
R2408 vdd.n3481 vdd.n639 146.341
R2409 vdd.n3481 vdd.n632 146.341
R2410 vdd.n3491 vdd.n632 146.341
R2411 vdd.n3492 vdd.n3491 146.341
R2412 vdd.n3492 vdd.n341 146.341
R2413 vdd.n342 vdd.n341 146.341
R2414 vdd.n343 vdd.n342 146.341
R2415 vdd.n3499 vdd.n343 146.341
R2416 vdd.n3499 vdd.n351 146.341
R2417 vdd.n352 vdd.n351 146.341
R2418 vdd.n353 vdd.n352 146.341
R2419 vdd.n3506 vdd.n353 146.341
R2420 vdd.n3506 vdd.n362 146.341
R2421 vdd.n363 vdd.n362 146.341
R2422 vdd.n364 vdd.n363 146.341
R2423 vdd.n3514 vdd.n364 146.341
R2424 vdd.n3514 vdd.n372 146.341
R2425 vdd.n373 vdd.n372 146.341
R2426 vdd.n374 vdd.n373 146.341
R2427 vdd.n3521 vdd.n374 146.341
R2428 vdd.n3521 vdd.n383 146.341
R2429 vdd.n384 vdd.n383 146.341
R2430 vdd.n385 vdd.n384 146.341
R2431 vdd.n3528 vdd.n385 146.341
R2432 vdd.n3528 vdd.n393 146.341
R2433 vdd.n725 vdd.n724 146.341
R2434 vdd.n728 vdd.n724 146.341
R2435 vdd.n734 vdd.n733 146.341
R2436 vdd.n3394 vdd.n3393 146.341
R2437 vdd.n3390 vdd.n3389 146.341
R2438 vdd.n3386 vdd.n3385 146.341
R2439 vdd.n3382 vdd.n3381 146.341
R2440 vdd.n3378 vdd.n3377 146.341
R2441 vdd.n3374 vdd.n3373 146.341
R2442 vdd.n3370 vdd.n3369 146.341
R2443 vdd.n3361 vdd.n3360 146.341
R2444 vdd.n3358 vdd.n3357 146.341
R2445 vdd.n3354 vdd.n3353 146.341
R2446 vdd.n3350 vdd.n3349 146.341
R2447 vdd.n3346 vdd.n3345 146.341
R2448 vdd.n3342 vdd.n3341 146.341
R2449 vdd.n3338 vdd.n3337 146.341
R2450 vdd.n3334 vdd.n3333 146.341
R2451 vdd.n3330 vdd.n3329 146.341
R2452 vdd.n3326 vdd.n3325 146.341
R2453 vdd.n3322 vdd.n3321 146.341
R2454 vdd.n3315 vdd.n3314 146.341
R2455 vdd.n3312 vdd.n3311 146.341
R2456 vdd.n3308 vdd.n3307 146.341
R2457 vdd.n3304 vdd.n3303 146.341
R2458 vdd.n3300 vdd.n3299 146.341
R2459 vdd.n3296 vdd.n3295 146.341
R2460 vdd.n3292 vdd.n3291 146.341
R2461 vdd.n3288 vdd.n3287 146.341
R2462 vdd.n3284 vdd.n3283 146.341
R2463 vdd.n3280 vdd.n3279 146.341
R2464 vdd.n3406 vdd.n691 146.341
R2465 vdd.n3414 vdd.n684 146.341
R2466 vdd.n3414 vdd.n680 146.341
R2467 vdd.n3420 vdd.n680 146.341
R2468 vdd.n3420 vdd.n672 146.341
R2469 vdd.n3431 vdd.n672 146.341
R2470 vdd.n3431 vdd.n668 146.341
R2471 vdd.n3437 vdd.n668 146.341
R2472 vdd.n3437 vdd.n661 146.341
R2473 vdd.n3447 vdd.n661 146.341
R2474 vdd.n3447 vdd.n657 146.341
R2475 vdd.n3453 vdd.n657 146.341
R2476 vdd.n3453 vdd.n649 146.341
R2477 vdd.n3464 vdd.n649 146.341
R2478 vdd.n3464 vdd.n645 146.341
R2479 vdd.n3470 vdd.n645 146.341
R2480 vdd.n3470 vdd.n638 146.341
R2481 vdd.n3483 vdd.n638 146.341
R2482 vdd.n3483 vdd.n634 146.341
R2483 vdd.n3489 vdd.n634 146.341
R2484 vdd.n3489 vdd.n338 146.341
R2485 vdd.n3578 vdd.n338 146.341
R2486 vdd.n3578 vdd.n339 146.341
R2487 vdd.n3574 vdd.n339 146.341
R2488 vdd.n3574 vdd.n345 146.341
R2489 vdd.n3570 vdd.n345 146.341
R2490 vdd.n3570 vdd.n350 146.341
R2491 vdd.n3566 vdd.n350 146.341
R2492 vdd.n3566 vdd.n354 146.341
R2493 vdd.n3562 vdd.n354 146.341
R2494 vdd.n3562 vdd.n360 146.341
R2495 vdd.n3558 vdd.n360 146.341
R2496 vdd.n3558 vdd.n365 146.341
R2497 vdd.n3554 vdd.n365 146.341
R2498 vdd.n3554 vdd.n371 146.341
R2499 vdd.n3550 vdd.n371 146.341
R2500 vdd.n3550 vdd.n376 146.341
R2501 vdd.n3546 vdd.n376 146.341
R2502 vdd.n3546 vdd.n382 146.341
R2503 vdd.n3542 vdd.n382 146.341
R2504 vdd.n3542 vdd.n387 146.341
R2505 vdd.n3538 vdd.n387 146.341
R2506 vdd.n2189 vdd.n2188 146.341
R2507 vdd.n2186 vdd.n1983 146.341
R2508 vdd.n2179 vdd.n1989 146.341
R2509 vdd.n2177 vdd.n2176 146.341
R2510 vdd.n2174 vdd.n1991 146.341
R2511 vdd.n2170 vdd.n2169 146.341
R2512 vdd.n2167 vdd.n1998 146.341
R2513 vdd.n2163 vdd.n2162 146.341
R2514 vdd.n2160 vdd.n2005 146.341
R2515 vdd.n2016 vdd.n2013 146.341
R2516 vdd.n2152 vdd.n2151 146.341
R2517 vdd.n2149 vdd.n2018 146.341
R2518 vdd.n2145 vdd.n2144 146.341
R2519 vdd.n2142 vdd.n2024 146.341
R2520 vdd.n2138 vdd.n2137 146.341
R2521 vdd.n2135 vdd.n2031 146.341
R2522 vdd.n2131 vdd.n2130 146.341
R2523 vdd.n2128 vdd.n2038 146.341
R2524 vdd.n2124 vdd.n2123 146.341
R2525 vdd.n2121 vdd.n2045 146.341
R2526 vdd.n2056 vdd.n2053 146.341
R2527 vdd.n2113 vdd.n2112 146.341
R2528 vdd.n2110 vdd.n2058 146.341
R2529 vdd.n2106 vdd.n2105 146.341
R2530 vdd.n2103 vdd.n2064 146.341
R2531 vdd.n2099 vdd.n2098 146.341
R2532 vdd.n2096 vdd.n2071 146.341
R2533 vdd.n2092 vdd.n2091 146.341
R2534 vdd.n2089 vdd.n2086 146.341
R2535 vdd.n2084 vdd.n2081 146.341
R2536 vdd.n2079 vdd.n1149 146.341
R2537 vdd.n1508 vdd.n1268 146.341
R2538 vdd.n1508 vdd.n1264 146.341
R2539 vdd.n1514 vdd.n1264 146.341
R2540 vdd.n1514 vdd.n1256 146.341
R2541 vdd.n1525 vdd.n1256 146.341
R2542 vdd.n1525 vdd.n1252 146.341
R2543 vdd.n1531 vdd.n1252 146.341
R2544 vdd.n1531 vdd.n1246 146.341
R2545 vdd.n1542 vdd.n1246 146.341
R2546 vdd.n1542 vdd.n1242 146.341
R2547 vdd.n1548 vdd.n1242 146.341
R2548 vdd.n1548 vdd.n1233 146.341
R2549 vdd.n1558 vdd.n1233 146.341
R2550 vdd.n1558 vdd.n1229 146.341
R2551 vdd.n1564 vdd.n1229 146.341
R2552 vdd.n1564 vdd.n1222 146.341
R2553 vdd.n1575 vdd.n1222 146.341
R2554 vdd.n1575 vdd.n1218 146.341
R2555 vdd.n1581 vdd.n1218 146.341
R2556 vdd.n1581 vdd.n1211 146.341
R2557 vdd.n1898 vdd.n1211 146.341
R2558 vdd.n1898 vdd.n1207 146.341
R2559 vdd.n1904 vdd.n1207 146.341
R2560 vdd.n1904 vdd.n1199 146.341
R2561 vdd.n1915 vdd.n1199 146.341
R2562 vdd.n1915 vdd.n1195 146.341
R2563 vdd.n1921 vdd.n1195 146.341
R2564 vdd.n1921 vdd.n1189 146.341
R2565 vdd.n1932 vdd.n1189 146.341
R2566 vdd.n1932 vdd.n1185 146.341
R2567 vdd.n1938 vdd.n1185 146.341
R2568 vdd.n1938 vdd.n1176 146.341
R2569 vdd.n1948 vdd.n1176 146.341
R2570 vdd.n1948 vdd.n1172 146.341
R2571 vdd.n1954 vdd.n1172 146.341
R2572 vdd.n1954 vdd.n1166 146.341
R2573 vdd.n1965 vdd.n1166 146.341
R2574 vdd.n1965 vdd.n1161 146.341
R2575 vdd.n1973 vdd.n1161 146.341
R2576 vdd.n1973 vdd.n1151 146.341
R2577 vdd.n2197 vdd.n1151 146.341
R2578 vdd.n1497 vdd.n1273 146.341
R2579 vdd.n1497 vdd.n1306 146.341
R2580 vdd.n1310 vdd.n1309 146.341
R2581 vdd.n1312 vdd.n1311 146.341
R2582 vdd.n1316 vdd.n1315 146.341
R2583 vdd.n1318 vdd.n1317 146.341
R2584 vdd.n1322 vdd.n1321 146.341
R2585 vdd.n1324 vdd.n1323 146.341
R2586 vdd.n1328 vdd.n1327 146.341
R2587 vdd.n1330 vdd.n1329 146.341
R2588 vdd.n1336 vdd.n1335 146.341
R2589 vdd.n1338 vdd.n1337 146.341
R2590 vdd.n1342 vdd.n1341 146.341
R2591 vdd.n1344 vdd.n1343 146.341
R2592 vdd.n1348 vdd.n1347 146.341
R2593 vdd.n1350 vdd.n1349 146.341
R2594 vdd.n1354 vdd.n1353 146.341
R2595 vdd.n1356 vdd.n1355 146.341
R2596 vdd.n1360 vdd.n1359 146.341
R2597 vdd.n1362 vdd.n1361 146.341
R2598 vdd.n1434 vdd.n1365 146.341
R2599 vdd.n1367 vdd.n1366 146.341
R2600 vdd.n1371 vdd.n1370 146.341
R2601 vdd.n1373 vdd.n1372 146.341
R2602 vdd.n1377 vdd.n1376 146.341
R2603 vdd.n1379 vdd.n1378 146.341
R2604 vdd.n1383 vdd.n1382 146.341
R2605 vdd.n1385 vdd.n1384 146.341
R2606 vdd.n1389 vdd.n1388 146.341
R2607 vdd.n1391 vdd.n1390 146.341
R2608 vdd.n1395 vdd.n1394 146.341
R2609 vdd.n1396 vdd.n1304 146.341
R2610 vdd.n1506 vdd.n1269 146.341
R2611 vdd.n1506 vdd.n1262 146.341
R2612 vdd.n1517 vdd.n1262 146.341
R2613 vdd.n1517 vdd.n1258 146.341
R2614 vdd.n1523 vdd.n1258 146.341
R2615 vdd.n1523 vdd.n1251 146.341
R2616 vdd.n1534 vdd.n1251 146.341
R2617 vdd.n1534 vdd.n1247 146.341
R2618 vdd.n1540 vdd.n1247 146.341
R2619 vdd.n1540 vdd.n1240 146.341
R2620 vdd.n1550 vdd.n1240 146.341
R2621 vdd.n1550 vdd.n1236 146.341
R2622 vdd.n1556 vdd.n1236 146.341
R2623 vdd.n1556 vdd.n1228 146.341
R2624 vdd.n1567 vdd.n1228 146.341
R2625 vdd.n1567 vdd.n1224 146.341
R2626 vdd.n1573 vdd.n1224 146.341
R2627 vdd.n1573 vdd.n1217 146.341
R2628 vdd.n1583 vdd.n1217 146.341
R2629 vdd.n1583 vdd.n1213 146.341
R2630 vdd.n1896 vdd.n1213 146.341
R2631 vdd.n1896 vdd.n1205 146.341
R2632 vdd.n1907 vdd.n1205 146.341
R2633 vdd.n1907 vdd.n1201 146.341
R2634 vdd.n1913 vdd.n1201 146.341
R2635 vdd.n1913 vdd.n1194 146.341
R2636 vdd.n1924 vdd.n1194 146.341
R2637 vdd.n1924 vdd.n1190 146.341
R2638 vdd.n1930 vdd.n1190 146.341
R2639 vdd.n1930 vdd.n1183 146.341
R2640 vdd.n1940 vdd.n1183 146.341
R2641 vdd.n1940 vdd.n1179 146.341
R2642 vdd.n1946 vdd.n1179 146.341
R2643 vdd.n1946 vdd.n1171 146.341
R2644 vdd.n1957 vdd.n1171 146.341
R2645 vdd.n1957 vdd.n1167 146.341
R2646 vdd.n1963 vdd.n1167 146.341
R2647 vdd.n1963 vdd.n1159 146.341
R2648 vdd.n1976 vdd.n1159 146.341
R2649 vdd.n1976 vdd.n1154 146.341
R2650 vdd.n2195 vdd.n1154 146.341
R2651 vdd.n1136 vdd.t74 127.284
R2652 vdd.n997 vdd.t111 127.284
R2653 vdd.n1130 vdd.t138 127.284
R2654 vdd.n988 vdd.t134 127.284
R2655 vdd.n885 vdd.t84 127.284
R2656 vdd.n885 vdd.t85 127.284
R2657 vdd.n2761 vdd.t129 127.284
R2658 vdd.n832 vdd.t97 127.284
R2659 vdd.n2830 vdd.t116 127.284
R2660 vdd.n799 vdd.t69 127.284
R2661 vdd.n1058 vdd.t125 127.284
R2662 vdd.n1058 vdd.t126 127.284
R2663 vdd.n22 vdd.n20 117.314
R2664 vdd.n17 vdd.n15 117.314
R2665 vdd.n27 vdd.n26 116.927
R2666 vdd.n24 vdd.n23 116.927
R2667 vdd.n22 vdd.n21 116.927
R2668 vdd.n17 vdd.n16 116.927
R2669 vdd.n19 vdd.n18 116.927
R2670 vdd.n27 vdd.n25 116.927
R2671 vdd.n1137 vdd.t73 111.188
R2672 vdd.n998 vdd.t112 111.188
R2673 vdd.n1131 vdd.t137 111.188
R2674 vdd.n989 vdd.t135 111.188
R2675 vdd.n2762 vdd.t128 111.188
R2676 vdd.n833 vdd.t98 111.188
R2677 vdd.n2831 vdd.t115 111.188
R2678 vdd.n800 vdd.t70 111.188
R2679 vdd.n3016 vdd.n938 99.5127
R2680 vdd.n3024 vdd.n938 99.5127
R2681 vdd.n3024 vdd.n936 99.5127
R2682 vdd.n3028 vdd.n936 99.5127
R2683 vdd.n3028 vdd.n926 99.5127
R2684 vdd.n3036 vdd.n926 99.5127
R2685 vdd.n3036 vdd.n924 99.5127
R2686 vdd.n3040 vdd.n924 99.5127
R2687 vdd.n3040 vdd.n916 99.5127
R2688 vdd.n3048 vdd.n916 99.5127
R2689 vdd.n3048 vdd.n914 99.5127
R2690 vdd.n3052 vdd.n914 99.5127
R2691 vdd.n3052 vdd.n904 99.5127
R2692 vdd.n3060 vdd.n904 99.5127
R2693 vdd.n3060 vdd.n902 99.5127
R2694 vdd.n3064 vdd.n902 99.5127
R2695 vdd.n3064 vdd.n893 99.5127
R2696 vdd.n3072 vdd.n893 99.5127
R2697 vdd.n3072 vdd.n891 99.5127
R2698 vdd.n3076 vdd.n891 99.5127
R2699 vdd.n3076 vdd.n880 99.5127
R2700 vdd.n3085 vdd.n880 99.5127
R2701 vdd.n3085 vdd.n878 99.5127
R2702 vdd.n3089 vdd.n878 99.5127
R2703 vdd.n3089 vdd.n867 99.5127
R2704 vdd.n3097 vdd.n867 99.5127
R2705 vdd.n3097 vdd.n865 99.5127
R2706 vdd.n3101 vdd.n865 99.5127
R2707 vdd.n3101 vdd.n856 99.5127
R2708 vdd.n3109 vdd.n856 99.5127
R2709 vdd.n3109 vdd.n854 99.5127
R2710 vdd.n3113 vdd.n854 99.5127
R2711 vdd.n3113 vdd.n842 99.5127
R2712 vdd.n3166 vdd.n842 99.5127
R2713 vdd.n3166 vdd.n840 99.5127
R2714 vdd.n3170 vdd.n840 99.5127
R2715 vdd.n3170 vdd.n808 99.5127
R2716 vdd.n3240 vdd.n808 99.5127
R2717 vdd.n3236 vdd.n809 99.5127
R2718 vdd.n3234 vdd.n3233 99.5127
R2719 vdd.n3231 vdd.n813 99.5127
R2720 vdd.n3227 vdd.n3226 99.5127
R2721 vdd.n3224 vdd.n816 99.5127
R2722 vdd.n3220 vdd.n3219 99.5127
R2723 vdd.n3217 vdd.n819 99.5127
R2724 vdd.n3213 vdd.n3212 99.5127
R2725 vdd.n3210 vdd.n3208 99.5127
R2726 vdd.n3206 vdd.n822 99.5127
R2727 vdd.n3202 vdd.n3201 99.5127
R2728 vdd.n3199 vdd.n825 99.5127
R2729 vdd.n3195 vdd.n3194 99.5127
R2730 vdd.n3192 vdd.n828 99.5127
R2731 vdd.n3188 vdd.n3187 99.5127
R2732 vdd.n3185 vdd.n831 99.5127
R2733 vdd.n3180 vdd.n3179 99.5127
R2734 vdd.n2898 vdd.n944 99.5127
R2735 vdd.n2898 vdd.n939 99.5127
R2736 vdd.n3000 vdd.n939 99.5127
R2737 vdd.n3000 vdd.n934 99.5127
R2738 vdd.n2996 vdd.n934 99.5127
R2739 vdd.n2996 vdd.n928 99.5127
R2740 vdd.n2993 vdd.n928 99.5127
R2741 vdd.n2993 vdd.n922 99.5127
R2742 vdd.n2990 vdd.n922 99.5127
R2743 vdd.n2990 vdd.n917 99.5127
R2744 vdd.n2940 vdd.n917 99.5127
R2745 vdd.n2940 vdd.n912 99.5127
R2746 vdd.n2943 vdd.n912 99.5127
R2747 vdd.n2943 vdd.n906 99.5127
R2748 vdd.n2976 vdd.n906 99.5127
R2749 vdd.n2976 vdd.n899 99.5127
R2750 vdd.n2972 vdd.n899 99.5127
R2751 vdd.n2972 vdd.n894 99.5127
R2752 vdd.n2969 vdd.n894 99.5127
R2753 vdd.n2969 vdd.n889 99.5127
R2754 vdd.n2966 vdd.n889 99.5127
R2755 vdd.n2966 vdd.n882 99.5127
R2756 vdd.n2963 vdd.n882 99.5127
R2757 vdd.n2963 vdd.n875 99.5127
R2758 vdd.n2960 vdd.n875 99.5127
R2759 vdd.n2960 vdd.n868 99.5127
R2760 vdd.n2957 vdd.n868 99.5127
R2761 vdd.n2957 vdd.n862 99.5127
R2762 vdd.n2954 vdd.n862 99.5127
R2763 vdd.n2954 vdd.n857 99.5127
R2764 vdd.n2951 vdd.n857 99.5127
R2765 vdd.n2951 vdd.n852 99.5127
R2766 vdd.n2948 vdd.n852 99.5127
R2767 vdd.n2948 vdd.n844 99.5127
R2768 vdd.n844 vdd.n837 99.5127
R2769 vdd.n3172 vdd.n837 99.5127
R2770 vdd.n3173 vdd.n3172 99.5127
R2771 vdd.n3173 vdd.n806 99.5127
R2772 vdd.n3012 vdd.n949 99.5127
R2773 vdd.n2832 vdd.n949 99.5127
R2774 vdd.n2836 vdd.n2835 99.5127
R2775 vdd.n2840 vdd.n2839 99.5127
R2776 vdd.n2844 vdd.n2843 99.5127
R2777 vdd.n2848 vdd.n2847 99.5127
R2778 vdd.n2852 vdd.n2851 99.5127
R2779 vdd.n2856 vdd.n2855 99.5127
R2780 vdd.n2860 vdd.n2859 99.5127
R2781 vdd.n2864 vdd.n2863 99.5127
R2782 vdd.n2868 vdd.n2867 99.5127
R2783 vdd.n2872 vdd.n2871 99.5127
R2784 vdd.n2876 vdd.n2875 99.5127
R2785 vdd.n2880 vdd.n2879 99.5127
R2786 vdd.n2884 vdd.n2883 99.5127
R2787 vdd.n2888 vdd.n2887 99.5127
R2788 vdd.n2893 vdd.n2892 99.5127
R2789 vdd.n2725 vdd.n986 99.5127
R2790 vdd.n2721 vdd.n2720 99.5127
R2791 vdd.n2717 vdd.n2716 99.5127
R2792 vdd.n2713 vdd.n2712 99.5127
R2793 vdd.n2709 vdd.n2708 99.5127
R2794 vdd.n2705 vdd.n2704 99.5127
R2795 vdd.n2701 vdd.n2700 99.5127
R2796 vdd.n2697 vdd.n2696 99.5127
R2797 vdd.n2693 vdd.n2692 99.5127
R2798 vdd.n2689 vdd.n2688 99.5127
R2799 vdd.n2685 vdd.n2684 99.5127
R2800 vdd.n2681 vdd.n2680 99.5127
R2801 vdd.n2677 vdd.n2676 99.5127
R2802 vdd.n2673 vdd.n2672 99.5127
R2803 vdd.n2669 vdd.n2668 99.5127
R2804 vdd.n2665 vdd.n2664 99.5127
R2805 vdd.n2660 vdd.n2659 99.5127
R2806 vdd.n2392 vdd.n1111 99.5127
R2807 vdd.n2392 vdd.n1105 99.5127
R2808 vdd.n2389 vdd.n1105 99.5127
R2809 vdd.n2389 vdd.n1099 99.5127
R2810 vdd.n2386 vdd.n1099 99.5127
R2811 vdd.n2386 vdd.n1093 99.5127
R2812 vdd.n2383 vdd.n1093 99.5127
R2813 vdd.n2383 vdd.n1087 99.5127
R2814 vdd.n2380 vdd.n1087 99.5127
R2815 vdd.n2380 vdd.n1081 99.5127
R2816 vdd.n2377 vdd.n1081 99.5127
R2817 vdd.n2377 vdd.n1075 99.5127
R2818 vdd.n2374 vdd.n1075 99.5127
R2819 vdd.n2374 vdd.n1068 99.5127
R2820 vdd.n2371 vdd.n1068 99.5127
R2821 vdd.n2371 vdd.n1061 99.5127
R2822 vdd.n2368 vdd.n1061 99.5127
R2823 vdd.n2368 vdd.n1055 99.5127
R2824 vdd.n2365 vdd.n1055 99.5127
R2825 vdd.n2365 vdd.n1050 99.5127
R2826 vdd.n2362 vdd.n1050 99.5127
R2827 vdd.n2362 vdd.n1044 99.5127
R2828 vdd.n2359 vdd.n1044 99.5127
R2829 vdd.n2359 vdd.n1037 99.5127
R2830 vdd.n2326 vdd.n1037 99.5127
R2831 vdd.n2326 vdd.n1031 99.5127
R2832 vdd.n2329 vdd.n1031 99.5127
R2833 vdd.n2329 vdd.n1026 99.5127
R2834 vdd.n2345 vdd.n1026 99.5127
R2835 vdd.n2345 vdd.n1021 99.5127
R2836 vdd.n2341 vdd.n1021 99.5127
R2837 vdd.n2341 vdd.n1016 99.5127
R2838 vdd.n2338 vdd.n1016 99.5127
R2839 vdd.n2338 vdd.n1009 99.5127
R2840 vdd.n2335 vdd.n1009 99.5127
R2841 vdd.n2335 vdd.n1002 99.5127
R2842 vdd.n1002 vdd.n991 99.5127
R2843 vdd.n2655 vdd.n991 99.5127
R2844 vdd.n2462 vdd.n2460 99.5127
R2845 vdd.n2460 vdd.n2459 99.5127
R2846 vdd.n2456 vdd.n2455 99.5127
R2847 vdd.n2453 vdd.n1117 99.5127
R2848 vdd.n2449 vdd.n2447 99.5127
R2849 vdd.n2445 vdd.n1119 99.5127
R2850 vdd.n2441 vdd.n2439 99.5127
R2851 vdd.n2437 vdd.n1121 99.5127
R2852 vdd.n2433 vdd.n2431 99.5127
R2853 vdd.n2429 vdd.n1123 99.5127
R2854 vdd.n2425 vdd.n2423 99.5127
R2855 vdd.n2421 vdd.n1125 99.5127
R2856 vdd.n2417 vdd.n2415 99.5127
R2857 vdd.n2413 vdd.n1127 99.5127
R2858 vdd.n2409 vdd.n2407 99.5127
R2859 vdd.n2405 vdd.n1129 99.5127
R2860 vdd.n2400 vdd.n2398 99.5127
R2861 vdd.n2466 vdd.n1103 99.5127
R2862 vdd.n2474 vdd.n1103 99.5127
R2863 vdd.n2474 vdd.n1101 99.5127
R2864 vdd.n2478 vdd.n1101 99.5127
R2865 vdd.n2478 vdd.n1091 99.5127
R2866 vdd.n2486 vdd.n1091 99.5127
R2867 vdd.n2486 vdd.n1089 99.5127
R2868 vdd.n2490 vdd.n1089 99.5127
R2869 vdd.n2490 vdd.n1079 99.5127
R2870 vdd.n2498 vdd.n1079 99.5127
R2871 vdd.n2498 vdd.n1077 99.5127
R2872 vdd.n2502 vdd.n1077 99.5127
R2873 vdd.n2502 vdd.n1066 99.5127
R2874 vdd.n2510 vdd.n1066 99.5127
R2875 vdd.n2510 vdd.n1064 99.5127
R2876 vdd.n2514 vdd.n1064 99.5127
R2877 vdd.n2514 vdd.n1054 99.5127
R2878 vdd.n2523 vdd.n1054 99.5127
R2879 vdd.n2523 vdd.n1052 99.5127
R2880 vdd.n2527 vdd.n1052 99.5127
R2881 vdd.n2527 vdd.n1042 99.5127
R2882 vdd.n2535 vdd.n1042 99.5127
R2883 vdd.n2535 vdd.n1040 99.5127
R2884 vdd.n2539 vdd.n1040 99.5127
R2885 vdd.n2539 vdd.n1030 99.5127
R2886 vdd.n2547 vdd.n1030 99.5127
R2887 vdd.n2547 vdd.n1028 99.5127
R2888 vdd.n2551 vdd.n1028 99.5127
R2889 vdd.n2551 vdd.n1020 99.5127
R2890 vdd.n2559 vdd.n1020 99.5127
R2891 vdd.n2559 vdd.n1018 99.5127
R2892 vdd.n2563 vdd.n1018 99.5127
R2893 vdd.n2563 vdd.n1007 99.5127
R2894 vdd.n2573 vdd.n1007 99.5127
R2895 vdd.n2573 vdd.n1004 99.5127
R2896 vdd.n2578 vdd.n1004 99.5127
R2897 vdd.n2578 vdd.n1005 99.5127
R2898 vdd.n1005 vdd.n985 99.5127
R2899 vdd.n3156 vdd.n3155 99.5127
R2900 vdd.n3153 vdd.n3119 99.5127
R2901 vdd.n3149 vdd.n3148 99.5127
R2902 vdd.n3146 vdd.n3122 99.5127
R2903 vdd.n3142 vdd.n3141 99.5127
R2904 vdd.n3139 vdd.n3125 99.5127
R2905 vdd.n3135 vdd.n3134 99.5127
R2906 vdd.n3132 vdd.n3129 99.5127
R2907 vdd.n3273 vdd.n787 99.5127
R2908 vdd.n3271 vdd.n3270 99.5127
R2909 vdd.n3268 vdd.n789 99.5127
R2910 vdd.n3264 vdd.n3263 99.5127
R2911 vdd.n3261 vdd.n792 99.5127
R2912 vdd.n3257 vdd.n3256 99.5127
R2913 vdd.n3254 vdd.n795 99.5127
R2914 vdd.n3250 vdd.n3249 99.5127
R2915 vdd.n3247 vdd.n798 99.5127
R2916 vdd.n3005 vdd.n945 99.5127
R2917 vdd.n3005 vdd.n940 99.5127
R2918 vdd.n3002 vdd.n940 99.5127
R2919 vdd.n3002 vdd.n935 99.5127
R2920 vdd.n2902 vdd.n935 99.5127
R2921 vdd.n2902 vdd.n929 99.5127
R2922 vdd.n2905 vdd.n929 99.5127
R2923 vdd.n2905 vdd.n923 99.5127
R2924 vdd.n2988 vdd.n923 99.5127
R2925 vdd.n2988 vdd.n918 99.5127
R2926 vdd.n2984 vdd.n918 99.5127
R2927 vdd.n2984 vdd.n913 99.5127
R2928 vdd.n2981 vdd.n913 99.5127
R2929 vdd.n2981 vdd.n907 99.5127
R2930 vdd.n2978 vdd.n907 99.5127
R2931 vdd.n2978 vdd.n900 99.5127
R2932 vdd.n2937 vdd.n900 99.5127
R2933 vdd.n2937 vdd.n895 99.5127
R2934 vdd.n2934 vdd.n895 99.5127
R2935 vdd.n2934 vdd.n890 99.5127
R2936 vdd.n2931 vdd.n890 99.5127
R2937 vdd.n2931 vdd.n883 99.5127
R2938 vdd.n2928 vdd.n883 99.5127
R2939 vdd.n2928 vdd.n876 99.5127
R2940 vdd.n2925 vdd.n876 99.5127
R2941 vdd.n2925 vdd.n869 99.5127
R2942 vdd.n2922 vdd.n869 99.5127
R2943 vdd.n2922 vdd.n863 99.5127
R2944 vdd.n2919 vdd.n863 99.5127
R2945 vdd.n2919 vdd.n858 99.5127
R2946 vdd.n2916 vdd.n858 99.5127
R2947 vdd.n2916 vdd.n853 99.5127
R2948 vdd.n2913 vdd.n853 99.5127
R2949 vdd.n2913 vdd.n845 99.5127
R2950 vdd.n2910 vdd.n845 99.5127
R2951 vdd.n2910 vdd.n838 99.5127
R2952 vdd.n838 vdd.n804 99.5127
R2953 vdd.n3242 vdd.n804 99.5127
R2954 vdd.n2766 vdd.n2765 99.5127
R2955 vdd.n2770 vdd.n2769 99.5127
R2956 vdd.n2774 vdd.n2773 99.5127
R2957 vdd.n2778 vdd.n2777 99.5127
R2958 vdd.n2782 vdd.n2781 99.5127
R2959 vdd.n2786 vdd.n2785 99.5127
R2960 vdd.n2790 vdd.n2789 99.5127
R2961 vdd.n2794 vdd.n2793 99.5127
R2962 vdd.n2798 vdd.n2797 99.5127
R2963 vdd.n2802 vdd.n2801 99.5127
R2964 vdd.n2806 vdd.n2805 99.5127
R2965 vdd.n2810 vdd.n2809 99.5127
R2966 vdd.n2814 vdd.n2813 99.5127
R2967 vdd.n2818 vdd.n2817 99.5127
R2968 vdd.n2822 vdd.n2821 99.5127
R2969 vdd.n2826 vdd.n2825 99.5127
R2970 vdd.n3009 vdd.n2760 99.5127
R2971 vdd.n3018 vdd.n941 99.5127
R2972 vdd.n3022 vdd.n941 99.5127
R2973 vdd.n3022 vdd.n933 99.5127
R2974 vdd.n3030 vdd.n933 99.5127
R2975 vdd.n3030 vdd.n931 99.5127
R2976 vdd.n3034 vdd.n931 99.5127
R2977 vdd.n3034 vdd.n921 99.5127
R2978 vdd.n3042 vdd.n921 99.5127
R2979 vdd.n3042 vdd.n919 99.5127
R2980 vdd.n3046 vdd.n919 99.5127
R2981 vdd.n3046 vdd.n910 99.5127
R2982 vdd.n3054 vdd.n910 99.5127
R2983 vdd.n3054 vdd.n908 99.5127
R2984 vdd.n3058 vdd.n908 99.5127
R2985 vdd.n3058 vdd.n898 99.5127
R2986 vdd.n3066 vdd.n898 99.5127
R2987 vdd.n3066 vdd.n896 99.5127
R2988 vdd.n3070 vdd.n896 99.5127
R2989 vdd.n3070 vdd.n887 99.5127
R2990 vdd.n3078 vdd.n887 99.5127
R2991 vdd.n3078 vdd.n884 99.5127
R2992 vdd.n3083 vdd.n884 99.5127
R2993 vdd.n3083 vdd.n873 99.5127
R2994 vdd.n3091 vdd.n873 99.5127
R2995 vdd.n3091 vdd.n871 99.5127
R2996 vdd.n3095 vdd.n871 99.5127
R2997 vdd.n3095 vdd.n861 99.5127
R2998 vdd.n3103 vdd.n861 99.5127
R2999 vdd.n3103 vdd.n859 99.5127
R3000 vdd.n3107 vdd.n859 99.5127
R3001 vdd.n3107 vdd.n850 99.5127
R3002 vdd.n3115 vdd.n850 99.5127
R3003 vdd.n3115 vdd.n847 99.5127
R3004 vdd.n3164 vdd.n847 99.5127
R3005 vdd.n3164 vdd.n848 99.5127
R3006 vdd.n848 vdd.n839 99.5127
R3007 vdd.n3159 vdd.n839 99.5127
R3008 vdd.n3159 vdd.n807 99.5127
R3009 vdd.n2649 vdd.n2648 99.5127
R3010 vdd.n2645 vdd.n2644 99.5127
R3011 vdd.n2641 vdd.n2640 99.5127
R3012 vdd.n2637 vdd.n2636 99.5127
R3013 vdd.n2633 vdd.n2632 99.5127
R3014 vdd.n2629 vdd.n2628 99.5127
R3015 vdd.n2625 vdd.n2624 99.5127
R3016 vdd.n2621 vdd.n2620 99.5127
R3017 vdd.n2617 vdd.n2616 99.5127
R3018 vdd.n2613 vdd.n2612 99.5127
R3019 vdd.n2609 vdd.n2608 99.5127
R3020 vdd.n2605 vdd.n2604 99.5127
R3021 vdd.n2601 vdd.n2600 99.5127
R3022 vdd.n2597 vdd.n2596 99.5127
R3023 vdd.n2593 vdd.n2592 99.5127
R3024 vdd.n2589 vdd.n2588 99.5127
R3025 vdd.n2585 vdd.n967 99.5127
R3026 vdd.n2285 vdd.n1112 99.5127
R3027 vdd.n2285 vdd.n1106 99.5127
R3028 vdd.n2288 vdd.n1106 99.5127
R3029 vdd.n2288 vdd.n1100 99.5127
R3030 vdd.n2291 vdd.n1100 99.5127
R3031 vdd.n2291 vdd.n1094 99.5127
R3032 vdd.n2294 vdd.n1094 99.5127
R3033 vdd.n2294 vdd.n1088 99.5127
R3034 vdd.n2297 vdd.n1088 99.5127
R3035 vdd.n2297 vdd.n1082 99.5127
R3036 vdd.n2300 vdd.n1082 99.5127
R3037 vdd.n2300 vdd.n1076 99.5127
R3038 vdd.n2303 vdd.n1076 99.5127
R3039 vdd.n2303 vdd.n1069 99.5127
R3040 vdd.n2306 vdd.n1069 99.5127
R3041 vdd.n2306 vdd.n1062 99.5127
R3042 vdd.n2309 vdd.n1062 99.5127
R3043 vdd.n2309 vdd.n1056 99.5127
R3044 vdd.n2312 vdd.n1056 99.5127
R3045 vdd.n2312 vdd.n1051 99.5127
R3046 vdd.n2315 vdd.n1051 99.5127
R3047 vdd.n2315 vdd.n1045 99.5127
R3048 vdd.n2357 vdd.n1045 99.5127
R3049 vdd.n2357 vdd.n1038 99.5127
R3050 vdd.n2353 vdd.n1038 99.5127
R3051 vdd.n2353 vdd.n1032 99.5127
R3052 vdd.n2350 vdd.n1032 99.5127
R3053 vdd.n2350 vdd.n1027 99.5127
R3054 vdd.n2347 vdd.n1027 99.5127
R3055 vdd.n2347 vdd.n1022 99.5127
R3056 vdd.n2323 vdd.n1022 99.5127
R3057 vdd.n2323 vdd.n1017 99.5127
R3058 vdd.n2320 vdd.n1017 99.5127
R3059 vdd.n2320 vdd.n1010 99.5127
R3060 vdd.n1010 vdd.n1001 99.5127
R3061 vdd.n2580 vdd.n1001 99.5127
R3062 vdd.n2581 vdd.n2580 99.5127
R3063 vdd.n2581 vdd.n993 99.5127
R3064 vdd.n2218 vdd.n2216 99.5127
R3065 vdd.n2222 vdd.n2213 99.5127
R3066 vdd.n2226 vdd.n2224 99.5127
R3067 vdd.n2230 vdd.n2211 99.5127
R3068 vdd.n2234 vdd.n2232 99.5127
R3069 vdd.n2238 vdd.n2209 99.5127
R3070 vdd.n2242 vdd.n2240 99.5127
R3071 vdd.n2246 vdd.n2207 99.5127
R3072 vdd.n2250 vdd.n2248 99.5127
R3073 vdd.n2254 vdd.n1143 99.5127
R3074 vdd.n2258 vdd.n2256 99.5127
R3075 vdd.n2262 vdd.n1141 99.5127
R3076 vdd.n2266 vdd.n2264 99.5127
R3077 vdd.n2270 vdd.n1139 99.5127
R3078 vdd.n2274 vdd.n2272 99.5127
R3079 vdd.n2279 vdd.n1135 99.5127
R3080 vdd.n2282 vdd.n2281 99.5127
R3081 vdd.n2468 vdd.n1107 99.5127
R3082 vdd.n2472 vdd.n1107 99.5127
R3083 vdd.n2472 vdd.n1097 99.5127
R3084 vdd.n2480 vdd.n1097 99.5127
R3085 vdd.n2480 vdd.n1095 99.5127
R3086 vdd.n2484 vdd.n1095 99.5127
R3087 vdd.n2484 vdd.n1085 99.5127
R3088 vdd.n2492 vdd.n1085 99.5127
R3089 vdd.n2492 vdd.n1083 99.5127
R3090 vdd.n2496 vdd.n1083 99.5127
R3091 vdd.n2496 vdd.n1073 99.5127
R3092 vdd.n2504 vdd.n1073 99.5127
R3093 vdd.n2504 vdd.n1071 99.5127
R3094 vdd.n2508 vdd.n1071 99.5127
R3095 vdd.n2508 vdd.n1060 99.5127
R3096 vdd.n2516 vdd.n1060 99.5127
R3097 vdd.n2516 vdd.n1057 99.5127
R3098 vdd.n2521 vdd.n1057 99.5127
R3099 vdd.n2521 vdd.n1048 99.5127
R3100 vdd.n2529 vdd.n1048 99.5127
R3101 vdd.n2529 vdd.n1046 99.5127
R3102 vdd.n2533 vdd.n1046 99.5127
R3103 vdd.n2533 vdd.n1036 99.5127
R3104 vdd.n2541 vdd.n1036 99.5127
R3105 vdd.n2541 vdd.n1034 99.5127
R3106 vdd.n2545 vdd.n1034 99.5127
R3107 vdd.n2545 vdd.n1025 99.5127
R3108 vdd.n2553 vdd.n1025 99.5127
R3109 vdd.n2553 vdd.n1023 99.5127
R3110 vdd.n2557 vdd.n1023 99.5127
R3111 vdd.n2557 vdd.n1014 99.5127
R3112 vdd.n2565 vdd.n1014 99.5127
R3113 vdd.n2565 vdd.n1011 99.5127
R3114 vdd.n2571 vdd.n1011 99.5127
R3115 vdd.n2571 vdd.n1012 99.5127
R3116 vdd.n1012 vdd.n1003 99.5127
R3117 vdd.n1003 vdd.n994 99.5127
R3118 vdd.n2653 vdd.n994 99.5127
R3119 vdd.n9 vdd.n7 98.9633
R3120 vdd.n2 vdd.n0 98.9633
R3121 vdd.n9 vdd.n8 98.6055
R3122 vdd.n11 vdd.n10 98.6055
R3123 vdd.n13 vdd.n12 98.6055
R3124 vdd.n6 vdd.n5 98.6055
R3125 vdd.n4 vdd.n3 98.6055
R3126 vdd.n2 vdd.n1 98.6055
R3127 vdd.t142 vdd.n303 85.8723
R3128 vdd.t219 vdd.n244 85.8723
R3129 vdd.t145 vdd.n201 85.8723
R3130 vdd.t199 vdd.n142 85.8723
R3131 vdd.t244 vdd.n100 85.8723
R3132 vdd.t268 vdd.n41 85.8723
R3133 vdd.t298 vdd.n1802 85.8723
R3134 vdd.t249 vdd.n1861 85.8723
R3135 vdd.t282 vdd.n1700 85.8723
R3136 vdd.t235 vdd.n1759 85.8723
R3137 vdd.t239 vdd.n1599 85.8723
R3138 vdd.t246 vdd.n1658 85.8723
R3139 vdd.n3080 vdd.n885 78.546
R3140 vdd.n2519 vdd.n1058 78.546
R3141 vdd.n290 vdd.n289 75.1835
R3142 vdd.n288 vdd.n287 75.1835
R3143 vdd.n286 vdd.n285 75.1835
R3144 vdd.n284 vdd.n283 75.1835
R3145 vdd.n282 vdd.n281 75.1835
R3146 vdd.n280 vdd.n279 75.1835
R3147 vdd.n278 vdd.n277 75.1835
R3148 vdd.n276 vdd.n275 75.1835
R3149 vdd.n274 vdd.n273 75.1835
R3150 vdd.n188 vdd.n187 75.1835
R3151 vdd.n186 vdd.n185 75.1835
R3152 vdd.n184 vdd.n183 75.1835
R3153 vdd.n182 vdd.n181 75.1835
R3154 vdd.n180 vdd.n179 75.1835
R3155 vdd.n178 vdd.n177 75.1835
R3156 vdd.n176 vdd.n175 75.1835
R3157 vdd.n174 vdd.n173 75.1835
R3158 vdd.n172 vdd.n171 75.1835
R3159 vdd.n87 vdd.n86 75.1835
R3160 vdd.n85 vdd.n84 75.1835
R3161 vdd.n83 vdd.n82 75.1835
R3162 vdd.n81 vdd.n80 75.1835
R3163 vdd.n79 vdd.n78 75.1835
R3164 vdd.n77 vdd.n76 75.1835
R3165 vdd.n75 vdd.n74 75.1835
R3166 vdd.n73 vdd.n72 75.1835
R3167 vdd.n71 vdd.n70 75.1835
R3168 vdd.n1832 vdd.n1831 75.1835
R3169 vdd.n1834 vdd.n1833 75.1835
R3170 vdd.n1836 vdd.n1835 75.1835
R3171 vdd.n1838 vdd.n1837 75.1835
R3172 vdd.n1840 vdd.n1839 75.1835
R3173 vdd.n1842 vdd.n1841 75.1835
R3174 vdd.n1844 vdd.n1843 75.1835
R3175 vdd.n1846 vdd.n1845 75.1835
R3176 vdd.n1848 vdd.n1847 75.1835
R3177 vdd.n1730 vdd.n1729 75.1835
R3178 vdd.n1732 vdd.n1731 75.1835
R3179 vdd.n1734 vdd.n1733 75.1835
R3180 vdd.n1736 vdd.n1735 75.1835
R3181 vdd.n1738 vdd.n1737 75.1835
R3182 vdd.n1740 vdd.n1739 75.1835
R3183 vdd.n1742 vdd.n1741 75.1835
R3184 vdd.n1744 vdd.n1743 75.1835
R3185 vdd.n1746 vdd.n1745 75.1835
R3186 vdd.n1629 vdd.n1628 75.1835
R3187 vdd.n1631 vdd.n1630 75.1835
R3188 vdd.n1633 vdd.n1632 75.1835
R3189 vdd.n1635 vdd.n1634 75.1835
R3190 vdd.n1637 vdd.n1636 75.1835
R3191 vdd.n1639 vdd.n1638 75.1835
R3192 vdd.n1641 vdd.n1640 75.1835
R3193 vdd.n1643 vdd.n1642 75.1835
R3194 vdd.n1645 vdd.n1644 75.1835
R3195 vdd.n3010 vdd.n2743 72.8958
R3196 vdd.n3010 vdd.n2744 72.8958
R3197 vdd.n3010 vdd.n2745 72.8958
R3198 vdd.n3010 vdd.n2746 72.8958
R3199 vdd.n3010 vdd.n2747 72.8958
R3200 vdd.n3010 vdd.n2748 72.8958
R3201 vdd.n3010 vdd.n2749 72.8958
R3202 vdd.n3010 vdd.n2750 72.8958
R3203 vdd.n3010 vdd.n2751 72.8958
R3204 vdd.n3010 vdd.n2752 72.8958
R3205 vdd.n3010 vdd.n2753 72.8958
R3206 vdd.n3010 vdd.n2754 72.8958
R3207 vdd.n3010 vdd.n2755 72.8958
R3208 vdd.n3010 vdd.n2756 72.8958
R3209 vdd.n3010 vdd.n2757 72.8958
R3210 vdd.n3010 vdd.n2758 72.8958
R3211 vdd.n3010 vdd.n2759 72.8958
R3212 vdd.n803 vdd.n692 72.8958
R3213 vdd.n3248 vdd.n692 72.8958
R3214 vdd.n797 vdd.n692 72.8958
R3215 vdd.n3255 vdd.n692 72.8958
R3216 vdd.n794 vdd.n692 72.8958
R3217 vdd.n3262 vdd.n692 72.8958
R3218 vdd.n791 vdd.n692 72.8958
R3219 vdd.n3269 vdd.n692 72.8958
R3220 vdd.n3272 vdd.n692 72.8958
R3221 vdd.n3128 vdd.n692 72.8958
R3222 vdd.n3133 vdd.n692 72.8958
R3223 vdd.n3127 vdd.n692 72.8958
R3224 vdd.n3140 vdd.n692 72.8958
R3225 vdd.n3124 vdd.n692 72.8958
R3226 vdd.n3147 vdd.n692 72.8958
R3227 vdd.n3121 vdd.n692 72.8958
R3228 vdd.n3154 vdd.n692 72.8958
R3229 vdd.n2461 vdd.n1110 72.8958
R3230 vdd.n1115 vdd.n1110 72.8958
R3231 vdd.n2454 vdd.n1110 72.8958
R3232 vdd.n2448 vdd.n1110 72.8958
R3233 vdd.n2446 vdd.n1110 72.8958
R3234 vdd.n2440 vdd.n1110 72.8958
R3235 vdd.n2438 vdd.n1110 72.8958
R3236 vdd.n2432 vdd.n1110 72.8958
R3237 vdd.n2430 vdd.n1110 72.8958
R3238 vdd.n2424 vdd.n1110 72.8958
R3239 vdd.n2422 vdd.n1110 72.8958
R3240 vdd.n2416 vdd.n1110 72.8958
R3241 vdd.n2414 vdd.n1110 72.8958
R3242 vdd.n2408 vdd.n1110 72.8958
R3243 vdd.n2406 vdd.n1110 72.8958
R3244 vdd.n2399 vdd.n1110 72.8958
R3245 vdd.n2397 vdd.n1110 72.8958
R3246 vdd.n2726 vdd.n968 72.8958
R3247 vdd.n2726 vdd.n969 72.8958
R3248 vdd.n2726 vdd.n970 72.8958
R3249 vdd.n2726 vdd.n971 72.8958
R3250 vdd.n2726 vdd.n972 72.8958
R3251 vdd.n2726 vdd.n973 72.8958
R3252 vdd.n2726 vdd.n974 72.8958
R3253 vdd.n2726 vdd.n975 72.8958
R3254 vdd.n2726 vdd.n976 72.8958
R3255 vdd.n2726 vdd.n977 72.8958
R3256 vdd.n2726 vdd.n978 72.8958
R3257 vdd.n2726 vdd.n979 72.8958
R3258 vdd.n2726 vdd.n980 72.8958
R3259 vdd.n2726 vdd.n981 72.8958
R3260 vdd.n2726 vdd.n982 72.8958
R3261 vdd.n2726 vdd.n983 72.8958
R3262 vdd.n2726 vdd.n984 72.8958
R3263 vdd.n3011 vdd.n3010 72.8958
R3264 vdd.n3010 vdd.n2727 72.8958
R3265 vdd.n3010 vdd.n2728 72.8958
R3266 vdd.n3010 vdd.n2729 72.8958
R3267 vdd.n3010 vdd.n2730 72.8958
R3268 vdd.n3010 vdd.n2731 72.8958
R3269 vdd.n3010 vdd.n2732 72.8958
R3270 vdd.n3010 vdd.n2733 72.8958
R3271 vdd.n3010 vdd.n2734 72.8958
R3272 vdd.n3010 vdd.n2735 72.8958
R3273 vdd.n3010 vdd.n2736 72.8958
R3274 vdd.n3010 vdd.n2737 72.8958
R3275 vdd.n3010 vdd.n2738 72.8958
R3276 vdd.n3010 vdd.n2739 72.8958
R3277 vdd.n3010 vdd.n2740 72.8958
R3278 vdd.n3010 vdd.n2741 72.8958
R3279 vdd.n3010 vdd.n2742 72.8958
R3280 vdd.n3178 vdd.n692 72.8958
R3281 vdd.n835 vdd.n692 72.8958
R3282 vdd.n3186 vdd.n692 72.8958
R3283 vdd.n830 vdd.n692 72.8958
R3284 vdd.n3193 vdd.n692 72.8958
R3285 vdd.n827 vdd.n692 72.8958
R3286 vdd.n3200 vdd.n692 72.8958
R3287 vdd.n824 vdd.n692 72.8958
R3288 vdd.n3207 vdd.n692 72.8958
R3289 vdd.n3211 vdd.n692 72.8958
R3290 vdd.n821 vdd.n692 72.8958
R3291 vdd.n3218 vdd.n692 72.8958
R3292 vdd.n818 vdd.n692 72.8958
R3293 vdd.n3225 vdd.n692 72.8958
R3294 vdd.n815 vdd.n692 72.8958
R3295 vdd.n3232 vdd.n692 72.8958
R3296 vdd.n3235 vdd.n692 72.8958
R3297 vdd.n2726 vdd.n966 72.8958
R3298 vdd.n2726 vdd.n965 72.8958
R3299 vdd.n2726 vdd.n964 72.8958
R3300 vdd.n2726 vdd.n963 72.8958
R3301 vdd.n2726 vdd.n962 72.8958
R3302 vdd.n2726 vdd.n961 72.8958
R3303 vdd.n2726 vdd.n960 72.8958
R3304 vdd.n2726 vdd.n959 72.8958
R3305 vdd.n2726 vdd.n958 72.8958
R3306 vdd.n2726 vdd.n957 72.8958
R3307 vdd.n2726 vdd.n956 72.8958
R3308 vdd.n2726 vdd.n955 72.8958
R3309 vdd.n2726 vdd.n954 72.8958
R3310 vdd.n2726 vdd.n953 72.8958
R3311 vdd.n2726 vdd.n952 72.8958
R3312 vdd.n2726 vdd.n951 72.8958
R3313 vdd.n2726 vdd.n950 72.8958
R3314 vdd.n2215 vdd.n1110 72.8958
R3315 vdd.n2217 vdd.n1110 72.8958
R3316 vdd.n2223 vdd.n1110 72.8958
R3317 vdd.n2225 vdd.n1110 72.8958
R3318 vdd.n2231 vdd.n1110 72.8958
R3319 vdd.n2233 vdd.n1110 72.8958
R3320 vdd.n2239 vdd.n1110 72.8958
R3321 vdd.n2241 vdd.n1110 72.8958
R3322 vdd.n2247 vdd.n1110 72.8958
R3323 vdd.n2249 vdd.n1110 72.8958
R3324 vdd.n2255 vdd.n1110 72.8958
R3325 vdd.n2257 vdd.n1110 72.8958
R3326 vdd.n2263 vdd.n1110 72.8958
R3327 vdd.n2265 vdd.n1110 72.8958
R3328 vdd.n2271 vdd.n1110 72.8958
R3329 vdd.n2273 vdd.n1110 72.8958
R3330 vdd.n2280 vdd.n1110 72.8958
R3331 vdd.n1499 vdd.n1498 66.2847
R3332 vdd.n1498 vdd.n1274 66.2847
R3333 vdd.n1498 vdd.n1275 66.2847
R3334 vdd.n1498 vdd.n1276 66.2847
R3335 vdd.n1498 vdd.n1277 66.2847
R3336 vdd.n1498 vdd.n1278 66.2847
R3337 vdd.n1498 vdd.n1279 66.2847
R3338 vdd.n1498 vdd.n1280 66.2847
R3339 vdd.n1498 vdd.n1281 66.2847
R3340 vdd.n1498 vdd.n1282 66.2847
R3341 vdd.n1498 vdd.n1283 66.2847
R3342 vdd.n1498 vdd.n1284 66.2847
R3343 vdd.n1498 vdd.n1285 66.2847
R3344 vdd.n1498 vdd.n1286 66.2847
R3345 vdd.n1498 vdd.n1287 66.2847
R3346 vdd.n1498 vdd.n1288 66.2847
R3347 vdd.n1498 vdd.n1289 66.2847
R3348 vdd.n1498 vdd.n1290 66.2847
R3349 vdd.n1498 vdd.n1291 66.2847
R3350 vdd.n1498 vdd.n1292 66.2847
R3351 vdd.n1498 vdd.n1293 66.2847
R3352 vdd.n1498 vdd.n1294 66.2847
R3353 vdd.n1498 vdd.n1295 66.2847
R3354 vdd.n1498 vdd.n1296 66.2847
R3355 vdd.n1498 vdd.n1297 66.2847
R3356 vdd.n1498 vdd.n1298 66.2847
R3357 vdd.n1498 vdd.n1299 66.2847
R3358 vdd.n1498 vdd.n1300 66.2847
R3359 vdd.n1498 vdd.n1301 66.2847
R3360 vdd.n1498 vdd.n1302 66.2847
R3361 vdd.n1498 vdd.n1303 66.2847
R3362 vdd.n1153 vdd.n1150 66.2847
R3363 vdd.n2080 vdd.n1153 66.2847
R3364 vdd.n2085 vdd.n1153 66.2847
R3365 vdd.n2090 vdd.n1153 66.2847
R3366 vdd.n2078 vdd.n1153 66.2847
R3367 vdd.n2097 vdd.n1153 66.2847
R3368 vdd.n2070 vdd.n1153 66.2847
R3369 vdd.n2104 vdd.n1153 66.2847
R3370 vdd.n2063 vdd.n1153 66.2847
R3371 vdd.n2111 vdd.n1153 66.2847
R3372 vdd.n2057 vdd.n1153 66.2847
R3373 vdd.n2052 vdd.n1153 66.2847
R3374 vdd.n2122 vdd.n1153 66.2847
R3375 vdd.n2044 vdd.n1153 66.2847
R3376 vdd.n2129 vdd.n1153 66.2847
R3377 vdd.n2037 vdd.n1153 66.2847
R3378 vdd.n2136 vdd.n1153 66.2847
R3379 vdd.n2030 vdd.n1153 66.2847
R3380 vdd.n2143 vdd.n1153 66.2847
R3381 vdd.n2023 vdd.n1153 66.2847
R3382 vdd.n2150 vdd.n1153 66.2847
R3383 vdd.n2017 vdd.n1153 66.2847
R3384 vdd.n2012 vdd.n1153 66.2847
R3385 vdd.n2161 vdd.n1153 66.2847
R3386 vdd.n2004 vdd.n1153 66.2847
R3387 vdd.n2168 vdd.n1153 66.2847
R3388 vdd.n1997 vdd.n1153 66.2847
R3389 vdd.n2175 vdd.n1153 66.2847
R3390 vdd.n2178 vdd.n1153 66.2847
R3391 vdd.n1988 vdd.n1153 66.2847
R3392 vdd.n2187 vdd.n1153 66.2847
R3393 vdd.n1982 vdd.n1153 66.2847
R3394 vdd.n3405 vdd.n3404 66.2847
R3395 vdd.n3405 vdd.n693 66.2847
R3396 vdd.n3405 vdd.n694 66.2847
R3397 vdd.n3405 vdd.n695 66.2847
R3398 vdd.n3405 vdd.n696 66.2847
R3399 vdd.n3405 vdd.n697 66.2847
R3400 vdd.n3405 vdd.n698 66.2847
R3401 vdd.n3405 vdd.n699 66.2847
R3402 vdd.n3405 vdd.n700 66.2847
R3403 vdd.n3405 vdd.n701 66.2847
R3404 vdd.n3405 vdd.n702 66.2847
R3405 vdd.n3405 vdd.n703 66.2847
R3406 vdd.n3405 vdd.n704 66.2847
R3407 vdd.n3405 vdd.n705 66.2847
R3408 vdd.n3405 vdd.n706 66.2847
R3409 vdd.n3405 vdd.n707 66.2847
R3410 vdd.n3405 vdd.n708 66.2847
R3411 vdd.n3405 vdd.n709 66.2847
R3412 vdd.n3405 vdd.n710 66.2847
R3413 vdd.n3405 vdd.n711 66.2847
R3414 vdd.n3405 vdd.n712 66.2847
R3415 vdd.n3405 vdd.n713 66.2847
R3416 vdd.n3405 vdd.n714 66.2847
R3417 vdd.n3405 vdd.n715 66.2847
R3418 vdd.n3405 vdd.n716 66.2847
R3419 vdd.n3405 vdd.n717 66.2847
R3420 vdd.n3405 vdd.n718 66.2847
R3421 vdd.n3405 vdd.n719 66.2847
R3422 vdd.n3405 vdd.n720 66.2847
R3423 vdd.n3405 vdd.n721 66.2847
R3424 vdd.n3405 vdd.n722 66.2847
R3425 vdd.n3536 vdd.n3535 66.2847
R3426 vdd.n3536 vdd.n424 66.2847
R3427 vdd.n3536 vdd.n423 66.2847
R3428 vdd.n3536 vdd.n422 66.2847
R3429 vdd.n3536 vdd.n421 66.2847
R3430 vdd.n3536 vdd.n420 66.2847
R3431 vdd.n3536 vdd.n419 66.2847
R3432 vdd.n3536 vdd.n418 66.2847
R3433 vdd.n3536 vdd.n417 66.2847
R3434 vdd.n3536 vdd.n416 66.2847
R3435 vdd.n3536 vdd.n415 66.2847
R3436 vdd.n3536 vdd.n414 66.2847
R3437 vdd.n3536 vdd.n413 66.2847
R3438 vdd.n3536 vdd.n412 66.2847
R3439 vdd.n3536 vdd.n411 66.2847
R3440 vdd.n3536 vdd.n410 66.2847
R3441 vdd.n3536 vdd.n409 66.2847
R3442 vdd.n3536 vdd.n408 66.2847
R3443 vdd.n3536 vdd.n407 66.2847
R3444 vdd.n3536 vdd.n406 66.2847
R3445 vdd.n3536 vdd.n405 66.2847
R3446 vdd.n3536 vdd.n404 66.2847
R3447 vdd.n3536 vdd.n403 66.2847
R3448 vdd.n3536 vdd.n402 66.2847
R3449 vdd.n3536 vdd.n401 66.2847
R3450 vdd.n3536 vdd.n400 66.2847
R3451 vdd.n3536 vdd.n399 66.2847
R3452 vdd.n3536 vdd.n398 66.2847
R3453 vdd.n3536 vdd.n397 66.2847
R3454 vdd.n3536 vdd.n396 66.2847
R3455 vdd.n3536 vdd.n395 66.2847
R3456 vdd.n3536 vdd.n394 66.2847
R3457 vdd.n467 vdd.n394 52.4337
R3458 vdd.n473 vdd.n395 52.4337
R3459 vdd.n477 vdd.n396 52.4337
R3460 vdd.n483 vdd.n397 52.4337
R3461 vdd.n487 vdd.n398 52.4337
R3462 vdd.n493 vdd.n399 52.4337
R3463 vdd.n497 vdd.n400 52.4337
R3464 vdd.n503 vdd.n401 52.4337
R3465 vdd.n507 vdd.n402 52.4337
R3466 vdd.n513 vdd.n403 52.4337
R3467 vdd.n517 vdd.n404 52.4337
R3468 vdd.n523 vdd.n405 52.4337
R3469 vdd.n527 vdd.n406 52.4337
R3470 vdd.n533 vdd.n407 52.4337
R3471 vdd.n537 vdd.n408 52.4337
R3472 vdd.n543 vdd.n409 52.4337
R3473 vdd.n547 vdd.n410 52.4337
R3474 vdd.n553 vdd.n411 52.4337
R3475 vdd.n557 vdd.n412 52.4337
R3476 vdd.n563 vdd.n413 52.4337
R3477 vdd.n567 vdd.n414 52.4337
R3478 vdd.n573 vdd.n415 52.4337
R3479 vdd.n577 vdd.n416 52.4337
R3480 vdd.n583 vdd.n417 52.4337
R3481 vdd.n587 vdd.n418 52.4337
R3482 vdd.n593 vdd.n419 52.4337
R3483 vdd.n597 vdd.n420 52.4337
R3484 vdd.n603 vdd.n421 52.4337
R3485 vdd.n607 vdd.n422 52.4337
R3486 vdd.n613 vdd.n423 52.4337
R3487 vdd.n616 vdd.n424 52.4337
R3488 vdd.n3535 vdd.n3534 52.4337
R3489 vdd.n3404 vdd.n3403 52.4337
R3490 vdd.n728 vdd.n693 52.4337
R3491 vdd.n734 vdd.n694 52.4337
R3492 vdd.n3393 vdd.n695 52.4337
R3493 vdd.n3389 vdd.n696 52.4337
R3494 vdd.n3385 vdd.n697 52.4337
R3495 vdd.n3381 vdd.n698 52.4337
R3496 vdd.n3377 vdd.n699 52.4337
R3497 vdd.n3373 vdd.n700 52.4337
R3498 vdd.n3369 vdd.n701 52.4337
R3499 vdd.n3361 vdd.n702 52.4337
R3500 vdd.n3357 vdd.n703 52.4337
R3501 vdd.n3353 vdd.n704 52.4337
R3502 vdd.n3349 vdd.n705 52.4337
R3503 vdd.n3345 vdd.n706 52.4337
R3504 vdd.n3341 vdd.n707 52.4337
R3505 vdd.n3337 vdd.n708 52.4337
R3506 vdd.n3333 vdd.n709 52.4337
R3507 vdd.n3329 vdd.n710 52.4337
R3508 vdd.n3325 vdd.n711 52.4337
R3509 vdd.n3321 vdd.n712 52.4337
R3510 vdd.n3315 vdd.n713 52.4337
R3511 vdd.n3311 vdd.n714 52.4337
R3512 vdd.n3307 vdd.n715 52.4337
R3513 vdd.n3303 vdd.n716 52.4337
R3514 vdd.n3299 vdd.n717 52.4337
R3515 vdd.n3295 vdd.n718 52.4337
R3516 vdd.n3291 vdd.n719 52.4337
R3517 vdd.n3287 vdd.n720 52.4337
R3518 vdd.n3283 vdd.n721 52.4337
R3519 vdd.n3279 vdd.n722 52.4337
R3520 vdd.n2189 vdd.n1982 52.4337
R3521 vdd.n2187 vdd.n2186 52.4337
R3522 vdd.n1989 vdd.n1988 52.4337
R3523 vdd.n2178 vdd.n2177 52.4337
R3524 vdd.n2175 vdd.n2174 52.4337
R3525 vdd.n2170 vdd.n1997 52.4337
R3526 vdd.n2168 vdd.n2167 52.4337
R3527 vdd.n2163 vdd.n2004 52.4337
R3528 vdd.n2161 vdd.n2160 52.4337
R3529 vdd.n2013 vdd.n2012 52.4337
R3530 vdd.n2152 vdd.n2017 52.4337
R3531 vdd.n2150 vdd.n2149 52.4337
R3532 vdd.n2145 vdd.n2023 52.4337
R3533 vdd.n2143 vdd.n2142 52.4337
R3534 vdd.n2138 vdd.n2030 52.4337
R3535 vdd.n2136 vdd.n2135 52.4337
R3536 vdd.n2131 vdd.n2037 52.4337
R3537 vdd.n2129 vdd.n2128 52.4337
R3538 vdd.n2124 vdd.n2044 52.4337
R3539 vdd.n2122 vdd.n2121 52.4337
R3540 vdd.n2053 vdd.n2052 52.4337
R3541 vdd.n2113 vdd.n2057 52.4337
R3542 vdd.n2111 vdd.n2110 52.4337
R3543 vdd.n2106 vdd.n2063 52.4337
R3544 vdd.n2104 vdd.n2103 52.4337
R3545 vdd.n2099 vdd.n2070 52.4337
R3546 vdd.n2097 vdd.n2096 52.4337
R3547 vdd.n2092 vdd.n2078 52.4337
R3548 vdd.n2090 vdd.n2089 52.4337
R3549 vdd.n2085 vdd.n2084 52.4337
R3550 vdd.n2080 vdd.n2079 52.4337
R3551 vdd.n2198 vdd.n1150 52.4337
R3552 vdd.n1500 vdd.n1499 52.4337
R3553 vdd.n1306 vdd.n1274 52.4337
R3554 vdd.n1310 vdd.n1275 52.4337
R3555 vdd.n1312 vdd.n1276 52.4337
R3556 vdd.n1316 vdd.n1277 52.4337
R3557 vdd.n1318 vdd.n1278 52.4337
R3558 vdd.n1322 vdd.n1279 52.4337
R3559 vdd.n1324 vdd.n1280 52.4337
R3560 vdd.n1328 vdd.n1281 52.4337
R3561 vdd.n1330 vdd.n1282 52.4337
R3562 vdd.n1336 vdd.n1283 52.4337
R3563 vdd.n1338 vdd.n1284 52.4337
R3564 vdd.n1342 vdd.n1285 52.4337
R3565 vdd.n1344 vdd.n1286 52.4337
R3566 vdd.n1348 vdd.n1287 52.4337
R3567 vdd.n1350 vdd.n1288 52.4337
R3568 vdd.n1354 vdd.n1289 52.4337
R3569 vdd.n1356 vdd.n1290 52.4337
R3570 vdd.n1360 vdd.n1291 52.4337
R3571 vdd.n1362 vdd.n1292 52.4337
R3572 vdd.n1434 vdd.n1293 52.4337
R3573 vdd.n1367 vdd.n1294 52.4337
R3574 vdd.n1371 vdd.n1295 52.4337
R3575 vdd.n1373 vdd.n1296 52.4337
R3576 vdd.n1377 vdd.n1297 52.4337
R3577 vdd.n1379 vdd.n1298 52.4337
R3578 vdd.n1383 vdd.n1299 52.4337
R3579 vdd.n1385 vdd.n1300 52.4337
R3580 vdd.n1389 vdd.n1301 52.4337
R3581 vdd.n1391 vdd.n1302 52.4337
R3582 vdd.n1395 vdd.n1303 52.4337
R3583 vdd.n1499 vdd.n1273 52.4337
R3584 vdd.n1309 vdd.n1274 52.4337
R3585 vdd.n1311 vdd.n1275 52.4337
R3586 vdd.n1315 vdd.n1276 52.4337
R3587 vdd.n1317 vdd.n1277 52.4337
R3588 vdd.n1321 vdd.n1278 52.4337
R3589 vdd.n1323 vdd.n1279 52.4337
R3590 vdd.n1327 vdd.n1280 52.4337
R3591 vdd.n1329 vdd.n1281 52.4337
R3592 vdd.n1335 vdd.n1282 52.4337
R3593 vdd.n1337 vdd.n1283 52.4337
R3594 vdd.n1341 vdd.n1284 52.4337
R3595 vdd.n1343 vdd.n1285 52.4337
R3596 vdd.n1347 vdd.n1286 52.4337
R3597 vdd.n1349 vdd.n1287 52.4337
R3598 vdd.n1353 vdd.n1288 52.4337
R3599 vdd.n1355 vdd.n1289 52.4337
R3600 vdd.n1359 vdd.n1290 52.4337
R3601 vdd.n1361 vdd.n1291 52.4337
R3602 vdd.n1365 vdd.n1292 52.4337
R3603 vdd.n1366 vdd.n1293 52.4337
R3604 vdd.n1370 vdd.n1294 52.4337
R3605 vdd.n1372 vdd.n1295 52.4337
R3606 vdd.n1376 vdd.n1296 52.4337
R3607 vdd.n1378 vdd.n1297 52.4337
R3608 vdd.n1382 vdd.n1298 52.4337
R3609 vdd.n1384 vdd.n1299 52.4337
R3610 vdd.n1388 vdd.n1300 52.4337
R3611 vdd.n1390 vdd.n1301 52.4337
R3612 vdd.n1394 vdd.n1302 52.4337
R3613 vdd.n1396 vdd.n1303 52.4337
R3614 vdd.n1150 vdd.n1149 52.4337
R3615 vdd.n2081 vdd.n2080 52.4337
R3616 vdd.n2086 vdd.n2085 52.4337
R3617 vdd.n2091 vdd.n2090 52.4337
R3618 vdd.n2078 vdd.n2071 52.4337
R3619 vdd.n2098 vdd.n2097 52.4337
R3620 vdd.n2070 vdd.n2064 52.4337
R3621 vdd.n2105 vdd.n2104 52.4337
R3622 vdd.n2063 vdd.n2058 52.4337
R3623 vdd.n2112 vdd.n2111 52.4337
R3624 vdd.n2057 vdd.n2056 52.4337
R3625 vdd.n2052 vdd.n2045 52.4337
R3626 vdd.n2123 vdd.n2122 52.4337
R3627 vdd.n2044 vdd.n2038 52.4337
R3628 vdd.n2130 vdd.n2129 52.4337
R3629 vdd.n2037 vdd.n2031 52.4337
R3630 vdd.n2137 vdd.n2136 52.4337
R3631 vdd.n2030 vdd.n2024 52.4337
R3632 vdd.n2144 vdd.n2143 52.4337
R3633 vdd.n2023 vdd.n2018 52.4337
R3634 vdd.n2151 vdd.n2150 52.4337
R3635 vdd.n2017 vdd.n2016 52.4337
R3636 vdd.n2012 vdd.n2005 52.4337
R3637 vdd.n2162 vdd.n2161 52.4337
R3638 vdd.n2004 vdd.n1998 52.4337
R3639 vdd.n2169 vdd.n2168 52.4337
R3640 vdd.n1997 vdd.n1991 52.4337
R3641 vdd.n2176 vdd.n2175 52.4337
R3642 vdd.n2179 vdd.n2178 52.4337
R3643 vdd.n1988 vdd.n1983 52.4337
R3644 vdd.n2188 vdd.n2187 52.4337
R3645 vdd.n1982 vdd.n1155 52.4337
R3646 vdd.n3404 vdd.n725 52.4337
R3647 vdd.n733 vdd.n693 52.4337
R3648 vdd.n3394 vdd.n694 52.4337
R3649 vdd.n3390 vdd.n695 52.4337
R3650 vdd.n3386 vdd.n696 52.4337
R3651 vdd.n3382 vdd.n697 52.4337
R3652 vdd.n3378 vdd.n698 52.4337
R3653 vdd.n3374 vdd.n699 52.4337
R3654 vdd.n3370 vdd.n700 52.4337
R3655 vdd.n3360 vdd.n701 52.4337
R3656 vdd.n3358 vdd.n702 52.4337
R3657 vdd.n3354 vdd.n703 52.4337
R3658 vdd.n3350 vdd.n704 52.4337
R3659 vdd.n3346 vdd.n705 52.4337
R3660 vdd.n3342 vdd.n706 52.4337
R3661 vdd.n3338 vdd.n707 52.4337
R3662 vdd.n3334 vdd.n708 52.4337
R3663 vdd.n3330 vdd.n709 52.4337
R3664 vdd.n3326 vdd.n710 52.4337
R3665 vdd.n3322 vdd.n711 52.4337
R3666 vdd.n3314 vdd.n712 52.4337
R3667 vdd.n3312 vdd.n713 52.4337
R3668 vdd.n3308 vdd.n714 52.4337
R3669 vdd.n3304 vdd.n715 52.4337
R3670 vdd.n3300 vdd.n716 52.4337
R3671 vdd.n3296 vdd.n717 52.4337
R3672 vdd.n3292 vdd.n718 52.4337
R3673 vdd.n3288 vdd.n719 52.4337
R3674 vdd.n3284 vdd.n720 52.4337
R3675 vdd.n3280 vdd.n721 52.4337
R3676 vdd.n722 vdd.n691 52.4337
R3677 vdd.n3535 vdd.n425 52.4337
R3678 vdd.n614 vdd.n424 52.4337
R3679 vdd.n608 vdd.n423 52.4337
R3680 vdd.n604 vdd.n422 52.4337
R3681 vdd.n598 vdd.n421 52.4337
R3682 vdd.n594 vdd.n420 52.4337
R3683 vdd.n588 vdd.n419 52.4337
R3684 vdd.n584 vdd.n418 52.4337
R3685 vdd.n578 vdd.n417 52.4337
R3686 vdd.n574 vdd.n416 52.4337
R3687 vdd.n568 vdd.n415 52.4337
R3688 vdd.n564 vdd.n414 52.4337
R3689 vdd.n558 vdd.n413 52.4337
R3690 vdd.n554 vdd.n412 52.4337
R3691 vdd.n548 vdd.n411 52.4337
R3692 vdd.n544 vdd.n410 52.4337
R3693 vdd.n538 vdd.n409 52.4337
R3694 vdd.n534 vdd.n408 52.4337
R3695 vdd.n528 vdd.n407 52.4337
R3696 vdd.n524 vdd.n406 52.4337
R3697 vdd.n518 vdd.n405 52.4337
R3698 vdd.n514 vdd.n404 52.4337
R3699 vdd.n508 vdd.n403 52.4337
R3700 vdd.n504 vdd.n402 52.4337
R3701 vdd.n498 vdd.n401 52.4337
R3702 vdd.n494 vdd.n400 52.4337
R3703 vdd.n488 vdd.n399 52.4337
R3704 vdd.n484 vdd.n398 52.4337
R3705 vdd.n478 vdd.n397 52.4337
R3706 vdd.n474 vdd.n396 52.4337
R3707 vdd.n468 vdd.n395 52.4337
R3708 vdd.n394 vdd.n392 52.4337
R3709 vdd.t0 vdd.t10 51.4683
R3710 vdd.n274 vdd.n272 42.0461
R3711 vdd.n172 vdd.n170 42.0461
R3712 vdd.n71 vdd.n69 42.0461
R3713 vdd.n1832 vdd.n1830 42.0461
R3714 vdd.n1730 vdd.n1728 42.0461
R3715 vdd.n1629 vdd.n1627 42.0461
R3716 vdd.n332 vdd.n331 41.6884
R3717 vdd.n230 vdd.n229 41.6884
R3718 vdd.n129 vdd.n128 41.6884
R3719 vdd.n1890 vdd.n1889 41.6884
R3720 vdd.n1788 vdd.n1787 41.6884
R3721 vdd.n1687 vdd.n1686 41.6884
R3722 vdd.n1399 vdd.n1398 41.1157
R3723 vdd.n1437 vdd.n1436 41.1157
R3724 vdd.n1333 vdd.n1332 41.1157
R3725 vdd.n428 vdd.n427 41.1157
R3726 vdd.n566 vdd.n441 41.1157
R3727 vdd.n454 vdd.n453 41.1157
R3728 vdd.n3235 vdd.n3234 39.2114
R3729 vdd.n3232 vdd.n3231 39.2114
R3730 vdd.n3227 vdd.n815 39.2114
R3731 vdd.n3225 vdd.n3224 39.2114
R3732 vdd.n3220 vdd.n818 39.2114
R3733 vdd.n3218 vdd.n3217 39.2114
R3734 vdd.n3213 vdd.n821 39.2114
R3735 vdd.n3211 vdd.n3210 39.2114
R3736 vdd.n3207 vdd.n3206 39.2114
R3737 vdd.n3202 vdd.n824 39.2114
R3738 vdd.n3200 vdd.n3199 39.2114
R3739 vdd.n3195 vdd.n827 39.2114
R3740 vdd.n3193 vdd.n3192 39.2114
R3741 vdd.n3188 vdd.n830 39.2114
R3742 vdd.n3186 vdd.n3185 39.2114
R3743 vdd.n3180 vdd.n835 39.2114
R3744 vdd.n3178 vdd.n3177 39.2114
R3745 vdd.n3011 vdd.n947 39.2114
R3746 vdd.n2832 vdd.n2727 39.2114
R3747 vdd.n2836 vdd.n2728 39.2114
R3748 vdd.n2840 vdd.n2729 39.2114
R3749 vdd.n2844 vdd.n2730 39.2114
R3750 vdd.n2848 vdd.n2731 39.2114
R3751 vdd.n2852 vdd.n2732 39.2114
R3752 vdd.n2856 vdd.n2733 39.2114
R3753 vdd.n2860 vdd.n2734 39.2114
R3754 vdd.n2864 vdd.n2735 39.2114
R3755 vdd.n2868 vdd.n2736 39.2114
R3756 vdd.n2872 vdd.n2737 39.2114
R3757 vdd.n2876 vdd.n2738 39.2114
R3758 vdd.n2880 vdd.n2739 39.2114
R3759 vdd.n2884 vdd.n2740 39.2114
R3760 vdd.n2888 vdd.n2741 39.2114
R3761 vdd.n2893 vdd.n2742 39.2114
R3762 vdd.n2721 vdd.n984 39.2114
R3763 vdd.n2717 vdd.n983 39.2114
R3764 vdd.n2713 vdd.n982 39.2114
R3765 vdd.n2709 vdd.n981 39.2114
R3766 vdd.n2705 vdd.n980 39.2114
R3767 vdd.n2701 vdd.n979 39.2114
R3768 vdd.n2697 vdd.n978 39.2114
R3769 vdd.n2693 vdd.n977 39.2114
R3770 vdd.n2689 vdd.n976 39.2114
R3771 vdd.n2685 vdd.n975 39.2114
R3772 vdd.n2681 vdd.n974 39.2114
R3773 vdd.n2677 vdd.n973 39.2114
R3774 vdd.n2673 vdd.n972 39.2114
R3775 vdd.n2669 vdd.n971 39.2114
R3776 vdd.n2665 vdd.n970 39.2114
R3777 vdd.n2660 vdd.n969 39.2114
R3778 vdd.n2656 vdd.n968 39.2114
R3779 vdd.n2461 vdd.n1113 39.2114
R3780 vdd.n2459 vdd.n1115 39.2114
R3781 vdd.n2455 vdd.n2454 39.2114
R3782 vdd.n2448 vdd.n1117 39.2114
R3783 vdd.n2447 vdd.n2446 39.2114
R3784 vdd.n2440 vdd.n1119 39.2114
R3785 vdd.n2439 vdd.n2438 39.2114
R3786 vdd.n2432 vdd.n1121 39.2114
R3787 vdd.n2431 vdd.n2430 39.2114
R3788 vdd.n2424 vdd.n1123 39.2114
R3789 vdd.n2423 vdd.n2422 39.2114
R3790 vdd.n2416 vdd.n1125 39.2114
R3791 vdd.n2415 vdd.n2414 39.2114
R3792 vdd.n2408 vdd.n1127 39.2114
R3793 vdd.n2407 vdd.n2406 39.2114
R3794 vdd.n2399 vdd.n1129 39.2114
R3795 vdd.n2398 vdd.n2397 39.2114
R3796 vdd.n3154 vdd.n3153 39.2114
R3797 vdd.n3149 vdd.n3121 39.2114
R3798 vdd.n3147 vdd.n3146 39.2114
R3799 vdd.n3142 vdd.n3124 39.2114
R3800 vdd.n3140 vdd.n3139 39.2114
R3801 vdd.n3135 vdd.n3127 39.2114
R3802 vdd.n3133 vdd.n3132 39.2114
R3803 vdd.n3128 vdd.n787 39.2114
R3804 vdd.n3272 vdd.n3271 39.2114
R3805 vdd.n3269 vdd.n3268 39.2114
R3806 vdd.n3264 vdd.n791 39.2114
R3807 vdd.n3262 vdd.n3261 39.2114
R3808 vdd.n3257 vdd.n794 39.2114
R3809 vdd.n3255 vdd.n3254 39.2114
R3810 vdd.n3250 vdd.n797 39.2114
R3811 vdd.n3248 vdd.n3247 39.2114
R3812 vdd.n3243 vdd.n803 39.2114
R3813 vdd.n2743 vdd.n943 39.2114
R3814 vdd.n2766 vdd.n2744 39.2114
R3815 vdd.n2770 vdd.n2745 39.2114
R3816 vdd.n2774 vdd.n2746 39.2114
R3817 vdd.n2778 vdd.n2747 39.2114
R3818 vdd.n2782 vdd.n2748 39.2114
R3819 vdd.n2786 vdd.n2749 39.2114
R3820 vdd.n2790 vdd.n2750 39.2114
R3821 vdd.n2794 vdd.n2751 39.2114
R3822 vdd.n2798 vdd.n2752 39.2114
R3823 vdd.n2802 vdd.n2753 39.2114
R3824 vdd.n2806 vdd.n2754 39.2114
R3825 vdd.n2810 vdd.n2755 39.2114
R3826 vdd.n2814 vdd.n2756 39.2114
R3827 vdd.n2818 vdd.n2757 39.2114
R3828 vdd.n2822 vdd.n2758 39.2114
R3829 vdd.n2826 vdd.n2759 39.2114
R3830 vdd.n2765 vdd.n2743 39.2114
R3831 vdd.n2769 vdd.n2744 39.2114
R3832 vdd.n2773 vdd.n2745 39.2114
R3833 vdd.n2777 vdd.n2746 39.2114
R3834 vdd.n2781 vdd.n2747 39.2114
R3835 vdd.n2785 vdd.n2748 39.2114
R3836 vdd.n2789 vdd.n2749 39.2114
R3837 vdd.n2793 vdd.n2750 39.2114
R3838 vdd.n2797 vdd.n2751 39.2114
R3839 vdd.n2801 vdd.n2752 39.2114
R3840 vdd.n2805 vdd.n2753 39.2114
R3841 vdd.n2809 vdd.n2754 39.2114
R3842 vdd.n2813 vdd.n2755 39.2114
R3843 vdd.n2817 vdd.n2756 39.2114
R3844 vdd.n2821 vdd.n2757 39.2114
R3845 vdd.n2825 vdd.n2758 39.2114
R3846 vdd.n2760 vdd.n2759 39.2114
R3847 vdd.n803 vdd.n798 39.2114
R3848 vdd.n3249 vdd.n3248 39.2114
R3849 vdd.n797 vdd.n795 39.2114
R3850 vdd.n3256 vdd.n3255 39.2114
R3851 vdd.n794 vdd.n792 39.2114
R3852 vdd.n3263 vdd.n3262 39.2114
R3853 vdd.n791 vdd.n789 39.2114
R3854 vdd.n3270 vdd.n3269 39.2114
R3855 vdd.n3273 vdd.n3272 39.2114
R3856 vdd.n3129 vdd.n3128 39.2114
R3857 vdd.n3134 vdd.n3133 39.2114
R3858 vdd.n3127 vdd.n3125 39.2114
R3859 vdd.n3141 vdd.n3140 39.2114
R3860 vdd.n3124 vdd.n3122 39.2114
R3861 vdd.n3148 vdd.n3147 39.2114
R3862 vdd.n3121 vdd.n3119 39.2114
R3863 vdd.n3155 vdd.n3154 39.2114
R3864 vdd.n2462 vdd.n2461 39.2114
R3865 vdd.n2456 vdd.n1115 39.2114
R3866 vdd.n2454 vdd.n2453 39.2114
R3867 vdd.n2449 vdd.n2448 39.2114
R3868 vdd.n2446 vdd.n2445 39.2114
R3869 vdd.n2441 vdd.n2440 39.2114
R3870 vdd.n2438 vdd.n2437 39.2114
R3871 vdd.n2433 vdd.n2432 39.2114
R3872 vdd.n2430 vdd.n2429 39.2114
R3873 vdd.n2425 vdd.n2424 39.2114
R3874 vdd.n2422 vdd.n2421 39.2114
R3875 vdd.n2417 vdd.n2416 39.2114
R3876 vdd.n2414 vdd.n2413 39.2114
R3877 vdd.n2409 vdd.n2408 39.2114
R3878 vdd.n2406 vdd.n2405 39.2114
R3879 vdd.n2400 vdd.n2399 39.2114
R3880 vdd.n2397 vdd.n2396 39.2114
R3881 vdd.n2659 vdd.n968 39.2114
R3882 vdd.n2664 vdd.n969 39.2114
R3883 vdd.n2668 vdd.n970 39.2114
R3884 vdd.n2672 vdd.n971 39.2114
R3885 vdd.n2676 vdd.n972 39.2114
R3886 vdd.n2680 vdd.n973 39.2114
R3887 vdd.n2684 vdd.n974 39.2114
R3888 vdd.n2688 vdd.n975 39.2114
R3889 vdd.n2692 vdd.n976 39.2114
R3890 vdd.n2696 vdd.n977 39.2114
R3891 vdd.n2700 vdd.n978 39.2114
R3892 vdd.n2704 vdd.n979 39.2114
R3893 vdd.n2708 vdd.n980 39.2114
R3894 vdd.n2712 vdd.n981 39.2114
R3895 vdd.n2716 vdd.n982 39.2114
R3896 vdd.n2720 vdd.n983 39.2114
R3897 vdd.n986 vdd.n984 39.2114
R3898 vdd.n3012 vdd.n3011 39.2114
R3899 vdd.n2835 vdd.n2727 39.2114
R3900 vdd.n2839 vdd.n2728 39.2114
R3901 vdd.n2843 vdd.n2729 39.2114
R3902 vdd.n2847 vdd.n2730 39.2114
R3903 vdd.n2851 vdd.n2731 39.2114
R3904 vdd.n2855 vdd.n2732 39.2114
R3905 vdd.n2859 vdd.n2733 39.2114
R3906 vdd.n2863 vdd.n2734 39.2114
R3907 vdd.n2867 vdd.n2735 39.2114
R3908 vdd.n2871 vdd.n2736 39.2114
R3909 vdd.n2875 vdd.n2737 39.2114
R3910 vdd.n2879 vdd.n2738 39.2114
R3911 vdd.n2883 vdd.n2739 39.2114
R3912 vdd.n2887 vdd.n2740 39.2114
R3913 vdd.n2892 vdd.n2741 39.2114
R3914 vdd.n2895 vdd.n2742 39.2114
R3915 vdd.n3179 vdd.n3178 39.2114
R3916 vdd.n835 vdd.n831 39.2114
R3917 vdd.n3187 vdd.n3186 39.2114
R3918 vdd.n830 vdd.n828 39.2114
R3919 vdd.n3194 vdd.n3193 39.2114
R3920 vdd.n827 vdd.n825 39.2114
R3921 vdd.n3201 vdd.n3200 39.2114
R3922 vdd.n824 vdd.n822 39.2114
R3923 vdd.n3208 vdd.n3207 39.2114
R3924 vdd.n3212 vdd.n3211 39.2114
R3925 vdd.n821 vdd.n819 39.2114
R3926 vdd.n3219 vdd.n3218 39.2114
R3927 vdd.n818 vdd.n816 39.2114
R3928 vdd.n3226 vdd.n3225 39.2114
R3929 vdd.n815 vdd.n813 39.2114
R3930 vdd.n3233 vdd.n3232 39.2114
R3931 vdd.n3236 vdd.n3235 39.2114
R3932 vdd.n995 vdd.n950 39.2114
R3933 vdd.n2648 vdd.n951 39.2114
R3934 vdd.n2644 vdd.n952 39.2114
R3935 vdd.n2640 vdd.n953 39.2114
R3936 vdd.n2636 vdd.n954 39.2114
R3937 vdd.n2632 vdd.n955 39.2114
R3938 vdd.n2628 vdd.n956 39.2114
R3939 vdd.n2624 vdd.n957 39.2114
R3940 vdd.n2620 vdd.n958 39.2114
R3941 vdd.n2616 vdd.n959 39.2114
R3942 vdd.n2612 vdd.n960 39.2114
R3943 vdd.n2608 vdd.n961 39.2114
R3944 vdd.n2604 vdd.n962 39.2114
R3945 vdd.n2600 vdd.n963 39.2114
R3946 vdd.n2596 vdd.n964 39.2114
R3947 vdd.n2592 vdd.n965 39.2114
R3948 vdd.n2588 vdd.n966 39.2114
R3949 vdd.n2215 vdd.n1109 39.2114
R3950 vdd.n2218 vdd.n2217 39.2114
R3951 vdd.n2223 vdd.n2222 39.2114
R3952 vdd.n2226 vdd.n2225 39.2114
R3953 vdd.n2231 vdd.n2230 39.2114
R3954 vdd.n2234 vdd.n2233 39.2114
R3955 vdd.n2239 vdd.n2238 39.2114
R3956 vdd.n2242 vdd.n2241 39.2114
R3957 vdd.n2247 vdd.n2246 39.2114
R3958 vdd.n2250 vdd.n2249 39.2114
R3959 vdd.n2255 vdd.n2254 39.2114
R3960 vdd.n2258 vdd.n2257 39.2114
R3961 vdd.n2263 vdd.n2262 39.2114
R3962 vdd.n2266 vdd.n2265 39.2114
R3963 vdd.n2271 vdd.n2270 39.2114
R3964 vdd.n2274 vdd.n2273 39.2114
R3965 vdd.n2280 vdd.n2279 39.2114
R3966 vdd.n2585 vdd.n966 39.2114
R3967 vdd.n2589 vdd.n965 39.2114
R3968 vdd.n2593 vdd.n964 39.2114
R3969 vdd.n2597 vdd.n963 39.2114
R3970 vdd.n2601 vdd.n962 39.2114
R3971 vdd.n2605 vdd.n961 39.2114
R3972 vdd.n2609 vdd.n960 39.2114
R3973 vdd.n2613 vdd.n959 39.2114
R3974 vdd.n2617 vdd.n958 39.2114
R3975 vdd.n2621 vdd.n957 39.2114
R3976 vdd.n2625 vdd.n956 39.2114
R3977 vdd.n2629 vdd.n955 39.2114
R3978 vdd.n2633 vdd.n954 39.2114
R3979 vdd.n2637 vdd.n953 39.2114
R3980 vdd.n2641 vdd.n952 39.2114
R3981 vdd.n2645 vdd.n951 39.2114
R3982 vdd.n2649 vdd.n950 39.2114
R3983 vdd.n2216 vdd.n2215 39.2114
R3984 vdd.n2217 vdd.n2213 39.2114
R3985 vdd.n2224 vdd.n2223 39.2114
R3986 vdd.n2225 vdd.n2211 39.2114
R3987 vdd.n2232 vdd.n2231 39.2114
R3988 vdd.n2233 vdd.n2209 39.2114
R3989 vdd.n2240 vdd.n2239 39.2114
R3990 vdd.n2241 vdd.n2207 39.2114
R3991 vdd.n2248 vdd.n2247 39.2114
R3992 vdd.n2249 vdd.n1143 39.2114
R3993 vdd.n2256 vdd.n2255 39.2114
R3994 vdd.n2257 vdd.n1141 39.2114
R3995 vdd.n2264 vdd.n2263 39.2114
R3996 vdd.n2265 vdd.n1139 39.2114
R3997 vdd.n2272 vdd.n2271 39.2114
R3998 vdd.n2273 vdd.n1135 39.2114
R3999 vdd.n2281 vdd.n2280 39.2114
R4000 vdd.n2202 vdd.n2201 37.2369
R4001 vdd.n2118 vdd.n2051 37.2369
R4002 vdd.n2157 vdd.n2011 37.2369
R4003 vdd.n3320 vdd.n769 37.2369
R4004 vdd.n3368 vdd.n3367 37.2369
R4005 vdd.n690 vdd.n689 37.2369
R4006 vdd.n2277 vdd.n1137 30.449
R4007 vdd.n999 vdd.n998 30.449
R4008 vdd.n2402 vdd.n1131 30.449
R4009 vdd.n2662 vdd.n989 30.449
R4010 vdd.n2763 vdd.n2762 30.449
R4011 vdd.n3182 vdd.n833 30.449
R4012 vdd.n2890 vdd.n2831 30.449
R4013 vdd.n801 vdd.n800 30.449
R4014 vdd.n2465 vdd.n2464 30.4395
R4015 vdd.n2724 vdd.n987 30.4395
R4016 vdd.n2657 vdd.n990 30.4395
R4017 vdd.n2395 vdd.n2394 30.4395
R4018 vdd.n2897 vdd.n2896 30.4395
R4019 vdd.n3176 vdd.n3175 30.4395
R4020 vdd.n3015 vdd.n3014 30.4395
R4021 vdd.n3239 vdd.n3238 30.4395
R4022 vdd.n3158 vdd.n3157 30.4395
R4023 vdd.n3244 vdd.n802 30.4395
R4024 vdd.n3008 vdd.n3007 30.4395
R4025 vdd.n3019 vdd.n942 30.4395
R4026 vdd.n2469 vdd.n1108 30.4395
R4027 vdd.n2652 vdd.n2651 30.4395
R4028 vdd.n2584 vdd.n2583 30.4395
R4029 vdd.n2284 vdd.n2283 30.4395
R4030 vdd.n1498 vdd.n1305 22.2201
R4031 vdd.n2196 vdd.n1153 22.2201
R4032 vdd.n3405 vdd.n723 22.2201
R4033 vdd.n3537 vdd.n3536 22.2201
R4034 vdd.n1509 vdd.n1267 19.3944
R4035 vdd.n1509 vdd.n1265 19.3944
R4036 vdd.n1513 vdd.n1265 19.3944
R4037 vdd.n1513 vdd.n1255 19.3944
R4038 vdd.n1526 vdd.n1255 19.3944
R4039 vdd.n1526 vdd.n1253 19.3944
R4040 vdd.n1530 vdd.n1253 19.3944
R4041 vdd.n1530 vdd.n1245 19.3944
R4042 vdd.n1543 vdd.n1245 19.3944
R4043 vdd.n1543 vdd.n1243 19.3944
R4044 vdd.n1547 vdd.n1243 19.3944
R4045 vdd.n1547 vdd.n1232 19.3944
R4046 vdd.n1559 vdd.n1232 19.3944
R4047 vdd.n1559 vdd.n1230 19.3944
R4048 vdd.n1563 vdd.n1230 19.3944
R4049 vdd.n1563 vdd.n1221 19.3944
R4050 vdd.n1576 vdd.n1221 19.3944
R4051 vdd.n1576 vdd.n1219 19.3944
R4052 vdd.n1580 vdd.n1219 19.3944
R4053 vdd.n1580 vdd.n1210 19.3944
R4054 vdd.n1899 vdd.n1210 19.3944
R4055 vdd.n1899 vdd.n1208 19.3944
R4056 vdd.n1903 vdd.n1208 19.3944
R4057 vdd.n1903 vdd.n1198 19.3944
R4058 vdd.n1916 vdd.n1198 19.3944
R4059 vdd.n1916 vdd.n1196 19.3944
R4060 vdd.n1920 vdd.n1196 19.3944
R4061 vdd.n1920 vdd.n1188 19.3944
R4062 vdd.n1933 vdd.n1188 19.3944
R4063 vdd.n1933 vdd.n1186 19.3944
R4064 vdd.n1937 vdd.n1186 19.3944
R4065 vdd.n1937 vdd.n1175 19.3944
R4066 vdd.n1949 vdd.n1175 19.3944
R4067 vdd.n1949 vdd.n1173 19.3944
R4068 vdd.n1953 vdd.n1173 19.3944
R4069 vdd.n1953 vdd.n1165 19.3944
R4070 vdd.n1966 vdd.n1165 19.3944
R4071 vdd.n1966 vdd.n1162 19.3944
R4072 vdd.n1972 vdd.n1162 19.3944
R4073 vdd.n1972 vdd.n1163 19.3944
R4074 vdd.n1163 vdd.n1152 19.3944
R4075 vdd.n1433 vdd.n1368 19.3944
R4076 vdd.n1429 vdd.n1368 19.3944
R4077 vdd.n1429 vdd.n1428 19.3944
R4078 vdd.n1428 vdd.n1427 19.3944
R4079 vdd.n1427 vdd.n1374 19.3944
R4080 vdd.n1423 vdd.n1374 19.3944
R4081 vdd.n1423 vdd.n1422 19.3944
R4082 vdd.n1422 vdd.n1421 19.3944
R4083 vdd.n1421 vdd.n1380 19.3944
R4084 vdd.n1417 vdd.n1380 19.3944
R4085 vdd.n1417 vdd.n1416 19.3944
R4086 vdd.n1416 vdd.n1415 19.3944
R4087 vdd.n1415 vdd.n1386 19.3944
R4088 vdd.n1411 vdd.n1386 19.3944
R4089 vdd.n1411 vdd.n1410 19.3944
R4090 vdd.n1410 vdd.n1409 19.3944
R4091 vdd.n1409 vdd.n1392 19.3944
R4092 vdd.n1405 vdd.n1392 19.3944
R4093 vdd.n1405 vdd.n1404 19.3944
R4094 vdd.n1404 vdd.n1403 19.3944
R4095 vdd.n1468 vdd.n1467 19.3944
R4096 vdd.n1467 vdd.n1466 19.3944
R4097 vdd.n1466 vdd.n1339 19.3944
R4098 vdd.n1462 vdd.n1339 19.3944
R4099 vdd.n1462 vdd.n1461 19.3944
R4100 vdd.n1461 vdd.n1460 19.3944
R4101 vdd.n1460 vdd.n1345 19.3944
R4102 vdd.n1456 vdd.n1345 19.3944
R4103 vdd.n1456 vdd.n1455 19.3944
R4104 vdd.n1455 vdd.n1454 19.3944
R4105 vdd.n1454 vdd.n1351 19.3944
R4106 vdd.n1450 vdd.n1351 19.3944
R4107 vdd.n1450 vdd.n1449 19.3944
R4108 vdd.n1449 vdd.n1448 19.3944
R4109 vdd.n1448 vdd.n1357 19.3944
R4110 vdd.n1444 vdd.n1357 19.3944
R4111 vdd.n1444 vdd.n1443 19.3944
R4112 vdd.n1443 vdd.n1442 19.3944
R4113 vdd.n1442 vdd.n1363 19.3944
R4114 vdd.n1438 vdd.n1363 19.3944
R4115 vdd.n1501 vdd.n1272 19.3944
R4116 vdd.n1496 vdd.n1272 19.3944
R4117 vdd.n1496 vdd.n1307 19.3944
R4118 vdd.n1492 vdd.n1307 19.3944
R4119 vdd.n1492 vdd.n1491 19.3944
R4120 vdd.n1491 vdd.n1490 19.3944
R4121 vdd.n1490 vdd.n1313 19.3944
R4122 vdd.n1486 vdd.n1313 19.3944
R4123 vdd.n1486 vdd.n1485 19.3944
R4124 vdd.n1485 vdd.n1484 19.3944
R4125 vdd.n1484 vdd.n1319 19.3944
R4126 vdd.n1480 vdd.n1319 19.3944
R4127 vdd.n1480 vdd.n1479 19.3944
R4128 vdd.n1479 vdd.n1478 19.3944
R4129 vdd.n1478 vdd.n1325 19.3944
R4130 vdd.n1474 vdd.n1325 19.3944
R4131 vdd.n1474 vdd.n1473 19.3944
R4132 vdd.n1473 vdd.n1472 19.3944
R4133 vdd.n2114 vdd.n2049 19.3944
R4134 vdd.n2114 vdd.n2055 19.3944
R4135 vdd.n2109 vdd.n2055 19.3944
R4136 vdd.n2109 vdd.n2108 19.3944
R4137 vdd.n2108 vdd.n2107 19.3944
R4138 vdd.n2107 vdd.n2062 19.3944
R4139 vdd.n2102 vdd.n2062 19.3944
R4140 vdd.n2102 vdd.n2101 19.3944
R4141 vdd.n2101 vdd.n2100 19.3944
R4142 vdd.n2100 vdd.n2069 19.3944
R4143 vdd.n2095 vdd.n2069 19.3944
R4144 vdd.n2095 vdd.n2094 19.3944
R4145 vdd.n2094 vdd.n2093 19.3944
R4146 vdd.n2093 vdd.n2077 19.3944
R4147 vdd.n2088 vdd.n2077 19.3944
R4148 vdd.n2088 vdd.n2087 19.3944
R4149 vdd.n2083 vdd.n2082 19.3944
R4150 vdd.n2203 vdd.n1148 19.3944
R4151 vdd.n2153 vdd.n2009 19.3944
R4152 vdd.n2153 vdd.n2015 19.3944
R4153 vdd.n2148 vdd.n2015 19.3944
R4154 vdd.n2148 vdd.n2147 19.3944
R4155 vdd.n2147 vdd.n2146 19.3944
R4156 vdd.n2146 vdd.n2022 19.3944
R4157 vdd.n2141 vdd.n2022 19.3944
R4158 vdd.n2141 vdd.n2140 19.3944
R4159 vdd.n2140 vdd.n2139 19.3944
R4160 vdd.n2139 vdd.n2029 19.3944
R4161 vdd.n2134 vdd.n2029 19.3944
R4162 vdd.n2134 vdd.n2133 19.3944
R4163 vdd.n2133 vdd.n2132 19.3944
R4164 vdd.n2132 vdd.n2036 19.3944
R4165 vdd.n2127 vdd.n2036 19.3944
R4166 vdd.n2127 vdd.n2126 19.3944
R4167 vdd.n2126 vdd.n2125 19.3944
R4168 vdd.n2125 vdd.n2043 19.3944
R4169 vdd.n2120 vdd.n2043 19.3944
R4170 vdd.n2120 vdd.n2119 19.3944
R4171 vdd.n2191 vdd.n2190 19.3944
R4172 vdd.n2190 vdd.n1981 19.3944
R4173 vdd.n2185 vdd.n2184 19.3944
R4174 vdd.n2180 vdd.n1985 19.3944
R4175 vdd.n2180 vdd.n1987 19.3944
R4176 vdd.n1990 vdd.n1987 19.3944
R4177 vdd.n2173 vdd.n1990 19.3944
R4178 vdd.n2173 vdd.n2172 19.3944
R4179 vdd.n2172 vdd.n2171 19.3944
R4180 vdd.n2171 vdd.n1996 19.3944
R4181 vdd.n2166 vdd.n1996 19.3944
R4182 vdd.n2166 vdd.n2165 19.3944
R4183 vdd.n2165 vdd.n2164 19.3944
R4184 vdd.n2164 vdd.n2003 19.3944
R4185 vdd.n2159 vdd.n2003 19.3944
R4186 vdd.n2159 vdd.n2158 19.3944
R4187 vdd.n1505 vdd.n1270 19.3944
R4188 vdd.n1505 vdd.n1261 19.3944
R4189 vdd.n1518 vdd.n1261 19.3944
R4190 vdd.n1518 vdd.n1259 19.3944
R4191 vdd.n1522 vdd.n1259 19.3944
R4192 vdd.n1522 vdd.n1250 19.3944
R4193 vdd.n1535 vdd.n1250 19.3944
R4194 vdd.n1535 vdd.n1248 19.3944
R4195 vdd.n1539 vdd.n1248 19.3944
R4196 vdd.n1539 vdd.n1239 19.3944
R4197 vdd.n1551 vdd.n1239 19.3944
R4198 vdd.n1551 vdd.n1237 19.3944
R4199 vdd.n1555 vdd.n1237 19.3944
R4200 vdd.n1555 vdd.n1227 19.3944
R4201 vdd.n1568 vdd.n1227 19.3944
R4202 vdd.n1568 vdd.n1225 19.3944
R4203 vdd.n1572 vdd.n1225 19.3944
R4204 vdd.n1572 vdd.n1216 19.3944
R4205 vdd.n1584 vdd.n1216 19.3944
R4206 vdd.n1584 vdd.n1214 19.3944
R4207 vdd.n1895 vdd.n1214 19.3944
R4208 vdd.n1895 vdd.n1204 19.3944
R4209 vdd.n1908 vdd.n1204 19.3944
R4210 vdd.n1908 vdd.n1202 19.3944
R4211 vdd.n1912 vdd.n1202 19.3944
R4212 vdd.n1912 vdd.n1193 19.3944
R4213 vdd.n1925 vdd.n1193 19.3944
R4214 vdd.n1925 vdd.n1191 19.3944
R4215 vdd.n1929 vdd.n1191 19.3944
R4216 vdd.n1929 vdd.n1182 19.3944
R4217 vdd.n1941 vdd.n1182 19.3944
R4218 vdd.n1941 vdd.n1180 19.3944
R4219 vdd.n1945 vdd.n1180 19.3944
R4220 vdd.n1945 vdd.n1170 19.3944
R4221 vdd.n1958 vdd.n1170 19.3944
R4222 vdd.n1958 vdd.n1168 19.3944
R4223 vdd.n1962 vdd.n1168 19.3944
R4224 vdd.n1962 vdd.n1158 19.3944
R4225 vdd.n1977 vdd.n1158 19.3944
R4226 vdd.n1977 vdd.n1156 19.3944
R4227 vdd.n2194 vdd.n1156 19.3944
R4228 vdd.n3411 vdd.n686 19.3944
R4229 vdd.n3411 vdd.n676 19.3944
R4230 vdd.n3423 vdd.n676 19.3944
R4231 vdd.n3423 vdd.n674 19.3944
R4232 vdd.n3427 vdd.n674 19.3944
R4233 vdd.n3427 vdd.n666 19.3944
R4234 vdd.n3440 vdd.n666 19.3944
R4235 vdd.n3440 vdd.n664 19.3944
R4236 vdd.n3444 vdd.n664 19.3944
R4237 vdd.n3444 vdd.n653 19.3944
R4238 vdd.n3456 vdd.n653 19.3944
R4239 vdd.n3456 vdd.n651 19.3944
R4240 vdd.n3460 vdd.n651 19.3944
R4241 vdd.n3460 vdd.n642 19.3944
R4242 vdd.n3473 vdd.n642 19.3944
R4243 vdd.n3473 vdd.n640 19.3944
R4244 vdd.n3480 vdd.n640 19.3944
R4245 vdd.n3480 vdd.n3479 19.3944
R4246 vdd.n3479 vdd.n631 19.3944
R4247 vdd.n3493 vdd.n631 19.3944
R4248 vdd.n3494 vdd.n3493 19.3944
R4249 vdd.n3494 vdd.n629 19.3944
R4250 vdd.n3498 vdd.n629 19.3944
R4251 vdd.n3500 vdd.n3498 19.3944
R4252 vdd.n3501 vdd.n3500 19.3944
R4253 vdd.n3501 vdd.n627 19.3944
R4254 vdd.n3505 vdd.n627 19.3944
R4255 vdd.n3507 vdd.n3505 19.3944
R4256 vdd.n3508 vdd.n3507 19.3944
R4257 vdd.n3508 vdd.n625 19.3944
R4258 vdd.n3512 vdd.n625 19.3944
R4259 vdd.n3515 vdd.n3512 19.3944
R4260 vdd.n3516 vdd.n3515 19.3944
R4261 vdd.n3516 vdd.n623 19.3944
R4262 vdd.n3520 vdd.n623 19.3944
R4263 vdd.n3522 vdd.n3520 19.3944
R4264 vdd.n3523 vdd.n3522 19.3944
R4265 vdd.n3523 vdd.n621 19.3944
R4266 vdd.n3527 vdd.n621 19.3944
R4267 vdd.n3529 vdd.n3527 19.3944
R4268 vdd.n3530 vdd.n3529 19.3944
R4269 vdd.n569 vdd.n438 19.3944
R4270 vdd.n575 vdd.n438 19.3944
R4271 vdd.n576 vdd.n575 19.3944
R4272 vdd.n579 vdd.n576 19.3944
R4273 vdd.n579 vdd.n436 19.3944
R4274 vdd.n585 vdd.n436 19.3944
R4275 vdd.n586 vdd.n585 19.3944
R4276 vdd.n589 vdd.n586 19.3944
R4277 vdd.n589 vdd.n434 19.3944
R4278 vdd.n595 vdd.n434 19.3944
R4279 vdd.n596 vdd.n595 19.3944
R4280 vdd.n599 vdd.n596 19.3944
R4281 vdd.n599 vdd.n432 19.3944
R4282 vdd.n605 vdd.n432 19.3944
R4283 vdd.n606 vdd.n605 19.3944
R4284 vdd.n609 vdd.n606 19.3944
R4285 vdd.n609 vdd.n430 19.3944
R4286 vdd.n615 vdd.n430 19.3944
R4287 vdd.n617 vdd.n615 19.3944
R4288 vdd.n618 vdd.n617 19.3944
R4289 vdd.n516 vdd.n515 19.3944
R4290 vdd.n519 vdd.n516 19.3944
R4291 vdd.n519 vdd.n450 19.3944
R4292 vdd.n525 vdd.n450 19.3944
R4293 vdd.n526 vdd.n525 19.3944
R4294 vdd.n529 vdd.n526 19.3944
R4295 vdd.n529 vdd.n448 19.3944
R4296 vdd.n535 vdd.n448 19.3944
R4297 vdd.n536 vdd.n535 19.3944
R4298 vdd.n539 vdd.n536 19.3944
R4299 vdd.n539 vdd.n446 19.3944
R4300 vdd.n545 vdd.n446 19.3944
R4301 vdd.n546 vdd.n545 19.3944
R4302 vdd.n549 vdd.n546 19.3944
R4303 vdd.n549 vdd.n444 19.3944
R4304 vdd.n555 vdd.n444 19.3944
R4305 vdd.n556 vdd.n555 19.3944
R4306 vdd.n559 vdd.n556 19.3944
R4307 vdd.n559 vdd.n442 19.3944
R4308 vdd.n565 vdd.n442 19.3944
R4309 vdd.n466 vdd.n465 19.3944
R4310 vdd.n469 vdd.n466 19.3944
R4311 vdd.n469 vdd.n462 19.3944
R4312 vdd.n475 vdd.n462 19.3944
R4313 vdd.n476 vdd.n475 19.3944
R4314 vdd.n479 vdd.n476 19.3944
R4315 vdd.n479 vdd.n460 19.3944
R4316 vdd.n485 vdd.n460 19.3944
R4317 vdd.n486 vdd.n485 19.3944
R4318 vdd.n489 vdd.n486 19.3944
R4319 vdd.n489 vdd.n458 19.3944
R4320 vdd.n495 vdd.n458 19.3944
R4321 vdd.n496 vdd.n495 19.3944
R4322 vdd.n499 vdd.n496 19.3944
R4323 vdd.n499 vdd.n456 19.3944
R4324 vdd.n505 vdd.n456 19.3944
R4325 vdd.n506 vdd.n505 19.3944
R4326 vdd.n509 vdd.n506 19.3944
R4327 vdd.n3415 vdd.n683 19.3944
R4328 vdd.n3415 vdd.n681 19.3944
R4329 vdd.n3419 vdd.n681 19.3944
R4330 vdd.n3419 vdd.n671 19.3944
R4331 vdd.n3432 vdd.n671 19.3944
R4332 vdd.n3432 vdd.n669 19.3944
R4333 vdd.n3436 vdd.n669 19.3944
R4334 vdd.n3436 vdd.n660 19.3944
R4335 vdd.n3448 vdd.n660 19.3944
R4336 vdd.n3448 vdd.n658 19.3944
R4337 vdd.n3452 vdd.n658 19.3944
R4338 vdd.n3452 vdd.n648 19.3944
R4339 vdd.n3465 vdd.n648 19.3944
R4340 vdd.n3465 vdd.n646 19.3944
R4341 vdd.n3469 vdd.n646 19.3944
R4342 vdd.n3469 vdd.n637 19.3944
R4343 vdd.n3484 vdd.n637 19.3944
R4344 vdd.n3484 vdd.n635 19.3944
R4345 vdd.n3488 vdd.n635 19.3944
R4346 vdd.n3488 vdd.n336 19.3944
R4347 vdd.n3579 vdd.n336 19.3944
R4348 vdd.n3579 vdd.n337 19.3944
R4349 vdd.n3573 vdd.n337 19.3944
R4350 vdd.n3573 vdd.n3572 19.3944
R4351 vdd.n3572 vdd.n3571 19.3944
R4352 vdd.n3571 vdd.n349 19.3944
R4353 vdd.n3565 vdd.n349 19.3944
R4354 vdd.n3565 vdd.n3564 19.3944
R4355 vdd.n3564 vdd.n3563 19.3944
R4356 vdd.n3563 vdd.n359 19.3944
R4357 vdd.n3557 vdd.n359 19.3944
R4358 vdd.n3557 vdd.n3556 19.3944
R4359 vdd.n3556 vdd.n3555 19.3944
R4360 vdd.n3555 vdd.n370 19.3944
R4361 vdd.n3549 vdd.n370 19.3944
R4362 vdd.n3549 vdd.n3548 19.3944
R4363 vdd.n3548 vdd.n3547 19.3944
R4364 vdd.n3547 vdd.n381 19.3944
R4365 vdd.n3541 vdd.n381 19.3944
R4366 vdd.n3541 vdd.n3540 19.3944
R4367 vdd.n3540 vdd.n3539 19.3944
R4368 vdd.n3362 vdd.n747 19.3944
R4369 vdd.n3362 vdd.n3359 19.3944
R4370 vdd.n3359 vdd.n3356 19.3944
R4371 vdd.n3356 vdd.n3355 19.3944
R4372 vdd.n3355 vdd.n3352 19.3944
R4373 vdd.n3352 vdd.n3351 19.3944
R4374 vdd.n3351 vdd.n3348 19.3944
R4375 vdd.n3348 vdd.n3347 19.3944
R4376 vdd.n3347 vdd.n3344 19.3944
R4377 vdd.n3344 vdd.n3343 19.3944
R4378 vdd.n3343 vdd.n3340 19.3944
R4379 vdd.n3340 vdd.n3339 19.3944
R4380 vdd.n3339 vdd.n3336 19.3944
R4381 vdd.n3336 vdd.n3335 19.3944
R4382 vdd.n3335 vdd.n3332 19.3944
R4383 vdd.n3332 vdd.n3331 19.3944
R4384 vdd.n3331 vdd.n3328 19.3944
R4385 vdd.n3328 vdd.n3327 19.3944
R4386 vdd.n3327 vdd.n3324 19.3944
R4387 vdd.n3324 vdd.n3323 19.3944
R4388 vdd.n3402 vdd.n3401 19.3944
R4389 vdd.n3401 vdd.n3400 19.3944
R4390 vdd.n732 vdd.n729 19.3944
R4391 vdd.n3396 vdd.n3395 19.3944
R4392 vdd.n3395 vdd.n3392 19.3944
R4393 vdd.n3392 vdd.n3391 19.3944
R4394 vdd.n3391 vdd.n3388 19.3944
R4395 vdd.n3388 vdd.n3387 19.3944
R4396 vdd.n3387 vdd.n3384 19.3944
R4397 vdd.n3384 vdd.n3383 19.3944
R4398 vdd.n3383 vdd.n3380 19.3944
R4399 vdd.n3380 vdd.n3379 19.3944
R4400 vdd.n3379 vdd.n3376 19.3944
R4401 vdd.n3376 vdd.n3375 19.3944
R4402 vdd.n3375 vdd.n3372 19.3944
R4403 vdd.n3372 vdd.n3371 19.3944
R4404 vdd.n3316 vdd.n767 19.3944
R4405 vdd.n3316 vdd.n3313 19.3944
R4406 vdd.n3313 vdd.n3310 19.3944
R4407 vdd.n3310 vdd.n3309 19.3944
R4408 vdd.n3309 vdd.n3306 19.3944
R4409 vdd.n3306 vdd.n3305 19.3944
R4410 vdd.n3305 vdd.n3302 19.3944
R4411 vdd.n3302 vdd.n3301 19.3944
R4412 vdd.n3301 vdd.n3298 19.3944
R4413 vdd.n3298 vdd.n3297 19.3944
R4414 vdd.n3297 vdd.n3294 19.3944
R4415 vdd.n3294 vdd.n3293 19.3944
R4416 vdd.n3293 vdd.n3290 19.3944
R4417 vdd.n3290 vdd.n3289 19.3944
R4418 vdd.n3289 vdd.n3286 19.3944
R4419 vdd.n3286 vdd.n3285 19.3944
R4420 vdd.n3282 vdd.n3281 19.3944
R4421 vdd.n3278 vdd.n3277 19.3944
R4422 vdd.n1437 vdd.n1433 19.0066
R4423 vdd.n2118 vdd.n2049 19.0066
R4424 vdd.n569 vdd.n566 19.0066
R4425 vdd.n3320 vdd.n767 19.0066
R4426 vdd.n1137 vdd.n1136 16.0975
R4427 vdd.n998 vdd.n997 16.0975
R4428 vdd.n1398 vdd.n1397 16.0975
R4429 vdd.n1436 vdd.n1435 16.0975
R4430 vdd.n1332 vdd.n1331 16.0975
R4431 vdd.n2201 vdd.n2200 16.0975
R4432 vdd.n2051 vdd.n2050 16.0975
R4433 vdd.n2011 vdd.n2010 16.0975
R4434 vdd.n1131 vdd.n1130 16.0975
R4435 vdd.n989 vdd.n988 16.0975
R4436 vdd.n2762 vdd.n2761 16.0975
R4437 vdd.n427 vdd.n426 16.0975
R4438 vdd.n441 vdd.n440 16.0975
R4439 vdd.n453 vdd.n452 16.0975
R4440 vdd.n769 vdd.n768 16.0975
R4441 vdd.n3367 vdd.n3366 16.0975
R4442 vdd.n833 vdd.n832 16.0975
R4443 vdd.n2831 vdd.n2830 16.0975
R4444 vdd.n689 vdd.n688 16.0975
R4445 vdd.n800 vdd.n799 16.0975
R4446 vdd.t10 vdd.n2726 15.4182
R4447 vdd.n3010 vdd.t0 15.4182
R4448 vdd.n28 vdd.n27 14.5035
R4449 vdd.n2467 vdd.n1110 13.6043
R4450 vdd.n3241 vdd.n692 13.6043
R4451 vdd.n328 vdd.n293 13.1884
R4452 vdd.n269 vdd.n234 13.1884
R4453 vdd.n226 vdd.n191 13.1884
R4454 vdd.n167 vdd.n132 13.1884
R4455 vdd.n125 vdd.n90 13.1884
R4456 vdd.n66 vdd.n31 13.1884
R4457 vdd.n1827 vdd.n1792 13.1884
R4458 vdd.n1886 vdd.n1851 13.1884
R4459 vdd.n1725 vdd.n1690 13.1884
R4460 vdd.n1784 vdd.n1749 13.1884
R4461 vdd.n1624 vdd.n1589 13.1884
R4462 vdd.n1683 vdd.n1648 13.1884
R4463 vdd.n1468 vdd.n1333 12.9944
R4464 vdd.n1472 vdd.n1333 12.9944
R4465 vdd.n2157 vdd.n2009 12.9944
R4466 vdd.n2158 vdd.n2157 12.9944
R4467 vdd.n515 vdd.n454 12.9944
R4468 vdd.n509 vdd.n454 12.9944
R4469 vdd.n3368 vdd.n747 12.9944
R4470 vdd.n3371 vdd.n3368 12.9944
R4471 vdd.n329 vdd.n291 12.8005
R4472 vdd.n324 vdd.n295 12.8005
R4473 vdd.n270 vdd.n232 12.8005
R4474 vdd.n265 vdd.n236 12.8005
R4475 vdd.n227 vdd.n189 12.8005
R4476 vdd.n222 vdd.n193 12.8005
R4477 vdd.n168 vdd.n130 12.8005
R4478 vdd.n163 vdd.n134 12.8005
R4479 vdd.n126 vdd.n88 12.8005
R4480 vdd.n121 vdd.n92 12.8005
R4481 vdd.n67 vdd.n29 12.8005
R4482 vdd.n62 vdd.n33 12.8005
R4483 vdd.n1828 vdd.n1790 12.8005
R4484 vdd.n1823 vdd.n1794 12.8005
R4485 vdd.n1887 vdd.n1849 12.8005
R4486 vdd.n1882 vdd.n1853 12.8005
R4487 vdd.n1726 vdd.n1688 12.8005
R4488 vdd.n1721 vdd.n1692 12.8005
R4489 vdd.n1785 vdd.n1747 12.8005
R4490 vdd.n1780 vdd.n1751 12.8005
R4491 vdd.n1625 vdd.n1587 12.8005
R4492 vdd.n1620 vdd.n1591 12.8005
R4493 vdd.n1684 vdd.n1646 12.8005
R4494 vdd.n1679 vdd.n1650 12.8005
R4495 vdd.n323 vdd.n296 12.0247
R4496 vdd.n264 vdd.n237 12.0247
R4497 vdd.n221 vdd.n194 12.0247
R4498 vdd.n162 vdd.n135 12.0247
R4499 vdd.n120 vdd.n93 12.0247
R4500 vdd.n61 vdd.n34 12.0247
R4501 vdd.n1822 vdd.n1795 12.0247
R4502 vdd.n1881 vdd.n1854 12.0247
R4503 vdd.n1720 vdd.n1693 12.0247
R4504 vdd.n1779 vdd.n1752 12.0247
R4505 vdd.n1619 vdd.n1592 12.0247
R4506 vdd.n1678 vdd.n1651 12.0247
R4507 vdd.n1507 vdd.n1263 11.337
R4508 vdd.n1516 vdd.n1263 11.337
R4509 vdd.n1516 vdd.n1515 11.337
R4510 vdd.n1524 vdd.n1257 11.337
R4511 vdd.n1533 vdd.n1532 11.337
R4512 vdd.n1549 vdd.n1241 11.337
R4513 vdd.n1557 vdd.n1234 11.337
R4514 vdd.n1566 vdd.n1565 11.337
R4515 vdd.n1574 vdd.n1223 11.337
R4516 vdd.n1897 vdd.n1212 11.337
R4517 vdd.n1906 vdd.n1206 11.337
R4518 vdd.n1914 vdd.n1200 11.337
R4519 vdd.n1923 vdd.n1922 11.337
R4520 vdd.n1939 vdd.n1184 11.337
R4521 vdd.n1947 vdd.n1177 11.337
R4522 vdd.n1956 vdd.n1955 11.337
R4523 vdd.n1964 vdd.n1160 11.337
R4524 vdd.n1975 vdd.n1160 11.337
R4525 vdd.n1975 vdd.n1974 11.337
R4526 vdd.n3413 vdd.n678 11.337
R4527 vdd.n3421 vdd.n678 11.337
R4528 vdd.n3421 vdd.n679 11.337
R4529 vdd.n3430 vdd.n3429 11.337
R4530 vdd.n3446 vdd.n662 11.337
R4531 vdd.n3454 vdd.n655 11.337
R4532 vdd.n3463 vdd.n3462 11.337
R4533 vdd.n3471 vdd.n644 11.337
R4534 vdd.n3490 vdd.n633 11.337
R4535 vdd.n3577 vdd.n340 11.337
R4536 vdd.n3575 vdd.n344 11.337
R4537 vdd.n3569 vdd.n3568 11.337
R4538 vdd.n3561 vdd.n361 11.337
R4539 vdd.n3560 vdd.n3559 11.337
R4540 vdd.n3553 vdd.n3552 11.337
R4541 vdd.n3551 vdd.n375 11.337
R4542 vdd.n3545 vdd.n3544 11.337
R4543 vdd.n3544 vdd.n3543 11.337
R4544 vdd.n3543 vdd.n386 11.337
R4545 vdd.n320 vdd.n319 11.249
R4546 vdd.n261 vdd.n260 11.249
R4547 vdd.n218 vdd.n217 11.249
R4548 vdd.n159 vdd.n158 11.249
R4549 vdd.n117 vdd.n116 11.249
R4550 vdd.n58 vdd.n57 11.249
R4551 vdd.n1819 vdd.n1818 11.249
R4552 vdd.n1878 vdd.n1877 11.249
R4553 vdd.n1717 vdd.n1716 11.249
R4554 vdd.n1776 vdd.n1775 11.249
R4555 vdd.n1616 vdd.n1615 11.249
R4556 vdd.n1675 vdd.n1674 11.249
R4557 vdd.n1305 vdd.t106 11.2237
R4558 vdd.n3537 vdd.t76 11.2237
R4559 vdd.t202 vdd.n1178 10.7702
R4560 vdd.n3438 vdd.t185 10.7702
R4561 vdd.n305 vdd.n304 10.7238
R4562 vdd.n246 vdd.n245 10.7238
R4563 vdd.n203 vdd.n202 10.7238
R4564 vdd.n144 vdd.n143 10.7238
R4565 vdd.n102 vdd.n101 10.7238
R4566 vdd.n43 vdd.n42 10.7238
R4567 vdd.n1804 vdd.n1803 10.7238
R4568 vdd.n1863 vdd.n1862 10.7238
R4569 vdd.n1702 vdd.n1701 10.7238
R4570 vdd.n1761 vdd.n1760 10.7238
R4571 vdd.n1601 vdd.n1600 10.7238
R4572 vdd.n1660 vdd.n1659 10.7238
R4573 vdd.n2465 vdd.n1102 10.6151
R4574 vdd.n2475 vdd.n1102 10.6151
R4575 vdd.n2476 vdd.n2475 10.6151
R4576 vdd.n2477 vdd.n2476 10.6151
R4577 vdd.n2477 vdd.n1090 10.6151
R4578 vdd.n2487 vdd.n1090 10.6151
R4579 vdd.n2488 vdd.n2487 10.6151
R4580 vdd.n2489 vdd.n2488 10.6151
R4581 vdd.n2489 vdd.n1078 10.6151
R4582 vdd.n2499 vdd.n1078 10.6151
R4583 vdd.n2500 vdd.n2499 10.6151
R4584 vdd.n2501 vdd.n2500 10.6151
R4585 vdd.n2501 vdd.n1065 10.6151
R4586 vdd.n2511 vdd.n1065 10.6151
R4587 vdd.n2512 vdd.n2511 10.6151
R4588 vdd.n2513 vdd.n2512 10.6151
R4589 vdd.n2513 vdd.n1053 10.6151
R4590 vdd.n2524 vdd.n1053 10.6151
R4591 vdd.n2525 vdd.n2524 10.6151
R4592 vdd.n2526 vdd.n2525 10.6151
R4593 vdd.n2526 vdd.n1041 10.6151
R4594 vdd.n2536 vdd.n1041 10.6151
R4595 vdd.n2537 vdd.n2536 10.6151
R4596 vdd.n2538 vdd.n2537 10.6151
R4597 vdd.n2538 vdd.n1029 10.6151
R4598 vdd.n2548 vdd.n1029 10.6151
R4599 vdd.n2549 vdd.n2548 10.6151
R4600 vdd.n2550 vdd.n2549 10.6151
R4601 vdd.n2550 vdd.n1019 10.6151
R4602 vdd.n2560 vdd.n1019 10.6151
R4603 vdd.n2561 vdd.n2560 10.6151
R4604 vdd.n2562 vdd.n2561 10.6151
R4605 vdd.n2562 vdd.n1006 10.6151
R4606 vdd.n2574 vdd.n1006 10.6151
R4607 vdd.n2575 vdd.n2574 10.6151
R4608 vdd.n2577 vdd.n2575 10.6151
R4609 vdd.n2577 vdd.n2576 10.6151
R4610 vdd.n2576 vdd.n987 10.6151
R4611 vdd.n2724 vdd.n2723 10.6151
R4612 vdd.n2723 vdd.n2722 10.6151
R4613 vdd.n2722 vdd.n2719 10.6151
R4614 vdd.n2719 vdd.n2718 10.6151
R4615 vdd.n2718 vdd.n2715 10.6151
R4616 vdd.n2715 vdd.n2714 10.6151
R4617 vdd.n2714 vdd.n2711 10.6151
R4618 vdd.n2711 vdd.n2710 10.6151
R4619 vdd.n2710 vdd.n2707 10.6151
R4620 vdd.n2707 vdd.n2706 10.6151
R4621 vdd.n2706 vdd.n2703 10.6151
R4622 vdd.n2703 vdd.n2702 10.6151
R4623 vdd.n2702 vdd.n2699 10.6151
R4624 vdd.n2699 vdd.n2698 10.6151
R4625 vdd.n2698 vdd.n2695 10.6151
R4626 vdd.n2695 vdd.n2694 10.6151
R4627 vdd.n2694 vdd.n2691 10.6151
R4628 vdd.n2691 vdd.n2690 10.6151
R4629 vdd.n2690 vdd.n2687 10.6151
R4630 vdd.n2687 vdd.n2686 10.6151
R4631 vdd.n2686 vdd.n2683 10.6151
R4632 vdd.n2683 vdd.n2682 10.6151
R4633 vdd.n2682 vdd.n2679 10.6151
R4634 vdd.n2679 vdd.n2678 10.6151
R4635 vdd.n2678 vdd.n2675 10.6151
R4636 vdd.n2675 vdd.n2674 10.6151
R4637 vdd.n2674 vdd.n2671 10.6151
R4638 vdd.n2671 vdd.n2670 10.6151
R4639 vdd.n2670 vdd.n2667 10.6151
R4640 vdd.n2667 vdd.n2666 10.6151
R4641 vdd.n2666 vdd.n2663 10.6151
R4642 vdd.n2661 vdd.n2658 10.6151
R4643 vdd.n2658 vdd.n2657 10.6151
R4644 vdd.n2394 vdd.n2393 10.6151
R4645 vdd.n2393 vdd.n2391 10.6151
R4646 vdd.n2391 vdd.n2390 10.6151
R4647 vdd.n2390 vdd.n2388 10.6151
R4648 vdd.n2388 vdd.n2387 10.6151
R4649 vdd.n2387 vdd.n2385 10.6151
R4650 vdd.n2385 vdd.n2384 10.6151
R4651 vdd.n2384 vdd.n2382 10.6151
R4652 vdd.n2382 vdd.n2381 10.6151
R4653 vdd.n2381 vdd.n2379 10.6151
R4654 vdd.n2379 vdd.n2378 10.6151
R4655 vdd.n2378 vdd.n2376 10.6151
R4656 vdd.n2376 vdd.n2375 10.6151
R4657 vdd.n2375 vdd.n2373 10.6151
R4658 vdd.n2373 vdd.n2372 10.6151
R4659 vdd.n2372 vdd.n2370 10.6151
R4660 vdd.n2370 vdd.n2369 10.6151
R4661 vdd.n2369 vdd.n2367 10.6151
R4662 vdd.n2367 vdd.n2366 10.6151
R4663 vdd.n2366 vdd.n2364 10.6151
R4664 vdd.n2364 vdd.n2363 10.6151
R4665 vdd.n2363 vdd.n2361 10.6151
R4666 vdd.n2361 vdd.n2360 10.6151
R4667 vdd.n2360 vdd.n1133 10.6151
R4668 vdd.n2327 vdd.n1133 10.6151
R4669 vdd.n2328 vdd.n2327 10.6151
R4670 vdd.n2330 vdd.n2328 10.6151
R4671 vdd.n2331 vdd.n2330 10.6151
R4672 vdd.n2344 vdd.n2331 10.6151
R4673 vdd.n2344 vdd.n2343 10.6151
R4674 vdd.n2343 vdd.n2342 10.6151
R4675 vdd.n2342 vdd.n2340 10.6151
R4676 vdd.n2340 vdd.n2339 10.6151
R4677 vdd.n2339 vdd.n2337 10.6151
R4678 vdd.n2337 vdd.n2336 10.6151
R4679 vdd.n2336 vdd.n2333 10.6151
R4680 vdd.n2333 vdd.n2332 10.6151
R4681 vdd.n2332 vdd.n990 10.6151
R4682 vdd.n2464 vdd.n2463 10.6151
R4683 vdd.n2463 vdd.n1114 10.6151
R4684 vdd.n2458 vdd.n1114 10.6151
R4685 vdd.n2458 vdd.n2457 10.6151
R4686 vdd.n2457 vdd.n1116 10.6151
R4687 vdd.n2452 vdd.n1116 10.6151
R4688 vdd.n2452 vdd.n2451 10.6151
R4689 vdd.n2451 vdd.n2450 10.6151
R4690 vdd.n2450 vdd.n1118 10.6151
R4691 vdd.n2444 vdd.n1118 10.6151
R4692 vdd.n2444 vdd.n2443 10.6151
R4693 vdd.n2443 vdd.n2442 10.6151
R4694 vdd.n2442 vdd.n1120 10.6151
R4695 vdd.n2436 vdd.n1120 10.6151
R4696 vdd.n2436 vdd.n2435 10.6151
R4697 vdd.n2435 vdd.n2434 10.6151
R4698 vdd.n2434 vdd.n1122 10.6151
R4699 vdd.n2428 vdd.n1122 10.6151
R4700 vdd.n2428 vdd.n2427 10.6151
R4701 vdd.n2427 vdd.n2426 10.6151
R4702 vdd.n2426 vdd.n1124 10.6151
R4703 vdd.n2420 vdd.n1124 10.6151
R4704 vdd.n2420 vdd.n2419 10.6151
R4705 vdd.n2419 vdd.n2418 10.6151
R4706 vdd.n2418 vdd.n1126 10.6151
R4707 vdd.n2412 vdd.n1126 10.6151
R4708 vdd.n2412 vdd.n2411 10.6151
R4709 vdd.n2411 vdd.n2410 10.6151
R4710 vdd.n2410 vdd.n1128 10.6151
R4711 vdd.n2404 vdd.n1128 10.6151
R4712 vdd.n2404 vdd.n2403 10.6151
R4713 vdd.n2401 vdd.n1132 10.6151
R4714 vdd.n2395 vdd.n1132 10.6151
R4715 vdd.n2899 vdd.n2897 10.6151
R4716 vdd.n2900 vdd.n2899 10.6151
R4717 vdd.n2999 vdd.n2900 10.6151
R4718 vdd.n2999 vdd.n2998 10.6151
R4719 vdd.n2998 vdd.n2997 10.6151
R4720 vdd.n2997 vdd.n2995 10.6151
R4721 vdd.n2995 vdd.n2994 10.6151
R4722 vdd.n2994 vdd.n2992 10.6151
R4723 vdd.n2992 vdd.n2991 10.6151
R4724 vdd.n2991 vdd.n2901 10.6151
R4725 vdd.n2941 vdd.n2901 10.6151
R4726 vdd.n2942 vdd.n2941 10.6151
R4727 vdd.n2944 vdd.n2942 10.6151
R4728 vdd.n2945 vdd.n2944 10.6151
R4729 vdd.n2975 vdd.n2945 10.6151
R4730 vdd.n2975 vdd.n2974 10.6151
R4731 vdd.n2974 vdd.n2973 10.6151
R4732 vdd.n2973 vdd.n2971 10.6151
R4733 vdd.n2971 vdd.n2970 10.6151
R4734 vdd.n2970 vdd.n2968 10.6151
R4735 vdd.n2968 vdd.n2967 10.6151
R4736 vdd.n2967 vdd.n2965 10.6151
R4737 vdd.n2965 vdd.n2964 10.6151
R4738 vdd.n2964 vdd.n2962 10.6151
R4739 vdd.n2962 vdd.n2961 10.6151
R4740 vdd.n2961 vdd.n2959 10.6151
R4741 vdd.n2959 vdd.n2958 10.6151
R4742 vdd.n2958 vdd.n2956 10.6151
R4743 vdd.n2956 vdd.n2955 10.6151
R4744 vdd.n2955 vdd.n2953 10.6151
R4745 vdd.n2953 vdd.n2952 10.6151
R4746 vdd.n2952 vdd.n2950 10.6151
R4747 vdd.n2950 vdd.n2949 10.6151
R4748 vdd.n2949 vdd.n2947 10.6151
R4749 vdd.n2947 vdd.n2946 10.6151
R4750 vdd.n2946 vdd.n836 10.6151
R4751 vdd.n3174 vdd.n836 10.6151
R4752 vdd.n3175 vdd.n3174 10.6151
R4753 vdd.n3014 vdd.n3013 10.6151
R4754 vdd.n3013 vdd.n948 10.6151
R4755 vdd.n2833 vdd.n948 10.6151
R4756 vdd.n2834 vdd.n2833 10.6151
R4757 vdd.n2837 vdd.n2834 10.6151
R4758 vdd.n2838 vdd.n2837 10.6151
R4759 vdd.n2841 vdd.n2838 10.6151
R4760 vdd.n2842 vdd.n2841 10.6151
R4761 vdd.n2845 vdd.n2842 10.6151
R4762 vdd.n2846 vdd.n2845 10.6151
R4763 vdd.n2849 vdd.n2846 10.6151
R4764 vdd.n2850 vdd.n2849 10.6151
R4765 vdd.n2853 vdd.n2850 10.6151
R4766 vdd.n2854 vdd.n2853 10.6151
R4767 vdd.n2857 vdd.n2854 10.6151
R4768 vdd.n2858 vdd.n2857 10.6151
R4769 vdd.n2861 vdd.n2858 10.6151
R4770 vdd.n2862 vdd.n2861 10.6151
R4771 vdd.n2865 vdd.n2862 10.6151
R4772 vdd.n2866 vdd.n2865 10.6151
R4773 vdd.n2869 vdd.n2866 10.6151
R4774 vdd.n2870 vdd.n2869 10.6151
R4775 vdd.n2873 vdd.n2870 10.6151
R4776 vdd.n2874 vdd.n2873 10.6151
R4777 vdd.n2877 vdd.n2874 10.6151
R4778 vdd.n2878 vdd.n2877 10.6151
R4779 vdd.n2881 vdd.n2878 10.6151
R4780 vdd.n2882 vdd.n2881 10.6151
R4781 vdd.n2885 vdd.n2882 10.6151
R4782 vdd.n2886 vdd.n2885 10.6151
R4783 vdd.n2889 vdd.n2886 10.6151
R4784 vdd.n2894 vdd.n2891 10.6151
R4785 vdd.n2896 vdd.n2894 10.6151
R4786 vdd.n3015 vdd.n937 10.6151
R4787 vdd.n3025 vdd.n937 10.6151
R4788 vdd.n3026 vdd.n3025 10.6151
R4789 vdd.n3027 vdd.n3026 10.6151
R4790 vdd.n3027 vdd.n925 10.6151
R4791 vdd.n3037 vdd.n925 10.6151
R4792 vdd.n3038 vdd.n3037 10.6151
R4793 vdd.n3039 vdd.n3038 10.6151
R4794 vdd.n3039 vdd.n915 10.6151
R4795 vdd.n3049 vdd.n915 10.6151
R4796 vdd.n3050 vdd.n3049 10.6151
R4797 vdd.n3051 vdd.n3050 10.6151
R4798 vdd.n3051 vdd.n903 10.6151
R4799 vdd.n3061 vdd.n903 10.6151
R4800 vdd.n3062 vdd.n3061 10.6151
R4801 vdd.n3063 vdd.n3062 10.6151
R4802 vdd.n3063 vdd.n892 10.6151
R4803 vdd.n3073 vdd.n892 10.6151
R4804 vdd.n3074 vdd.n3073 10.6151
R4805 vdd.n3075 vdd.n3074 10.6151
R4806 vdd.n3075 vdd.n879 10.6151
R4807 vdd.n3086 vdd.n879 10.6151
R4808 vdd.n3087 vdd.n3086 10.6151
R4809 vdd.n3088 vdd.n3087 10.6151
R4810 vdd.n3088 vdd.n866 10.6151
R4811 vdd.n3098 vdd.n866 10.6151
R4812 vdd.n3099 vdd.n3098 10.6151
R4813 vdd.n3100 vdd.n3099 10.6151
R4814 vdd.n3100 vdd.n855 10.6151
R4815 vdd.n3110 vdd.n855 10.6151
R4816 vdd.n3111 vdd.n3110 10.6151
R4817 vdd.n3112 vdd.n3111 10.6151
R4818 vdd.n3112 vdd.n841 10.6151
R4819 vdd.n3167 vdd.n841 10.6151
R4820 vdd.n3168 vdd.n3167 10.6151
R4821 vdd.n3169 vdd.n3168 10.6151
R4822 vdd.n3169 vdd.n810 10.6151
R4823 vdd.n3239 vdd.n810 10.6151
R4824 vdd.n3238 vdd.n3237 10.6151
R4825 vdd.n3237 vdd.n811 10.6151
R4826 vdd.n812 vdd.n811 10.6151
R4827 vdd.n3230 vdd.n812 10.6151
R4828 vdd.n3230 vdd.n3229 10.6151
R4829 vdd.n3229 vdd.n3228 10.6151
R4830 vdd.n3228 vdd.n814 10.6151
R4831 vdd.n3223 vdd.n814 10.6151
R4832 vdd.n3223 vdd.n3222 10.6151
R4833 vdd.n3222 vdd.n3221 10.6151
R4834 vdd.n3221 vdd.n817 10.6151
R4835 vdd.n3216 vdd.n817 10.6151
R4836 vdd.n3216 vdd.n3215 10.6151
R4837 vdd.n3215 vdd.n3214 10.6151
R4838 vdd.n3214 vdd.n820 10.6151
R4839 vdd.n3209 vdd.n820 10.6151
R4840 vdd.n3209 vdd.n731 10.6151
R4841 vdd.n3205 vdd.n731 10.6151
R4842 vdd.n3205 vdd.n3204 10.6151
R4843 vdd.n3204 vdd.n3203 10.6151
R4844 vdd.n3203 vdd.n823 10.6151
R4845 vdd.n3198 vdd.n823 10.6151
R4846 vdd.n3198 vdd.n3197 10.6151
R4847 vdd.n3197 vdd.n3196 10.6151
R4848 vdd.n3196 vdd.n826 10.6151
R4849 vdd.n3191 vdd.n826 10.6151
R4850 vdd.n3191 vdd.n3190 10.6151
R4851 vdd.n3190 vdd.n3189 10.6151
R4852 vdd.n3189 vdd.n829 10.6151
R4853 vdd.n3184 vdd.n829 10.6151
R4854 vdd.n3184 vdd.n3183 10.6151
R4855 vdd.n3181 vdd.n834 10.6151
R4856 vdd.n3176 vdd.n834 10.6151
R4857 vdd.n3157 vdd.n3118 10.6151
R4858 vdd.n3152 vdd.n3118 10.6151
R4859 vdd.n3152 vdd.n3151 10.6151
R4860 vdd.n3151 vdd.n3150 10.6151
R4861 vdd.n3150 vdd.n3120 10.6151
R4862 vdd.n3145 vdd.n3120 10.6151
R4863 vdd.n3145 vdd.n3144 10.6151
R4864 vdd.n3144 vdd.n3143 10.6151
R4865 vdd.n3143 vdd.n3123 10.6151
R4866 vdd.n3138 vdd.n3123 10.6151
R4867 vdd.n3138 vdd.n3137 10.6151
R4868 vdd.n3137 vdd.n3136 10.6151
R4869 vdd.n3136 vdd.n3126 10.6151
R4870 vdd.n3131 vdd.n3126 10.6151
R4871 vdd.n3131 vdd.n3130 10.6151
R4872 vdd.n3130 vdd.n785 10.6151
R4873 vdd.n3274 vdd.n785 10.6151
R4874 vdd.n3274 vdd.n786 10.6151
R4875 vdd.n788 vdd.n786 10.6151
R4876 vdd.n3267 vdd.n788 10.6151
R4877 vdd.n3267 vdd.n3266 10.6151
R4878 vdd.n3266 vdd.n3265 10.6151
R4879 vdd.n3265 vdd.n790 10.6151
R4880 vdd.n3260 vdd.n790 10.6151
R4881 vdd.n3260 vdd.n3259 10.6151
R4882 vdd.n3259 vdd.n3258 10.6151
R4883 vdd.n3258 vdd.n793 10.6151
R4884 vdd.n3253 vdd.n793 10.6151
R4885 vdd.n3253 vdd.n3252 10.6151
R4886 vdd.n3252 vdd.n3251 10.6151
R4887 vdd.n3251 vdd.n796 10.6151
R4888 vdd.n3246 vdd.n3245 10.6151
R4889 vdd.n3245 vdd.n3244 10.6151
R4890 vdd.n3007 vdd.n3006 10.6151
R4891 vdd.n3006 vdd.n3004 10.6151
R4892 vdd.n3004 vdd.n3003 10.6151
R4893 vdd.n3003 vdd.n2829 10.6151
R4894 vdd.n2903 vdd.n2829 10.6151
R4895 vdd.n2904 vdd.n2903 10.6151
R4896 vdd.n2906 vdd.n2904 10.6151
R4897 vdd.n2907 vdd.n2906 10.6151
R4898 vdd.n2987 vdd.n2907 10.6151
R4899 vdd.n2987 vdd.n2986 10.6151
R4900 vdd.n2986 vdd.n2985 10.6151
R4901 vdd.n2985 vdd.n2983 10.6151
R4902 vdd.n2983 vdd.n2982 10.6151
R4903 vdd.n2982 vdd.n2980 10.6151
R4904 vdd.n2980 vdd.n2979 10.6151
R4905 vdd.n2979 vdd.n2939 10.6151
R4906 vdd.n2939 vdd.n2938 10.6151
R4907 vdd.n2938 vdd.n2936 10.6151
R4908 vdd.n2936 vdd.n2935 10.6151
R4909 vdd.n2935 vdd.n2933 10.6151
R4910 vdd.n2933 vdd.n2932 10.6151
R4911 vdd.n2932 vdd.n2930 10.6151
R4912 vdd.n2930 vdd.n2929 10.6151
R4913 vdd.n2929 vdd.n2927 10.6151
R4914 vdd.n2927 vdd.n2926 10.6151
R4915 vdd.n2926 vdd.n2924 10.6151
R4916 vdd.n2924 vdd.n2923 10.6151
R4917 vdd.n2923 vdd.n2921 10.6151
R4918 vdd.n2921 vdd.n2920 10.6151
R4919 vdd.n2920 vdd.n2918 10.6151
R4920 vdd.n2918 vdd.n2917 10.6151
R4921 vdd.n2917 vdd.n2915 10.6151
R4922 vdd.n2915 vdd.n2914 10.6151
R4923 vdd.n2914 vdd.n2912 10.6151
R4924 vdd.n2912 vdd.n2911 10.6151
R4925 vdd.n2911 vdd.n2909 10.6151
R4926 vdd.n2909 vdd.n2908 10.6151
R4927 vdd.n2908 vdd.n802 10.6151
R4928 vdd.n2764 vdd.n942 10.6151
R4929 vdd.n2767 vdd.n2764 10.6151
R4930 vdd.n2768 vdd.n2767 10.6151
R4931 vdd.n2771 vdd.n2768 10.6151
R4932 vdd.n2772 vdd.n2771 10.6151
R4933 vdd.n2775 vdd.n2772 10.6151
R4934 vdd.n2776 vdd.n2775 10.6151
R4935 vdd.n2779 vdd.n2776 10.6151
R4936 vdd.n2780 vdd.n2779 10.6151
R4937 vdd.n2783 vdd.n2780 10.6151
R4938 vdd.n2784 vdd.n2783 10.6151
R4939 vdd.n2787 vdd.n2784 10.6151
R4940 vdd.n2788 vdd.n2787 10.6151
R4941 vdd.n2791 vdd.n2788 10.6151
R4942 vdd.n2792 vdd.n2791 10.6151
R4943 vdd.n2795 vdd.n2792 10.6151
R4944 vdd.n2796 vdd.n2795 10.6151
R4945 vdd.n2799 vdd.n2796 10.6151
R4946 vdd.n2800 vdd.n2799 10.6151
R4947 vdd.n2803 vdd.n2800 10.6151
R4948 vdd.n2804 vdd.n2803 10.6151
R4949 vdd.n2807 vdd.n2804 10.6151
R4950 vdd.n2808 vdd.n2807 10.6151
R4951 vdd.n2811 vdd.n2808 10.6151
R4952 vdd.n2812 vdd.n2811 10.6151
R4953 vdd.n2815 vdd.n2812 10.6151
R4954 vdd.n2816 vdd.n2815 10.6151
R4955 vdd.n2819 vdd.n2816 10.6151
R4956 vdd.n2820 vdd.n2819 10.6151
R4957 vdd.n2823 vdd.n2820 10.6151
R4958 vdd.n2824 vdd.n2823 10.6151
R4959 vdd.n2828 vdd.n2827 10.6151
R4960 vdd.n3008 vdd.n2828 10.6151
R4961 vdd.n3020 vdd.n3019 10.6151
R4962 vdd.n3021 vdd.n3020 10.6151
R4963 vdd.n3021 vdd.n932 10.6151
R4964 vdd.n3031 vdd.n932 10.6151
R4965 vdd.n3032 vdd.n3031 10.6151
R4966 vdd.n3033 vdd.n3032 10.6151
R4967 vdd.n3033 vdd.n920 10.6151
R4968 vdd.n3043 vdd.n920 10.6151
R4969 vdd.n3044 vdd.n3043 10.6151
R4970 vdd.n3045 vdd.n3044 10.6151
R4971 vdd.n3045 vdd.n909 10.6151
R4972 vdd.n3055 vdd.n909 10.6151
R4973 vdd.n3056 vdd.n3055 10.6151
R4974 vdd.n3057 vdd.n3056 10.6151
R4975 vdd.n3057 vdd.n897 10.6151
R4976 vdd.n3067 vdd.n897 10.6151
R4977 vdd.n3068 vdd.n3067 10.6151
R4978 vdd.n3069 vdd.n3068 10.6151
R4979 vdd.n3069 vdd.n886 10.6151
R4980 vdd.n3079 vdd.n886 10.6151
R4981 vdd.n3082 vdd.n3081 10.6151
R4982 vdd.n3082 vdd.n872 10.6151
R4983 vdd.n3092 vdd.n872 10.6151
R4984 vdd.n3093 vdd.n3092 10.6151
R4985 vdd.n3094 vdd.n3093 10.6151
R4986 vdd.n3094 vdd.n860 10.6151
R4987 vdd.n3104 vdd.n860 10.6151
R4988 vdd.n3105 vdd.n3104 10.6151
R4989 vdd.n3106 vdd.n3105 10.6151
R4990 vdd.n3106 vdd.n849 10.6151
R4991 vdd.n3116 vdd.n849 10.6151
R4992 vdd.n3117 vdd.n3116 10.6151
R4993 vdd.n3163 vdd.n3117 10.6151
R4994 vdd.n3163 vdd.n3162 10.6151
R4995 vdd.n3162 vdd.n3161 10.6151
R4996 vdd.n3161 vdd.n3160 10.6151
R4997 vdd.n3160 vdd.n3158 10.6151
R4998 vdd.n2470 vdd.n2469 10.6151
R4999 vdd.n2471 vdd.n2470 10.6151
R5000 vdd.n2471 vdd.n1096 10.6151
R5001 vdd.n2481 vdd.n1096 10.6151
R5002 vdd.n2482 vdd.n2481 10.6151
R5003 vdd.n2483 vdd.n2482 10.6151
R5004 vdd.n2483 vdd.n1084 10.6151
R5005 vdd.n2493 vdd.n1084 10.6151
R5006 vdd.n2494 vdd.n2493 10.6151
R5007 vdd.n2495 vdd.n2494 10.6151
R5008 vdd.n2495 vdd.n1072 10.6151
R5009 vdd.n2505 vdd.n1072 10.6151
R5010 vdd.n2506 vdd.n2505 10.6151
R5011 vdd.n2507 vdd.n2506 10.6151
R5012 vdd.n2507 vdd.n1059 10.6151
R5013 vdd.n2517 vdd.n1059 10.6151
R5014 vdd.n2518 vdd.n2517 10.6151
R5015 vdd.n2520 vdd.n1047 10.6151
R5016 vdd.n2530 vdd.n1047 10.6151
R5017 vdd.n2531 vdd.n2530 10.6151
R5018 vdd.n2532 vdd.n2531 10.6151
R5019 vdd.n2532 vdd.n1035 10.6151
R5020 vdd.n2542 vdd.n1035 10.6151
R5021 vdd.n2543 vdd.n2542 10.6151
R5022 vdd.n2544 vdd.n2543 10.6151
R5023 vdd.n2544 vdd.n1024 10.6151
R5024 vdd.n2554 vdd.n1024 10.6151
R5025 vdd.n2555 vdd.n2554 10.6151
R5026 vdd.n2556 vdd.n2555 10.6151
R5027 vdd.n2556 vdd.n1013 10.6151
R5028 vdd.n2566 vdd.n1013 10.6151
R5029 vdd.n2567 vdd.n2566 10.6151
R5030 vdd.n2570 vdd.n2567 10.6151
R5031 vdd.n2570 vdd.n2569 10.6151
R5032 vdd.n2569 vdd.n2568 10.6151
R5033 vdd.n2568 vdd.n996 10.6151
R5034 vdd.n2652 vdd.n996 10.6151
R5035 vdd.n2651 vdd.n2650 10.6151
R5036 vdd.n2650 vdd.n2647 10.6151
R5037 vdd.n2647 vdd.n2646 10.6151
R5038 vdd.n2646 vdd.n2643 10.6151
R5039 vdd.n2643 vdd.n2642 10.6151
R5040 vdd.n2642 vdd.n2639 10.6151
R5041 vdd.n2639 vdd.n2638 10.6151
R5042 vdd.n2638 vdd.n2635 10.6151
R5043 vdd.n2635 vdd.n2634 10.6151
R5044 vdd.n2634 vdd.n2631 10.6151
R5045 vdd.n2631 vdd.n2630 10.6151
R5046 vdd.n2630 vdd.n2627 10.6151
R5047 vdd.n2627 vdd.n2626 10.6151
R5048 vdd.n2626 vdd.n2623 10.6151
R5049 vdd.n2623 vdd.n2622 10.6151
R5050 vdd.n2622 vdd.n2619 10.6151
R5051 vdd.n2619 vdd.n2618 10.6151
R5052 vdd.n2618 vdd.n2615 10.6151
R5053 vdd.n2615 vdd.n2614 10.6151
R5054 vdd.n2614 vdd.n2611 10.6151
R5055 vdd.n2611 vdd.n2610 10.6151
R5056 vdd.n2610 vdd.n2607 10.6151
R5057 vdd.n2607 vdd.n2606 10.6151
R5058 vdd.n2606 vdd.n2603 10.6151
R5059 vdd.n2603 vdd.n2602 10.6151
R5060 vdd.n2602 vdd.n2599 10.6151
R5061 vdd.n2599 vdd.n2598 10.6151
R5062 vdd.n2598 vdd.n2595 10.6151
R5063 vdd.n2595 vdd.n2594 10.6151
R5064 vdd.n2594 vdd.n2591 10.6151
R5065 vdd.n2591 vdd.n2590 10.6151
R5066 vdd.n2587 vdd.n2586 10.6151
R5067 vdd.n2586 vdd.n2584 10.6151
R5068 vdd.n2286 vdd.n2284 10.6151
R5069 vdd.n2287 vdd.n2286 10.6151
R5070 vdd.n2289 vdd.n2287 10.6151
R5071 vdd.n2290 vdd.n2289 10.6151
R5072 vdd.n2292 vdd.n2290 10.6151
R5073 vdd.n2293 vdd.n2292 10.6151
R5074 vdd.n2295 vdd.n2293 10.6151
R5075 vdd.n2296 vdd.n2295 10.6151
R5076 vdd.n2298 vdd.n2296 10.6151
R5077 vdd.n2299 vdd.n2298 10.6151
R5078 vdd.n2301 vdd.n2299 10.6151
R5079 vdd.n2302 vdd.n2301 10.6151
R5080 vdd.n2304 vdd.n2302 10.6151
R5081 vdd.n2305 vdd.n2304 10.6151
R5082 vdd.n2307 vdd.n2305 10.6151
R5083 vdd.n2308 vdd.n2307 10.6151
R5084 vdd.n2310 vdd.n2308 10.6151
R5085 vdd.n2311 vdd.n2310 10.6151
R5086 vdd.n2313 vdd.n2311 10.6151
R5087 vdd.n2314 vdd.n2313 10.6151
R5088 vdd.n2316 vdd.n2314 10.6151
R5089 vdd.n2317 vdd.n2316 10.6151
R5090 vdd.n2356 vdd.n2317 10.6151
R5091 vdd.n2356 vdd.n2355 10.6151
R5092 vdd.n2355 vdd.n2354 10.6151
R5093 vdd.n2354 vdd.n2352 10.6151
R5094 vdd.n2352 vdd.n2351 10.6151
R5095 vdd.n2351 vdd.n2349 10.6151
R5096 vdd.n2349 vdd.n2348 10.6151
R5097 vdd.n2348 vdd.n2325 10.6151
R5098 vdd.n2325 vdd.n2324 10.6151
R5099 vdd.n2324 vdd.n2322 10.6151
R5100 vdd.n2322 vdd.n2321 10.6151
R5101 vdd.n2321 vdd.n2319 10.6151
R5102 vdd.n2319 vdd.n2318 10.6151
R5103 vdd.n2318 vdd.n1000 10.6151
R5104 vdd.n2582 vdd.n1000 10.6151
R5105 vdd.n2583 vdd.n2582 10.6151
R5106 vdd.n2214 vdd.n1108 10.6151
R5107 vdd.n2219 vdd.n2214 10.6151
R5108 vdd.n2220 vdd.n2219 10.6151
R5109 vdd.n2221 vdd.n2220 10.6151
R5110 vdd.n2221 vdd.n2212 10.6151
R5111 vdd.n2227 vdd.n2212 10.6151
R5112 vdd.n2228 vdd.n2227 10.6151
R5113 vdd.n2229 vdd.n2228 10.6151
R5114 vdd.n2229 vdd.n2210 10.6151
R5115 vdd.n2235 vdd.n2210 10.6151
R5116 vdd.n2236 vdd.n2235 10.6151
R5117 vdd.n2237 vdd.n2236 10.6151
R5118 vdd.n2237 vdd.n2208 10.6151
R5119 vdd.n2243 vdd.n2208 10.6151
R5120 vdd.n2244 vdd.n2243 10.6151
R5121 vdd.n2245 vdd.n2244 10.6151
R5122 vdd.n2245 vdd.n2206 10.6151
R5123 vdd.n2251 vdd.n2206 10.6151
R5124 vdd.n2252 vdd.n2251 10.6151
R5125 vdd.n2253 vdd.n2252 10.6151
R5126 vdd.n2253 vdd.n1142 10.6151
R5127 vdd.n2259 vdd.n1142 10.6151
R5128 vdd.n2260 vdd.n2259 10.6151
R5129 vdd.n2261 vdd.n2260 10.6151
R5130 vdd.n2261 vdd.n1140 10.6151
R5131 vdd.n2267 vdd.n1140 10.6151
R5132 vdd.n2268 vdd.n2267 10.6151
R5133 vdd.n2269 vdd.n2268 10.6151
R5134 vdd.n2269 vdd.n1138 10.6151
R5135 vdd.n2275 vdd.n1138 10.6151
R5136 vdd.n2276 vdd.n2275 10.6151
R5137 vdd.n2278 vdd.n1134 10.6151
R5138 vdd.n2283 vdd.n1134 10.6151
R5139 vdd.n1931 vdd.t232 10.5435
R5140 vdd.n656 vdd.t190 10.5435
R5141 vdd.n316 vdd.n298 10.4732
R5142 vdd.n257 vdd.n239 10.4732
R5143 vdd.n214 vdd.n196 10.4732
R5144 vdd.n155 vdd.n137 10.4732
R5145 vdd.n113 vdd.n95 10.4732
R5146 vdd.n54 vdd.n36 10.4732
R5147 vdd.n1815 vdd.n1797 10.4732
R5148 vdd.n1874 vdd.n1856 10.4732
R5149 vdd.n1713 vdd.n1695 10.4732
R5150 vdd.n1772 vdd.n1754 10.4732
R5151 vdd.n1612 vdd.n1594 10.4732
R5152 vdd.n1671 vdd.n1653 10.4732
R5153 vdd.t175 vdd.n1905 10.3167
R5154 vdd.n3482 vdd.t254 10.3167
R5155 vdd.n2654 vdd.t39 10.2034
R5156 vdd.n3017 vdd.t31 10.2034
R5157 vdd.n1582 vdd.t148 10.09
R5158 vdd.n3576 vdd.t208 10.09
R5159 vdd.n2182 vdd.n1122 9.88581
R5160 vdd.n3398 vdd.n731 9.88581
R5161 vdd.n3275 vdd.n3274 9.88581
R5162 vdd.n2206 vdd.n2205 9.88581
R5163 vdd.t139 vdd.n1235 9.86327
R5164 vdd.n3567 vdd.t258 9.86327
R5165 vdd.n315 vdd.n300 9.69747
R5166 vdd.n256 vdd.n241 9.69747
R5167 vdd.n213 vdd.n198 9.69747
R5168 vdd.n154 vdd.n139 9.69747
R5169 vdd.n112 vdd.n97 9.69747
R5170 vdd.n53 vdd.n38 9.69747
R5171 vdd.n1814 vdd.n1799 9.69747
R5172 vdd.n1873 vdd.n1858 9.69747
R5173 vdd.n1712 vdd.n1697 9.69747
R5174 vdd.n1771 vdd.n1756 9.69747
R5175 vdd.n1611 vdd.n1596 9.69747
R5176 vdd.n1670 vdd.n1655 9.69747
R5177 vdd.n1541 vdd.t220 9.63654
R5178 vdd.n3513 vdd.t217 9.63654
R5179 vdd.n331 vdd.n330 9.45567
R5180 vdd.n272 vdd.n271 9.45567
R5181 vdd.n229 vdd.n228 9.45567
R5182 vdd.n170 vdd.n169 9.45567
R5183 vdd.n128 vdd.n127 9.45567
R5184 vdd.n69 vdd.n68 9.45567
R5185 vdd.n1830 vdd.n1829 9.45567
R5186 vdd.n1889 vdd.n1888 9.45567
R5187 vdd.n1728 vdd.n1727 9.45567
R5188 vdd.n1787 vdd.n1786 9.45567
R5189 vdd.n1627 vdd.n1626 9.45567
R5190 vdd.n1686 vdd.n1685 9.45567
R5191 vdd.n1515 vdd.t234 9.40981
R5192 vdd.n3545 vdd.t141 9.40981
R5193 vdd.n2155 vdd.n2009 9.3005
R5194 vdd.n2154 vdd.n2153 9.3005
R5195 vdd.n2015 vdd.n2014 9.3005
R5196 vdd.n2148 vdd.n2019 9.3005
R5197 vdd.n2147 vdd.n2020 9.3005
R5198 vdd.n2146 vdd.n2021 9.3005
R5199 vdd.n2025 vdd.n2022 9.3005
R5200 vdd.n2141 vdd.n2026 9.3005
R5201 vdd.n2140 vdd.n2027 9.3005
R5202 vdd.n2139 vdd.n2028 9.3005
R5203 vdd.n2032 vdd.n2029 9.3005
R5204 vdd.n2134 vdd.n2033 9.3005
R5205 vdd.n2133 vdd.n2034 9.3005
R5206 vdd.n2132 vdd.n2035 9.3005
R5207 vdd.n2039 vdd.n2036 9.3005
R5208 vdd.n2127 vdd.n2040 9.3005
R5209 vdd.n2126 vdd.n2041 9.3005
R5210 vdd.n2125 vdd.n2042 9.3005
R5211 vdd.n2046 vdd.n2043 9.3005
R5212 vdd.n2120 vdd.n2047 9.3005
R5213 vdd.n2119 vdd.n2048 9.3005
R5214 vdd.n2118 vdd.n2117 9.3005
R5215 vdd.n2116 vdd.n2049 9.3005
R5216 vdd.n2115 vdd.n2114 9.3005
R5217 vdd.n2055 vdd.n2054 9.3005
R5218 vdd.n2109 vdd.n2059 9.3005
R5219 vdd.n2108 vdd.n2060 9.3005
R5220 vdd.n2107 vdd.n2061 9.3005
R5221 vdd.n2065 vdd.n2062 9.3005
R5222 vdd.n2102 vdd.n2066 9.3005
R5223 vdd.n2101 vdd.n2067 9.3005
R5224 vdd.n2100 vdd.n2068 9.3005
R5225 vdd.n2072 vdd.n2069 9.3005
R5226 vdd.n2095 vdd.n2073 9.3005
R5227 vdd.n2094 vdd.n2074 9.3005
R5228 vdd.n2093 vdd.n2075 9.3005
R5229 vdd.n2077 vdd.n2076 9.3005
R5230 vdd.n2088 vdd.n1144 9.3005
R5231 vdd.n2157 vdd.n2156 9.3005
R5232 vdd.n2181 vdd.n2180 9.3005
R5233 vdd.n1987 vdd.n1986 9.3005
R5234 vdd.n1992 vdd.n1990 9.3005
R5235 vdd.n2173 vdd.n1993 9.3005
R5236 vdd.n2172 vdd.n1994 9.3005
R5237 vdd.n2171 vdd.n1995 9.3005
R5238 vdd.n1999 vdd.n1996 9.3005
R5239 vdd.n2166 vdd.n2000 9.3005
R5240 vdd.n2165 vdd.n2001 9.3005
R5241 vdd.n2164 vdd.n2002 9.3005
R5242 vdd.n2006 vdd.n2003 9.3005
R5243 vdd.n2159 vdd.n2007 9.3005
R5244 vdd.n2158 vdd.n2008 9.3005
R5245 vdd.n2190 vdd.n1980 9.3005
R5246 vdd.n2192 vdd.n2191 9.3005
R5247 vdd.n1895 vdd.n1894 9.3005
R5248 vdd.n1204 vdd.n1203 9.3005
R5249 vdd.n1909 vdd.n1908 9.3005
R5250 vdd.n1910 vdd.n1202 9.3005
R5251 vdd.n1912 vdd.n1911 9.3005
R5252 vdd.n1193 vdd.n1192 9.3005
R5253 vdd.n1926 vdd.n1925 9.3005
R5254 vdd.n1927 vdd.n1191 9.3005
R5255 vdd.n1929 vdd.n1928 9.3005
R5256 vdd.n1182 vdd.n1181 9.3005
R5257 vdd.n1942 vdd.n1941 9.3005
R5258 vdd.n1943 vdd.n1180 9.3005
R5259 vdd.n1945 vdd.n1944 9.3005
R5260 vdd.n1170 vdd.n1169 9.3005
R5261 vdd.n1959 vdd.n1958 9.3005
R5262 vdd.n1960 vdd.n1168 9.3005
R5263 vdd.n1962 vdd.n1961 9.3005
R5264 vdd.n1158 vdd.n1157 9.3005
R5265 vdd.n1978 vdd.n1977 9.3005
R5266 vdd.n1979 vdd.n1156 9.3005
R5267 vdd.n2194 vdd.n2193 9.3005
R5268 vdd.n307 vdd.n306 9.3005
R5269 vdd.n302 vdd.n301 9.3005
R5270 vdd.n313 vdd.n312 9.3005
R5271 vdd.n315 vdd.n314 9.3005
R5272 vdd.n298 vdd.n297 9.3005
R5273 vdd.n321 vdd.n320 9.3005
R5274 vdd.n323 vdd.n322 9.3005
R5275 vdd.n295 vdd.n292 9.3005
R5276 vdd.n330 vdd.n329 9.3005
R5277 vdd.n248 vdd.n247 9.3005
R5278 vdd.n243 vdd.n242 9.3005
R5279 vdd.n254 vdd.n253 9.3005
R5280 vdd.n256 vdd.n255 9.3005
R5281 vdd.n239 vdd.n238 9.3005
R5282 vdd.n262 vdd.n261 9.3005
R5283 vdd.n264 vdd.n263 9.3005
R5284 vdd.n236 vdd.n233 9.3005
R5285 vdd.n271 vdd.n270 9.3005
R5286 vdd.n205 vdd.n204 9.3005
R5287 vdd.n200 vdd.n199 9.3005
R5288 vdd.n211 vdd.n210 9.3005
R5289 vdd.n213 vdd.n212 9.3005
R5290 vdd.n196 vdd.n195 9.3005
R5291 vdd.n219 vdd.n218 9.3005
R5292 vdd.n221 vdd.n220 9.3005
R5293 vdd.n193 vdd.n190 9.3005
R5294 vdd.n228 vdd.n227 9.3005
R5295 vdd.n146 vdd.n145 9.3005
R5296 vdd.n141 vdd.n140 9.3005
R5297 vdd.n152 vdd.n151 9.3005
R5298 vdd.n154 vdd.n153 9.3005
R5299 vdd.n137 vdd.n136 9.3005
R5300 vdd.n160 vdd.n159 9.3005
R5301 vdd.n162 vdd.n161 9.3005
R5302 vdd.n134 vdd.n131 9.3005
R5303 vdd.n169 vdd.n168 9.3005
R5304 vdd.n104 vdd.n103 9.3005
R5305 vdd.n99 vdd.n98 9.3005
R5306 vdd.n110 vdd.n109 9.3005
R5307 vdd.n112 vdd.n111 9.3005
R5308 vdd.n95 vdd.n94 9.3005
R5309 vdd.n118 vdd.n117 9.3005
R5310 vdd.n120 vdd.n119 9.3005
R5311 vdd.n92 vdd.n89 9.3005
R5312 vdd.n127 vdd.n126 9.3005
R5313 vdd.n45 vdd.n44 9.3005
R5314 vdd.n40 vdd.n39 9.3005
R5315 vdd.n51 vdd.n50 9.3005
R5316 vdd.n53 vdd.n52 9.3005
R5317 vdd.n36 vdd.n35 9.3005
R5318 vdd.n59 vdd.n58 9.3005
R5319 vdd.n61 vdd.n60 9.3005
R5320 vdd.n33 vdd.n30 9.3005
R5321 vdd.n68 vdd.n67 9.3005
R5322 vdd.n3320 vdd.n3319 9.3005
R5323 vdd.n3323 vdd.n766 9.3005
R5324 vdd.n3324 vdd.n765 9.3005
R5325 vdd.n3327 vdd.n764 9.3005
R5326 vdd.n3328 vdd.n763 9.3005
R5327 vdd.n3331 vdd.n762 9.3005
R5328 vdd.n3332 vdd.n761 9.3005
R5329 vdd.n3335 vdd.n760 9.3005
R5330 vdd.n3336 vdd.n759 9.3005
R5331 vdd.n3339 vdd.n758 9.3005
R5332 vdd.n3340 vdd.n757 9.3005
R5333 vdd.n3343 vdd.n756 9.3005
R5334 vdd.n3344 vdd.n755 9.3005
R5335 vdd.n3347 vdd.n754 9.3005
R5336 vdd.n3348 vdd.n753 9.3005
R5337 vdd.n3351 vdd.n752 9.3005
R5338 vdd.n3352 vdd.n751 9.3005
R5339 vdd.n3355 vdd.n750 9.3005
R5340 vdd.n3356 vdd.n749 9.3005
R5341 vdd.n3359 vdd.n748 9.3005
R5342 vdd.n3363 vdd.n3362 9.3005
R5343 vdd.n3364 vdd.n747 9.3005
R5344 vdd.n3368 vdd.n3365 9.3005
R5345 vdd.n3371 vdd.n746 9.3005
R5346 vdd.n3372 vdd.n745 9.3005
R5347 vdd.n3375 vdd.n744 9.3005
R5348 vdd.n3376 vdd.n743 9.3005
R5349 vdd.n3379 vdd.n742 9.3005
R5350 vdd.n3380 vdd.n741 9.3005
R5351 vdd.n3383 vdd.n740 9.3005
R5352 vdd.n3384 vdd.n739 9.3005
R5353 vdd.n3387 vdd.n738 9.3005
R5354 vdd.n3388 vdd.n737 9.3005
R5355 vdd.n3391 vdd.n736 9.3005
R5356 vdd.n3392 vdd.n735 9.3005
R5357 vdd.n3395 vdd.n730 9.3005
R5358 vdd.n3401 vdd.n727 9.3005
R5359 vdd.n3402 vdd.n726 9.3005
R5360 vdd.n3416 vdd.n3415 9.3005
R5361 vdd.n3417 vdd.n681 9.3005
R5362 vdd.n3419 vdd.n3418 9.3005
R5363 vdd.n671 vdd.n670 9.3005
R5364 vdd.n3433 vdd.n3432 9.3005
R5365 vdd.n3434 vdd.n669 9.3005
R5366 vdd.n3436 vdd.n3435 9.3005
R5367 vdd.n660 vdd.n659 9.3005
R5368 vdd.n3449 vdd.n3448 9.3005
R5369 vdd.n3450 vdd.n658 9.3005
R5370 vdd.n3452 vdd.n3451 9.3005
R5371 vdd.n648 vdd.n647 9.3005
R5372 vdd.n3466 vdd.n3465 9.3005
R5373 vdd.n3467 vdd.n646 9.3005
R5374 vdd.n3469 vdd.n3468 9.3005
R5375 vdd.n637 vdd.n636 9.3005
R5376 vdd.n3485 vdd.n3484 9.3005
R5377 vdd.n3486 vdd.n635 9.3005
R5378 vdd.n3488 vdd.n3487 9.3005
R5379 vdd.n336 vdd.n334 9.3005
R5380 vdd.n683 vdd.n682 9.3005
R5381 vdd.n3580 vdd.n3579 9.3005
R5382 vdd.n337 vdd.n335 9.3005
R5383 vdd.n3573 vdd.n346 9.3005
R5384 vdd.n3572 vdd.n347 9.3005
R5385 vdd.n3571 vdd.n348 9.3005
R5386 vdd.n355 vdd.n349 9.3005
R5387 vdd.n3565 vdd.n356 9.3005
R5388 vdd.n3564 vdd.n357 9.3005
R5389 vdd.n3563 vdd.n358 9.3005
R5390 vdd.n366 vdd.n359 9.3005
R5391 vdd.n3557 vdd.n367 9.3005
R5392 vdd.n3556 vdd.n368 9.3005
R5393 vdd.n3555 vdd.n369 9.3005
R5394 vdd.n377 vdd.n370 9.3005
R5395 vdd.n3549 vdd.n378 9.3005
R5396 vdd.n3548 vdd.n379 9.3005
R5397 vdd.n3547 vdd.n380 9.3005
R5398 vdd.n388 vdd.n381 9.3005
R5399 vdd.n3541 vdd.n389 9.3005
R5400 vdd.n3540 vdd.n390 9.3005
R5401 vdd.n3539 vdd.n391 9.3005
R5402 vdd.n466 vdd.n463 9.3005
R5403 vdd.n470 vdd.n469 9.3005
R5404 vdd.n471 vdd.n462 9.3005
R5405 vdd.n475 vdd.n472 9.3005
R5406 vdd.n476 vdd.n461 9.3005
R5407 vdd.n480 vdd.n479 9.3005
R5408 vdd.n481 vdd.n460 9.3005
R5409 vdd.n485 vdd.n482 9.3005
R5410 vdd.n486 vdd.n459 9.3005
R5411 vdd.n490 vdd.n489 9.3005
R5412 vdd.n491 vdd.n458 9.3005
R5413 vdd.n495 vdd.n492 9.3005
R5414 vdd.n496 vdd.n457 9.3005
R5415 vdd.n500 vdd.n499 9.3005
R5416 vdd.n501 vdd.n456 9.3005
R5417 vdd.n505 vdd.n502 9.3005
R5418 vdd.n506 vdd.n455 9.3005
R5419 vdd.n510 vdd.n509 9.3005
R5420 vdd.n511 vdd.n454 9.3005
R5421 vdd.n515 vdd.n512 9.3005
R5422 vdd.n516 vdd.n451 9.3005
R5423 vdd.n520 vdd.n519 9.3005
R5424 vdd.n521 vdd.n450 9.3005
R5425 vdd.n525 vdd.n522 9.3005
R5426 vdd.n526 vdd.n449 9.3005
R5427 vdd.n530 vdd.n529 9.3005
R5428 vdd.n531 vdd.n448 9.3005
R5429 vdd.n535 vdd.n532 9.3005
R5430 vdd.n536 vdd.n447 9.3005
R5431 vdd.n540 vdd.n539 9.3005
R5432 vdd.n541 vdd.n446 9.3005
R5433 vdd.n545 vdd.n542 9.3005
R5434 vdd.n546 vdd.n445 9.3005
R5435 vdd.n550 vdd.n549 9.3005
R5436 vdd.n551 vdd.n444 9.3005
R5437 vdd.n555 vdd.n552 9.3005
R5438 vdd.n556 vdd.n443 9.3005
R5439 vdd.n560 vdd.n559 9.3005
R5440 vdd.n561 vdd.n442 9.3005
R5441 vdd.n565 vdd.n562 9.3005
R5442 vdd.n566 vdd.n439 9.3005
R5443 vdd.n570 vdd.n569 9.3005
R5444 vdd.n571 vdd.n438 9.3005
R5445 vdd.n575 vdd.n572 9.3005
R5446 vdd.n576 vdd.n437 9.3005
R5447 vdd.n580 vdd.n579 9.3005
R5448 vdd.n581 vdd.n436 9.3005
R5449 vdd.n585 vdd.n582 9.3005
R5450 vdd.n586 vdd.n435 9.3005
R5451 vdd.n590 vdd.n589 9.3005
R5452 vdd.n591 vdd.n434 9.3005
R5453 vdd.n595 vdd.n592 9.3005
R5454 vdd.n596 vdd.n433 9.3005
R5455 vdd.n600 vdd.n599 9.3005
R5456 vdd.n601 vdd.n432 9.3005
R5457 vdd.n605 vdd.n602 9.3005
R5458 vdd.n606 vdd.n431 9.3005
R5459 vdd.n610 vdd.n609 9.3005
R5460 vdd.n611 vdd.n430 9.3005
R5461 vdd.n615 vdd.n612 9.3005
R5462 vdd.n617 vdd.n429 9.3005
R5463 vdd.n619 vdd.n618 9.3005
R5464 vdd.n3533 vdd.n3532 9.3005
R5465 vdd.n465 vdd.n464 9.3005
R5466 vdd.n3411 vdd.n3410 9.3005
R5467 vdd.n676 vdd.n675 9.3005
R5468 vdd.n3424 vdd.n3423 9.3005
R5469 vdd.n3425 vdd.n674 9.3005
R5470 vdd.n3427 vdd.n3426 9.3005
R5471 vdd.n666 vdd.n665 9.3005
R5472 vdd.n3441 vdd.n3440 9.3005
R5473 vdd.n3442 vdd.n664 9.3005
R5474 vdd.n3444 vdd.n3443 9.3005
R5475 vdd.n653 vdd.n652 9.3005
R5476 vdd.n3457 vdd.n3456 9.3005
R5477 vdd.n3458 vdd.n651 9.3005
R5478 vdd.n3460 vdd.n3459 9.3005
R5479 vdd.n642 vdd.n641 9.3005
R5480 vdd.n3474 vdd.n3473 9.3005
R5481 vdd.n3475 vdd.n640 9.3005
R5482 vdd.n3480 vdd.n3476 9.3005
R5483 vdd.n3479 vdd.n3478 9.3005
R5484 vdd.n3477 vdd.n631 9.3005
R5485 vdd.n3493 vdd.n630 9.3005
R5486 vdd.n3495 vdd.n3494 9.3005
R5487 vdd.n3496 vdd.n629 9.3005
R5488 vdd.n3498 vdd.n3497 9.3005
R5489 vdd.n3500 vdd.n628 9.3005
R5490 vdd.n3502 vdd.n3501 9.3005
R5491 vdd.n3503 vdd.n627 9.3005
R5492 vdd.n3505 vdd.n3504 9.3005
R5493 vdd.n3507 vdd.n626 9.3005
R5494 vdd.n3509 vdd.n3508 9.3005
R5495 vdd.n3510 vdd.n625 9.3005
R5496 vdd.n3512 vdd.n3511 9.3005
R5497 vdd.n3515 vdd.n624 9.3005
R5498 vdd.n3517 vdd.n3516 9.3005
R5499 vdd.n3518 vdd.n623 9.3005
R5500 vdd.n3520 vdd.n3519 9.3005
R5501 vdd.n3522 vdd.n622 9.3005
R5502 vdd.n3524 vdd.n3523 9.3005
R5503 vdd.n3525 vdd.n621 9.3005
R5504 vdd.n3527 vdd.n3526 9.3005
R5505 vdd.n3529 vdd.n620 9.3005
R5506 vdd.n3531 vdd.n3530 9.3005
R5507 vdd.n3409 vdd.n686 9.3005
R5508 vdd.n3408 vdd.n3407 9.3005
R5509 vdd.n3277 vdd.n687 9.3005
R5510 vdd.n3286 vdd.n783 9.3005
R5511 vdd.n3289 vdd.n782 9.3005
R5512 vdd.n3290 vdd.n781 9.3005
R5513 vdd.n3293 vdd.n780 9.3005
R5514 vdd.n3294 vdd.n779 9.3005
R5515 vdd.n3297 vdd.n778 9.3005
R5516 vdd.n3298 vdd.n777 9.3005
R5517 vdd.n3301 vdd.n776 9.3005
R5518 vdd.n3302 vdd.n775 9.3005
R5519 vdd.n3305 vdd.n774 9.3005
R5520 vdd.n3306 vdd.n773 9.3005
R5521 vdd.n3309 vdd.n772 9.3005
R5522 vdd.n3310 vdd.n771 9.3005
R5523 vdd.n3313 vdd.n770 9.3005
R5524 vdd.n3317 vdd.n3316 9.3005
R5525 vdd.n3318 vdd.n767 9.3005
R5526 vdd.n2204 vdd.n2203 9.3005
R5527 vdd.n2199 vdd.n1147 9.3005
R5528 vdd.n1510 vdd.n1509 9.3005
R5529 vdd.n1511 vdd.n1265 9.3005
R5530 vdd.n1513 vdd.n1512 9.3005
R5531 vdd.n1255 vdd.n1254 9.3005
R5532 vdd.n1527 vdd.n1526 9.3005
R5533 vdd.n1528 vdd.n1253 9.3005
R5534 vdd.n1530 vdd.n1529 9.3005
R5535 vdd.n1245 vdd.n1244 9.3005
R5536 vdd.n1544 vdd.n1543 9.3005
R5537 vdd.n1545 vdd.n1243 9.3005
R5538 vdd.n1547 vdd.n1546 9.3005
R5539 vdd.n1232 vdd.n1231 9.3005
R5540 vdd.n1560 vdd.n1559 9.3005
R5541 vdd.n1561 vdd.n1230 9.3005
R5542 vdd.n1563 vdd.n1562 9.3005
R5543 vdd.n1221 vdd.n1220 9.3005
R5544 vdd.n1577 vdd.n1576 9.3005
R5545 vdd.n1578 vdd.n1219 9.3005
R5546 vdd.n1580 vdd.n1579 9.3005
R5547 vdd.n1210 vdd.n1209 9.3005
R5548 vdd.n1900 vdd.n1899 9.3005
R5549 vdd.n1901 vdd.n1208 9.3005
R5550 vdd.n1903 vdd.n1902 9.3005
R5551 vdd.n1198 vdd.n1197 9.3005
R5552 vdd.n1917 vdd.n1916 9.3005
R5553 vdd.n1918 vdd.n1196 9.3005
R5554 vdd.n1920 vdd.n1919 9.3005
R5555 vdd.n1188 vdd.n1187 9.3005
R5556 vdd.n1934 vdd.n1933 9.3005
R5557 vdd.n1935 vdd.n1186 9.3005
R5558 vdd.n1937 vdd.n1936 9.3005
R5559 vdd.n1175 vdd.n1174 9.3005
R5560 vdd.n1950 vdd.n1949 9.3005
R5561 vdd.n1951 vdd.n1173 9.3005
R5562 vdd.n1953 vdd.n1952 9.3005
R5563 vdd.n1165 vdd.n1164 9.3005
R5564 vdd.n1967 vdd.n1966 9.3005
R5565 vdd.n1968 vdd.n1162 9.3005
R5566 vdd.n1972 vdd.n1971 9.3005
R5567 vdd.n1970 vdd.n1163 9.3005
R5568 vdd.n1969 vdd.n1152 9.3005
R5569 vdd.n1267 vdd.n1266 9.3005
R5570 vdd.n1403 vdd.n1402 9.3005
R5571 vdd.n1404 vdd.n1393 9.3005
R5572 vdd.n1406 vdd.n1405 9.3005
R5573 vdd.n1407 vdd.n1392 9.3005
R5574 vdd.n1409 vdd.n1408 9.3005
R5575 vdd.n1410 vdd.n1387 9.3005
R5576 vdd.n1412 vdd.n1411 9.3005
R5577 vdd.n1413 vdd.n1386 9.3005
R5578 vdd.n1415 vdd.n1414 9.3005
R5579 vdd.n1416 vdd.n1381 9.3005
R5580 vdd.n1418 vdd.n1417 9.3005
R5581 vdd.n1419 vdd.n1380 9.3005
R5582 vdd.n1421 vdd.n1420 9.3005
R5583 vdd.n1422 vdd.n1375 9.3005
R5584 vdd.n1424 vdd.n1423 9.3005
R5585 vdd.n1425 vdd.n1374 9.3005
R5586 vdd.n1427 vdd.n1426 9.3005
R5587 vdd.n1428 vdd.n1369 9.3005
R5588 vdd.n1430 vdd.n1429 9.3005
R5589 vdd.n1431 vdd.n1368 9.3005
R5590 vdd.n1433 vdd.n1432 9.3005
R5591 vdd.n1437 vdd.n1364 9.3005
R5592 vdd.n1439 vdd.n1438 9.3005
R5593 vdd.n1440 vdd.n1363 9.3005
R5594 vdd.n1442 vdd.n1441 9.3005
R5595 vdd.n1443 vdd.n1358 9.3005
R5596 vdd.n1445 vdd.n1444 9.3005
R5597 vdd.n1446 vdd.n1357 9.3005
R5598 vdd.n1448 vdd.n1447 9.3005
R5599 vdd.n1449 vdd.n1352 9.3005
R5600 vdd.n1451 vdd.n1450 9.3005
R5601 vdd.n1452 vdd.n1351 9.3005
R5602 vdd.n1454 vdd.n1453 9.3005
R5603 vdd.n1455 vdd.n1346 9.3005
R5604 vdd.n1457 vdd.n1456 9.3005
R5605 vdd.n1458 vdd.n1345 9.3005
R5606 vdd.n1460 vdd.n1459 9.3005
R5607 vdd.n1461 vdd.n1340 9.3005
R5608 vdd.n1463 vdd.n1462 9.3005
R5609 vdd.n1464 vdd.n1339 9.3005
R5610 vdd.n1466 vdd.n1465 9.3005
R5611 vdd.n1467 vdd.n1334 9.3005
R5612 vdd.n1469 vdd.n1468 9.3005
R5613 vdd.n1470 vdd.n1333 9.3005
R5614 vdd.n1472 vdd.n1471 9.3005
R5615 vdd.n1473 vdd.n1326 9.3005
R5616 vdd.n1475 vdd.n1474 9.3005
R5617 vdd.n1476 vdd.n1325 9.3005
R5618 vdd.n1478 vdd.n1477 9.3005
R5619 vdd.n1479 vdd.n1320 9.3005
R5620 vdd.n1481 vdd.n1480 9.3005
R5621 vdd.n1482 vdd.n1319 9.3005
R5622 vdd.n1484 vdd.n1483 9.3005
R5623 vdd.n1485 vdd.n1314 9.3005
R5624 vdd.n1487 vdd.n1486 9.3005
R5625 vdd.n1488 vdd.n1313 9.3005
R5626 vdd.n1490 vdd.n1489 9.3005
R5627 vdd.n1491 vdd.n1308 9.3005
R5628 vdd.n1493 vdd.n1492 9.3005
R5629 vdd.n1494 vdd.n1307 9.3005
R5630 vdd.n1496 vdd.n1495 9.3005
R5631 vdd.n1272 vdd.n1271 9.3005
R5632 vdd.n1502 vdd.n1501 9.3005
R5633 vdd.n1401 vdd.n1400 9.3005
R5634 vdd.n1505 vdd.n1504 9.3005
R5635 vdd.n1261 vdd.n1260 9.3005
R5636 vdd.n1519 vdd.n1518 9.3005
R5637 vdd.n1520 vdd.n1259 9.3005
R5638 vdd.n1522 vdd.n1521 9.3005
R5639 vdd.n1250 vdd.n1249 9.3005
R5640 vdd.n1536 vdd.n1535 9.3005
R5641 vdd.n1537 vdd.n1248 9.3005
R5642 vdd.n1539 vdd.n1538 9.3005
R5643 vdd.n1239 vdd.n1238 9.3005
R5644 vdd.n1552 vdd.n1551 9.3005
R5645 vdd.n1553 vdd.n1237 9.3005
R5646 vdd.n1555 vdd.n1554 9.3005
R5647 vdd.n1227 vdd.n1226 9.3005
R5648 vdd.n1569 vdd.n1568 9.3005
R5649 vdd.n1570 vdd.n1225 9.3005
R5650 vdd.n1572 vdd.n1571 9.3005
R5651 vdd.n1216 vdd.n1215 9.3005
R5652 vdd.n1585 vdd.n1584 9.3005
R5653 vdd.n1586 vdd.n1214 9.3005
R5654 vdd.n1503 vdd.n1270 9.3005
R5655 vdd.n1806 vdd.n1805 9.3005
R5656 vdd.n1801 vdd.n1800 9.3005
R5657 vdd.n1812 vdd.n1811 9.3005
R5658 vdd.n1814 vdd.n1813 9.3005
R5659 vdd.n1797 vdd.n1796 9.3005
R5660 vdd.n1820 vdd.n1819 9.3005
R5661 vdd.n1822 vdd.n1821 9.3005
R5662 vdd.n1794 vdd.n1791 9.3005
R5663 vdd.n1829 vdd.n1828 9.3005
R5664 vdd.n1865 vdd.n1864 9.3005
R5665 vdd.n1860 vdd.n1859 9.3005
R5666 vdd.n1871 vdd.n1870 9.3005
R5667 vdd.n1873 vdd.n1872 9.3005
R5668 vdd.n1856 vdd.n1855 9.3005
R5669 vdd.n1879 vdd.n1878 9.3005
R5670 vdd.n1881 vdd.n1880 9.3005
R5671 vdd.n1853 vdd.n1850 9.3005
R5672 vdd.n1888 vdd.n1887 9.3005
R5673 vdd.n1704 vdd.n1703 9.3005
R5674 vdd.n1699 vdd.n1698 9.3005
R5675 vdd.n1710 vdd.n1709 9.3005
R5676 vdd.n1712 vdd.n1711 9.3005
R5677 vdd.n1695 vdd.n1694 9.3005
R5678 vdd.n1718 vdd.n1717 9.3005
R5679 vdd.n1720 vdd.n1719 9.3005
R5680 vdd.n1692 vdd.n1689 9.3005
R5681 vdd.n1727 vdd.n1726 9.3005
R5682 vdd.n1763 vdd.n1762 9.3005
R5683 vdd.n1758 vdd.n1757 9.3005
R5684 vdd.n1769 vdd.n1768 9.3005
R5685 vdd.n1771 vdd.n1770 9.3005
R5686 vdd.n1754 vdd.n1753 9.3005
R5687 vdd.n1777 vdd.n1776 9.3005
R5688 vdd.n1779 vdd.n1778 9.3005
R5689 vdd.n1751 vdd.n1748 9.3005
R5690 vdd.n1786 vdd.n1785 9.3005
R5691 vdd.n1603 vdd.n1602 9.3005
R5692 vdd.n1598 vdd.n1597 9.3005
R5693 vdd.n1609 vdd.n1608 9.3005
R5694 vdd.n1611 vdd.n1610 9.3005
R5695 vdd.n1594 vdd.n1593 9.3005
R5696 vdd.n1617 vdd.n1616 9.3005
R5697 vdd.n1619 vdd.n1618 9.3005
R5698 vdd.n1591 vdd.n1588 9.3005
R5699 vdd.n1626 vdd.n1625 9.3005
R5700 vdd.n1662 vdd.n1661 9.3005
R5701 vdd.n1657 vdd.n1656 9.3005
R5702 vdd.n1668 vdd.n1667 9.3005
R5703 vdd.n1670 vdd.n1669 9.3005
R5704 vdd.n1653 vdd.n1652 9.3005
R5705 vdd.n1676 vdd.n1675 9.3005
R5706 vdd.n1678 vdd.n1677 9.3005
R5707 vdd.n1650 vdd.n1647 9.3005
R5708 vdd.n1685 vdd.n1684 9.3005
R5709 vdd.n1541 vdd.t240 9.18308
R5710 vdd.n3513 vdd.t187 9.18308
R5711 vdd.n1235 vdd.t230 8.95635
R5712 vdd.n2196 vdd.t90 8.95635
R5713 vdd.n723 vdd.t64 8.95635
R5714 vdd.t196 vdd.n3567 8.95635
R5715 vdd.n312 vdd.n311 8.92171
R5716 vdd.n253 vdd.n252 8.92171
R5717 vdd.n210 vdd.n209 8.92171
R5718 vdd.n151 vdd.n150 8.92171
R5719 vdd.n109 vdd.n108 8.92171
R5720 vdd.n50 vdd.n49 8.92171
R5721 vdd.n1811 vdd.n1810 8.92171
R5722 vdd.n1870 vdd.n1869 8.92171
R5723 vdd.n1709 vdd.n1708 8.92171
R5724 vdd.n1768 vdd.n1767 8.92171
R5725 vdd.n1608 vdd.n1607 8.92171
R5726 vdd.n1667 vdd.n1666 8.92171
R5727 vdd.n231 vdd.n129 8.81535
R5728 vdd.n1789 vdd.n1687 8.81535
R5729 vdd.n1582 vdd.t146 8.72962
R5730 vdd.t223 vdd.n3576 8.72962
R5731 vdd.n1905 vdd.t143 8.50289
R5732 vdd.n3482 vdd.t168 8.50289
R5733 vdd.n28 vdd.n14 8.42249
R5734 vdd.n1931 vdd.t179 8.27616
R5735 vdd.t225 vdd.n656 8.27616
R5736 vdd.n3582 vdd.n3581 8.16225
R5737 vdd.n1893 vdd.n1892 8.16225
R5738 vdd.n308 vdd.n302 8.14595
R5739 vdd.n249 vdd.n243 8.14595
R5740 vdd.n206 vdd.n200 8.14595
R5741 vdd.n147 vdd.n141 8.14595
R5742 vdd.n105 vdd.n99 8.14595
R5743 vdd.n46 vdd.n40 8.14595
R5744 vdd.n1807 vdd.n1801 8.14595
R5745 vdd.n1866 vdd.n1860 8.14595
R5746 vdd.n1705 vdd.n1699 8.14595
R5747 vdd.n1764 vdd.n1758 8.14595
R5748 vdd.n1604 vdd.n1598 8.14595
R5749 vdd.n1663 vdd.n1657 8.14595
R5750 vdd.n1178 vdd.t155 8.04943
R5751 vdd.n3438 vdd.t152 8.04943
R5752 vdd.n2467 vdd.n1104 7.70933
R5753 vdd.n2473 vdd.n1104 7.70933
R5754 vdd.n2479 vdd.n1098 7.70933
R5755 vdd.n2479 vdd.n1092 7.70933
R5756 vdd.n2485 vdd.n1092 7.70933
R5757 vdd.n2485 vdd.n1086 7.70933
R5758 vdd.n2491 vdd.n1086 7.70933
R5759 vdd.n2497 vdd.n1080 7.70933
R5760 vdd.n2503 vdd.n1074 7.70933
R5761 vdd.n2509 vdd.n1067 7.70933
R5762 vdd.n2509 vdd.n1070 7.70933
R5763 vdd.n2515 vdd.n1063 7.70933
R5764 vdd.n2522 vdd.n1049 7.70933
R5765 vdd.n2528 vdd.n1049 7.70933
R5766 vdd.n2534 vdd.n1043 7.70933
R5767 vdd.n2540 vdd.n1039 7.70933
R5768 vdd.n2546 vdd.n1033 7.70933
R5769 vdd.n2564 vdd.n1015 7.70933
R5770 vdd.n2564 vdd.n1008 7.70933
R5771 vdd.n2572 vdd.n1008 7.70933
R5772 vdd.n2654 vdd.n992 7.70933
R5773 vdd.n3017 vdd.n946 7.70933
R5774 vdd.n3029 vdd.n927 7.70933
R5775 vdd.n3035 vdd.n927 7.70933
R5776 vdd.n3035 vdd.n930 7.70933
R5777 vdd.n3053 vdd.n911 7.70933
R5778 vdd.n3059 vdd.n905 7.70933
R5779 vdd.n3065 vdd.n901 7.70933
R5780 vdd.n3071 vdd.n888 7.70933
R5781 vdd.n3077 vdd.n888 7.70933
R5782 vdd.n3084 vdd.n881 7.70933
R5783 vdd.n3090 vdd.n874 7.70933
R5784 vdd.n3090 vdd.n877 7.70933
R5785 vdd.n3096 vdd.n870 7.70933
R5786 vdd.n3102 vdd.n864 7.70933
R5787 vdd.n3108 vdd.n851 7.70933
R5788 vdd.n3114 vdd.n851 7.70933
R5789 vdd.n3114 vdd.n843 7.70933
R5790 vdd.n3165 vdd.n843 7.70933
R5791 vdd.n3165 vdd.n846 7.70933
R5792 vdd.n3171 vdd.n805 7.70933
R5793 vdd.n3241 vdd.n805 7.70933
R5794 vdd.t17 vdd.n1080 7.59597
R5795 vdd.n2346 vdd.t44 7.59597
R5796 vdd.n2989 vdd.t46 7.59597
R5797 vdd.n864 vdd.t19 7.59597
R5798 vdd.n307 vdd.n304 7.3702
R5799 vdd.n248 vdd.n245 7.3702
R5800 vdd.n205 vdd.n202 7.3702
R5801 vdd.n146 vdd.n143 7.3702
R5802 vdd.n104 vdd.n101 7.3702
R5803 vdd.n45 vdd.n42 7.3702
R5804 vdd.n1806 vdd.n1803 7.3702
R5805 vdd.n1865 vdd.n1862 7.3702
R5806 vdd.n1704 vdd.n1701 7.3702
R5807 vdd.n1763 vdd.n1760 7.3702
R5808 vdd.n1603 vdd.n1600 7.3702
R5809 vdd.n1662 vdd.n1659 7.3702
R5810 vdd.n1964 vdd.t238 7.1425
R5811 vdd.n679 vdd.t198 7.1425
R5812 vdd.n1438 vdd.n1437 6.98232
R5813 vdd.n2119 vdd.n2118 6.98232
R5814 vdd.n566 vdd.n565 6.98232
R5815 vdd.n3323 vdd.n3320 6.98232
R5816 vdd.t166 vdd.n1177 6.91577
R5817 vdd.n2503 vdd.t45 6.91577
R5818 vdd.n3096 vdd.t43 6.91577
R5819 vdd.n3446 vdd.t163 6.91577
R5820 vdd.n3081 vdd.n3080 6.86879
R5821 vdd.n2519 vdd.n2518 6.86879
R5822 vdd.n2579 vdd.t37 6.80241
R5823 vdd.n3023 vdd.t29 6.80241
R5824 vdd.n1923 vdd.t236 6.68904
R5825 vdd.n3462 vdd.t161 6.68904
R5826 vdd.t177 vdd.n1206 6.46231
R5827 vdd.n3490 vdd.t157 6.46231
R5828 vdd.n3582 vdd.n333 6.38151
R5829 vdd.n1892 vdd.n1891 6.38151
R5830 vdd.n2346 vdd.t47 6.34895
R5831 vdd.n2989 vdd.t33 6.34895
R5832 vdd.n1574 vdd.t204 6.23558
R5833 vdd.t150 vdd.n344 6.23558
R5834 vdd.t192 vdd.n1234 6.00885
R5835 vdd.t24 vdd.n1043 6.00885
R5836 vdd.n901 vdd.t13 6.00885
R5837 vdd.n3561 vdd.t159 6.00885
R5838 vdd.n308 vdd.n307 5.81868
R5839 vdd.n249 vdd.n248 5.81868
R5840 vdd.n206 vdd.n205 5.81868
R5841 vdd.n147 vdd.n146 5.81868
R5842 vdd.n105 vdd.n104 5.81868
R5843 vdd.n46 vdd.n45 5.81868
R5844 vdd.n1807 vdd.n1806 5.81868
R5845 vdd.n1866 vdd.n1865 5.81868
R5846 vdd.n1705 vdd.n1704 5.81868
R5847 vdd.n1764 vdd.n1763 5.81868
R5848 vdd.n1604 vdd.n1603 5.81868
R5849 vdd.n1663 vdd.n1662 5.81868
R5850 vdd.n1533 vdd.t181 5.78212
R5851 vdd.n3552 vdd.t278 5.78212
R5852 vdd.n2662 vdd.n2661 5.77611
R5853 vdd.n2402 vdd.n2401 5.77611
R5854 vdd.n2891 vdd.n2890 5.77611
R5855 vdd.n3182 vdd.n3181 5.77611
R5856 vdd.n3246 vdd.n801 5.77611
R5857 vdd.n2827 vdd.n2763 5.77611
R5858 vdd.n2587 vdd.n999 5.77611
R5859 vdd.n2278 vdd.n2277 5.77611
R5860 vdd.n1400 vdd.n1399 5.62474
R5861 vdd.n2202 vdd.n2199 5.62474
R5862 vdd.n3533 vdd.n428 5.62474
R5863 vdd.n3407 vdd.n690 5.62474
R5864 vdd.n1257 vdd.t181 5.55539
R5865 vdd.t278 vdd.n3551 5.55539
R5866 vdd.n2540 vdd.t35 5.44203
R5867 vdd.n3059 vdd.t5 5.44203
R5868 vdd.n1549 vdd.t192 5.32866
R5869 vdd.t159 vdd.n3560 5.32866
R5870 vdd.n1565 vdd.t204 5.10193
R5871 vdd.n2515 vdd.t41 5.10193
R5872 vdd.n2534 vdd.t42 5.10193
R5873 vdd.n3065 vdd.t18 5.10193
R5874 vdd.n3084 vdd.t299 5.10193
R5875 vdd.n3569 vdd.t150 5.10193
R5876 vdd.n311 vdd.n302 5.04292
R5877 vdd.n252 vdd.n243 5.04292
R5878 vdd.n209 vdd.n200 5.04292
R5879 vdd.n150 vdd.n141 5.04292
R5880 vdd.n108 vdd.n99 5.04292
R5881 vdd.n49 vdd.n40 5.04292
R5882 vdd.n1810 vdd.n1801 5.04292
R5883 vdd.n1869 vdd.n1860 5.04292
R5884 vdd.n1708 vdd.n1699 5.04292
R5885 vdd.n1767 vdd.n1758 5.04292
R5886 vdd.n1607 vdd.n1598 5.04292
R5887 vdd.n1666 vdd.n1657 5.04292
R5888 vdd.n1063 vdd.t124 4.98857
R5889 vdd.t83 vdd.n881 4.98857
R5890 vdd.n1897 vdd.t177 4.8752
R5891 vdd.t72 vdd.n1098 4.8752
R5892 vdd.t7 vdd.t22 4.8752
R5893 vdd.n2334 vdd.t110 4.8752
R5894 vdd.n3001 vdd.t114 4.8752
R5895 vdd.t49 vdd.t9 4.8752
R5896 vdd.n846 vdd.t68 4.8752
R5897 vdd.t157 vdd.n340 4.8752
R5898 vdd.n2663 vdd.n2662 4.83952
R5899 vdd.n2403 vdd.n2402 4.83952
R5900 vdd.n2890 vdd.n2889 4.83952
R5901 vdd.n3183 vdd.n3182 4.83952
R5902 vdd.n801 vdd.n796 4.83952
R5903 vdd.n2824 vdd.n2763 4.83952
R5904 vdd.n2590 vdd.n999 4.83952
R5905 vdd.n2277 vdd.n2276 4.83952
R5906 vdd.n2558 vdd.t14 4.76184
R5907 vdd.n3041 vdd.t20 4.76184
R5908 vdd.n2087 vdd.n1145 4.74817
R5909 vdd.n2082 vdd.n1146 4.74817
R5910 vdd.n1984 vdd.n1981 4.74817
R5911 vdd.n2183 vdd.n1985 4.74817
R5912 vdd.n2185 vdd.n1984 4.74817
R5913 vdd.n2184 vdd.n2183 4.74817
R5914 vdd.n3400 vdd.n3399 4.74817
R5915 vdd.n3397 vdd.n3396 4.74817
R5916 vdd.n3397 vdd.n732 4.74817
R5917 vdd.n3399 vdd.n729 4.74817
R5918 vdd.n3282 vdd.n784 4.74817
R5919 vdd.n3278 vdd.n3276 4.74817
R5920 vdd.n3281 vdd.n3276 4.74817
R5921 vdd.n3285 vdd.n784 4.74817
R5922 vdd.n2083 vdd.n1145 4.74817
R5923 vdd.n1148 vdd.n1146 4.74817
R5924 vdd.n333 vdd.n332 4.7074
R5925 vdd.n231 vdd.n230 4.7074
R5926 vdd.n1891 vdd.n1890 4.7074
R5927 vdd.n1789 vdd.n1788 4.7074
R5928 vdd.n1200 vdd.t236 4.64847
R5929 vdd.n3471 vdd.t161 4.64847
R5930 vdd.n1939 vdd.t166 4.42174
R5931 vdd.t163 vdd.n655 4.42174
R5932 vdd.n2334 vdd.t3 4.30838
R5933 vdd.n3001 vdd.t302 4.30838
R5934 vdd.n312 vdd.n300 4.26717
R5935 vdd.n253 vdd.n241 4.26717
R5936 vdd.n210 vdd.n198 4.26717
R5937 vdd.n151 vdd.n139 4.26717
R5938 vdd.n109 vdd.n97 4.26717
R5939 vdd.n50 vdd.n38 4.26717
R5940 vdd.n1811 vdd.n1799 4.26717
R5941 vdd.n1870 vdd.n1858 4.26717
R5942 vdd.n1709 vdd.n1697 4.26717
R5943 vdd.n1768 vdd.n1756 4.26717
R5944 vdd.n1608 vdd.n1596 4.26717
R5945 vdd.n1667 vdd.n1655 4.26717
R5946 vdd.n1955 vdd.t238 4.19501
R5947 vdd.t2 vdd.n1074 4.19501
R5948 vdd.n1033 vdd.t12 4.19501
R5949 vdd.t8 vdd.n911 4.19501
R5950 vdd.n870 vdd.t16 4.19501
R5951 vdd.n3430 vdd.t198 4.19501
R5952 vdd.n333 vdd.n231 4.10845
R5953 vdd.n1891 vdd.n1789 4.10845
R5954 vdd.n289 vdd.t251 4.06363
R5955 vdd.n289 vdd.t291 4.06363
R5956 vdd.n287 vdd.t160 4.06363
R5957 vdd.n287 vdd.t213 4.06363
R5958 vdd.n285 vdd.t216 4.06363
R5959 vdd.n285 vdd.t269 4.06363
R5960 vdd.n283 vdd.t271 4.06363
R5961 vdd.n283 vdd.t151 4.06363
R5962 vdd.n281 vdd.t174 4.06363
R5963 vdd.n281 vdd.t245 4.06363
R5964 vdd.n279 vdd.t272 4.06363
R5965 vdd.n279 vdd.t287 4.06363
R5966 vdd.n277 vdd.t290 4.06363
R5967 vdd.n277 vdd.t183 4.06363
R5968 vdd.n275 vdd.t214 4.06363
R5969 vdd.n275 vdd.t289 4.06363
R5970 vdd.n273 vdd.t295 4.06363
R5971 vdd.n273 vdd.t212 4.06363
R5972 vdd.n187 vdd.t243 4.06363
R5973 vdd.n187 vdd.t279 4.06363
R5974 vdd.n185 vdd.t296 4.06363
R5975 vdd.n185 vdd.t188 4.06363
R5976 vdd.n183 vdd.t197 4.06363
R5977 vdd.n183 vdd.t259 4.06363
R5978 vdd.n181 vdd.t260 4.06363
R5979 vdd.n181 vdd.t288 4.06363
R5980 vdd.n179 vdd.t158 4.06363
R5981 vdd.n179 vdd.t224 4.06363
R5982 vdd.n177 vdd.t263 4.06363
R5983 vdd.n177 vdd.t273 4.06363
R5984 vdd.n175 vdd.t281 4.06363
R5985 vdd.n175 vdd.t162 4.06363
R5986 vdd.n173 vdd.t189 4.06363
R5987 vdd.n173 vdd.t280 4.06363
R5988 vdd.n171 vdd.t284 4.06363
R5989 vdd.n171 vdd.t186 4.06363
R5990 vdd.n86 vdd.t218 4.06363
R5991 vdd.n86 vdd.t292 4.06363
R5992 vdd.n84 vdd.t194 4.06363
R5993 vdd.n84 vdd.t276 4.06363
R5994 vdd.n82 vdd.t229 4.06363
R5995 vdd.n82 vdd.t261 4.06363
R5996 vdd.n80 vdd.t209 4.06363
R5997 vdd.n80 vdd.t285 4.06363
R5998 vdd.n78 vdd.t173 4.06363
R5999 vdd.n78 vdd.t270 4.06363
R6000 vdd.n76 vdd.t169 4.06363
R6001 vdd.n76 vdd.t255 4.06363
R6002 vdd.n74 vdd.t191 4.06363
R6003 vdd.n74 vdd.t274 4.06363
R6004 vdd.n72 vdd.t164 4.06363
R6005 vdd.n72 vdd.t226 4.06363
R6006 vdd.n70 vdd.t153 4.06363
R6007 vdd.n70 vdd.t200 4.06363
R6008 vdd.n1831 vdd.t264 4.06363
R6009 vdd.n1831 vdd.t211 4.06363
R6010 vdd.n1833 vdd.t206 4.06363
R6011 vdd.n1833 vdd.t266 4.06363
R6012 vdd.n1835 vdd.t250 4.06363
R6013 vdd.n1835 vdd.t248 4.06363
R6014 vdd.n1837 vdd.t201 4.06363
R6015 vdd.n1837 vdd.t172 4.06363
R6016 vdd.n1839 vdd.t170 4.06363
R6017 vdd.n1839 vdd.t247 4.06363
R6018 vdd.n1841 vdd.t222 4.06363
R6019 vdd.n1841 vdd.t171 4.06363
R6020 vdd.n1843 vdd.t165 4.06363
R6021 vdd.n1843 vdd.t267 4.06363
R6022 vdd.n1845 vdd.t265 4.06363
R6023 vdd.n1845 vdd.t215 4.06363
R6024 vdd.n1847 vdd.t207 4.06363
R6025 vdd.n1847 vdd.t294 4.06363
R6026 vdd.n1729 vdd.t252 4.06363
R6027 vdd.n1729 vdd.t184 4.06363
R6028 vdd.n1731 vdd.t180 4.06363
R6029 vdd.n1731 vdd.t253 4.06363
R6030 vdd.n1733 vdd.t237 4.06363
R6031 vdd.n1733 vdd.t233 4.06363
R6032 vdd.n1735 vdd.t176 4.06363
R6033 vdd.n1735 vdd.t154 4.06363
R6034 vdd.n1737 vdd.t147 4.06363
R6035 vdd.n1737 vdd.t228 4.06363
R6036 vdd.n1739 vdd.t205 4.06363
R6037 vdd.n1739 vdd.t149 4.06363
R6038 vdd.n1741 vdd.t140 4.06363
R6039 vdd.n1741 vdd.t257 4.06363
R6040 vdd.n1743 vdd.t241 4.06363
R6041 vdd.n1743 vdd.t195 4.06363
R6042 vdd.n1745 vdd.t182 4.06363
R6043 vdd.n1745 vdd.t283 4.06363
R6044 vdd.n1628 vdd.t203 4.06363
R6045 vdd.n1628 vdd.t156 4.06363
R6046 vdd.n1630 vdd.t227 4.06363
R6047 vdd.n1630 vdd.t167 4.06363
R6048 vdd.n1632 vdd.t275 4.06363
R6049 vdd.n1632 vdd.t297 4.06363
R6050 vdd.n1634 vdd.t256 4.06363
R6051 vdd.n1634 vdd.t144 4.06363
R6052 vdd.n1636 vdd.t242 4.06363
R6053 vdd.n1636 vdd.t178 4.06363
R6054 vdd.n1638 vdd.t286 4.06363
R6055 vdd.n1638 vdd.t210 4.06363
R6056 vdd.n1640 vdd.t262 4.06363
R6057 vdd.n1640 vdd.t231 4.06363
R6058 vdd.n1642 vdd.t277 4.06363
R6059 vdd.n1642 vdd.t193 4.06363
R6060 vdd.n1644 vdd.t293 4.06363
R6061 vdd.n1644 vdd.t221 4.06363
R6062 vdd.n26 vdd.t55 3.9605
R6063 vdd.n26 vdd.t59 3.9605
R6064 vdd.n23 vdd.t60 3.9605
R6065 vdd.n23 vdd.t61 3.9605
R6066 vdd.n21 vdd.t58 3.9605
R6067 vdd.n21 vdd.t57 3.9605
R6068 vdd.n20 vdd.t54 3.9605
R6069 vdd.n20 vdd.t28 3.9605
R6070 vdd.n15 vdd.t51 3.9605
R6071 vdd.n15 vdd.t56 3.9605
R6072 vdd.n16 vdd.t62 3.9605
R6073 vdd.n16 vdd.t27 3.9605
R6074 vdd.n18 vdd.t53 3.9605
R6075 vdd.n18 vdd.t300 3.9605
R6076 vdd.n25 vdd.t301 3.9605
R6077 vdd.n25 vdd.t52 3.9605
R6078 vdd.n3080 vdd.n3079 3.74684
R6079 vdd.n2520 vdd.n2519 3.74684
R6080 vdd.n7 vdd.t50 3.61217
R6081 vdd.n7 vdd.t6 3.61217
R6082 vdd.n8 vdd.t21 3.61217
R6083 vdd.n8 vdd.t34 3.61217
R6084 vdd.n10 vdd.t30 3.61217
R6085 vdd.n10 vdd.t303 3.61217
R6086 vdd.n12 vdd.t1 3.61217
R6087 vdd.n12 vdd.t32 3.61217
R6088 vdd.n5 vdd.t40 3.61217
R6089 vdd.n5 vdd.t11 3.61217
R6090 vdd.n3 vdd.t4 3.61217
R6091 vdd.n3 vdd.t38 3.61217
R6092 vdd.n1 vdd.t48 3.61217
R6093 vdd.n1 vdd.t15 3.61217
R6094 vdd.n0 vdd.t36 3.61217
R6095 vdd.n0 vdd.t23 3.61217
R6096 vdd.n2497 vdd.t2 3.51482
R6097 vdd.n2552 vdd.t12 3.51482
R6098 vdd.n3047 vdd.t8 3.51482
R6099 vdd.n3102 vdd.t16 3.51482
R6100 vdd.n316 vdd.n315 3.49141
R6101 vdd.n257 vdd.n256 3.49141
R6102 vdd.n214 vdd.n213 3.49141
R6103 vdd.n155 vdd.n154 3.49141
R6104 vdd.n113 vdd.n112 3.49141
R6105 vdd.n54 vdd.n53 3.49141
R6106 vdd.n1815 vdd.n1814 3.49141
R6107 vdd.n1874 vdd.n1873 3.49141
R6108 vdd.n1713 vdd.n1712 3.49141
R6109 vdd.n1772 vdd.n1771 3.49141
R6110 vdd.n1612 vdd.n1611 3.49141
R6111 vdd.n1671 vdd.n1670 3.49141
R6112 vdd.n2572 vdd.t3 3.40145
R6113 vdd.n2726 vdd.t39 3.40145
R6114 vdd.n3010 vdd.t31 3.40145
R6115 vdd.n3029 vdd.t302 3.40145
R6116 vdd.n1956 vdd.t155 3.28809
R6117 vdd.n3429 vdd.t152 3.28809
R6118 vdd.t179 vdd.n1184 3.06136
R6119 vdd.n3454 vdd.t225 3.06136
R6120 vdd.t14 vdd.n1015 2.94799
R6121 vdd.n930 vdd.t20 2.94799
R6122 vdd.n1914 vdd.t143 2.83463
R6123 vdd.n2473 vdd.t72 2.83463
R6124 vdd.n2579 vdd.t110 2.83463
R6125 vdd.n3023 vdd.t114 2.83463
R6126 vdd.n3171 vdd.t68 2.83463
R6127 vdd.n644 vdd.t168 2.83463
R6128 vdd.n319 vdd.n298 2.71565
R6129 vdd.n260 vdd.n239 2.71565
R6130 vdd.n217 vdd.n196 2.71565
R6131 vdd.n158 vdd.n137 2.71565
R6132 vdd.n116 vdd.n95 2.71565
R6133 vdd.n57 vdd.n36 2.71565
R6134 vdd.n1818 vdd.n1797 2.71565
R6135 vdd.n1877 vdd.n1856 2.71565
R6136 vdd.n1716 vdd.n1695 2.71565
R6137 vdd.n1775 vdd.n1754 2.71565
R6138 vdd.n1615 vdd.n1594 2.71565
R6139 vdd.n1674 vdd.n1653 2.71565
R6140 vdd.t146 vdd.n1212 2.6079
R6141 vdd.n1070 vdd.t41 2.6079
R6142 vdd.n2358 vdd.t42 2.6079
R6143 vdd.n2977 vdd.t18 2.6079
R6144 vdd.t299 vdd.n874 2.6079
R6145 vdd.n3577 vdd.t223 2.6079
R6146 vdd.n306 vdd.n305 2.4129
R6147 vdd.n247 vdd.n246 2.4129
R6148 vdd.n204 vdd.n203 2.4129
R6149 vdd.n145 vdd.n144 2.4129
R6150 vdd.n103 vdd.n102 2.4129
R6151 vdd.n44 vdd.n43 2.4129
R6152 vdd.n1805 vdd.n1804 2.4129
R6153 vdd.n1864 vdd.n1863 2.4129
R6154 vdd.n1703 vdd.n1702 2.4129
R6155 vdd.n1762 vdd.n1761 2.4129
R6156 vdd.n1602 vdd.n1601 2.4129
R6157 vdd.n1661 vdd.n1660 2.4129
R6158 vdd.n1566 vdd.t230 2.38117
R6159 vdd.n1974 vdd.t90 2.38117
R6160 vdd.n3413 vdd.t64 2.38117
R6161 vdd.n3568 vdd.t196 2.38117
R6162 vdd.n2182 vdd.n1984 2.27742
R6163 vdd.n2183 vdd.n2182 2.27742
R6164 vdd.n3398 vdd.n3397 2.27742
R6165 vdd.n3399 vdd.n3398 2.27742
R6166 vdd.n3276 vdd.n3275 2.27742
R6167 vdd.n3275 vdd.n784 2.27742
R6168 vdd.n2205 vdd.n1145 2.27742
R6169 vdd.n2205 vdd.n1146 2.27742
R6170 vdd.n2358 vdd.t35 2.2678
R6171 vdd.n2977 vdd.t5 2.2678
R6172 vdd.t240 vdd.n1241 2.15444
R6173 vdd.n3559 vdd.t187 2.15444
R6174 vdd.n2546 vdd.t22 2.04107
R6175 vdd.n3053 vdd.t49 2.04107
R6176 vdd.n320 vdd.n296 1.93989
R6177 vdd.n261 vdd.n237 1.93989
R6178 vdd.n218 vdd.n194 1.93989
R6179 vdd.n159 vdd.n135 1.93989
R6180 vdd.n117 vdd.n93 1.93989
R6181 vdd.n58 vdd.n34 1.93989
R6182 vdd.n1819 vdd.n1795 1.93989
R6183 vdd.n1878 vdd.n1854 1.93989
R6184 vdd.n1717 vdd.n1693 1.93989
R6185 vdd.n1776 vdd.n1752 1.93989
R6186 vdd.n1616 vdd.n1592 1.93989
R6187 vdd.n1675 vdd.n1651 1.93989
R6188 vdd.n1524 vdd.t234 1.92771
R6189 vdd.t141 vdd.n375 1.92771
R6190 vdd.n1532 vdd.t220 1.70098
R6191 vdd.n2522 vdd.t26 1.70098
R6192 vdd.n2528 vdd.t24 1.70098
R6193 vdd.n3071 vdd.t13 1.70098
R6194 vdd.n3077 vdd.t25 1.70098
R6195 vdd.n3553 vdd.t217 1.70098
R6196 vdd.n1557 vdd.t139 1.47425
R6197 vdd.n361 vdd.t258 1.47425
R6198 vdd.n2552 vdd.t47 1.36088
R6199 vdd.n3047 vdd.t33 1.36088
R6200 vdd.n1223 vdd.t148 1.24752
R6201 vdd.t208 vdd.n3575 1.24752
R6202 vdd.n331 vdd.n291 1.16414
R6203 vdd.n324 vdd.n323 1.16414
R6204 vdd.n272 vdd.n232 1.16414
R6205 vdd.n265 vdd.n264 1.16414
R6206 vdd.n229 vdd.n189 1.16414
R6207 vdd.n222 vdd.n221 1.16414
R6208 vdd.n170 vdd.n130 1.16414
R6209 vdd.n163 vdd.n162 1.16414
R6210 vdd.n128 vdd.n88 1.16414
R6211 vdd.n121 vdd.n120 1.16414
R6212 vdd.n69 vdd.n29 1.16414
R6213 vdd.n62 vdd.n61 1.16414
R6214 vdd.n1830 vdd.n1790 1.16414
R6215 vdd.n1823 vdd.n1822 1.16414
R6216 vdd.n1889 vdd.n1849 1.16414
R6217 vdd.n1882 vdd.n1881 1.16414
R6218 vdd.n1728 vdd.n1688 1.16414
R6219 vdd.n1721 vdd.n1720 1.16414
R6220 vdd.n1787 vdd.n1747 1.16414
R6221 vdd.n1780 vdd.n1779 1.16414
R6222 vdd.n1627 vdd.n1587 1.16414
R6223 vdd.n1620 vdd.n1619 1.16414
R6224 vdd.n1686 vdd.n1646 1.16414
R6225 vdd.n1679 vdd.n1678 1.16414
R6226 vdd.n1892 vdd.n28 1.11236
R6227 vdd vdd.n3582 1.10453
R6228 vdd.n1906 vdd.t175 1.02079
R6229 vdd.t124 vdd.t26 1.02079
R6230 vdd.t25 vdd.t83 1.02079
R6231 vdd.t254 vdd.n633 1.02079
R6232 vdd.n1403 vdd.n1399 0.970197
R6233 vdd.n2203 vdd.n2202 0.970197
R6234 vdd.n618 vdd.n428 0.970197
R6235 vdd.n3277 vdd.n690 0.970197
R6236 vdd.t37 vdd.n992 0.907421
R6237 vdd.n946 vdd.t29 0.907421
R6238 vdd.n1922 vdd.t232 0.794056
R6239 vdd.t45 vdd.n1067 0.794056
R6240 vdd.n1039 vdd.t7 0.794056
R6241 vdd.t9 vdd.n905 0.794056
R6242 vdd.n877 vdd.t43 0.794056
R6243 vdd.n3463 vdd.t190 0.794056
R6244 vdd.n1947 vdd.t202 0.567326
R6245 vdd.t185 vdd.n662 0.567326
R6246 vdd.n2193 vdd.n2192 0.530988
R6247 vdd.n726 vdd.n682 0.530988
R6248 vdd.n464 vdd.n391 0.530988
R6249 vdd.n3532 vdd.n3531 0.530988
R6250 vdd.n3409 vdd.n3408 0.530988
R6251 vdd.n1969 vdd.n1147 0.530988
R6252 vdd.n1401 vdd.n1266 0.530988
R6253 vdd.n1503 vdd.n1502 0.530988
R6254 vdd.n4 vdd.n2 0.459552
R6255 vdd.n11 vdd.n9 0.459552
R6256 vdd.n329 vdd.n328 0.388379
R6257 vdd.n295 vdd.n293 0.388379
R6258 vdd.n270 vdd.n269 0.388379
R6259 vdd.n236 vdd.n234 0.388379
R6260 vdd.n227 vdd.n226 0.388379
R6261 vdd.n193 vdd.n191 0.388379
R6262 vdd.n168 vdd.n167 0.388379
R6263 vdd.n134 vdd.n132 0.388379
R6264 vdd.n126 vdd.n125 0.388379
R6265 vdd.n92 vdd.n90 0.388379
R6266 vdd.n67 vdd.n66 0.388379
R6267 vdd.n33 vdd.n31 0.388379
R6268 vdd.n1828 vdd.n1827 0.388379
R6269 vdd.n1794 vdd.n1792 0.388379
R6270 vdd.n1887 vdd.n1886 0.388379
R6271 vdd.n1853 vdd.n1851 0.388379
R6272 vdd.n1726 vdd.n1725 0.388379
R6273 vdd.n1692 vdd.n1690 0.388379
R6274 vdd.n1785 vdd.n1784 0.388379
R6275 vdd.n1751 vdd.n1749 0.388379
R6276 vdd.n1625 vdd.n1624 0.388379
R6277 vdd.n1591 vdd.n1589 0.388379
R6278 vdd.n1684 vdd.n1683 0.388379
R6279 vdd.n1650 vdd.n1648 0.388379
R6280 vdd.n19 vdd.n17 0.387128
R6281 vdd.n24 vdd.n22 0.387128
R6282 vdd.n6 vdd.n4 0.358259
R6283 vdd.n13 vdd.n11 0.358259
R6284 vdd.n276 vdd.n274 0.358259
R6285 vdd.n278 vdd.n276 0.358259
R6286 vdd.n280 vdd.n278 0.358259
R6287 vdd.n282 vdd.n280 0.358259
R6288 vdd.n284 vdd.n282 0.358259
R6289 vdd.n286 vdd.n284 0.358259
R6290 vdd.n288 vdd.n286 0.358259
R6291 vdd.n290 vdd.n288 0.358259
R6292 vdd.n332 vdd.n290 0.358259
R6293 vdd.n174 vdd.n172 0.358259
R6294 vdd.n176 vdd.n174 0.358259
R6295 vdd.n178 vdd.n176 0.358259
R6296 vdd.n180 vdd.n178 0.358259
R6297 vdd.n182 vdd.n180 0.358259
R6298 vdd.n184 vdd.n182 0.358259
R6299 vdd.n186 vdd.n184 0.358259
R6300 vdd.n188 vdd.n186 0.358259
R6301 vdd.n230 vdd.n188 0.358259
R6302 vdd.n73 vdd.n71 0.358259
R6303 vdd.n75 vdd.n73 0.358259
R6304 vdd.n77 vdd.n75 0.358259
R6305 vdd.n79 vdd.n77 0.358259
R6306 vdd.n81 vdd.n79 0.358259
R6307 vdd.n83 vdd.n81 0.358259
R6308 vdd.n85 vdd.n83 0.358259
R6309 vdd.n87 vdd.n85 0.358259
R6310 vdd.n129 vdd.n87 0.358259
R6311 vdd.n1890 vdd.n1848 0.358259
R6312 vdd.n1848 vdd.n1846 0.358259
R6313 vdd.n1846 vdd.n1844 0.358259
R6314 vdd.n1844 vdd.n1842 0.358259
R6315 vdd.n1842 vdd.n1840 0.358259
R6316 vdd.n1840 vdd.n1838 0.358259
R6317 vdd.n1838 vdd.n1836 0.358259
R6318 vdd.n1836 vdd.n1834 0.358259
R6319 vdd.n1834 vdd.n1832 0.358259
R6320 vdd.n1788 vdd.n1746 0.358259
R6321 vdd.n1746 vdd.n1744 0.358259
R6322 vdd.n1744 vdd.n1742 0.358259
R6323 vdd.n1742 vdd.n1740 0.358259
R6324 vdd.n1740 vdd.n1738 0.358259
R6325 vdd.n1738 vdd.n1736 0.358259
R6326 vdd.n1736 vdd.n1734 0.358259
R6327 vdd.n1734 vdd.n1732 0.358259
R6328 vdd.n1732 vdd.n1730 0.358259
R6329 vdd.n1687 vdd.n1645 0.358259
R6330 vdd.n1645 vdd.n1643 0.358259
R6331 vdd.n1643 vdd.n1641 0.358259
R6332 vdd.n1641 vdd.n1639 0.358259
R6333 vdd.n1639 vdd.n1637 0.358259
R6334 vdd.n1637 vdd.n1635 0.358259
R6335 vdd.n1635 vdd.n1633 0.358259
R6336 vdd.n1633 vdd.n1631 0.358259
R6337 vdd.n1631 vdd.n1629 0.358259
R6338 vdd.n14 vdd.n6 0.334552
R6339 vdd.n14 vdd.n13 0.334552
R6340 vdd.n27 vdd.n19 0.21707
R6341 vdd.n27 vdd.n24 0.21707
R6342 vdd.n330 vdd.n292 0.155672
R6343 vdd.n322 vdd.n292 0.155672
R6344 vdd.n322 vdd.n321 0.155672
R6345 vdd.n321 vdd.n297 0.155672
R6346 vdd.n314 vdd.n297 0.155672
R6347 vdd.n314 vdd.n313 0.155672
R6348 vdd.n313 vdd.n301 0.155672
R6349 vdd.n306 vdd.n301 0.155672
R6350 vdd.n271 vdd.n233 0.155672
R6351 vdd.n263 vdd.n233 0.155672
R6352 vdd.n263 vdd.n262 0.155672
R6353 vdd.n262 vdd.n238 0.155672
R6354 vdd.n255 vdd.n238 0.155672
R6355 vdd.n255 vdd.n254 0.155672
R6356 vdd.n254 vdd.n242 0.155672
R6357 vdd.n247 vdd.n242 0.155672
R6358 vdd.n228 vdd.n190 0.155672
R6359 vdd.n220 vdd.n190 0.155672
R6360 vdd.n220 vdd.n219 0.155672
R6361 vdd.n219 vdd.n195 0.155672
R6362 vdd.n212 vdd.n195 0.155672
R6363 vdd.n212 vdd.n211 0.155672
R6364 vdd.n211 vdd.n199 0.155672
R6365 vdd.n204 vdd.n199 0.155672
R6366 vdd.n169 vdd.n131 0.155672
R6367 vdd.n161 vdd.n131 0.155672
R6368 vdd.n161 vdd.n160 0.155672
R6369 vdd.n160 vdd.n136 0.155672
R6370 vdd.n153 vdd.n136 0.155672
R6371 vdd.n153 vdd.n152 0.155672
R6372 vdd.n152 vdd.n140 0.155672
R6373 vdd.n145 vdd.n140 0.155672
R6374 vdd.n127 vdd.n89 0.155672
R6375 vdd.n119 vdd.n89 0.155672
R6376 vdd.n119 vdd.n118 0.155672
R6377 vdd.n118 vdd.n94 0.155672
R6378 vdd.n111 vdd.n94 0.155672
R6379 vdd.n111 vdd.n110 0.155672
R6380 vdd.n110 vdd.n98 0.155672
R6381 vdd.n103 vdd.n98 0.155672
R6382 vdd.n68 vdd.n30 0.155672
R6383 vdd.n60 vdd.n30 0.155672
R6384 vdd.n60 vdd.n59 0.155672
R6385 vdd.n59 vdd.n35 0.155672
R6386 vdd.n52 vdd.n35 0.155672
R6387 vdd.n52 vdd.n51 0.155672
R6388 vdd.n51 vdd.n39 0.155672
R6389 vdd.n44 vdd.n39 0.155672
R6390 vdd.n1829 vdd.n1791 0.155672
R6391 vdd.n1821 vdd.n1791 0.155672
R6392 vdd.n1821 vdd.n1820 0.155672
R6393 vdd.n1820 vdd.n1796 0.155672
R6394 vdd.n1813 vdd.n1796 0.155672
R6395 vdd.n1813 vdd.n1812 0.155672
R6396 vdd.n1812 vdd.n1800 0.155672
R6397 vdd.n1805 vdd.n1800 0.155672
R6398 vdd.n1888 vdd.n1850 0.155672
R6399 vdd.n1880 vdd.n1850 0.155672
R6400 vdd.n1880 vdd.n1879 0.155672
R6401 vdd.n1879 vdd.n1855 0.155672
R6402 vdd.n1872 vdd.n1855 0.155672
R6403 vdd.n1872 vdd.n1871 0.155672
R6404 vdd.n1871 vdd.n1859 0.155672
R6405 vdd.n1864 vdd.n1859 0.155672
R6406 vdd.n1727 vdd.n1689 0.155672
R6407 vdd.n1719 vdd.n1689 0.155672
R6408 vdd.n1719 vdd.n1718 0.155672
R6409 vdd.n1718 vdd.n1694 0.155672
R6410 vdd.n1711 vdd.n1694 0.155672
R6411 vdd.n1711 vdd.n1710 0.155672
R6412 vdd.n1710 vdd.n1698 0.155672
R6413 vdd.n1703 vdd.n1698 0.155672
R6414 vdd.n1786 vdd.n1748 0.155672
R6415 vdd.n1778 vdd.n1748 0.155672
R6416 vdd.n1778 vdd.n1777 0.155672
R6417 vdd.n1777 vdd.n1753 0.155672
R6418 vdd.n1770 vdd.n1753 0.155672
R6419 vdd.n1770 vdd.n1769 0.155672
R6420 vdd.n1769 vdd.n1757 0.155672
R6421 vdd.n1762 vdd.n1757 0.155672
R6422 vdd.n1626 vdd.n1588 0.155672
R6423 vdd.n1618 vdd.n1588 0.155672
R6424 vdd.n1618 vdd.n1617 0.155672
R6425 vdd.n1617 vdd.n1593 0.155672
R6426 vdd.n1610 vdd.n1593 0.155672
R6427 vdd.n1610 vdd.n1609 0.155672
R6428 vdd.n1609 vdd.n1597 0.155672
R6429 vdd.n1602 vdd.n1597 0.155672
R6430 vdd.n1685 vdd.n1647 0.155672
R6431 vdd.n1677 vdd.n1647 0.155672
R6432 vdd.n1677 vdd.n1676 0.155672
R6433 vdd.n1676 vdd.n1652 0.155672
R6434 vdd.n1669 vdd.n1652 0.155672
R6435 vdd.n1669 vdd.n1668 0.155672
R6436 vdd.n1668 vdd.n1656 0.155672
R6437 vdd.n1661 vdd.n1656 0.155672
R6438 vdd.n2181 vdd.n1986 0.152939
R6439 vdd.n1992 vdd.n1986 0.152939
R6440 vdd.n1993 vdd.n1992 0.152939
R6441 vdd.n1994 vdd.n1993 0.152939
R6442 vdd.n1995 vdd.n1994 0.152939
R6443 vdd.n1999 vdd.n1995 0.152939
R6444 vdd.n2000 vdd.n1999 0.152939
R6445 vdd.n2001 vdd.n2000 0.152939
R6446 vdd.n2002 vdd.n2001 0.152939
R6447 vdd.n2006 vdd.n2002 0.152939
R6448 vdd.n2007 vdd.n2006 0.152939
R6449 vdd.n2008 vdd.n2007 0.152939
R6450 vdd.n2156 vdd.n2008 0.152939
R6451 vdd.n2156 vdd.n2155 0.152939
R6452 vdd.n2155 vdd.n2154 0.152939
R6453 vdd.n2154 vdd.n2014 0.152939
R6454 vdd.n2019 vdd.n2014 0.152939
R6455 vdd.n2020 vdd.n2019 0.152939
R6456 vdd.n2021 vdd.n2020 0.152939
R6457 vdd.n2025 vdd.n2021 0.152939
R6458 vdd.n2026 vdd.n2025 0.152939
R6459 vdd.n2027 vdd.n2026 0.152939
R6460 vdd.n2028 vdd.n2027 0.152939
R6461 vdd.n2032 vdd.n2028 0.152939
R6462 vdd.n2033 vdd.n2032 0.152939
R6463 vdd.n2034 vdd.n2033 0.152939
R6464 vdd.n2035 vdd.n2034 0.152939
R6465 vdd.n2039 vdd.n2035 0.152939
R6466 vdd.n2040 vdd.n2039 0.152939
R6467 vdd.n2041 vdd.n2040 0.152939
R6468 vdd.n2042 vdd.n2041 0.152939
R6469 vdd.n2046 vdd.n2042 0.152939
R6470 vdd.n2047 vdd.n2046 0.152939
R6471 vdd.n2048 vdd.n2047 0.152939
R6472 vdd.n2117 vdd.n2048 0.152939
R6473 vdd.n2117 vdd.n2116 0.152939
R6474 vdd.n2116 vdd.n2115 0.152939
R6475 vdd.n2115 vdd.n2054 0.152939
R6476 vdd.n2059 vdd.n2054 0.152939
R6477 vdd.n2060 vdd.n2059 0.152939
R6478 vdd.n2061 vdd.n2060 0.152939
R6479 vdd.n2065 vdd.n2061 0.152939
R6480 vdd.n2066 vdd.n2065 0.152939
R6481 vdd.n2067 vdd.n2066 0.152939
R6482 vdd.n2068 vdd.n2067 0.152939
R6483 vdd.n2072 vdd.n2068 0.152939
R6484 vdd.n2073 vdd.n2072 0.152939
R6485 vdd.n2074 vdd.n2073 0.152939
R6486 vdd.n2075 vdd.n2074 0.152939
R6487 vdd.n2076 vdd.n2075 0.152939
R6488 vdd.n2076 vdd.n1144 0.152939
R6489 vdd.n2192 vdd.n1980 0.152939
R6490 vdd.n1894 vdd.n1203 0.152939
R6491 vdd.n1909 vdd.n1203 0.152939
R6492 vdd.n1910 vdd.n1909 0.152939
R6493 vdd.n1911 vdd.n1910 0.152939
R6494 vdd.n1911 vdd.n1192 0.152939
R6495 vdd.n1926 vdd.n1192 0.152939
R6496 vdd.n1927 vdd.n1926 0.152939
R6497 vdd.n1928 vdd.n1927 0.152939
R6498 vdd.n1928 vdd.n1181 0.152939
R6499 vdd.n1942 vdd.n1181 0.152939
R6500 vdd.n1943 vdd.n1942 0.152939
R6501 vdd.n1944 vdd.n1943 0.152939
R6502 vdd.n1944 vdd.n1169 0.152939
R6503 vdd.n1959 vdd.n1169 0.152939
R6504 vdd.n1960 vdd.n1959 0.152939
R6505 vdd.n1961 vdd.n1960 0.152939
R6506 vdd.n1961 vdd.n1157 0.152939
R6507 vdd.n1978 vdd.n1157 0.152939
R6508 vdd.n1979 vdd.n1978 0.152939
R6509 vdd.n2193 vdd.n1979 0.152939
R6510 vdd.n735 vdd.n730 0.152939
R6511 vdd.n736 vdd.n735 0.152939
R6512 vdd.n737 vdd.n736 0.152939
R6513 vdd.n738 vdd.n737 0.152939
R6514 vdd.n739 vdd.n738 0.152939
R6515 vdd.n740 vdd.n739 0.152939
R6516 vdd.n741 vdd.n740 0.152939
R6517 vdd.n742 vdd.n741 0.152939
R6518 vdd.n743 vdd.n742 0.152939
R6519 vdd.n744 vdd.n743 0.152939
R6520 vdd.n745 vdd.n744 0.152939
R6521 vdd.n746 vdd.n745 0.152939
R6522 vdd.n3365 vdd.n746 0.152939
R6523 vdd.n3365 vdd.n3364 0.152939
R6524 vdd.n3364 vdd.n3363 0.152939
R6525 vdd.n3363 vdd.n748 0.152939
R6526 vdd.n749 vdd.n748 0.152939
R6527 vdd.n750 vdd.n749 0.152939
R6528 vdd.n751 vdd.n750 0.152939
R6529 vdd.n752 vdd.n751 0.152939
R6530 vdd.n753 vdd.n752 0.152939
R6531 vdd.n754 vdd.n753 0.152939
R6532 vdd.n755 vdd.n754 0.152939
R6533 vdd.n756 vdd.n755 0.152939
R6534 vdd.n757 vdd.n756 0.152939
R6535 vdd.n758 vdd.n757 0.152939
R6536 vdd.n759 vdd.n758 0.152939
R6537 vdd.n760 vdd.n759 0.152939
R6538 vdd.n761 vdd.n760 0.152939
R6539 vdd.n762 vdd.n761 0.152939
R6540 vdd.n763 vdd.n762 0.152939
R6541 vdd.n764 vdd.n763 0.152939
R6542 vdd.n765 vdd.n764 0.152939
R6543 vdd.n766 vdd.n765 0.152939
R6544 vdd.n3319 vdd.n766 0.152939
R6545 vdd.n3319 vdd.n3318 0.152939
R6546 vdd.n3318 vdd.n3317 0.152939
R6547 vdd.n3317 vdd.n770 0.152939
R6548 vdd.n771 vdd.n770 0.152939
R6549 vdd.n772 vdd.n771 0.152939
R6550 vdd.n773 vdd.n772 0.152939
R6551 vdd.n774 vdd.n773 0.152939
R6552 vdd.n775 vdd.n774 0.152939
R6553 vdd.n776 vdd.n775 0.152939
R6554 vdd.n777 vdd.n776 0.152939
R6555 vdd.n778 vdd.n777 0.152939
R6556 vdd.n779 vdd.n778 0.152939
R6557 vdd.n780 vdd.n779 0.152939
R6558 vdd.n781 vdd.n780 0.152939
R6559 vdd.n782 vdd.n781 0.152939
R6560 vdd.n783 vdd.n782 0.152939
R6561 vdd.n727 vdd.n726 0.152939
R6562 vdd.n3416 vdd.n682 0.152939
R6563 vdd.n3417 vdd.n3416 0.152939
R6564 vdd.n3418 vdd.n3417 0.152939
R6565 vdd.n3418 vdd.n670 0.152939
R6566 vdd.n3433 vdd.n670 0.152939
R6567 vdd.n3434 vdd.n3433 0.152939
R6568 vdd.n3435 vdd.n3434 0.152939
R6569 vdd.n3435 vdd.n659 0.152939
R6570 vdd.n3449 vdd.n659 0.152939
R6571 vdd.n3450 vdd.n3449 0.152939
R6572 vdd.n3451 vdd.n3450 0.152939
R6573 vdd.n3451 vdd.n647 0.152939
R6574 vdd.n3466 vdd.n647 0.152939
R6575 vdd.n3467 vdd.n3466 0.152939
R6576 vdd.n3468 vdd.n3467 0.152939
R6577 vdd.n3468 vdd.n636 0.152939
R6578 vdd.n3485 vdd.n636 0.152939
R6579 vdd.n3486 vdd.n3485 0.152939
R6580 vdd.n3487 vdd.n3486 0.152939
R6581 vdd.n3487 vdd.n334 0.152939
R6582 vdd.n3580 vdd.n335 0.152939
R6583 vdd.n346 vdd.n335 0.152939
R6584 vdd.n347 vdd.n346 0.152939
R6585 vdd.n348 vdd.n347 0.152939
R6586 vdd.n355 vdd.n348 0.152939
R6587 vdd.n356 vdd.n355 0.152939
R6588 vdd.n357 vdd.n356 0.152939
R6589 vdd.n358 vdd.n357 0.152939
R6590 vdd.n366 vdd.n358 0.152939
R6591 vdd.n367 vdd.n366 0.152939
R6592 vdd.n368 vdd.n367 0.152939
R6593 vdd.n369 vdd.n368 0.152939
R6594 vdd.n377 vdd.n369 0.152939
R6595 vdd.n378 vdd.n377 0.152939
R6596 vdd.n379 vdd.n378 0.152939
R6597 vdd.n380 vdd.n379 0.152939
R6598 vdd.n388 vdd.n380 0.152939
R6599 vdd.n389 vdd.n388 0.152939
R6600 vdd.n390 vdd.n389 0.152939
R6601 vdd.n391 vdd.n390 0.152939
R6602 vdd.n464 vdd.n463 0.152939
R6603 vdd.n470 vdd.n463 0.152939
R6604 vdd.n471 vdd.n470 0.152939
R6605 vdd.n472 vdd.n471 0.152939
R6606 vdd.n472 vdd.n461 0.152939
R6607 vdd.n480 vdd.n461 0.152939
R6608 vdd.n481 vdd.n480 0.152939
R6609 vdd.n482 vdd.n481 0.152939
R6610 vdd.n482 vdd.n459 0.152939
R6611 vdd.n490 vdd.n459 0.152939
R6612 vdd.n491 vdd.n490 0.152939
R6613 vdd.n492 vdd.n491 0.152939
R6614 vdd.n492 vdd.n457 0.152939
R6615 vdd.n500 vdd.n457 0.152939
R6616 vdd.n501 vdd.n500 0.152939
R6617 vdd.n502 vdd.n501 0.152939
R6618 vdd.n502 vdd.n455 0.152939
R6619 vdd.n510 vdd.n455 0.152939
R6620 vdd.n511 vdd.n510 0.152939
R6621 vdd.n512 vdd.n511 0.152939
R6622 vdd.n512 vdd.n451 0.152939
R6623 vdd.n520 vdd.n451 0.152939
R6624 vdd.n521 vdd.n520 0.152939
R6625 vdd.n522 vdd.n521 0.152939
R6626 vdd.n522 vdd.n449 0.152939
R6627 vdd.n530 vdd.n449 0.152939
R6628 vdd.n531 vdd.n530 0.152939
R6629 vdd.n532 vdd.n531 0.152939
R6630 vdd.n532 vdd.n447 0.152939
R6631 vdd.n540 vdd.n447 0.152939
R6632 vdd.n541 vdd.n540 0.152939
R6633 vdd.n542 vdd.n541 0.152939
R6634 vdd.n542 vdd.n445 0.152939
R6635 vdd.n550 vdd.n445 0.152939
R6636 vdd.n551 vdd.n550 0.152939
R6637 vdd.n552 vdd.n551 0.152939
R6638 vdd.n552 vdd.n443 0.152939
R6639 vdd.n560 vdd.n443 0.152939
R6640 vdd.n561 vdd.n560 0.152939
R6641 vdd.n562 vdd.n561 0.152939
R6642 vdd.n562 vdd.n439 0.152939
R6643 vdd.n570 vdd.n439 0.152939
R6644 vdd.n571 vdd.n570 0.152939
R6645 vdd.n572 vdd.n571 0.152939
R6646 vdd.n572 vdd.n437 0.152939
R6647 vdd.n580 vdd.n437 0.152939
R6648 vdd.n581 vdd.n580 0.152939
R6649 vdd.n582 vdd.n581 0.152939
R6650 vdd.n582 vdd.n435 0.152939
R6651 vdd.n590 vdd.n435 0.152939
R6652 vdd.n591 vdd.n590 0.152939
R6653 vdd.n592 vdd.n591 0.152939
R6654 vdd.n592 vdd.n433 0.152939
R6655 vdd.n600 vdd.n433 0.152939
R6656 vdd.n601 vdd.n600 0.152939
R6657 vdd.n602 vdd.n601 0.152939
R6658 vdd.n602 vdd.n431 0.152939
R6659 vdd.n610 vdd.n431 0.152939
R6660 vdd.n611 vdd.n610 0.152939
R6661 vdd.n612 vdd.n611 0.152939
R6662 vdd.n612 vdd.n429 0.152939
R6663 vdd.n619 vdd.n429 0.152939
R6664 vdd.n3532 vdd.n619 0.152939
R6665 vdd.n3410 vdd.n3409 0.152939
R6666 vdd.n3410 vdd.n675 0.152939
R6667 vdd.n3424 vdd.n675 0.152939
R6668 vdd.n3425 vdd.n3424 0.152939
R6669 vdd.n3426 vdd.n3425 0.152939
R6670 vdd.n3426 vdd.n665 0.152939
R6671 vdd.n3441 vdd.n665 0.152939
R6672 vdd.n3442 vdd.n3441 0.152939
R6673 vdd.n3443 vdd.n3442 0.152939
R6674 vdd.n3443 vdd.n652 0.152939
R6675 vdd.n3457 vdd.n652 0.152939
R6676 vdd.n3458 vdd.n3457 0.152939
R6677 vdd.n3459 vdd.n3458 0.152939
R6678 vdd.n3459 vdd.n641 0.152939
R6679 vdd.n3474 vdd.n641 0.152939
R6680 vdd.n3475 vdd.n3474 0.152939
R6681 vdd.n3476 vdd.n3475 0.152939
R6682 vdd.n3478 vdd.n3476 0.152939
R6683 vdd.n3478 vdd.n3477 0.152939
R6684 vdd.n3477 vdd.n630 0.152939
R6685 vdd.n3495 vdd.n630 0.152939
R6686 vdd.n3496 vdd.n3495 0.152939
R6687 vdd.n3497 vdd.n3496 0.152939
R6688 vdd.n3497 vdd.n628 0.152939
R6689 vdd.n3502 vdd.n628 0.152939
R6690 vdd.n3503 vdd.n3502 0.152939
R6691 vdd.n3504 vdd.n3503 0.152939
R6692 vdd.n3504 vdd.n626 0.152939
R6693 vdd.n3509 vdd.n626 0.152939
R6694 vdd.n3510 vdd.n3509 0.152939
R6695 vdd.n3511 vdd.n3510 0.152939
R6696 vdd.n3511 vdd.n624 0.152939
R6697 vdd.n3517 vdd.n624 0.152939
R6698 vdd.n3518 vdd.n3517 0.152939
R6699 vdd.n3519 vdd.n3518 0.152939
R6700 vdd.n3519 vdd.n622 0.152939
R6701 vdd.n3524 vdd.n622 0.152939
R6702 vdd.n3525 vdd.n3524 0.152939
R6703 vdd.n3526 vdd.n3525 0.152939
R6704 vdd.n3526 vdd.n620 0.152939
R6705 vdd.n3531 vdd.n620 0.152939
R6706 vdd.n3408 vdd.n687 0.152939
R6707 vdd.n2204 vdd.n1147 0.152939
R6708 vdd.n1510 vdd.n1266 0.152939
R6709 vdd.n1511 vdd.n1510 0.152939
R6710 vdd.n1512 vdd.n1511 0.152939
R6711 vdd.n1512 vdd.n1254 0.152939
R6712 vdd.n1527 vdd.n1254 0.152939
R6713 vdd.n1528 vdd.n1527 0.152939
R6714 vdd.n1529 vdd.n1528 0.152939
R6715 vdd.n1529 vdd.n1244 0.152939
R6716 vdd.n1544 vdd.n1244 0.152939
R6717 vdd.n1545 vdd.n1544 0.152939
R6718 vdd.n1546 vdd.n1545 0.152939
R6719 vdd.n1546 vdd.n1231 0.152939
R6720 vdd.n1560 vdd.n1231 0.152939
R6721 vdd.n1561 vdd.n1560 0.152939
R6722 vdd.n1562 vdd.n1561 0.152939
R6723 vdd.n1562 vdd.n1220 0.152939
R6724 vdd.n1577 vdd.n1220 0.152939
R6725 vdd.n1578 vdd.n1577 0.152939
R6726 vdd.n1579 vdd.n1578 0.152939
R6727 vdd.n1579 vdd.n1209 0.152939
R6728 vdd.n1900 vdd.n1209 0.152939
R6729 vdd.n1901 vdd.n1900 0.152939
R6730 vdd.n1902 vdd.n1901 0.152939
R6731 vdd.n1902 vdd.n1197 0.152939
R6732 vdd.n1917 vdd.n1197 0.152939
R6733 vdd.n1918 vdd.n1917 0.152939
R6734 vdd.n1919 vdd.n1918 0.152939
R6735 vdd.n1919 vdd.n1187 0.152939
R6736 vdd.n1934 vdd.n1187 0.152939
R6737 vdd.n1935 vdd.n1934 0.152939
R6738 vdd.n1936 vdd.n1935 0.152939
R6739 vdd.n1936 vdd.n1174 0.152939
R6740 vdd.n1950 vdd.n1174 0.152939
R6741 vdd.n1951 vdd.n1950 0.152939
R6742 vdd.n1952 vdd.n1951 0.152939
R6743 vdd.n1952 vdd.n1164 0.152939
R6744 vdd.n1967 vdd.n1164 0.152939
R6745 vdd.n1968 vdd.n1967 0.152939
R6746 vdd.n1971 vdd.n1968 0.152939
R6747 vdd.n1971 vdd.n1970 0.152939
R6748 vdd.n1970 vdd.n1969 0.152939
R6749 vdd.n1502 vdd.n1271 0.152939
R6750 vdd.n1495 vdd.n1271 0.152939
R6751 vdd.n1495 vdd.n1494 0.152939
R6752 vdd.n1494 vdd.n1493 0.152939
R6753 vdd.n1493 vdd.n1308 0.152939
R6754 vdd.n1489 vdd.n1308 0.152939
R6755 vdd.n1489 vdd.n1488 0.152939
R6756 vdd.n1488 vdd.n1487 0.152939
R6757 vdd.n1487 vdd.n1314 0.152939
R6758 vdd.n1483 vdd.n1314 0.152939
R6759 vdd.n1483 vdd.n1482 0.152939
R6760 vdd.n1482 vdd.n1481 0.152939
R6761 vdd.n1481 vdd.n1320 0.152939
R6762 vdd.n1477 vdd.n1320 0.152939
R6763 vdd.n1477 vdd.n1476 0.152939
R6764 vdd.n1476 vdd.n1475 0.152939
R6765 vdd.n1475 vdd.n1326 0.152939
R6766 vdd.n1471 vdd.n1326 0.152939
R6767 vdd.n1471 vdd.n1470 0.152939
R6768 vdd.n1470 vdd.n1469 0.152939
R6769 vdd.n1469 vdd.n1334 0.152939
R6770 vdd.n1465 vdd.n1334 0.152939
R6771 vdd.n1465 vdd.n1464 0.152939
R6772 vdd.n1464 vdd.n1463 0.152939
R6773 vdd.n1463 vdd.n1340 0.152939
R6774 vdd.n1459 vdd.n1340 0.152939
R6775 vdd.n1459 vdd.n1458 0.152939
R6776 vdd.n1458 vdd.n1457 0.152939
R6777 vdd.n1457 vdd.n1346 0.152939
R6778 vdd.n1453 vdd.n1346 0.152939
R6779 vdd.n1453 vdd.n1452 0.152939
R6780 vdd.n1452 vdd.n1451 0.152939
R6781 vdd.n1451 vdd.n1352 0.152939
R6782 vdd.n1447 vdd.n1352 0.152939
R6783 vdd.n1447 vdd.n1446 0.152939
R6784 vdd.n1446 vdd.n1445 0.152939
R6785 vdd.n1445 vdd.n1358 0.152939
R6786 vdd.n1441 vdd.n1358 0.152939
R6787 vdd.n1441 vdd.n1440 0.152939
R6788 vdd.n1440 vdd.n1439 0.152939
R6789 vdd.n1439 vdd.n1364 0.152939
R6790 vdd.n1432 vdd.n1364 0.152939
R6791 vdd.n1432 vdd.n1431 0.152939
R6792 vdd.n1431 vdd.n1430 0.152939
R6793 vdd.n1430 vdd.n1369 0.152939
R6794 vdd.n1426 vdd.n1369 0.152939
R6795 vdd.n1426 vdd.n1425 0.152939
R6796 vdd.n1425 vdd.n1424 0.152939
R6797 vdd.n1424 vdd.n1375 0.152939
R6798 vdd.n1420 vdd.n1375 0.152939
R6799 vdd.n1420 vdd.n1419 0.152939
R6800 vdd.n1419 vdd.n1418 0.152939
R6801 vdd.n1418 vdd.n1381 0.152939
R6802 vdd.n1414 vdd.n1381 0.152939
R6803 vdd.n1414 vdd.n1413 0.152939
R6804 vdd.n1413 vdd.n1412 0.152939
R6805 vdd.n1412 vdd.n1387 0.152939
R6806 vdd.n1408 vdd.n1387 0.152939
R6807 vdd.n1408 vdd.n1407 0.152939
R6808 vdd.n1407 vdd.n1406 0.152939
R6809 vdd.n1406 vdd.n1393 0.152939
R6810 vdd.n1402 vdd.n1393 0.152939
R6811 vdd.n1402 vdd.n1401 0.152939
R6812 vdd.n1504 vdd.n1503 0.152939
R6813 vdd.n1504 vdd.n1260 0.152939
R6814 vdd.n1519 vdd.n1260 0.152939
R6815 vdd.n1520 vdd.n1519 0.152939
R6816 vdd.n1521 vdd.n1520 0.152939
R6817 vdd.n1521 vdd.n1249 0.152939
R6818 vdd.n1536 vdd.n1249 0.152939
R6819 vdd.n1537 vdd.n1536 0.152939
R6820 vdd.n1538 vdd.n1537 0.152939
R6821 vdd.n1538 vdd.n1238 0.152939
R6822 vdd.n1552 vdd.n1238 0.152939
R6823 vdd.n1553 vdd.n1552 0.152939
R6824 vdd.n1554 vdd.n1553 0.152939
R6825 vdd.n1554 vdd.n1226 0.152939
R6826 vdd.n1569 vdd.n1226 0.152939
R6827 vdd.n1570 vdd.n1569 0.152939
R6828 vdd.n1571 vdd.n1570 0.152939
R6829 vdd.n1571 vdd.n1215 0.152939
R6830 vdd.n1585 vdd.n1215 0.152939
R6831 vdd.n1586 vdd.n1585 0.152939
R6832 vdd.n1507 vdd.t106 0.113865
R6833 vdd.n2491 vdd.t17 0.113865
R6834 vdd.n2558 vdd.t44 0.113865
R6835 vdd.n3041 vdd.t46 0.113865
R6836 vdd.n3108 vdd.t19 0.113865
R6837 vdd.t76 vdd.n386 0.113865
R6838 vdd.n2182 vdd.n1980 0.110256
R6839 vdd.n3398 vdd.n727 0.110256
R6840 vdd.n3275 vdd.n687 0.110256
R6841 vdd.n2205 vdd.n2204 0.110256
R6842 vdd.n1894 vdd.n1893 0.0695946
R6843 vdd.n3581 vdd.n334 0.0695946
R6844 vdd.n3581 vdd.n3580 0.0695946
R6845 vdd.n1893 vdd.n1586 0.0695946
R6846 vdd.n2182 vdd.n2181 0.0431829
R6847 vdd.n2205 vdd.n1144 0.0431829
R6848 vdd.n3398 vdd.n730 0.0431829
R6849 vdd.n3275 vdd.n783 0.0431829
R6850 vdd vdd.n28 0.00833333
R6851 CSoutput.n19 CSoutput.t202 184.661
R6852 CSoutput.n78 CSoutput.n77 165.8
R6853 CSoutput.n76 CSoutput.n0 165.8
R6854 CSoutput.n75 CSoutput.n74 165.8
R6855 CSoutput.n73 CSoutput.n72 165.8
R6856 CSoutput.n71 CSoutput.n2 165.8
R6857 CSoutput.n69 CSoutput.n68 165.8
R6858 CSoutput.n67 CSoutput.n3 165.8
R6859 CSoutput.n66 CSoutput.n65 165.8
R6860 CSoutput.n63 CSoutput.n4 165.8
R6861 CSoutput.n61 CSoutput.n60 165.8
R6862 CSoutput.n59 CSoutput.n5 165.8
R6863 CSoutput.n58 CSoutput.n57 165.8
R6864 CSoutput.n55 CSoutput.n6 165.8
R6865 CSoutput.n54 CSoutput.n53 165.8
R6866 CSoutput.n52 CSoutput.n51 165.8
R6867 CSoutput.n50 CSoutput.n8 165.8
R6868 CSoutput.n48 CSoutput.n47 165.8
R6869 CSoutput.n46 CSoutput.n9 165.8
R6870 CSoutput.n45 CSoutput.n44 165.8
R6871 CSoutput.n42 CSoutput.n10 165.8
R6872 CSoutput.n41 CSoutput.n40 165.8
R6873 CSoutput.n39 CSoutput.n38 165.8
R6874 CSoutput.n37 CSoutput.n12 165.8
R6875 CSoutput.n35 CSoutput.n34 165.8
R6876 CSoutput.n33 CSoutput.n13 165.8
R6877 CSoutput.n32 CSoutput.n31 165.8
R6878 CSoutput.n29 CSoutput.n14 165.8
R6879 CSoutput.n28 CSoutput.n27 165.8
R6880 CSoutput.n26 CSoutput.n25 165.8
R6881 CSoutput.n24 CSoutput.n16 165.8
R6882 CSoutput.n22 CSoutput.n21 165.8
R6883 CSoutput.n20 CSoutput.n17 165.8
R6884 CSoutput.n77 CSoutput.t204 162.194
R6885 CSoutput.n18 CSoutput.t197 120.501
R6886 CSoutput.n23 CSoutput.t192 120.501
R6887 CSoutput.n15 CSoutput.t205 120.501
R6888 CSoutput.n30 CSoutput.t198 120.501
R6889 CSoutput.n36 CSoutput.t200 120.501
R6890 CSoutput.n11 CSoutput.t209 120.501
R6891 CSoutput.n43 CSoutput.t211 120.501
R6892 CSoutput.n49 CSoutput.t203 120.501
R6893 CSoutput.n7 CSoutput.t193 120.501
R6894 CSoutput.n56 CSoutput.t212 120.501
R6895 CSoutput.n62 CSoutput.t208 120.501
R6896 CSoutput.n64 CSoutput.t201 120.501
R6897 CSoutput.n70 CSoutput.t195 120.501
R6898 CSoutput.n1 CSoutput.t210 120.501
R6899 CSoutput.n330 CSoutput.n328 103.469
R6900 CSoutput.n310 CSoutput.n308 103.469
R6901 CSoutput.n291 CSoutput.n289 103.469
R6902 CSoutput.n120 CSoutput.n118 103.469
R6903 CSoutput.n100 CSoutput.n98 103.469
R6904 CSoutput.n81 CSoutput.n79 103.469
R6905 CSoutput.n344 CSoutput.n343 103.111
R6906 CSoutput.n342 CSoutput.n341 103.111
R6907 CSoutput.n340 CSoutput.n339 103.111
R6908 CSoutput.n338 CSoutput.n337 103.111
R6909 CSoutput.n336 CSoutput.n335 103.111
R6910 CSoutput.n334 CSoutput.n333 103.111
R6911 CSoutput.n332 CSoutput.n331 103.111
R6912 CSoutput.n330 CSoutput.n329 103.111
R6913 CSoutput.n326 CSoutput.n325 103.111
R6914 CSoutput.n324 CSoutput.n323 103.111
R6915 CSoutput.n322 CSoutput.n321 103.111
R6916 CSoutput.n320 CSoutput.n319 103.111
R6917 CSoutput.n318 CSoutput.n317 103.111
R6918 CSoutput.n316 CSoutput.n315 103.111
R6919 CSoutput.n314 CSoutput.n313 103.111
R6920 CSoutput.n312 CSoutput.n311 103.111
R6921 CSoutput.n310 CSoutput.n309 103.111
R6922 CSoutput.n307 CSoutput.n306 103.111
R6923 CSoutput.n305 CSoutput.n304 103.111
R6924 CSoutput.n303 CSoutput.n302 103.111
R6925 CSoutput.n301 CSoutput.n300 103.111
R6926 CSoutput.n299 CSoutput.n298 103.111
R6927 CSoutput.n297 CSoutput.n296 103.111
R6928 CSoutput.n295 CSoutput.n294 103.111
R6929 CSoutput.n293 CSoutput.n292 103.111
R6930 CSoutput.n291 CSoutput.n290 103.111
R6931 CSoutput.n120 CSoutput.n119 103.111
R6932 CSoutput.n122 CSoutput.n121 103.111
R6933 CSoutput.n124 CSoutput.n123 103.111
R6934 CSoutput.n126 CSoutput.n125 103.111
R6935 CSoutput.n128 CSoutput.n127 103.111
R6936 CSoutput.n130 CSoutput.n129 103.111
R6937 CSoutput.n132 CSoutput.n131 103.111
R6938 CSoutput.n134 CSoutput.n133 103.111
R6939 CSoutput.n136 CSoutput.n135 103.111
R6940 CSoutput.n100 CSoutput.n99 103.111
R6941 CSoutput.n102 CSoutput.n101 103.111
R6942 CSoutput.n104 CSoutput.n103 103.111
R6943 CSoutput.n106 CSoutput.n105 103.111
R6944 CSoutput.n108 CSoutput.n107 103.111
R6945 CSoutput.n110 CSoutput.n109 103.111
R6946 CSoutput.n112 CSoutput.n111 103.111
R6947 CSoutput.n114 CSoutput.n113 103.111
R6948 CSoutput.n116 CSoutput.n115 103.111
R6949 CSoutput.n81 CSoutput.n80 103.111
R6950 CSoutput.n83 CSoutput.n82 103.111
R6951 CSoutput.n85 CSoutput.n84 103.111
R6952 CSoutput.n87 CSoutput.n86 103.111
R6953 CSoutput.n89 CSoutput.n88 103.111
R6954 CSoutput.n91 CSoutput.n90 103.111
R6955 CSoutput.n93 CSoutput.n92 103.111
R6956 CSoutput.n95 CSoutput.n94 103.111
R6957 CSoutput.n97 CSoutput.n96 103.111
R6958 CSoutput.n346 CSoutput.n345 103.111
R6959 CSoutput.n374 CSoutput.n372 81.5057
R6960 CSoutput.n362 CSoutput.n360 81.5057
R6961 CSoutput.n351 CSoutput.n349 81.5057
R6962 CSoutput.n410 CSoutput.n408 81.5057
R6963 CSoutput.n398 CSoutput.n396 81.5057
R6964 CSoutput.n387 CSoutput.n385 81.5057
R6965 CSoutput.n382 CSoutput.n381 80.9324
R6966 CSoutput.n380 CSoutput.n379 80.9324
R6967 CSoutput.n378 CSoutput.n377 80.9324
R6968 CSoutput.n376 CSoutput.n375 80.9324
R6969 CSoutput.n374 CSoutput.n373 80.9324
R6970 CSoutput.n370 CSoutput.n369 80.9324
R6971 CSoutput.n368 CSoutput.n367 80.9324
R6972 CSoutput.n366 CSoutput.n365 80.9324
R6973 CSoutput.n364 CSoutput.n363 80.9324
R6974 CSoutput.n362 CSoutput.n361 80.9324
R6975 CSoutput.n359 CSoutput.n358 80.9324
R6976 CSoutput.n357 CSoutput.n356 80.9324
R6977 CSoutput.n355 CSoutput.n354 80.9324
R6978 CSoutput.n353 CSoutput.n352 80.9324
R6979 CSoutput.n351 CSoutput.n350 80.9324
R6980 CSoutput.n410 CSoutput.n409 80.9324
R6981 CSoutput.n412 CSoutput.n411 80.9324
R6982 CSoutput.n414 CSoutput.n413 80.9324
R6983 CSoutput.n416 CSoutput.n415 80.9324
R6984 CSoutput.n418 CSoutput.n417 80.9324
R6985 CSoutput.n398 CSoutput.n397 80.9324
R6986 CSoutput.n400 CSoutput.n399 80.9324
R6987 CSoutput.n402 CSoutput.n401 80.9324
R6988 CSoutput.n404 CSoutput.n403 80.9324
R6989 CSoutput.n406 CSoutput.n405 80.9324
R6990 CSoutput.n387 CSoutput.n386 80.9324
R6991 CSoutput.n389 CSoutput.n388 80.9324
R6992 CSoutput.n391 CSoutput.n390 80.9324
R6993 CSoutput.n393 CSoutput.n392 80.9324
R6994 CSoutput.n395 CSoutput.n394 80.9324
R6995 CSoutput.n25 CSoutput.n24 48.1486
R6996 CSoutput.n69 CSoutput.n3 48.1486
R6997 CSoutput.n38 CSoutput.n37 48.1486
R6998 CSoutput.n42 CSoutput.n41 48.1486
R6999 CSoutput.n51 CSoutput.n50 48.1486
R7000 CSoutput.n55 CSoutput.n54 48.1486
R7001 CSoutput.n22 CSoutput.n17 46.462
R7002 CSoutput.n72 CSoutput.n71 46.462
R7003 CSoutput.n20 CSoutput.n19 44.9055
R7004 CSoutput.n29 CSoutput.n28 43.7635
R7005 CSoutput.n65 CSoutput.n63 43.7635
R7006 CSoutput.n35 CSoutput.n13 41.7396
R7007 CSoutput.n57 CSoutput.n5 41.7396
R7008 CSoutput.n44 CSoutput.n9 37.0171
R7009 CSoutput.n48 CSoutput.n9 37.0171
R7010 CSoutput.n76 CSoutput.n75 34.9932
R7011 CSoutput.n31 CSoutput.n13 32.2947
R7012 CSoutput.n61 CSoutput.n5 32.2947
R7013 CSoutput.n30 CSoutput.n29 29.6014
R7014 CSoutput.n63 CSoutput.n62 29.6014
R7015 CSoutput.n19 CSoutput.n18 28.4085
R7016 CSoutput.n18 CSoutput.n17 25.1176
R7017 CSoutput.n72 CSoutput.n1 25.1176
R7018 CSoutput.n43 CSoutput.n42 22.0922
R7019 CSoutput.n50 CSoutput.n49 22.0922
R7020 CSoutput.n77 CSoutput.n76 21.8586
R7021 CSoutput.n37 CSoutput.n36 18.9681
R7022 CSoutput.n56 CSoutput.n55 18.9681
R7023 CSoutput.n25 CSoutput.n15 17.6292
R7024 CSoutput.n64 CSoutput.n3 17.6292
R7025 CSoutput.n24 CSoutput.n23 15.844
R7026 CSoutput.n70 CSoutput.n69 15.844
R7027 CSoutput.n38 CSoutput.n11 14.5051
R7028 CSoutput.n54 CSoutput.n7 14.5051
R7029 CSoutput.n421 CSoutput.n78 11.4997
R7030 CSoutput.n41 CSoutput.n11 11.3811
R7031 CSoutput.n51 CSoutput.n7 11.3811
R7032 CSoutput.n23 CSoutput.n22 10.0422
R7033 CSoutput.n71 CSoutput.n70 10.0422
R7034 CSoutput.n327 CSoutput.n307 9.25285
R7035 CSoutput.n117 CSoutput.n97 9.25285
R7036 CSoutput.n371 CSoutput.n359 8.98182
R7037 CSoutput.n407 CSoutput.n395 8.98182
R7038 CSoutput.n384 CSoutput.n348 8.61339
R7039 CSoutput.n28 CSoutput.n15 8.25698
R7040 CSoutput.n65 CSoutput.n64 8.25698
R7041 CSoutput.n348 CSoutput.n347 7.12641
R7042 CSoutput.n138 CSoutput.n137 7.12641
R7043 CSoutput.n36 CSoutput.n35 6.91809
R7044 CSoutput.n57 CSoutput.n56 6.91809
R7045 CSoutput.n384 CSoutput.n383 6.02792
R7046 CSoutput.n420 CSoutput.n419 6.02792
R7047 CSoutput.n383 CSoutput.n382 5.25266
R7048 CSoutput.n371 CSoutput.n370 5.25266
R7049 CSoutput.n419 CSoutput.n418 5.25266
R7050 CSoutput.n407 CSoutput.n406 5.25266
R7051 CSoutput.n347 CSoutput.n346 5.1449
R7052 CSoutput.n327 CSoutput.n326 5.1449
R7053 CSoutput.n137 CSoutput.n136 5.1449
R7054 CSoutput.n117 CSoutput.n116 5.1449
R7055 CSoutput.n421 CSoutput.n138 4.91834
R7056 CSoutput.n229 CSoutput.n182 4.5005
R7057 CSoutput.n198 CSoutput.n182 4.5005
R7058 CSoutput.n193 CSoutput.n177 4.5005
R7059 CSoutput.n193 CSoutput.n179 4.5005
R7060 CSoutput.n193 CSoutput.n176 4.5005
R7061 CSoutput.n193 CSoutput.n180 4.5005
R7062 CSoutput.n193 CSoutput.n175 4.5005
R7063 CSoutput.n193 CSoutput.t206 4.5005
R7064 CSoutput.n193 CSoutput.n174 4.5005
R7065 CSoutput.n193 CSoutput.n181 4.5005
R7066 CSoutput.n193 CSoutput.n182 4.5005
R7067 CSoutput.n191 CSoutput.n177 4.5005
R7068 CSoutput.n191 CSoutput.n179 4.5005
R7069 CSoutput.n191 CSoutput.n176 4.5005
R7070 CSoutput.n191 CSoutput.n180 4.5005
R7071 CSoutput.n191 CSoutput.n175 4.5005
R7072 CSoutput.n191 CSoutput.t206 4.5005
R7073 CSoutput.n191 CSoutput.n174 4.5005
R7074 CSoutput.n191 CSoutput.n181 4.5005
R7075 CSoutput.n191 CSoutput.n182 4.5005
R7076 CSoutput.n190 CSoutput.n177 4.5005
R7077 CSoutput.n190 CSoutput.n179 4.5005
R7078 CSoutput.n190 CSoutput.n176 4.5005
R7079 CSoutput.n190 CSoutput.n180 4.5005
R7080 CSoutput.n190 CSoutput.n175 4.5005
R7081 CSoutput.n190 CSoutput.t206 4.5005
R7082 CSoutput.n190 CSoutput.n174 4.5005
R7083 CSoutput.n190 CSoutput.n181 4.5005
R7084 CSoutput.n190 CSoutput.n182 4.5005
R7085 CSoutput.n275 CSoutput.n177 4.5005
R7086 CSoutput.n275 CSoutput.n179 4.5005
R7087 CSoutput.n275 CSoutput.n176 4.5005
R7088 CSoutput.n275 CSoutput.n180 4.5005
R7089 CSoutput.n275 CSoutput.n175 4.5005
R7090 CSoutput.n275 CSoutput.t206 4.5005
R7091 CSoutput.n275 CSoutput.n174 4.5005
R7092 CSoutput.n275 CSoutput.n181 4.5005
R7093 CSoutput.n275 CSoutput.n182 4.5005
R7094 CSoutput.n273 CSoutput.n177 4.5005
R7095 CSoutput.n273 CSoutput.n179 4.5005
R7096 CSoutput.n273 CSoutput.n176 4.5005
R7097 CSoutput.n273 CSoutput.n180 4.5005
R7098 CSoutput.n273 CSoutput.n175 4.5005
R7099 CSoutput.n273 CSoutput.t206 4.5005
R7100 CSoutput.n273 CSoutput.n174 4.5005
R7101 CSoutput.n273 CSoutput.n181 4.5005
R7102 CSoutput.n271 CSoutput.n177 4.5005
R7103 CSoutput.n271 CSoutput.n179 4.5005
R7104 CSoutput.n271 CSoutput.n176 4.5005
R7105 CSoutput.n271 CSoutput.n180 4.5005
R7106 CSoutput.n271 CSoutput.n175 4.5005
R7107 CSoutput.n271 CSoutput.t206 4.5005
R7108 CSoutput.n271 CSoutput.n174 4.5005
R7109 CSoutput.n271 CSoutput.n181 4.5005
R7110 CSoutput.n201 CSoutput.n177 4.5005
R7111 CSoutput.n201 CSoutput.n179 4.5005
R7112 CSoutput.n201 CSoutput.n176 4.5005
R7113 CSoutput.n201 CSoutput.n180 4.5005
R7114 CSoutput.n201 CSoutput.n175 4.5005
R7115 CSoutput.n201 CSoutput.t206 4.5005
R7116 CSoutput.n201 CSoutput.n174 4.5005
R7117 CSoutput.n201 CSoutput.n181 4.5005
R7118 CSoutput.n201 CSoutput.n182 4.5005
R7119 CSoutput.n200 CSoutput.n177 4.5005
R7120 CSoutput.n200 CSoutput.n179 4.5005
R7121 CSoutput.n200 CSoutput.n176 4.5005
R7122 CSoutput.n200 CSoutput.n180 4.5005
R7123 CSoutput.n200 CSoutput.n175 4.5005
R7124 CSoutput.n200 CSoutput.t206 4.5005
R7125 CSoutput.n200 CSoutput.n174 4.5005
R7126 CSoutput.n200 CSoutput.n181 4.5005
R7127 CSoutput.n200 CSoutput.n182 4.5005
R7128 CSoutput.n204 CSoutput.n177 4.5005
R7129 CSoutput.n204 CSoutput.n179 4.5005
R7130 CSoutput.n204 CSoutput.n176 4.5005
R7131 CSoutput.n204 CSoutput.n180 4.5005
R7132 CSoutput.n204 CSoutput.n175 4.5005
R7133 CSoutput.n204 CSoutput.t206 4.5005
R7134 CSoutput.n204 CSoutput.n174 4.5005
R7135 CSoutput.n204 CSoutput.n181 4.5005
R7136 CSoutput.n204 CSoutput.n182 4.5005
R7137 CSoutput.n203 CSoutput.n177 4.5005
R7138 CSoutput.n203 CSoutput.n179 4.5005
R7139 CSoutput.n203 CSoutput.n176 4.5005
R7140 CSoutput.n203 CSoutput.n180 4.5005
R7141 CSoutput.n203 CSoutput.n175 4.5005
R7142 CSoutput.n203 CSoutput.t206 4.5005
R7143 CSoutput.n203 CSoutput.n174 4.5005
R7144 CSoutput.n203 CSoutput.n181 4.5005
R7145 CSoutput.n203 CSoutput.n182 4.5005
R7146 CSoutput.n186 CSoutput.n177 4.5005
R7147 CSoutput.n186 CSoutput.n179 4.5005
R7148 CSoutput.n186 CSoutput.n176 4.5005
R7149 CSoutput.n186 CSoutput.n180 4.5005
R7150 CSoutput.n186 CSoutput.n175 4.5005
R7151 CSoutput.n186 CSoutput.t206 4.5005
R7152 CSoutput.n186 CSoutput.n174 4.5005
R7153 CSoutput.n186 CSoutput.n181 4.5005
R7154 CSoutput.n186 CSoutput.n182 4.5005
R7155 CSoutput.n278 CSoutput.n177 4.5005
R7156 CSoutput.n278 CSoutput.n179 4.5005
R7157 CSoutput.n278 CSoutput.n176 4.5005
R7158 CSoutput.n278 CSoutput.n180 4.5005
R7159 CSoutput.n278 CSoutput.n175 4.5005
R7160 CSoutput.n278 CSoutput.t206 4.5005
R7161 CSoutput.n278 CSoutput.n174 4.5005
R7162 CSoutput.n278 CSoutput.n181 4.5005
R7163 CSoutput.n278 CSoutput.n182 4.5005
R7164 CSoutput.n265 CSoutput.n236 4.5005
R7165 CSoutput.n265 CSoutput.n242 4.5005
R7166 CSoutput.n223 CSoutput.n212 4.5005
R7167 CSoutput.n223 CSoutput.n214 4.5005
R7168 CSoutput.n223 CSoutput.n211 4.5005
R7169 CSoutput.n223 CSoutput.n215 4.5005
R7170 CSoutput.n223 CSoutput.n210 4.5005
R7171 CSoutput.n223 CSoutput.t196 4.5005
R7172 CSoutput.n223 CSoutput.n209 4.5005
R7173 CSoutput.n223 CSoutput.n216 4.5005
R7174 CSoutput.n265 CSoutput.n223 4.5005
R7175 CSoutput.n244 CSoutput.n212 4.5005
R7176 CSoutput.n244 CSoutput.n214 4.5005
R7177 CSoutput.n244 CSoutput.n211 4.5005
R7178 CSoutput.n244 CSoutput.n215 4.5005
R7179 CSoutput.n244 CSoutput.n210 4.5005
R7180 CSoutput.n244 CSoutput.t196 4.5005
R7181 CSoutput.n244 CSoutput.n209 4.5005
R7182 CSoutput.n244 CSoutput.n216 4.5005
R7183 CSoutput.n265 CSoutput.n244 4.5005
R7184 CSoutput.n222 CSoutput.n212 4.5005
R7185 CSoutput.n222 CSoutput.n214 4.5005
R7186 CSoutput.n222 CSoutput.n211 4.5005
R7187 CSoutput.n222 CSoutput.n215 4.5005
R7188 CSoutput.n222 CSoutput.n210 4.5005
R7189 CSoutput.n222 CSoutput.t196 4.5005
R7190 CSoutput.n222 CSoutput.n209 4.5005
R7191 CSoutput.n222 CSoutput.n216 4.5005
R7192 CSoutput.n265 CSoutput.n222 4.5005
R7193 CSoutput.n246 CSoutput.n212 4.5005
R7194 CSoutput.n246 CSoutput.n214 4.5005
R7195 CSoutput.n246 CSoutput.n211 4.5005
R7196 CSoutput.n246 CSoutput.n215 4.5005
R7197 CSoutput.n246 CSoutput.n210 4.5005
R7198 CSoutput.n246 CSoutput.t196 4.5005
R7199 CSoutput.n246 CSoutput.n209 4.5005
R7200 CSoutput.n246 CSoutput.n216 4.5005
R7201 CSoutput.n265 CSoutput.n246 4.5005
R7202 CSoutput.n212 CSoutput.n207 4.5005
R7203 CSoutput.n214 CSoutput.n207 4.5005
R7204 CSoutput.n211 CSoutput.n207 4.5005
R7205 CSoutput.n215 CSoutput.n207 4.5005
R7206 CSoutput.n210 CSoutput.n207 4.5005
R7207 CSoutput.t196 CSoutput.n207 4.5005
R7208 CSoutput.n209 CSoutput.n207 4.5005
R7209 CSoutput.n216 CSoutput.n207 4.5005
R7210 CSoutput.n268 CSoutput.n212 4.5005
R7211 CSoutput.n268 CSoutput.n214 4.5005
R7212 CSoutput.n268 CSoutput.n211 4.5005
R7213 CSoutput.n268 CSoutput.n215 4.5005
R7214 CSoutput.n268 CSoutput.n210 4.5005
R7215 CSoutput.n268 CSoutput.t196 4.5005
R7216 CSoutput.n268 CSoutput.n209 4.5005
R7217 CSoutput.n268 CSoutput.n216 4.5005
R7218 CSoutput.n266 CSoutput.n212 4.5005
R7219 CSoutput.n266 CSoutput.n214 4.5005
R7220 CSoutput.n266 CSoutput.n211 4.5005
R7221 CSoutput.n266 CSoutput.n215 4.5005
R7222 CSoutput.n266 CSoutput.n210 4.5005
R7223 CSoutput.n266 CSoutput.t196 4.5005
R7224 CSoutput.n266 CSoutput.n209 4.5005
R7225 CSoutput.n266 CSoutput.n216 4.5005
R7226 CSoutput.n266 CSoutput.n265 4.5005
R7227 CSoutput.n248 CSoutput.n212 4.5005
R7228 CSoutput.n248 CSoutput.n214 4.5005
R7229 CSoutput.n248 CSoutput.n211 4.5005
R7230 CSoutput.n248 CSoutput.n215 4.5005
R7231 CSoutput.n248 CSoutput.n210 4.5005
R7232 CSoutput.n248 CSoutput.t196 4.5005
R7233 CSoutput.n248 CSoutput.n209 4.5005
R7234 CSoutput.n248 CSoutput.n216 4.5005
R7235 CSoutput.n265 CSoutput.n248 4.5005
R7236 CSoutput.n220 CSoutput.n212 4.5005
R7237 CSoutput.n220 CSoutput.n214 4.5005
R7238 CSoutput.n220 CSoutput.n211 4.5005
R7239 CSoutput.n220 CSoutput.n215 4.5005
R7240 CSoutput.n220 CSoutput.n210 4.5005
R7241 CSoutput.n220 CSoutput.t196 4.5005
R7242 CSoutput.n220 CSoutput.n209 4.5005
R7243 CSoutput.n220 CSoutput.n216 4.5005
R7244 CSoutput.n265 CSoutput.n220 4.5005
R7245 CSoutput.n250 CSoutput.n212 4.5005
R7246 CSoutput.n250 CSoutput.n214 4.5005
R7247 CSoutput.n250 CSoutput.n211 4.5005
R7248 CSoutput.n250 CSoutput.n215 4.5005
R7249 CSoutput.n250 CSoutput.n210 4.5005
R7250 CSoutput.n250 CSoutput.t196 4.5005
R7251 CSoutput.n250 CSoutput.n209 4.5005
R7252 CSoutput.n250 CSoutput.n216 4.5005
R7253 CSoutput.n265 CSoutput.n250 4.5005
R7254 CSoutput.n219 CSoutput.n212 4.5005
R7255 CSoutput.n219 CSoutput.n214 4.5005
R7256 CSoutput.n219 CSoutput.n211 4.5005
R7257 CSoutput.n219 CSoutput.n215 4.5005
R7258 CSoutput.n219 CSoutput.n210 4.5005
R7259 CSoutput.n219 CSoutput.t196 4.5005
R7260 CSoutput.n219 CSoutput.n209 4.5005
R7261 CSoutput.n219 CSoutput.n216 4.5005
R7262 CSoutput.n265 CSoutput.n219 4.5005
R7263 CSoutput.n264 CSoutput.n212 4.5005
R7264 CSoutput.n264 CSoutput.n214 4.5005
R7265 CSoutput.n264 CSoutput.n211 4.5005
R7266 CSoutput.n264 CSoutput.n215 4.5005
R7267 CSoutput.n264 CSoutput.n210 4.5005
R7268 CSoutput.n264 CSoutput.t196 4.5005
R7269 CSoutput.n264 CSoutput.n209 4.5005
R7270 CSoutput.n264 CSoutput.n216 4.5005
R7271 CSoutput.n265 CSoutput.n264 4.5005
R7272 CSoutput.n263 CSoutput.n148 4.5005
R7273 CSoutput.n164 CSoutput.n148 4.5005
R7274 CSoutput.n159 CSoutput.n143 4.5005
R7275 CSoutput.n159 CSoutput.n145 4.5005
R7276 CSoutput.n159 CSoutput.n142 4.5005
R7277 CSoutput.n159 CSoutput.n146 4.5005
R7278 CSoutput.n159 CSoutput.n141 4.5005
R7279 CSoutput.n159 CSoutput.t199 4.5005
R7280 CSoutput.n159 CSoutput.n140 4.5005
R7281 CSoutput.n159 CSoutput.n147 4.5005
R7282 CSoutput.n159 CSoutput.n148 4.5005
R7283 CSoutput.n157 CSoutput.n143 4.5005
R7284 CSoutput.n157 CSoutput.n145 4.5005
R7285 CSoutput.n157 CSoutput.n142 4.5005
R7286 CSoutput.n157 CSoutput.n146 4.5005
R7287 CSoutput.n157 CSoutput.n141 4.5005
R7288 CSoutput.n157 CSoutput.t199 4.5005
R7289 CSoutput.n157 CSoutput.n140 4.5005
R7290 CSoutput.n157 CSoutput.n147 4.5005
R7291 CSoutput.n157 CSoutput.n148 4.5005
R7292 CSoutput.n156 CSoutput.n143 4.5005
R7293 CSoutput.n156 CSoutput.n145 4.5005
R7294 CSoutput.n156 CSoutput.n142 4.5005
R7295 CSoutput.n156 CSoutput.n146 4.5005
R7296 CSoutput.n156 CSoutput.n141 4.5005
R7297 CSoutput.n156 CSoutput.t199 4.5005
R7298 CSoutput.n156 CSoutput.n140 4.5005
R7299 CSoutput.n156 CSoutput.n147 4.5005
R7300 CSoutput.n156 CSoutput.n148 4.5005
R7301 CSoutput.n285 CSoutput.n143 4.5005
R7302 CSoutput.n285 CSoutput.n145 4.5005
R7303 CSoutput.n285 CSoutput.n142 4.5005
R7304 CSoutput.n285 CSoutput.n146 4.5005
R7305 CSoutput.n285 CSoutput.n141 4.5005
R7306 CSoutput.n285 CSoutput.t199 4.5005
R7307 CSoutput.n285 CSoutput.n140 4.5005
R7308 CSoutput.n285 CSoutput.n147 4.5005
R7309 CSoutput.n285 CSoutput.n148 4.5005
R7310 CSoutput.n283 CSoutput.n143 4.5005
R7311 CSoutput.n283 CSoutput.n145 4.5005
R7312 CSoutput.n283 CSoutput.n142 4.5005
R7313 CSoutput.n283 CSoutput.n146 4.5005
R7314 CSoutput.n283 CSoutput.n141 4.5005
R7315 CSoutput.n283 CSoutput.t199 4.5005
R7316 CSoutput.n283 CSoutput.n140 4.5005
R7317 CSoutput.n283 CSoutput.n147 4.5005
R7318 CSoutput.n281 CSoutput.n143 4.5005
R7319 CSoutput.n281 CSoutput.n145 4.5005
R7320 CSoutput.n281 CSoutput.n142 4.5005
R7321 CSoutput.n281 CSoutput.n146 4.5005
R7322 CSoutput.n281 CSoutput.n141 4.5005
R7323 CSoutput.n281 CSoutput.t199 4.5005
R7324 CSoutput.n281 CSoutput.n140 4.5005
R7325 CSoutput.n281 CSoutput.n147 4.5005
R7326 CSoutput.n167 CSoutput.n143 4.5005
R7327 CSoutput.n167 CSoutput.n145 4.5005
R7328 CSoutput.n167 CSoutput.n142 4.5005
R7329 CSoutput.n167 CSoutput.n146 4.5005
R7330 CSoutput.n167 CSoutput.n141 4.5005
R7331 CSoutput.n167 CSoutput.t199 4.5005
R7332 CSoutput.n167 CSoutput.n140 4.5005
R7333 CSoutput.n167 CSoutput.n147 4.5005
R7334 CSoutput.n167 CSoutput.n148 4.5005
R7335 CSoutput.n166 CSoutput.n143 4.5005
R7336 CSoutput.n166 CSoutput.n145 4.5005
R7337 CSoutput.n166 CSoutput.n142 4.5005
R7338 CSoutput.n166 CSoutput.n146 4.5005
R7339 CSoutput.n166 CSoutput.n141 4.5005
R7340 CSoutput.n166 CSoutput.t199 4.5005
R7341 CSoutput.n166 CSoutput.n140 4.5005
R7342 CSoutput.n166 CSoutput.n147 4.5005
R7343 CSoutput.n166 CSoutput.n148 4.5005
R7344 CSoutput.n170 CSoutput.n143 4.5005
R7345 CSoutput.n170 CSoutput.n145 4.5005
R7346 CSoutput.n170 CSoutput.n142 4.5005
R7347 CSoutput.n170 CSoutput.n146 4.5005
R7348 CSoutput.n170 CSoutput.n141 4.5005
R7349 CSoutput.n170 CSoutput.t199 4.5005
R7350 CSoutput.n170 CSoutput.n140 4.5005
R7351 CSoutput.n170 CSoutput.n147 4.5005
R7352 CSoutput.n170 CSoutput.n148 4.5005
R7353 CSoutput.n169 CSoutput.n143 4.5005
R7354 CSoutput.n169 CSoutput.n145 4.5005
R7355 CSoutput.n169 CSoutput.n142 4.5005
R7356 CSoutput.n169 CSoutput.n146 4.5005
R7357 CSoutput.n169 CSoutput.n141 4.5005
R7358 CSoutput.n169 CSoutput.t199 4.5005
R7359 CSoutput.n169 CSoutput.n140 4.5005
R7360 CSoutput.n169 CSoutput.n147 4.5005
R7361 CSoutput.n169 CSoutput.n148 4.5005
R7362 CSoutput.n152 CSoutput.n143 4.5005
R7363 CSoutput.n152 CSoutput.n145 4.5005
R7364 CSoutput.n152 CSoutput.n142 4.5005
R7365 CSoutput.n152 CSoutput.n146 4.5005
R7366 CSoutput.n152 CSoutput.n141 4.5005
R7367 CSoutput.n152 CSoutput.t199 4.5005
R7368 CSoutput.n152 CSoutput.n140 4.5005
R7369 CSoutput.n152 CSoutput.n147 4.5005
R7370 CSoutput.n152 CSoutput.n148 4.5005
R7371 CSoutput.n288 CSoutput.n143 4.5005
R7372 CSoutput.n288 CSoutput.n145 4.5005
R7373 CSoutput.n288 CSoutput.n142 4.5005
R7374 CSoutput.n288 CSoutput.n146 4.5005
R7375 CSoutput.n288 CSoutput.n141 4.5005
R7376 CSoutput.n288 CSoutput.t199 4.5005
R7377 CSoutput.n288 CSoutput.n140 4.5005
R7378 CSoutput.n288 CSoutput.n147 4.5005
R7379 CSoutput.n288 CSoutput.n148 4.5005
R7380 CSoutput.n347 CSoutput.n327 4.10845
R7381 CSoutput.n137 CSoutput.n117 4.10845
R7382 CSoutput.n345 CSoutput.t170 4.06363
R7383 CSoutput.n345 CSoutput.t82 4.06363
R7384 CSoutput.n343 CSoutput.t106 4.06363
R7385 CSoutput.n343 CSoutput.t133 4.06363
R7386 CSoutput.n341 CSoutput.t150 4.06363
R7387 CSoutput.n341 CSoutput.t67 4.06363
R7388 CSoutput.n339 CSoutput.t61 4.06363
R7389 CSoutput.n339 CSoutput.t109 4.06363
R7390 CSoutput.n337 CSoutput.t127 4.06363
R7391 CSoutput.n337 CSoutput.t152 4.06363
R7392 CSoutput.n335 CSoutput.t167 4.06363
R7393 CSoutput.n335 CSoutput.t79 4.06363
R7394 CSoutput.n333 CSoutput.t85 4.06363
R7395 CSoutput.n333 CSoutput.t153 4.06363
R7396 CSoutput.n331 CSoutput.t169 4.06363
R7397 CSoutput.n331 CSoutput.t171 4.06363
R7398 CSoutput.n329 CSoutput.t105 4.06363
R7399 CSoutput.n329 CSoutput.t107 4.06363
R7400 CSoutput.n328 CSoutput.t111 4.06363
R7401 CSoutput.n328 CSoutput.t175 4.06363
R7402 CSoutput.n325 CSoutput.t159 4.06363
R7403 CSoutput.n325 CSoutput.t68 4.06363
R7404 CSoutput.n323 CSoutput.t88 4.06363
R7405 CSoutput.n323 CSoutput.t125 4.06363
R7406 CSoutput.n321 CSoutput.t140 4.06363
R7407 CSoutput.n321 CSoutput.t176 4.06363
R7408 CSoutput.n319 CSoutput.t168 4.06363
R7409 CSoutput.n319 CSoutput.t94 4.06363
R7410 CSoutput.n317 CSoutput.t114 4.06363
R7411 CSoutput.n317 CSoutput.t141 4.06363
R7412 CSoutput.n315 CSoutput.t154 4.06363
R7413 CSoutput.n315 CSoutput.t66 4.06363
R7414 CSoutput.n313 CSoutput.t69 4.06363
R7415 CSoutput.n313 CSoutput.t144 4.06363
R7416 CSoutput.n311 CSoutput.t160 4.06363
R7417 CSoutput.n311 CSoutput.t161 4.06363
R7418 CSoutput.n309 CSoutput.t87 4.06363
R7419 CSoutput.n309 CSoutput.t89 4.06363
R7420 CSoutput.n308 CSoutput.t95 4.06363
R7421 CSoutput.n308 CSoutput.t163 4.06363
R7422 CSoutput.n306 CSoutput.t172 4.06363
R7423 CSoutput.n306 CSoutput.t126 4.06363
R7424 CSoutput.n304 CSoutput.t157 4.06363
R7425 CSoutput.n304 CSoutput.t110 4.06363
R7426 CSoutput.n302 CSoutput.t142 4.06363
R7427 CSoutput.n302 CSoutput.t92 4.06363
R7428 CSoutput.n300 CSoutput.t164 4.06363
R7429 CSoutput.n300 CSoutput.t118 4.06363
R7430 CSoutput.n298 CSoutput.t151 4.06363
R7431 CSoutput.n298 CSoutput.t102 4.06363
R7432 CSoutput.n296 CSoutput.t137 4.06363
R7433 CSoutput.n296 CSoutput.t78 4.06363
R7434 CSoutput.n294 CSoutput.t155 4.06363
R7435 CSoutput.n294 CSoutput.t73 4.06363
R7436 CSoutput.n292 CSoutput.t115 4.06363
R7437 CSoutput.n292 CSoutput.t90 4.06363
R7438 CSoutput.n290 CSoutput.t96 4.06363
R7439 CSoutput.n290 CSoutput.t70 4.06363
R7440 CSoutput.n289 CSoutput.t149 4.06363
R7441 CSoutput.n289 CSoutput.t63 4.06363
R7442 CSoutput.n118 CSoutput.t104 4.06363
R7443 CSoutput.n118 CSoutput.t178 4.06363
R7444 CSoutput.n119 CSoutput.t147 4.06363
R7445 CSoutput.n119 CSoutput.t145 4.06363
R7446 CSoutput.n121 CSoutput.t130 4.06363
R7447 CSoutput.n121 CSoutput.t100 4.06363
R7448 CSoutput.n123 CSoutput.t77 4.06363
R7449 CSoutput.n123 CSoutput.t132 4.06363
R7450 CSoutput.n125 CSoutput.t129 4.06363
R7451 CSoutput.n125 CSoutput.t97 4.06363
R7452 CSoutput.n127 CSoutput.t76 4.06363
R7453 CSoutput.n127 CSoutput.t75 4.06363
R7454 CSoutput.n129 CSoutput.t148 4.06363
R7455 CSoutput.n129 CSoutput.t113 4.06363
R7456 CSoutput.n131 CSoutput.t108 4.06363
R7457 CSoutput.n131 CSoutput.t71 4.06363
R7458 CSoutput.n133 CSoutput.t174 4.06363
R7459 CSoutput.n133 CSoutput.t146 4.06363
R7460 CSoutput.n135 CSoutput.t131 4.06363
R7461 CSoutput.n135 CSoutput.t101 4.06363
R7462 CSoutput.n98 CSoutput.t86 4.06363
R7463 CSoutput.n98 CSoutput.t166 4.06363
R7464 CSoutput.n99 CSoutput.t136 4.06363
R7465 CSoutput.n99 CSoutput.t134 4.06363
R7466 CSoutput.n101 CSoutput.t120 4.06363
R7467 CSoutput.n101 CSoutput.t83 4.06363
R7468 CSoutput.n103 CSoutput.t64 4.06363
R7469 CSoutput.n103 CSoutput.t122 4.06363
R7470 CSoutput.n105 CSoutput.t117 4.06363
R7471 CSoutput.n105 CSoutput.t80 4.06363
R7472 CSoutput.n107 CSoutput.t62 4.06363
R7473 CSoutput.n107 CSoutput.t60 4.06363
R7474 CSoutput.n109 CSoutput.t139 4.06363
R7475 CSoutput.n109 CSoutput.t99 4.06363
R7476 CSoutput.n111 CSoutput.t93 4.06363
R7477 CSoutput.n111 CSoutput.t59 4.06363
R7478 CSoutput.n113 CSoutput.t162 4.06363
R7479 CSoutput.n113 CSoutput.t135 4.06363
R7480 CSoutput.n115 CSoutput.t121 4.06363
R7481 CSoutput.n115 CSoutput.t84 4.06363
R7482 CSoutput.n79 CSoutput.t65 4.06363
R7483 CSoutput.n79 CSoutput.t123 4.06363
R7484 CSoutput.n80 CSoutput.t72 4.06363
R7485 CSoutput.n80 CSoutput.t98 4.06363
R7486 CSoutput.n82 CSoutput.t177 4.06363
R7487 CSoutput.n82 CSoutput.t116 4.06363
R7488 CSoutput.n84 CSoutput.t74 4.06363
R7489 CSoutput.n84 CSoutput.t156 4.06363
R7490 CSoutput.n86 CSoutput.t81 4.06363
R7491 CSoutput.n86 CSoutput.t138 4.06363
R7492 CSoutput.n88 CSoutput.t103 4.06363
R7493 CSoutput.n88 CSoutput.t124 4.06363
R7494 CSoutput.n90 CSoutput.t119 4.06363
R7495 CSoutput.n90 CSoutput.t165 4.06363
R7496 CSoutput.n92 CSoutput.t91 4.06363
R7497 CSoutput.n92 CSoutput.t143 4.06363
R7498 CSoutput.n94 CSoutput.t112 4.06363
R7499 CSoutput.n94 CSoutput.t158 4.06363
R7500 CSoutput.n96 CSoutput.t128 4.06363
R7501 CSoutput.n96 CSoutput.t173 4.06363
R7502 CSoutput.n44 CSoutput.n43 3.79402
R7503 CSoutput.n49 CSoutput.n48 3.79402
R7504 CSoutput.n383 CSoutput.n371 3.72967
R7505 CSoutput.n419 CSoutput.n407 3.72967
R7506 CSoutput.n421 CSoutput.n420 3.67605
R7507 CSoutput.n348 CSoutput.n138 2.99158
R7508 CSoutput.n381 CSoutput.t28 2.82907
R7509 CSoutput.n381 CSoutput.t27 2.82907
R7510 CSoutput.n379 CSoutput.t26 2.82907
R7511 CSoutput.n379 CSoutput.t41 2.82907
R7512 CSoutput.n377 CSoutput.t37 2.82907
R7513 CSoutput.n377 CSoutput.t3 2.82907
R7514 CSoutput.n375 CSoutput.t188 2.82907
R7515 CSoutput.n375 CSoutput.t7 2.82907
R7516 CSoutput.n373 CSoutput.t9 2.82907
R7517 CSoutput.n373 CSoutput.t44 2.82907
R7518 CSoutput.n372 CSoutput.t185 2.82907
R7519 CSoutput.n372 CSoutput.t0 2.82907
R7520 CSoutput.n369 CSoutput.t189 2.82907
R7521 CSoutput.n369 CSoutput.t2 2.82907
R7522 CSoutput.n367 CSoutput.t22 2.82907
R7523 CSoutput.n367 CSoutput.t56 2.82907
R7524 CSoutput.n365 CSoutput.t183 2.82907
R7525 CSoutput.n365 CSoutput.t5 2.82907
R7526 CSoutput.n363 CSoutput.t187 2.82907
R7527 CSoutput.n363 CSoutput.t23 2.82907
R7528 CSoutput.n361 CSoutput.t14 2.82907
R7529 CSoutput.n361 CSoutput.t29 2.82907
R7530 CSoutput.n360 CSoutput.t6 2.82907
R7531 CSoutput.n360 CSoutput.t47 2.82907
R7532 CSoutput.n358 CSoutput.t57 2.82907
R7533 CSoutput.n358 CSoutput.t12 2.82907
R7534 CSoutput.n356 CSoutput.t35 2.82907
R7535 CSoutput.n356 CSoutput.t36 2.82907
R7536 CSoutput.n354 CSoutput.t1 2.82907
R7537 CSoutput.n354 CSoutput.t52 2.82907
R7538 CSoutput.n352 CSoutput.t25 2.82907
R7539 CSoutput.n352 CSoutput.t34 2.82907
R7540 CSoutput.n350 CSoutput.t53 2.82907
R7541 CSoutput.n350 CSoutput.t39 2.82907
R7542 CSoutput.n349 CSoutput.t38 2.82907
R7543 CSoutput.n349 CSoutput.t10 2.82907
R7544 CSoutput.n408 CSoutput.t58 2.82907
R7545 CSoutput.n408 CSoutput.t31 2.82907
R7546 CSoutput.n409 CSoutput.t24 2.82907
R7547 CSoutput.n409 CSoutput.t40 2.82907
R7548 CSoutput.n411 CSoutput.t33 2.82907
R7549 CSoutput.n411 CSoutput.t13 2.82907
R7550 CSoutput.n413 CSoutput.t42 2.82907
R7551 CSoutput.n413 CSoutput.t55 2.82907
R7552 CSoutput.n415 CSoutput.t16 2.82907
R7553 CSoutput.n415 CSoutput.t18 2.82907
R7554 CSoutput.n417 CSoutput.t46 2.82907
R7555 CSoutput.n417 CSoutput.t45 2.82907
R7556 CSoutput.n396 CSoutput.t20 2.82907
R7557 CSoutput.n396 CSoutput.t186 2.82907
R7558 CSoutput.n397 CSoutput.t30 2.82907
R7559 CSoutput.n397 CSoutput.t50 2.82907
R7560 CSoutput.n399 CSoutput.t51 2.82907
R7561 CSoutput.n399 CSoutput.t17 2.82907
R7562 CSoutput.n401 CSoutput.t180 2.82907
R7563 CSoutput.n401 CSoutput.t19 2.82907
R7564 CSoutput.n403 CSoutput.t190 2.82907
R7565 CSoutput.n403 CSoutput.t21 2.82907
R7566 CSoutput.n405 CSoutput.t182 2.82907
R7567 CSoutput.n405 CSoutput.t15 2.82907
R7568 CSoutput.n385 CSoutput.t49 2.82907
R7569 CSoutput.n385 CSoutput.t181 2.82907
R7570 CSoutput.n386 CSoutput.t191 2.82907
R7571 CSoutput.n386 CSoutput.t32 2.82907
R7572 CSoutput.n388 CSoutput.t8 2.82907
R7573 CSoutput.n388 CSoutput.t43 2.82907
R7574 CSoutput.n390 CSoutput.t54 2.82907
R7575 CSoutput.n390 CSoutput.t184 2.82907
R7576 CSoutput.n392 CSoutput.t179 2.82907
R7577 CSoutput.n392 CSoutput.t48 2.82907
R7578 CSoutput.n394 CSoutput.t4 2.82907
R7579 CSoutput.n394 CSoutput.t11 2.82907
R7580 CSoutput.n420 CSoutput.n384 2.75627
R7581 CSoutput.n75 CSoutput.n1 2.45513
R7582 CSoutput.n229 CSoutput.n227 2.251
R7583 CSoutput.n229 CSoutput.n226 2.251
R7584 CSoutput.n229 CSoutput.n225 2.251
R7585 CSoutput.n229 CSoutput.n224 2.251
R7586 CSoutput.n198 CSoutput.n197 2.251
R7587 CSoutput.n198 CSoutput.n196 2.251
R7588 CSoutput.n198 CSoutput.n195 2.251
R7589 CSoutput.n198 CSoutput.n194 2.251
R7590 CSoutput.n271 CSoutput.n270 2.251
R7591 CSoutput.n236 CSoutput.n234 2.251
R7592 CSoutput.n236 CSoutput.n233 2.251
R7593 CSoutput.n236 CSoutput.n232 2.251
R7594 CSoutput.n254 CSoutput.n236 2.251
R7595 CSoutput.n242 CSoutput.n241 2.251
R7596 CSoutput.n242 CSoutput.n240 2.251
R7597 CSoutput.n242 CSoutput.n239 2.251
R7598 CSoutput.n242 CSoutput.n238 2.251
R7599 CSoutput.n268 CSoutput.n208 2.251
R7600 CSoutput.n263 CSoutput.n261 2.251
R7601 CSoutput.n263 CSoutput.n260 2.251
R7602 CSoutput.n263 CSoutput.n259 2.251
R7603 CSoutput.n263 CSoutput.n258 2.251
R7604 CSoutput.n164 CSoutput.n163 2.251
R7605 CSoutput.n164 CSoutput.n162 2.251
R7606 CSoutput.n164 CSoutput.n161 2.251
R7607 CSoutput.n164 CSoutput.n160 2.251
R7608 CSoutput.n281 CSoutput.n280 2.251
R7609 CSoutput.n198 CSoutput.n178 2.2505
R7610 CSoutput.n193 CSoutput.n178 2.2505
R7611 CSoutput.n191 CSoutput.n178 2.2505
R7612 CSoutput.n190 CSoutput.n178 2.2505
R7613 CSoutput.n275 CSoutput.n178 2.2505
R7614 CSoutput.n273 CSoutput.n178 2.2505
R7615 CSoutput.n271 CSoutput.n178 2.2505
R7616 CSoutput.n201 CSoutput.n178 2.2505
R7617 CSoutput.n200 CSoutput.n178 2.2505
R7618 CSoutput.n204 CSoutput.n178 2.2505
R7619 CSoutput.n203 CSoutput.n178 2.2505
R7620 CSoutput.n186 CSoutput.n178 2.2505
R7621 CSoutput.n278 CSoutput.n178 2.2505
R7622 CSoutput.n278 CSoutput.n277 2.2505
R7623 CSoutput.n242 CSoutput.n213 2.2505
R7624 CSoutput.n223 CSoutput.n213 2.2505
R7625 CSoutput.n244 CSoutput.n213 2.2505
R7626 CSoutput.n222 CSoutput.n213 2.2505
R7627 CSoutput.n246 CSoutput.n213 2.2505
R7628 CSoutput.n213 CSoutput.n207 2.2505
R7629 CSoutput.n268 CSoutput.n213 2.2505
R7630 CSoutput.n266 CSoutput.n213 2.2505
R7631 CSoutput.n248 CSoutput.n213 2.2505
R7632 CSoutput.n220 CSoutput.n213 2.2505
R7633 CSoutput.n250 CSoutput.n213 2.2505
R7634 CSoutput.n219 CSoutput.n213 2.2505
R7635 CSoutput.n264 CSoutput.n213 2.2505
R7636 CSoutput.n264 CSoutput.n217 2.2505
R7637 CSoutput.n164 CSoutput.n144 2.2505
R7638 CSoutput.n159 CSoutput.n144 2.2505
R7639 CSoutput.n157 CSoutput.n144 2.2505
R7640 CSoutput.n156 CSoutput.n144 2.2505
R7641 CSoutput.n285 CSoutput.n144 2.2505
R7642 CSoutput.n283 CSoutput.n144 2.2505
R7643 CSoutput.n281 CSoutput.n144 2.2505
R7644 CSoutput.n167 CSoutput.n144 2.2505
R7645 CSoutput.n166 CSoutput.n144 2.2505
R7646 CSoutput.n170 CSoutput.n144 2.2505
R7647 CSoutput.n169 CSoutput.n144 2.2505
R7648 CSoutput.n152 CSoutput.n144 2.2505
R7649 CSoutput.n288 CSoutput.n144 2.2505
R7650 CSoutput.n288 CSoutput.n287 2.2505
R7651 CSoutput.n206 CSoutput.n199 2.25024
R7652 CSoutput.n206 CSoutput.n192 2.25024
R7653 CSoutput.n274 CSoutput.n206 2.25024
R7654 CSoutput.n206 CSoutput.n202 2.25024
R7655 CSoutput.n206 CSoutput.n205 2.25024
R7656 CSoutput.n206 CSoutput.n173 2.25024
R7657 CSoutput.n256 CSoutput.n253 2.25024
R7658 CSoutput.n256 CSoutput.n252 2.25024
R7659 CSoutput.n256 CSoutput.n251 2.25024
R7660 CSoutput.n256 CSoutput.n218 2.25024
R7661 CSoutput.n256 CSoutput.n255 2.25024
R7662 CSoutput.n257 CSoutput.n256 2.25024
R7663 CSoutput.n172 CSoutput.n165 2.25024
R7664 CSoutput.n172 CSoutput.n158 2.25024
R7665 CSoutput.n284 CSoutput.n172 2.25024
R7666 CSoutput.n172 CSoutput.n168 2.25024
R7667 CSoutput.n172 CSoutput.n171 2.25024
R7668 CSoutput.n172 CSoutput.n139 2.25024
R7669 CSoutput.n273 CSoutput.n183 1.50111
R7670 CSoutput.n221 CSoutput.n207 1.50111
R7671 CSoutput.n283 CSoutput.n149 1.50111
R7672 CSoutput.n229 CSoutput.n228 1.501
R7673 CSoutput.n236 CSoutput.n235 1.501
R7674 CSoutput.n263 CSoutput.n262 1.501
R7675 CSoutput.n277 CSoutput.n188 1.12536
R7676 CSoutput.n277 CSoutput.n189 1.12536
R7677 CSoutput.n277 CSoutput.n276 1.12536
R7678 CSoutput.n237 CSoutput.n217 1.12536
R7679 CSoutput.n243 CSoutput.n217 1.12536
R7680 CSoutput.n245 CSoutput.n217 1.12536
R7681 CSoutput.n287 CSoutput.n154 1.12536
R7682 CSoutput.n287 CSoutput.n155 1.12536
R7683 CSoutput.n287 CSoutput.n286 1.12536
R7684 CSoutput.n277 CSoutput.n184 1.12536
R7685 CSoutput.n277 CSoutput.n185 1.12536
R7686 CSoutput.n277 CSoutput.n187 1.12536
R7687 CSoutput.n267 CSoutput.n217 1.12536
R7688 CSoutput.n247 CSoutput.n217 1.12536
R7689 CSoutput.n249 CSoutput.n217 1.12536
R7690 CSoutput.n287 CSoutput.n150 1.12536
R7691 CSoutput.n287 CSoutput.n151 1.12536
R7692 CSoutput.n287 CSoutput.n153 1.12536
R7693 CSoutput.n31 CSoutput.n30 0.669944
R7694 CSoutput.n62 CSoutput.n61 0.669944
R7695 CSoutput.n376 CSoutput.n374 0.573776
R7696 CSoutput.n378 CSoutput.n376 0.573776
R7697 CSoutput.n380 CSoutput.n378 0.573776
R7698 CSoutput.n382 CSoutput.n380 0.573776
R7699 CSoutput.n364 CSoutput.n362 0.573776
R7700 CSoutput.n366 CSoutput.n364 0.573776
R7701 CSoutput.n368 CSoutput.n366 0.573776
R7702 CSoutput.n370 CSoutput.n368 0.573776
R7703 CSoutput.n353 CSoutput.n351 0.573776
R7704 CSoutput.n355 CSoutput.n353 0.573776
R7705 CSoutput.n357 CSoutput.n355 0.573776
R7706 CSoutput.n359 CSoutput.n357 0.573776
R7707 CSoutput.n418 CSoutput.n416 0.573776
R7708 CSoutput.n416 CSoutput.n414 0.573776
R7709 CSoutput.n414 CSoutput.n412 0.573776
R7710 CSoutput.n412 CSoutput.n410 0.573776
R7711 CSoutput.n406 CSoutput.n404 0.573776
R7712 CSoutput.n404 CSoutput.n402 0.573776
R7713 CSoutput.n402 CSoutput.n400 0.573776
R7714 CSoutput.n400 CSoutput.n398 0.573776
R7715 CSoutput.n395 CSoutput.n393 0.573776
R7716 CSoutput.n393 CSoutput.n391 0.573776
R7717 CSoutput.n391 CSoutput.n389 0.573776
R7718 CSoutput.n389 CSoutput.n387 0.573776
R7719 CSoutput.n421 CSoutput.n288 0.534538
R7720 CSoutput.n332 CSoutput.n330 0.358259
R7721 CSoutput.n334 CSoutput.n332 0.358259
R7722 CSoutput.n336 CSoutput.n334 0.358259
R7723 CSoutput.n338 CSoutput.n336 0.358259
R7724 CSoutput.n340 CSoutput.n338 0.358259
R7725 CSoutput.n342 CSoutput.n340 0.358259
R7726 CSoutput.n344 CSoutput.n342 0.358259
R7727 CSoutput.n346 CSoutput.n344 0.358259
R7728 CSoutput.n312 CSoutput.n310 0.358259
R7729 CSoutput.n314 CSoutput.n312 0.358259
R7730 CSoutput.n316 CSoutput.n314 0.358259
R7731 CSoutput.n318 CSoutput.n316 0.358259
R7732 CSoutput.n320 CSoutput.n318 0.358259
R7733 CSoutput.n322 CSoutput.n320 0.358259
R7734 CSoutput.n324 CSoutput.n322 0.358259
R7735 CSoutput.n326 CSoutput.n324 0.358259
R7736 CSoutput.n293 CSoutput.n291 0.358259
R7737 CSoutput.n295 CSoutput.n293 0.358259
R7738 CSoutput.n297 CSoutput.n295 0.358259
R7739 CSoutput.n299 CSoutput.n297 0.358259
R7740 CSoutput.n301 CSoutput.n299 0.358259
R7741 CSoutput.n303 CSoutput.n301 0.358259
R7742 CSoutput.n305 CSoutput.n303 0.358259
R7743 CSoutput.n307 CSoutput.n305 0.358259
R7744 CSoutput.n136 CSoutput.n134 0.358259
R7745 CSoutput.n134 CSoutput.n132 0.358259
R7746 CSoutput.n132 CSoutput.n130 0.358259
R7747 CSoutput.n130 CSoutput.n128 0.358259
R7748 CSoutput.n128 CSoutput.n126 0.358259
R7749 CSoutput.n126 CSoutput.n124 0.358259
R7750 CSoutput.n124 CSoutput.n122 0.358259
R7751 CSoutput.n122 CSoutput.n120 0.358259
R7752 CSoutput.n116 CSoutput.n114 0.358259
R7753 CSoutput.n114 CSoutput.n112 0.358259
R7754 CSoutput.n112 CSoutput.n110 0.358259
R7755 CSoutput.n110 CSoutput.n108 0.358259
R7756 CSoutput.n108 CSoutput.n106 0.358259
R7757 CSoutput.n106 CSoutput.n104 0.358259
R7758 CSoutput.n104 CSoutput.n102 0.358259
R7759 CSoutput.n102 CSoutput.n100 0.358259
R7760 CSoutput.n97 CSoutput.n95 0.358259
R7761 CSoutput.n95 CSoutput.n93 0.358259
R7762 CSoutput.n93 CSoutput.n91 0.358259
R7763 CSoutput.n91 CSoutput.n89 0.358259
R7764 CSoutput.n89 CSoutput.n87 0.358259
R7765 CSoutput.n87 CSoutput.n85 0.358259
R7766 CSoutput.n85 CSoutput.n83 0.358259
R7767 CSoutput.n83 CSoutput.n81 0.358259
R7768 CSoutput.n21 CSoutput.n20 0.169105
R7769 CSoutput.n21 CSoutput.n16 0.169105
R7770 CSoutput.n26 CSoutput.n16 0.169105
R7771 CSoutput.n27 CSoutput.n26 0.169105
R7772 CSoutput.n27 CSoutput.n14 0.169105
R7773 CSoutput.n32 CSoutput.n14 0.169105
R7774 CSoutput.n33 CSoutput.n32 0.169105
R7775 CSoutput.n34 CSoutput.n33 0.169105
R7776 CSoutput.n34 CSoutput.n12 0.169105
R7777 CSoutput.n39 CSoutput.n12 0.169105
R7778 CSoutput.n40 CSoutput.n39 0.169105
R7779 CSoutput.n40 CSoutput.n10 0.169105
R7780 CSoutput.n45 CSoutput.n10 0.169105
R7781 CSoutput.n46 CSoutput.n45 0.169105
R7782 CSoutput.n47 CSoutput.n46 0.169105
R7783 CSoutput.n47 CSoutput.n8 0.169105
R7784 CSoutput.n52 CSoutput.n8 0.169105
R7785 CSoutput.n53 CSoutput.n52 0.169105
R7786 CSoutput.n53 CSoutput.n6 0.169105
R7787 CSoutput.n58 CSoutput.n6 0.169105
R7788 CSoutput.n59 CSoutput.n58 0.169105
R7789 CSoutput.n60 CSoutput.n59 0.169105
R7790 CSoutput.n60 CSoutput.n4 0.169105
R7791 CSoutput.n66 CSoutput.n4 0.169105
R7792 CSoutput.n67 CSoutput.n66 0.169105
R7793 CSoutput.n68 CSoutput.n67 0.169105
R7794 CSoutput.n68 CSoutput.n2 0.169105
R7795 CSoutput.n73 CSoutput.n2 0.169105
R7796 CSoutput.n74 CSoutput.n73 0.169105
R7797 CSoutput.n74 CSoutput.n0 0.169105
R7798 CSoutput.n78 CSoutput.n0 0.169105
R7799 CSoutput.n231 CSoutput.n230 0.0910737
R7800 CSoutput.n282 CSoutput.n279 0.0723685
R7801 CSoutput.n236 CSoutput.n231 0.0522944
R7802 CSoutput.n279 CSoutput.n278 0.0499135
R7803 CSoutput.n230 CSoutput.n229 0.0499135
R7804 CSoutput.n264 CSoutput.n263 0.0464294
R7805 CSoutput.n272 CSoutput.n269 0.0391444
R7806 CSoutput.n231 CSoutput.t207 0.023435
R7807 CSoutput.n279 CSoutput.t194 0.02262
R7808 CSoutput.n230 CSoutput.t213 0.02262
R7809 CSoutput CSoutput.n421 0.0052
R7810 CSoutput.n201 CSoutput.n184 0.00365111
R7811 CSoutput.n204 CSoutput.n185 0.00365111
R7812 CSoutput.n187 CSoutput.n186 0.00365111
R7813 CSoutput.n229 CSoutput.n188 0.00365111
R7814 CSoutput.n193 CSoutput.n189 0.00365111
R7815 CSoutput.n276 CSoutput.n190 0.00365111
R7816 CSoutput.n267 CSoutput.n266 0.00365111
R7817 CSoutput.n247 CSoutput.n220 0.00365111
R7818 CSoutput.n249 CSoutput.n219 0.00365111
R7819 CSoutput.n237 CSoutput.n236 0.00365111
R7820 CSoutput.n243 CSoutput.n223 0.00365111
R7821 CSoutput.n245 CSoutput.n222 0.00365111
R7822 CSoutput.n167 CSoutput.n150 0.00365111
R7823 CSoutput.n170 CSoutput.n151 0.00365111
R7824 CSoutput.n153 CSoutput.n152 0.00365111
R7825 CSoutput.n263 CSoutput.n154 0.00365111
R7826 CSoutput.n159 CSoutput.n155 0.00365111
R7827 CSoutput.n286 CSoutput.n156 0.00365111
R7828 CSoutput.n198 CSoutput.n188 0.00340054
R7829 CSoutput.n191 CSoutput.n189 0.00340054
R7830 CSoutput.n276 CSoutput.n275 0.00340054
R7831 CSoutput.n271 CSoutput.n184 0.00340054
R7832 CSoutput.n200 CSoutput.n185 0.00340054
R7833 CSoutput.n203 CSoutput.n187 0.00340054
R7834 CSoutput.n242 CSoutput.n237 0.00340054
R7835 CSoutput.n244 CSoutput.n243 0.00340054
R7836 CSoutput.n246 CSoutput.n245 0.00340054
R7837 CSoutput.n268 CSoutput.n267 0.00340054
R7838 CSoutput.n248 CSoutput.n247 0.00340054
R7839 CSoutput.n250 CSoutput.n249 0.00340054
R7840 CSoutput.n164 CSoutput.n154 0.00340054
R7841 CSoutput.n157 CSoutput.n155 0.00340054
R7842 CSoutput.n286 CSoutput.n285 0.00340054
R7843 CSoutput.n281 CSoutput.n150 0.00340054
R7844 CSoutput.n166 CSoutput.n151 0.00340054
R7845 CSoutput.n169 CSoutput.n153 0.00340054
R7846 CSoutput.n199 CSoutput.n193 0.00252698
R7847 CSoutput.n192 CSoutput.n190 0.00252698
R7848 CSoutput.n274 CSoutput.n273 0.00252698
R7849 CSoutput.n202 CSoutput.n200 0.00252698
R7850 CSoutput.n205 CSoutput.n203 0.00252698
R7851 CSoutput.n278 CSoutput.n173 0.00252698
R7852 CSoutput.n199 CSoutput.n198 0.00252698
R7853 CSoutput.n192 CSoutput.n191 0.00252698
R7854 CSoutput.n275 CSoutput.n274 0.00252698
R7855 CSoutput.n202 CSoutput.n201 0.00252698
R7856 CSoutput.n205 CSoutput.n204 0.00252698
R7857 CSoutput.n186 CSoutput.n173 0.00252698
R7858 CSoutput.n253 CSoutput.n223 0.00252698
R7859 CSoutput.n252 CSoutput.n222 0.00252698
R7860 CSoutput.n251 CSoutput.n207 0.00252698
R7861 CSoutput.n248 CSoutput.n218 0.00252698
R7862 CSoutput.n255 CSoutput.n250 0.00252698
R7863 CSoutput.n264 CSoutput.n257 0.00252698
R7864 CSoutput.n253 CSoutput.n242 0.00252698
R7865 CSoutput.n252 CSoutput.n244 0.00252698
R7866 CSoutput.n251 CSoutput.n246 0.00252698
R7867 CSoutput.n266 CSoutput.n218 0.00252698
R7868 CSoutput.n255 CSoutput.n220 0.00252698
R7869 CSoutput.n257 CSoutput.n219 0.00252698
R7870 CSoutput.n165 CSoutput.n159 0.00252698
R7871 CSoutput.n158 CSoutput.n156 0.00252698
R7872 CSoutput.n284 CSoutput.n283 0.00252698
R7873 CSoutput.n168 CSoutput.n166 0.00252698
R7874 CSoutput.n171 CSoutput.n169 0.00252698
R7875 CSoutput.n288 CSoutput.n139 0.00252698
R7876 CSoutput.n165 CSoutput.n164 0.00252698
R7877 CSoutput.n158 CSoutput.n157 0.00252698
R7878 CSoutput.n285 CSoutput.n284 0.00252698
R7879 CSoutput.n168 CSoutput.n167 0.00252698
R7880 CSoutput.n171 CSoutput.n170 0.00252698
R7881 CSoutput.n152 CSoutput.n139 0.00252698
R7882 CSoutput.n273 CSoutput.n272 0.0020275
R7883 CSoutput.n272 CSoutput.n271 0.0020275
R7884 CSoutput.n269 CSoutput.n207 0.0020275
R7885 CSoutput.n269 CSoutput.n268 0.0020275
R7886 CSoutput.n283 CSoutput.n282 0.0020275
R7887 CSoutput.n282 CSoutput.n281 0.0020275
R7888 CSoutput.n183 CSoutput.n182 0.00166668
R7889 CSoutput.n265 CSoutput.n221 0.00166668
R7890 CSoutput.n149 CSoutput.n148 0.00166668
R7891 CSoutput.n287 CSoutput.n149 0.00133328
R7892 CSoutput.n221 CSoutput.n217 0.00133328
R7893 CSoutput.n277 CSoutput.n183 0.00133328
R7894 CSoutput.n280 CSoutput.n172 0.001
R7895 CSoutput.n258 CSoutput.n172 0.001
R7896 CSoutput.n160 CSoutput.n140 0.001
R7897 CSoutput.n259 CSoutput.n140 0.001
R7898 CSoutput.n161 CSoutput.n141 0.001
R7899 CSoutput.n260 CSoutput.n141 0.001
R7900 CSoutput.n162 CSoutput.n142 0.001
R7901 CSoutput.n261 CSoutput.n142 0.001
R7902 CSoutput.n163 CSoutput.n143 0.001
R7903 CSoutput.n262 CSoutput.n143 0.001
R7904 CSoutput.n256 CSoutput.n208 0.001
R7905 CSoutput.n256 CSoutput.n254 0.001
R7906 CSoutput.n238 CSoutput.n209 0.001
R7907 CSoutput.n232 CSoutput.n209 0.001
R7908 CSoutput.n239 CSoutput.n210 0.001
R7909 CSoutput.n233 CSoutput.n210 0.001
R7910 CSoutput.n240 CSoutput.n211 0.001
R7911 CSoutput.n234 CSoutput.n211 0.001
R7912 CSoutput.n241 CSoutput.n212 0.001
R7913 CSoutput.n235 CSoutput.n212 0.001
R7914 CSoutput.n270 CSoutput.n206 0.001
R7915 CSoutput.n224 CSoutput.n206 0.001
R7916 CSoutput.n194 CSoutput.n174 0.001
R7917 CSoutput.n225 CSoutput.n174 0.001
R7918 CSoutput.n195 CSoutput.n175 0.001
R7919 CSoutput.n226 CSoutput.n175 0.001
R7920 CSoutput.n196 CSoutput.n176 0.001
R7921 CSoutput.n227 CSoutput.n176 0.001
R7922 CSoutput.n197 CSoutput.n177 0.001
R7923 CSoutput.n228 CSoutput.n177 0.001
R7924 CSoutput.n228 CSoutput.n178 0.001
R7925 CSoutput.n227 CSoutput.n179 0.001
R7926 CSoutput.n226 CSoutput.n180 0.001
R7927 CSoutput.n225 CSoutput.t206 0.001
R7928 CSoutput.n224 CSoutput.n181 0.001
R7929 CSoutput.n197 CSoutput.n179 0.001
R7930 CSoutput.n196 CSoutput.n180 0.001
R7931 CSoutput.n195 CSoutput.t206 0.001
R7932 CSoutput.n194 CSoutput.n181 0.001
R7933 CSoutput.n270 CSoutput.n182 0.001
R7934 CSoutput.n235 CSoutput.n213 0.001
R7935 CSoutput.n234 CSoutput.n214 0.001
R7936 CSoutput.n233 CSoutput.n215 0.001
R7937 CSoutput.n232 CSoutput.t196 0.001
R7938 CSoutput.n254 CSoutput.n216 0.001
R7939 CSoutput.n241 CSoutput.n214 0.001
R7940 CSoutput.n240 CSoutput.n215 0.001
R7941 CSoutput.n239 CSoutput.t196 0.001
R7942 CSoutput.n238 CSoutput.n216 0.001
R7943 CSoutput.n265 CSoutput.n208 0.001
R7944 CSoutput.n262 CSoutput.n144 0.001
R7945 CSoutput.n261 CSoutput.n145 0.001
R7946 CSoutput.n260 CSoutput.n146 0.001
R7947 CSoutput.n259 CSoutput.t199 0.001
R7948 CSoutput.n258 CSoutput.n147 0.001
R7949 CSoutput.n163 CSoutput.n145 0.001
R7950 CSoutput.n162 CSoutput.n146 0.001
R7951 CSoutput.n161 CSoutput.t199 0.001
R7952 CSoutput.n160 CSoutput.n147 0.001
R7953 CSoutput.n280 CSoutput.n148 0.001
R7954 commonsourceibias.n25 commonsourceibias.t30 230.006
R7955 commonsourceibias.n91 commonsourceibias.t73 230.006
R7956 commonsourceibias.n218 commonsourceibias.t98 230.006
R7957 commonsourceibias.n154 commonsourceibias.t70 230.006
R7958 commonsourceibias.n322 commonsourceibias.t4 230.006
R7959 commonsourceibias.n281 commonsourceibias.t111 230.006
R7960 commonsourceibias.n483 commonsourceibias.t113 230.006
R7961 commonsourceibias.n419 commonsourceibias.t52 230.006
R7962 commonsourceibias.n70 commonsourceibias.t6 207.983
R7963 commonsourceibias.n136 commonsourceibias.t89 207.983
R7964 commonsourceibias.n263 commonsourceibias.t109 207.983
R7965 commonsourceibias.n199 commonsourceibias.t54 207.983
R7966 commonsourceibias.n368 commonsourceibias.t34 207.983
R7967 commonsourceibias.n402 commonsourceibias.t69 207.983
R7968 commonsourceibias.n529 commonsourceibias.t63 207.983
R7969 commonsourceibias.n465 commonsourceibias.t112 207.983
R7970 commonsourceibias.n10 commonsourceibias.t24 168.701
R7971 commonsourceibias.n63 commonsourceibias.t20 168.701
R7972 commonsourceibias.n57 commonsourceibias.t42 168.701
R7973 commonsourceibias.n16 commonsourceibias.t10 168.701
R7974 commonsourceibias.n49 commonsourceibias.t40 168.701
R7975 commonsourceibias.n43 commonsourceibias.t28 168.701
R7976 commonsourceibias.n19 commonsourceibias.t46 168.701
R7977 commonsourceibias.n21 commonsourceibias.t16 168.701
R7978 commonsourceibias.n23 commonsourceibias.t26 168.701
R7979 commonsourceibias.n26 commonsourceibias.t0 168.701
R7980 commonsourceibias.n1 commonsourceibias.t51 168.701
R7981 commonsourceibias.n129 commonsourceibias.t95 168.701
R7982 commonsourceibias.n123 commonsourceibias.t90 168.701
R7983 commonsourceibias.n7 commonsourceibias.t101 168.701
R7984 commonsourceibias.n115 commonsourceibias.t86 168.701
R7985 commonsourceibias.n109 commonsourceibias.t77 168.701
R7986 commonsourceibias.n85 commonsourceibias.t94 168.701
R7987 commonsourceibias.n87 commonsourceibias.t87 168.701
R7988 commonsourceibias.n89 commonsourceibias.t58 168.701
R7989 commonsourceibias.n92 commonsourceibias.t80 168.701
R7990 commonsourceibias.n219 commonsourceibias.t102 168.701
R7991 commonsourceibias.n216 commonsourceibias.t48 168.701
R7992 commonsourceibias.n214 commonsourceibias.t103 168.701
R7993 commonsourceibias.n212 commonsourceibias.t108 168.701
R7994 commonsourceibias.n236 commonsourceibias.t88 168.701
R7995 commonsourceibias.n242 commonsourceibias.t68 168.701
R7996 commonsourceibias.n209 commonsourceibias.t115 168.701
R7997 commonsourceibias.n250 commonsourceibias.t93 168.701
R7998 commonsourceibias.n256 commonsourceibias.t96 168.701
R7999 commonsourceibias.n203 commonsourceibias.t57 168.701
R8000 commonsourceibias.n139 commonsourceibias.t119 168.701
R8001 commonsourceibias.n192 commonsourceibias.t110 168.701
R8002 commonsourceibias.n186 commonsourceibias.t60 168.701
R8003 commonsourceibias.n145 commonsourceibias.t117 168.701
R8004 commonsourceibias.n178 commonsourceibias.t65 168.701
R8005 commonsourceibias.n172 commonsourceibias.t59 168.701
R8006 commonsourceibias.n148 commonsourceibias.t118 168.701
R8007 commonsourceibias.n150 commonsourceibias.t71 168.701
R8008 commonsourceibias.n152 commonsourceibias.t83 168.701
R8009 commonsourceibias.n155 commonsourceibias.t116 168.701
R8010 commonsourceibias.n323 commonsourceibias.t38 168.701
R8011 commonsourceibias.n320 commonsourceibias.t12 168.701
R8012 commonsourceibias.n318 commonsourceibias.t36 168.701
R8013 commonsourceibias.n316 commonsourceibias.t2 168.701
R8014 commonsourceibias.n340 commonsourceibias.t44 168.701
R8015 commonsourceibias.n346 commonsourceibias.t22 168.701
R8016 commonsourceibias.n348 commonsourceibias.t18 168.701
R8017 commonsourceibias.n355 commonsourceibias.t32 168.701
R8018 commonsourceibias.n361 commonsourceibias.t14 168.701
R8019 commonsourceibias.n308 commonsourceibias.t8 168.701
R8020 commonsourceibias.n267 commonsourceibias.t99 168.701
R8021 commonsourceibias.n395 commonsourceibias.t84 168.701
R8022 commonsourceibias.n389 commonsourceibias.t72 168.701
R8023 commonsourceibias.n382 commonsourceibias.t92 168.701
R8024 commonsourceibias.n380 commonsourceibias.t66 168.701
R8025 commonsourceibias.n282 commonsourceibias.t64 168.701
R8026 commonsourceibias.n279 commonsourceibias.t104 168.701
R8027 commonsourceibias.n277 commonsourceibias.t67 168.701
R8028 commonsourceibias.n275 commonsourceibias.t79 168.701
R8029 commonsourceibias.n299 commonsourceibias.t56 168.701
R8030 commonsourceibias.n484 commonsourceibias.t97 168.701
R8031 commonsourceibias.n481 commonsourceibias.t78 168.701
R8032 commonsourceibias.n479 commonsourceibias.t53 168.701
R8033 commonsourceibias.n477 commonsourceibias.t62 168.701
R8034 commonsourceibias.n501 commonsourceibias.t82 168.701
R8035 commonsourceibias.n507 commonsourceibias.t85 168.701
R8036 commonsourceibias.n509 commonsourceibias.t76 168.701
R8037 commonsourceibias.n516 commonsourceibias.t100 168.701
R8038 commonsourceibias.n522 commonsourceibias.t91 168.701
R8039 commonsourceibias.n469 commonsourceibias.t81 168.701
R8040 commonsourceibias.n420 commonsourceibias.t61 168.701
R8041 commonsourceibias.n417 commonsourceibias.t75 168.701
R8042 commonsourceibias.n415 commonsourceibias.t55 168.701
R8043 commonsourceibias.n413 commonsourceibias.t105 168.701
R8044 commonsourceibias.n437 commonsourceibias.t74 168.701
R8045 commonsourceibias.n443 commonsourceibias.t49 168.701
R8046 commonsourceibias.n445 commonsourceibias.t106 168.701
R8047 commonsourceibias.n452 commonsourceibias.t114 168.701
R8048 commonsourceibias.n458 commonsourceibias.t50 168.701
R8049 commonsourceibias.n405 commonsourceibias.t107 168.701
R8050 commonsourceibias.n27 commonsourceibias.n24 161.3
R8051 commonsourceibias.n29 commonsourceibias.n28 161.3
R8052 commonsourceibias.n31 commonsourceibias.n30 161.3
R8053 commonsourceibias.n32 commonsourceibias.n22 161.3
R8054 commonsourceibias.n34 commonsourceibias.n33 161.3
R8055 commonsourceibias.n36 commonsourceibias.n35 161.3
R8056 commonsourceibias.n37 commonsourceibias.n20 161.3
R8057 commonsourceibias.n39 commonsourceibias.n38 161.3
R8058 commonsourceibias.n41 commonsourceibias.n40 161.3
R8059 commonsourceibias.n42 commonsourceibias.n18 161.3
R8060 commonsourceibias.n45 commonsourceibias.n44 161.3
R8061 commonsourceibias.n46 commonsourceibias.n17 161.3
R8062 commonsourceibias.n48 commonsourceibias.n47 161.3
R8063 commonsourceibias.n50 commonsourceibias.n15 161.3
R8064 commonsourceibias.n52 commonsourceibias.n51 161.3
R8065 commonsourceibias.n53 commonsourceibias.n14 161.3
R8066 commonsourceibias.n55 commonsourceibias.n54 161.3
R8067 commonsourceibias.n56 commonsourceibias.n13 161.3
R8068 commonsourceibias.n59 commonsourceibias.n58 161.3
R8069 commonsourceibias.n60 commonsourceibias.n12 161.3
R8070 commonsourceibias.n62 commonsourceibias.n61 161.3
R8071 commonsourceibias.n64 commonsourceibias.n11 161.3
R8072 commonsourceibias.n66 commonsourceibias.n65 161.3
R8073 commonsourceibias.n68 commonsourceibias.n67 161.3
R8074 commonsourceibias.n69 commonsourceibias.n9 161.3
R8075 commonsourceibias.n93 commonsourceibias.n90 161.3
R8076 commonsourceibias.n95 commonsourceibias.n94 161.3
R8077 commonsourceibias.n97 commonsourceibias.n96 161.3
R8078 commonsourceibias.n98 commonsourceibias.n88 161.3
R8079 commonsourceibias.n100 commonsourceibias.n99 161.3
R8080 commonsourceibias.n102 commonsourceibias.n101 161.3
R8081 commonsourceibias.n103 commonsourceibias.n86 161.3
R8082 commonsourceibias.n105 commonsourceibias.n104 161.3
R8083 commonsourceibias.n107 commonsourceibias.n106 161.3
R8084 commonsourceibias.n108 commonsourceibias.n84 161.3
R8085 commonsourceibias.n111 commonsourceibias.n110 161.3
R8086 commonsourceibias.n112 commonsourceibias.n8 161.3
R8087 commonsourceibias.n114 commonsourceibias.n113 161.3
R8088 commonsourceibias.n116 commonsourceibias.n6 161.3
R8089 commonsourceibias.n118 commonsourceibias.n117 161.3
R8090 commonsourceibias.n119 commonsourceibias.n5 161.3
R8091 commonsourceibias.n121 commonsourceibias.n120 161.3
R8092 commonsourceibias.n122 commonsourceibias.n4 161.3
R8093 commonsourceibias.n125 commonsourceibias.n124 161.3
R8094 commonsourceibias.n126 commonsourceibias.n3 161.3
R8095 commonsourceibias.n128 commonsourceibias.n127 161.3
R8096 commonsourceibias.n130 commonsourceibias.n2 161.3
R8097 commonsourceibias.n132 commonsourceibias.n131 161.3
R8098 commonsourceibias.n134 commonsourceibias.n133 161.3
R8099 commonsourceibias.n135 commonsourceibias.n0 161.3
R8100 commonsourceibias.n262 commonsourceibias.n202 161.3
R8101 commonsourceibias.n261 commonsourceibias.n260 161.3
R8102 commonsourceibias.n259 commonsourceibias.n258 161.3
R8103 commonsourceibias.n257 commonsourceibias.n204 161.3
R8104 commonsourceibias.n255 commonsourceibias.n254 161.3
R8105 commonsourceibias.n253 commonsourceibias.n205 161.3
R8106 commonsourceibias.n252 commonsourceibias.n251 161.3
R8107 commonsourceibias.n249 commonsourceibias.n206 161.3
R8108 commonsourceibias.n248 commonsourceibias.n247 161.3
R8109 commonsourceibias.n246 commonsourceibias.n207 161.3
R8110 commonsourceibias.n245 commonsourceibias.n244 161.3
R8111 commonsourceibias.n243 commonsourceibias.n208 161.3
R8112 commonsourceibias.n241 commonsourceibias.n240 161.3
R8113 commonsourceibias.n239 commonsourceibias.n210 161.3
R8114 commonsourceibias.n238 commonsourceibias.n237 161.3
R8115 commonsourceibias.n235 commonsourceibias.n211 161.3
R8116 commonsourceibias.n234 commonsourceibias.n233 161.3
R8117 commonsourceibias.n232 commonsourceibias.n231 161.3
R8118 commonsourceibias.n230 commonsourceibias.n213 161.3
R8119 commonsourceibias.n229 commonsourceibias.n228 161.3
R8120 commonsourceibias.n227 commonsourceibias.n226 161.3
R8121 commonsourceibias.n225 commonsourceibias.n215 161.3
R8122 commonsourceibias.n224 commonsourceibias.n223 161.3
R8123 commonsourceibias.n222 commonsourceibias.n221 161.3
R8124 commonsourceibias.n220 commonsourceibias.n217 161.3
R8125 commonsourceibias.n156 commonsourceibias.n153 161.3
R8126 commonsourceibias.n158 commonsourceibias.n157 161.3
R8127 commonsourceibias.n160 commonsourceibias.n159 161.3
R8128 commonsourceibias.n161 commonsourceibias.n151 161.3
R8129 commonsourceibias.n163 commonsourceibias.n162 161.3
R8130 commonsourceibias.n165 commonsourceibias.n164 161.3
R8131 commonsourceibias.n166 commonsourceibias.n149 161.3
R8132 commonsourceibias.n168 commonsourceibias.n167 161.3
R8133 commonsourceibias.n170 commonsourceibias.n169 161.3
R8134 commonsourceibias.n171 commonsourceibias.n147 161.3
R8135 commonsourceibias.n174 commonsourceibias.n173 161.3
R8136 commonsourceibias.n175 commonsourceibias.n146 161.3
R8137 commonsourceibias.n177 commonsourceibias.n176 161.3
R8138 commonsourceibias.n179 commonsourceibias.n144 161.3
R8139 commonsourceibias.n181 commonsourceibias.n180 161.3
R8140 commonsourceibias.n182 commonsourceibias.n143 161.3
R8141 commonsourceibias.n184 commonsourceibias.n183 161.3
R8142 commonsourceibias.n185 commonsourceibias.n142 161.3
R8143 commonsourceibias.n188 commonsourceibias.n187 161.3
R8144 commonsourceibias.n189 commonsourceibias.n141 161.3
R8145 commonsourceibias.n191 commonsourceibias.n190 161.3
R8146 commonsourceibias.n193 commonsourceibias.n140 161.3
R8147 commonsourceibias.n195 commonsourceibias.n194 161.3
R8148 commonsourceibias.n197 commonsourceibias.n196 161.3
R8149 commonsourceibias.n198 commonsourceibias.n138 161.3
R8150 commonsourceibias.n367 commonsourceibias.n307 161.3
R8151 commonsourceibias.n366 commonsourceibias.n365 161.3
R8152 commonsourceibias.n364 commonsourceibias.n363 161.3
R8153 commonsourceibias.n362 commonsourceibias.n309 161.3
R8154 commonsourceibias.n360 commonsourceibias.n359 161.3
R8155 commonsourceibias.n358 commonsourceibias.n310 161.3
R8156 commonsourceibias.n357 commonsourceibias.n356 161.3
R8157 commonsourceibias.n354 commonsourceibias.n311 161.3
R8158 commonsourceibias.n353 commonsourceibias.n352 161.3
R8159 commonsourceibias.n351 commonsourceibias.n312 161.3
R8160 commonsourceibias.n350 commonsourceibias.n349 161.3
R8161 commonsourceibias.n347 commonsourceibias.n313 161.3
R8162 commonsourceibias.n345 commonsourceibias.n344 161.3
R8163 commonsourceibias.n343 commonsourceibias.n314 161.3
R8164 commonsourceibias.n342 commonsourceibias.n341 161.3
R8165 commonsourceibias.n339 commonsourceibias.n315 161.3
R8166 commonsourceibias.n338 commonsourceibias.n337 161.3
R8167 commonsourceibias.n336 commonsourceibias.n335 161.3
R8168 commonsourceibias.n334 commonsourceibias.n317 161.3
R8169 commonsourceibias.n333 commonsourceibias.n332 161.3
R8170 commonsourceibias.n331 commonsourceibias.n330 161.3
R8171 commonsourceibias.n329 commonsourceibias.n319 161.3
R8172 commonsourceibias.n328 commonsourceibias.n327 161.3
R8173 commonsourceibias.n326 commonsourceibias.n325 161.3
R8174 commonsourceibias.n324 commonsourceibias.n321 161.3
R8175 commonsourceibias.n301 commonsourceibias.n300 161.3
R8176 commonsourceibias.n298 commonsourceibias.n274 161.3
R8177 commonsourceibias.n297 commonsourceibias.n296 161.3
R8178 commonsourceibias.n295 commonsourceibias.n294 161.3
R8179 commonsourceibias.n293 commonsourceibias.n276 161.3
R8180 commonsourceibias.n292 commonsourceibias.n291 161.3
R8181 commonsourceibias.n290 commonsourceibias.n289 161.3
R8182 commonsourceibias.n288 commonsourceibias.n278 161.3
R8183 commonsourceibias.n287 commonsourceibias.n286 161.3
R8184 commonsourceibias.n285 commonsourceibias.n284 161.3
R8185 commonsourceibias.n283 commonsourceibias.n280 161.3
R8186 commonsourceibias.n377 commonsourceibias.n273 161.3
R8187 commonsourceibias.n401 commonsourceibias.n266 161.3
R8188 commonsourceibias.n400 commonsourceibias.n399 161.3
R8189 commonsourceibias.n398 commonsourceibias.n397 161.3
R8190 commonsourceibias.n396 commonsourceibias.n268 161.3
R8191 commonsourceibias.n394 commonsourceibias.n393 161.3
R8192 commonsourceibias.n392 commonsourceibias.n269 161.3
R8193 commonsourceibias.n391 commonsourceibias.n390 161.3
R8194 commonsourceibias.n388 commonsourceibias.n270 161.3
R8195 commonsourceibias.n387 commonsourceibias.n386 161.3
R8196 commonsourceibias.n385 commonsourceibias.n271 161.3
R8197 commonsourceibias.n384 commonsourceibias.n383 161.3
R8198 commonsourceibias.n381 commonsourceibias.n272 161.3
R8199 commonsourceibias.n379 commonsourceibias.n378 161.3
R8200 commonsourceibias.n528 commonsourceibias.n468 161.3
R8201 commonsourceibias.n527 commonsourceibias.n526 161.3
R8202 commonsourceibias.n525 commonsourceibias.n524 161.3
R8203 commonsourceibias.n523 commonsourceibias.n470 161.3
R8204 commonsourceibias.n521 commonsourceibias.n520 161.3
R8205 commonsourceibias.n519 commonsourceibias.n471 161.3
R8206 commonsourceibias.n518 commonsourceibias.n517 161.3
R8207 commonsourceibias.n515 commonsourceibias.n472 161.3
R8208 commonsourceibias.n514 commonsourceibias.n513 161.3
R8209 commonsourceibias.n512 commonsourceibias.n473 161.3
R8210 commonsourceibias.n511 commonsourceibias.n510 161.3
R8211 commonsourceibias.n508 commonsourceibias.n474 161.3
R8212 commonsourceibias.n506 commonsourceibias.n505 161.3
R8213 commonsourceibias.n504 commonsourceibias.n475 161.3
R8214 commonsourceibias.n503 commonsourceibias.n502 161.3
R8215 commonsourceibias.n500 commonsourceibias.n476 161.3
R8216 commonsourceibias.n499 commonsourceibias.n498 161.3
R8217 commonsourceibias.n497 commonsourceibias.n496 161.3
R8218 commonsourceibias.n495 commonsourceibias.n478 161.3
R8219 commonsourceibias.n494 commonsourceibias.n493 161.3
R8220 commonsourceibias.n492 commonsourceibias.n491 161.3
R8221 commonsourceibias.n490 commonsourceibias.n480 161.3
R8222 commonsourceibias.n489 commonsourceibias.n488 161.3
R8223 commonsourceibias.n487 commonsourceibias.n486 161.3
R8224 commonsourceibias.n485 commonsourceibias.n482 161.3
R8225 commonsourceibias.n464 commonsourceibias.n404 161.3
R8226 commonsourceibias.n463 commonsourceibias.n462 161.3
R8227 commonsourceibias.n461 commonsourceibias.n460 161.3
R8228 commonsourceibias.n459 commonsourceibias.n406 161.3
R8229 commonsourceibias.n457 commonsourceibias.n456 161.3
R8230 commonsourceibias.n455 commonsourceibias.n407 161.3
R8231 commonsourceibias.n454 commonsourceibias.n453 161.3
R8232 commonsourceibias.n451 commonsourceibias.n408 161.3
R8233 commonsourceibias.n450 commonsourceibias.n449 161.3
R8234 commonsourceibias.n448 commonsourceibias.n409 161.3
R8235 commonsourceibias.n447 commonsourceibias.n446 161.3
R8236 commonsourceibias.n444 commonsourceibias.n410 161.3
R8237 commonsourceibias.n442 commonsourceibias.n441 161.3
R8238 commonsourceibias.n440 commonsourceibias.n411 161.3
R8239 commonsourceibias.n439 commonsourceibias.n438 161.3
R8240 commonsourceibias.n436 commonsourceibias.n412 161.3
R8241 commonsourceibias.n435 commonsourceibias.n434 161.3
R8242 commonsourceibias.n433 commonsourceibias.n432 161.3
R8243 commonsourceibias.n431 commonsourceibias.n414 161.3
R8244 commonsourceibias.n430 commonsourceibias.n429 161.3
R8245 commonsourceibias.n428 commonsourceibias.n427 161.3
R8246 commonsourceibias.n426 commonsourceibias.n416 161.3
R8247 commonsourceibias.n425 commonsourceibias.n424 161.3
R8248 commonsourceibias.n423 commonsourceibias.n422 161.3
R8249 commonsourceibias.n421 commonsourceibias.n418 161.3
R8250 commonsourceibias.n80 commonsourceibias.n78 81.5057
R8251 commonsourceibias.n304 commonsourceibias.n302 81.5057
R8252 commonsourceibias.n80 commonsourceibias.n79 80.9324
R8253 commonsourceibias.n82 commonsourceibias.n81 80.9324
R8254 commonsourceibias.n77 commonsourceibias.n76 80.9324
R8255 commonsourceibias.n75 commonsourceibias.n74 80.9324
R8256 commonsourceibias.n73 commonsourceibias.n72 80.9324
R8257 commonsourceibias.n371 commonsourceibias.n370 80.9324
R8258 commonsourceibias.n373 commonsourceibias.n372 80.9324
R8259 commonsourceibias.n375 commonsourceibias.n374 80.9324
R8260 commonsourceibias.n306 commonsourceibias.n305 80.9324
R8261 commonsourceibias.n304 commonsourceibias.n303 80.9324
R8262 commonsourceibias.n71 commonsourceibias.n70 80.6037
R8263 commonsourceibias.n137 commonsourceibias.n136 80.6037
R8264 commonsourceibias.n264 commonsourceibias.n263 80.6037
R8265 commonsourceibias.n200 commonsourceibias.n199 80.6037
R8266 commonsourceibias.n369 commonsourceibias.n368 80.6037
R8267 commonsourceibias.n403 commonsourceibias.n402 80.6037
R8268 commonsourceibias.n530 commonsourceibias.n529 80.6037
R8269 commonsourceibias.n466 commonsourceibias.n465 80.6037
R8270 commonsourceibias.n65 commonsourceibias.n64 56.5617
R8271 commonsourceibias.n51 commonsourceibias.n50 56.5617
R8272 commonsourceibias.n42 commonsourceibias.n41 56.5617
R8273 commonsourceibias.n28 commonsourceibias.n27 56.5617
R8274 commonsourceibias.n131 commonsourceibias.n130 56.5617
R8275 commonsourceibias.n117 commonsourceibias.n116 56.5617
R8276 commonsourceibias.n108 commonsourceibias.n107 56.5617
R8277 commonsourceibias.n94 commonsourceibias.n93 56.5617
R8278 commonsourceibias.n221 commonsourceibias.n220 56.5617
R8279 commonsourceibias.n235 commonsourceibias.n234 56.5617
R8280 commonsourceibias.n244 commonsourceibias.n243 56.5617
R8281 commonsourceibias.n258 commonsourceibias.n257 56.5617
R8282 commonsourceibias.n194 commonsourceibias.n193 56.5617
R8283 commonsourceibias.n180 commonsourceibias.n179 56.5617
R8284 commonsourceibias.n171 commonsourceibias.n170 56.5617
R8285 commonsourceibias.n157 commonsourceibias.n156 56.5617
R8286 commonsourceibias.n325 commonsourceibias.n324 56.5617
R8287 commonsourceibias.n339 commonsourceibias.n338 56.5617
R8288 commonsourceibias.n349 commonsourceibias.n347 56.5617
R8289 commonsourceibias.n363 commonsourceibias.n362 56.5617
R8290 commonsourceibias.n397 commonsourceibias.n396 56.5617
R8291 commonsourceibias.n383 commonsourceibias.n381 56.5617
R8292 commonsourceibias.n284 commonsourceibias.n283 56.5617
R8293 commonsourceibias.n298 commonsourceibias.n297 56.5617
R8294 commonsourceibias.n486 commonsourceibias.n485 56.5617
R8295 commonsourceibias.n500 commonsourceibias.n499 56.5617
R8296 commonsourceibias.n510 commonsourceibias.n508 56.5617
R8297 commonsourceibias.n524 commonsourceibias.n523 56.5617
R8298 commonsourceibias.n422 commonsourceibias.n421 56.5617
R8299 commonsourceibias.n436 commonsourceibias.n435 56.5617
R8300 commonsourceibias.n446 commonsourceibias.n444 56.5617
R8301 commonsourceibias.n460 commonsourceibias.n459 56.5617
R8302 commonsourceibias.n56 commonsourceibias.n55 56.0773
R8303 commonsourceibias.n37 commonsourceibias.n36 56.0773
R8304 commonsourceibias.n122 commonsourceibias.n121 56.0773
R8305 commonsourceibias.n103 commonsourceibias.n102 56.0773
R8306 commonsourceibias.n230 commonsourceibias.n229 56.0773
R8307 commonsourceibias.n249 commonsourceibias.n248 56.0773
R8308 commonsourceibias.n185 commonsourceibias.n184 56.0773
R8309 commonsourceibias.n166 commonsourceibias.n165 56.0773
R8310 commonsourceibias.n334 commonsourceibias.n333 56.0773
R8311 commonsourceibias.n354 commonsourceibias.n353 56.0773
R8312 commonsourceibias.n388 commonsourceibias.n387 56.0773
R8313 commonsourceibias.n293 commonsourceibias.n292 56.0773
R8314 commonsourceibias.n495 commonsourceibias.n494 56.0773
R8315 commonsourceibias.n515 commonsourceibias.n514 56.0773
R8316 commonsourceibias.n431 commonsourceibias.n430 56.0773
R8317 commonsourceibias.n451 commonsourceibias.n450 56.0773
R8318 commonsourceibias.n70 commonsourceibias.n69 46.0096
R8319 commonsourceibias.n136 commonsourceibias.n135 46.0096
R8320 commonsourceibias.n263 commonsourceibias.n262 46.0096
R8321 commonsourceibias.n199 commonsourceibias.n198 46.0096
R8322 commonsourceibias.n368 commonsourceibias.n367 46.0096
R8323 commonsourceibias.n402 commonsourceibias.n401 46.0096
R8324 commonsourceibias.n529 commonsourceibias.n528 46.0096
R8325 commonsourceibias.n465 commonsourceibias.n464 46.0096
R8326 commonsourceibias.n58 commonsourceibias.n12 41.5458
R8327 commonsourceibias.n33 commonsourceibias.n32 41.5458
R8328 commonsourceibias.n124 commonsourceibias.n3 41.5458
R8329 commonsourceibias.n99 commonsourceibias.n98 41.5458
R8330 commonsourceibias.n226 commonsourceibias.n225 41.5458
R8331 commonsourceibias.n251 commonsourceibias.n205 41.5458
R8332 commonsourceibias.n187 commonsourceibias.n141 41.5458
R8333 commonsourceibias.n162 commonsourceibias.n161 41.5458
R8334 commonsourceibias.n330 commonsourceibias.n329 41.5458
R8335 commonsourceibias.n356 commonsourceibias.n310 41.5458
R8336 commonsourceibias.n390 commonsourceibias.n269 41.5458
R8337 commonsourceibias.n289 commonsourceibias.n288 41.5458
R8338 commonsourceibias.n491 commonsourceibias.n490 41.5458
R8339 commonsourceibias.n517 commonsourceibias.n471 41.5458
R8340 commonsourceibias.n427 commonsourceibias.n426 41.5458
R8341 commonsourceibias.n453 commonsourceibias.n407 41.5458
R8342 commonsourceibias.n48 commonsourceibias.n17 40.577
R8343 commonsourceibias.n44 commonsourceibias.n17 40.577
R8344 commonsourceibias.n114 commonsourceibias.n8 40.577
R8345 commonsourceibias.n110 commonsourceibias.n8 40.577
R8346 commonsourceibias.n237 commonsourceibias.n210 40.577
R8347 commonsourceibias.n241 commonsourceibias.n210 40.577
R8348 commonsourceibias.n177 commonsourceibias.n146 40.577
R8349 commonsourceibias.n173 commonsourceibias.n146 40.577
R8350 commonsourceibias.n341 commonsourceibias.n314 40.577
R8351 commonsourceibias.n345 commonsourceibias.n314 40.577
R8352 commonsourceibias.n379 commonsourceibias.n273 40.577
R8353 commonsourceibias.n300 commonsourceibias.n273 40.577
R8354 commonsourceibias.n502 commonsourceibias.n475 40.577
R8355 commonsourceibias.n506 commonsourceibias.n475 40.577
R8356 commonsourceibias.n438 commonsourceibias.n411 40.577
R8357 commonsourceibias.n442 commonsourceibias.n411 40.577
R8358 commonsourceibias.n62 commonsourceibias.n12 39.6083
R8359 commonsourceibias.n32 commonsourceibias.n31 39.6083
R8360 commonsourceibias.n128 commonsourceibias.n3 39.6083
R8361 commonsourceibias.n98 commonsourceibias.n97 39.6083
R8362 commonsourceibias.n225 commonsourceibias.n224 39.6083
R8363 commonsourceibias.n255 commonsourceibias.n205 39.6083
R8364 commonsourceibias.n191 commonsourceibias.n141 39.6083
R8365 commonsourceibias.n161 commonsourceibias.n160 39.6083
R8366 commonsourceibias.n329 commonsourceibias.n328 39.6083
R8367 commonsourceibias.n360 commonsourceibias.n310 39.6083
R8368 commonsourceibias.n394 commonsourceibias.n269 39.6083
R8369 commonsourceibias.n288 commonsourceibias.n287 39.6083
R8370 commonsourceibias.n490 commonsourceibias.n489 39.6083
R8371 commonsourceibias.n521 commonsourceibias.n471 39.6083
R8372 commonsourceibias.n426 commonsourceibias.n425 39.6083
R8373 commonsourceibias.n457 commonsourceibias.n407 39.6083
R8374 commonsourceibias.n26 commonsourceibias.n25 33.0515
R8375 commonsourceibias.n92 commonsourceibias.n91 33.0515
R8376 commonsourceibias.n155 commonsourceibias.n154 33.0515
R8377 commonsourceibias.n219 commonsourceibias.n218 33.0515
R8378 commonsourceibias.n323 commonsourceibias.n322 33.0515
R8379 commonsourceibias.n282 commonsourceibias.n281 33.0515
R8380 commonsourceibias.n484 commonsourceibias.n483 33.0515
R8381 commonsourceibias.n420 commonsourceibias.n419 33.0515
R8382 commonsourceibias.n25 commonsourceibias.n24 28.5514
R8383 commonsourceibias.n91 commonsourceibias.n90 28.5514
R8384 commonsourceibias.n218 commonsourceibias.n217 28.5514
R8385 commonsourceibias.n154 commonsourceibias.n153 28.5514
R8386 commonsourceibias.n322 commonsourceibias.n321 28.5514
R8387 commonsourceibias.n281 commonsourceibias.n280 28.5514
R8388 commonsourceibias.n483 commonsourceibias.n482 28.5514
R8389 commonsourceibias.n419 commonsourceibias.n418 28.5514
R8390 commonsourceibias.n69 commonsourceibias.n68 26.0455
R8391 commonsourceibias.n135 commonsourceibias.n134 26.0455
R8392 commonsourceibias.n262 commonsourceibias.n261 26.0455
R8393 commonsourceibias.n198 commonsourceibias.n197 26.0455
R8394 commonsourceibias.n367 commonsourceibias.n366 26.0455
R8395 commonsourceibias.n401 commonsourceibias.n400 26.0455
R8396 commonsourceibias.n528 commonsourceibias.n527 26.0455
R8397 commonsourceibias.n464 commonsourceibias.n463 26.0455
R8398 commonsourceibias.n55 commonsourceibias.n14 25.0767
R8399 commonsourceibias.n38 commonsourceibias.n37 25.0767
R8400 commonsourceibias.n121 commonsourceibias.n5 25.0767
R8401 commonsourceibias.n104 commonsourceibias.n103 25.0767
R8402 commonsourceibias.n231 commonsourceibias.n230 25.0767
R8403 commonsourceibias.n248 commonsourceibias.n207 25.0767
R8404 commonsourceibias.n184 commonsourceibias.n143 25.0767
R8405 commonsourceibias.n167 commonsourceibias.n166 25.0767
R8406 commonsourceibias.n335 commonsourceibias.n334 25.0767
R8407 commonsourceibias.n353 commonsourceibias.n312 25.0767
R8408 commonsourceibias.n387 commonsourceibias.n271 25.0767
R8409 commonsourceibias.n294 commonsourceibias.n293 25.0767
R8410 commonsourceibias.n496 commonsourceibias.n495 25.0767
R8411 commonsourceibias.n514 commonsourceibias.n473 25.0767
R8412 commonsourceibias.n432 commonsourceibias.n431 25.0767
R8413 commonsourceibias.n450 commonsourceibias.n409 25.0767
R8414 commonsourceibias.n51 commonsourceibias.n16 24.3464
R8415 commonsourceibias.n41 commonsourceibias.n19 24.3464
R8416 commonsourceibias.n117 commonsourceibias.n7 24.3464
R8417 commonsourceibias.n107 commonsourceibias.n85 24.3464
R8418 commonsourceibias.n234 commonsourceibias.n212 24.3464
R8419 commonsourceibias.n244 commonsourceibias.n209 24.3464
R8420 commonsourceibias.n180 commonsourceibias.n145 24.3464
R8421 commonsourceibias.n170 commonsourceibias.n148 24.3464
R8422 commonsourceibias.n338 commonsourceibias.n316 24.3464
R8423 commonsourceibias.n349 commonsourceibias.n348 24.3464
R8424 commonsourceibias.n383 commonsourceibias.n382 24.3464
R8425 commonsourceibias.n297 commonsourceibias.n275 24.3464
R8426 commonsourceibias.n499 commonsourceibias.n477 24.3464
R8427 commonsourceibias.n510 commonsourceibias.n509 24.3464
R8428 commonsourceibias.n435 commonsourceibias.n413 24.3464
R8429 commonsourceibias.n446 commonsourceibias.n445 24.3464
R8430 commonsourceibias.n65 commonsourceibias.n10 23.8546
R8431 commonsourceibias.n27 commonsourceibias.n26 23.8546
R8432 commonsourceibias.n131 commonsourceibias.n1 23.8546
R8433 commonsourceibias.n93 commonsourceibias.n92 23.8546
R8434 commonsourceibias.n220 commonsourceibias.n219 23.8546
R8435 commonsourceibias.n258 commonsourceibias.n203 23.8546
R8436 commonsourceibias.n194 commonsourceibias.n139 23.8546
R8437 commonsourceibias.n156 commonsourceibias.n155 23.8546
R8438 commonsourceibias.n324 commonsourceibias.n323 23.8546
R8439 commonsourceibias.n363 commonsourceibias.n308 23.8546
R8440 commonsourceibias.n397 commonsourceibias.n267 23.8546
R8441 commonsourceibias.n283 commonsourceibias.n282 23.8546
R8442 commonsourceibias.n485 commonsourceibias.n484 23.8546
R8443 commonsourceibias.n524 commonsourceibias.n469 23.8546
R8444 commonsourceibias.n421 commonsourceibias.n420 23.8546
R8445 commonsourceibias.n460 commonsourceibias.n405 23.8546
R8446 commonsourceibias.n64 commonsourceibias.n63 16.9689
R8447 commonsourceibias.n28 commonsourceibias.n23 16.9689
R8448 commonsourceibias.n130 commonsourceibias.n129 16.9689
R8449 commonsourceibias.n94 commonsourceibias.n89 16.9689
R8450 commonsourceibias.n221 commonsourceibias.n216 16.9689
R8451 commonsourceibias.n257 commonsourceibias.n256 16.9689
R8452 commonsourceibias.n193 commonsourceibias.n192 16.9689
R8453 commonsourceibias.n157 commonsourceibias.n152 16.9689
R8454 commonsourceibias.n325 commonsourceibias.n320 16.9689
R8455 commonsourceibias.n362 commonsourceibias.n361 16.9689
R8456 commonsourceibias.n396 commonsourceibias.n395 16.9689
R8457 commonsourceibias.n284 commonsourceibias.n279 16.9689
R8458 commonsourceibias.n486 commonsourceibias.n481 16.9689
R8459 commonsourceibias.n523 commonsourceibias.n522 16.9689
R8460 commonsourceibias.n422 commonsourceibias.n417 16.9689
R8461 commonsourceibias.n459 commonsourceibias.n458 16.9689
R8462 commonsourceibias.n50 commonsourceibias.n49 16.477
R8463 commonsourceibias.n43 commonsourceibias.n42 16.477
R8464 commonsourceibias.n116 commonsourceibias.n115 16.477
R8465 commonsourceibias.n109 commonsourceibias.n108 16.477
R8466 commonsourceibias.n236 commonsourceibias.n235 16.477
R8467 commonsourceibias.n243 commonsourceibias.n242 16.477
R8468 commonsourceibias.n179 commonsourceibias.n178 16.477
R8469 commonsourceibias.n172 commonsourceibias.n171 16.477
R8470 commonsourceibias.n340 commonsourceibias.n339 16.477
R8471 commonsourceibias.n347 commonsourceibias.n346 16.477
R8472 commonsourceibias.n381 commonsourceibias.n380 16.477
R8473 commonsourceibias.n299 commonsourceibias.n298 16.477
R8474 commonsourceibias.n501 commonsourceibias.n500 16.477
R8475 commonsourceibias.n508 commonsourceibias.n507 16.477
R8476 commonsourceibias.n437 commonsourceibias.n436 16.477
R8477 commonsourceibias.n444 commonsourceibias.n443 16.477
R8478 commonsourceibias.n57 commonsourceibias.n56 15.9852
R8479 commonsourceibias.n36 commonsourceibias.n21 15.9852
R8480 commonsourceibias.n123 commonsourceibias.n122 15.9852
R8481 commonsourceibias.n102 commonsourceibias.n87 15.9852
R8482 commonsourceibias.n229 commonsourceibias.n214 15.9852
R8483 commonsourceibias.n250 commonsourceibias.n249 15.9852
R8484 commonsourceibias.n186 commonsourceibias.n185 15.9852
R8485 commonsourceibias.n165 commonsourceibias.n150 15.9852
R8486 commonsourceibias.n333 commonsourceibias.n318 15.9852
R8487 commonsourceibias.n355 commonsourceibias.n354 15.9852
R8488 commonsourceibias.n389 commonsourceibias.n388 15.9852
R8489 commonsourceibias.n292 commonsourceibias.n277 15.9852
R8490 commonsourceibias.n494 commonsourceibias.n479 15.9852
R8491 commonsourceibias.n516 commonsourceibias.n515 15.9852
R8492 commonsourceibias.n430 commonsourceibias.n415 15.9852
R8493 commonsourceibias.n452 commonsourceibias.n451 15.9852
R8494 commonsourceibias.n73 commonsourceibias.n71 13.2057
R8495 commonsourceibias.n371 commonsourceibias.n369 13.2057
R8496 commonsourceibias.n532 commonsourceibias.n265 10.122
R8497 commonsourceibias.n112 commonsourceibias.n83 9.50363
R8498 commonsourceibias.n377 commonsourceibias.n376 9.50363
R8499 commonsourceibias.n201 commonsourceibias.n137 8.7339
R8500 commonsourceibias.n467 commonsourceibias.n403 8.7339
R8501 commonsourceibias.n58 commonsourceibias.n57 8.60764
R8502 commonsourceibias.n33 commonsourceibias.n21 8.60764
R8503 commonsourceibias.n124 commonsourceibias.n123 8.60764
R8504 commonsourceibias.n99 commonsourceibias.n87 8.60764
R8505 commonsourceibias.n226 commonsourceibias.n214 8.60764
R8506 commonsourceibias.n251 commonsourceibias.n250 8.60764
R8507 commonsourceibias.n187 commonsourceibias.n186 8.60764
R8508 commonsourceibias.n162 commonsourceibias.n150 8.60764
R8509 commonsourceibias.n330 commonsourceibias.n318 8.60764
R8510 commonsourceibias.n356 commonsourceibias.n355 8.60764
R8511 commonsourceibias.n390 commonsourceibias.n389 8.60764
R8512 commonsourceibias.n289 commonsourceibias.n277 8.60764
R8513 commonsourceibias.n491 commonsourceibias.n479 8.60764
R8514 commonsourceibias.n517 commonsourceibias.n516 8.60764
R8515 commonsourceibias.n427 commonsourceibias.n415 8.60764
R8516 commonsourceibias.n453 commonsourceibias.n452 8.60764
R8517 commonsourceibias.n532 commonsourceibias.n531 8.46921
R8518 commonsourceibias.n49 commonsourceibias.n48 8.11581
R8519 commonsourceibias.n44 commonsourceibias.n43 8.11581
R8520 commonsourceibias.n115 commonsourceibias.n114 8.11581
R8521 commonsourceibias.n110 commonsourceibias.n109 8.11581
R8522 commonsourceibias.n237 commonsourceibias.n236 8.11581
R8523 commonsourceibias.n242 commonsourceibias.n241 8.11581
R8524 commonsourceibias.n178 commonsourceibias.n177 8.11581
R8525 commonsourceibias.n173 commonsourceibias.n172 8.11581
R8526 commonsourceibias.n341 commonsourceibias.n340 8.11581
R8527 commonsourceibias.n346 commonsourceibias.n345 8.11581
R8528 commonsourceibias.n380 commonsourceibias.n379 8.11581
R8529 commonsourceibias.n300 commonsourceibias.n299 8.11581
R8530 commonsourceibias.n502 commonsourceibias.n501 8.11581
R8531 commonsourceibias.n507 commonsourceibias.n506 8.11581
R8532 commonsourceibias.n438 commonsourceibias.n437 8.11581
R8533 commonsourceibias.n443 commonsourceibias.n442 8.11581
R8534 commonsourceibias.n63 commonsourceibias.n62 7.62397
R8535 commonsourceibias.n31 commonsourceibias.n23 7.62397
R8536 commonsourceibias.n129 commonsourceibias.n128 7.62397
R8537 commonsourceibias.n97 commonsourceibias.n89 7.62397
R8538 commonsourceibias.n224 commonsourceibias.n216 7.62397
R8539 commonsourceibias.n256 commonsourceibias.n255 7.62397
R8540 commonsourceibias.n192 commonsourceibias.n191 7.62397
R8541 commonsourceibias.n160 commonsourceibias.n152 7.62397
R8542 commonsourceibias.n328 commonsourceibias.n320 7.62397
R8543 commonsourceibias.n361 commonsourceibias.n360 7.62397
R8544 commonsourceibias.n395 commonsourceibias.n394 7.62397
R8545 commonsourceibias.n287 commonsourceibias.n279 7.62397
R8546 commonsourceibias.n489 commonsourceibias.n481 7.62397
R8547 commonsourceibias.n522 commonsourceibias.n521 7.62397
R8548 commonsourceibias.n425 commonsourceibias.n417 7.62397
R8549 commonsourceibias.n458 commonsourceibias.n457 7.62397
R8550 commonsourceibias.n265 commonsourceibias.n264 5.00473
R8551 commonsourceibias.n201 commonsourceibias.n200 5.00473
R8552 commonsourceibias.n531 commonsourceibias.n530 5.00473
R8553 commonsourceibias.n467 commonsourceibias.n466 5.00473
R8554 commonsourceibias commonsourceibias.n532 3.97901
R8555 commonsourceibias.n265 commonsourceibias.n201 3.72967
R8556 commonsourceibias.n531 commonsourceibias.n467 3.72967
R8557 commonsourceibias.n78 commonsourceibias.t1 2.82907
R8558 commonsourceibias.n78 commonsourceibias.t31 2.82907
R8559 commonsourceibias.n79 commonsourceibias.t17 2.82907
R8560 commonsourceibias.n79 commonsourceibias.t27 2.82907
R8561 commonsourceibias.n81 commonsourceibias.t29 2.82907
R8562 commonsourceibias.n81 commonsourceibias.t47 2.82907
R8563 commonsourceibias.n76 commonsourceibias.t11 2.82907
R8564 commonsourceibias.n76 commonsourceibias.t41 2.82907
R8565 commonsourceibias.n74 commonsourceibias.t21 2.82907
R8566 commonsourceibias.n74 commonsourceibias.t43 2.82907
R8567 commonsourceibias.n72 commonsourceibias.t7 2.82907
R8568 commonsourceibias.n72 commonsourceibias.t25 2.82907
R8569 commonsourceibias.n370 commonsourceibias.t9 2.82907
R8570 commonsourceibias.n370 commonsourceibias.t35 2.82907
R8571 commonsourceibias.n372 commonsourceibias.t33 2.82907
R8572 commonsourceibias.n372 commonsourceibias.t15 2.82907
R8573 commonsourceibias.n374 commonsourceibias.t23 2.82907
R8574 commonsourceibias.n374 commonsourceibias.t19 2.82907
R8575 commonsourceibias.n305 commonsourceibias.t3 2.82907
R8576 commonsourceibias.n305 commonsourceibias.t45 2.82907
R8577 commonsourceibias.n303 commonsourceibias.t13 2.82907
R8578 commonsourceibias.n303 commonsourceibias.t37 2.82907
R8579 commonsourceibias.n302 commonsourceibias.t5 2.82907
R8580 commonsourceibias.n302 commonsourceibias.t39 2.82907
R8581 commonsourceibias.n68 commonsourceibias.n10 0.738255
R8582 commonsourceibias.n134 commonsourceibias.n1 0.738255
R8583 commonsourceibias.n261 commonsourceibias.n203 0.738255
R8584 commonsourceibias.n197 commonsourceibias.n139 0.738255
R8585 commonsourceibias.n366 commonsourceibias.n308 0.738255
R8586 commonsourceibias.n400 commonsourceibias.n267 0.738255
R8587 commonsourceibias.n527 commonsourceibias.n469 0.738255
R8588 commonsourceibias.n463 commonsourceibias.n405 0.738255
R8589 commonsourceibias.n75 commonsourceibias.n73 0.573776
R8590 commonsourceibias.n77 commonsourceibias.n75 0.573776
R8591 commonsourceibias.n82 commonsourceibias.n80 0.573776
R8592 commonsourceibias.n306 commonsourceibias.n304 0.573776
R8593 commonsourceibias.n375 commonsourceibias.n373 0.573776
R8594 commonsourceibias.n373 commonsourceibias.n371 0.573776
R8595 commonsourceibias.n83 commonsourceibias.n77 0.287138
R8596 commonsourceibias.n83 commonsourceibias.n82 0.287138
R8597 commonsourceibias.n376 commonsourceibias.n306 0.287138
R8598 commonsourceibias.n376 commonsourceibias.n375 0.287138
R8599 commonsourceibias.n71 commonsourceibias.n9 0.285035
R8600 commonsourceibias.n137 commonsourceibias.n0 0.285035
R8601 commonsourceibias.n264 commonsourceibias.n202 0.285035
R8602 commonsourceibias.n200 commonsourceibias.n138 0.285035
R8603 commonsourceibias.n369 commonsourceibias.n307 0.285035
R8604 commonsourceibias.n403 commonsourceibias.n266 0.285035
R8605 commonsourceibias.n530 commonsourceibias.n468 0.285035
R8606 commonsourceibias.n466 commonsourceibias.n404 0.285035
R8607 commonsourceibias.n16 commonsourceibias.n14 0.246418
R8608 commonsourceibias.n38 commonsourceibias.n19 0.246418
R8609 commonsourceibias.n7 commonsourceibias.n5 0.246418
R8610 commonsourceibias.n104 commonsourceibias.n85 0.246418
R8611 commonsourceibias.n231 commonsourceibias.n212 0.246418
R8612 commonsourceibias.n209 commonsourceibias.n207 0.246418
R8613 commonsourceibias.n145 commonsourceibias.n143 0.246418
R8614 commonsourceibias.n167 commonsourceibias.n148 0.246418
R8615 commonsourceibias.n335 commonsourceibias.n316 0.246418
R8616 commonsourceibias.n348 commonsourceibias.n312 0.246418
R8617 commonsourceibias.n382 commonsourceibias.n271 0.246418
R8618 commonsourceibias.n294 commonsourceibias.n275 0.246418
R8619 commonsourceibias.n496 commonsourceibias.n477 0.246418
R8620 commonsourceibias.n509 commonsourceibias.n473 0.246418
R8621 commonsourceibias.n432 commonsourceibias.n413 0.246418
R8622 commonsourceibias.n445 commonsourceibias.n409 0.246418
R8623 commonsourceibias.n67 commonsourceibias.n9 0.189894
R8624 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8625 commonsourceibias.n66 commonsourceibias.n11 0.189894
R8626 commonsourceibias.n61 commonsourceibias.n11 0.189894
R8627 commonsourceibias.n61 commonsourceibias.n60 0.189894
R8628 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8629 commonsourceibias.n59 commonsourceibias.n13 0.189894
R8630 commonsourceibias.n54 commonsourceibias.n13 0.189894
R8631 commonsourceibias.n54 commonsourceibias.n53 0.189894
R8632 commonsourceibias.n53 commonsourceibias.n52 0.189894
R8633 commonsourceibias.n52 commonsourceibias.n15 0.189894
R8634 commonsourceibias.n47 commonsourceibias.n15 0.189894
R8635 commonsourceibias.n47 commonsourceibias.n46 0.189894
R8636 commonsourceibias.n46 commonsourceibias.n45 0.189894
R8637 commonsourceibias.n45 commonsourceibias.n18 0.189894
R8638 commonsourceibias.n40 commonsourceibias.n18 0.189894
R8639 commonsourceibias.n40 commonsourceibias.n39 0.189894
R8640 commonsourceibias.n39 commonsourceibias.n20 0.189894
R8641 commonsourceibias.n35 commonsourceibias.n20 0.189894
R8642 commonsourceibias.n35 commonsourceibias.n34 0.189894
R8643 commonsourceibias.n34 commonsourceibias.n22 0.189894
R8644 commonsourceibias.n30 commonsourceibias.n22 0.189894
R8645 commonsourceibias.n30 commonsourceibias.n29 0.189894
R8646 commonsourceibias.n29 commonsourceibias.n24 0.189894
R8647 commonsourceibias.n111 commonsourceibias.n84 0.189894
R8648 commonsourceibias.n106 commonsourceibias.n84 0.189894
R8649 commonsourceibias.n106 commonsourceibias.n105 0.189894
R8650 commonsourceibias.n105 commonsourceibias.n86 0.189894
R8651 commonsourceibias.n101 commonsourceibias.n86 0.189894
R8652 commonsourceibias.n101 commonsourceibias.n100 0.189894
R8653 commonsourceibias.n100 commonsourceibias.n88 0.189894
R8654 commonsourceibias.n96 commonsourceibias.n88 0.189894
R8655 commonsourceibias.n96 commonsourceibias.n95 0.189894
R8656 commonsourceibias.n95 commonsourceibias.n90 0.189894
R8657 commonsourceibias.n133 commonsourceibias.n0 0.189894
R8658 commonsourceibias.n133 commonsourceibias.n132 0.189894
R8659 commonsourceibias.n132 commonsourceibias.n2 0.189894
R8660 commonsourceibias.n127 commonsourceibias.n2 0.189894
R8661 commonsourceibias.n127 commonsourceibias.n126 0.189894
R8662 commonsourceibias.n126 commonsourceibias.n125 0.189894
R8663 commonsourceibias.n125 commonsourceibias.n4 0.189894
R8664 commonsourceibias.n120 commonsourceibias.n4 0.189894
R8665 commonsourceibias.n120 commonsourceibias.n119 0.189894
R8666 commonsourceibias.n119 commonsourceibias.n118 0.189894
R8667 commonsourceibias.n118 commonsourceibias.n6 0.189894
R8668 commonsourceibias.n113 commonsourceibias.n6 0.189894
R8669 commonsourceibias.n260 commonsourceibias.n202 0.189894
R8670 commonsourceibias.n260 commonsourceibias.n259 0.189894
R8671 commonsourceibias.n259 commonsourceibias.n204 0.189894
R8672 commonsourceibias.n254 commonsourceibias.n204 0.189894
R8673 commonsourceibias.n254 commonsourceibias.n253 0.189894
R8674 commonsourceibias.n253 commonsourceibias.n252 0.189894
R8675 commonsourceibias.n252 commonsourceibias.n206 0.189894
R8676 commonsourceibias.n247 commonsourceibias.n206 0.189894
R8677 commonsourceibias.n247 commonsourceibias.n246 0.189894
R8678 commonsourceibias.n246 commonsourceibias.n245 0.189894
R8679 commonsourceibias.n245 commonsourceibias.n208 0.189894
R8680 commonsourceibias.n240 commonsourceibias.n208 0.189894
R8681 commonsourceibias.n240 commonsourceibias.n239 0.189894
R8682 commonsourceibias.n239 commonsourceibias.n238 0.189894
R8683 commonsourceibias.n238 commonsourceibias.n211 0.189894
R8684 commonsourceibias.n233 commonsourceibias.n211 0.189894
R8685 commonsourceibias.n233 commonsourceibias.n232 0.189894
R8686 commonsourceibias.n232 commonsourceibias.n213 0.189894
R8687 commonsourceibias.n228 commonsourceibias.n213 0.189894
R8688 commonsourceibias.n228 commonsourceibias.n227 0.189894
R8689 commonsourceibias.n227 commonsourceibias.n215 0.189894
R8690 commonsourceibias.n223 commonsourceibias.n215 0.189894
R8691 commonsourceibias.n223 commonsourceibias.n222 0.189894
R8692 commonsourceibias.n222 commonsourceibias.n217 0.189894
R8693 commonsourceibias.n196 commonsourceibias.n138 0.189894
R8694 commonsourceibias.n196 commonsourceibias.n195 0.189894
R8695 commonsourceibias.n195 commonsourceibias.n140 0.189894
R8696 commonsourceibias.n190 commonsourceibias.n140 0.189894
R8697 commonsourceibias.n190 commonsourceibias.n189 0.189894
R8698 commonsourceibias.n189 commonsourceibias.n188 0.189894
R8699 commonsourceibias.n188 commonsourceibias.n142 0.189894
R8700 commonsourceibias.n183 commonsourceibias.n142 0.189894
R8701 commonsourceibias.n183 commonsourceibias.n182 0.189894
R8702 commonsourceibias.n182 commonsourceibias.n181 0.189894
R8703 commonsourceibias.n181 commonsourceibias.n144 0.189894
R8704 commonsourceibias.n176 commonsourceibias.n144 0.189894
R8705 commonsourceibias.n176 commonsourceibias.n175 0.189894
R8706 commonsourceibias.n175 commonsourceibias.n174 0.189894
R8707 commonsourceibias.n174 commonsourceibias.n147 0.189894
R8708 commonsourceibias.n169 commonsourceibias.n147 0.189894
R8709 commonsourceibias.n169 commonsourceibias.n168 0.189894
R8710 commonsourceibias.n168 commonsourceibias.n149 0.189894
R8711 commonsourceibias.n164 commonsourceibias.n149 0.189894
R8712 commonsourceibias.n164 commonsourceibias.n163 0.189894
R8713 commonsourceibias.n163 commonsourceibias.n151 0.189894
R8714 commonsourceibias.n159 commonsourceibias.n151 0.189894
R8715 commonsourceibias.n159 commonsourceibias.n158 0.189894
R8716 commonsourceibias.n158 commonsourceibias.n153 0.189894
R8717 commonsourceibias.n326 commonsourceibias.n321 0.189894
R8718 commonsourceibias.n327 commonsourceibias.n326 0.189894
R8719 commonsourceibias.n327 commonsourceibias.n319 0.189894
R8720 commonsourceibias.n331 commonsourceibias.n319 0.189894
R8721 commonsourceibias.n332 commonsourceibias.n331 0.189894
R8722 commonsourceibias.n332 commonsourceibias.n317 0.189894
R8723 commonsourceibias.n336 commonsourceibias.n317 0.189894
R8724 commonsourceibias.n337 commonsourceibias.n336 0.189894
R8725 commonsourceibias.n337 commonsourceibias.n315 0.189894
R8726 commonsourceibias.n342 commonsourceibias.n315 0.189894
R8727 commonsourceibias.n343 commonsourceibias.n342 0.189894
R8728 commonsourceibias.n344 commonsourceibias.n343 0.189894
R8729 commonsourceibias.n344 commonsourceibias.n313 0.189894
R8730 commonsourceibias.n350 commonsourceibias.n313 0.189894
R8731 commonsourceibias.n351 commonsourceibias.n350 0.189894
R8732 commonsourceibias.n352 commonsourceibias.n351 0.189894
R8733 commonsourceibias.n352 commonsourceibias.n311 0.189894
R8734 commonsourceibias.n357 commonsourceibias.n311 0.189894
R8735 commonsourceibias.n358 commonsourceibias.n357 0.189894
R8736 commonsourceibias.n359 commonsourceibias.n358 0.189894
R8737 commonsourceibias.n359 commonsourceibias.n309 0.189894
R8738 commonsourceibias.n364 commonsourceibias.n309 0.189894
R8739 commonsourceibias.n365 commonsourceibias.n364 0.189894
R8740 commonsourceibias.n365 commonsourceibias.n307 0.189894
R8741 commonsourceibias.n285 commonsourceibias.n280 0.189894
R8742 commonsourceibias.n286 commonsourceibias.n285 0.189894
R8743 commonsourceibias.n286 commonsourceibias.n278 0.189894
R8744 commonsourceibias.n290 commonsourceibias.n278 0.189894
R8745 commonsourceibias.n291 commonsourceibias.n290 0.189894
R8746 commonsourceibias.n291 commonsourceibias.n276 0.189894
R8747 commonsourceibias.n295 commonsourceibias.n276 0.189894
R8748 commonsourceibias.n296 commonsourceibias.n295 0.189894
R8749 commonsourceibias.n296 commonsourceibias.n274 0.189894
R8750 commonsourceibias.n301 commonsourceibias.n274 0.189894
R8751 commonsourceibias.n378 commonsourceibias.n272 0.189894
R8752 commonsourceibias.n384 commonsourceibias.n272 0.189894
R8753 commonsourceibias.n385 commonsourceibias.n384 0.189894
R8754 commonsourceibias.n386 commonsourceibias.n385 0.189894
R8755 commonsourceibias.n386 commonsourceibias.n270 0.189894
R8756 commonsourceibias.n391 commonsourceibias.n270 0.189894
R8757 commonsourceibias.n392 commonsourceibias.n391 0.189894
R8758 commonsourceibias.n393 commonsourceibias.n392 0.189894
R8759 commonsourceibias.n393 commonsourceibias.n268 0.189894
R8760 commonsourceibias.n398 commonsourceibias.n268 0.189894
R8761 commonsourceibias.n399 commonsourceibias.n398 0.189894
R8762 commonsourceibias.n399 commonsourceibias.n266 0.189894
R8763 commonsourceibias.n487 commonsourceibias.n482 0.189894
R8764 commonsourceibias.n488 commonsourceibias.n487 0.189894
R8765 commonsourceibias.n488 commonsourceibias.n480 0.189894
R8766 commonsourceibias.n492 commonsourceibias.n480 0.189894
R8767 commonsourceibias.n493 commonsourceibias.n492 0.189894
R8768 commonsourceibias.n493 commonsourceibias.n478 0.189894
R8769 commonsourceibias.n497 commonsourceibias.n478 0.189894
R8770 commonsourceibias.n498 commonsourceibias.n497 0.189894
R8771 commonsourceibias.n498 commonsourceibias.n476 0.189894
R8772 commonsourceibias.n503 commonsourceibias.n476 0.189894
R8773 commonsourceibias.n504 commonsourceibias.n503 0.189894
R8774 commonsourceibias.n505 commonsourceibias.n504 0.189894
R8775 commonsourceibias.n505 commonsourceibias.n474 0.189894
R8776 commonsourceibias.n511 commonsourceibias.n474 0.189894
R8777 commonsourceibias.n512 commonsourceibias.n511 0.189894
R8778 commonsourceibias.n513 commonsourceibias.n512 0.189894
R8779 commonsourceibias.n513 commonsourceibias.n472 0.189894
R8780 commonsourceibias.n518 commonsourceibias.n472 0.189894
R8781 commonsourceibias.n519 commonsourceibias.n518 0.189894
R8782 commonsourceibias.n520 commonsourceibias.n519 0.189894
R8783 commonsourceibias.n520 commonsourceibias.n470 0.189894
R8784 commonsourceibias.n525 commonsourceibias.n470 0.189894
R8785 commonsourceibias.n526 commonsourceibias.n525 0.189894
R8786 commonsourceibias.n526 commonsourceibias.n468 0.189894
R8787 commonsourceibias.n423 commonsourceibias.n418 0.189894
R8788 commonsourceibias.n424 commonsourceibias.n423 0.189894
R8789 commonsourceibias.n424 commonsourceibias.n416 0.189894
R8790 commonsourceibias.n428 commonsourceibias.n416 0.189894
R8791 commonsourceibias.n429 commonsourceibias.n428 0.189894
R8792 commonsourceibias.n429 commonsourceibias.n414 0.189894
R8793 commonsourceibias.n433 commonsourceibias.n414 0.189894
R8794 commonsourceibias.n434 commonsourceibias.n433 0.189894
R8795 commonsourceibias.n434 commonsourceibias.n412 0.189894
R8796 commonsourceibias.n439 commonsourceibias.n412 0.189894
R8797 commonsourceibias.n440 commonsourceibias.n439 0.189894
R8798 commonsourceibias.n441 commonsourceibias.n440 0.189894
R8799 commonsourceibias.n441 commonsourceibias.n410 0.189894
R8800 commonsourceibias.n447 commonsourceibias.n410 0.189894
R8801 commonsourceibias.n448 commonsourceibias.n447 0.189894
R8802 commonsourceibias.n449 commonsourceibias.n448 0.189894
R8803 commonsourceibias.n449 commonsourceibias.n408 0.189894
R8804 commonsourceibias.n454 commonsourceibias.n408 0.189894
R8805 commonsourceibias.n455 commonsourceibias.n454 0.189894
R8806 commonsourceibias.n456 commonsourceibias.n455 0.189894
R8807 commonsourceibias.n456 commonsourceibias.n406 0.189894
R8808 commonsourceibias.n461 commonsourceibias.n406 0.189894
R8809 commonsourceibias.n462 commonsourceibias.n461 0.189894
R8810 commonsourceibias.n462 commonsourceibias.n404 0.189894
R8811 commonsourceibias.n112 commonsourceibias.n111 0.170955
R8812 commonsourceibias.n113 commonsourceibias.n112 0.170955
R8813 commonsourceibias.n377 commonsourceibias.n301 0.170955
R8814 commonsourceibias.n378 commonsourceibias.n377 0.170955
R8815 gnd.n6891 gnd.n6890 1779.25
R8816 gnd.n6232 gnd.n2304 928.563
R8817 gnd.n7345 gnd.n171 838.452
R8818 gnd.n7332 gnd.n169 838.452
R8819 gnd.n2821 gnd.n2744 838.452
R8820 gnd.n5806 gnd.n5317 838.452
R8821 gnd.n6085 gnd.n2536 838.452
R8822 gnd.n3670 gnd.n2534 838.452
R8823 gnd.n3844 gnd.n2324 838.452
R8824 gnd.n3891 gnd.n2326 838.452
R8825 gnd.n7347 gnd.n166 783.196
R8826 gnd.n7207 gnd.n168 783.196
R8827 gnd.n5808 gnd.n2818 783.196
R8828 gnd.n5925 gnd.n2748 783.196
R8829 gnd.n6087 gnd.n2531 783.196
R8830 gnd.n4425 gnd.n2533 783.196
R8831 gnd.n4103 gnd.n2323 783.196
R8832 gnd.n6214 gnd.n2327 783.196
R8833 gnd.n3578 gnd.n2573 771.183
R8834 gnd.n5188 gnd.n5187 771.183
R8835 gnd.n6070 gnd.n2548 771.183
R8836 gnd.n5935 gnd.n2682 771.183
R8837 gnd.n2212 gnd.n843 766.379
R8838 gnd.n2215 gnd.n2214 766.379
R8839 gnd.n1452 gnd.n1355 766.379
R8840 gnd.n1448 gnd.n1353 766.379
R8841 gnd.n2303 gnd.n865 756.769
R8842 gnd.n2206 gnd.n2205 756.769
R8843 gnd.n1545 gnd.n1262 756.769
R8844 gnd.n1543 gnd.n1265 756.769
R8845 gnd.n6401 gnd.n671 703.915
R8846 gnd.n6892 gnd.n381 703.915
R8847 gnd.n7102 gnd.n251 703.915
R8848 gnd.n6233 gnd.n841 703.915
R8849 gnd.n6402 gnd.n6401 585
R8850 gnd.n6401 gnd.n6400 585
R8851 gnd.n675 gnd.n674 585
R8852 gnd.n6399 gnd.n675 585
R8853 gnd.n6397 gnd.n6396 585
R8854 gnd.n6398 gnd.n6397 585
R8855 gnd.n6395 gnd.n677 585
R8856 gnd.n677 gnd.n676 585
R8857 gnd.n6394 gnd.n6393 585
R8858 gnd.n6393 gnd.n6392 585
R8859 gnd.n682 gnd.n681 585
R8860 gnd.n6391 gnd.n682 585
R8861 gnd.n6389 gnd.n6388 585
R8862 gnd.n6390 gnd.n6389 585
R8863 gnd.n6387 gnd.n684 585
R8864 gnd.n684 gnd.n683 585
R8865 gnd.n6386 gnd.n6385 585
R8866 gnd.n6385 gnd.n6384 585
R8867 gnd.n690 gnd.n689 585
R8868 gnd.n6383 gnd.n690 585
R8869 gnd.n6381 gnd.n6380 585
R8870 gnd.n6382 gnd.n6381 585
R8871 gnd.n6379 gnd.n692 585
R8872 gnd.n692 gnd.n691 585
R8873 gnd.n6378 gnd.n6377 585
R8874 gnd.n6377 gnd.n6376 585
R8875 gnd.n698 gnd.n697 585
R8876 gnd.n6375 gnd.n698 585
R8877 gnd.n6373 gnd.n6372 585
R8878 gnd.n6374 gnd.n6373 585
R8879 gnd.n6371 gnd.n700 585
R8880 gnd.n700 gnd.n699 585
R8881 gnd.n6370 gnd.n6369 585
R8882 gnd.n6369 gnd.n6368 585
R8883 gnd.n706 gnd.n705 585
R8884 gnd.n6367 gnd.n706 585
R8885 gnd.n6365 gnd.n6364 585
R8886 gnd.n6366 gnd.n6365 585
R8887 gnd.n6363 gnd.n708 585
R8888 gnd.n708 gnd.n707 585
R8889 gnd.n6362 gnd.n6361 585
R8890 gnd.n6361 gnd.n6360 585
R8891 gnd.n714 gnd.n713 585
R8892 gnd.n6359 gnd.n714 585
R8893 gnd.n6357 gnd.n6356 585
R8894 gnd.n6358 gnd.n6357 585
R8895 gnd.n6355 gnd.n716 585
R8896 gnd.n716 gnd.n715 585
R8897 gnd.n6354 gnd.n6353 585
R8898 gnd.n6353 gnd.n6352 585
R8899 gnd.n722 gnd.n721 585
R8900 gnd.n6351 gnd.n722 585
R8901 gnd.n6349 gnd.n6348 585
R8902 gnd.n6350 gnd.n6349 585
R8903 gnd.n6347 gnd.n724 585
R8904 gnd.n724 gnd.n723 585
R8905 gnd.n6346 gnd.n6345 585
R8906 gnd.n6345 gnd.n6344 585
R8907 gnd.n730 gnd.n729 585
R8908 gnd.n6343 gnd.n730 585
R8909 gnd.n6341 gnd.n6340 585
R8910 gnd.n6342 gnd.n6341 585
R8911 gnd.n6339 gnd.n732 585
R8912 gnd.n732 gnd.n731 585
R8913 gnd.n6338 gnd.n6337 585
R8914 gnd.n6337 gnd.n6336 585
R8915 gnd.n738 gnd.n737 585
R8916 gnd.n6335 gnd.n738 585
R8917 gnd.n6333 gnd.n6332 585
R8918 gnd.n6334 gnd.n6333 585
R8919 gnd.n6331 gnd.n740 585
R8920 gnd.n740 gnd.n739 585
R8921 gnd.n6330 gnd.n6329 585
R8922 gnd.n6329 gnd.n6328 585
R8923 gnd.n746 gnd.n745 585
R8924 gnd.n6327 gnd.n746 585
R8925 gnd.n6325 gnd.n6324 585
R8926 gnd.n6326 gnd.n6325 585
R8927 gnd.n6323 gnd.n748 585
R8928 gnd.n748 gnd.n747 585
R8929 gnd.n6322 gnd.n6321 585
R8930 gnd.n6321 gnd.n6320 585
R8931 gnd.n754 gnd.n753 585
R8932 gnd.n6319 gnd.n754 585
R8933 gnd.n6317 gnd.n6316 585
R8934 gnd.n6318 gnd.n6317 585
R8935 gnd.n6315 gnd.n756 585
R8936 gnd.n756 gnd.n755 585
R8937 gnd.n6314 gnd.n6313 585
R8938 gnd.n6313 gnd.n6312 585
R8939 gnd.n762 gnd.n761 585
R8940 gnd.n6311 gnd.n762 585
R8941 gnd.n6309 gnd.n6308 585
R8942 gnd.n6310 gnd.n6309 585
R8943 gnd.n6307 gnd.n764 585
R8944 gnd.n764 gnd.n763 585
R8945 gnd.n6306 gnd.n6305 585
R8946 gnd.n6305 gnd.n6304 585
R8947 gnd.n770 gnd.n769 585
R8948 gnd.n6303 gnd.n770 585
R8949 gnd.n6301 gnd.n6300 585
R8950 gnd.n6302 gnd.n6301 585
R8951 gnd.n6299 gnd.n772 585
R8952 gnd.n772 gnd.n771 585
R8953 gnd.n6298 gnd.n6297 585
R8954 gnd.n6297 gnd.n6296 585
R8955 gnd.n778 gnd.n777 585
R8956 gnd.n6295 gnd.n778 585
R8957 gnd.n6293 gnd.n6292 585
R8958 gnd.n6294 gnd.n6293 585
R8959 gnd.n6291 gnd.n780 585
R8960 gnd.n780 gnd.n779 585
R8961 gnd.n6290 gnd.n6289 585
R8962 gnd.n6289 gnd.n6288 585
R8963 gnd.n786 gnd.n785 585
R8964 gnd.n6287 gnd.n786 585
R8965 gnd.n6285 gnd.n6284 585
R8966 gnd.n6286 gnd.n6285 585
R8967 gnd.n6283 gnd.n788 585
R8968 gnd.n788 gnd.n787 585
R8969 gnd.n6282 gnd.n6281 585
R8970 gnd.n6281 gnd.n6280 585
R8971 gnd.n794 gnd.n793 585
R8972 gnd.n6279 gnd.n794 585
R8973 gnd.n6277 gnd.n6276 585
R8974 gnd.n6278 gnd.n6277 585
R8975 gnd.n6275 gnd.n796 585
R8976 gnd.n796 gnd.n795 585
R8977 gnd.n6274 gnd.n6273 585
R8978 gnd.n6273 gnd.n6272 585
R8979 gnd.n802 gnd.n801 585
R8980 gnd.n6271 gnd.n802 585
R8981 gnd.n6269 gnd.n6268 585
R8982 gnd.n6270 gnd.n6269 585
R8983 gnd.n6267 gnd.n804 585
R8984 gnd.n804 gnd.n803 585
R8985 gnd.n6266 gnd.n6265 585
R8986 gnd.n6265 gnd.n6264 585
R8987 gnd.n810 gnd.n809 585
R8988 gnd.n6263 gnd.n810 585
R8989 gnd.n6261 gnd.n6260 585
R8990 gnd.n6262 gnd.n6261 585
R8991 gnd.n6259 gnd.n812 585
R8992 gnd.n812 gnd.n811 585
R8993 gnd.n6258 gnd.n6257 585
R8994 gnd.n6257 gnd.n6256 585
R8995 gnd.n818 gnd.n817 585
R8996 gnd.n6255 gnd.n818 585
R8997 gnd.n6253 gnd.n6252 585
R8998 gnd.n6254 gnd.n6253 585
R8999 gnd.n6251 gnd.n820 585
R9000 gnd.n820 gnd.n819 585
R9001 gnd.n6250 gnd.n6249 585
R9002 gnd.n6249 gnd.n6248 585
R9003 gnd.n826 gnd.n825 585
R9004 gnd.n6247 gnd.n826 585
R9005 gnd.n6245 gnd.n6244 585
R9006 gnd.n6246 gnd.n6245 585
R9007 gnd.n6243 gnd.n828 585
R9008 gnd.n828 gnd.n827 585
R9009 gnd.n6242 gnd.n6241 585
R9010 gnd.n6241 gnd.n6240 585
R9011 gnd.n834 gnd.n833 585
R9012 gnd.n6239 gnd.n834 585
R9013 gnd.n6237 gnd.n6236 585
R9014 gnd.n6238 gnd.n6237 585
R9015 gnd.n6235 gnd.n836 585
R9016 gnd.n836 gnd.n835 585
R9017 gnd.n672 gnd.n671 585
R9018 gnd.n671 gnd.n670 585
R9019 gnd.n6407 gnd.n6406 585
R9020 gnd.n6408 gnd.n6407 585
R9021 gnd.n669 gnd.n668 585
R9022 gnd.n6409 gnd.n669 585
R9023 gnd.n6412 gnd.n6411 585
R9024 gnd.n6411 gnd.n6410 585
R9025 gnd.n666 gnd.n665 585
R9026 gnd.n665 gnd.n664 585
R9027 gnd.n6417 gnd.n6416 585
R9028 gnd.n6418 gnd.n6417 585
R9029 gnd.n663 gnd.n662 585
R9030 gnd.n6419 gnd.n663 585
R9031 gnd.n6422 gnd.n6421 585
R9032 gnd.n6421 gnd.n6420 585
R9033 gnd.n660 gnd.n659 585
R9034 gnd.n659 gnd.n658 585
R9035 gnd.n6427 gnd.n6426 585
R9036 gnd.n6428 gnd.n6427 585
R9037 gnd.n657 gnd.n656 585
R9038 gnd.n6429 gnd.n657 585
R9039 gnd.n6432 gnd.n6431 585
R9040 gnd.n6431 gnd.n6430 585
R9041 gnd.n654 gnd.n653 585
R9042 gnd.n653 gnd.n652 585
R9043 gnd.n6437 gnd.n6436 585
R9044 gnd.n6438 gnd.n6437 585
R9045 gnd.n651 gnd.n650 585
R9046 gnd.n6439 gnd.n651 585
R9047 gnd.n6442 gnd.n6441 585
R9048 gnd.n6441 gnd.n6440 585
R9049 gnd.n648 gnd.n647 585
R9050 gnd.n647 gnd.n646 585
R9051 gnd.n6447 gnd.n6446 585
R9052 gnd.n6448 gnd.n6447 585
R9053 gnd.n645 gnd.n644 585
R9054 gnd.n6449 gnd.n645 585
R9055 gnd.n6452 gnd.n6451 585
R9056 gnd.n6451 gnd.n6450 585
R9057 gnd.n642 gnd.n641 585
R9058 gnd.n641 gnd.n640 585
R9059 gnd.n6457 gnd.n6456 585
R9060 gnd.n6458 gnd.n6457 585
R9061 gnd.n639 gnd.n638 585
R9062 gnd.n6459 gnd.n639 585
R9063 gnd.n6462 gnd.n6461 585
R9064 gnd.n6461 gnd.n6460 585
R9065 gnd.n636 gnd.n635 585
R9066 gnd.n635 gnd.n634 585
R9067 gnd.n6467 gnd.n6466 585
R9068 gnd.n6468 gnd.n6467 585
R9069 gnd.n633 gnd.n632 585
R9070 gnd.n6469 gnd.n633 585
R9071 gnd.n6472 gnd.n6471 585
R9072 gnd.n6471 gnd.n6470 585
R9073 gnd.n630 gnd.n629 585
R9074 gnd.n629 gnd.n628 585
R9075 gnd.n6477 gnd.n6476 585
R9076 gnd.n6478 gnd.n6477 585
R9077 gnd.n627 gnd.n626 585
R9078 gnd.n6479 gnd.n627 585
R9079 gnd.n6482 gnd.n6481 585
R9080 gnd.n6481 gnd.n6480 585
R9081 gnd.n624 gnd.n623 585
R9082 gnd.n623 gnd.n622 585
R9083 gnd.n6487 gnd.n6486 585
R9084 gnd.n6488 gnd.n6487 585
R9085 gnd.n621 gnd.n620 585
R9086 gnd.n6489 gnd.n621 585
R9087 gnd.n6492 gnd.n6491 585
R9088 gnd.n6491 gnd.n6490 585
R9089 gnd.n618 gnd.n617 585
R9090 gnd.n617 gnd.n616 585
R9091 gnd.n6497 gnd.n6496 585
R9092 gnd.n6498 gnd.n6497 585
R9093 gnd.n615 gnd.n614 585
R9094 gnd.n6499 gnd.n615 585
R9095 gnd.n6502 gnd.n6501 585
R9096 gnd.n6501 gnd.n6500 585
R9097 gnd.n612 gnd.n611 585
R9098 gnd.n611 gnd.n610 585
R9099 gnd.n6507 gnd.n6506 585
R9100 gnd.n6508 gnd.n6507 585
R9101 gnd.n609 gnd.n608 585
R9102 gnd.n6509 gnd.n609 585
R9103 gnd.n6512 gnd.n6511 585
R9104 gnd.n6511 gnd.n6510 585
R9105 gnd.n606 gnd.n605 585
R9106 gnd.n605 gnd.n604 585
R9107 gnd.n6517 gnd.n6516 585
R9108 gnd.n6518 gnd.n6517 585
R9109 gnd.n603 gnd.n602 585
R9110 gnd.n6519 gnd.n603 585
R9111 gnd.n6522 gnd.n6521 585
R9112 gnd.n6521 gnd.n6520 585
R9113 gnd.n600 gnd.n599 585
R9114 gnd.n599 gnd.n598 585
R9115 gnd.n6527 gnd.n6526 585
R9116 gnd.n6528 gnd.n6527 585
R9117 gnd.n597 gnd.n596 585
R9118 gnd.n6529 gnd.n597 585
R9119 gnd.n6532 gnd.n6531 585
R9120 gnd.n6531 gnd.n6530 585
R9121 gnd.n594 gnd.n593 585
R9122 gnd.n593 gnd.n592 585
R9123 gnd.n6537 gnd.n6536 585
R9124 gnd.n6538 gnd.n6537 585
R9125 gnd.n591 gnd.n590 585
R9126 gnd.n6539 gnd.n591 585
R9127 gnd.n6542 gnd.n6541 585
R9128 gnd.n6541 gnd.n6540 585
R9129 gnd.n588 gnd.n587 585
R9130 gnd.n587 gnd.n586 585
R9131 gnd.n6547 gnd.n6546 585
R9132 gnd.n6548 gnd.n6547 585
R9133 gnd.n585 gnd.n584 585
R9134 gnd.n6549 gnd.n585 585
R9135 gnd.n6552 gnd.n6551 585
R9136 gnd.n6551 gnd.n6550 585
R9137 gnd.n582 gnd.n581 585
R9138 gnd.n581 gnd.n580 585
R9139 gnd.n6557 gnd.n6556 585
R9140 gnd.n6558 gnd.n6557 585
R9141 gnd.n579 gnd.n578 585
R9142 gnd.n6559 gnd.n579 585
R9143 gnd.n6562 gnd.n6561 585
R9144 gnd.n6561 gnd.n6560 585
R9145 gnd.n576 gnd.n575 585
R9146 gnd.n575 gnd.n574 585
R9147 gnd.n6567 gnd.n6566 585
R9148 gnd.n6568 gnd.n6567 585
R9149 gnd.n573 gnd.n572 585
R9150 gnd.n6569 gnd.n573 585
R9151 gnd.n6572 gnd.n6571 585
R9152 gnd.n6571 gnd.n6570 585
R9153 gnd.n570 gnd.n569 585
R9154 gnd.n569 gnd.n568 585
R9155 gnd.n6577 gnd.n6576 585
R9156 gnd.n6578 gnd.n6577 585
R9157 gnd.n567 gnd.n566 585
R9158 gnd.n6579 gnd.n567 585
R9159 gnd.n6582 gnd.n6581 585
R9160 gnd.n6581 gnd.n6580 585
R9161 gnd.n564 gnd.n563 585
R9162 gnd.n563 gnd.n562 585
R9163 gnd.n6587 gnd.n6586 585
R9164 gnd.n6588 gnd.n6587 585
R9165 gnd.n561 gnd.n560 585
R9166 gnd.n6589 gnd.n561 585
R9167 gnd.n6592 gnd.n6591 585
R9168 gnd.n6591 gnd.n6590 585
R9169 gnd.n558 gnd.n557 585
R9170 gnd.n557 gnd.n556 585
R9171 gnd.n6597 gnd.n6596 585
R9172 gnd.n6598 gnd.n6597 585
R9173 gnd.n555 gnd.n554 585
R9174 gnd.n6599 gnd.n555 585
R9175 gnd.n6602 gnd.n6601 585
R9176 gnd.n6601 gnd.n6600 585
R9177 gnd.n552 gnd.n551 585
R9178 gnd.n551 gnd.n550 585
R9179 gnd.n6607 gnd.n6606 585
R9180 gnd.n6608 gnd.n6607 585
R9181 gnd.n549 gnd.n548 585
R9182 gnd.n6609 gnd.n549 585
R9183 gnd.n6612 gnd.n6611 585
R9184 gnd.n6611 gnd.n6610 585
R9185 gnd.n546 gnd.n545 585
R9186 gnd.n545 gnd.n544 585
R9187 gnd.n6617 gnd.n6616 585
R9188 gnd.n6618 gnd.n6617 585
R9189 gnd.n543 gnd.n542 585
R9190 gnd.n6619 gnd.n543 585
R9191 gnd.n6622 gnd.n6621 585
R9192 gnd.n6621 gnd.n6620 585
R9193 gnd.n540 gnd.n539 585
R9194 gnd.n539 gnd.n538 585
R9195 gnd.n6627 gnd.n6626 585
R9196 gnd.n6628 gnd.n6627 585
R9197 gnd.n537 gnd.n536 585
R9198 gnd.n6629 gnd.n537 585
R9199 gnd.n6632 gnd.n6631 585
R9200 gnd.n6631 gnd.n6630 585
R9201 gnd.n534 gnd.n533 585
R9202 gnd.n533 gnd.n532 585
R9203 gnd.n6637 gnd.n6636 585
R9204 gnd.n6638 gnd.n6637 585
R9205 gnd.n531 gnd.n530 585
R9206 gnd.n6639 gnd.n531 585
R9207 gnd.n6642 gnd.n6641 585
R9208 gnd.n6641 gnd.n6640 585
R9209 gnd.n528 gnd.n527 585
R9210 gnd.n527 gnd.n526 585
R9211 gnd.n6647 gnd.n6646 585
R9212 gnd.n6648 gnd.n6647 585
R9213 gnd.n525 gnd.n524 585
R9214 gnd.n6649 gnd.n525 585
R9215 gnd.n6652 gnd.n6651 585
R9216 gnd.n6651 gnd.n6650 585
R9217 gnd.n522 gnd.n521 585
R9218 gnd.n521 gnd.n520 585
R9219 gnd.n6657 gnd.n6656 585
R9220 gnd.n6658 gnd.n6657 585
R9221 gnd.n519 gnd.n518 585
R9222 gnd.n6659 gnd.n519 585
R9223 gnd.n6662 gnd.n6661 585
R9224 gnd.n6661 gnd.n6660 585
R9225 gnd.n516 gnd.n515 585
R9226 gnd.n515 gnd.n514 585
R9227 gnd.n6667 gnd.n6666 585
R9228 gnd.n6668 gnd.n6667 585
R9229 gnd.n513 gnd.n512 585
R9230 gnd.n6669 gnd.n513 585
R9231 gnd.n6672 gnd.n6671 585
R9232 gnd.n6671 gnd.n6670 585
R9233 gnd.n510 gnd.n509 585
R9234 gnd.n509 gnd.n508 585
R9235 gnd.n6677 gnd.n6676 585
R9236 gnd.n6678 gnd.n6677 585
R9237 gnd.n507 gnd.n506 585
R9238 gnd.n6679 gnd.n507 585
R9239 gnd.n6682 gnd.n6681 585
R9240 gnd.n6681 gnd.n6680 585
R9241 gnd.n504 gnd.n503 585
R9242 gnd.n503 gnd.n502 585
R9243 gnd.n6687 gnd.n6686 585
R9244 gnd.n6688 gnd.n6687 585
R9245 gnd.n501 gnd.n500 585
R9246 gnd.n6689 gnd.n501 585
R9247 gnd.n6692 gnd.n6691 585
R9248 gnd.n6691 gnd.n6690 585
R9249 gnd.n498 gnd.n497 585
R9250 gnd.n497 gnd.n496 585
R9251 gnd.n6697 gnd.n6696 585
R9252 gnd.n6698 gnd.n6697 585
R9253 gnd.n495 gnd.n494 585
R9254 gnd.n6699 gnd.n495 585
R9255 gnd.n6702 gnd.n6701 585
R9256 gnd.n6701 gnd.n6700 585
R9257 gnd.n492 gnd.n491 585
R9258 gnd.n491 gnd.n490 585
R9259 gnd.n6707 gnd.n6706 585
R9260 gnd.n6708 gnd.n6707 585
R9261 gnd.n489 gnd.n488 585
R9262 gnd.n6709 gnd.n489 585
R9263 gnd.n6712 gnd.n6711 585
R9264 gnd.n6711 gnd.n6710 585
R9265 gnd.n486 gnd.n485 585
R9266 gnd.n485 gnd.n484 585
R9267 gnd.n6717 gnd.n6716 585
R9268 gnd.n6718 gnd.n6717 585
R9269 gnd.n483 gnd.n482 585
R9270 gnd.n6719 gnd.n483 585
R9271 gnd.n6722 gnd.n6721 585
R9272 gnd.n6721 gnd.n6720 585
R9273 gnd.n480 gnd.n479 585
R9274 gnd.n479 gnd.n478 585
R9275 gnd.n6727 gnd.n6726 585
R9276 gnd.n6728 gnd.n6727 585
R9277 gnd.n477 gnd.n476 585
R9278 gnd.n6729 gnd.n477 585
R9279 gnd.n6732 gnd.n6731 585
R9280 gnd.n6731 gnd.n6730 585
R9281 gnd.n474 gnd.n473 585
R9282 gnd.n473 gnd.n472 585
R9283 gnd.n6737 gnd.n6736 585
R9284 gnd.n6738 gnd.n6737 585
R9285 gnd.n471 gnd.n470 585
R9286 gnd.n6739 gnd.n471 585
R9287 gnd.n6742 gnd.n6741 585
R9288 gnd.n6741 gnd.n6740 585
R9289 gnd.n468 gnd.n467 585
R9290 gnd.n467 gnd.n466 585
R9291 gnd.n6747 gnd.n6746 585
R9292 gnd.n6748 gnd.n6747 585
R9293 gnd.n465 gnd.n464 585
R9294 gnd.n6749 gnd.n465 585
R9295 gnd.n6752 gnd.n6751 585
R9296 gnd.n6751 gnd.n6750 585
R9297 gnd.n462 gnd.n461 585
R9298 gnd.n461 gnd.n460 585
R9299 gnd.n6757 gnd.n6756 585
R9300 gnd.n6758 gnd.n6757 585
R9301 gnd.n459 gnd.n458 585
R9302 gnd.n6759 gnd.n459 585
R9303 gnd.n6762 gnd.n6761 585
R9304 gnd.n6761 gnd.n6760 585
R9305 gnd.n456 gnd.n455 585
R9306 gnd.n455 gnd.n454 585
R9307 gnd.n6767 gnd.n6766 585
R9308 gnd.n6768 gnd.n6767 585
R9309 gnd.n453 gnd.n452 585
R9310 gnd.n6769 gnd.n453 585
R9311 gnd.n6772 gnd.n6771 585
R9312 gnd.n6771 gnd.n6770 585
R9313 gnd.n450 gnd.n449 585
R9314 gnd.n449 gnd.n448 585
R9315 gnd.n6777 gnd.n6776 585
R9316 gnd.n6778 gnd.n6777 585
R9317 gnd.n447 gnd.n446 585
R9318 gnd.n6779 gnd.n447 585
R9319 gnd.n6782 gnd.n6781 585
R9320 gnd.n6781 gnd.n6780 585
R9321 gnd.n444 gnd.n443 585
R9322 gnd.n443 gnd.n442 585
R9323 gnd.n6787 gnd.n6786 585
R9324 gnd.n6788 gnd.n6787 585
R9325 gnd.n441 gnd.n440 585
R9326 gnd.n6789 gnd.n441 585
R9327 gnd.n6792 gnd.n6791 585
R9328 gnd.n6791 gnd.n6790 585
R9329 gnd.n438 gnd.n437 585
R9330 gnd.n437 gnd.n436 585
R9331 gnd.n6797 gnd.n6796 585
R9332 gnd.n6798 gnd.n6797 585
R9333 gnd.n435 gnd.n434 585
R9334 gnd.n6799 gnd.n435 585
R9335 gnd.n6802 gnd.n6801 585
R9336 gnd.n6801 gnd.n6800 585
R9337 gnd.n432 gnd.n431 585
R9338 gnd.n431 gnd.n430 585
R9339 gnd.n6807 gnd.n6806 585
R9340 gnd.n6808 gnd.n6807 585
R9341 gnd.n429 gnd.n428 585
R9342 gnd.n6809 gnd.n429 585
R9343 gnd.n6812 gnd.n6811 585
R9344 gnd.n6811 gnd.n6810 585
R9345 gnd.n426 gnd.n425 585
R9346 gnd.n425 gnd.n424 585
R9347 gnd.n6817 gnd.n6816 585
R9348 gnd.n6818 gnd.n6817 585
R9349 gnd.n423 gnd.n422 585
R9350 gnd.n6819 gnd.n423 585
R9351 gnd.n6822 gnd.n6821 585
R9352 gnd.n6821 gnd.n6820 585
R9353 gnd.n420 gnd.n419 585
R9354 gnd.n419 gnd.n418 585
R9355 gnd.n6827 gnd.n6826 585
R9356 gnd.n6828 gnd.n6827 585
R9357 gnd.n417 gnd.n416 585
R9358 gnd.n6829 gnd.n417 585
R9359 gnd.n6832 gnd.n6831 585
R9360 gnd.n6831 gnd.n6830 585
R9361 gnd.n414 gnd.n413 585
R9362 gnd.n413 gnd.n412 585
R9363 gnd.n6837 gnd.n6836 585
R9364 gnd.n6838 gnd.n6837 585
R9365 gnd.n411 gnd.n410 585
R9366 gnd.n6839 gnd.n411 585
R9367 gnd.n6842 gnd.n6841 585
R9368 gnd.n6841 gnd.n6840 585
R9369 gnd.n408 gnd.n407 585
R9370 gnd.n407 gnd.n406 585
R9371 gnd.n6847 gnd.n6846 585
R9372 gnd.n6848 gnd.n6847 585
R9373 gnd.n405 gnd.n404 585
R9374 gnd.n6849 gnd.n405 585
R9375 gnd.n6852 gnd.n6851 585
R9376 gnd.n6851 gnd.n6850 585
R9377 gnd.n402 gnd.n401 585
R9378 gnd.n401 gnd.n400 585
R9379 gnd.n6857 gnd.n6856 585
R9380 gnd.n6858 gnd.n6857 585
R9381 gnd.n399 gnd.n398 585
R9382 gnd.n6859 gnd.n399 585
R9383 gnd.n6862 gnd.n6861 585
R9384 gnd.n6861 gnd.n6860 585
R9385 gnd.n396 gnd.n395 585
R9386 gnd.n395 gnd.n394 585
R9387 gnd.n6867 gnd.n6866 585
R9388 gnd.n6868 gnd.n6867 585
R9389 gnd.n393 gnd.n392 585
R9390 gnd.n6869 gnd.n393 585
R9391 gnd.n6872 gnd.n6871 585
R9392 gnd.n6871 gnd.n6870 585
R9393 gnd.n390 gnd.n389 585
R9394 gnd.n389 gnd.n388 585
R9395 gnd.n6877 gnd.n6876 585
R9396 gnd.n6878 gnd.n6877 585
R9397 gnd.n387 gnd.n386 585
R9398 gnd.n6879 gnd.n387 585
R9399 gnd.n6882 gnd.n6881 585
R9400 gnd.n6881 gnd.n6880 585
R9401 gnd.n384 gnd.n383 585
R9402 gnd.n383 gnd.n382 585
R9403 gnd.n6888 gnd.n6887 585
R9404 gnd.n6889 gnd.n6888 585
R9405 gnd.n6886 gnd.n381 585
R9406 gnd.n6890 gnd.n381 585
R9407 gnd.n256 gnd.n255 585
R9408 gnd.n7100 gnd.n256 585
R9409 gnd.n7098 gnd.n7097 585
R9410 gnd.n7099 gnd.n7098 585
R9411 gnd.n259 gnd.n258 585
R9412 gnd.n258 gnd.n257 585
R9413 gnd.n7093 gnd.n7092 585
R9414 gnd.n7092 gnd.n7091 585
R9415 gnd.n262 gnd.n261 585
R9416 gnd.n7090 gnd.n262 585
R9417 gnd.n7088 gnd.n7087 585
R9418 gnd.n7089 gnd.n7088 585
R9419 gnd.n265 gnd.n264 585
R9420 gnd.n264 gnd.n263 585
R9421 gnd.n7083 gnd.n7082 585
R9422 gnd.n7082 gnd.n7081 585
R9423 gnd.n268 gnd.n267 585
R9424 gnd.n7080 gnd.n268 585
R9425 gnd.n7078 gnd.n7077 585
R9426 gnd.n7079 gnd.n7078 585
R9427 gnd.n271 gnd.n270 585
R9428 gnd.n270 gnd.n269 585
R9429 gnd.n7073 gnd.n7072 585
R9430 gnd.n7072 gnd.n7071 585
R9431 gnd.n274 gnd.n273 585
R9432 gnd.n7070 gnd.n274 585
R9433 gnd.n7068 gnd.n7067 585
R9434 gnd.n7069 gnd.n7068 585
R9435 gnd.n277 gnd.n276 585
R9436 gnd.n276 gnd.n275 585
R9437 gnd.n7063 gnd.n7062 585
R9438 gnd.n7062 gnd.n7061 585
R9439 gnd.n280 gnd.n279 585
R9440 gnd.n7060 gnd.n280 585
R9441 gnd.n7058 gnd.n7057 585
R9442 gnd.n7059 gnd.n7058 585
R9443 gnd.n283 gnd.n282 585
R9444 gnd.n282 gnd.n281 585
R9445 gnd.n7053 gnd.n7052 585
R9446 gnd.n7052 gnd.n7051 585
R9447 gnd.n286 gnd.n285 585
R9448 gnd.n7050 gnd.n286 585
R9449 gnd.n7048 gnd.n7047 585
R9450 gnd.n7049 gnd.n7048 585
R9451 gnd.n289 gnd.n288 585
R9452 gnd.n288 gnd.n287 585
R9453 gnd.n7043 gnd.n7042 585
R9454 gnd.n7042 gnd.n7041 585
R9455 gnd.n292 gnd.n291 585
R9456 gnd.n7040 gnd.n292 585
R9457 gnd.n7038 gnd.n7037 585
R9458 gnd.n7039 gnd.n7038 585
R9459 gnd.n295 gnd.n294 585
R9460 gnd.n294 gnd.n293 585
R9461 gnd.n7033 gnd.n7032 585
R9462 gnd.n7032 gnd.n7031 585
R9463 gnd.n298 gnd.n297 585
R9464 gnd.n7030 gnd.n298 585
R9465 gnd.n7028 gnd.n7027 585
R9466 gnd.n7029 gnd.n7028 585
R9467 gnd.n301 gnd.n300 585
R9468 gnd.n300 gnd.n299 585
R9469 gnd.n7023 gnd.n7022 585
R9470 gnd.n7022 gnd.n7021 585
R9471 gnd.n304 gnd.n303 585
R9472 gnd.n7020 gnd.n304 585
R9473 gnd.n7018 gnd.n7017 585
R9474 gnd.n7019 gnd.n7018 585
R9475 gnd.n307 gnd.n306 585
R9476 gnd.n306 gnd.n305 585
R9477 gnd.n7013 gnd.n7012 585
R9478 gnd.n7012 gnd.n7011 585
R9479 gnd.n310 gnd.n309 585
R9480 gnd.n7010 gnd.n310 585
R9481 gnd.n7008 gnd.n7007 585
R9482 gnd.n7009 gnd.n7008 585
R9483 gnd.n313 gnd.n312 585
R9484 gnd.n312 gnd.n311 585
R9485 gnd.n7003 gnd.n7002 585
R9486 gnd.n7002 gnd.n7001 585
R9487 gnd.n316 gnd.n315 585
R9488 gnd.n7000 gnd.n316 585
R9489 gnd.n6998 gnd.n6997 585
R9490 gnd.n6999 gnd.n6998 585
R9491 gnd.n319 gnd.n318 585
R9492 gnd.n318 gnd.n317 585
R9493 gnd.n6993 gnd.n6992 585
R9494 gnd.n6992 gnd.n6991 585
R9495 gnd.n322 gnd.n321 585
R9496 gnd.n6990 gnd.n322 585
R9497 gnd.n6988 gnd.n6987 585
R9498 gnd.n6989 gnd.n6988 585
R9499 gnd.n325 gnd.n324 585
R9500 gnd.n324 gnd.n323 585
R9501 gnd.n6983 gnd.n6982 585
R9502 gnd.n6982 gnd.n6981 585
R9503 gnd.n328 gnd.n327 585
R9504 gnd.n6980 gnd.n328 585
R9505 gnd.n6978 gnd.n6977 585
R9506 gnd.n6979 gnd.n6978 585
R9507 gnd.n331 gnd.n330 585
R9508 gnd.n330 gnd.n329 585
R9509 gnd.n6973 gnd.n6972 585
R9510 gnd.n6972 gnd.n6971 585
R9511 gnd.n334 gnd.n333 585
R9512 gnd.n6970 gnd.n334 585
R9513 gnd.n6968 gnd.n6967 585
R9514 gnd.n6969 gnd.n6968 585
R9515 gnd.n337 gnd.n336 585
R9516 gnd.n336 gnd.n335 585
R9517 gnd.n6963 gnd.n6962 585
R9518 gnd.n6962 gnd.n6961 585
R9519 gnd.n340 gnd.n339 585
R9520 gnd.n6960 gnd.n340 585
R9521 gnd.n6958 gnd.n6957 585
R9522 gnd.n6959 gnd.n6958 585
R9523 gnd.n343 gnd.n342 585
R9524 gnd.n342 gnd.n341 585
R9525 gnd.n6953 gnd.n6952 585
R9526 gnd.n6952 gnd.n6951 585
R9527 gnd.n346 gnd.n345 585
R9528 gnd.n6950 gnd.n346 585
R9529 gnd.n6948 gnd.n6947 585
R9530 gnd.n6949 gnd.n6948 585
R9531 gnd.n349 gnd.n348 585
R9532 gnd.n348 gnd.n347 585
R9533 gnd.n6943 gnd.n6942 585
R9534 gnd.n6942 gnd.n6941 585
R9535 gnd.n352 gnd.n351 585
R9536 gnd.n6940 gnd.n352 585
R9537 gnd.n6938 gnd.n6937 585
R9538 gnd.n6939 gnd.n6938 585
R9539 gnd.n355 gnd.n354 585
R9540 gnd.n354 gnd.n353 585
R9541 gnd.n6933 gnd.n6932 585
R9542 gnd.n6932 gnd.n6931 585
R9543 gnd.n358 gnd.n357 585
R9544 gnd.n6930 gnd.n358 585
R9545 gnd.n6928 gnd.n6927 585
R9546 gnd.n6929 gnd.n6928 585
R9547 gnd.n361 gnd.n360 585
R9548 gnd.n360 gnd.n359 585
R9549 gnd.n6923 gnd.n6922 585
R9550 gnd.n6922 gnd.n6921 585
R9551 gnd.n364 gnd.n363 585
R9552 gnd.n6920 gnd.n364 585
R9553 gnd.n6918 gnd.n6917 585
R9554 gnd.n6919 gnd.n6918 585
R9555 gnd.n367 gnd.n366 585
R9556 gnd.n366 gnd.n365 585
R9557 gnd.n6913 gnd.n6912 585
R9558 gnd.n6912 gnd.n6911 585
R9559 gnd.n370 gnd.n369 585
R9560 gnd.n6910 gnd.n370 585
R9561 gnd.n6908 gnd.n6907 585
R9562 gnd.n6909 gnd.n6908 585
R9563 gnd.n373 gnd.n372 585
R9564 gnd.n372 gnd.n371 585
R9565 gnd.n6903 gnd.n6902 585
R9566 gnd.n6902 gnd.n6901 585
R9567 gnd.n376 gnd.n375 585
R9568 gnd.n6900 gnd.n376 585
R9569 gnd.n6898 gnd.n6897 585
R9570 gnd.n6899 gnd.n6898 585
R9571 gnd.n379 gnd.n378 585
R9572 gnd.n378 gnd.n377 585
R9573 gnd.n6893 gnd.n6892 585
R9574 gnd.n6892 gnd.n6891 585
R9575 gnd.n6085 gnd.n6084 585
R9576 gnd.n6086 gnd.n6085 585
R9577 gnd.n2522 gnd.n2521 585
R9578 gnd.n6079 gnd.n2522 585
R9579 gnd.n6094 gnd.n6093 585
R9580 gnd.n6093 gnd.n6092 585
R9581 gnd.n6095 gnd.n2517 585
R9582 gnd.n4228 gnd.n2517 585
R9583 gnd.n6097 gnd.n6096 585
R9584 gnd.n6098 gnd.n6097 585
R9585 gnd.n2501 gnd.n2500 585
R9586 gnd.n4222 gnd.n2501 585
R9587 gnd.n6106 gnd.n6105 585
R9588 gnd.n6105 gnd.n6104 585
R9589 gnd.n6107 gnd.n2496 585
R9590 gnd.n4217 gnd.n2496 585
R9591 gnd.n6109 gnd.n6108 585
R9592 gnd.n6110 gnd.n6109 585
R9593 gnd.n2480 gnd.n2479 585
R9594 gnd.n4213 gnd.n2480 585
R9595 gnd.n6118 gnd.n6117 585
R9596 gnd.n6117 gnd.n6116 585
R9597 gnd.n6119 gnd.n2475 585
R9598 gnd.n4245 gnd.n2475 585
R9599 gnd.n6121 gnd.n6120 585
R9600 gnd.n6122 gnd.n6121 585
R9601 gnd.n2460 gnd.n2459 585
R9602 gnd.n4206 gnd.n2460 585
R9603 gnd.n6130 gnd.n6129 585
R9604 gnd.n6129 gnd.n6128 585
R9605 gnd.n6131 gnd.n2455 585
R9606 gnd.n4198 gnd.n2455 585
R9607 gnd.n6133 gnd.n6132 585
R9608 gnd.n6134 gnd.n6133 585
R9609 gnd.n2442 gnd.n2441 585
R9610 gnd.n4192 gnd.n2442 585
R9611 gnd.n6143 gnd.n6142 585
R9612 gnd.n6142 gnd.n6141 585
R9613 gnd.n6144 gnd.n2437 585
R9614 gnd.n4184 gnd.n2437 585
R9615 gnd.n6146 gnd.n6145 585
R9616 gnd.n6147 gnd.n6146 585
R9617 gnd.n2425 gnd.n2424 585
R9618 gnd.n4178 gnd.n2425 585
R9619 gnd.n6156 gnd.n6155 585
R9620 gnd.n6155 gnd.n6154 585
R9621 gnd.n6157 gnd.n2420 585
R9622 gnd.n4170 gnd.n2420 585
R9623 gnd.n6159 gnd.n6158 585
R9624 gnd.n6160 gnd.n6159 585
R9625 gnd.n2406 gnd.n2405 585
R9626 gnd.n4164 gnd.n2406 585
R9627 gnd.n6169 gnd.n6168 585
R9628 gnd.n6168 gnd.n6167 585
R9629 gnd.n6170 gnd.n2401 585
R9630 gnd.n4156 gnd.n2401 585
R9631 gnd.n6172 gnd.n6171 585
R9632 gnd.n6173 gnd.n6172 585
R9633 gnd.n2386 gnd.n2385 585
R9634 gnd.n4150 gnd.n2386 585
R9635 gnd.n6181 gnd.n6180 585
R9636 gnd.n6180 gnd.n6179 585
R9637 gnd.n6182 gnd.n2381 585
R9638 gnd.n4142 gnd.n2381 585
R9639 gnd.n6184 gnd.n6183 585
R9640 gnd.n6185 gnd.n6184 585
R9641 gnd.n2365 gnd.n2364 585
R9642 gnd.n4136 gnd.n2365 585
R9643 gnd.n6193 gnd.n6192 585
R9644 gnd.n6192 gnd.n6191 585
R9645 gnd.n6194 gnd.n2360 585
R9646 gnd.n4128 gnd.n2360 585
R9647 gnd.n6196 gnd.n6195 585
R9648 gnd.n6197 gnd.n6196 585
R9649 gnd.n2345 gnd.n2344 585
R9650 gnd.n4122 gnd.n2345 585
R9651 gnd.n6205 gnd.n6204 585
R9652 gnd.n6204 gnd.n6203 585
R9653 gnd.n6206 gnd.n2339 585
R9654 gnd.n4114 gnd.n2339 585
R9655 gnd.n6208 gnd.n6207 585
R9656 gnd.n6209 gnd.n6208 585
R9657 gnd.n2340 gnd.n2338 585
R9658 gnd.n3848 gnd.n2338 585
R9659 gnd.n4107 gnd.n2326 585
R9660 gnd.n6215 gnd.n2326 585
R9661 gnd.n3892 gnd.n3891 585
R9662 gnd.n3889 gnd.n3821 585
R9663 gnd.n3888 gnd.n3887 585
R9664 gnd.n3886 gnd.n3885 585
R9665 gnd.n3884 gnd.n3825 585
R9666 gnd.n3882 gnd.n3881 585
R9667 gnd.n3880 gnd.n3826 585
R9668 gnd.n3879 gnd.n3878 585
R9669 gnd.n3876 gnd.n3831 585
R9670 gnd.n3874 gnd.n3873 585
R9671 gnd.n3872 gnd.n3832 585
R9672 gnd.n3871 gnd.n3870 585
R9673 gnd.n3868 gnd.n3837 585
R9674 gnd.n3866 gnd.n3865 585
R9675 gnd.n3864 gnd.n3838 585
R9676 gnd.n3863 gnd.n3862 585
R9677 gnd.n3860 gnd.n3843 585
R9678 gnd.n3858 gnd.n3857 585
R9679 gnd.n3845 gnd.n3844 585
R9680 gnd.n3844 gnd.n2314 585
R9681 gnd.n3670 gnd.n3669 585
R9682 gnd.n3668 gnd.n3375 585
R9683 gnd.n3377 gnd.n3376 585
R9684 gnd.n3657 gnd.n3656 585
R9685 gnd.n3655 gnd.n3654 585
R9686 gnd.n3643 gnd.n3387 585
R9687 gnd.n3645 gnd.n3644 585
R9688 gnd.n3642 gnd.n3393 585
R9689 gnd.n3392 gnd.n3391 585
R9690 gnd.n3633 gnd.n3632 585
R9691 gnd.n3631 gnd.n3630 585
R9692 gnd.n3619 gnd.n3399 585
R9693 gnd.n3621 gnd.n3620 585
R9694 gnd.n3618 gnd.n3405 585
R9695 gnd.n3404 gnd.n3403 585
R9696 gnd.n3609 gnd.n3608 585
R9697 gnd.n3607 gnd.n3606 585
R9698 gnd.n3412 gnd.n3411 585
R9699 gnd.n3597 gnd.n2536 585
R9700 gnd.n4372 gnd.n2536 585
R9701 gnd.n2542 gnd.n2534 585
R9702 gnd.n6086 gnd.n2534 585
R9703 gnd.n6078 gnd.n6077 585
R9704 gnd.n6079 gnd.n6078 585
R9705 gnd.n2541 gnd.n2525 585
R9706 gnd.n6092 gnd.n2525 585
R9707 gnd.n4231 gnd.n4229 585
R9708 gnd.n4229 gnd.n4228 585
R9709 gnd.n4232 gnd.n2515 585
R9710 gnd.n6098 gnd.n2515 585
R9711 gnd.n4233 gnd.n3698 585
R9712 gnd.n4222 gnd.n3698 585
R9713 gnd.n3696 gnd.n2504 585
R9714 gnd.n6104 gnd.n2504 585
R9715 gnd.n4237 gnd.n3695 585
R9716 gnd.n4217 gnd.n3695 585
R9717 gnd.n4238 gnd.n2494 585
R9718 gnd.n6110 gnd.n2494 585
R9719 gnd.n4239 gnd.n3694 585
R9720 gnd.n4213 gnd.n3694 585
R9721 gnd.n3691 gnd.n2483 585
R9722 gnd.n6116 gnd.n2483 585
R9723 gnd.n4244 gnd.n4243 585
R9724 gnd.n4245 gnd.n4244 585
R9725 gnd.n3690 gnd.n2474 585
R9726 gnd.n6122 gnd.n2474 585
R9727 gnd.n4205 gnd.n4204 585
R9728 gnd.n4206 gnd.n4205 585
R9729 gnd.n3701 gnd.n2463 585
R9730 gnd.n6128 gnd.n2463 585
R9731 gnd.n4200 gnd.n4199 585
R9732 gnd.n4199 gnd.n4198 585
R9733 gnd.n3703 gnd.n2453 585
R9734 gnd.n6134 gnd.n2453 585
R9735 gnd.n4191 gnd.n4190 585
R9736 gnd.n4192 gnd.n4191 585
R9737 gnd.n3706 gnd.n2445 585
R9738 gnd.n6141 gnd.n2445 585
R9739 gnd.n4186 gnd.n4185 585
R9740 gnd.n4185 gnd.n4184 585
R9741 gnd.n3708 gnd.n2436 585
R9742 gnd.n6147 gnd.n2436 585
R9743 gnd.n4177 gnd.n4176 585
R9744 gnd.n4178 gnd.n4177 585
R9745 gnd.n3712 gnd.n2428 585
R9746 gnd.n6154 gnd.n2428 585
R9747 gnd.n4172 gnd.n4171 585
R9748 gnd.n4171 gnd.n4170 585
R9749 gnd.n3714 gnd.n2418 585
R9750 gnd.n6160 gnd.n2418 585
R9751 gnd.n4163 gnd.n4162 585
R9752 gnd.n4164 gnd.n4163 585
R9753 gnd.n3717 gnd.n2409 585
R9754 gnd.n6167 gnd.n2409 585
R9755 gnd.n4158 gnd.n4157 585
R9756 gnd.n4157 gnd.n4156 585
R9757 gnd.n3719 gnd.n2400 585
R9758 gnd.n6173 gnd.n2400 585
R9759 gnd.n4149 gnd.n4148 585
R9760 gnd.n4150 gnd.n4149 585
R9761 gnd.n3723 gnd.n2389 585
R9762 gnd.n6179 gnd.n2389 585
R9763 gnd.n4144 gnd.n4143 585
R9764 gnd.n4143 gnd.n4142 585
R9765 gnd.n3725 gnd.n2379 585
R9766 gnd.n6185 gnd.n2379 585
R9767 gnd.n4135 gnd.n4134 585
R9768 gnd.n4136 gnd.n4135 585
R9769 gnd.n3728 gnd.n2368 585
R9770 gnd.n6191 gnd.n2368 585
R9771 gnd.n4130 gnd.n4129 585
R9772 gnd.n4129 gnd.n4128 585
R9773 gnd.n3730 gnd.n2359 585
R9774 gnd.n6197 gnd.n2359 585
R9775 gnd.n4121 gnd.n4120 585
R9776 gnd.n4122 gnd.n4121 585
R9777 gnd.n3815 gnd.n2348 585
R9778 gnd.n6203 gnd.n2348 585
R9779 gnd.n4116 gnd.n4115 585
R9780 gnd.n4115 gnd.n4114 585
R9781 gnd.n3817 gnd.n2336 585
R9782 gnd.n6209 gnd.n2336 585
R9783 gnd.n3850 gnd.n3849 585
R9784 gnd.n3849 gnd.n3848 585
R9785 gnd.n3851 gnd.n2324 585
R9786 gnd.n6215 gnd.n2324 585
R9787 gnd.n2212 gnd.n2211 585
R9788 gnd.n2213 gnd.n2212 585
R9789 gnd.n918 gnd.n917 585
R9790 gnd.n924 gnd.n917 585
R9791 gnd.n2187 gnd.n936 585
R9792 gnd.n936 gnd.n923 585
R9793 gnd.n2189 gnd.n2188 585
R9794 gnd.n2190 gnd.n2189 585
R9795 gnd.n937 gnd.n935 585
R9796 gnd.n935 gnd.n931 585
R9797 gnd.n1921 gnd.n1920 585
R9798 gnd.n1920 gnd.n1919 585
R9799 gnd.n942 gnd.n941 585
R9800 gnd.n1890 gnd.n942 585
R9801 gnd.n1910 gnd.n1909 585
R9802 gnd.n1909 gnd.n1908 585
R9803 gnd.n949 gnd.n948 585
R9804 gnd.n1896 gnd.n949 585
R9805 gnd.n1866 gnd.n969 585
R9806 gnd.n969 gnd.n968 585
R9807 gnd.n1868 gnd.n1867 585
R9808 gnd.n1869 gnd.n1868 585
R9809 gnd.n970 gnd.n967 585
R9810 gnd.n978 gnd.n967 585
R9811 gnd.n1844 gnd.n990 585
R9812 gnd.n990 gnd.n977 585
R9813 gnd.n1846 gnd.n1845 585
R9814 gnd.n1847 gnd.n1846 585
R9815 gnd.n991 gnd.n989 585
R9816 gnd.n989 gnd.n985 585
R9817 gnd.n1832 gnd.n1831 585
R9818 gnd.n1831 gnd.n1830 585
R9819 gnd.n996 gnd.n995 585
R9820 gnd.n1006 gnd.n996 585
R9821 gnd.n1821 gnd.n1820 585
R9822 gnd.n1820 gnd.n1819 585
R9823 gnd.n1003 gnd.n1002 585
R9824 gnd.n1807 gnd.n1003 585
R9825 gnd.n1779 gnd.n1023 585
R9826 gnd.n1023 gnd.n1013 585
R9827 gnd.n1781 gnd.n1780 585
R9828 gnd.n1782 gnd.n1781 585
R9829 gnd.n1024 gnd.n1022 585
R9830 gnd.n1032 gnd.n1022 585
R9831 gnd.n1757 gnd.n1044 585
R9832 gnd.n1044 gnd.n1031 585
R9833 gnd.n1759 gnd.n1758 585
R9834 gnd.n1760 gnd.n1759 585
R9835 gnd.n1045 gnd.n1043 585
R9836 gnd.n1043 gnd.n1039 585
R9837 gnd.n1745 gnd.n1744 585
R9838 gnd.n1744 gnd.n1743 585
R9839 gnd.n1050 gnd.n1049 585
R9840 gnd.n1059 gnd.n1050 585
R9841 gnd.n1734 gnd.n1733 585
R9842 gnd.n1733 gnd.n1732 585
R9843 gnd.n1057 gnd.n1056 585
R9844 gnd.n1720 gnd.n1057 585
R9845 gnd.n1158 gnd.n1157 585
R9846 gnd.n1158 gnd.n1066 585
R9847 gnd.n1677 gnd.n1676 585
R9848 gnd.n1676 gnd.n1675 585
R9849 gnd.n1678 gnd.n1152 585
R9850 gnd.n1163 gnd.n1152 585
R9851 gnd.n1680 gnd.n1679 585
R9852 gnd.n1681 gnd.n1680 585
R9853 gnd.n1153 gnd.n1151 585
R9854 gnd.n1176 gnd.n1151 585
R9855 gnd.n1136 gnd.n1135 585
R9856 gnd.n1139 gnd.n1136 585
R9857 gnd.n1691 gnd.n1690 585
R9858 gnd.n1690 gnd.n1689 585
R9859 gnd.n1692 gnd.n1130 585
R9860 gnd.n1651 gnd.n1130 585
R9861 gnd.n1694 gnd.n1693 585
R9862 gnd.n1695 gnd.n1694 585
R9863 gnd.n1131 gnd.n1129 585
R9864 gnd.n1190 gnd.n1129 585
R9865 gnd.n1643 gnd.n1642 585
R9866 gnd.n1642 gnd.n1641 585
R9867 gnd.n1187 gnd.n1186 585
R9868 gnd.n1625 gnd.n1187 585
R9869 gnd.n1612 gnd.n1206 585
R9870 gnd.n1206 gnd.n1205 585
R9871 gnd.n1614 gnd.n1613 585
R9872 gnd.n1615 gnd.n1614 585
R9873 gnd.n1207 gnd.n1204 585
R9874 gnd.n1213 gnd.n1204 585
R9875 gnd.n1593 gnd.n1592 585
R9876 gnd.n1594 gnd.n1593 585
R9877 gnd.n1224 gnd.n1223 585
R9878 gnd.n1223 gnd.n1219 585
R9879 gnd.n1583 gnd.n1582 585
R9880 gnd.n1584 gnd.n1583 585
R9881 gnd.n1234 gnd.n1233 585
R9882 gnd.n1239 gnd.n1233 585
R9883 gnd.n1561 gnd.n1252 585
R9884 gnd.n1252 gnd.n1238 585
R9885 gnd.n1563 gnd.n1562 585
R9886 gnd.n1564 gnd.n1563 585
R9887 gnd.n1253 gnd.n1251 585
R9888 gnd.n1251 gnd.n1247 585
R9889 gnd.n1552 gnd.n1551 585
R9890 gnd.n1553 gnd.n1552 585
R9891 gnd.n1260 gnd.n1259 585
R9892 gnd.n1264 gnd.n1259 585
R9893 gnd.n1529 gnd.n1281 585
R9894 gnd.n1281 gnd.n1263 585
R9895 gnd.n1531 gnd.n1530 585
R9896 gnd.n1532 gnd.n1531 585
R9897 gnd.n1282 gnd.n1280 585
R9898 gnd.n1280 gnd.n1271 585
R9899 gnd.n1524 gnd.n1523 585
R9900 gnd.n1523 gnd.n1522 585
R9901 gnd.n1329 gnd.n1328 585
R9902 gnd.n1330 gnd.n1329 585
R9903 gnd.n1483 gnd.n1482 585
R9904 gnd.n1484 gnd.n1483 585
R9905 gnd.n1339 gnd.n1338 585
R9906 gnd.n1338 gnd.n1337 585
R9907 gnd.n1478 gnd.n1477 585
R9908 gnd.n1477 gnd.n1476 585
R9909 gnd.n1342 gnd.n1341 585
R9910 gnd.n1343 gnd.n1342 585
R9911 gnd.n1467 gnd.n1466 585
R9912 gnd.n1468 gnd.n1467 585
R9913 gnd.n1350 gnd.n1349 585
R9914 gnd.n1459 gnd.n1349 585
R9915 gnd.n1462 gnd.n1461 585
R9916 gnd.n1461 gnd.n1460 585
R9917 gnd.n1353 gnd.n1352 585
R9918 gnd.n1354 gnd.n1353 585
R9919 gnd.n1448 gnd.n1447 585
R9920 gnd.n1446 gnd.n1372 585
R9921 gnd.n1445 gnd.n1371 585
R9922 gnd.n1450 gnd.n1371 585
R9923 gnd.n1444 gnd.n1443 585
R9924 gnd.n1442 gnd.n1441 585
R9925 gnd.n1440 gnd.n1439 585
R9926 gnd.n1438 gnd.n1437 585
R9927 gnd.n1436 gnd.n1435 585
R9928 gnd.n1434 gnd.n1433 585
R9929 gnd.n1432 gnd.n1431 585
R9930 gnd.n1430 gnd.n1429 585
R9931 gnd.n1428 gnd.n1427 585
R9932 gnd.n1426 gnd.n1425 585
R9933 gnd.n1424 gnd.n1423 585
R9934 gnd.n1422 gnd.n1421 585
R9935 gnd.n1420 gnd.n1419 585
R9936 gnd.n1418 gnd.n1417 585
R9937 gnd.n1416 gnd.n1415 585
R9938 gnd.n1414 gnd.n1413 585
R9939 gnd.n1412 gnd.n1411 585
R9940 gnd.n1410 gnd.n1409 585
R9941 gnd.n1408 gnd.n1407 585
R9942 gnd.n1406 gnd.n1405 585
R9943 gnd.n1404 gnd.n1403 585
R9944 gnd.n1402 gnd.n1401 585
R9945 gnd.n1359 gnd.n1358 585
R9946 gnd.n1453 gnd.n1452 585
R9947 gnd.n2216 gnd.n2215 585
R9948 gnd.n2218 gnd.n2217 585
R9949 gnd.n2220 gnd.n2219 585
R9950 gnd.n2222 gnd.n2221 585
R9951 gnd.n2224 gnd.n2223 585
R9952 gnd.n2226 gnd.n2225 585
R9953 gnd.n2228 gnd.n2227 585
R9954 gnd.n2230 gnd.n2229 585
R9955 gnd.n2232 gnd.n2231 585
R9956 gnd.n2234 gnd.n2233 585
R9957 gnd.n2236 gnd.n2235 585
R9958 gnd.n2238 gnd.n2237 585
R9959 gnd.n2240 gnd.n2239 585
R9960 gnd.n2242 gnd.n2241 585
R9961 gnd.n2244 gnd.n2243 585
R9962 gnd.n2246 gnd.n2245 585
R9963 gnd.n2248 gnd.n2247 585
R9964 gnd.n2250 gnd.n2249 585
R9965 gnd.n2252 gnd.n2251 585
R9966 gnd.n2254 gnd.n2253 585
R9967 gnd.n2256 gnd.n2255 585
R9968 gnd.n2258 gnd.n2257 585
R9969 gnd.n2260 gnd.n2259 585
R9970 gnd.n2262 gnd.n2261 585
R9971 gnd.n2264 gnd.n2263 585
R9972 gnd.n2265 gnd.n885 585
R9973 gnd.n2266 gnd.n843 585
R9974 gnd.n2304 gnd.n843 585
R9975 gnd.n2214 gnd.n915 585
R9976 gnd.n2214 gnd.n2213 585
R9977 gnd.n1883 gnd.n914 585
R9978 gnd.n924 gnd.n914 585
R9979 gnd.n1885 gnd.n1884 585
R9980 gnd.n1884 gnd.n923 585
R9981 gnd.n1886 gnd.n933 585
R9982 gnd.n2190 gnd.n933 585
R9983 gnd.n1888 gnd.n1887 585
R9984 gnd.n1887 gnd.n931 585
R9985 gnd.n1889 gnd.n944 585
R9986 gnd.n1919 gnd.n944 585
R9987 gnd.n1892 gnd.n1891 585
R9988 gnd.n1891 gnd.n1890 585
R9989 gnd.n1893 gnd.n951 585
R9990 gnd.n1908 gnd.n951 585
R9991 gnd.n1895 gnd.n1894 585
R9992 gnd.n1896 gnd.n1895 585
R9993 gnd.n961 gnd.n960 585
R9994 gnd.n968 gnd.n960 585
R9995 gnd.n1871 gnd.n1870 585
R9996 gnd.n1870 gnd.n1869 585
R9997 gnd.n964 gnd.n963 585
R9998 gnd.n978 gnd.n964 585
R9999 gnd.n1795 gnd.n1794 585
R10000 gnd.n1794 gnd.n977 585
R10001 gnd.n1796 gnd.n987 585
R10002 gnd.n1847 gnd.n987 585
R10003 gnd.n1798 gnd.n1797 585
R10004 gnd.n1797 gnd.n985 585
R10005 gnd.n1799 gnd.n998 585
R10006 gnd.n1830 gnd.n998 585
R10007 gnd.n1801 gnd.n1800 585
R10008 gnd.n1800 gnd.n1006 585
R10009 gnd.n1802 gnd.n1005 585
R10010 gnd.n1819 gnd.n1005 585
R10011 gnd.n1804 gnd.n1803 585
R10012 gnd.n1807 gnd.n1804 585
R10013 gnd.n1016 gnd.n1015 585
R10014 gnd.n1015 gnd.n1013 585
R10015 gnd.n1784 gnd.n1783 585
R10016 gnd.n1783 gnd.n1782 585
R10017 gnd.n1019 gnd.n1018 585
R10018 gnd.n1032 gnd.n1019 585
R10019 gnd.n1708 gnd.n1707 585
R10020 gnd.n1707 gnd.n1031 585
R10021 gnd.n1709 gnd.n1041 585
R10022 gnd.n1760 gnd.n1041 585
R10023 gnd.n1711 gnd.n1710 585
R10024 gnd.n1710 gnd.n1039 585
R10025 gnd.n1712 gnd.n1052 585
R10026 gnd.n1743 gnd.n1052 585
R10027 gnd.n1714 gnd.n1713 585
R10028 gnd.n1713 gnd.n1059 585
R10029 gnd.n1715 gnd.n1058 585
R10030 gnd.n1732 gnd.n1058 585
R10031 gnd.n1717 gnd.n1716 585
R10032 gnd.n1720 gnd.n1717 585
R10033 gnd.n1069 gnd.n1068 585
R10034 gnd.n1068 gnd.n1066 585
R10035 gnd.n1160 gnd.n1159 585
R10036 gnd.n1675 gnd.n1159 585
R10037 gnd.n1162 gnd.n1161 585
R10038 gnd.n1163 gnd.n1162 585
R10039 gnd.n1173 gnd.n1149 585
R10040 gnd.n1681 gnd.n1149 585
R10041 gnd.n1175 gnd.n1174 585
R10042 gnd.n1176 gnd.n1175 585
R10043 gnd.n1172 gnd.n1171 585
R10044 gnd.n1172 gnd.n1139 585
R10045 gnd.n1170 gnd.n1137 585
R10046 gnd.n1689 gnd.n1137 585
R10047 gnd.n1126 gnd.n1124 585
R10048 gnd.n1651 gnd.n1126 585
R10049 gnd.n1697 gnd.n1696 585
R10050 gnd.n1696 gnd.n1695 585
R10051 gnd.n1125 gnd.n1123 585
R10052 gnd.n1190 gnd.n1125 585
R10053 gnd.n1622 gnd.n1189 585
R10054 gnd.n1641 gnd.n1189 585
R10055 gnd.n1624 gnd.n1623 585
R10056 gnd.n1625 gnd.n1624 585
R10057 gnd.n1199 gnd.n1198 585
R10058 gnd.n1205 gnd.n1198 585
R10059 gnd.n1617 gnd.n1616 585
R10060 gnd.n1616 gnd.n1615 585
R10061 gnd.n1202 gnd.n1201 585
R10062 gnd.n1213 gnd.n1202 585
R10063 gnd.n1502 gnd.n1221 585
R10064 gnd.n1594 gnd.n1221 585
R10065 gnd.n1504 gnd.n1503 585
R10066 gnd.n1503 gnd.n1219 585
R10067 gnd.n1505 gnd.n1232 585
R10068 gnd.n1584 gnd.n1232 585
R10069 gnd.n1507 gnd.n1506 585
R10070 gnd.n1507 gnd.n1239 585
R10071 gnd.n1509 gnd.n1508 585
R10072 gnd.n1508 gnd.n1238 585
R10073 gnd.n1510 gnd.n1249 585
R10074 gnd.n1564 gnd.n1249 585
R10075 gnd.n1512 gnd.n1511 585
R10076 gnd.n1511 gnd.n1247 585
R10077 gnd.n1513 gnd.n1258 585
R10078 gnd.n1553 gnd.n1258 585
R10079 gnd.n1515 gnd.n1514 585
R10080 gnd.n1515 gnd.n1264 585
R10081 gnd.n1517 gnd.n1516 585
R10082 gnd.n1516 gnd.n1263 585
R10083 gnd.n1518 gnd.n1279 585
R10084 gnd.n1532 gnd.n1279 585
R10085 gnd.n1519 gnd.n1332 585
R10086 gnd.n1332 gnd.n1271 585
R10087 gnd.n1521 gnd.n1520 585
R10088 gnd.n1522 gnd.n1521 585
R10089 gnd.n1333 gnd.n1331 585
R10090 gnd.n1331 gnd.n1330 585
R10091 gnd.n1486 gnd.n1485 585
R10092 gnd.n1485 gnd.n1484 585
R10093 gnd.n1336 gnd.n1335 585
R10094 gnd.n1337 gnd.n1336 585
R10095 gnd.n1475 gnd.n1474 585
R10096 gnd.n1476 gnd.n1475 585
R10097 gnd.n1345 gnd.n1344 585
R10098 gnd.n1344 gnd.n1343 585
R10099 gnd.n1470 gnd.n1469 585
R10100 gnd.n1469 gnd.n1468 585
R10101 gnd.n1348 gnd.n1347 585
R10102 gnd.n1459 gnd.n1348 585
R10103 gnd.n1458 gnd.n1457 585
R10104 gnd.n1460 gnd.n1458 585
R10105 gnd.n1356 gnd.n1355 585
R10106 gnd.n1355 gnd.n1354 585
R10107 gnd.n7345 gnd.n7344 585
R10108 gnd.n7346 gnd.n7345 585
R10109 gnd.n156 gnd.n155 585
R10110 gnd.n7339 gnd.n156 585
R10111 gnd.n7354 gnd.n7353 585
R10112 gnd.n7353 gnd.n7352 585
R10113 gnd.n7355 gnd.n151 585
R10114 gnd.n5636 gnd.n151 585
R10115 gnd.n7357 gnd.n7356 585
R10116 gnd.n7358 gnd.n7357 585
R10117 gnd.n136 gnd.n135 585
R10118 gnd.n5642 gnd.n136 585
R10119 gnd.n7366 gnd.n7365 585
R10120 gnd.n7365 gnd.n7364 585
R10121 gnd.n7367 gnd.n131 585
R10122 gnd.n5695 gnd.n131 585
R10123 gnd.n7369 gnd.n7368 585
R10124 gnd.n7370 gnd.n7369 585
R10125 gnd.n115 gnd.n114 585
R10126 gnd.n5701 gnd.n115 585
R10127 gnd.n7378 gnd.n7377 585
R10128 gnd.n7377 gnd.n7376 585
R10129 gnd.n7379 gnd.n110 585
R10130 gnd.n5707 gnd.n110 585
R10131 gnd.n7381 gnd.n7380 585
R10132 gnd.n7382 gnd.n7381 585
R10133 gnd.n96 gnd.n95 585
R10134 gnd.n5713 gnd.n96 585
R10135 gnd.n7390 gnd.n7389 585
R10136 gnd.n7389 gnd.n7388 585
R10137 gnd.n7391 gnd.n90 585
R10138 gnd.n5719 gnd.n90 585
R10139 gnd.n7393 gnd.n7392 585
R10140 gnd.n7394 gnd.n7393 585
R10141 gnd.n91 gnd.n89 585
R10142 gnd.n5610 gnd.n89 585
R10143 gnd.n5731 gnd.n5730 585
R10144 gnd.n5730 gnd.n5729 585
R10145 gnd.n5732 gnd.n71 585
R10146 gnd.n7402 gnd.n71 585
R10147 gnd.n5733 gnd.n5419 585
R10148 gnd.n5599 gnd.n5419 585
R10149 gnd.n5735 gnd.n5734 585
R10150 gnd.n5742 gnd.n5735 585
R10151 gnd.n5420 gnd.n5418 585
R10152 gnd.n5418 gnd.n5414 585
R10153 gnd.n5587 gnd.n5586 585
R10154 gnd.n5586 gnd.n5407 585
R10155 gnd.n5399 gnd.n5398 585
R10156 gnd.n5751 gnd.n5399 585
R10157 gnd.n5758 gnd.n5757 585
R10158 gnd.n5757 gnd.n5756 585
R10159 gnd.n5759 gnd.n5394 585
R10160 gnd.n5580 gnd.n5394 585
R10161 gnd.n5761 gnd.n5760 585
R10162 gnd.n5762 gnd.n5761 585
R10163 gnd.n5380 gnd.n5379 585
R10164 gnd.n5564 gnd.n5380 585
R10165 gnd.n5770 gnd.n5769 585
R10166 gnd.n5769 gnd.n5768 585
R10167 gnd.n5771 gnd.n5375 585
R10168 gnd.n5525 gnd.n5375 585
R10169 gnd.n5773 gnd.n5772 585
R10170 gnd.n5774 gnd.n5773 585
R10171 gnd.n5360 gnd.n5359 585
R10172 gnd.n5516 gnd.n5360 585
R10173 gnd.n5782 gnd.n5781 585
R10174 gnd.n5781 gnd.n5780 585
R10175 gnd.n5783 gnd.n5355 585
R10176 gnd.n5510 gnd.n5355 585
R10177 gnd.n5785 gnd.n5784 585
R10178 gnd.n5786 gnd.n5785 585
R10179 gnd.n5340 gnd.n5339 585
R10180 gnd.n5539 gnd.n5340 585
R10181 gnd.n5794 gnd.n5793 585
R10182 gnd.n5793 gnd.n5792 585
R10183 gnd.n5795 gnd.n5334 585
R10184 gnd.n5503 gnd.n5334 585
R10185 gnd.n5797 gnd.n5796 585
R10186 gnd.n5798 gnd.n5797 585
R10187 gnd.n5335 gnd.n5318 585
R10188 gnd.n5495 gnd.n5318 585
R10189 gnd.n5805 gnd.n5319 585
R10190 gnd.n5805 gnd.n5804 585
R10191 gnd.n5806 gnd.n2815 585
R10192 gnd.n5807 gnd.n5806 585
R10193 gnd.n5317 gnd.n5316 585
R10194 gnd.n5315 gnd.n2824 585
R10195 gnd.n2826 gnd.n2825 585
R10196 gnd.n5308 gnd.n5215 585
R10197 gnd.n5307 gnd.n5216 585
R10198 gnd.n5223 gnd.n5217 585
R10199 gnd.n5300 gnd.n5224 585
R10200 gnd.n5299 gnd.n5225 585
R10201 gnd.n5227 gnd.n5226 585
R10202 gnd.n5292 gnd.n5235 585
R10203 gnd.n5291 gnd.n5236 585
R10204 gnd.n5243 gnd.n5237 585
R10205 gnd.n5284 gnd.n5244 585
R10206 gnd.n5283 gnd.n5245 585
R10207 gnd.n5247 gnd.n5246 585
R10208 gnd.n5276 gnd.n5255 585
R10209 gnd.n5275 gnd.n5256 585
R10210 gnd.n5260 gnd.n5257 585
R10211 gnd.n5268 gnd.n2744 585
R10212 gnd.n5927 gnd.n2744 585
R10213 gnd.n7333 gnd.n7332 585
R10214 gnd.n181 gnd.n180 585
R10215 gnd.n239 gnd.n238 585
R10216 gnd.n191 gnd.n190 585
R10217 gnd.n234 gnd.n233 585
R10218 gnd.n232 gnd.n231 585
R10219 gnd.n230 gnd.n229 585
R10220 gnd.n223 gnd.n193 585
R10221 gnd.n225 gnd.n224 585
R10222 gnd.n222 gnd.n221 585
R10223 gnd.n220 gnd.n219 585
R10224 gnd.n213 gnd.n195 585
R10225 gnd.n215 gnd.n214 585
R10226 gnd.n212 gnd.n211 585
R10227 gnd.n210 gnd.n209 585
R10228 gnd.n203 gnd.n197 585
R10229 gnd.n205 gnd.n204 585
R10230 gnd.n202 gnd.n201 585
R10231 gnd.n200 gnd.n171 585
R10232 gnd.n7330 gnd.n171 585
R10233 gnd.n7336 gnd.n169 585
R10234 gnd.n7346 gnd.n169 585
R10235 gnd.n7338 gnd.n7337 585
R10236 gnd.n7339 gnd.n7338 585
R10237 gnd.n175 gnd.n159 585
R10238 gnd.n7352 gnd.n159 585
R10239 gnd.n5635 gnd.n5634 585
R10240 gnd.n5636 gnd.n5635 585
R10241 gnd.n5629 gnd.n149 585
R10242 gnd.n7358 gnd.n149 585
R10243 gnd.n5644 gnd.n5643 585
R10244 gnd.n5643 gnd.n5642 585
R10245 gnd.n5645 gnd.n138 585
R10246 gnd.n7364 gnd.n138 585
R10247 gnd.n5647 gnd.n5646 585
R10248 gnd.n5695 gnd.n5647 585
R10249 gnd.n5622 gnd.n129 585
R10250 gnd.n7370 gnd.n129 585
R10251 gnd.n5703 gnd.n5702 585
R10252 gnd.n5702 gnd.n5701 585
R10253 gnd.n5704 gnd.n118 585
R10254 gnd.n7376 gnd.n118 585
R10255 gnd.n5706 gnd.n5705 585
R10256 gnd.n5707 gnd.n5706 585
R10257 gnd.n5437 gnd.n108 585
R10258 gnd.n7382 gnd.n108 585
R10259 gnd.n5715 gnd.n5714 585
R10260 gnd.n5714 gnd.n5713 585
R10261 gnd.n5716 gnd.n98 585
R10262 gnd.n7388 gnd.n98 585
R10263 gnd.n5718 gnd.n5717 585
R10264 gnd.n5719 gnd.n5718 585
R10265 gnd.n5433 gnd.n87 585
R10266 gnd.n7394 gnd.n87 585
R10267 gnd.n5609 gnd.n5608 585
R10268 gnd.n5610 gnd.n5609 585
R10269 gnd.n68 gnd.n67 585
R10270 gnd.n5729 gnd.n68 585
R10271 gnd.n7404 gnd.n7403 585
R10272 gnd.n7403 gnd.n7402 585
R10273 gnd.n7405 gnd.n66 585
R10274 gnd.n5599 gnd.n66 585
R10275 gnd.n5416 gnd.n64 585
R10276 gnd.n5742 gnd.n5416 585
R10277 gnd.n5572 gnd.n5571 585
R10278 gnd.n5571 gnd.n5414 585
R10279 gnd.n5573 gnd.n5570 585
R10280 gnd.n5570 gnd.n5407 585
R10281 gnd.n5574 gnd.n5406 585
R10282 gnd.n5751 gnd.n5406 585
R10283 gnd.n5441 gnd.n5402 585
R10284 gnd.n5756 gnd.n5402 585
R10285 gnd.n5579 gnd.n5578 585
R10286 gnd.n5580 gnd.n5579 585
R10287 gnd.n5440 gnd.n5392 585
R10288 gnd.n5762 gnd.n5392 585
R10289 gnd.n5566 gnd.n5565 585
R10290 gnd.n5565 gnd.n5564 585
R10291 gnd.n5443 gnd.n5383 585
R10292 gnd.n5768 gnd.n5383 585
R10293 gnd.n5527 gnd.n5526 585
R10294 gnd.n5526 gnd.n5525 585
R10295 gnd.n5485 gnd.n5373 585
R10296 gnd.n5774 gnd.n5373 585
R10297 gnd.n5531 gnd.n5484 585
R10298 gnd.n5516 gnd.n5484 585
R10299 gnd.n5532 gnd.n5363 585
R10300 gnd.n5780 gnd.n5363 585
R10301 gnd.n5533 gnd.n5483 585
R10302 gnd.n5510 gnd.n5483 585
R10303 gnd.n5480 gnd.n5353 585
R10304 gnd.n5786 gnd.n5353 585
R10305 gnd.n5538 gnd.n5537 585
R10306 gnd.n5539 gnd.n5538 585
R10307 gnd.n5479 gnd.n5343 585
R10308 gnd.n5792 gnd.n5343 585
R10309 gnd.n5502 gnd.n5501 585
R10310 gnd.n5503 gnd.n5502 585
R10311 gnd.n5487 gnd.n5332 585
R10312 gnd.n5798 gnd.n5332 585
R10313 gnd.n5497 gnd.n5496 585
R10314 gnd.n5496 gnd.n5495 585
R10315 gnd.n5491 gnd.n5320 585
R10316 gnd.n5804 gnd.n5320 585
R10317 gnd.n5490 gnd.n2821 585
R10318 gnd.n5807 gnd.n2821 585
R10319 gnd.n2199 gnd.n865 585
R10320 gnd.n865 gnd.n842 585
R10321 gnd.n2200 gnd.n926 585
R10322 gnd.n926 gnd.n916 585
R10323 gnd.n2202 gnd.n2201 585
R10324 gnd.n2203 gnd.n2202 585
R10325 gnd.n927 gnd.n925 585
R10326 gnd.n934 gnd.n925 585
R10327 gnd.n2193 gnd.n2192 585
R10328 gnd.n2192 gnd.n2191 585
R10329 gnd.n930 gnd.n929 585
R10330 gnd.n1918 gnd.n930 585
R10331 gnd.n1904 gnd.n953 585
R10332 gnd.n953 gnd.n943 585
R10333 gnd.n1906 gnd.n1905 585
R10334 gnd.n1907 gnd.n1906 585
R10335 gnd.n954 gnd.n952 585
R10336 gnd.n952 gnd.n950 585
R10337 gnd.n1899 gnd.n1898 585
R10338 gnd.n1898 gnd.n1897 585
R10339 gnd.n957 gnd.n956 585
R10340 gnd.n966 gnd.n957 585
R10341 gnd.n1855 gnd.n980 585
R10342 gnd.n980 gnd.n965 585
R10343 gnd.n1857 gnd.n1856 585
R10344 gnd.n1858 gnd.n1857 585
R10345 gnd.n981 gnd.n979 585
R10346 gnd.n988 gnd.n979 585
R10347 gnd.n1850 gnd.n1849 585
R10348 gnd.n1849 gnd.n1848 585
R10349 gnd.n984 gnd.n983 585
R10350 gnd.n1829 gnd.n984 585
R10351 gnd.n1815 gnd.n1008 585
R10352 gnd.n1008 gnd.n997 585
R10353 gnd.n1817 gnd.n1816 585
R10354 gnd.n1818 gnd.n1817 585
R10355 gnd.n1009 gnd.n1007 585
R10356 gnd.n1806 gnd.n1007 585
R10357 gnd.n1810 gnd.n1809 585
R10358 gnd.n1809 gnd.n1808 585
R10359 gnd.n1012 gnd.n1011 585
R10360 gnd.n1021 gnd.n1012 585
R10361 gnd.n1768 gnd.n1034 585
R10362 gnd.n1034 gnd.n1020 585
R10363 gnd.n1770 gnd.n1769 585
R10364 gnd.n1771 gnd.n1770 585
R10365 gnd.n1035 gnd.n1033 585
R10366 gnd.n1042 gnd.n1033 585
R10367 gnd.n1763 gnd.n1762 585
R10368 gnd.n1762 gnd.n1761 585
R10369 gnd.n1038 gnd.n1037 585
R10370 gnd.n1742 gnd.n1038 585
R10371 gnd.n1728 gnd.n1061 585
R10372 gnd.n1061 gnd.n1051 585
R10373 gnd.n1730 gnd.n1729 585
R10374 gnd.n1731 gnd.n1730 585
R10375 gnd.n1062 gnd.n1060 585
R10376 gnd.n1719 gnd.n1060 585
R10377 gnd.n1723 gnd.n1722 585
R10378 gnd.n1722 gnd.n1721 585
R10379 gnd.n1065 gnd.n1064 585
R10380 gnd.n1674 gnd.n1065 585
R10381 gnd.n1167 gnd.n1166 585
R10382 gnd.n1168 gnd.n1167 585
R10383 gnd.n1147 gnd.n1146 585
R10384 gnd.n1150 gnd.n1147 585
R10385 gnd.n1684 gnd.n1683 585
R10386 gnd.n1683 gnd.n1682 585
R10387 gnd.n1685 gnd.n1141 585
R10388 gnd.n1177 gnd.n1141 585
R10389 gnd.n1687 gnd.n1686 585
R10390 gnd.n1688 gnd.n1687 585
R10391 gnd.n1142 gnd.n1140 585
R10392 gnd.n1652 gnd.n1140 585
R10393 gnd.n1636 gnd.n1635 585
R10394 gnd.n1635 gnd.n1128 585
R10395 gnd.n1637 gnd.n1192 585
R10396 gnd.n1192 gnd.n1127 585
R10397 gnd.n1639 gnd.n1638 585
R10398 gnd.n1640 gnd.n1639 585
R10399 gnd.n1193 gnd.n1191 585
R10400 gnd.n1191 gnd.n1188 585
R10401 gnd.n1628 gnd.n1627 585
R10402 gnd.n1627 gnd.n1626 585
R10403 gnd.n1196 gnd.n1195 585
R10404 gnd.n1203 gnd.n1196 585
R10405 gnd.n1602 gnd.n1601 585
R10406 gnd.n1603 gnd.n1602 585
R10407 gnd.n1215 gnd.n1214 585
R10408 gnd.n1222 gnd.n1214 585
R10409 gnd.n1597 gnd.n1596 585
R10410 gnd.n1596 gnd.n1595 585
R10411 gnd.n1218 gnd.n1217 585
R10412 gnd.n1585 gnd.n1218 585
R10413 gnd.n1572 gnd.n1242 585
R10414 gnd.n1242 gnd.n1241 585
R10415 gnd.n1574 gnd.n1573 585
R10416 gnd.n1575 gnd.n1574 585
R10417 gnd.n1243 gnd.n1240 585
R10418 gnd.n1250 gnd.n1240 585
R10419 gnd.n1567 gnd.n1566 585
R10420 gnd.n1566 gnd.n1565 585
R10421 gnd.n1246 gnd.n1245 585
R10422 gnd.n1554 gnd.n1246 585
R10423 gnd.n1541 gnd.n1267 585
R10424 gnd.n1267 gnd.n1266 585
R10425 gnd.n1543 gnd.n1542 585
R10426 gnd.n1544 gnd.n1543 585
R10427 gnd.n1537 gnd.n1265 585
R10428 gnd.n1536 gnd.n1535 585
R10429 gnd.n1270 gnd.n1269 585
R10430 gnd.n1533 gnd.n1270 585
R10431 gnd.n1292 gnd.n1291 585
R10432 gnd.n1295 gnd.n1294 585
R10433 gnd.n1293 gnd.n1288 585
R10434 gnd.n1300 gnd.n1299 585
R10435 gnd.n1302 gnd.n1301 585
R10436 gnd.n1305 gnd.n1304 585
R10437 gnd.n1303 gnd.n1286 585
R10438 gnd.n1310 gnd.n1309 585
R10439 gnd.n1312 gnd.n1311 585
R10440 gnd.n1315 gnd.n1314 585
R10441 gnd.n1313 gnd.n1284 585
R10442 gnd.n1320 gnd.n1319 585
R10443 gnd.n1324 gnd.n1321 585
R10444 gnd.n1325 gnd.n1262 585
R10445 gnd.n2205 gnd.n880 585
R10446 gnd.n2272 gnd.n2271 585
R10447 gnd.n2274 gnd.n2273 585
R10448 gnd.n2276 gnd.n2275 585
R10449 gnd.n2278 gnd.n2277 585
R10450 gnd.n2280 gnd.n2279 585
R10451 gnd.n2282 gnd.n2281 585
R10452 gnd.n2284 gnd.n2283 585
R10453 gnd.n2286 gnd.n2285 585
R10454 gnd.n2288 gnd.n2287 585
R10455 gnd.n2290 gnd.n2289 585
R10456 gnd.n2292 gnd.n2291 585
R10457 gnd.n2294 gnd.n2293 585
R10458 gnd.n2297 gnd.n2296 585
R10459 gnd.n2295 gnd.n868 585
R10460 gnd.n2301 gnd.n866 585
R10461 gnd.n2303 gnd.n2302 585
R10462 gnd.n2304 gnd.n2303 585
R10463 gnd.n2206 gnd.n921 585
R10464 gnd.n2206 gnd.n842 585
R10465 gnd.n2208 gnd.n2207 585
R10466 gnd.n2207 gnd.n916 585
R10467 gnd.n2204 gnd.n920 585
R10468 gnd.n2204 gnd.n2203 585
R10469 gnd.n2183 gnd.n922 585
R10470 gnd.n934 gnd.n922 585
R10471 gnd.n2182 gnd.n932 585
R10472 gnd.n2191 gnd.n932 585
R10473 gnd.n1917 gnd.n939 585
R10474 gnd.n1918 gnd.n1917 585
R10475 gnd.n1916 gnd.n1915 585
R10476 gnd.n1916 gnd.n943 585
R10477 gnd.n1914 gnd.n945 585
R10478 gnd.n1907 gnd.n945 585
R10479 gnd.n958 gnd.n946 585
R10480 gnd.n958 gnd.n950 585
R10481 gnd.n1863 gnd.n959 585
R10482 gnd.n1897 gnd.n959 585
R10483 gnd.n1862 gnd.n1861 585
R10484 gnd.n1861 gnd.n966 585
R10485 gnd.n1860 gnd.n974 585
R10486 gnd.n1860 gnd.n965 585
R10487 gnd.n1859 gnd.n976 585
R10488 gnd.n1859 gnd.n1858 585
R10489 gnd.n1838 gnd.n975 585
R10490 gnd.n988 gnd.n975 585
R10491 gnd.n1837 gnd.n986 585
R10492 gnd.n1848 gnd.n986 585
R10493 gnd.n1828 gnd.n993 585
R10494 gnd.n1829 gnd.n1828 585
R10495 gnd.n1827 gnd.n1826 585
R10496 gnd.n1827 gnd.n997 585
R10497 gnd.n1825 gnd.n999 585
R10498 gnd.n1818 gnd.n999 585
R10499 gnd.n1805 gnd.n1000 585
R10500 gnd.n1806 gnd.n1805 585
R10501 gnd.n1776 gnd.n1014 585
R10502 gnd.n1808 gnd.n1014 585
R10503 gnd.n1775 gnd.n1774 585
R10504 gnd.n1774 gnd.n1021 585
R10505 gnd.n1773 gnd.n1028 585
R10506 gnd.n1773 gnd.n1020 585
R10507 gnd.n1772 gnd.n1030 585
R10508 gnd.n1772 gnd.n1771 585
R10509 gnd.n1751 gnd.n1029 585
R10510 gnd.n1042 gnd.n1029 585
R10511 gnd.n1750 gnd.n1040 585
R10512 gnd.n1761 gnd.n1040 585
R10513 gnd.n1741 gnd.n1047 585
R10514 gnd.n1742 gnd.n1741 585
R10515 gnd.n1740 gnd.n1739 585
R10516 gnd.n1740 gnd.n1051 585
R10517 gnd.n1738 gnd.n1053 585
R10518 gnd.n1731 gnd.n1053 585
R10519 gnd.n1718 gnd.n1054 585
R10520 gnd.n1719 gnd.n1718 585
R10521 gnd.n1671 gnd.n1067 585
R10522 gnd.n1721 gnd.n1067 585
R10523 gnd.n1673 gnd.n1672 585
R10524 gnd.n1674 gnd.n1673 585
R10525 gnd.n1666 gnd.n1169 585
R10526 gnd.n1169 gnd.n1168 585
R10527 gnd.n1664 gnd.n1663 585
R10528 gnd.n1663 gnd.n1150 585
R10529 gnd.n1661 gnd.n1148 585
R10530 gnd.n1682 gnd.n1148 585
R10531 gnd.n1179 gnd.n1178 585
R10532 gnd.n1178 gnd.n1177 585
R10533 gnd.n1655 gnd.n1138 585
R10534 gnd.n1688 gnd.n1138 585
R10535 gnd.n1654 gnd.n1653 585
R10536 gnd.n1653 gnd.n1652 585
R10537 gnd.n1650 gnd.n1181 585
R10538 gnd.n1650 gnd.n1128 585
R10539 gnd.n1649 gnd.n1648 585
R10540 gnd.n1649 gnd.n1127 585
R10541 gnd.n1184 gnd.n1183 585
R10542 gnd.n1640 gnd.n1183 585
R10543 gnd.n1608 gnd.n1607 585
R10544 gnd.n1607 gnd.n1188 585
R10545 gnd.n1609 gnd.n1197 585
R10546 gnd.n1626 gnd.n1197 585
R10547 gnd.n1606 gnd.n1605 585
R10548 gnd.n1605 gnd.n1203 585
R10549 gnd.n1604 gnd.n1211 585
R10550 gnd.n1604 gnd.n1603 585
R10551 gnd.n1589 gnd.n1212 585
R10552 gnd.n1222 gnd.n1212 585
R10553 gnd.n1588 gnd.n1220 585
R10554 gnd.n1595 gnd.n1220 585
R10555 gnd.n1587 gnd.n1586 585
R10556 gnd.n1586 gnd.n1585 585
R10557 gnd.n1231 gnd.n1228 585
R10558 gnd.n1241 gnd.n1231 585
R10559 gnd.n1577 gnd.n1576 585
R10560 gnd.n1576 gnd.n1575 585
R10561 gnd.n1237 gnd.n1236 585
R10562 gnd.n1250 gnd.n1237 585
R10563 gnd.n1557 gnd.n1248 585
R10564 gnd.n1565 gnd.n1248 585
R10565 gnd.n1556 gnd.n1555 585
R10566 gnd.n1555 gnd.n1554 585
R10567 gnd.n1257 gnd.n1255 585
R10568 gnd.n1266 gnd.n1257 585
R10569 gnd.n1546 gnd.n1545 585
R10570 gnd.n1545 gnd.n1544 585
R10571 gnd.n5126 gnd.n5125 585
R10572 gnd.n5127 gnd.n5126 585
R10573 gnd.n2891 gnd.n2889 585
R10574 gnd.n2889 gnd.n2885 585
R10575 gnd.n4999 gnd.n4998 585
R10576 gnd.n5000 gnd.n4999 585
R10577 gnd.n4997 gnd.n2964 585
R10578 gnd.n2969 gnd.n2964 585
R10579 gnd.n4996 gnd.n4995 585
R10580 gnd.n4995 gnd.n4994 585
R10581 gnd.n2966 gnd.n2965 585
R10582 gnd.n4971 gnd.n2966 585
R10583 gnd.n4983 gnd.n4982 585
R10584 gnd.n4984 gnd.n4983 585
R10585 gnd.n4981 gnd.n2980 585
R10586 gnd.n2980 gnd.n2976 585
R10587 gnd.n4980 gnd.n4979 585
R10588 gnd.n4979 gnd.n4978 585
R10589 gnd.n2982 gnd.n2981 585
R10590 gnd.n4911 gnd.n2982 585
R10591 gnd.n4964 gnd.n4963 585
R10592 gnd.n4965 gnd.n4964 585
R10593 gnd.n4962 gnd.n2989 585
R10594 gnd.n2989 gnd.n2988 585
R10595 gnd.n4961 gnd.n4960 585
R10596 gnd.n4960 gnd.n4959 585
R10597 gnd.n2991 gnd.n2990 585
R10598 gnd.n3004 gnd.n2991 585
R10599 gnd.n4946 gnd.n4945 585
R10600 gnd.n4947 gnd.n4946 585
R10601 gnd.n4944 gnd.n3005 585
R10602 gnd.n3005 gnd.n3001 585
R10603 gnd.n4943 gnd.n4942 585
R10604 gnd.n4942 gnd.n4941 585
R10605 gnd.n3007 gnd.n3006 585
R10606 gnd.n4819 gnd.n3007 585
R10607 gnd.n4886 gnd.n4885 585
R10608 gnd.n4886 gnd.n3015 585
R10609 gnd.n4888 gnd.n4887 585
R10610 gnd.n4887 gnd.t133 585
R10611 gnd.n4889 gnd.n3028 585
R10612 gnd.n3028 gnd.n3026 585
R10613 gnd.n4891 gnd.n4890 585
R10614 gnd.n4892 gnd.n4891 585
R10615 gnd.n4884 gnd.n3027 585
R10616 gnd.n3027 gnd.n3022 585
R10617 gnd.n4883 gnd.n4882 585
R10618 gnd.n4882 gnd.n4881 585
R10619 gnd.n3030 gnd.n3029 585
R10620 gnd.n4815 gnd.n3030 585
R10621 gnd.n4854 gnd.n4853 585
R10622 gnd.n4854 gnd.n3039 585
R10623 gnd.n4856 gnd.n4855 585
R10624 gnd.n4855 gnd.n3038 585
R10625 gnd.n4857 gnd.n3052 585
R10626 gnd.n4842 gnd.n3052 585
R10627 gnd.n4859 gnd.n4858 585
R10628 gnd.n4860 gnd.n4859 585
R10629 gnd.n4852 gnd.n3051 585
R10630 gnd.n3051 gnd.n3046 585
R10631 gnd.n4851 gnd.n4850 585
R10632 gnd.n4850 gnd.n4849 585
R10633 gnd.n3054 gnd.n3053 585
R10634 gnd.n3061 gnd.n3054 585
R10635 gnd.n4808 gnd.n4807 585
R10636 gnd.n4809 gnd.n4808 585
R10637 gnd.n4806 gnd.n3063 585
R10638 gnd.n3063 gnd.n3060 585
R10639 gnd.n4805 gnd.n4804 585
R10640 gnd.n4804 gnd.n4803 585
R10641 gnd.n3065 gnd.n3064 585
R10642 gnd.n3079 gnd.n3065 585
R10643 gnd.n4790 gnd.n4789 585
R10644 gnd.n4791 gnd.n4790 585
R10645 gnd.n4788 gnd.n3080 585
R10646 gnd.n3080 gnd.n3076 585
R10647 gnd.n4787 gnd.n4786 585
R10648 gnd.n4786 gnd.n4785 585
R10649 gnd.n3082 gnd.n3081 585
R10650 gnd.n3083 gnd.n3082 585
R10651 gnd.n4745 gnd.n4744 585
R10652 gnd.n4745 gnd.n3092 585
R10653 gnd.n4747 gnd.n4746 585
R10654 gnd.n4746 gnd.n3091 585
R10655 gnd.n4748 gnd.n3106 585
R10656 gnd.n3106 gnd.n3104 585
R10657 gnd.n4750 gnd.n4749 585
R10658 gnd.n4751 gnd.n4750 585
R10659 gnd.n4743 gnd.n3105 585
R10660 gnd.n4737 gnd.n3105 585
R10661 gnd.n4742 gnd.n4741 585
R10662 gnd.n4741 gnd.n4740 585
R10663 gnd.n3108 gnd.n3107 585
R10664 gnd.n3109 gnd.n3108 585
R10665 gnd.n4713 gnd.n4712 585
R10666 gnd.n4714 gnd.n4713 585
R10667 gnd.n4711 gnd.n3115 585
R10668 gnd.n4707 gnd.n3115 585
R10669 gnd.n4710 gnd.n4709 585
R10670 gnd.n4709 gnd.n4708 585
R10671 gnd.n3117 gnd.n3116 585
R10672 gnd.n4694 gnd.n3117 585
R10673 gnd.n4683 gnd.n3134 585
R10674 gnd.n3134 gnd.n3127 585
R10675 gnd.n4685 gnd.n4684 585
R10676 gnd.n4686 gnd.n4685 585
R10677 gnd.n4682 gnd.n3133 585
R10678 gnd.n3139 gnd.n3133 585
R10679 gnd.n4681 gnd.n4680 585
R10680 gnd.n4680 gnd.n4679 585
R10681 gnd.n3136 gnd.n3135 585
R10682 gnd.n4655 gnd.n3136 585
R10683 gnd.n4667 gnd.n4666 585
R10684 gnd.n4668 gnd.n4667 585
R10685 gnd.n4665 gnd.n3149 585
R10686 gnd.n3149 gnd.n3145 585
R10687 gnd.n4664 gnd.n4663 585
R10688 gnd.n4663 gnd.n4662 585
R10689 gnd.n3151 gnd.n3150 585
R10690 gnd.n3158 gnd.n3151 585
R10691 gnd.n4649 gnd.n4648 585
R10692 gnd.n4650 gnd.n4649 585
R10693 gnd.n4647 gnd.n3160 585
R10694 gnd.n3160 gnd.n3157 585
R10695 gnd.n4646 gnd.n4645 585
R10696 gnd.n4645 gnd.t6 585
R10697 gnd.n3162 gnd.n3161 585
R10698 gnd.n3175 gnd.n3162 585
R10699 gnd.n4632 gnd.n4631 585
R10700 gnd.n4633 gnd.n4632 585
R10701 gnd.n4630 gnd.n3176 585
R10702 gnd.n4625 gnd.n3176 585
R10703 gnd.n4629 gnd.n4628 585
R10704 gnd.n4628 gnd.n4627 585
R10705 gnd.n3178 gnd.n3177 585
R10706 gnd.n4615 gnd.n3178 585
R10707 gnd.n4613 gnd.n4612 585
R10708 gnd.n4614 gnd.n4613 585
R10709 gnd.n4611 gnd.n3186 585
R10710 gnd.n4577 gnd.n3186 585
R10711 gnd.n4610 gnd.n4609 585
R10712 gnd.n4609 gnd.n4608 585
R10713 gnd.n3188 gnd.n3187 585
R10714 gnd.n3189 gnd.n3188 585
R10715 gnd.n4592 gnd.n4591 585
R10716 gnd.n4593 gnd.n4592 585
R10717 gnd.n4590 gnd.n3201 585
R10718 gnd.n3201 gnd.n3198 585
R10719 gnd.n4589 gnd.n4588 585
R10720 gnd.n4588 gnd.n4587 585
R10721 gnd.n3203 gnd.n3202 585
R10722 gnd.n3492 gnd.n3203 585
R10723 gnd.n4572 gnd.n4571 585
R10724 gnd.n4573 gnd.n4572 585
R10725 gnd.n4570 gnd.n3209 585
R10726 gnd.n3215 gnd.n3209 585
R10727 gnd.n4569 gnd.n4568 585
R10728 gnd.n4568 gnd.n4567 585
R10729 gnd.n3211 gnd.n3210 585
R10730 gnd.n3289 gnd.n3211 585
R10731 gnd.n4553 gnd.n4552 585
R10732 gnd.n4554 gnd.n4553 585
R10733 gnd.n4551 gnd.n3225 585
R10734 gnd.n3225 gnd.n3222 585
R10735 gnd.n4549 gnd.n4548 585
R10736 gnd.n3247 gnd.n3246 585
R10737 gnd.n4545 gnd.n4544 585
R10738 gnd.n4546 gnd.n4545 585
R10739 gnd.n4543 gnd.n3282 585
R10740 gnd.n4542 gnd.n4541 585
R10741 gnd.n4540 gnd.n4539 585
R10742 gnd.n4538 gnd.n4537 585
R10743 gnd.n4536 gnd.n4535 585
R10744 gnd.n4534 gnd.n4533 585
R10745 gnd.n4532 gnd.n4531 585
R10746 gnd.n4530 gnd.n4529 585
R10747 gnd.n4528 gnd.n4527 585
R10748 gnd.n4526 gnd.n4525 585
R10749 gnd.n4524 gnd.n4523 585
R10750 gnd.n4522 gnd.n4521 585
R10751 gnd.n4520 gnd.n4519 585
R10752 gnd.n4518 gnd.n4517 585
R10753 gnd.n4516 gnd.n4515 585
R10754 gnd.n4514 gnd.n4513 585
R10755 gnd.n4512 gnd.n4511 585
R10756 gnd.n4510 gnd.n4509 585
R10757 gnd.n4508 gnd.n4507 585
R10758 gnd.n4506 gnd.n4505 585
R10759 gnd.n4504 gnd.n4503 585
R10760 gnd.n4502 gnd.n4501 585
R10761 gnd.n4500 gnd.n4499 585
R10762 gnd.n4498 gnd.n4497 585
R10763 gnd.n4496 gnd.n4495 585
R10764 gnd.n4494 gnd.n4493 585
R10765 gnd.n4492 gnd.n4491 585
R10766 gnd.n4490 gnd.n4489 585
R10767 gnd.n4488 gnd.n4487 585
R10768 gnd.n4486 gnd.n4485 585
R10769 gnd.n4484 gnd.n3358 585
R10770 gnd.n3357 gnd.n3356 585
R10771 gnd.n3355 gnd.n3354 585
R10772 gnd.n3352 gnd.n3351 585
R10773 gnd.n3350 gnd.n3349 585
R10774 gnd.n3348 gnd.n3347 585
R10775 gnd.n3346 gnd.n3345 585
R10776 gnd.n3344 gnd.n3343 585
R10777 gnd.n3342 gnd.n3341 585
R10778 gnd.n3340 gnd.n3339 585
R10779 gnd.n3338 gnd.n3337 585
R10780 gnd.n3336 gnd.n3335 585
R10781 gnd.n3334 gnd.n3333 585
R10782 gnd.n3332 gnd.n3331 585
R10783 gnd.n3330 gnd.n3329 585
R10784 gnd.n3328 gnd.n3327 585
R10785 gnd.n3326 gnd.n3325 585
R10786 gnd.n3324 gnd.n3323 585
R10787 gnd.n3322 gnd.n3321 585
R10788 gnd.n3320 gnd.n3319 585
R10789 gnd.n3318 gnd.n3317 585
R10790 gnd.n3316 gnd.n3315 585
R10791 gnd.n3314 gnd.n3313 585
R10792 gnd.n3312 gnd.n3311 585
R10793 gnd.n3310 gnd.n3309 585
R10794 gnd.n3308 gnd.n3307 585
R10795 gnd.n3306 gnd.n3305 585
R10796 gnd.n3304 gnd.n3303 585
R10797 gnd.n3302 gnd.n3301 585
R10798 gnd.n3300 gnd.n3299 585
R10799 gnd.n3298 gnd.n3297 585
R10800 gnd.n3296 gnd.n3295 585
R10801 gnd.n5007 gnd.n5006 585
R10802 gnd.n5008 gnd.n2960 585
R10803 gnd.n5010 gnd.n5009 585
R10804 gnd.n5012 gnd.n2958 585
R10805 gnd.n5014 gnd.n5013 585
R10806 gnd.n5015 gnd.n2957 585
R10807 gnd.n5017 gnd.n5016 585
R10808 gnd.n5019 gnd.n2955 585
R10809 gnd.n5021 gnd.n5020 585
R10810 gnd.n5022 gnd.n2954 585
R10811 gnd.n5024 gnd.n5023 585
R10812 gnd.n5026 gnd.n2952 585
R10813 gnd.n5028 gnd.n5027 585
R10814 gnd.n5029 gnd.n2951 585
R10815 gnd.n5031 gnd.n5030 585
R10816 gnd.n5033 gnd.n2949 585
R10817 gnd.n5035 gnd.n5034 585
R10818 gnd.n5036 gnd.n2948 585
R10819 gnd.n5038 gnd.n5037 585
R10820 gnd.n5040 gnd.n2946 585
R10821 gnd.n5042 gnd.n5041 585
R10822 gnd.n5043 gnd.n2945 585
R10823 gnd.n5045 gnd.n5044 585
R10824 gnd.n5047 gnd.n2943 585
R10825 gnd.n5049 gnd.n5048 585
R10826 gnd.n5050 gnd.n2942 585
R10827 gnd.n5052 gnd.n5051 585
R10828 gnd.n5054 gnd.n2940 585
R10829 gnd.n5056 gnd.n5055 585
R10830 gnd.n5058 gnd.n2937 585
R10831 gnd.n5060 gnd.n5059 585
R10832 gnd.n5062 gnd.n2936 585
R10833 gnd.n5063 gnd.n2877 585
R10834 gnd.n5066 gnd.n2777 585
R10835 gnd.n5068 gnd.n5067 585
R10836 gnd.n5070 gnd.n2934 585
R10837 gnd.n5072 gnd.n5071 585
R10838 gnd.n5074 gnd.n2931 585
R10839 gnd.n5076 gnd.n5075 585
R10840 gnd.n5078 gnd.n2929 585
R10841 gnd.n5080 gnd.n5079 585
R10842 gnd.n5081 gnd.n2928 585
R10843 gnd.n5083 gnd.n5082 585
R10844 gnd.n5085 gnd.n2926 585
R10845 gnd.n5087 gnd.n5086 585
R10846 gnd.n5088 gnd.n2925 585
R10847 gnd.n5090 gnd.n5089 585
R10848 gnd.n5092 gnd.n2923 585
R10849 gnd.n5094 gnd.n5093 585
R10850 gnd.n5095 gnd.n2922 585
R10851 gnd.n5097 gnd.n5096 585
R10852 gnd.n5099 gnd.n2920 585
R10853 gnd.n5101 gnd.n5100 585
R10854 gnd.n5102 gnd.n2919 585
R10855 gnd.n5104 gnd.n5103 585
R10856 gnd.n5106 gnd.n2917 585
R10857 gnd.n5108 gnd.n5107 585
R10858 gnd.n5109 gnd.n2916 585
R10859 gnd.n5111 gnd.n5110 585
R10860 gnd.n5113 gnd.n2914 585
R10861 gnd.n5115 gnd.n5114 585
R10862 gnd.n5116 gnd.n2913 585
R10863 gnd.n5118 gnd.n5117 585
R10864 gnd.n5120 gnd.n2911 585
R10865 gnd.n5122 gnd.n5121 585
R10866 gnd.n5123 gnd.n2890 585
R10867 gnd.n5004 gnd.n2887 585
R10868 gnd.n5127 gnd.n2887 585
R10869 gnd.n5003 gnd.n5002 585
R10870 gnd.n5002 gnd.n2885 585
R10871 gnd.n5001 gnd.n2961 585
R10872 gnd.n5001 gnd.n5000 585
R10873 gnd.n4969 gnd.n2962 585
R10874 gnd.n2969 gnd.n2962 585
R10875 gnd.n4970 gnd.n2967 585
R10876 gnd.n4994 gnd.n2967 585
R10877 gnd.n4973 gnd.n4972 585
R10878 gnd.n4972 gnd.n4971 585
R10879 gnd.n4974 gnd.n2978 585
R10880 gnd.n4984 gnd.n2978 585
R10881 gnd.n4975 gnd.n2985 585
R10882 gnd.n2985 gnd.n2976 585
R10883 gnd.n4977 gnd.n4976 585
R10884 gnd.n4978 gnd.n4977 585
R10885 gnd.n4968 gnd.n2984 585
R10886 gnd.n4911 gnd.n2984 585
R10887 gnd.n4967 gnd.n4966 585
R10888 gnd.n4966 gnd.n4965 585
R10889 gnd.n2987 gnd.n2986 585
R10890 gnd.n2988 gnd.n2987 585
R10891 gnd.n4821 gnd.n2993 585
R10892 gnd.n4959 gnd.n2993 585
R10893 gnd.n4823 gnd.n4822 585
R10894 gnd.n4822 gnd.n3004 585
R10895 gnd.n4824 gnd.n3003 585
R10896 gnd.n4947 gnd.n3003 585
R10897 gnd.n4826 gnd.n4825 585
R10898 gnd.n4825 gnd.n3001 585
R10899 gnd.n4827 gnd.n3008 585
R10900 gnd.n4941 gnd.n3008 585
R10901 gnd.n4828 gnd.n4820 585
R10902 gnd.n4820 gnd.n4819 585
R10903 gnd.n4830 gnd.n4829 585
R10904 gnd.n4830 gnd.n3015 585
R10905 gnd.n4831 gnd.n4817 585
R10906 gnd.n4831 gnd.t133 585
R10907 gnd.n4833 gnd.n4832 585
R10908 gnd.n4832 gnd.n3026 585
R10909 gnd.n4834 gnd.n3024 585
R10910 gnd.n4892 gnd.n3024 585
R10911 gnd.n4836 gnd.n4835 585
R10912 gnd.n4835 gnd.n3022 585
R10913 gnd.n4837 gnd.n3031 585
R10914 gnd.n4881 gnd.n3031 585
R10915 gnd.n4838 gnd.n4816 585
R10916 gnd.n4816 gnd.n4815 585
R10917 gnd.n4840 gnd.n4839 585
R10918 gnd.n4840 gnd.n3039 585
R10919 gnd.n4841 gnd.n4813 585
R10920 gnd.n4841 gnd.n3038 585
R10921 gnd.n4844 gnd.n4843 585
R10922 gnd.n4843 gnd.n4842 585
R10923 gnd.n4845 gnd.n3048 585
R10924 gnd.n4860 gnd.n3048 585
R10925 gnd.n4846 gnd.n3057 585
R10926 gnd.n3057 gnd.n3046 585
R10927 gnd.n4848 gnd.n4847 585
R10928 gnd.n4849 gnd.n4848 585
R10929 gnd.n4812 gnd.n3056 585
R10930 gnd.n3061 gnd.n3056 585
R10931 gnd.n4811 gnd.n4810 585
R10932 gnd.n4810 gnd.n4809 585
R10933 gnd.n3059 gnd.n3058 585
R10934 gnd.n3060 gnd.n3059 585
R10935 gnd.n4721 gnd.n3067 585
R10936 gnd.n4803 gnd.n3067 585
R10937 gnd.n4723 gnd.n4722 585
R10938 gnd.n4722 gnd.n3079 585
R10939 gnd.n4724 gnd.n3078 585
R10940 gnd.n4791 gnd.n3078 585
R10941 gnd.n4726 gnd.n4725 585
R10942 gnd.n4725 gnd.n3076 585
R10943 gnd.n4727 gnd.n3084 585
R10944 gnd.n4785 gnd.n3084 585
R10945 gnd.n4728 gnd.n4720 585
R10946 gnd.n4720 gnd.n3083 585
R10947 gnd.n4730 gnd.n4729 585
R10948 gnd.n4730 gnd.n3092 585
R10949 gnd.n4731 gnd.n4719 585
R10950 gnd.n4731 gnd.n3091 585
R10951 gnd.n4733 gnd.n4732 585
R10952 gnd.n4732 gnd.n3104 585
R10953 gnd.n4734 gnd.n3102 585
R10954 gnd.n4751 gnd.n3102 585
R10955 gnd.n4736 gnd.n4735 585
R10956 gnd.n4737 gnd.n4736 585
R10957 gnd.n4718 gnd.n3110 585
R10958 gnd.n4740 gnd.n3110 585
R10959 gnd.n4717 gnd.n4716 585
R10960 gnd.n4716 gnd.n3109 585
R10961 gnd.n4715 gnd.n3112 585
R10962 gnd.n4715 gnd.n4714 585
R10963 gnd.n4690 gnd.n3113 585
R10964 gnd.n4707 gnd.n3113 585
R10965 gnd.n4691 gnd.n3119 585
R10966 gnd.n4708 gnd.n3119 585
R10967 gnd.n4693 gnd.n4692 585
R10968 gnd.n4694 gnd.n4693 585
R10969 gnd.n4689 gnd.n3129 585
R10970 gnd.n3129 gnd.n3127 585
R10971 gnd.n4688 gnd.n4687 585
R10972 gnd.n4687 gnd.n4686 585
R10973 gnd.n3131 gnd.n3130 585
R10974 gnd.n3139 gnd.n3131 585
R10975 gnd.n4654 gnd.n3137 585
R10976 gnd.n4679 gnd.n3137 585
R10977 gnd.n4657 gnd.n4656 585
R10978 gnd.n4656 gnd.n4655 585
R10979 gnd.n4658 gnd.n3147 585
R10980 gnd.n4668 gnd.n3147 585
R10981 gnd.n4659 gnd.n3154 585
R10982 gnd.n3154 gnd.n3145 585
R10983 gnd.n4661 gnd.n4660 585
R10984 gnd.n4662 gnd.n4661 585
R10985 gnd.n4653 gnd.n3153 585
R10986 gnd.n3158 gnd.n3153 585
R10987 gnd.n4652 gnd.n4651 585
R10988 gnd.n4651 gnd.n4650 585
R10989 gnd.n3156 gnd.n3155 585
R10990 gnd.n3157 gnd.n3156 585
R10991 gnd.n4619 gnd.n3165 585
R10992 gnd.t6 gnd.n3165 585
R10993 gnd.n4621 gnd.n4620 585
R10994 gnd.n4620 gnd.n3175 585
R10995 gnd.n4622 gnd.n3174 585
R10996 gnd.n4633 gnd.n3174 585
R10997 gnd.n4624 gnd.n4623 585
R10998 gnd.n4625 gnd.n4624 585
R10999 gnd.n4618 gnd.n3180 585
R11000 gnd.n4627 gnd.n3180 585
R11001 gnd.n4617 gnd.n4616 585
R11002 gnd.n4616 gnd.n4615 585
R11003 gnd.n3183 gnd.n3182 585
R11004 gnd.n4614 gnd.n3183 585
R11005 gnd.n4579 gnd.n4578 585
R11006 gnd.n4578 gnd.n4577 585
R11007 gnd.n4580 gnd.n3190 585
R11008 gnd.n4608 gnd.n3190 585
R11009 gnd.n4582 gnd.n4581 585
R11010 gnd.n4581 gnd.n3189 585
R11011 gnd.n4583 gnd.n3200 585
R11012 gnd.n4593 gnd.n3200 585
R11013 gnd.n4584 gnd.n3205 585
R11014 gnd.n3205 gnd.n3198 585
R11015 gnd.n4586 gnd.n4585 585
R11016 gnd.n4587 gnd.n4586 585
R11017 gnd.n4576 gnd.n3204 585
R11018 gnd.n3492 gnd.n3204 585
R11019 gnd.n4575 gnd.n4574 585
R11020 gnd.n4574 gnd.n4573 585
R11021 gnd.n3207 gnd.n3206 585
R11022 gnd.n3215 gnd.n3207 585
R11023 gnd.n3288 gnd.n3213 585
R11024 gnd.n4567 gnd.n3213 585
R11025 gnd.n3291 gnd.n3290 585
R11026 gnd.n3290 gnd.n3289 585
R11027 gnd.n3292 gnd.n3224 585
R11028 gnd.n4554 gnd.n3224 585
R11029 gnd.n3294 gnd.n3293 585
R11030 gnd.n3294 gnd.n3222 585
R11031 gnd.n6088 gnd.n6087 585
R11032 gnd.n6087 gnd.n6086 585
R11033 gnd.n6089 gnd.n2526 585
R11034 gnd.n6079 gnd.n2526 585
R11035 gnd.n6091 gnd.n6090 585
R11036 gnd.n6092 gnd.n6091 585
R11037 gnd.n2512 gnd.n2511 585
R11038 gnd.n4228 gnd.n2512 585
R11039 gnd.n6100 gnd.n6099 585
R11040 gnd.n6099 gnd.n6098 585
R11041 gnd.n6101 gnd.n2506 585
R11042 gnd.n4222 gnd.n2506 585
R11043 gnd.n6103 gnd.n6102 585
R11044 gnd.n6104 gnd.n6103 585
R11045 gnd.n2491 gnd.n2490 585
R11046 gnd.n4217 gnd.n2491 585
R11047 gnd.n6112 gnd.n6111 585
R11048 gnd.n6111 gnd.n6110 585
R11049 gnd.n6113 gnd.n2485 585
R11050 gnd.n4213 gnd.n2485 585
R11051 gnd.n6115 gnd.n6114 585
R11052 gnd.n6116 gnd.n6115 585
R11053 gnd.n2471 gnd.n2470 585
R11054 gnd.n4245 gnd.n2471 585
R11055 gnd.n6124 gnd.n6123 585
R11056 gnd.n6123 gnd.n6122 585
R11057 gnd.n6125 gnd.n2465 585
R11058 gnd.n4206 gnd.n2465 585
R11059 gnd.n6127 gnd.n6126 585
R11060 gnd.n6128 gnd.n6127 585
R11061 gnd.n2450 gnd.n2449 585
R11062 gnd.n4198 gnd.n2450 585
R11063 gnd.n6136 gnd.n6135 585
R11064 gnd.n6135 gnd.n6134 585
R11065 gnd.n6137 gnd.n2447 585
R11066 gnd.n4192 gnd.n2447 585
R11067 gnd.n6140 gnd.n6139 585
R11068 gnd.n6141 gnd.n6140 585
R11069 gnd.n2448 gnd.n2433 585
R11070 gnd.n4184 gnd.n2433 585
R11071 gnd.n6149 gnd.n6148 585
R11072 gnd.n6148 gnd.n6147 585
R11073 gnd.n6150 gnd.n2430 585
R11074 gnd.n4178 gnd.n2430 585
R11075 gnd.n6153 gnd.n6152 585
R11076 gnd.n6154 gnd.n6153 585
R11077 gnd.n2431 gnd.n2415 585
R11078 gnd.n4170 gnd.n2415 585
R11079 gnd.n6162 gnd.n6161 585
R11080 gnd.n6161 gnd.n6160 585
R11081 gnd.n6163 gnd.n2411 585
R11082 gnd.n4164 gnd.n2411 585
R11083 gnd.n6166 gnd.n6165 585
R11084 gnd.n6167 gnd.n6166 585
R11085 gnd.n2397 gnd.n2396 585
R11086 gnd.n4156 gnd.n2397 585
R11087 gnd.n6175 gnd.n6174 585
R11088 gnd.n6174 gnd.n6173 585
R11089 gnd.n6176 gnd.n2391 585
R11090 gnd.n4150 gnd.n2391 585
R11091 gnd.n6178 gnd.n6177 585
R11092 gnd.n6179 gnd.n6178 585
R11093 gnd.n2376 gnd.n2375 585
R11094 gnd.n4142 gnd.n2376 585
R11095 gnd.n6187 gnd.n6186 585
R11096 gnd.n6186 gnd.n6185 585
R11097 gnd.n6188 gnd.n2370 585
R11098 gnd.n4136 gnd.n2370 585
R11099 gnd.n6190 gnd.n6189 585
R11100 gnd.n6191 gnd.n6190 585
R11101 gnd.n2356 gnd.n2355 585
R11102 gnd.n4128 gnd.n2356 585
R11103 gnd.n6199 gnd.n6198 585
R11104 gnd.n6198 gnd.n6197 585
R11105 gnd.n6200 gnd.n2350 585
R11106 gnd.n4122 gnd.n2350 585
R11107 gnd.n6202 gnd.n6201 585
R11108 gnd.n6203 gnd.n6202 585
R11109 gnd.n2333 gnd.n2332 585
R11110 gnd.n4114 gnd.n2333 585
R11111 gnd.n6211 gnd.n6210 585
R11112 gnd.n6210 gnd.n6209 585
R11113 gnd.n6212 gnd.n2328 585
R11114 gnd.n3848 gnd.n2328 585
R11115 gnd.n6214 gnd.n6213 585
R11116 gnd.n6215 gnd.n6214 585
R11117 gnd.n3957 gnd.n2327 585
R11118 gnd.n3960 gnd.n3959 585
R11119 gnd.n3955 gnd.n3954 585
R11120 gnd.n3954 gnd.n2314 585
R11121 gnd.n3965 gnd.n3964 585
R11122 gnd.n3967 gnd.n3953 585
R11123 gnd.n3970 gnd.n3969 585
R11124 gnd.n3951 gnd.n3950 585
R11125 gnd.n3975 gnd.n3974 585
R11126 gnd.n3977 gnd.n3949 585
R11127 gnd.n3980 gnd.n3979 585
R11128 gnd.n3947 gnd.n3946 585
R11129 gnd.n3985 gnd.n3984 585
R11130 gnd.n3987 gnd.n3945 585
R11131 gnd.n3990 gnd.n3989 585
R11132 gnd.n3943 gnd.n3942 585
R11133 gnd.n3995 gnd.n3994 585
R11134 gnd.n3997 gnd.n3938 585
R11135 gnd.n4000 gnd.n3999 585
R11136 gnd.n3936 gnd.n3935 585
R11137 gnd.n4005 gnd.n4004 585
R11138 gnd.n4007 gnd.n3934 585
R11139 gnd.n4010 gnd.n4009 585
R11140 gnd.n3932 gnd.n3931 585
R11141 gnd.n4015 gnd.n4014 585
R11142 gnd.n4017 gnd.n3930 585
R11143 gnd.n4020 gnd.n4019 585
R11144 gnd.n3928 gnd.n3927 585
R11145 gnd.n4025 gnd.n4024 585
R11146 gnd.n4027 gnd.n3926 585
R11147 gnd.n4030 gnd.n4029 585
R11148 gnd.n3924 gnd.n3923 585
R11149 gnd.n4035 gnd.n4034 585
R11150 gnd.n4037 gnd.n3922 585
R11151 gnd.n4040 gnd.n4039 585
R11152 gnd.n3920 gnd.n3919 585
R11153 gnd.n4045 gnd.n4044 585
R11154 gnd.n4047 gnd.n3918 585
R11155 gnd.n4052 gnd.n4049 585
R11156 gnd.n3916 gnd.n3915 585
R11157 gnd.n4057 gnd.n4056 585
R11158 gnd.n4059 gnd.n3914 585
R11159 gnd.n4062 gnd.n4061 585
R11160 gnd.n3912 gnd.n3911 585
R11161 gnd.n4067 gnd.n4066 585
R11162 gnd.n4069 gnd.n3910 585
R11163 gnd.n4072 gnd.n4071 585
R11164 gnd.n3908 gnd.n3907 585
R11165 gnd.n4077 gnd.n4076 585
R11166 gnd.n4079 gnd.n3906 585
R11167 gnd.n4082 gnd.n4081 585
R11168 gnd.n3904 gnd.n3903 585
R11169 gnd.n4087 gnd.n4086 585
R11170 gnd.n4089 gnd.n3902 585
R11171 gnd.n4092 gnd.n4091 585
R11172 gnd.n3900 gnd.n3899 585
R11173 gnd.n4098 gnd.n4097 585
R11174 gnd.n4100 gnd.n3898 585
R11175 gnd.n4101 gnd.n3897 585
R11176 gnd.n4104 gnd.n4103 585
R11177 gnd.n4425 gnd.n4424 585
R11178 gnd.n4427 gnd.n4420 585
R11179 gnd.n4429 gnd.n4428 585
R11180 gnd.n4430 gnd.n4413 585
R11181 gnd.n4432 gnd.n4431 585
R11182 gnd.n4434 gnd.n4411 585
R11183 gnd.n4436 gnd.n4435 585
R11184 gnd.n4437 gnd.n4406 585
R11185 gnd.n4439 gnd.n4438 585
R11186 gnd.n4441 gnd.n4404 585
R11187 gnd.n4443 gnd.n4442 585
R11188 gnd.n4444 gnd.n4399 585
R11189 gnd.n4446 gnd.n4445 585
R11190 gnd.n4448 gnd.n4397 585
R11191 gnd.n4450 gnd.n4449 585
R11192 gnd.n4451 gnd.n4392 585
R11193 gnd.n4453 gnd.n4452 585
R11194 gnd.n4455 gnd.n4391 585
R11195 gnd.n4456 gnd.n4388 585
R11196 gnd.n4459 gnd.n4458 585
R11197 gnd.n4390 gnd.n4384 585
R11198 gnd.n4463 gnd.n4381 585
R11199 gnd.n4465 gnd.n4464 585
R11200 gnd.n4467 gnd.n4379 585
R11201 gnd.n4469 gnd.n4468 585
R11202 gnd.n4470 gnd.n4374 585
R11203 gnd.n4472 gnd.n4471 585
R11204 gnd.n4474 gnd.n4373 585
R11205 gnd.n4475 gnd.n3364 585
R11206 gnd.n4478 gnd.n4477 585
R11207 gnd.n3365 gnd.n3359 585
R11208 gnd.n4324 gnd.n3360 585
R11209 gnd.n4326 gnd.n4325 585
R11210 gnd.n4328 gnd.n4327 585
R11211 gnd.n4330 gnd.n4329 585
R11212 gnd.n4332 gnd.n4331 585
R11213 gnd.n4334 gnd.n4333 585
R11214 gnd.n4336 gnd.n4335 585
R11215 gnd.n4338 gnd.n4337 585
R11216 gnd.n4341 gnd.n4340 585
R11217 gnd.n4343 gnd.n4342 585
R11218 gnd.n4345 gnd.n4344 585
R11219 gnd.n4347 gnd.n4346 585
R11220 gnd.n4349 gnd.n4348 585
R11221 gnd.n4351 gnd.n4350 585
R11222 gnd.n4353 gnd.n4352 585
R11223 gnd.n4355 gnd.n4354 585
R11224 gnd.n4357 gnd.n4356 585
R11225 gnd.n4359 gnd.n4358 585
R11226 gnd.n4361 gnd.n4360 585
R11227 gnd.n4363 gnd.n4362 585
R11228 gnd.n4365 gnd.n4364 585
R11229 gnd.n4367 gnd.n4366 585
R11230 gnd.n4368 gnd.n4294 585
R11231 gnd.n4370 gnd.n4369 585
R11232 gnd.n4295 gnd.n4293 585
R11233 gnd.n4296 gnd.n2531 585
R11234 gnd.n4372 gnd.n2531 585
R11235 gnd.n6082 gnd.n2533 585
R11236 gnd.n6086 gnd.n2533 585
R11237 gnd.n6081 gnd.n6080 585
R11238 gnd.n6080 gnd.n6079 585
R11239 gnd.n2539 gnd.n2524 585
R11240 gnd.n6092 gnd.n2524 585
R11241 gnd.n4227 gnd.n4226 585
R11242 gnd.n4228 gnd.n4227 585
R11243 gnd.n4225 gnd.n2514 585
R11244 gnd.n6098 gnd.n2514 585
R11245 gnd.n4224 gnd.n4223 585
R11246 gnd.n4223 gnd.n4222 585
R11247 gnd.n4220 gnd.n2503 585
R11248 gnd.n6104 gnd.n2503 585
R11249 gnd.n4219 gnd.n4218 585
R11250 gnd.n4218 gnd.n4217 585
R11251 gnd.n4216 gnd.n2493 585
R11252 gnd.n6110 gnd.n2493 585
R11253 gnd.n4215 gnd.n4214 585
R11254 gnd.n4214 gnd.n4213 585
R11255 gnd.n4211 gnd.n2482 585
R11256 gnd.n6116 gnd.n2482 585
R11257 gnd.n4210 gnd.n3689 585
R11258 gnd.n4245 gnd.n3689 585
R11259 gnd.n4209 gnd.n2473 585
R11260 gnd.n6122 gnd.n2473 585
R11261 gnd.n4208 gnd.n4207 585
R11262 gnd.n4207 gnd.n4206 585
R11263 gnd.n3699 gnd.n2462 585
R11264 gnd.n6128 gnd.n2462 585
R11265 gnd.n4197 gnd.n4196 585
R11266 gnd.n4198 gnd.n4197 585
R11267 gnd.n4195 gnd.n2452 585
R11268 gnd.n6134 gnd.n2452 585
R11269 gnd.n4194 gnd.n4193 585
R11270 gnd.n4193 gnd.n4192 585
R11271 gnd.n3704 gnd.n2444 585
R11272 gnd.n6141 gnd.n2444 585
R11273 gnd.n4183 gnd.n4182 585
R11274 gnd.n4184 gnd.n4183 585
R11275 gnd.n4181 gnd.n2435 585
R11276 gnd.n6147 gnd.n2435 585
R11277 gnd.n4180 gnd.n4179 585
R11278 gnd.n4179 gnd.n4178 585
R11279 gnd.n3710 gnd.n2427 585
R11280 gnd.n6154 gnd.n2427 585
R11281 gnd.n4169 gnd.n4168 585
R11282 gnd.n4170 gnd.n4169 585
R11283 gnd.n4167 gnd.n2417 585
R11284 gnd.n6160 gnd.n2417 585
R11285 gnd.n4166 gnd.n4165 585
R11286 gnd.n4165 gnd.n4164 585
R11287 gnd.n3715 gnd.n2408 585
R11288 gnd.n6167 gnd.n2408 585
R11289 gnd.n4155 gnd.n4154 585
R11290 gnd.n4156 gnd.n4155 585
R11291 gnd.n4153 gnd.n2399 585
R11292 gnd.n6173 gnd.n2399 585
R11293 gnd.n4152 gnd.n4151 585
R11294 gnd.n4151 gnd.n4150 585
R11295 gnd.n3721 gnd.n2388 585
R11296 gnd.n6179 gnd.n2388 585
R11297 gnd.n4141 gnd.n4140 585
R11298 gnd.n4142 gnd.n4141 585
R11299 gnd.n4139 gnd.n2378 585
R11300 gnd.n6185 gnd.n2378 585
R11301 gnd.n4138 gnd.n4137 585
R11302 gnd.n4137 gnd.n4136 585
R11303 gnd.n3726 gnd.n2367 585
R11304 gnd.n6191 gnd.n2367 585
R11305 gnd.n4127 gnd.n4126 585
R11306 gnd.n4128 gnd.n4127 585
R11307 gnd.n4125 gnd.n2358 585
R11308 gnd.n6197 gnd.n2358 585
R11309 gnd.n4124 gnd.n4123 585
R11310 gnd.n4123 gnd.n4122 585
R11311 gnd.n3813 gnd.n2347 585
R11312 gnd.n6203 gnd.n2347 585
R11313 gnd.n4113 gnd.n4112 585
R11314 gnd.n4114 gnd.n4113 585
R11315 gnd.n4111 gnd.n2335 585
R11316 gnd.n6209 gnd.n2335 585
R11317 gnd.n4110 gnd.n3819 585
R11318 gnd.n3848 gnd.n3819 585
R11319 gnd.n3818 gnd.n2323 585
R11320 gnd.n6215 gnd.n2323 585
R11321 gnd.n7348 gnd.n7347 585
R11322 gnd.n7347 gnd.n7346 585
R11323 gnd.n7349 gnd.n161 585
R11324 gnd.n7339 gnd.n161 585
R11325 gnd.n7351 gnd.n7350 585
R11326 gnd.n7352 gnd.n7351 585
R11327 gnd.n146 gnd.n145 585
R11328 gnd.n5636 gnd.n146 585
R11329 gnd.n7360 gnd.n7359 585
R11330 gnd.n7359 gnd.n7358 585
R11331 gnd.n7361 gnd.n140 585
R11332 gnd.n5642 gnd.n140 585
R11333 gnd.n7363 gnd.n7362 585
R11334 gnd.n7364 gnd.n7363 585
R11335 gnd.n126 gnd.n125 585
R11336 gnd.n5695 gnd.n126 585
R11337 gnd.n7372 gnd.n7371 585
R11338 gnd.n7371 gnd.n7370 585
R11339 gnd.n7373 gnd.n120 585
R11340 gnd.n5701 gnd.n120 585
R11341 gnd.n7375 gnd.n7374 585
R11342 gnd.n7376 gnd.n7375 585
R11343 gnd.n105 gnd.n104 585
R11344 gnd.n5707 gnd.n105 585
R11345 gnd.n7384 gnd.n7383 585
R11346 gnd.n7383 gnd.n7382 585
R11347 gnd.n7385 gnd.n100 585
R11348 gnd.n5713 gnd.n100 585
R11349 gnd.n7387 gnd.n7386 585
R11350 gnd.n7388 gnd.n7387 585
R11351 gnd.n84 gnd.n82 585
R11352 gnd.n5719 gnd.n84 585
R11353 gnd.n7396 gnd.n7395 585
R11354 gnd.n7395 gnd.n7394 585
R11355 gnd.n83 gnd.n75 585
R11356 gnd.n5610 gnd.n83 585
R11357 gnd.n7399 gnd.n73 585
R11358 gnd.n5729 gnd.n73 585
R11359 gnd.n7401 gnd.n7400 585
R11360 gnd.n7402 gnd.n7401 585
R11361 gnd.n5739 gnd.n72 585
R11362 gnd.n5599 gnd.n72 585
R11363 gnd.n5741 gnd.n5740 585
R11364 gnd.n5742 gnd.n5741 585
R11365 gnd.n5738 gnd.n5737 585
R11366 gnd.n5738 gnd.n5414 585
R11367 gnd.n5736 gnd.n5403 585
R11368 gnd.n5407 gnd.n5403 585
R11369 gnd.n5753 gnd.n5752 585
R11370 gnd.n5752 gnd.n5751 585
R11371 gnd.n5755 gnd.n5754 585
R11372 gnd.n5756 gnd.n5755 585
R11373 gnd.n5390 gnd.n5389 585
R11374 gnd.n5580 gnd.n5390 585
R11375 gnd.n5764 gnd.n5763 585
R11376 gnd.n5763 gnd.n5762 585
R11377 gnd.n5765 gnd.n5385 585
R11378 gnd.n5564 gnd.n5385 585
R11379 gnd.n5767 gnd.n5766 585
R11380 gnd.n5768 gnd.n5767 585
R11381 gnd.n5370 gnd.n5369 585
R11382 gnd.n5525 gnd.n5370 585
R11383 gnd.n5776 gnd.n5775 585
R11384 gnd.n5775 gnd.n5774 585
R11385 gnd.n5777 gnd.n5364 585
R11386 gnd.n5516 gnd.n5364 585
R11387 gnd.n5779 gnd.n5778 585
R11388 gnd.n5780 gnd.n5779 585
R11389 gnd.n5351 gnd.n5350 585
R11390 gnd.n5510 gnd.n5351 585
R11391 gnd.n5788 gnd.n5787 585
R11392 gnd.n5787 gnd.n5786 585
R11393 gnd.n5789 gnd.n5345 585
R11394 gnd.n5539 gnd.n5345 585
R11395 gnd.n5791 gnd.n5790 585
R11396 gnd.n5792 gnd.n5791 585
R11397 gnd.n5329 gnd.n5328 585
R11398 gnd.n5503 gnd.n5329 585
R11399 gnd.n5800 gnd.n5799 585
R11400 gnd.n5799 gnd.n5798 585
R11401 gnd.n5801 gnd.n5322 585
R11402 gnd.n5495 gnd.n5322 585
R11403 gnd.n5803 gnd.n5802 585
R11404 gnd.n5804 gnd.n5803 585
R11405 gnd.n5323 gnd.n2748 585
R11406 gnd.n5807 gnd.n2748 585
R11407 gnd.n5925 gnd.n5924 585
R11408 gnd.n5923 gnd.n2747 585
R11409 gnd.n5922 gnd.n2746 585
R11410 gnd.n5927 gnd.n2746 585
R11411 gnd.n5921 gnd.n5920 585
R11412 gnd.n5919 gnd.n5918 585
R11413 gnd.n5917 gnd.n5916 585
R11414 gnd.n5915 gnd.n5914 585
R11415 gnd.n5913 gnd.n5912 585
R11416 gnd.n5911 gnd.n5910 585
R11417 gnd.n5909 gnd.n5908 585
R11418 gnd.n5907 gnd.n5906 585
R11419 gnd.n5905 gnd.n5904 585
R11420 gnd.n5903 gnd.n5902 585
R11421 gnd.n5901 gnd.n5900 585
R11422 gnd.n5899 gnd.n5898 585
R11423 gnd.n5897 gnd.n5896 585
R11424 gnd.n5895 gnd.n5894 585
R11425 gnd.n5893 gnd.n5892 585
R11426 gnd.n5890 gnd.n5889 585
R11427 gnd.n5888 gnd.n5887 585
R11428 gnd.n5886 gnd.n5885 585
R11429 gnd.n5884 gnd.n5883 585
R11430 gnd.n5882 gnd.n5881 585
R11431 gnd.n5880 gnd.n5879 585
R11432 gnd.n5878 gnd.n5877 585
R11433 gnd.n5876 gnd.n5875 585
R11434 gnd.n5873 gnd.n5872 585
R11435 gnd.n5871 gnd.n5870 585
R11436 gnd.n5869 gnd.n5868 585
R11437 gnd.n5867 gnd.n5866 585
R11438 gnd.n5865 gnd.n5864 585
R11439 gnd.n5863 gnd.n5862 585
R11440 gnd.n5861 gnd.n5860 585
R11441 gnd.n5859 gnd.n5858 585
R11442 gnd.n5857 gnd.n5856 585
R11443 gnd.n5855 gnd.n5854 585
R11444 gnd.n5853 gnd.n5852 585
R11445 gnd.n5851 gnd.n5850 585
R11446 gnd.n5849 gnd.n5848 585
R11447 gnd.n5847 gnd.n5846 585
R11448 gnd.n5845 gnd.n5844 585
R11449 gnd.n5843 gnd.n5842 585
R11450 gnd.n5841 gnd.n5840 585
R11451 gnd.n5839 gnd.n5838 585
R11452 gnd.n5837 gnd.n5836 585
R11453 gnd.n5835 gnd.n5834 585
R11454 gnd.n5833 gnd.n5832 585
R11455 gnd.n5831 gnd.n5830 585
R11456 gnd.n5829 gnd.n5828 585
R11457 gnd.n5827 gnd.n5826 585
R11458 gnd.n5825 gnd.n5824 585
R11459 gnd.n5823 gnd.n5822 585
R11460 gnd.n5821 gnd.n5820 585
R11461 gnd.n5819 gnd.n5818 585
R11462 gnd.n5817 gnd.n5816 585
R11463 gnd.n5815 gnd.n5814 585
R11464 gnd.n2818 gnd.n2811 585
R11465 gnd.n7208 gnd.n7207 585
R11466 gnd.n7214 gnd.n7213 585
R11467 gnd.n7216 gnd.n7215 585
R11468 gnd.n7218 gnd.n7217 585
R11469 gnd.n7220 gnd.n7219 585
R11470 gnd.n7222 gnd.n7221 585
R11471 gnd.n7224 gnd.n7223 585
R11472 gnd.n7226 gnd.n7225 585
R11473 gnd.n7228 gnd.n7227 585
R11474 gnd.n7230 gnd.n7229 585
R11475 gnd.n7232 gnd.n7231 585
R11476 gnd.n7234 gnd.n7233 585
R11477 gnd.n7236 gnd.n7235 585
R11478 gnd.n7238 gnd.n7237 585
R11479 gnd.n7240 gnd.n7239 585
R11480 gnd.n7242 gnd.n7241 585
R11481 gnd.n7244 gnd.n7243 585
R11482 gnd.n7246 gnd.n7245 585
R11483 gnd.n7248 gnd.n7247 585
R11484 gnd.n7251 gnd.n7250 585
R11485 gnd.n7249 gnd.n7187 585
R11486 gnd.n7256 gnd.n7255 585
R11487 gnd.n7258 gnd.n7257 585
R11488 gnd.n7260 gnd.n7259 585
R11489 gnd.n7262 gnd.n7261 585
R11490 gnd.n7264 gnd.n7263 585
R11491 gnd.n7266 gnd.n7265 585
R11492 gnd.n7268 gnd.n7267 585
R11493 gnd.n7270 gnd.n7269 585
R11494 gnd.n7272 gnd.n7271 585
R11495 gnd.n7274 gnd.n7273 585
R11496 gnd.n7276 gnd.n7275 585
R11497 gnd.n7278 gnd.n7277 585
R11498 gnd.n7280 gnd.n7279 585
R11499 gnd.n7282 gnd.n7281 585
R11500 gnd.n7284 gnd.n7283 585
R11501 gnd.n7286 gnd.n7285 585
R11502 gnd.n7288 gnd.n7287 585
R11503 gnd.n7290 gnd.n7289 585
R11504 gnd.n7292 gnd.n7291 585
R11505 gnd.n7294 gnd.n7293 585
R11506 gnd.n7299 gnd.n7298 585
R11507 gnd.n7301 gnd.n7300 585
R11508 gnd.n7303 gnd.n7302 585
R11509 gnd.n7305 gnd.n7304 585
R11510 gnd.n7307 gnd.n7306 585
R11511 gnd.n7309 gnd.n7308 585
R11512 gnd.n7311 gnd.n7310 585
R11513 gnd.n7313 gnd.n7312 585
R11514 gnd.n7315 gnd.n7314 585
R11515 gnd.n7317 gnd.n7316 585
R11516 gnd.n7319 gnd.n7318 585
R11517 gnd.n7321 gnd.n7320 585
R11518 gnd.n7323 gnd.n7322 585
R11519 gnd.n7325 gnd.n7324 585
R11520 gnd.n7326 gnd.n7147 585
R11521 gnd.n7328 gnd.n7327 585
R11522 gnd.n7148 gnd.n7146 585
R11523 gnd.n7149 gnd.n166 585
R11524 gnd.n7330 gnd.n166 585
R11525 gnd.n7342 gnd.n168 585
R11526 gnd.n7346 gnd.n168 585
R11527 gnd.n7341 gnd.n7340 585
R11528 gnd.n7340 gnd.n7339 585
R11529 gnd.n174 gnd.n158 585
R11530 gnd.n7352 gnd.n158 585
R11531 gnd.n5638 gnd.n5637 585
R11532 gnd.n5637 gnd.n5636 585
R11533 gnd.n5639 gnd.n148 585
R11534 gnd.n7358 gnd.n148 585
R11535 gnd.n5641 gnd.n5640 585
R11536 gnd.n5642 gnd.n5641 585
R11537 gnd.n5624 gnd.n137 585
R11538 gnd.n7364 gnd.n137 585
R11539 gnd.n5697 gnd.n5696 585
R11540 gnd.n5696 gnd.n5695 585
R11541 gnd.n5698 gnd.n128 585
R11542 gnd.n7370 gnd.n128 585
R11543 gnd.n5700 gnd.n5699 585
R11544 gnd.n5701 gnd.n5700 585
R11545 gnd.n5617 gnd.n117 585
R11546 gnd.n7376 gnd.n117 585
R11547 gnd.n5709 gnd.n5708 585
R11548 gnd.n5708 gnd.n5707 585
R11549 gnd.n5710 gnd.n107 585
R11550 gnd.n7382 gnd.n107 585
R11551 gnd.n5712 gnd.n5711 585
R11552 gnd.n5713 gnd.n5712 585
R11553 gnd.n5615 gnd.n97 585
R11554 gnd.n7388 gnd.n97 585
R11555 gnd.n5614 gnd.n5432 585
R11556 gnd.n5719 gnd.n5432 585
R11557 gnd.n5613 gnd.n86 585
R11558 gnd.n7394 gnd.n86 585
R11559 gnd.n5612 gnd.n5611 585
R11560 gnd.n5611 gnd.n5610 585
R11561 gnd.n5603 gnd.n5425 585
R11562 gnd.n5729 gnd.n5425 585
R11563 gnd.n5602 gnd.n69 585
R11564 gnd.n7402 gnd.n69 585
R11565 gnd.n5601 gnd.n5600 585
R11566 gnd.n5600 gnd.n5599 585
R11567 gnd.n5593 gnd.n5415 585
R11568 gnd.n5742 gnd.n5415 585
R11569 gnd.n5592 gnd.n5591 585
R11570 gnd.n5591 gnd.n5414 585
R11571 gnd.n5590 gnd.n5438 585
R11572 gnd.n5590 gnd.n5407 585
R11573 gnd.n5584 gnd.n5405 585
R11574 gnd.n5751 gnd.n5405 585
R11575 gnd.n5583 gnd.n5401 585
R11576 gnd.n5756 gnd.n5401 585
R11577 gnd.n5582 gnd.n5581 585
R11578 gnd.n5581 gnd.n5580 585
R11579 gnd.n5439 gnd.n5391 585
R11580 gnd.n5762 gnd.n5391 585
R11581 gnd.n5521 gnd.n5444 585
R11582 gnd.n5564 gnd.n5444 585
R11583 gnd.n5522 gnd.n5382 585
R11584 gnd.n5768 gnd.n5382 585
R11585 gnd.n5524 gnd.n5523 585
R11586 gnd.n5525 gnd.n5524 585
R11587 gnd.n5519 gnd.n5372 585
R11588 gnd.n5774 gnd.n5372 585
R11589 gnd.n5518 gnd.n5517 585
R11590 gnd.n5517 gnd.n5516 585
R11591 gnd.n5513 gnd.n5362 585
R11592 gnd.n5780 gnd.n5362 585
R11593 gnd.n5512 gnd.n5511 585
R11594 gnd.n5511 gnd.n5510 585
R11595 gnd.n5509 gnd.n5352 585
R11596 gnd.n5786 gnd.n5352 585
R11597 gnd.n5508 gnd.n5478 585
R11598 gnd.n5539 gnd.n5478 585
R11599 gnd.n5506 gnd.n5342 585
R11600 gnd.n5792 gnd.n5342 585
R11601 gnd.n5505 gnd.n5504 585
R11602 gnd.n5504 gnd.n5503 585
R11603 gnd.n5486 gnd.n5331 585
R11604 gnd.n5798 gnd.n5331 585
R11605 gnd.n5494 gnd.n5493 585
R11606 gnd.n5495 gnd.n5494 585
R11607 gnd.n2819 gnd.n2817 585
R11608 gnd.n5804 gnd.n2819 585
R11609 gnd.n5809 gnd.n5808 585
R11610 gnd.n5808 gnd.n5807 585
R11611 gnd.n6234 gnd.n6233 585
R11612 gnd.n6233 gnd.n6232 585
R11613 gnd.n7103 gnd.n7102 585
R11614 gnd.n7102 gnd.n7101 585
R11615 gnd.n7106 gnd.n251 585
R11616 gnd.n251 gnd.n250 585
R11617 gnd.n7108 gnd.n7107 585
R11618 gnd.n7109 gnd.n7108 585
R11619 gnd.n249 gnd.n248 585
R11620 gnd.n7110 gnd.n249 585
R11621 gnd.n7113 gnd.n7112 585
R11622 gnd.n7112 gnd.n7111 585
R11623 gnd.n7114 gnd.n243 585
R11624 gnd.n243 gnd.n241 585
R11625 gnd.n7116 gnd.n7115 585
R11626 gnd.n7117 gnd.n7116 585
R11627 gnd.n244 gnd.n242 585
R11628 gnd.n242 gnd.n182 585
R11629 gnd.n5682 gnd.n5681 585
R11630 gnd.n5682 gnd.n170 585
R11631 gnd.n5684 gnd.n5683 585
R11632 gnd.n5683 gnd.n167 585
R11633 gnd.n5685 gnd.n5674 585
R11634 gnd.n5674 gnd.n160 585
R11635 gnd.n5687 gnd.n5686 585
R11636 gnd.n5687 gnd.n157 585
R11637 gnd.n5688 gnd.n5673 585
R11638 gnd.n5688 gnd.n150 585
R11639 gnd.n5690 gnd.n5689 585
R11640 gnd.n5689 gnd.n147 585
R11641 gnd.n5691 gnd.n5649 585
R11642 gnd.n5649 gnd.n139 585
R11643 gnd.n5693 gnd.n5692 585
R11644 gnd.n5694 gnd.n5693 585
R11645 gnd.n5650 gnd.n5648 585
R11646 gnd.n5648 gnd.n130 585
R11647 gnd.n5667 gnd.n5666 585
R11648 gnd.n5666 gnd.n127 585
R11649 gnd.n5665 gnd.n5652 585
R11650 gnd.n5665 gnd.n119 585
R11651 gnd.n5664 gnd.n5663 585
R11652 gnd.n5664 gnd.n116 585
R11653 gnd.n5654 gnd.n5653 585
R11654 gnd.n5653 gnd.n109 585
R11655 gnd.n5659 gnd.n5658 585
R11656 gnd.n5658 gnd.n106 585
R11657 gnd.n5657 gnd.n5431 585
R11658 gnd.n5431 gnd.n99 585
R11659 gnd.n5721 gnd.n5430 585
R11660 gnd.n5721 gnd.n5720 585
R11661 gnd.n5723 gnd.n5722 585
R11662 gnd.n5722 gnd.n88 585
R11663 gnd.n5724 gnd.n5427 585
R11664 gnd.n5427 gnd.n85 585
R11665 gnd.n5727 gnd.n5726 585
R11666 gnd.n5728 gnd.n5727 585
R11667 gnd.n5428 gnd.n5426 585
R11668 gnd.n5426 gnd.n70 585
R11669 gnd.n5597 gnd.n5596 585
R11670 gnd.n5598 gnd.n5597 585
R11671 gnd.n5594 gnd.n5412 585
R11672 gnd.n5417 gnd.n5412 585
R11673 gnd.n5745 gnd.n5744 585
R11674 gnd.n5744 gnd.n5743 585
R11675 gnd.n5746 gnd.n5409 585
R11676 gnd.n5413 gnd.n5409 585
R11677 gnd.n5749 gnd.n5748 585
R11678 gnd.n5750 gnd.n5749 585
R11679 gnd.n5410 gnd.n5408 585
R11680 gnd.n5408 gnd.n5404 585
R11681 gnd.n5559 gnd.n5558 585
R11682 gnd.n5558 gnd.n5400 585
R11683 gnd.n5560 gnd.n5446 585
R11684 gnd.n5446 gnd.n5393 585
R11685 gnd.n5562 gnd.n5561 585
R11686 gnd.n5563 gnd.n5562 585
R11687 gnd.n5447 gnd.n5445 585
R11688 gnd.n5445 gnd.n5384 585
R11689 gnd.n5552 gnd.n5551 585
R11690 gnd.n5551 gnd.n5381 585
R11691 gnd.n5550 gnd.n5449 585
R11692 gnd.n5550 gnd.n5374 585
R11693 gnd.n5549 gnd.n5548 585
R11694 gnd.n5549 gnd.n5371 585
R11695 gnd.n5451 gnd.n5450 585
R11696 gnd.n5515 gnd.n5450 585
R11697 gnd.n5544 gnd.n5543 585
R11698 gnd.n5543 gnd.n5361 585
R11699 gnd.n5542 gnd.n5453 585
R11700 gnd.n5542 gnd.n5354 585
R11701 gnd.n5541 gnd.n5477 585
R11702 gnd.n5541 gnd.n5540 585
R11703 gnd.n5455 gnd.n5454 585
R11704 gnd.n5454 gnd.n5344 585
R11705 gnd.n5473 gnd.n5472 585
R11706 gnd.n5472 gnd.n5341 585
R11707 gnd.n5471 gnd.n5457 585
R11708 gnd.n5471 gnd.n5333 585
R11709 gnd.n5470 gnd.n5469 585
R11710 gnd.n5470 gnd.n5330 585
R11711 gnd.n5459 gnd.n5458 585
R11712 gnd.n5458 gnd.n5321 585
R11713 gnd.n5465 gnd.n5464 585
R11714 gnd.n5464 gnd.n2822 585
R11715 gnd.n5463 gnd.n5462 585
R11716 gnd.n5463 gnd.n2820 585
R11717 gnd.n2706 gnd.n2705 585
R11718 gnd.n2745 gnd.n2706 585
R11719 gnd.n5930 gnd.n5929 585
R11720 gnd.n5929 gnd.n5928 585
R11721 gnd.n5931 gnd.n2700 585
R11722 gnd.n2700 gnd.n2698 585
R11723 gnd.n5933 gnd.n5932 585
R11724 gnd.n5934 gnd.n5933 585
R11725 gnd.n2701 gnd.n2699 585
R11726 gnd.n2699 gnd.n2683 585
R11727 gnd.n5185 gnd.n5184 585
R11728 gnd.n5186 gnd.n5185 585
R11729 gnd.n2841 gnd.n2840 585
R11730 gnd.n2840 gnd.n2839 585
R11731 gnd.n5179 gnd.n5178 585
R11732 gnd.n5178 gnd.n5177 585
R11733 gnd.n2844 gnd.n2843 585
R11734 gnd.n2845 gnd.n2844 585
R11735 gnd.n5167 gnd.n5166 585
R11736 gnd.n5168 gnd.n5167 585
R11737 gnd.n2855 gnd.n2854 585
R11738 gnd.n2854 gnd.n2852 585
R11739 gnd.n5162 gnd.n5161 585
R11740 gnd.n5161 gnd.n5160 585
R11741 gnd.n2858 gnd.n2857 585
R11742 gnd.n2865 gnd.n2858 585
R11743 gnd.n5151 gnd.n5150 585
R11744 gnd.n5152 gnd.n5151 585
R11745 gnd.n2868 gnd.n2867 585
R11746 gnd.n2867 gnd.n2864 585
R11747 gnd.n5146 gnd.n5145 585
R11748 gnd.n5145 gnd.n5144 585
R11749 gnd.n2871 gnd.n2870 585
R11750 gnd.n2878 gnd.n2871 585
R11751 gnd.n5135 gnd.n5134 585
R11752 gnd.n5136 gnd.n5135 585
R11753 gnd.n2881 gnd.n2880 585
R11754 gnd.n2888 gnd.n2880 585
R11755 gnd.n5130 gnd.n5129 585
R11756 gnd.n5129 gnd.n5128 585
R11757 gnd.n2884 gnd.n2883 585
R11758 gnd.n2963 gnd.n2884 585
R11759 gnd.n4992 gnd.n4991 585
R11760 gnd.n4993 gnd.n4992 585
R11761 gnd.n2972 gnd.n2971 585
R11762 gnd.n2979 gnd.n2971 585
R11763 gnd.n4987 gnd.n4986 585
R11764 gnd.n4986 gnd.n4985 585
R11765 gnd.n2975 gnd.n2974 585
R11766 gnd.n2983 gnd.n2975 585
R11767 gnd.n4955 gnd.n2996 585
R11768 gnd.n4913 gnd.n2996 585
R11769 gnd.n4957 gnd.n4956 585
R11770 gnd.n4958 gnd.n4957 585
R11771 gnd.n2997 gnd.n2995 585
R11772 gnd.n2995 gnd.n2992 585
R11773 gnd.n4950 gnd.n4949 585
R11774 gnd.n4949 gnd.n4948 585
R11775 gnd.n3000 gnd.n2999 585
R11776 gnd.n4940 gnd.n3000 585
R11777 gnd.n4901 gnd.n3017 585
R11778 gnd.n4818 gnd.n3017 585
R11779 gnd.n4903 gnd.n4902 585
R11780 gnd.n4904 gnd.n4903 585
R11781 gnd.n3018 gnd.n3016 585
R11782 gnd.n3025 gnd.n3016 585
R11783 gnd.n4896 gnd.n4895 585
R11784 gnd.n4895 gnd.n4894 585
R11785 gnd.n3021 gnd.n3020 585
R11786 gnd.n4880 gnd.n3021 585
R11787 gnd.n4868 gnd.n3041 585
R11788 gnd.n4814 gnd.n3041 585
R11789 gnd.n4870 gnd.n4869 585
R11790 gnd.n4871 gnd.n4870 585
R11791 gnd.n3042 gnd.n3040 585
R11792 gnd.n3050 gnd.n3040 585
R11793 gnd.n4863 gnd.n4862 585
R11794 gnd.n4862 gnd.n4861 585
R11795 gnd.n3045 gnd.n3044 585
R11796 gnd.n3055 gnd.n3045 585
R11797 gnd.n4799 gnd.n3071 585
R11798 gnd.n3071 gnd.n3062 585
R11799 gnd.n4801 gnd.n4800 585
R11800 gnd.n4802 gnd.n4801 585
R11801 gnd.n3072 gnd.n3070 585
R11802 gnd.n3070 gnd.n3066 585
R11803 gnd.n4794 gnd.n4793 585
R11804 gnd.n4793 gnd.n4792 585
R11805 gnd.n3075 gnd.n3074 585
R11806 gnd.n4784 gnd.n3075 585
R11807 gnd.n4759 gnd.n3096 585
R11808 gnd.n3096 gnd.n3095 585
R11809 gnd.n4761 gnd.n4760 585
R11810 gnd.n4762 gnd.n4761 585
R11811 gnd.n3097 gnd.n3093 585
R11812 gnd.n3103 gnd.n3093 585
R11813 gnd.n4754 gnd.n4753 585
R11814 gnd.n4753 gnd.n4752 585
R11815 gnd.n3100 gnd.n3099 585
R11816 gnd.n4739 gnd.n3100 585
R11817 gnd.n4703 gnd.n3122 585
R11818 gnd.n3122 gnd.n3114 585
R11819 gnd.n4705 gnd.n4704 585
R11820 gnd.n4706 gnd.n4705 585
R11821 gnd.n3123 gnd.n3121 585
R11822 gnd.n3121 gnd.n3118 585
R11823 gnd.n4698 gnd.n4697 585
R11824 gnd.n4697 gnd.n4696 585
R11825 gnd.n3126 gnd.n3125 585
R11826 gnd.n3132 gnd.n3126 585
R11827 gnd.n4677 gnd.n4676 585
R11828 gnd.n4678 gnd.n4677 585
R11829 gnd.n3141 gnd.n3140 585
R11830 gnd.n3148 gnd.n3140 585
R11831 gnd.n4672 gnd.n4671 585
R11832 gnd.n4671 gnd.n4670 585
R11833 gnd.n3144 gnd.n3143 585
R11834 gnd.n3152 gnd.n3144 585
R11835 gnd.n4641 gnd.n3168 585
R11836 gnd.n3168 gnd.n3159 585
R11837 gnd.n4643 gnd.n4642 585
R11838 gnd.n4644 gnd.n4643 585
R11839 gnd.n3169 gnd.n3167 585
R11840 gnd.n3167 gnd.n3164 585
R11841 gnd.n4636 gnd.n4635 585
R11842 gnd.n4635 gnd.n4634 585
R11843 gnd.n3172 gnd.n3171 585
R11844 gnd.n4626 gnd.n3172 585
R11845 gnd.n4603 gnd.n4602 585
R11846 gnd.n4602 gnd.n3179 585
R11847 gnd.n4604 gnd.n3193 585
R11848 gnd.n3193 gnd.n3185 585
R11849 gnd.n4606 gnd.n4605 585
R11850 gnd.n4607 gnd.n4606 585
R11851 gnd.n3194 gnd.n3192 585
R11852 gnd.n3498 gnd.n3192 585
R11853 gnd.n4596 gnd.n4595 585
R11854 gnd.n4595 gnd.n4594 585
R11855 gnd.n3197 gnd.n3196 585
R11856 gnd.n3494 gnd.n3197 585
R11857 gnd.n4563 gnd.n3217 585
R11858 gnd.n3217 gnd.n3208 585
R11859 gnd.n4565 gnd.n4564 585
R11860 gnd.n4566 gnd.n4565 585
R11861 gnd.n3218 gnd.n3216 585
R11862 gnd.n3216 gnd.n3212 585
R11863 gnd.n4558 gnd.n4557 585
R11864 gnd.n4557 gnd.n4556 585
R11865 gnd.n3221 gnd.n3220 585
R11866 gnd.n3281 gnd.n3221 585
R11867 gnd.n3481 gnd.n3438 585
R11868 gnd.n3438 gnd.n3248 585
R11869 gnd.n3483 gnd.n3482 585
R11870 gnd.n3484 gnd.n3483 585
R11871 gnd.n3439 gnd.n3437 585
R11872 gnd.n3473 gnd.n3437 585
R11873 gnd.n3476 gnd.n3475 585
R11874 gnd.n3475 gnd.n3474 585
R11875 gnd.n3442 gnd.n3441 585
R11876 gnd.n3471 gnd.n3442 585
R11877 gnd.n3469 gnd.n3468 585
R11878 gnd.n3470 gnd.n3469 585
R11879 gnd.n3445 gnd.n3444 585
R11880 gnd.n3461 gnd.n3444 585
R11881 gnd.n3464 gnd.n3463 585
R11882 gnd.n3463 gnd.n3462 585
R11883 gnd.n3448 gnd.n3447 585
R11884 gnd.n3459 gnd.n3448 585
R11885 gnd.n3457 gnd.n3456 585
R11886 gnd.n3458 gnd.n3457 585
R11887 gnd.n3452 gnd.n3451 585
R11888 gnd.n3451 gnd.n3449 585
R11889 gnd.n2572 gnd.n2571 585
R11890 gnd.n6062 gnd.n2572 585
R11891 gnd.n6065 gnd.n6064 585
R11892 gnd.n6064 gnd.n6063 585
R11893 gnd.n6066 gnd.n2566 585
R11894 gnd.n2566 gnd.n2564 585
R11895 gnd.n6068 gnd.n6067 585
R11896 gnd.n6069 gnd.n6068 585
R11897 gnd.n2567 gnd.n2565 585
R11898 gnd.n2565 gnd.n2549 585
R11899 gnd.n4278 gnd.n4277 585
R11900 gnd.n4279 gnd.n4278 585
R11901 gnd.n3673 gnd.n3672 585
R11902 gnd.n3672 gnd.n3366 585
R11903 gnd.n4272 gnd.n4271 585
R11904 gnd.n4271 gnd.n2535 585
R11905 gnd.n4270 gnd.n3675 585
R11906 gnd.n4270 gnd.n2532 585
R11907 gnd.n4269 gnd.n4268 585
R11908 gnd.n4269 gnd.n2540 585
R11909 gnd.n3677 gnd.n3676 585
R11910 gnd.n3676 gnd.n2523 585
R11911 gnd.n4264 gnd.n4263 585
R11912 gnd.n4263 gnd.n2516 585
R11913 gnd.n4262 gnd.n3679 585
R11914 gnd.n4262 gnd.n2513 585
R11915 gnd.n4261 gnd.n4260 585
R11916 gnd.n4261 gnd.n2505 585
R11917 gnd.n3681 gnd.n3680 585
R11918 gnd.n3680 gnd.n2502 585
R11919 gnd.n4256 gnd.n4255 585
R11920 gnd.n4255 gnd.n2495 585
R11921 gnd.n4254 gnd.n3683 585
R11922 gnd.n4254 gnd.n2492 585
R11923 gnd.n4253 gnd.n4252 585
R11924 gnd.n4253 gnd.n2484 585
R11925 gnd.n3685 gnd.n3684 585
R11926 gnd.n3684 gnd.n2481 585
R11927 gnd.n4248 gnd.n4247 585
R11928 gnd.n4247 gnd.n4246 585
R11929 gnd.n3688 gnd.n3687 585
R11930 gnd.n3688 gnd.n2472 585
R11931 gnd.n3774 gnd.n3773 585
R11932 gnd.n3774 gnd.n2464 585
R11933 gnd.n3776 gnd.n3775 585
R11934 gnd.n3775 gnd.n2461 585
R11935 gnd.n3777 gnd.n3770 585
R11936 gnd.n3770 gnd.n2454 585
R11937 gnd.n3779 gnd.n3778 585
R11938 gnd.n3779 gnd.n2451 585
R11939 gnd.n3781 gnd.n3780 585
R11940 gnd.n3780 gnd.n2446 585
R11941 gnd.n3783 gnd.n3782 585
R11942 gnd.n3783 gnd.n2443 585
R11943 gnd.n3785 gnd.n3784 585
R11944 gnd.n3784 gnd.n3709 585
R11945 gnd.n3787 gnd.n3786 585
R11946 gnd.n3787 gnd.n2434 585
R11947 gnd.n3789 gnd.n3788 585
R11948 gnd.n3789 gnd.n2429 585
R11949 gnd.n3790 gnd.n3768 585
R11950 gnd.n3790 gnd.n2426 585
R11951 gnd.n3792 gnd.n3791 585
R11952 gnd.n3791 gnd.n2419 585
R11953 gnd.n3769 gnd.n3763 585
R11954 gnd.n3769 gnd.n2416 585
R11955 gnd.n3796 gnd.n3762 585
R11956 gnd.n3762 gnd.n2410 585
R11957 gnd.n3797 gnd.n3758 585
R11958 gnd.n3758 gnd.n2407 585
R11959 gnd.n3799 gnd.n3798 585
R11960 gnd.n3799 gnd.n3720 585
R11961 gnd.n3800 gnd.n3757 585
R11962 gnd.n3800 gnd.n2398 585
R11963 gnd.n3802 gnd.n3801 585
R11964 gnd.n3801 gnd.n2390 585
R11965 gnd.n3803 gnd.n3752 585
R11966 gnd.n3752 gnd.n2387 585
R11967 gnd.n3805 gnd.n3804 585
R11968 gnd.n3805 gnd.n2380 585
R11969 gnd.n3806 gnd.n3751 585
R11970 gnd.n3806 gnd.n2377 585
R11971 gnd.n3808 gnd.n3807 585
R11972 gnd.n3807 gnd.n2369 585
R11973 gnd.n3809 gnd.n3732 585
R11974 gnd.n3732 gnd.n2366 585
R11975 gnd.n3811 gnd.n3810 585
R11976 gnd.n3812 gnd.n3811 585
R11977 gnd.n3733 gnd.n3731 585
R11978 gnd.n3731 gnd.n2357 585
R11979 gnd.n3745 gnd.n3744 585
R11980 gnd.n3744 gnd.n2349 585
R11981 gnd.n3743 gnd.n3735 585
R11982 gnd.n3743 gnd.n2346 585
R11983 gnd.n3742 gnd.n3741 585
R11984 gnd.n3742 gnd.n2337 585
R11985 gnd.n3737 gnd.n3736 585
R11986 gnd.n3736 gnd.n2334 585
R11987 gnd.n2321 gnd.n2320 585
R11988 gnd.n2325 gnd.n2321 585
R11989 gnd.n6218 gnd.n6217 585
R11990 gnd.n6217 gnd.n6216 585
R11991 gnd.n6219 gnd.n2315 585
R11992 gnd.n2322 gnd.n2315 585
R11993 gnd.n6221 gnd.n6220 585
R11994 gnd.n6222 gnd.n6221 585
R11995 gnd.n2313 gnd.n2312 585
R11996 gnd.n6223 gnd.n2313 585
R11997 gnd.n6226 gnd.n6225 585
R11998 gnd.n6225 gnd.n6224 585
R11999 gnd.n6227 gnd.n2306 585
R12000 gnd.n2306 gnd.n2305 585
R12001 gnd.n6229 gnd.n6228 585
R12002 gnd.n6230 gnd.n6229 585
R12003 gnd.n2307 gnd.n841 585
R12004 gnd.n6231 gnd.n841 585
R12005 gnd.n5187 gnd.n2838 585
R12006 gnd.n5187 gnd.n5186 585
R12007 gnd.n2848 gnd.n2837 585
R12008 gnd.n2839 gnd.n2837 585
R12009 gnd.n5176 gnd.n5175 585
R12010 gnd.n5177 gnd.n5176 585
R12011 gnd.n2847 gnd.n2846 585
R12012 gnd.n2846 gnd.n2845 585
R12013 gnd.n5170 gnd.n5169 585
R12014 gnd.n5169 gnd.n5168 585
R12015 gnd.n2851 gnd.n2850 585
R12016 gnd.n2852 gnd.n2851 585
R12017 gnd.n5159 gnd.n5158 585
R12018 gnd.n5160 gnd.n5159 585
R12019 gnd.n2860 gnd.n2859 585
R12020 gnd.n2865 gnd.n2859 585
R12021 gnd.n5154 gnd.n5153 585
R12022 gnd.n5153 gnd.n5152 585
R12023 gnd.n2863 gnd.n2862 585
R12024 gnd.n2864 gnd.n2863 585
R12025 gnd.n5143 gnd.n5142 585
R12026 gnd.n5144 gnd.n5143 585
R12027 gnd.n2873 gnd.n2872 585
R12028 gnd.n2878 gnd.n2872 585
R12029 gnd.n5138 gnd.n5137 585
R12030 gnd.n5137 gnd.n5136 585
R12031 gnd.n2876 gnd.n2875 585
R12032 gnd.n2888 gnd.n2876 585
R12033 gnd.n4921 gnd.n2886 585
R12034 gnd.n5128 gnd.n2886 585
R12035 gnd.n4920 gnd.n4919 585
R12036 gnd.n4919 gnd.n2963 585
R12037 gnd.n4925 gnd.n2968 585
R12038 gnd.n4993 gnd.n2968 585
R12039 gnd.n4926 gnd.n4918 585
R12040 gnd.n4918 gnd.n2979 585
R12041 gnd.n4927 gnd.n2977 585
R12042 gnd.n4985 gnd.n2977 585
R12043 gnd.n4916 gnd.n4915 585
R12044 gnd.n4915 gnd.n2983 585
R12045 gnd.n4931 gnd.n4914 585
R12046 gnd.n4914 gnd.n4913 585
R12047 gnd.n4932 gnd.n2994 585
R12048 gnd.n4958 gnd.n2994 585
R12049 gnd.n4933 gnd.n4910 585
R12050 gnd.n4910 gnd.n2992 585
R12051 gnd.n3011 gnd.n3002 585
R12052 gnd.n4948 gnd.n3002 585
R12053 gnd.n4938 gnd.n4937 585
R12054 gnd.n4940 gnd.n4938 585
R12055 gnd.n3010 gnd.n3009 585
R12056 gnd.n4818 gnd.n3009 585
R12057 gnd.n4906 gnd.n4905 585
R12058 gnd.n4905 gnd.n4904 585
R12059 gnd.n3014 gnd.n3013 585
R12060 gnd.n3025 gnd.n3014 585
R12061 gnd.n3034 gnd.n3023 585
R12062 gnd.n4894 gnd.n3023 585
R12063 gnd.n4879 gnd.n4878 585
R12064 gnd.n4880 gnd.n4879 585
R12065 gnd.n3033 gnd.n3032 585
R12066 gnd.n4814 gnd.n3032 585
R12067 gnd.n4873 gnd.n4872 585
R12068 gnd.n4872 gnd.n4871 585
R12069 gnd.n3037 gnd.n3036 585
R12070 gnd.n3050 gnd.n3037 585
R12071 gnd.n4772 gnd.n3047 585
R12072 gnd.n4861 gnd.n3047 585
R12073 gnd.n4771 gnd.n4770 585
R12074 gnd.n4770 gnd.n3055 585
R12075 gnd.n4776 gnd.n4769 585
R12076 gnd.n4769 gnd.n3062 585
R12077 gnd.n4777 gnd.n3068 585
R12078 gnd.n4802 gnd.n3068 585
R12079 gnd.n4778 gnd.n4768 585
R12080 gnd.n4768 gnd.n3066 585
R12081 gnd.n3087 gnd.n3077 585
R12082 gnd.n4792 gnd.n3077 585
R12083 gnd.n4783 gnd.n4782 585
R12084 gnd.n4784 gnd.n4783 585
R12085 gnd.n3086 gnd.n3085 585
R12086 gnd.n3095 gnd.n3085 585
R12087 gnd.n4764 gnd.n4763 585
R12088 gnd.n4763 gnd.n4762 585
R12089 gnd.n3090 gnd.n3089 585
R12090 gnd.n3103 gnd.n3090 585
R12091 gnd.n3517 gnd.n3101 585
R12092 gnd.n4752 gnd.n3101 585
R12093 gnd.n3520 gnd.n3111 585
R12094 gnd.n4739 gnd.n3111 585
R12095 gnd.n3521 gnd.n3516 585
R12096 gnd.n3516 gnd.n3114 585
R12097 gnd.n3522 gnd.n3120 585
R12098 gnd.n4706 gnd.n3120 585
R12099 gnd.n3514 gnd.n3513 585
R12100 gnd.n3513 gnd.n3118 585
R12101 gnd.n3526 gnd.n3128 585
R12102 gnd.n4696 gnd.n3128 585
R12103 gnd.n3527 gnd.n3512 585
R12104 gnd.n3512 gnd.n3132 585
R12105 gnd.n3528 gnd.n3138 585
R12106 gnd.n4678 gnd.n3138 585
R12107 gnd.n3510 gnd.n3509 585
R12108 gnd.n3509 gnd.n3148 585
R12109 gnd.n3532 gnd.n3146 585
R12110 gnd.n4670 gnd.n3146 585
R12111 gnd.n3533 gnd.n3508 585
R12112 gnd.n3508 gnd.n3152 585
R12113 gnd.n3534 gnd.n3507 585
R12114 gnd.n3507 gnd.n3159 585
R12115 gnd.n3505 gnd.n3166 585
R12116 gnd.n4644 gnd.n3166 585
R12117 gnd.n3538 gnd.n3504 585
R12118 gnd.n3504 gnd.n3164 585
R12119 gnd.n3539 gnd.n3173 585
R12120 gnd.n4634 gnd.n3173 585
R12121 gnd.n3540 gnd.n3181 585
R12122 gnd.n4626 gnd.n3181 585
R12123 gnd.n3502 gnd.n3501 585
R12124 gnd.n3501 gnd.n3179 585
R12125 gnd.n3544 gnd.n3500 585
R12126 gnd.n3500 gnd.n3185 585
R12127 gnd.n3545 gnd.n3191 585
R12128 gnd.n4607 gnd.n3191 585
R12129 gnd.n3546 gnd.n3499 585
R12130 gnd.n3499 gnd.n3498 585
R12131 gnd.n3496 gnd.n3199 585
R12132 gnd.n4594 gnd.n3199 585
R12133 gnd.n3550 gnd.n3495 585
R12134 gnd.n3495 gnd.n3494 585
R12135 gnd.n3551 gnd.n3491 585
R12136 gnd.n3491 gnd.n3208 585
R12137 gnd.n3552 gnd.n3214 585
R12138 gnd.n4566 gnd.n3214 585
R12139 gnd.n3489 gnd.n3488 585
R12140 gnd.n3488 gnd.n3212 585
R12141 gnd.n3556 gnd.n3223 585
R12142 gnd.n4556 gnd.n3223 585
R12143 gnd.n3557 gnd.n3487 585
R12144 gnd.n3487 gnd.n3281 585
R12145 gnd.n3558 gnd.n3486 585
R12146 gnd.n3486 gnd.n3248 585
R12147 gnd.n3485 gnd.n3435 585
R12148 gnd.n3485 gnd.n3484 585
R12149 gnd.n3562 gnd.n3434 585
R12150 gnd.n3473 gnd.n3434 585
R12151 gnd.n3563 gnd.n3433 585
R12152 gnd.n3474 gnd.n3433 585
R12153 gnd.n3564 gnd.n3432 585
R12154 gnd.n3471 gnd.n3432 585
R12155 gnd.n3443 gnd.n3430 585
R12156 gnd.n3470 gnd.n3443 585
R12157 gnd.n3568 gnd.n3429 585
R12158 gnd.n3461 gnd.n3429 585
R12159 gnd.n3569 gnd.n3428 585
R12160 gnd.n3462 gnd.n3428 585
R12161 gnd.n3570 gnd.n3427 585
R12162 gnd.n3459 gnd.n3427 585
R12163 gnd.n3450 gnd.n3425 585
R12164 gnd.n3458 gnd.n3450 585
R12165 gnd.n3574 gnd.n3424 585
R12166 gnd.n3449 gnd.n3424 585
R12167 gnd.n3575 gnd.n2574 585
R12168 gnd.n6062 gnd.n2574 585
R12169 gnd.n3576 gnd.n2573 585
R12170 gnd.n6063 gnd.n2573 585
R12171 gnd.n3579 gnd.n3578 585
R12172 gnd.n3421 gnd.n3420 585
R12173 gnd.n3583 gnd.n3422 585
R12174 gnd.n3585 gnd.n3584 585
R12175 gnd.n3587 gnd.n3586 585
R12176 gnd.n3417 gnd.n3416 585
R12177 gnd.n3591 gnd.n3418 585
R12178 gnd.n3594 gnd.n3593 585
R12179 gnd.n3592 gnd.n3414 585
R12180 gnd.n3601 gnd.n3600 585
R12181 gnd.n3603 gnd.n3602 585
R12182 gnd.n3408 gnd.n3407 585
R12183 gnd.n3612 gnd.n3409 585
R12184 gnd.n3615 gnd.n3614 585
R12185 gnd.n3613 gnd.n3401 585
R12186 gnd.n3625 gnd.n3624 585
R12187 gnd.n3627 gnd.n3626 585
R12188 gnd.n3396 gnd.n3395 585
R12189 gnd.n3636 gnd.n3397 585
R12190 gnd.n3639 gnd.n3638 585
R12191 gnd.n3637 gnd.n3389 585
R12192 gnd.n3649 gnd.n3648 585
R12193 gnd.n3651 gnd.n3650 585
R12194 gnd.n3384 gnd.n3383 585
R12195 gnd.n3660 gnd.n3385 585
R12196 gnd.n3664 gnd.n3663 585
R12197 gnd.n3662 gnd.n2546 585
R12198 gnd.n6072 gnd.n2547 585
R12199 gnd.n6071 gnd.n6070 585
R12200 gnd.n6070 gnd.n6069 585
R12201 gnd.n2682 gnd.n2678 585
R12202 gnd.n5186 gnd.n2682 585
R12203 gnd.n5940 gnd.n2677 585
R12204 gnd.n2839 gnd.n2677 585
R12205 gnd.n5941 gnd.n2676 585
R12206 gnd.n5177 gnd.n2676 585
R12207 gnd.n5942 gnd.n2675 585
R12208 gnd.n2845 gnd.n2675 585
R12209 gnd.n2853 gnd.n2673 585
R12210 gnd.n5168 gnd.n2853 585
R12211 gnd.n5946 gnd.n2672 585
R12212 gnd.n2852 gnd.n2672 585
R12213 gnd.n5947 gnd.n2671 585
R12214 gnd.n5160 gnd.n2671 585
R12215 gnd.n5948 gnd.n2670 585
R12216 gnd.n2865 gnd.n2670 585
R12217 gnd.n2866 gnd.n2668 585
R12218 gnd.n5152 gnd.n2866 585
R12219 gnd.n5952 gnd.n2667 585
R12220 gnd.n2864 gnd.n2667 585
R12221 gnd.n5953 gnd.n2666 585
R12222 gnd.n5144 gnd.n2666 585
R12223 gnd.n5954 gnd.n2665 585
R12224 gnd.n2878 gnd.n2665 585
R12225 gnd.n2879 gnd.n2663 585
R12226 gnd.n5136 gnd.n2879 585
R12227 gnd.n5958 gnd.n2662 585
R12228 gnd.n2888 gnd.n2662 585
R12229 gnd.n5959 gnd.n2661 585
R12230 gnd.n5128 gnd.n2661 585
R12231 gnd.n5960 gnd.n2660 585
R12232 gnd.n2963 gnd.n2660 585
R12233 gnd.n2970 gnd.n2658 585
R12234 gnd.n4993 gnd.n2970 585
R12235 gnd.n5964 gnd.n2657 585
R12236 gnd.n2979 gnd.n2657 585
R12237 gnd.n5965 gnd.n2656 585
R12238 gnd.n4985 gnd.n2656 585
R12239 gnd.n5966 gnd.n2655 585
R12240 gnd.n2983 gnd.n2655 585
R12241 gnd.n4912 gnd.n2653 585
R12242 gnd.n4913 gnd.n4912 585
R12243 gnd.n5970 gnd.n2652 585
R12244 gnd.n4958 gnd.n2652 585
R12245 gnd.n5971 gnd.n2651 585
R12246 gnd.n2992 gnd.n2651 585
R12247 gnd.n5972 gnd.n2650 585
R12248 gnd.n4948 gnd.n2650 585
R12249 gnd.n4939 gnd.n2648 585
R12250 gnd.n4940 gnd.n4939 585
R12251 gnd.n5976 gnd.n2647 585
R12252 gnd.n4818 gnd.n2647 585
R12253 gnd.n5977 gnd.n2646 585
R12254 gnd.n4904 gnd.n2646 585
R12255 gnd.n5978 gnd.n2645 585
R12256 gnd.n3025 gnd.n2645 585
R12257 gnd.n4893 gnd.n2643 585
R12258 gnd.n4894 gnd.n4893 585
R12259 gnd.n5982 gnd.n2642 585
R12260 gnd.n4880 gnd.n2642 585
R12261 gnd.n5983 gnd.n2641 585
R12262 gnd.n4814 gnd.n2641 585
R12263 gnd.n5984 gnd.n2640 585
R12264 gnd.n4871 gnd.n2640 585
R12265 gnd.n3049 gnd.n2638 585
R12266 gnd.n3050 gnd.n3049 585
R12267 gnd.n5988 gnd.n2637 585
R12268 gnd.n4861 gnd.n2637 585
R12269 gnd.n5989 gnd.n2636 585
R12270 gnd.n3055 gnd.n2636 585
R12271 gnd.n5990 gnd.n2635 585
R12272 gnd.n3062 gnd.n2635 585
R12273 gnd.n3069 gnd.n2633 585
R12274 gnd.n4802 gnd.n3069 585
R12275 gnd.n5994 gnd.n2632 585
R12276 gnd.n3066 gnd.n2632 585
R12277 gnd.n5995 gnd.n2631 585
R12278 gnd.n4792 gnd.n2631 585
R12279 gnd.n5996 gnd.n2630 585
R12280 gnd.n4784 gnd.n2630 585
R12281 gnd.n3094 gnd.n2628 585
R12282 gnd.n3095 gnd.n3094 585
R12283 gnd.n6000 gnd.n2627 585
R12284 gnd.n4762 gnd.n2627 585
R12285 gnd.n6001 gnd.n2626 585
R12286 gnd.n3103 gnd.n2626 585
R12287 gnd.n6002 gnd.n2625 585
R12288 gnd.n4752 gnd.n2625 585
R12289 gnd.n4738 gnd.n2623 585
R12290 gnd.n4739 gnd.n4738 585
R12291 gnd.n6006 gnd.n2622 585
R12292 gnd.n3114 gnd.n2622 585
R12293 gnd.n6007 gnd.n2621 585
R12294 gnd.n4706 gnd.n2621 585
R12295 gnd.n6008 gnd.n2620 585
R12296 gnd.n3118 gnd.n2620 585
R12297 gnd.n4695 gnd.n2618 585
R12298 gnd.n4696 gnd.n4695 585
R12299 gnd.n6012 gnd.n2617 585
R12300 gnd.n3132 gnd.n2617 585
R12301 gnd.n6013 gnd.n2616 585
R12302 gnd.n4678 gnd.n2616 585
R12303 gnd.n6014 gnd.n2615 585
R12304 gnd.n3148 gnd.n2615 585
R12305 gnd.n4669 gnd.n2613 585
R12306 gnd.n4670 gnd.n4669 585
R12307 gnd.n6018 gnd.n2612 585
R12308 gnd.n3152 gnd.n2612 585
R12309 gnd.n6019 gnd.n2611 585
R12310 gnd.n3159 gnd.n2611 585
R12311 gnd.n6020 gnd.n2610 585
R12312 gnd.n4644 gnd.n2610 585
R12313 gnd.n3163 gnd.n2608 585
R12314 gnd.n3164 gnd.n3163 585
R12315 gnd.n6024 gnd.n2607 585
R12316 gnd.n4634 gnd.n2607 585
R12317 gnd.n6025 gnd.n2606 585
R12318 gnd.n4626 gnd.n2606 585
R12319 gnd.n6026 gnd.n2605 585
R12320 gnd.n3179 gnd.n2605 585
R12321 gnd.n3184 gnd.n2603 585
R12322 gnd.n3185 gnd.n3184 585
R12323 gnd.n6030 gnd.n2602 585
R12324 gnd.n4607 gnd.n2602 585
R12325 gnd.n6031 gnd.n2601 585
R12326 gnd.n3498 gnd.n2601 585
R12327 gnd.n6032 gnd.n2600 585
R12328 gnd.n4594 gnd.n2600 585
R12329 gnd.n3493 gnd.n2598 585
R12330 gnd.n3494 gnd.n3493 585
R12331 gnd.n6036 gnd.n2597 585
R12332 gnd.n3208 gnd.n2597 585
R12333 gnd.n6037 gnd.n2596 585
R12334 gnd.n4566 gnd.n2596 585
R12335 gnd.n6038 gnd.n2595 585
R12336 gnd.n3212 gnd.n2595 585
R12337 gnd.n4555 gnd.n2593 585
R12338 gnd.n4556 gnd.n4555 585
R12339 gnd.n6042 gnd.n2592 585
R12340 gnd.n3281 gnd.n2592 585
R12341 gnd.n6043 gnd.n2591 585
R12342 gnd.n3248 gnd.n2591 585
R12343 gnd.n6044 gnd.n2590 585
R12344 gnd.n3484 gnd.n2590 585
R12345 gnd.n3472 gnd.n2588 585
R12346 gnd.n3473 gnd.n3472 585
R12347 gnd.n6048 gnd.n2587 585
R12348 gnd.n3474 gnd.n2587 585
R12349 gnd.n6049 gnd.n2586 585
R12350 gnd.n3471 gnd.n2586 585
R12351 gnd.n6050 gnd.n2585 585
R12352 gnd.n3470 gnd.n2585 585
R12353 gnd.n3460 gnd.n2583 585
R12354 gnd.n3461 gnd.n3460 585
R12355 gnd.n6054 gnd.n2582 585
R12356 gnd.n3462 gnd.n2582 585
R12357 gnd.n6055 gnd.n2581 585
R12358 gnd.n3459 gnd.n2581 585
R12359 gnd.n6056 gnd.n2580 585
R12360 gnd.n3458 gnd.n2580 585
R12361 gnd.n2577 gnd.n2575 585
R12362 gnd.n3449 gnd.n2575 585
R12363 gnd.n6061 gnd.n6060 585
R12364 gnd.n6062 gnd.n6061 585
R12365 gnd.n2576 gnd.n2548 585
R12366 gnd.n6063 gnd.n2548 585
R12367 gnd.n5253 gnd.n5252 585
R12368 gnd.n5279 gnd.n5251 585
R12369 gnd.n5280 gnd.n5250 585
R12370 gnd.n5249 gnd.n5241 585
R12371 gnd.n5287 gnd.n5240 585
R12372 gnd.n5288 gnd.n5239 585
R12373 gnd.n5233 gnd.n5232 585
R12374 gnd.n5295 gnd.n5231 585
R12375 gnd.n5296 gnd.n5230 585
R12376 gnd.n5229 gnd.n5221 585
R12377 gnd.n5303 gnd.n5220 585
R12378 gnd.n5304 gnd.n5219 585
R12379 gnd.n5213 gnd.n5212 585
R12380 gnd.n5311 gnd.n5211 585
R12381 gnd.n5312 gnd.n5210 585
R12382 gnd.n5209 gnd.n5208 585
R12383 gnd.n5207 gnd.n5204 585
R12384 gnd.n5203 gnd.n5202 585
R12385 gnd.n5201 gnd.n2831 585
R12386 gnd.n2830 gnd.n2829 585
R12387 gnd.n5197 gnd.n5196 585
R12388 gnd.n5195 gnd.n5194 585
R12389 gnd.n5193 gnd.n2835 585
R12390 gnd.n2834 gnd.n2833 585
R12391 gnd.n5189 gnd.n5188 585
R12392 gnd.n5936 gnd.n5935 585
R12393 gnd.n5935 gnd.n5934 585
R12394 gnd.n2681 gnd.n2680 585
R12395 gnd.n5271 gnd.n5266 585
R12396 gnd.n5272 gnd.n5265 585
R12397 gnd.n5126 gnd.n2890 511.721
R12398 gnd.n5006 gnd.n2887 511.721
R12399 gnd.n3295 gnd.n3294 511.721
R12400 gnd.n4548 gnd.n3225 511.721
R12401 gnd.n6400 gnd.n670 508.505
R12402 gnd.n3286 gnd.t251 389.64
R12403 gnd.n2938 gnd.t207 389.64
R12404 gnd.n3283 gnd.t171 389.64
R12405 gnd.n2932 gnd.t257 389.64
R12406 gnd.n3381 gnd.t241 371.625
R12407 gnd.n5258 gnd.t269 371.625
R12408 gnd.n3378 gnd.t281 371.625
R12409 gnd.n2767 gnd.t266 371.625
R12410 gnd.n2790 gnd.t254 371.625
R12411 gnd.n2812 gnd.t197 371.625
R12412 gnd.n7209 gnd.t201 371.625
R12413 gnd.n7188 gnd.t193 371.625
R12414 gnd.n7295 gnd.t260 371.625
R12415 gnd.n178 gnd.t275 371.625
R12416 gnd.n3939 gnd.t232 371.625
R12417 gnd.n4050 gnd.t211 371.625
R12418 gnd.n3895 gnd.t235 371.625
R12419 gnd.n3855 gnd.t189 371.625
R12420 gnd.n4315 gnd.t272 371.625
R12421 gnd.n4418 gnd.t218 371.625
R12422 gnd.n4385 gnd.t238 371.625
R12423 gnd.n5262 gnd.t222 371.625
R12424 gnd.n7101 gnd.n7100 368.44
R12425 gnd.n1322 gnd.t284 323.425
R12426 gnd.n881 gnd.t179 323.425
R12427 gnd.n6891 gnd.n377 301.784
R12428 gnd.n6899 gnd.n377 301.784
R12429 gnd.n6900 gnd.n6899 301.784
R12430 gnd.n6901 gnd.n6900 301.784
R12431 gnd.n6901 gnd.n371 301.784
R12432 gnd.n6909 gnd.n371 301.784
R12433 gnd.n6910 gnd.n6909 301.784
R12434 gnd.n6911 gnd.n6910 301.784
R12435 gnd.n6911 gnd.n365 301.784
R12436 gnd.n6919 gnd.n365 301.784
R12437 gnd.n6920 gnd.n6919 301.784
R12438 gnd.n6921 gnd.n6920 301.784
R12439 gnd.n6921 gnd.n359 301.784
R12440 gnd.n6929 gnd.n359 301.784
R12441 gnd.n6930 gnd.n6929 301.784
R12442 gnd.n6931 gnd.n6930 301.784
R12443 gnd.n6931 gnd.n353 301.784
R12444 gnd.n6939 gnd.n353 301.784
R12445 gnd.n6940 gnd.n6939 301.784
R12446 gnd.n6941 gnd.n6940 301.784
R12447 gnd.n6941 gnd.n347 301.784
R12448 gnd.n6949 gnd.n347 301.784
R12449 gnd.n6950 gnd.n6949 301.784
R12450 gnd.n6951 gnd.n6950 301.784
R12451 gnd.n6951 gnd.n341 301.784
R12452 gnd.n6959 gnd.n341 301.784
R12453 gnd.n6960 gnd.n6959 301.784
R12454 gnd.n6961 gnd.n6960 301.784
R12455 gnd.n6961 gnd.n335 301.784
R12456 gnd.n6969 gnd.n335 301.784
R12457 gnd.n6970 gnd.n6969 301.784
R12458 gnd.n6971 gnd.n6970 301.784
R12459 gnd.n6971 gnd.n329 301.784
R12460 gnd.n6979 gnd.n329 301.784
R12461 gnd.n6980 gnd.n6979 301.784
R12462 gnd.n6981 gnd.n6980 301.784
R12463 gnd.n6981 gnd.n323 301.784
R12464 gnd.n6989 gnd.n323 301.784
R12465 gnd.n6990 gnd.n6989 301.784
R12466 gnd.n6991 gnd.n6990 301.784
R12467 gnd.n6991 gnd.n317 301.784
R12468 gnd.n6999 gnd.n317 301.784
R12469 gnd.n7000 gnd.n6999 301.784
R12470 gnd.n7001 gnd.n7000 301.784
R12471 gnd.n7001 gnd.n311 301.784
R12472 gnd.n7009 gnd.n311 301.784
R12473 gnd.n7010 gnd.n7009 301.784
R12474 gnd.n7011 gnd.n7010 301.784
R12475 gnd.n7011 gnd.n305 301.784
R12476 gnd.n7019 gnd.n305 301.784
R12477 gnd.n7020 gnd.n7019 301.784
R12478 gnd.n7021 gnd.n7020 301.784
R12479 gnd.n7021 gnd.n299 301.784
R12480 gnd.n7029 gnd.n299 301.784
R12481 gnd.n7030 gnd.n7029 301.784
R12482 gnd.n7031 gnd.n7030 301.784
R12483 gnd.n7031 gnd.n293 301.784
R12484 gnd.n7039 gnd.n293 301.784
R12485 gnd.n7040 gnd.n7039 301.784
R12486 gnd.n7041 gnd.n7040 301.784
R12487 gnd.n7041 gnd.n287 301.784
R12488 gnd.n7049 gnd.n287 301.784
R12489 gnd.n7050 gnd.n7049 301.784
R12490 gnd.n7051 gnd.n7050 301.784
R12491 gnd.n7051 gnd.n281 301.784
R12492 gnd.n7059 gnd.n281 301.784
R12493 gnd.n7060 gnd.n7059 301.784
R12494 gnd.n7061 gnd.n7060 301.784
R12495 gnd.n7061 gnd.n275 301.784
R12496 gnd.n7069 gnd.n275 301.784
R12497 gnd.n7070 gnd.n7069 301.784
R12498 gnd.n7071 gnd.n7070 301.784
R12499 gnd.n7071 gnd.n269 301.784
R12500 gnd.n7079 gnd.n269 301.784
R12501 gnd.n7080 gnd.n7079 301.784
R12502 gnd.n7081 gnd.n7080 301.784
R12503 gnd.n7081 gnd.n263 301.784
R12504 gnd.n7089 gnd.n263 301.784
R12505 gnd.n7090 gnd.n7089 301.784
R12506 gnd.n7091 gnd.n7090 301.784
R12507 gnd.n7091 gnd.n257 301.784
R12508 gnd.n7099 gnd.n257 301.784
R12509 gnd.n7100 gnd.n7099 301.784
R12510 gnd.n2172 gnd.n2146 289.615
R12511 gnd.n2140 gnd.n2114 289.615
R12512 gnd.n2108 gnd.n2082 289.615
R12513 gnd.n2077 gnd.n2051 289.615
R12514 gnd.n2045 gnd.n2019 289.615
R12515 gnd.n2013 gnd.n1987 289.615
R12516 gnd.n1981 gnd.n1955 289.615
R12517 gnd.n1950 gnd.n1924 289.615
R12518 gnd.n1396 gnd.t175 279.217
R12519 gnd.n907 gnd.t214 279.217
R12520 gnd.n3232 gnd.t188 260.649
R12521 gnd.n2903 gnd.t228 260.649
R12522 gnd.n4547 gnd.n4546 256.663
R12523 gnd.n4546 gnd.n3249 256.663
R12524 gnd.n4546 gnd.n3250 256.663
R12525 gnd.n4546 gnd.n3251 256.663
R12526 gnd.n4546 gnd.n3252 256.663
R12527 gnd.n4546 gnd.n3253 256.663
R12528 gnd.n4546 gnd.n3254 256.663
R12529 gnd.n4546 gnd.n3255 256.663
R12530 gnd.n4546 gnd.n3256 256.663
R12531 gnd.n4546 gnd.n3257 256.663
R12532 gnd.n4546 gnd.n3258 256.663
R12533 gnd.n4546 gnd.n3259 256.663
R12534 gnd.n4546 gnd.n3260 256.663
R12535 gnd.n4546 gnd.n3261 256.663
R12536 gnd.n4546 gnd.n3262 256.663
R12537 gnd.n4546 gnd.n3263 256.663
R12538 gnd.n4486 gnd.n4483 256.663
R12539 gnd.n4546 gnd.n3264 256.663
R12540 gnd.n4546 gnd.n3265 256.663
R12541 gnd.n4546 gnd.n3266 256.663
R12542 gnd.n4546 gnd.n3267 256.663
R12543 gnd.n4546 gnd.n3268 256.663
R12544 gnd.n4546 gnd.n3269 256.663
R12545 gnd.n4546 gnd.n3270 256.663
R12546 gnd.n4546 gnd.n3271 256.663
R12547 gnd.n4546 gnd.n3272 256.663
R12548 gnd.n4546 gnd.n3273 256.663
R12549 gnd.n4546 gnd.n3274 256.663
R12550 gnd.n4546 gnd.n3275 256.663
R12551 gnd.n4546 gnd.n3276 256.663
R12552 gnd.n4546 gnd.n3277 256.663
R12553 gnd.n4546 gnd.n3278 256.663
R12554 gnd.n4546 gnd.n3279 256.663
R12555 gnd.n4546 gnd.n3280 256.663
R12556 gnd.n5005 gnd.n2877 256.663
R12557 gnd.n5011 gnd.n2877 256.663
R12558 gnd.n2959 gnd.n2877 256.663
R12559 gnd.n5018 gnd.n2877 256.663
R12560 gnd.n2956 gnd.n2877 256.663
R12561 gnd.n5025 gnd.n2877 256.663
R12562 gnd.n2953 gnd.n2877 256.663
R12563 gnd.n5032 gnd.n2877 256.663
R12564 gnd.n2950 gnd.n2877 256.663
R12565 gnd.n5039 gnd.n2877 256.663
R12566 gnd.n2947 gnd.n2877 256.663
R12567 gnd.n5046 gnd.n2877 256.663
R12568 gnd.n2944 gnd.n2877 256.663
R12569 gnd.n5053 gnd.n2877 256.663
R12570 gnd.n2941 gnd.n2877 256.663
R12571 gnd.n5061 gnd.n2877 256.663
R12572 gnd.n5064 gnd.n2777 256.663
R12573 gnd.n5065 gnd.n2877 256.663
R12574 gnd.n5069 gnd.n2877 256.663
R12575 gnd.n2935 gnd.n2877 256.663
R12576 gnd.n5077 gnd.n2877 256.663
R12577 gnd.n2930 gnd.n2877 256.663
R12578 gnd.n5084 gnd.n2877 256.663
R12579 gnd.n2927 gnd.n2877 256.663
R12580 gnd.n5091 gnd.n2877 256.663
R12581 gnd.n2924 gnd.n2877 256.663
R12582 gnd.n5098 gnd.n2877 256.663
R12583 gnd.n2921 gnd.n2877 256.663
R12584 gnd.n5105 gnd.n2877 256.663
R12585 gnd.n2918 gnd.n2877 256.663
R12586 gnd.n5112 gnd.n2877 256.663
R12587 gnd.n2915 gnd.n2877 256.663
R12588 gnd.n5119 gnd.n2877 256.663
R12589 gnd.n2912 gnd.n2877 256.663
R12590 gnd.n3890 gnd.n2314 242.672
R12591 gnd.n3822 gnd.n2314 242.672
R12592 gnd.n3883 gnd.n2314 242.672
R12593 gnd.n3877 gnd.n2314 242.672
R12594 gnd.n3875 gnd.n2314 242.672
R12595 gnd.n3869 gnd.n2314 242.672
R12596 gnd.n3867 gnd.n2314 242.672
R12597 gnd.n3861 gnd.n2314 242.672
R12598 gnd.n3859 gnd.n2314 242.672
R12599 gnd.n4372 gnd.n3671 242.672
R12600 gnd.n4372 gnd.n3374 242.672
R12601 gnd.n4372 gnd.n3373 242.672
R12602 gnd.n4372 gnd.n3372 242.672
R12603 gnd.n4372 gnd.n3371 242.672
R12604 gnd.n4372 gnd.n3370 242.672
R12605 gnd.n4372 gnd.n3369 242.672
R12606 gnd.n4372 gnd.n3368 242.672
R12607 gnd.n4372 gnd.n3367 242.672
R12608 gnd.n1450 gnd.n1449 242.672
R12609 gnd.n1450 gnd.n1360 242.672
R12610 gnd.n1450 gnd.n1361 242.672
R12611 gnd.n1450 gnd.n1362 242.672
R12612 gnd.n1450 gnd.n1363 242.672
R12613 gnd.n1450 gnd.n1364 242.672
R12614 gnd.n1450 gnd.n1365 242.672
R12615 gnd.n1450 gnd.n1366 242.672
R12616 gnd.n1450 gnd.n1367 242.672
R12617 gnd.n1450 gnd.n1368 242.672
R12618 gnd.n1450 gnd.n1369 242.672
R12619 gnd.n1450 gnd.n1370 242.672
R12620 gnd.n1451 gnd.n1450 242.672
R12621 gnd.n2304 gnd.n856 242.672
R12622 gnd.n2304 gnd.n855 242.672
R12623 gnd.n2304 gnd.n854 242.672
R12624 gnd.n2304 gnd.n853 242.672
R12625 gnd.n2304 gnd.n852 242.672
R12626 gnd.n2304 gnd.n851 242.672
R12627 gnd.n2304 gnd.n850 242.672
R12628 gnd.n2304 gnd.n849 242.672
R12629 gnd.n2304 gnd.n848 242.672
R12630 gnd.n2304 gnd.n847 242.672
R12631 gnd.n2304 gnd.n846 242.672
R12632 gnd.n2304 gnd.n845 242.672
R12633 gnd.n2304 gnd.n844 242.672
R12634 gnd.n5927 gnd.n2735 242.672
R12635 gnd.n5927 gnd.n2736 242.672
R12636 gnd.n5927 gnd.n2737 242.672
R12637 gnd.n5927 gnd.n2738 242.672
R12638 gnd.n5927 gnd.n2739 242.672
R12639 gnd.n5927 gnd.n2740 242.672
R12640 gnd.n5927 gnd.n2741 242.672
R12641 gnd.n5927 gnd.n2742 242.672
R12642 gnd.n5927 gnd.n2743 242.672
R12643 gnd.n7331 gnd.n7330 242.672
R12644 gnd.n7330 gnd.n240 242.672
R12645 gnd.n7330 gnd.n189 242.672
R12646 gnd.n7330 gnd.n188 242.672
R12647 gnd.n7330 gnd.n187 242.672
R12648 gnd.n7330 gnd.n186 242.672
R12649 gnd.n7330 gnd.n185 242.672
R12650 gnd.n7330 gnd.n184 242.672
R12651 gnd.n7330 gnd.n183 242.672
R12652 gnd.n1534 gnd.n1533 242.672
R12653 gnd.n1533 gnd.n1272 242.672
R12654 gnd.n1533 gnd.n1273 242.672
R12655 gnd.n1533 gnd.n1274 242.672
R12656 gnd.n1533 gnd.n1275 242.672
R12657 gnd.n1533 gnd.n1276 242.672
R12658 gnd.n1533 gnd.n1277 242.672
R12659 gnd.n1533 gnd.n1278 242.672
R12660 gnd.n2304 gnd.n857 242.672
R12661 gnd.n2304 gnd.n858 242.672
R12662 gnd.n2304 gnd.n859 242.672
R12663 gnd.n2304 gnd.n860 242.672
R12664 gnd.n2304 gnd.n861 242.672
R12665 gnd.n2304 gnd.n862 242.672
R12666 gnd.n2304 gnd.n863 242.672
R12667 gnd.n2304 gnd.n864 242.672
R12668 gnd.n3958 gnd.n2314 242.672
R12669 gnd.n3966 gnd.n2314 242.672
R12670 gnd.n3968 gnd.n2314 242.672
R12671 gnd.n3976 gnd.n2314 242.672
R12672 gnd.n3978 gnd.n2314 242.672
R12673 gnd.n3986 gnd.n2314 242.672
R12674 gnd.n3988 gnd.n2314 242.672
R12675 gnd.n3996 gnd.n2314 242.672
R12676 gnd.n3998 gnd.n2314 242.672
R12677 gnd.n4006 gnd.n2314 242.672
R12678 gnd.n4008 gnd.n2314 242.672
R12679 gnd.n4016 gnd.n2314 242.672
R12680 gnd.n4018 gnd.n2314 242.672
R12681 gnd.n4026 gnd.n2314 242.672
R12682 gnd.n4028 gnd.n2314 242.672
R12683 gnd.n4036 gnd.n2314 242.672
R12684 gnd.n4038 gnd.n2314 242.672
R12685 gnd.n4046 gnd.n2314 242.672
R12686 gnd.n4048 gnd.n2314 242.672
R12687 gnd.n4058 gnd.n2314 242.672
R12688 gnd.n4060 gnd.n2314 242.672
R12689 gnd.n4068 gnd.n2314 242.672
R12690 gnd.n4070 gnd.n2314 242.672
R12691 gnd.n4078 gnd.n2314 242.672
R12692 gnd.n4080 gnd.n2314 242.672
R12693 gnd.n4088 gnd.n2314 242.672
R12694 gnd.n4090 gnd.n2314 242.672
R12695 gnd.n4099 gnd.n2314 242.672
R12696 gnd.n4102 gnd.n2314 242.672
R12697 gnd.n4426 gnd.n4372 242.672
R12698 gnd.n4421 gnd.n4372 242.672
R12699 gnd.n4433 gnd.n4372 242.672
R12700 gnd.n4412 gnd.n4372 242.672
R12701 gnd.n4440 gnd.n4372 242.672
R12702 gnd.n4405 gnd.n4372 242.672
R12703 gnd.n4447 gnd.n4372 242.672
R12704 gnd.n4398 gnd.n4372 242.672
R12705 gnd.n4454 gnd.n4372 242.672
R12706 gnd.n4457 gnd.n4372 242.672
R12707 gnd.n4389 gnd.n4372 242.672
R12708 gnd.n4466 gnd.n4372 242.672
R12709 gnd.n4380 gnd.n4372 242.672
R12710 gnd.n4473 gnd.n4372 242.672
R12711 gnd.n4476 gnd.n4372 242.672
R12712 gnd.n4372 gnd.n4280 242.672
R12713 gnd.n4482 gnd.n3361 242.672
R12714 gnd.n4372 gnd.n4281 242.672
R12715 gnd.n4372 gnd.n4282 242.672
R12716 gnd.n4372 gnd.n4283 242.672
R12717 gnd.n4372 gnd.n4284 242.672
R12718 gnd.n4372 gnd.n4285 242.672
R12719 gnd.n4372 gnd.n4286 242.672
R12720 gnd.n4372 gnd.n4287 242.672
R12721 gnd.n4372 gnd.n4288 242.672
R12722 gnd.n4372 gnd.n4289 242.672
R12723 gnd.n4372 gnd.n4290 242.672
R12724 gnd.n4372 gnd.n4291 242.672
R12725 gnd.n4372 gnd.n4292 242.672
R12726 gnd.n4372 gnd.n4371 242.672
R12727 gnd.n5927 gnd.n5926 242.672
R12728 gnd.n5927 gnd.n2707 242.672
R12729 gnd.n5927 gnd.n2708 242.672
R12730 gnd.n5927 gnd.n2709 242.672
R12731 gnd.n5927 gnd.n2710 242.672
R12732 gnd.n5927 gnd.n2711 242.672
R12733 gnd.n5927 gnd.n2712 242.672
R12734 gnd.n5927 gnd.n2713 242.672
R12735 gnd.n5927 gnd.n2714 242.672
R12736 gnd.n5927 gnd.n2715 242.672
R12737 gnd.n5927 gnd.n2716 242.672
R12738 gnd.n5927 gnd.n2717 242.672
R12739 gnd.n5927 gnd.n2718 242.672
R12740 gnd.n5874 gnd.n2778 242.672
R12741 gnd.n5927 gnd.n2719 242.672
R12742 gnd.n5927 gnd.n2720 242.672
R12743 gnd.n5927 gnd.n2721 242.672
R12744 gnd.n5927 gnd.n2722 242.672
R12745 gnd.n5927 gnd.n2723 242.672
R12746 gnd.n5927 gnd.n2724 242.672
R12747 gnd.n5927 gnd.n2725 242.672
R12748 gnd.n5927 gnd.n2726 242.672
R12749 gnd.n5927 gnd.n2727 242.672
R12750 gnd.n5927 gnd.n2728 242.672
R12751 gnd.n5927 gnd.n2729 242.672
R12752 gnd.n5927 gnd.n2730 242.672
R12753 gnd.n5927 gnd.n2731 242.672
R12754 gnd.n5927 gnd.n2732 242.672
R12755 gnd.n5927 gnd.n2733 242.672
R12756 gnd.n5927 gnd.n2734 242.672
R12757 gnd.n7330 gnd.n7118 242.672
R12758 gnd.n7330 gnd.n7119 242.672
R12759 gnd.n7330 gnd.n7120 242.672
R12760 gnd.n7330 gnd.n7121 242.672
R12761 gnd.n7330 gnd.n7122 242.672
R12762 gnd.n7330 gnd.n7123 242.672
R12763 gnd.n7330 gnd.n7124 242.672
R12764 gnd.n7330 gnd.n7125 242.672
R12765 gnd.n7330 gnd.n7126 242.672
R12766 gnd.n7330 gnd.n7127 242.672
R12767 gnd.n7330 gnd.n7128 242.672
R12768 gnd.n7330 gnd.n7129 242.672
R12769 gnd.n7330 gnd.n7130 242.672
R12770 gnd.n7330 gnd.n7131 242.672
R12771 gnd.n7330 gnd.n7132 242.672
R12772 gnd.n7330 gnd.n7133 242.672
R12773 gnd.n7330 gnd.n7134 242.672
R12774 gnd.n7330 gnd.n7135 242.672
R12775 gnd.n7330 gnd.n7136 242.672
R12776 gnd.n7330 gnd.n7137 242.672
R12777 gnd.n7330 gnd.n7138 242.672
R12778 gnd.n7330 gnd.n7139 242.672
R12779 gnd.n7330 gnd.n7140 242.672
R12780 gnd.n7330 gnd.n7141 242.672
R12781 gnd.n7330 gnd.n7142 242.672
R12782 gnd.n7330 gnd.n7143 242.672
R12783 gnd.n7330 gnd.n7144 242.672
R12784 gnd.n7330 gnd.n7145 242.672
R12785 gnd.n7330 gnd.n7329 242.672
R12786 gnd.n6069 gnd.n2550 242.672
R12787 gnd.n6069 gnd.n2551 242.672
R12788 gnd.n6069 gnd.n2552 242.672
R12789 gnd.n6069 gnd.n2553 242.672
R12790 gnd.n6069 gnd.n2554 242.672
R12791 gnd.n6069 gnd.n2555 242.672
R12792 gnd.n6069 gnd.n2556 242.672
R12793 gnd.n6069 gnd.n2557 242.672
R12794 gnd.n6069 gnd.n2558 242.672
R12795 gnd.n6069 gnd.n2559 242.672
R12796 gnd.n6069 gnd.n2560 242.672
R12797 gnd.n6069 gnd.n2561 242.672
R12798 gnd.n6069 gnd.n2562 242.672
R12799 gnd.n6069 gnd.n2563 242.672
R12800 gnd.n5934 gnd.n2696 242.672
R12801 gnd.n5934 gnd.n2695 242.672
R12802 gnd.n5934 gnd.n2694 242.672
R12803 gnd.n5934 gnd.n2693 242.672
R12804 gnd.n5934 gnd.n2692 242.672
R12805 gnd.n5934 gnd.n2691 242.672
R12806 gnd.n5934 gnd.n2690 242.672
R12807 gnd.n5934 gnd.n2689 242.672
R12808 gnd.n5934 gnd.n2688 242.672
R12809 gnd.n5934 gnd.n2687 242.672
R12810 gnd.n5934 gnd.n2686 242.672
R12811 gnd.n5934 gnd.n2685 242.672
R12812 gnd.n5934 gnd.n2684 242.672
R12813 gnd.n5934 gnd.n2697 242.672
R12814 gnd.n7146 gnd.n166 240.244
R12815 gnd.n7328 gnd.n7147 240.244
R12816 gnd.n7324 gnd.n7323 240.244
R12817 gnd.n7320 gnd.n7319 240.244
R12818 gnd.n7316 gnd.n7315 240.244
R12819 gnd.n7312 gnd.n7311 240.244
R12820 gnd.n7308 gnd.n7307 240.244
R12821 gnd.n7304 gnd.n7303 240.244
R12822 gnd.n7300 gnd.n7299 240.244
R12823 gnd.n7293 gnd.n7292 240.244
R12824 gnd.n7289 gnd.n7288 240.244
R12825 gnd.n7285 gnd.n7284 240.244
R12826 gnd.n7281 gnd.n7280 240.244
R12827 gnd.n7277 gnd.n7276 240.244
R12828 gnd.n7273 gnd.n7272 240.244
R12829 gnd.n7269 gnd.n7268 240.244
R12830 gnd.n7265 gnd.n7264 240.244
R12831 gnd.n7261 gnd.n7260 240.244
R12832 gnd.n7257 gnd.n7256 240.244
R12833 gnd.n7250 gnd.n7249 240.244
R12834 gnd.n7247 gnd.n7246 240.244
R12835 gnd.n7243 gnd.n7242 240.244
R12836 gnd.n7239 gnd.n7238 240.244
R12837 gnd.n7235 gnd.n7234 240.244
R12838 gnd.n7231 gnd.n7230 240.244
R12839 gnd.n7227 gnd.n7226 240.244
R12840 gnd.n7223 gnd.n7222 240.244
R12841 gnd.n7219 gnd.n7218 240.244
R12842 gnd.n7215 gnd.n7214 240.244
R12843 gnd.n5808 gnd.n2819 240.244
R12844 gnd.n5494 gnd.n2819 240.244
R12845 gnd.n5494 gnd.n5331 240.244
R12846 gnd.n5504 gnd.n5331 240.244
R12847 gnd.n5504 gnd.n5342 240.244
R12848 gnd.n5478 gnd.n5342 240.244
R12849 gnd.n5478 gnd.n5352 240.244
R12850 gnd.n5511 gnd.n5352 240.244
R12851 gnd.n5511 gnd.n5362 240.244
R12852 gnd.n5517 gnd.n5362 240.244
R12853 gnd.n5517 gnd.n5372 240.244
R12854 gnd.n5524 gnd.n5372 240.244
R12855 gnd.n5524 gnd.n5382 240.244
R12856 gnd.n5444 gnd.n5382 240.244
R12857 gnd.n5444 gnd.n5391 240.244
R12858 gnd.n5581 gnd.n5391 240.244
R12859 gnd.n5581 gnd.n5401 240.244
R12860 gnd.n5405 gnd.n5401 240.244
R12861 gnd.n5590 gnd.n5405 240.244
R12862 gnd.n5591 gnd.n5590 240.244
R12863 gnd.n5591 gnd.n5415 240.244
R12864 gnd.n5600 gnd.n5415 240.244
R12865 gnd.n5600 gnd.n69 240.244
R12866 gnd.n5425 gnd.n69 240.244
R12867 gnd.n5611 gnd.n5425 240.244
R12868 gnd.n5611 gnd.n86 240.244
R12869 gnd.n5432 gnd.n86 240.244
R12870 gnd.n5432 gnd.n97 240.244
R12871 gnd.n5712 gnd.n97 240.244
R12872 gnd.n5712 gnd.n107 240.244
R12873 gnd.n5708 gnd.n107 240.244
R12874 gnd.n5708 gnd.n117 240.244
R12875 gnd.n5700 gnd.n117 240.244
R12876 gnd.n5700 gnd.n128 240.244
R12877 gnd.n5696 gnd.n128 240.244
R12878 gnd.n5696 gnd.n137 240.244
R12879 gnd.n5641 gnd.n137 240.244
R12880 gnd.n5641 gnd.n148 240.244
R12881 gnd.n5637 gnd.n148 240.244
R12882 gnd.n5637 gnd.n158 240.244
R12883 gnd.n7340 gnd.n158 240.244
R12884 gnd.n7340 gnd.n168 240.244
R12885 gnd.n2747 gnd.n2746 240.244
R12886 gnd.n5920 gnd.n2746 240.244
R12887 gnd.n5918 gnd.n5917 240.244
R12888 gnd.n5914 gnd.n5913 240.244
R12889 gnd.n5910 gnd.n5909 240.244
R12890 gnd.n5906 gnd.n5905 240.244
R12891 gnd.n5902 gnd.n5901 240.244
R12892 gnd.n5898 gnd.n5897 240.244
R12893 gnd.n5894 gnd.n5893 240.244
R12894 gnd.n5889 gnd.n5888 240.244
R12895 gnd.n5885 gnd.n5884 240.244
R12896 gnd.n5881 gnd.n5880 240.244
R12897 gnd.n5877 gnd.n5876 240.244
R12898 gnd.n5872 gnd.n5871 240.244
R12899 gnd.n5868 gnd.n5867 240.244
R12900 gnd.n5864 gnd.n5863 240.244
R12901 gnd.n5860 gnd.n5859 240.244
R12902 gnd.n5856 gnd.n5855 240.244
R12903 gnd.n5852 gnd.n5851 240.244
R12904 gnd.n5848 gnd.n5847 240.244
R12905 gnd.n5844 gnd.n5843 240.244
R12906 gnd.n5840 gnd.n5839 240.244
R12907 gnd.n5836 gnd.n5835 240.244
R12908 gnd.n5832 gnd.n5831 240.244
R12909 gnd.n5828 gnd.n5827 240.244
R12910 gnd.n5824 gnd.n5823 240.244
R12911 gnd.n5820 gnd.n5819 240.244
R12912 gnd.n5816 gnd.n5815 240.244
R12913 gnd.n5803 gnd.n2748 240.244
R12914 gnd.n5803 gnd.n5322 240.244
R12915 gnd.n5799 gnd.n5322 240.244
R12916 gnd.n5799 gnd.n5329 240.244
R12917 gnd.n5791 gnd.n5329 240.244
R12918 gnd.n5791 gnd.n5345 240.244
R12919 gnd.n5787 gnd.n5345 240.244
R12920 gnd.n5787 gnd.n5351 240.244
R12921 gnd.n5779 gnd.n5351 240.244
R12922 gnd.n5779 gnd.n5364 240.244
R12923 gnd.n5775 gnd.n5364 240.244
R12924 gnd.n5775 gnd.n5370 240.244
R12925 gnd.n5767 gnd.n5370 240.244
R12926 gnd.n5767 gnd.n5385 240.244
R12927 gnd.n5763 gnd.n5385 240.244
R12928 gnd.n5763 gnd.n5390 240.244
R12929 gnd.n5755 gnd.n5390 240.244
R12930 gnd.n5755 gnd.n5752 240.244
R12931 gnd.n5752 gnd.n5403 240.244
R12932 gnd.n5738 gnd.n5403 240.244
R12933 gnd.n5741 gnd.n5738 240.244
R12934 gnd.n5741 gnd.n72 240.244
R12935 gnd.n7401 gnd.n72 240.244
R12936 gnd.n7401 gnd.n73 240.244
R12937 gnd.n83 gnd.n73 240.244
R12938 gnd.n7395 gnd.n83 240.244
R12939 gnd.n7395 gnd.n84 240.244
R12940 gnd.n7387 gnd.n84 240.244
R12941 gnd.n7387 gnd.n100 240.244
R12942 gnd.n7383 gnd.n100 240.244
R12943 gnd.n7383 gnd.n105 240.244
R12944 gnd.n7375 gnd.n105 240.244
R12945 gnd.n7375 gnd.n120 240.244
R12946 gnd.n7371 gnd.n120 240.244
R12947 gnd.n7371 gnd.n126 240.244
R12948 gnd.n7363 gnd.n126 240.244
R12949 gnd.n7363 gnd.n140 240.244
R12950 gnd.n7359 gnd.n140 240.244
R12951 gnd.n7359 gnd.n146 240.244
R12952 gnd.n7351 gnd.n146 240.244
R12953 gnd.n7351 gnd.n161 240.244
R12954 gnd.n7347 gnd.n161 240.244
R12955 gnd.n4293 gnd.n2531 240.244
R12956 gnd.n4370 gnd.n4294 240.244
R12957 gnd.n4366 gnd.n4365 240.244
R12958 gnd.n4362 gnd.n4361 240.244
R12959 gnd.n4358 gnd.n4357 240.244
R12960 gnd.n4354 gnd.n4353 240.244
R12961 gnd.n4350 gnd.n4349 240.244
R12962 gnd.n4346 gnd.n4345 240.244
R12963 gnd.n4342 gnd.n4341 240.244
R12964 gnd.n4337 gnd.n4336 240.244
R12965 gnd.n4333 gnd.n4332 240.244
R12966 gnd.n4329 gnd.n4328 240.244
R12967 gnd.n4325 gnd.n4324 240.244
R12968 gnd.n4477 gnd.n3365 240.244
R12969 gnd.n4475 gnd.n4474 240.244
R12970 gnd.n4472 gnd.n4374 240.244
R12971 gnd.n4468 gnd.n4467 240.244
R12972 gnd.n4465 gnd.n4381 240.244
R12973 gnd.n4458 gnd.n4390 240.244
R12974 gnd.n4456 gnd.n4455 240.244
R12975 gnd.n4453 gnd.n4392 240.244
R12976 gnd.n4449 gnd.n4448 240.244
R12977 gnd.n4446 gnd.n4399 240.244
R12978 gnd.n4442 gnd.n4441 240.244
R12979 gnd.n4439 gnd.n4406 240.244
R12980 gnd.n4435 gnd.n4434 240.244
R12981 gnd.n4432 gnd.n4413 240.244
R12982 gnd.n4428 gnd.n4427 240.244
R12983 gnd.n3819 gnd.n2323 240.244
R12984 gnd.n3819 gnd.n2335 240.244
R12985 gnd.n4113 gnd.n2335 240.244
R12986 gnd.n4113 gnd.n2347 240.244
R12987 gnd.n4123 gnd.n2347 240.244
R12988 gnd.n4123 gnd.n2358 240.244
R12989 gnd.n4127 gnd.n2358 240.244
R12990 gnd.n4127 gnd.n2367 240.244
R12991 gnd.n4137 gnd.n2367 240.244
R12992 gnd.n4137 gnd.n2378 240.244
R12993 gnd.n4141 gnd.n2378 240.244
R12994 gnd.n4141 gnd.n2388 240.244
R12995 gnd.n4151 gnd.n2388 240.244
R12996 gnd.n4151 gnd.n2399 240.244
R12997 gnd.n4155 gnd.n2399 240.244
R12998 gnd.n4155 gnd.n2408 240.244
R12999 gnd.n4165 gnd.n2408 240.244
R13000 gnd.n4165 gnd.n2417 240.244
R13001 gnd.n4169 gnd.n2417 240.244
R13002 gnd.n4169 gnd.n2427 240.244
R13003 gnd.n4179 gnd.n2427 240.244
R13004 gnd.n4179 gnd.n2435 240.244
R13005 gnd.n4183 gnd.n2435 240.244
R13006 gnd.n4183 gnd.n2444 240.244
R13007 gnd.n4193 gnd.n2444 240.244
R13008 gnd.n4193 gnd.n2452 240.244
R13009 gnd.n4197 gnd.n2452 240.244
R13010 gnd.n4197 gnd.n2462 240.244
R13011 gnd.n4207 gnd.n2462 240.244
R13012 gnd.n4207 gnd.n2473 240.244
R13013 gnd.n3689 gnd.n2473 240.244
R13014 gnd.n3689 gnd.n2482 240.244
R13015 gnd.n4214 gnd.n2482 240.244
R13016 gnd.n4214 gnd.n2493 240.244
R13017 gnd.n4218 gnd.n2493 240.244
R13018 gnd.n4218 gnd.n2503 240.244
R13019 gnd.n4223 gnd.n2503 240.244
R13020 gnd.n4223 gnd.n2514 240.244
R13021 gnd.n4227 gnd.n2514 240.244
R13022 gnd.n4227 gnd.n2524 240.244
R13023 gnd.n6080 gnd.n2524 240.244
R13024 gnd.n6080 gnd.n2533 240.244
R13025 gnd.n3959 gnd.n3954 240.244
R13026 gnd.n3965 gnd.n3954 240.244
R13027 gnd.n3969 gnd.n3967 240.244
R13028 gnd.n3975 gnd.n3950 240.244
R13029 gnd.n3979 gnd.n3977 240.244
R13030 gnd.n3985 gnd.n3946 240.244
R13031 gnd.n3989 gnd.n3987 240.244
R13032 gnd.n3995 gnd.n3942 240.244
R13033 gnd.n3999 gnd.n3997 240.244
R13034 gnd.n4005 gnd.n3935 240.244
R13035 gnd.n4009 gnd.n4007 240.244
R13036 gnd.n4015 gnd.n3931 240.244
R13037 gnd.n4019 gnd.n4017 240.244
R13038 gnd.n4025 gnd.n3927 240.244
R13039 gnd.n4029 gnd.n4027 240.244
R13040 gnd.n4035 gnd.n3923 240.244
R13041 gnd.n4039 gnd.n4037 240.244
R13042 gnd.n4045 gnd.n3919 240.244
R13043 gnd.n4049 gnd.n4047 240.244
R13044 gnd.n4057 gnd.n3915 240.244
R13045 gnd.n4061 gnd.n4059 240.244
R13046 gnd.n4067 gnd.n3911 240.244
R13047 gnd.n4071 gnd.n4069 240.244
R13048 gnd.n4077 gnd.n3907 240.244
R13049 gnd.n4081 gnd.n4079 240.244
R13050 gnd.n4087 gnd.n3903 240.244
R13051 gnd.n4091 gnd.n4089 240.244
R13052 gnd.n4098 gnd.n3899 240.244
R13053 gnd.n4101 gnd.n4100 240.244
R13054 gnd.n6214 gnd.n2328 240.244
R13055 gnd.n6210 gnd.n2328 240.244
R13056 gnd.n6210 gnd.n2333 240.244
R13057 gnd.n6202 gnd.n2333 240.244
R13058 gnd.n6202 gnd.n2350 240.244
R13059 gnd.n6198 gnd.n2350 240.244
R13060 gnd.n6198 gnd.n2356 240.244
R13061 gnd.n6190 gnd.n2356 240.244
R13062 gnd.n6190 gnd.n2370 240.244
R13063 gnd.n6186 gnd.n2370 240.244
R13064 gnd.n6186 gnd.n2376 240.244
R13065 gnd.n6178 gnd.n2376 240.244
R13066 gnd.n6178 gnd.n2391 240.244
R13067 gnd.n6174 gnd.n2391 240.244
R13068 gnd.n6174 gnd.n2397 240.244
R13069 gnd.n6166 gnd.n2397 240.244
R13070 gnd.n6166 gnd.n2411 240.244
R13071 gnd.n6161 gnd.n2411 240.244
R13072 gnd.n6161 gnd.n2415 240.244
R13073 gnd.n6153 gnd.n2415 240.244
R13074 gnd.n6153 gnd.n2430 240.244
R13075 gnd.n6148 gnd.n2430 240.244
R13076 gnd.n6148 gnd.n2433 240.244
R13077 gnd.n6140 gnd.n2433 240.244
R13078 gnd.n6140 gnd.n2447 240.244
R13079 gnd.n6135 gnd.n2447 240.244
R13080 gnd.n6135 gnd.n2450 240.244
R13081 gnd.n6127 gnd.n2450 240.244
R13082 gnd.n6127 gnd.n2465 240.244
R13083 gnd.n6123 gnd.n2465 240.244
R13084 gnd.n6123 gnd.n2471 240.244
R13085 gnd.n6115 gnd.n2471 240.244
R13086 gnd.n6115 gnd.n2485 240.244
R13087 gnd.n6111 gnd.n2485 240.244
R13088 gnd.n6111 gnd.n2491 240.244
R13089 gnd.n6103 gnd.n2491 240.244
R13090 gnd.n6103 gnd.n2506 240.244
R13091 gnd.n6099 gnd.n2506 240.244
R13092 gnd.n6099 gnd.n2512 240.244
R13093 gnd.n6091 gnd.n2512 240.244
R13094 gnd.n6091 gnd.n2526 240.244
R13095 gnd.n6087 gnd.n2526 240.244
R13096 gnd.n2303 gnd.n866 240.244
R13097 gnd.n2296 gnd.n2295 240.244
R13098 gnd.n2293 gnd.n2292 240.244
R13099 gnd.n2289 gnd.n2288 240.244
R13100 gnd.n2285 gnd.n2284 240.244
R13101 gnd.n2281 gnd.n2280 240.244
R13102 gnd.n2277 gnd.n2276 240.244
R13103 gnd.n2273 gnd.n2272 240.244
R13104 gnd.n1545 gnd.n1257 240.244
R13105 gnd.n1555 gnd.n1257 240.244
R13106 gnd.n1555 gnd.n1248 240.244
R13107 gnd.n1248 gnd.n1237 240.244
R13108 gnd.n1576 gnd.n1237 240.244
R13109 gnd.n1576 gnd.n1231 240.244
R13110 gnd.n1586 gnd.n1231 240.244
R13111 gnd.n1586 gnd.n1220 240.244
R13112 gnd.n1220 gnd.n1212 240.244
R13113 gnd.n1604 gnd.n1212 240.244
R13114 gnd.n1605 gnd.n1604 240.244
R13115 gnd.n1605 gnd.n1197 240.244
R13116 gnd.n1607 gnd.n1197 240.244
R13117 gnd.n1607 gnd.n1183 240.244
R13118 gnd.n1649 gnd.n1183 240.244
R13119 gnd.n1650 gnd.n1649 240.244
R13120 gnd.n1653 gnd.n1650 240.244
R13121 gnd.n1653 gnd.n1138 240.244
R13122 gnd.n1178 gnd.n1138 240.244
R13123 gnd.n1178 gnd.n1148 240.244
R13124 gnd.n1663 gnd.n1148 240.244
R13125 gnd.n1663 gnd.n1169 240.244
R13126 gnd.n1673 gnd.n1169 240.244
R13127 gnd.n1673 gnd.n1067 240.244
R13128 gnd.n1718 gnd.n1067 240.244
R13129 gnd.n1718 gnd.n1053 240.244
R13130 gnd.n1740 gnd.n1053 240.244
R13131 gnd.n1741 gnd.n1740 240.244
R13132 gnd.n1741 gnd.n1040 240.244
R13133 gnd.n1040 gnd.n1029 240.244
R13134 gnd.n1772 gnd.n1029 240.244
R13135 gnd.n1773 gnd.n1772 240.244
R13136 gnd.n1774 gnd.n1773 240.244
R13137 gnd.n1774 gnd.n1014 240.244
R13138 gnd.n1805 gnd.n1014 240.244
R13139 gnd.n1805 gnd.n999 240.244
R13140 gnd.n1827 gnd.n999 240.244
R13141 gnd.n1828 gnd.n1827 240.244
R13142 gnd.n1828 gnd.n986 240.244
R13143 gnd.n986 gnd.n975 240.244
R13144 gnd.n1859 gnd.n975 240.244
R13145 gnd.n1860 gnd.n1859 240.244
R13146 gnd.n1861 gnd.n1860 240.244
R13147 gnd.n1861 gnd.n959 240.244
R13148 gnd.n959 gnd.n958 240.244
R13149 gnd.n958 gnd.n945 240.244
R13150 gnd.n1916 gnd.n945 240.244
R13151 gnd.n1917 gnd.n1916 240.244
R13152 gnd.n1917 gnd.n932 240.244
R13153 gnd.n932 gnd.n922 240.244
R13154 gnd.n2204 gnd.n922 240.244
R13155 gnd.n2207 gnd.n2204 240.244
R13156 gnd.n2207 gnd.n2206 240.244
R13157 gnd.n1535 gnd.n1270 240.244
R13158 gnd.n1291 gnd.n1270 240.244
R13159 gnd.n1294 gnd.n1293 240.244
R13160 gnd.n1301 gnd.n1300 240.244
R13161 gnd.n1304 gnd.n1303 240.244
R13162 gnd.n1311 gnd.n1310 240.244
R13163 gnd.n1314 gnd.n1313 240.244
R13164 gnd.n1321 gnd.n1320 240.244
R13165 gnd.n1543 gnd.n1267 240.244
R13166 gnd.n1267 gnd.n1246 240.244
R13167 gnd.n1566 gnd.n1246 240.244
R13168 gnd.n1566 gnd.n1240 240.244
R13169 gnd.n1574 gnd.n1240 240.244
R13170 gnd.n1574 gnd.n1242 240.244
R13171 gnd.n1242 gnd.n1218 240.244
R13172 gnd.n1596 gnd.n1218 240.244
R13173 gnd.n1596 gnd.n1214 240.244
R13174 gnd.n1602 gnd.n1214 240.244
R13175 gnd.n1602 gnd.n1196 240.244
R13176 gnd.n1627 gnd.n1196 240.244
R13177 gnd.n1627 gnd.n1191 240.244
R13178 gnd.n1639 gnd.n1191 240.244
R13179 gnd.n1639 gnd.n1192 240.244
R13180 gnd.n1635 gnd.n1192 240.244
R13181 gnd.n1635 gnd.n1140 240.244
R13182 gnd.n1687 gnd.n1140 240.244
R13183 gnd.n1687 gnd.n1141 240.244
R13184 gnd.n1683 gnd.n1141 240.244
R13185 gnd.n1683 gnd.n1147 240.244
R13186 gnd.n1167 gnd.n1147 240.244
R13187 gnd.n1167 gnd.n1065 240.244
R13188 gnd.n1722 gnd.n1065 240.244
R13189 gnd.n1722 gnd.n1060 240.244
R13190 gnd.n1730 gnd.n1060 240.244
R13191 gnd.n1730 gnd.n1061 240.244
R13192 gnd.n1061 gnd.n1038 240.244
R13193 gnd.n1762 gnd.n1038 240.244
R13194 gnd.n1762 gnd.n1033 240.244
R13195 gnd.n1770 gnd.n1033 240.244
R13196 gnd.n1770 gnd.n1034 240.244
R13197 gnd.n1034 gnd.n1012 240.244
R13198 gnd.n1809 gnd.n1012 240.244
R13199 gnd.n1809 gnd.n1007 240.244
R13200 gnd.n1817 gnd.n1007 240.244
R13201 gnd.n1817 gnd.n1008 240.244
R13202 gnd.n1008 gnd.n984 240.244
R13203 gnd.n1849 gnd.n984 240.244
R13204 gnd.n1849 gnd.n979 240.244
R13205 gnd.n1857 gnd.n979 240.244
R13206 gnd.n1857 gnd.n980 240.244
R13207 gnd.n980 gnd.n957 240.244
R13208 gnd.n1898 gnd.n957 240.244
R13209 gnd.n1898 gnd.n952 240.244
R13210 gnd.n1906 gnd.n952 240.244
R13211 gnd.n1906 gnd.n953 240.244
R13212 gnd.n953 gnd.n930 240.244
R13213 gnd.n2192 gnd.n930 240.244
R13214 gnd.n2192 gnd.n925 240.244
R13215 gnd.n2202 gnd.n925 240.244
R13216 gnd.n2202 gnd.n926 240.244
R13217 gnd.n926 gnd.n865 240.244
R13218 gnd.n201 gnd.n171 240.244
R13219 gnd.n204 gnd.n203 240.244
R13220 gnd.n211 gnd.n210 240.244
R13221 gnd.n214 gnd.n213 240.244
R13222 gnd.n221 gnd.n220 240.244
R13223 gnd.n224 gnd.n223 240.244
R13224 gnd.n231 gnd.n230 240.244
R13225 gnd.n233 gnd.n190 240.244
R13226 gnd.n239 gnd.n181 240.244
R13227 gnd.n5320 gnd.n2821 240.244
R13228 gnd.n5496 gnd.n5320 240.244
R13229 gnd.n5496 gnd.n5332 240.244
R13230 gnd.n5502 gnd.n5332 240.244
R13231 gnd.n5502 gnd.n5343 240.244
R13232 gnd.n5538 gnd.n5343 240.244
R13233 gnd.n5538 gnd.n5353 240.244
R13234 gnd.n5483 gnd.n5353 240.244
R13235 gnd.n5483 gnd.n5363 240.244
R13236 gnd.n5484 gnd.n5363 240.244
R13237 gnd.n5484 gnd.n5373 240.244
R13238 gnd.n5526 gnd.n5373 240.244
R13239 gnd.n5526 gnd.n5383 240.244
R13240 gnd.n5565 gnd.n5383 240.244
R13241 gnd.n5565 gnd.n5392 240.244
R13242 gnd.n5579 gnd.n5392 240.244
R13243 gnd.n5579 gnd.n5402 240.244
R13244 gnd.n5406 gnd.n5402 240.244
R13245 gnd.n5570 gnd.n5406 240.244
R13246 gnd.n5571 gnd.n5570 240.244
R13247 gnd.n5571 gnd.n5416 240.244
R13248 gnd.n5416 gnd.n66 240.244
R13249 gnd.n7403 gnd.n66 240.244
R13250 gnd.n7403 gnd.n68 240.244
R13251 gnd.n5609 gnd.n68 240.244
R13252 gnd.n5609 gnd.n87 240.244
R13253 gnd.n5718 gnd.n87 240.244
R13254 gnd.n5718 gnd.n98 240.244
R13255 gnd.n5714 gnd.n98 240.244
R13256 gnd.n5714 gnd.n108 240.244
R13257 gnd.n5706 gnd.n108 240.244
R13258 gnd.n5706 gnd.n118 240.244
R13259 gnd.n5702 gnd.n118 240.244
R13260 gnd.n5702 gnd.n129 240.244
R13261 gnd.n5647 gnd.n129 240.244
R13262 gnd.n5647 gnd.n138 240.244
R13263 gnd.n5643 gnd.n138 240.244
R13264 gnd.n5643 gnd.n149 240.244
R13265 gnd.n5635 gnd.n149 240.244
R13266 gnd.n5635 gnd.n159 240.244
R13267 gnd.n7338 gnd.n159 240.244
R13268 gnd.n7338 gnd.n169 240.244
R13269 gnd.n2825 gnd.n2824 240.244
R13270 gnd.n5216 gnd.n5215 240.244
R13271 gnd.n5224 gnd.n5223 240.244
R13272 gnd.n5226 gnd.n5225 240.244
R13273 gnd.n5236 gnd.n5235 240.244
R13274 gnd.n5244 gnd.n5243 240.244
R13275 gnd.n5246 gnd.n5245 240.244
R13276 gnd.n5256 gnd.n5255 240.244
R13277 gnd.n5257 gnd.n2744 240.244
R13278 gnd.n5806 gnd.n5805 240.244
R13279 gnd.n5805 gnd.n5318 240.244
R13280 gnd.n5797 gnd.n5318 240.244
R13281 gnd.n5797 gnd.n5334 240.244
R13282 gnd.n5793 gnd.n5334 240.244
R13283 gnd.n5793 gnd.n5340 240.244
R13284 gnd.n5785 gnd.n5340 240.244
R13285 gnd.n5785 gnd.n5355 240.244
R13286 gnd.n5781 gnd.n5355 240.244
R13287 gnd.n5781 gnd.n5360 240.244
R13288 gnd.n5773 gnd.n5360 240.244
R13289 gnd.n5773 gnd.n5375 240.244
R13290 gnd.n5769 gnd.n5375 240.244
R13291 gnd.n5769 gnd.n5380 240.244
R13292 gnd.n5761 gnd.n5380 240.244
R13293 gnd.n5761 gnd.n5394 240.244
R13294 gnd.n5757 gnd.n5394 240.244
R13295 gnd.n5757 gnd.n5399 240.244
R13296 gnd.n5586 gnd.n5399 240.244
R13297 gnd.n5586 gnd.n5418 240.244
R13298 gnd.n5735 gnd.n5418 240.244
R13299 gnd.n5735 gnd.n5419 240.244
R13300 gnd.n5419 gnd.n71 240.244
R13301 gnd.n5730 gnd.n71 240.244
R13302 gnd.n5730 gnd.n89 240.244
R13303 gnd.n7393 gnd.n89 240.244
R13304 gnd.n7393 gnd.n90 240.244
R13305 gnd.n7389 gnd.n90 240.244
R13306 gnd.n7389 gnd.n96 240.244
R13307 gnd.n7381 gnd.n96 240.244
R13308 gnd.n7381 gnd.n110 240.244
R13309 gnd.n7377 gnd.n110 240.244
R13310 gnd.n7377 gnd.n115 240.244
R13311 gnd.n7369 gnd.n115 240.244
R13312 gnd.n7369 gnd.n131 240.244
R13313 gnd.n7365 gnd.n131 240.244
R13314 gnd.n7365 gnd.n136 240.244
R13315 gnd.n7357 gnd.n136 240.244
R13316 gnd.n7357 gnd.n151 240.244
R13317 gnd.n7353 gnd.n151 240.244
R13318 gnd.n7353 gnd.n156 240.244
R13319 gnd.n7345 gnd.n156 240.244
R13320 gnd.n885 gnd.n843 240.244
R13321 gnd.n2263 gnd.n2262 240.244
R13322 gnd.n2259 gnd.n2258 240.244
R13323 gnd.n2255 gnd.n2254 240.244
R13324 gnd.n2251 gnd.n2250 240.244
R13325 gnd.n2247 gnd.n2246 240.244
R13326 gnd.n2243 gnd.n2242 240.244
R13327 gnd.n2239 gnd.n2238 240.244
R13328 gnd.n2235 gnd.n2234 240.244
R13329 gnd.n2231 gnd.n2230 240.244
R13330 gnd.n2227 gnd.n2226 240.244
R13331 gnd.n2223 gnd.n2222 240.244
R13332 gnd.n2219 gnd.n2218 240.244
R13333 gnd.n1458 gnd.n1355 240.244
R13334 gnd.n1458 gnd.n1348 240.244
R13335 gnd.n1469 gnd.n1348 240.244
R13336 gnd.n1469 gnd.n1344 240.244
R13337 gnd.n1475 gnd.n1344 240.244
R13338 gnd.n1475 gnd.n1336 240.244
R13339 gnd.n1485 gnd.n1336 240.244
R13340 gnd.n1485 gnd.n1331 240.244
R13341 gnd.n1521 gnd.n1331 240.244
R13342 gnd.n1521 gnd.n1332 240.244
R13343 gnd.n1332 gnd.n1279 240.244
R13344 gnd.n1516 gnd.n1279 240.244
R13345 gnd.n1516 gnd.n1515 240.244
R13346 gnd.n1515 gnd.n1258 240.244
R13347 gnd.n1511 gnd.n1258 240.244
R13348 gnd.n1511 gnd.n1249 240.244
R13349 gnd.n1508 gnd.n1249 240.244
R13350 gnd.n1508 gnd.n1507 240.244
R13351 gnd.n1507 gnd.n1232 240.244
R13352 gnd.n1503 gnd.n1232 240.244
R13353 gnd.n1503 gnd.n1221 240.244
R13354 gnd.n1221 gnd.n1202 240.244
R13355 gnd.n1616 gnd.n1202 240.244
R13356 gnd.n1616 gnd.n1198 240.244
R13357 gnd.n1624 gnd.n1198 240.244
R13358 gnd.n1624 gnd.n1189 240.244
R13359 gnd.n1189 gnd.n1125 240.244
R13360 gnd.n1696 gnd.n1125 240.244
R13361 gnd.n1696 gnd.n1126 240.244
R13362 gnd.n1137 gnd.n1126 240.244
R13363 gnd.n1172 gnd.n1137 240.244
R13364 gnd.n1175 gnd.n1172 240.244
R13365 gnd.n1175 gnd.n1149 240.244
R13366 gnd.n1162 gnd.n1149 240.244
R13367 gnd.n1162 gnd.n1159 240.244
R13368 gnd.n1159 gnd.n1068 240.244
R13369 gnd.n1717 gnd.n1068 240.244
R13370 gnd.n1717 gnd.n1058 240.244
R13371 gnd.n1713 gnd.n1058 240.244
R13372 gnd.n1713 gnd.n1052 240.244
R13373 gnd.n1710 gnd.n1052 240.244
R13374 gnd.n1710 gnd.n1041 240.244
R13375 gnd.n1707 gnd.n1041 240.244
R13376 gnd.n1707 gnd.n1019 240.244
R13377 gnd.n1783 gnd.n1019 240.244
R13378 gnd.n1783 gnd.n1015 240.244
R13379 gnd.n1804 gnd.n1015 240.244
R13380 gnd.n1804 gnd.n1005 240.244
R13381 gnd.n1800 gnd.n1005 240.244
R13382 gnd.n1800 gnd.n998 240.244
R13383 gnd.n1797 gnd.n998 240.244
R13384 gnd.n1797 gnd.n987 240.244
R13385 gnd.n1794 gnd.n987 240.244
R13386 gnd.n1794 gnd.n964 240.244
R13387 gnd.n1870 gnd.n964 240.244
R13388 gnd.n1870 gnd.n960 240.244
R13389 gnd.n1895 gnd.n960 240.244
R13390 gnd.n1895 gnd.n951 240.244
R13391 gnd.n1891 gnd.n951 240.244
R13392 gnd.n1891 gnd.n944 240.244
R13393 gnd.n1887 gnd.n944 240.244
R13394 gnd.n1887 gnd.n933 240.244
R13395 gnd.n1884 gnd.n933 240.244
R13396 gnd.n1884 gnd.n914 240.244
R13397 gnd.n2214 gnd.n914 240.244
R13398 gnd.n1372 gnd.n1371 240.244
R13399 gnd.n1443 gnd.n1371 240.244
R13400 gnd.n1441 gnd.n1440 240.244
R13401 gnd.n1437 gnd.n1436 240.244
R13402 gnd.n1433 gnd.n1432 240.244
R13403 gnd.n1429 gnd.n1428 240.244
R13404 gnd.n1425 gnd.n1424 240.244
R13405 gnd.n1421 gnd.n1420 240.244
R13406 gnd.n1417 gnd.n1416 240.244
R13407 gnd.n1413 gnd.n1412 240.244
R13408 gnd.n1409 gnd.n1408 240.244
R13409 gnd.n1405 gnd.n1404 240.244
R13410 gnd.n1401 gnd.n1359 240.244
R13411 gnd.n1461 gnd.n1353 240.244
R13412 gnd.n1461 gnd.n1349 240.244
R13413 gnd.n1467 gnd.n1349 240.244
R13414 gnd.n1467 gnd.n1342 240.244
R13415 gnd.n1477 gnd.n1342 240.244
R13416 gnd.n1477 gnd.n1338 240.244
R13417 gnd.n1483 gnd.n1338 240.244
R13418 gnd.n1483 gnd.n1329 240.244
R13419 gnd.n1523 gnd.n1329 240.244
R13420 gnd.n1523 gnd.n1280 240.244
R13421 gnd.n1531 gnd.n1280 240.244
R13422 gnd.n1531 gnd.n1281 240.244
R13423 gnd.n1281 gnd.n1259 240.244
R13424 gnd.n1552 gnd.n1259 240.244
R13425 gnd.n1552 gnd.n1251 240.244
R13426 gnd.n1563 gnd.n1251 240.244
R13427 gnd.n1563 gnd.n1252 240.244
R13428 gnd.n1252 gnd.n1233 240.244
R13429 gnd.n1583 gnd.n1233 240.244
R13430 gnd.n1583 gnd.n1223 240.244
R13431 gnd.n1593 gnd.n1223 240.244
R13432 gnd.n1593 gnd.n1204 240.244
R13433 gnd.n1614 gnd.n1204 240.244
R13434 gnd.n1614 gnd.n1206 240.244
R13435 gnd.n1206 gnd.n1187 240.244
R13436 gnd.n1642 gnd.n1187 240.244
R13437 gnd.n1642 gnd.n1129 240.244
R13438 gnd.n1694 gnd.n1129 240.244
R13439 gnd.n1694 gnd.n1130 240.244
R13440 gnd.n1690 gnd.n1130 240.244
R13441 gnd.n1690 gnd.n1136 240.244
R13442 gnd.n1151 gnd.n1136 240.244
R13443 gnd.n1680 gnd.n1151 240.244
R13444 gnd.n1680 gnd.n1152 240.244
R13445 gnd.n1676 gnd.n1152 240.244
R13446 gnd.n1676 gnd.n1158 240.244
R13447 gnd.n1158 gnd.n1057 240.244
R13448 gnd.n1733 gnd.n1057 240.244
R13449 gnd.n1733 gnd.n1050 240.244
R13450 gnd.n1744 gnd.n1050 240.244
R13451 gnd.n1744 gnd.n1043 240.244
R13452 gnd.n1759 gnd.n1043 240.244
R13453 gnd.n1759 gnd.n1044 240.244
R13454 gnd.n1044 gnd.n1022 240.244
R13455 gnd.n1781 gnd.n1022 240.244
R13456 gnd.n1781 gnd.n1023 240.244
R13457 gnd.n1023 gnd.n1003 240.244
R13458 gnd.n1820 gnd.n1003 240.244
R13459 gnd.n1820 gnd.n996 240.244
R13460 gnd.n1831 gnd.n996 240.244
R13461 gnd.n1831 gnd.n989 240.244
R13462 gnd.n1846 gnd.n989 240.244
R13463 gnd.n1846 gnd.n990 240.244
R13464 gnd.n990 gnd.n967 240.244
R13465 gnd.n1868 gnd.n967 240.244
R13466 gnd.n1868 gnd.n969 240.244
R13467 gnd.n969 gnd.n949 240.244
R13468 gnd.n1909 gnd.n949 240.244
R13469 gnd.n1909 gnd.n942 240.244
R13470 gnd.n1920 gnd.n942 240.244
R13471 gnd.n1920 gnd.n935 240.244
R13472 gnd.n2189 gnd.n935 240.244
R13473 gnd.n2189 gnd.n936 240.244
R13474 gnd.n936 gnd.n917 240.244
R13475 gnd.n2212 gnd.n917 240.244
R13476 gnd.n3411 gnd.n2536 240.244
R13477 gnd.n3608 gnd.n3607 240.244
R13478 gnd.n3405 gnd.n3404 240.244
R13479 gnd.n3620 gnd.n3619 240.244
R13480 gnd.n3632 gnd.n3631 240.244
R13481 gnd.n3393 gnd.n3392 240.244
R13482 gnd.n3644 gnd.n3643 240.244
R13483 gnd.n3656 gnd.n3655 240.244
R13484 gnd.n3376 gnd.n3375 240.244
R13485 gnd.n3849 gnd.n2324 240.244
R13486 gnd.n3849 gnd.n2336 240.244
R13487 gnd.n4115 gnd.n2336 240.244
R13488 gnd.n4115 gnd.n2348 240.244
R13489 gnd.n4121 gnd.n2348 240.244
R13490 gnd.n4121 gnd.n2359 240.244
R13491 gnd.n4129 gnd.n2359 240.244
R13492 gnd.n4129 gnd.n2368 240.244
R13493 gnd.n4135 gnd.n2368 240.244
R13494 gnd.n4135 gnd.n2379 240.244
R13495 gnd.n4143 gnd.n2379 240.244
R13496 gnd.n4143 gnd.n2389 240.244
R13497 gnd.n4149 gnd.n2389 240.244
R13498 gnd.n4149 gnd.n2400 240.244
R13499 gnd.n4157 gnd.n2400 240.244
R13500 gnd.n4157 gnd.n2409 240.244
R13501 gnd.n4163 gnd.n2409 240.244
R13502 gnd.n4163 gnd.n2418 240.244
R13503 gnd.n4171 gnd.n2418 240.244
R13504 gnd.n4171 gnd.n2428 240.244
R13505 gnd.n4177 gnd.n2428 240.244
R13506 gnd.n4177 gnd.n2436 240.244
R13507 gnd.n4185 gnd.n2436 240.244
R13508 gnd.n4185 gnd.n2445 240.244
R13509 gnd.n4191 gnd.n2445 240.244
R13510 gnd.n4191 gnd.n2453 240.244
R13511 gnd.n4199 gnd.n2453 240.244
R13512 gnd.n4199 gnd.n2463 240.244
R13513 gnd.n4205 gnd.n2463 240.244
R13514 gnd.n4205 gnd.n2474 240.244
R13515 gnd.n4244 gnd.n2474 240.244
R13516 gnd.n4244 gnd.n2483 240.244
R13517 gnd.n3694 gnd.n2483 240.244
R13518 gnd.n3694 gnd.n2494 240.244
R13519 gnd.n3695 gnd.n2494 240.244
R13520 gnd.n3695 gnd.n2504 240.244
R13521 gnd.n3698 gnd.n2504 240.244
R13522 gnd.n3698 gnd.n2515 240.244
R13523 gnd.n4229 gnd.n2515 240.244
R13524 gnd.n4229 gnd.n2525 240.244
R13525 gnd.n6078 gnd.n2525 240.244
R13526 gnd.n6078 gnd.n2534 240.244
R13527 gnd.n3889 gnd.n3888 240.244
R13528 gnd.n3885 gnd.n3884 240.244
R13529 gnd.n3882 gnd.n3826 240.244
R13530 gnd.n3878 gnd.n3876 240.244
R13531 gnd.n3874 gnd.n3832 240.244
R13532 gnd.n3870 gnd.n3868 240.244
R13533 gnd.n3866 gnd.n3838 240.244
R13534 gnd.n3862 gnd.n3860 240.244
R13535 gnd.n3858 gnd.n3844 240.244
R13536 gnd.n2338 gnd.n2326 240.244
R13537 gnd.n6208 gnd.n2338 240.244
R13538 gnd.n6208 gnd.n2339 240.244
R13539 gnd.n6204 gnd.n2339 240.244
R13540 gnd.n6204 gnd.n2345 240.244
R13541 gnd.n6196 gnd.n2345 240.244
R13542 gnd.n6196 gnd.n2360 240.244
R13543 gnd.n6192 gnd.n2360 240.244
R13544 gnd.n6192 gnd.n2365 240.244
R13545 gnd.n6184 gnd.n2365 240.244
R13546 gnd.n6184 gnd.n2381 240.244
R13547 gnd.n6180 gnd.n2381 240.244
R13548 gnd.n6180 gnd.n2386 240.244
R13549 gnd.n6172 gnd.n2386 240.244
R13550 gnd.n6172 gnd.n2401 240.244
R13551 gnd.n6168 gnd.n2401 240.244
R13552 gnd.n6168 gnd.n2406 240.244
R13553 gnd.n6159 gnd.n2406 240.244
R13554 gnd.n6159 gnd.n2420 240.244
R13555 gnd.n6155 gnd.n2420 240.244
R13556 gnd.n6155 gnd.n2425 240.244
R13557 gnd.n6146 gnd.n2425 240.244
R13558 gnd.n6146 gnd.n2437 240.244
R13559 gnd.n6142 gnd.n2437 240.244
R13560 gnd.n6142 gnd.n2442 240.244
R13561 gnd.n6133 gnd.n2442 240.244
R13562 gnd.n6133 gnd.n2455 240.244
R13563 gnd.n6129 gnd.n2455 240.244
R13564 gnd.n6129 gnd.n2460 240.244
R13565 gnd.n6121 gnd.n2460 240.244
R13566 gnd.n6121 gnd.n2475 240.244
R13567 gnd.n6117 gnd.n2475 240.244
R13568 gnd.n6117 gnd.n2480 240.244
R13569 gnd.n6109 gnd.n2480 240.244
R13570 gnd.n6109 gnd.n2496 240.244
R13571 gnd.n6105 gnd.n2496 240.244
R13572 gnd.n6105 gnd.n2501 240.244
R13573 gnd.n6097 gnd.n2501 240.244
R13574 gnd.n6097 gnd.n2517 240.244
R13575 gnd.n6093 gnd.n2517 240.244
R13576 gnd.n6093 gnd.n2522 240.244
R13577 gnd.n6085 gnd.n2522 240.244
R13578 gnd.n6407 gnd.n671 240.244
R13579 gnd.n6407 gnd.n669 240.244
R13580 gnd.n6411 gnd.n669 240.244
R13581 gnd.n6411 gnd.n665 240.244
R13582 gnd.n6417 gnd.n665 240.244
R13583 gnd.n6417 gnd.n663 240.244
R13584 gnd.n6421 gnd.n663 240.244
R13585 gnd.n6421 gnd.n659 240.244
R13586 gnd.n6427 gnd.n659 240.244
R13587 gnd.n6427 gnd.n657 240.244
R13588 gnd.n6431 gnd.n657 240.244
R13589 gnd.n6431 gnd.n653 240.244
R13590 gnd.n6437 gnd.n653 240.244
R13591 gnd.n6437 gnd.n651 240.244
R13592 gnd.n6441 gnd.n651 240.244
R13593 gnd.n6441 gnd.n647 240.244
R13594 gnd.n6447 gnd.n647 240.244
R13595 gnd.n6447 gnd.n645 240.244
R13596 gnd.n6451 gnd.n645 240.244
R13597 gnd.n6451 gnd.n641 240.244
R13598 gnd.n6457 gnd.n641 240.244
R13599 gnd.n6457 gnd.n639 240.244
R13600 gnd.n6461 gnd.n639 240.244
R13601 gnd.n6461 gnd.n635 240.244
R13602 gnd.n6467 gnd.n635 240.244
R13603 gnd.n6467 gnd.n633 240.244
R13604 gnd.n6471 gnd.n633 240.244
R13605 gnd.n6471 gnd.n629 240.244
R13606 gnd.n6477 gnd.n629 240.244
R13607 gnd.n6477 gnd.n627 240.244
R13608 gnd.n6481 gnd.n627 240.244
R13609 gnd.n6481 gnd.n623 240.244
R13610 gnd.n6487 gnd.n623 240.244
R13611 gnd.n6487 gnd.n621 240.244
R13612 gnd.n6491 gnd.n621 240.244
R13613 gnd.n6491 gnd.n617 240.244
R13614 gnd.n6497 gnd.n617 240.244
R13615 gnd.n6497 gnd.n615 240.244
R13616 gnd.n6501 gnd.n615 240.244
R13617 gnd.n6501 gnd.n611 240.244
R13618 gnd.n6507 gnd.n611 240.244
R13619 gnd.n6507 gnd.n609 240.244
R13620 gnd.n6511 gnd.n609 240.244
R13621 gnd.n6511 gnd.n605 240.244
R13622 gnd.n6517 gnd.n605 240.244
R13623 gnd.n6517 gnd.n603 240.244
R13624 gnd.n6521 gnd.n603 240.244
R13625 gnd.n6521 gnd.n599 240.244
R13626 gnd.n6527 gnd.n599 240.244
R13627 gnd.n6527 gnd.n597 240.244
R13628 gnd.n6531 gnd.n597 240.244
R13629 gnd.n6531 gnd.n593 240.244
R13630 gnd.n6537 gnd.n593 240.244
R13631 gnd.n6537 gnd.n591 240.244
R13632 gnd.n6541 gnd.n591 240.244
R13633 gnd.n6541 gnd.n587 240.244
R13634 gnd.n6547 gnd.n587 240.244
R13635 gnd.n6547 gnd.n585 240.244
R13636 gnd.n6551 gnd.n585 240.244
R13637 gnd.n6551 gnd.n581 240.244
R13638 gnd.n6557 gnd.n581 240.244
R13639 gnd.n6557 gnd.n579 240.244
R13640 gnd.n6561 gnd.n579 240.244
R13641 gnd.n6561 gnd.n575 240.244
R13642 gnd.n6567 gnd.n575 240.244
R13643 gnd.n6567 gnd.n573 240.244
R13644 gnd.n6571 gnd.n573 240.244
R13645 gnd.n6571 gnd.n569 240.244
R13646 gnd.n6577 gnd.n569 240.244
R13647 gnd.n6577 gnd.n567 240.244
R13648 gnd.n6581 gnd.n567 240.244
R13649 gnd.n6581 gnd.n563 240.244
R13650 gnd.n6587 gnd.n563 240.244
R13651 gnd.n6587 gnd.n561 240.244
R13652 gnd.n6591 gnd.n561 240.244
R13653 gnd.n6591 gnd.n557 240.244
R13654 gnd.n6597 gnd.n557 240.244
R13655 gnd.n6597 gnd.n555 240.244
R13656 gnd.n6601 gnd.n555 240.244
R13657 gnd.n6601 gnd.n551 240.244
R13658 gnd.n6607 gnd.n551 240.244
R13659 gnd.n6607 gnd.n549 240.244
R13660 gnd.n6611 gnd.n549 240.244
R13661 gnd.n6611 gnd.n545 240.244
R13662 gnd.n6617 gnd.n545 240.244
R13663 gnd.n6617 gnd.n543 240.244
R13664 gnd.n6621 gnd.n543 240.244
R13665 gnd.n6621 gnd.n539 240.244
R13666 gnd.n6627 gnd.n539 240.244
R13667 gnd.n6627 gnd.n537 240.244
R13668 gnd.n6631 gnd.n537 240.244
R13669 gnd.n6631 gnd.n533 240.244
R13670 gnd.n6637 gnd.n533 240.244
R13671 gnd.n6637 gnd.n531 240.244
R13672 gnd.n6641 gnd.n531 240.244
R13673 gnd.n6641 gnd.n527 240.244
R13674 gnd.n6647 gnd.n527 240.244
R13675 gnd.n6647 gnd.n525 240.244
R13676 gnd.n6651 gnd.n525 240.244
R13677 gnd.n6651 gnd.n521 240.244
R13678 gnd.n6657 gnd.n521 240.244
R13679 gnd.n6657 gnd.n519 240.244
R13680 gnd.n6661 gnd.n519 240.244
R13681 gnd.n6661 gnd.n515 240.244
R13682 gnd.n6667 gnd.n515 240.244
R13683 gnd.n6667 gnd.n513 240.244
R13684 gnd.n6671 gnd.n513 240.244
R13685 gnd.n6671 gnd.n509 240.244
R13686 gnd.n6677 gnd.n509 240.244
R13687 gnd.n6677 gnd.n507 240.244
R13688 gnd.n6681 gnd.n507 240.244
R13689 gnd.n6681 gnd.n503 240.244
R13690 gnd.n6687 gnd.n503 240.244
R13691 gnd.n6687 gnd.n501 240.244
R13692 gnd.n6691 gnd.n501 240.244
R13693 gnd.n6691 gnd.n497 240.244
R13694 gnd.n6697 gnd.n497 240.244
R13695 gnd.n6697 gnd.n495 240.244
R13696 gnd.n6701 gnd.n495 240.244
R13697 gnd.n6701 gnd.n491 240.244
R13698 gnd.n6707 gnd.n491 240.244
R13699 gnd.n6707 gnd.n489 240.244
R13700 gnd.n6711 gnd.n489 240.244
R13701 gnd.n6711 gnd.n485 240.244
R13702 gnd.n6717 gnd.n485 240.244
R13703 gnd.n6717 gnd.n483 240.244
R13704 gnd.n6721 gnd.n483 240.244
R13705 gnd.n6721 gnd.n479 240.244
R13706 gnd.n6727 gnd.n479 240.244
R13707 gnd.n6727 gnd.n477 240.244
R13708 gnd.n6731 gnd.n477 240.244
R13709 gnd.n6731 gnd.n473 240.244
R13710 gnd.n6737 gnd.n473 240.244
R13711 gnd.n6737 gnd.n471 240.244
R13712 gnd.n6741 gnd.n471 240.244
R13713 gnd.n6741 gnd.n467 240.244
R13714 gnd.n6747 gnd.n467 240.244
R13715 gnd.n6747 gnd.n465 240.244
R13716 gnd.n6751 gnd.n465 240.244
R13717 gnd.n6751 gnd.n461 240.244
R13718 gnd.n6757 gnd.n461 240.244
R13719 gnd.n6757 gnd.n459 240.244
R13720 gnd.n6761 gnd.n459 240.244
R13721 gnd.n6761 gnd.n455 240.244
R13722 gnd.n6767 gnd.n455 240.244
R13723 gnd.n6767 gnd.n453 240.244
R13724 gnd.n6771 gnd.n453 240.244
R13725 gnd.n6771 gnd.n449 240.244
R13726 gnd.n6777 gnd.n449 240.244
R13727 gnd.n6777 gnd.n447 240.244
R13728 gnd.n6781 gnd.n447 240.244
R13729 gnd.n6781 gnd.n443 240.244
R13730 gnd.n6787 gnd.n443 240.244
R13731 gnd.n6787 gnd.n441 240.244
R13732 gnd.n6791 gnd.n441 240.244
R13733 gnd.n6791 gnd.n437 240.244
R13734 gnd.n6797 gnd.n437 240.244
R13735 gnd.n6797 gnd.n435 240.244
R13736 gnd.n6801 gnd.n435 240.244
R13737 gnd.n6801 gnd.n431 240.244
R13738 gnd.n6807 gnd.n431 240.244
R13739 gnd.n6807 gnd.n429 240.244
R13740 gnd.n6811 gnd.n429 240.244
R13741 gnd.n6811 gnd.n425 240.244
R13742 gnd.n6817 gnd.n425 240.244
R13743 gnd.n6817 gnd.n423 240.244
R13744 gnd.n6821 gnd.n423 240.244
R13745 gnd.n6821 gnd.n419 240.244
R13746 gnd.n6827 gnd.n419 240.244
R13747 gnd.n6827 gnd.n417 240.244
R13748 gnd.n6831 gnd.n417 240.244
R13749 gnd.n6831 gnd.n413 240.244
R13750 gnd.n6837 gnd.n413 240.244
R13751 gnd.n6837 gnd.n411 240.244
R13752 gnd.n6841 gnd.n411 240.244
R13753 gnd.n6841 gnd.n407 240.244
R13754 gnd.n6847 gnd.n407 240.244
R13755 gnd.n6847 gnd.n405 240.244
R13756 gnd.n6851 gnd.n405 240.244
R13757 gnd.n6851 gnd.n401 240.244
R13758 gnd.n6857 gnd.n401 240.244
R13759 gnd.n6857 gnd.n399 240.244
R13760 gnd.n6861 gnd.n399 240.244
R13761 gnd.n6861 gnd.n395 240.244
R13762 gnd.n6867 gnd.n395 240.244
R13763 gnd.n6867 gnd.n393 240.244
R13764 gnd.n6871 gnd.n393 240.244
R13765 gnd.n6871 gnd.n389 240.244
R13766 gnd.n6877 gnd.n389 240.244
R13767 gnd.n6877 gnd.n387 240.244
R13768 gnd.n6881 gnd.n387 240.244
R13769 gnd.n6881 gnd.n383 240.244
R13770 gnd.n6888 gnd.n383 240.244
R13771 gnd.n6888 gnd.n381 240.244
R13772 gnd.n6892 gnd.n378 240.244
R13773 gnd.n6898 gnd.n378 240.244
R13774 gnd.n6898 gnd.n376 240.244
R13775 gnd.n6902 gnd.n376 240.244
R13776 gnd.n6902 gnd.n372 240.244
R13777 gnd.n6908 gnd.n372 240.244
R13778 gnd.n6908 gnd.n370 240.244
R13779 gnd.n6912 gnd.n370 240.244
R13780 gnd.n6912 gnd.n366 240.244
R13781 gnd.n6918 gnd.n366 240.244
R13782 gnd.n6918 gnd.n364 240.244
R13783 gnd.n6922 gnd.n364 240.244
R13784 gnd.n6922 gnd.n360 240.244
R13785 gnd.n6928 gnd.n360 240.244
R13786 gnd.n6928 gnd.n358 240.244
R13787 gnd.n6932 gnd.n358 240.244
R13788 gnd.n6932 gnd.n354 240.244
R13789 gnd.n6938 gnd.n354 240.244
R13790 gnd.n6938 gnd.n352 240.244
R13791 gnd.n6942 gnd.n352 240.244
R13792 gnd.n6942 gnd.n348 240.244
R13793 gnd.n6948 gnd.n348 240.244
R13794 gnd.n6948 gnd.n346 240.244
R13795 gnd.n6952 gnd.n346 240.244
R13796 gnd.n6952 gnd.n342 240.244
R13797 gnd.n6958 gnd.n342 240.244
R13798 gnd.n6958 gnd.n340 240.244
R13799 gnd.n6962 gnd.n340 240.244
R13800 gnd.n6962 gnd.n336 240.244
R13801 gnd.n6968 gnd.n336 240.244
R13802 gnd.n6968 gnd.n334 240.244
R13803 gnd.n6972 gnd.n334 240.244
R13804 gnd.n6972 gnd.n330 240.244
R13805 gnd.n6978 gnd.n330 240.244
R13806 gnd.n6978 gnd.n328 240.244
R13807 gnd.n6982 gnd.n328 240.244
R13808 gnd.n6982 gnd.n324 240.244
R13809 gnd.n6988 gnd.n324 240.244
R13810 gnd.n6988 gnd.n322 240.244
R13811 gnd.n6992 gnd.n322 240.244
R13812 gnd.n6992 gnd.n318 240.244
R13813 gnd.n6998 gnd.n318 240.244
R13814 gnd.n6998 gnd.n316 240.244
R13815 gnd.n7002 gnd.n316 240.244
R13816 gnd.n7002 gnd.n312 240.244
R13817 gnd.n7008 gnd.n312 240.244
R13818 gnd.n7008 gnd.n310 240.244
R13819 gnd.n7012 gnd.n310 240.244
R13820 gnd.n7012 gnd.n306 240.244
R13821 gnd.n7018 gnd.n306 240.244
R13822 gnd.n7018 gnd.n304 240.244
R13823 gnd.n7022 gnd.n304 240.244
R13824 gnd.n7022 gnd.n300 240.244
R13825 gnd.n7028 gnd.n300 240.244
R13826 gnd.n7028 gnd.n298 240.244
R13827 gnd.n7032 gnd.n298 240.244
R13828 gnd.n7032 gnd.n294 240.244
R13829 gnd.n7038 gnd.n294 240.244
R13830 gnd.n7038 gnd.n292 240.244
R13831 gnd.n7042 gnd.n292 240.244
R13832 gnd.n7042 gnd.n288 240.244
R13833 gnd.n7048 gnd.n288 240.244
R13834 gnd.n7048 gnd.n286 240.244
R13835 gnd.n7052 gnd.n286 240.244
R13836 gnd.n7052 gnd.n282 240.244
R13837 gnd.n7058 gnd.n282 240.244
R13838 gnd.n7058 gnd.n280 240.244
R13839 gnd.n7062 gnd.n280 240.244
R13840 gnd.n7062 gnd.n276 240.244
R13841 gnd.n7068 gnd.n276 240.244
R13842 gnd.n7068 gnd.n274 240.244
R13843 gnd.n7072 gnd.n274 240.244
R13844 gnd.n7072 gnd.n270 240.244
R13845 gnd.n7078 gnd.n270 240.244
R13846 gnd.n7078 gnd.n268 240.244
R13847 gnd.n7082 gnd.n268 240.244
R13848 gnd.n7082 gnd.n264 240.244
R13849 gnd.n7088 gnd.n264 240.244
R13850 gnd.n7088 gnd.n262 240.244
R13851 gnd.n7092 gnd.n262 240.244
R13852 gnd.n7092 gnd.n258 240.244
R13853 gnd.n7098 gnd.n258 240.244
R13854 gnd.n7098 gnd.n256 240.244
R13855 gnd.n7102 gnd.n256 240.244
R13856 gnd.n6229 gnd.n841 240.244
R13857 gnd.n6229 gnd.n2306 240.244
R13858 gnd.n6225 gnd.n2306 240.244
R13859 gnd.n6225 gnd.n2313 240.244
R13860 gnd.n6221 gnd.n2313 240.244
R13861 gnd.n6221 gnd.n2315 240.244
R13862 gnd.n6217 gnd.n2315 240.244
R13863 gnd.n6217 gnd.n2321 240.244
R13864 gnd.n3736 gnd.n2321 240.244
R13865 gnd.n3742 gnd.n3736 240.244
R13866 gnd.n3743 gnd.n3742 240.244
R13867 gnd.n3744 gnd.n3743 240.244
R13868 gnd.n3744 gnd.n3731 240.244
R13869 gnd.n3811 gnd.n3731 240.244
R13870 gnd.n3811 gnd.n3732 240.244
R13871 gnd.n3807 gnd.n3732 240.244
R13872 gnd.n3807 gnd.n3806 240.244
R13873 gnd.n3806 gnd.n3805 240.244
R13874 gnd.n3805 gnd.n3752 240.244
R13875 gnd.n3801 gnd.n3752 240.244
R13876 gnd.n3801 gnd.n3800 240.244
R13877 gnd.n3800 gnd.n3799 240.244
R13878 gnd.n3799 gnd.n3758 240.244
R13879 gnd.n3762 gnd.n3758 240.244
R13880 gnd.n3769 gnd.n3762 240.244
R13881 gnd.n3791 gnd.n3769 240.244
R13882 gnd.n3791 gnd.n3790 240.244
R13883 gnd.n3790 gnd.n3789 240.244
R13884 gnd.n3789 gnd.n3787 240.244
R13885 gnd.n3787 gnd.n3784 240.244
R13886 gnd.n3784 gnd.n3783 240.244
R13887 gnd.n3783 gnd.n3780 240.244
R13888 gnd.n3780 gnd.n3779 240.244
R13889 gnd.n3779 gnd.n3770 240.244
R13890 gnd.n3775 gnd.n3770 240.244
R13891 gnd.n3775 gnd.n3774 240.244
R13892 gnd.n3774 gnd.n3688 240.244
R13893 gnd.n4247 gnd.n3688 240.244
R13894 gnd.n4247 gnd.n3684 240.244
R13895 gnd.n4253 gnd.n3684 240.244
R13896 gnd.n4254 gnd.n4253 240.244
R13897 gnd.n4255 gnd.n4254 240.244
R13898 gnd.n4255 gnd.n3680 240.244
R13899 gnd.n4261 gnd.n3680 240.244
R13900 gnd.n4262 gnd.n4261 240.244
R13901 gnd.n4263 gnd.n4262 240.244
R13902 gnd.n4263 gnd.n3676 240.244
R13903 gnd.n4269 gnd.n3676 240.244
R13904 gnd.n4270 gnd.n4269 240.244
R13905 gnd.n4271 gnd.n4270 240.244
R13906 gnd.n4271 gnd.n3672 240.244
R13907 gnd.n4278 gnd.n3672 240.244
R13908 gnd.n4278 gnd.n2565 240.244
R13909 gnd.n6068 gnd.n2565 240.244
R13910 gnd.n6068 gnd.n2566 240.244
R13911 gnd.n6064 gnd.n2566 240.244
R13912 gnd.n6064 gnd.n2572 240.244
R13913 gnd.n3451 gnd.n2572 240.244
R13914 gnd.n3457 gnd.n3451 240.244
R13915 gnd.n3457 gnd.n3448 240.244
R13916 gnd.n3463 gnd.n3448 240.244
R13917 gnd.n3463 gnd.n3444 240.244
R13918 gnd.n3469 gnd.n3444 240.244
R13919 gnd.n3469 gnd.n3442 240.244
R13920 gnd.n3475 gnd.n3442 240.244
R13921 gnd.n3475 gnd.n3437 240.244
R13922 gnd.n3483 gnd.n3437 240.244
R13923 gnd.n3483 gnd.n3438 240.244
R13924 gnd.n3438 gnd.n3221 240.244
R13925 gnd.n4557 gnd.n3221 240.244
R13926 gnd.n4557 gnd.n3216 240.244
R13927 gnd.n4565 gnd.n3216 240.244
R13928 gnd.n4565 gnd.n3217 240.244
R13929 gnd.n3217 gnd.n3197 240.244
R13930 gnd.n4595 gnd.n3197 240.244
R13931 gnd.n4595 gnd.n3192 240.244
R13932 gnd.n4606 gnd.n3192 240.244
R13933 gnd.n4606 gnd.n3193 240.244
R13934 gnd.n4602 gnd.n3193 240.244
R13935 gnd.n4602 gnd.n3172 240.244
R13936 gnd.n4635 gnd.n3172 240.244
R13937 gnd.n4635 gnd.n3167 240.244
R13938 gnd.n4643 gnd.n3167 240.244
R13939 gnd.n4643 gnd.n3168 240.244
R13940 gnd.n3168 gnd.n3144 240.244
R13941 gnd.n4671 gnd.n3144 240.244
R13942 gnd.n4671 gnd.n3140 240.244
R13943 gnd.n4677 gnd.n3140 240.244
R13944 gnd.n4677 gnd.n3126 240.244
R13945 gnd.n4697 gnd.n3126 240.244
R13946 gnd.n4697 gnd.n3121 240.244
R13947 gnd.n4705 gnd.n3121 240.244
R13948 gnd.n4705 gnd.n3122 240.244
R13949 gnd.n3122 gnd.n3100 240.244
R13950 gnd.n4753 gnd.n3100 240.244
R13951 gnd.n4753 gnd.n3093 240.244
R13952 gnd.n4761 gnd.n3093 240.244
R13953 gnd.n4761 gnd.n3096 240.244
R13954 gnd.n3096 gnd.n3075 240.244
R13955 gnd.n4793 gnd.n3075 240.244
R13956 gnd.n4793 gnd.n3070 240.244
R13957 gnd.n4801 gnd.n3070 240.244
R13958 gnd.n4801 gnd.n3071 240.244
R13959 gnd.n3071 gnd.n3045 240.244
R13960 gnd.n4862 gnd.n3045 240.244
R13961 gnd.n4862 gnd.n3040 240.244
R13962 gnd.n4870 gnd.n3040 240.244
R13963 gnd.n4870 gnd.n3041 240.244
R13964 gnd.n3041 gnd.n3021 240.244
R13965 gnd.n4895 gnd.n3021 240.244
R13966 gnd.n4895 gnd.n3016 240.244
R13967 gnd.n4903 gnd.n3016 240.244
R13968 gnd.n4903 gnd.n3017 240.244
R13969 gnd.n3017 gnd.n3000 240.244
R13970 gnd.n4949 gnd.n3000 240.244
R13971 gnd.n4949 gnd.n2995 240.244
R13972 gnd.n4957 gnd.n2995 240.244
R13973 gnd.n4957 gnd.n2996 240.244
R13974 gnd.n2996 gnd.n2975 240.244
R13975 gnd.n4986 gnd.n2975 240.244
R13976 gnd.n4986 gnd.n2971 240.244
R13977 gnd.n4992 gnd.n2971 240.244
R13978 gnd.n4992 gnd.n2884 240.244
R13979 gnd.n5129 gnd.n2884 240.244
R13980 gnd.n5129 gnd.n2880 240.244
R13981 gnd.n5135 gnd.n2880 240.244
R13982 gnd.n5135 gnd.n2871 240.244
R13983 gnd.n5145 gnd.n2871 240.244
R13984 gnd.n5145 gnd.n2867 240.244
R13985 gnd.n5151 gnd.n2867 240.244
R13986 gnd.n5151 gnd.n2858 240.244
R13987 gnd.n5161 gnd.n2858 240.244
R13988 gnd.n5161 gnd.n2854 240.244
R13989 gnd.n5167 gnd.n2854 240.244
R13990 gnd.n5167 gnd.n2844 240.244
R13991 gnd.n5178 gnd.n2844 240.244
R13992 gnd.n5178 gnd.n2840 240.244
R13993 gnd.n5185 gnd.n2840 240.244
R13994 gnd.n5185 gnd.n2699 240.244
R13995 gnd.n5933 gnd.n2699 240.244
R13996 gnd.n5933 gnd.n2700 240.244
R13997 gnd.n5929 gnd.n2700 240.244
R13998 gnd.n5929 gnd.n2706 240.244
R13999 gnd.n5463 gnd.n2706 240.244
R14000 gnd.n5464 gnd.n5463 240.244
R14001 gnd.n5464 gnd.n5458 240.244
R14002 gnd.n5470 gnd.n5458 240.244
R14003 gnd.n5471 gnd.n5470 240.244
R14004 gnd.n5472 gnd.n5471 240.244
R14005 gnd.n5472 gnd.n5454 240.244
R14006 gnd.n5541 gnd.n5454 240.244
R14007 gnd.n5542 gnd.n5541 240.244
R14008 gnd.n5543 gnd.n5542 240.244
R14009 gnd.n5543 gnd.n5450 240.244
R14010 gnd.n5549 gnd.n5450 240.244
R14011 gnd.n5550 gnd.n5549 240.244
R14012 gnd.n5551 gnd.n5550 240.244
R14013 gnd.n5551 gnd.n5445 240.244
R14014 gnd.n5562 gnd.n5445 240.244
R14015 gnd.n5562 gnd.n5446 240.244
R14016 gnd.n5558 gnd.n5446 240.244
R14017 gnd.n5558 gnd.n5408 240.244
R14018 gnd.n5749 gnd.n5408 240.244
R14019 gnd.n5749 gnd.n5409 240.244
R14020 gnd.n5744 gnd.n5409 240.244
R14021 gnd.n5744 gnd.n5412 240.244
R14022 gnd.n5597 gnd.n5412 240.244
R14023 gnd.n5597 gnd.n5426 240.244
R14024 gnd.n5727 gnd.n5426 240.244
R14025 gnd.n5727 gnd.n5427 240.244
R14026 gnd.n5722 gnd.n5427 240.244
R14027 gnd.n5722 gnd.n5721 240.244
R14028 gnd.n5721 gnd.n5431 240.244
R14029 gnd.n5658 gnd.n5431 240.244
R14030 gnd.n5658 gnd.n5653 240.244
R14031 gnd.n5664 gnd.n5653 240.244
R14032 gnd.n5665 gnd.n5664 240.244
R14033 gnd.n5666 gnd.n5665 240.244
R14034 gnd.n5666 gnd.n5648 240.244
R14035 gnd.n5693 gnd.n5648 240.244
R14036 gnd.n5693 gnd.n5649 240.244
R14037 gnd.n5689 gnd.n5649 240.244
R14038 gnd.n5689 gnd.n5688 240.244
R14039 gnd.n5688 gnd.n5687 240.244
R14040 gnd.n5687 gnd.n5674 240.244
R14041 gnd.n5683 gnd.n5674 240.244
R14042 gnd.n5683 gnd.n5682 240.244
R14043 gnd.n5682 gnd.n242 240.244
R14044 gnd.n7116 gnd.n242 240.244
R14045 gnd.n7116 gnd.n243 240.244
R14046 gnd.n7112 gnd.n243 240.244
R14047 gnd.n7112 gnd.n249 240.244
R14048 gnd.n7108 gnd.n249 240.244
R14049 gnd.n7108 gnd.n251 240.244
R14050 gnd.n6401 gnd.n675 240.244
R14051 gnd.n6397 gnd.n675 240.244
R14052 gnd.n6397 gnd.n677 240.244
R14053 gnd.n6393 gnd.n677 240.244
R14054 gnd.n6393 gnd.n682 240.244
R14055 gnd.n6389 gnd.n682 240.244
R14056 gnd.n6389 gnd.n684 240.244
R14057 gnd.n6385 gnd.n684 240.244
R14058 gnd.n6385 gnd.n690 240.244
R14059 gnd.n6381 gnd.n690 240.244
R14060 gnd.n6381 gnd.n692 240.244
R14061 gnd.n6377 gnd.n692 240.244
R14062 gnd.n6377 gnd.n698 240.244
R14063 gnd.n6373 gnd.n698 240.244
R14064 gnd.n6373 gnd.n700 240.244
R14065 gnd.n6369 gnd.n700 240.244
R14066 gnd.n6369 gnd.n706 240.244
R14067 gnd.n6365 gnd.n706 240.244
R14068 gnd.n6365 gnd.n708 240.244
R14069 gnd.n6361 gnd.n708 240.244
R14070 gnd.n6361 gnd.n714 240.244
R14071 gnd.n6357 gnd.n714 240.244
R14072 gnd.n6357 gnd.n716 240.244
R14073 gnd.n6353 gnd.n716 240.244
R14074 gnd.n6353 gnd.n722 240.244
R14075 gnd.n6349 gnd.n722 240.244
R14076 gnd.n6349 gnd.n724 240.244
R14077 gnd.n6345 gnd.n724 240.244
R14078 gnd.n6345 gnd.n730 240.244
R14079 gnd.n6341 gnd.n730 240.244
R14080 gnd.n6341 gnd.n732 240.244
R14081 gnd.n6337 gnd.n732 240.244
R14082 gnd.n6337 gnd.n738 240.244
R14083 gnd.n6333 gnd.n738 240.244
R14084 gnd.n6333 gnd.n740 240.244
R14085 gnd.n6329 gnd.n740 240.244
R14086 gnd.n6329 gnd.n746 240.244
R14087 gnd.n6325 gnd.n746 240.244
R14088 gnd.n6325 gnd.n748 240.244
R14089 gnd.n6321 gnd.n748 240.244
R14090 gnd.n6321 gnd.n754 240.244
R14091 gnd.n6317 gnd.n754 240.244
R14092 gnd.n6317 gnd.n756 240.244
R14093 gnd.n6313 gnd.n756 240.244
R14094 gnd.n6313 gnd.n762 240.244
R14095 gnd.n6309 gnd.n762 240.244
R14096 gnd.n6309 gnd.n764 240.244
R14097 gnd.n6305 gnd.n764 240.244
R14098 gnd.n6305 gnd.n770 240.244
R14099 gnd.n6301 gnd.n770 240.244
R14100 gnd.n6301 gnd.n772 240.244
R14101 gnd.n6297 gnd.n772 240.244
R14102 gnd.n6297 gnd.n778 240.244
R14103 gnd.n6293 gnd.n778 240.244
R14104 gnd.n6293 gnd.n780 240.244
R14105 gnd.n6289 gnd.n780 240.244
R14106 gnd.n6289 gnd.n786 240.244
R14107 gnd.n6285 gnd.n786 240.244
R14108 gnd.n6285 gnd.n788 240.244
R14109 gnd.n6281 gnd.n788 240.244
R14110 gnd.n6281 gnd.n794 240.244
R14111 gnd.n6277 gnd.n794 240.244
R14112 gnd.n6277 gnd.n796 240.244
R14113 gnd.n6273 gnd.n796 240.244
R14114 gnd.n6273 gnd.n802 240.244
R14115 gnd.n6269 gnd.n802 240.244
R14116 gnd.n6269 gnd.n804 240.244
R14117 gnd.n6265 gnd.n804 240.244
R14118 gnd.n6265 gnd.n810 240.244
R14119 gnd.n6261 gnd.n810 240.244
R14120 gnd.n6261 gnd.n812 240.244
R14121 gnd.n6257 gnd.n812 240.244
R14122 gnd.n6257 gnd.n818 240.244
R14123 gnd.n6253 gnd.n818 240.244
R14124 gnd.n6253 gnd.n820 240.244
R14125 gnd.n6249 gnd.n820 240.244
R14126 gnd.n6249 gnd.n826 240.244
R14127 gnd.n6245 gnd.n826 240.244
R14128 gnd.n6245 gnd.n828 240.244
R14129 gnd.n6241 gnd.n828 240.244
R14130 gnd.n6241 gnd.n834 240.244
R14131 gnd.n6237 gnd.n834 240.244
R14132 gnd.n6237 gnd.n836 240.244
R14133 gnd.n6233 gnd.n836 240.244
R14134 gnd.n2574 gnd.n2573 240.244
R14135 gnd.n3424 gnd.n2574 240.244
R14136 gnd.n3450 gnd.n3424 240.244
R14137 gnd.n3450 gnd.n3427 240.244
R14138 gnd.n3428 gnd.n3427 240.244
R14139 gnd.n3429 gnd.n3428 240.244
R14140 gnd.n3443 gnd.n3429 240.244
R14141 gnd.n3443 gnd.n3432 240.244
R14142 gnd.n3433 gnd.n3432 240.244
R14143 gnd.n3434 gnd.n3433 240.244
R14144 gnd.n3485 gnd.n3434 240.244
R14145 gnd.n3486 gnd.n3485 240.244
R14146 gnd.n3487 gnd.n3486 240.244
R14147 gnd.n3487 gnd.n3223 240.244
R14148 gnd.n3488 gnd.n3223 240.244
R14149 gnd.n3488 gnd.n3214 240.244
R14150 gnd.n3491 gnd.n3214 240.244
R14151 gnd.n3495 gnd.n3491 240.244
R14152 gnd.n3495 gnd.n3199 240.244
R14153 gnd.n3499 gnd.n3199 240.244
R14154 gnd.n3499 gnd.n3191 240.244
R14155 gnd.n3500 gnd.n3191 240.244
R14156 gnd.n3501 gnd.n3500 240.244
R14157 gnd.n3501 gnd.n3181 240.244
R14158 gnd.n3181 gnd.n3173 240.244
R14159 gnd.n3504 gnd.n3173 240.244
R14160 gnd.n3504 gnd.n3166 240.244
R14161 gnd.n3507 gnd.n3166 240.244
R14162 gnd.n3508 gnd.n3507 240.244
R14163 gnd.n3508 gnd.n3146 240.244
R14164 gnd.n3509 gnd.n3146 240.244
R14165 gnd.n3509 gnd.n3138 240.244
R14166 gnd.n3512 gnd.n3138 240.244
R14167 gnd.n3512 gnd.n3128 240.244
R14168 gnd.n3513 gnd.n3128 240.244
R14169 gnd.n3513 gnd.n3120 240.244
R14170 gnd.n3516 gnd.n3120 240.244
R14171 gnd.n3516 gnd.n3111 240.244
R14172 gnd.n3111 gnd.n3101 240.244
R14173 gnd.n3101 gnd.n3090 240.244
R14174 gnd.n4763 gnd.n3090 240.244
R14175 gnd.n4763 gnd.n3085 240.244
R14176 gnd.n4783 gnd.n3085 240.244
R14177 gnd.n4783 gnd.n3077 240.244
R14178 gnd.n4768 gnd.n3077 240.244
R14179 gnd.n4768 gnd.n3068 240.244
R14180 gnd.n4769 gnd.n3068 240.244
R14181 gnd.n4770 gnd.n4769 240.244
R14182 gnd.n4770 gnd.n3047 240.244
R14183 gnd.n3047 gnd.n3037 240.244
R14184 gnd.n4872 gnd.n3037 240.244
R14185 gnd.n4872 gnd.n3032 240.244
R14186 gnd.n4879 gnd.n3032 240.244
R14187 gnd.n4879 gnd.n3023 240.244
R14188 gnd.n3023 gnd.n3014 240.244
R14189 gnd.n4905 gnd.n3014 240.244
R14190 gnd.n4905 gnd.n3009 240.244
R14191 gnd.n4938 gnd.n3009 240.244
R14192 gnd.n4938 gnd.n3002 240.244
R14193 gnd.n4910 gnd.n3002 240.244
R14194 gnd.n4910 gnd.n2994 240.244
R14195 gnd.n4914 gnd.n2994 240.244
R14196 gnd.n4915 gnd.n4914 240.244
R14197 gnd.n4915 gnd.n2977 240.244
R14198 gnd.n4918 gnd.n2977 240.244
R14199 gnd.n4918 gnd.n2968 240.244
R14200 gnd.n4919 gnd.n2968 240.244
R14201 gnd.n4919 gnd.n2886 240.244
R14202 gnd.n2886 gnd.n2876 240.244
R14203 gnd.n5137 gnd.n2876 240.244
R14204 gnd.n5137 gnd.n2872 240.244
R14205 gnd.n5143 gnd.n2872 240.244
R14206 gnd.n5143 gnd.n2863 240.244
R14207 gnd.n5153 gnd.n2863 240.244
R14208 gnd.n5153 gnd.n2859 240.244
R14209 gnd.n5159 gnd.n2859 240.244
R14210 gnd.n5159 gnd.n2851 240.244
R14211 gnd.n5169 gnd.n2851 240.244
R14212 gnd.n5169 gnd.n2846 240.244
R14213 gnd.n5176 gnd.n2846 240.244
R14214 gnd.n5176 gnd.n2837 240.244
R14215 gnd.n5187 gnd.n2837 240.244
R14216 gnd.n3422 gnd.n3421 240.244
R14217 gnd.n3586 gnd.n3585 240.244
R14218 gnd.n3418 gnd.n3417 240.244
R14219 gnd.n3593 gnd.n3592 240.244
R14220 gnd.n3602 gnd.n3601 240.244
R14221 gnd.n3409 gnd.n3408 240.244
R14222 gnd.n3614 gnd.n3613 240.244
R14223 gnd.n3626 gnd.n3625 240.244
R14224 gnd.n3397 gnd.n3396 240.244
R14225 gnd.n3638 gnd.n3637 240.244
R14226 gnd.n3650 gnd.n3649 240.244
R14227 gnd.n3385 gnd.n3384 240.244
R14228 gnd.n3663 gnd.n3662 240.244
R14229 gnd.n6070 gnd.n2547 240.244
R14230 gnd.n6061 gnd.n2548 240.244
R14231 gnd.n6061 gnd.n2575 240.244
R14232 gnd.n2580 gnd.n2575 240.244
R14233 gnd.n2581 gnd.n2580 240.244
R14234 gnd.n2582 gnd.n2581 240.244
R14235 gnd.n3460 gnd.n2582 240.244
R14236 gnd.n3460 gnd.n2585 240.244
R14237 gnd.n2586 gnd.n2585 240.244
R14238 gnd.n2587 gnd.n2586 240.244
R14239 gnd.n3472 gnd.n2587 240.244
R14240 gnd.n3472 gnd.n2590 240.244
R14241 gnd.n2591 gnd.n2590 240.244
R14242 gnd.n2592 gnd.n2591 240.244
R14243 gnd.n4555 gnd.n2592 240.244
R14244 gnd.n4555 gnd.n2595 240.244
R14245 gnd.n2596 gnd.n2595 240.244
R14246 gnd.n2597 gnd.n2596 240.244
R14247 gnd.n3493 gnd.n2597 240.244
R14248 gnd.n3493 gnd.n2600 240.244
R14249 gnd.n2601 gnd.n2600 240.244
R14250 gnd.n2602 gnd.n2601 240.244
R14251 gnd.n3184 gnd.n2602 240.244
R14252 gnd.n3184 gnd.n2605 240.244
R14253 gnd.n2606 gnd.n2605 240.244
R14254 gnd.n2607 gnd.n2606 240.244
R14255 gnd.n3163 gnd.n2607 240.244
R14256 gnd.n3163 gnd.n2610 240.244
R14257 gnd.n2611 gnd.n2610 240.244
R14258 gnd.n2612 gnd.n2611 240.244
R14259 gnd.n4669 gnd.n2612 240.244
R14260 gnd.n4669 gnd.n2615 240.244
R14261 gnd.n2616 gnd.n2615 240.244
R14262 gnd.n2617 gnd.n2616 240.244
R14263 gnd.n4695 gnd.n2617 240.244
R14264 gnd.n4695 gnd.n2620 240.244
R14265 gnd.n2621 gnd.n2620 240.244
R14266 gnd.n2622 gnd.n2621 240.244
R14267 gnd.n4738 gnd.n2622 240.244
R14268 gnd.n4738 gnd.n2625 240.244
R14269 gnd.n2626 gnd.n2625 240.244
R14270 gnd.n2627 gnd.n2626 240.244
R14271 gnd.n3094 gnd.n2627 240.244
R14272 gnd.n3094 gnd.n2630 240.244
R14273 gnd.n2631 gnd.n2630 240.244
R14274 gnd.n2632 gnd.n2631 240.244
R14275 gnd.n3069 gnd.n2632 240.244
R14276 gnd.n3069 gnd.n2635 240.244
R14277 gnd.n2636 gnd.n2635 240.244
R14278 gnd.n2637 gnd.n2636 240.244
R14279 gnd.n3049 gnd.n2637 240.244
R14280 gnd.n3049 gnd.n2640 240.244
R14281 gnd.n2641 gnd.n2640 240.244
R14282 gnd.n2642 gnd.n2641 240.244
R14283 gnd.n4893 gnd.n2642 240.244
R14284 gnd.n4893 gnd.n2645 240.244
R14285 gnd.n2646 gnd.n2645 240.244
R14286 gnd.n2647 gnd.n2646 240.244
R14287 gnd.n4939 gnd.n2647 240.244
R14288 gnd.n4939 gnd.n2650 240.244
R14289 gnd.n2651 gnd.n2650 240.244
R14290 gnd.n2652 gnd.n2651 240.244
R14291 gnd.n4912 gnd.n2652 240.244
R14292 gnd.n4912 gnd.n2655 240.244
R14293 gnd.n2656 gnd.n2655 240.244
R14294 gnd.n2657 gnd.n2656 240.244
R14295 gnd.n2970 gnd.n2657 240.244
R14296 gnd.n2970 gnd.n2660 240.244
R14297 gnd.n2661 gnd.n2660 240.244
R14298 gnd.n2662 gnd.n2661 240.244
R14299 gnd.n2879 gnd.n2662 240.244
R14300 gnd.n2879 gnd.n2665 240.244
R14301 gnd.n2666 gnd.n2665 240.244
R14302 gnd.n2667 gnd.n2666 240.244
R14303 gnd.n2866 gnd.n2667 240.244
R14304 gnd.n2866 gnd.n2670 240.244
R14305 gnd.n2671 gnd.n2670 240.244
R14306 gnd.n2672 gnd.n2671 240.244
R14307 gnd.n2853 gnd.n2672 240.244
R14308 gnd.n2853 gnd.n2675 240.244
R14309 gnd.n2676 gnd.n2675 240.244
R14310 gnd.n2677 gnd.n2676 240.244
R14311 gnd.n2682 gnd.n2677 240.244
R14312 gnd.n2835 gnd.n2834 240.244
R14313 gnd.n5196 gnd.n5195 240.244
R14314 gnd.n2831 gnd.n2830 240.244
R14315 gnd.n5204 gnd.n5203 240.244
R14316 gnd.n5210 gnd.n5209 240.244
R14317 gnd.n5212 gnd.n5211 240.244
R14318 gnd.n5220 gnd.n5219 240.244
R14319 gnd.n5230 gnd.n5229 240.244
R14320 gnd.n5232 gnd.n5231 240.244
R14321 gnd.n5240 gnd.n5239 240.244
R14322 gnd.n5250 gnd.n5249 240.244
R14323 gnd.n5252 gnd.n5251 240.244
R14324 gnd.n5266 gnd.n5265 240.244
R14325 gnd.n5935 gnd.n2681 240.244
R14326 gnd.n3232 gnd.n3231 240.132
R14327 gnd.n2903 gnd.n2902 240.132
R14328 gnd.n6408 gnd.n670 225.874
R14329 gnd.n6409 gnd.n6408 225.874
R14330 gnd.n6410 gnd.n6409 225.874
R14331 gnd.n6410 gnd.n664 225.874
R14332 gnd.n6418 gnd.n664 225.874
R14333 gnd.n6419 gnd.n6418 225.874
R14334 gnd.n6420 gnd.n6419 225.874
R14335 gnd.n6420 gnd.n658 225.874
R14336 gnd.n6428 gnd.n658 225.874
R14337 gnd.n6429 gnd.n6428 225.874
R14338 gnd.n6430 gnd.n6429 225.874
R14339 gnd.n6430 gnd.n652 225.874
R14340 gnd.n6438 gnd.n652 225.874
R14341 gnd.n6439 gnd.n6438 225.874
R14342 gnd.n6440 gnd.n6439 225.874
R14343 gnd.n6440 gnd.n646 225.874
R14344 gnd.n6448 gnd.n646 225.874
R14345 gnd.n6449 gnd.n6448 225.874
R14346 gnd.n6450 gnd.n6449 225.874
R14347 gnd.n6450 gnd.n640 225.874
R14348 gnd.n6458 gnd.n640 225.874
R14349 gnd.n6459 gnd.n6458 225.874
R14350 gnd.n6460 gnd.n6459 225.874
R14351 gnd.n6460 gnd.n634 225.874
R14352 gnd.n6468 gnd.n634 225.874
R14353 gnd.n6469 gnd.n6468 225.874
R14354 gnd.n6470 gnd.n6469 225.874
R14355 gnd.n6470 gnd.n628 225.874
R14356 gnd.n6478 gnd.n628 225.874
R14357 gnd.n6479 gnd.n6478 225.874
R14358 gnd.n6480 gnd.n6479 225.874
R14359 gnd.n6480 gnd.n622 225.874
R14360 gnd.n6488 gnd.n622 225.874
R14361 gnd.n6489 gnd.n6488 225.874
R14362 gnd.n6490 gnd.n6489 225.874
R14363 gnd.n6490 gnd.n616 225.874
R14364 gnd.n6498 gnd.n616 225.874
R14365 gnd.n6499 gnd.n6498 225.874
R14366 gnd.n6500 gnd.n6499 225.874
R14367 gnd.n6500 gnd.n610 225.874
R14368 gnd.n6508 gnd.n610 225.874
R14369 gnd.n6509 gnd.n6508 225.874
R14370 gnd.n6510 gnd.n6509 225.874
R14371 gnd.n6510 gnd.n604 225.874
R14372 gnd.n6518 gnd.n604 225.874
R14373 gnd.n6519 gnd.n6518 225.874
R14374 gnd.n6520 gnd.n6519 225.874
R14375 gnd.n6520 gnd.n598 225.874
R14376 gnd.n6528 gnd.n598 225.874
R14377 gnd.n6529 gnd.n6528 225.874
R14378 gnd.n6530 gnd.n6529 225.874
R14379 gnd.n6530 gnd.n592 225.874
R14380 gnd.n6538 gnd.n592 225.874
R14381 gnd.n6539 gnd.n6538 225.874
R14382 gnd.n6540 gnd.n6539 225.874
R14383 gnd.n6540 gnd.n586 225.874
R14384 gnd.n6548 gnd.n586 225.874
R14385 gnd.n6549 gnd.n6548 225.874
R14386 gnd.n6550 gnd.n6549 225.874
R14387 gnd.n6550 gnd.n580 225.874
R14388 gnd.n6558 gnd.n580 225.874
R14389 gnd.n6559 gnd.n6558 225.874
R14390 gnd.n6560 gnd.n6559 225.874
R14391 gnd.n6560 gnd.n574 225.874
R14392 gnd.n6568 gnd.n574 225.874
R14393 gnd.n6569 gnd.n6568 225.874
R14394 gnd.n6570 gnd.n6569 225.874
R14395 gnd.n6570 gnd.n568 225.874
R14396 gnd.n6578 gnd.n568 225.874
R14397 gnd.n6579 gnd.n6578 225.874
R14398 gnd.n6580 gnd.n6579 225.874
R14399 gnd.n6580 gnd.n562 225.874
R14400 gnd.n6588 gnd.n562 225.874
R14401 gnd.n6589 gnd.n6588 225.874
R14402 gnd.n6590 gnd.n6589 225.874
R14403 gnd.n6590 gnd.n556 225.874
R14404 gnd.n6598 gnd.n556 225.874
R14405 gnd.n6599 gnd.n6598 225.874
R14406 gnd.n6600 gnd.n6599 225.874
R14407 gnd.n6600 gnd.n550 225.874
R14408 gnd.n6608 gnd.n550 225.874
R14409 gnd.n6609 gnd.n6608 225.874
R14410 gnd.n6610 gnd.n6609 225.874
R14411 gnd.n6610 gnd.n544 225.874
R14412 gnd.n6618 gnd.n544 225.874
R14413 gnd.n6619 gnd.n6618 225.874
R14414 gnd.n6620 gnd.n6619 225.874
R14415 gnd.n6620 gnd.n538 225.874
R14416 gnd.n6628 gnd.n538 225.874
R14417 gnd.n6629 gnd.n6628 225.874
R14418 gnd.n6630 gnd.n6629 225.874
R14419 gnd.n6630 gnd.n532 225.874
R14420 gnd.n6638 gnd.n532 225.874
R14421 gnd.n6639 gnd.n6638 225.874
R14422 gnd.n6640 gnd.n6639 225.874
R14423 gnd.n6640 gnd.n526 225.874
R14424 gnd.n6648 gnd.n526 225.874
R14425 gnd.n6649 gnd.n6648 225.874
R14426 gnd.n6650 gnd.n6649 225.874
R14427 gnd.n6650 gnd.n520 225.874
R14428 gnd.n6658 gnd.n520 225.874
R14429 gnd.n6659 gnd.n6658 225.874
R14430 gnd.n6660 gnd.n6659 225.874
R14431 gnd.n6660 gnd.n514 225.874
R14432 gnd.n6668 gnd.n514 225.874
R14433 gnd.n6669 gnd.n6668 225.874
R14434 gnd.n6670 gnd.n6669 225.874
R14435 gnd.n6670 gnd.n508 225.874
R14436 gnd.n6678 gnd.n508 225.874
R14437 gnd.n6679 gnd.n6678 225.874
R14438 gnd.n6680 gnd.n6679 225.874
R14439 gnd.n6680 gnd.n502 225.874
R14440 gnd.n6688 gnd.n502 225.874
R14441 gnd.n6689 gnd.n6688 225.874
R14442 gnd.n6690 gnd.n6689 225.874
R14443 gnd.n6690 gnd.n496 225.874
R14444 gnd.n6698 gnd.n496 225.874
R14445 gnd.n6699 gnd.n6698 225.874
R14446 gnd.n6700 gnd.n6699 225.874
R14447 gnd.n6700 gnd.n490 225.874
R14448 gnd.n6708 gnd.n490 225.874
R14449 gnd.n6709 gnd.n6708 225.874
R14450 gnd.n6710 gnd.n6709 225.874
R14451 gnd.n6710 gnd.n484 225.874
R14452 gnd.n6718 gnd.n484 225.874
R14453 gnd.n6719 gnd.n6718 225.874
R14454 gnd.n6720 gnd.n6719 225.874
R14455 gnd.n6720 gnd.n478 225.874
R14456 gnd.n6728 gnd.n478 225.874
R14457 gnd.n6729 gnd.n6728 225.874
R14458 gnd.n6730 gnd.n6729 225.874
R14459 gnd.n6730 gnd.n472 225.874
R14460 gnd.n6738 gnd.n472 225.874
R14461 gnd.n6739 gnd.n6738 225.874
R14462 gnd.n6740 gnd.n6739 225.874
R14463 gnd.n6740 gnd.n466 225.874
R14464 gnd.n6748 gnd.n466 225.874
R14465 gnd.n6749 gnd.n6748 225.874
R14466 gnd.n6750 gnd.n6749 225.874
R14467 gnd.n6750 gnd.n460 225.874
R14468 gnd.n6758 gnd.n460 225.874
R14469 gnd.n6759 gnd.n6758 225.874
R14470 gnd.n6760 gnd.n6759 225.874
R14471 gnd.n6760 gnd.n454 225.874
R14472 gnd.n6768 gnd.n454 225.874
R14473 gnd.n6769 gnd.n6768 225.874
R14474 gnd.n6770 gnd.n6769 225.874
R14475 gnd.n6770 gnd.n448 225.874
R14476 gnd.n6778 gnd.n448 225.874
R14477 gnd.n6779 gnd.n6778 225.874
R14478 gnd.n6780 gnd.n6779 225.874
R14479 gnd.n6780 gnd.n442 225.874
R14480 gnd.n6788 gnd.n442 225.874
R14481 gnd.n6789 gnd.n6788 225.874
R14482 gnd.n6790 gnd.n6789 225.874
R14483 gnd.n6790 gnd.n436 225.874
R14484 gnd.n6798 gnd.n436 225.874
R14485 gnd.n6799 gnd.n6798 225.874
R14486 gnd.n6800 gnd.n6799 225.874
R14487 gnd.n6800 gnd.n430 225.874
R14488 gnd.n6808 gnd.n430 225.874
R14489 gnd.n6809 gnd.n6808 225.874
R14490 gnd.n6810 gnd.n6809 225.874
R14491 gnd.n6810 gnd.n424 225.874
R14492 gnd.n6818 gnd.n424 225.874
R14493 gnd.n6819 gnd.n6818 225.874
R14494 gnd.n6820 gnd.n6819 225.874
R14495 gnd.n6820 gnd.n418 225.874
R14496 gnd.n6828 gnd.n418 225.874
R14497 gnd.n6829 gnd.n6828 225.874
R14498 gnd.n6830 gnd.n6829 225.874
R14499 gnd.n6830 gnd.n412 225.874
R14500 gnd.n6838 gnd.n412 225.874
R14501 gnd.n6839 gnd.n6838 225.874
R14502 gnd.n6840 gnd.n6839 225.874
R14503 gnd.n6840 gnd.n406 225.874
R14504 gnd.n6848 gnd.n406 225.874
R14505 gnd.n6849 gnd.n6848 225.874
R14506 gnd.n6850 gnd.n6849 225.874
R14507 gnd.n6850 gnd.n400 225.874
R14508 gnd.n6858 gnd.n400 225.874
R14509 gnd.n6859 gnd.n6858 225.874
R14510 gnd.n6860 gnd.n6859 225.874
R14511 gnd.n6860 gnd.n394 225.874
R14512 gnd.n6868 gnd.n394 225.874
R14513 gnd.n6869 gnd.n6868 225.874
R14514 gnd.n6870 gnd.n6869 225.874
R14515 gnd.n6870 gnd.n388 225.874
R14516 gnd.n6878 gnd.n388 225.874
R14517 gnd.n6879 gnd.n6878 225.874
R14518 gnd.n6880 gnd.n6879 225.874
R14519 gnd.n6880 gnd.n382 225.874
R14520 gnd.n6889 gnd.n382 225.874
R14521 gnd.n6890 gnd.n6889 225.874
R14522 gnd.n1396 gnd.t178 224.174
R14523 gnd.n907 gnd.t216 224.174
R14524 gnd.n2778 gnd.n2718 199.319
R14525 gnd.n2778 gnd.n2719 199.319
R14526 gnd.n4281 gnd.n3361 199.319
R14527 gnd.n4280 gnd.n3361 199.319
R14528 gnd.n3233 gnd.n3230 186.49
R14529 gnd.n2904 gnd.n2901 186.49
R14530 gnd.n2173 gnd.n2172 185
R14531 gnd.n2171 gnd.n2170 185
R14532 gnd.n2150 gnd.n2149 185
R14533 gnd.n2165 gnd.n2164 185
R14534 gnd.n2163 gnd.n2162 185
R14535 gnd.n2154 gnd.n2153 185
R14536 gnd.n2157 gnd.n2156 185
R14537 gnd.n2141 gnd.n2140 185
R14538 gnd.n2139 gnd.n2138 185
R14539 gnd.n2118 gnd.n2117 185
R14540 gnd.n2133 gnd.n2132 185
R14541 gnd.n2131 gnd.n2130 185
R14542 gnd.n2122 gnd.n2121 185
R14543 gnd.n2125 gnd.n2124 185
R14544 gnd.n2109 gnd.n2108 185
R14545 gnd.n2107 gnd.n2106 185
R14546 gnd.n2086 gnd.n2085 185
R14547 gnd.n2101 gnd.n2100 185
R14548 gnd.n2099 gnd.n2098 185
R14549 gnd.n2090 gnd.n2089 185
R14550 gnd.n2093 gnd.n2092 185
R14551 gnd.n2078 gnd.n2077 185
R14552 gnd.n2076 gnd.n2075 185
R14553 gnd.n2055 gnd.n2054 185
R14554 gnd.n2070 gnd.n2069 185
R14555 gnd.n2068 gnd.n2067 185
R14556 gnd.n2059 gnd.n2058 185
R14557 gnd.n2062 gnd.n2061 185
R14558 gnd.n2046 gnd.n2045 185
R14559 gnd.n2044 gnd.n2043 185
R14560 gnd.n2023 gnd.n2022 185
R14561 gnd.n2038 gnd.n2037 185
R14562 gnd.n2036 gnd.n2035 185
R14563 gnd.n2027 gnd.n2026 185
R14564 gnd.n2030 gnd.n2029 185
R14565 gnd.n2014 gnd.n2013 185
R14566 gnd.n2012 gnd.n2011 185
R14567 gnd.n1991 gnd.n1990 185
R14568 gnd.n2006 gnd.n2005 185
R14569 gnd.n2004 gnd.n2003 185
R14570 gnd.n1995 gnd.n1994 185
R14571 gnd.n1998 gnd.n1997 185
R14572 gnd.n1982 gnd.n1981 185
R14573 gnd.n1980 gnd.n1979 185
R14574 gnd.n1959 gnd.n1958 185
R14575 gnd.n1974 gnd.n1973 185
R14576 gnd.n1972 gnd.n1971 185
R14577 gnd.n1963 gnd.n1962 185
R14578 gnd.n1966 gnd.n1965 185
R14579 gnd.n1951 gnd.n1950 185
R14580 gnd.n1949 gnd.n1948 185
R14581 gnd.n1928 gnd.n1927 185
R14582 gnd.n1943 gnd.n1942 185
R14583 gnd.n1941 gnd.n1940 185
R14584 gnd.n1932 gnd.n1931 185
R14585 gnd.n1935 gnd.n1934 185
R14586 gnd.n1397 gnd.t177 178.987
R14587 gnd.n908 gnd.t217 178.987
R14588 gnd.n1 gnd.t157 170.774
R14589 gnd.n7 gnd.t147 170.103
R14590 gnd.n6 gnd.t312 170.103
R14591 gnd.n5 gnd.t149 170.103
R14592 gnd.n4 gnd.t135 170.103
R14593 gnd.n3 gnd.t314 170.103
R14594 gnd.n2 gnd.t137 170.103
R14595 gnd.n1 gnd.t161 170.103
R14596 gnd.n5121 gnd.n5120 163.367
R14597 gnd.n5118 gnd.n2913 163.367
R14598 gnd.n5114 gnd.n5113 163.367
R14599 gnd.n5111 gnd.n2916 163.367
R14600 gnd.n5107 gnd.n5106 163.367
R14601 gnd.n5104 gnd.n2919 163.367
R14602 gnd.n5100 gnd.n5099 163.367
R14603 gnd.n5097 gnd.n2922 163.367
R14604 gnd.n5093 gnd.n5092 163.367
R14605 gnd.n5090 gnd.n2925 163.367
R14606 gnd.n5086 gnd.n5085 163.367
R14607 gnd.n5083 gnd.n2928 163.367
R14608 gnd.n5079 gnd.n5078 163.367
R14609 gnd.n5076 gnd.n2931 163.367
R14610 gnd.n5071 gnd.n5070 163.367
R14611 gnd.n5068 gnd.n5066 163.367
R14612 gnd.n5063 gnd.n5062 163.367
R14613 gnd.n5060 gnd.n2937 163.367
R14614 gnd.n5055 gnd.n5054 163.367
R14615 gnd.n5052 gnd.n2942 163.367
R14616 gnd.n5048 gnd.n5047 163.367
R14617 gnd.n5045 gnd.n2945 163.367
R14618 gnd.n5041 gnd.n5040 163.367
R14619 gnd.n5038 gnd.n2948 163.367
R14620 gnd.n5034 gnd.n5033 163.367
R14621 gnd.n5031 gnd.n2951 163.367
R14622 gnd.n5027 gnd.n5026 163.367
R14623 gnd.n5024 gnd.n2954 163.367
R14624 gnd.n5020 gnd.n5019 163.367
R14625 gnd.n5017 gnd.n2957 163.367
R14626 gnd.n5013 gnd.n5012 163.367
R14627 gnd.n5010 gnd.n2960 163.367
R14628 gnd.n3294 gnd.n3224 163.367
R14629 gnd.n3290 gnd.n3224 163.367
R14630 gnd.n3290 gnd.n3213 163.367
R14631 gnd.n3213 gnd.n3207 163.367
R14632 gnd.n4574 gnd.n3207 163.367
R14633 gnd.n4574 gnd.n3204 163.367
R14634 gnd.n4586 gnd.n3204 163.367
R14635 gnd.n4586 gnd.n3205 163.367
R14636 gnd.n3205 gnd.n3200 163.367
R14637 gnd.n4581 gnd.n3200 163.367
R14638 gnd.n4581 gnd.n3190 163.367
R14639 gnd.n4578 gnd.n3190 163.367
R14640 gnd.n4578 gnd.n3183 163.367
R14641 gnd.n4616 gnd.n3183 163.367
R14642 gnd.n4616 gnd.n3180 163.367
R14643 gnd.n4624 gnd.n3180 163.367
R14644 gnd.n4624 gnd.n3174 163.367
R14645 gnd.n4620 gnd.n3174 163.367
R14646 gnd.n4620 gnd.n3165 163.367
R14647 gnd.n3165 gnd.n3156 163.367
R14648 gnd.n4651 gnd.n3156 163.367
R14649 gnd.n4651 gnd.n3153 163.367
R14650 gnd.n4661 gnd.n3153 163.367
R14651 gnd.n4661 gnd.n3154 163.367
R14652 gnd.n3154 gnd.n3147 163.367
R14653 gnd.n4656 gnd.n3147 163.367
R14654 gnd.n4656 gnd.n3137 163.367
R14655 gnd.n3137 gnd.n3131 163.367
R14656 gnd.n4687 gnd.n3131 163.367
R14657 gnd.n4687 gnd.n3129 163.367
R14658 gnd.n4693 gnd.n3129 163.367
R14659 gnd.n4693 gnd.n3119 163.367
R14660 gnd.n3119 gnd.n3113 163.367
R14661 gnd.n4715 gnd.n3113 163.367
R14662 gnd.n4716 gnd.n4715 163.367
R14663 gnd.n4716 gnd.n3110 163.367
R14664 gnd.n4736 gnd.n3110 163.367
R14665 gnd.n4736 gnd.n3102 163.367
R14666 gnd.n4732 gnd.n3102 163.367
R14667 gnd.n4732 gnd.n4731 163.367
R14668 gnd.n4731 gnd.n4730 163.367
R14669 gnd.n4730 gnd.n4720 163.367
R14670 gnd.n4720 gnd.n3084 163.367
R14671 gnd.n4725 gnd.n3084 163.367
R14672 gnd.n4725 gnd.n3078 163.367
R14673 gnd.n4722 gnd.n3078 163.367
R14674 gnd.n4722 gnd.n3067 163.367
R14675 gnd.n3067 gnd.n3059 163.367
R14676 gnd.n4810 gnd.n3059 163.367
R14677 gnd.n4810 gnd.n3056 163.367
R14678 gnd.n4848 gnd.n3056 163.367
R14679 gnd.n4848 gnd.n3057 163.367
R14680 gnd.n3057 gnd.n3048 163.367
R14681 gnd.n4843 gnd.n3048 163.367
R14682 gnd.n4843 gnd.n4841 163.367
R14683 gnd.n4841 gnd.n4840 163.367
R14684 gnd.n4840 gnd.n4816 163.367
R14685 gnd.n4816 gnd.n3031 163.367
R14686 gnd.n4835 gnd.n3031 163.367
R14687 gnd.n4835 gnd.n3024 163.367
R14688 gnd.n4832 gnd.n3024 163.367
R14689 gnd.n4832 gnd.n4831 163.367
R14690 gnd.n4831 gnd.n4830 163.367
R14691 gnd.n4830 gnd.n4820 163.367
R14692 gnd.n4820 gnd.n3008 163.367
R14693 gnd.n4825 gnd.n3008 163.367
R14694 gnd.n4825 gnd.n3003 163.367
R14695 gnd.n4822 gnd.n3003 163.367
R14696 gnd.n4822 gnd.n2993 163.367
R14697 gnd.n2993 gnd.n2987 163.367
R14698 gnd.n4966 gnd.n2987 163.367
R14699 gnd.n4966 gnd.n2984 163.367
R14700 gnd.n4977 gnd.n2984 163.367
R14701 gnd.n4977 gnd.n2985 163.367
R14702 gnd.n2985 gnd.n2978 163.367
R14703 gnd.n4972 gnd.n2978 163.367
R14704 gnd.n4972 gnd.n2967 163.367
R14705 gnd.n2967 gnd.n2962 163.367
R14706 gnd.n5001 gnd.n2962 163.367
R14707 gnd.n5002 gnd.n5001 163.367
R14708 gnd.n5002 gnd.n2887 163.367
R14709 gnd.n4545 gnd.n3247 163.367
R14710 gnd.n4545 gnd.n3282 163.367
R14711 gnd.n4541 gnd.n4540 163.367
R14712 gnd.n4537 gnd.n4536 163.367
R14713 gnd.n4533 gnd.n4532 163.367
R14714 gnd.n4529 gnd.n4528 163.367
R14715 gnd.n4525 gnd.n4524 163.367
R14716 gnd.n4521 gnd.n4520 163.367
R14717 gnd.n4517 gnd.n4516 163.367
R14718 gnd.n4513 gnd.n4512 163.367
R14719 gnd.n4509 gnd.n4508 163.367
R14720 gnd.n4505 gnd.n4504 163.367
R14721 gnd.n4501 gnd.n4500 163.367
R14722 gnd.n4497 gnd.n4496 163.367
R14723 gnd.n4493 gnd.n4492 163.367
R14724 gnd.n4489 gnd.n4488 163.367
R14725 gnd.n4485 gnd.n4484 163.367
R14726 gnd.n3356 gnd.n3355 163.367
R14727 gnd.n3351 gnd.n3350 163.367
R14728 gnd.n3347 gnd.n3346 163.367
R14729 gnd.n3343 gnd.n3342 163.367
R14730 gnd.n3339 gnd.n3338 163.367
R14731 gnd.n3335 gnd.n3334 163.367
R14732 gnd.n3331 gnd.n3330 163.367
R14733 gnd.n3327 gnd.n3326 163.367
R14734 gnd.n3323 gnd.n3322 163.367
R14735 gnd.n3319 gnd.n3318 163.367
R14736 gnd.n3315 gnd.n3314 163.367
R14737 gnd.n3311 gnd.n3310 163.367
R14738 gnd.n3307 gnd.n3306 163.367
R14739 gnd.n3303 gnd.n3302 163.367
R14740 gnd.n3299 gnd.n3298 163.367
R14741 gnd.n4553 gnd.n3225 163.367
R14742 gnd.n4553 gnd.n3211 163.367
R14743 gnd.n4568 gnd.n3211 163.367
R14744 gnd.n4568 gnd.n3209 163.367
R14745 gnd.n4572 gnd.n3209 163.367
R14746 gnd.n4572 gnd.n3203 163.367
R14747 gnd.n4588 gnd.n3203 163.367
R14748 gnd.n4588 gnd.n3201 163.367
R14749 gnd.n4592 gnd.n3201 163.367
R14750 gnd.n4592 gnd.n3188 163.367
R14751 gnd.n4609 gnd.n3188 163.367
R14752 gnd.n4609 gnd.n3186 163.367
R14753 gnd.n4613 gnd.n3186 163.367
R14754 gnd.n4613 gnd.n3178 163.367
R14755 gnd.n4628 gnd.n3178 163.367
R14756 gnd.n4628 gnd.n3176 163.367
R14757 gnd.n4632 gnd.n3176 163.367
R14758 gnd.n4632 gnd.n3162 163.367
R14759 gnd.n4645 gnd.n3162 163.367
R14760 gnd.n4645 gnd.n3160 163.367
R14761 gnd.n4649 gnd.n3160 163.367
R14762 gnd.n4649 gnd.n3151 163.367
R14763 gnd.n4663 gnd.n3151 163.367
R14764 gnd.n4663 gnd.n3149 163.367
R14765 gnd.n4667 gnd.n3149 163.367
R14766 gnd.n4667 gnd.n3136 163.367
R14767 gnd.n4680 gnd.n3136 163.367
R14768 gnd.n4680 gnd.n3133 163.367
R14769 gnd.n4685 gnd.n3133 163.367
R14770 gnd.n4685 gnd.n3134 163.367
R14771 gnd.n3134 gnd.n3117 163.367
R14772 gnd.n4709 gnd.n3117 163.367
R14773 gnd.n4709 gnd.n3115 163.367
R14774 gnd.n4713 gnd.n3115 163.367
R14775 gnd.n4713 gnd.n3108 163.367
R14776 gnd.n4741 gnd.n3108 163.367
R14777 gnd.n4741 gnd.n3105 163.367
R14778 gnd.n4750 gnd.n3105 163.367
R14779 gnd.n4750 gnd.n3106 163.367
R14780 gnd.n4746 gnd.n3106 163.367
R14781 gnd.n4746 gnd.n4745 163.367
R14782 gnd.n4745 gnd.n3082 163.367
R14783 gnd.n4786 gnd.n3082 163.367
R14784 gnd.n4786 gnd.n3080 163.367
R14785 gnd.n4790 gnd.n3080 163.367
R14786 gnd.n4790 gnd.n3065 163.367
R14787 gnd.n4804 gnd.n3065 163.367
R14788 gnd.n4804 gnd.n3063 163.367
R14789 gnd.n4808 gnd.n3063 163.367
R14790 gnd.n4808 gnd.n3054 163.367
R14791 gnd.n4850 gnd.n3054 163.367
R14792 gnd.n4850 gnd.n3051 163.367
R14793 gnd.n4859 gnd.n3051 163.367
R14794 gnd.n4859 gnd.n3052 163.367
R14795 gnd.n4855 gnd.n3052 163.367
R14796 gnd.n4855 gnd.n4854 163.367
R14797 gnd.n4854 gnd.n3030 163.367
R14798 gnd.n4882 gnd.n3030 163.367
R14799 gnd.n4882 gnd.n3027 163.367
R14800 gnd.n4891 gnd.n3027 163.367
R14801 gnd.n4891 gnd.n3028 163.367
R14802 gnd.n4887 gnd.n3028 163.367
R14803 gnd.n4887 gnd.n4886 163.367
R14804 gnd.n4886 gnd.n3007 163.367
R14805 gnd.n4942 gnd.n3007 163.367
R14806 gnd.n4942 gnd.n3005 163.367
R14807 gnd.n4946 gnd.n3005 163.367
R14808 gnd.n4946 gnd.n2991 163.367
R14809 gnd.n4960 gnd.n2991 163.367
R14810 gnd.n4960 gnd.n2989 163.367
R14811 gnd.n4964 gnd.n2989 163.367
R14812 gnd.n4964 gnd.n2982 163.367
R14813 gnd.n4979 gnd.n2982 163.367
R14814 gnd.n4979 gnd.n2980 163.367
R14815 gnd.n4983 gnd.n2980 163.367
R14816 gnd.n4983 gnd.n2966 163.367
R14817 gnd.n4995 gnd.n2966 163.367
R14818 gnd.n4995 gnd.n2964 163.367
R14819 gnd.n4999 gnd.n2964 163.367
R14820 gnd.n4999 gnd.n2889 163.367
R14821 gnd.n5126 gnd.n2889 163.367
R14822 gnd.n2910 gnd.n2909 156.462
R14823 gnd.n2113 gnd.n2081 153.042
R14824 gnd.n2177 gnd.n2176 152.079
R14825 gnd.n2145 gnd.n2144 152.079
R14826 gnd.n2113 gnd.n2112 152.079
R14827 gnd.n3238 gnd.n3237 152
R14828 gnd.n3239 gnd.n3228 152
R14829 gnd.n3241 gnd.n3240 152
R14830 gnd.n3243 gnd.n3226 152
R14831 gnd.n3245 gnd.n3244 152
R14832 gnd.n2908 gnd.n2892 152
R14833 gnd.n2900 gnd.n2893 152
R14834 gnd.n2899 gnd.n2898 152
R14835 gnd.n2897 gnd.n2894 152
R14836 gnd.n2895 gnd.t226 150.546
R14837 gnd.t144 gnd.n2155 147.661
R14838 gnd.t142 gnd.n2123 147.661
R14839 gnd.t316 gnd.n2091 147.661
R14840 gnd.t319 gnd.n2060 147.661
R14841 gnd.t159 gnd.n2028 147.661
R14842 gnd.t151 gnd.n1996 147.661
R14843 gnd.t154 gnd.n1964 147.661
R14844 gnd.t308 gnd.n1933 147.661
R14845 gnd.n5065 gnd.n5064 143.351
R14846 gnd.n4483 gnd.n3263 143.351
R14847 gnd.n4483 gnd.n3264 143.351
R14848 gnd.n3235 gnd.t278 130.484
R14849 gnd.n3244 gnd.t186 126.766
R14850 gnd.n3242 gnd.t248 126.766
R14851 gnd.n3228 gnd.t204 126.766
R14852 gnd.n3236 gnd.t229 126.766
R14853 gnd.n2896 gnd.t288 126.766
R14854 gnd.n2898 gnd.t245 126.766
R14855 gnd.n2907 gnd.t183 126.766
R14856 gnd.n2909 gnd.t263 126.766
R14857 gnd.n5874 gnd.n2777 108.609
R14858 gnd.n4486 gnd.n4482 108.609
R14859 gnd.n2172 gnd.n2171 104.615
R14860 gnd.n2171 gnd.n2149 104.615
R14861 gnd.n2164 gnd.n2149 104.615
R14862 gnd.n2164 gnd.n2163 104.615
R14863 gnd.n2163 gnd.n2153 104.615
R14864 gnd.n2156 gnd.n2153 104.615
R14865 gnd.n2140 gnd.n2139 104.615
R14866 gnd.n2139 gnd.n2117 104.615
R14867 gnd.n2132 gnd.n2117 104.615
R14868 gnd.n2132 gnd.n2131 104.615
R14869 gnd.n2131 gnd.n2121 104.615
R14870 gnd.n2124 gnd.n2121 104.615
R14871 gnd.n2108 gnd.n2107 104.615
R14872 gnd.n2107 gnd.n2085 104.615
R14873 gnd.n2100 gnd.n2085 104.615
R14874 gnd.n2100 gnd.n2099 104.615
R14875 gnd.n2099 gnd.n2089 104.615
R14876 gnd.n2092 gnd.n2089 104.615
R14877 gnd.n2077 gnd.n2076 104.615
R14878 gnd.n2076 gnd.n2054 104.615
R14879 gnd.n2069 gnd.n2054 104.615
R14880 gnd.n2069 gnd.n2068 104.615
R14881 gnd.n2068 gnd.n2058 104.615
R14882 gnd.n2061 gnd.n2058 104.615
R14883 gnd.n2045 gnd.n2044 104.615
R14884 gnd.n2044 gnd.n2022 104.615
R14885 gnd.n2037 gnd.n2022 104.615
R14886 gnd.n2037 gnd.n2036 104.615
R14887 gnd.n2036 gnd.n2026 104.615
R14888 gnd.n2029 gnd.n2026 104.615
R14889 gnd.n2013 gnd.n2012 104.615
R14890 gnd.n2012 gnd.n1990 104.615
R14891 gnd.n2005 gnd.n1990 104.615
R14892 gnd.n2005 gnd.n2004 104.615
R14893 gnd.n2004 gnd.n1994 104.615
R14894 gnd.n1997 gnd.n1994 104.615
R14895 gnd.n1981 gnd.n1980 104.615
R14896 gnd.n1980 gnd.n1958 104.615
R14897 gnd.n1973 gnd.n1958 104.615
R14898 gnd.n1973 gnd.n1972 104.615
R14899 gnd.n1972 gnd.n1962 104.615
R14900 gnd.n1965 gnd.n1962 104.615
R14901 gnd.n1950 gnd.n1949 104.615
R14902 gnd.n1949 gnd.n1927 104.615
R14903 gnd.n1942 gnd.n1927 104.615
R14904 gnd.n1942 gnd.n1941 104.615
R14905 gnd.n1941 gnd.n1931 104.615
R14906 gnd.n1934 gnd.n1931 104.615
R14907 gnd.n1322 gnd.t287 100.632
R14908 gnd.n881 gnd.t181 100.632
R14909 gnd.n7329 gnd.n7328 99.6594
R14910 gnd.n7324 gnd.n7145 99.6594
R14911 gnd.n7320 gnd.n7144 99.6594
R14912 gnd.n7316 gnd.n7143 99.6594
R14913 gnd.n7312 gnd.n7142 99.6594
R14914 gnd.n7308 gnd.n7141 99.6594
R14915 gnd.n7304 gnd.n7140 99.6594
R14916 gnd.n7300 gnd.n7139 99.6594
R14917 gnd.n7293 gnd.n7138 99.6594
R14918 gnd.n7289 gnd.n7137 99.6594
R14919 gnd.n7285 gnd.n7136 99.6594
R14920 gnd.n7281 gnd.n7135 99.6594
R14921 gnd.n7277 gnd.n7134 99.6594
R14922 gnd.n7273 gnd.n7133 99.6594
R14923 gnd.n7269 gnd.n7132 99.6594
R14924 gnd.n7265 gnd.n7131 99.6594
R14925 gnd.n7261 gnd.n7130 99.6594
R14926 gnd.n7257 gnd.n7129 99.6594
R14927 gnd.n7249 gnd.n7128 99.6594
R14928 gnd.n7247 gnd.n7127 99.6594
R14929 gnd.n7243 gnd.n7126 99.6594
R14930 gnd.n7239 gnd.n7125 99.6594
R14931 gnd.n7235 gnd.n7124 99.6594
R14932 gnd.n7231 gnd.n7123 99.6594
R14933 gnd.n7227 gnd.n7122 99.6594
R14934 gnd.n7223 gnd.n7121 99.6594
R14935 gnd.n7219 gnd.n7120 99.6594
R14936 gnd.n7215 gnd.n7119 99.6594
R14937 gnd.n7207 gnd.n7118 99.6594
R14938 gnd.n5926 gnd.n5925 99.6594
R14939 gnd.n5920 gnd.n2707 99.6594
R14940 gnd.n5917 gnd.n2708 99.6594
R14941 gnd.n5913 gnd.n2709 99.6594
R14942 gnd.n5909 gnd.n2710 99.6594
R14943 gnd.n5905 gnd.n2711 99.6594
R14944 gnd.n5901 gnd.n2712 99.6594
R14945 gnd.n5897 gnd.n2713 99.6594
R14946 gnd.n5893 gnd.n2714 99.6594
R14947 gnd.n5888 gnd.n2715 99.6594
R14948 gnd.n5884 gnd.n2716 99.6594
R14949 gnd.n5880 gnd.n2717 99.6594
R14950 gnd.n5876 gnd.n2718 99.6594
R14951 gnd.n5871 gnd.n2720 99.6594
R14952 gnd.n5867 gnd.n2721 99.6594
R14953 gnd.n5863 gnd.n2722 99.6594
R14954 gnd.n5859 gnd.n2723 99.6594
R14955 gnd.n5855 gnd.n2724 99.6594
R14956 gnd.n5851 gnd.n2725 99.6594
R14957 gnd.n5847 gnd.n2726 99.6594
R14958 gnd.n5843 gnd.n2727 99.6594
R14959 gnd.n5839 gnd.n2728 99.6594
R14960 gnd.n5835 gnd.n2729 99.6594
R14961 gnd.n5831 gnd.n2730 99.6594
R14962 gnd.n5827 gnd.n2731 99.6594
R14963 gnd.n5823 gnd.n2732 99.6594
R14964 gnd.n5819 gnd.n2733 99.6594
R14965 gnd.n5815 gnd.n2734 99.6594
R14966 gnd.n4371 gnd.n4370 99.6594
R14967 gnd.n4366 gnd.n4292 99.6594
R14968 gnd.n4362 gnd.n4291 99.6594
R14969 gnd.n4358 gnd.n4290 99.6594
R14970 gnd.n4354 gnd.n4289 99.6594
R14971 gnd.n4350 gnd.n4288 99.6594
R14972 gnd.n4346 gnd.n4287 99.6594
R14973 gnd.n4342 gnd.n4286 99.6594
R14974 gnd.n4337 gnd.n4285 99.6594
R14975 gnd.n4333 gnd.n4284 99.6594
R14976 gnd.n4329 gnd.n4283 99.6594
R14977 gnd.n4325 gnd.n4282 99.6594
R14978 gnd.n4280 gnd.n3365 99.6594
R14979 gnd.n4476 gnd.n4475 99.6594
R14980 gnd.n4473 gnd.n4472 99.6594
R14981 gnd.n4468 gnd.n4380 99.6594
R14982 gnd.n4466 gnd.n4465 99.6594
R14983 gnd.n4390 gnd.n4389 99.6594
R14984 gnd.n4457 gnd.n4456 99.6594
R14985 gnd.n4454 gnd.n4453 99.6594
R14986 gnd.n4449 gnd.n4398 99.6594
R14987 gnd.n4447 gnd.n4446 99.6594
R14988 gnd.n4442 gnd.n4405 99.6594
R14989 gnd.n4440 gnd.n4439 99.6594
R14990 gnd.n4435 gnd.n4412 99.6594
R14991 gnd.n4433 gnd.n4432 99.6594
R14992 gnd.n4428 gnd.n4421 99.6594
R14993 gnd.n4426 gnd.n4425 99.6594
R14994 gnd.n3958 gnd.n2327 99.6594
R14995 gnd.n3966 gnd.n3965 99.6594
R14996 gnd.n3969 gnd.n3968 99.6594
R14997 gnd.n3976 gnd.n3975 99.6594
R14998 gnd.n3979 gnd.n3978 99.6594
R14999 gnd.n3986 gnd.n3985 99.6594
R15000 gnd.n3989 gnd.n3988 99.6594
R15001 gnd.n3996 gnd.n3995 99.6594
R15002 gnd.n3999 gnd.n3998 99.6594
R15003 gnd.n4006 gnd.n4005 99.6594
R15004 gnd.n4009 gnd.n4008 99.6594
R15005 gnd.n4016 gnd.n4015 99.6594
R15006 gnd.n4019 gnd.n4018 99.6594
R15007 gnd.n4026 gnd.n4025 99.6594
R15008 gnd.n4029 gnd.n4028 99.6594
R15009 gnd.n4036 gnd.n4035 99.6594
R15010 gnd.n4039 gnd.n4038 99.6594
R15011 gnd.n4046 gnd.n4045 99.6594
R15012 gnd.n4049 gnd.n4048 99.6594
R15013 gnd.n4058 gnd.n4057 99.6594
R15014 gnd.n4061 gnd.n4060 99.6594
R15015 gnd.n4068 gnd.n4067 99.6594
R15016 gnd.n4071 gnd.n4070 99.6594
R15017 gnd.n4078 gnd.n4077 99.6594
R15018 gnd.n4081 gnd.n4080 99.6594
R15019 gnd.n4088 gnd.n4087 99.6594
R15020 gnd.n4091 gnd.n4090 99.6594
R15021 gnd.n4099 gnd.n4098 99.6594
R15022 gnd.n4102 gnd.n4101 99.6594
R15023 gnd.n2295 gnd.n864 99.6594
R15024 gnd.n2293 gnd.n863 99.6594
R15025 gnd.n2289 gnd.n862 99.6594
R15026 gnd.n2285 gnd.n861 99.6594
R15027 gnd.n2281 gnd.n860 99.6594
R15028 gnd.n2277 gnd.n859 99.6594
R15029 gnd.n2273 gnd.n858 99.6594
R15030 gnd.n2205 gnd.n857 99.6594
R15031 gnd.n1534 gnd.n1265 99.6594
R15032 gnd.n1291 gnd.n1272 99.6594
R15033 gnd.n1293 gnd.n1273 99.6594
R15034 gnd.n1301 gnd.n1274 99.6594
R15035 gnd.n1303 gnd.n1275 99.6594
R15036 gnd.n1311 gnd.n1276 99.6594
R15037 gnd.n1313 gnd.n1277 99.6594
R15038 gnd.n1321 gnd.n1278 99.6594
R15039 gnd.n204 gnd.n183 99.6594
R15040 gnd.n210 gnd.n184 99.6594
R15041 gnd.n214 gnd.n185 99.6594
R15042 gnd.n220 gnd.n186 99.6594
R15043 gnd.n224 gnd.n187 99.6594
R15044 gnd.n230 gnd.n188 99.6594
R15045 gnd.n233 gnd.n189 99.6594
R15046 gnd.n240 gnd.n239 99.6594
R15047 gnd.n7332 gnd.n7331 99.6594
R15048 gnd.n5317 gnd.n2735 99.6594
R15049 gnd.n2825 gnd.n2736 99.6594
R15050 gnd.n5216 gnd.n2737 99.6594
R15051 gnd.n5224 gnd.n2738 99.6594
R15052 gnd.n5226 gnd.n2739 99.6594
R15053 gnd.n5236 gnd.n2740 99.6594
R15054 gnd.n5244 gnd.n2741 99.6594
R15055 gnd.n5246 gnd.n2742 99.6594
R15056 gnd.n5256 gnd.n2743 99.6594
R15057 gnd.n2263 gnd.n844 99.6594
R15058 gnd.n2259 gnd.n845 99.6594
R15059 gnd.n2255 gnd.n846 99.6594
R15060 gnd.n2251 gnd.n847 99.6594
R15061 gnd.n2247 gnd.n848 99.6594
R15062 gnd.n2243 gnd.n849 99.6594
R15063 gnd.n2239 gnd.n850 99.6594
R15064 gnd.n2235 gnd.n851 99.6594
R15065 gnd.n2231 gnd.n852 99.6594
R15066 gnd.n2227 gnd.n853 99.6594
R15067 gnd.n2223 gnd.n854 99.6594
R15068 gnd.n2219 gnd.n855 99.6594
R15069 gnd.n2215 gnd.n856 99.6594
R15070 gnd.n1449 gnd.n1448 99.6594
R15071 gnd.n1443 gnd.n1360 99.6594
R15072 gnd.n1440 gnd.n1361 99.6594
R15073 gnd.n1436 gnd.n1362 99.6594
R15074 gnd.n1432 gnd.n1363 99.6594
R15075 gnd.n1428 gnd.n1364 99.6594
R15076 gnd.n1424 gnd.n1365 99.6594
R15077 gnd.n1420 gnd.n1366 99.6594
R15078 gnd.n1416 gnd.n1367 99.6594
R15079 gnd.n1412 gnd.n1368 99.6594
R15080 gnd.n1408 gnd.n1369 99.6594
R15081 gnd.n1404 gnd.n1370 99.6594
R15082 gnd.n1451 gnd.n1359 99.6594
R15083 gnd.n3607 gnd.n3367 99.6594
R15084 gnd.n3404 gnd.n3368 99.6594
R15085 gnd.n3620 gnd.n3369 99.6594
R15086 gnd.n3631 gnd.n3370 99.6594
R15087 gnd.n3392 gnd.n3371 99.6594
R15088 gnd.n3644 gnd.n3372 99.6594
R15089 gnd.n3655 gnd.n3373 99.6594
R15090 gnd.n3376 gnd.n3374 99.6594
R15091 gnd.n3671 gnd.n3670 99.6594
R15092 gnd.n3891 gnd.n3890 99.6594
R15093 gnd.n3888 gnd.n3822 99.6594
R15094 gnd.n3884 gnd.n3883 99.6594
R15095 gnd.n3877 gnd.n3826 99.6594
R15096 gnd.n3876 gnd.n3875 99.6594
R15097 gnd.n3869 gnd.n3832 99.6594
R15098 gnd.n3868 gnd.n3867 99.6594
R15099 gnd.n3861 gnd.n3838 99.6594
R15100 gnd.n3860 gnd.n3859 99.6594
R15101 gnd.n3890 gnd.n3889 99.6594
R15102 gnd.n3885 gnd.n3822 99.6594
R15103 gnd.n3883 gnd.n3882 99.6594
R15104 gnd.n3878 gnd.n3877 99.6594
R15105 gnd.n3875 gnd.n3874 99.6594
R15106 gnd.n3870 gnd.n3869 99.6594
R15107 gnd.n3867 gnd.n3866 99.6594
R15108 gnd.n3862 gnd.n3861 99.6594
R15109 gnd.n3859 gnd.n3858 99.6594
R15110 gnd.n3671 gnd.n3375 99.6594
R15111 gnd.n3656 gnd.n3374 99.6594
R15112 gnd.n3643 gnd.n3373 99.6594
R15113 gnd.n3393 gnd.n3372 99.6594
R15114 gnd.n3632 gnd.n3371 99.6594
R15115 gnd.n3619 gnd.n3370 99.6594
R15116 gnd.n3405 gnd.n3369 99.6594
R15117 gnd.n3608 gnd.n3368 99.6594
R15118 gnd.n3411 gnd.n3367 99.6594
R15119 gnd.n1449 gnd.n1372 99.6594
R15120 gnd.n1441 gnd.n1360 99.6594
R15121 gnd.n1437 gnd.n1361 99.6594
R15122 gnd.n1433 gnd.n1362 99.6594
R15123 gnd.n1429 gnd.n1363 99.6594
R15124 gnd.n1425 gnd.n1364 99.6594
R15125 gnd.n1421 gnd.n1365 99.6594
R15126 gnd.n1417 gnd.n1366 99.6594
R15127 gnd.n1413 gnd.n1367 99.6594
R15128 gnd.n1409 gnd.n1368 99.6594
R15129 gnd.n1405 gnd.n1369 99.6594
R15130 gnd.n1401 gnd.n1370 99.6594
R15131 gnd.n1452 gnd.n1451 99.6594
R15132 gnd.n2218 gnd.n856 99.6594
R15133 gnd.n2222 gnd.n855 99.6594
R15134 gnd.n2226 gnd.n854 99.6594
R15135 gnd.n2230 gnd.n853 99.6594
R15136 gnd.n2234 gnd.n852 99.6594
R15137 gnd.n2238 gnd.n851 99.6594
R15138 gnd.n2242 gnd.n850 99.6594
R15139 gnd.n2246 gnd.n849 99.6594
R15140 gnd.n2250 gnd.n848 99.6594
R15141 gnd.n2254 gnd.n847 99.6594
R15142 gnd.n2258 gnd.n846 99.6594
R15143 gnd.n2262 gnd.n845 99.6594
R15144 gnd.n885 gnd.n844 99.6594
R15145 gnd.n2824 gnd.n2735 99.6594
R15146 gnd.n5215 gnd.n2736 99.6594
R15147 gnd.n5223 gnd.n2737 99.6594
R15148 gnd.n5225 gnd.n2738 99.6594
R15149 gnd.n5235 gnd.n2739 99.6594
R15150 gnd.n5243 gnd.n2740 99.6594
R15151 gnd.n5245 gnd.n2741 99.6594
R15152 gnd.n5255 gnd.n2742 99.6594
R15153 gnd.n5257 gnd.n2743 99.6594
R15154 gnd.n7331 gnd.n181 99.6594
R15155 gnd.n240 gnd.n190 99.6594
R15156 gnd.n231 gnd.n189 99.6594
R15157 gnd.n223 gnd.n188 99.6594
R15158 gnd.n221 gnd.n187 99.6594
R15159 gnd.n213 gnd.n186 99.6594
R15160 gnd.n211 gnd.n185 99.6594
R15161 gnd.n203 gnd.n184 99.6594
R15162 gnd.n201 gnd.n183 99.6594
R15163 gnd.n1535 gnd.n1534 99.6594
R15164 gnd.n1294 gnd.n1272 99.6594
R15165 gnd.n1300 gnd.n1273 99.6594
R15166 gnd.n1304 gnd.n1274 99.6594
R15167 gnd.n1310 gnd.n1275 99.6594
R15168 gnd.n1314 gnd.n1276 99.6594
R15169 gnd.n1320 gnd.n1277 99.6594
R15170 gnd.n1278 gnd.n1262 99.6594
R15171 gnd.n2272 gnd.n857 99.6594
R15172 gnd.n2276 gnd.n858 99.6594
R15173 gnd.n2280 gnd.n859 99.6594
R15174 gnd.n2284 gnd.n860 99.6594
R15175 gnd.n2288 gnd.n861 99.6594
R15176 gnd.n2292 gnd.n862 99.6594
R15177 gnd.n2296 gnd.n863 99.6594
R15178 gnd.n866 gnd.n864 99.6594
R15179 gnd.n3959 gnd.n3958 99.6594
R15180 gnd.n3967 gnd.n3966 99.6594
R15181 gnd.n3968 gnd.n3950 99.6594
R15182 gnd.n3977 gnd.n3976 99.6594
R15183 gnd.n3978 gnd.n3946 99.6594
R15184 gnd.n3987 gnd.n3986 99.6594
R15185 gnd.n3988 gnd.n3942 99.6594
R15186 gnd.n3997 gnd.n3996 99.6594
R15187 gnd.n3998 gnd.n3935 99.6594
R15188 gnd.n4007 gnd.n4006 99.6594
R15189 gnd.n4008 gnd.n3931 99.6594
R15190 gnd.n4017 gnd.n4016 99.6594
R15191 gnd.n4018 gnd.n3927 99.6594
R15192 gnd.n4027 gnd.n4026 99.6594
R15193 gnd.n4028 gnd.n3923 99.6594
R15194 gnd.n4037 gnd.n4036 99.6594
R15195 gnd.n4038 gnd.n3919 99.6594
R15196 gnd.n4047 gnd.n4046 99.6594
R15197 gnd.n4048 gnd.n3915 99.6594
R15198 gnd.n4059 gnd.n4058 99.6594
R15199 gnd.n4060 gnd.n3911 99.6594
R15200 gnd.n4069 gnd.n4068 99.6594
R15201 gnd.n4070 gnd.n3907 99.6594
R15202 gnd.n4079 gnd.n4078 99.6594
R15203 gnd.n4080 gnd.n3903 99.6594
R15204 gnd.n4089 gnd.n4088 99.6594
R15205 gnd.n4090 gnd.n3899 99.6594
R15206 gnd.n4100 gnd.n4099 99.6594
R15207 gnd.n4103 gnd.n4102 99.6594
R15208 gnd.n4427 gnd.n4426 99.6594
R15209 gnd.n4421 gnd.n4413 99.6594
R15210 gnd.n4434 gnd.n4433 99.6594
R15211 gnd.n4412 gnd.n4406 99.6594
R15212 gnd.n4441 gnd.n4440 99.6594
R15213 gnd.n4405 gnd.n4399 99.6594
R15214 gnd.n4448 gnd.n4447 99.6594
R15215 gnd.n4398 gnd.n4392 99.6594
R15216 gnd.n4455 gnd.n4454 99.6594
R15217 gnd.n4458 gnd.n4457 99.6594
R15218 gnd.n4389 gnd.n4381 99.6594
R15219 gnd.n4467 gnd.n4466 99.6594
R15220 gnd.n4380 gnd.n4374 99.6594
R15221 gnd.n4474 gnd.n4473 99.6594
R15222 gnd.n4477 gnd.n4476 99.6594
R15223 gnd.n4324 gnd.n4281 99.6594
R15224 gnd.n4328 gnd.n4282 99.6594
R15225 gnd.n4332 gnd.n4283 99.6594
R15226 gnd.n4336 gnd.n4284 99.6594
R15227 gnd.n4341 gnd.n4285 99.6594
R15228 gnd.n4345 gnd.n4286 99.6594
R15229 gnd.n4349 gnd.n4287 99.6594
R15230 gnd.n4353 gnd.n4288 99.6594
R15231 gnd.n4357 gnd.n4289 99.6594
R15232 gnd.n4361 gnd.n4290 99.6594
R15233 gnd.n4365 gnd.n4291 99.6594
R15234 gnd.n4294 gnd.n4292 99.6594
R15235 gnd.n4371 gnd.n4293 99.6594
R15236 gnd.n5926 gnd.n2747 99.6594
R15237 gnd.n5918 gnd.n2707 99.6594
R15238 gnd.n5914 gnd.n2708 99.6594
R15239 gnd.n5910 gnd.n2709 99.6594
R15240 gnd.n5906 gnd.n2710 99.6594
R15241 gnd.n5902 gnd.n2711 99.6594
R15242 gnd.n5898 gnd.n2712 99.6594
R15243 gnd.n5894 gnd.n2713 99.6594
R15244 gnd.n5889 gnd.n2714 99.6594
R15245 gnd.n5885 gnd.n2715 99.6594
R15246 gnd.n5881 gnd.n2716 99.6594
R15247 gnd.n5877 gnd.n2717 99.6594
R15248 gnd.n5872 gnd.n2719 99.6594
R15249 gnd.n5868 gnd.n2720 99.6594
R15250 gnd.n5864 gnd.n2721 99.6594
R15251 gnd.n5860 gnd.n2722 99.6594
R15252 gnd.n5856 gnd.n2723 99.6594
R15253 gnd.n5852 gnd.n2724 99.6594
R15254 gnd.n5848 gnd.n2725 99.6594
R15255 gnd.n5844 gnd.n2726 99.6594
R15256 gnd.n5840 gnd.n2727 99.6594
R15257 gnd.n5836 gnd.n2728 99.6594
R15258 gnd.n5832 gnd.n2729 99.6594
R15259 gnd.n5828 gnd.n2730 99.6594
R15260 gnd.n5824 gnd.n2731 99.6594
R15261 gnd.n5820 gnd.n2732 99.6594
R15262 gnd.n5816 gnd.n2733 99.6594
R15263 gnd.n2818 gnd.n2734 99.6594
R15264 gnd.n7214 gnd.n7118 99.6594
R15265 gnd.n7218 gnd.n7119 99.6594
R15266 gnd.n7222 gnd.n7120 99.6594
R15267 gnd.n7226 gnd.n7121 99.6594
R15268 gnd.n7230 gnd.n7122 99.6594
R15269 gnd.n7234 gnd.n7123 99.6594
R15270 gnd.n7238 gnd.n7124 99.6594
R15271 gnd.n7242 gnd.n7125 99.6594
R15272 gnd.n7246 gnd.n7126 99.6594
R15273 gnd.n7250 gnd.n7127 99.6594
R15274 gnd.n7256 gnd.n7128 99.6594
R15275 gnd.n7260 gnd.n7129 99.6594
R15276 gnd.n7264 gnd.n7130 99.6594
R15277 gnd.n7268 gnd.n7131 99.6594
R15278 gnd.n7272 gnd.n7132 99.6594
R15279 gnd.n7276 gnd.n7133 99.6594
R15280 gnd.n7280 gnd.n7134 99.6594
R15281 gnd.n7284 gnd.n7135 99.6594
R15282 gnd.n7288 gnd.n7136 99.6594
R15283 gnd.n7292 gnd.n7137 99.6594
R15284 gnd.n7299 gnd.n7138 99.6594
R15285 gnd.n7303 gnd.n7139 99.6594
R15286 gnd.n7307 gnd.n7140 99.6594
R15287 gnd.n7311 gnd.n7141 99.6594
R15288 gnd.n7315 gnd.n7142 99.6594
R15289 gnd.n7319 gnd.n7143 99.6594
R15290 gnd.n7323 gnd.n7144 99.6594
R15291 gnd.n7147 gnd.n7145 99.6594
R15292 gnd.n7329 gnd.n7146 99.6594
R15293 gnd.n3578 gnd.n2550 99.6594
R15294 gnd.n3422 gnd.n2551 99.6594
R15295 gnd.n3586 gnd.n2552 99.6594
R15296 gnd.n3418 gnd.n2553 99.6594
R15297 gnd.n3592 gnd.n2554 99.6594
R15298 gnd.n3602 gnd.n2555 99.6594
R15299 gnd.n3409 gnd.n2556 99.6594
R15300 gnd.n3613 gnd.n2557 99.6594
R15301 gnd.n3626 gnd.n2558 99.6594
R15302 gnd.n3397 gnd.n2559 99.6594
R15303 gnd.n3637 gnd.n2560 99.6594
R15304 gnd.n3650 gnd.n2561 99.6594
R15305 gnd.n3385 gnd.n2562 99.6594
R15306 gnd.n3662 gnd.n2563 99.6594
R15307 gnd.n3421 gnd.n2550 99.6594
R15308 gnd.n3585 gnd.n2551 99.6594
R15309 gnd.n3417 gnd.n2552 99.6594
R15310 gnd.n3593 gnd.n2553 99.6594
R15311 gnd.n3601 gnd.n2554 99.6594
R15312 gnd.n3408 gnd.n2555 99.6594
R15313 gnd.n3614 gnd.n2556 99.6594
R15314 gnd.n3625 gnd.n2557 99.6594
R15315 gnd.n3396 gnd.n2558 99.6594
R15316 gnd.n3638 gnd.n2559 99.6594
R15317 gnd.n3649 gnd.n2560 99.6594
R15318 gnd.n3384 gnd.n2561 99.6594
R15319 gnd.n3663 gnd.n2562 99.6594
R15320 gnd.n2563 gnd.n2547 99.6594
R15321 gnd.n5188 gnd.n2684 99.6594
R15322 gnd.n2835 gnd.n2685 99.6594
R15323 gnd.n5196 gnd.n2686 99.6594
R15324 gnd.n2831 gnd.n2687 99.6594
R15325 gnd.n5204 gnd.n2688 99.6594
R15326 gnd.n5210 gnd.n2689 99.6594
R15327 gnd.n5212 gnd.n2690 99.6594
R15328 gnd.n5220 gnd.n2691 99.6594
R15329 gnd.n5230 gnd.n2692 99.6594
R15330 gnd.n5232 gnd.n2693 99.6594
R15331 gnd.n5240 gnd.n2694 99.6594
R15332 gnd.n5250 gnd.n2695 99.6594
R15333 gnd.n5252 gnd.n2696 99.6594
R15334 gnd.n5266 gnd.n2697 99.6594
R15335 gnd.n5251 gnd.n2695 99.6594
R15336 gnd.n5249 gnd.n2694 99.6594
R15337 gnd.n5239 gnd.n2693 99.6594
R15338 gnd.n5231 gnd.n2692 99.6594
R15339 gnd.n5229 gnd.n2691 99.6594
R15340 gnd.n5219 gnd.n2690 99.6594
R15341 gnd.n5211 gnd.n2689 99.6594
R15342 gnd.n5209 gnd.n2688 99.6594
R15343 gnd.n5203 gnd.n2687 99.6594
R15344 gnd.n2830 gnd.n2686 99.6594
R15345 gnd.n5195 gnd.n2685 99.6594
R15346 gnd.n2834 gnd.n2684 99.6594
R15347 gnd.n2697 gnd.n2681 99.6594
R15348 gnd.n5265 gnd.n2696 99.6594
R15349 gnd.n3381 gnd.t244 98.63
R15350 gnd.n5258 gnd.t271 98.63
R15351 gnd.n3378 gnd.t282 98.63
R15352 gnd.n2767 gnd.t268 98.63
R15353 gnd.n2790 gnd.t256 98.63
R15354 gnd.n2812 gnd.t200 98.63
R15355 gnd.n7209 gnd.t202 98.63
R15356 gnd.n7188 gnd.t195 98.63
R15357 gnd.n7295 gnd.t261 98.63
R15358 gnd.n178 gnd.t276 98.63
R15359 gnd.n3939 gnd.t234 98.63
R15360 gnd.n4050 gnd.t213 98.63
R15361 gnd.n3895 gnd.t237 98.63
R15362 gnd.n3855 gnd.t192 98.63
R15363 gnd.n4315 gnd.t273 98.63
R15364 gnd.n4418 gnd.t220 98.63
R15365 gnd.n4385 gnd.t239 98.63
R15366 gnd.n5262 gnd.t224 98.63
R15367 gnd.n3286 gnd.t253 96.6984
R15368 gnd.n2938 gnd.t209 96.6984
R15369 gnd.n3283 gnd.t174 96.6906
R15370 gnd.n2932 gnd.t258 96.6906
R15371 gnd.n3235 gnd.n3234 81.8399
R15372 gnd.n1323 gnd.t286 74.8376
R15373 gnd.n882 gnd.t182 74.8376
R15374 gnd.n3287 gnd.t252 72.8438
R15375 gnd.n2939 gnd.t210 72.8438
R15376 gnd.n3236 gnd.n3229 72.8411
R15377 gnd.n3242 gnd.n3227 72.8411
R15378 gnd.n2907 gnd.n2906 72.8411
R15379 gnd.n3382 gnd.t243 72.836
R15380 gnd.n3284 gnd.t173 72.836
R15381 gnd.n2933 gnd.t259 72.836
R15382 gnd.n5259 gnd.t270 72.836
R15383 gnd.n3379 gnd.t283 72.836
R15384 gnd.n2768 gnd.t267 72.836
R15385 gnd.n2791 gnd.t255 72.836
R15386 gnd.n2813 gnd.t199 72.836
R15387 gnd.n7210 gnd.t203 72.836
R15388 gnd.n7189 gnd.t196 72.836
R15389 gnd.n7296 gnd.t262 72.836
R15390 gnd.n179 gnd.t277 72.836
R15391 gnd.n3940 gnd.t233 72.836
R15392 gnd.n4051 gnd.t212 72.836
R15393 gnd.n3896 gnd.t236 72.836
R15394 gnd.n3856 gnd.t191 72.836
R15395 gnd.n4316 gnd.t274 72.836
R15396 gnd.n4419 gnd.t221 72.836
R15397 gnd.n4386 gnd.t240 72.836
R15398 gnd.n5263 gnd.t225 72.836
R15399 gnd.n5121 gnd.n2912 71.676
R15400 gnd.n5119 gnd.n5118 71.676
R15401 gnd.n5114 gnd.n2915 71.676
R15402 gnd.n5112 gnd.n5111 71.676
R15403 gnd.n5107 gnd.n2918 71.676
R15404 gnd.n5105 gnd.n5104 71.676
R15405 gnd.n5100 gnd.n2921 71.676
R15406 gnd.n5098 gnd.n5097 71.676
R15407 gnd.n5093 gnd.n2924 71.676
R15408 gnd.n5091 gnd.n5090 71.676
R15409 gnd.n5086 gnd.n2927 71.676
R15410 gnd.n5084 gnd.n5083 71.676
R15411 gnd.n5079 gnd.n2930 71.676
R15412 gnd.n5077 gnd.n5076 71.676
R15413 gnd.n5071 gnd.n2935 71.676
R15414 gnd.n5069 gnd.n5068 71.676
R15415 gnd.n5064 gnd.n5063 71.676
R15416 gnd.n5061 gnd.n5060 71.676
R15417 gnd.n5055 gnd.n2941 71.676
R15418 gnd.n5053 gnd.n5052 71.676
R15419 gnd.n5048 gnd.n2944 71.676
R15420 gnd.n5046 gnd.n5045 71.676
R15421 gnd.n5041 gnd.n2947 71.676
R15422 gnd.n5039 gnd.n5038 71.676
R15423 gnd.n5034 gnd.n2950 71.676
R15424 gnd.n5032 gnd.n5031 71.676
R15425 gnd.n5027 gnd.n2953 71.676
R15426 gnd.n5025 gnd.n5024 71.676
R15427 gnd.n5020 gnd.n2956 71.676
R15428 gnd.n5018 gnd.n5017 71.676
R15429 gnd.n5013 gnd.n2959 71.676
R15430 gnd.n5011 gnd.n5010 71.676
R15431 gnd.n5006 gnd.n5005 71.676
R15432 gnd.n4548 gnd.n4547 71.676
R15433 gnd.n3282 gnd.n3249 71.676
R15434 gnd.n4540 gnd.n3250 71.676
R15435 gnd.n4536 gnd.n3251 71.676
R15436 gnd.n4532 gnd.n3252 71.676
R15437 gnd.n4528 gnd.n3253 71.676
R15438 gnd.n4524 gnd.n3254 71.676
R15439 gnd.n4520 gnd.n3255 71.676
R15440 gnd.n4516 gnd.n3256 71.676
R15441 gnd.n4512 gnd.n3257 71.676
R15442 gnd.n4508 gnd.n3258 71.676
R15443 gnd.n4504 gnd.n3259 71.676
R15444 gnd.n4500 gnd.n3260 71.676
R15445 gnd.n4496 gnd.n3261 71.676
R15446 gnd.n4492 gnd.n3262 71.676
R15447 gnd.n4488 gnd.n3263 71.676
R15448 gnd.n4484 gnd.n3265 71.676
R15449 gnd.n3355 gnd.n3266 71.676
R15450 gnd.n3350 gnd.n3267 71.676
R15451 gnd.n3346 gnd.n3268 71.676
R15452 gnd.n3342 gnd.n3269 71.676
R15453 gnd.n3338 gnd.n3270 71.676
R15454 gnd.n3334 gnd.n3271 71.676
R15455 gnd.n3330 gnd.n3272 71.676
R15456 gnd.n3326 gnd.n3273 71.676
R15457 gnd.n3322 gnd.n3274 71.676
R15458 gnd.n3318 gnd.n3275 71.676
R15459 gnd.n3314 gnd.n3276 71.676
R15460 gnd.n3310 gnd.n3277 71.676
R15461 gnd.n3306 gnd.n3278 71.676
R15462 gnd.n3302 gnd.n3279 71.676
R15463 gnd.n3298 gnd.n3280 71.676
R15464 gnd.n4547 gnd.n3247 71.676
R15465 gnd.n4541 gnd.n3249 71.676
R15466 gnd.n4537 gnd.n3250 71.676
R15467 gnd.n4533 gnd.n3251 71.676
R15468 gnd.n4529 gnd.n3252 71.676
R15469 gnd.n4525 gnd.n3253 71.676
R15470 gnd.n4521 gnd.n3254 71.676
R15471 gnd.n4517 gnd.n3255 71.676
R15472 gnd.n4513 gnd.n3256 71.676
R15473 gnd.n4509 gnd.n3257 71.676
R15474 gnd.n4505 gnd.n3258 71.676
R15475 gnd.n4501 gnd.n3259 71.676
R15476 gnd.n4497 gnd.n3260 71.676
R15477 gnd.n4493 gnd.n3261 71.676
R15478 gnd.n4489 gnd.n3262 71.676
R15479 gnd.n4485 gnd.n3264 71.676
R15480 gnd.n3356 gnd.n3265 71.676
R15481 gnd.n3351 gnd.n3266 71.676
R15482 gnd.n3347 gnd.n3267 71.676
R15483 gnd.n3343 gnd.n3268 71.676
R15484 gnd.n3339 gnd.n3269 71.676
R15485 gnd.n3335 gnd.n3270 71.676
R15486 gnd.n3331 gnd.n3271 71.676
R15487 gnd.n3327 gnd.n3272 71.676
R15488 gnd.n3323 gnd.n3273 71.676
R15489 gnd.n3319 gnd.n3274 71.676
R15490 gnd.n3315 gnd.n3275 71.676
R15491 gnd.n3311 gnd.n3276 71.676
R15492 gnd.n3307 gnd.n3277 71.676
R15493 gnd.n3303 gnd.n3278 71.676
R15494 gnd.n3299 gnd.n3279 71.676
R15495 gnd.n3295 gnd.n3280 71.676
R15496 gnd.n5005 gnd.n2960 71.676
R15497 gnd.n5012 gnd.n5011 71.676
R15498 gnd.n2959 gnd.n2957 71.676
R15499 gnd.n5019 gnd.n5018 71.676
R15500 gnd.n2956 gnd.n2954 71.676
R15501 gnd.n5026 gnd.n5025 71.676
R15502 gnd.n2953 gnd.n2951 71.676
R15503 gnd.n5033 gnd.n5032 71.676
R15504 gnd.n2950 gnd.n2948 71.676
R15505 gnd.n5040 gnd.n5039 71.676
R15506 gnd.n2947 gnd.n2945 71.676
R15507 gnd.n5047 gnd.n5046 71.676
R15508 gnd.n2944 gnd.n2942 71.676
R15509 gnd.n5054 gnd.n5053 71.676
R15510 gnd.n2941 gnd.n2937 71.676
R15511 gnd.n5062 gnd.n5061 71.676
R15512 gnd.n5066 gnd.n5065 71.676
R15513 gnd.n5070 gnd.n5069 71.676
R15514 gnd.n2935 gnd.n2931 71.676
R15515 gnd.n5078 gnd.n5077 71.676
R15516 gnd.n2930 gnd.n2928 71.676
R15517 gnd.n5085 gnd.n5084 71.676
R15518 gnd.n2927 gnd.n2925 71.676
R15519 gnd.n5092 gnd.n5091 71.676
R15520 gnd.n2924 gnd.n2922 71.676
R15521 gnd.n5099 gnd.n5098 71.676
R15522 gnd.n2921 gnd.n2919 71.676
R15523 gnd.n5106 gnd.n5105 71.676
R15524 gnd.n2918 gnd.n2916 71.676
R15525 gnd.n5113 gnd.n5112 71.676
R15526 gnd.n2915 gnd.n2913 71.676
R15527 gnd.n5120 gnd.n5119 71.676
R15528 gnd.n2912 gnd.n2890 71.676
R15529 gnd.n8 gnd.t132 69.1507
R15530 gnd.n14 gnd.t310 68.4792
R15531 gnd.n13 gnd.t170 68.4792
R15532 gnd.n12 gnd.t168 68.4792
R15533 gnd.n11 gnd.t163 68.4792
R15534 gnd.n10 gnd.t1 68.4792
R15535 gnd.n9 gnd.t9 68.4792
R15536 gnd.n8 gnd.t140 68.4792
R15537 gnd.n1450 gnd.n1354 64.369
R15538 gnd.n3353 gnd.n3287 59.5399
R15539 gnd.n5057 gnd.n2939 59.5399
R15540 gnd.n3285 gnd.n3284 59.5399
R15541 gnd.n5073 gnd.n2933 59.5399
R15542 gnd.n4550 gnd.n3245 59.1804
R15543 gnd.n2304 gnd.n842 57.3586
R15544 gnd.n1109 gnd.t68 56.407
R15545 gnd.n1074 gnd.t115 56.407
R15546 gnd.n1085 gnd.t27 56.407
R15547 gnd.n1097 gnd.t108 56.407
R15548 gnd.n52 gnd.t43 56.407
R15549 gnd.n17 gnd.t34 56.407
R15550 gnd.n28 gnd.t124 56.407
R15551 gnd.n40 gnd.t83 56.407
R15552 gnd.n1118 gnd.t94 55.8337
R15553 gnd.n1083 gnd.t23 55.8337
R15554 gnd.n1094 gnd.t126 55.8337
R15555 gnd.n1106 gnd.t28 55.8337
R15556 gnd.n61 gnd.t66 55.8337
R15557 gnd.n26 gnd.t59 55.8337
R15558 gnd.n37 gnd.t107 55.8337
R15559 gnd.n49 gnd.t104 55.8337
R15560 gnd.n6232 gnd.n6231 55.128
R15561 gnd.n7101 gnd.n250 55.128
R15562 gnd.n3233 gnd.n3232 54.358
R15563 gnd.n2904 gnd.n2903 54.358
R15564 gnd.n1109 gnd.n1108 53.0052
R15565 gnd.n1111 gnd.n1110 53.0052
R15566 gnd.n1113 gnd.n1112 53.0052
R15567 gnd.n1115 gnd.n1114 53.0052
R15568 gnd.n1117 gnd.n1116 53.0052
R15569 gnd.n1074 gnd.n1073 53.0052
R15570 gnd.n1076 gnd.n1075 53.0052
R15571 gnd.n1078 gnd.n1077 53.0052
R15572 gnd.n1080 gnd.n1079 53.0052
R15573 gnd.n1082 gnd.n1081 53.0052
R15574 gnd.n1085 gnd.n1084 53.0052
R15575 gnd.n1087 gnd.n1086 53.0052
R15576 gnd.n1089 gnd.n1088 53.0052
R15577 gnd.n1091 gnd.n1090 53.0052
R15578 gnd.n1093 gnd.n1092 53.0052
R15579 gnd.n1097 gnd.n1096 53.0052
R15580 gnd.n1099 gnd.n1098 53.0052
R15581 gnd.n1101 gnd.n1100 53.0052
R15582 gnd.n1103 gnd.n1102 53.0052
R15583 gnd.n1105 gnd.n1104 53.0052
R15584 gnd.n60 gnd.n59 53.0052
R15585 gnd.n58 gnd.n57 53.0052
R15586 gnd.n56 gnd.n55 53.0052
R15587 gnd.n54 gnd.n53 53.0052
R15588 gnd.n52 gnd.n51 53.0052
R15589 gnd.n25 gnd.n24 53.0052
R15590 gnd.n23 gnd.n22 53.0052
R15591 gnd.n21 gnd.n20 53.0052
R15592 gnd.n19 gnd.n18 53.0052
R15593 gnd.n17 gnd.n16 53.0052
R15594 gnd.n36 gnd.n35 53.0052
R15595 gnd.n34 gnd.n33 53.0052
R15596 gnd.n32 gnd.n31 53.0052
R15597 gnd.n30 gnd.n29 53.0052
R15598 gnd.n28 gnd.n27 53.0052
R15599 gnd.n48 gnd.n47 53.0052
R15600 gnd.n46 gnd.n45 53.0052
R15601 gnd.n44 gnd.n43 53.0052
R15602 gnd.n42 gnd.n41 53.0052
R15603 gnd.n40 gnd.n39 53.0052
R15604 gnd.n2895 gnd.n2894 52.4801
R15605 gnd.n2156 gnd.t144 52.3082
R15606 gnd.n2124 gnd.t142 52.3082
R15607 gnd.n2092 gnd.t316 52.3082
R15608 gnd.n2061 gnd.t319 52.3082
R15609 gnd.n2029 gnd.t159 52.3082
R15610 gnd.n1997 gnd.t151 52.3082
R15611 gnd.n1965 gnd.t154 52.3082
R15612 gnd.n1934 gnd.t308 52.3082
R15613 gnd.n1986 gnd.n1954 51.4173
R15614 gnd.n2050 gnd.n2049 50.455
R15615 gnd.n2018 gnd.n2017 50.455
R15616 gnd.n1986 gnd.n1985 50.455
R15617 gnd.n1397 gnd.n1396 45.1884
R15618 gnd.n908 gnd.n907 45.1884
R15619 gnd.n5124 gnd.n2910 44.3322
R15620 gnd.n3236 gnd.n3235 44.3189
R15621 gnd.n6400 gnd.n6399 43.8864
R15622 gnd.n6399 gnd.n6398 43.8864
R15623 gnd.n6398 gnd.n676 43.8864
R15624 gnd.n6392 gnd.n676 43.8864
R15625 gnd.n6392 gnd.n6391 43.8864
R15626 gnd.n6391 gnd.n6390 43.8864
R15627 gnd.n6390 gnd.n683 43.8864
R15628 gnd.n6384 gnd.n683 43.8864
R15629 gnd.n6384 gnd.n6383 43.8864
R15630 gnd.n6383 gnd.n6382 43.8864
R15631 gnd.n6382 gnd.n691 43.8864
R15632 gnd.n6376 gnd.n691 43.8864
R15633 gnd.n6376 gnd.n6375 43.8864
R15634 gnd.n6375 gnd.n6374 43.8864
R15635 gnd.n6374 gnd.n699 43.8864
R15636 gnd.n6368 gnd.n699 43.8864
R15637 gnd.n6368 gnd.n6367 43.8864
R15638 gnd.n6367 gnd.n6366 43.8864
R15639 gnd.n6366 gnd.n707 43.8864
R15640 gnd.n6360 gnd.n707 43.8864
R15641 gnd.n6360 gnd.n6359 43.8864
R15642 gnd.n6359 gnd.n6358 43.8864
R15643 gnd.n6358 gnd.n715 43.8864
R15644 gnd.n6352 gnd.n715 43.8864
R15645 gnd.n6352 gnd.n6351 43.8864
R15646 gnd.n6351 gnd.n6350 43.8864
R15647 gnd.n6350 gnd.n723 43.8864
R15648 gnd.n6344 gnd.n723 43.8864
R15649 gnd.n6344 gnd.n6343 43.8864
R15650 gnd.n6343 gnd.n6342 43.8864
R15651 gnd.n6342 gnd.n731 43.8864
R15652 gnd.n6336 gnd.n731 43.8864
R15653 gnd.n6336 gnd.n6335 43.8864
R15654 gnd.n6335 gnd.n6334 43.8864
R15655 gnd.n6334 gnd.n739 43.8864
R15656 gnd.n6328 gnd.n739 43.8864
R15657 gnd.n6328 gnd.n6327 43.8864
R15658 gnd.n6327 gnd.n6326 43.8864
R15659 gnd.n6326 gnd.n747 43.8864
R15660 gnd.n6320 gnd.n747 43.8864
R15661 gnd.n6320 gnd.n6319 43.8864
R15662 gnd.n6319 gnd.n6318 43.8864
R15663 gnd.n6318 gnd.n755 43.8864
R15664 gnd.n6312 gnd.n755 43.8864
R15665 gnd.n6312 gnd.n6311 43.8864
R15666 gnd.n6311 gnd.n6310 43.8864
R15667 gnd.n6310 gnd.n763 43.8864
R15668 gnd.n6304 gnd.n763 43.8864
R15669 gnd.n6304 gnd.n6303 43.8864
R15670 gnd.n6303 gnd.n6302 43.8864
R15671 gnd.n6302 gnd.n771 43.8864
R15672 gnd.n6296 gnd.n771 43.8864
R15673 gnd.n6296 gnd.n6295 43.8864
R15674 gnd.n6295 gnd.n6294 43.8864
R15675 gnd.n6294 gnd.n779 43.8864
R15676 gnd.n6288 gnd.n779 43.8864
R15677 gnd.n6288 gnd.n6287 43.8864
R15678 gnd.n6287 gnd.n6286 43.8864
R15679 gnd.n6286 gnd.n787 43.8864
R15680 gnd.n6280 gnd.n787 43.8864
R15681 gnd.n6280 gnd.n6279 43.8864
R15682 gnd.n6279 gnd.n6278 43.8864
R15683 gnd.n6278 gnd.n795 43.8864
R15684 gnd.n6272 gnd.n795 43.8864
R15685 gnd.n6272 gnd.n6271 43.8864
R15686 gnd.n6271 gnd.n6270 43.8864
R15687 gnd.n6270 gnd.n803 43.8864
R15688 gnd.n6264 gnd.n803 43.8864
R15689 gnd.n6264 gnd.n6263 43.8864
R15690 gnd.n6263 gnd.n6262 43.8864
R15691 gnd.n6262 gnd.n811 43.8864
R15692 gnd.n6256 gnd.n811 43.8864
R15693 gnd.n6256 gnd.n6255 43.8864
R15694 gnd.n6255 gnd.n6254 43.8864
R15695 gnd.n6254 gnd.n819 43.8864
R15696 gnd.n6248 gnd.n819 43.8864
R15697 gnd.n6248 gnd.n6247 43.8864
R15698 gnd.n6247 gnd.n6246 43.8864
R15699 gnd.n6246 gnd.n827 43.8864
R15700 gnd.n6240 gnd.n827 43.8864
R15701 gnd.n6240 gnd.n6239 43.8864
R15702 gnd.n6239 gnd.n6238 43.8864
R15703 gnd.n6238 gnd.n835 43.8864
R15704 gnd.n3661 gnd.n3382 42.2793
R15705 gnd.n5260 gnd.n5259 42.2793
R15706 gnd.n1398 gnd.n1397 42.2793
R15707 gnd.n909 gnd.n908 42.2793
R15708 gnd.n1324 gnd.n1323 42.2793
R15709 gnd.n2271 gnd.n882 42.2793
R15710 gnd.n3668 gnd.n3379 42.2793
R15711 gnd.n5891 gnd.n2768 42.2793
R15712 gnd.n5854 gnd.n2791 42.2793
R15713 gnd.n5814 gnd.n2813 42.2793
R15714 gnd.n7213 gnd.n7210 42.2793
R15715 gnd.n7255 gnd.n7189 42.2793
R15716 gnd.n7297 gnd.n7296 42.2793
R15717 gnd.n180 gnd.n179 42.2793
R15718 gnd.n3941 gnd.n3940 42.2793
R15719 gnd.n4052 gnd.n4051 42.2793
R15720 gnd.n3897 gnd.n3896 42.2793
R15721 gnd.n3857 gnd.n3856 42.2793
R15722 gnd.n4339 gnd.n4316 42.2793
R15723 gnd.n4420 gnd.n4419 42.2793
R15724 gnd.n4463 gnd.n4386 42.2793
R15725 gnd.n5264 gnd.n5263 42.2793
R15726 gnd.n3234 gnd.n3233 41.6274
R15727 gnd.n2905 gnd.n2904 41.6274
R15728 gnd.n3243 gnd.n3242 40.8975
R15729 gnd.n2908 gnd.n2907 40.8975
R15730 gnd.n3242 gnd.n3241 35.055
R15731 gnd.n3237 gnd.n3236 35.055
R15732 gnd.n2897 gnd.n2896 35.055
R15733 gnd.n2907 gnd.n2893 35.055
R15734 gnd.n5007 gnd.n5004 33.2493
R15735 gnd.n3296 gnd.n3293 33.2493
R15736 gnd.n1460 gnd.n1354 31.8661
R15737 gnd.n1460 gnd.n1459 31.8661
R15738 gnd.n1468 gnd.n1343 31.8661
R15739 gnd.n1476 gnd.n1343 31.8661
R15740 gnd.n1476 gnd.n1337 31.8661
R15741 gnd.n1484 gnd.n1337 31.8661
R15742 gnd.n1484 gnd.n1330 31.8661
R15743 gnd.n1522 gnd.n1330 31.8661
R15744 gnd.n1532 gnd.n1263 31.8661
R15745 gnd.n6231 gnd.n6230 31.8661
R15746 gnd.n6230 gnd.n2305 31.8661
R15747 gnd.n6224 gnd.n2305 31.8661
R15748 gnd.n6224 gnd.n6223 31.8661
R15749 gnd.n6223 gnd.n6222 31.8661
R15750 gnd.n6216 gnd.n2322 31.8661
R15751 gnd.n3366 gnd.n2535 31.8661
R15752 gnd.n4279 gnd.n2549 31.8661
R15753 gnd.n6069 gnd.n2549 31.8661
R15754 gnd.n6069 gnd.n2564 31.8661
R15755 gnd.n6063 gnd.n2564 31.8661
R15756 gnd.n6063 gnd.n6062 31.8661
R15757 gnd.n3458 gnd.n3449 31.8661
R15758 gnd.n3459 gnd.n3458 31.8661
R15759 gnd.n3462 gnd.n3459 31.8661
R15760 gnd.n3462 gnd.n3461 31.8661
R15761 gnd.n3471 gnd.n3470 31.8661
R15762 gnd.n3474 gnd.n3471 31.8661
R15763 gnd.n3474 gnd.n3473 31.8661
R15764 gnd.n3484 gnd.n3248 31.8661
R15765 gnd.n5144 gnd.n2864 31.8661
R15766 gnd.n5152 gnd.n2864 31.8661
R15767 gnd.n5152 gnd.n2865 31.8661
R15768 gnd.n5160 gnd.n2852 31.8661
R15769 gnd.n5168 gnd.n2852 31.8661
R15770 gnd.n5168 gnd.n2845 31.8661
R15771 gnd.n5177 gnd.n2845 31.8661
R15772 gnd.n5186 gnd.n2839 31.8661
R15773 gnd.n5186 gnd.n2683 31.8661
R15774 gnd.n5934 gnd.n2683 31.8661
R15775 gnd.n5934 gnd.n2698 31.8661
R15776 gnd.n5928 gnd.n2698 31.8661
R15777 gnd.n2820 gnd.n2745 31.8661
R15778 gnd.n182 gnd.n170 31.8661
R15779 gnd.n7117 gnd.n241 31.8661
R15780 gnd.n7111 gnd.n241 31.8661
R15781 gnd.n7111 gnd.n7110 31.8661
R15782 gnd.n7110 gnd.n7109 31.8661
R15783 gnd.n7109 gnd.n250 31.8661
R15784 gnd.n3473 gnd.t131 30.9101
R15785 gnd.n5144 gnd.t146 30.9101
R15786 gnd.t264 gnd.n2878 30.5915
R15787 gnd.n4546 gnd.n3281 28.3609
R15788 gnd.n2888 gnd.n2877 28.3609
R15789 gnd.n4372 gnd.n4279 27.4049
R15790 gnd.n5928 gnd.n5927 27.4049
R15791 gnd.n6215 gnd.n2325 26.7676
R15792 gnd.n6209 gnd.n2337 26.7676
R15793 gnd.n4114 gnd.n2346 26.7676
R15794 gnd.n6203 gnd.n2349 26.7676
R15795 gnd.n4122 gnd.n2357 26.7676
R15796 gnd.n4128 gnd.n2366 26.7676
R15797 gnd.n6191 gnd.n2369 26.7676
R15798 gnd.n6185 gnd.n2380 26.7676
R15799 gnd.n6179 gnd.n2390 26.7676
R15800 gnd.n4150 gnd.n2398 26.7676
R15801 gnd.n4156 gnd.n2407 26.7676
R15802 gnd.n6167 gnd.n2410 26.7676
R15803 gnd.n6160 gnd.n2419 26.7676
R15804 gnd.n6154 gnd.n2429 26.7676
R15805 gnd.n4178 gnd.n2434 26.7676
R15806 gnd.n4184 gnd.n2443 26.7676
R15807 gnd.n6141 gnd.n2446 26.7676
R15808 gnd.n4192 gnd.n2451 26.7676
R15809 gnd.n6134 gnd.n2454 26.7676
R15810 gnd.n6128 gnd.n2464 26.7676
R15811 gnd.n4206 gnd.n2472 26.7676
R15812 gnd.n4245 gnd.n2481 26.7676
R15813 gnd.n6116 gnd.n2484 26.7676
R15814 gnd.n4213 gnd.n2492 26.7676
R15815 gnd.n6110 gnd.n2495 26.7676
R15816 gnd.n6104 gnd.n2505 26.7676
R15817 gnd.n4222 gnd.n2513 26.7676
R15818 gnd.n6098 gnd.n2516 26.7676
R15819 gnd.n4228 gnd.n2523 26.7676
R15820 gnd.n6079 gnd.n2532 26.7676
R15821 gnd.n6086 gnd.n2535 26.7676
R15822 gnd.n5807 gnd.n2820 26.7676
R15823 gnd.n5804 gnd.n2822 26.7676
R15824 gnd.n5798 gnd.n5330 26.7676
R15825 gnd.n5503 gnd.n5333 26.7676
R15826 gnd.n5792 gnd.n5341 26.7676
R15827 gnd.n5539 gnd.n5344 26.7676
R15828 gnd.n5510 gnd.n5354 26.7676
R15829 gnd.n5780 gnd.n5361 26.7676
R15830 gnd.n5516 gnd.n5515 26.7676
R15831 gnd.n5774 gnd.n5371 26.7676
R15832 gnd.n5768 gnd.n5381 26.7676
R15833 gnd.n5564 gnd.n5384 26.7676
R15834 gnd.n5580 gnd.n5393 26.7676
R15835 gnd.n5756 gnd.n5400 26.7676
R15836 gnd.n5751 gnd.n5404 26.7676
R15837 gnd.n5750 gnd.n5407 26.7676
R15838 gnd.n5743 gnd.n5742 26.7676
R15839 gnd.n5599 gnd.n5417 26.7676
R15840 gnd.n5729 gnd.n70 26.7676
R15841 gnd.n7394 gnd.n85 26.7676
R15842 gnd.n5719 gnd.n88 26.7676
R15843 gnd.n5713 gnd.n99 26.7676
R15844 gnd.n7382 gnd.n106 26.7676
R15845 gnd.n7376 gnd.n116 26.7676
R15846 gnd.n7370 gnd.n127 26.7676
R15847 gnd.n5695 gnd.n130 26.7676
R15848 gnd.n5642 gnd.n139 26.7676
R15849 gnd.n7358 gnd.n147 26.7676
R15850 gnd.n5636 gnd.n150 26.7676
R15851 gnd.n7352 gnd.n157 26.7676
R15852 gnd.n7346 gnd.n167 26.7676
R15853 gnd.t39 gnd.n2416 26.4489
R15854 gnd.n5728 gnd.t13 26.4489
R15855 gnd.n1004 gnd.n835 26.332
R15856 gnd.n2322 gnd.n2314 26.1303
R15857 gnd.n7330 gnd.n182 26.1303
R15858 gnd.t60 gnd.n2377 25.8116
R15859 gnd.t17 gnd.n119 25.8116
R15860 gnd.n3382 gnd.n3381 25.7944
R15861 gnd.n5259 gnd.n5258 25.7944
R15862 gnd.n1323 gnd.n1322 25.7944
R15863 gnd.n882 gnd.n881 25.7944
R15864 gnd.n3379 gnd.n3378 25.7944
R15865 gnd.n2768 gnd.n2767 25.7944
R15866 gnd.n2791 gnd.n2790 25.7944
R15867 gnd.n2813 gnd.n2812 25.7944
R15868 gnd.n7210 gnd.n7209 25.7944
R15869 gnd.n7189 gnd.n7188 25.7944
R15870 gnd.n7296 gnd.n7295 25.7944
R15871 gnd.n179 gnd.n178 25.7944
R15872 gnd.n3940 gnd.n3939 25.7944
R15873 gnd.n4051 gnd.n4050 25.7944
R15874 gnd.n3896 gnd.n3895 25.7944
R15875 gnd.n3856 gnd.n3855 25.7944
R15876 gnd.n4316 gnd.n4315 25.7944
R15877 gnd.n4419 gnd.n4418 25.7944
R15878 gnd.n4386 gnd.n4385 25.7944
R15879 gnd.n5263 gnd.n5262 25.7944
R15880 gnd.n1544 gnd.n1264 24.8557
R15881 gnd.n1554 gnd.n1247 24.8557
R15882 gnd.n1250 gnd.n1238 24.8557
R15883 gnd.n1575 gnd.n1239 24.8557
R15884 gnd.n1585 gnd.n1219 24.8557
R15885 gnd.n1595 gnd.n1594 24.8557
R15886 gnd.n1205 gnd.n1203 24.8557
R15887 gnd.n1626 gnd.n1625 24.8557
R15888 gnd.n1641 gnd.n1188 24.8557
R15889 gnd.n1695 gnd.n1127 24.8557
R15890 gnd.n1651 gnd.n1128 24.8557
R15891 gnd.n1688 gnd.n1139 24.8557
R15892 gnd.n1177 gnd.n1176 24.8557
R15893 gnd.n1682 gnd.n1681 24.8557
R15894 gnd.n1163 gnd.n1150 24.8557
R15895 gnd.n1721 gnd.n1720 24.8557
R15896 gnd.n1731 gnd.n1059 24.8557
R15897 gnd.n1743 gnd.n1051 24.8557
R15898 gnd.n1742 gnd.n1039 24.8557
R15899 gnd.n1761 gnd.n1760 24.8557
R15900 gnd.n1771 gnd.n1032 24.8557
R15901 gnd.n1782 gnd.n1020 24.8557
R15902 gnd.n1808 gnd.n1807 24.8557
R15903 gnd.n1818 gnd.n1006 24.8557
R15904 gnd.n1830 gnd.n997 24.8557
R15905 gnd.n1848 gnd.n1847 24.8557
R15906 gnd.n988 gnd.n977 24.8557
R15907 gnd.n1869 gnd.n965 24.8557
R15908 gnd.n1897 gnd.n1896 24.8557
R15909 gnd.n1908 gnd.n950 24.8557
R15910 gnd.n1919 gnd.n943 24.8557
R15911 gnd.n1918 gnd.n931 24.8557
R15912 gnd.n2191 gnd.n2190 24.8557
R15913 gnd.n2213 gnd.n916 24.8557
R15914 gnd.n3287 gnd.n3286 23.855
R15915 gnd.n2939 gnd.n2938 23.855
R15916 gnd.n3284 gnd.n3283 23.855
R15917 gnd.n2933 gnd.n2932 23.855
R15918 gnd.n1565 gnd.t307 23.2624
R15919 gnd.n1266 gnd.t285 22.6251
R15920 gnd.n4142 gnd.t46 21.9878
R15921 gnd.n5707 gnd.t80 21.9878
R15922 gnd.n4587 gnd.n3198 21.6691
R15923 gnd.n4608 gnd.n3189 21.6691
R15924 gnd.n4615 gnd.n4614 21.6691
R15925 gnd.n4633 gnd.n3175 21.6691
R15926 gnd.n4650 gnd.n3157 21.6691
R15927 gnd.n4708 gnd.n4707 21.6691
R15928 gnd.n4740 gnd.n3109 21.6691
R15929 gnd.n4751 gnd.n3104 21.6691
R15930 gnd.n4785 gnd.n3083 21.6691
R15931 gnd.n4791 gnd.n3079 21.6691
R15932 gnd.n4809 gnd.n3060 21.6691
R15933 gnd.n4892 gnd.n3026 21.6691
R15934 gnd.n4819 gnd.n3015 21.6691
R15935 gnd.n4947 gnd.n3004 21.6691
R15936 gnd.n4965 gnd.n2988 21.6691
R15937 gnd.n5000 gnd.n2885 21.6691
R15938 gnd.t318 gnd.n1271 21.3504
R15939 gnd.n4170 gnd.t84 21.3504
R15940 gnd.n7402 gnd.t63 21.3504
R15941 gnd.n4551 gnd.n4550 21.0737
R15942 gnd.n5125 gnd.n5124 21.0737
R15943 gnd.n4627 gnd.n3179 21.0318
R15944 gnd.n3103 gnd.n3091 21.0318
R15945 gnd.n3095 gnd.n3092 21.0318
R15946 gnd.n4948 gnd.n3001 21.0318
R15947 gnd.t304 gnd.n978 20.7131
R15948 gnd.n4198 gnd.t20 20.7131
R15949 gnd.n3470 gnd.t156 20.7131
R15950 gnd.n2865 gnd.t309 20.7131
R15951 gnd.n5762 gnd.t41 20.7131
R15952 gnd.n4994 gnd.t208 20.3945
R15953 gnd.t291 gnd.n1013 20.0758
R15954 gnd.n4217 gnd.t26 20.0758
R15955 gnd.n5786 gnd.t33 20.0758
R15956 gnd.n3231 gnd.t250 19.8005
R15957 gnd.n3231 gnd.t206 19.8005
R15958 gnd.n3230 gnd.t231 19.8005
R15959 gnd.n3230 gnd.t280 19.8005
R15960 gnd.n2902 gnd.t290 19.8005
R15961 gnd.n2902 gnd.t247 19.8005
R15962 gnd.n2901 gnd.t185 19.8005
R15963 gnd.n2901 gnd.t265 19.8005
R15964 gnd.n4554 gnd.t249 19.7572
R15965 gnd.t6 gnd.n4644 19.7572
R15966 gnd.n4739 gnd.n4737 19.7572
R15967 gnd.n4792 gnd.n3076 19.7572
R15968 gnd.n3025 gnd.t133 19.7572
R15969 gnd.n3227 gnd.n3226 19.5087
R15970 gnd.n3240 gnd.n3227 19.5087
R15971 gnd.n3238 gnd.n3229 19.5087
R15972 gnd.n2906 gnd.n2900 19.5087
R15973 gnd.n1732 gnd.t292 19.4385
R15974 gnd.n6060 gnd.n2576 19.3944
R15975 gnd.n6060 gnd.n2577 19.3944
R15976 gnd.n6056 gnd.n2577 19.3944
R15977 gnd.n6056 gnd.n6055 19.3944
R15978 gnd.n6055 gnd.n6054 19.3944
R15979 gnd.n6054 gnd.n2583 19.3944
R15980 gnd.n6050 gnd.n2583 19.3944
R15981 gnd.n6050 gnd.n6049 19.3944
R15982 gnd.n6049 gnd.n6048 19.3944
R15983 gnd.n6048 gnd.n2588 19.3944
R15984 gnd.n6044 gnd.n2588 19.3944
R15985 gnd.n6044 gnd.n6043 19.3944
R15986 gnd.n6043 gnd.n6042 19.3944
R15987 gnd.n6042 gnd.n2593 19.3944
R15988 gnd.n6038 gnd.n2593 19.3944
R15989 gnd.n6038 gnd.n6037 19.3944
R15990 gnd.n6037 gnd.n6036 19.3944
R15991 gnd.n6036 gnd.n2598 19.3944
R15992 gnd.n6032 gnd.n2598 19.3944
R15993 gnd.n6032 gnd.n6031 19.3944
R15994 gnd.n6031 gnd.n6030 19.3944
R15995 gnd.n6030 gnd.n2603 19.3944
R15996 gnd.n6026 gnd.n2603 19.3944
R15997 gnd.n6026 gnd.n6025 19.3944
R15998 gnd.n6025 gnd.n6024 19.3944
R15999 gnd.n6024 gnd.n2608 19.3944
R16000 gnd.n6020 gnd.n2608 19.3944
R16001 gnd.n6020 gnd.n6019 19.3944
R16002 gnd.n6019 gnd.n6018 19.3944
R16003 gnd.n6018 gnd.n2613 19.3944
R16004 gnd.n6014 gnd.n2613 19.3944
R16005 gnd.n6014 gnd.n6013 19.3944
R16006 gnd.n6013 gnd.n6012 19.3944
R16007 gnd.n6012 gnd.n2618 19.3944
R16008 gnd.n6008 gnd.n2618 19.3944
R16009 gnd.n6008 gnd.n6007 19.3944
R16010 gnd.n6007 gnd.n6006 19.3944
R16011 gnd.n6006 gnd.n2623 19.3944
R16012 gnd.n6002 gnd.n2623 19.3944
R16013 gnd.n6002 gnd.n6001 19.3944
R16014 gnd.n6001 gnd.n6000 19.3944
R16015 gnd.n6000 gnd.n2628 19.3944
R16016 gnd.n5996 gnd.n2628 19.3944
R16017 gnd.n5996 gnd.n5995 19.3944
R16018 gnd.n5995 gnd.n5994 19.3944
R16019 gnd.n5994 gnd.n2633 19.3944
R16020 gnd.n5990 gnd.n2633 19.3944
R16021 gnd.n5990 gnd.n5989 19.3944
R16022 gnd.n5989 gnd.n5988 19.3944
R16023 gnd.n5988 gnd.n2638 19.3944
R16024 gnd.n5984 gnd.n2638 19.3944
R16025 gnd.n5984 gnd.n5983 19.3944
R16026 gnd.n5983 gnd.n5982 19.3944
R16027 gnd.n5982 gnd.n2643 19.3944
R16028 gnd.n5978 gnd.n2643 19.3944
R16029 gnd.n5978 gnd.n5977 19.3944
R16030 gnd.n5977 gnd.n5976 19.3944
R16031 gnd.n5976 gnd.n2648 19.3944
R16032 gnd.n5972 gnd.n2648 19.3944
R16033 gnd.n5972 gnd.n5971 19.3944
R16034 gnd.n5971 gnd.n5970 19.3944
R16035 gnd.n5970 gnd.n2653 19.3944
R16036 gnd.n5966 gnd.n2653 19.3944
R16037 gnd.n5966 gnd.n5965 19.3944
R16038 gnd.n5965 gnd.n5964 19.3944
R16039 gnd.n5964 gnd.n2658 19.3944
R16040 gnd.n5960 gnd.n2658 19.3944
R16041 gnd.n5960 gnd.n5959 19.3944
R16042 gnd.n5959 gnd.n5958 19.3944
R16043 gnd.n5958 gnd.n2663 19.3944
R16044 gnd.n5954 gnd.n2663 19.3944
R16045 gnd.n5954 gnd.n5953 19.3944
R16046 gnd.n5953 gnd.n5952 19.3944
R16047 gnd.n5952 gnd.n2668 19.3944
R16048 gnd.n5948 gnd.n2668 19.3944
R16049 gnd.n5948 gnd.n5947 19.3944
R16050 gnd.n5947 gnd.n5946 19.3944
R16051 gnd.n5946 gnd.n2673 19.3944
R16052 gnd.n5942 gnd.n2673 19.3944
R16053 gnd.n5942 gnd.n5941 19.3944
R16054 gnd.n5941 gnd.n5940 19.3944
R16055 gnd.n5940 gnd.n2678 19.3944
R16056 gnd.n3664 gnd.n2546 19.3944
R16057 gnd.n6072 gnd.n2546 19.3944
R16058 gnd.n6072 gnd.n6071 19.3944
R16059 gnd.n3579 gnd.n3420 19.3944
R16060 gnd.n3583 gnd.n3420 19.3944
R16061 gnd.n3584 gnd.n3583 19.3944
R16062 gnd.n3587 gnd.n3584 19.3944
R16063 gnd.n3587 gnd.n3416 19.3944
R16064 gnd.n3591 gnd.n3416 19.3944
R16065 gnd.n3594 gnd.n3591 19.3944
R16066 gnd.n3594 gnd.n3414 19.3944
R16067 gnd.n3600 gnd.n3414 19.3944
R16068 gnd.n3603 gnd.n3600 19.3944
R16069 gnd.n3603 gnd.n3407 19.3944
R16070 gnd.n3612 gnd.n3407 19.3944
R16071 gnd.n3615 gnd.n3612 19.3944
R16072 gnd.n3615 gnd.n3401 19.3944
R16073 gnd.n3624 gnd.n3401 19.3944
R16074 gnd.n3627 gnd.n3624 19.3944
R16075 gnd.n3627 gnd.n3395 19.3944
R16076 gnd.n3636 gnd.n3395 19.3944
R16077 gnd.n3639 gnd.n3636 19.3944
R16078 gnd.n3639 gnd.n3389 19.3944
R16079 gnd.n3648 gnd.n3389 19.3944
R16080 gnd.n3651 gnd.n3648 19.3944
R16081 gnd.n3651 gnd.n3383 19.3944
R16082 gnd.n3660 gnd.n3383 19.3944
R16083 gnd.n5316 gnd.n5315 19.3944
R16084 gnd.n5315 gnd.n2826 19.3944
R16085 gnd.n5308 gnd.n2826 19.3944
R16086 gnd.n5308 gnd.n5307 19.3944
R16087 gnd.n5307 gnd.n5217 19.3944
R16088 gnd.n5300 gnd.n5217 19.3944
R16089 gnd.n5300 gnd.n5299 19.3944
R16090 gnd.n5299 gnd.n5227 19.3944
R16091 gnd.n5292 gnd.n5227 19.3944
R16092 gnd.n5292 gnd.n5291 19.3944
R16093 gnd.n5291 gnd.n5237 19.3944
R16094 gnd.n5284 gnd.n5237 19.3944
R16095 gnd.n5284 gnd.n5283 19.3944
R16096 gnd.n5283 gnd.n5247 19.3944
R16097 gnd.n5276 gnd.n5247 19.3944
R16098 gnd.n5276 gnd.n5275 19.3944
R16099 gnd.n1447 gnd.n1446 19.3944
R16100 gnd.n1446 gnd.n1445 19.3944
R16101 gnd.n1445 gnd.n1444 19.3944
R16102 gnd.n1444 gnd.n1442 19.3944
R16103 gnd.n1442 gnd.n1439 19.3944
R16104 gnd.n1439 gnd.n1438 19.3944
R16105 gnd.n1438 gnd.n1435 19.3944
R16106 gnd.n1435 gnd.n1434 19.3944
R16107 gnd.n1434 gnd.n1431 19.3944
R16108 gnd.n1431 gnd.n1430 19.3944
R16109 gnd.n1430 gnd.n1427 19.3944
R16110 gnd.n1427 gnd.n1426 19.3944
R16111 gnd.n1426 gnd.n1423 19.3944
R16112 gnd.n1423 gnd.n1422 19.3944
R16113 gnd.n1422 gnd.n1419 19.3944
R16114 gnd.n1419 gnd.n1418 19.3944
R16115 gnd.n1418 gnd.n1415 19.3944
R16116 gnd.n1415 gnd.n1414 19.3944
R16117 gnd.n1414 gnd.n1411 19.3944
R16118 gnd.n1411 gnd.n1410 19.3944
R16119 gnd.n1410 gnd.n1407 19.3944
R16120 gnd.n1407 gnd.n1406 19.3944
R16121 gnd.n1403 gnd.n1402 19.3944
R16122 gnd.n1402 gnd.n1358 19.3944
R16123 gnd.n1453 gnd.n1358 19.3944
R16124 gnd.n2221 gnd.n2220 19.3944
R16125 gnd.n2220 gnd.n2217 19.3944
R16126 gnd.n2217 gnd.n2216 19.3944
R16127 gnd.n2266 gnd.n2265 19.3944
R16128 gnd.n2265 gnd.n2264 19.3944
R16129 gnd.n2264 gnd.n2261 19.3944
R16130 gnd.n2261 gnd.n2260 19.3944
R16131 gnd.n2260 gnd.n2257 19.3944
R16132 gnd.n2257 gnd.n2256 19.3944
R16133 gnd.n2256 gnd.n2253 19.3944
R16134 gnd.n2253 gnd.n2252 19.3944
R16135 gnd.n2252 gnd.n2249 19.3944
R16136 gnd.n2249 gnd.n2248 19.3944
R16137 gnd.n2248 gnd.n2245 19.3944
R16138 gnd.n2245 gnd.n2244 19.3944
R16139 gnd.n2244 gnd.n2241 19.3944
R16140 gnd.n2241 gnd.n2240 19.3944
R16141 gnd.n2240 gnd.n2237 19.3944
R16142 gnd.n2237 gnd.n2236 19.3944
R16143 gnd.n2236 gnd.n2233 19.3944
R16144 gnd.n2233 gnd.n2232 19.3944
R16145 gnd.n2232 gnd.n2229 19.3944
R16146 gnd.n2229 gnd.n2228 19.3944
R16147 gnd.n2228 gnd.n2225 19.3944
R16148 gnd.n2225 gnd.n2224 19.3944
R16149 gnd.n1546 gnd.n1255 19.3944
R16150 gnd.n1556 gnd.n1255 19.3944
R16151 gnd.n1557 gnd.n1556 19.3944
R16152 gnd.n1557 gnd.n1236 19.3944
R16153 gnd.n1577 gnd.n1236 19.3944
R16154 gnd.n1577 gnd.n1228 19.3944
R16155 gnd.n1587 gnd.n1228 19.3944
R16156 gnd.n1588 gnd.n1587 19.3944
R16157 gnd.n1589 gnd.n1588 19.3944
R16158 gnd.n1589 gnd.n1211 19.3944
R16159 gnd.n1606 gnd.n1211 19.3944
R16160 gnd.n1609 gnd.n1606 19.3944
R16161 gnd.n1609 gnd.n1608 19.3944
R16162 gnd.n1608 gnd.n1184 19.3944
R16163 gnd.n1648 gnd.n1184 19.3944
R16164 gnd.n1648 gnd.n1181 19.3944
R16165 gnd.n1654 gnd.n1181 19.3944
R16166 gnd.n1655 gnd.n1654 19.3944
R16167 gnd.n1655 gnd.n1179 19.3944
R16168 gnd.n1661 gnd.n1179 19.3944
R16169 gnd.n1664 gnd.n1661 19.3944
R16170 gnd.n1666 gnd.n1664 19.3944
R16171 gnd.n1672 gnd.n1666 19.3944
R16172 gnd.n1672 gnd.n1671 19.3944
R16173 gnd.n1671 gnd.n1054 19.3944
R16174 gnd.n1738 gnd.n1054 19.3944
R16175 gnd.n1739 gnd.n1738 19.3944
R16176 gnd.n1739 gnd.n1047 19.3944
R16177 gnd.n1750 gnd.n1047 19.3944
R16178 gnd.n1751 gnd.n1750 19.3944
R16179 gnd.n1751 gnd.n1030 19.3944
R16180 gnd.n1030 gnd.n1028 19.3944
R16181 gnd.n1775 gnd.n1028 19.3944
R16182 gnd.n1776 gnd.n1775 19.3944
R16183 gnd.n1776 gnd.n1000 19.3944
R16184 gnd.n1825 gnd.n1000 19.3944
R16185 gnd.n1826 gnd.n1825 19.3944
R16186 gnd.n1826 gnd.n993 19.3944
R16187 gnd.n1837 gnd.n993 19.3944
R16188 gnd.n1838 gnd.n1837 19.3944
R16189 gnd.n1838 gnd.n976 19.3944
R16190 gnd.n976 gnd.n974 19.3944
R16191 gnd.n1862 gnd.n974 19.3944
R16192 gnd.n1863 gnd.n1862 19.3944
R16193 gnd.n1863 gnd.n946 19.3944
R16194 gnd.n1914 gnd.n946 19.3944
R16195 gnd.n1915 gnd.n1914 19.3944
R16196 gnd.n1915 gnd.n939 19.3944
R16197 gnd.n2182 gnd.n939 19.3944
R16198 gnd.n2183 gnd.n2182 19.3944
R16199 gnd.n2183 gnd.n920 19.3944
R16200 gnd.n2208 gnd.n920 19.3944
R16201 gnd.n2208 gnd.n921 19.3944
R16202 gnd.n1537 gnd.n1536 19.3944
R16203 gnd.n1536 gnd.n1269 19.3944
R16204 gnd.n1292 gnd.n1269 19.3944
R16205 gnd.n1295 gnd.n1292 19.3944
R16206 gnd.n1295 gnd.n1288 19.3944
R16207 gnd.n1299 gnd.n1288 19.3944
R16208 gnd.n1302 gnd.n1299 19.3944
R16209 gnd.n1305 gnd.n1302 19.3944
R16210 gnd.n1305 gnd.n1286 19.3944
R16211 gnd.n1309 gnd.n1286 19.3944
R16212 gnd.n1312 gnd.n1309 19.3944
R16213 gnd.n1315 gnd.n1312 19.3944
R16214 gnd.n1315 gnd.n1284 19.3944
R16215 gnd.n1319 gnd.n1284 19.3944
R16216 gnd.n1542 gnd.n1541 19.3944
R16217 gnd.n1541 gnd.n1245 19.3944
R16218 gnd.n1567 gnd.n1245 19.3944
R16219 gnd.n1567 gnd.n1243 19.3944
R16220 gnd.n1573 gnd.n1243 19.3944
R16221 gnd.n1573 gnd.n1572 19.3944
R16222 gnd.n1572 gnd.n1217 19.3944
R16223 gnd.n1597 gnd.n1217 19.3944
R16224 gnd.n1597 gnd.n1215 19.3944
R16225 gnd.n1601 gnd.n1215 19.3944
R16226 gnd.n1601 gnd.n1195 19.3944
R16227 gnd.n1628 gnd.n1195 19.3944
R16228 gnd.n1628 gnd.n1193 19.3944
R16229 gnd.n1638 gnd.n1193 19.3944
R16230 gnd.n1638 gnd.n1637 19.3944
R16231 gnd.n1637 gnd.n1636 19.3944
R16232 gnd.n1636 gnd.n1142 19.3944
R16233 gnd.n1686 gnd.n1142 19.3944
R16234 gnd.n1686 gnd.n1685 19.3944
R16235 gnd.n1685 gnd.n1684 19.3944
R16236 gnd.n1684 gnd.n1146 19.3944
R16237 gnd.n1166 gnd.n1146 19.3944
R16238 gnd.n1166 gnd.n1064 19.3944
R16239 gnd.n1723 gnd.n1064 19.3944
R16240 gnd.n1723 gnd.n1062 19.3944
R16241 gnd.n1729 gnd.n1062 19.3944
R16242 gnd.n1729 gnd.n1728 19.3944
R16243 gnd.n1728 gnd.n1037 19.3944
R16244 gnd.n1763 gnd.n1037 19.3944
R16245 gnd.n1763 gnd.n1035 19.3944
R16246 gnd.n1769 gnd.n1035 19.3944
R16247 gnd.n1769 gnd.n1768 19.3944
R16248 gnd.n1768 gnd.n1011 19.3944
R16249 gnd.n1810 gnd.n1011 19.3944
R16250 gnd.n1810 gnd.n1009 19.3944
R16251 gnd.n1816 gnd.n1009 19.3944
R16252 gnd.n1816 gnd.n1815 19.3944
R16253 gnd.n1815 gnd.n983 19.3944
R16254 gnd.n1850 gnd.n983 19.3944
R16255 gnd.n1850 gnd.n981 19.3944
R16256 gnd.n1856 gnd.n981 19.3944
R16257 gnd.n1856 gnd.n1855 19.3944
R16258 gnd.n1855 gnd.n956 19.3944
R16259 gnd.n1899 gnd.n956 19.3944
R16260 gnd.n1899 gnd.n954 19.3944
R16261 gnd.n1905 gnd.n954 19.3944
R16262 gnd.n1905 gnd.n1904 19.3944
R16263 gnd.n1904 gnd.n929 19.3944
R16264 gnd.n2193 gnd.n929 19.3944
R16265 gnd.n2193 gnd.n927 19.3944
R16266 gnd.n2201 gnd.n927 19.3944
R16267 gnd.n2201 gnd.n2200 19.3944
R16268 gnd.n2200 gnd.n2199 19.3944
R16269 gnd.n2302 gnd.n2301 19.3944
R16270 gnd.n2301 gnd.n868 19.3944
R16271 gnd.n2297 gnd.n868 19.3944
R16272 gnd.n2297 gnd.n2294 19.3944
R16273 gnd.n2294 gnd.n2291 19.3944
R16274 gnd.n2291 gnd.n2290 19.3944
R16275 gnd.n2290 gnd.n2287 19.3944
R16276 gnd.n2287 gnd.n2286 19.3944
R16277 gnd.n2286 gnd.n2283 19.3944
R16278 gnd.n2283 gnd.n2282 19.3944
R16279 gnd.n2282 gnd.n2279 19.3944
R16280 gnd.n2279 gnd.n2278 19.3944
R16281 gnd.n2278 gnd.n2275 19.3944
R16282 gnd.n2275 gnd.n2274 19.3944
R16283 gnd.n1457 gnd.n1356 19.3944
R16284 gnd.n1457 gnd.n1347 19.3944
R16285 gnd.n1470 gnd.n1347 19.3944
R16286 gnd.n1470 gnd.n1345 19.3944
R16287 gnd.n1474 gnd.n1345 19.3944
R16288 gnd.n1474 gnd.n1335 19.3944
R16289 gnd.n1486 gnd.n1335 19.3944
R16290 gnd.n1486 gnd.n1333 19.3944
R16291 gnd.n1520 gnd.n1333 19.3944
R16292 gnd.n1520 gnd.n1519 19.3944
R16293 gnd.n1519 gnd.n1518 19.3944
R16294 gnd.n1518 gnd.n1517 19.3944
R16295 gnd.n1517 gnd.n1514 19.3944
R16296 gnd.n1514 gnd.n1513 19.3944
R16297 gnd.n1513 gnd.n1512 19.3944
R16298 gnd.n1512 gnd.n1510 19.3944
R16299 gnd.n1510 gnd.n1509 19.3944
R16300 gnd.n1509 gnd.n1506 19.3944
R16301 gnd.n1506 gnd.n1505 19.3944
R16302 gnd.n1505 gnd.n1504 19.3944
R16303 gnd.n1504 gnd.n1502 19.3944
R16304 gnd.n1502 gnd.n1201 19.3944
R16305 gnd.n1617 gnd.n1201 19.3944
R16306 gnd.n1617 gnd.n1199 19.3944
R16307 gnd.n1623 gnd.n1199 19.3944
R16308 gnd.n1623 gnd.n1622 19.3944
R16309 gnd.n1622 gnd.n1123 19.3944
R16310 gnd.n1697 gnd.n1123 19.3944
R16311 gnd.n1697 gnd.n1124 19.3944
R16312 gnd.n1171 gnd.n1170 19.3944
R16313 gnd.n1174 gnd.n1173 19.3944
R16314 gnd.n1161 gnd.n1160 19.3944
R16315 gnd.n1716 gnd.n1069 19.3944
R16316 gnd.n1716 gnd.n1715 19.3944
R16317 gnd.n1715 gnd.n1714 19.3944
R16318 gnd.n1714 gnd.n1712 19.3944
R16319 gnd.n1712 gnd.n1711 19.3944
R16320 gnd.n1711 gnd.n1709 19.3944
R16321 gnd.n1709 gnd.n1708 19.3944
R16322 gnd.n1708 gnd.n1018 19.3944
R16323 gnd.n1784 gnd.n1018 19.3944
R16324 gnd.n1784 gnd.n1016 19.3944
R16325 gnd.n1803 gnd.n1016 19.3944
R16326 gnd.n1803 gnd.n1802 19.3944
R16327 gnd.n1802 gnd.n1801 19.3944
R16328 gnd.n1801 gnd.n1799 19.3944
R16329 gnd.n1799 gnd.n1798 19.3944
R16330 gnd.n1798 gnd.n1796 19.3944
R16331 gnd.n1796 gnd.n1795 19.3944
R16332 gnd.n1795 gnd.n963 19.3944
R16333 gnd.n1871 gnd.n963 19.3944
R16334 gnd.n1871 gnd.n961 19.3944
R16335 gnd.n1894 gnd.n961 19.3944
R16336 gnd.n1894 gnd.n1893 19.3944
R16337 gnd.n1893 gnd.n1892 19.3944
R16338 gnd.n1892 gnd.n1889 19.3944
R16339 gnd.n1889 gnd.n1888 19.3944
R16340 gnd.n1888 gnd.n1886 19.3944
R16341 gnd.n1886 gnd.n1885 19.3944
R16342 gnd.n1885 gnd.n1883 19.3944
R16343 gnd.n1883 gnd.n915 19.3944
R16344 gnd.n1462 gnd.n1352 19.3944
R16345 gnd.n1462 gnd.n1350 19.3944
R16346 gnd.n1466 gnd.n1350 19.3944
R16347 gnd.n1466 gnd.n1341 19.3944
R16348 gnd.n1478 gnd.n1341 19.3944
R16349 gnd.n1478 gnd.n1339 19.3944
R16350 gnd.n1482 gnd.n1339 19.3944
R16351 gnd.n1482 gnd.n1328 19.3944
R16352 gnd.n1524 gnd.n1328 19.3944
R16353 gnd.n1524 gnd.n1282 19.3944
R16354 gnd.n1530 gnd.n1282 19.3944
R16355 gnd.n1530 gnd.n1529 19.3944
R16356 gnd.n1529 gnd.n1260 19.3944
R16357 gnd.n1551 gnd.n1260 19.3944
R16358 gnd.n1551 gnd.n1253 19.3944
R16359 gnd.n1562 gnd.n1253 19.3944
R16360 gnd.n1562 gnd.n1561 19.3944
R16361 gnd.n1561 gnd.n1234 19.3944
R16362 gnd.n1582 gnd.n1234 19.3944
R16363 gnd.n1582 gnd.n1224 19.3944
R16364 gnd.n1592 gnd.n1224 19.3944
R16365 gnd.n1592 gnd.n1207 19.3944
R16366 gnd.n1613 gnd.n1207 19.3944
R16367 gnd.n1613 gnd.n1612 19.3944
R16368 gnd.n1612 gnd.n1186 19.3944
R16369 gnd.n1643 gnd.n1186 19.3944
R16370 gnd.n1643 gnd.n1131 19.3944
R16371 gnd.n1693 gnd.n1131 19.3944
R16372 gnd.n1693 gnd.n1692 19.3944
R16373 gnd.n1692 gnd.n1691 19.3944
R16374 gnd.n1691 gnd.n1135 19.3944
R16375 gnd.n1153 gnd.n1135 19.3944
R16376 gnd.n1679 gnd.n1153 19.3944
R16377 gnd.n1679 gnd.n1678 19.3944
R16378 gnd.n1678 gnd.n1677 19.3944
R16379 gnd.n1677 gnd.n1157 19.3944
R16380 gnd.n1157 gnd.n1056 19.3944
R16381 gnd.n1734 gnd.n1056 19.3944
R16382 gnd.n1734 gnd.n1049 19.3944
R16383 gnd.n1745 gnd.n1049 19.3944
R16384 gnd.n1745 gnd.n1045 19.3944
R16385 gnd.n1758 gnd.n1045 19.3944
R16386 gnd.n1758 gnd.n1757 19.3944
R16387 gnd.n1757 gnd.n1024 19.3944
R16388 gnd.n1780 gnd.n1024 19.3944
R16389 gnd.n1780 gnd.n1779 19.3944
R16390 gnd.n1779 gnd.n1002 19.3944
R16391 gnd.n1821 gnd.n1002 19.3944
R16392 gnd.n1821 gnd.n995 19.3944
R16393 gnd.n1832 gnd.n995 19.3944
R16394 gnd.n1832 gnd.n991 19.3944
R16395 gnd.n1845 gnd.n991 19.3944
R16396 gnd.n1845 gnd.n1844 19.3944
R16397 gnd.n1844 gnd.n970 19.3944
R16398 gnd.n1867 gnd.n970 19.3944
R16399 gnd.n1867 gnd.n1866 19.3944
R16400 gnd.n1866 gnd.n948 19.3944
R16401 gnd.n1910 gnd.n948 19.3944
R16402 gnd.n1910 gnd.n941 19.3944
R16403 gnd.n1921 gnd.n941 19.3944
R16404 gnd.n1921 gnd.n937 19.3944
R16405 gnd.n2188 gnd.n937 19.3944
R16406 gnd.n2188 gnd.n2187 19.3944
R16407 gnd.n2187 gnd.n918 19.3944
R16408 gnd.n2211 gnd.n918 19.3944
R16409 gnd.n3597 gnd.n3412 19.3944
R16410 gnd.n3606 gnd.n3412 19.3944
R16411 gnd.n3609 gnd.n3606 19.3944
R16412 gnd.n3609 gnd.n3403 19.3944
R16413 gnd.n3618 gnd.n3403 19.3944
R16414 gnd.n3621 gnd.n3618 19.3944
R16415 gnd.n3621 gnd.n3399 19.3944
R16416 gnd.n3630 gnd.n3399 19.3944
R16417 gnd.n3633 gnd.n3630 19.3944
R16418 gnd.n3633 gnd.n3391 19.3944
R16419 gnd.n3642 gnd.n3391 19.3944
R16420 gnd.n3645 gnd.n3642 19.3944
R16421 gnd.n3645 gnd.n3387 19.3944
R16422 gnd.n3654 gnd.n3387 19.3944
R16423 gnd.n3657 gnd.n3654 19.3944
R16424 gnd.n3657 gnd.n3377 19.3944
R16425 gnd.n6893 gnd.n379 19.3944
R16426 gnd.n6897 gnd.n379 19.3944
R16427 gnd.n6897 gnd.n375 19.3944
R16428 gnd.n6903 gnd.n375 19.3944
R16429 gnd.n6903 gnd.n373 19.3944
R16430 gnd.n6907 gnd.n373 19.3944
R16431 gnd.n6907 gnd.n369 19.3944
R16432 gnd.n6913 gnd.n369 19.3944
R16433 gnd.n6913 gnd.n367 19.3944
R16434 gnd.n6917 gnd.n367 19.3944
R16435 gnd.n6917 gnd.n363 19.3944
R16436 gnd.n6923 gnd.n363 19.3944
R16437 gnd.n6923 gnd.n361 19.3944
R16438 gnd.n6927 gnd.n361 19.3944
R16439 gnd.n6927 gnd.n357 19.3944
R16440 gnd.n6933 gnd.n357 19.3944
R16441 gnd.n6933 gnd.n355 19.3944
R16442 gnd.n6937 gnd.n355 19.3944
R16443 gnd.n6937 gnd.n351 19.3944
R16444 gnd.n6943 gnd.n351 19.3944
R16445 gnd.n6943 gnd.n349 19.3944
R16446 gnd.n6947 gnd.n349 19.3944
R16447 gnd.n6947 gnd.n345 19.3944
R16448 gnd.n6953 gnd.n345 19.3944
R16449 gnd.n6953 gnd.n343 19.3944
R16450 gnd.n6957 gnd.n343 19.3944
R16451 gnd.n6957 gnd.n339 19.3944
R16452 gnd.n6963 gnd.n339 19.3944
R16453 gnd.n6963 gnd.n337 19.3944
R16454 gnd.n6967 gnd.n337 19.3944
R16455 gnd.n6967 gnd.n333 19.3944
R16456 gnd.n6973 gnd.n333 19.3944
R16457 gnd.n6973 gnd.n331 19.3944
R16458 gnd.n6977 gnd.n331 19.3944
R16459 gnd.n6977 gnd.n327 19.3944
R16460 gnd.n6983 gnd.n327 19.3944
R16461 gnd.n6983 gnd.n325 19.3944
R16462 gnd.n6987 gnd.n325 19.3944
R16463 gnd.n6987 gnd.n321 19.3944
R16464 gnd.n6993 gnd.n321 19.3944
R16465 gnd.n6993 gnd.n319 19.3944
R16466 gnd.n6997 gnd.n319 19.3944
R16467 gnd.n6997 gnd.n315 19.3944
R16468 gnd.n7003 gnd.n315 19.3944
R16469 gnd.n7003 gnd.n313 19.3944
R16470 gnd.n7007 gnd.n313 19.3944
R16471 gnd.n7007 gnd.n309 19.3944
R16472 gnd.n7013 gnd.n309 19.3944
R16473 gnd.n7013 gnd.n307 19.3944
R16474 gnd.n7017 gnd.n307 19.3944
R16475 gnd.n7017 gnd.n303 19.3944
R16476 gnd.n7023 gnd.n303 19.3944
R16477 gnd.n7023 gnd.n301 19.3944
R16478 gnd.n7027 gnd.n301 19.3944
R16479 gnd.n7027 gnd.n297 19.3944
R16480 gnd.n7033 gnd.n297 19.3944
R16481 gnd.n7033 gnd.n295 19.3944
R16482 gnd.n7037 gnd.n295 19.3944
R16483 gnd.n7037 gnd.n291 19.3944
R16484 gnd.n7043 gnd.n291 19.3944
R16485 gnd.n7043 gnd.n289 19.3944
R16486 gnd.n7047 gnd.n289 19.3944
R16487 gnd.n7047 gnd.n285 19.3944
R16488 gnd.n7053 gnd.n285 19.3944
R16489 gnd.n7053 gnd.n283 19.3944
R16490 gnd.n7057 gnd.n283 19.3944
R16491 gnd.n7057 gnd.n279 19.3944
R16492 gnd.n7063 gnd.n279 19.3944
R16493 gnd.n7063 gnd.n277 19.3944
R16494 gnd.n7067 gnd.n277 19.3944
R16495 gnd.n7067 gnd.n273 19.3944
R16496 gnd.n7073 gnd.n273 19.3944
R16497 gnd.n7073 gnd.n271 19.3944
R16498 gnd.n7077 gnd.n271 19.3944
R16499 gnd.n7077 gnd.n267 19.3944
R16500 gnd.n7083 gnd.n267 19.3944
R16501 gnd.n7083 gnd.n265 19.3944
R16502 gnd.n7087 gnd.n265 19.3944
R16503 gnd.n7087 gnd.n261 19.3944
R16504 gnd.n7093 gnd.n261 19.3944
R16505 gnd.n7093 gnd.n259 19.3944
R16506 gnd.n7097 gnd.n259 19.3944
R16507 gnd.n7097 gnd.n255 19.3944
R16508 gnd.n7103 gnd.n255 19.3944
R16509 gnd.n6406 gnd.n672 19.3944
R16510 gnd.n6406 gnd.n668 19.3944
R16511 gnd.n6412 gnd.n668 19.3944
R16512 gnd.n6412 gnd.n666 19.3944
R16513 gnd.n6416 gnd.n666 19.3944
R16514 gnd.n6416 gnd.n662 19.3944
R16515 gnd.n6422 gnd.n662 19.3944
R16516 gnd.n6422 gnd.n660 19.3944
R16517 gnd.n6426 gnd.n660 19.3944
R16518 gnd.n6426 gnd.n656 19.3944
R16519 gnd.n6432 gnd.n656 19.3944
R16520 gnd.n6432 gnd.n654 19.3944
R16521 gnd.n6436 gnd.n654 19.3944
R16522 gnd.n6436 gnd.n650 19.3944
R16523 gnd.n6442 gnd.n650 19.3944
R16524 gnd.n6442 gnd.n648 19.3944
R16525 gnd.n6446 gnd.n648 19.3944
R16526 gnd.n6446 gnd.n644 19.3944
R16527 gnd.n6452 gnd.n644 19.3944
R16528 gnd.n6452 gnd.n642 19.3944
R16529 gnd.n6456 gnd.n642 19.3944
R16530 gnd.n6456 gnd.n638 19.3944
R16531 gnd.n6462 gnd.n638 19.3944
R16532 gnd.n6462 gnd.n636 19.3944
R16533 gnd.n6466 gnd.n636 19.3944
R16534 gnd.n6466 gnd.n632 19.3944
R16535 gnd.n6472 gnd.n632 19.3944
R16536 gnd.n6472 gnd.n630 19.3944
R16537 gnd.n6476 gnd.n630 19.3944
R16538 gnd.n6476 gnd.n626 19.3944
R16539 gnd.n6482 gnd.n626 19.3944
R16540 gnd.n6482 gnd.n624 19.3944
R16541 gnd.n6486 gnd.n624 19.3944
R16542 gnd.n6486 gnd.n620 19.3944
R16543 gnd.n6492 gnd.n620 19.3944
R16544 gnd.n6492 gnd.n618 19.3944
R16545 gnd.n6496 gnd.n618 19.3944
R16546 gnd.n6496 gnd.n614 19.3944
R16547 gnd.n6502 gnd.n614 19.3944
R16548 gnd.n6502 gnd.n612 19.3944
R16549 gnd.n6506 gnd.n612 19.3944
R16550 gnd.n6506 gnd.n608 19.3944
R16551 gnd.n6512 gnd.n608 19.3944
R16552 gnd.n6512 gnd.n606 19.3944
R16553 gnd.n6516 gnd.n606 19.3944
R16554 gnd.n6516 gnd.n602 19.3944
R16555 gnd.n6522 gnd.n602 19.3944
R16556 gnd.n6522 gnd.n600 19.3944
R16557 gnd.n6526 gnd.n600 19.3944
R16558 gnd.n6526 gnd.n596 19.3944
R16559 gnd.n6532 gnd.n596 19.3944
R16560 gnd.n6532 gnd.n594 19.3944
R16561 gnd.n6536 gnd.n594 19.3944
R16562 gnd.n6536 gnd.n590 19.3944
R16563 gnd.n6542 gnd.n590 19.3944
R16564 gnd.n6542 gnd.n588 19.3944
R16565 gnd.n6546 gnd.n588 19.3944
R16566 gnd.n6546 gnd.n584 19.3944
R16567 gnd.n6552 gnd.n584 19.3944
R16568 gnd.n6552 gnd.n582 19.3944
R16569 gnd.n6556 gnd.n582 19.3944
R16570 gnd.n6556 gnd.n578 19.3944
R16571 gnd.n6562 gnd.n578 19.3944
R16572 gnd.n6562 gnd.n576 19.3944
R16573 gnd.n6566 gnd.n576 19.3944
R16574 gnd.n6566 gnd.n572 19.3944
R16575 gnd.n6572 gnd.n572 19.3944
R16576 gnd.n6572 gnd.n570 19.3944
R16577 gnd.n6576 gnd.n570 19.3944
R16578 gnd.n6576 gnd.n566 19.3944
R16579 gnd.n6582 gnd.n566 19.3944
R16580 gnd.n6582 gnd.n564 19.3944
R16581 gnd.n6586 gnd.n564 19.3944
R16582 gnd.n6586 gnd.n560 19.3944
R16583 gnd.n6592 gnd.n560 19.3944
R16584 gnd.n6592 gnd.n558 19.3944
R16585 gnd.n6596 gnd.n558 19.3944
R16586 gnd.n6596 gnd.n554 19.3944
R16587 gnd.n6602 gnd.n554 19.3944
R16588 gnd.n6602 gnd.n552 19.3944
R16589 gnd.n6606 gnd.n552 19.3944
R16590 gnd.n6606 gnd.n548 19.3944
R16591 gnd.n6612 gnd.n548 19.3944
R16592 gnd.n6612 gnd.n546 19.3944
R16593 gnd.n6616 gnd.n546 19.3944
R16594 gnd.n6616 gnd.n542 19.3944
R16595 gnd.n6622 gnd.n542 19.3944
R16596 gnd.n6622 gnd.n540 19.3944
R16597 gnd.n6626 gnd.n540 19.3944
R16598 gnd.n6626 gnd.n536 19.3944
R16599 gnd.n6632 gnd.n536 19.3944
R16600 gnd.n6632 gnd.n534 19.3944
R16601 gnd.n6636 gnd.n534 19.3944
R16602 gnd.n6636 gnd.n530 19.3944
R16603 gnd.n6642 gnd.n530 19.3944
R16604 gnd.n6642 gnd.n528 19.3944
R16605 gnd.n6646 gnd.n528 19.3944
R16606 gnd.n6646 gnd.n524 19.3944
R16607 gnd.n6652 gnd.n524 19.3944
R16608 gnd.n6652 gnd.n522 19.3944
R16609 gnd.n6656 gnd.n522 19.3944
R16610 gnd.n6656 gnd.n518 19.3944
R16611 gnd.n6662 gnd.n518 19.3944
R16612 gnd.n6662 gnd.n516 19.3944
R16613 gnd.n6666 gnd.n516 19.3944
R16614 gnd.n6666 gnd.n512 19.3944
R16615 gnd.n6672 gnd.n512 19.3944
R16616 gnd.n6672 gnd.n510 19.3944
R16617 gnd.n6676 gnd.n510 19.3944
R16618 gnd.n6676 gnd.n506 19.3944
R16619 gnd.n6682 gnd.n506 19.3944
R16620 gnd.n6682 gnd.n504 19.3944
R16621 gnd.n6686 gnd.n504 19.3944
R16622 gnd.n6686 gnd.n500 19.3944
R16623 gnd.n6692 gnd.n500 19.3944
R16624 gnd.n6692 gnd.n498 19.3944
R16625 gnd.n6696 gnd.n498 19.3944
R16626 gnd.n6696 gnd.n494 19.3944
R16627 gnd.n6702 gnd.n494 19.3944
R16628 gnd.n6702 gnd.n492 19.3944
R16629 gnd.n6706 gnd.n492 19.3944
R16630 gnd.n6706 gnd.n488 19.3944
R16631 gnd.n6712 gnd.n488 19.3944
R16632 gnd.n6712 gnd.n486 19.3944
R16633 gnd.n6716 gnd.n486 19.3944
R16634 gnd.n6716 gnd.n482 19.3944
R16635 gnd.n6722 gnd.n482 19.3944
R16636 gnd.n6722 gnd.n480 19.3944
R16637 gnd.n6726 gnd.n480 19.3944
R16638 gnd.n6726 gnd.n476 19.3944
R16639 gnd.n6732 gnd.n476 19.3944
R16640 gnd.n6732 gnd.n474 19.3944
R16641 gnd.n6736 gnd.n474 19.3944
R16642 gnd.n6736 gnd.n470 19.3944
R16643 gnd.n6742 gnd.n470 19.3944
R16644 gnd.n6742 gnd.n468 19.3944
R16645 gnd.n6746 gnd.n468 19.3944
R16646 gnd.n6746 gnd.n464 19.3944
R16647 gnd.n6752 gnd.n464 19.3944
R16648 gnd.n6752 gnd.n462 19.3944
R16649 gnd.n6756 gnd.n462 19.3944
R16650 gnd.n6756 gnd.n458 19.3944
R16651 gnd.n6762 gnd.n458 19.3944
R16652 gnd.n6762 gnd.n456 19.3944
R16653 gnd.n6766 gnd.n456 19.3944
R16654 gnd.n6766 gnd.n452 19.3944
R16655 gnd.n6772 gnd.n452 19.3944
R16656 gnd.n6772 gnd.n450 19.3944
R16657 gnd.n6776 gnd.n450 19.3944
R16658 gnd.n6776 gnd.n446 19.3944
R16659 gnd.n6782 gnd.n446 19.3944
R16660 gnd.n6782 gnd.n444 19.3944
R16661 gnd.n6786 gnd.n444 19.3944
R16662 gnd.n6786 gnd.n440 19.3944
R16663 gnd.n6792 gnd.n440 19.3944
R16664 gnd.n6792 gnd.n438 19.3944
R16665 gnd.n6796 gnd.n438 19.3944
R16666 gnd.n6796 gnd.n434 19.3944
R16667 gnd.n6802 gnd.n434 19.3944
R16668 gnd.n6802 gnd.n432 19.3944
R16669 gnd.n6806 gnd.n432 19.3944
R16670 gnd.n6806 gnd.n428 19.3944
R16671 gnd.n6812 gnd.n428 19.3944
R16672 gnd.n6812 gnd.n426 19.3944
R16673 gnd.n6816 gnd.n426 19.3944
R16674 gnd.n6816 gnd.n422 19.3944
R16675 gnd.n6822 gnd.n422 19.3944
R16676 gnd.n6822 gnd.n420 19.3944
R16677 gnd.n6826 gnd.n420 19.3944
R16678 gnd.n6826 gnd.n416 19.3944
R16679 gnd.n6832 gnd.n416 19.3944
R16680 gnd.n6832 gnd.n414 19.3944
R16681 gnd.n6836 gnd.n414 19.3944
R16682 gnd.n6836 gnd.n410 19.3944
R16683 gnd.n6842 gnd.n410 19.3944
R16684 gnd.n6842 gnd.n408 19.3944
R16685 gnd.n6846 gnd.n408 19.3944
R16686 gnd.n6846 gnd.n404 19.3944
R16687 gnd.n6852 gnd.n404 19.3944
R16688 gnd.n6852 gnd.n402 19.3944
R16689 gnd.n6856 gnd.n402 19.3944
R16690 gnd.n6856 gnd.n398 19.3944
R16691 gnd.n6862 gnd.n398 19.3944
R16692 gnd.n6862 gnd.n396 19.3944
R16693 gnd.n6866 gnd.n396 19.3944
R16694 gnd.n6866 gnd.n392 19.3944
R16695 gnd.n6872 gnd.n392 19.3944
R16696 gnd.n6872 gnd.n390 19.3944
R16697 gnd.n6876 gnd.n390 19.3944
R16698 gnd.n6876 gnd.n386 19.3944
R16699 gnd.n6882 gnd.n386 19.3944
R16700 gnd.n6882 gnd.n384 19.3944
R16701 gnd.n6887 gnd.n384 19.3944
R16702 gnd.n6887 gnd.n6886 19.3944
R16703 gnd.n5924 gnd.n5923 19.3944
R16704 gnd.n5923 gnd.n5922 19.3944
R16705 gnd.n5922 gnd.n5921 19.3944
R16706 gnd.n5921 gnd.n5919 19.3944
R16707 gnd.n5919 gnd.n5916 19.3944
R16708 gnd.n5916 gnd.n5915 19.3944
R16709 gnd.n5915 gnd.n5912 19.3944
R16710 gnd.n5912 gnd.n5911 19.3944
R16711 gnd.n5911 gnd.n5908 19.3944
R16712 gnd.n5908 gnd.n5907 19.3944
R16713 gnd.n5907 gnd.n5904 19.3944
R16714 gnd.n5904 gnd.n5903 19.3944
R16715 gnd.n5903 gnd.n5900 19.3944
R16716 gnd.n5900 gnd.n5899 19.3944
R16717 gnd.n5899 gnd.n5896 19.3944
R16718 gnd.n5896 gnd.n5895 19.3944
R16719 gnd.n5895 gnd.n5892 19.3944
R16720 gnd.n5890 gnd.n5887 19.3944
R16721 gnd.n5887 gnd.n5886 19.3944
R16722 gnd.n5886 gnd.n5883 19.3944
R16723 gnd.n5883 gnd.n5882 19.3944
R16724 gnd.n5882 gnd.n5879 19.3944
R16725 gnd.n5879 gnd.n5878 19.3944
R16726 gnd.n5878 gnd.n5875 19.3944
R16727 gnd.n5873 gnd.n5870 19.3944
R16728 gnd.n5870 gnd.n5869 19.3944
R16729 gnd.n5869 gnd.n5866 19.3944
R16730 gnd.n5866 gnd.n5865 19.3944
R16731 gnd.n5865 gnd.n5862 19.3944
R16732 gnd.n5862 gnd.n5861 19.3944
R16733 gnd.n5861 gnd.n5858 19.3944
R16734 gnd.n5858 gnd.n5857 19.3944
R16735 gnd.n5853 gnd.n5850 19.3944
R16736 gnd.n5850 gnd.n5849 19.3944
R16737 gnd.n5849 gnd.n5846 19.3944
R16738 gnd.n5846 gnd.n5845 19.3944
R16739 gnd.n5845 gnd.n5842 19.3944
R16740 gnd.n5842 gnd.n5841 19.3944
R16741 gnd.n5841 gnd.n5838 19.3944
R16742 gnd.n5838 gnd.n5837 19.3944
R16743 gnd.n5837 gnd.n5834 19.3944
R16744 gnd.n5834 gnd.n5833 19.3944
R16745 gnd.n5833 gnd.n5830 19.3944
R16746 gnd.n5830 gnd.n5829 19.3944
R16747 gnd.n5829 gnd.n5826 19.3944
R16748 gnd.n5826 gnd.n5825 19.3944
R16749 gnd.n5825 gnd.n5822 19.3944
R16750 gnd.n5822 gnd.n5821 19.3944
R16751 gnd.n5821 gnd.n5818 19.3944
R16752 gnd.n5818 gnd.n5817 19.3944
R16753 gnd.n5809 gnd.n2817 19.3944
R16754 gnd.n5493 gnd.n2817 19.3944
R16755 gnd.n5493 gnd.n5486 19.3944
R16756 gnd.n5505 gnd.n5486 19.3944
R16757 gnd.n5506 gnd.n5505 19.3944
R16758 gnd.n5508 gnd.n5506 19.3944
R16759 gnd.n5509 gnd.n5508 19.3944
R16760 gnd.n5512 gnd.n5509 19.3944
R16761 gnd.n5513 gnd.n5512 19.3944
R16762 gnd.n5518 gnd.n5513 19.3944
R16763 gnd.n5519 gnd.n5518 19.3944
R16764 gnd.n5523 gnd.n5519 19.3944
R16765 gnd.n5523 gnd.n5522 19.3944
R16766 gnd.n5522 gnd.n5521 19.3944
R16767 gnd.n5521 gnd.n5439 19.3944
R16768 gnd.n5582 gnd.n5439 19.3944
R16769 gnd.n5583 gnd.n5582 19.3944
R16770 gnd.n5584 gnd.n5583 19.3944
R16771 gnd.n5584 gnd.n5438 19.3944
R16772 gnd.n5592 gnd.n5438 19.3944
R16773 gnd.n5593 gnd.n5592 19.3944
R16774 gnd.n5601 gnd.n5593 19.3944
R16775 gnd.n5602 gnd.n5601 19.3944
R16776 gnd.n5603 gnd.n5602 19.3944
R16777 gnd.n5612 gnd.n5603 19.3944
R16778 gnd.n5613 gnd.n5612 19.3944
R16779 gnd.n5614 gnd.n5613 19.3944
R16780 gnd.n5615 gnd.n5614 19.3944
R16781 gnd.n5711 gnd.n5615 19.3944
R16782 gnd.n5711 gnd.n5710 19.3944
R16783 gnd.n5710 gnd.n5709 19.3944
R16784 gnd.n5709 gnd.n5617 19.3944
R16785 gnd.n5699 gnd.n5617 19.3944
R16786 gnd.n5699 gnd.n5698 19.3944
R16787 gnd.n5698 gnd.n5697 19.3944
R16788 gnd.n5697 gnd.n5624 19.3944
R16789 gnd.n5640 gnd.n5624 19.3944
R16790 gnd.n5640 gnd.n5639 19.3944
R16791 gnd.n5639 gnd.n5638 19.3944
R16792 gnd.n5638 gnd.n174 19.3944
R16793 gnd.n7341 gnd.n174 19.3944
R16794 gnd.n7342 gnd.n7341 19.3944
R16795 gnd.n5319 gnd.n2815 19.3944
R16796 gnd.n5335 gnd.n5319 19.3944
R16797 gnd.n5796 gnd.n5335 19.3944
R16798 gnd.n5796 gnd.n5795 19.3944
R16799 gnd.n5795 gnd.n5794 19.3944
R16800 gnd.n5794 gnd.n5339 19.3944
R16801 gnd.n5784 gnd.n5339 19.3944
R16802 gnd.n5784 gnd.n5783 19.3944
R16803 gnd.n5783 gnd.n5782 19.3944
R16804 gnd.n5782 gnd.n5359 19.3944
R16805 gnd.n5772 gnd.n5359 19.3944
R16806 gnd.n5772 gnd.n5771 19.3944
R16807 gnd.n5771 gnd.n5770 19.3944
R16808 gnd.n5770 gnd.n5379 19.3944
R16809 gnd.n5760 gnd.n5379 19.3944
R16810 gnd.n5760 gnd.n5759 19.3944
R16811 gnd.n5759 gnd.n5758 19.3944
R16812 gnd.n5758 gnd.n5398 19.3944
R16813 gnd.n5587 gnd.n5398 19.3944
R16814 gnd.n5587 gnd.n5420 19.3944
R16815 gnd.n5734 gnd.n5420 19.3944
R16816 gnd.n5734 gnd.n5733 19.3944
R16817 gnd.n5733 gnd.n5732 19.3944
R16818 gnd.n5732 gnd.n5731 19.3944
R16819 gnd.n5731 gnd.n91 19.3944
R16820 gnd.n7392 gnd.n91 19.3944
R16821 gnd.n7392 gnd.n7391 19.3944
R16822 gnd.n7391 gnd.n7390 19.3944
R16823 gnd.n7390 gnd.n95 19.3944
R16824 gnd.n7380 gnd.n95 19.3944
R16825 gnd.n7380 gnd.n7379 19.3944
R16826 gnd.n7379 gnd.n7378 19.3944
R16827 gnd.n7378 gnd.n114 19.3944
R16828 gnd.n7368 gnd.n114 19.3944
R16829 gnd.n7368 gnd.n7367 19.3944
R16830 gnd.n7367 gnd.n7366 19.3944
R16831 gnd.n7366 gnd.n135 19.3944
R16832 gnd.n7356 gnd.n135 19.3944
R16833 gnd.n7356 gnd.n7355 19.3944
R16834 gnd.n7355 gnd.n7354 19.3944
R16835 gnd.n7354 gnd.n155 19.3944
R16836 gnd.n7344 gnd.n155 19.3944
R16837 gnd.n7251 gnd.n7187 19.3944
R16838 gnd.n7251 gnd.n7248 19.3944
R16839 gnd.n7248 gnd.n7245 19.3944
R16840 gnd.n7245 gnd.n7244 19.3944
R16841 gnd.n7244 gnd.n7241 19.3944
R16842 gnd.n7241 gnd.n7240 19.3944
R16843 gnd.n7240 gnd.n7237 19.3944
R16844 gnd.n7237 gnd.n7236 19.3944
R16845 gnd.n7236 gnd.n7233 19.3944
R16846 gnd.n7233 gnd.n7232 19.3944
R16847 gnd.n7232 gnd.n7229 19.3944
R16848 gnd.n7229 gnd.n7228 19.3944
R16849 gnd.n7228 gnd.n7225 19.3944
R16850 gnd.n7225 gnd.n7224 19.3944
R16851 gnd.n7224 gnd.n7221 19.3944
R16852 gnd.n7221 gnd.n7220 19.3944
R16853 gnd.n7220 gnd.n7217 19.3944
R16854 gnd.n7217 gnd.n7216 19.3944
R16855 gnd.n7294 gnd.n7291 19.3944
R16856 gnd.n7291 gnd.n7290 19.3944
R16857 gnd.n7290 gnd.n7287 19.3944
R16858 gnd.n7287 gnd.n7286 19.3944
R16859 gnd.n7286 gnd.n7283 19.3944
R16860 gnd.n7283 gnd.n7282 19.3944
R16861 gnd.n7282 gnd.n7279 19.3944
R16862 gnd.n7279 gnd.n7278 19.3944
R16863 gnd.n7278 gnd.n7275 19.3944
R16864 gnd.n7275 gnd.n7274 19.3944
R16865 gnd.n7274 gnd.n7271 19.3944
R16866 gnd.n7271 gnd.n7270 19.3944
R16867 gnd.n7270 gnd.n7267 19.3944
R16868 gnd.n7267 gnd.n7266 19.3944
R16869 gnd.n7266 gnd.n7263 19.3944
R16870 gnd.n7263 gnd.n7262 19.3944
R16871 gnd.n7262 gnd.n7259 19.3944
R16872 gnd.n7259 gnd.n7258 19.3944
R16873 gnd.n7149 gnd.n7148 19.3944
R16874 gnd.n7327 gnd.n7148 19.3944
R16875 gnd.n7327 gnd.n7326 19.3944
R16876 gnd.n7326 gnd.n7325 19.3944
R16877 gnd.n7325 gnd.n7322 19.3944
R16878 gnd.n7322 gnd.n7321 19.3944
R16879 gnd.n7321 gnd.n7318 19.3944
R16880 gnd.n7318 gnd.n7317 19.3944
R16881 gnd.n7317 gnd.n7314 19.3944
R16882 gnd.n7314 gnd.n7313 19.3944
R16883 gnd.n7313 gnd.n7310 19.3944
R16884 gnd.n7310 gnd.n7309 19.3944
R16885 gnd.n7309 gnd.n7306 19.3944
R16886 gnd.n7306 gnd.n7305 19.3944
R16887 gnd.n7305 gnd.n7302 19.3944
R16888 gnd.n7302 gnd.n7301 19.3944
R16889 gnd.n7301 gnd.n7298 19.3944
R16890 gnd.n202 gnd.n200 19.3944
R16891 gnd.n205 gnd.n202 19.3944
R16892 gnd.n205 gnd.n197 19.3944
R16893 gnd.n209 gnd.n197 19.3944
R16894 gnd.n212 gnd.n209 19.3944
R16895 gnd.n215 gnd.n212 19.3944
R16896 gnd.n215 gnd.n195 19.3944
R16897 gnd.n219 gnd.n195 19.3944
R16898 gnd.n222 gnd.n219 19.3944
R16899 gnd.n225 gnd.n222 19.3944
R16900 gnd.n225 gnd.n193 19.3944
R16901 gnd.n229 gnd.n193 19.3944
R16902 gnd.n232 gnd.n229 19.3944
R16903 gnd.n234 gnd.n232 19.3944
R16904 gnd.n234 gnd.n191 19.3944
R16905 gnd.n238 gnd.n191 19.3944
R16906 gnd.n5491 gnd.n5490 19.3944
R16907 gnd.n5497 gnd.n5491 19.3944
R16908 gnd.n5497 gnd.n5487 19.3944
R16909 gnd.n5501 gnd.n5487 19.3944
R16910 gnd.n5501 gnd.n5479 19.3944
R16911 gnd.n5537 gnd.n5479 19.3944
R16912 gnd.n5537 gnd.n5480 19.3944
R16913 gnd.n5533 gnd.n5480 19.3944
R16914 gnd.n5533 gnd.n5532 19.3944
R16915 gnd.n5532 gnd.n5531 19.3944
R16916 gnd.n5531 gnd.n5485 19.3944
R16917 gnd.n5527 gnd.n5485 19.3944
R16918 gnd.n5527 gnd.n5443 19.3944
R16919 gnd.n5566 gnd.n5443 19.3944
R16920 gnd.n5566 gnd.n5440 19.3944
R16921 gnd.n5578 gnd.n5440 19.3944
R16922 gnd.n5578 gnd.n5441 19.3944
R16923 gnd.n5574 gnd.n5441 19.3944
R16924 gnd.n5574 gnd.n5573 19.3944
R16925 gnd.n5573 gnd.n5572 19.3944
R16926 gnd.n5572 gnd.n64 19.3944
R16927 gnd.n7405 gnd.n64 19.3944
R16928 gnd.n7405 gnd.n7404 19.3944
R16929 gnd.n7404 gnd.n67 19.3944
R16930 gnd.n5608 gnd.n67 19.3944
R16931 gnd.n5608 gnd.n5433 19.3944
R16932 gnd.n5717 gnd.n5433 19.3944
R16933 gnd.n5717 gnd.n5716 19.3944
R16934 gnd.n5716 gnd.n5715 19.3944
R16935 gnd.n5715 gnd.n5437 19.3944
R16936 gnd.n5705 gnd.n5437 19.3944
R16937 gnd.n5705 gnd.n5704 19.3944
R16938 gnd.n5704 gnd.n5703 19.3944
R16939 gnd.n5703 gnd.n5622 19.3944
R16940 gnd.n5646 gnd.n5622 19.3944
R16941 gnd.n5646 gnd.n5645 19.3944
R16942 gnd.n5645 gnd.n5644 19.3944
R16943 gnd.n5644 gnd.n5629 19.3944
R16944 gnd.n5634 gnd.n5629 19.3944
R16945 gnd.n5634 gnd.n175 19.3944
R16946 gnd.n7337 gnd.n175 19.3944
R16947 gnd.n7337 gnd.n7336 19.3944
R16948 gnd.n5802 gnd.n5323 19.3944
R16949 gnd.n5802 gnd.n5801 19.3944
R16950 gnd.n5801 gnd.n5800 19.3944
R16951 gnd.n5800 gnd.n5328 19.3944
R16952 gnd.n5790 gnd.n5328 19.3944
R16953 gnd.n5790 gnd.n5789 19.3944
R16954 gnd.n5789 gnd.n5788 19.3944
R16955 gnd.n5788 gnd.n5350 19.3944
R16956 gnd.n5778 gnd.n5350 19.3944
R16957 gnd.n5778 gnd.n5777 19.3944
R16958 gnd.n5777 gnd.n5776 19.3944
R16959 gnd.n5776 gnd.n5369 19.3944
R16960 gnd.n5766 gnd.n5369 19.3944
R16961 gnd.n5766 gnd.n5765 19.3944
R16962 gnd.n5765 gnd.n5764 19.3944
R16963 gnd.n5764 gnd.n5389 19.3944
R16964 gnd.n5754 gnd.n5753 19.3944
R16965 gnd.n5737 gnd.n5736 19.3944
R16966 gnd.n5740 gnd.n5739 19.3944
R16967 gnd.n7400 gnd.n7399 19.3944
R16968 gnd.n7396 gnd.n75 19.3944
R16969 gnd.n7396 gnd.n82 19.3944
R16970 gnd.n7386 gnd.n82 19.3944
R16971 gnd.n7386 gnd.n7385 19.3944
R16972 gnd.n7385 gnd.n7384 19.3944
R16973 gnd.n7384 gnd.n104 19.3944
R16974 gnd.n7374 gnd.n104 19.3944
R16975 gnd.n7374 gnd.n7373 19.3944
R16976 gnd.n7373 gnd.n7372 19.3944
R16977 gnd.n7372 gnd.n125 19.3944
R16978 gnd.n7362 gnd.n125 19.3944
R16979 gnd.n7362 gnd.n7361 19.3944
R16980 gnd.n7361 gnd.n7360 19.3944
R16981 gnd.n7360 gnd.n145 19.3944
R16982 gnd.n7350 gnd.n145 19.3944
R16983 gnd.n7350 gnd.n7349 19.3944
R16984 gnd.n7349 gnd.n7348 19.3944
R16985 gnd.n6228 gnd.n2307 19.3944
R16986 gnd.n6228 gnd.n6227 19.3944
R16987 gnd.n6227 gnd.n6226 19.3944
R16988 gnd.n6226 gnd.n2312 19.3944
R16989 gnd.n6220 gnd.n2312 19.3944
R16990 gnd.n6220 gnd.n6219 19.3944
R16991 gnd.n6219 gnd.n6218 19.3944
R16992 gnd.n6218 gnd.n2320 19.3944
R16993 gnd.n3737 gnd.n2320 19.3944
R16994 gnd.n3741 gnd.n3737 19.3944
R16995 gnd.n3741 gnd.n3735 19.3944
R16996 gnd.n3745 gnd.n3735 19.3944
R16997 gnd.n3745 gnd.n3733 19.3944
R16998 gnd.n3810 gnd.n3733 19.3944
R16999 gnd.n3810 gnd.n3809 19.3944
R17000 gnd.n3809 gnd.n3808 19.3944
R17001 gnd.n3808 gnd.n3751 19.3944
R17002 gnd.n3804 gnd.n3751 19.3944
R17003 gnd.n3804 gnd.n3803 19.3944
R17004 gnd.n3803 gnd.n3802 19.3944
R17005 gnd.n3802 gnd.n3757 19.3944
R17006 gnd.n3798 gnd.n3757 19.3944
R17007 gnd.n3798 gnd.n3797 19.3944
R17008 gnd.n3797 gnd.n3796 19.3944
R17009 gnd.n3792 gnd.n3763 19.3944
R17010 gnd.n3788 gnd.n3768 19.3944
R17011 gnd.n3786 gnd.n3785 19.3944
R17012 gnd.n3782 gnd.n3781 19.3944
R17013 gnd.n3778 gnd.n3777 19.3944
R17014 gnd.n3777 gnd.n3776 19.3944
R17015 gnd.n3776 gnd.n3773 19.3944
R17016 gnd.n3773 gnd.n3687 19.3944
R17017 gnd.n4248 gnd.n3687 19.3944
R17018 gnd.n4248 gnd.n3685 19.3944
R17019 gnd.n4252 gnd.n3685 19.3944
R17020 gnd.n4252 gnd.n3683 19.3944
R17021 gnd.n4256 gnd.n3683 19.3944
R17022 gnd.n4256 gnd.n3681 19.3944
R17023 gnd.n4260 gnd.n3681 19.3944
R17024 gnd.n4260 gnd.n3679 19.3944
R17025 gnd.n4264 gnd.n3679 19.3944
R17026 gnd.n4264 gnd.n3677 19.3944
R17027 gnd.n4268 gnd.n3677 19.3944
R17028 gnd.n4268 gnd.n3675 19.3944
R17029 gnd.n4272 gnd.n3675 19.3944
R17030 gnd.n4272 gnd.n3673 19.3944
R17031 gnd.n4277 gnd.n3673 19.3944
R17032 gnd.n4277 gnd.n2567 19.3944
R17033 gnd.n6067 gnd.n2567 19.3944
R17034 gnd.n6067 gnd.n6066 19.3944
R17035 gnd.n6066 gnd.n6065 19.3944
R17036 gnd.n6065 gnd.n2571 19.3944
R17037 gnd.n3452 gnd.n2571 19.3944
R17038 gnd.n3456 gnd.n3452 19.3944
R17039 gnd.n3456 gnd.n3447 19.3944
R17040 gnd.n3464 gnd.n3447 19.3944
R17041 gnd.n3464 gnd.n3445 19.3944
R17042 gnd.n3468 gnd.n3445 19.3944
R17043 gnd.n3468 gnd.n3441 19.3944
R17044 gnd.n3476 gnd.n3441 19.3944
R17045 gnd.n3476 gnd.n3439 19.3944
R17046 gnd.n3482 gnd.n3439 19.3944
R17047 gnd.n3482 gnd.n3481 19.3944
R17048 gnd.n3481 gnd.n3220 19.3944
R17049 gnd.n4558 gnd.n3220 19.3944
R17050 gnd.n4558 gnd.n3218 19.3944
R17051 gnd.n4564 gnd.n3218 19.3944
R17052 gnd.n4564 gnd.n4563 19.3944
R17053 gnd.n4563 gnd.n3196 19.3944
R17054 gnd.n4596 gnd.n3196 19.3944
R17055 gnd.n4596 gnd.n3194 19.3944
R17056 gnd.n4605 gnd.n3194 19.3944
R17057 gnd.n4605 gnd.n4604 19.3944
R17058 gnd.n4604 gnd.n4603 19.3944
R17059 gnd.n4603 gnd.n3171 19.3944
R17060 gnd.n4636 gnd.n3171 19.3944
R17061 gnd.n4636 gnd.n3169 19.3944
R17062 gnd.n4642 gnd.n3169 19.3944
R17063 gnd.n4642 gnd.n4641 19.3944
R17064 gnd.n4641 gnd.n3143 19.3944
R17065 gnd.n4672 gnd.n3143 19.3944
R17066 gnd.n4672 gnd.n3141 19.3944
R17067 gnd.n4676 gnd.n3141 19.3944
R17068 gnd.n4676 gnd.n3125 19.3944
R17069 gnd.n4698 gnd.n3125 19.3944
R17070 gnd.n4698 gnd.n3123 19.3944
R17071 gnd.n4704 gnd.n3123 19.3944
R17072 gnd.n4704 gnd.n4703 19.3944
R17073 gnd.n4703 gnd.n3099 19.3944
R17074 gnd.n4754 gnd.n3099 19.3944
R17075 gnd.n4754 gnd.n3097 19.3944
R17076 gnd.n4760 gnd.n3097 19.3944
R17077 gnd.n4760 gnd.n4759 19.3944
R17078 gnd.n4759 gnd.n3074 19.3944
R17079 gnd.n4794 gnd.n3074 19.3944
R17080 gnd.n4794 gnd.n3072 19.3944
R17081 gnd.n4800 gnd.n3072 19.3944
R17082 gnd.n4800 gnd.n4799 19.3944
R17083 gnd.n4799 gnd.n3044 19.3944
R17084 gnd.n4863 gnd.n3044 19.3944
R17085 gnd.n4863 gnd.n3042 19.3944
R17086 gnd.n4869 gnd.n3042 19.3944
R17087 gnd.n4869 gnd.n4868 19.3944
R17088 gnd.n4868 gnd.n3020 19.3944
R17089 gnd.n4896 gnd.n3020 19.3944
R17090 gnd.n4896 gnd.n3018 19.3944
R17091 gnd.n4902 gnd.n3018 19.3944
R17092 gnd.n4902 gnd.n4901 19.3944
R17093 gnd.n4901 gnd.n2999 19.3944
R17094 gnd.n4950 gnd.n2999 19.3944
R17095 gnd.n4950 gnd.n2997 19.3944
R17096 gnd.n4956 gnd.n2997 19.3944
R17097 gnd.n4956 gnd.n4955 19.3944
R17098 gnd.n4955 gnd.n2974 19.3944
R17099 gnd.n4987 gnd.n2974 19.3944
R17100 gnd.n4987 gnd.n2972 19.3944
R17101 gnd.n4991 gnd.n2972 19.3944
R17102 gnd.n4991 gnd.n2883 19.3944
R17103 gnd.n5130 gnd.n2883 19.3944
R17104 gnd.n5130 gnd.n2881 19.3944
R17105 gnd.n5134 gnd.n2881 19.3944
R17106 gnd.n5134 gnd.n2870 19.3944
R17107 gnd.n5146 gnd.n2870 19.3944
R17108 gnd.n5146 gnd.n2868 19.3944
R17109 gnd.n5150 gnd.n2868 19.3944
R17110 gnd.n5150 gnd.n2857 19.3944
R17111 gnd.n5162 gnd.n2857 19.3944
R17112 gnd.n5162 gnd.n2855 19.3944
R17113 gnd.n5166 gnd.n2855 19.3944
R17114 gnd.n5166 gnd.n2843 19.3944
R17115 gnd.n5179 gnd.n2843 19.3944
R17116 gnd.n5179 gnd.n2841 19.3944
R17117 gnd.n5184 gnd.n2841 19.3944
R17118 gnd.n5184 gnd.n2701 19.3944
R17119 gnd.n5932 gnd.n2701 19.3944
R17120 gnd.n5932 gnd.n5931 19.3944
R17121 gnd.n5931 gnd.n5930 19.3944
R17122 gnd.n5930 gnd.n2705 19.3944
R17123 gnd.n5462 gnd.n2705 19.3944
R17124 gnd.n5465 gnd.n5462 19.3944
R17125 gnd.n5465 gnd.n5459 19.3944
R17126 gnd.n5469 gnd.n5459 19.3944
R17127 gnd.n5469 gnd.n5457 19.3944
R17128 gnd.n5473 gnd.n5457 19.3944
R17129 gnd.n5473 gnd.n5455 19.3944
R17130 gnd.n5477 gnd.n5455 19.3944
R17131 gnd.n5477 gnd.n5453 19.3944
R17132 gnd.n5544 gnd.n5453 19.3944
R17133 gnd.n5544 gnd.n5451 19.3944
R17134 gnd.n5548 gnd.n5451 19.3944
R17135 gnd.n5548 gnd.n5449 19.3944
R17136 gnd.n5552 gnd.n5449 19.3944
R17137 gnd.n5552 gnd.n5447 19.3944
R17138 gnd.n5561 gnd.n5447 19.3944
R17139 gnd.n5561 gnd.n5560 19.3944
R17140 gnd.n5560 gnd.n5559 19.3944
R17141 gnd.n5748 gnd.n5410 19.3944
R17142 gnd.n5746 gnd.n5745 19.3944
R17143 gnd.n5596 gnd.n5594 19.3944
R17144 gnd.n5726 gnd.n5428 19.3944
R17145 gnd.n5724 gnd.n5723 19.3944
R17146 gnd.n5723 gnd.n5430 19.3944
R17147 gnd.n5657 gnd.n5430 19.3944
R17148 gnd.n5659 gnd.n5657 19.3944
R17149 gnd.n5659 gnd.n5654 19.3944
R17150 gnd.n5663 gnd.n5654 19.3944
R17151 gnd.n5663 gnd.n5652 19.3944
R17152 gnd.n5667 gnd.n5652 19.3944
R17153 gnd.n5667 gnd.n5650 19.3944
R17154 gnd.n5692 gnd.n5650 19.3944
R17155 gnd.n5692 gnd.n5691 19.3944
R17156 gnd.n5691 gnd.n5690 19.3944
R17157 gnd.n5690 gnd.n5673 19.3944
R17158 gnd.n5686 gnd.n5673 19.3944
R17159 gnd.n5686 gnd.n5685 19.3944
R17160 gnd.n5685 gnd.n5684 19.3944
R17161 gnd.n5684 gnd.n5681 19.3944
R17162 gnd.n5681 gnd.n244 19.3944
R17163 gnd.n7115 gnd.n244 19.3944
R17164 gnd.n7115 gnd.n7114 19.3944
R17165 gnd.n7114 gnd.n7113 19.3944
R17166 gnd.n7113 gnd.n248 19.3944
R17167 gnd.n7107 gnd.n248 19.3944
R17168 gnd.n7107 gnd.n7106 19.3944
R17169 gnd.n3960 gnd.n3957 19.3944
R17170 gnd.n3960 gnd.n3955 19.3944
R17171 gnd.n3964 gnd.n3955 19.3944
R17172 gnd.n3964 gnd.n3953 19.3944
R17173 gnd.n3970 gnd.n3953 19.3944
R17174 gnd.n3970 gnd.n3951 19.3944
R17175 gnd.n3974 gnd.n3951 19.3944
R17176 gnd.n3974 gnd.n3949 19.3944
R17177 gnd.n3980 gnd.n3949 19.3944
R17178 gnd.n3980 gnd.n3947 19.3944
R17179 gnd.n3984 gnd.n3947 19.3944
R17180 gnd.n3984 gnd.n3945 19.3944
R17181 gnd.n3990 gnd.n3945 19.3944
R17182 gnd.n3990 gnd.n3943 19.3944
R17183 gnd.n3994 gnd.n3943 19.3944
R17184 gnd.n3994 gnd.n3938 19.3944
R17185 gnd.n4000 gnd.n3938 19.3944
R17186 gnd.n4004 gnd.n3936 19.3944
R17187 gnd.n4004 gnd.n3934 19.3944
R17188 gnd.n4010 gnd.n3934 19.3944
R17189 gnd.n4010 gnd.n3932 19.3944
R17190 gnd.n4014 gnd.n3932 19.3944
R17191 gnd.n4014 gnd.n3930 19.3944
R17192 gnd.n4020 gnd.n3930 19.3944
R17193 gnd.n4020 gnd.n3928 19.3944
R17194 gnd.n4024 gnd.n3928 19.3944
R17195 gnd.n4024 gnd.n3926 19.3944
R17196 gnd.n4030 gnd.n3926 19.3944
R17197 gnd.n4030 gnd.n3924 19.3944
R17198 gnd.n4034 gnd.n3924 19.3944
R17199 gnd.n4034 gnd.n3922 19.3944
R17200 gnd.n4040 gnd.n3922 19.3944
R17201 gnd.n4040 gnd.n3920 19.3944
R17202 gnd.n4044 gnd.n3920 19.3944
R17203 gnd.n4044 gnd.n3918 19.3944
R17204 gnd.n4056 gnd.n3916 19.3944
R17205 gnd.n4056 gnd.n3914 19.3944
R17206 gnd.n4062 gnd.n3914 19.3944
R17207 gnd.n4062 gnd.n3912 19.3944
R17208 gnd.n4066 gnd.n3912 19.3944
R17209 gnd.n4066 gnd.n3910 19.3944
R17210 gnd.n4072 gnd.n3910 19.3944
R17211 gnd.n4072 gnd.n3908 19.3944
R17212 gnd.n4076 gnd.n3908 19.3944
R17213 gnd.n4076 gnd.n3906 19.3944
R17214 gnd.n4082 gnd.n3906 19.3944
R17215 gnd.n4082 gnd.n3904 19.3944
R17216 gnd.n4086 gnd.n3904 19.3944
R17217 gnd.n4086 gnd.n3902 19.3944
R17218 gnd.n4092 gnd.n3902 19.3944
R17219 gnd.n4092 gnd.n3900 19.3944
R17220 gnd.n4097 gnd.n3900 19.3944
R17221 gnd.n4097 gnd.n3898 19.3944
R17222 gnd.n3892 gnd.n3821 19.3944
R17223 gnd.n3887 gnd.n3821 19.3944
R17224 gnd.n3887 gnd.n3886 19.3944
R17225 gnd.n3886 gnd.n3825 19.3944
R17226 gnd.n3881 gnd.n3825 19.3944
R17227 gnd.n3881 gnd.n3880 19.3944
R17228 gnd.n3880 gnd.n3879 19.3944
R17229 gnd.n3879 gnd.n3831 19.3944
R17230 gnd.n3873 gnd.n3831 19.3944
R17231 gnd.n3873 gnd.n3872 19.3944
R17232 gnd.n3872 gnd.n3871 19.3944
R17233 gnd.n3871 gnd.n3837 19.3944
R17234 gnd.n3865 gnd.n3837 19.3944
R17235 gnd.n3865 gnd.n3864 19.3944
R17236 gnd.n3864 gnd.n3863 19.3944
R17237 gnd.n3863 gnd.n3843 19.3944
R17238 gnd.n3851 gnd.n3850 19.3944
R17239 gnd.n3850 gnd.n3817 19.3944
R17240 gnd.n4116 gnd.n3817 19.3944
R17241 gnd.n4116 gnd.n3815 19.3944
R17242 gnd.n4120 gnd.n3815 19.3944
R17243 gnd.n4120 gnd.n3730 19.3944
R17244 gnd.n4130 gnd.n3730 19.3944
R17245 gnd.n4130 gnd.n3728 19.3944
R17246 gnd.n4134 gnd.n3728 19.3944
R17247 gnd.n4134 gnd.n3725 19.3944
R17248 gnd.n4144 gnd.n3725 19.3944
R17249 gnd.n4144 gnd.n3723 19.3944
R17250 gnd.n4148 gnd.n3723 19.3944
R17251 gnd.n4148 gnd.n3719 19.3944
R17252 gnd.n4158 gnd.n3719 19.3944
R17253 gnd.n4158 gnd.n3717 19.3944
R17254 gnd.n4162 gnd.n3717 19.3944
R17255 gnd.n4162 gnd.n3714 19.3944
R17256 gnd.n4172 gnd.n3714 19.3944
R17257 gnd.n4172 gnd.n3712 19.3944
R17258 gnd.n4176 gnd.n3712 19.3944
R17259 gnd.n4176 gnd.n3708 19.3944
R17260 gnd.n4186 gnd.n3708 19.3944
R17261 gnd.n4186 gnd.n3706 19.3944
R17262 gnd.n4190 gnd.n3706 19.3944
R17263 gnd.n4190 gnd.n3703 19.3944
R17264 gnd.n4200 gnd.n3703 19.3944
R17265 gnd.n4200 gnd.n3701 19.3944
R17266 gnd.n4204 gnd.n3701 19.3944
R17267 gnd.n4204 gnd.n3690 19.3944
R17268 gnd.n4243 gnd.n3690 19.3944
R17269 gnd.n4243 gnd.n3691 19.3944
R17270 gnd.n4239 gnd.n3691 19.3944
R17271 gnd.n4239 gnd.n4238 19.3944
R17272 gnd.n4238 gnd.n4237 19.3944
R17273 gnd.n4237 gnd.n3696 19.3944
R17274 gnd.n4233 gnd.n3696 19.3944
R17275 gnd.n4233 gnd.n4232 19.3944
R17276 gnd.n4232 gnd.n4231 19.3944
R17277 gnd.n4231 gnd.n2541 19.3944
R17278 gnd.n6077 gnd.n2541 19.3944
R17279 gnd.n6077 gnd.n2542 19.3944
R17280 gnd.n4110 gnd.n3818 19.3944
R17281 gnd.n4111 gnd.n4110 19.3944
R17282 gnd.n4112 gnd.n4111 19.3944
R17283 gnd.n4112 gnd.n3813 19.3944
R17284 gnd.n4124 gnd.n3813 19.3944
R17285 gnd.n4125 gnd.n4124 19.3944
R17286 gnd.n4126 gnd.n4125 19.3944
R17287 gnd.n4126 gnd.n3726 19.3944
R17288 gnd.n4138 gnd.n3726 19.3944
R17289 gnd.n4139 gnd.n4138 19.3944
R17290 gnd.n4140 gnd.n4139 19.3944
R17291 gnd.n4140 gnd.n3721 19.3944
R17292 gnd.n4152 gnd.n3721 19.3944
R17293 gnd.n4153 gnd.n4152 19.3944
R17294 gnd.n4154 gnd.n4153 19.3944
R17295 gnd.n4154 gnd.n3715 19.3944
R17296 gnd.n4166 gnd.n3715 19.3944
R17297 gnd.n4167 gnd.n4166 19.3944
R17298 gnd.n4168 gnd.n4167 19.3944
R17299 gnd.n4168 gnd.n3710 19.3944
R17300 gnd.n4180 gnd.n3710 19.3944
R17301 gnd.n4181 gnd.n4180 19.3944
R17302 gnd.n4182 gnd.n4181 19.3944
R17303 gnd.n4182 gnd.n3704 19.3944
R17304 gnd.n4194 gnd.n3704 19.3944
R17305 gnd.n4195 gnd.n4194 19.3944
R17306 gnd.n4196 gnd.n4195 19.3944
R17307 gnd.n4196 gnd.n3699 19.3944
R17308 gnd.n4208 gnd.n3699 19.3944
R17309 gnd.n4209 gnd.n4208 19.3944
R17310 gnd.n4210 gnd.n4209 19.3944
R17311 gnd.n4211 gnd.n4210 19.3944
R17312 gnd.n4215 gnd.n4211 19.3944
R17313 gnd.n4216 gnd.n4215 19.3944
R17314 gnd.n4219 gnd.n4216 19.3944
R17315 gnd.n4220 gnd.n4219 19.3944
R17316 gnd.n4224 gnd.n4220 19.3944
R17317 gnd.n4225 gnd.n4224 19.3944
R17318 gnd.n4226 gnd.n4225 19.3944
R17319 gnd.n4226 gnd.n2539 19.3944
R17320 gnd.n6081 gnd.n2539 19.3944
R17321 gnd.n6082 gnd.n6081 19.3944
R17322 gnd.n4107 gnd.n2340 19.3944
R17323 gnd.n6207 gnd.n2340 19.3944
R17324 gnd.n6207 gnd.n6206 19.3944
R17325 gnd.n6206 gnd.n6205 19.3944
R17326 gnd.n6205 gnd.n2344 19.3944
R17327 gnd.n6195 gnd.n2344 19.3944
R17328 gnd.n6195 gnd.n6194 19.3944
R17329 gnd.n6194 gnd.n6193 19.3944
R17330 gnd.n6193 gnd.n2364 19.3944
R17331 gnd.n6183 gnd.n2364 19.3944
R17332 gnd.n6183 gnd.n6182 19.3944
R17333 gnd.n6182 gnd.n6181 19.3944
R17334 gnd.n6181 gnd.n2385 19.3944
R17335 gnd.n6171 gnd.n2385 19.3944
R17336 gnd.n6171 gnd.n6170 19.3944
R17337 gnd.n6170 gnd.n6169 19.3944
R17338 gnd.n6169 gnd.n2405 19.3944
R17339 gnd.n6158 gnd.n2405 19.3944
R17340 gnd.n6158 gnd.n6157 19.3944
R17341 gnd.n6157 gnd.n6156 19.3944
R17342 gnd.n6156 gnd.n2424 19.3944
R17343 gnd.n6145 gnd.n2424 19.3944
R17344 gnd.n6145 gnd.n6144 19.3944
R17345 gnd.n6144 gnd.n6143 19.3944
R17346 gnd.n6143 gnd.n2441 19.3944
R17347 gnd.n6132 gnd.n2441 19.3944
R17348 gnd.n6132 gnd.n6131 19.3944
R17349 gnd.n6131 gnd.n6130 19.3944
R17350 gnd.n6130 gnd.n2459 19.3944
R17351 gnd.n6120 gnd.n2459 19.3944
R17352 gnd.n6120 gnd.n6119 19.3944
R17353 gnd.n6119 gnd.n6118 19.3944
R17354 gnd.n6118 gnd.n2479 19.3944
R17355 gnd.n6108 gnd.n2479 19.3944
R17356 gnd.n6108 gnd.n6107 19.3944
R17357 gnd.n6107 gnd.n6106 19.3944
R17358 gnd.n6106 gnd.n2500 19.3944
R17359 gnd.n6096 gnd.n2500 19.3944
R17360 gnd.n6096 gnd.n6095 19.3944
R17361 gnd.n6095 gnd.n6094 19.3944
R17362 gnd.n6094 gnd.n2521 19.3944
R17363 gnd.n6084 gnd.n2521 19.3944
R17364 gnd.n4296 gnd.n4295 19.3944
R17365 gnd.n4369 gnd.n4295 19.3944
R17366 gnd.n4369 gnd.n4368 19.3944
R17367 gnd.n4368 gnd.n4367 19.3944
R17368 gnd.n4367 gnd.n4364 19.3944
R17369 gnd.n4364 gnd.n4363 19.3944
R17370 gnd.n4363 gnd.n4360 19.3944
R17371 gnd.n4360 gnd.n4359 19.3944
R17372 gnd.n4359 gnd.n4356 19.3944
R17373 gnd.n4356 gnd.n4355 19.3944
R17374 gnd.n4355 gnd.n4352 19.3944
R17375 gnd.n4352 gnd.n4351 19.3944
R17376 gnd.n4351 gnd.n4348 19.3944
R17377 gnd.n4348 gnd.n4347 19.3944
R17378 gnd.n4347 gnd.n4344 19.3944
R17379 gnd.n4344 gnd.n4343 19.3944
R17380 gnd.n4343 gnd.n4340 19.3944
R17381 gnd.n4459 gnd.n4384 19.3944
R17382 gnd.n4459 gnd.n4388 19.3944
R17383 gnd.n4391 gnd.n4388 19.3944
R17384 gnd.n4452 gnd.n4391 19.3944
R17385 gnd.n4452 gnd.n4451 19.3944
R17386 gnd.n4451 gnd.n4450 19.3944
R17387 gnd.n4450 gnd.n4397 19.3944
R17388 gnd.n4445 gnd.n4397 19.3944
R17389 gnd.n4445 gnd.n4444 19.3944
R17390 gnd.n4444 gnd.n4443 19.3944
R17391 gnd.n4443 gnd.n4404 19.3944
R17392 gnd.n4438 gnd.n4404 19.3944
R17393 gnd.n4438 gnd.n4437 19.3944
R17394 gnd.n4437 gnd.n4436 19.3944
R17395 gnd.n4436 gnd.n4411 19.3944
R17396 gnd.n4431 gnd.n4411 19.3944
R17397 gnd.n4431 gnd.n4430 19.3944
R17398 gnd.n4430 gnd.n4429 19.3944
R17399 gnd.n4478 gnd.n3359 19.3944
R17400 gnd.n4478 gnd.n3364 19.3944
R17401 gnd.n4373 gnd.n3364 19.3944
R17402 gnd.n4471 gnd.n4373 19.3944
R17403 gnd.n4471 gnd.n4470 19.3944
R17404 gnd.n4470 gnd.n4469 19.3944
R17405 gnd.n4469 gnd.n4379 19.3944
R17406 gnd.n4464 gnd.n4379 19.3944
R17407 gnd.n4338 gnd.n4335 19.3944
R17408 gnd.n4335 gnd.n4334 19.3944
R17409 gnd.n4334 gnd.n4331 19.3944
R17410 gnd.n4331 gnd.n4330 19.3944
R17411 gnd.n4330 gnd.n4327 19.3944
R17412 gnd.n4327 gnd.n4326 19.3944
R17413 gnd.n4326 gnd.n3360 19.3944
R17414 gnd.n6213 gnd.n6212 19.3944
R17415 gnd.n6212 gnd.n6211 19.3944
R17416 gnd.n6211 gnd.n2332 19.3944
R17417 gnd.n6201 gnd.n2332 19.3944
R17418 gnd.n6201 gnd.n6200 19.3944
R17419 gnd.n6200 gnd.n6199 19.3944
R17420 gnd.n6199 gnd.n2355 19.3944
R17421 gnd.n6189 gnd.n2355 19.3944
R17422 gnd.n6189 gnd.n6188 19.3944
R17423 gnd.n6188 gnd.n6187 19.3944
R17424 gnd.n6187 gnd.n2375 19.3944
R17425 gnd.n6177 gnd.n2375 19.3944
R17426 gnd.n6177 gnd.n6176 19.3944
R17427 gnd.n6176 gnd.n6175 19.3944
R17428 gnd.n6175 gnd.n2396 19.3944
R17429 gnd.n6165 gnd.n2396 19.3944
R17430 gnd.n6163 gnd.n6162 19.3944
R17431 gnd.n6152 gnd.n2431 19.3944
R17432 gnd.n6150 gnd.n6149 19.3944
R17433 gnd.n6139 gnd.n2448 19.3944
R17434 gnd.n6137 gnd.n6136 19.3944
R17435 gnd.n6136 gnd.n2449 19.3944
R17436 gnd.n6126 gnd.n2449 19.3944
R17437 gnd.n6126 gnd.n6125 19.3944
R17438 gnd.n6125 gnd.n6124 19.3944
R17439 gnd.n6124 gnd.n2470 19.3944
R17440 gnd.n6114 gnd.n2470 19.3944
R17441 gnd.n6114 gnd.n6113 19.3944
R17442 gnd.n6113 gnd.n6112 19.3944
R17443 gnd.n6112 gnd.n2490 19.3944
R17444 gnd.n6102 gnd.n2490 19.3944
R17445 gnd.n6102 gnd.n6101 19.3944
R17446 gnd.n6101 gnd.n6100 19.3944
R17447 gnd.n6100 gnd.n2511 19.3944
R17448 gnd.n6090 gnd.n2511 19.3944
R17449 gnd.n6090 gnd.n6089 19.3944
R17450 gnd.n6089 gnd.n6088 19.3944
R17451 gnd.n6402 gnd.n674 19.3944
R17452 gnd.n6396 gnd.n674 19.3944
R17453 gnd.n6396 gnd.n6395 19.3944
R17454 gnd.n6395 gnd.n6394 19.3944
R17455 gnd.n6394 gnd.n681 19.3944
R17456 gnd.n6388 gnd.n681 19.3944
R17457 gnd.n6388 gnd.n6387 19.3944
R17458 gnd.n6387 gnd.n6386 19.3944
R17459 gnd.n6386 gnd.n689 19.3944
R17460 gnd.n6380 gnd.n689 19.3944
R17461 gnd.n6380 gnd.n6379 19.3944
R17462 gnd.n6379 gnd.n6378 19.3944
R17463 gnd.n6378 gnd.n697 19.3944
R17464 gnd.n6372 gnd.n697 19.3944
R17465 gnd.n6372 gnd.n6371 19.3944
R17466 gnd.n6371 gnd.n6370 19.3944
R17467 gnd.n6370 gnd.n705 19.3944
R17468 gnd.n6364 gnd.n705 19.3944
R17469 gnd.n6364 gnd.n6363 19.3944
R17470 gnd.n6363 gnd.n6362 19.3944
R17471 gnd.n6362 gnd.n713 19.3944
R17472 gnd.n6356 gnd.n713 19.3944
R17473 gnd.n6356 gnd.n6355 19.3944
R17474 gnd.n6355 gnd.n6354 19.3944
R17475 gnd.n6354 gnd.n721 19.3944
R17476 gnd.n6348 gnd.n721 19.3944
R17477 gnd.n6348 gnd.n6347 19.3944
R17478 gnd.n6347 gnd.n6346 19.3944
R17479 gnd.n6346 gnd.n729 19.3944
R17480 gnd.n6340 gnd.n729 19.3944
R17481 gnd.n6340 gnd.n6339 19.3944
R17482 gnd.n6339 gnd.n6338 19.3944
R17483 gnd.n6338 gnd.n737 19.3944
R17484 gnd.n6332 gnd.n737 19.3944
R17485 gnd.n6332 gnd.n6331 19.3944
R17486 gnd.n6331 gnd.n6330 19.3944
R17487 gnd.n6330 gnd.n745 19.3944
R17488 gnd.n6324 gnd.n745 19.3944
R17489 gnd.n6324 gnd.n6323 19.3944
R17490 gnd.n6323 gnd.n6322 19.3944
R17491 gnd.n6322 gnd.n753 19.3944
R17492 gnd.n6316 gnd.n753 19.3944
R17493 gnd.n6316 gnd.n6315 19.3944
R17494 gnd.n6315 gnd.n6314 19.3944
R17495 gnd.n6314 gnd.n761 19.3944
R17496 gnd.n6308 gnd.n761 19.3944
R17497 gnd.n6308 gnd.n6307 19.3944
R17498 gnd.n6307 gnd.n6306 19.3944
R17499 gnd.n6306 gnd.n769 19.3944
R17500 gnd.n6300 gnd.n769 19.3944
R17501 gnd.n6300 gnd.n6299 19.3944
R17502 gnd.n6299 gnd.n6298 19.3944
R17503 gnd.n6298 gnd.n777 19.3944
R17504 gnd.n6292 gnd.n777 19.3944
R17505 gnd.n6292 gnd.n6291 19.3944
R17506 gnd.n6291 gnd.n6290 19.3944
R17507 gnd.n6290 gnd.n785 19.3944
R17508 gnd.n6284 gnd.n785 19.3944
R17509 gnd.n6284 gnd.n6283 19.3944
R17510 gnd.n6283 gnd.n6282 19.3944
R17511 gnd.n6282 gnd.n793 19.3944
R17512 gnd.n6276 gnd.n793 19.3944
R17513 gnd.n6276 gnd.n6275 19.3944
R17514 gnd.n6275 gnd.n6274 19.3944
R17515 gnd.n6274 gnd.n801 19.3944
R17516 gnd.n6268 gnd.n801 19.3944
R17517 gnd.n6268 gnd.n6267 19.3944
R17518 gnd.n6267 gnd.n6266 19.3944
R17519 gnd.n6266 gnd.n809 19.3944
R17520 gnd.n6260 gnd.n809 19.3944
R17521 gnd.n6260 gnd.n6259 19.3944
R17522 gnd.n6259 gnd.n6258 19.3944
R17523 gnd.n6258 gnd.n817 19.3944
R17524 gnd.n6252 gnd.n817 19.3944
R17525 gnd.n6252 gnd.n6251 19.3944
R17526 gnd.n6251 gnd.n6250 19.3944
R17527 gnd.n6250 gnd.n825 19.3944
R17528 gnd.n6244 gnd.n825 19.3944
R17529 gnd.n6244 gnd.n6243 19.3944
R17530 gnd.n6243 gnd.n6242 19.3944
R17531 gnd.n6242 gnd.n833 19.3944
R17532 gnd.n6236 gnd.n833 19.3944
R17533 gnd.n6236 gnd.n6235 19.3944
R17534 gnd.n6235 gnd.n6234 19.3944
R17535 gnd.n3576 gnd.n3575 19.3944
R17536 gnd.n3575 gnd.n3574 19.3944
R17537 gnd.n3574 gnd.n3425 19.3944
R17538 gnd.n3570 gnd.n3425 19.3944
R17539 gnd.n3570 gnd.n3569 19.3944
R17540 gnd.n3569 gnd.n3568 19.3944
R17541 gnd.n3568 gnd.n3430 19.3944
R17542 gnd.n3564 gnd.n3430 19.3944
R17543 gnd.n3564 gnd.n3563 19.3944
R17544 gnd.n3563 gnd.n3562 19.3944
R17545 gnd.n3562 gnd.n3435 19.3944
R17546 gnd.n3558 gnd.n3435 19.3944
R17547 gnd.n3558 gnd.n3557 19.3944
R17548 gnd.n3557 gnd.n3556 19.3944
R17549 gnd.n3556 gnd.n3489 19.3944
R17550 gnd.n3552 gnd.n3489 19.3944
R17551 gnd.n3552 gnd.n3551 19.3944
R17552 gnd.n3551 gnd.n3550 19.3944
R17553 gnd.n3550 gnd.n3496 19.3944
R17554 gnd.n3546 gnd.n3496 19.3944
R17555 gnd.n3546 gnd.n3545 19.3944
R17556 gnd.n3545 gnd.n3544 19.3944
R17557 gnd.n3544 gnd.n3502 19.3944
R17558 gnd.n3540 gnd.n3502 19.3944
R17559 gnd.n3540 gnd.n3539 19.3944
R17560 gnd.n3539 gnd.n3538 19.3944
R17561 gnd.n3538 gnd.n3505 19.3944
R17562 gnd.n3534 gnd.n3505 19.3944
R17563 gnd.n3534 gnd.n3533 19.3944
R17564 gnd.n3533 gnd.n3532 19.3944
R17565 gnd.n3532 gnd.n3510 19.3944
R17566 gnd.n3528 gnd.n3510 19.3944
R17567 gnd.n3528 gnd.n3527 19.3944
R17568 gnd.n3527 gnd.n3526 19.3944
R17569 gnd.n3526 gnd.n3514 19.3944
R17570 gnd.n3522 gnd.n3514 19.3944
R17571 gnd.n3522 gnd.n3521 19.3944
R17572 gnd.n3521 gnd.n3520 19.3944
R17573 gnd.n3520 gnd.n3517 19.3944
R17574 gnd.n3517 gnd.n3089 19.3944
R17575 gnd.n4764 gnd.n3089 19.3944
R17576 gnd.n4764 gnd.n3086 19.3944
R17577 gnd.n4782 gnd.n3086 19.3944
R17578 gnd.n4782 gnd.n3087 19.3944
R17579 gnd.n4778 gnd.n3087 19.3944
R17580 gnd.n4778 gnd.n4777 19.3944
R17581 gnd.n4777 gnd.n4776 19.3944
R17582 gnd.n4776 gnd.n4771 19.3944
R17583 gnd.n4772 gnd.n4771 19.3944
R17584 gnd.n4772 gnd.n3036 19.3944
R17585 gnd.n4873 gnd.n3036 19.3944
R17586 gnd.n4873 gnd.n3033 19.3944
R17587 gnd.n4878 gnd.n3033 19.3944
R17588 gnd.n4878 gnd.n3034 19.3944
R17589 gnd.n3034 gnd.n3013 19.3944
R17590 gnd.n4906 gnd.n3013 19.3944
R17591 gnd.n4906 gnd.n3010 19.3944
R17592 gnd.n4937 gnd.n3010 19.3944
R17593 gnd.n4937 gnd.n3011 19.3944
R17594 gnd.n4933 gnd.n3011 19.3944
R17595 gnd.n4933 gnd.n4932 19.3944
R17596 gnd.n4932 gnd.n4931 19.3944
R17597 gnd.n4931 gnd.n4916 19.3944
R17598 gnd.n4927 gnd.n4916 19.3944
R17599 gnd.n4927 gnd.n4926 19.3944
R17600 gnd.n4926 gnd.n4925 19.3944
R17601 gnd.n4925 gnd.n4920 19.3944
R17602 gnd.n4921 gnd.n4920 19.3944
R17603 gnd.n4921 gnd.n2875 19.3944
R17604 gnd.n5138 gnd.n2875 19.3944
R17605 gnd.n5138 gnd.n2873 19.3944
R17606 gnd.n5142 gnd.n2873 19.3944
R17607 gnd.n5142 gnd.n2862 19.3944
R17608 gnd.n5154 gnd.n2862 19.3944
R17609 gnd.n5154 gnd.n2860 19.3944
R17610 gnd.n5158 gnd.n2860 19.3944
R17611 gnd.n5158 gnd.n2850 19.3944
R17612 gnd.n5170 gnd.n2850 19.3944
R17613 gnd.n5170 gnd.n2847 19.3944
R17614 gnd.n5175 gnd.n2847 19.3944
R17615 gnd.n5175 gnd.n2848 19.3944
R17616 gnd.n2848 gnd.n2838 19.3944
R17617 gnd.n5189 gnd.n2833 19.3944
R17618 gnd.n5193 gnd.n2833 19.3944
R17619 gnd.n5194 gnd.n5193 19.3944
R17620 gnd.n5197 gnd.n5194 19.3944
R17621 gnd.n5197 gnd.n2829 19.3944
R17622 gnd.n5201 gnd.n2829 19.3944
R17623 gnd.n5202 gnd.n5201 19.3944
R17624 gnd.n5207 gnd.n5202 19.3944
R17625 gnd.n5208 gnd.n5207 19.3944
R17626 gnd.n5312 gnd.n5208 19.3944
R17627 gnd.n5312 gnd.n5311 19.3944
R17628 gnd.n5311 gnd.n5213 19.3944
R17629 gnd.n5304 gnd.n5213 19.3944
R17630 gnd.n5304 gnd.n5303 19.3944
R17631 gnd.n5303 gnd.n5221 19.3944
R17632 gnd.n5296 gnd.n5221 19.3944
R17633 gnd.n5296 gnd.n5295 19.3944
R17634 gnd.n5295 gnd.n5233 19.3944
R17635 gnd.n5288 gnd.n5233 19.3944
R17636 gnd.n5288 gnd.n5287 19.3944
R17637 gnd.n5287 gnd.n5241 19.3944
R17638 gnd.n5280 gnd.n5241 19.3944
R17639 gnd.n5280 gnd.n5279 19.3944
R17640 gnd.n5279 gnd.n5253 19.3944
R17641 gnd.n5272 gnd.n5271 19.3944
R17642 gnd.n5271 gnd.n2680 19.3944
R17643 gnd.n5936 gnd.n2680 19.3944
R17644 gnd.n1689 gnd.t302 18.8012
R17645 gnd.n1674 gnd.t141 18.8012
R17646 gnd.n1533 gnd.n1532 18.4825
R17647 gnd.n4594 gnd.n4593 18.4825
R17648 gnd.n4686 gnd.t165 18.4825
R17649 gnd.t2 gnd.n3046 18.4825
R17650 gnd.n4911 gnd.n2983 18.4825
R17651 gnd.n5875 gnd.n5874 18.4247
R17652 gnd.n4482 gnd.n3360 18.4247
R17653 gnd.n5275 gnd.n5260 18.2308
R17654 gnd.n3668 gnd.n3377 18.2308
R17655 gnd.n238 gnd.n180 18.2308
R17656 gnd.n3857 gnd.n3843 18.2308
R17657 gnd.t303 gnd.n1213 18.1639
R17658 gnd.n1819 gnd.n1004 17.8452
R17659 gnd.n1241 gnd.t299 17.5266
R17660 gnd.n4556 gnd.n3222 17.2079
R17661 gnd.n3492 gnd.n3208 17.2079
R17662 gnd.n4668 gnd.n3148 17.2079
R17663 gnd.n4871 gnd.n3039 17.2079
R17664 gnd.n4984 gnd.n2979 17.2079
R17665 gnd.n1640 gnd.t296 16.8893
R17666 gnd.n3848 gnd.t190 16.8893
R17667 gnd.n4246 gnd.t52 16.8893
R17668 gnd.t24 gnd.n5374 16.8893
R17669 gnd.n7339 gnd.t194 16.8893
R17670 gnd.n5857 gnd.n5854 16.6793
R17671 gnd.n7258 gnd.n7255 16.6793
R17672 gnd.n4052 gnd.n3918 16.6793
R17673 gnd.n4464 gnd.n4463 16.6793
R17674 gnd.n4679 gnd.t152 16.5706
R17675 gnd.n4842 gnd.t164 16.5706
R17676 gnd.n1468 gnd.t176 16.2519
R17677 gnd.n1168 gnd.t294 16.2519
R17678 gnd.n3709 gnd.t73 16.2519
R17679 gnd.n6062 gnd.t242 16.2519
R17680 gnd.t223 gnd.n2839 16.2519
R17681 gnd.t48 gnd.n5413 16.2519
R17682 gnd.n4567 gnd.n3212 15.9333
R17683 gnd.n4678 gnd.n3139 15.9333
R17684 gnd.n3139 gnd.n3132 15.9333
R17685 gnd.n4861 gnd.n4860 15.9333
R17686 gnd.n4860 gnd.n3050 15.9333
R17687 gnd.n2157 gnd.n2155 15.6674
R17688 gnd.n2125 gnd.n2123 15.6674
R17689 gnd.n2093 gnd.n2091 15.6674
R17690 gnd.n2062 gnd.n2060 15.6674
R17691 gnd.n2030 gnd.n2028 15.6674
R17692 gnd.n1998 gnd.n1996 15.6674
R17693 gnd.n1966 gnd.n1964 15.6674
R17694 gnd.n1935 gnd.n1933 15.6674
R17695 gnd.n1459 gnd.t176 15.6146
R17696 gnd.t215 gnd.n923 15.6146
R17697 gnd.t180 gnd.n924 15.6146
R17698 gnd.n3720 gnd.t70 15.6146
R17699 gnd.n3449 gnd.t242 15.6146
R17700 gnd.n4625 gnd.t136 15.6146
R17701 gnd.n4941 gnd.t167 15.6146
R17702 gnd.n5177 gnd.t223 15.6146
R17703 gnd.n5720 gnd.t44 15.6146
R17704 gnd.n5814 gnd.n2811 15.3217
R17705 gnd.n7213 gnd.n7208 15.3217
R17706 gnd.n4104 gnd.n3897 15.3217
R17707 gnd.n4424 gnd.n4420 15.3217
R17708 gnd.n2896 gnd.n2895 15.0827
R17709 gnd.n3234 gnd.n3229 15.0481
R17710 gnd.n2906 gnd.n2905 15.0481
R17711 gnd.n1829 gnd.t300 14.9773
R17712 gnd.n3812 gnd.t22 14.9773
R17713 gnd.n6092 gnd.t219 14.9773
R17714 gnd.t313 gnd.n4694 14.9773
R17715 gnd.n3061 gnd.t162 14.9773
R17716 gnd.n5495 gnd.t198 14.9773
R17717 gnd.n5694 gnd.t58 14.9773
R17718 gnd.n3494 gnd.n3492 14.6587
R17719 gnd.n4607 gnd.t155 14.6587
R17720 gnd.n4670 gnd.n4668 14.6587
R17721 gnd.n4694 gnd.n3118 14.6587
R17722 gnd.n3062 gnd.n3061 14.6587
R17723 gnd.n4814 gnd.n3039 14.6587
R17724 gnd.t7 gnd.n4958 14.6587
R17725 gnd.n4985 gnd.n4984 14.6587
R17726 gnd.n5127 gnd.n2888 14.6587
R17727 gnd.t158 gnd.n966 14.34
R17728 gnd.n1907 gnd.t297 14.34
R17729 gnd.n1615 gnd.t315 13.7027
R17730 gnd.n1325 gnd.n1324 13.5763
R17731 gnd.n2271 gnd.n880 13.5763
R17732 gnd.n1533 gnd.n1271 13.384
R17733 gnd.n3159 gnd.n3158 13.384
R17734 gnd.n3158 gnd.t166 13.384
R17735 gnd.n4714 gnd.n3114 13.384
R17736 gnd.n4803 gnd.n3066 13.384
R17737 gnd.t145 gnd.n3022 13.384
R17738 gnd.n4894 gnd.n3022 13.384
R17739 gnd.n4913 gnd.n4911 13.384
R17740 gnd.n3245 gnd.n3226 13.1884
R17741 gnd.n3240 gnd.n3239 13.1884
R17742 gnd.n3239 gnd.n3238 13.1884
R17743 gnd.n2899 gnd.n2894 13.1884
R17744 gnd.n2900 gnd.n2899 13.1884
R17745 gnd.n3241 gnd.n3228 13.146
R17746 gnd.n3237 gnd.n3228 13.146
R17747 gnd.n2898 gnd.n2897 13.146
R17748 gnd.n2898 gnd.n2893 13.146
R17749 gnd.t160 gnd.n4566 13.0654
R17750 gnd.n4993 gnd.t169 13.0654
R17751 gnd.n2158 gnd.n2154 12.8005
R17752 gnd.n2126 gnd.n2122 12.8005
R17753 gnd.n2094 gnd.n2090 12.8005
R17754 gnd.n2063 gnd.n2059 12.8005
R17755 gnd.n2031 gnd.n2027 12.8005
R17756 gnd.n1999 gnd.n1995 12.8005
R17757 gnd.n1967 gnd.n1963 12.8005
R17758 gnd.n1936 gnd.n1932 12.8005
R17759 gnd.t205 gnd.t172 12.7467
R17760 gnd.n1324 gnd.n1319 12.4126
R17761 gnd.n2274 gnd.n2271 12.4126
R17762 gnd.n4550 gnd.n4549 12.1761
R17763 gnd.n5124 gnd.n5123 12.1761
R17764 gnd.n4577 gnd.n3185 12.1094
R17765 gnd.t6 gnd.n3164 12.1094
R17766 gnd.n4904 gnd.t133 12.1094
R17767 gnd.n4959 gnd.n2992 12.1094
R17768 gnd.t227 gnd.n2976 12.1094
R17769 gnd.n5128 gnd.t184 12.1094
R17770 gnd.n2162 gnd.n2161 12.0247
R17771 gnd.n2130 gnd.n2129 12.0247
R17772 gnd.n2098 gnd.n2097 12.0247
R17773 gnd.n2067 gnd.n2066 12.0247
R17774 gnd.n2035 gnd.n2034 12.0247
R17775 gnd.n2003 gnd.n2002 12.0247
R17776 gnd.n1971 gnd.n1970 12.0247
R17777 gnd.n1940 gnd.n1939 12.0247
R17778 gnd.n6197 gnd.t22 11.7908
R17779 gnd.n2540 gnd.t219 11.7908
R17780 gnd.t198 gnd.n5321 11.7908
R17781 gnd.n7364 gnd.t58 11.7908
R17782 gnd.t187 gnd.n3222 11.4721
R17783 gnd.n4714 gnd.t3 11.4721
R17784 gnd.n4803 gnd.t10 11.4721
R17785 gnd.n2165 gnd.n2152 11.249
R17786 gnd.n2133 gnd.n2120 11.249
R17787 gnd.n2101 gnd.n2088 11.249
R17788 gnd.n2070 gnd.n2057 11.249
R17789 gnd.n2038 gnd.n2025 11.249
R17790 gnd.n2006 gnd.n1993 11.249
R17791 gnd.n1974 gnd.n1961 11.249
R17792 gnd.n1943 gnd.n1930 11.249
R17793 gnd.n1603 gnd.t315 11.1535
R17794 gnd.n6173 gnd.t70 11.1535
R17795 gnd.n3461 gnd.t156 11.1535
R17796 gnd.n4662 gnd.t8 11.1535
R17797 gnd.n4881 gnd.t148 11.1535
R17798 gnd.n5160 gnd.t309 11.1535
R17799 gnd.n7388 gnd.t44 11.1535
R17800 gnd.n4626 gnd.n4625 10.8348
R17801 gnd.n4762 gnd.n3091 10.8348
R17802 gnd.n4762 gnd.n3092 10.8348
R17803 gnd.n4941 gnd.n4940 10.8348
R17804 gnd.n5817 gnd.n5814 10.6672
R17805 gnd.n7216 gnd.n7213 10.6672
R17806 gnd.n3898 gnd.n3897 10.6672
R17807 gnd.n4429 gnd.n4420 10.6672
R17808 gnd.n5059 gnd.n2936 10.6151
R17809 gnd.n5059 gnd.n5058 10.6151
R17810 gnd.n5056 gnd.n2940 10.6151
R17811 gnd.n5051 gnd.n2940 10.6151
R17812 gnd.n5051 gnd.n5050 10.6151
R17813 gnd.n5050 gnd.n5049 10.6151
R17814 gnd.n5049 gnd.n2943 10.6151
R17815 gnd.n5044 gnd.n2943 10.6151
R17816 gnd.n5044 gnd.n5043 10.6151
R17817 gnd.n5043 gnd.n5042 10.6151
R17818 gnd.n5042 gnd.n2946 10.6151
R17819 gnd.n5037 gnd.n2946 10.6151
R17820 gnd.n5037 gnd.n5036 10.6151
R17821 gnd.n5036 gnd.n5035 10.6151
R17822 gnd.n5035 gnd.n2949 10.6151
R17823 gnd.n5030 gnd.n2949 10.6151
R17824 gnd.n5030 gnd.n5029 10.6151
R17825 gnd.n5029 gnd.n5028 10.6151
R17826 gnd.n5028 gnd.n2952 10.6151
R17827 gnd.n5023 gnd.n2952 10.6151
R17828 gnd.n5023 gnd.n5022 10.6151
R17829 gnd.n5022 gnd.n5021 10.6151
R17830 gnd.n5021 gnd.n2955 10.6151
R17831 gnd.n5016 gnd.n2955 10.6151
R17832 gnd.n5016 gnd.n5015 10.6151
R17833 gnd.n5015 gnd.n5014 10.6151
R17834 gnd.n5014 gnd.n2958 10.6151
R17835 gnd.n5009 gnd.n2958 10.6151
R17836 gnd.n5009 gnd.n5008 10.6151
R17837 gnd.n5008 gnd.n5007 10.6151
R17838 gnd.n3293 gnd.n3292 10.6151
R17839 gnd.n3292 gnd.n3291 10.6151
R17840 gnd.n3291 gnd.n3288 10.6151
R17841 gnd.n3288 gnd.n3206 10.6151
R17842 gnd.n4575 gnd.n3206 10.6151
R17843 gnd.n4576 gnd.n4575 10.6151
R17844 gnd.n4585 gnd.n4576 10.6151
R17845 gnd.n4585 gnd.n4584 10.6151
R17846 gnd.n4584 gnd.n4583 10.6151
R17847 gnd.n4583 gnd.n4582 10.6151
R17848 gnd.n4582 gnd.n4580 10.6151
R17849 gnd.n4580 gnd.n4579 10.6151
R17850 gnd.n4579 gnd.n3182 10.6151
R17851 gnd.n4617 gnd.n3182 10.6151
R17852 gnd.n4618 gnd.n4617 10.6151
R17853 gnd.n4623 gnd.n4618 10.6151
R17854 gnd.n4623 gnd.n4622 10.6151
R17855 gnd.n4622 gnd.n4621 10.6151
R17856 gnd.n4621 gnd.n4619 10.6151
R17857 gnd.n4619 gnd.n3155 10.6151
R17858 gnd.n4652 gnd.n3155 10.6151
R17859 gnd.n4653 gnd.n4652 10.6151
R17860 gnd.n4660 gnd.n4653 10.6151
R17861 gnd.n4660 gnd.n4659 10.6151
R17862 gnd.n4659 gnd.n4658 10.6151
R17863 gnd.n4658 gnd.n4657 10.6151
R17864 gnd.n4657 gnd.n4654 10.6151
R17865 gnd.n4654 gnd.n3130 10.6151
R17866 gnd.n4688 gnd.n3130 10.6151
R17867 gnd.n4689 gnd.n4688 10.6151
R17868 gnd.n4692 gnd.n4689 10.6151
R17869 gnd.n4692 gnd.n4691 10.6151
R17870 gnd.n4691 gnd.n4690 10.6151
R17871 gnd.n4690 gnd.n3112 10.6151
R17872 gnd.n4717 gnd.n3112 10.6151
R17873 gnd.n4718 gnd.n4717 10.6151
R17874 gnd.n4735 gnd.n4718 10.6151
R17875 gnd.n4735 gnd.n4734 10.6151
R17876 gnd.n4734 gnd.n4733 10.6151
R17877 gnd.n4733 gnd.n4719 10.6151
R17878 gnd.n4729 gnd.n4719 10.6151
R17879 gnd.n4729 gnd.n4728 10.6151
R17880 gnd.n4728 gnd.n4727 10.6151
R17881 gnd.n4727 gnd.n4726 10.6151
R17882 gnd.n4726 gnd.n4724 10.6151
R17883 gnd.n4724 gnd.n4723 10.6151
R17884 gnd.n4723 gnd.n4721 10.6151
R17885 gnd.n4721 gnd.n3058 10.6151
R17886 gnd.n4811 gnd.n3058 10.6151
R17887 gnd.n4812 gnd.n4811 10.6151
R17888 gnd.n4847 gnd.n4812 10.6151
R17889 gnd.n4847 gnd.n4846 10.6151
R17890 gnd.n4846 gnd.n4845 10.6151
R17891 gnd.n4845 gnd.n4844 10.6151
R17892 gnd.n4844 gnd.n4813 10.6151
R17893 gnd.n4839 gnd.n4813 10.6151
R17894 gnd.n4839 gnd.n4838 10.6151
R17895 gnd.n4838 gnd.n4837 10.6151
R17896 gnd.n4837 gnd.n4836 10.6151
R17897 gnd.n4836 gnd.n4834 10.6151
R17898 gnd.n4834 gnd.n4833 10.6151
R17899 gnd.n4833 gnd.n4817 10.6151
R17900 gnd.n4829 gnd.n4817 10.6151
R17901 gnd.n4829 gnd.n4828 10.6151
R17902 gnd.n4828 gnd.n4827 10.6151
R17903 gnd.n4827 gnd.n4826 10.6151
R17904 gnd.n4826 gnd.n4824 10.6151
R17905 gnd.n4824 gnd.n4823 10.6151
R17906 gnd.n4823 gnd.n4821 10.6151
R17907 gnd.n4821 gnd.n2986 10.6151
R17908 gnd.n4967 gnd.n2986 10.6151
R17909 gnd.n4968 gnd.n4967 10.6151
R17910 gnd.n4976 gnd.n4968 10.6151
R17911 gnd.n4976 gnd.n4975 10.6151
R17912 gnd.n4975 gnd.n4974 10.6151
R17913 gnd.n4974 gnd.n4973 10.6151
R17914 gnd.n4973 gnd.n4970 10.6151
R17915 gnd.n4970 gnd.n4969 10.6151
R17916 gnd.n4969 gnd.n2961 10.6151
R17917 gnd.n5003 gnd.n2961 10.6151
R17918 gnd.n5004 gnd.n5003 10.6151
R17919 gnd.n3358 gnd.n3357 10.6151
R17920 gnd.n3357 gnd.n3354 10.6151
R17921 gnd.n3352 gnd.n3349 10.6151
R17922 gnd.n3349 gnd.n3348 10.6151
R17923 gnd.n3348 gnd.n3345 10.6151
R17924 gnd.n3345 gnd.n3344 10.6151
R17925 gnd.n3344 gnd.n3341 10.6151
R17926 gnd.n3341 gnd.n3340 10.6151
R17927 gnd.n3340 gnd.n3337 10.6151
R17928 gnd.n3337 gnd.n3336 10.6151
R17929 gnd.n3336 gnd.n3333 10.6151
R17930 gnd.n3333 gnd.n3332 10.6151
R17931 gnd.n3332 gnd.n3329 10.6151
R17932 gnd.n3329 gnd.n3328 10.6151
R17933 gnd.n3328 gnd.n3325 10.6151
R17934 gnd.n3325 gnd.n3324 10.6151
R17935 gnd.n3324 gnd.n3321 10.6151
R17936 gnd.n3321 gnd.n3320 10.6151
R17937 gnd.n3320 gnd.n3317 10.6151
R17938 gnd.n3317 gnd.n3316 10.6151
R17939 gnd.n3316 gnd.n3313 10.6151
R17940 gnd.n3313 gnd.n3312 10.6151
R17941 gnd.n3312 gnd.n3309 10.6151
R17942 gnd.n3309 gnd.n3308 10.6151
R17943 gnd.n3308 gnd.n3305 10.6151
R17944 gnd.n3305 gnd.n3304 10.6151
R17945 gnd.n3304 gnd.n3301 10.6151
R17946 gnd.n3301 gnd.n3300 10.6151
R17947 gnd.n3300 gnd.n3297 10.6151
R17948 gnd.n3297 gnd.n3296 10.6151
R17949 gnd.n4549 gnd.n3246 10.6151
R17950 gnd.n4544 gnd.n3246 10.6151
R17951 gnd.n4544 gnd.n4543 10.6151
R17952 gnd.n4543 gnd.n4542 10.6151
R17953 gnd.n4542 gnd.n4539 10.6151
R17954 gnd.n4539 gnd.n4538 10.6151
R17955 gnd.n4538 gnd.n4535 10.6151
R17956 gnd.n4535 gnd.n4534 10.6151
R17957 gnd.n4534 gnd.n4531 10.6151
R17958 gnd.n4531 gnd.n4530 10.6151
R17959 gnd.n4530 gnd.n4527 10.6151
R17960 gnd.n4527 gnd.n4526 10.6151
R17961 gnd.n4526 gnd.n4523 10.6151
R17962 gnd.n4523 gnd.n4522 10.6151
R17963 gnd.n4522 gnd.n4519 10.6151
R17964 gnd.n4519 gnd.n4518 10.6151
R17965 gnd.n4518 gnd.n4515 10.6151
R17966 gnd.n4515 gnd.n4514 10.6151
R17967 gnd.n4514 gnd.n4511 10.6151
R17968 gnd.n4511 gnd.n4510 10.6151
R17969 gnd.n4510 gnd.n4507 10.6151
R17970 gnd.n4507 gnd.n4506 10.6151
R17971 gnd.n4506 gnd.n4503 10.6151
R17972 gnd.n4503 gnd.n4502 10.6151
R17973 gnd.n4502 gnd.n4499 10.6151
R17974 gnd.n4499 gnd.n4498 10.6151
R17975 gnd.n4498 gnd.n4495 10.6151
R17976 gnd.n4495 gnd.n4494 10.6151
R17977 gnd.n4491 gnd.n4490 10.6151
R17978 gnd.n4490 gnd.n4487 10.6151
R17979 gnd.n5123 gnd.n5122 10.6151
R17980 gnd.n5122 gnd.n2911 10.6151
R17981 gnd.n5117 gnd.n2911 10.6151
R17982 gnd.n5117 gnd.n5116 10.6151
R17983 gnd.n5116 gnd.n5115 10.6151
R17984 gnd.n5115 gnd.n2914 10.6151
R17985 gnd.n5110 gnd.n2914 10.6151
R17986 gnd.n5110 gnd.n5109 10.6151
R17987 gnd.n5109 gnd.n5108 10.6151
R17988 gnd.n5108 gnd.n2917 10.6151
R17989 gnd.n5103 gnd.n2917 10.6151
R17990 gnd.n5103 gnd.n5102 10.6151
R17991 gnd.n5102 gnd.n5101 10.6151
R17992 gnd.n5101 gnd.n2920 10.6151
R17993 gnd.n5096 gnd.n2920 10.6151
R17994 gnd.n5096 gnd.n5095 10.6151
R17995 gnd.n5095 gnd.n5094 10.6151
R17996 gnd.n5094 gnd.n2923 10.6151
R17997 gnd.n5089 gnd.n2923 10.6151
R17998 gnd.n5089 gnd.n5088 10.6151
R17999 gnd.n5088 gnd.n5087 10.6151
R18000 gnd.n5087 gnd.n2926 10.6151
R18001 gnd.n5082 gnd.n2926 10.6151
R18002 gnd.n5082 gnd.n5081 10.6151
R18003 gnd.n5081 gnd.n5080 10.6151
R18004 gnd.n5080 gnd.n2929 10.6151
R18005 gnd.n5075 gnd.n2929 10.6151
R18006 gnd.n5075 gnd.n5074 10.6151
R18007 gnd.n5072 gnd.n2934 10.6151
R18008 gnd.n5067 gnd.n2934 10.6151
R18009 gnd.n4552 gnd.n4551 10.6151
R18010 gnd.n4552 gnd.n3210 10.6151
R18011 gnd.n4569 gnd.n3210 10.6151
R18012 gnd.n4570 gnd.n4569 10.6151
R18013 gnd.n4571 gnd.n4570 10.6151
R18014 gnd.n4571 gnd.n3202 10.6151
R18015 gnd.n4589 gnd.n3202 10.6151
R18016 gnd.n4590 gnd.n4589 10.6151
R18017 gnd.n4591 gnd.n4590 10.6151
R18018 gnd.n4591 gnd.n3187 10.6151
R18019 gnd.n4610 gnd.n3187 10.6151
R18020 gnd.n4611 gnd.n4610 10.6151
R18021 gnd.n4612 gnd.n4611 10.6151
R18022 gnd.n4612 gnd.n3177 10.6151
R18023 gnd.n4629 gnd.n3177 10.6151
R18024 gnd.n4630 gnd.n4629 10.6151
R18025 gnd.n4631 gnd.n4630 10.6151
R18026 gnd.n4631 gnd.n3161 10.6151
R18027 gnd.n4646 gnd.n3161 10.6151
R18028 gnd.n4647 gnd.n4646 10.6151
R18029 gnd.n4648 gnd.n4647 10.6151
R18030 gnd.n4648 gnd.n3150 10.6151
R18031 gnd.n4664 gnd.n3150 10.6151
R18032 gnd.n4665 gnd.n4664 10.6151
R18033 gnd.n4666 gnd.n4665 10.6151
R18034 gnd.n4666 gnd.n3135 10.6151
R18035 gnd.n4681 gnd.n3135 10.6151
R18036 gnd.n4682 gnd.n4681 10.6151
R18037 gnd.n4684 gnd.n4682 10.6151
R18038 gnd.n4684 gnd.n4683 10.6151
R18039 gnd.n4683 gnd.n3116 10.6151
R18040 gnd.n4710 gnd.n3116 10.6151
R18041 gnd.n4711 gnd.n4710 10.6151
R18042 gnd.n4712 gnd.n4711 10.6151
R18043 gnd.n4712 gnd.n3107 10.6151
R18044 gnd.n4742 gnd.n3107 10.6151
R18045 gnd.n4743 gnd.n4742 10.6151
R18046 gnd.n4749 gnd.n4743 10.6151
R18047 gnd.n4749 gnd.n4748 10.6151
R18048 gnd.n4748 gnd.n4747 10.6151
R18049 gnd.n4747 gnd.n4744 10.6151
R18050 gnd.n4744 gnd.n3081 10.6151
R18051 gnd.n4787 gnd.n3081 10.6151
R18052 gnd.n4788 gnd.n4787 10.6151
R18053 gnd.n4789 gnd.n4788 10.6151
R18054 gnd.n4789 gnd.n3064 10.6151
R18055 gnd.n4805 gnd.n3064 10.6151
R18056 gnd.n4806 gnd.n4805 10.6151
R18057 gnd.n4807 gnd.n4806 10.6151
R18058 gnd.n4807 gnd.n3053 10.6151
R18059 gnd.n4851 gnd.n3053 10.6151
R18060 gnd.n4852 gnd.n4851 10.6151
R18061 gnd.n4858 gnd.n4852 10.6151
R18062 gnd.n4858 gnd.n4857 10.6151
R18063 gnd.n4857 gnd.n4856 10.6151
R18064 gnd.n4856 gnd.n4853 10.6151
R18065 gnd.n4853 gnd.n3029 10.6151
R18066 gnd.n4883 gnd.n3029 10.6151
R18067 gnd.n4884 gnd.n4883 10.6151
R18068 gnd.n4890 gnd.n4884 10.6151
R18069 gnd.n4890 gnd.n4889 10.6151
R18070 gnd.n4889 gnd.n4888 10.6151
R18071 gnd.n4888 gnd.n4885 10.6151
R18072 gnd.n4885 gnd.n3006 10.6151
R18073 gnd.n4943 gnd.n3006 10.6151
R18074 gnd.n4944 gnd.n4943 10.6151
R18075 gnd.n4945 gnd.n4944 10.6151
R18076 gnd.n4945 gnd.n2990 10.6151
R18077 gnd.n4961 gnd.n2990 10.6151
R18078 gnd.n4962 gnd.n4961 10.6151
R18079 gnd.n4963 gnd.n4962 10.6151
R18080 gnd.n4963 gnd.n2981 10.6151
R18081 gnd.n4980 gnd.n2981 10.6151
R18082 gnd.n4981 gnd.n4980 10.6151
R18083 gnd.n4982 gnd.n4981 10.6151
R18084 gnd.n4982 gnd.n2965 10.6151
R18085 gnd.n4996 gnd.n2965 10.6151
R18086 gnd.n4997 gnd.n4996 10.6151
R18087 gnd.n4998 gnd.n4997 10.6151
R18088 gnd.n4998 gnd.n2891 10.6151
R18089 gnd.n5125 gnd.n2891 10.6151
R18090 gnd.n1522 gnd.t318 10.5161
R18091 gnd.n968 gnd.t158 10.5161
R18092 gnd.n1890 gnd.t297 10.5161
R18093 gnd.n6147 gnd.t73 10.5161
R18094 gnd.t8 gnd.n3145 10.5161
R18095 gnd.n4815 gnd.t148 10.5161
R18096 gnd.n5414 gnd.t48 10.5161
R18097 gnd.n2166 gnd.n2150 10.4732
R18098 gnd.n2134 gnd.n2118 10.4732
R18099 gnd.n2102 gnd.n2086 10.4732
R18100 gnd.n2071 gnd.n2055 10.4732
R18101 gnd.n2039 gnd.n2023 10.4732
R18102 gnd.n2007 gnd.n1991 10.4732
R18103 gnd.n1975 gnd.n1959 10.4732
R18104 gnd.n1944 gnd.n1928 10.4732
R18105 gnd.t300 gnd.n985 9.87883
R18106 gnd.t190 gnd.n2334 9.87883
R18107 gnd.n6122 gnd.t52 9.87883
R18108 gnd.n4752 gnd.t0 9.87883
R18109 gnd.n4784 gnd.t134 9.87883
R18110 gnd.n5525 gnd.t24 9.87883
R18111 gnd.t194 gnd.n160 9.87883
R18112 gnd.n2170 gnd.n2169 9.69747
R18113 gnd.n2138 gnd.n2137 9.69747
R18114 gnd.n2106 gnd.n2105 9.69747
R18115 gnd.n2075 gnd.n2074 9.69747
R18116 gnd.n2043 gnd.n2042 9.69747
R18117 gnd.n2011 gnd.n2010 9.69747
R18118 gnd.n1979 gnd.n1978 9.69747
R18119 gnd.n1948 gnd.n1947 9.69747
R18120 gnd.n4614 gnd.n3185 9.56018
R18121 gnd.n3175 gnd.n3164 9.56018
R18122 gnd.n4752 gnd.n4751 9.56018
R18123 gnd.n4785 gnd.n4784 9.56018
R18124 gnd.n4904 gnd.n3015 9.56018
R18125 gnd.n3004 gnd.n2992 9.56018
R18126 gnd.n4978 gnd.t227 9.56018
R18127 gnd.n2176 gnd.n2175 9.45567
R18128 gnd.n2144 gnd.n2143 9.45567
R18129 gnd.n2112 gnd.n2111 9.45567
R18130 gnd.n2081 gnd.n2080 9.45567
R18131 gnd.n2049 gnd.n2048 9.45567
R18132 gnd.n2017 gnd.n2016 9.45567
R18133 gnd.n1985 gnd.n1984 9.45567
R18134 gnd.n1954 gnd.n1953 9.45567
R18135 gnd.n5854 gnd.n5853 9.30959
R18136 gnd.n7255 gnd.n7187 9.30959
R18137 gnd.n4052 gnd.n3916 9.30959
R18138 gnd.n4463 gnd.n4384 9.30959
R18139 gnd.n2175 gnd.n2174 9.3005
R18140 gnd.n2148 gnd.n2147 9.3005
R18141 gnd.n2169 gnd.n2168 9.3005
R18142 gnd.n2167 gnd.n2166 9.3005
R18143 gnd.n2152 gnd.n2151 9.3005
R18144 gnd.n2161 gnd.n2160 9.3005
R18145 gnd.n2159 gnd.n2158 9.3005
R18146 gnd.n2143 gnd.n2142 9.3005
R18147 gnd.n2116 gnd.n2115 9.3005
R18148 gnd.n2137 gnd.n2136 9.3005
R18149 gnd.n2135 gnd.n2134 9.3005
R18150 gnd.n2120 gnd.n2119 9.3005
R18151 gnd.n2129 gnd.n2128 9.3005
R18152 gnd.n2127 gnd.n2126 9.3005
R18153 gnd.n2111 gnd.n2110 9.3005
R18154 gnd.n2084 gnd.n2083 9.3005
R18155 gnd.n2105 gnd.n2104 9.3005
R18156 gnd.n2103 gnd.n2102 9.3005
R18157 gnd.n2088 gnd.n2087 9.3005
R18158 gnd.n2097 gnd.n2096 9.3005
R18159 gnd.n2095 gnd.n2094 9.3005
R18160 gnd.n2080 gnd.n2079 9.3005
R18161 gnd.n2053 gnd.n2052 9.3005
R18162 gnd.n2074 gnd.n2073 9.3005
R18163 gnd.n2072 gnd.n2071 9.3005
R18164 gnd.n2057 gnd.n2056 9.3005
R18165 gnd.n2066 gnd.n2065 9.3005
R18166 gnd.n2064 gnd.n2063 9.3005
R18167 gnd.n2048 gnd.n2047 9.3005
R18168 gnd.n2021 gnd.n2020 9.3005
R18169 gnd.n2042 gnd.n2041 9.3005
R18170 gnd.n2040 gnd.n2039 9.3005
R18171 gnd.n2025 gnd.n2024 9.3005
R18172 gnd.n2034 gnd.n2033 9.3005
R18173 gnd.n2032 gnd.n2031 9.3005
R18174 gnd.n2016 gnd.n2015 9.3005
R18175 gnd.n1989 gnd.n1988 9.3005
R18176 gnd.n2010 gnd.n2009 9.3005
R18177 gnd.n2008 gnd.n2007 9.3005
R18178 gnd.n1993 gnd.n1992 9.3005
R18179 gnd.n2002 gnd.n2001 9.3005
R18180 gnd.n2000 gnd.n1999 9.3005
R18181 gnd.n1984 gnd.n1983 9.3005
R18182 gnd.n1957 gnd.n1956 9.3005
R18183 gnd.n1978 gnd.n1977 9.3005
R18184 gnd.n1976 gnd.n1975 9.3005
R18185 gnd.n1961 gnd.n1960 9.3005
R18186 gnd.n1970 gnd.n1969 9.3005
R18187 gnd.n1968 gnd.n1967 9.3005
R18188 gnd.n1953 gnd.n1952 9.3005
R18189 gnd.n1926 gnd.n1925 9.3005
R18190 gnd.n1947 gnd.n1946 9.3005
R18191 gnd.n1945 gnd.n1944 9.3005
R18192 gnd.n1930 gnd.n1929 9.3005
R18193 gnd.n1939 gnd.n1938 9.3005
R18194 gnd.n1937 gnd.n1936 9.3005
R18195 gnd.n2301 gnd.n2300 9.3005
R18196 gnd.n2299 gnd.n868 9.3005
R18197 gnd.n2298 gnd.n2297 9.3005
R18198 gnd.n2294 gnd.n869 9.3005
R18199 gnd.n2291 gnd.n870 9.3005
R18200 gnd.n2290 gnd.n871 9.3005
R18201 gnd.n2287 gnd.n872 9.3005
R18202 gnd.n2286 gnd.n873 9.3005
R18203 gnd.n2283 gnd.n874 9.3005
R18204 gnd.n2282 gnd.n875 9.3005
R18205 gnd.n2279 gnd.n876 9.3005
R18206 gnd.n2278 gnd.n877 9.3005
R18207 gnd.n2275 gnd.n878 9.3005
R18208 gnd.n2274 gnd.n879 9.3005
R18209 gnd.n2271 gnd.n2270 9.3005
R18210 gnd.n2269 gnd.n880 9.3005
R18211 gnd.n2302 gnd.n867 9.3005
R18212 gnd.n1541 gnd.n1540 9.3005
R18213 gnd.n1245 gnd.n1244 9.3005
R18214 gnd.n1568 gnd.n1567 9.3005
R18215 gnd.n1569 gnd.n1243 9.3005
R18216 gnd.n1573 gnd.n1570 9.3005
R18217 gnd.n1572 gnd.n1571 9.3005
R18218 gnd.n1217 gnd.n1216 9.3005
R18219 gnd.n1598 gnd.n1597 9.3005
R18220 gnd.n1599 gnd.n1215 9.3005
R18221 gnd.n1601 gnd.n1600 9.3005
R18222 gnd.n1195 gnd.n1194 9.3005
R18223 gnd.n1629 gnd.n1628 9.3005
R18224 gnd.n1630 gnd.n1193 9.3005
R18225 gnd.n1638 gnd.n1631 9.3005
R18226 gnd.n1637 gnd.n1632 9.3005
R18227 gnd.n1636 gnd.n1634 9.3005
R18228 gnd.n1633 gnd.n1142 9.3005
R18229 gnd.n1686 gnd.n1143 9.3005
R18230 gnd.n1685 gnd.n1144 9.3005
R18231 gnd.n1684 gnd.n1145 9.3005
R18232 gnd.n1164 gnd.n1146 9.3005
R18233 gnd.n1166 gnd.n1165 9.3005
R18234 gnd.n1064 gnd.n1063 9.3005
R18235 gnd.n1724 gnd.n1723 9.3005
R18236 gnd.n1725 gnd.n1062 9.3005
R18237 gnd.n1729 gnd.n1726 9.3005
R18238 gnd.n1728 gnd.n1727 9.3005
R18239 gnd.n1037 gnd.n1036 9.3005
R18240 gnd.n1764 gnd.n1763 9.3005
R18241 gnd.n1765 gnd.n1035 9.3005
R18242 gnd.n1769 gnd.n1766 9.3005
R18243 gnd.n1768 gnd.n1767 9.3005
R18244 gnd.n1011 gnd.n1010 9.3005
R18245 gnd.n1811 gnd.n1810 9.3005
R18246 gnd.n1812 gnd.n1009 9.3005
R18247 gnd.n1816 gnd.n1813 9.3005
R18248 gnd.n1815 gnd.n1814 9.3005
R18249 gnd.n983 gnd.n982 9.3005
R18250 gnd.n1851 gnd.n1850 9.3005
R18251 gnd.n1852 gnd.n981 9.3005
R18252 gnd.n1856 gnd.n1853 9.3005
R18253 gnd.n1855 gnd.n1854 9.3005
R18254 gnd.n956 gnd.n955 9.3005
R18255 gnd.n1900 gnd.n1899 9.3005
R18256 gnd.n1901 gnd.n954 9.3005
R18257 gnd.n1905 gnd.n1902 9.3005
R18258 gnd.n1904 gnd.n1903 9.3005
R18259 gnd.n929 gnd.n928 9.3005
R18260 gnd.n2194 gnd.n2193 9.3005
R18261 gnd.n2195 gnd.n927 9.3005
R18262 gnd.n2201 gnd.n2196 9.3005
R18263 gnd.n2200 gnd.n2197 9.3005
R18264 gnd.n2199 gnd.n2198 9.3005
R18265 gnd.n1542 gnd.n1539 9.3005
R18266 gnd.n1324 gnd.n1283 9.3005
R18267 gnd.n1319 gnd.n1318 9.3005
R18268 gnd.n1317 gnd.n1284 9.3005
R18269 gnd.n1316 gnd.n1315 9.3005
R18270 gnd.n1312 gnd.n1285 9.3005
R18271 gnd.n1309 gnd.n1308 9.3005
R18272 gnd.n1307 gnd.n1286 9.3005
R18273 gnd.n1306 gnd.n1305 9.3005
R18274 gnd.n1302 gnd.n1287 9.3005
R18275 gnd.n1299 gnd.n1298 9.3005
R18276 gnd.n1297 gnd.n1288 9.3005
R18277 gnd.n1296 gnd.n1295 9.3005
R18278 gnd.n1292 gnd.n1290 9.3005
R18279 gnd.n1289 gnd.n1269 9.3005
R18280 gnd.n1536 gnd.n1268 9.3005
R18281 gnd.n1538 gnd.n1537 9.3005
R18282 gnd.n1326 gnd.n1325 9.3005
R18283 gnd.n1549 gnd.n1255 9.3005
R18284 gnd.n1556 gnd.n1256 9.3005
R18285 gnd.n1558 gnd.n1557 9.3005
R18286 gnd.n1559 gnd.n1236 9.3005
R18287 gnd.n1578 gnd.n1577 9.3005
R18288 gnd.n1580 gnd.n1228 9.3005
R18289 gnd.n1587 gnd.n1230 9.3005
R18290 gnd.n1588 gnd.n1225 9.3005
R18291 gnd.n1590 gnd.n1589 9.3005
R18292 gnd.n1226 gnd.n1211 9.3005
R18293 gnd.n1606 gnd.n1209 9.3005
R18294 gnd.n1610 gnd.n1609 9.3005
R18295 gnd.n1608 gnd.n1185 9.3005
R18296 gnd.n1645 gnd.n1184 9.3005
R18297 gnd.n1648 gnd.n1647 9.3005
R18298 gnd.n1181 gnd.n1180 9.3005
R18299 gnd.n1654 gnd.n1182 9.3005
R18300 gnd.n1656 gnd.n1655 9.3005
R18301 gnd.n1658 gnd.n1179 9.3005
R18302 gnd.n1661 gnd.n1660 9.3005
R18303 gnd.n1664 gnd.n1662 9.3005
R18304 gnd.n1666 gnd.n1665 9.3005
R18305 gnd.n1672 gnd.n1667 9.3005
R18306 gnd.n1671 gnd.n1670 9.3005
R18307 gnd.n1055 gnd.n1054 9.3005
R18308 gnd.n1738 gnd.n1737 9.3005
R18309 gnd.n1739 gnd.n1048 9.3005
R18310 gnd.n1747 gnd.n1047 9.3005
R18311 gnd.n1750 gnd.n1749 9.3005
R18312 gnd.n1752 gnd.n1751 9.3005
R18313 gnd.n1755 gnd.n1030 9.3005
R18314 gnd.n1753 gnd.n1028 9.3005
R18315 gnd.n1775 gnd.n1026 9.3005
R18316 gnd.n1777 gnd.n1776 9.3005
R18317 gnd.n1001 gnd.n1000 9.3005
R18318 gnd.n1825 gnd.n1824 9.3005
R18319 gnd.n1826 gnd.n994 9.3005
R18320 gnd.n1834 gnd.n993 9.3005
R18321 gnd.n1837 gnd.n1836 9.3005
R18322 gnd.n1839 gnd.n1838 9.3005
R18323 gnd.n1842 gnd.n976 9.3005
R18324 gnd.n1840 gnd.n974 9.3005
R18325 gnd.n1862 gnd.n972 9.3005
R18326 gnd.n1864 gnd.n1863 9.3005
R18327 gnd.n947 gnd.n946 9.3005
R18328 gnd.n1914 gnd.n1913 9.3005
R18329 gnd.n1915 gnd.n940 9.3005
R18330 gnd.n1923 gnd.n939 9.3005
R18331 gnd.n2182 gnd.n2181 9.3005
R18332 gnd.n2184 gnd.n2183 9.3005
R18333 gnd.n2185 gnd.n920 9.3005
R18334 gnd.n2209 gnd.n2208 9.3005
R18335 gnd.n921 gnd.n883 9.3005
R18336 gnd.n1547 gnd.n1546 9.3005
R18337 gnd.n2265 gnd.n884 9.3005
R18338 gnd.n2264 gnd.n886 9.3005
R18339 gnd.n2261 gnd.n887 9.3005
R18340 gnd.n2260 gnd.n888 9.3005
R18341 gnd.n2257 gnd.n889 9.3005
R18342 gnd.n2256 gnd.n890 9.3005
R18343 gnd.n2253 gnd.n891 9.3005
R18344 gnd.n2252 gnd.n892 9.3005
R18345 gnd.n2249 gnd.n893 9.3005
R18346 gnd.n2248 gnd.n894 9.3005
R18347 gnd.n2245 gnd.n895 9.3005
R18348 gnd.n2244 gnd.n896 9.3005
R18349 gnd.n2241 gnd.n897 9.3005
R18350 gnd.n2240 gnd.n898 9.3005
R18351 gnd.n2237 gnd.n899 9.3005
R18352 gnd.n2236 gnd.n900 9.3005
R18353 gnd.n2233 gnd.n901 9.3005
R18354 gnd.n2232 gnd.n902 9.3005
R18355 gnd.n2229 gnd.n903 9.3005
R18356 gnd.n2228 gnd.n904 9.3005
R18357 gnd.n2225 gnd.n905 9.3005
R18358 gnd.n2224 gnd.n906 9.3005
R18359 gnd.n2221 gnd.n910 9.3005
R18360 gnd.n2220 gnd.n911 9.3005
R18361 gnd.n2217 gnd.n912 9.3005
R18362 gnd.n2216 gnd.n913 9.3005
R18363 gnd.n2267 gnd.n2266 9.3005
R18364 gnd.n1716 gnd.n1700 9.3005
R18365 gnd.n1715 gnd.n1701 9.3005
R18366 gnd.n1714 gnd.n1702 9.3005
R18367 gnd.n1712 gnd.n1703 9.3005
R18368 gnd.n1711 gnd.n1704 9.3005
R18369 gnd.n1709 gnd.n1705 9.3005
R18370 gnd.n1708 gnd.n1706 9.3005
R18371 gnd.n1018 gnd.n1017 9.3005
R18372 gnd.n1785 gnd.n1784 9.3005
R18373 gnd.n1786 gnd.n1016 9.3005
R18374 gnd.n1803 gnd.n1787 9.3005
R18375 gnd.n1802 gnd.n1788 9.3005
R18376 gnd.n1801 gnd.n1789 9.3005
R18377 gnd.n1799 gnd.n1790 9.3005
R18378 gnd.n1798 gnd.n1791 9.3005
R18379 gnd.n1796 gnd.n1792 9.3005
R18380 gnd.n1795 gnd.n1793 9.3005
R18381 gnd.n963 gnd.n962 9.3005
R18382 gnd.n1872 gnd.n1871 9.3005
R18383 gnd.n1873 gnd.n961 9.3005
R18384 gnd.n1894 gnd.n1874 9.3005
R18385 gnd.n1893 gnd.n1875 9.3005
R18386 gnd.n1892 gnd.n1876 9.3005
R18387 gnd.n1889 gnd.n1877 9.3005
R18388 gnd.n1888 gnd.n1878 9.3005
R18389 gnd.n1886 gnd.n1879 9.3005
R18390 gnd.n1885 gnd.n1880 9.3005
R18391 gnd.n1883 gnd.n1882 9.3005
R18392 gnd.n1881 gnd.n915 9.3005
R18393 gnd.n1457 gnd.n1456 9.3005
R18394 gnd.n1347 gnd.n1346 9.3005
R18395 gnd.n1471 gnd.n1470 9.3005
R18396 gnd.n1472 gnd.n1345 9.3005
R18397 gnd.n1474 gnd.n1473 9.3005
R18398 gnd.n1335 gnd.n1334 9.3005
R18399 gnd.n1487 gnd.n1486 9.3005
R18400 gnd.n1488 gnd.n1333 9.3005
R18401 gnd.n1520 gnd.n1489 9.3005
R18402 gnd.n1519 gnd.n1490 9.3005
R18403 gnd.n1518 gnd.n1491 9.3005
R18404 gnd.n1517 gnd.n1492 9.3005
R18405 gnd.n1514 gnd.n1493 9.3005
R18406 gnd.n1513 gnd.n1494 9.3005
R18407 gnd.n1512 gnd.n1495 9.3005
R18408 gnd.n1510 gnd.n1496 9.3005
R18409 gnd.n1509 gnd.n1497 9.3005
R18410 gnd.n1506 gnd.n1498 9.3005
R18411 gnd.n1505 gnd.n1499 9.3005
R18412 gnd.n1504 gnd.n1500 9.3005
R18413 gnd.n1502 gnd.n1501 9.3005
R18414 gnd.n1201 gnd.n1200 9.3005
R18415 gnd.n1618 gnd.n1617 9.3005
R18416 gnd.n1619 gnd.n1199 9.3005
R18417 gnd.n1623 gnd.n1620 9.3005
R18418 gnd.n1622 gnd.n1621 9.3005
R18419 gnd.n1123 gnd.n1122 9.3005
R18420 gnd.n1698 gnd.n1697 9.3005
R18421 gnd.n1455 gnd.n1356 9.3005
R18422 gnd.n1358 gnd.n1357 9.3005
R18423 gnd.n1402 gnd.n1400 9.3005
R18424 gnd.n1403 gnd.n1399 9.3005
R18425 gnd.n1406 gnd.n1395 9.3005
R18426 gnd.n1407 gnd.n1394 9.3005
R18427 gnd.n1410 gnd.n1393 9.3005
R18428 gnd.n1411 gnd.n1392 9.3005
R18429 gnd.n1414 gnd.n1391 9.3005
R18430 gnd.n1415 gnd.n1390 9.3005
R18431 gnd.n1418 gnd.n1389 9.3005
R18432 gnd.n1419 gnd.n1388 9.3005
R18433 gnd.n1422 gnd.n1387 9.3005
R18434 gnd.n1423 gnd.n1386 9.3005
R18435 gnd.n1426 gnd.n1385 9.3005
R18436 gnd.n1427 gnd.n1384 9.3005
R18437 gnd.n1430 gnd.n1383 9.3005
R18438 gnd.n1431 gnd.n1382 9.3005
R18439 gnd.n1434 gnd.n1381 9.3005
R18440 gnd.n1435 gnd.n1380 9.3005
R18441 gnd.n1438 gnd.n1379 9.3005
R18442 gnd.n1439 gnd.n1378 9.3005
R18443 gnd.n1442 gnd.n1377 9.3005
R18444 gnd.n1444 gnd.n1376 9.3005
R18445 gnd.n1445 gnd.n1375 9.3005
R18446 gnd.n1446 gnd.n1374 9.3005
R18447 gnd.n1447 gnd.n1373 9.3005
R18448 gnd.n1454 gnd.n1453 9.3005
R18449 gnd.n1463 gnd.n1462 9.3005
R18450 gnd.n1464 gnd.n1350 9.3005
R18451 gnd.n1466 gnd.n1465 9.3005
R18452 gnd.n1341 gnd.n1340 9.3005
R18453 gnd.n1479 gnd.n1478 9.3005
R18454 gnd.n1480 gnd.n1339 9.3005
R18455 gnd.n1482 gnd.n1481 9.3005
R18456 gnd.n1328 gnd.n1327 9.3005
R18457 gnd.n1525 gnd.n1524 9.3005
R18458 gnd.n1526 gnd.n1282 9.3005
R18459 gnd.n1530 gnd.n1528 9.3005
R18460 gnd.n1529 gnd.n1261 9.3005
R18461 gnd.n1548 gnd.n1260 9.3005
R18462 gnd.n1551 gnd.n1550 9.3005
R18463 gnd.n1254 gnd.n1253 9.3005
R18464 gnd.n1562 gnd.n1560 9.3005
R18465 gnd.n1561 gnd.n1235 9.3005
R18466 gnd.n1579 gnd.n1234 9.3005
R18467 gnd.n1582 gnd.n1581 9.3005
R18468 gnd.n1229 gnd.n1224 9.3005
R18469 gnd.n1592 gnd.n1591 9.3005
R18470 gnd.n1227 gnd.n1207 9.3005
R18471 gnd.n1613 gnd.n1208 9.3005
R18472 gnd.n1612 gnd.n1611 9.3005
R18473 gnd.n1210 gnd.n1186 9.3005
R18474 gnd.n1644 gnd.n1643 9.3005
R18475 gnd.n1646 gnd.n1131 9.3005
R18476 gnd.n1693 gnd.n1132 9.3005
R18477 gnd.n1692 gnd.n1133 9.3005
R18478 gnd.n1691 gnd.n1134 9.3005
R18479 gnd.n1657 gnd.n1135 9.3005
R18480 gnd.n1659 gnd.n1153 9.3005
R18481 gnd.n1679 gnd.n1154 9.3005
R18482 gnd.n1678 gnd.n1155 9.3005
R18483 gnd.n1677 gnd.n1156 9.3005
R18484 gnd.n1668 gnd.n1157 9.3005
R18485 gnd.n1669 gnd.n1056 9.3005
R18486 gnd.n1735 gnd.n1734 9.3005
R18487 gnd.n1736 gnd.n1049 9.3005
R18488 gnd.n1746 gnd.n1745 9.3005
R18489 gnd.n1748 gnd.n1045 9.3005
R18490 gnd.n1758 gnd.n1046 9.3005
R18491 gnd.n1757 gnd.n1756 9.3005
R18492 gnd.n1754 gnd.n1024 9.3005
R18493 gnd.n1780 gnd.n1025 9.3005
R18494 gnd.n1779 gnd.n1778 9.3005
R18495 gnd.n1027 gnd.n1002 9.3005
R18496 gnd.n1822 gnd.n1821 9.3005
R18497 gnd.n1823 gnd.n995 9.3005
R18498 gnd.n1833 gnd.n1832 9.3005
R18499 gnd.n1835 gnd.n991 9.3005
R18500 gnd.n1845 gnd.n992 9.3005
R18501 gnd.n1844 gnd.n1843 9.3005
R18502 gnd.n1841 gnd.n970 9.3005
R18503 gnd.n1867 gnd.n971 9.3005
R18504 gnd.n1866 gnd.n1865 9.3005
R18505 gnd.n973 gnd.n948 9.3005
R18506 gnd.n1911 gnd.n1910 9.3005
R18507 gnd.n1912 gnd.n941 9.3005
R18508 gnd.n1922 gnd.n1921 9.3005
R18509 gnd.n2180 gnd.n937 9.3005
R18510 gnd.n2188 gnd.n938 9.3005
R18511 gnd.n2187 gnd.n2186 9.3005
R18512 gnd.n919 gnd.n918 9.3005
R18513 gnd.n2211 gnd.n2210 9.3005
R18514 gnd.n1352 gnd.n1351 9.3005
R18515 gnd.n6404 gnd.n672 9.3005
R18516 gnd.n6406 gnd.n6405 9.3005
R18517 gnd.n668 gnd.n667 9.3005
R18518 gnd.n6413 gnd.n6412 9.3005
R18519 gnd.n6414 gnd.n666 9.3005
R18520 gnd.n6416 gnd.n6415 9.3005
R18521 gnd.n662 gnd.n661 9.3005
R18522 gnd.n6423 gnd.n6422 9.3005
R18523 gnd.n6424 gnd.n660 9.3005
R18524 gnd.n6426 gnd.n6425 9.3005
R18525 gnd.n656 gnd.n655 9.3005
R18526 gnd.n6433 gnd.n6432 9.3005
R18527 gnd.n6434 gnd.n654 9.3005
R18528 gnd.n6436 gnd.n6435 9.3005
R18529 gnd.n650 gnd.n649 9.3005
R18530 gnd.n6443 gnd.n6442 9.3005
R18531 gnd.n6444 gnd.n648 9.3005
R18532 gnd.n6446 gnd.n6445 9.3005
R18533 gnd.n644 gnd.n643 9.3005
R18534 gnd.n6453 gnd.n6452 9.3005
R18535 gnd.n6454 gnd.n642 9.3005
R18536 gnd.n6456 gnd.n6455 9.3005
R18537 gnd.n638 gnd.n637 9.3005
R18538 gnd.n6463 gnd.n6462 9.3005
R18539 gnd.n6464 gnd.n636 9.3005
R18540 gnd.n6466 gnd.n6465 9.3005
R18541 gnd.n632 gnd.n631 9.3005
R18542 gnd.n6473 gnd.n6472 9.3005
R18543 gnd.n6474 gnd.n630 9.3005
R18544 gnd.n6476 gnd.n6475 9.3005
R18545 gnd.n626 gnd.n625 9.3005
R18546 gnd.n6483 gnd.n6482 9.3005
R18547 gnd.n6484 gnd.n624 9.3005
R18548 gnd.n6486 gnd.n6485 9.3005
R18549 gnd.n620 gnd.n619 9.3005
R18550 gnd.n6493 gnd.n6492 9.3005
R18551 gnd.n6494 gnd.n618 9.3005
R18552 gnd.n6496 gnd.n6495 9.3005
R18553 gnd.n614 gnd.n613 9.3005
R18554 gnd.n6503 gnd.n6502 9.3005
R18555 gnd.n6504 gnd.n612 9.3005
R18556 gnd.n6506 gnd.n6505 9.3005
R18557 gnd.n608 gnd.n607 9.3005
R18558 gnd.n6513 gnd.n6512 9.3005
R18559 gnd.n6514 gnd.n606 9.3005
R18560 gnd.n6516 gnd.n6515 9.3005
R18561 gnd.n602 gnd.n601 9.3005
R18562 gnd.n6523 gnd.n6522 9.3005
R18563 gnd.n6524 gnd.n600 9.3005
R18564 gnd.n6526 gnd.n6525 9.3005
R18565 gnd.n596 gnd.n595 9.3005
R18566 gnd.n6533 gnd.n6532 9.3005
R18567 gnd.n6534 gnd.n594 9.3005
R18568 gnd.n6536 gnd.n6535 9.3005
R18569 gnd.n590 gnd.n589 9.3005
R18570 gnd.n6543 gnd.n6542 9.3005
R18571 gnd.n6544 gnd.n588 9.3005
R18572 gnd.n6546 gnd.n6545 9.3005
R18573 gnd.n584 gnd.n583 9.3005
R18574 gnd.n6553 gnd.n6552 9.3005
R18575 gnd.n6554 gnd.n582 9.3005
R18576 gnd.n6556 gnd.n6555 9.3005
R18577 gnd.n578 gnd.n577 9.3005
R18578 gnd.n6563 gnd.n6562 9.3005
R18579 gnd.n6564 gnd.n576 9.3005
R18580 gnd.n6566 gnd.n6565 9.3005
R18581 gnd.n572 gnd.n571 9.3005
R18582 gnd.n6573 gnd.n6572 9.3005
R18583 gnd.n6574 gnd.n570 9.3005
R18584 gnd.n6576 gnd.n6575 9.3005
R18585 gnd.n566 gnd.n565 9.3005
R18586 gnd.n6583 gnd.n6582 9.3005
R18587 gnd.n6584 gnd.n564 9.3005
R18588 gnd.n6586 gnd.n6585 9.3005
R18589 gnd.n560 gnd.n559 9.3005
R18590 gnd.n6593 gnd.n6592 9.3005
R18591 gnd.n6594 gnd.n558 9.3005
R18592 gnd.n6596 gnd.n6595 9.3005
R18593 gnd.n554 gnd.n553 9.3005
R18594 gnd.n6603 gnd.n6602 9.3005
R18595 gnd.n6604 gnd.n552 9.3005
R18596 gnd.n6606 gnd.n6605 9.3005
R18597 gnd.n548 gnd.n547 9.3005
R18598 gnd.n6613 gnd.n6612 9.3005
R18599 gnd.n6614 gnd.n546 9.3005
R18600 gnd.n6616 gnd.n6615 9.3005
R18601 gnd.n542 gnd.n541 9.3005
R18602 gnd.n6623 gnd.n6622 9.3005
R18603 gnd.n6624 gnd.n540 9.3005
R18604 gnd.n6626 gnd.n6625 9.3005
R18605 gnd.n536 gnd.n535 9.3005
R18606 gnd.n6633 gnd.n6632 9.3005
R18607 gnd.n6634 gnd.n534 9.3005
R18608 gnd.n6636 gnd.n6635 9.3005
R18609 gnd.n530 gnd.n529 9.3005
R18610 gnd.n6643 gnd.n6642 9.3005
R18611 gnd.n6644 gnd.n528 9.3005
R18612 gnd.n6646 gnd.n6645 9.3005
R18613 gnd.n524 gnd.n523 9.3005
R18614 gnd.n6653 gnd.n6652 9.3005
R18615 gnd.n6654 gnd.n522 9.3005
R18616 gnd.n6656 gnd.n6655 9.3005
R18617 gnd.n518 gnd.n517 9.3005
R18618 gnd.n6663 gnd.n6662 9.3005
R18619 gnd.n6664 gnd.n516 9.3005
R18620 gnd.n6666 gnd.n6665 9.3005
R18621 gnd.n512 gnd.n511 9.3005
R18622 gnd.n6673 gnd.n6672 9.3005
R18623 gnd.n6674 gnd.n510 9.3005
R18624 gnd.n6676 gnd.n6675 9.3005
R18625 gnd.n506 gnd.n505 9.3005
R18626 gnd.n6683 gnd.n6682 9.3005
R18627 gnd.n6684 gnd.n504 9.3005
R18628 gnd.n6686 gnd.n6685 9.3005
R18629 gnd.n500 gnd.n499 9.3005
R18630 gnd.n6693 gnd.n6692 9.3005
R18631 gnd.n6694 gnd.n498 9.3005
R18632 gnd.n6696 gnd.n6695 9.3005
R18633 gnd.n494 gnd.n493 9.3005
R18634 gnd.n6703 gnd.n6702 9.3005
R18635 gnd.n6704 gnd.n492 9.3005
R18636 gnd.n6706 gnd.n6705 9.3005
R18637 gnd.n488 gnd.n487 9.3005
R18638 gnd.n6713 gnd.n6712 9.3005
R18639 gnd.n6714 gnd.n486 9.3005
R18640 gnd.n6716 gnd.n6715 9.3005
R18641 gnd.n482 gnd.n481 9.3005
R18642 gnd.n6723 gnd.n6722 9.3005
R18643 gnd.n6724 gnd.n480 9.3005
R18644 gnd.n6726 gnd.n6725 9.3005
R18645 gnd.n476 gnd.n475 9.3005
R18646 gnd.n6733 gnd.n6732 9.3005
R18647 gnd.n6734 gnd.n474 9.3005
R18648 gnd.n6736 gnd.n6735 9.3005
R18649 gnd.n470 gnd.n469 9.3005
R18650 gnd.n6743 gnd.n6742 9.3005
R18651 gnd.n6744 gnd.n468 9.3005
R18652 gnd.n6746 gnd.n6745 9.3005
R18653 gnd.n464 gnd.n463 9.3005
R18654 gnd.n6753 gnd.n6752 9.3005
R18655 gnd.n6754 gnd.n462 9.3005
R18656 gnd.n6756 gnd.n6755 9.3005
R18657 gnd.n458 gnd.n457 9.3005
R18658 gnd.n6763 gnd.n6762 9.3005
R18659 gnd.n6764 gnd.n456 9.3005
R18660 gnd.n6766 gnd.n6765 9.3005
R18661 gnd.n452 gnd.n451 9.3005
R18662 gnd.n6773 gnd.n6772 9.3005
R18663 gnd.n6774 gnd.n450 9.3005
R18664 gnd.n6776 gnd.n6775 9.3005
R18665 gnd.n446 gnd.n445 9.3005
R18666 gnd.n6783 gnd.n6782 9.3005
R18667 gnd.n6784 gnd.n444 9.3005
R18668 gnd.n6786 gnd.n6785 9.3005
R18669 gnd.n440 gnd.n439 9.3005
R18670 gnd.n6793 gnd.n6792 9.3005
R18671 gnd.n6794 gnd.n438 9.3005
R18672 gnd.n6796 gnd.n6795 9.3005
R18673 gnd.n434 gnd.n433 9.3005
R18674 gnd.n6803 gnd.n6802 9.3005
R18675 gnd.n6804 gnd.n432 9.3005
R18676 gnd.n6806 gnd.n6805 9.3005
R18677 gnd.n428 gnd.n427 9.3005
R18678 gnd.n6813 gnd.n6812 9.3005
R18679 gnd.n6814 gnd.n426 9.3005
R18680 gnd.n6816 gnd.n6815 9.3005
R18681 gnd.n422 gnd.n421 9.3005
R18682 gnd.n6823 gnd.n6822 9.3005
R18683 gnd.n6824 gnd.n420 9.3005
R18684 gnd.n6826 gnd.n6825 9.3005
R18685 gnd.n416 gnd.n415 9.3005
R18686 gnd.n6833 gnd.n6832 9.3005
R18687 gnd.n6834 gnd.n414 9.3005
R18688 gnd.n6836 gnd.n6835 9.3005
R18689 gnd.n410 gnd.n409 9.3005
R18690 gnd.n6843 gnd.n6842 9.3005
R18691 gnd.n6844 gnd.n408 9.3005
R18692 gnd.n6846 gnd.n6845 9.3005
R18693 gnd.n404 gnd.n403 9.3005
R18694 gnd.n6853 gnd.n6852 9.3005
R18695 gnd.n6854 gnd.n402 9.3005
R18696 gnd.n6856 gnd.n6855 9.3005
R18697 gnd.n398 gnd.n397 9.3005
R18698 gnd.n6863 gnd.n6862 9.3005
R18699 gnd.n6864 gnd.n396 9.3005
R18700 gnd.n6866 gnd.n6865 9.3005
R18701 gnd.n392 gnd.n391 9.3005
R18702 gnd.n6873 gnd.n6872 9.3005
R18703 gnd.n6874 gnd.n390 9.3005
R18704 gnd.n6876 gnd.n6875 9.3005
R18705 gnd.n386 gnd.n385 9.3005
R18706 gnd.n6883 gnd.n6882 9.3005
R18707 gnd.n6884 gnd.n384 9.3005
R18708 gnd.n6887 gnd.n6885 9.3005
R18709 gnd.n6886 gnd.n380 9.3005
R18710 gnd.n6895 gnd.n379 9.3005
R18711 gnd.n6897 gnd.n6896 9.3005
R18712 gnd.n375 gnd.n374 9.3005
R18713 gnd.n6904 gnd.n6903 9.3005
R18714 gnd.n6905 gnd.n373 9.3005
R18715 gnd.n6907 gnd.n6906 9.3005
R18716 gnd.n369 gnd.n368 9.3005
R18717 gnd.n6914 gnd.n6913 9.3005
R18718 gnd.n6915 gnd.n367 9.3005
R18719 gnd.n6917 gnd.n6916 9.3005
R18720 gnd.n363 gnd.n362 9.3005
R18721 gnd.n6924 gnd.n6923 9.3005
R18722 gnd.n6925 gnd.n361 9.3005
R18723 gnd.n6927 gnd.n6926 9.3005
R18724 gnd.n357 gnd.n356 9.3005
R18725 gnd.n6934 gnd.n6933 9.3005
R18726 gnd.n6935 gnd.n355 9.3005
R18727 gnd.n6937 gnd.n6936 9.3005
R18728 gnd.n351 gnd.n350 9.3005
R18729 gnd.n6944 gnd.n6943 9.3005
R18730 gnd.n6945 gnd.n349 9.3005
R18731 gnd.n6947 gnd.n6946 9.3005
R18732 gnd.n345 gnd.n344 9.3005
R18733 gnd.n6954 gnd.n6953 9.3005
R18734 gnd.n6955 gnd.n343 9.3005
R18735 gnd.n6957 gnd.n6956 9.3005
R18736 gnd.n339 gnd.n338 9.3005
R18737 gnd.n6964 gnd.n6963 9.3005
R18738 gnd.n6965 gnd.n337 9.3005
R18739 gnd.n6967 gnd.n6966 9.3005
R18740 gnd.n333 gnd.n332 9.3005
R18741 gnd.n6974 gnd.n6973 9.3005
R18742 gnd.n6975 gnd.n331 9.3005
R18743 gnd.n6977 gnd.n6976 9.3005
R18744 gnd.n327 gnd.n326 9.3005
R18745 gnd.n6984 gnd.n6983 9.3005
R18746 gnd.n6985 gnd.n325 9.3005
R18747 gnd.n6987 gnd.n6986 9.3005
R18748 gnd.n321 gnd.n320 9.3005
R18749 gnd.n6994 gnd.n6993 9.3005
R18750 gnd.n6995 gnd.n319 9.3005
R18751 gnd.n6997 gnd.n6996 9.3005
R18752 gnd.n315 gnd.n314 9.3005
R18753 gnd.n7004 gnd.n7003 9.3005
R18754 gnd.n7005 gnd.n313 9.3005
R18755 gnd.n7007 gnd.n7006 9.3005
R18756 gnd.n309 gnd.n308 9.3005
R18757 gnd.n7014 gnd.n7013 9.3005
R18758 gnd.n7015 gnd.n307 9.3005
R18759 gnd.n7017 gnd.n7016 9.3005
R18760 gnd.n303 gnd.n302 9.3005
R18761 gnd.n7024 gnd.n7023 9.3005
R18762 gnd.n7025 gnd.n301 9.3005
R18763 gnd.n7027 gnd.n7026 9.3005
R18764 gnd.n297 gnd.n296 9.3005
R18765 gnd.n7034 gnd.n7033 9.3005
R18766 gnd.n7035 gnd.n295 9.3005
R18767 gnd.n7037 gnd.n7036 9.3005
R18768 gnd.n291 gnd.n290 9.3005
R18769 gnd.n7044 gnd.n7043 9.3005
R18770 gnd.n7045 gnd.n289 9.3005
R18771 gnd.n7047 gnd.n7046 9.3005
R18772 gnd.n285 gnd.n284 9.3005
R18773 gnd.n7054 gnd.n7053 9.3005
R18774 gnd.n7055 gnd.n283 9.3005
R18775 gnd.n7057 gnd.n7056 9.3005
R18776 gnd.n279 gnd.n278 9.3005
R18777 gnd.n7064 gnd.n7063 9.3005
R18778 gnd.n7065 gnd.n277 9.3005
R18779 gnd.n7067 gnd.n7066 9.3005
R18780 gnd.n273 gnd.n272 9.3005
R18781 gnd.n7074 gnd.n7073 9.3005
R18782 gnd.n7075 gnd.n271 9.3005
R18783 gnd.n7077 gnd.n7076 9.3005
R18784 gnd.n267 gnd.n266 9.3005
R18785 gnd.n7084 gnd.n7083 9.3005
R18786 gnd.n7085 gnd.n265 9.3005
R18787 gnd.n7087 gnd.n7086 9.3005
R18788 gnd.n261 gnd.n260 9.3005
R18789 gnd.n7094 gnd.n7093 9.3005
R18790 gnd.n7095 gnd.n259 9.3005
R18791 gnd.n7097 gnd.n7096 9.3005
R18792 gnd.n255 gnd.n254 9.3005
R18793 gnd.n7104 gnd.n7103 9.3005
R18794 gnd.n6894 gnd.n6893 9.3005
R18795 gnd.n7406 gnd.n7405 9.3005
R18796 gnd.n7404 gnd.n65 9.3005
R18797 gnd.n5605 gnd.n67 9.3005
R18798 gnd.n5608 gnd.n5607 9.3005
R18799 gnd.n5606 gnd.n5433 9.3005
R18800 gnd.n5717 gnd.n5434 9.3005
R18801 gnd.n5716 gnd.n5435 9.3005
R18802 gnd.n5715 gnd.n5436 9.3005
R18803 gnd.n5618 gnd.n5437 9.3005
R18804 gnd.n5705 gnd.n5619 9.3005
R18805 gnd.n5704 gnd.n5620 9.3005
R18806 gnd.n5703 gnd.n5621 9.3005
R18807 gnd.n5625 gnd.n5622 9.3005
R18808 gnd.n5646 gnd.n5626 9.3005
R18809 gnd.n5645 gnd.n5627 9.3005
R18810 gnd.n5644 gnd.n5628 9.3005
R18811 gnd.n5631 gnd.n5629 9.3005
R18812 gnd.n5634 gnd.n5633 9.3005
R18813 gnd.n5632 gnd.n175 9.3005
R18814 gnd.n7337 gnd.n176 9.3005
R18815 gnd.n7336 gnd.n7335 9.3005
R18816 gnd.n202 gnd.n198 9.3005
R18817 gnd.n206 gnd.n205 9.3005
R18818 gnd.n207 gnd.n197 9.3005
R18819 gnd.n209 gnd.n208 9.3005
R18820 gnd.n212 gnd.n196 9.3005
R18821 gnd.n216 gnd.n215 9.3005
R18822 gnd.n217 gnd.n195 9.3005
R18823 gnd.n219 gnd.n218 9.3005
R18824 gnd.n222 gnd.n194 9.3005
R18825 gnd.n226 gnd.n225 9.3005
R18826 gnd.n227 gnd.n193 9.3005
R18827 gnd.n229 gnd.n228 9.3005
R18828 gnd.n232 gnd.n192 9.3005
R18829 gnd.n235 gnd.n234 9.3005
R18830 gnd.n236 gnd.n191 9.3005
R18831 gnd.n238 gnd.n237 9.3005
R18832 gnd.n180 gnd.n177 9.3005
R18833 gnd.n7334 gnd.n7333 9.3005
R18834 gnd.n200 gnd.n199 9.3005
R18835 gnd.n7151 gnd.n7148 9.3005
R18836 gnd.n7327 gnd.n7152 9.3005
R18837 gnd.n7326 gnd.n7153 9.3005
R18838 gnd.n7325 gnd.n7154 9.3005
R18839 gnd.n7322 gnd.n7155 9.3005
R18840 gnd.n7321 gnd.n7156 9.3005
R18841 gnd.n7318 gnd.n7157 9.3005
R18842 gnd.n7317 gnd.n7158 9.3005
R18843 gnd.n7314 gnd.n7159 9.3005
R18844 gnd.n7313 gnd.n7160 9.3005
R18845 gnd.n7310 gnd.n7161 9.3005
R18846 gnd.n7309 gnd.n7162 9.3005
R18847 gnd.n7306 gnd.n7163 9.3005
R18848 gnd.n7305 gnd.n7164 9.3005
R18849 gnd.n7302 gnd.n7165 9.3005
R18850 gnd.n7301 gnd.n7166 9.3005
R18851 gnd.n7298 gnd.n7167 9.3005
R18852 gnd.n7294 gnd.n7168 9.3005
R18853 gnd.n7291 gnd.n7169 9.3005
R18854 gnd.n7290 gnd.n7170 9.3005
R18855 gnd.n7287 gnd.n7171 9.3005
R18856 gnd.n7286 gnd.n7172 9.3005
R18857 gnd.n7283 gnd.n7173 9.3005
R18858 gnd.n7282 gnd.n7174 9.3005
R18859 gnd.n7279 gnd.n7175 9.3005
R18860 gnd.n7278 gnd.n7176 9.3005
R18861 gnd.n7275 gnd.n7177 9.3005
R18862 gnd.n7274 gnd.n7178 9.3005
R18863 gnd.n7271 gnd.n7179 9.3005
R18864 gnd.n7270 gnd.n7180 9.3005
R18865 gnd.n7267 gnd.n7181 9.3005
R18866 gnd.n7266 gnd.n7182 9.3005
R18867 gnd.n7263 gnd.n7183 9.3005
R18868 gnd.n7262 gnd.n7184 9.3005
R18869 gnd.n7259 gnd.n7185 9.3005
R18870 gnd.n7258 gnd.n7186 9.3005
R18871 gnd.n7255 gnd.n7254 9.3005
R18872 gnd.n7253 gnd.n7187 9.3005
R18873 gnd.n7252 gnd.n7251 9.3005
R18874 gnd.n7248 gnd.n7190 9.3005
R18875 gnd.n7245 gnd.n7191 9.3005
R18876 gnd.n7244 gnd.n7192 9.3005
R18877 gnd.n7241 gnd.n7193 9.3005
R18878 gnd.n7240 gnd.n7194 9.3005
R18879 gnd.n7237 gnd.n7195 9.3005
R18880 gnd.n7236 gnd.n7196 9.3005
R18881 gnd.n7233 gnd.n7197 9.3005
R18882 gnd.n7232 gnd.n7198 9.3005
R18883 gnd.n7229 gnd.n7199 9.3005
R18884 gnd.n7228 gnd.n7200 9.3005
R18885 gnd.n7225 gnd.n7201 9.3005
R18886 gnd.n7224 gnd.n7202 9.3005
R18887 gnd.n7221 gnd.n7203 9.3005
R18888 gnd.n7220 gnd.n7204 9.3005
R18889 gnd.n7217 gnd.n7205 9.3005
R18890 gnd.n7216 gnd.n7206 9.3005
R18891 gnd.n7213 gnd.n7212 9.3005
R18892 gnd.n7211 gnd.n7208 9.3005
R18893 gnd.n7150 gnd.n7149 9.3005
R18894 gnd.n5319 gnd.n2816 9.3005
R18895 gnd.n5492 gnd.n5335 9.3005
R18896 gnd.n5796 gnd.n5336 9.3005
R18897 gnd.n5795 gnd.n5337 9.3005
R18898 gnd.n5794 gnd.n5338 9.3005
R18899 gnd.n5507 gnd.n5339 9.3005
R18900 gnd.n5784 gnd.n5356 9.3005
R18901 gnd.n5783 gnd.n5357 9.3005
R18902 gnd.n5782 gnd.n5358 9.3005
R18903 gnd.n5514 gnd.n5359 9.3005
R18904 gnd.n5772 gnd.n5376 9.3005
R18905 gnd.n5771 gnd.n5377 9.3005
R18906 gnd.n5770 gnd.n5378 9.3005
R18907 gnd.n5520 gnd.n5379 9.3005
R18908 gnd.n5760 gnd.n5395 9.3005
R18909 gnd.n5759 gnd.n5396 9.3005
R18910 gnd.n5758 gnd.n5397 9.3005
R18911 gnd.n5585 gnd.n5398 9.3005
R18912 gnd.n5588 gnd.n5587 9.3005
R18913 gnd.n5589 gnd.n5420 9.3005
R18914 gnd.n5734 gnd.n5421 9.3005
R18915 gnd.n5733 gnd.n5422 9.3005
R18916 gnd.n5732 gnd.n5423 9.3005
R18917 gnd.n5731 gnd.n5424 9.3005
R18918 gnd.n5604 gnd.n91 9.3005
R18919 gnd.n7392 gnd.n92 9.3005
R18920 gnd.n7391 gnd.n93 9.3005
R18921 gnd.n7390 gnd.n94 9.3005
R18922 gnd.n5616 gnd.n95 9.3005
R18923 gnd.n7380 gnd.n111 9.3005
R18924 gnd.n7379 gnd.n112 9.3005
R18925 gnd.n7378 gnd.n113 9.3005
R18926 gnd.n5623 gnd.n114 9.3005
R18927 gnd.n7368 gnd.n132 9.3005
R18928 gnd.n7367 gnd.n133 9.3005
R18929 gnd.n7366 gnd.n134 9.3005
R18930 gnd.n5630 gnd.n135 9.3005
R18931 gnd.n7356 gnd.n152 9.3005
R18932 gnd.n7355 gnd.n153 9.3005
R18933 gnd.n7354 gnd.n154 9.3005
R18934 gnd.n172 gnd.n155 9.3005
R18935 gnd.n7344 gnd.n7343 9.3005
R18936 gnd.n5810 gnd.n2815 9.3005
R18937 gnd.n2817 gnd.n2816 9.3005
R18938 gnd.n5493 gnd.n5492 9.3005
R18939 gnd.n5486 gnd.n5336 9.3005
R18940 gnd.n5505 gnd.n5337 9.3005
R18941 gnd.n5506 gnd.n5338 9.3005
R18942 gnd.n5508 gnd.n5507 9.3005
R18943 gnd.n5509 gnd.n5356 9.3005
R18944 gnd.n5512 gnd.n5357 9.3005
R18945 gnd.n5513 gnd.n5358 9.3005
R18946 gnd.n5518 gnd.n5514 9.3005
R18947 gnd.n5519 gnd.n5376 9.3005
R18948 gnd.n5523 gnd.n5377 9.3005
R18949 gnd.n5522 gnd.n5378 9.3005
R18950 gnd.n5521 gnd.n5520 9.3005
R18951 gnd.n5439 gnd.n5395 9.3005
R18952 gnd.n5582 gnd.n5396 9.3005
R18953 gnd.n5583 gnd.n5397 9.3005
R18954 gnd.n5585 gnd.n5584 9.3005
R18955 gnd.n5588 gnd.n5438 9.3005
R18956 gnd.n5592 gnd.n5589 9.3005
R18957 gnd.n5593 gnd.n5421 9.3005
R18958 gnd.n5601 gnd.n5422 9.3005
R18959 gnd.n5602 gnd.n5423 9.3005
R18960 gnd.n5603 gnd.n5424 9.3005
R18961 gnd.n5612 gnd.n5604 9.3005
R18962 gnd.n5613 gnd.n92 9.3005
R18963 gnd.n5614 gnd.n93 9.3005
R18964 gnd.n5615 gnd.n94 9.3005
R18965 gnd.n5711 gnd.n5616 9.3005
R18966 gnd.n5710 gnd.n111 9.3005
R18967 gnd.n5709 gnd.n112 9.3005
R18968 gnd.n5617 gnd.n113 9.3005
R18969 gnd.n5699 gnd.n5623 9.3005
R18970 gnd.n5698 gnd.n132 9.3005
R18971 gnd.n5697 gnd.n133 9.3005
R18972 gnd.n5624 gnd.n134 9.3005
R18973 gnd.n5640 gnd.n5630 9.3005
R18974 gnd.n5639 gnd.n152 9.3005
R18975 gnd.n5638 gnd.n153 9.3005
R18976 gnd.n174 gnd.n154 9.3005
R18977 gnd.n7341 gnd.n172 9.3005
R18978 gnd.n7343 gnd.n7342 9.3005
R18979 gnd.n5810 gnd.n5809 9.3005
R18980 gnd.n5814 gnd.n5813 9.3005
R18981 gnd.n5817 gnd.n2810 9.3005
R18982 gnd.n5818 gnd.n2809 9.3005
R18983 gnd.n5821 gnd.n2808 9.3005
R18984 gnd.n5822 gnd.n2807 9.3005
R18985 gnd.n5825 gnd.n2806 9.3005
R18986 gnd.n5826 gnd.n2805 9.3005
R18987 gnd.n5829 gnd.n2804 9.3005
R18988 gnd.n5830 gnd.n2803 9.3005
R18989 gnd.n5833 gnd.n2802 9.3005
R18990 gnd.n5834 gnd.n2801 9.3005
R18991 gnd.n5837 gnd.n2800 9.3005
R18992 gnd.n5838 gnd.n2799 9.3005
R18993 gnd.n5841 gnd.n2798 9.3005
R18994 gnd.n5842 gnd.n2797 9.3005
R18995 gnd.n5845 gnd.n2796 9.3005
R18996 gnd.n5846 gnd.n2795 9.3005
R18997 gnd.n5849 gnd.n2794 9.3005
R18998 gnd.n5850 gnd.n2793 9.3005
R18999 gnd.n5853 gnd.n2792 9.3005
R19000 gnd.n5857 gnd.n2788 9.3005
R19001 gnd.n5858 gnd.n2787 9.3005
R19002 gnd.n5861 gnd.n2786 9.3005
R19003 gnd.n5862 gnd.n2785 9.3005
R19004 gnd.n5865 gnd.n2784 9.3005
R19005 gnd.n5866 gnd.n2783 9.3005
R19006 gnd.n5869 gnd.n2782 9.3005
R19007 gnd.n5870 gnd.n2781 9.3005
R19008 gnd.n5873 gnd.n2780 9.3005
R19009 gnd.n5875 gnd.n2776 9.3005
R19010 gnd.n5878 gnd.n2775 9.3005
R19011 gnd.n5879 gnd.n2774 9.3005
R19012 gnd.n5882 gnd.n2773 9.3005
R19013 gnd.n5883 gnd.n2772 9.3005
R19014 gnd.n5886 gnd.n2771 9.3005
R19015 gnd.n5887 gnd.n2770 9.3005
R19016 gnd.n5890 gnd.n2769 9.3005
R19017 gnd.n5892 gnd.n2766 9.3005
R19018 gnd.n5895 gnd.n2765 9.3005
R19019 gnd.n5896 gnd.n2764 9.3005
R19020 gnd.n5899 gnd.n2763 9.3005
R19021 gnd.n5900 gnd.n2762 9.3005
R19022 gnd.n5903 gnd.n2761 9.3005
R19023 gnd.n5904 gnd.n2760 9.3005
R19024 gnd.n5907 gnd.n2759 9.3005
R19025 gnd.n5908 gnd.n2758 9.3005
R19026 gnd.n5911 gnd.n2757 9.3005
R19027 gnd.n5912 gnd.n2756 9.3005
R19028 gnd.n5915 gnd.n2755 9.3005
R19029 gnd.n5916 gnd.n2754 9.3005
R19030 gnd.n5919 gnd.n2753 9.3005
R19031 gnd.n5921 gnd.n2752 9.3005
R19032 gnd.n5922 gnd.n2751 9.3005
R19033 gnd.n5923 gnd.n2750 9.3005
R19034 gnd.n5924 gnd.n2749 9.3005
R19035 gnd.n5854 gnd.n2789 9.3005
R19036 gnd.n5812 gnd.n2811 9.3005
R19037 gnd.n5802 gnd.n5325 9.3005
R19038 gnd.n5801 gnd.n5326 9.3005
R19039 gnd.n5800 gnd.n5327 9.3005
R19040 gnd.n5346 gnd.n5328 9.3005
R19041 gnd.n5790 gnd.n5347 9.3005
R19042 gnd.n5789 gnd.n5348 9.3005
R19043 gnd.n5788 gnd.n5349 9.3005
R19044 gnd.n5365 gnd.n5350 9.3005
R19045 gnd.n5778 gnd.n5366 9.3005
R19046 gnd.n5777 gnd.n5367 9.3005
R19047 gnd.n5776 gnd.n5368 9.3005
R19048 gnd.n5386 gnd.n5369 9.3005
R19049 gnd.n5766 gnd.n5387 9.3005
R19050 gnd.n5765 gnd.n5388 9.3005
R19051 gnd.n5764 gnd.n77 9.3005
R19052 gnd.n82 gnd.n76 9.3005
R19053 gnd.n7386 gnd.n101 9.3005
R19054 gnd.n7385 gnd.n102 9.3005
R19055 gnd.n7384 gnd.n103 9.3005
R19056 gnd.n121 gnd.n104 9.3005
R19057 gnd.n7374 gnd.n122 9.3005
R19058 gnd.n7373 gnd.n123 9.3005
R19059 gnd.n7372 gnd.n124 9.3005
R19060 gnd.n141 gnd.n125 9.3005
R19061 gnd.n7362 gnd.n142 9.3005
R19062 gnd.n7361 gnd.n143 9.3005
R19063 gnd.n7360 gnd.n144 9.3005
R19064 gnd.n162 gnd.n145 9.3005
R19065 gnd.n7350 gnd.n163 9.3005
R19066 gnd.n7349 gnd.n164 9.3005
R19067 gnd.n7348 gnd.n165 9.3005
R19068 gnd.n5324 gnd.n5323 9.3005
R19069 gnd.n7397 gnd.n7396 9.3005
R19070 gnd.n3777 gnd.n3764 9.3005
R19071 gnd.n3776 gnd.n3771 9.3005
R19072 gnd.n3773 gnd.n3772 9.3005
R19073 gnd.n3687 gnd.n3686 9.3005
R19074 gnd.n4249 gnd.n4248 9.3005
R19075 gnd.n4250 gnd.n3685 9.3005
R19076 gnd.n4252 gnd.n4251 9.3005
R19077 gnd.n3683 gnd.n3682 9.3005
R19078 gnd.n4257 gnd.n4256 9.3005
R19079 gnd.n4258 gnd.n3681 9.3005
R19080 gnd.n4260 gnd.n4259 9.3005
R19081 gnd.n3679 gnd.n3678 9.3005
R19082 gnd.n4265 gnd.n4264 9.3005
R19083 gnd.n4266 gnd.n3677 9.3005
R19084 gnd.n4268 gnd.n4267 9.3005
R19085 gnd.n3675 gnd.n3674 9.3005
R19086 gnd.n4273 gnd.n4272 9.3005
R19087 gnd.n4274 gnd.n3673 9.3005
R19088 gnd.n4277 gnd.n4276 9.3005
R19089 gnd.n4275 gnd.n2567 9.3005
R19090 gnd.n6067 gnd.n2568 9.3005
R19091 gnd.n6066 gnd.n2569 9.3005
R19092 gnd.n6065 gnd.n2570 9.3005
R19093 gnd.n3453 gnd.n2571 9.3005
R19094 gnd.n3454 gnd.n3452 9.3005
R19095 gnd.n3456 gnd.n3455 9.3005
R19096 gnd.n3447 gnd.n3446 9.3005
R19097 gnd.n3465 gnd.n3464 9.3005
R19098 gnd.n3466 gnd.n3445 9.3005
R19099 gnd.n3468 gnd.n3467 9.3005
R19100 gnd.n3441 gnd.n3440 9.3005
R19101 gnd.n3477 gnd.n3476 9.3005
R19102 gnd.n3478 gnd.n3439 9.3005
R19103 gnd.n3482 gnd.n3479 9.3005
R19104 gnd.n3481 gnd.n3480 9.3005
R19105 gnd.n3220 gnd.n3219 9.3005
R19106 gnd.n4559 gnd.n4558 9.3005
R19107 gnd.n4560 gnd.n3218 9.3005
R19108 gnd.n4564 gnd.n4561 9.3005
R19109 gnd.n4563 gnd.n4562 9.3005
R19110 gnd.n3196 gnd.n3195 9.3005
R19111 gnd.n4597 gnd.n4596 9.3005
R19112 gnd.n4598 gnd.n3194 9.3005
R19113 gnd.n4605 gnd.n4599 9.3005
R19114 gnd.n4604 gnd.n4600 9.3005
R19115 gnd.n4603 gnd.n4601 9.3005
R19116 gnd.n3171 gnd.n3170 9.3005
R19117 gnd.n4637 gnd.n4636 9.3005
R19118 gnd.n4638 gnd.n3169 9.3005
R19119 gnd.n4642 gnd.n4639 9.3005
R19120 gnd.n4641 gnd.n4640 9.3005
R19121 gnd.n3143 gnd.n3142 9.3005
R19122 gnd.n4673 gnd.n4672 9.3005
R19123 gnd.n4674 gnd.n3141 9.3005
R19124 gnd.n4676 gnd.n4675 9.3005
R19125 gnd.n3125 gnd.n3124 9.3005
R19126 gnd.n4699 gnd.n4698 9.3005
R19127 gnd.n4700 gnd.n3123 9.3005
R19128 gnd.n4704 gnd.n4701 9.3005
R19129 gnd.n4703 gnd.n4702 9.3005
R19130 gnd.n3099 gnd.n3098 9.3005
R19131 gnd.n4755 gnd.n4754 9.3005
R19132 gnd.n4756 gnd.n3097 9.3005
R19133 gnd.n4760 gnd.n4757 9.3005
R19134 gnd.n4759 gnd.n4758 9.3005
R19135 gnd.n3074 gnd.n3073 9.3005
R19136 gnd.n4795 gnd.n4794 9.3005
R19137 gnd.n4796 gnd.n3072 9.3005
R19138 gnd.n4800 gnd.n4797 9.3005
R19139 gnd.n4799 gnd.n4798 9.3005
R19140 gnd.n3044 gnd.n3043 9.3005
R19141 gnd.n4864 gnd.n4863 9.3005
R19142 gnd.n4865 gnd.n3042 9.3005
R19143 gnd.n4869 gnd.n4866 9.3005
R19144 gnd.n4868 gnd.n4867 9.3005
R19145 gnd.n3020 gnd.n3019 9.3005
R19146 gnd.n4897 gnd.n4896 9.3005
R19147 gnd.n4898 gnd.n3018 9.3005
R19148 gnd.n4902 gnd.n4899 9.3005
R19149 gnd.n4901 gnd.n4900 9.3005
R19150 gnd.n2999 gnd.n2998 9.3005
R19151 gnd.n4951 gnd.n4950 9.3005
R19152 gnd.n4952 gnd.n2997 9.3005
R19153 gnd.n4956 gnd.n4953 9.3005
R19154 gnd.n4955 gnd.n4954 9.3005
R19155 gnd.n2974 gnd.n2973 9.3005
R19156 gnd.n4988 gnd.n4987 9.3005
R19157 gnd.n4989 gnd.n2972 9.3005
R19158 gnd.n4991 gnd.n4990 9.3005
R19159 gnd.n2883 gnd.n2882 9.3005
R19160 gnd.n5131 gnd.n5130 9.3005
R19161 gnd.n5132 gnd.n2881 9.3005
R19162 gnd.n5134 gnd.n5133 9.3005
R19163 gnd.n2870 gnd.n2869 9.3005
R19164 gnd.n5147 gnd.n5146 9.3005
R19165 gnd.n5148 gnd.n2868 9.3005
R19166 gnd.n5150 gnd.n5149 9.3005
R19167 gnd.n2857 gnd.n2856 9.3005
R19168 gnd.n5163 gnd.n5162 9.3005
R19169 gnd.n5164 gnd.n2855 9.3005
R19170 gnd.n5166 gnd.n5165 9.3005
R19171 gnd.n2843 gnd.n2842 9.3005
R19172 gnd.n5180 gnd.n5179 9.3005
R19173 gnd.n5181 gnd.n2841 9.3005
R19174 gnd.n5184 gnd.n5183 9.3005
R19175 gnd.n5182 gnd.n2701 9.3005
R19176 gnd.n5932 gnd.n2702 9.3005
R19177 gnd.n5931 gnd.n2703 9.3005
R19178 gnd.n5930 gnd.n2704 9.3005
R19179 gnd.n5460 gnd.n2705 9.3005
R19180 gnd.n5462 gnd.n5461 9.3005
R19181 gnd.n5466 gnd.n5465 9.3005
R19182 gnd.n5467 gnd.n5459 9.3005
R19183 gnd.n5469 gnd.n5468 9.3005
R19184 gnd.n5457 gnd.n5456 9.3005
R19185 gnd.n5474 gnd.n5473 9.3005
R19186 gnd.n5475 gnd.n5455 9.3005
R19187 gnd.n5477 gnd.n5476 9.3005
R19188 gnd.n5453 gnd.n5452 9.3005
R19189 gnd.n5545 gnd.n5544 9.3005
R19190 gnd.n5546 gnd.n5451 9.3005
R19191 gnd.n5548 gnd.n5547 9.3005
R19192 gnd.n5449 gnd.n5448 9.3005
R19193 gnd.n5553 gnd.n5552 9.3005
R19194 gnd.n5554 gnd.n5447 9.3005
R19195 gnd.n5561 gnd.n5555 9.3005
R19196 gnd.n5560 gnd.n5556 9.3005
R19197 gnd.n5723 gnd.n5429 9.3005
R19198 gnd.n5655 gnd.n5430 9.3005
R19199 gnd.n5657 gnd.n5656 9.3005
R19200 gnd.n5660 gnd.n5659 9.3005
R19201 gnd.n5661 gnd.n5654 9.3005
R19202 gnd.n5663 gnd.n5662 9.3005
R19203 gnd.n5652 gnd.n5651 9.3005
R19204 gnd.n5668 gnd.n5667 9.3005
R19205 gnd.n5669 gnd.n5650 9.3005
R19206 gnd.n5692 gnd.n5670 9.3005
R19207 gnd.n5691 gnd.n5671 9.3005
R19208 gnd.n5690 gnd.n5672 9.3005
R19209 gnd.n5675 gnd.n5673 9.3005
R19210 gnd.n5686 gnd.n5676 9.3005
R19211 gnd.n5685 gnd.n5677 9.3005
R19212 gnd.n5684 gnd.n5678 9.3005
R19213 gnd.n5681 gnd.n5680 9.3005
R19214 gnd.n5679 gnd.n244 9.3005
R19215 gnd.n7115 gnd.n245 9.3005
R19216 gnd.n7114 gnd.n246 9.3005
R19217 gnd.n7113 gnd.n247 9.3005
R19218 gnd.n252 gnd.n248 9.3005
R19219 gnd.n7107 gnd.n253 9.3005
R19220 gnd.n7106 gnd.n7105 9.3005
R19221 gnd.n4176 gnd.n4175 9.3005
R19222 gnd.n3850 gnd.n3847 9.3005
R19223 gnd.n3817 gnd.n3816 9.3005
R19224 gnd.n4117 gnd.n4116 9.3005
R19225 gnd.n4118 gnd.n3815 9.3005
R19226 gnd.n4120 gnd.n4119 9.3005
R19227 gnd.n3730 gnd.n3729 9.3005
R19228 gnd.n4131 gnd.n4130 9.3005
R19229 gnd.n4132 gnd.n3728 9.3005
R19230 gnd.n4134 gnd.n4133 9.3005
R19231 gnd.n3725 gnd.n3724 9.3005
R19232 gnd.n4145 gnd.n4144 9.3005
R19233 gnd.n4146 gnd.n3723 9.3005
R19234 gnd.n4148 gnd.n4147 9.3005
R19235 gnd.n3719 gnd.n3718 9.3005
R19236 gnd.n4159 gnd.n4158 9.3005
R19237 gnd.n4160 gnd.n3717 9.3005
R19238 gnd.n4162 gnd.n4161 9.3005
R19239 gnd.n3714 gnd.n3713 9.3005
R19240 gnd.n4173 gnd.n4172 9.3005
R19241 gnd.n4174 gnd.n3712 9.3005
R19242 gnd.n3852 gnd.n3851 9.3005
R19243 gnd.n3846 gnd.n3843 9.3005
R19244 gnd.n3863 gnd.n3842 9.3005
R19245 gnd.n3864 gnd.n3841 9.3005
R19246 gnd.n3865 gnd.n3840 9.3005
R19247 gnd.n3839 gnd.n3837 9.3005
R19248 gnd.n3871 gnd.n3836 9.3005
R19249 gnd.n3872 gnd.n3835 9.3005
R19250 gnd.n3873 gnd.n3834 9.3005
R19251 gnd.n3833 gnd.n3831 9.3005
R19252 gnd.n3879 gnd.n3830 9.3005
R19253 gnd.n3880 gnd.n3829 9.3005
R19254 gnd.n3881 gnd.n3828 9.3005
R19255 gnd.n3827 gnd.n3825 9.3005
R19256 gnd.n3886 gnd.n3824 9.3005
R19257 gnd.n3887 gnd.n3823 9.3005
R19258 gnd.n3821 gnd.n3820 9.3005
R19259 gnd.n3893 gnd.n3892 9.3005
R19260 gnd.n3857 gnd.n3854 9.3005
R19261 gnd.n3853 gnd.n3845 9.3005
R19262 gnd.n3362 gnd.n3360 9.3005
R19263 gnd.n4326 gnd.n4323 9.3005
R19264 gnd.n4327 gnd.n4322 9.3005
R19265 gnd.n4330 gnd.n4321 9.3005
R19266 gnd.n4331 gnd.n4320 9.3005
R19267 gnd.n4334 gnd.n4319 9.3005
R19268 gnd.n4335 gnd.n4318 9.3005
R19269 gnd.n4338 gnd.n4317 9.3005
R19270 gnd.n4340 gnd.n4314 9.3005
R19271 gnd.n4343 gnd.n4313 9.3005
R19272 gnd.n4344 gnd.n4312 9.3005
R19273 gnd.n4347 gnd.n4311 9.3005
R19274 gnd.n4348 gnd.n4310 9.3005
R19275 gnd.n4351 gnd.n4309 9.3005
R19276 gnd.n4352 gnd.n4308 9.3005
R19277 gnd.n4355 gnd.n4307 9.3005
R19278 gnd.n4356 gnd.n4306 9.3005
R19279 gnd.n4359 gnd.n4305 9.3005
R19280 gnd.n4360 gnd.n4304 9.3005
R19281 gnd.n4363 gnd.n4303 9.3005
R19282 gnd.n4364 gnd.n4302 9.3005
R19283 gnd.n4367 gnd.n4301 9.3005
R19284 gnd.n4368 gnd.n4300 9.3005
R19285 gnd.n4369 gnd.n4299 9.3005
R19286 gnd.n4298 gnd.n4295 9.3005
R19287 gnd.n4297 gnd.n4296 9.3005
R19288 gnd.n4479 gnd.n4478 9.3005
R19289 gnd.n3364 gnd.n3363 9.3005
R19290 gnd.n4375 gnd.n4373 9.3005
R19291 gnd.n4471 gnd.n4376 9.3005
R19292 gnd.n4470 gnd.n4377 9.3005
R19293 gnd.n4469 gnd.n4378 9.3005
R19294 gnd.n4382 gnd.n4379 9.3005
R19295 gnd.n4464 gnd.n4383 9.3005
R19296 gnd.n4463 gnd.n4462 9.3005
R19297 gnd.n4461 gnd.n4384 9.3005
R19298 gnd.n4460 gnd.n4459 9.3005
R19299 gnd.n4388 gnd.n4387 9.3005
R19300 gnd.n4393 gnd.n4391 9.3005
R19301 gnd.n4452 gnd.n4394 9.3005
R19302 gnd.n4451 gnd.n4395 9.3005
R19303 gnd.n4450 gnd.n4396 9.3005
R19304 gnd.n4400 gnd.n4397 9.3005
R19305 gnd.n4445 gnd.n4401 9.3005
R19306 gnd.n4444 gnd.n4402 9.3005
R19307 gnd.n4443 gnd.n4403 9.3005
R19308 gnd.n4407 gnd.n4404 9.3005
R19309 gnd.n4438 gnd.n4408 9.3005
R19310 gnd.n4437 gnd.n4409 9.3005
R19311 gnd.n4436 gnd.n4410 9.3005
R19312 gnd.n4414 gnd.n4411 9.3005
R19313 gnd.n4431 gnd.n4415 9.3005
R19314 gnd.n4430 gnd.n4416 9.3005
R19315 gnd.n4429 gnd.n4417 9.3005
R19316 gnd.n4422 gnd.n4420 9.3005
R19317 gnd.n4424 gnd.n4423 9.3005
R19318 gnd.n4480 gnd.n3359 9.3005
R19319 gnd.n4109 gnd.n2340 9.3005
R19320 gnd.n6207 gnd.n2341 9.3005
R19321 gnd.n6206 gnd.n2342 9.3005
R19322 gnd.n6205 gnd.n2343 9.3005
R19323 gnd.n3814 gnd.n2344 9.3005
R19324 gnd.n6195 gnd.n2361 9.3005
R19325 gnd.n6194 gnd.n2362 9.3005
R19326 gnd.n6193 gnd.n2363 9.3005
R19327 gnd.n3727 gnd.n2364 9.3005
R19328 gnd.n6183 gnd.n2382 9.3005
R19329 gnd.n6182 gnd.n2383 9.3005
R19330 gnd.n6181 gnd.n2384 9.3005
R19331 gnd.n3722 gnd.n2385 9.3005
R19332 gnd.n6171 gnd.n2402 9.3005
R19333 gnd.n6170 gnd.n2403 9.3005
R19334 gnd.n6169 gnd.n2404 9.3005
R19335 gnd.n3716 gnd.n2405 9.3005
R19336 gnd.n6158 gnd.n2421 9.3005
R19337 gnd.n6157 gnd.n2422 9.3005
R19338 gnd.n6156 gnd.n2423 9.3005
R19339 gnd.n3711 gnd.n2424 9.3005
R19340 gnd.n6145 gnd.n2438 9.3005
R19341 gnd.n6144 gnd.n2439 9.3005
R19342 gnd.n6143 gnd.n2440 9.3005
R19343 gnd.n3705 gnd.n2441 9.3005
R19344 gnd.n6132 gnd.n2456 9.3005
R19345 gnd.n6131 gnd.n2457 9.3005
R19346 gnd.n6130 gnd.n2458 9.3005
R19347 gnd.n3700 gnd.n2459 9.3005
R19348 gnd.n6120 gnd.n2476 9.3005
R19349 gnd.n6119 gnd.n2477 9.3005
R19350 gnd.n6118 gnd.n2478 9.3005
R19351 gnd.n4212 gnd.n2479 9.3005
R19352 gnd.n6108 gnd.n2497 9.3005
R19353 gnd.n6107 gnd.n2498 9.3005
R19354 gnd.n6106 gnd.n2499 9.3005
R19355 gnd.n4221 gnd.n2500 9.3005
R19356 gnd.n6096 gnd.n2518 9.3005
R19357 gnd.n6095 gnd.n2519 9.3005
R19358 gnd.n6094 gnd.n2520 9.3005
R19359 gnd.n2537 gnd.n2521 9.3005
R19360 gnd.n6084 gnd.n6083 9.3005
R19361 gnd.n4108 gnd.n4107 9.3005
R19362 gnd.n4110 gnd.n4109 9.3005
R19363 gnd.n4111 gnd.n2341 9.3005
R19364 gnd.n4112 gnd.n2342 9.3005
R19365 gnd.n3813 gnd.n2343 9.3005
R19366 gnd.n4124 gnd.n3814 9.3005
R19367 gnd.n4125 gnd.n2361 9.3005
R19368 gnd.n4126 gnd.n2362 9.3005
R19369 gnd.n3726 gnd.n2363 9.3005
R19370 gnd.n4138 gnd.n3727 9.3005
R19371 gnd.n4139 gnd.n2382 9.3005
R19372 gnd.n4140 gnd.n2383 9.3005
R19373 gnd.n3721 gnd.n2384 9.3005
R19374 gnd.n4152 gnd.n3722 9.3005
R19375 gnd.n4153 gnd.n2402 9.3005
R19376 gnd.n4154 gnd.n2403 9.3005
R19377 gnd.n3715 gnd.n2404 9.3005
R19378 gnd.n4166 gnd.n3716 9.3005
R19379 gnd.n4167 gnd.n2421 9.3005
R19380 gnd.n4168 gnd.n2422 9.3005
R19381 gnd.n3710 gnd.n2423 9.3005
R19382 gnd.n4180 gnd.n3711 9.3005
R19383 gnd.n4181 gnd.n2438 9.3005
R19384 gnd.n4182 gnd.n2439 9.3005
R19385 gnd.n3704 gnd.n2440 9.3005
R19386 gnd.n4194 gnd.n3705 9.3005
R19387 gnd.n4195 gnd.n2456 9.3005
R19388 gnd.n4196 gnd.n2457 9.3005
R19389 gnd.n3699 gnd.n2458 9.3005
R19390 gnd.n4208 gnd.n3700 9.3005
R19391 gnd.n4209 gnd.n2476 9.3005
R19392 gnd.n4210 gnd.n2477 9.3005
R19393 gnd.n4211 gnd.n2478 9.3005
R19394 gnd.n4215 gnd.n4212 9.3005
R19395 gnd.n4216 gnd.n2497 9.3005
R19396 gnd.n4219 gnd.n2498 9.3005
R19397 gnd.n4220 gnd.n2499 9.3005
R19398 gnd.n4224 gnd.n4221 9.3005
R19399 gnd.n4225 gnd.n2518 9.3005
R19400 gnd.n4226 gnd.n2519 9.3005
R19401 gnd.n2539 gnd.n2520 9.3005
R19402 gnd.n6081 gnd.n2537 9.3005
R19403 gnd.n6083 gnd.n6082 9.3005
R19404 gnd.n4108 gnd.n3818 9.3005
R19405 gnd.n3897 gnd.n3894 9.3005
R19406 gnd.n4095 gnd.n3898 9.3005
R19407 gnd.n4097 gnd.n4096 9.3005
R19408 gnd.n4094 gnd.n3900 9.3005
R19409 gnd.n4093 gnd.n4092 9.3005
R19410 gnd.n3902 gnd.n3901 9.3005
R19411 gnd.n4086 gnd.n4085 9.3005
R19412 gnd.n4084 gnd.n3904 9.3005
R19413 gnd.n4083 gnd.n4082 9.3005
R19414 gnd.n3906 gnd.n3905 9.3005
R19415 gnd.n4076 gnd.n4075 9.3005
R19416 gnd.n4074 gnd.n3908 9.3005
R19417 gnd.n4073 gnd.n4072 9.3005
R19418 gnd.n3910 gnd.n3909 9.3005
R19419 gnd.n4066 gnd.n4065 9.3005
R19420 gnd.n4064 gnd.n3912 9.3005
R19421 gnd.n4063 gnd.n4062 9.3005
R19422 gnd.n3914 gnd.n3913 9.3005
R19423 gnd.n4056 gnd.n4055 9.3005
R19424 gnd.n4054 gnd.n3916 9.3005
R19425 gnd.n3918 gnd.n3917 9.3005
R19426 gnd.n4044 gnd.n4043 9.3005
R19427 gnd.n4042 gnd.n3920 9.3005
R19428 gnd.n4041 gnd.n4040 9.3005
R19429 gnd.n3922 gnd.n3921 9.3005
R19430 gnd.n4034 gnd.n4033 9.3005
R19431 gnd.n4032 gnd.n3924 9.3005
R19432 gnd.n4031 gnd.n4030 9.3005
R19433 gnd.n3926 gnd.n3925 9.3005
R19434 gnd.n4024 gnd.n4023 9.3005
R19435 gnd.n4022 gnd.n3928 9.3005
R19436 gnd.n4021 gnd.n4020 9.3005
R19437 gnd.n3930 gnd.n3929 9.3005
R19438 gnd.n4014 gnd.n4013 9.3005
R19439 gnd.n4012 gnd.n3932 9.3005
R19440 gnd.n4011 gnd.n4010 9.3005
R19441 gnd.n3934 gnd.n3933 9.3005
R19442 gnd.n4004 gnd.n4003 9.3005
R19443 gnd.n4002 gnd.n3936 9.3005
R19444 gnd.n4001 gnd.n4000 9.3005
R19445 gnd.n3938 gnd.n3937 9.3005
R19446 gnd.n3994 gnd.n3993 9.3005
R19447 gnd.n3992 gnd.n3943 9.3005
R19448 gnd.n3991 gnd.n3990 9.3005
R19449 gnd.n3945 gnd.n3944 9.3005
R19450 gnd.n3984 gnd.n3983 9.3005
R19451 gnd.n3982 gnd.n3947 9.3005
R19452 gnd.n3981 gnd.n3980 9.3005
R19453 gnd.n3949 gnd.n3948 9.3005
R19454 gnd.n3974 gnd.n3973 9.3005
R19455 gnd.n3972 gnd.n3951 9.3005
R19456 gnd.n3971 gnd.n3970 9.3005
R19457 gnd.n3953 gnd.n3952 9.3005
R19458 gnd.n3964 gnd.n3963 9.3005
R19459 gnd.n3962 gnd.n3955 9.3005
R19460 gnd.n3961 gnd.n3960 9.3005
R19461 gnd.n3957 gnd.n3956 9.3005
R19462 gnd.n4053 gnd.n4052 9.3005
R19463 gnd.n4105 gnd.n4104 9.3005
R19464 gnd.n6212 gnd.n2330 9.3005
R19465 gnd.n6211 gnd.n2331 9.3005
R19466 gnd.n2351 gnd.n2332 9.3005
R19467 gnd.n6201 gnd.n2352 9.3005
R19468 gnd.n6200 gnd.n2353 9.3005
R19469 gnd.n6199 gnd.n2354 9.3005
R19470 gnd.n2371 gnd.n2355 9.3005
R19471 gnd.n6189 gnd.n2372 9.3005
R19472 gnd.n6188 gnd.n2373 9.3005
R19473 gnd.n6187 gnd.n2374 9.3005
R19474 gnd.n2392 gnd.n2375 9.3005
R19475 gnd.n6177 gnd.n2393 9.3005
R19476 gnd.n6176 gnd.n2394 9.3005
R19477 gnd.n6175 gnd.n2395 9.3005
R19478 gnd.n2412 gnd.n2396 9.3005
R19479 gnd.n2466 gnd.n2449 9.3005
R19480 gnd.n6126 gnd.n2467 9.3005
R19481 gnd.n6125 gnd.n2468 9.3005
R19482 gnd.n6124 gnd.n2469 9.3005
R19483 gnd.n2486 gnd.n2470 9.3005
R19484 gnd.n6114 gnd.n2487 9.3005
R19485 gnd.n6113 gnd.n2488 9.3005
R19486 gnd.n6112 gnd.n2489 9.3005
R19487 gnd.n2507 gnd.n2490 9.3005
R19488 gnd.n6102 gnd.n2508 9.3005
R19489 gnd.n6101 gnd.n2509 9.3005
R19490 gnd.n6100 gnd.n2510 9.3005
R19491 gnd.n2527 gnd.n2511 9.3005
R19492 gnd.n6090 gnd.n2528 9.3005
R19493 gnd.n6089 gnd.n2529 9.3005
R19494 gnd.n6088 gnd.n2530 9.3005
R19495 gnd.n6213 gnd.n2329 9.3005
R19496 gnd.n6136 gnd.n2413 9.3005
R19497 gnd.n6228 gnd.n2309 9.3005
R19498 gnd.n6227 gnd.n2310 9.3005
R19499 gnd.n6226 gnd.n2311 9.3005
R19500 gnd.n2316 gnd.n2312 9.3005
R19501 gnd.n6220 gnd.n2317 9.3005
R19502 gnd.n6219 gnd.n2318 9.3005
R19503 gnd.n6218 gnd.n2319 9.3005
R19504 gnd.n3738 gnd.n2320 9.3005
R19505 gnd.n3739 gnd.n3737 9.3005
R19506 gnd.n3741 gnd.n3740 9.3005
R19507 gnd.n3735 gnd.n3734 9.3005
R19508 gnd.n3746 gnd.n3745 9.3005
R19509 gnd.n3747 gnd.n3733 9.3005
R19510 gnd.n3810 gnd.n3748 9.3005
R19511 gnd.n3809 gnd.n3749 9.3005
R19512 gnd.n3808 gnd.n3750 9.3005
R19513 gnd.n3753 gnd.n3751 9.3005
R19514 gnd.n3804 gnd.n3754 9.3005
R19515 gnd.n3803 gnd.n3755 9.3005
R19516 gnd.n3802 gnd.n3756 9.3005
R19517 gnd.n3759 gnd.n3757 9.3005
R19518 gnd.n3798 gnd.n3760 9.3005
R19519 gnd.n3797 gnd.n3761 9.3005
R19520 gnd.n2308 gnd.n2307 9.3005
R19521 gnd.n6235 gnd.n839 9.3005
R19522 gnd.n6236 gnd.n838 9.3005
R19523 gnd.n837 gnd.n833 9.3005
R19524 gnd.n6242 gnd.n832 9.3005
R19525 gnd.n6243 gnd.n831 9.3005
R19526 gnd.n6244 gnd.n830 9.3005
R19527 gnd.n829 gnd.n825 9.3005
R19528 gnd.n6250 gnd.n824 9.3005
R19529 gnd.n6251 gnd.n823 9.3005
R19530 gnd.n6252 gnd.n822 9.3005
R19531 gnd.n821 gnd.n817 9.3005
R19532 gnd.n6258 gnd.n816 9.3005
R19533 gnd.n6259 gnd.n815 9.3005
R19534 gnd.n6260 gnd.n814 9.3005
R19535 gnd.n813 gnd.n809 9.3005
R19536 gnd.n6266 gnd.n808 9.3005
R19537 gnd.n6267 gnd.n807 9.3005
R19538 gnd.n6268 gnd.n806 9.3005
R19539 gnd.n805 gnd.n801 9.3005
R19540 gnd.n6274 gnd.n800 9.3005
R19541 gnd.n6275 gnd.n799 9.3005
R19542 gnd.n6276 gnd.n798 9.3005
R19543 gnd.n797 gnd.n793 9.3005
R19544 gnd.n6282 gnd.n792 9.3005
R19545 gnd.n6283 gnd.n791 9.3005
R19546 gnd.n6284 gnd.n790 9.3005
R19547 gnd.n789 gnd.n785 9.3005
R19548 gnd.n6290 gnd.n784 9.3005
R19549 gnd.n6291 gnd.n783 9.3005
R19550 gnd.n6292 gnd.n782 9.3005
R19551 gnd.n781 gnd.n777 9.3005
R19552 gnd.n6298 gnd.n776 9.3005
R19553 gnd.n6299 gnd.n775 9.3005
R19554 gnd.n6300 gnd.n774 9.3005
R19555 gnd.n773 gnd.n769 9.3005
R19556 gnd.n6306 gnd.n768 9.3005
R19557 gnd.n6307 gnd.n767 9.3005
R19558 gnd.n6308 gnd.n766 9.3005
R19559 gnd.n765 gnd.n761 9.3005
R19560 gnd.n6314 gnd.n760 9.3005
R19561 gnd.n6315 gnd.n759 9.3005
R19562 gnd.n6316 gnd.n758 9.3005
R19563 gnd.n757 gnd.n753 9.3005
R19564 gnd.n6322 gnd.n752 9.3005
R19565 gnd.n6323 gnd.n751 9.3005
R19566 gnd.n6324 gnd.n750 9.3005
R19567 gnd.n749 gnd.n745 9.3005
R19568 gnd.n6330 gnd.n744 9.3005
R19569 gnd.n6331 gnd.n743 9.3005
R19570 gnd.n6332 gnd.n742 9.3005
R19571 gnd.n741 gnd.n737 9.3005
R19572 gnd.n6338 gnd.n736 9.3005
R19573 gnd.n6339 gnd.n735 9.3005
R19574 gnd.n6340 gnd.n734 9.3005
R19575 gnd.n733 gnd.n729 9.3005
R19576 gnd.n6346 gnd.n728 9.3005
R19577 gnd.n6347 gnd.n727 9.3005
R19578 gnd.n6348 gnd.n726 9.3005
R19579 gnd.n725 gnd.n721 9.3005
R19580 gnd.n6354 gnd.n720 9.3005
R19581 gnd.n6355 gnd.n719 9.3005
R19582 gnd.n6356 gnd.n718 9.3005
R19583 gnd.n717 gnd.n713 9.3005
R19584 gnd.n6362 gnd.n712 9.3005
R19585 gnd.n6363 gnd.n711 9.3005
R19586 gnd.n6364 gnd.n710 9.3005
R19587 gnd.n709 gnd.n705 9.3005
R19588 gnd.n6370 gnd.n704 9.3005
R19589 gnd.n6371 gnd.n703 9.3005
R19590 gnd.n6372 gnd.n702 9.3005
R19591 gnd.n701 gnd.n697 9.3005
R19592 gnd.n6378 gnd.n696 9.3005
R19593 gnd.n6379 gnd.n695 9.3005
R19594 gnd.n6380 gnd.n694 9.3005
R19595 gnd.n693 gnd.n689 9.3005
R19596 gnd.n6386 gnd.n688 9.3005
R19597 gnd.n6387 gnd.n687 9.3005
R19598 gnd.n6388 gnd.n686 9.3005
R19599 gnd.n685 gnd.n681 9.3005
R19600 gnd.n6394 gnd.n680 9.3005
R19601 gnd.n6395 gnd.n679 9.3005
R19602 gnd.n6396 gnd.n678 9.3005
R19603 gnd.n674 gnd.n673 9.3005
R19604 gnd.n6403 gnd.n6402 9.3005
R19605 gnd.n6234 gnd.n840 9.3005
R19606 gnd.n5937 gnd.n5936 9.3005
R19607 gnd.n6060 gnd.n6059 9.3005
R19608 gnd.n6058 gnd.n2577 9.3005
R19609 gnd.n6057 gnd.n6056 9.3005
R19610 gnd.n6055 gnd.n2579 9.3005
R19611 gnd.n6054 gnd.n6053 9.3005
R19612 gnd.n6052 gnd.n2583 9.3005
R19613 gnd.n6051 gnd.n6050 9.3005
R19614 gnd.n6049 gnd.n2584 9.3005
R19615 gnd.n6048 gnd.n6047 9.3005
R19616 gnd.n6046 gnd.n2588 9.3005
R19617 gnd.n6045 gnd.n6044 9.3005
R19618 gnd.n6043 gnd.n2589 9.3005
R19619 gnd.n6042 gnd.n6041 9.3005
R19620 gnd.n6040 gnd.n2593 9.3005
R19621 gnd.n6039 gnd.n6038 9.3005
R19622 gnd.n6037 gnd.n2594 9.3005
R19623 gnd.n6036 gnd.n6035 9.3005
R19624 gnd.n6034 gnd.n2598 9.3005
R19625 gnd.n6033 gnd.n6032 9.3005
R19626 gnd.n6031 gnd.n2599 9.3005
R19627 gnd.n6030 gnd.n6029 9.3005
R19628 gnd.n6028 gnd.n2603 9.3005
R19629 gnd.n6027 gnd.n6026 9.3005
R19630 gnd.n6025 gnd.n2604 9.3005
R19631 gnd.n6024 gnd.n6023 9.3005
R19632 gnd.n6022 gnd.n2608 9.3005
R19633 gnd.n6021 gnd.n6020 9.3005
R19634 gnd.n6019 gnd.n2609 9.3005
R19635 gnd.n6018 gnd.n6017 9.3005
R19636 gnd.n6016 gnd.n2613 9.3005
R19637 gnd.n6015 gnd.n6014 9.3005
R19638 gnd.n6013 gnd.n2614 9.3005
R19639 gnd.n6012 gnd.n6011 9.3005
R19640 gnd.n6010 gnd.n2618 9.3005
R19641 gnd.n6009 gnd.n6008 9.3005
R19642 gnd.n6007 gnd.n2619 9.3005
R19643 gnd.n6006 gnd.n6005 9.3005
R19644 gnd.n6004 gnd.n2623 9.3005
R19645 gnd.n6003 gnd.n6002 9.3005
R19646 gnd.n6001 gnd.n2624 9.3005
R19647 gnd.n6000 gnd.n5999 9.3005
R19648 gnd.n5998 gnd.n2628 9.3005
R19649 gnd.n5997 gnd.n5996 9.3005
R19650 gnd.n5995 gnd.n2629 9.3005
R19651 gnd.n5994 gnd.n5993 9.3005
R19652 gnd.n5992 gnd.n2633 9.3005
R19653 gnd.n5991 gnd.n5990 9.3005
R19654 gnd.n5989 gnd.n2634 9.3005
R19655 gnd.n5988 gnd.n5987 9.3005
R19656 gnd.n5986 gnd.n2638 9.3005
R19657 gnd.n5985 gnd.n5984 9.3005
R19658 gnd.n5983 gnd.n2639 9.3005
R19659 gnd.n5982 gnd.n5981 9.3005
R19660 gnd.n5980 gnd.n2643 9.3005
R19661 gnd.n5979 gnd.n5978 9.3005
R19662 gnd.n5977 gnd.n2644 9.3005
R19663 gnd.n5976 gnd.n5975 9.3005
R19664 gnd.n5974 gnd.n2648 9.3005
R19665 gnd.n5973 gnd.n5972 9.3005
R19666 gnd.n5971 gnd.n2649 9.3005
R19667 gnd.n5970 gnd.n5969 9.3005
R19668 gnd.n5968 gnd.n2653 9.3005
R19669 gnd.n5967 gnd.n5966 9.3005
R19670 gnd.n5965 gnd.n2654 9.3005
R19671 gnd.n5964 gnd.n5963 9.3005
R19672 gnd.n5962 gnd.n2658 9.3005
R19673 gnd.n5961 gnd.n5960 9.3005
R19674 gnd.n5959 gnd.n2659 9.3005
R19675 gnd.n5958 gnd.n5957 9.3005
R19676 gnd.n5956 gnd.n2663 9.3005
R19677 gnd.n5955 gnd.n5954 9.3005
R19678 gnd.n5953 gnd.n2664 9.3005
R19679 gnd.n5952 gnd.n5951 9.3005
R19680 gnd.n5950 gnd.n2668 9.3005
R19681 gnd.n5949 gnd.n5948 9.3005
R19682 gnd.n5947 gnd.n2669 9.3005
R19683 gnd.n5946 gnd.n5945 9.3005
R19684 gnd.n5944 gnd.n2673 9.3005
R19685 gnd.n5943 gnd.n5942 9.3005
R19686 gnd.n5941 gnd.n2674 9.3005
R19687 gnd.n5940 gnd.n5939 9.3005
R19688 gnd.n5938 gnd.n2678 9.3005
R19689 gnd.n2578 gnd.n2576 9.3005
R19690 gnd.n6071 gnd.n2544 9.3005
R19691 gnd.n3708 gnd.n3707 9.3005
R19692 gnd.n4187 gnd.n4186 9.3005
R19693 gnd.n4188 gnd.n3706 9.3005
R19694 gnd.n4190 gnd.n4189 9.3005
R19695 gnd.n3703 gnd.n3702 9.3005
R19696 gnd.n4201 gnd.n4200 9.3005
R19697 gnd.n4202 gnd.n3701 9.3005
R19698 gnd.n4204 gnd.n4203 9.3005
R19699 gnd.n3692 gnd.n3690 9.3005
R19700 gnd.n4243 gnd.n4242 9.3005
R19701 gnd.n4241 gnd.n3691 9.3005
R19702 gnd.n4240 gnd.n4239 9.3005
R19703 gnd.n4238 gnd.n3693 9.3005
R19704 gnd.n4237 gnd.n4236 9.3005
R19705 gnd.n4235 gnd.n3696 9.3005
R19706 gnd.n4234 gnd.n4233 9.3005
R19707 gnd.n4232 gnd.n3697 9.3005
R19708 gnd.n4231 gnd.n4230 9.3005
R19709 gnd.n2543 gnd.n2541 9.3005
R19710 gnd.n6077 gnd.n6076 9.3005
R19711 gnd.n6075 gnd.n2542 9.3005
R19712 gnd.n3413 gnd.n3412 9.3005
R19713 gnd.n3606 gnd.n3605 9.3005
R19714 gnd.n3610 gnd.n3609 9.3005
R19715 gnd.n3406 gnd.n3403 9.3005
R19716 gnd.n3618 gnd.n3617 9.3005
R19717 gnd.n3622 gnd.n3621 9.3005
R19718 gnd.n3400 gnd.n3399 9.3005
R19719 gnd.n3630 gnd.n3629 9.3005
R19720 gnd.n3634 gnd.n3633 9.3005
R19721 gnd.n3394 gnd.n3391 9.3005
R19722 gnd.n3642 gnd.n3641 9.3005
R19723 gnd.n3646 gnd.n3645 9.3005
R19724 gnd.n3388 gnd.n3387 9.3005
R19725 gnd.n3654 gnd.n3653 9.3005
R19726 gnd.n3658 gnd.n3657 9.3005
R19727 gnd.n3380 gnd.n3377 9.3005
R19728 gnd.n3668 gnd.n3667 9.3005
R19729 gnd.n3669 gnd.n2545 9.3005
R19730 gnd.n3598 gnd.n3597 9.3005
R19731 gnd.n6073 gnd.n6072 9.3005
R19732 gnd.n3666 gnd.n2546 9.3005
R19733 gnd.n3665 gnd.n3664 9.3005
R19734 gnd.n3660 gnd.n3659 9.3005
R19735 gnd.n3386 gnd.n3383 9.3005
R19736 gnd.n3652 gnd.n3651 9.3005
R19737 gnd.n3648 gnd.n3647 9.3005
R19738 gnd.n3390 gnd.n3389 9.3005
R19739 gnd.n3640 gnd.n3639 9.3005
R19740 gnd.n3636 gnd.n3635 9.3005
R19741 gnd.n3398 gnd.n3395 9.3005
R19742 gnd.n3628 gnd.n3627 9.3005
R19743 gnd.n3624 gnd.n3623 9.3005
R19744 gnd.n3402 gnd.n3401 9.3005
R19745 gnd.n3616 gnd.n3615 9.3005
R19746 gnd.n3612 gnd.n3611 9.3005
R19747 gnd.n3410 gnd.n3407 9.3005
R19748 gnd.n3604 gnd.n3603 9.3005
R19749 gnd.n3600 gnd.n3599 9.3005
R19750 gnd.n3596 gnd.n3414 9.3005
R19751 gnd.n3595 gnd.n3594 9.3005
R19752 gnd.n3591 gnd.n3590 9.3005
R19753 gnd.n3589 gnd.n3416 9.3005
R19754 gnd.n3588 gnd.n3587 9.3005
R19755 gnd.n3584 gnd.n3419 9.3005
R19756 gnd.n3583 gnd.n3582 9.3005
R19757 gnd.n3581 gnd.n3420 9.3005
R19758 gnd.n3580 gnd.n3579 9.3005
R19759 gnd.n3575 gnd.n3423 9.3005
R19760 gnd.n3574 gnd.n3573 9.3005
R19761 gnd.n3572 gnd.n3425 9.3005
R19762 gnd.n3571 gnd.n3570 9.3005
R19763 gnd.n3569 gnd.n3426 9.3005
R19764 gnd.n3568 gnd.n3567 9.3005
R19765 gnd.n3566 gnd.n3430 9.3005
R19766 gnd.n3565 gnd.n3564 9.3005
R19767 gnd.n3563 gnd.n3431 9.3005
R19768 gnd.n3562 gnd.n3561 9.3005
R19769 gnd.n3560 gnd.n3435 9.3005
R19770 gnd.n3559 gnd.n3558 9.3005
R19771 gnd.n3557 gnd.n3436 9.3005
R19772 gnd.n3556 gnd.n3555 9.3005
R19773 gnd.n3554 gnd.n3489 9.3005
R19774 gnd.n3553 gnd.n3552 9.3005
R19775 gnd.n3551 gnd.n3490 9.3005
R19776 gnd.n3550 gnd.n3549 9.3005
R19777 gnd.n3548 gnd.n3496 9.3005
R19778 gnd.n3547 gnd.n3546 9.3005
R19779 gnd.n3545 gnd.n3497 9.3005
R19780 gnd.n3544 gnd.n3543 9.3005
R19781 gnd.n3542 gnd.n3502 9.3005
R19782 gnd.n3541 gnd.n3540 9.3005
R19783 gnd.n3539 gnd.n3503 9.3005
R19784 gnd.n3538 gnd.n3537 9.3005
R19785 gnd.n3536 gnd.n3505 9.3005
R19786 gnd.n3535 gnd.n3534 9.3005
R19787 gnd.n3533 gnd.n3506 9.3005
R19788 gnd.n3532 gnd.n3531 9.3005
R19789 gnd.n3530 gnd.n3510 9.3005
R19790 gnd.n3529 gnd.n3528 9.3005
R19791 gnd.n3527 gnd.n3511 9.3005
R19792 gnd.n3526 gnd.n3525 9.3005
R19793 gnd.n3524 gnd.n3514 9.3005
R19794 gnd.n3523 gnd.n3522 9.3005
R19795 gnd.n3521 gnd.n3515 9.3005
R19796 gnd.n3520 gnd.n3519 9.3005
R19797 gnd.n3518 gnd.n3517 9.3005
R19798 gnd.n3089 gnd.n3088 9.3005
R19799 gnd.n4765 gnd.n4764 9.3005
R19800 gnd.n4766 gnd.n3086 9.3005
R19801 gnd.n4782 gnd.n4781 9.3005
R19802 gnd.n4780 gnd.n3087 9.3005
R19803 gnd.n4779 gnd.n4778 9.3005
R19804 gnd.n4777 gnd.n4767 9.3005
R19805 gnd.n4776 gnd.n4775 9.3005
R19806 gnd.n4774 gnd.n4771 9.3005
R19807 gnd.n4773 gnd.n4772 9.3005
R19808 gnd.n3036 gnd.n3035 9.3005
R19809 gnd.n4874 gnd.n4873 9.3005
R19810 gnd.n4875 gnd.n3033 9.3005
R19811 gnd.n4878 gnd.n4877 9.3005
R19812 gnd.n4876 gnd.n3034 9.3005
R19813 gnd.n3013 gnd.n3012 9.3005
R19814 gnd.n4907 gnd.n4906 9.3005
R19815 gnd.n4908 gnd.n3010 9.3005
R19816 gnd.n4937 gnd.n4936 9.3005
R19817 gnd.n4935 gnd.n3011 9.3005
R19818 gnd.n4934 gnd.n4933 9.3005
R19819 gnd.n4932 gnd.n4909 9.3005
R19820 gnd.n4931 gnd.n4930 9.3005
R19821 gnd.n4929 gnd.n4916 9.3005
R19822 gnd.n4928 gnd.n4927 9.3005
R19823 gnd.n4926 gnd.n4917 9.3005
R19824 gnd.n4925 gnd.n4924 9.3005
R19825 gnd.n4923 gnd.n4920 9.3005
R19826 gnd.n4922 gnd.n4921 9.3005
R19827 gnd.n2875 gnd.n2874 9.3005
R19828 gnd.n5139 gnd.n5138 9.3005
R19829 gnd.n5140 gnd.n2873 9.3005
R19830 gnd.n5142 gnd.n5141 9.3005
R19831 gnd.n2862 gnd.n2861 9.3005
R19832 gnd.n5155 gnd.n5154 9.3005
R19833 gnd.n5156 gnd.n2860 9.3005
R19834 gnd.n5158 gnd.n5157 9.3005
R19835 gnd.n2850 gnd.n2849 9.3005
R19836 gnd.n5171 gnd.n5170 9.3005
R19837 gnd.n5172 gnd.n2847 9.3005
R19838 gnd.n5175 gnd.n5174 9.3005
R19839 gnd.n5173 gnd.n2848 9.3005
R19840 gnd.n2838 gnd.n2836 9.3005
R19841 gnd.n3577 gnd.n3576 9.3005
R19842 gnd.n5191 gnd.n2833 9.3005
R19843 gnd.n5193 gnd.n5192 9.3005
R19844 gnd.n5194 gnd.n2832 9.3005
R19845 gnd.n5198 gnd.n5197 9.3005
R19846 gnd.n5199 gnd.n2829 9.3005
R19847 gnd.n5201 gnd.n5200 9.3005
R19848 gnd.n5190 gnd.n5189 9.3005
R19849 gnd.n5275 gnd.n5274 9.3005
R19850 gnd.n5277 gnd.n5276 9.3005
R19851 gnd.n5248 gnd.n5247 9.3005
R19852 gnd.n5283 gnd.n5282 9.3005
R19853 gnd.n5285 gnd.n5284 9.3005
R19854 gnd.n5238 gnd.n5237 9.3005
R19855 gnd.n5291 gnd.n5290 9.3005
R19856 gnd.n5293 gnd.n5292 9.3005
R19857 gnd.n5228 gnd.n5227 9.3005
R19858 gnd.n5299 gnd.n5298 9.3005
R19859 gnd.n5301 gnd.n5300 9.3005
R19860 gnd.n5218 gnd.n5217 9.3005
R19861 gnd.n5307 gnd.n5306 9.3005
R19862 gnd.n5309 gnd.n5308 9.3005
R19863 gnd.n2828 gnd.n2826 9.3005
R19864 gnd.n5315 gnd.n5314 9.3005
R19865 gnd.n5316 gnd.n2823 9.3005
R19866 gnd.n5261 gnd.n5260 9.3005
R19867 gnd.n5269 gnd.n5268 9.3005
R19868 gnd.n5205 gnd.n5202 9.3005
R19869 gnd.n5207 gnd.n5206 9.3005
R19870 gnd.n5208 gnd.n2827 9.3005
R19871 gnd.n5313 gnd.n5312 9.3005
R19872 gnd.n5311 gnd.n5310 9.3005
R19873 gnd.n5214 gnd.n5213 9.3005
R19874 gnd.n5305 gnd.n5304 9.3005
R19875 gnd.n5303 gnd.n5302 9.3005
R19876 gnd.n5222 gnd.n5221 9.3005
R19877 gnd.n5297 gnd.n5296 9.3005
R19878 gnd.n5295 gnd.n5294 9.3005
R19879 gnd.n5234 gnd.n5233 9.3005
R19880 gnd.n5289 gnd.n5288 9.3005
R19881 gnd.n5287 gnd.n5286 9.3005
R19882 gnd.n5242 gnd.n5241 9.3005
R19883 gnd.n5281 gnd.n5280 9.3005
R19884 gnd.n5279 gnd.n5278 9.3005
R19885 gnd.n5254 gnd.n5253 9.3005
R19886 gnd.n5273 gnd.n5272 9.3005
R19887 gnd.n5271 gnd.n5270 9.3005
R19888 gnd.n5267 gnd.n2680 9.3005
R19889 gnd.n5491 gnd.n5488 9.3005
R19890 gnd.n5498 gnd.n5497 9.3005
R19891 gnd.n5499 gnd.n5487 9.3005
R19892 gnd.n5501 gnd.n5500 9.3005
R19893 gnd.n5481 gnd.n5479 9.3005
R19894 gnd.n5537 gnd.n5536 9.3005
R19895 gnd.n5535 gnd.n5480 9.3005
R19896 gnd.n5534 gnd.n5533 9.3005
R19897 gnd.n5532 gnd.n5482 9.3005
R19898 gnd.n5531 gnd.n5530 9.3005
R19899 gnd.n5529 gnd.n5485 9.3005
R19900 gnd.n5528 gnd.n5527 9.3005
R19901 gnd.n5443 gnd.n5442 9.3005
R19902 gnd.n5567 gnd.n5566 9.3005
R19903 gnd.n5568 gnd.n5440 9.3005
R19904 gnd.n5578 gnd.n5577 9.3005
R19905 gnd.n5576 gnd.n5441 9.3005
R19906 gnd.n5575 gnd.n5574 9.3005
R19907 gnd.n5573 gnd.n5569 9.3005
R19908 gnd.n5572 gnd.n63 9.3005
R19909 gnd.n5490 gnd.n5489 9.3005
R19910 gnd.n7407 gnd.n64 9.3005
R19911 gnd.t305 gnd.n1031 9.24152
R19912 gnd.n934 gnd.t215 9.24152
R19913 gnd.n2203 gnd.t180 9.24152
R19914 gnd.t150 gnd.t305 8.92286
R19915 gnd.t246 gnd.n2963 8.92286
R19916 gnd.n2173 gnd.n2148 8.92171
R19917 gnd.n2141 gnd.n2116 8.92171
R19918 gnd.n2109 gnd.n2084 8.92171
R19919 gnd.n2078 gnd.n2053 8.92171
R19920 gnd.n2046 gnd.n2021 8.92171
R19921 gnd.n2014 gnd.n1989 8.92171
R19922 gnd.n1982 gnd.n1957 8.92171
R19923 gnd.n1951 gnd.n1926 8.92171
R19924 gnd.n2910 gnd.n2892 8.72777
R19925 gnd.n1675 gnd.t294 8.60421
R19926 gnd.n1095 gnd.n1083 8.43656
R19927 gnd.n38 gnd.n26 8.43656
R19928 gnd.n3498 gnd.t279 8.28555
R19929 gnd.n4627 gnd.t5 8.28555
R19930 gnd.n4650 gnd.n3159 8.28555
R19931 gnd.n3114 gnd.n3109 8.28555
R19932 gnd.n3079 gnd.n3066 8.28555
R19933 gnd.n4894 gnd.n4892 8.28555
R19934 gnd.t4 gnd.n3001 8.28555
R19935 gnd.n2174 gnd.n2146 8.14595
R19936 gnd.n2142 gnd.n2114 8.14595
R19937 gnd.n2110 gnd.n2082 8.14595
R19938 gnd.n2079 gnd.n2051 8.14595
R19939 gnd.n2047 gnd.n2019 8.14595
R19940 gnd.n2015 gnd.n1987 8.14595
R19941 gnd.n1983 gnd.n1955 8.14595
R19942 gnd.n1952 gnd.n1924 8.14595
R19943 gnd.n4175 gnd.n0 8.10675
R19944 gnd.n7408 gnd.n7407 8.10675
R19945 gnd.n2179 gnd.n2178 7.97301
R19946 gnd.t296 gnd.n1190 7.9669
R19947 gnd.n7408 gnd.n62 7.78567
R19948 gnd.n5268 gnd.n5260 7.75808
R19949 gnd.n3669 gnd.n3668 7.75808
R19950 gnd.n7333 gnd.n180 7.75808
R19951 gnd.n3857 gnd.n3845 7.75808
R19952 gnd.n3215 gnd.t205 7.64824
R19953 gnd.n1120 gnd.n1119 7.53171
R19954 gnd.n1584 gnd.t299 7.32958
R19955 gnd.n3244 gnd.n3243 7.30353
R19956 gnd.n2909 gnd.n2908 7.30353
R19957 gnd.n1544 gnd.n1263 7.01093
R19958 gnd.n1266 gnd.n1264 7.01093
R19959 gnd.n1554 gnd.n1553 7.01093
R19960 gnd.n1565 gnd.n1247 7.01093
R19961 gnd.n1564 gnd.n1250 7.01093
R19962 gnd.n1575 gnd.n1238 7.01093
R19963 gnd.n1241 gnd.n1239 7.01093
R19964 gnd.n1585 gnd.n1584 7.01093
R19965 gnd.n1595 gnd.n1219 7.01093
R19966 gnd.n1594 gnd.n1222 7.01093
R19967 gnd.n1603 gnd.n1213 7.01093
R19968 gnd.n1615 gnd.n1203 7.01093
R19969 gnd.n1625 gnd.n1188 7.01093
R19970 gnd.n1641 gnd.n1640 7.01093
R19971 gnd.n1190 gnd.n1127 7.01093
R19972 gnd.n1695 gnd.n1128 7.01093
R19973 gnd.n1689 gnd.n1688 7.01093
R19974 gnd.n1177 gnd.n1139 7.01093
R19975 gnd.n1681 gnd.n1150 7.01093
R19976 gnd.n1168 gnd.n1163 7.01093
R19977 gnd.n1675 gnd.n1674 7.01093
R19978 gnd.n1721 gnd.n1066 7.01093
R19979 gnd.n1720 gnd.n1719 7.01093
R19980 gnd.n1732 gnd.n1731 7.01093
R19981 gnd.n1059 gnd.n1051 7.01093
R19982 gnd.n1761 gnd.n1039 7.01093
R19983 gnd.n1760 gnd.n1042 7.01093
R19984 gnd.n1771 gnd.n1031 7.01093
R19985 gnd.n1032 gnd.n1020 7.01093
R19986 gnd.n1782 gnd.n1021 7.01093
R19987 gnd.n1808 gnd.n1013 7.01093
R19988 gnd.n1807 gnd.n1806 7.01093
R19989 gnd.n1806 gnd.n1004 7.01093
R19990 gnd.n1830 gnd.n1829 7.01093
R19991 gnd.n1848 gnd.n985 7.01093
R19992 gnd.n1847 gnd.n988 7.01093
R19993 gnd.n1858 gnd.n977 7.01093
R19994 gnd.n978 gnd.n965 7.01093
R19995 gnd.n1869 gnd.n966 7.01093
R19996 gnd.n1896 gnd.n950 7.01093
R19997 gnd.n1908 gnd.n1907 7.01093
R19998 gnd.n1890 gnd.n943 7.01093
R19999 gnd.n1919 gnd.n1918 7.01093
R20000 gnd.n2191 gnd.n931 7.01093
R20001 gnd.n2190 gnd.n934 7.01093
R20002 gnd.n2203 gnd.n923 7.01093
R20003 gnd.n924 gnd.n916 7.01093
R20004 gnd.n2213 gnd.n842 7.01093
R20005 gnd.n4670 gnd.n3145 7.01093
R20006 gnd.n4708 gnd.n3118 7.01093
R20007 gnd.n4706 gnd.t3 7.01093
R20008 gnd.t10 gnd.n4802 7.01093
R20009 gnd.n4809 gnd.n3062 7.01093
R20010 gnd.n4815 gnd.n4814 7.01093
R20011 gnd.n4985 gnd.n2976 7.01093
R20012 gnd.n2969 gnd.t246 7.01093
R20013 gnd.n1222 gnd.t303 6.69227
R20014 gnd.n1042 gnd.t150 6.69227
R20015 gnd.n1897 gnd.t293 6.69227
R20016 gnd.t26 gnd.n2502 6.69227
R20017 gnd.n3498 gnd.t139 6.69227
R20018 gnd.n4913 gnd.t311 6.69227
R20019 gnd.n5540 gnd.t33 6.69227
R20020 gnd.n5058 gnd.n5057 6.5566
R20021 gnd.n3354 gnd.n3353 6.5566
R20022 gnd.n4491 gnd.n3285 6.5566
R20023 gnd.n5073 gnd.n5072 6.5566
R20024 gnd.n3664 gnd.n3661 6.20656
R20025 gnd.n5272 gnd.n5264 6.20656
R20026 gnd.t153 gnd.n1651 6.05496
R20027 gnd.n1652 gnd.t302 6.05496
R20028 gnd.t141 gnd.n1066 6.05496
R20029 gnd.t295 gnd.n1818 6.05496
R20030 gnd.t20 gnd.n2461 6.05496
R20031 gnd.n5563 gnd.t41 6.05496
R20032 gnd.n2176 gnd.n2146 5.81868
R20033 gnd.n2144 gnd.n2114 5.81868
R20034 gnd.n2112 gnd.n2082 5.81868
R20035 gnd.n2081 gnd.n2051 5.81868
R20036 gnd.n2049 gnd.n2019 5.81868
R20037 gnd.n2017 gnd.n1987 5.81868
R20038 gnd.n1985 gnd.n1955 5.81868
R20039 gnd.n1954 gnd.n1924 5.81868
R20040 gnd.n6222 gnd.n2314 5.73631
R20041 gnd.n3289 gnd.n3212 5.73631
R20042 gnd.n4566 gnd.n3215 5.73631
R20043 gnd.n4679 gnd.n4678 5.73631
R20044 gnd.n4686 gnd.n3132 5.73631
R20045 gnd.n4861 gnd.n3046 5.73631
R20046 gnd.n4842 gnd.n3050 5.73631
R20047 gnd.n4994 gnd.n4993 5.73631
R20048 gnd.n5000 gnd.n2963 5.73631
R20049 gnd.n7330 gnd.n7117 5.73631
R20050 gnd.n2936 gnd.n2777 5.62001
R20051 gnd.n4486 gnd.n3358 5.62001
R20052 gnd.n4487 gnd.n4486 5.62001
R20053 gnd.n5067 gnd.n2777 5.62001
R20054 gnd.n1403 gnd.n1398 5.4308
R20055 gnd.n2221 gnd.n909 5.4308
R20056 gnd.n1719 gnd.t292 5.41765
R20057 gnd.t298 gnd.n1742 5.41765
R20058 gnd.t143 gnd.n997 5.41765
R20059 gnd.t84 gnd.n2426 5.41765
R20060 gnd.n4634 gnd.t136 5.41765
R20061 gnd.n4818 gnd.t167 5.41765
R20062 gnd.n5598 gnd.t63 5.41765
R20063 gnd.n6216 gnd.n6215 5.09899
R20064 gnd.n3848 gnd.n2325 5.09899
R20065 gnd.n6209 gnd.n2334 5.09899
R20066 gnd.n4114 gnd.n2337 5.09899
R20067 gnd.n6203 gnd.n2346 5.09899
R20068 gnd.n4122 gnd.n2349 5.09899
R20069 gnd.n6197 gnd.n2357 5.09899
R20070 gnd.n4128 gnd.n3812 5.09899
R20071 gnd.n6191 gnd.n2366 5.09899
R20072 gnd.n4136 gnd.n2369 5.09899
R20073 gnd.n6185 gnd.n2377 5.09899
R20074 gnd.n4142 gnd.n2380 5.09899
R20075 gnd.n6179 gnd.n2387 5.09899
R20076 gnd.n4150 gnd.n2390 5.09899
R20077 gnd.n6173 gnd.n2398 5.09899
R20078 gnd.n4156 gnd.n3720 5.09899
R20079 gnd.n6167 gnd.n2407 5.09899
R20080 gnd.n4164 gnd.n2410 5.09899
R20081 gnd.n6160 gnd.n2416 5.09899
R20082 gnd.n4170 gnd.n2419 5.09899
R20083 gnd.n6154 gnd.n2426 5.09899
R20084 gnd.n4178 gnd.n2429 5.09899
R20085 gnd.n6147 gnd.n2434 5.09899
R20086 gnd.n4184 gnd.n3709 5.09899
R20087 gnd.n6141 gnd.n2443 5.09899
R20088 gnd.n6134 gnd.n2451 5.09899
R20089 gnd.n4198 gnd.n2454 5.09899
R20090 gnd.n6128 gnd.n2461 5.09899
R20091 gnd.n4206 gnd.n2464 5.09899
R20092 gnd.n6122 gnd.n2472 5.09899
R20093 gnd.n4246 gnd.n4245 5.09899
R20094 gnd.n6116 gnd.n2481 5.09899
R20095 gnd.n6110 gnd.n2492 5.09899
R20096 gnd.n4217 gnd.n2495 5.09899
R20097 gnd.n6104 gnd.n2502 5.09899
R20098 gnd.n4222 gnd.n2505 5.09899
R20099 gnd.n6098 gnd.n2513 5.09899
R20100 gnd.n4228 gnd.n2516 5.09899
R20101 gnd.n6092 gnd.n2523 5.09899
R20102 gnd.n6079 gnd.n2540 5.09899
R20103 gnd.n6086 gnd.n2532 5.09899
R20104 gnd.n4593 gnd.t279 5.09899
R20105 gnd.n4577 gnd.t155 5.09899
R20106 gnd.t166 gnd.n3152 5.09899
R20107 gnd.n4655 gnd.t152 5.09899
R20108 gnd.t164 gnd.n3038 5.09899
R20109 gnd.n4880 gnd.t145 5.09899
R20110 gnd.n4959 gnd.t7 5.09899
R20111 gnd.t184 gnd.n5127 5.09899
R20112 gnd.n5807 gnd.n2822 5.09899
R20113 gnd.n5804 gnd.n5321 5.09899
R20114 gnd.n5495 gnd.n5330 5.09899
R20115 gnd.n5798 gnd.n5333 5.09899
R20116 gnd.n5503 gnd.n5341 5.09899
R20117 gnd.n5792 gnd.n5344 5.09899
R20118 gnd.n5540 gnd.n5539 5.09899
R20119 gnd.n5786 gnd.n5354 5.09899
R20120 gnd.n5510 gnd.n5361 5.09899
R20121 gnd.n5516 gnd.n5371 5.09899
R20122 gnd.n5774 gnd.n5374 5.09899
R20123 gnd.n5525 gnd.n5381 5.09899
R20124 gnd.n5768 gnd.n5384 5.09899
R20125 gnd.n5564 gnd.n5563 5.09899
R20126 gnd.n5762 gnd.n5393 5.09899
R20127 gnd.n5580 gnd.n5400 5.09899
R20128 gnd.n5751 gnd.n5750 5.09899
R20129 gnd.n5413 gnd.n5407 5.09899
R20130 gnd.n5743 gnd.n5414 5.09899
R20131 gnd.n5742 gnd.n5417 5.09899
R20132 gnd.n5599 gnd.n5598 5.09899
R20133 gnd.n7402 gnd.n70 5.09899
R20134 gnd.n5729 gnd.n5728 5.09899
R20135 gnd.n5610 gnd.n85 5.09899
R20136 gnd.n7394 gnd.n88 5.09899
R20137 gnd.n5720 gnd.n5719 5.09899
R20138 gnd.n7388 gnd.n99 5.09899
R20139 gnd.n5713 gnd.n106 5.09899
R20140 gnd.n7382 gnd.n109 5.09899
R20141 gnd.n5707 gnd.n116 5.09899
R20142 gnd.n7376 gnd.n119 5.09899
R20143 gnd.n5701 gnd.n127 5.09899
R20144 gnd.n7370 gnd.n130 5.09899
R20145 gnd.n5695 gnd.n5694 5.09899
R20146 gnd.n7364 gnd.n139 5.09899
R20147 gnd.n5642 gnd.n147 5.09899
R20148 gnd.n7358 gnd.n150 5.09899
R20149 gnd.n5636 gnd.n157 5.09899
R20150 gnd.n7352 gnd.n160 5.09899
R20151 gnd.n7339 gnd.n167 5.09899
R20152 gnd.n7346 gnd.n170 5.09899
R20153 gnd.n2174 gnd.n2173 5.04292
R20154 gnd.n2142 gnd.n2141 5.04292
R20155 gnd.n2110 gnd.n2109 5.04292
R20156 gnd.n2079 gnd.n2078 5.04292
R20157 gnd.n2047 gnd.n2046 5.04292
R20158 gnd.n2015 gnd.n2014 5.04292
R20159 gnd.n1983 gnd.n1982 5.04292
R20160 gnd.n1952 gnd.n1951 5.04292
R20161 gnd.n1682 gnd.t301 4.78034
R20162 gnd.n1021 gnd.t291 4.78034
R20163 gnd.t46 gnd.n2387 4.78034
R20164 gnd.t31 gnd.n2446 4.78034
R20165 gnd.n5404 gnd.t15 4.78034
R20166 gnd.t80 gnd.n109 4.78034
R20167 gnd.n1124 gnd.n1121 4.74817
R20168 gnd.n1174 gnd.n1072 4.74817
R20169 gnd.n1161 gnd.n1071 4.74817
R20170 gnd.n1070 gnd.n1069 4.74817
R20171 gnd.n1170 gnd.n1121 4.74817
R20172 gnd.n1171 gnd.n1072 4.74817
R20173 gnd.n1173 gnd.n1071 4.74817
R20174 gnd.n1160 gnd.n1070 4.74817
R20175 gnd.n5754 gnd.n81 4.74817
R20176 gnd.n5736 gnd.n80 4.74817
R20177 gnd.n5740 gnd.n79 4.74817
R20178 gnd.n7400 gnd.n74 4.74817
R20179 gnd.n7398 gnd.n75 4.74817
R20180 gnd.n5389 gnd.n81 4.74817
R20181 gnd.n5753 gnd.n80 4.74817
R20182 gnd.n5737 gnd.n79 4.74817
R20183 gnd.n5739 gnd.n74 4.74817
R20184 gnd.n7399 gnd.n7398 4.74817
R20185 gnd.n3796 gnd.n3795 4.74817
R20186 gnd.n3793 gnd.n3768 4.74817
R20187 gnd.n3786 gnd.n3767 4.74817
R20188 gnd.n3782 gnd.n3766 4.74817
R20189 gnd.n3778 gnd.n3765 4.74817
R20190 gnd.n5557 gnd.n5410 4.74817
R20191 gnd.n5747 gnd.n5746 4.74817
R20192 gnd.n5594 gnd.n5411 4.74817
R20193 gnd.n5595 gnd.n5428 4.74817
R20194 gnd.n5725 gnd.n5724 4.74817
R20195 gnd.n5559 gnd.n5557 4.74817
R20196 gnd.n5748 gnd.n5747 4.74817
R20197 gnd.n5745 gnd.n5411 4.74817
R20198 gnd.n5596 gnd.n5595 4.74817
R20199 gnd.n5726 gnd.n5725 4.74817
R20200 gnd.n6164 gnd.n6163 4.74817
R20201 gnd.n2431 gnd.n2414 4.74817
R20202 gnd.n6151 gnd.n6150 4.74817
R20203 gnd.n2448 gnd.n2432 4.74817
R20204 gnd.n6138 gnd.n6137 4.74817
R20205 gnd.n6165 gnd.n6164 4.74817
R20206 gnd.n6162 gnd.n2414 4.74817
R20207 gnd.n6152 gnd.n6151 4.74817
R20208 gnd.n6149 gnd.n2432 4.74817
R20209 gnd.n6139 gnd.n6138 4.74817
R20210 gnd.n3795 gnd.n3763 4.74817
R20211 gnd.n3793 gnd.n3792 4.74817
R20212 gnd.n3788 gnd.n3767 4.74817
R20213 gnd.n3785 gnd.n3766 4.74817
R20214 gnd.n3781 gnd.n3765 4.74817
R20215 gnd.n1119 gnd.n1118 4.74296
R20216 gnd.n62 gnd.n61 4.74296
R20217 gnd.n1095 gnd.n1094 4.7074
R20218 gnd.n1107 gnd.n1106 4.7074
R20219 gnd.n38 gnd.n37 4.7074
R20220 gnd.n50 gnd.n49 4.7074
R20221 gnd.n1119 gnd.n1107 4.65959
R20222 gnd.n62 gnd.n50 4.65959
R20223 gnd.n5874 gnd.n2779 4.6132
R20224 gnd.n4482 gnd.n4481 4.6132
R20225 gnd.n4372 gnd.n3366 4.46168
R20226 gnd.n4556 gnd.n4554 4.46168
R20227 gnd.n4573 gnd.n3208 4.46168
R20228 gnd.n4587 gnd.t230 4.46168
R20229 gnd.n4655 gnd.n3148 4.46168
R20230 gnd.n4696 gnd.n3127 4.46168
R20231 gnd.n4849 gnd.n3055 4.46168
R20232 gnd.n4871 gnd.n3038 4.46168
R20233 gnd.n5128 gnd.n2885 4.46168
R20234 gnd.n5927 gnd.n2745 4.46168
R20235 gnd.n2905 gnd.n2892 4.46111
R20236 gnd.n2159 gnd.n2155 4.38594
R20237 gnd.n2127 gnd.n2123 4.38594
R20238 gnd.n2095 gnd.n2091 4.38594
R20239 gnd.n2064 gnd.n2060 4.38594
R20240 gnd.n2032 gnd.n2028 4.38594
R20241 gnd.n2000 gnd.n1996 4.38594
R20242 gnd.n1968 gnd.n1964 4.38594
R20243 gnd.n1937 gnd.n1933 4.38594
R20244 gnd.n2170 gnd.n2148 4.26717
R20245 gnd.n2138 gnd.n2116 4.26717
R20246 gnd.n2106 gnd.n2084 4.26717
R20247 gnd.n2075 gnd.n2053 4.26717
R20248 gnd.n2043 gnd.n2021 4.26717
R20249 gnd.n2011 gnd.n1989 4.26717
R20250 gnd.n1979 gnd.n1957 4.26717
R20251 gnd.n1948 gnd.n1926 4.26717
R20252 gnd.n1626 gnd.t306 4.14303
R20253 gnd.n1858 gnd.t304 4.14303
R20254 gnd.t36 gnd.n2484 4.14303
R20255 gnd.n5515 gnd.t11 4.14303
R20256 gnd.n2178 gnd.n2177 4.08274
R20257 gnd.n5057 gnd.n5056 4.05904
R20258 gnd.n3353 gnd.n3352 4.05904
R20259 gnd.n4494 gnd.n3285 4.05904
R20260 gnd.n5074 gnd.n5073 4.05904
R20261 gnd.n15 gnd.n7 3.99943
R20262 gnd.n1699 gnd.n1120 3.86464
R20263 gnd.n1107 gnd.n1095 3.72967
R20264 gnd.n50 gnd.n38 3.72967
R20265 gnd.n2178 gnd.n2050 3.70378
R20266 gnd.n15 gnd.n14 3.60163
R20267 gnd.n4546 gnd.n3248 3.50571
R20268 gnd.n5136 gnd.n2877 3.50571
R20269 gnd.n2169 gnd.n2150 3.49141
R20270 gnd.n2137 gnd.n2118 3.49141
R20271 gnd.n2105 gnd.n2086 3.49141
R20272 gnd.n2074 gnd.n2055 3.49141
R20273 gnd.n2042 gnd.n2023 3.49141
R20274 gnd.n2010 gnd.n1991 3.49141
R20275 gnd.n1978 gnd.n1959 3.49141
R20276 gnd.n1947 gnd.n1928 3.49141
R20277 gnd.n5892 gnd.n5891 3.29747
R20278 gnd.n5891 gnd.n5890 3.29747
R20279 gnd.n7297 gnd.n7294 3.29747
R20280 gnd.n7298 gnd.n7297 3.29747
R20281 gnd.n4000 gnd.n3941 3.29747
R20282 gnd.n3941 gnd.n3936 3.29747
R20283 gnd.n4340 gnd.n4339 3.29747
R20284 gnd.n4339 gnd.n4338 3.29747
R20285 gnd.n3281 gnd.t187 3.18706
R20286 gnd.n4594 gnd.n3198 3.18706
R20287 gnd.n4662 gnd.n3152 3.18706
R20288 gnd.t165 gnd.n3127 3.18706
R20289 gnd.n4707 gnd.n4706 3.18706
R20290 gnd.n4802 gnd.n3060 3.18706
R20291 gnd.n4849 gnd.t2 3.18706
R20292 gnd.n4881 gnd.n4880 3.18706
R20293 gnd.n4978 gnd.n2983 3.18706
R20294 gnd.n1205 gnd.t306 2.8684
R20295 gnd.n4567 gnd.t160 2.8684
R20296 gnd.t169 gnd.n2969 2.8684
R20297 gnd.n1108 gnd.t53 2.82907
R20298 gnd.n1108 gnd.t114 2.82907
R20299 gnd.n1110 gnd.t32 2.82907
R20300 gnd.n1110 gnd.t67 2.82907
R20301 gnd.n1112 gnd.t85 2.82907
R20302 gnd.n1112 gnd.t74 2.82907
R20303 gnd.n1114 gnd.t71 2.82907
R20304 gnd.n1114 gnd.t62 2.82907
R20305 gnd.n1116 gnd.t72 2.82907
R20306 gnd.n1116 gnd.t103 2.82907
R20307 gnd.n1073 gnd.t78 2.82907
R20308 gnd.n1073 gnd.t93 2.82907
R20309 gnd.n1075 gnd.t100 2.82907
R20310 gnd.n1075 gnd.t56 2.82907
R20311 gnd.n1077 gnd.t92 2.82907
R20312 gnd.n1077 gnd.t89 2.82907
R20313 gnd.n1079 gnd.t125 2.82907
R20314 gnd.n1079 gnd.t116 2.82907
R20315 gnd.n1081 gnd.t61 2.82907
R20316 gnd.n1081 gnd.t97 2.82907
R20317 gnd.n1084 gnd.t128 2.82907
R20318 gnd.n1084 gnd.t37 2.82907
R20319 gnd.n1086 gnd.t38 2.82907
R20320 gnd.n1086 gnd.t21 2.82907
R20321 gnd.n1088 gnd.t102 2.82907
R20322 gnd.n1088 gnd.t129 2.82907
R20323 gnd.n1090 gnd.t123 2.82907
R20324 gnd.n1090 gnd.t40 2.82907
R20325 gnd.n1092 gnd.t117 2.82907
R20326 gnd.n1092 gnd.t101 2.82907
R20327 gnd.n1096 gnd.t90 2.82907
R20328 gnd.n1096 gnd.t57 2.82907
R20329 gnd.n1098 gnd.t77 2.82907
R20330 gnd.n1098 gnd.t105 2.82907
R20331 gnd.n1100 gnd.t122 2.82907
R20332 gnd.n1100 gnd.t111 2.82907
R20333 gnd.n1102 gnd.t110 2.82907
R20334 gnd.n1102 gnd.t96 2.82907
R20335 gnd.n1104 gnd.t113 2.82907
R20336 gnd.n1104 gnd.t47 2.82907
R20337 gnd.n59 gnd.t81 2.82907
R20338 gnd.n59 gnd.t55 2.82907
R20339 gnd.n57 gnd.t29 2.82907
R20340 gnd.n57 gnd.t45 2.82907
R20341 gnd.n55 gnd.t49 2.82907
R20342 gnd.n55 gnd.t64 2.82907
R20343 gnd.n53 gnd.t42 2.82907
R20344 gnd.n53 gnd.t99 2.82907
R20345 gnd.n51 gnd.t79 2.82907
R20346 gnd.n51 gnd.t25 2.82907
R20347 gnd.n24 gnd.t130 2.82907
R20348 gnd.n24 gnd.t51 2.82907
R20349 gnd.n22 gnd.t35 2.82907
R20350 gnd.n22 gnd.t50 2.82907
R20351 gnd.n20 gnd.t109 2.82907
R20352 gnd.n20 gnd.t86 2.82907
R20353 gnd.n18 gnd.t76 2.82907
R20354 gnd.n18 gnd.t19 2.82907
R20355 gnd.n16 gnd.t121 2.82907
R20356 gnd.n16 gnd.t65 2.82907
R20357 gnd.n35 gnd.t91 2.82907
R20358 gnd.n35 gnd.t18 2.82907
R20359 gnd.n33 gnd.t14 2.82907
R20360 gnd.n33 gnd.t106 2.82907
R20361 gnd.n31 gnd.t112 2.82907
R20362 gnd.n31 gnd.t119 2.82907
R20363 gnd.n29 gnd.t118 2.82907
R20364 gnd.n29 gnd.t16 2.82907
R20365 gnd.n27 gnd.t12 2.82907
R20366 gnd.n27 gnd.t30 2.82907
R20367 gnd.n47 gnd.t120 2.82907
R20368 gnd.n47 gnd.t95 2.82907
R20369 gnd.n45 gnd.t75 2.82907
R20370 gnd.n45 gnd.t87 2.82907
R20371 gnd.n43 gnd.t88 2.82907
R20372 gnd.n43 gnd.t98 2.82907
R20373 gnd.n41 gnd.t82 2.82907
R20374 gnd.n41 gnd.t54 2.82907
R20375 gnd.n39 gnd.t127 2.82907
R20376 gnd.n39 gnd.t69 2.82907
R20377 gnd.n2166 gnd.n2165 2.71565
R20378 gnd.n2134 gnd.n2133 2.71565
R20379 gnd.n2102 gnd.n2101 2.71565
R20380 gnd.n2071 gnd.n2070 2.71565
R20381 gnd.n2039 gnd.n2038 2.71565
R20382 gnd.n2007 gnd.n2006 2.71565
R20383 gnd.n1975 gnd.n1974 2.71565
R20384 gnd.n1944 gnd.n1943 2.71565
R20385 gnd.n3494 gnd.t230 2.54975
R20386 gnd.t5 gnd.n4626 2.54975
R20387 gnd.n4940 gnd.t4 2.54975
R20388 gnd.n4971 gnd.t289 2.54975
R20389 gnd.n1699 gnd.n1121 2.27742
R20390 gnd.n1699 gnd.n1072 2.27742
R20391 gnd.n1699 gnd.n1071 2.27742
R20392 gnd.n1699 gnd.n1070 2.27742
R20393 gnd.n7397 gnd.n81 2.27742
R20394 gnd.n7397 gnd.n80 2.27742
R20395 gnd.n7397 gnd.n79 2.27742
R20396 gnd.n7397 gnd.n74 2.27742
R20397 gnd.n7398 gnd.n7397 2.27742
R20398 gnd.n5557 gnd.n78 2.27742
R20399 gnd.n5747 gnd.n78 2.27742
R20400 gnd.n5411 gnd.n78 2.27742
R20401 gnd.n5595 gnd.n78 2.27742
R20402 gnd.n5725 gnd.n78 2.27742
R20403 gnd.n6164 gnd.n2413 2.27742
R20404 gnd.n2414 gnd.n2413 2.27742
R20405 gnd.n6151 gnd.n2413 2.27742
R20406 gnd.n2432 gnd.n2413 2.27742
R20407 gnd.n6138 gnd.n2413 2.27742
R20408 gnd.n3795 gnd.n3794 2.27742
R20409 gnd.n3794 gnd.n3793 2.27742
R20410 gnd.n3794 gnd.n3767 2.27742
R20411 gnd.n3794 gnd.n3766 2.27742
R20412 gnd.n3794 gnd.n3765 2.27742
R20413 gnd.n1553 gnd.t285 2.23109
R20414 gnd.n1176 gnd.t301 2.23109
R20415 gnd.n4696 gnd.t313 2.23109
R20416 gnd.t162 gnd.n3055 2.23109
R20417 gnd.n2162 gnd.n2152 1.93989
R20418 gnd.n2130 gnd.n2120 1.93989
R20419 gnd.n2098 gnd.n2088 1.93989
R20420 gnd.n2067 gnd.n2057 1.93989
R20421 gnd.n2035 gnd.n2025 1.93989
R20422 gnd.n2003 gnd.n1993 1.93989
R20423 gnd.n1971 gnd.n1961 1.93989
R20424 gnd.n1940 gnd.n1930 1.93989
R20425 gnd.n3289 gnd.t249 1.91244
R20426 gnd.n4608 gnd.n4607 1.91244
R20427 gnd.n4644 gnd.n3157 1.91244
R20428 gnd.n4740 gnd.n4739 1.91244
R20429 gnd.n4737 gnd.t138 1.91244
R20430 gnd.t317 gnd.n3076 1.91244
R20431 gnd.n4792 gnd.n4791 1.91244
R20432 gnd.n3026 gnd.n3025 1.91244
R20433 gnd.n4958 gnd.n2988 1.91244
R20434 gnd.t289 gnd.n2979 1.91244
R20435 gnd.t307 gnd.n1564 1.59378
R20436 gnd.n1743 gnd.t298 1.59378
R20437 gnd.n1006 gnd.t143 1.59378
R20438 gnd.t139 gnd.n3189 1.59378
R20439 gnd.n4965 gnd.t311 1.59378
R20440 gnd.n4573 gnd.t172 1.27512
R20441 gnd.n4971 gnd.t208 1.27512
R20442 gnd.n5136 gnd.t264 1.27512
R20443 gnd.n1406 gnd.n1398 1.16414
R20444 gnd.n2224 gnd.n909 1.16414
R20445 gnd.n2161 gnd.n2154 1.16414
R20446 gnd.n2129 gnd.n2122 1.16414
R20447 gnd.n2097 gnd.n2090 1.16414
R20448 gnd.n2066 gnd.n2059 1.16414
R20449 gnd.n2034 gnd.n2027 1.16414
R20450 gnd.n2002 gnd.n1995 1.16414
R20451 gnd.n1970 gnd.n1963 1.16414
R20452 gnd.n1939 gnd.n1932 1.16414
R20453 gnd.n5874 gnd.n5873 0.970197
R20454 gnd.n4482 gnd.n3359 0.970197
R20455 gnd.n2145 gnd.n2113 0.962709
R20456 gnd.n2177 gnd.n2145 0.962709
R20457 gnd.n2018 gnd.n1986 0.962709
R20458 gnd.n2050 gnd.n2018 0.962709
R20459 gnd.n1652 gnd.t153 0.956468
R20460 gnd.n1819 gnd.t295 0.956468
R20461 gnd.n4136 gnd.t60 0.956468
R20462 gnd.n4213 gnd.t36 0.956468
R20463 gnd.n3484 gnd.t131 0.956468
R20464 gnd.n2878 gnd.t146 0.956468
R20465 gnd.n5780 gnd.t11 0.956468
R20466 gnd.n5701 gnd.t17 0.956468
R20467 gnd.n2 gnd.n1 0.672012
R20468 gnd.n3 gnd.n2 0.672012
R20469 gnd.n4 gnd.n3 0.672012
R20470 gnd.n5 gnd.n4 0.672012
R20471 gnd.n6 gnd.n5 0.672012
R20472 gnd.n7 gnd.n6 0.672012
R20473 gnd.n9 gnd.n8 0.672012
R20474 gnd.n10 gnd.n9 0.672012
R20475 gnd.n11 gnd.n10 0.672012
R20476 gnd.n12 gnd.n11 0.672012
R20477 gnd.n13 gnd.n12 0.672012
R20478 gnd.n14 gnd.n13 0.672012
R20479 gnd.n4615 gnd.n3179 0.637812
R20480 gnd.n4634 gnd.n4633 0.637812
R20481 gnd.n3104 gnd.n3103 0.637812
R20482 gnd.n3095 gnd.n3083 0.637812
R20483 gnd.n4819 gnd.n4818 0.637812
R20484 gnd.n4948 gnd.n4947 0.637812
R20485 gnd.n1118 gnd.n1117 0.573776
R20486 gnd.n1117 gnd.n1115 0.573776
R20487 gnd.n1115 gnd.n1113 0.573776
R20488 gnd.n1113 gnd.n1111 0.573776
R20489 gnd.n1111 gnd.n1109 0.573776
R20490 gnd.n1083 gnd.n1082 0.573776
R20491 gnd.n1082 gnd.n1080 0.573776
R20492 gnd.n1080 gnd.n1078 0.573776
R20493 gnd.n1078 gnd.n1076 0.573776
R20494 gnd.n1076 gnd.n1074 0.573776
R20495 gnd.n1094 gnd.n1093 0.573776
R20496 gnd.n1093 gnd.n1091 0.573776
R20497 gnd.n1091 gnd.n1089 0.573776
R20498 gnd.n1089 gnd.n1087 0.573776
R20499 gnd.n1087 gnd.n1085 0.573776
R20500 gnd.n1106 gnd.n1105 0.573776
R20501 gnd.n1105 gnd.n1103 0.573776
R20502 gnd.n1103 gnd.n1101 0.573776
R20503 gnd.n1101 gnd.n1099 0.573776
R20504 gnd.n1099 gnd.n1097 0.573776
R20505 gnd.n54 gnd.n52 0.573776
R20506 gnd.n56 gnd.n54 0.573776
R20507 gnd.n58 gnd.n56 0.573776
R20508 gnd.n60 gnd.n58 0.573776
R20509 gnd.n61 gnd.n60 0.573776
R20510 gnd.n19 gnd.n17 0.573776
R20511 gnd.n21 gnd.n19 0.573776
R20512 gnd.n23 gnd.n21 0.573776
R20513 gnd.n25 gnd.n23 0.573776
R20514 gnd.n26 gnd.n25 0.573776
R20515 gnd.n30 gnd.n28 0.573776
R20516 gnd.n32 gnd.n30 0.573776
R20517 gnd.n34 gnd.n32 0.573776
R20518 gnd.n36 gnd.n34 0.573776
R20519 gnd.n37 gnd.n36 0.573776
R20520 gnd.n42 gnd.n40 0.573776
R20521 gnd.n44 gnd.n42 0.573776
R20522 gnd.n46 gnd.n44 0.573776
R20523 gnd.n48 gnd.n46 0.573776
R20524 gnd.n49 gnd.n48 0.573776
R20525 gnd gnd.n0 0.551497
R20526 gnd.n7335 gnd.n7334 0.532512
R20527 gnd.n3853 gnd.n3852 0.532512
R20528 gnd.n7150 gnd.n165 0.497451
R20529 gnd.n4297 gnd.n2530 0.497451
R20530 gnd.n5324 gnd.n2749 0.497451
R20531 gnd.n3956 gnd.n2329 0.497451
R20532 gnd.n5938 gnd.n5937 0.489829
R20533 gnd.n2578 gnd.n2544 0.489829
R20534 gnd.n3580 gnd.n3577 0.489829
R20535 gnd.n5190 gnd.n2836 0.489829
R20536 gnd.n1881 gnd.n913 0.486781
R20537 gnd.n1455 gnd.n1454 0.48678
R20538 gnd.n2198 gnd.n867 0.480683
R20539 gnd.n1539 gnd.n1538 0.480683
R20540 gnd.n7409 gnd.n7408 0.470187
R20541 gnd.n6404 gnd.n6403 0.447146
R20542 gnd.n6894 gnd.n380 0.447146
R20543 gnd.n7105 gnd.n7104 0.447146
R20544 gnd.n2308 gnd.n840 0.447146
R20545 gnd.n7397 gnd.n78 0.4255
R20546 gnd.n3794 gnd.n2413 0.4255
R20547 gnd.n3661 gnd.n3660 0.388379
R20548 gnd.n2158 gnd.n2157 0.388379
R20549 gnd.n2126 gnd.n2125 0.388379
R20550 gnd.n2094 gnd.n2093 0.388379
R20551 gnd.n2063 gnd.n2062 0.388379
R20552 gnd.n2031 gnd.n2030 0.388379
R20553 gnd.n1999 gnd.n1998 0.388379
R20554 gnd.n1967 gnd.n1966 0.388379
R20555 gnd.n1936 gnd.n1935 0.388379
R20556 gnd.n5264 gnd.n5253 0.388379
R20557 gnd.n7409 gnd.n15 0.374463
R20558 gnd.n968 gnd.t293 0.319156
R20559 gnd.n4164 gnd.t39 0.319156
R20560 gnd.n4192 gnd.t31 0.319156
R20561 gnd.t138 gnd.t0 0.319156
R20562 gnd.t134 gnd.t317 0.319156
R20563 gnd.n5756 gnd.t15 0.319156
R20564 gnd.n5610 gnd.t13 0.319156
R20565 gnd.n1373 gnd.n1351 0.311721
R20566 gnd.n6075 gnd.n6074 0.302329
R20567 gnd.n5489 gnd.n2679 0.302329
R20568 gnd gnd.n7409 0.295112
R20569 gnd.n199 gnd.n173 0.293183
R20570 gnd.n4106 gnd.n3893 0.293183
R20571 gnd.n2269 gnd.n2268 0.268793
R20572 gnd.n7211 gnd.n173 0.258122
R20573 gnd.n5812 gnd.n5811 0.258122
R20574 gnd.n4423 gnd.n2538 0.258122
R20575 gnd.n4106 gnd.n4105 0.258122
R20576 gnd.n2268 gnd.n2267 0.241354
R20577 gnd.n2779 gnd.n2776 0.229039
R20578 gnd.n2780 gnd.n2779 0.229039
R20579 gnd.n4481 gnd.n3362 0.229039
R20580 gnd.n4481 gnd.n4480 0.229039
R20581 gnd.n1527 gnd.n1326 0.206293
R20582 gnd.n2175 gnd.n2147 0.155672
R20583 gnd.n2168 gnd.n2147 0.155672
R20584 gnd.n2168 gnd.n2167 0.155672
R20585 gnd.n2167 gnd.n2151 0.155672
R20586 gnd.n2160 gnd.n2151 0.155672
R20587 gnd.n2160 gnd.n2159 0.155672
R20588 gnd.n2143 gnd.n2115 0.155672
R20589 gnd.n2136 gnd.n2115 0.155672
R20590 gnd.n2136 gnd.n2135 0.155672
R20591 gnd.n2135 gnd.n2119 0.155672
R20592 gnd.n2128 gnd.n2119 0.155672
R20593 gnd.n2128 gnd.n2127 0.155672
R20594 gnd.n2111 gnd.n2083 0.155672
R20595 gnd.n2104 gnd.n2083 0.155672
R20596 gnd.n2104 gnd.n2103 0.155672
R20597 gnd.n2103 gnd.n2087 0.155672
R20598 gnd.n2096 gnd.n2087 0.155672
R20599 gnd.n2096 gnd.n2095 0.155672
R20600 gnd.n2080 gnd.n2052 0.155672
R20601 gnd.n2073 gnd.n2052 0.155672
R20602 gnd.n2073 gnd.n2072 0.155672
R20603 gnd.n2072 gnd.n2056 0.155672
R20604 gnd.n2065 gnd.n2056 0.155672
R20605 gnd.n2065 gnd.n2064 0.155672
R20606 gnd.n2048 gnd.n2020 0.155672
R20607 gnd.n2041 gnd.n2020 0.155672
R20608 gnd.n2041 gnd.n2040 0.155672
R20609 gnd.n2040 gnd.n2024 0.155672
R20610 gnd.n2033 gnd.n2024 0.155672
R20611 gnd.n2033 gnd.n2032 0.155672
R20612 gnd.n2016 gnd.n1988 0.155672
R20613 gnd.n2009 gnd.n1988 0.155672
R20614 gnd.n2009 gnd.n2008 0.155672
R20615 gnd.n2008 gnd.n1992 0.155672
R20616 gnd.n2001 gnd.n1992 0.155672
R20617 gnd.n2001 gnd.n2000 0.155672
R20618 gnd.n1984 gnd.n1956 0.155672
R20619 gnd.n1977 gnd.n1956 0.155672
R20620 gnd.n1977 gnd.n1976 0.155672
R20621 gnd.n1976 gnd.n1960 0.155672
R20622 gnd.n1969 gnd.n1960 0.155672
R20623 gnd.n1969 gnd.n1968 0.155672
R20624 gnd.n1953 gnd.n1925 0.155672
R20625 gnd.n1946 gnd.n1925 0.155672
R20626 gnd.n1946 gnd.n1945 0.155672
R20627 gnd.n1945 gnd.n1929 0.155672
R20628 gnd.n1938 gnd.n1929 0.155672
R20629 gnd.n1938 gnd.n1937 0.155672
R20630 gnd.n2300 gnd.n867 0.152939
R20631 gnd.n2300 gnd.n2299 0.152939
R20632 gnd.n2299 gnd.n2298 0.152939
R20633 gnd.n2298 gnd.n869 0.152939
R20634 gnd.n870 gnd.n869 0.152939
R20635 gnd.n871 gnd.n870 0.152939
R20636 gnd.n872 gnd.n871 0.152939
R20637 gnd.n873 gnd.n872 0.152939
R20638 gnd.n874 gnd.n873 0.152939
R20639 gnd.n875 gnd.n874 0.152939
R20640 gnd.n876 gnd.n875 0.152939
R20641 gnd.n877 gnd.n876 0.152939
R20642 gnd.n878 gnd.n877 0.152939
R20643 gnd.n879 gnd.n878 0.152939
R20644 gnd.n2270 gnd.n879 0.152939
R20645 gnd.n2270 gnd.n2269 0.152939
R20646 gnd.n1540 gnd.n1539 0.152939
R20647 gnd.n1540 gnd.n1244 0.152939
R20648 gnd.n1568 gnd.n1244 0.152939
R20649 gnd.n1569 gnd.n1568 0.152939
R20650 gnd.n1570 gnd.n1569 0.152939
R20651 gnd.n1571 gnd.n1570 0.152939
R20652 gnd.n1571 gnd.n1216 0.152939
R20653 gnd.n1598 gnd.n1216 0.152939
R20654 gnd.n1599 gnd.n1598 0.152939
R20655 gnd.n1600 gnd.n1599 0.152939
R20656 gnd.n1600 gnd.n1194 0.152939
R20657 gnd.n1629 gnd.n1194 0.152939
R20658 gnd.n1630 gnd.n1629 0.152939
R20659 gnd.n1631 gnd.n1630 0.152939
R20660 gnd.n1632 gnd.n1631 0.152939
R20661 gnd.n1634 gnd.n1632 0.152939
R20662 gnd.n1634 gnd.n1633 0.152939
R20663 gnd.n1633 gnd.n1143 0.152939
R20664 gnd.n1144 gnd.n1143 0.152939
R20665 gnd.n1145 gnd.n1144 0.152939
R20666 gnd.n1164 gnd.n1145 0.152939
R20667 gnd.n1165 gnd.n1164 0.152939
R20668 gnd.n1165 gnd.n1063 0.152939
R20669 gnd.n1724 gnd.n1063 0.152939
R20670 gnd.n1725 gnd.n1724 0.152939
R20671 gnd.n1726 gnd.n1725 0.152939
R20672 gnd.n1727 gnd.n1726 0.152939
R20673 gnd.n1727 gnd.n1036 0.152939
R20674 gnd.n1764 gnd.n1036 0.152939
R20675 gnd.n1765 gnd.n1764 0.152939
R20676 gnd.n1766 gnd.n1765 0.152939
R20677 gnd.n1767 gnd.n1766 0.152939
R20678 gnd.n1767 gnd.n1010 0.152939
R20679 gnd.n1811 gnd.n1010 0.152939
R20680 gnd.n1812 gnd.n1811 0.152939
R20681 gnd.n1813 gnd.n1812 0.152939
R20682 gnd.n1814 gnd.n1813 0.152939
R20683 gnd.n1814 gnd.n982 0.152939
R20684 gnd.n1851 gnd.n982 0.152939
R20685 gnd.n1852 gnd.n1851 0.152939
R20686 gnd.n1853 gnd.n1852 0.152939
R20687 gnd.n1854 gnd.n1853 0.152939
R20688 gnd.n1854 gnd.n955 0.152939
R20689 gnd.n1900 gnd.n955 0.152939
R20690 gnd.n1901 gnd.n1900 0.152939
R20691 gnd.n1902 gnd.n1901 0.152939
R20692 gnd.n1903 gnd.n1902 0.152939
R20693 gnd.n1903 gnd.n928 0.152939
R20694 gnd.n2194 gnd.n928 0.152939
R20695 gnd.n2195 gnd.n2194 0.152939
R20696 gnd.n2196 gnd.n2195 0.152939
R20697 gnd.n2197 gnd.n2196 0.152939
R20698 gnd.n2198 gnd.n2197 0.152939
R20699 gnd.n1538 gnd.n1268 0.152939
R20700 gnd.n1289 gnd.n1268 0.152939
R20701 gnd.n1290 gnd.n1289 0.152939
R20702 gnd.n1296 gnd.n1290 0.152939
R20703 gnd.n1297 gnd.n1296 0.152939
R20704 gnd.n1298 gnd.n1297 0.152939
R20705 gnd.n1298 gnd.n1287 0.152939
R20706 gnd.n1306 gnd.n1287 0.152939
R20707 gnd.n1307 gnd.n1306 0.152939
R20708 gnd.n1308 gnd.n1307 0.152939
R20709 gnd.n1308 gnd.n1285 0.152939
R20710 gnd.n1316 gnd.n1285 0.152939
R20711 gnd.n1317 gnd.n1316 0.152939
R20712 gnd.n1318 gnd.n1317 0.152939
R20713 gnd.n1318 gnd.n1283 0.152939
R20714 gnd.n1326 gnd.n1283 0.152939
R20715 gnd.n2267 gnd.n884 0.152939
R20716 gnd.n886 gnd.n884 0.152939
R20717 gnd.n887 gnd.n886 0.152939
R20718 gnd.n888 gnd.n887 0.152939
R20719 gnd.n889 gnd.n888 0.152939
R20720 gnd.n890 gnd.n889 0.152939
R20721 gnd.n891 gnd.n890 0.152939
R20722 gnd.n892 gnd.n891 0.152939
R20723 gnd.n893 gnd.n892 0.152939
R20724 gnd.n894 gnd.n893 0.152939
R20725 gnd.n895 gnd.n894 0.152939
R20726 gnd.n896 gnd.n895 0.152939
R20727 gnd.n897 gnd.n896 0.152939
R20728 gnd.n898 gnd.n897 0.152939
R20729 gnd.n899 gnd.n898 0.152939
R20730 gnd.n900 gnd.n899 0.152939
R20731 gnd.n901 gnd.n900 0.152939
R20732 gnd.n902 gnd.n901 0.152939
R20733 gnd.n903 gnd.n902 0.152939
R20734 gnd.n904 gnd.n903 0.152939
R20735 gnd.n905 gnd.n904 0.152939
R20736 gnd.n906 gnd.n905 0.152939
R20737 gnd.n910 gnd.n906 0.152939
R20738 gnd.n911 gnd.n910 0.152939
R20739 gnd.n912 gnd.n911 0.152939
R20740 gnd.n913 gnd.n912 0.152939
R20741 gnd.n1701 gnd.n1700 0.152939
R20742 gnd.n1702 gnd.n1701 0.152939
R20743 gnd.n1703 gnd.n1702 0.152939
R20744 gnd.n1704 gnd.n1703 0.152939
R20745 gnd.n1705 gnd.n1704 0.152939
R20746 gnd.n1706 gnd.n1705 0.152939
R20747 gnd.n1706 gnd.n1017 0.152939
R20748 gnd.n1785 gnd.n1017 0.152939
R20749 gnd.n1786 gnd.n1785 0.152939
R20750 gnd.n1787 gnd.n1786 0.152939
R20751 gnd.n1788 gnd.n1787 0.152939
R20752 gnd.n1789 gnd.n1788 0.152939
R20753 gnd.n1790 gnd.n1789 0.152939
R20754 gnd.n1791 gnd.n1790 0.152939
R20755 gnd.n1792 gnd.n1791 0.152939
R20756 gnd.n1793 gnd.n1792 0.152939
R20757 gnd.n1793 gnd.n962 0.152939
R20758 gnd.n1872 gnd.n962 0.152939
R20759 gnd.n1873 gnd.n1872 0.152939
R20760 gnd.n1874 gnd.n1873 0.152939
R20761 gnd.n1875 gnd.n1874 0.152939
R20762 gnd.n1876 gnd.n1875 0.152939
R20763 gnd.n1877 gnd.n1876 0.152939
R20764 gnd.n1878 gnd.n1877 0.152939
R20765 gnd.n1879 gnd.n1878 0.152939
R20766 gnd.n1880 gnd.n1879 0.152939
R20767 gnd.n1882 gnd.n1880 0.152939
R20768 gnd.n1882 gnd.n1881 0.152939
R20769 gnd.n1456 gnd.n1455 0.152939
R20770 gnd.n1456 gnd.n1346 0.152939
R20771 gnd.n1471 gnd.n1346 0.152939
R20772 gnd.n1472 gnd.n1471 0.152939
R20773 gnd.n1473 gnd.n1472 0.152939
R20774 gnd.n1473 gnd.n1334 0.152939
R20775 gnd.n1487 gnd.n1334 0.152939
R20776 gnd.n1488 gnd.n1487 0.152939
R20777 gnd.n1489 gnd.n1488 0.152939
R20778 gnd.n1490 gnd.n1489 0.152939
R20779 gnd.n1491 gnd.n1490 0.152939
R20780 gnd.n1492 gnd.n1491 0.152939
R20781 gnd.n1493 gnd.n1492 0.152939
R20782 gnd.n1494 gnd.n1493 0.152939
R20783 gnd.n1495 gnd.n1494 0.152939
R20784 gnd.n1496 gnd.n1495 0.152939
R20785 gnd.n1497 gnd.n1496 0.152939
R20786 gnd.n1498 gnd.n1497 0.152939
R20787 gnd.n1499 gnd.n1498 0.152939
R20788 gnd.n1500 gnd.n1499 0.152939
R20789 gnd.n1501 gnd.n1500 0.152939
R20790 gnd.n1501 gnd.n1200 0.152939
R20791 gnd.n1618 gnd.n1200 0.152939
R20792 gnd.n1619 gnd.n1618 0.152939
R20793 gnd.n1620 gnd.n1619 0.152939
R20794 gnd.n1621 gnd.n1620 0.152939
R20795 gnd.n1621 gnd.n1122 0.152939
R20796 gnd.n1698 gnd.n1122 0.152939
R20797 gnd.n1374 gnd.n1373 0.152939
R20798 gnd.n1375 gnd.n1374 0.152939
R20799 gnd.n1376 gnd.n1375 0.152939
R20800 gnd.n1377 gnd.n1376 0.152939
R20801 gnd.n1378 gnd.n1377 0.152939
R20802 gnd.n1379 gnd.n1378 0.152939
R20803 gnd.n1380 gnd.n1379 0.152939
R20804 gnd.n1381 gnd.n1380 0.152939
R20805 gnd.n1382 gnd.n1381 0.152939
R20806 gnd.n1383 gnd.n1382 0.152939
R20807 gnd.n1384 gnd.n1383 0.152939
R20808 gnd.n1385 gnd.n1384 0.152939
R20809 gnd.n1386 gnd.n1385 0.152939
R20810 gnd.n1387 gnd.n1386 0.152939
R20811 gnd.n1388 gnd.n1387 0.152939
R20812 gnd.n1389 gnd.n1388 0.152939
R20813 gnd.n1390 gnd.n1389 0.152939
R20814 gnd.n1391 gnd.n1390 0.152939
R20815 gnd.n1392 gnd.n1391 0.152939
R20816 gnd.n1393 gnd.n1392 0.152939
R20817 gnd.n1394 gnd.n1393 0.152939
R20818 gnd.n1395 gnd.n1394 0.152939
R20819 gnd.n1399 gnd.n1395 0.152939
R20820 gnd.n1400 gnd.n1399 0.152939
R20821 gnd.n1400 gnd.n1357 0.152939
R20822 gnd.n1454 gnd.n1357 0.152939
R20823 gnd.n6405 gnd.n6404 0.152939
R20824 gnd.n6405 gnd.n667 0.152939
R20825 gnd.n6413 gnd.n667 0.152939
R20826 gnd.n6414 gnd.n6413 0.152939
R20827 gnd.n6415 gnd.n6414 0.152939
R20828 gnd.n6415 gnd.n661 0.152939
R20829 gnd.n6423 gnd.n661 0.152939
R20830 gnd.n6424 gnd.n6423 0.152939
R20831 gnd.n6425 gnd.n6424 0.152939
R20832 gnd.n6425 gnd.n655 0.152939
R20833 gnd.n6433 gnd.n655 0.152939
R20834 gnd.n6434 gnd.n6433 0.152939
R20835 gnd.n6435 gnd.n6434 0.152939
R20836 gnd.n6435 gnd.n649 0.152939
R20837 gnd.n6443 gnd.n649 0.152939
R20838 gnd.n6444 gnd.n6443 0.152939
R20839 gnd.n6445 gnd.n6444 0.152939
R20840 gnd.n6445 gnd.n643 0.152939
R20841 gnd.n6453 gnd.n643 0.152939
R20842 gnd.n6454 gnd.n6453 0.152939
R20843 gnd.n6455 gnd.n6454 0.152939
R20844 gnd.n6455 gnd.n637 0.152939
R20845 gnd.n6463 gnd.n637 0.152939
R20846 gnd.n6464 gnd.n6463 0.152939
R20847 gnd.n6465 gnd.n6464 0.152939
R20848 gnd.n6465 gnd.n631 0.152939
R20849 gnd.n6473 gnd.n631 0.152939
R20850 gnd.n6474 gnd.n6473 0.152939
R20851 gnd.n6475 gnd.n6474 0.152939
R20852 gnd.n6475 gnd.n625 0.152939
R20853 gnd.n6483 gnd.n625 0.152939
R20854 gnd.n6484 gnd.n6483 0.152939
R20855 gnd.n6485 gnd.n6484 0.152939
R20856 gnd.n6485 gnd.n619 0.152939
R20857 gnd.n6493 gnd.n619 0.152939
R20858 gnd.n6494 gnd.n6493 0.152939
R20859 gnd.n6495 gnd.n6494 0.152939
R20860 gnd.n6495 gnd.n613 0.152939
R20861 gnd.n6503 gnd.n613 0.152939
R20862 gnd.n6504 gnd.n6503 0.152939
R20863 gnd.n6505 gnd.n6504 0.152939
R20864 gnd.n6505 gnd.n607 0.152939
R20865 gnd.n6513 gnd.n607 0.152939
R20866 gnd.n6514 gnd.n6513 0.152939
R20867 gnd.n6515 gnd.n6514 0.152939
R20868 gnd.n6515 gnd.n601 0.152939
R20869 gnd.n6523 gnd.n601 0.152939
R20870 gnd.n6524 gnd.n6523 0.152939
R20871 gnd.n6525 gnd.n6524 0.152939
R20872 gnd.n6525 gnd.n595 0.152939
R20873 gnd.n6533 gnd.n595 0.152939
R20874 gnd.n6534 gnd.n6533 0.152939
R20875 gnd.n6535 gnd.n6534 0.152939
R20876 gnd.n6535 gnd.n589 0.152939
R20877 gnd.n6543 gnd.n589 0.152939
R20878 gnd.n6544 gnd.n6543 0.152939
R20879 gnd.n6545 gnd.n6544 0.152939
R20880 gnd.n6545 gnd.n583 0.152939
R20881 gnd.n6553 gnd.n583 0.152939
R20882 gnd.n6554 gnd.n6553 0.152939
R20883 gnd.n6555 gnd.n6554 0.152939
R20884 gnd.n6555 gnd.n577 0.152939
R20885 gnd.n6563 gnd.n577 0.152939
R20886 gnd.n6564 gnd.n6563 0.152939
R20887 gnd.n6565 gnd.n6564 0.152939
R20888 gnd.n6565 gnd.n571 0.152939
R20889 gnd.n6573 gnd.n571 0.152939
R20890 gnd.n6574 gnd.n6573 0.152939
R20891 gnd.n6575 gnd.n6574 0.152939
R20892 gnd.n6575 gnd.n565 0.152939
R20893 gnd.n6583 gnd.n565 0.152939
R20894 gnd.n6584 gnd.n6583 0.152939
R20895 gnd.n6585 gnd.n6584 0.152939
R20896 gnd.n6585 gnd.n559 0.152939
R20897 gnd.n6593 gnd.n559 0.152939
R20898 gnd.n6594 gnd.n6593 0.152939
R20899 gnd.n6595 gnd.n6594 0.152939
R20900 gnd.n6595 gnd.n553 0.152939
R20901 gnd.n6603 gnd.n553 0.152939
R20902 gnd.n6604 gnd.n6603 0.152939
R20903 gnd.n6605 gnd.n6604 0.152939
R20904 gnd.n6605 gnd.n547 0.152939
R20905 gnd.n6613 gnd.n547 0.152939
R20906 gnd.n6614 gnd.n6613 0.152939
R20907 gnd.n6615 gnd.n6614 0.152939
R20908 gnd.n6615 gnd.n541 0.152939
R20909 gnd.n6623 gnd.n541 0.152939
R20910 gnd.n6624 gnd.n6623 0.152939
R20911 gnd.n6625 gnd.n6624 0.152939
R20912 gnd.n6625 gnd.n535 0.152939
R20913 gnd.n6633 gnd.n535 0.152939
R20914 gnd.n6634 gnd.n6633 0.152939
R20915 gnd.n6635 gnd.n6634 0.152939
R20916 gnd.n6635 gnd.n529 0.152939
R20917 gnd.n6643 gnd.n529 0.152939
R20918 gnd.n6644 gnd.n6643 0.152939
R20919 gnd.n6645 gnd.n6644 0.152939
R20920 gnd.n6645 gnd.n523 0.152939
R20921 gnd.n6653 gnd.n523 0.152939
R20922 gnd.n6654 gnd.n6653 0.152939
R20923 gnd.n6655 gnd.n6654 0.152939
R20924 gnd.n6655 gnd.n517 0.152939
R20925 gnd.n6663 gnd.n517 0.152939
R20926 gnd.n6664 gnd.n6663 0.152939
R20927 gnd.n6665 gnd.n6664 0.152939
R20928 gnd.n6665 gnd.n511 0.152939
R20929 gnd.n6673 gnd.n511 0.152939
R20930 gnd.n6674 gnd.n6673 0.152939
R20931 gnd.n6675 gnd.n6674 0.152939
R20932 gnd.n6675 gnd.n505 0.152939
R20933 gnd.n6683 gnd.n505 0.152939
R20934 gnd.n6684 gnd.n6683 0.152939
R20935 gnd.n6685 gnd.n6684 0.152939
R20936 gnd.n6685 gnd.n499 0.152939
R20937 gnd.n6693 gnd.n499 0.152939
R20938 gnd.n6694 gnd.n6693 0.152939
R20939 gnd.n6695 gnd.n6694 0.152939
R20940 gnd.n6695 gnd.n493 0.152939
R20941 gnd.n6703 gnd.n493 0.152939
R20942 gnd.n6704 gnd.n6703 0.152939
R20943 gnd.n6705 gnd.n6704 0.152939
R20944 gnd.n6705 gnd.n487 0.152939
R20945 gnd.n6713 gnd.n487 0.152939
R20946 gnd.n6714 gnd.n6713 0.152939
R20947 gnd.n6715 gnd.n6714 0.152939
R20948 gnd.n6715 gnd.n481 0.152939
R20949 gnd.n6723 gnd.n481 0.152939
R20950 gnd.n6724 gnd.n6723 0.152939
R20951 gnd.n6725 gnd.n6724 0.152939
R20952 gnd.n6725 gnd.n475 0.152939
R20953 gnd.n6733 gnd.n475 0.152939
R20954 gnd.n6734 gnd.n6733 0.152939
R20955 gnd.n6735 gnd.n6734 0.152939
R20956 gnd.n6735 gnd.n469 0.152939
R20957 gnd.n6743 gnd.n469 0.152939
R20958 gnd.n6744 gnd.n6743 0.152939
R20959 gnd.n6745 gnd.n6744 0.152939
R20960 gnd.n6745 gnd.n463 0.152939
R20961 gnd.n6753 gnd.n463 0.152939
R20962 gnd.n6754 gnd.n6753 0.152939
R20963 gnd.n6755 gnd.n6754 0.152939
R20964 gnd.n6755 gnd.n457 0.152939
R20965 gnd.n6763 gnd.n457 0.152939
R20966 gnd.n6764 gnd.n6763 0.152939
R20967 gnd.n6765 gnd.n6764 0.152939
R20968 gnd.n6765 gnd.n451 0.152939
R20969 gnd.n6773 gnd.n451 0.152939
R20970 gnd.n6774 gnd.n6773 0.152939
R20971 gnd.n6775 gnd.n6774 0.152939
R20972 gnd.n6775 gnd.n445 0.152939
R20973 gnd.n6783 gnd.n445 0.152939
R20974 gnd.n6784 gnd.n6783 0.152939
R20975 gnd.n6785 gnd.n6784 0.152939
R20976 gnd.n6785 gnd.n439 0.152939
R20977 gnd.n6793 gnd.n439 0.152939
R20978 gnd.n6794 gnd.n6793 0.152939
R20979 gnd.n6795 gnd.n6794 0.152939
R20980 gnd.n6795 gnd.n433 0.152939
R20981 gnd.n6803 gnd.n433 0.152939
R20982 gnd.n6804 gnd.n6803 0.152939
R20983 gnd.n6805 gnd.n6804 0.152939
R20984 gnd.n6805 gnd.n427 0.152939
R20985 gnd.n6813 gnd.n427 0.152939
R20986 gnd.n6814 gnd.n6813 0.152939
R20987 gnd.n6815 gnd.n6814 0.152939
R20988 gnd.n6815 gnd.n421 0.152939
R20989 gnd.n6823 gnd.n421 0.152939
R20990 gnd.n6824 gnd.n6823 0.152939
R20991 gnd.n6825 gnd.n6824 0.152939
R20992 gnd.n6825 gnd.n415 0.152939
R20993 gnd.n6833 gnd.n415 0.152939
R20994 gnd.n6834 gnd.n6833 0.152939
R20995 gnd.n6835 gnd.n6834 0.152939
R20996 gnd.n6835 gnd.n409 0.152939
R20997 gnd.n6843 gnd.n409 0.152939
R20998 gnd.n6844 gnd.n6843 0.152939
R20999 gnd.n6845 gnd.n6844 0.152939
R21000 gnd.n6845 gnd.n403 0.152939
R21001 gnd.n6853 gnd.n403 0.152939
R21002 gnd.n6854 gnd.n6853 0.152939
R21003 gnd.n6855 gnd.n6854 0.152939
R21004 gnd.n6855 gnd.n397 0.152939
R21005 gnd.n6863 gnd.n397 0.152939
R21006 gnd.n6864 gnd.n6863 0.152939
R21007 gnd.n6865 gnd.n6864 0.152939
R21008 gnd.n6865 gnd.n391 0.152939
R21009 gnd.n6873 gnd.n391 0.152939
R21010 gnd.n6874 gnd.n6873 0.152939
R21011 gnd.n6875 gnd.n6874 0.152939
R21012 gnd.n6875 gnd.n385 0.152939
R21013 gnd.n6883 gnd.n385 0.152939
R21014 gnd.n6884 gnd.n6883 0.152939
R21015 gnd.n6885 gnd.n6884 0.152939
R21016 gnd.n6885 gnd.n380 0.152939
R21017 gnd.n6895 gnd.n6894 0.152939
R21018 gnd.n6896 gnd.n6895 0.152939
R21019 gnd.n6896 gnd.n374 0.152939
R21020 gnd.n6904 gnd.n374 0.152939
R21021 gnd.n6905 gnd.n6904 0.152939
R21022 gnd.n6906 gnd.n6905 0.152939
R21023 gnd.n6906 gnd.n368 0.152939
R21024 gnd.n6914 gnd.n368 0.152939
R21025 gnd.n6915 gnd.n6914 0.152939
R21026 gnd.n6916 gnd.n6915 0.152939
R21027 gnd.n6916 gnd.n362 0.152939
R21028 gnd.n6924 gnd.n362 0.152939
R21029 gnd.n6925 gnd.n6924 0.152939
R21030 gnd.n6926 gnd.n6925 0.152939
R21031 gnd.n6926 gnd.n356 0.152939
R21032 gnd.n6934 gnd.n356 0.152939
R21033 gnd.n6935 gnd.n6934 0.152939
R21034 gnd.n6936 gnd.n6935 0.152939
R21035 gnd.n6936 gnd.n350 0.152939
R21036 gnd.n6944 gnd.n350 0.152939
R21037 gnd.n6945 gnd.n6944 0.152939
R21038 gnd.n6946 gnd.n6945 0.152939
R21039 gnd.n6946 gnd.n344 0.152939
R21040 gnd.n6954 gnd.n344 0.152939
R21041 gnd.n6955 gnd.n6954 0.152939
R21042 gnd.n6956 gnd.n6955 0.152939
R21043 gnd.n6956 gnd.n338 0.152939
R21044 gnd.n6964 gnd.n338 0.152939
R21045 gnd.n6965 gnd.n6964 0.152939
R21046 gnd.n6966 gnd.n6965 0.152939
R21047 gnd.n6966 gnd.n332 0.152939
R21048 gnd.n6974 gnd.n332 0.152939
R21049 gnd.n6975 gnd.n6974 0.152939
R21050 gnd.n6976 gnd.n6975 0.152939
R21051 gnd.n6976 gnd.n326 0.152939
R21052 gnd.n6984 gnd.n326 0.152939
R21053 gnd.n6985 gnd.n6984 0.152939
R21054 gnd.n6986 gnd.n6985 0.152939
R21055 gnd.n6986 gnd.n320 0.152939
R21056 gnd.n6994 gnd.n320 0.152939
R21057 gnd.n6995 gnd.n6994 0.152939
R21058 gnd.n6996 gnd.n6995 0.152939
R21059 gnd.n6996 gnd.n314 0.152939
R21060 gnd.n7004 gnd.n314 0.152939
R21061 gnd.n7005 gnd.n7004 0.152939
R21062 gnd.n7006 gnd.n7005 0.152939
R21063 gnd.n7006 gnd.n308 0.152939
R21064 gnd.n7014 gnd.n308 0.152939
R21065 gnd.n7015 gnd.n7014 0.152939
R21066 gnd.n7016 gnd.n7015 0.152939
R21067 gnd.n7016 gnd.n302 0.152939
R21068 gnd.n7024 gnd.n302 0.152939
R21069 gnd.n7025 gnd.n7024 0.152939
R21070 gnd.n7026 gnd.n7025 0.152939
R21071 gnd.n7026 gnd.n296 0.152939
R21072 gnd.n7034 gnd.n296 0.152939
R21073 gnd.n7035 gnd.n7034 0.152939
R21074 gnd.n7036 gnd.n7035 0.152939
R21075 gnd.n7036 gnd.n290 0.152939
R21076 gnd.n7044 gnd.n290 0.152939
R21077 gnd.n7045 gnd.n7044 0.152939
R21078 gnd.n7046 gnd.n7045 0.152939
R21079 gnd.n7046 gnd.n284 0.152939
R21080 gnd.n7054 gnd.n284 0.152939
R21081 gnd.n7055 gnd.n7054 0.152939
R21082 gnd.n7056 gnd.n7055 0.152939
R21083 gnd.n7056 gnd.n278 0.152939
R21084 gnd.n7064 gnd.n278 0.152939
R21085 gnd.n7065 gnd.n7064 0.152939
R21086 gnd.n7066 gnd.n7065 0.152939
R21087 gnd.n7066 gnd.n272 0.152939
R21088 gnd.n7074 gnd.n272 0.152939
R21089 gnd.n7075 gnd.n7074 0.152939
R21090 gnd.n7076 gnd.n7075 0.152939
R21091 gnd.n7076 gnd.n266 0.152939
R21092 gnd.n7084 gnd.n266 0.152939
R21093 gnd.n7085 gnd.n7084 0.152939
R21094 gnd.n7086 gnd.n7085 0.152939
R21095 gnd.n7086 gnd.n260 0.152939
R21096 gnd.n7094 gnd.n260 0.152939
R21097 gnd.n7095 gnd.n7094 0.152939
R21098 gnd.n7096 gnd.n7095 0.152939
R21099 gnd.n7096 gnd.n254 0.152939
R21100 gnd.n7104 gnd.n254 0.152939
R21101 gnd.n5655 gnd.n5429 0.152939
R21102 gnd.n5656 gnd.n5655 0.152939
R21103 gnd.n5660 gnd.n5656 0.152939
R21104 gnd.n5661 gnd.n5660 0.152939
R21105 gnd.n5662 gnd.n5661 0.152939
R21106 gnd.n5662 gnd.n5651 0.152939
R21107 gnd.n5668 gnd.n5651 0.152939
R21108 gnd.n5669 gnd.n5668 0.152939
R21109 gnd.n5670 gnd.n5669 0.152939
R21110 gnd.n5671 gnd.n5670 0.152939
R21111 gnd.n5672 gnd.n5671 0.152939
R21112 gnd.n5675 gnd.n5672 0.152939
R21113 gnd.n5676 gnd.n5675 0.152939
R21114 gnd.n5677 gnd.n5676 0.152939
R21115 gnd.n5678 gnd.n5677 0.152939
R21116 gnd.n5680 gnd.n5678 0.152939
R21117 gnd.n5680 gnd.n5679 0.152939
R21118 gnd.n5679 gnd.n245 0.152939
R21119 gnd.n246 gnd.n245 0.152939
R21120 gnd.n247 gnd.n246 0.152939
R21121 gnd.n252 gnd.n247 0.152939
R21122 gnd.n253 gnd.n252 0.152939
R21123 gnd.n7105 gnd.n253 0.152939
R21124 gnd.n7397 gnd.n76 0.152939
R21125 gnd.n101 gnd.n76 0.152939
R21126 gnd.n102 gnd.n101 0.152939
R21127 gnd.n103 gnd.n102 0.152939
R21128 gnd.n121 gnd.n103 0.152939
R21129 gnd.n122 gnd.n121 0.152939
R21130 gnd.n123 gnd.n122 0.152939
R21131 gnd.n124 gnd.n123 0.152939
R21132 gnd.n141 gnd.n124 0.152939
R21133 gnd.n142 gnd.n141 0.152939
R21134 gnd.n143 gnd.n142 0.152939
R21135 gnd.n144 gnd.n143 0.152939
R21136 gnd.n162 gnd.n144 0.152939
R21137 gnd.n163 gnd.n162 0.152939
R21138 gnd.n164 gnd.n163 0.152939
R21139 gnd.n165 gnd.n164 0.152939
R21140 gnd.n7406 gnd.n65 0.152939
R21141 gnd.n5605 gnd.n65 0.152939
R21142 gnd.n5607 gnd.n5605 0.152939
R21143 gnd.n5607 gnd.n5606 0.152939
R21144 gnd.n5606 gnd.n5434 0.152939
R21145 gnd.n5435 gnd.n5434 0.152939
R21146 gnd.n5436 gnd.n5435 0.152939
R21147 gnd.n5618 gnd.n5436 0.152939
R21148 gnd.n5619 gnd.n5618 0.152939
R21149 gnd.n5620 gnd.n5619 0.152939
R21150 gnd.n5621 gnd.n5620 0.152939
R21151 gnd.n5625 gnd.n5621 0.152939
R21152 gnd.n5626 gnd.n5625 0.152939
R21153 gnd.n5627 gnd.n5626 0.152939
R21154 gnd.n5628 gnd.n5627 0.152939
R21155 gnd.n5631 gnd.n5628 0.152939
R21156 gnd.n5633 gnd.n5631 0.152939
R21157 gnd.n5633 gnd.n5632 0.152939
R21158 gnd.n5632 gnd.n176 0.152939
R21159 gnd.n7335 gnd.n176 0.152939
R21160 gnd.n199 gnd.n198 0.152939
R21161 gnd.n206 gnd.n198 0.152939
R21162 gnd.n207 gnd.n206 0.152939
R21163 gnd.n208 gnd.n207 0.152939
R21164 gnd.n208 gnd.n196 0.152939
R21165 gnd.n216 gnd.n196 0.152939
R21166 gnd.n217 gnd.n216 0.152939
R21167 gnd.n218 gnd.n217 0.152939
R21168 gnd.n218 gnd.n194 0.152939
R21169 gnd.n226 gnd.n194 0.152939
R21170 gnd.n227 gnd.n226 0.152939
R21171 gnd.n228 gnd.n227 0.152939
R21172 gnd.n228 gnd.n192 0.152939
R21173 gnd.n235 gnd.n192 0.152939
R21174 gnd.n236 gnd.n235 0.152939
R21175 gnd.n237 gnd.n236 0.152939
R21176 gnd.n237 gnd.n177 0.152939
R21177 gnd.n7334 gnd.n177 0.152939
R21178 gnd.n7151 gnd.n7150 0.152939
R21179 gnd.n7152 gnd.n7151 0.152939
R21180 gnd.n7153 gnd.n7152 0.152939
R21181 gnd.n7154 gnd.n7153 0.152939
R21182 gnd.n7155 gnd.n7154 0.152939
R21183 gnd.n7156 gnd.n7155 0.152939
R21184 gnd.n7157 gnd.n7156 0.152939
R21185 gnd.n7158 gnd.n7157 0.152939
R21186 gnd.n7159 gnd.n7158 0.152939
R21187 gnd.n7160 gnd.n7159 0.152939
R21188 gnd.n7161 gnd.n7160 0.152939
R21189 gnd.n7162 gnd.n7161 0.152939
R21190 gnd.n7163 gnd.n7162 0.152939
R21191 gnd.n7164 gnd.n7163 0.152939
R21192 gnd.n7165 gnd.n7164 0.152939
R21193 gnd.n7166 gnd.n7165 0.152939
R21194 gnd.n7167 gnd.n7166 0.152939
R21195 gnd.n7168 gnd.n7167 0.152939
R21196 gnd.n7169 gnd.n7168 0.152939
R21197 gnd.n7170 gnd.n7169 0.152939
R21198 gnd.n7171 gnd.n7170 0.152939
R21199 gnd.n7172 gnd.n7171 0.152939
R21200 gnd.n7173 gnd.n7172 0.152939
R21201 gnd.n7174 gnd.n7173 0.152939
R21202 gnd.n7175 gnd.n7174 0.152939
R21203 gnd.n7176 gnd.n7175 0.152939
R21204 gnd.n7177 gnd.n7176 0.152939
R21205 gnd.n7178 gnd.n7177 0.152939
R21206 gnd.n7179 gnd.n7178 0.152939
R21207 gnd.n7180 gnd.n7179 0.152939
R21208 gnd.n7181 gnd.n7180 0.152939
R21209 gnd.n7182 gnd.n7181 0.152939
R21210 gnd.n7183 gnd.n7182 0.152939
R21211 gnd.n7184 gnd.n7183 0.152939
R21212 gnd.n7185 gnd.n7184 0.152939
R21213 gnd.n7186 gnd.n7185 0.152939
R21214 gnd.n7254 gnd.n7186 0.152939
R21215 gnd.n7254 gnd.n7253 0.152939
R21216 gnd.n7253 gnd.n7252 0.152939
R21217 gnd.n7252 gnd.n7190 0.152939
R21218 gnd.n7191 gnd.n7190 0.152939
R21219 gnd.n7192 gnd.n7191 0.152939
R21220 gnd.n7193 gnd.n7192 0.152939
R21221 gnd.n7194 gnd.n7193 0.152939
R21222 gnd.n7195 gnd.n7194 0.152939
R21223 gnd.n7196 gnd.n7195 0.152939
R21224 gnd.n7197 gnd.n7196 0.152939
R21225 gnd.n7198 gnd.n7197 0.152939
R21226 gnd.n7199 gnd.n7198 0.152939
R21227 gnd.n7200 gnd.n7199 0.152939
R21228 gnd.n7201 gnd.n7200 0.152939
R21229 gnd.n7202 gnd.n7201 0.152939
R21230 gnd.n7203 gnd.n7202 0.152939
R21231 gnd.n7204 gnd.n7203 0.152939
R21232 gnd.n7205 gnd.n7204 0.152939
R21233 gnd.n7206 gnd.n7205 0.152939
R21234 gnd.n7212 gnd.n7206 0.152939
R21235 gnd.n7212 gnd.n7211 0.152939
R21236 gnd.n2750 gnd.n2749 0.152939
R21237 gnd.n2751 gnd.n2750 0.152939
R21238 gnd.n2752 gnd.n2751 0.152939
R21239 gnd.n2753 gnd.n2752 0.152939
R21240 gnd.n2754 gnd.n2753 0.152939
R21241 gnd.n2755 gnd.n2754 0.152939
R21242 gnd.n2756 gnd.n2755 0.152939
R21243 gnd.n2757 gnd.n2756 0.152939
R21244 gnd.n2758 gnd.n2757 0.152939
R21245 gnd.n2759 gnd.n2758 0.152939
R21246 gnd.n2760 gnd.n2759 0.152939
R21247 gnd.n2761 gnd.n2760 0.152939
R21248 gnd.n2762 gnd.n2761 0.152939
R21249 gnd.n2763 gnd.n2762 0.152939
R21250 gnd.n2764 gnd.n2763 0.152939
R21251 gnd.n2765 gnd.n2764 0.152939
R21252 gnd.n2766 gnd.n2765 0.152939
R21253 gnd.n2769 gnd.n2766 0.152939
R21254 gnd.n2770 gnd.n2769 0.152939
R21255 gnd.n2771 gnd.n2770 0.152939
R21256 gnd.n2772 gnd.n2771 0.152939
R21257 gnd.n2773 gnd.n2772 0.152939
R21258 gnd.n2774 gnd.n2773 0.152939
R21259 gnd.n2775 gnd.n2774 0.152939
R21260 gnd.n2776 gnd.n2775 0.152939
R21261 gnd.n2781 gnd.n2780 0.152939
R21262 gnd.n2782 gnd.n2781 0.152939
R21263 gnd.n2783 gnd.n2782 0.152939
R21264 gnd.n2784 gnd.n2783 0.152939
R21265 gnd.n2785 gnd.n2784 0.152939
R21266 gnd.n2786 gnd.n2785 0.152939
R21267 gnd.n2787 gnd.n2786 0.152939
R21268 gnd.n2788 gnd.n2787 0.152939
R21269 gnd.n2789 gnd.n2788 0.152939
R21270 gnd.n2792 gnd.n2789 0.152939
R21271 gnd.n2793 gnd.n2792 0.152939
R21272 gnd.n2794 gnd.n2793 0.152939
R21273 gnd.n2795 gnd.n2794 0.152939
R21274 gnd.n2796 gnd.n2795 0.152939
R21275 gnd.n2797 gnd.n2796 0.152939
R21276 gnd.n2798 gnd.n2797 0.152939
R21277 gnd.n2799 gnd.n2798 0.152939
R21278 gnd.n2800 gnd.n2799 0.152939
R21279 gnd.n2801 gnd.n2800 0.152939
R21280 gnd.n2802 gnd.n2801 0.152939
R21281 gnd.n2803 gnd.n2802 0.152939
R21282 gnd.n2804 gnd.n2803 0.152939
R21283 gnd.n2805 gnd.n2804 0.152939
R21284 gnd.n2806 gnd.n2805 0.152939
R21285 gnd.n2807 gnd.n2806 0.152939
R21286 gnd.n2808 gnd.n2807 0.152939
R21287 gnd.n2809 gnd.n2808 0.152939
R21288 gnd.n2810 gnd.n2809 0.152939
R21289 gnd.n5813 gnd.n2810 0.152939
R21290 gnd.n5813 gnd.n5812 0.152939
R21291 gnd.n5325 gnd.n5324 0.152939
R21292 gnd.n5326 gnd.n5325 0.152939
R21293 gnd.n5327 gnd.n5326 0.152939
R21294 gnd.n5346 gnd.n5327 0.152939
R21295 gnd.n5347 gnd.n5346 0.152939
R21296 gnd.n5348 gnd.n5347 0.152939
R21297 gnd.n5349 gnd.n5348 0.152939
R21298 gnd.n5365 gnd.n5349 0.152939
R21299 gnd.n5366 gnd.n5365 0.152939
R21300 gnd.n5367 gnd.n5366 0.152939
R21301 gnd.n5368 gnd.n5367 0.152939
R21302 gnd.n5386 gnd.n5368 0.152939
R21303 gnd.n5387 gnd.n5386 0.152939
R21304 gnd.n5388 gnd.n5387 0.152939
R21305 gnd.n5388 gnd.n77 0.152939
R21306 gnd.n7397 gnd.n77 0.152939
R21307 gnd.n3771 gnd.n3764 0.152939
R21308 gnd.n3772 gnd.n3771 0.152939
R21309 gnd.n3772 gnd.n3686 0.152939
R21310 gnd.n4249 gnd.n3686 0.152939
R21311 gnd.n4250 gnd.n4249 0.152939
R21312 gnd.n4251 gnd.n4250 0.152939
R21313 gnd.n4251 gnd.n3682 0.152939
R21314 gnd.n4257 gnd.n3682 0.152939
R21315 gnd.n4258 gnd.n4257 0.152939
R21316 gnd.n4259 gnd.n4258 0.152939
R21317 gnd.n4259 gnd.n3678 0.152939
R21318 gnd.n4265 gnd.n3678 0.152939
R21319 gnd.n4266 gnd.n4265 0.152939
R21320 gnd.n4267 gnd.n4266 0.152939
R21321 gnd.n4267 gnd.n3674 0.152939
R21322 gnd.n4273 gnd.n3674 0.152939
R21323 gnd.n4274 gnd.n4273 0.152939
R21324 gnd.n4276 gnd.n4274 0.152939
R21325 gnd.n4276 gnd.n4275 0.152939
R21326 gnd.n4275 gnd.n2568 0.152939
R21327 gnd.n2569 gnd.n2568 0.152939
R21328 gnd.n2570 gnd.n2569 0.152939
R21329 gnd.n3453 gnd.n2570 0.152939
R21330 gnd.n3454 gnd.n3453 0.152939
R21331 gnd.n3455 gnd.n3454 0.152939
R21332 gnd.n3455 gnd.n3446 0.152939
R21333 gnd.n3465 gnd.n3446 0.152939
R21334 gnd.n3466 gnd.n3465 0.152939
R21335 gnd.n3467 gnd.n3466 0.152939
R21336 gnd.n3467 gnd.n3440 0.152939
R21337 gnd.n3477 gnd.n3440 0.152939
R21338 gnd.n3478 gnd.n3477 0.152939
R21339 gnd.n3479 gnd.n3478 0.152939
R21340 gnd.n3480 gnd.n3479 0.152939
R21341 gnd.n3480 gnd.n3219 0.152939
R21342 gnd.n4559 gnd.n3219 0.152939
R21343 gnd.n4560 gnd.n4559 0.152939
R21344 gnd.n4561 gnd.n4560 0.152939
R21345 gnd.n4562 gnd.n4561 0.152939
R21346 gnd.n4562 gnd.n3195 0.152939
R21347 gnd.n4597 gnd.n3195 0.152939
R21348 gnd.n4598 gnd.n4597 0.152939
R21349 gnd.n4599 gnd.n4598 0.152939
R21350 gnd.n4600 gnd.n4599 0.152939
R21351 gnd.n4601 gnd.n4600 0.152939
R21352 gnd.n4601 gnd.n3170 0.152939
R21353 gnd.n4637 gnd.n3170 0.152939
R21354 gnd.n4638 gnd.n4637 0.152939
R21355 gnd.n4639 gnd.n4638 0.152939
R21356 gnd.n4640 gnd.n4639 0.152939
R21357 gnd.n4640 gnd.n3142 0.152939
R21358 gnd.n4673 gnd.n3142 0.152939
R21359 gnd.n4674 gnd.n4673 0.152939
R21360 gnd.n4675 gnd.n4674 0.152939
R21361 gnd.n4675 gnd.n3124 0.152939
R21362 gnd.n4699 gnd.n3124 0.152939
R21363 gnd.n4700 gnd.n4699 0.152939
R21364 gnd.n4701 gnd.n4700 0.152939
R21365 gnd.n4702 gnd.n4701 0.152939
R21366 gnd.n4702 gnd.n3098 0.152939
R21367 gnd.n4755 gnd.n3098 0.152939
R21368 gnd.n4756 gnd.n4755 0.152939
R21369 gnd.n4757 gnd.n4756 0.152939
R21370 gnd.n4758 gnd.n4757 0.152939
R21371 gnd.n4758 gnd.n3073 0.152939
R21372 gnd.n4795 gnd.n3073 0.152939
R21373 gnd.n4796 gnd.n4795 0.152939
R21374 gnd.n4797 gnd.n4796 0.152939
R21375 gnd.n4798 gnd.n4797 0.152939
R21376 gnd.n4798 gnd.n3043 0.152939
R21377 gnd.n4864 gnd.n3043 0.152939
R21378 gnd.n4865 gnd.n4864 0.152939
R21379 gnd.n4866 gnd.n4865 0.152939
R21380 gnd.n4867 gnd.n4866 0.152939
R21381 gnd.n4867 gnd.n3019 0.152939
R21382 gnd.n4897 gnd.n3019 0.152939
R21383 gnd.n4898 gnd.n4897 0.152939
R21384 gnd.n4899 gnd.n4898 0.152939
R21385 gnd.n4900 gnd.n4899 0.152939
R21386 gnd.n4900 gnd.n2998 0.152939
R21387 gnd.n4951 gnd.n2998 0.152939
R21388 gnd.n4952 gnd.n4951 0.152939
R21389 gnd.n4953 gnd.n4952 0.152939
R21390 gnd.n4954 gnd.n4953 0.152939
R21391 gnd.n4954 gnd.n2973 0.152939
R21392 gnd.n4988 gnd.n2973 0.152939
R21393 gnd.n4989 gnd.n4988 0.152939
R21394 gnd.n4990 gnd.n4989 0.152939
R21395 gnd.n4990 gnd.n2882 0.152939
R21396 gnd.n5131 gnd.n2882 0.152939
R21397 gnd.n5132 gnd.n5131 0.152939
R21398 gnd.n5133 gnd.n5132 0.152939
R21399 gnd.n5133 gnd.n2869 0.152939
R21400 gnd.n5147 gnd.n2869 0.152939
R21401 gnd.n5148 gnd.n5147 0.152939
R21402 gnd.n5149 gnd.n5148 0.152939
R21403 gnd.n5149 gnd.n2856 0.152939
R21404 gnd.n5163 gnd.n2856 0.152939
R21405 gnd.n5164 gnd.n5163 0.152939
R21406 gnd.n5165 gnd.n5164 0.152939
R21407 gnd.n5165 gnd.n2842 0.152939
R21408 gnd.n5180 gnd.n2842 0.152939
R21409 gnd.n5181 gnd.n5180 0.152939
R21410 gnd.n5183 gnd.n5181 0.152939
R21411 gnd.n5183 gnd.n5182 0.152939
R21412 gnd.n5182 gnd.n2702 0.152939
R21413 gnd.n2703 gnd.n2702 0.152939
R21414 gnd.n2704 gnd.n2703 0.152939
R21415 gnd.n5460 gnd.n2704 0.152939
R21416 gnd.n5461 gnd.n5460 0.152939
R21417 gnd.n5466 gnd.n5461 0.152939
R21418 gnd.n5467 gnd.n5466 0.152939
R21419 gnd.n5468 gnd.n5467 0.152939
R21420 gnd.n5468 gnd.n5456 0.152939
R21421 gnd.n5474 gnd.n5456 0.152939
R21422 gnd.n5475 gnd.n5474 0.152939
R21423 gnd.n5476 gnd.n5475 0.152939
R21424 gnd.n5476 gnd.n5452 0.152939
R21425 gnd.n5545 gnd.n5452 0.152939
R21426 gnd.n5546 gnd.n5545 0.152939
R21427 gnd.n5547 gnd.n5546 0.152939
R21428 gnd.n5547 gnd.n5448 0.152939
R21429 gnd.n5553 gnd.n5448 0.152939
R21430 gnd.n5554 gnd.n5553 0.152939
R21431 gnd.n5555 gnd.n5554 0.152939
R21432 gnd.n5556 gnd.n5555 0.152939
R21433 gnd.n3852 gnd.n3847 0.152939
R21434 gnd.n3847 gnd.n3816 0.152939
R21435 gnd.n4117 gnd.n3816 0.152939
R21436 gnd.n4118 gnd.n4117 0.152939
R21437 gnd.n4119 gnd.n4118 0.152939
R21438 gnd.n4119 gnd.n3729 0.152939
R21439 gnd.n4131 gnd.n3729 0.152939
R21440 gnd.n4132 gnd.n4131 0.152939
R21441 gnd.n4133 gnd.n4132 0.152939
R21442 gnd.n4133 gnd.n3724 0.152939
R21443 gnd.n4145 gnd.n3724 0.152939
R21444 gnd.n4146 gnd.n4145 0.152939
R21445 gnd.n4147 gnd.n4146 0.152939
R21446 gnd.n4147 gnd.n3718 0.152939
R21447 gnd.n4159 gnd.n3718 0.152939
R21448 gnd.n4160 gnd.n4159 0.152939
R21449 gnd.n4161 gnd.n4160 0.152939
R21450 gnd.n4161 gnd.n3713 0.152939
R21451 gnd.n4173 gnd.n3713 0.152939
R21452 gnd.n4174 gnd.n4173 0.152939
R21453 gnd.n3893 gnd.n3820 0.152939
R21454 gnd.n3823 gnd.n3820 0.152939
R21455 gnd.n3824 gnd.n3823 0.152939
R21456 gnd.n3827 gnd.n3824 0.152939
R21457 gnd.n3828 gnd.n3827 0.152939
R21458 gnd.n3829 gnd.n3828 0.152939
R21459 gnd.n3830 gnd.n3829 0.152939
R21460 gnd.n3833 gnd.n3830 0.152939
R21461 gnd.n3834 gnd.n3833 0.152939
R21462 gnd.n3835 gnd.n3834 0.152939
R21463 gnd.n3836 gnd.n3835 0.152939
R21464 gnd.n3839 gnd.n3836 0.152939
R21465 gnd.n3840 gnd.n3839 0.152939
R21466 gnd.n3841 gnd.n3840 0.152939
R21467 gnd.n3842 gnd.n3841 0.152939
R21468 gnd.n3846 gnd.n3842 0.152939
R21469 gnd.n3854 gnd.n3846 0.152939
R21470 gnd.n3854 gnd.n3853 0.152939
R21471 gnd.n2466 gnd.n2413 0.152939
R21472 gnd.n2467 gnd.n2466 0.152939
R21473 gnd.n2468 gnd.n2467 0.152939
R21474 gnd.n2469 gnd.n2468 0.152939
R21475 gnd.n2486 gnd.n2469 0.152939
R21476 gnd.n2487 gnd.n2486 0.152939
R21477 gnd.n2488 gnd.n2487 0.152939
R21478 gnd.n2489 gnd.n2488 0.152939
R21479 gnd.n2507 gnd.n2489 0.152939
R21480 gnd.n2508 gnd.n2507 0.152939
R21481 gnd.n2509 gnd.n2508 0.152939
R21482 gnd.n2510 gnd.n2509 0.152939
R21483 gnd.n2527 gnd.n2510 0.152939
R21484 gnd.n2528 gnd.n2527 0.152939
R21485 gnd.n2529 gnd.n2528 0.152939
R21486 gnd.n2530 gnd.n2529 0.152939
R21487 gnd.n4298 gnd.n4297 0.152939
R21488 gnd.n4299 gnd.n4298 0.152939
R21489 gnd.n4300 gnd.n4299 0.152939
R21490 gnd.n4301 gnd.n4300 0.152939
R21491 gnd.n4302 gnd.n4301 0.152939
R21492 gnd.n4303 gnd.n4302 0.152939
R21493 gnd.n4304 gnd.n4303 0.152939
R21494 gnd.n4305 gnd.n4304 0.152939
R21495 gnd.n4306 gnd.n4305 0.152939
R21496 gnd.n4307 gnd.n4306 0.152939
R21497 gnd.n4308 gnd.n4307 0.152939
R21498 gnd.n4309 gnd.n4308 0.152939
R21499 gnd.n4310 gnd.n4309 0.152939
R21500 gnd.n4311 gnd.n4310 0.152939
R21501 gnd.n4312 gnd.n4311 0.152939
R21502 gnd.n4313 gnd.n4312 0.152939
R21503 gnd.n4314 gnd.n4313 0.152939
R21504 gnd.n4317 gnd.n4314 0.152939
R21505 gnd.n4318 gnd.n4317 0.152939
R21506 gnd.n4319 gnd.n4318 0.152939
R21507 gnd.n4320 gnd.n4319 0.152939
R21508 gnd.n4321 gnd.n4320 0.152939
R21509 gnd.n4322 gnd.n4321 0.152939
R21510 gnd.n4323 gnd.n4322 0.152939
R21511 gnd.n4323 gnd.n3362 0.152939
R21512 gnd.n4480 gnd.n4479 0.152939
R21513 gnd.n4479 gnd.n3363 0.152939
R21514 gnd.n4375 gnd.n3363 0.152939
R21515 gnd.n4376 gnd.n4375 0.152939
R21516 gnd.n4377 gnd.n4376 0.152939
R21517 gnd.n4378 gnd.n4377 0.152939
R21518 gnd.n4382 gnd.n4378 0.152939
R21519 gnd.n4383 gnd.n4382 0.152939
R21520 gnd.n4462 gnd.n4383 0.152939
R21521 gnd.n4462 gnd.n4461 0.152939
R21522 gnd.n4461 gnd.n4460 0.152939
R21523 gnd.n4460 gnd.n4387 0.152939
R21524 gnd.n4393 gnd.n4387 0.152939
R21525 gnd.n4394 gnd.n4393 0.152939
R21526 gnd.n4395 gnd.n4394 0.152939
R21527 gnd.n4396 gnd.n4395 0.152939
R21528 gnd.n4400 gnd.n4396 0.152939
R21529 gnd.n4401 gnd.n4400 0.152939
R21530 gnd.n4402 gnd.n4401 0.152939
R21531 gnd.n4403 gnd.n4402 0.152939
R21532 gnd.n4407 gnd.n4403 0.152939
R21533 gnd.n4408 gnd.n4407 0.152939
R21534 gnd.n4409 gnd.n4408 0.152939
R21535 gnd.n4410 gnd.n4409 0.152939
R21536 gnd.n4414 gnd.n4410 0.152939
R21537 gnd.n4415 gnd.n4414 0.152939
R21538 gnd.n4416 gnd.n4415 0.152939
R21539 gnd.n4417 gnd.n4416 0.152939
R21540 gnd.n4422 gnd.n4417 0.152939
R21541 gnd.n4423 gnd.n4422 0.152939
R21542 gnd.n3961 gnd.n3956 0.152939
R21543 gnd.n3962 gnd.n3961 0.152939
R21544 gnd.n3963 gnd.n3962 0.152939
R21545 gnd.n3963 gnd.n3952 0.152939
R21546 gnd.n3971 gnd.n3952 0.152939
R21547 gnd.n3972 gnd.n3971 0.152939
R21548 gnd.n3973 gnd.n3972 0.152939
R21549 gnd.n3973 gnd.n3948 0.152939
R21550 gnd.n3981 gnd.n3948 0.152939
R21551 gnd.n3982 gnd.n3981 0.152939
R21552 gnd.n3983 gnd.n3982 0.152939
R21553 gnd.n3983 gnd.n3944 0.152939
R21554 gnd.n3991 gnd.n3944 0.152939
R21555 gnd.n3992 gnd.n3991 0.152939
R21556 gnd.n3993 gnd.n3992 0.152939
R21557 gnd.n3993 gnd.n3937 0.152939
R21558 gnd.n4001 gnd.n3937 0.152939
R21559 gnd.n4002 gnd.n4001 0.152939
R21560 gnd.n4003 gnd.n4002 0.152939
R21561 gnd.n4003 gnd.n3933 0.152939
R21562 gnd.n4011 gnd.n3933 0.152939
R21563 gnd.n4012 gnd.n4011 0.152939
R21564 gnd.n4013 gnd.n4012 0.152939
R21565 gnd.n4013 gnd.n3929 0.152939
R21566 gnd.n4021 gnd.n3929 0.152939
R21567 gnd.n4022 gnd.n4021 0.152939
R21568 gnd.n4023 gnd.n4022 0.152939
R21569 gnd.n4023 gnd.n3925 0.152939
R21570 gnd.n4031 gnd.n3925 0.152939
R21571 gnd.n4032 gnd.n4031 0.152939
R21572 gnd.n4033 gnd.n4032 0.152939
R21573 gnd.n4033 gnd.n3921 0.152939
R21574 gnd.n4041 gnd.n3921 0.152939
R21575 gnd.n4042 gnd.n4041 0.152939
R21576 gnd.n4043 gnd.n4042 0.152939
R21577 gnd.n4043 gnd.n3917 0.152939
R21578 gnd.n4053 gnd.n3917 0.152939
R21579 gnd.n4054 gnd.n4053 0.152939
R21580 gnd.n4055 gnd.n4054 0.152939
R21581 gnd.n4055 gnd.n3913 0.152939
R21582 gnd.n4063 gnd.n3913 0.152939
R21583 gnd.n4064 gnd.n4063 0.152939
R21584 gnd.n4065 gnd.n4064 0.152939
R21585 gnd.n4065 gnd.n3909 0.152939
R21586 gnd.n4073 gnd.n3909 0.152939
R21587 gnd.n4074 gnd.n4073 0.152939
R21588 gnd.n4075 gnd.n4074 0.152939
R21589 gnd.n4075 gnd.n3905 0.152939
R21590 gnd.n4083 gnd.n3905 0.152939
R21591 gnd.n4084 gnd.n4083 0.152939
R21592 gnd.n4085 gnd.n4084 0.152939
R21593 gnd.n4085 gnd.n3901 0.152939
R21594 gnd.n4093 gnd.n3901 0.152939
R21595 gnd.n4094 gnd.n4093 0.152939
R21596 gnd.n4096 gnd.n4094 0.152939
R21597 gnd.n4096 gnd.n4095 0.152939
R21598 gnd.n4095 gnd.n3894 0.152939
R21599 gnd.n4105 gnd.n3894 0.152939
R21600 gnd.n2330 gnd.n2329 0.152939
R21601 gnd.n2331 gnd.n2330 0.152939
R21602 gnd.n2351 gnd.n2331 0.152939
R21603 gnd.n2352 gnd.n2351 0.152939
R21604 gnd.n2353 gnd.n2352 0.152939
R21605 gnd.n2354 gnd.n2353 0.152939
R21606 gnd.n2371 gnd.n2354 0.152939
R21607 gnd.n2372 gnd.n2371 0.152939
R21608 gnd.n2373 gnd.n2372 0.152939
R21609 gnd.n2374 gnd.n2373 0.152939
R21610 gnd.n2392 gnd.n2374 0.152939
R21611 gnd.n2393 gnd.n2392 0.152939
R21612 gnd.n2394 gnd.n2393 0.152939
R21613 gnd.n2395 gnd.n2394 0.152939
R21614 gnd.n2412 gnd.n2395 0.152939
R21615 gnd.n2413 gnd.n2412 0.152939
R21616 gnd.n2309 gnd.n2308 0.152939
R21617 gnd.n2310 gnd.n2309 0.152939
R21618 gnd.n2311 gnd.n2310 0.152939
R21619 gnd.n2316 gnd.n2311 0.152939
R21620 gnd.n2317 gnd.n2316 0.152939
R21621 gnd.n2318 gnd.n2317 0.152939
R21622 gnd.n2319 gnd.n2318 0.152939
R21623 gnd.n3738 gnd.n2319 0.152939
R21624 gnd.n3739 gnd.n3738 0.152939
R21625 gnd.n3740 gnd.n3739 0.152939
R21626 gnd.n3740 gnd.n3734 0.152939
R21627 gnd.n3746 gnd.n3734 0.152939
R21628 gnd.n3747 gnd.n3746 0.152939
R21629 gnd.n3748 gnd.n3747 0.152939
R21630 gnd.n3749 gnd.n3748 0.152939
R21631 gnd.n3750 gnd.n3749 0.152939
R21632 gnd.n3753 gnd.n3750 0.152939
R21633 gnd.n3754 gnd.n3753 0.152939
R21634 gnd.n3755 gnd.n3754 0.152939
R21635 gnd.n3756 gnd.n3755 0.152939
R21636 gnd.n3759 gnd.n3756 0.152939
R21637 gnd.n3760 gnd.n3759 0.152939
R21638 gnd.n3761 gnd.n3760 0.152939
R21639 gnd.n6403 gnd.n673 0.152939
R21640 gnd.n678 gnd.n673 0.152939
R21641 gnd.n679 gnd.n678 0.152939
R21642 gnd.n680 gnd.n679 0.152939
R21643 gnd.n685 gnd.n680 0.152939
R21644 gnd.n686 gnd.n685 0.152939
R21645 gnd.n687 gnd.n686 0.152939
R21646 gnd.n688 gnd.n687 0.152939
R21647 gnd.n693 gnd.n688 0.152939
R21648 gnd.n694 gnd.n693 0.152939
R21649 gnd.n695 gnd.n694 0.152939
R21650 gnd.n696 gnd.n695 0.152939
R21651 gnd.n701 gnd.n696 0.152939
R21652 gnd.n702 gnd.n701 0.152939
R21653 gnd.n703 gnd.n702 0.152939
R21654 gnd.n704 gnd.n703 0.152939
R21655 gnd.n709 gnd.n704 0.152939
R21656 gnd.n710 gnd.n709 0.152939
R21657 gnd.n711 gnd.n710 0.152939
R21658 gnd.n712 gnd.n711 0.152939
R21659 gnd.n717 gnd.n712 0.152939
R21660 gnd.n718 gnd.n717 0.152939
R21661 gnd.n719 gnd.n718 0.152939
R21662 gnd.n720 gnd.n719 0.152939
R21663 gnd.n725 gnd.n720 0.152939
R21664 gnd.n726 gnd.n725 0.152939
R21665 gnd.n727 gnd.n726 0.152939
R21666 gnd.n728 gnd.n727 0.152939
R21667 gnd.n733 gnd.n728 0.152939
R21668 gnd.n734 gnd.n733 0.152939
R21669 gnd.n735 gnd.n734 0.152939
R21670 gnd.n736 gnd.n735 0.152939
R21671 gnd.n741 gnd.n736 0.152939
R21672 gnd.n742 gnd.n741 0.152939
R21673 gnd.n743 gnd.n742 0.152939
R21674 gnd.n744 gnd.n743 0.152939
R21675 gnd.n749 gnd.n744 0.152939
R21676 gnd.n750 gnd.n749 0.152939
R21677 gnd.n751 gnd.n750 0.152939
R21678 gnd.n752 gnd.n751 0.152939
R21679 gnd.n757 gnd.n752 0.152939
R21680 gnd.n758 gnd.n757 0.152939
R21681 gnd.n759 gnd.n758 0.152939
R21682 gnd.n760 gnd.n759 0.152939
R21683 gnd.n765 gnd.n760 0.152939
R21684 gnd.n766 gnd.n765 0.152939
R21685 gnd.n767 gnd.n766 0.152939
R21686 gnd.n768 gnd.n767 0.152939
R21687 gnd.n773 gnd.n768 0.152939
R21688 gnd.n774 gnd.n773 0.152939
R21689 gnd.n775 gnd.n774 0.152939
R21690 gnd.n776 gnd.n775 0.152939
R21691 gnd.n781 gnd.n776 0.152939
R21692 gnd.n782 gnd.n781 0.152939
R21693 gnd.n783 gnd.n782 0.152939
R21694 gnd.n784 gnd.n783 0.152939
R21695 gnd.n789 gnd.n784 0.152939
R21696 gnd.n790 gnd.n789 0.152939
R21697 gnd.n791 gnd.n790 0.152939
R21698 gnd.n792 gnd.n791 0.152939
R21699 gnd.n797 gnd.n792 0.152939
R21700 gnd.n798 gnd.n797 0.152939
R21701 gnd.n799 gnd.n798 0.152939
R21702 gnd.n800 gnd.n799 0.152939
R21703 gnd.n805 gnd.n800 0.152939
R21704 gnd.n806 gnd.n805 0.152939
R21705 gnd.n807 gnd.n806 0.152939
R21706 gnd.n808 gnd.n807 0.152939
R21707 gnd.n813 gnd.n808 0.152939
R21708 gnd.n814 gnd.n813 0.152939
R21709 gnd.n815 gnd.n814 0.152939
R21710 gnd.n816 gnd.n815 0.152939
R21711 gnd.n821 gnd.n816 0.152939
R21712 gnd.n822 gnd.n821 0.152939
R21713 gnd.n823 gnd.n822 0.152939
R21714 gnd.n824 gnd.n823 0.152939
R21715 gnd.n829 gnd.n824 0.152939
R21716 gnd.n830 gnd.n829 0.152939
R21717 gnd.n831 gnd.n830 0.152939
R21718 gnd.n832 gnd.n831 0.152939
R21719 gnd.n837 gnd.n832 0.152939
R21720 gnd.n838 gnd.n837 0.152939
R21721 gnd.n839 gnd.n838 0.152939
R21722 gnd.n840 gnd.n839 0.152939
R21723 gnd.n6059 gnd.n2578 0.152939
R21724 gnd.n6059 gnd.n6058 0.152939
R21725 gnd.n6058 gnd.n6057 0.152939
R21726 gnd.n6057 gnd.n2579 0.152939
R21727 gnd.n6053 gnd.n2579 0.152939
R21728 gnd.n6053 gnd.n6052 0.152939
R21729 gnd.n6052 gnd.n6051 0.152939
R21730 gnd.n6051 gnd.n2584 0.152939
R21731 gnd.n6047 gnd.n2584 0.152939
R21732 gnd.n6047 gnd.n6046 0.152939
R21733 gnd.n6046 gnd.n6045 0.152939
R21734 gnd.n6045 gnd.n2589 0.152939
R21735 gnd.n6041 gnd.n2589 0.152939
R21736 gnd.n6041 gnd.n6040 0.152939
R21737 gnd.n6040 gnd.n6039 0.152939
R21738 gnd.n6039 gnd.n2594 0.152939
R21739 gnd.n6035 gnd.n2594 0.152939
R21740 gnd.n6035 gnd.n6034 0.152939
R21741 gnd.n6034 gnd.n6033 0.152939
R21742 gnd.n6033 gnd.n2599 0.152939
R21743 gnd.n6029 gnd.n2599 0.152939
R21744 gnd.n6029 gnd.n6028 0.152939
R21745 gnd.n6028 gnd.n6027 0.152939
R21746 gnd.n6027 gnd.n2604 0.152939
R21747 gnd.n6023 gnd.n2604 0.152939
R21748 gnd.n6023 gnd.n6022 0.152939
R21749 gnd.n6022 gnd.n6021 0.152939
R21750 gnd.n6021 gnd.n2609 0.152939
R21751 gnd.n6017 gnd.n2609 0.152939
R21752 gnd.n6017 gnd.n6016 0.152939
R21753 gnd.n6016 gnd.n6015 0.152939
R21754 gnd.n6015 gnd.n2614 0.152939
R21755 gnd.n6011 gnd.n2614 0.152939
R21756 gnd.n6011 gnd.n6010 0.152939
R21757 gnd.n6010 gnd.n6009 0.152939
R21758 gnd.n6009 gnd.n2619 0.152939
R21759 gnd.n6005 gnd.n2619 0.152939
R21760 gnd.n6005 gnd.n6004 0.152939
R21761 gnd.n6004 gnd.n6003 0.152939
R21762 gnd.n6003 gnd.n2624 0.152939
R21763 gnd.n5999 gnd.n2624 0.152939
R21764 gnd.n5999 gnd.n5998 0.152939
R21765 gnd.n5998 gnd.n5997 0.152939
R21766 gnd.n5997 gnd.n2629 0.152939
R21767 gnd.n5993 gnd.n2629 0.152939
R21768 gnd.n5993 gnd.n5992 0.152939
R21769 gnd.n5992 gnd.n5991 0.152939
R21770 gnd.n5991 gnd.n2634 0.152939
R21771 gnd.n5987 gnd.n2634 0.152939
R21772 gnd.n5987 gnd.n5986 0.152939
R21773 gnd.n5986 gnd.n5985 0.152939
R21774 gnd.n5985 gnd.n2639 0.152939
R21775 gnd.n5981 gnd.n2639 0.152939
R21776 gnd.n5981 gnd.n5980 0.152939
R21777 gnd.n5980 gnd.n5979 0.152939
R21778 gnd.n5979 gnd.n2644 0.152939
R21779 gnd.n5975 gnd.n2644 0.152939
R21780 gnd.n5975 gnd.n5974 0.152939
R21781 gnd.n5974 gnd.n5973 0.152939
R21782 gnd.n5973 gnd.n2649 0.152939
R21783 gnd.n5969 gnd.n2649 0.152939
R21784 gnd.n5969 gnd.n5968 0.152939
R21785 gnd.n5968 gnd.n5967 0.152939
R21786 gnd.n5967 gnd.n2654 0.152939
R21787 gnd.n5963 gnd.n2654 0.152939
R21788 gnd.n5963 gnd.n5962 0.152939
R21789 gnd.n5962 gnd.n5961 0.152939
R21790 gnd.n5961 gnd.n2659 0.152939
R21791 gnd.n5957 gnd.n2659 0.152939
R21792 gnd.n5957 gnd.n5956 0.152939
R21793 gnd.n5956 gnd.n5955 0.152939
R21794 gnd.n5955 gnd.n2664 0.152939
R21795 gnd.n5951 gnd.n2664 0.152939
R21796 gnd.n5951 gnd.n5950 0.152939
R21797 gnd.n5950 gnd.n5949 0.152939
R21798 gnd.n5949 gnd.n2669 0.152939
R21799 gnd.n5945 gnd.n2669 0.152939
R21800 gnd.n5945 gnd.n5944 0.152939
R21801 gnd.n5944 gnd.n5943 0.152939
R21802 gnd.n5943 gnd.n2674 0.152939
R21803 gnd.n5939 gnd.n2674 0.152939
R21804 gnd.n5939 gnd.n5938 0.152939
R21805 gnd.n4187 gnd.n3707 0.152939
R21806 gnd.n4188 gnd.n4187 0.152939
R21807 gnd.n4189 gnd.n4188 0.152939
R21808 gnd.n4189 gnd.n3702 0.152939
R21809 gnd.n4201 gnd.n3702 0.152939
R21810 gnd.n4202 gnd.n4201 0.152939
R21811 gnd.n4203 gnd.n4202 0.152939
R21812 gnd.n4203 gnd.n3692 0.152939
R21813 gnd.n4242 gnd.n3692 0.152939
R21814 gnd.n4242 gnd.n4241 0.152939
R21815 gnd.n4241 gnd.n4240 0.152939
R21816 gnd.n4240 gnd.n3693 0.152939
R21817 gnd.n4236 gnd.n3693 0.152939
R21818 gnd.n4236 gnd.n4235 0.152939
R21819 gnd.n4235 gnd.n4234 0.152939
R21820 gnd.n4234 gnd.n3697 0.152939
R21821 gnd.n4230 gnd.n3697 0.152939
R21822 gnd.n4230 gnd.n2543 0.152939
R21823 gnd.n6076 gnd.n2543 0.152939
R21824 gnd.n6076 gnd.n6075 0.152939
R21825 gnd.n3581 gnd.n3580 0.152939
R21826 gnd.n3582 gnd.n3581 0.152939
R21827 gnd.n3582 gnd.n3419 0.152939
R21828 gnd.n3588 gnd.n3419 0.152939
R21829 gnd.n3589 gnd.n3588 0.152939
R21830 gnd.n3590 gnd.n3589 0.152939
R21831 gnd.n3577 gnd.n3423 0.152939
R21832 gnd.n3573 gnd.n3423 0.152939
R21833 gnd.n3573 gnd.n3572 0.152939
R21834 gnd.n3572 gnd.n3571 0.152939
R21835 gnd.n3571 gnd.n3426 0.152939
R21836 gnd.n3567 gnd.n3426 0.152939
R21837 gnd.n3567 gnd.n3566 0.152939
R21838 gnd.n3566 gnd.n3565 0.152939
R21839 gnd.n3565 gnd.n3431 0.152939
R21840 gnd.n3561 gnd.n3431 0.152939
R21841 gnd.n3561 gnd.n3560 0.152939
R21842 gnd.n3560 gnd.n3559 0.152939
R21843 gnd.n3559 gnd.n3436 0.152939
R21844 gnd.n3555 gnd.n3436 0.152939
R21845 gnd.n3555 gnd.n3554 0.152939
R21846 gnd.n3554 gnd.n3553 0.152939
R21847 gnd.n3553 gnd.n3490 0.152939
R21848 gnd.n3549 gnd.n3490 0.152939
R21849 gnd.n3549 gnd.n3548 0.152939
R21850 gnd.n3548 gnd.n3547 0.152939
R21851 gnd.n3547 gnd.n3497 0.152939
R21852 gnd.n3543 gnd.n3497 0.152939
R21853 gnd.n3543 gnd.n3542 0.152939
R21854 gnd.n3542 gnd.n3541 0.152939
R21855 gnd.n3541 gnd.n3503 0.152939
R21856 gnd.n3537 gnd.n3503 0.152939
R21857 gnd.n3537 gnd.n3536 0.152939
R21858 gnd.n3536 gnd.n3535 0.152939
R21859 gnd.n3535 gnd.n3506 0.152939
R21860 gnd.n3531 gnd.n3506 0.152939
R21861 gnd.n3531 gnd.n3530 0.152939
R21862 gnd.n3530 gnd.n3529 0.152939
R21863 gnd.n3529 gnd.n3511 0.152939
R21864 gnd.n3525 gnd.n3511 0.152939
R21865 gnd.n3525 gnd.n3524 0.152939
R21866 gnd.n3524 gnd.n3523 0.152939
R21867 gnd.n3523 gnd.n3515 0.152939
R21868 gnd.n3519 gnd.n3515 0.152939
R21869 gnd.n3519 gnd.n3518 0.152939
R21870 gnd.n3518 gnd.n3088 0.152939
R21871 gnd.n4765 gnd.n3088 0.152939
R21872 gnd.n4766 gnd.n4765 0.152939
R21873 gnd.n4781 gnd.n4766 0.152939
R21874 gnd.n4781 gnd.n4780 0.152939
R21875 gnd.n4780 gnd.n4779 0.152939
R21876 gnd.n4779 gnd.n4767 0.152939
R21877 gnd.n4775 gnd.n4767 0.152939
R21878 gnd.n4775 gnd.n4774 0.152939
R21879 gnd.n4774 gnd.n4773 0.152939
R21880 gnd.n4773 gnd.n3035 0.152939
R21881 gnd.n4874 gnd.n3035 0.152939
R21882 gnd.n4875 gnd.n4874 0.152939
R21883 gnd.n4877 gnd.n4875 0.152939
R21884 gnd.n4877 gnd.n4876 0.152939
R21885 gnd.n4876 gnd.n3012 0.152939
R21886 gnd.n4907 gnd.n3012 0.152939
R21887 gnd.n4908 gnd.n4907 0.152939
R21888 gnd.n4936 gnd.n4908 0.152939
R21889 gnd.n4936 gnd.n4935 0.152939
R21890 gnd.n4935 gnd.n4934 0.152939
R21891 gnd.n4934 gnd.n4909 0.152939
R21892 gnd.n4930 gnd.n4909 0.152939
R21893 gnd.n4930 gnd.n4929 0.152939
R21894 gnd.n4929 gnd.n4928 0.152939
R21895 gnd.n4928 gnd.n4917 0.152939
R21896 gnd.n4924 gnd.n4917 0.152939
R21897 gnd.n4924 gnd.n4923 0.152939
R21898 gnd.n4923 gnd.n4922 0.152939
R21899 gnd.n4922 gnd.n2874 0.152939
R21900 gnd.n5139 gnd.n2874 0.152939
R21901 gnd.n5140 gnd.n5139 0.152939
R21902 gnd.n5141 gnd.n5140 0.152939
R21903 gnd.n5141 gnd.n2861 0.152939
R21904 gnd.n5155 gnd.n2861 0.152939
R21905 gnd.n5156 gnd.n5155 0.152939
R21906 gnd.n5157 gnd.n5156 0.152939
R21907 gnd.n5157 gnd.n2849 0.152939
R21908 gnd.n5171 gnd.n2849 0.152939
R21909 gnd.n5172 gnd.n5171 0.152939
R21910 gnd.n5174 gnd.n5172 0.152939
R21911 gnd.n5174 gnd.n5173 0.152939
R21912 gnd.n5173 gnd.n2836 0.152939
R21913 gnd.n5191 gnd.n5190 0.152939
R21914 gnd.n5192 gnd.n5191 0.152939
R21915 gnd.n5192 gnd.n2832 0.152939
R21916 gnd.n5198 gnd.n2832 0.152939
R21917 gnd.n5199 gnd.n5198 0.152939
R21918 gnd.n5200 gnd.n5199 0.152939
R21919 gnd.n5489 gnd.n5488 0.152939
R21920 gnd.n5498 gnd.n5488 0.152939
R21921 gnd.n5499 gnd.n5498 0.152939
R21922 gnd.n5500 gnd.n5499 0.152939
R21923 gnd.n5500 gnd.n5481 0.152939
R21924 gnd.n5536 gnd.n5481 0.152939
R21925 gnd.n5536 gnd.n5535 0.152939
R21926 gnd.n5535 gnd.n5534 0.152939
R21927 gnd.n5534 gnd.n5482 0.152939
R21928 gnd.n5530 gnd.n5482 0.152939
R21929 gnd.n5530 gnd.n5529 0.152939
R21930 gnd.n5529 gnd.n5528 0.152939
R21931 gnd.n5528 gnd.n5442 0.152939
R21932 gnd.n5567 gnd.n5442 0.152939
R21933 gnd.n5568 gnd.n5567 0.152939
R21934 gnd.n5577 gnd.n5568 0.152939
R21935 gnd.n5577 gnd.n5576 0.152939
R21936 gnd.n5576 gnd.n5575 0.152939
R21937 gnd.n5575 gnd.n5569 0.152939
R21938 gnd.n5569 gnd.n63 0.152939
R21939 gnd.n7407 gnd.n7406 0.145814
R21940 gnd.n4175 gnd.n4174 0.145814
R21941 gnd.n4175 gnd.n3707 0.145814
R21942 gnd.n7407 gnd.n63 0.145814
R21943 gnd.n3794 gnd.n3764 0.128549
R21944 gnd.n5556 gnd.n78 0.128549
R21945 gnd.n3590 gnd.n3415 0.128549
R21946 gnd.n5200 gnd.n2814 0.128549
R21947 gnd.n1120 gnd.n0 0.127478
R21948 gnd.n1700 gnd.n1699 0.0767195
R21949 gnd.n1699 gnd.n1698 0.0767195
R21950 gnd.n3415 gnd.n2538 0.063
R21951 gnd.n5811 gnd.n2814 0.063
R21952 gnd.n5811 gnd.n5810 0.0538288
R21953 gnd.n7343 gnd.n173 0.0538288
R21954 gnd.n4108 gnd.n4106 0.0538288
R21955 gnd.n6083 gnd.n2538 0.0538288
R21956 gnd.n2268 gnd.n883 0.0477147
R21957 gnd.n1463 gnd.n1351 0.0442063
R21958 gnd.n1464 gnd.n1463 0.0442063
R21959 gnd.n1465 gnd.n1464 0.0442063
R21960 gnd.n1465 gnd.n1340 0.0442063
R21961 gnd.n1479 gnd.n1340 0.0442063
R21962 gnd.n1480 gnd.n1479 0.0442063
R21963 gnd.n1481 gnd.n1480 0.0442063
R21964 gnd.n1481 gnd.n1327 0.0442063
R21965 gnd.n1525 gnd.n1327 0.0442063
R21966 gnd.n1526 gnd.n1525 0.0442063
R21967 gnd.n1528 gnd.n1261 0.0344674
R21968 gnd.n5810 gnd.n2816 0.0344674
R21969 gnd.n5492 gnd.n2816 0.0344674
R21970 gnd.n5492 gnd.n5336 0.0344674
R21971 gnd.n5337 gnd.n5336 0.0344674
R21972 gnd.n5338 gnd.n5337 0.0344674
R21973 gnd.n5507 gnd.n5338 0.0344674
R21974 gnd.n5507 gnd.n5356 0.0344674
R21975 gnd.n5357 gnd.n5356 0.0344674
R21976 gnd.n5358 gnd.n5357 0.0344674
R21977 gnd.n5514 gnd.n5358 0.0344674
R21978 gnd.n5514 gnd.n5376 0.0344674
R21979 gnd.n5377 gnd.n5376 0.0344674
R21980 gnd.n5378 gnd.n5377 0.0344674
R21981 gnd.n5520 gnd.n5378 0.0344674
R21982 gnd.n5520 gnd.n5395 0.0344674
R21983 gnd.n5396 gnd.n5395 0.0344674
R21984 gnd.n5397 gnd.n5396 0.0344674
R21985 gnd.n5585 gnd.n5397 0.0344674
R21986 gnd.n5588 gnd.n5585 0.0344674
R21987 gnd.n5589 gnd.n5588 0.0344674
R21988 gnd.n5589 gnd.n5421 0.0344674
R21989 gnd.n5422 gnd.n5421 0.0344674
R21990 gnd.n5423 gnd.n5422 0.0344674
R21991 gnd.n5424 gnd.n5423 0.0344674
R21992 gnd.n5604 gnd.n5424 0.0344674
R21993 gnd.n5604 gnd.n92 0.0344674
R21994 gnd.n93 gnd.n92 0.0344674
R21995 gnd.n94 gnd.n93 0.0344674
R21996 gnd.n5616 gnd.n94 0.0344674
R21997 gnd.n5616 gnd.n111 0.0344674
R21998 gnd.n112 gnd.n111 0.0344674
R21999 gnd.n113 gnd.n112 0.0344674
R22000 gnd.n5623 gnd.n113 0.0344674
R22001 gnd.n5623 gnd.n132 0.0344674
R22002 gnd.n133 gnd.n132 0.0344674
R22003 gnd.n134 gnd.n133 0.0344674
R22004 gnd.n5630 gnd.n134 0.0344674
R22005 gnd.n5630 gnd.n152 0.0344674
R22006 gnd.n153 gnd.n152 0.0344674
R22007 gnd.n154 gnd.n153 0.0344674
R22008 gnd.n172 gnd.n154 0.0344674
R22009 gnd.n7343 gnd.n172 0.0344674
R22010 gnd.n4109 gnd.n4108 0.0344674
R22011 gnd.n4109 gnd.n2341 0.0344674
R22012 gnd.n2342 gnd.n2341 0.0344674
R22013 gnd.n2343 gnd.n2342 0.0344674
R22014 gnd.n3814 gnd.n2343 0.0344674
R22015 gnd.n3814 gnd.n2361 0.0344674
R22016 gnd.n2362 gnd.n2361 0.0344674
R22017 gnd.n2363 gnd.n2362 0.0344674
R22018 gnd.n3727 gnd.n2363 0.0344674
R22019 gnd.n3727 gnd.n2382 0.0344674
R22020 gnd.n2383 gnd.n2382 0.0344674
R22021 gnd.n2384 gnd.n2383 0.0344674
R22022 gnd.n3722 gnd.n2384 0.0344674
R22023 gnd.n3722 gnd.n2402 0.0344674
R22024 gnd.n2403 gnd.n2402 0.0344674
R22025 gnd.n2404 gnd.n2403 0.0344674
R22026 gnd.n3716 gnd.n2404 0.0344674
R22027 gnd.n3716 gnd.n2421 0.0344674
R22028 gnd.n2422 gnd.n2421 0.0344674
R22029 gnd.n2423 gnd.n2422 0.0344674
R22030 gnd.n3711 gnd.n2423 0.0344674
R22031 gnd.n3711 gnd.n2438 0.0344674
R22032 gnd.n2439 gnd.n2438 0.0344674
R22033 gnd.n2440 gnd.n2439 0.0344674
R22034 gnd.n3705 gnd.n2440 0.0344674
R22035 gnd.n3705 gnd.n2456 0.0344674
R22036 gnd.n2457 gnd.n2456 0.0344674
R22037 gnd.n2458 gnd.n2457 0.0344674
R22038 gnd.n3700 gnd.n2458 0.0344674
R22039 gnd.n3700 gnd.n2476 0.0344674
R22040 gnd.n2477 gnd.n2476 0.0344674
R22041 gnd.n2478 gnd.n2477 0.0344674
R22042 gnd.n4212 gnd.n2478 0.0344674
R22043 gnd.n4212 gnd.n2497 0.0344674
R22044 gnd.n2498 gnd.n2497 0.0344674
R22045 gnd.n2499 gnd.n2498 0.0344674
R22046 gnd.n4221 gnd.n2499 0.0344674
R22047 gnd.n4221 gnd.n2518 0.0344674
R22048 gnd.n2519 gnd.n2518 0.0344674
R22049 gnd.n2520 gnd.n2519 0.0344674
R22050 gnd.n2537 gnd.n2520 0.0344674
R22051 gnd.n6083 gnd.n2537 0.0344674
R22052 gnd.n3596 gnd.n3595 0.0344674
R22053 gnd.n5206 gnd.n5205 0.0344674
R22054 gnd.n6074 gnd.n6073 0.029712
R22055 gnd.n5267 gnd.n2679 0.029712
R22056 gnd.n1548 gnd.n1547 0.0269946
R22057 gnd.n1550 gnd.n1549 0.0269946
R22058 gnd.n1256 gnd.n1254 0.0269946
R22059 gnd.n1560 gnd.n1558 0.0269946
R22060 gnd.n1559 gnd.n1235 0.0269946
R22061 gnd.n1579 gnd.n1578 0.0269946
R22062 gnd.n1581 gnd.n1580 0.0269946
R22063 gnd.n1230 gnd.n1229 0.0269946
R22064 gnd.n1591 gnd.n1225 0.0269946
R22065 gnd.n1590 gnd.n1227 0.0269946
R22066 gnd.n1226 gnd.n1208 0.0269946
R22067 gnd.n1611 gnd.n1209 0.0269946
R22068 gnd.n1610 gnd.n1210 0.0269946
R22069 gnd.n1644 gnd.n1185 0.0269946
R22070 gnd.n1646 gnd.n1645 0.0269946
R22071 gnd.n1647 gnd.n1132 0.0269946
R22072 gnd.n1180 gnd.n1133 0.0269946
R22073 gnd.n1182 gnd.n1134 0.0269946
R22074 gnd.n1657 gnd.n1656 0.0269946
R22075 gnd.n1659 gnd.n1658 0.0269946
R22076 gnd.n1660 gnd.n1154 0.0269946
R22077 gnd.n1662 gnd.n1155 0.0269946
R22078 gnd.n1665 gnd.n1156 0.0269946
R22079 gnd.n1668 gnd.n1667 0.0269946
R22080 gnd.n1670 gnd.n1669 0.0269946
R22081 gnd.n1735 gnd.n1055 0.0269946
R22082 gnd.n1737 gnd.n1736 0.0269946
R22083 gnd.n1746 gnd.n1048 0.0269946
R22084 gnd.n1748 gnd.n1747 0.0269946
R22085 gnd.n1749 gnd.n1046 0.0269946
R22086 gnd.n1756 gnd.n1752 0.0269946
R22087 gnd.n1755 gnd.n1754 0.0269946
R22088 gnd.n1753 gnd.n1025 0.0269946
R22089 gnd.n1778 gnd.n1026 0.0269946
R22090 gnd.n1777 gnd.n1027 0.0269946
R22091 gnd.n1822 gnd.n1001 0.0269946
R22092 gnd.n1824 gnd.n1823 0.0269946
R22093 gnd.n1833 gnd.n994 0.0269946
R22094 gnd.n1835 gnd.n1834 0.0269946
R22095 gnd.n1836 gnd.n992 0.0269946
R22096 gnd.n1843 gnd.n1839 0.0269946
R22097 gnd.n1842 gnd.n1841 0.0269946
R22098 gnd.n1840 gnd.n971 0.0269946
R22099 gnd.n1865 gnd.n972 0.0269946
R22100 gnd.n1864 gnd.n973 0.0269946
R22101 gnd.n1911 gnd.n947 0.0269946
R22102 gnd.n1913 gnd.n1912 0.0269946
R22103 gnd.n1922 gnd.n940 0.0269946
R22104 gnd.n2181 gnd.n938 0.0269946
R22105 gnd.n2186 gnd.n2184 0.0269946
R22106 gnd.n2185 gnd.n919 0.0269946
R22107 gnd.n2210 gnd.n2209 0.0269946
R22108 gnd.n5429 gnd.n78 0.0248902
R22109 gnd.n3794 gnd.n3761 0.0248902
R22110 gnd.n3599 gnd.n3598 0.0225788
R22111 gnd.n3604 gnd.n3413 0.0225788
R22112 gnd.n3605 gnd.n3410 0.0225788
R22113 gnd.n3611 gnd.n3610 0.0225788
R22114 gnd.n3616 gnd.n3406 0.0225788
R22115 gnd.n3617 gnd.n3402 0.0225788
R22116 gnd.n3623 gnd.n3622 0.0225788
R22117 gnd.n3628 gnd.n3400 0.0225788
R22118 gnd.n3629 gnd.n3398 0.0225788
R22119 gnd.n3635 gnd.n3634 0.0225788
R22120 gnd.n3640 gnd.n3394 0.0225788
R22121 gnd.n3641 gnd.n3390 0.0225788
R22122 gnd.n3647 gnd.n3646 0.0225788
R22123 gnd.n3652 gnd.n3388 0.0225788
R22124 gnd.n3653 gnd.n3386 0.0225788
R22125 gnd.n3659 gnd.n3658 0.0225788
R22126 gnd.n3665 gnd.n3380 0.0225788
R22127 gnd.n3667 gnd.n3666 0.0225788
R22128 gnd.n6073 gnd.n2545 0.0225788
R22129 gnd.n2827 gnd.n2823 0.0225788
R22130 gnd.n5314 gnd.n5313 0.0225788
R22131 gnd.n5310 gnd.n2828 0.0225788
R22132 gnd.n5309 gnd.n5214 0.0225788
R22133 gnd.n5306 gnd.n5305 0.0225788
R22134 gnd.n5302 gnd.n5218 0.0225788
R22135 gnd.n5301 gnd.n5222 0.0225788
R22136 gnd.n5298 gnd.n5297 0.0225788
R22137 gnd.n5294 gnd.n5228 0.0225788
R22138 gnd.n5293 gnd.n5234 0.0225788
R22139 gnd.n5290 gnd.n5289 0.0225788
R22140 gnd.n5286 gnd.n5238 0.0225788
R22141 gnd.n5285 gnd.n5242 0.0225788
R22142 gnd.n5282 gnd.n5281 0.0225788
R22143 gnd.n5278 gnd.n5248 0.0225788
R22144 gnd.n5277 gnd.n5254 0.0225788
R22145 gnd.n5274 gnd.n5273 0.0225788
R22146 gnd.n5270 gnd.n5261 0.0225788
R22147 gnd.n5269 gnd.n5267 0.0225788
R22148 gnd.n5937 gnd.n2679 0.0218415
R22149 gnd.n6074 gnd.n2544 0.0218415
R22150 gnd.n1528 gnd.n1527 0.0202011
R22151 gnd.n1527 gnd.n1526 0.0148637
R22152 gnd.n2179 gnd.n1923 0.0144266
R22153 gnd.n2180 gnd.n2179 0.0130679
R22154 gnd.n3598 gnd.n3596 0.0123886
R22155 gnd.n3599 gnd.n3413 0.0123886
R22156 gnd.n3605 gnd.n3604 0.0123886
R22157 gnd.n3610 gnd.n3410 0.0123886
R22158 gnd.n3611 gnd.n3406 0.0123886
R22159 gnd.n3617 gnd.n3616 0.0123886
R22160 gnd.n3622 gnd.n3402 0.0123886
R22161 gnd.n3623 gnd.n3400 0.0123886
R22162 gnd.n3629 gnd.n3628 0.0123886
R22163 gnd.n3634 gnd.n3398 0.0123886
R22164 gnd.n3635 gnd.n3394 0.0123886
R22165 gnd.n3641 gnd.n3640 0.0123886
R22166 gnd.n3646 gnd.n3390 0.0123886
R22167 gnd.n3647 gnd.n3388 0.0123886
R22168 gnd.n3653 gnd.n3652 0.0123886
R22169 gnd.n3658 gnd.n3386 0.0123886
R22170 gnd.n3659 gnd.n3380 0.0123886
R22171 gnd.n3667 gnd.n3665 0.0123886
R22172 gnd.n3666 gnd.n2545 0.0123886
R22173 gnd.n5206 gnd.n2823 0.0123886
R22174 gnd.n5314 gnd.n2827 0.0123886
R22175 gnd.n5313 gnd.n2828 0.0123886
R22176 gnd.n5310 gnd.n5309 0.0123886
R22177 gnd.n5306 gnd.n5214 0.0123886
R22178 gnd.n5305 gnd.n5218 0.0123886
R22179 gnd.n5302 gnd.n5301 0.0123886
R22180 gnd.n5298 gnd.n5222 0.0123886
R22181 gnd.n5297 gnd.n5228 0.0123886
R22182 gnd.n5294 gnd.n5293 0.0123886
R22183 gnd.n5290 gnd.n5234 0.0123886
R22184 gnd.n5289 gnd.n5238 0.0123886
R22185 gnd.n5286 gnd.n5285 0.0123886
R22186 gnd.n5282 gnd.n5242 0.0123886
R22187 gnd.n5281 gnd.n5248 0.0123886
R22188 gnd.n5278 gnd.n5277 0.0123886
R22189 gnd.n5274 gnd.n5254 0.0123886
R22190 gnd.n5273 gnd.n5261 0.0123886
R22191 gnd.n5270 gnd.n5269 0.0123886
R22192 gnd.n1547 gnd.n1261 0.00797283
R22193 gnd.n1549 gnd.n1548 0.00797283
R22194 gnd.n1550 gnd.n1256 0.00797283
R22195 gnd.n1558 gnd.n1254 0.00797283
R22196 gnd.n1560 gnd.n1559 0.00797283
R22197 gnd.n1578 gnd.n1235 0.00797283
R22198 gnd.n1580 gnd.n1579 0.00797283
R22199 gnd.n1581 gnd.n1230 0.00797283
R22200 gnd.n1229 gnd.n1225 0.00797283
R22201 gnd.n1591 gnd.n1590 0.00797283
R22202 gnd.n1227 gnd.n1226 0.00797283
R22203 gnd.n1209 gnd.n1208 0.00797283
R22204 gnd.n1611 gnd.n1610 0.00797283
R22205 gnd.n1210 gnd.n1185 0.00797283
R22206 gnd.n1645 gnd.n1644 0.00797283
R22207 gnd.n1647 gnd.n1646 0.00797283
R22208 gnd.n1180 gnd.n1132 0.00797283
R22209 gnd.n1182 gnd.n1133 0.00797283
R22210 gnd.n1656 gnd.n1134 0.00797283
R22211 gnd.n1658 gnd.n1657 0.00797283
R22212 gnd.n1660 gnd.n1659 0.00797283
R22213 gnd.n1662 gnd.n1154 0.00797283
R22214 gnd.n1665 gnd.n1155 0.00797283
R22215 gnd.n1667 gnd.n1156 0.00797283
R22216 gnd.n1670 gnd.n1668 0.00797283
R22217 gnd.n1669 gnd.n1055 0.00797283
R22218 gnd.n1737 gnd.n1735 0.00797283
R22219 gnd.n1736 gnd.n1048 0.00797283
R22220 gnd.n1747 gnd.n1746 0.00797283
R22221 gnd.n1749 gnd.n1748 0.00797283
R22222 gnd.n1752 gnd.n1046 0.00797283
R22223 gnd.n1756 gnd.n1755 0.00797283
R22224 gnd.n1754 gnd.n1753 0.00797283
R22225 gnd.n1026 gnd.n1025 0.00797283
R22226 gnd.n1778 gnd.n1777 0.00797283
R22227 gnd.n1027 gnd.n1001 0.00797283
R22228 gnd.n1824 gnd.n1822 0.00797283
R22229 gnd.n1823 gnd.n994 0.00797283
R22230 gnd.n1834 gnd.n1833 0.00797283
R22231 gnd.n1836 gnd.n1835 0.00797283
R22232 gnd.n1839 gnd.n992 0.00797283
R22233 gnd.n1843 gnd.n1842 0.00797283
R22234 gnd.n1841 gnd.n1840 0.00797283
R22235 gnd.n972 gnd.n971 0.00797283
R22236 gnd.n1865 gnd.n1864 0.00797283
R22237 gnd.n973 gnd.n947 0.00797283
R22238 gnd.n1913 gnd.n1911 0.00797283
R22239 gnd.n1912 gnd.n940 0.00797283
R22240 gnd.n1923 gnd.n1922 0.00797283
R22241 gnd.n2181 gnd.n2180 0.00797283
R22242 gnd.n2184 gnd.n938 0.00797283
R22243 gnd.n2186 gnd.n2185 0.00797283
R22244 gnd.n2209 gnd.n919 0.00797283
R22245 gnd.n2210 gnd.n883 0.00797283
R22246 gnd.n3595 gnd.n3415 0.00593478
R22247 gnd.n5205 gnd.n2814 0.00593478
R22248 a_n2650_13878.n131 a_n2650_13878.t6 512.366
R22249 a_n2650_13878.n130 a_n2650_13878.t30 512.366
R22250 a_n2650_13878.n70 a_n2650_13878.t42 512.366
R22251 a_n2650_13878.n129 a_n2650_13878.t4 512.366
R22252 a_n2650_13878.n128 a_n2650_13878.t24 512.366
R22253 a_n2650_13878.n71 a_n2650_13878.t32 512.366
R22254 a_n2650_13878.n127 a_n2650_13878.t10 512.366
R22255 a_n2650_13878.n126 a_n2650_13878.t8 512.366
R22256 a_n2650_13878.n72 a_n2650_13878.t38 512.366
R22257 a_n2650_13878.n117 a_n2650_13878.t90 512.366
R22258 a_n2650_13878.n116 a_n2650_13878.t69 512.366
R22259 a_n2650_13878.n73 a_n2650_13878.t74 512.366
R22260 a_n2650_13878.n115 a_n2650_13878.t63 512.366
R22261 a_n2650_13878.n114 a_n2650_13878.t79 512.366
R22262 a_n2650_13878.n74 a_n2650_13878.t87 512.366
R22263 a_n2650_13878.n113 a_n2650_13878.t88 512.366
R22264 a_n2650_13878.n112 a_n2650_13878.t58 512.366
R22265 a_n2650_13878.n75 a_n2650_13878.t71 512.366
R22266 a_n2650_13878.n91 a_n2650_13878.t14 512.366
R22267 a_n2650_13878.n92 a_n2650_13878.t26 512.366
R22268 a_n2650_13878.n81 a_n2650_13878.t40 512.366
R22269 a_n2650_13878.n93 a_n2650_13878.t36 512.366
R22270 a_n2650_13878.n94 a_n2650_13878.t18 512.366
R22271 a_n2650_13878.n95 a_n2650_13878.t28 512.366
R22272 a_n2650_13878.n96 a_n2650_13878.t22 512.366
R22273 a_n2650_13878.n80 a_n2650_13878.t20 512.366
R22274 a_n2650_13878.n97 a_n2650_13878.t12 512.366
R22275 a_n2650_13878.n84 a_n2650_13878.t62 512.366
R22276 a_n2650_13878.n85 a_n2650_13878.t85 512.366
R22277 a_n2650_13878.n83 a_n2650_13878.t86 512.366
R22278 a_n2650_13878.n86 a_n2650_13878.t60 512.366
R22279 a_n2650_13878.n87 a_n2650_13878.t82 512.366
R22280 a_n2650_13878.n88 a_n2650_13878.t83 512.366
R22281 a_n2650_13878.n89 a_n2650_13878.t57 512.366
R22282 a_n2650_13878.n82 a_n2650_13878.t68 512.366
R22283 a_n2650_13878.n90 a_n2650_13878.t78 512.366
R22284 a_n2650_13878.n109 a_n2650_13878.t76 512.366
R22285 a_n2650_13878.n99 a_n2650_13878.t66 512.366
R22286 a_n2650_13878.n110 a_n2650_13878.t56 512.366
R22287 a_n2650_13878.n107 a_n2650_13878.t84 512.366
R22288 a_n2650_13878.n100 a_n2650_13878.t73 512.366
R22289 a_n2650_13878.n108 a_n2650_13878.t72 512.366
R22290 a_n2650_13878.n105 a_n2650_13878.t80 512.366
R22291 a_n2650_13878.n101 a_n2650_13878.t64 512.366
R22292 a_n2650_13878.n106 a_n2650_13878.t65 512.366
R22293 a_n2650_13878.n103 a_n2650_13878.t67 512.366
R22294 a_n2650_13878.n102 a_n2650_13878.t77 512.366
R22295 a_n2650_13878.n104 a_n2650_13878.t91 512.366
R22296 a_n2650_13878.n33 a_n2650_13878.n69 70.1674
R22297 a_n2650_13878.n7 a_n2650_13878.n62 70.1674
R22298 a_n2650_13878.n20 a_n2650_13878.n47 70.1674
R22299 a_n2650_13878.n24 a_n2650_13878.n40 70.1674
R22300 a_n2650_13878.n90 a_n2650_13878.n40 20.9683
R22301 a_n2650_13878.n39 a_n2650_13878.n24 74.73
R22302 a_n2650_13878.n39 a_n2650_13878.n82 11.843
R22303 a_n2650_13878.n23 a_n2650_13878.n38 80.4688
R22304 a_n2650_13878.n89 a_n2650_13878.n38 0.365327
R22305 a_n2650_13878.n37 a_n2650_13878.n23 75.0448
R22306 a_n2650_13878.n25 a_n2650_13878.n36 70.1674
R22307 a_n2650_13878.n86 a_n2650_13878.n36 20.9683
R22308 a_n2650_13878.n35 a_n2650_13878.n25 70.3058
R22309 a_n2650_13878.n35 a_n2650_13878.n83 20.6913
R22310 a_n2650_13878.n26 a_n2650_13878.n34 75.3623
R22311 a_n2650_13878.n85 a_n2650_13878.n34 10.5784
R22312 a_n2650_13878.n84 a_n2650_13878.n26 161.3
R22313 a_n2650_13878.n97 a_n2650_13878.n47 20.9683
R22314 a_n2650_13878.n46 a_n2650_13878.n20 74.73
R22315 a_n2650_13878.n46 a_n2650_13878.n80 11.843
R22316 a_n2650_13878.n19 a_n2650_13878.n45 80.4688
R22317 a_n2650_13878.n96 a_n2650_13878.n45 0.365327
R22318 a_n2650_13878.n44 a_n2650_13878.n19 75.0448
R22319 a_n2650_13878.n21 a_n2650_13878.n43 70.1674
R22320 a_n2650_13878.n93 a_n2650_13878.n43 20.9683
R22321 a_n2650_13878.n42 a_n2650_13878.n21 70.3058
R22322 a_n2650_13878.n42 a_n2650_13878.n81 20.6913
R22323 a_n2650_13878.n22 a_n2650_13878.n41 75.3623
R22324 a_n2650_13878.n92 a_n2650_13878.n41 10.5784
R22325 a_n2650_13878.n91 a_n2650_13878.n22 161.3
R22326 a_n2650_13878.n10 a_n2650_13878.n55 70.1674
R22327 a_n2650_13878.n12 a_n2650_13878.n53 70.1674
R22328 a_n2650_13878.n14 a_n2650_13878.n51 70.1674
R22329 a_n2650_13878.n17 a_n2650_13878.n49 70.1674
R22330 a_n2650_13878.n104 a_n2650_13878.n49 20.9683
R22331 a_n2650_13878.n48 a_n2650_13878.n18 75.0448
R22332 a_n2650_13878.n48 a_n2650_13878.n102 11.2134
R22333 a_n2650_13878.n18 a_n2650_13878.n103 161.3
R22334 a_n2650_13878.n106 a_n2650_13878.n51 20.9683
R22335 a_n2650_13878.n50 a_n2650_13878.n15 75.0448
R22336 a_n2650_13878.n50 a_n2650_13878.n101 11.2134
R22337 a_n2650_13878.n15 a_n2650_13878.n105 161.3
R22338 a_n2650_13878.n108 a_n2650_13878.n53 20.9683
R22339 a_n2650_13878.n52 a_n2650_13878.n13 75.0448
R22340 a_n2650_13878.n52 a_n2650_13878.n100 11.2134
R22341 a_n2650_13878.n13 a_n2650_13878.n107 161.3
R22342 a_n2650_13878.n110 a_n2650_13878.n55 20.9683
R22343 a_n2650_13878.n54 a_n2650_13878.n11 75.0448
R22344 a_n2650_13878.n54 a_n2650_13878.n99 11.2134
R22345 a_n2650_13878.n11 a_n2650_13878.n109 161.3
R22346 a_n2650_13878.n62 a_n2650_13878.n75 20.9683
R22347 a_n2650_13878.n61 a_n2650_13878.n7 74.73
R22348 a_n2650_13878.n112 a_n2650_13878.n61 11.843
R22349 a_n2650_13878.n60 a_n2650_13878.n6 80.4688
R22350 a_n2650_13878.n60 a_n2650_13878.n113 0.365327
R22351 a_n2650_13878.n6 a_n2650_13878.n59 75.0448
R22352 a_n2650_13878.n58 a_n2650_13878.n8 70.1674
R22353 a_n2650_13878.n115 a_n2650_13878.n58 20.9683
R22354 a_n2650_13878.n8 a_n2650_13878.n57 70.3058
R22355 a_n2650_13878.n57 a_n2650_13878.n73 20.6913
R22356 a_n2650_13878.n56 a_n2650_13878.n9 75.3623
R22357 a_n2650_13878.n116 a_n2650_13878.n56 10.5784
R22358 a_n2650_13878.n9 a_n2650_13878.n117 161.3
R22359 a_n2650_13878.n69 a_n2650_13878.n72 20.9683
R22360 a_n2650_13878.n68 a_n2650_13878.n33 74.73
R22361 a_n2650_13878.n126 a_n2650_13878.n68 11.843
R22362 a_n2650_13878.n67 a_n2650_13878.n4 80.4688
R22363 a_n2650_13878.n67 a_n2650_13878.n127 0.365327
R22364 a_n2650_13878.n4 a_n2650_13878.n66 75.0448
R22365 a_n2650_13878.n65 a_n2650_13878.n3 70.1674
R22366 a_n2650_13878.n129 a_n2650_13878.n65 20.9683
R22367 a_n2650_13878.n3 a_n2650_13878.n64 70.3058
R22368 a_n2650_13878.n64 a_n2650_13878.n70 20.6913
R22369 a_n2650_13878.n63 a_n2650_13878.n5 75.3623
R22370 a_n2650_13878.n130 a_n2650_13878.n63 10.5784
R22371 a_n2650_13878.n5 a_n2650_13878.n131 161.3
R22372 a_n2650_13878.n1 a_n2650_13878.n124 81.4626
R22373 a_n2650_13878.n2 a_n2650_13878.n120 81.4626
R22374 a_n2650_13878.n2 a_n2650_13878.n118 81.4626
R22375 a_n2650_13878.n1 a_n2650_13878.n125 80.9324
R22376 a_n2650_13878.n1 a_n2650_13878.n123 80.9324
R22377 a_n2650_13878.n0 a_n2650_13878.n122 80.9324
R22378 a_n2650_13878.n2 a_n2650_13878.n121 80.9324
R22379 a_n2650_13878.n2 a_n2650_13878.n119 80.9324
R22380 a_n2650_13878.n30 a_n2650_13878.t17 74.6477
R22381 a_n2650_13878.n27 a_n2650_13878.t15 74.6477
R22382 a_n2650_13878.n31 a_n2650_13878.t7 74.2899
R22383 a_n2650_13878.n29 a_n2650_13878.t35 74.2897
R22384 a_n2650_13878.n30 a_n2650_13878.n134 70.6783
R22385 a_n2650_13878.n30 a_n2650_13878.n135 70.6783
R22386 a_n2650_13878.n32 a_n2650_13878.n133 70.6783
R22387 a_n2650_13878.n29 a_n2650_13878.n79 70.6783
R22388 a_n2650_13878.n28 a_n2650_13878.n78 70.6783
R22389 a_n2650_13878.n28 a_n2650_13878.n77 70.6783
R22390 a_n2650_13878.n27 a_n2650_13878.n76 70.6783
R22391 a_n2650_13878.n136 a_n2650_13878.n32 70.6782
R22392 a_n2650_13878.n131 a_n2650_13878.n130 48.2005
R22393 a_n2650_13878.n65 a_n2650_13878.n128 20.9683
R22394 a_n2650_13878.n127 a_n2650_13878.n71 48.2005
R22395 a_n2650_13878.t16 a_n2650_13878.n69 533.335
R22396 a_n2650_13878.n117 a_n2650_13878.n116 48.2005
R22397 a_n2650_13878.n58 a_n2650_13878.n114 20.9683
R22398 a_n2650_13878.n113 a_n2650_13878.n74 48.2005
R22399 a_n2650_13878.t61 a_n2650_13878.n62 533.335
R22400 a_n2650_13878.n92 a_n2650_13878.n91 48.2005
R22401 a_n2650_13878.n94 a_n2650_13878.n43 20.9683
R22402 a_n2650_13878.n96 a_n2650_13878.n95 48.2005
R22403 a_n2650_13878.t34 a_n2650_13878.n47 533.335
R22404 a_n2650_13878.n85 a_n2650_13878.n84 48.2005
R22405 a_n2650_13878.n87 a_n2650_13878.n36 20.9683
R22406 a_n2650_13878.n89 a_n2650_13878.n88 48.2005
R22407 a_n2650_13878.t59 a_n2650_13878.n40 533.335
R22408 a_n2650_13878.n109 a_n2650_13878.n99 48.2005
R22409 a_n2650_13878.t81 a_n2650_13878.n55 533.335
R22410 a_n2650_13878.n107 a_n2650_13878.n100 48.2005
R22411 a_n2650_13878.t89 a_n2650_13878.n53 533.335
R22412 a_n2650_13878.n105 a_n2650_13878.n101 48.2005
R22413 a_n2650_13878.t75 a_n2650_13878.n51 533.335
R22414 a_n2650_13878.n103 a_n2650_13878.n102 48.2005
R22415 a_n2650_13878.t70 a_n2650_13878.n49 533.335
R22416 a_n2650_13878.n129 a_n2650_13878.n64 21.4216
R22417 a_n2650_13878.n115 a_n2650_13878.n57 21.4216
R22418 a_n2650_13878.n93 a_n2650_13878.n42 21.4216
R22419 a_n2650_13878.n86 a_n2650_13878.n35 21.4216
R22420 a_n2650_13878.n68 a_n2650_13878.n72 34.4824
R22421 a_n2650_13878.n61 a_n2650_13878.n75 34.4824
R22422 a_n2650_13878.n97 a_n2650_13878.n46 34.4824
R22423 a_n2650_13878.n90 a_n2650_13878.n39 34.4824
R22424 a_n2650_13878.n128 a_n2650_13878.n66 35.3134
R22425 a_n2650_13878.n66 a_n2650_13878.n71 11.2134
R22426 a_n2650_13878.n114 a_n2650_13878.n59 35.3134
R22427 a_n2650_13878.n59 a_n2650_13878.n74 11.2134
R22428 a_n2650_13878.n94 a_n2650_13878.n44 35.3134
R22429 a_n2650_13878.n95 a_n2650_13878.n44 11.2134
R22430 a_n2650_13878.n87 a_n2650_13878.n37 35.3134
R22431 a_n2650_13878.n88 a_n2650_13878.n37 11.2134
R22432 a_n2650_13878.n110 a_n2650_13878.n54 35.3134
R22433 a_n2650_13878.n108 a_n2650_13878.n52 35.3134
R22434 a_n2650_13878.n106 a_n2650_13878.n50 35.3134
R22435 a_n2650_13878.n104 a_n2650_13878.n48 35.3134
R22436 a_n2650_13878.n33 a_n2650_13878.n1 23.891
R22437 a_n2650_13878.n63 a_n2650_13878.n70 36.139
R22438 a_n2650_13878.n56 a_n2650_13878.n73 36.139
R22439 a_n2650_13878.n81 a_n2650_13878.n41 36.139
R22440 a_n2650_13878.n83 a_n2650_13878.n34 36.139
R22441 a_n2650_13878.n26 a_n2650_13878.n16 13.3641
R22442 a_n2650_13878.n7 a_n2650_13878.n111 13.1596
R22443 a_n2650_13878.n132 a_n2650_13878.n5 11.8547
R22444 a_n2650_13878.n98 a_n2650_13878.n29 10.2167
R22445 a_n2650_13878.n18 a_n2650_13878.n16 9.99103
R22446 a_n2650_13878.n111 a_n2650_13878.n10 9.99103
R22447 a_n2650_13878.n98 a_n2650_13878.n20 8.01944
R22448 a_n2650_13878.n31 a_n2650_13878.n132 6.37334
R22449 a_n2650_13878.n111 a_n2650_13878.n98 5.3452
R22450 a_n2650_13878.n22 a_n2650_13878.n24 4.07247
R22451 a_n2650_13878.n33 a_n2650_13878.n9 4.06146
R22452 a_n2650_13878.n134 a_n2650_13878.t9 3.61217
R22453 a_n2650_13878.n134 a_n2650_13878.t39 3.61217
R22454 a_n2650_13878.n135 a_n2650_13878.t33 3.61217
R22455 a_n2650_13878.n135 a_n2650_13878.t11 3.61217
R22456 a_n2650_13878.n133 a_n2650_13878.t31 3.61217
R22457 a_n2650_13878.n133 a_n2650_13878.t43 3.61217
R22458 a_n2650_13878.n79 a_n2650_13878.t21 3.61217
R22459 a_n2650_13878.n79 a_n2650_13878.t13 3.61217
R22460 a_n2650_13878.n78 a_n2650_13878.t29 3.61217
R22461 a_n2650_13878.n78 a_n2650_13878.t23 3.61217
R22462 a_n2650_13878.n77 a_n2650_13878.t37 3.61217
R22463 a_n2650_13878.n77 a_n2650_13878.t19 3.61217
R22464 a_n2650_13878.n76 a_n2650_13878.t27 3.61217
R22465 a_n2650_13878.n76 a_n2650_13878.t41 3.61217
R22466 a_n2650_13878.t5 a_n2650_13878.n136 3.61217
R22467 a_n2650_13878.n136 a_n2650_13878.t25 3.61217
R22468 a_n2650_13878.n124 a_n2650_13878.t1 2.82907
R22469 a_n2650_13878.n124 a_n2650_13878.t50 2.82907
R22470 a_n2650_13878.n125 a_n2650_13878.t46 2.82907
R22471 a_n2650_13878.n125 a_n2650_13878.t51 2.82907
R22472 a_n2650_13878.n123 a_n2650_13878.t2 2.82907
R22473 a_n2650_13878.n123 a_n2650_13878.t52 2.82907
R22474 a_n2650_13878.n122 a_n2650_13878.t48 2.82907
R22475 a_n2650_13878.n122 a_n2650_13878.t53 2.82907
R22476 a_n2650_13878.n120 a_n2650_13878.t47 2.82907
R22477 a_n2650_13878.n120 a_n2650_13878.t3 2.82907
R22478 a_n2650_13878.n121 a_n2650_13878.t45 2.82907
R22479 a_n2650_13878.n121 a_n2650_13878.t44 2.82907
R22480 a_n2650_13878.n119 a_n2650_13878.t0 2.82907
R22481 a_n2650_13878.n119 a_n2650_13878.t49 2.82907
R22482 a_n2650_13878.n118 a_n2650_13878.t55 2.82907
R22483 a_n2650_13878.n118 a_n2650_13878.t54 2.82907
R22484 a_n2650_13878.n132 a_n2650_13878.n16 1.30542
R22485 a_n2650_13878.n13 a_n2650_13878.n14 1.04595
R22486 a_n2650_13878.n67 a_n2650_13878.n126 47.835
R22487 a_n2650_13878.n60 a_n2650_13878.n112 47.835
R22488 a_n2650_13878.n80 a_n2650_13878.n45 47.835
R22489 a_n2650_13878.n82 a_n2650_13878.n38 47.835
R22490 a_n2650_13878.n0 a_n2650_13878.n2 32.5247
R22491 a_n2650_13878.n24 a_n2650_13878.n23 1.13686
R22492 a_n2650_13878.n20 a_n2650_13878.n19 1.13686
R22493 a_n2650_13878.n7 a_n2650_13878.n6 1.13686
R22494 a_n2650_13878.n33 a_n2650_13878.n4 1.11
R22495 a_n2650_13878.n1 a_n2650_13878.n0 1.06084
R22496 a_n2650_13878.n25 a_n2650_13878.n26 0.758076
R22497 a_n2650_13878.n23 a_n2650_13878.n25 0.758076
R22498 a_n2650_13878.n21 a_n2650_13878.n22 0.758076
R22499 a_n2650_13878.n19 a_n2650_13878.n21 0.758076
R22500 a_n2650_13878.n18 a_n2650_13878.n17 0.758076
R22501 a_n2650_13878.n15 a_n2650_13878.n14 0.758076
R22502 a_n2650_13878.n13 a_n2650_13878.n12 0.758076
R22503 a_n2650_13878.n11 a_n2650_13878.n10 0.758076
R22504 a_n2650_13878.n9 a_n2650_13878.n8 0.758076
R22505 a_n2650_13878.n6 a_n2650_13878.n8 0.758076
R22506 a_n2650_13878.n5 a_n2650_13878.n3 0.758076
R22507 a_n2650_13878.n4 a_n2650_13878.n3 0.758076
R22508 a_n2650_13878.n32 a_n2650_13878.n30 0.716017
R22509 a_n2650_13878.n32 a_n2650_13878.n31 0.716017
R22510 a_n2650_13878.n29 a_n2650_13878.n28 0.716017
R22511 a_n2650_13878.n28 a_n2650_13878.n27 0.716017
R22512 a_n2650_13878.n15 a_n2650_13878.n17 0.67853
R22513 a_n2650_13878.n11 a_n2650_13878.n12 0.67853
R22514 a_n2472_13878.n25 a_n2472_13878.n24 98.9632
R22515 a_n2472_13878.n2 a_n2472_13878.n0 98.7517
R22516 a_n2472_13878.n20 a_n2472_13878.n19 98.6055
R22517 a_n2472_13878.n22 a_n2472_13878.n21 98.6055
R22518 a_n2472_13878.n24 a_n2472_13878.n23 98.6055
R22519 a_n2472_13878.n8 a_n2472_13878.n7 98.6055
R22520 a_n2472_13878.n6 a_n2472_13878.n5 98.6055
R22521 a_n2472_13878.n4 a_n2472_13878.n3 98.6055
R22522 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R22523 a_n2472_13878.n18 a_n2472_13878.n17 98.6054
R22524 a_n2472_13878.n10 a_n2472_13878.t21 74.6477
R22525 a_n2472_13878.n15 a_n2472_13878.t22 74.2899
R22526 a_n2472_13878.n12 a_n2472_13878.t23 74.2899
R22527 a_n2472_13878.n11 a_n2472_13878.t20 74.2899
R22528 a_n2472_13878.n14 a_n2472_13878.n13 70.6783
R22529 a_n2472_13878.n10 a_n2472_13878.n9 70.6783
R22530 a_n2472_13878.n16 a_n2472_13878.n8 15.0004
R22531 a_n2472_13878.n18 a_n2472_13878.n16 12.2917
R22532 a_n2472_13878.n16 a_n2472_13878.n15 7.67184
R22533 a_n2472_13878.n17 a_n2472_13878.t16 3.61217
R22534 a_n2472_13878.n17 a_n2472_13878.t5 3.61217
R22535 a_n2472_13878.n19 a_n2472_13878.t8 3.61217
R22536 a_n2472_13878.n19 a_n2472_13878.t9 3.61217
R22537 a_n2472_13878.n21 a_n2472_13878.t17 3.61217
R22538 a_n2472_13878.n21 a_n2472_13878.t18 3.61217
R22539 a_n2472_13878.n23 a_n2472_13878.t0 3.61217
R22540 a_n2472_13878.n23 a_n2472_13878.t10 3.61217
R22541 a_n2472_13878.n13 a_n2472_13878.t26 3.61217
R22542 a_n2472_13878.n13 a_n2472_13878.t27 3.61217
R22543 a_n2472_13878.n9 a_n2472_13878.t24 3.61217
R22544 a_n2472_13878.n9 a_n2472_13878.t25 3.61217
R22545 a_n2472_13878.n7 a_n2472_13878.t11 3.61217
R22546 a_n2472_13878.n7 a_n2472_13878.t1 3.61217
R22547 a_n2472_13878.n5 a_n2472_13878.t14 3.61217
R22548 a_n2472_13878.n5 a_n2472_13878.t3 3.61217
R22549 a_n2472_13878.n3 a_n2472_13878.t2 3.61217
R22550 a_n2472_13878.n3 a_n2472_13878.t4 3.61217
R22551 a_n2472_13878.n1 a_n2472_13878.t12 3.61217
R22552 a_n2472_13878.n1 a_n2472_13878.t6 3.61217
R22553 a_n2472_13878.n0 a_n2472_13878.t15 3.61217
R22554 a_n2472_13878.n0 a_n2472_13878.t7 3.61217
R22555 a_n2472_13878.n25 a_n2472_13878.t13 3.61217
R22556 a_n2472_13878.t19 a_n2472_13878.n25 3.61217
R22557 a_n2472_13878.n11 a_n2472_13878.n10 0.358259
R22558 a_n2472_13878.n14 a_n2472_13878.n12 0.358259
R22559 a_n2472_13878.n15 a_n2472_13878.n14 0.358259
R22560 a_n2472_13878.n24 a_n2472_13878.n22 0.358259
R22561 a_n2472_13878.n22 a_n2472_13878.n20 0.358259
R22562 a_n2472_13878.n20 a_n2472_13878.n18 0.358259
R22563 a_n2472_13878.n4 a_n2472_13878.n2 0.146627
R22564 a_n2472_13878.n6 a_n2472_13878.n4 0.146627
R22565 a_n2472_13878.n8 a_n2472_13878.n6 0.146627
R22566 a_n2472_13878.n12 a_n2472_13878.n11 0.101793
R22567 output.n41 output.n15 289.615
R22568 output.n72 output.n46 289.615
R22569 output.n104 output.n78 289.615
R22570 output.n136 output.n110 289.615
R22571 output.n77 output.n45 197.26
R22572 output.n77 output.n76 196.298
R22573 output.n109 output.n108 196.298
R22574 output.n141 output.n140 196.298
R22575 output.n42 output.n41 185
R22576 output.n40 output.n39 185
R22577 output.n19 output.n18 185
R22578 output.n34 output.n33 185
R22579 output.n32 output.n31 185
R22580 output.n23 output.n22 185
R22581 output.n26 output.n25 185
R22582 output.n73 output.n72 185
R22583 output.n71 output.n70 185
R22584 output.n50 output.n49 185
R22585 output.n65 output.n64 185
R22586 output.n63 output.n62 185
R22587 output.n54 output.n53 185
R22588 output.n57 output.n56 185
R22589 output.n105 output.n104 185
R22590 output.n103 output.n102 185
R22591 output.n82 output.n81 185
R22592 output.n97 output.n96 185
R22593 output.n95 output.n94 185
R22594 output.n86 output.n85 185
R22595 output.n89 output.n88 185
R22596 output.n137 output.n136 185
R22597 output.n135 output.n134 185
R22598 output.n114 output.n113 185
R22599 output.n129 output.n128 185
R22600 output.n127 output.n126 185
R22601 output.n118 output.n117 185
R22602 output.n121 output.n120 185
R22603 output.t1 output.n24 147.661
R22604 output.t0 output.n55 147.661
R22605 output.t18 output.n87 147.661
R22606 output.t19 output.n119 147.661
R22607 output.n41 output.n40 104.615
R22608 output.n40 output.n18 104.615
R22609 output.n33 output.n18 104.615
R22610 output.n33 output.n32 104.615
R22611 output.n32 output.n22 104.615
R22612 output.n25 output.n22 104.615
R22613 output.n72 output.n71 104.615
R22614 output.n71 output.n49 104.615
R22615 output.n64 output.n49 104.615
R22616 output.n64 output.n63 104.615
R22617 output.n63 output.n53 104.615
R22618 output.n56 output.n53 104.615
R22619 output.n104 output.n103 104.615
R22620 output.n103 output.n81 104.615
R22621 output.n96 output.n81 104.615
R22622 output.n96 output.n95 104.615
R22623 output.n95 output.n85 104.615
R22624 output.n88 output.n85 104.615
R22625 output.n136 output.n135 104.615
R22626 output.n135 output.n113 104.615
R22627 output.n128 output.n113 104.615
R22628 output.n128 output.n127 104.615
R22629 output.n127 output.n117 104.615
R22630 output.n120 output.n117 104.615
R22631 output.n1 output.t8 77.056
R22632 output.n14 output.t10 76.6694
R22633 output.n1 output.n0 72.7095
R22634 output.n3 output.n2 72.7095
R22635 output.n5 output.n4 72.7095
R22636 output.n7 output.n6 72.7095
R22637 output.n9 output.n8 72.7095
R22638 output.n11 output.n10 72.7095
R22639 output.n13 output.n12 72.7095
R22640 output.n25 output.t1 52.3082
R22641 output.n56 output.t0 52.3082
R22642 output.n88 output.t18 52.3082
R22643 output.n120 output.t19 52.3082
R22644 output.n26 output.n24 15.6674
R22645 output.n57 output.n55 15.6674
R22646 output.n89 output.n87 15.6674
R22647 output.n121 output.n119 15.6674
R22648 output.n27 output.n23 12.8005
R22649 output.n58 output.n54 12.8005
R22650 output.n90 output.n86 12.8005
R22651 output.n122 output.n118 12.8005
R22652 output.n31 output.n30 12.0247
R22653 output.n62 output.n61 12.0247
R22654 output.n94 output.n93 12.0247
R22655 output.n126 output.n125 12.0247
R22656 output.n34 output.n21 11.249
R22657 output.n65 output.n52 11.249
R22658 output.n97 output.n84 11.249
R22659 output.n129 output.n116 11.249
R22660 output.n35 output.n19 10.4732
R22661 output.n66 output.n50 10.4732
R22662 output.n98 output.n82 10.4732
R22663 output.n130 output.n114 10.4732
R22664 output.n39 output.n38 9.69747
R22665 output.n70 output.n69 9.69747
R22666 output.n102 output.n101 9.69747
R22667 output.n134 output.n133 9.69747
R22668 output.n45 output.n44 9.45567
R22669 output.n76 output.n75 9.45567
R22670 output.n108 output.n107 9.45567
R22671 output.n140 output.n139 9.45567
R22672 output.n44 output.n43 9.3005
R22673 output.n17 output.n16 9.3005
R22674 output.n38 output.n37 9.3005
R22675 output.n36 output.n35 9.3005
R22676 output.n21 output.n20 9.3005
R22677 output.n30 output.n29 9.3005
R22678 output.n28 output.n27 9.3005
R22679 output.n75 output.n74 9.3005
R22680 output.n48 output.n47 9.3005
R22681 output.n69 output.n68 9.3005
R22682 output.n67 output.n66 9.3005
R22683 output.n52 output.n51 9.3005
R22684 output.n61 output.n60 9.3005
R22685 output.n59 output.n58 9.3005
R22686 output.n107 output.n106 9.3005
R22687 output.n80 output.n79 9.3005
R22688 output.n101 output.n100 9.3005
R22689 output.n99 output.n98 9.3005
R22690 output.n84 output.n83 9.3005
R22691 output.n93 output.n92 9.3005
R22692 output.n91 output.n90 9.3005
R22693 output.n139 output.n138 9.3005
R22694 output.n112 output.n111 9.3005
R22695 output.n133 output.n132 9.3005
R22696 output.n131 output.n130 9.3005
R22697 output.n116 output.n115 9.3005
R22698 output.n125 output.n124 9.3005
R22699 output.n123 output.n122 9.3005
R22700 output.n42 output.n17 8.92171
R22701 output.n73 output.n48 8.92171
R22702 output.n105 output.n80 8.92171
R22703 output.n137 output.n112 8.92171
R22704 output output.n141 8.15037
R22705 output.n43 output.n15 8.14595
R22706 output.n74 output.n46 8.14595
R22707 output.n106 output.n78 8.14595
R22708 output.n138 output.n110 8.14595
R22709 output.n45 output.n15 5.81868
R22710 output.n76 output.n46 5.81868
R22711 output.n108 output.n78 5.81868
R22712 output.n140 output.n110 5.81868
R22713 output.n43 output.n42 5.04292
R22714 output.n74 output.n73 5.04292
R22715 output.n106 output.n105 5.04292
R22716 output.n138 output.n137 5.04292
R22717 output.n28 output.n24 4.38594
R22718 output.n59 output.n55 4.38594
R22719 output.n91 output.n87 4.38594
R22720 output.n123 output.n119 4.38594
R22721 output.n39 output.n17 4.26717
R22722 output.n70 output.n48 4.26717
R22723 output.n102 output.n80 4.26717
R22724 output.n134 output.n112 4.26717
R22725 output.n0 output.t15 3.9605
R22726 output.n0 output.t4 3.9605
R22727 output.n2 output.t6 3.9605
R22728 output.n2 output.t11 3.9605
R22729 output.n4 output.t16 3.9605
R22730 output.n4 output.t2 3.9605
R22731 output.n6 output.t3 3.9605
R22732 output.n6 output.t9 3.9605
R22733 output.n8 output.t12 3.9605
R22734 output.n8 output.t5 3.9605
R22735 output.n10 output.t7 3.9605
R22736 output.n10 output.t13 3.9605
R22737 output.n12 output.t14 3.9605
R22738 output.n12 output.t17 3.9605
R22739 output.n38 output.n19 3.49141
R22740 output.n69 output.n50 3.49141
R22741 output.n101 output.n82 3.49141
R22742 output.n133 output.n114 3.49141
R22743 output.n35 output.n34 2.71565
R22744 output.n66 output.n65 2.71565
R22745 output.n98 output.n97 2.71565
R22746 output.n130 output.n129 2.71565
R22747 output.n31 output.n21 1.93989
R22748 output.n62 output.n52 1.93989
R22749 output.n94 output.n84 1.93989
R22750 output.n126 output.n116 1.93989
R22751 output.n30 output.n23 1.16414
R22752 output.n61 output.n54 1.16414
R22753 output.n93 output.n86 1.16414
R22754 output.n125 output.n118 1.16414
R22755 output.n141 output.n109 0.962709
R22756 output.n109 output.n77 0.962709
R22757 output.n27 output.n26 0.388379
R22758 output.n58 output.n57 0.388379
R22759 output.n90 output.n89 0.388379
R22760 output.n122 output.n121 0.388379
R22761 output.n14 output.n13 0.387128
R22762 output.n13 output.n11 0.387128
R22763 output.n11 output.n9 0.387128
R22764 output.n9 output.n7 0.387128
R22765 output.n7 output.n5 0.387128
R22766 output.n5 output.n3 0.387128
R22767 output.n3 output.n1 0.387128
R22768 output.n44 output.n16 0.155672
R22769 output.n37 output.n16 0.155672
R22770 output.n37 output.n36 0.155672
R22771 output.n36 output.n20 0.155672
R22772 output.n29 output.n20 0.155672
R22773 output.n29 output.n28 0.155672
R22774 output.n75 output.n47 0.155672
R22775 output.n68 output.n47 0.155672
R22776 output.n68 output.n67 0.155672
R22777 output.n67 output.n51 0.155672
R22778 output.n60 output.n51 0.155672
R22779 output.n60 output.n59 0.155672
R22780 output.n107 output.n79 0.155672
R22781 output.n100 output.n79 0.155672
R22782 output.n100 output.n99 0.155672
R22783 output.n99 output.n83 0.155672
R22784 output.n92 output.n83 0.155672
R22785 output.n92 output.n91 0.155672
R22786 output.n139 output.n111 0.155672
R22787 output.n132 output.n111 0.155672
R22788 output.n132 output.n131 0.155672
R22789 output.n131 output.n115 0.155672
R22790 output.n124 output.n115 0.155672
R22791 output.n124 output.n123 0.155672
R22792 output output.n14 0.126227
R22793 plus.n46 plus.t9 252.611
R22794 plus.n9 plus.t11 252.611
R22795 plus.n76 plus.t4 243.97
R22796 plus.n72 plus.t12 231.093
R22797 plus.n35 plus.t7 231.093
R22798 plus.n76 plus.n75 223.454
R22799 plus.n78 plus.n77 223.454
R22800 plus.n47 plus.t5 187.445
R22801 plus.n44 plus.t18 187.445
R22802 plus.n42 plus.t17 187.445
R22803 plus.n59 plus.t13 187.445
R22804 plus.n65 plus.t14 187.445
R22805 plus.n38 plus.t10 187.445
R22806 plus.n1 plus.t6 187.445
R22807 plus.n28 plus.t16 187.445
R22808 plus.n22 plus.t15 187.445
R22809 plus.n5 plus.t20 187.445
R22810 plus.n7 plus.t19 187.445
R22811 plus.n10 plus.t8 187.445
R22812 plus.n73 plus.n72 161.3
R22813 plus.n71 plus.n37 161.3
R22814 plus.n70 plus.n69 161.3
R22815 plus.n68 plus.n67 161.3
R22816 plus.n66 plus.n39 161.3
R22817 plus.n64 plus.n63 161.3
R22818 plus.n62 plus.n40 161.3
R22819 plus.n61 plus.n60 161.3
R22820 plus.n58 plus.n41 161.3
R22821 plus.n57 plus.n56 161.3
R22822 plus.n55 plus.n54 161.3
R22823 plus.n53 plus.n43 161.3
R22824 plus.n52 plus.n51 161.3
R22825 plus.n50 plus.n49 161.3
R22826 plus.n48 plus.n45 161.3
R22827 plus.n11 plus.n8 161.3
R22828 plus.n13 plus.n12 161.3
R22829 plus.n15 plus.n14 161.3
R22830 plus.n16 plus.n6 161.3
R22831 plus.n18 plus.n17 161.3
R22832 plus.n20 plus.n19 161.3
R22833 plus.n21 plus.n4 161.3
R22834 plus.n24 plus.n23 161.3
R22835 plus.n25 plus.n3 161.3
R22836 plus.n27 plus.n26 161.3
R22837 plus.n29 plus.n2 161.3
R22838 plus.n31 plus.n30 161.3
R22839 plus.n33 plus.n32 161.3
R22840 plus.n34 plus.n0 161.3
R22841 plus.n36 plus.n35 161.3
R22842 plus.n49 plus.n48 56.5617
R22843 plus.n58 plus.n57 56.5617
R22844 plus.n67 plus.n66 56.5617
R22845 plus.n30 plus.n29 56.5617
R22846 plus.n21 plus.n20 56.5617
R22847 plus.n12 plus.n11 56.5617
R22848 plus.n71 plus.n70 46.3896
R22849 plus.n34 plus.n33 46.3896
R22850 plus.n46 plus.n45 42.8164
R22851 plus.n9 plus.n8 42.8164
R22852 plus.n54 plus.n53 42.5146
R22853 plus.n60 plus.n40 42.5146
R22854 plus.n23 plus.n3 42.5146
R22855 plus.n17 plus.n16 42.5146
R22856 plus.n53 plus.n52 38.6395
R22857 plus.n64 plus.n40 38.6395
R22858 plus.n27 plus.n3 38.6395
R22859 plus.n16 plus.n15 38.6395
R22860 plus.n47 plus.n46 38.2514
R22861 plus.n10 plus.n9 38.2514
R22862 plus.n74 plus.n73 31.491
R22863 plus.n49 plus.n44 19.9199
R22864 plus.n66 plus.n65 19.9199
R22865 plus.n29 plus.n28 19.9199
R22866 plus.n12 plus.n7 19.9199
R22867 plus.n75 plus.t1 19.8005
R22868 plus.n75 plus.t2 19.8005
R22869 plus.n77 plus.t0 19.8005
R22870 plus.n77 plus.t3 19.8005
R22871 plus.n57 plus.n42 17.9525
R22872 plus.n59 plus.n58 17.9525
R22873 plus.n22 plus.n21 17.9525
R22874 plus.n20 plus.n5 17.9525
R22875 plus.n48 plus.n47 15.9852
R22876 plus.n67 plus.n38 15.9852
R22877 plus.n30 plus.n1 15.9852
R22878 plus.n11 plus.n10 15.9852
R22879 plus.n72 plus.n71 15.3369
R22880 plus.n35 plus.n34 15.3369
R22881 plus plus.n79 14.3006
R22882 plus.n74 plus.n36 11.9494
R22883 plus.n70 plus.n38 8.60764
R22884 plus.n33 plus.n1 8.60764
R22885 plus.n54 plus.n42 6.6403
R22886 plus.n60 plus.n59 6.6403
R22887 plus.n23 plus.n22 6.6403
R22888 plus.n17 plus.n5 6.6403
R22889 plus.n79 plus.n78 5.40567
R22890 plus.n52 plus.n44 4.67295
R22891 plus.n65 plus.n64 4.67295
R22892 plus.n28 plus.n27 4.67295
R22893 plus.n15 plus.n7 4.67295
R22894 plus.n79 plus.n74 1.188
R22895 plus.n78 plus.n76 0.716017
R22896 plus.n50 plus.n45 0.189894
R22897 plus.n51 plus.n50 0.189894
R22898 plus.n51 plus.n43 0.189894
R22899 plus.n55 plus.n43 0.189894
R22900 plus.n56 plus.n55 0.189894
R22901 plus.n56 plus.n41 0.189894
R22902 plus.n61 plus.n41 0.189894
R22903 plus.n62 plus.n61 0.189894
R22904 plus.n63 plus.n62 0.189894
R22905 plus.n63 plus.n39 0.189894
R22906 plus.n68 plus.n39 0.189894
R22907 plus.n69 plus.n68 0.189894
R22908 plus.n69 plus.n37 0.189894
R22909 plus.n73 plus.n37 0.189894
R22910 plus.n36 plus.n0 0.189894
R22911 plus.n32 plus.n0 0.189894
R22912 plus.n32 plus.n31 0.189894
R22913 plus.n31 plus.n2 0.189894
R22914 plus.n26 plus.n2 0.189894
R22915 plus.n26 plus.n25 0.189894
R22916 plus.n25 plus.n24 0.189894
R22917 plus.n24 plus.n4 0.189894
R22918 plus.n19 plus.n4 0.189894
R22919 plus.n19 plus.n18 0.189894
R22920 plus.n18 plus.n6 0.189894
R22921 plus.n14 plus.n6 0.189894
R22922 plus.n14 plus.n13 0.189894
R22923 plus.n13 plus.n8 0.189894
R22924 a_n2903_n3924.n0 a_n2903_n3924.t27 214.981
R22925 a_n2903_n3924.n2 a_n2903_n3924.t24 214.452
R22926 a_n2903_n3924.n11 a_n2903_n3924.t36 214.321
R22927 a_n2903_n3924.n12 a_n2903_n3924.t25 214.321
R22928 a_n2903_n3924.n13 a_n2903_n3924.t20 214.321
R22929 a_n2903_n3924.n14 a_n2903_n3924.t37 214.321
R22930 a_n2903_n3924.n15 a_n2903_n3924.t21 214.321
R22931 a_n2903_n3924.n0 a_n2903_n3924.t30 214.321
R22932 a_n2903_n3924.n1 a_n2903_n3924.t15 55.8337
R22933 a_n2903_n3924.n3 a_n2903_n3924.t32 55.8337
R22934 a_n2903_n3924.n10 a_n2903_n3924.t29 55.8337
R22935 a_n2903_n3924.n34 a_n2903_n3924.t12 55.8335
R22936 a_n2903_n3924.n32 a_n2903_n3924.t3 55.8335
R22937 a_n2903_n3924.n25 a_n2903_n3924.t39 55.8335
R22938 a_n2903_n3924.n24 a_n2903_n3924.t13 55.8335
R22939 a_n2903_n3924.n17 a_n2903_n3924.t17 55.8335
R22940 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0052
R22941 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0052
R22942 a_n2903_n3924.n5 a_n2903_n3924.n4 53.0052
R22943 a_n2903_n3924.n7 a_n2903_n3924.n6 53.0052
R22944 a_n2903_n3924.n9 a_n2903_n3924.n8 53.0052
R22945 a_n2903_n3924.n31 a_n2903_n3924.n30 53.0051
R22946 a_n2903_n3924.n29 a_n2903_n3924.n28 53.0051
R22947 a_n2903_n3924.n27 a_n2903_n3924.n26 53.0051
R22948 a_n2903_n3924.n23 a_n2903_n3924.n22 53.0051
R22949 a_n2903_n3924.n21 a_n2903_n3924.n20 53.0051
R22950 a_n2903_n3924.n19 a_n2903_n3924.n18 53.0051
R22951 a_n2903_n3924.n40 a_n2903_n3924.n39 53.0051
R22952 a_n2903_n3924.n16 a_n2903_n3924.n10 12.2417
R22953 a_n2903_n3924.n34 a_n2903_n3924.n33 12.2417
R22954 a_n2903_n3924.n17 a_n2903_n3924.n16 5.16214
R22955 a_n2903_n3924.n33 a_n2903_n3924.n32 5.16214
R22956 a_n2903_n3924.n35 a_n2903_n3924.t10 2.82907
R22957 a_n2903_n3924.n35 a_n2903_n3924.t14 2.82907
R22958 a_n2903_n3924.n37 a_n2903_n3924.t7 2.82907
R22959 a_n2903_n3924.n37 a_n2903_n3924.t11 2.82907
R22960 a_n2903_n3924.n4 a_n2903_n3924.t33 2.82907
R22961 a_n2903_n3924.n4 a_n2903_n3924.t1 2.82907
R22962 a_n2903_n3924.n6 a_n2903_n3924.t34 2.82907
R22963 a_n2903_n3924.n6 a_n2903_n3924.t26 2.82907
R22964 a_n2903_n3924.n8 a_n2903_n3924.t35 2.82907
R22965 a_n2903_n3924.n8 a_n2903_n3924.t2 2.82907
R22966 a_n2903_n3924.n30 a_n2903_n3924.t22 2.82907
R22967 a_n2903_n3924.n30 a_n2903_n3924.t28 2.82907
R22968 a_n2903_n3924.n28 a_n2903_n3924.t31 2.82907
R22969 a_n2903_n3924.n28 a_n2903_n3924.t23 2.82907
R22970 a_n2903_n3924.n26 a_n2903_n3924.t38 2.82907
R22971 a_n2903_n3924.n26 a_n2903_n3924.t0 2.82907
R22972 a_n2903_n3924.n22 a_n2903_n3924.t5 2.82907
R22973 a_n2903_n3924.n22 a_n2903_n3924.t16 2.82907
R22974 a_n2903_n3924.n20 a_n2903_n3924.t9 2.82907
R22975 a_n2903_n3924.n20 a_n2903_n3924.t4 2.82907
R22976 a_n2903_n3924.n18 a_n2903_n3924.t18 2.82907
R22977 a_n2903_n3924.n18 a_n2903_n3924.t8 2.82907
R22978 a_n2903_n3924.t19 a_n2903_n3924.n40 2.82907
R22979 a_n2903_n3924.n40 a_n2903_n3924.t6 2.82907
R22980 a_n2903_n3924.n33 a_n2903_n3924.n2 1.95694
R22981 a_n2903_n3924.n16 a_n2903_n3924.n0 1.95694
R22982 a_n2903_n3924.n0 a_n2903_n3924.n15 0.684366
R22983 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R22984 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R22985 a_n2903_n3924.n13 a_n2903_n3924.n12 0.672012
R22986 a_n2903_n3924.n12 a_n2903_n3924.n11 0.672012
R22987 a_n2903_n3924.n11 a_n2903_n3924.n2 0.541924
R22988 a_n2903_n3924.n19 a_n2903_n3924.n17 0.530672
R22989 a_n2903_n3924.n21 a_n2903_n3924.n19 0.530672
R22990 a_n2903_n3924.n23 a_n2903_n3924.n21 0.530672
R22991 a_n2903_n3924.n24 a_n2903_n3924.n23 0.530672
R22992 a_n2903_n3924.n27 a_n2903_n3924.n25 0.530672
R22993 a_n2903_n3924.n29 a_n2903_n3924.n27 0.530672
R22994 a_n2903_n3924.n31 a_n2903_n3924.n29 0.530672
R22995 a_n2903_n3924.n32 a_n2903_n3924.n31 0.530672
R22996 a_n2903_n3924.n10 a_n2903_n3924.n9 0.530672
R22997 a_n2903_n3924.n9 a_n2903_n3924.n7 0.530672
R22998 a_n2903_n3924.n7 a_n2903_n3924.n5 0.530672
R22999 a_n2903_n3924.n5 a_n2903_n3924.n3 0.530672
R23000 a_n2903_n3924.n39 a_n2903_n3924.n1 0.530672
R23001 a_n2903_n3924.n39 a_n2903_n3924.n38 0.530672
R23002 a_n2903_n3924.n38 a_n2903_n3924.n36 0.530672
R23003 a_n2903_n3924.n36 a_n2903_n3924.n34 0.530672
R23004 a_n2903_n3924.n25 a_n2903_n3924.n24 0.235414
R23005 a_n2903_n3924.n3 a_n2903_n3924.n1 0.235414
R23006 minus.n46 minus.t20 252.611
R23007 minus.n9 minus.t13 252.611
R23008 minus.n78 minus.t3 243.255
R23009 minus.n72 minus.t15 231.093
R23010 minus.n35 minus.t17 231.093
R23011 minus.n77 minus.n75 224.169
R23012 minus.n77 minus.n76 223.454
R23013 minus.n38 minus.t12 187.445
R23014 minus.n65 minus.t7 187.445
R23015 minus.n59 minus.t6 187.445
R23016 minus.n42 minus.t11 187.445
R23017 minus.n44 minus.t10 187.445
R23018 minus.n47 minus.t16 187.445
R23019 minus.n10 minus.t9 187.445
R23020 minus.n7 minus.t8 187.445
R23021 minus.n5 minus.t5 187.445
R23022 minus.n22 minus.t18 187.445
R23023 minus.n28 minus.t19 187.445
R23024 minus.n1 minus.t14 187.445
R23025 minus.n48 minus.n45 161.3
R23026 minus.n50 minus.n49 161.3
R23027 minus.n52 minus.n51 161.3
R23028 minus.n53 minus.n43 161.3
R23029 minus.n55 minus.n54 161.3
R23030 minus.n57 minus.n56 161.3
R23031 minus.n58 minus.n41 161.3
R23032 minus.n61 minus.n60 161.3
R23033 minus.n62 minus.n40 161.3
R23034 minus.n64 minus.n63 161.3
R23035 minus.n66 minus.n39 161.3
R23036 minus.n68 minus.n67 161.3
R23037 minus.n70 minus.n69 161.3
R23038 minus.n71 minus.n37 161.3
R23039 minus.n73 minus.n72 161.3
R23040 minus.n36 minus.n35 161.3
R23041 minus.n34 minus.n0 161.3
R23042 minus.n33 minus.n32 161.3
R23043 minus.n31 minus.n30 161.3
R23044 minus.n29 minus.n2 161.3
R23045 minus.n27 minus.n26 161.3
R23046 minus.n25 minus.n3 161.3
R23047 minus.n24 minus.n23 161.3
R23048 minus.n21 minus.n4 161.3
R23049 minus.n20 minus.n19 161.3
R23050 minus.n18 minus.n17 161.3
R23051 minus.n16 minus.n6 161.3
R23052 minus.n15 minus.n14 161.3
R23053 minus.n13 minus.n12 161.3
R23054 minus.n11 minus.n8 161.3
R23055 minus.n67 minus.n66 56.5617
R23056 minus.n58 minus.n57 56.5617
R23057 minus.n49 minus.n48 56.5617
R23058 minus.n12 minus.n11 56.5617
R23059 minus.n21 minus.n20 56.5617
R23060 minus.n30 minus.n29 56.5617
R23061 minus.n71 minus.n70 46.3896
R23062 minus.n34 minus.n33 46.3896
R23063 minus.n46 minus.n45 42.8164
R23064 minus.n9 minus.n8 42.8164
R23065 minus.n60 minus.n40 42.5146
R23066 minus.n54 minus.n53 42.5146
R23067 minus.n17 minus.n16 42.5146
R23068 minus.n23 minus.n3 42.5146
R23069 minus.n64 minus.n40 38.6395
R23070 minus.n53 minus.n52 38.6395
R23071 minus.n16 minus.n15 38.6395
R23072 minus.n27 minus.n3 38.6395
R23073 minus.n47 minus.n46 38.2514
R23074 minus.n10 minus.n9 38.2514
R23075 minus.n74 minus.n73 31.7069
R23076 minus.n66 minus.n65 19.9199
R23077 minus.n49 minus.n44 19.9199
R23078 minus.n12 minus.n7 19.9199
R23079 minus.n29 minus.n28 19.9199
R23080 minus.n76 minus.t2 19.8005
R23081 minus.n76 minus.t0 19.8005
R23082 minus.n75 minus.t1 19.8005
R23083 minus.n75 minus.t4 19.8005
R23084 minus.n59 minus.n58 17.9525
R23085 minus.n57 minus.n42 17.9525
R23086 minus.n20 minus.n5 17.9525
R23087 minus.n22 minus.n21 17.9525
R23088 minus.n67 minus.n38 15.9852
R23089 minus.n48 minus.n47 15.9852
R23090 minus.n11 minus.n10 15.9852
R23091 minus.n30 minus.n1 15.9852
R23092 minus.n72 minus.n71 15.3369
R23093 minus.n35 minus.n34 15.3369
R23094 minus.n74 minus.n36 12.1653
R23095 minus minus.n79 11.4284
R23096 minus.n70 minus.n38 8.60764
R23097 minus.n33 minus.n1 8.60764
R23098 minus.n60 minus.n59 6.6403
R23099 minus.n54 minus.n42 6.6403
R23100 minus.n17 minus.n5 6.6403
R23101 minus.n23 minus.n22 6.6403
R23102 minus.n79 minus.n78 4.80222
R23103 minus.n65 minus.n64 4.67295
R23104 minus.n52 minus.n44 4.67295
R23105 minus.n15 minus.n7 4.67295
R23106 minus.n28 minus.n27 4.67295
R23107 minus.n79 minus.n74 0.972091
R23108 minus.n78 minus.n77 0.716017
R23109 minus.n73 minus.n37 0.189894
R23110 minus.n69 minus.n37 0.189894
R23111 minus.n69 minus.n68 0.189894
R23112 minus.n68 minus.n39 0.189894
R23113 minus.n63 minus.n39 0.189894
R23114 minus.n63 minus.n62 0.189894
R23115 minus.n62 minus.n61 0.189894
R23116 minus.n61 minus.n41 0.189894
R23117 minus.n56 minus.n41 0.189894
R23118 minus.n56 minus.n55 0.189894
R23119 minus.n55 minus.n43 0.189894
R23120 minus.n51 minus.n43 0.189894
R23121 minus.n51 minus.n50 0.189894
R23122 minus.n50 minus.n45 0.189894
R23123 minus.n13 minus.n8 0.189894
R23124 minus.n14 minus.n13 0.189894
R23125 minus.n14 minus.n6 0.189894
R23126 minus.n18 minus.n6 0.189894
R23127 minus.n19 minus.n18 0.189894
R23128 minus.n19 minus.n4 0.189894
R23129 minus.n24 minus.n4 0.189894
R23130 minus.n25 minus.n24 0.189894
R23131 minus.n26 minus.n25 0.189894
R23132 minus.n26 minus.n2 0.189894
R23133 minus.n31 minus.n2 0.189894
R23134 minus.n32 minus.n31 0.189894
R23135 minus.n32 minus.n0 0.189894
R23136 minus.n36 minus.n0 0.189894
R23137 a_n2650_8322.n10 a_n2650_8322.t3 74.6477
R23138 a_n2650_8322.n1 a_n2650_8322.t23 74.6477
R23139 a_n2650_8322.n24 a_n2650_8322.t25 74.6474
R23140 a_n2650_8322.n18 a_n2650_8322.t22 74.2899
R23141 a_n2650_8322.n11 a_n2650_8322.t1 74.2899
R23142 a_n2650_8322.n12 a_n2650_8322.t4 74.2899
R23143 a_n2650_8322.n15 a_n2650_8322.t5 74.2899
R23144 a_n2650_8322.n8 a_n2650_8322.t8 74.2899
R23145 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R23146 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R23147 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R23148 a_n2650_8322.n10 a_n2650_8322.n9 70.6783
R23149 a_n2650_8322.n14 a_n2650_8322.n13 70.6783
R23150 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R23151 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R23152 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R23153 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R23154 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R23155 a_n2650_8322.n16 a_n2650_8322.n8 24.1867
R23156 a_n2650_8322.n17 a_n2650_8322.t29 9.69192
R23157 a_n2650_8322.n16 a_n2650_8322.n15 7.67184
R23158 a_n2650_8322.n18 a_n2650_8322.n17 6.55222
R23159 a_n2650_8322.n17 a_n2650_8322.n16 5.3452
R23160 a_n2650_8322.n23 a_n2650_8322.t20 3.61217
R23161 a_n2650_8322.n23 a_n2650_8322.t16 3.61217
R23162 a_n2650_8322.n21 a_n2650_8322.t24 3.61217
R23163 a_n2650_8322.n21 a_n2650_8322.t14 3.61217
R23164 a_n2650_8322.n19 a_n2650_8322.t12 3.61217
R23165 a_n2650_8322.n19 a_n2650_8322.t11 3.61217
R23166 a_n2650_8322.n9 a_n2650_8322.t7 3.61217
R23167 a_n2650_8322.n9 a_n2650_8322.t6 3.61217
R23168 a_n2650_8322.n13 a_n2650_8322.t2 3.61217
R23169 a_n2650_8322.n13 a_n2650_8322.t0 3.61217
R23170 a_n2650_8322.n0 a_n2650_8322.t26 3.61217
R23171 a_n2650_8322.n0 a_n2650_8322.t18 3.61217
R23172 a_n2650_8322.n2 a_n2650_8322.t10 3.61217
R23173 a_n2650_8322.n2 a_n2650_8322.t9 3.61217
R23174 a_n2650_8322.n4 a_n2650_8322.t21 3.61217
R23175 a_n2650_8322.n4 a_n2650_8322.t15 3.61217
R23176 a_n2650_8322.n6 a_n2650_8322.t19 3.61217
R23177 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R23178 a_n2650_8322.n26 a_n2650_8322.t13 3.61217
R23179 a_n2650_8322.t27 a_n2650_8322.n26 3.61217
R23180 a_n2650_8322.n15 a_n2650_8322.n14 0.358259
R23181 a_n2650_8322.n14 a_n2650_8322.n12 0.358259
R23182 a_n2650_8322.n11 a_n2650_8322.n10 0.358259
R23183 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R23184 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R23185 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R23186 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R23187 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R23188 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R23189 a_n2650_8322.n25 a_n2650_8322.n22 0.358259
R23190 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R23191 a_n2650_8322.n12 a_n2650_8322.n11 0.101793
R23192 a_n2650_8322.t33 a_n2650_8322.t31 0.0788333
R23193 a_n2650_8322.t30 a_n2650_8322.t32 0.0788333
R23194 a_n2650_8322.t29 a_n2650_8322.t28 0.0788333
R23195 a_n2650_8322.t30 a_n2650_8322.t33 0.0318333
R23196 a_n2650_8322.t29 a_n2650_8322.t32 0.0318333
R23197 a_n2650_8322.t31 a_n2650_8322.t32 0.0318333
R23198 a_n2650_8322.t28 a_n2650_8322.t30 0.0318333
R23199 diffpairibias.n0 diffpairibias.t18 436.822
R23200 diffpairibias.n21 diffpairibias.t19 435.479
R23201 diffpairibias.n20 diffpairibias.t16 435.479
R23202 diffpairibias.n19 diffpairibias.t17 435.479
R23203 diffpairibias.n18 diffpairibias.t21 435.479
R23204 diffpairibias.n0 diffpairibias.t22 435.479
R23205 diffpairibias.n1 diffpairibias.t20 435.479
R23206 diffpairibias.n2 diffpairibias.t23 435.479
R23207 diffpairibias.n10 diffpairibias.t0 377.536
R23208 diffpairibias.n10 diffpairibias.t8 376.193
R23209 diffpairibias.n11 diffpairibias.t10 376.193
R23210 diffpairibias.n12 diffpairibias.t6 376.193
R23211 diffpairibias.n13 diffpairibias.t2 376.193
R23212 diffpairibias.n14 diffpairibias.t12 376.193
R23213 diffpairibias.n15 diffpairibias.t4 376.193
R23214 diffpairibias.n16 diffpairibias.t14 376.193
R23215 diffpairibias.n3 diffpairibias.t1 113.368
R23216 diffpairibias.n3 diffpairibias.t9 112.698
R23217 diffpairibias.n4 diffpairibias.t11 112.698
R23218 diffpairibias.n5 diffpairibias.t7 112.698
R23219 diffpairibias.n6 diffpairibias.t3 112.698
R23220 diffpairibias.n7 diffpairibias.t13 112.698
R23221 diffpairibias.n8 diffpairibias.t5 112.698
R23222 diffpairibias.n9 diffpairibias.t15 112.698
R23223 diffpairibias.n17 diffpairibias.n16 4.77242
R23224 diffpairibias.n17 diffpairibias.n9 4.30807
R23225 diffpairibias.n18 diffpairibias.n17 4.13945
R23226 diffpairibias.n16 diffpairibias.n15 1.34352
R23227 diffpairibias.n15 diffpairibias.n14 1.34352
R23228 diffpairibias.n14 diffpairibias.n13 1.34352
R23229 diffpairibias.n13 diffpairibias.n12 1.34352
R23230 diffpairibias.n12 diffpairibias.n11 1.34352
R23231 diffpairibias.n11 diffpairibias.n10 1.34352
R23232 diffpairibias.n2 diffpairibias.n1 1.34352
R23233 diffpairibias.n1 diffpairibias.n0 1.34352
R23234 diffpairibias.n19 diffpairibias.n18 1.34352
R23235 diffpairibias.n20 diffpairibias.n19 1.34352
R23236 diffpairibias.n21 diffpairibias.n20 1.34352
R23237 diffpairibias.n22 diffpairibias.n21 0.862419
R23238 diffpairibias diffpairibias.n22 0.684875
R23239 diffpairibias.n9 diffpairibias.n8 0.672012
R23240 diffpairibias.n8 diffpairibias.n7 0.672012
R23241 diffpairibias.n7 diffpairibias.n6 0.672012
R23242 diffpairibias.n6 diffpairibias.n5 0.672012
R23243 diffpairibias.n5 diffpairibias.n4 0.672012
R23244 diffpairibias.n4 diffpairibias.n3 0.672012
R23245 diffpairibias.n22 diffpairibias.n2 0.190907
R23246 outputibias.n27 outputibias.n1 289.615
R23247 outputibias.n58 outputibias.n32 289.615
R23248 outputibias.n90 outputibias.n64 289.615
R23249 outputibias.n122 outputibias.n96 289.615
R23250 outputibias.n28 outputibias.n27 185
R23251 outputibias.n26 outputibias.n25 185
R23252 outputibias.n5 outputibias.n4 185
R23253 outputibias.n20 outputibias.n19 185
R23254 outputibias.n18 outputibias.n17 185
R23255 outputibias.n9 outputibias.n8 185
R23256 outputibias.n12 outputibias.n11 185
R23257 outputibias.n59 outputibias.n58 185
R23258 outputibias.n57 outputibias.n56 185
R23259 outputibias.n36 outputibias.n35 185
R23260 outputibias.n51 outputibias.n50 185
R23261 outputibias.n49 outputibias.n48 185
R23262 outputibias.n40 outputibias.n39 185
R23263 outputibias.n43 outputibias.n42 185
R23264 outputibias.n91 outputibias.n90 185
R23265 outputibias.n89 outputibias.n88 185
R23266 outputibias.n68 outputibias.n67 185
R23267 outputibias.n83 outputibias.n82 185
R23268 outputibias.n81 outputibias.n80 185
R23269 outputibias.n72 outputibias.n71 185
R23270 outputibias.n75 outputibias.n74 185
R23271 outputibias.n123 outputibias.n122 185
R23272 outputibias.n121 outputibias.n120 185
R23273 outputibias.n100 outputibias.n99 185
R23274 outputibias.n115 outputibias.n114 185
R23275 outputibias.n113 outputibias.n112 185
R23276 outputibias.n104 outputibias.n103 185
R23277 outputibias.n107 outputibias.n106 185
R23278 outputibias.n0 outputibias.t8 178.945
R23279 outputibias.n133 outputibias.t11 177.018
R23280 outputibias.n132 outputibias.t9 177.018
R23281 outputibias.n0 outputibias.t10 177.018
R23282 outputibias.t1 outputibias.n10 147.661
R23283 outputibias.t3 outputibias.n41 147.661
R23284 outputibias.t5 outputibias.n73 147.661
R23285 outputibias.t7 outputibias.n105 147.661
R23286 outputibias.n128 outputibias.t0 132.363
R23287 outputibias.n128 outputibias.t2 130.436
R23288 outputibias.n129 outputibias.t4 130.436
R23289 outputibias.n130 outputibias.t6 130.436
R23290 outputibias.n27 outputibias.n26 104.615
R23291 outputibias.n26 outputibias.n4 104.615
R23292 outputibias.n19 outputibias.n4 104.615
R23293 outputibias.n19 outputibias.n18 104.615
R23294 outputibias.n18 outputibias.n8 104.615
R23295 outputibias.n11 outputibias.n8 104.615
R23296 outputibias.n58 outputibias.n57 104.615
R23297 outputibias.n57 outputibias.n35 104.615
R23298 outputibias.n50 outputibias.n35 104.615
R23299 outputibias.n50 outputibias.n49 104.615
R23300 outputibias.n49 outputibias.n39 104.615
R23301 outputibias.n42 outputibias.n39 104.615
R23302 outputibias.n90 outputibias.n89 104.615
R23303 outputibias.n89 outputibias.n67 104.615
R23304 outputibias.n82 outputibias.n67 104.615
R23305 outputibias.n82 outputibias.n81 104.615
R23306 outputibias.n81 outputibias.n71 104.615
R23307 outputibias.n74 outputibias.n71 104.615
R23308 outputibias.n122 outputibias.n121 104.615
R23309 outputibias.n121 outputibias.n99 104.615
R23310 outputibias.n114 outputibias.n99 104.615
R23311 outputibias.n114 outputibias.n113 104.615
R23312 outputibias.n113 outputibias.n103 104.615
R23313 outputibias.n106 outputibias.n103 104.615
R23314 outputibias.n63 outputibias.n31 95.6354
R23315 outputibias.n63 outputibias.n62 94.6732
R23316 outputibias.n95 outputibias.n94 94.6732
R23317 outputibias.n127 outputibias.n126 94.6732
R23318 outputibias.n11 outputibias.t1 52.3082
R23319 outputibias.n42 outputibias.t3 52.3082
R23320 outputibias.n74 outputibias.t5 52.3082
R23321 outputibias.n106 outputibias.t7 52.3082
R23322 outputibias.n12 outputibias.n10 15.6674
R23323 outputibias.n43 outputibias.n41 15.6674
R23324 outputibias.n75 outputibias.n73 15.6674
R23325 outputibias.n107 outputibias.n105 15.6674
R23326 outputibias.n13 outputibias.n9 12.8005
R23327 outputibias.n44 outputibias.n40 12.8005
R23328 outputibias.n76 outputibias.n72 12.8005
R23329 outputibias.n108 outputibias.n104 12.8005
R23330 outputibias.n17 outputibias.n16 12.0247
R23331 outputibias.n48 outputibias.n47 12.0247
R23332 outputibias.n80 outputibias.n79 12.0247
R23333 outputibias.n112 outputibias.n111 12.0247
R23334 outputibias.n20 outputibias.n7 11.249
R23335 outputibias.n51 outputibias.n38 11.249
R23336 outputibias.n83 outputibias.n70 11.249
R23337 outputibias.n115 outputibias.n102 11.249
R23338 outputibias.n21 outputibias.n5 10.4732
R23339 outputibias.n52 outputibias.n36 10.4732
R23340 outputibias.n84 outputibias.n68 10.4732
R23341 outputibias.n116 outputibias.n100 10.4732
R23342 outputibias.n25 outputibias.n24 9.69747
R23343 outputibias.n56 outputibias.n55 9.69747
R23344 outputibias.n88 outputibias.n87 9.69747
R23345 outputibias.n120 outputibias.n119 9.69747
R23346 outputibias.n31 outputibias.n30 9.45567
R23347 outputibias.n62 outputibias.n61 9.45567
R23348 outputibias.n94 outputibias.n93 9.45567
R23349 outputibias.n126 outputibias.n125 9.45567
R23350 outputibias.n30 outputibias.n29 9.3005
R23351 outputibias.n3 outputibias.n2 9.3005
R23352 outputibias.n24 outputibias.n23 9.3005
R23353 outputibias.n22 outputibias.n21 9.3005
R23354 outputibias.n7 outputibias.n6 9.3005
R23355 outputibias.n16 outputibias.n15 9.3005
R23356 outputibias.n14 outputibias.n13 9.3005
R23357 outputibias.n61 outputibias.n60 9.3005
R23358 outputibias.n34 outputibias.n33 9.3005
R23359 outputibias.n55 outputibias.n54 9.3005
R23360 outputibias.n53 outputibias.n52 9.3005
R23361 outputibias.n38 outputibias.n37 9.3005
R23362 outputibias.n47 outputibias.n46 9.3005
R23363 outputibias.n45 outputibias.n44 9.3005
R23364 outputibias.n93 outputibias.n92 9.3005
R23365 outputibias.n66 outputibias.n65 9.3005
R23366 outputibias.n87 outputibias.n86 9.3005
R23367 outputibias.n85 outputibias.n84 9.3005
R23368 outputibias.n70 outputibias.n69 9.3005
R23369 outputibias.n79 outputibias.n78 9.3005
R23370 outputibias.n77 outputibias.n76 9.3005
R23371 outputibias.n125 outputibias.n124 9.3005
R23372 outputibias.n98 outputibias.n97 9.3005
R23373 outputibias.n119 outputibias.n118 9.3005
R23374 outputibias.n117 outputibias.n116 9.3005
R23375 outputibias.n102 outputibias.n101 9.3005
R23376 outputibias.n111 outputibias.n110 9.3005
R23377 outputibias.n109 outputibias.n108 9.3005
R23378 outputibias.n28 outputibias.n3 8.92171
R23379 outputibias.n59 outputibias.n34 8.92171
R23380 outputibias.n91 outputibias.n66 8.92171
R23381 outputibias.n123 outputibias.n98 8.92171
R23382 outputibias.n29 outputibias.n1 8.14595
R23383 outputibias.n60 outputibias.n32 8.14595
R23384 outputibias.n92 outputibias.n64 8.14595
R23385 outputibias.n124 outputibias.n96 8.14595
R23386 outputibias.n31 outputibias.n1 5.81868
R23387 outputibias.n62 outputibias.n32 5.81868
R23388 outputibias.n94 outputibias.n64 5.81868
R23389 outputibias.n126 outputibias.n96 5.81868
R23390 outputibias.n131 outputibias.n130 5.20947
R23391 outputibias.n29 outputibias.n28 5.04292
R23392 outputibias.n60 outputibias.n59 5.04292
R23393 outputibias.n92 outputibias.n91 5.04292
R23394 outputibias.n124 outputibias.n123 5.04292
R23395 outputibias.n131 outputibias.n127 4.42209
R23396 outputibias.n14 outputibias.n10 4.38594
R23397 outputibias.n45 outputibias.n41 4.38594
R23398 outputibias.n77 outputibias.n73 4.38594
R23399 outputibias.n109 outputibias.n105 4.38594
R23400 outputibias.n132 outputibias.n131 4.28454
R23401 outputibias.n25 outputibias.n3 4.26717
R23402 outputibias.n56 outputibias.n34 4.26717
R23403 outputibias.n88 outputibias.n66 4.26717
R23404 outputibias.n120 outputibias.n98 4.26717
R23405 outputibias.n24 outputibias.n5 3.49141
R23406 outputibias.n55 outputibias.n36 3.49141
R23407 outputibias.n87 outputibias.n68 3.49141
R23408 outputibias.n119 outputibias.n100 3.49141
R23409 outputibias.n21 outputibias.n20 2.71565
R23410 outputibias.n52 outputibias.n51 2.71565
R23411 outputibias.n84 outputibias.n83 2.71565
R23412 outputibias.n116 outputibias.n115 2.71565
R23413 outputibias.n17 outputibias.n7 1.93989
R23414 outputibias.n48 outputibias.n38 1.93989
R23415 outputibias.n80 outputibias.n70 1.93989
R23416 outputibias.n112 outputibias.n102 1.93989
R23417 outputibias.n130 outputibias.n129 1.9266
R23418 outputibias.n129 outputibias.n128 1.9266
R23419 outputibias.n133 outputibias.n132 1.92658
R23420 outputibias.n134 outputibias.n133 1.29913
R23421 outputibias.n16 outputibias.n9 1.16414
R23422 outputibias.n47 outputibias.n40 1.16414
R23423 outputibias.n79 outputibias.n72 1.16414
R23424 outputibias.n111 outputibias.n104 1.16414
R23425 outputibias.n127 outputibias.n95 0.962709
R23426 outputibias.n95 outputibias.n63 0.962709
R23427 outputibias.n13 outputibias.n12 0.388379
R23428 outputibias.n44 outputibias.n43 0.388379
R23429 outputibias.n76 outputibias.n75 0.388379
R23430 outputibias.n108 outputibias.n107 0.388379
R23431 outputibias.n134 outputibias.n0 0.337251
R23432 outputibias outputibias.n134 0.302375
R23433 outputibias.n30 outputibias.n2 0.155672
R23434 outputibias.n23 outputibias.n2 0.155672
R23435 outputibias.n23 outputibias.n22 0.155672
R23436 outputibias.n22 outputibias.n6 0.155672
R23437 outputibias.n15 outputibias.n6 0.155672
R23438 outputibias.n15 outputibias.n14 0.155672
R23439 outputibias.n61 outputibias.n33 0.155672
R23440 outputibias.n54 outputibias.n33 0.155672
R23441 outputibias.n54 outputibias.n53 0.155672
R23442 outputibias.n53 outputibias.n37 0.155672
R23443 outputibias.n46 outputibias.n37 0.155672
R23444 outputibias.n46 outputibias.n45 0.155672
R23445 outputibias.n93 outputibias.n65 0.155672
R23446 outputibias.n86 outputibias.n65 0.155672
R23447 outputibias.n86 outputibias.n85 0.155672
R23448 outputibias.n85 outputibias.n69 0.155672
R23449 outputibias.n78 outputibias.n69 0.155672
R23450 outputibias.n78 outputibias.n77 0.155672
R23451 outputibias.n125 outputibias.n97 0.155672
R23452 outputibias.n118 outputibias.n97 0.155672
R23453 outputibias.n118 outputibias.n117 0.155672
R23454 outputibias.n117 outputibias.n101 0.155672
R23455 outputibias.n110 outputibias.n101 0.155672
R23456 outputibias.n110 outputibias.n109 0.155672
C0 CSoutput minus 2.67006f
C1 vdd plus 0.096826f
C2 commonsourceibias outputibias 0.003761f
C3 plus diffpairibias 2.47e-19
C4 vdd commonsourceibias 0.004173f
C5 CSoutput plus 0.849267f
C6 commonsourceibias diffpairibias 0.06482f
C7 CSoutput commonsourceibias 41.993103f
C8 minus plus 9.025571f
C9 minus commonsourceibias 0.323289f
C10 plus commonsourceibias 0.277692f
C11 output outputibias 2.34152f
C12 vdd output 7.23429f
C13 CSoutput output 6.13881f
C14 CSoutput outputibias 0.032386f
C15 vdd CSoutput 0.142056p
C16 minus diffpairibias 3.46e-19
C17 commonsourceibias output 0.006787f
C18 diffpairibias gnd 48.980137f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.144689p
C22 plus gnd 32.34897f
C23 minus gnd 26.507359f
C24 CSoutput gnd 0.106601p
C25 vdd gnd 0.507681p
C26 outputibias.t10 gnd 0.11477f
C27 outputibias.t8 gnd 0.115567f
C28 outputibias.n0 gnd 0.130108f
C29 outputibias.n1 gnd 0.001372f
C30 outputibias.n2 gnd 9.76e-19
C31 outputibias.n3 gnd 5.24e-19
C32 outputibias.n4 gnd 0.001239f
C33 outputibias.n5 gnd 5.55e-19
C34 outputibias.n6 gnd 9.76e-19
C35 outputibias.n7 gnd 5.24e-19
C36 outputibias.n8 gnd 0.001239f
C37 outputibias.n9 gnd 5.55e-19
C38 outputibias.n10 gnd 0.004176f
C39 outputibias.t1 gnd 0.00202f
C40 outputibias.n11 gnd 9.3e-19
C41 outputibias.n12 gnd 7.32e-19
C42 outputibias.n13 gnd 5.24e-19
C43 outputibias.n14 gnd 0.02322f
C44 outputibias.n15 gnd 9.76e-19
C45 outputibias.n16 gnd 5.24e-19
C46 outputibias.n17 gnd 5.55e-19
C47 outputibias.n18 gnd 0.001239f
C48 outputibias.n19 gnd 0.001239f
C49 outputibias.n20 gnd 5.55e-19
C50 outputibias.n21 gnd 5.24e-19
C51 outputibias.n22 gnd 9.76e-19
C52 outputibias.n23 gnd 9.76e-19
C53 outputibias.n24 gnd 5.24e-19
C54 outputibias.n25 gnd 5.55e-19
C55 outputibias.n26 gnd 0.001239f
C56 outputibias.n27 gnd 0.002683f
C57 outputibias.n28 gnd 5.55e-19
C58 outputibias.n29 gnd 5.24e-19
C59 outputibias.n30 gnd 0.002256f
C60 outputibias.n31 gnd 0.005781f
C61 outputibias.n32 gnd 0.001372f
C62 outputibias.n33 gnd 9.76e-19
C63 outputibias.n34 gnd 5.24e-19
C64 outputibias.n35 gnd 0.001239f
C65 outputibias.n36 gnd 5.55e-19
C66 outputibias.n37 gnd 9.76e-19
C67 outputibias.n38 gnd 5.24e-19
C68 outputibias.n39 gnd 0.001239f
C69 outputibias.n40 gnd 5.55e-19
C70 outputibias.n41 gnd 0.004176f
C71 outputibias.t3 gnd 0.00202f
C72 outputibias.n42 gnd 9.3e-19
C73 outputibias.n43 gnd 7.32e-19
C74 outputibias.n44 gnd 5.24e-19
C75 outputibias.n45 gnd 0.02322f
C76 outputibias.n46 gnd 9.76e-19
C77 outputibias.n47 gnd 5.24e-19
C78 outputibias.n48 gnd 5.55e-19
C79 outputibias.n49 gnd 0.001239f
C80 outputibias.n50 gnd 0.001239f
C81 outputibias.n51 gnd 5.55e-19
C82 outputibias.n52 gnd 5.24e-19
C83 outputibias.n53 gnd 9.76e-19
C84 outputibias.n54 gnd 9.76e-19
C85 outputibias.n55 gnd 5.24e-19
C86 outputibias.n56 gnd 5.55e-19
C87 outputibias.n57 gnd 0.001239f
C88 outputibias.n58 gnd 0.002683f
C89 outputibias.n59 gnd 5.55e-19
C90 outputibias.n60 gnd 5.24e-19
C91 outputibias.n61 gnd 0.002256f
C92 outputibias.n62 gnd 0.005197f
C93 outputibias.n63 gnd 0.121892f
C94 outputibias.n64 gnd 0.001372f
C95 outputibias.n65 gnd 9.76e-19
C96 outputibias.n66 gnd 5.24e-19
C97 outputibias.n67 gnd 0.001239f
C98 outputibias.n68 gnd 5.55e-19
C99 outputibias.n69 gnd 9.76e-19
C100 outputibias.n70 gnd 5.24e-19
C101 outputibias.n71 gnd 0.001239f
C102 outputibias.n72 gnd 5.55e-19
C103 outputibias.n73 gnd 0.004176f
C104 outputibias.t5 gnd 0.00202f
C105 outputibias.n74 gnd 9.3e-19
C106 outputibias.n75 gnd 7.32e-19
C107 outputibias.n76 gnd 5.24e-19
C108 outputibias.n77 gnd 0.02322f
C109 outputibias.n78 gnd 9.76e-19
C110 outputibias.n79 gnd 5.24e-19
C111 outputibias.n80 gnd 5.55e-19
C112 outputibias.n81 gnd 0.001239f
C113 outputibias.n82 gnd 0.001239f
C114 outputibias.n83 gnd 5.55e-19
C115 outputibias.n84 gnd 5.24e-19
C116 outputibias.n85 gnd 9.76e-19
C117 outputibias.n86 gnd 9.76e-19
C118 outputibias.n87 gnd 5.24e-19
C119 outputibias.n88 gnd 5.55e-19
C120 outputibias.n89 gnd 0.001239f
C121 outputibias.n90 gnd 0.002683f
C122 outputibias.n91 gnd 5.55e-19
C123 outputibias.n92 gnd 5.24e-19
C124 outputibias.n93 gnd 0.002256f
C125 outputibias.n94 gnd 0.005197f
C126 outputibias.n95 gnd 0.064513f
C127 outputibias.n96 gnd 0.001372f
C128 outputibias.n97 gnd 9.76e-19
C129 outputibias.n98 gnd 5.24e-19
C130 outputibias.n99 gnd 0.001239f
C131 outputibias.n100 gnd 5.55e-19
C132 outputibias.n101 gnd 9.76e-19
C133 outputibias.n102 gnd 5.24e-19
C134 outputibias.n103 gnd 0.001239f
C135 outputibias.n104 gnd 5.55e-19
C136 outputibias.n105 gnd 0.004176f
C137 outputibias.t7 gnd 0.00202f
C138 outputibias.n106 gnd 9.3e-19
C139 outputibias.n107 gnd 7.32e-19
C140 outputibias.n108 gnd 5.24e-19
C141 outputibias.n109 gnd 0.02322f
C142 outputibias.n110 gnd 9.76e-19
C143 outputibias.n111 gnd 5.24e-19
C144 outputibias.n112 gnd 5.55e-19
C145 outputibias.n113 gnd 0.001239f
C146 outputibias.n114 gnd 0.001239f
C147 outputibias.n115 gnd 5.55e-19
C148 outputibias.n116 gnd 5.24e-19
C149 outputibias.n117 gnd 9.76e-19
C150 outputibias.n118 gnd 9.76e-19
C151 outputibias.n119 gnd 5.24e-19
C152 outputibias.n120 gnd 5.55e-19
C153 outputibias.n121 gnd 0.001239f
C154 outputibias.n122 gnd 0.002683f
C155 outputibias.n123 gnd 5.55e-19
C156 outputibias.n124 gnd 5.24e-19
C157 outputibias.n125 gnd 0.002256f
C158 outputibias.n126 gnd 0.005197f
C159 outputibias.n127 gnd 0.084814f
C160 outputibias.t6 gnd 0.108319f
C161 outputibias.t4 gnd 0.108319f
C162 outputibias.t2 gnd 0.108319f
C163 outputibias.t0 gnd 0.109238f
C164 outputibias.n128 gnd 0.134674f
C165 outputibias.n129 gnd 0.07244f
C166 outputibias.n130 gnd 0.079818f
C167 outputibias.n131 gnd 0.164901f
C168 outputibias.t9 gnd 0.11477f
C169 outputibias.n132 gnd 0.067481f
C170 outputibias.t11 gnd 0.11477f
C171 outputibias.n133 gnd 0.065115f
C172 outputibias.n134 gnd 0.029159f
C173 diffpairibias.t18 gnd 0.087401f
C174 diffpairibias.t22 gnd 0.087239f
C175 diffpairibias.n0 gnd 0.102784f
C176 diffpairibias.t20 gnd 0.087239f
C177 diffpairibias.n1 gnd 0.050171f
C178 diffpairibias.t23 gnd 0.087239f
C179 diffpairibias.n2 gnd 0.039841f
C180 diffpairibias.t1 gnd 0.083757f
C181 diffpairibias.t9 gnd 0.083392f
C182 diffpairibias.n3 gnd 0.131682f
C183 diffpairibias.t11 gnd 0.083392f
C184 diffpairibias.n4 gnd 0.07027f
C185 diffpairibias.t7 gnd 0.083392f
C186 diffpairibias.n5 gnd 0.07027f
C187 diffpairibias.t3 gnd 0.083392f
C188 diffpairibias.n6 gnd 0.07027f
C189 diffpairibias.t13 gnd 0.083392f
C190 diffpairibias.n7 gnd 0.07027f
C191 diffpairibias.t5 gnd 0.083392f
C192 diffpairibias.n8 gnd 0.07027f
C193 diffpairibias.t15 gnd 0.083392f
C194 diffpairibias.n9 gnd 0.099771f
C195 diffpairibias.t0 gnd 0.08427f
C196 diffpairibias.t8 gnd 0.084123f
C197 diffpairibias.n10 gnd 0.091784f
C198 diffpairibias.t10 gnd 0.084123f
C199 diffpairibias.n11 gnd 0.050681f
C200 diffpairibias.t6 gnd 0.084123f
C201 diffpairibias.n12 gnd 0.050681f
C202 diffpairibias.t2 gnd 0.084123f
C203 diffpairibias.n13 gnd 0.050681f
C204 diffpairibias.t12 gnd 0.084123f
C205 diffpairibias.n14 gnd 0.050681f
C206 diffpairibias.t4 gnd 0.084123f
C207 diffpairibias.n15 gnd 0.050681f
C208 diffpairibias.t14 gnd 0.084123f
C209 diffpairibias.n16 gnd 0.059977f
C210 diffpairibias.n17 gnd 0.226448f
C211 diffpairibias.t21 gnd 0.087239f
C212 diffpairibias.n18 gnd 0.050181f
C213 diffpairibias.t17 gnd 0.087239f
C214 diffpairibias.n19 gnd 0.050171f
C215 diffpairibias.t16 gnd 0.087239f
C216 diffpairibias.n20 gnd 0.050171f
C217 diffpairibias.t19 gnd 0.087239f
C218 diffpairibias.n21 gnd 0.045859f
C219 diffpairibias.n22 gnd 0.046268f
C220 a_n2650_8322.t13 gnd 0.098066f
C221 a_n2650_8322.t32 gnd 20.3446f
C222 a_n2650_8322.t31 gnd 20.202f
C223 a_n2650_8322.t33 gnd 20.202f
C224 a_n2650_8322.t30 gnd 20.3446f
C225 a_n2650_8322.t28 gnd 20.202f
C226 a_n2650_8322.t29 gnd 28.365099f
C227 a_n2650_8322.t23 gnd 0.918238f
C228 a_n2650_8322.t26 gnd 0.098066f
C229 a_n2650_8322.t18 gnd 0.098066f
C230 a_n2650_8322.n0 gnd 0.690775f
C231 a_n2650_8322.n1 gnd 0.771839f
C232 a_n2650_8322.t10 gnd 0.098066f
C233 a_n2650_8322.t9 gnd 0.098066f
C234 a_n2650_8322.n2 gnd 0.690775f
C235 a_n2650_8322.n3 gnd 0.392162f
C236 a_n2650_8322.t21 gnd 0.098066f
C237 a_n2650_8322.t15 gnd 0.098066f
C238 a_n2650_8322.n4 gnd 0.690775f
C239 a_n2650_8322.n5 gnd 0.392162f
C240 a_n2650_8322.t19 gnd 0.098066f
C241 a_n2650_8322.t17 gnd 0.098066f
C242 a_n2650_8322.n6 gnd 0.690775f
C243 a_n2650_8322.n7 gnd 0.392162f
C244 a_n2650_8322.t8 gnd 0.916409f
C245 a_n2650_8322.n8 gnd 1.71012f
C246 a_n2650_8322.t3 gnd 0.918238f
C247 a_n2650_8322.t7 gnd 0.098066f
C248 a_n2650_8322.t6 gnd 0.098066f
C249 a_n2650_8322.n9 gnd 0.690775f
C250 a_n2650_8322.n10 gnd 0.771839f
C251 a_n2650_8322.t1 gnd 0.916409f
C252 a_n2650_8322.n11 gnd 0.3884f
C253 a_n2650_8322.t4 gnd 0.916409f
C254 a_n2650_8322.n12 gnd 0.3884f
C255 a_n2650_8322.t2 gnd 0.098066f
C256 a_n2650_8322.t0 gnd 0.098066f
C257 a_n2650_8322.n13 gnd 0.690775f
C258 a_n2650_8322.n14 gnd 0.392162f
C259 a_n2650_8322.t5 gnd 0.916409f
C260 a_n2650_8322.n15 gnd 1.27428f
C261 a_n2650_8322.n16 gnd 2.08205f
C262 a_n2650_8322.n17 gnd 3.23313f
C263 a_n2650_8322.t22 gnd 0.916409f
C264 a_n2650_8322.n18 gnd 0.996789f
C265 a_n2650_8322.t12 gnd 0.098066f
C266 a_n2650_8322.t11 gnd 0.098066f
C267 a_n2650_8322.n19 gnd 0.690775f
C268 a_n2650_8322.n20 gnd 0.392162f
C269 a_n2650_8322.t24 gnd 0.098066f
C270 a_n2650_8322.t14 gnd 0.098066f
C271 a_n2650_8322.n21 gnd 0.690775f
C272 a_n2650_8322.n22 gnd 0.392162f
C273 a_n2650_8322.t25 gnd 0.918235f
C274 a_n2650_8322.t20 gnd 0.098066f
C275 a_n2650_8322.t16 gnd 0.098066f
C276 a_n2650_8322.n23 gnd 0.690775f
C277 a_n2650_8322.n24 gnd 0.771841f
C278 a_n2650_8322.n25 gnd 0.39216f
C279 a_n2650_8322.n26 gnd 0.690777f
C280 a_n2650_8322.t27 gnd 0.098066f
C281 minus.n0 gnd 0.030241f
C282 minus.t14 gnd 0.50849f
C283 minus.n1 gnd 0.205656f
C284 minus.n2 gnd 0.030241f
C285 minus.t19 gnd 0.50849f
C286 minus.n3 gnd 0.024579f
C287 minus.n4 gnd 0.030241f
C288 minus.t18 gnd 0.50849f
C289 minus.t5 gnd 0.50849f
C290 minus.n5 gnd 0.205656f
C291 minus.n6 gnd 0.030241f
C292 minus.t8 gnd 0.50849f
C293 minus.n7 gnd 0.205656f
C294 minus.n8 gnd 0.129811f
C295 minus.t9 gnd 0.50849f
C296 minus.t13 gnd 0.570901f
C297 minus.n9 gnd 0.238618f
C298 minus.n10 gnd 0.237501f
C299 minus.n11 gnd 0.037617f
C300 minus.n12 gnd 0.035353f
C301 minus.n13 gnd 0.030241f
C302 minus.n14 gnd 0.030241f
C303 minus.n15 gnd 0.037881f
C304 minus.n16 gnd 0.024579f
C305 minus.n17 gnd 0.038903f
C306 minus.n18 gnd 0.030241f
C307 minus.n19 gnd 0.030241f
C308 minus.n20 gnd 0.036485f
C309 minus.n21 gnd 0.036485f
C310 minus.n22 gnd 0.205656f
C311 minus.n23 gnd 0.038903f
C312 minus.n24 gnd 0.030241f
C313 minus.n25 gnd 0.030241f
C314 minus.n26 gnd 0.030241f
C315 minus.n27 gnd 0.037881f
C316 minus.n28 gnd 0.205656f
C317 minus.n29 gnd 0.035353f
C318 minus.n30 gnd 0.037617f
C319 minus.n31 gnd 0.030241f
C320 minus.n32 gnd 0.030241f
C321 minus.n33 gnd 0.039384f
C322 minus.n34 gnd 0.012525f
C323 minus.t17 gnd 0.549932f
C324 minus.n35 gnd 0.238861f
C325 minus.n36 gnd 0.355332f
C326 minus.n37 gnd 0.030241f
C327 minus.t15 gnd 0.549932f
C328 minus.t12 gnd 0.50849f
C329 minus.n38 gnd 0.205656f
C330 minus.n39 gnd 0.030241f
C331 minus.t7 gnd 0.50849f
C332 minus.n40 gnd 0.024579f
C333 minus.n41 gnd 0.030241f
C334 minus.t6 gnd 0.50849f
C335 minus.t11 gnd 0.50849f
C336 minus.n42 gnd 0.205656f
C337 minus.n43 gnd 0.030241f
C338 minus.t10 gnd 0.50849f
C339 minus.n44 gnd 0.205656f
C340 minus.n45 gnd 0.129811f
C341 minus.t16 gnd 0.50849f
C342 minus.t20 gnd 0.570901f
C343 minus.n46 gnd 0.238618f
C344 minus.n47 gnd 0.237501f
C345 minus.n48 gnd 0.037617f
C346 minus.n49 gnd 0.035353f
C347 minus.n50 gnd 0.030241f
C348 minus.n51 gnd 0.030241f
C349 minus.n52 gnd 0.037881f
C350 minus.n53 gnd 0.024579f
C351 minus.n54 gnd 0.038903f
C352 minus.n55 gnd 0.030241f
C353 minus.n56 gnd 0.030241f
C354 minus.n57 gnd 0.036485f
C355 minus.n58 gnd 0.036485f
C356 minus.n59 gnd 0.205656f
C357 minus.n60 gnd 0.038903f
C358 minus.n61 gnd 0.030241f
C359 minus.n62 gnd 0.030241f
C360 minus.n63 gnd 0.030241f
C361 minus.n64 gnd 0.037881f
C362 minus.n65 gnd 0.205656f
C363 minus.n66 gnd 0.035353f
C364 minus.n67 gnd 0.037617f
C365 minus.n68 gnd 0.030241f
C366 minus.n69 gnd 0.030241f
C367 minus.n70 gnd 0.039384f
C368 minus.n71 gnd 0.012525f
C369 minus.n72 gnd 0.238861f
C370 minus.n73 gnd 0.942282f
C371 minus.n74 gnd 1.41632f
C372 minus.t1 gnd 0.009322f
C373 minus.t4 gnd 0.009322f
C374 minus.n75 gnd 0.030654f
C375 minus.t2 gnd 0.009322f
C376 minus.t0 gnd 0.009322f
C377 minus.n76 gnd 0.030234f
C378 minus.n77 gnd 0.258032f
C379 minus.t3 gnd 0.051887f
C380 minus.n78 gnd 0.140806f
C381 minus.n79 gnd 1.82867f
C382 a_n2903_n3924.n0 gnd 1.45586f
C383 a_n2903_n3924.t6 gnd 0.088483f
C384 a_n2903_n3924.t15 gnd 0.919619f
C385 a_n2903_n3924.n1 gnd 0.347657f
C386 a_n2903_n3924.t24 gnd 1.14306f
C387 a_n2903_n3924.n2 gnd 1.19083f
C388 a_n2903_n3924.t32 gnd 0.919619f
C389 a_n2903_n3924.n3 gnd 0.347657f
C390 a_n2903_n3924.t33 gnd 0.088483f
C391 a_n2903_n3924.t1 gnd 0.088483f
C392 a_n2903_n3924.n4 gnd 0.722655f
C393 a_n2903_n3924.n5 gnd 0.364177f
C394 a_n2903_n3924.t34 gnd 0.088483f
C395 a_n2903_n3924.t26 gnd 0.088483f
C396 a_n2903_n3924.n6 gnd 0.722655f
C397 a_n2903_n3924.n7 gnd 0.364177f
C398 a_n2903_n3924.t35 gnd 0.088483f
C399 a_n2903_n3924.t2 gnd 0.088483f
C400 a_n2903_n3924.n8 gnd 0.722655f
C401 a_n2903_n3924.n9 gnd 0.364177f
C402 a_n2903_n3924.t29 gnd 0.919619f
C403 a_n2903_n3924.n10 gnd 0.860834f
C404 a_n2903_n3924.t27 gnd 1.14419f
C405 a_n2903_n3924.t36 gnd 1.14261f
C406 a_n2903_n3924.n11 gnd 0.745791f
C407 a_n2903_n3924.t25 gnd 1.14261f
C408 a_n2903_n3924.n12 gnd 0.804756f
C409 a_n2903_n3924.t20 gnd 1.14261f
C410 a_n2903_n3924.n13 gnd 0.804756f
C411 a_n2903_n3924.t37 gnd 1.14261f
C412 a_n2903_n3924.n14 gnd 0.804756f
C413 a_n2903_n3924.t21 gnd 1.14261f
C414 a_n2903_n3924.n15 gnd 0.804756f
C415 a_n2903_n3924.t30 gnd 1.14261f
C416 a_n2903_n3924.n16 gnd 0.834168f
C417 a_n2903_n3924.t17 gnd 0.919616f
C418 a_n2903_n3924.n17 gnd 0.571219f
C419 a_n2903_n3924.t18 gnd 0.088483f
C420 a_n2903_n3924.t8 gnd 0.088483f
C421 a_n2903_n3924.n18 gnd 0.722654f
C422 a_n2903_n3924.n19 gnd 0.364178f
C423 a_n2903_n3924.t9 gnd 0.088483f
C424 a_n2903_n3924.t4 gnd 0.088483f
C425 a_n2903_n3924.n20 gnd 0.722654f
C426 a_n2903_n3924.n21 gnd 0.364178f
C427 a_n2903_n3924.t5 gnd 0.088483f
C428 a_n2903_n3924.t16 gnd 0.088483f
C429 a_n2903_n3924.n22 gnd 0.722654f
C430 a_n2903_n3924.n23 gnd 0.364178f
C431 a_n2903_n3924.t13 gnd 0.919616f
C432 a_n2903_n3924.n24 gnd 0.347661f
C433 a_n2903_n3924.t39 gnd 0.919616f
C434 a_n2903_n3924.n25 gnd 0.347661f
C435 a_n2903_n3924.t38 gnd 0.088483f
C436 a_n2903_n3924.t0 gnd 0.088483f
C437 a_n2903_n3924.n26 gnd 0.722654f
C438 a_n2903_n3924.n27 gnd 0.364178f
C439 a_n2903_n3924.t31 gnd 0.088483f
C440 a_n2903_n3924.t23 gnd 0.088483f
C441 a_n2903_n3924.n28 gnd 0.722654f
C442 a_n2903_n3924.n29 gnd 0.364178f
C443 a_n2903_n3924.t22 gnd 0.088483f
C444 a_n2903_n3924.t28 gnd 0.088483f
C445 a_n2903_n3924.n30 gnd 0.722654f
C446 a_n2903_n3924.n31 gnd 0.364178f
C447 a_n2903_n3924.t3 gnd 0.919616f
C448 a_n2903_n3924.n32 gnd 0.571219f
C449 a_n2903_n3924.n33 gnd 0.834168f
C450 a_n2903_n3924.t12 gnd 0.919616f
C451 a_n2903_n3924.n34 gnd 0.860837f
C452 a_n2903_n3924.t10 gnd 0.088483f
C453 a_n2903_n3924.t14 gnd 0.088483f
C454 a_n2903_n3924.n35 gnd 0.722655f
C455 a_n2903_n3924.n36 gnd 0.364177f
C456 a_n2903_n3924.t7 gnd 0.088483f
C457 a_n2903_n3924.t11 gnd 0.088483f
C458 a_n2903_n3924.n37 gnd 0.722655f
C459 a_n2903_n3924.n38 gnd 0.364177f
C460 a_n2903_n3924.n39 gnd 0.364176f
C461 a_n2903_n3924.n40 gnd 0.722656f
C462 a_n2903_n3924.t19 gnd 0.088483f
C463 plus.n0 gnd 0.022174f
C464 plus.t7 gnd 0.40324f
C465 plus.t6 gnd 0.372852f
C466 plus.n1 gnd 0.150798f
C467 plus.n2 gnd 0.022174f
C468 plus.t16 gnd 0.372852f
C469 plus.n3 gnd 0.018023f
C470 plus.n4 gnd 0.022174f
C471 plus.t15 gnd 0.372852f
C472 plus.t20 gnd 0.372852f
C473 plus.n5 gnd 0.150798f
C474 plus.n6 gnd 0.022174f
C475 plus.t19 gnd 0.372852f
C476 plus.n7 gnd 0.150798f
C477 plus.n8 gnd 0.095184f
C478 plus.t8 gnd 0.372852f
C479 plus.t11 gnd 0.418615f
C480 plus.n9 gnd 0.174967f
C481 plus.n10 gnd 0.174148f
C482 plus.n11 gnd 0.027583f
C483 plus.n12 gnd 0.025922f
C484 plus.n13 gnd 0.022174f
C485 plus.n14 gnd 0.022174f
C486 plus.n15 gnd 0.027777f
C487 plus.n16 gnd 0.018023f
C488 plus.n17 gnd 0.028526f
C489 plus.n18 gnd 0.022174f
C490 plus.n19 gnd 0.022174f
C491 plus.n20 gnd 0.026752f
C492 plus.n21 gnd 0.026752f
C493 plus.n22 gnd 0.150798f
C494 plus.n23 gnd 0.028526f
C495 plus.n24 gnd 0.022174f
C496 plus.n25 gnd 0.022174f
C497 plus.n26 gnd 0.022174f
C498 plus.n27 gnd 0.027777f
C499 plus.n28 gnd 0.150798f
C500 plus.n29 gnd 0.025922f
C501 plus.n30 gnd 0.027583f
C502 plus.n31 gnd 0.022174f
C503 plus.n32 gnd 0.022174f
C504 plus.n33 gnd 0.028879f
C505 plus.n34 gnd 0.009184f
C506 plus.n35 gnd 0.175146f
C507 plus.n36 gnd 0.254846f
C508 plus.n37 gnd 0.022174f
C509 plus.t10 gnd 0.372852f
C510 plus.n38 gnd 0.150798f
C511 plus.n39 gnd 0.022174f
C512 plus.t14 gnd 0.372852f
C513 plus.n40 gnd 0.018023f
C514 plus.n41 gnd 0.022174f
C515 plus.t13 gnd 0.372852f
C516 plus.t17 gnd 0.372852f
C517 plus.n42 gnd 0.150798f
C518 plus.n43 gnd 0.022174f
C519 plus.t18 gnd 0.372852f
C520 plus.n44 gnd 0.150798f
C521 plus.n45 gnd 0.095184f
C522 plus.t5 gnd 0.372852f
C523 plus.t9 gnd 0.418615f
C524 plus.n46 gnd 0.174967f
C525 plus.n47 gnd 0.174148f
C526 plus.n48 gnd 0.027583f
C527 plus.n49 gnd 0.025922f
C528 plus.n50 gnd 0.022174f
C529 plus.n51 gnd 0.022174f
C530 plus.n52 gnd 0.027777f
C531 plus.n53 gnd 0.018023f
C532 plus.n54 gnd 0.028526f
C533 plus.n55 gnd 0.022174f
C534 plus.n56 gnd 0.022174f
C535 plus.n57 gnd 0.026752f
C536 plus.n58 gnd 0.026752f
C537 plus.n59 gnd 0.150798f
C538 plus.n60 gnd 0.028526f
C539 plus.n61 gnd 0.022174f
C540 plus.n62 gnd 0.022174f
C541 plus.n63 gnd 0.022174f
C542 plus.n64 gnd 0.027777f
C543 plus.n65 gnd 0.150798f
C544 plus.n66 gnd 0.025922f
C545 plus.n67 gnd 0.027583f
C546 plus.n68 gnd 0.022174f
C547 plus.n69 gnd 0.022174f
C548 plus.n70 gnd 0.028879f
C549 plus.n71 gnd 0.009184f
C550 plus.t12 gnd 0.40324f
C551 plus.n72 gnd 0.175146f
C552 plus.n73 gnd 0.682047f
C553 plus.n74 gnd 1.02974f
C554 plus.t4 gnd 0.038279f
C555 plus.t1 gnd 0.006836f
C556 plus.t2 gnd 0.006836f
C557 plus.n75 gnd 0.022169f
C558 plus.n76 gnd 0.1721f
C559 plus.t0 gnd 0.006836f
C560 plus.t3 gnd 0.006836f
C561 plus.n77 gnd 0.022169f
C562 plus.n78 gnd 0.129182f
C563 plus.n79 gnd 2.40955f
C564 output.t8 gnd 0.464308f
C565 output.t15 gnd 0.044422f
C566 output.t4 gnd 0.044422f
C567 output.n0 gnd 0.364624f
C568 output.n1 gnd 0.614102f
C569 output.t6 gnd 0.044422f
C570 output.t11 gnd 0.044422f
C571 output.n2 gnd 0.364624f
C572 output.n3 gnd 0.350265f
C573 output.t16 gnd 0.044422f
C574 output.t2 gnd 0.044422f
C575 output.n4 gnd 0.364624f
C576 output.n5 gnd 0.350265f
C577 output.t3 gnd 0.044422f
C578 output.t9 gnd 0.044422f
C579 output.n6 gnd 0.364624f
C580 output.n7 gnd 0.350265f
C581 output.t12 gnd 0.044422f
C582 output.t5 gnd 0.044422f
C583 output.n8 gnd 0.364624f
C584 output.n9 gnd 0.350265f
C585 output.t7 gnd 0.044422f
C586 output.t13 gnd 0.044422f
C587 output.n10 gnd 0.364624f
C588 output.n11 gnd 0.350265f
C589 output.t14 gnd 0.044422f
C590 output.t17 gnd 0.044422f
C591 output.n12 gnd 0.364624f
C592 output.n13 gnd 0.350265f
C593 output.t10 gnd 0.462979f
C594 output.n14 gnd 0.28994f
C595 output.n15 gnd 0.015803f
C596 output.n16 gnd 0.011243f
C597 output.n17 gnd 0.006041f
C598 output.n18 gnd 0.01428f
C599 output.n19 gnd 0.006397f
C600 output.n20 gnd 0.011243f
C601 output.n21 gnd 0.006041f
C602 output.n22 gnd 0.01428f
C603 output.n23 gnd 0.006397f
C604 output.n24 gnd 0.048111f
C605 output.t1 gnd 0.023274f
C606 output.n25 gnd 0.01071f
C607 output.n26 gnd 0.008435f
C608 output.n27 gnd 0.006041f
C609 output.n28 gnd 0.267512f
C610 output.n29 gnd 0.011243f
C611 output.n30 gnd 0.006041f
C612 output.n31 gnd 0.006397f
C613 output.n32 gnd 0.01428f
C614 output.n33 gnd 0.01428f
C615 output.n34 gnd 0.006397f
C616 output.n35 gnd 0.006041f
C617 output.n36 gnd 0.011243f
C618 output.n37 gnd 0.011243f
C619 output.n38 gnd 0.006041f
C620 output.n39 gnd 0.006397f
C621 output.n40 gnd 0.01428f
C622 output.n41 gnd 0.030913f
C623 output.n42 gnd 0.006397f
C624 output.n43 gnd 0.006041f
C625 output.n44 gnd 0.025987f
C626 output.n45 gnd 0.097665f
C627 output.n46 gnd 0.015803f
C628 output.n47 gnd 0.011243f
C629 output.n48 gnd 0.006041f
C630 output.n49 gnd 0.01428f
C631 output.n50 gnd 0.006397f
C632 output.n51 gnd 0.011243f
C633 output.n52 gnd 0.006041f
C634 output.n53 gnd 0.01428f
C635 output.n54 gnd 0.006397f
C636 output.n55 gnd 0.048111f
C637 output.t0 gnd 0.023274f
C638 output.n56 gnd 0.01071f
C639 output.n57 gnd 0.008435f
C640 output.n58 gnd 0.006041f
C641 output.n59 gnd 0.267512f
C642 output.n60 gnd 0.011243f
C643 output.n61 gnd 0.006041f
C644 output.n62 gnd 0.006397f
C645 output.n63 gnd 0.01428f
C646 output.n64 gnd 0.01428f
C647 output.n65 gnd 0.006397f
C648 output.n66 gnd 0.006041f
C649 output.n67 gnd 0.011243f
C650 output.n68 gnd 0.011243f
C651 output.n69 gnd 0.006041f
C652 output.n70 gnd 0.006397f
C653 output.n71 gnd 0.01428f
C654 output.n72 gnd 0.030913f
C655 output.n73 gnd 0.006397f
C656 output.n74 gnd 0.006041f
C657 output.n75 gnd 0.025987f
C658 output.n76 gnd 0.09306f
C659 output.n77 gnd 1.65264f
C660 output.n78 gnd 0.015803f
C661 output.n79 gnd 0.011243f
C662 output.n80 gnd 0.006041f
C663 output.n81 gnd 0.01428f
C664 output.n82 gnd 0.006397f
C665 output.n83 gnd 0.011243f
C666 output.n84 gnd 0.006041f
C667 output.n85 gnd 0.01428f
C668 output.n86 gnd 0.006397f
C669 output.n87 gnd 0.048111f
C670 output.t18 gnd 0.023274f
C671 output.n88 gnd 0.01071f
C672 output.n89 gnd 0.008435f
C673 output.n90 gnd 0.006041f
C674 output.n91 gnd 0.267512f
C675 output.n92 gnd 0.011243f
C676 output.n93 gnd 0.006041f
C677 output.n94 gnd 0.006397f
C678 output.n95 gnd 0.01428f
C679 output.n96 gnd 0.01428f
C680 output.n97 gnd 0.006397f
C681 output.n98 gnd 0.006041f
C682 output.n99 gnd 0.011243f
C683 output.n100 gnd 0.011243f
C684 output.n101 gnd 0.006041f
C685 output.n102 gnd 0.006397f
C686 output.n103 gnd 0.01428f
C687 output.n104 gnd 0.030913f
C688 output.n105 gnd 0.006397f
C689 output.n106 gnd 0.006041f
C690 output.n107 gnd 0.025987f
C691 output.n108 gnd 0.09306f
C692 output.n109 gnd 0.713089f
C693 output.n110 gnd 0.015803f
C694 output.n111 gnd 0.011243f
C695 output.n112 gnd 0.006041f
C696 output.n113 gnd 0.01428f
C697 output.n114 gnd 0.006397f
C698 output.n115 gnd 0.011243f
C699 output.n116 gnd 0.006041f
C700 output.n117 gnd 0.01428f
C701 output.n118 gnd 0.006397f
C702 output.n119 gnd 0.048111f
C703 output.t19 gnd 0.023274f
C704 output.n120 gnd 0.01071f
C705 output.n121 gnd 0.008435f
C706 output.n122 gnd 0.006041f
C707 output.n123 gnd 0.267512f
C708 output.n124 gnd 0.011243f
C709 output.n125 gnd 0.006041f
C710 output.n126 gnd 0.006397f
C711 output.n127 gnd 0.01428f
C712 output.n128 gnd 0.01428f
C713 output.n129 gnd 0.006397f
C714 output.n130 gnd 0.006041f
C715 output.n131 gnd 0.011243f
C716 output.n132 gnd 0.011243f
C717 output.n133 gnd 0.006041f
C718 output.n134 gnd 0.006397f
C719 output.n135 gnd 0.01428f
C720 output.n136 gnd 0.030913f
C721 output.n137 gnd 0.006397f
C722 output.n138 gnd 0.006041f
C723 output.n139 gnd 0.025987f
C724 output.n140 gnd 0.09306f
C725 output.n141 gnd 1.67353f
C726 a_n2472_13878.t13 gnd 0.187752f
C727 a_n2472_13878.t15 gnd 0.187752f
C728 a_n2472_13878.t7 gnd 0.187752f
C729 a_n2472_13878.n0 gnd 1.47995f
C730 a_n2472_13878.t12 gnd 0.187752f
C731 a_n2472_13878.t6 gnd 0.187752f
C732 a_n2472_13878.n1 gnd 1.47838f
C733 a_n2472_13878.n2 gnd 2.06575f
C734 a_n2472_13878.t2 gnd 0.187752f
C735 a_n2472_13878.t4 gnd 0.187752f
C736 a_n2472_13878.n3 gnd 1.47838f
C737 a_n2472_13878.n4 gnd 1.00763f
C738 a_n2472_13878.t14 gnd 0.187752f
C739 a_n2472_13878.t3 gnd 0.187752f
C740 a_n2472_13878.n5 gnd 1.47838f
C741 a_n2472_13878.n6 gnd 1.00763f
C742 a_n2472_13878.t11 gnd 0.187752f
C743 a_n2472_13878.t1 gnd 0.187752f
C744 a_n2472_13878.n7 gnd 1.47838f
C745 a_n2472_13878.n8 gnd 4.40971f
C746 a_n2472_13878.t21 gnd 1.75801f
C747 a_n2472_13878.t24 gnd 0.187752f
C748 a_n2472_13878.t25 gnd 0.187752f
C749 a_n2472_13878.n9 gnd 1.32252f
C750 a_n2472_13878.n10 gnd 1.47772f
C751 a_n2472_13878.t20 gnd 1.75451f
C752 a_n2472_13878.n11 gnd 0.743612f
C753 a_n2472_13878.t23 gnd 1.75451f
C754 a_n2472_13878.n12 gnd 0.743612f
C755 a_n2472_13878.t26 gnd 0.187752f
C756 a_n2472_13878.t27 gnd 0.187752f
C757 a_n2472_13878.n13 gnd 1.32252f
C758 a_n2472_13878.n14 gnd 0.750813f
C759 a_n2472_13878.t22 gnd 1.75451f
C760 a_n2472_13878.n15 gnd 2.43968f
C761 a_n2472_13878.n16 gnd 3.23176f
C762 a_n2472_13878.t16 gnd 0.187752f
C763 a_n2472_13878.t5 gnd 0.187752f
C764 a_n2472_13878.n17 gnd 1.47838f
C765 a_n2472_13878.n18 gnd 2.22265f
C766 a_n2472_13878.t8 gnd 0.187752f
C767 a_n2472_13878.t9 gnd 0.187752f
C768 a_n2472_13878.n19 gnd 1.47838f
C769 a_n2472_13878.n20 gnd 0.655033f
C770 a_n2472_13878.t17 gnd 0.187752f
C771 a_n2472_13878.t18 gnd 0.187752f
C772 a_n2472_13878.n21 gnd 1.47838f
C773 a_n2472_13878.n22 gnd 0.655033f
C774 a_n2472_13878.t0 gnd 0.187752f
C775 a_n2472_13878.t10 gnd 0.187752f
C776 a_n2472_13878.n23 gnd 1.47838f
C777 a_n2472_13878.n24 gnd 1.32888f
C778 a_n2472_13878.n25 gnd 1.48083f
C779 a_n2472_13878.t19 gnd 0.187752f
C780 a_n2650_13878.n0 gnd 2.71632f
C781 a_n2650_13878.n1 gnd 3.9242f
C782 a_n2650_13878.n2 gnd 3.79431f
C783 a_n2650_13878.n3 gnd 0.209626f
C784 a_n2650_13878.n4 gnd 0.209626f
C785 a_n2650_13878.n5 gnd 0.779569f
C786 a_n2650_13878.n6 gnd 0.209626f
C787 a_n2650_13878.n7 gnd 0.907703f
C788 a_n2650_13878.n8 gnd 0.209626f
C789 a_n2650_13878.n9 gnd 0.487486f
C790 a_n2650_13878.n10 gnd 0.779488f
C791 a_n2650_13878.n11 gnd 0.198901f
C792 a_n2650_13878.n12 gnd 0.146494f
C793 a_n2650_13878.n13 gnd 0.230242f
C794 a_n2650_13878.n14 gnd 0.177836f
C795 a_n2650_13878.n15 gnd 0.198901f
C796 a_n2650_13878.n16 gnd 1.20434f
C797 a_n2650_13878.n17 gnd 0.146494f
C798 a_n2650_13878.n18 gnd 0.831895f
C799 a_n2650_13878.n19 gnd 0.209626f
C800 a_n2650_13878.n20 gnd 0.676448f
C801 a_n2650_13878.n21 gnd 0.209626f
C802 a_n2650_13878.n22 gnd 0.488406f
C803 a_n2650_13878.n23 gnd 0.209626f
C804 a_n2650_13878.n24 gnd 0.540812f
C805 a_n2650_13878.n25 gnd 0.209626f
C806 a_n2650_13878.n26 gnd 0.867796f
C807 a_n2650_13878.n27 gnd 1.14438f
C808 a_n2650_13878.n28 gnd 1.16289f
C809 a_n2650_13878.n29 gnd 2.17246f
C810 a_n2650_13878.n30 gnd 1.72583f
C811 a_n2650_13878.n31 gnd 1.40392f
C812 a_n2650_13878.n32 gnd 1.16289f
C813 a_n2650_13878.n33 gnd 3.13153f
C814 a_n2650_13878.n34 gnd 0.008411f
C815 a_n2650_13878.n35 gnd 4.05e-19
C816 a_n2650_13878.n37 gnd 0.008116f
C817 a_n2650_13878.n38 gnd 0.011801f
C818 a_n2650_13878.n39 gnd 0.007808f
C819 a_n2650_13878.n40 gnd 0.276916f
C820 a_n2650_13878.n41 gnd 0.008411f
C821 a_n2650_13878.n42 gnd 4.05e-19
C822 a_n2650_13878.n44 gnd 0.008116f
C823 a_n2650_13878.n45 gnd 0.011801f
C824 a_n2650_13878.n46 gnd 0.007808f
C825 a_n2650_13878.n47 gnd 0.276916f
C826 a_n2650_13878.n48 gnd 0.008116f
C827 a_n2650_13878.n49 gnd 0.276916f
C828 a_n2650_13878.n50 gnd 0.008116f
C829 a_n2650_13878.n51 gnd 0.276916f
C830 a_n2650_13878.n52 gnd 0.008116f
C831 a_n2650_13878.n53 gnd 0.276916f
C832 a_n2650_13878.n54 gnd 0.008116f
C833 a_n2650_13878.n55 gnd 0.276916f
C834 a_n2650_13878.n56 gnd 0.008411f
C835 a_n2650_13878.n57 gnd 4.05e-19
C836 a_n2650_13878.n59 gnd 0.008116f
C837 a_n2650_13878.n60 gnd 0.011801f
C838 a_n2650_13878.n61 gnd 0.007808f
C839 a_n2650_13878.n62 gnd 0.276916f
C840 a_n2650_13878.n63 gnd 0.008411f
C841 a_n2650_13878.n64 gnd 4.05e-19
C842 a_n2650_13878.n66 gnd 0.008116f
C843 a_n2650_13878.n67 gnd 0.011801f
C844 a_n2650_13878.n68 gnd 0.007808f
C845 a_n2650_13878.n69 gnd 0.276916f
C846 a_n2650_13878.t25 gnd 0.145399f
C847 a_n2650_13878.t6 gnd 0.676325f
C848 a_n2650_13878.t30 gnd 0.676325f
C849 a_n2650_13878.t42 gnd 0.676325f
C850 a_n2650_13878.n70 gnd 0.297222f
C851 a_n2650_13878.t4 gnd 0.676325f
C852 a_n2650_13878.t24 gnd 0.676325f
C853 a_n2650_13878.t32 gnd 0.676325f
C854 a_n2650_13878.n71 gnd 0.293579f
C855 a_n2650_13878.t10 gnd 0.676325f
C856 a_n2650_13878.t8 gnd 0.676325f
C857 a_n2650_13878.t38 gnd 0.676325f
C858 a_n2650_13878.n72 gnd 0.29734f
C859 a_n2650_13878.t90 gnd 0.676325f
C860 a_n2650_13878.t69 gnd 0.676325f
C861 a_n2650_13878.t74 gnd 0.676325f
C862 a_n2650_13878.n73 gnd 0.297222f
C863 a_n2650_13878.t63 gnd 0.676325f
C864 a_n2650_13878.t79 gnd 0.676325f
C865 a_n2650_13878.t87 gnd 0.676325f
C866 a_n2650_13878.n74 gnd 0.293579f
C867 a_n2650_13878.t88 gnd 0.676325f
C868 a_n2650_13878.t58 gnd 0.676325f
C869 a_n2650_13878.t71 gnd 0.676325f
C870 a_n2650_13878.n75 gnd 0.29734f
C871 a_n2650_13878.t15 gnd 1.36144f
C872 a_n2650_13878.t27 gnd 0.145399f
C873 a_n2650_13878.t41 gnd 0.145399f
C874 a_n2650_13878.n76 gnd 1.02419f
C875 a_n2650_13878.t37 gnd 0.145399f
C876 a_n2650_13878.t19 gnd 0.145399f
C877 a_n2650_13878.n77 gnd 1.02419f
C878 a_n2650_13878.t29 gnd 0.145399f
C879 a_n2650_13878.t23 gnd 0.145399f
C880 a_n2650_13878.n78 gnd 1.02419f
C881 a_n2650_13878.t21 gnd 0.145399f
C882 a_n2650_13878.t13 gnd 0.145399f
C883 a_n2650_13878.n79 gnd 1.02419f
C884 a_n2650_13878.t35 gnd 1.35873f
C885 a_n2650_13878.t20 gnd 0.676325f
C886 a_n2650_13878.n80 gnd 0.293831f
C887 a_n2650_13878.t28 gnd 0.676325f
C888 a_n2650_13878.t40 gnd 0.676325f
C889 a_n2650_13878.n81 gnd 0.297222f
C890 a_n2650_13878.t14 gnd 0.676325f
C891 a_n2650_13878.t68 gnd 0.676325f
C892 a_n2650_13878.n82 gnd 0.293831f
C893 a_n2650_13878.t83 gnd 0.676325f
C894 a_n2650_13878.t86 gnd 0.676325f
C895 a_n2650_13878.n83 gnd 0.297222f
C896 a_n2650_13878.t62 gnd 0.676325f
C897 a_n2650_13878.n84 gnd 0.288248f
C898 a_n2650_13878.t85 gnd 0.676325f
C899 a_n2650_13878.n85 gnd 0.293256f
C900 a_n2650_13878.t60 gnd 0.676325f
C901 a_n2650_13878.n86 gnd 0.299896f
C902 a_n2650_13878.t82 gnd 0.676325f
C903 a_n2650_13878.n87 gnd 0.297355f
C904 a_n2650_13878.n88 gnd 0.293579f
C905 a_n2650_13878.t57 gnd 0.676325f
C906 a_n2650_13878.n89 gnd 0.288409f
C907 a_n2650_13878.t78 gnd 0.676325f
C908 a_n2650_13878.n90 gnd 0.29734f
C909 a_n2650_13878.t59 gnd 0.687657f
C910 a_n2650_13878.n91 gnd 0.288248f
C911 a_n2650_13878.t26 gnd 0.676325f
C912 a_n2650_13878.n92 gnd 0.293256f
C913 a_n2650_13878.t36 gnd 0.676325f
C914 a_n2650_13878.n93 gnd 0.299896f
C915 a_n2650_13878.t18 gnd 0.676325f
C916 a_n2650_13878.n94 gnd 0.297355f
C917 a_n2650_13878.n95 gnd 0.293579f
C918 a_n2650_13878.t22 gnd 0.676325f
C919 a_n2650_13878.n96 gnd 0.288409f
C920 a_n2650_13878.t12 gnd 0.676325f
C921 a_n2650_13878.n97 gnd 0.29734f
C922 a_n2650_13878.t34 gnd 0.687657f
C923 a_n2650_13878.n98 gnd 1.23608f
C924 a_n2650_13878.t66 gnd 0.676325f
C925 a_n2650_13878.n99 gnd 0.293579f
C926 a_n2650_13878.t73 gnd 0.676325f
C927 a_n2650_13878.n100 gnd 0.293579f
C928 a_n2650_13878.t64 gnd 0.676325f
C929 a_n2650_13878.n101 gnd 0.293579f
C930 a_n2650_13878.t77 gnd 0.676325f
C931 a_n2650_13878.n102 gnd 0.293579f
C932 a_n2650_13878.t67 gnd 0.676325f
C933 a_n2650_13878.n103 gnd 0.288248f
C934 a_n2650_13878.t91 gnd 0.676325f
C935 a_n2650_13878.n104 gnd 0.297355f
C936 a_n2650_13878.t70 gnd 0.687657f
C937 a_n2650_13878.t80 gnd 0.676325f
C938 a_n2650_13878.n105 gnd 0.288248f
C939 a_n2650_13878.t65 gnd 0.676325f
C940 a_n2650_13878.n106 gnd 0.297355f
C941 a_n2650_13878.t75 gnd 0.687657f
C942 a_n2650_13878.t84 gnd 0.676325f
C943 a_n2650_13878.n107 gnd 0.288248f
C944 a_n2650_13878.t72 gnd 0.676325f
C945 a_n2650_13878.n108 gnd 0.297355f
C946 a_n2650_13878.t89 gnd 0.687657f
C947 a_n2650_13878.t76 gnd 0.676325f
C948 a_n2650_13878.n109 gnd 0.288248f
C949 a_n2650_13878.t56 gnd 0.676325f
C950 a_n2650_13878.n110 gnd 0.297355f
C951 a_n2650_13878.t81 gnd 0.687657f
C952 a_n2650_13878.n111 gnd 1.52654f
C953 a_n2650_13878.t61 gnd 0.687657f
C954 a_n2650_13878.n112 gnd 0.293831f
C955 a_n2650_13878.n113 gnd 0.288409f
C956 a_n2650_13878.n114 gnd 0.297355f
C957 a_n2650_13878.n115 gnd 0.299896f
C958 a_n2650_13878.n116 gnd 0.293256f
C959 a_n2650_13878.n117 gnd 0.288248f
C960 a_n2650_13878.t16 gnd 0.687657f
C961 a_n2650_13878.t55 gnd 0.113088f
C962 a_n2650_13878.t54 gnd 0.113088f
C963 a_n2650_13878.n118 gnd 1.00223f
C964 a_n2650_13878.t0 gnd 0.113088f
C965 a_n2650_13878.t49 gnd 0.113088f
C966 a_n2650_13878.n119 gnd 0.999285f
C967 a_n2650_13878.t47 gnd 0.113088f
C968 a_n2650_13878.t3 gnd 0.113088f
C969 a_n2650_13878.n120 gnd 1.00223f
C970 a_n2650_13878.t45 gnd 0.113088f
C971 a_n2650_13878.t44 gnd 0.113088f
C972 a_n2650_13878.n121 gnd 0.999285f
C973 a_n2650_13878.t48 gnd 0.113088f
C974 a_n2650_13878.t53 gnd 0.113088f
C975 a_n2650_13878.n122 gnd 0.999285f
C976 a_n2650_13878.t2 gnd 0.113088f
C977 a_n2650_13878.t52 gnd 0.113088f
C978 a_n2650_13878.n123 gnd 0.999285f
C979 a_n2650_13878.t1 gnd 0.113088f
C980 a_n2650_13878.t50 gnd 0.113088f
C981 a_n2650_13878.n124 gnd 1.00223f
C982 a_n2650_13878.t46 gnd 0.113088f
C983 a_n2650_13878.t51 gnd 0.113088f
C984 a_n2650_13878.n125 gnd 0.999285f
C985 a_n2650_13878.n126 gnd 0.293831f
C986 a_n2650_13878.n127 gnd 0.288409f
C987 a_n2650_13878.n128 gnd 0.297355f
C988 a_n2650_13878.n129 gnd 0.299896f
C989 a_n2650_13878.n130 gnd 0.293256f
C990 a_n2650_13878.n131 gnd 0.288248f
C991 a_n2650_13878.n132 gnd 0.913993f
C992 a_n2650_13878.t7 gnd 1.35873f
C993 a_n2650_13878.t31 gnd 0.145399f
C994 a_n2650_13878.t43 gnd 0.145399f
C995 a_n2650_13878.n133 gnd 1.02419f
C996 a_n2650_13878.t17 gnd 1.36144f
C997 a_n2650_13878.t9 gnd 0.145399f
C998 a_n2650_13878.t39 gnd 0.145399f
C999 a_n2650_13878.n134 gnd 1.02419f
C1000 a_n2650_13878.t33 gnd 0.145399f
C1001 a_n2650_13878.t11 gnd 0.145399f
C1002 a_n2650_13878.n135 gnd 1.02419f
C1003 a_n2650_13878.n136 gnd 1.02419f
C1004 a_n2650_13878.t5 gnd 0.145399f
C1005 commonsourceibias.n0 gnd 0.012301f
C1006 commonsourceibias.t89 gnd 0.186271f
C1007 commonsourceibias.t51 gnd 0.172234f
C1008 commonsourceibias.n1 gnd 0.068721f
C1009 commonsourceibias.n2 gnd 0.009219f
C1010 commonsourceibias.t95 gnd 0.172234f
C1011 commonsourceibias.n3 gnd 0.007457f
C1012 commonsourceibias.n4 gnd 0.009219f
C1013 commonsourceibias.t90 gnd 0.172234f
C1014 commonsourceibias.n5 gnd 0.0089f
C1015 commonsourceibias.n6 gnd 0.009219f
C1016 commonsourceibias.t101 gnd 0.172234f
C1017 commonsourceibias.n7 gnd 0.068721f
C1018 commonsourceibias.t86 gnd 0.172234f
C1019 commonsourceibias.n8 gnd 0.007446f
C1020 commonsourceibias.n9 gnd 0.012301f
C1021 commonsourceibias.t6 gnd 0.186271f
C1022 commonsourceibias.t24 gnd 0.172234f
C1023 commonsourceibias.n10 gnd 0.068721f
C1024 commonsourceibias.n11 gnd 0.009219f
C1025 commonsourceibias.t20 gnd 0.172234f
C1026 commonsourceibias.n12 gnd 0.007457f
C1027 commonsourceibias.n13 gnd 0.009219f
C1028 commonsourceibias.t42 gnd 0.172234f
C1029 commonsourceibias.n14 gnd 0.0089f
C1030 commonsourceibias.n15 gnd 0.009219f
C1031 commonsourceibias.t10 gnd 0.172234f
C1032 commonsourceibias.n16 gnd 0.068721f
C1033 commonsourceibias.t40 gnd 0.172234f
C1034 commonsourceibias.n17 gnd 0.007446f
C1035 commonsourceibias.n18 gnd 0.009219f
C1036 commonsourceibias.t28 gnd 0.172234f
C1037 commonsourceibias.t46 gnd 0.172234f
C1038 commonsourceibias.n19 gnd 0.068721f
C1039 commonsourceibias.n20 gnd 0.009219f
C1040 commonsourceibias.t16 gnd 0.172234f
C1041 commonsourceibias.n21 gnd 0.068721f
C1042 commonsourceibias.n22 gnd 0.009219f
C1043 commonsourceibias.t26 gnd 0.172234f
C1044 commonsourceibias.n23 gnd 0.068721f
C1045 commonsourceibias.n24 gnd 0.046409f
C1046 commonsourceibias.t0 gnd 0.172234f
C1047 commonsourceibias.t30 gnd 0.194346f
C1048 commonsourceibias.n25 gnd 0.079751f
C1049 commonsourceibias.n26 gnd 0.082563f
C1050 commonsourceibias.n27 gnd 0.011362f
C1051 commonsourceibias.n28 gnd 0.01257f
C1052 commonsourceibias.n29 gnd 0.009219f
C1053 commonsourceibias.n30 gnd 0.009219f
C1054 commonsourceibias.n31 gnd 0.012488f
C1055 commonsourceibias.n32 gnd 0.007457f
C1056 commonsourceibias.n33 gnd 0.012643f
C1057 commonsourceibias.n34 gnd 0.009219f
C1058 commonsourceibias.n35 gnd 0.009219f
C1059 commonsourceibias.n36 gnd 0.01272f
C1060 commonsourceibias.n37 gnd 0.010968f
C1061 commonsourceibias.n38 gnd 0.0089f
C1062 commonsourceibias.n39 gnd 0.009219f
C1063 commonsourceibias.n40 gnd 0.009219f
C1064 commonsourceibias.n41 gnd 0.011276f
C1065 commonsourceibias.n42 gnd 0.012656f
C1066 commonsourceibias.n43 gnd 0.068721f
C1067 commonsourceibias.n44 gnd 0.012571f
C1068 commonsourceibias.n45 gnd 0.009219f
C1069 commonsourceibias.n46 gnd 0.009219f
C1070 commonsourceibias.n47 gnd 0.009219f
C1071 commonsourceibias.n48 gnd 0.012571f
C1072 commonsourceibias.n49 gnd 0.068721f
C1073 commonsourceibias.n50 gnd 0.012656f
C1074 commonsourceibias.n51 gnd 0.011276f
C1075 commonsourceibias.n52 gnd 0.009219f
C1076 commonsourceibias.n53 gnd 0.009219f
C1077 commonsourceibias.n54 gnd 0.009219f
C1078 commonsourceibias.n55 gnd 0.010968f
C1079 commonsourceibias.n56 gnd 0.01272f
C1080 commonsourceibias.n57 gnd 0.068721f
C1081 commonsourceibias.n58 gnd 0.012643f
C1082 commonsourceibias.n59 gnd 0.009219f
C1083 commonsourceibias.n60 gnd 0.009219f
C1084 commonsourceibias.n61 gnd 0.009219f
C1085 commonsourceibias.n62 gnd 0.012488f
C1086 commonsourceibias.n63 gnd 0.068721f
C1087 commonsourceibias.n64 gnd 0.01257f
C1088 commonsourceibias.n65 gnd 0.011362f
C1089 commonsourceibias.n66 gnd 0.009219f
C1090 commonsourceibias.n67 gnd 0.009219f
C1091 commonsourceibias.n68 gnd 0.009352f
C1092 commonsourceibias.n69 gnd 0.009668f
C1093 commonsourceibias.n70 gnd 0.082226f
C1094 commonsourceibias.n71 gnd 0.091217f
C1095 commonsourceibias.t7 gnd 0.019893f
C1096 commonsourceibias.t25 gnd 0.019893f
C1097 commonsourceibias.n72 gnd 0.175781f
C1098 commonsourceibias.n73 gnd 0.151888f
C1099 commonsourceibias.t21 gnd 0.019893f
C1100 commonsourceibias.t43 gnd 0.019893f
C1101 commonsourceibias.n74 gnd 0.175781f
C1102 commonsourceibias.n75 gnd 0.080743f
C1103 commonsourceibias.t11 gnd 0.019893f
C1104 commonsourceibias.t41 gnd 0.019893f
C1105 commonsourceibias.n76 gnd 0.175781f
C1106 commonsourceibias.n77 gnd 0.067457f
C1107 commonsourceibias.t1 gnd 0.019893f
C1108 commonsourceibias.t31 gnd 0.019893f
C1109 commonsourceibias.n78 gnd 0.17637f
C1110 commonsourceibias.t17 gnd 0.019893f
C1111 commonsourceibias.t27 gnd 0.019893f
C1112 commonsourceibias.n79 gnd 0.175781f
C1113 commonsourceibias.n80 gnd 0.163796f
C1114 commonsourceibias.t29 gnd 0.019893f
C1115 commonsourceibias.t47 gnd 0.019893f
C1116 commonsourceibias.n81 gnd 0.175781f
C1117 commonsourceibias.n82 gnd 0.067457f
C1118 commonsourceibias.n83 gnd 0.081684f
C1119 commonsourceibias.n84 gnd 0.009219f
C1120 commonsourceibias.t77 gnd 0.172234f
C1121 commonsourceibias.t94 gnd 0.172234f
C1122 commonsourceibias.n85 gnd 0.068721f
C1123 commonsourceibias.n86 gnd 0.009219f
C1124 commonsourceibias.t87 gnd 0.172234f
C1125 commonsourceibias.n87 gnd 0.068721f
C1126 commonsourceibias.n88 gnd 0.009219f
C1127 commonsourceibias.t58 gnd 0.172234f
C1128 commonsourceibias.n89 gnd 0.068721f
C1129 commonsourceibias.n90 gnd 0.046409f
C1130 commonsourceibias.t80 gnd 0.172234f
C1131 commonsourceibias.t73 gnd 0.194346f
C1132 commonsourceibias.n91 gnd 0.079751f
C1133 commonsourceibias.n92 gnd 0.082563f
C1134 commonsourceibias.n93 gnd 0.011362f
C1135 commonsourceibias.n94 gnd 0.01257f
C1136 commonsourceibias.n95 gnd 0.009219f
C1137 commonsourceibias.n96 gnd 0.009219f
C1138 commonsourceibias.n97 gnd 0.012488f
C1139 commonsourceibias.n98 gnd 0.007457f
C1140 commonsourceibias.n99 gnd 0.012643f
C1141 commonsourceibias.n100 gnd 0.009219f
C1142 commonsourceibias.n101 gnd 0.009219f
C1143 commonsourceibias.n102 gnd 0.01272f
C1144 commonsourceibias.n103 gnd 0.010968f
C1145 commonsourceibias.n104 gnd 0.0089f
C1146 commonsourceibias.n105 gnd 0.009219f
C1147 commonsourceibias.n106 gnd 0.009219f
C1148 commonsourceibias.n107 gnd 0.011276f
C1149 commonsourceibias.n108 gnd 0.012656f
C1150 commonsourceibias.n109 gnd 0.068721f
C1151 commonsourceibias.n110 gnd 0.012571f
C1152 commonsourceibias.n111 gnd 0.009174f
C1153 commonsourceibias.n112 gnd 0.06664f
C1154 commonsourceibias.n113 gnd 0.009174f
C1155 commonsourceibias.n114 gnd 0.012571f
C1156 commonsourceibias.n115 gnd 0.068721f
C1157 commonsourceibias.n116 gnd 0.012656f
C1158 commonsourceibias.n117 gnd 0.011276f
C1159 commonsourceibias.n118 gnd 0.009219f
C1160 commonsourceibias.n119 gnd 0.009219f
C1161 commonsourceibias.n120 gnd 0.009219f
C1162 commonsourceibias.n121 gnd 0.010968f
C1163 commonsourceibias.n122 gnd 0.01272f
C1164 commonsourceibias.n123 gnd 0.068721f
C1165 commonsourceibias.n124 gnd 0.012643f
C1166 commonsourceibias.n125 gnd 0.009219f
C1167 commonsourceibias.n126 gnd 0.009219f
C1168 commonsourceibias.n127 gnd 0.009219f
C1169 commonsourceibias.n128 gnd 0.012488f
C1170 commonsourceibias.n129 gnd 0.068721f
C1171 commonsourceibias.n130 gnd 0.01257f
C1172 commonsourceibias.n131 gnd 0.011362f
C1173 commonsourceibias.n132 gnd 0.009219f
C1174 commonsourceibias.n133 gnd 0.009219f
C1175 commonsourceibias.n134 gnd 0.009352f
C1176 commonsourceibias.n135 gnd 0.009668f
C1177 commonsourceibias.n136 gnd 0.082226f
C1178 commonsourceibias.n137 gnd 0.053232f
C1179 commonsourceibias.n138 gnd 0.012301f
C1180 commonsourceibias.t54 gnd 0.186271f
C1181 commonsourceibias.t119 gnd 0.172234f
C1182 commonsourceibias.n139 gnd 0.068721f
C1183 commonsourceibias.n140 gnd 0.009219f
C1184 commonsourceibias.t110 gnd 0.172234f
C1185 commonsourceibias.n141 gnd 0.007457f
C1186 commonsourceibias.n142 gnd 0.009219f
C1187 commonsourceibias.t60 gnd 0.172234f
C1188 commonsourceibias.n143 gnd 0.0089f
C1189 commonsourceibias.n144 gnd 0.009219f
C1190 commonsourceibias.t117 gnd 0.172234f
C1191 commonsourceibias.n145 gnd 0.068721f
C1192 commonsourceibias.t65 gnd 0.172234f
C1193 commonsourceibias.n146 gnd 0.007446f
C1194 commonsourceibias.n147 gnd 0.009219f
C1195 commonsourceibias.t59 gnd 0.172234f
C1196 commonsourceibias.t118 gnd 0.172234f
C1197 commonsourceibias.n148 gnd 0.068721f
C1198 commonsourceibias.n149 gnd 0.009219f
C1199 commonsourceibias.t71 gnd 0.172234f
C1200 commonsourceibias.n150 gnd 0.068721f
C1201 commonsourceibias.n151 gnd 0.009219f
C1202 commonsourceibias.t83 gnd 0.172234f
C1203 commonsourceibias.n152 gnd 0.068721f
C1204 commonsourceibias.n153 gnd 0.046409f
C1205 commonsourceibias.t116 gnd 0.172234f
C1206 commonsourceibias.t70 gnd 0.194346f
C1207 commonsourceibias.n154 gnd 0.079751f
C1208 commonsourceibias.n155 gnd 0.082563f
C1209 commonsourceibias.n156 gnd 0.011362f
C1210 commonsourceibias.n157 gnd 0.01257f
C1211 commonsourceibias.n158 gnd 0.009219f
C1212 commonsourceibias.n159 gnd 0.009219f
C1213 commonsourceibias.n160 gnd 0.012488f
C1214 commonsourceibias.n161 gnd 0.007457f
C1215 commonsourceibias.n162 gnd 0.012643f
C1216 commonsourceibias.n163 gnd 0.009219f
C1217 commonsourceibias.n164 gnd 0.009219f
C1218 commonsourceibias.n165 gnd 0.01272f
C1219 commonsourceibias.n166 gnd 0.010968f
C1220 commonsourceibias.n167 gnd 0.0089f
C1221 commonsourceibias.n168 gnd 0.009219f
C1222 commonsourceibias.n169 gnd 0.009219f
C1223 commonsourceibias.n170 gnd 0.011276f
C1224 commonsourceibias.n171 gnd 0.012656f
C1225 commonsourceibias.n172 gnd 0.068721f
C1226 commonsourceibias.n173 gnd 0.012571f
C1227 commonsourceibias.n174 gnd 0.009219f
C1228 commonsourceibias.n175 gnd 0.009219f
C1229 commonsourceibias.n176 gnd 0.009219f
C1230 commonsourceibias.n177 gnd 0.012571f
C1231 commonsourceibias.n178 gnd 0.068721f
C1232 commonsourceibias.n179 gnd 0.012656f
C1233 commonsourceibias.n180 gnd 0.011276f
C1234 commonsourceibias.n181 gnd 0.009219f
C1235 commonsourceibias.n182 gnd 0.009219f
C1236 commonsourceibias.n183 gnd 0.009219f
C1237 commonsourceibias.n184 gnd 0.010968f
C1238 commonsourceibias.n185 gnd 0.01272f
C1239 commonsourceibias.n186 gnd 0.068721f
C1240 commonsourceibias.n187 gnd 0.012643f
C1241 commonsourceibias.n188 gnd 0.009219f
C1242 commonsourceibias.n189 gnd 0.009219f
C1243 commonsourceibias.n190 gnd 0.009219f
C1244 commonsourceibias.n191 gnd 0.012488f
C1245 commonsourceibias.n192 gnd 0.068721f
C1246 commonsourceibias.n193 gnd 0.01257f
C1247 commonsourceibias.n194 gnd 0.011362f
C1248 commonsourceibias.n195 gnd 0.009219f
C1249 commonsourceibias.n196 gnd 0.009219f
C1250 commonsourceibias.n197 gnd 0.009352f
C1251 commonsourceibias.n198 gnd 0.009668f
C1252 commonsourceibias.n199 gnd 0.082226f
C1253 commonsourceibias.n200 gnd 0.027982f
C1254 commonsourceibias.n201 gnd 0.147096f
C1255 commonsourceibias.n202 gnd 0.012301f
C1256 commonsourceibias.t57 gnd 0.172234f
C1257 commonsourceibias.n203 gnd 0.068721f
C1258 commonsourceibias.n204 gnd 0.009219f
C1259 commonsourceibias.t96 gnd 0.172234f
C1260 commonsourceibias.n205 gnd 0.007457f
C1261 commonsourceibias.n206 gnd 0.009219f
C1262 commonsourceibias.t93 gnd 0.172234f
C1263 commonsourceibias.n207 gnd 0.0089f
C1264 commonsourceibias.n208 gnd 0.009219f
C1265 commonsourceibias.t115 gnd 0.172234f
C1266 commonsourceibias.n209 gnd 0.068721f
C1267 commonsourceibias.t68 gnd 0.172234f
C1268 commonsourceibias.n210 gnd 0.007446f
C1269 commonsourceibias.n211 gnd 0.009219f
C1270 commonsourceibias.t88 gnd 0.172234f
C1271 commonsourceibias.t108 gnd 0.172234f
C1272 commonsourceibias.n212 gnd 0.068721f
C1273 commonsourceibias.n213 gnd 0.009219f
C1274 commonsourceibias.t103 gnd 0.172234f
C1275 commonsourceibias.n214 gnd 0.068721f
C1276 commonsourceibias.n215 gnd 0.009219f
C1277 commonsourceibias.t48 gnd 0.172234f
C1278 commonsourceibias.n216 gnd 0.068721f
C1279 commonsourceibias.n217 gnd 0.046409f
C1280 commonsourceibias.t102 gnd 0.172234f
C1281 commonsourceibias.t98 gnd 0.194346f
C1282 commonsourceibias.n218 gnd 0.079751f
C1283 commonsourceibias.n219 gnd 0.082563f
C1284 commonsourceibias.n220 gnd 0.011362f
C1285 commonsourceibias.n221 gnd 0.01257f
C1286 commonsourceibias.n222 gnd 0.009219f
C1287 commonsourceibias.n223 gnd 0.009219f
C1288 commonsourceibias.n224 gnd 0.012488f
C1289 commonsourceibias.n225 gnd 0.007457f
C1290 commonsourceibias.n226 gnd 0.012643f
C1291 commonsourceibias.n227 gnd 0.009219f
C1292 commonsourceibias.n228 gnd 0.009219f
C1293 commonsourceibias.n229 gnd 0.01272f
C1294 commonsourceibias.n230 gnd 0.010968f
C1295 commonsourceibias.n231 gnd 0.0089f
C1296 commonsourceibias.n232 gnd 0.009219f
C1297 commonsourceibias.n233 gnd 0.009219f
C1298 commonsourceibias.n234 gnd 0.011276f
C1299 commonsourceibias.n235 gnd 0.012656f
C1300 commonsourceibias.n236 gnd 0.068721f
C1301 commonsourceibias.n237 gnd 0.012571f
C1302 commonsourceibias.n238 gnd 0.009219f
C1303 commonsourceibias.n239 gnd 0.009219f
C1304 commonsourceibias.n240 gnd 0.009219f
C1305 commonsourceibias.n241 gnd 0.012571f
C1306 commonsourceibias.n242 gnd 0.068721f
C1307 commonsourceibias.n243 gnd 0.012656f
C1308 commonsourceibias.n244 gnd 0.011276f
C1309 commonsourceibias.n245 gnd 0.009219f
C1310 commonsourceibias.n246 gnd 0.009219f
C1311 commonsourceibias.n247 gnd 0.009219f
C1312 commonsourceibias.n248 gnd 0.010968f
C1313 commonsourceibias.n249 gnd 0.01272f
C1314 commonsourceibias.n250 gnd 0.068721f
C1315 commonsourceibias.n251 gnd 0.012643f
C1316 commonsourceibias.n252 gnd 0.009219f
C1317 commonsourceibias.n253 gnd 0.009219f
C1318 commonsourceibias.n254 gnd 0.009219f
C1319 commonsourceibias.n255 gnd 0.012488f
C1320 commonsourceibias.n256 gnd 0.068721f
C1321 commonsourceibias.n257 gnd 0.01257f
C1322 commonsourceibias.n258 gnd 0.011362f
C1323 commonsourceibias.n259 gnd 0.009219f
C1324 commonsourceibias.n260 gnd 0.009219f
C1325 commonsourceibias.n261 gnd 0.009352f
C1326 commonsourceibias.n262 gnd 0.009668f
C1327 commonsourceibias.t109 gnd 0.186271f
C1328 commonsourceibias.n263 gnd 0.082226f
C1329 commonsourceibias.n264 gnd 0.027982f
C1330 commonsourceibias.n265 gnd 0.437947f
C1331 commonsourceibias.n266 gnd 0.012301f
C1332 commonsourceibias.t69 gnd 0.186271f
C1333 commonsourceibias.t99 gnd 0.172234f
C1334 commonsourceibias.n267 gnd 0.068721f
C1335 commonsourceibias.n268 gnd 0.009219f
C1336 commonsourceibias.t84 gnd 0.172234f
C1337 commonsourceibias.n269 gnd 0.007457f
C1338 commonsourceibias.n270 gnd 0.009219f
C1339 commonsourceibias.t72 gnd 0.172234f
C1340 commonsourceibias.n271 gnd 0.0089f
C1341 commonsourceibias.n272 gnd 0.009219f
C1342 commonsourceibias.t66 gnd 0.172234f
C1343 commonsourceibias.n273 gnd 0.007446f
C1344 commonsourceibias.n274 gnd 0.009219f
C1345 commonsourceibias.t56 gnd 0.172234f
C1346 commonsourceibias.t79 gnd 0.172234f
C1347 commonsourceibias.n275 gnd 0.068721f
C1348 commonsourceibias.n276 gnd 0.009219f
C1349 commonsourceibias.t67 gnd 0.172234f
C1350 commonsourceibias.n277 gnd 0.068721f
C1351 commonsourceibias.n278 gnd 0.009219f
C1352 commonsourceibias.t104 gnd 0.172234f
C1353 commonsourceibias.n279 gnd 0.068721f
C1354 commonsourceibias.n280 gnd 0.046409f
C1355 commonsourceibias.t64 gnd 0.172234f
C1356 commonsourceibias.t111 gnd 0.194346f
C1357 commonsourceibias.n281 gnd 0.079751f
C1358 commonsourceibias.n282 gnd 0.082563f
C1359 commonsourceibias.n283 gnd 0.011362f
C1360 commonsourceibias.n284 gnd 0.01257f
C1361 commonsourceibias.n285 gnd 0.009219f
C1362 commonsourceibias.n286 gnd 0.009219f
C1363 commonsourceibias.n287 gnd 0.012488f
C1364 commonsourceibias.n288 gnd 0.007457f
C1365 commonsourceibias.n289 gnd 0.012643f
C1366 commonsourceibias.n290 gnd 0.009219f
C1367 commonsourceibias.n291 gnd 0.009219f
C1368 commonsourceibias.n292 gnd 0.01272f
C1369 commonsourceibias.n293 gnd 0.010968f
C1370 commonsourceibias.n294 gnd 0.0089f
C1371 commonsourceibias.n295 gnd 0.009219f
C1372 commonsourceibias.n296 gnd 0.009219f
C1373 commonsourceibias.n297 gnd 0.011276f
C1374 commonsourceibias.n298 gnd 0.012656f
C1375 commonsourceibias.n299 gnd 0.068721f
C1376 commonsourceibias.n300 gnd 0.012571f
C1377 commonsourceibias.n301 gnd 0.009174f
C1378 commonsourceibias.t5 gnd 0.019893f
C1379 commonsourceibias.t39 gnd 0.019893f
C1380 commonsourceibias.n302 gnd 0.17637f
C1381 commonsourceibias.t13 gnd 0.019893f
C1382 commonsourceibias.t37 gnd 0.019893f
C1383 commonsourceibias.n303 gnd 0.175781f
C1384 commonsourceibias.n304 gnd 0.163796f
C1385 commonsourceibias.t3 gnd 0.019893f
C1386 commonsourceibias.t45 gnd 0.019893f
C1387 commonsourceibias.n305 gnd 0.175781f
C1388 commonsourceibias.n306 gnd 0.067457f
C1389 commonsourceibias.n307 gnd 0.012301f
C1390 commonsourceibias.t8 gnd 0.172234f
C1391 commonsourceibias.n308 gnd 0.068721f
C1392 commonsourceibias.n309 gnd 0.009219f
C1393 commonsourceibias.t14 gnd 0.172234f
C1394 commonsourceibias.n310 gnd 0.007457f
C1395 commonsourceibias.n311 gnd 0.009219f
C1396 commonsourceibias.t32 gnd 0.172234f
C1397 commonsourceibias.n312 gnd 0.0089f
C1398 commonsourceibias.n313 gnd 0.009219f
C1399 commonsourceibias.t22 gnd 0.172234f
C1400 commonsourceibias.n314 gnd 0.007446f
C1401 commonsourceibias.n315 gnd 0.009219f
C1402 commonsourceibias.t44 gnd 0.172234f
C1403 commonsourceibias.t2 gnd 0.172234f
C1404 commonsourceibias.n316 gnd 0.068721f
C1405 commonsourceibias.n317 gnd 0.009219f
C1406 commonsourceibias.t36 gnd 0.172234f
C1407 commonsourceibias.n318 gnd 0.068721f
C1408 commonsourceibias.n319 gnd 0.009219f
C1409 commonsourceibias.t12 gnd 0.172234f
C1410 commonsourceibias.n320 gnd 0.068721f
C1411 commonsourceibias.n321 gnd 0.046409f
C1412 commonsourceibias.t38 gnd 0.172234f
C1413 commonsourceibias.t4 gnd 0.194346f
C1414 commonsourceibias.n322 gnd 0.079751f
C1415 commonsourceibias.n323 gnd 0.082563f
C1416 commonsourceibias.n324 gnd 0.011362f
C1417 commonsourceibias.n325 gnd 0.01257f
C1418 commonsourceibias.n326 gnd 0.009219f
C1419 commonsourceibias.n327 gnd 0.009219f
C1420 commonsourceibias.n328 gnd 0.012488f
C1421 commonsourceibias.n329 gnd 0.007457f
C1422 commonsourceibias.n330 gnd 0.012643f
C1423 commonsourceibias.n331 gnd 0.009219f
C1424 commonsourceibias.n332 gnd 0.009219f
C1425 commonsourceibias.n333 gnd 0.01272f
C1426 commonsourceibias.n334 gnd 0.010968f
C1427 commonsourceibias.n335 gnd 0.0089f
C1428 commonsourceibias.n336 gnd 0.009219f
C1429 commonsourceibias.n337 gnd 0.009219f
C1430 commonsourceibias.n338 gnd 0.011276f
C1431 commonsourceibias.n339 gnd 0.012656f
C1432 commonsourceibias.n340 gnd 0.068721f
C1433 commonsourceibias.n341 gnd 0.012571f
C1434 commonsourceibias.n342 gnd 0.009219f
C1435 commonsourceibias.n343 gnd 0.009219f
C1436 commonsourceibias.n344 gnd 0.009219f
C1437 commonsourceibias.n345 gnd 0.012571f
C1438 commonsourceibias.n346 gnd 0.068721f
C1439 commonsourceibias.n347 gnd 0.012656f
C1440 commonsourceibias.t18 gnd 0.172234f
C1441 commonsourceibias.n348 gnd 0.068721f
C1442 commonsourceibias.n349 gnd 0.011276f
C1443 commonsourceibias.n350 gnd 0.009219f
C1444 commonsourceibias.n351 gnd 0.009219f
C1445 commonsourceibias.n352 gnd 0.009219f
C1446 commonsourceibias.n353 gnd 0.010968f
C1447 commonsourceibias.n354 gnd 0.01272f
C1448 commonsourceibias.n355 gnd 0.068721f
C1449 commonsourceibias.n356 gnd 0.012643f
C1450 commonsourceibias.n357 gnd 0.009219f
C1451 commonsourceibias.n358 gnd 0.009219f
C1452 commonsourceibias.n359 gnd 0.009219f
C1453 commonsourceibias.n360 gnd 0.012488f
C1454 commonsourceibias.n361 gnd 0.068721f
C1455 commonsourceibias.n362 gnd 0.01257f
C1456 commonsourceibias.n363 gnd 0.011362f
C1457 commonsourceibias.n364 gnd 0.009219f
C1458 commonsourceibias.n365 gnd 0.009219f
C1459 commonsourceibias.n366 gnd 0.009352f
C1460 commonsourceibias.n367 gnd 0.009668f
C1461 commonsourceibias.t34 gnd 0.186271f
C1462 commonsourceibias.n368 gnd 0.082226f
C1463 commonsourceibias.n369 gnd 0.091217f
C1464 commonsourceibias.t9 gnd 0.019893f
C1465 commonsourceibias.t35 gnd 0.019893f
C1466 commonsourceibias.n370 gnd 0.175781f
C1467 commonsourceibias.n371 gnd 0.151888f
C1468 commonsourceibias.t33 gnd 0.019893f
C1469 commonsourceibias.t15 gnd 0.019893f
C1470 commonsourceibias.n372 gnd 0.175781f
C1471 commonsourceibias.n373 gnd 0.080743f
C1472 commonsourceibias.t23 gnd 0.019893f
C1473 commonsourceibias.t19 gnd 0.019893f
C1474 commonsourceibias.n374 gnd 0.175781f
C1475 commonsourceibias.n375 gnd 0.067457f
C1476 commonsourceibias.n376 gnd 0.081684f
C1477 commonsourceibias.n377 gnd 0.06664f
C1478 commonsourceibias.n378 gnd 0.009174f
C1479 commonsourceibias.n379 gnd 0.012571f
C1480 commonsourceibias.n380 gnd 0.068721f
C1481 commonsourceibias.n381 gnd 0.012656f
C1482 commonsourceibias.t92 gnd 0.172234f
C1483 commonsourceibias.n382 gnd 0.068721f
C1484 commonsourceibias.n383 gnd 0.011276f
C1485 commonsourceibias.n384 gnd 0.009219f
C1486 commonsourceibias.n385 gnd 0.009219f
C1487 commonsourceibias.n386 gnd 0.009219f
C1488 commonsourceibias.n387 gnd 0.010968f
C1489 commonsourceibias.n388 gnd 0.01272f
C1490 commonsourceibias.n389 gnd 0.068721f
C1491 commonsourceibias.n390 gnd 0.012643f
C1492 commonsourceibias.n391 gnd 0.009219f
C1493 commonsourceibias.n392 gnd 0.009219f
C1494 commonsourceibias.n393 gnd 0.009219f
C1495 commonsourceibias.n394 gnd 0.012488f
C1496 commonsourceibias.n395 gnd 0.068721f
C1497 commonsourceibias.n396 gnd 0.01257f
C1498 commonsourceibias.n397 gnd 0.011362f
C1499 commonsourceibias.n398 gnd 0.009219f
C1500 commonsourceibias.n399 gnd 0.009219f
C1501 commonsourceibias.n400 gnd 0.009352f
C1502 commonsourceibias.n401 gnd 0.009668f
C1503 commonsourceibias.n402 gnd 0.082226f
C1504 commonsourceibias.n403 gnd 0.053232f
C1505 commonsourceibias.n404 gnd 0.012301f
C1506 commonsourceibias.t107 gnd 0.172234f
C1507 commonsourceibias.n405 gnd 0.068721f
C1508 commonsourceibias.n406 gnd 0.009219f
C1509 commonsourceibias.t50 gnd 0.172234f
C1510 commonsourceibias.n407 gnd 0.007457f
C1511 commonsourceibias.n408 gnd 0.009219f
C1512 commonsourceibias.t114 gnd 0.172234f
C1513 commonsourceibias.n409 gnd 0.0089f
C1514 commonsourceibias.n410 gnd 0.009219f
C1515 commonsourceibias.t49 gnd 0.172234f
C1516 commonsourceibias.n411 gnd 0.007446f
C1517 commonsourceibias.n412 gnd 0.009219f
C1518 commonsourceibias.t74 gnd 0.172234f
C1519 commonsourceibias.t105 gnd 0.172234f
C1520 commonsourceibias.n413 gnd 0.068721f
C1521 commonsourceibias.n414 gnd 0.009219f
C1522 commonsourceibias.t55 gnd 0.172234f
C1523 commonsourceibias.n415 gnd 0.068721f
C1524 commonsourceibias.n416 gnd 0.009219f
C1525 commonsourceibias.t75 gnd 0.172234f
C1526 commonsourceibias.n417 gnd 0.068721f
C1527 commonsourceibias.n418 gnd 0.046409f
C1528 commonsourceibias.t61 gnd 0.172234f
C1529 commonsourceibias.t52 gnd 0.194346f
C1530 commonsourceibias.n419 gnd 0.079751f
C1531 commonsourceibias.n420 gnd 0.082563f
C1532 commonsourceibias.n421 gnd 0.011362f
C1533 commonsourceibias.n422 gnd 0.01257f
C1534 commonsourceibias.n423 gnd 0.009219f
C1535 commonsourceibias.n424 gnd 0.009219f
C1536 commonsourceibias.n425 gnd 0.012488f
C1537 commonsourceibias.n426 gnd 0.007457f
C1538 commonsourceibias.n427 gnd 0.012643f
C1539 commonsourceibias.n428 gnd 0.009219f
C1540 commonsourceibias.n429 gnd 0.009219f
C1541 commonsourceibias.n430 gnd 0.01272f
C1542 commonsourceibias.n431 gnd 0.010968f
C1543 commonsourceibias.n432 gnd 0.0089f
C1544 commonsourceibias.n433 gnd 0.009219f
C1545 commonsourceibias.n434 gnd 0.009219f
C1546 commonsourceibias.n435 gnd 0.011276f
C1547 commonsourceibias.n436 gnd 0.012656f
C1548 commonsourceibias.n437 gnd 0.068721f
C1549 commonsourceibias.n438 gnd 0.012571f
C1550 commonsourceibias.n439 gnd 0.009219f
C1551 commonsourceibias.n440 gnd 0.009219f
C1552 commonsourceibias.n441 gnd 0.009219f
C1553 commonsourceibias.n442 gnd 0.012571f
C1554 commonsourceibias.n443 gnd 0.068721f
C1555 commonsourceibias.n444 gnd 0.012656f
C1556 commonsourceibias.t106 gnd 0.172234f
C1557 commonsourceibias.n445 gnd 0.068721f
C1558 commonsourceibias.n446 gnd 0.011276f
C1559 commonsourceibias.n447 gnd 0.009219f
C1560 commonsourceibias.n448 gnd 0.009219f
C1561 commonsourceibias.n449 gnd 0.009219f
C1562 commonsourceibias.n450 gnd 0.010968f
C1563 commonsourceibias.n451 gnd 0.01272f
C1564 commonsourceibias.n452 gnd 0.068721f
C1565 commonsourceibias.n453 gnd 0.012643f
C1566 commonsourceibias.n454 gnd 0.009219f
C1567 commonsourceibias.n455 gnd 0.009219f
C1568 commonsourceibias.n456 gnd 0.009219f
C1569 commonsourceibias.n457 gnd 0.012488f
C1570 commonsourceibias.n458 gnd 0.068721f
C1571 commonsourceibias.n459 gnd 0.01257f
C1572 commonsourceibias.n460 gnd 0.011362f
C1573 commonsourceibias.n461 gnd 0.009219f
C1574 commonsourceibias.n462 gnd 0.009219f
C1575 commonsourceibias.n463 gnd 0.009352f
C1576 commonsourceibias.n464 gnd 0.009668f
C1577 commonsourceibias.t112 gnd 0.186271f
C1578 commonsourceibias.n465 gnd 0.082226f
C1579 commonsourceibias.n466 gnd 0.027982f
C1580 commonsourceibias.n467 gnd 0.147096f
C1581 commonsourceibias.n468 gnd 0.012301f
C1582 commonsourceibias.t81 gnd 0.172234f
C1583 commonsourceibias.n469 gnd 0.068721f
C1584 commonsourceibias.n470 gnd 0.009219f
C1585 commonsourceibias.t91 gnd 0.172234f
C1586 commonsourceibias.n471 gnd 0.007457f
C1587 commonsourceibias.n472 gnd 0.009219f
C1588 commonsourceibias.t100 gnd 0.172234f
C1589 commonsourceibias.n473 gnd 0.0089f
C1590 commonsourceibias.n474 gnd 0.009219f
C1591 commonsourceibias.t85 gnd 0.172234f
C1592 commonsourceibias.n475 gnd 0.007446f
C1593 commonsourceibias.n476 gnd 0.009219f
C1594 commonsourceibias.t82 gnd 0.172234f
C1595 commonsourceibias.t62 gnd 0.172234f
C1596 commonsourceibias.n477 gnd 0.068721f
C1597 commonsourceibias.n478 gnd 0.009219f
C1598 commonsourceibias.t53 gnd 0.172234f
C1599 commonsourceibias.n479 gnd 0.068721f
C1600 commonsourceibias.n480 gnd 0.009219f
C1601 commonsourceibias.t78 gnd 0.172234f
C1602 commonsourceibias.n481 gnd 0.068721f
C1603 commonsourceibias.n482 gnd 0.046409f
C1604 commonsourceibias.t97 gnd 0.172234f
C1605 commonsourceibias.t113 gnd 0.194346f
C1606 commonsourceibias.n483 gnd 0.079751f
C1607 commonsourceibias.n484 gnd 0.082563f
C1608 commonsourceibias.n485 gnd 0.011362f
C1609 commonsourceibias.n486 gnd 0.01257f
C1610 commonsourceibias.n487 gnd 0.009219f
C1611 commonsourceibias.n488 gnd 0.009219f
C1612 commonsourceibias.n489 gnd 0.012488f
C1613 commonsourceibias.n490 gnd 0.007457f
C1614 commonsourceibias.n491 gnd 0.012643f
C1615 commonsourceibias.n492 gnd 0.009219f
C1616 commonsourceibias.n493 gnd 0.009219f
C1617 commonsourceibias.n494 gnd 0.01272f
C1618 commonsourceibias.n495 gnd 0.010968f
C1619 commonsourceibias.n496 gnd 0.0089f
C1620 commonsourceibias.n497 gnd 0.009219f
C1621 commonsourceibias.n498 gnd 0.009219f
C1622 commonsourceibias.n499 gnd 0.011276f
C1623 commonsourceibias.n500 gnd 0.012656f
C1624 commonsourceibias.n501 gnd 0.068721f
C1625 commonsourceibias.n502 gnd 0.012571f
C1626 commonsourceibias.n503 gnd 0.009219f
C1627 commonsourceibias.n504 gnd 0.009219f
C1628 commonsourceibias.n505 gnd 0.009219f
C1629 commonsourceibias.n506 gnd 0.012571f
C1630 commonsourceibias.n507 gnd 0.068721f
C1631 commonsourceibias.n508 gnd 0.012656f
C1632 commonsourceibias.t76 gnd 0.172234f
C1633 commonsourceibias.n509 gnd 0.068721f
C1634 commonsourceibias.n510 gnd 0.011276f
C1635 commonsourceibias.n511 gnd 0.009219f
C1636 commonsourceibias.n512 gnd 0.009219f
C1637 commonsourceibias.n513 gnd 0.009219f
C1638 commonsourceibias.n514 gnd 0.010968f
C1639 commonsourceibias.n515 gnd 0.01272f
C1640 commonsourceibias.n516 gnd 0.068721f
C1641 commonsourceibias.n517 gnd 0.012643f
C1642 commonsourceibias.n518 gnd 0.009219f
C1643 commonsourceibias.n519 gnd 0.009219f
C1644 commonsourceibias.n520 gnd 0.009219f
C1645 commonsourceibias.n521 gnd 0.012488f
C1646 commonsourceibias.n522 gnd 0.068721f
C1647 commonsourceibias.n523 gnd 0.01257f
C1648 commonsourceibias.n524 gnd 0.011362f
C1649 commonsourceibias.n525 gnd 0.009219f
C1650 commonsourceibias.n526 gnd 0.009219f
C1651 commonsourceibias.n527 gnd 0.009352f
C1652 commonsourceibias.n528 gnd 0.009668f
C1653 commonsourceibias.t63 gnd 0.186271f
C1654 commonsourceibias.n529 gnd 0.082226f
C1655 commonsourceibias.n530 gnd 0.027982f
C1656 commonsourceibias.n531 gnd 0.194316f
C1657 commonsourceibias.n532 gnd 4.81454f
C1658 CSoutput.n0 gnd 0.049132f
C1659 CSoutput.t210 gnd 0.324994f
C1660 CSoutput.n1 gnd 0.146751f
C1661 CSoutput.n2 gnd 0.049132f
C1662 CSoutput.t195 gnd 0.324994f
C1663 CSoutput.n3 gnd 0.038941f
C1664 CSoutput.n4 gnd 0.049132f
C1665 CSoutput.t208 gnd 0.324994f
C1666 CSoutput.n5 gnd 0.033579f
C1667 CSoutput.n6 gnd 0.049132f
C1668 CSoutput.t212 gnd 0.324994f
C1669 CSoutput.t193 gnd 0.324994f
C1670 CSoutput.n7 gnd 0.145152f
C1671 CSoutput.n8 gnd 0.049132f
C1672 CSoutput.t203 gnd 0.324994f
C1673 CSoutput.n9 gnd 0.032016f
C1674 CSoutput.n10 gnd 0.049132f
C1675 CSoutput.t211 gnd 0.324994f
C1676 CSoutput.t209 gnd 0.324994f
C1677 CSoutput.n11 gnd 0.145152f
C1678 CSoutput.n12 gnd 0.049132f
C1679 CSoutput.t200 gnd 0.324994f
C1680 CSoutput.n13 gnd 0.033579f
C1681 CSoutput.n14 gnd 0.049132f
C1682 CSoutput.t198 gnd 0.324994f
C1683 CSoutput.t205 gnd 0.324994f
C1684 CSoutput.n15 gnd 0.145152f
C1685 CSoutput.n16 gnd 0.049132f
C1686 CSoutput.t192 gnd 0.324994f
C1687 CSoutput.n17 gnd 0.035864f
C1688 CSoutput.t202 gnd 0.388377f
C1689 CSoutput.t197 gnd 0.324994f
C1690 CSoutput.n18 gnd 0.185302f
C1691 CSoutput.n19 gnd 0.179807f
C1692 CSoutput.n20 gnd 0.208598f
C1693 CSoutput.n21 gnd 0.049132f
C1694 CSoutput.n22 gnd 0.041006f
C1695 CSoutput.n23 gnd 0.145152f
C1696 CSoutput.n24 gnd 0.039528f
C1697 CSoutput.n25 gnd 0.038941f
C1698 CSoutput.n26 gnd 0.049132f
C1699 CSoutput.n27 gnd 0.049132f
C1700 CSoutput.n28 gnd 0.04069f
C1701 CSoutput.n29 gnd 0.034547f
C1702 CSoutput.n30 gnd 0.148383f
C1703 CSoutput.n31 gnd 0.035023f
C1704 CSoutput.n32 gnd 0.049132f
C1705 CSoutput.n33 gnd 0.049132f
C1706 CSoutput.n34 gnd 0.049132f
C1707 CSoutput.n35 gnd 0.040257f
C1708 CSoutput.n36 gnd 0.145152f
C1709 CSoutput.n37 gnd 0.0385f
C1710 CSoutput.n38 gnd 0.039969f
C1711 CSoutput.n39 gnd 0.049132f
C1712 CSoutput.n40 gnd 0.049132f
C1713 CSoutput.n41 gnd 0.040997f
C1714 CSoutput.n42 gnd 0.037472f
C1715 CSoutput.n43 gnd 0.145152f
C1716 CSoutput.n44 gnd 0.038422f
C1717 CSoutput.n45 gnd 0.049132f
C1718 CSoutput.n46 gnd 0.049132f
C1719 CSoutput.n47 gnd 0.049132f
C1720 CSoutput.n48 gnd 0.038422f
C1721 CSoutput.n49 gnd 0.145152f
C1722 CSoutput.n50 gnd 0.037472f
C1723 CSoutput.n51 gnd 0.040997f
C1724 CSoutput.n52 gnd 0.049132f
C1725 CSoutput.n53 gnd 0.049132f
C1726 CSoutput.n54 gnd 0.039969f
C1727 CSoutput.n55 gnd 0.0385f
C1728 CSoutput.n56 gnd 0.145152f
C1729 CSoutput.n57 gnd 0.040257f
C1730 CSoutput.n58 gnd 0.049132f
C1731 CSoutput.n59 gnd 0.049132f
C1732 CSoutput.n60 gnd 0.049132f
C1733 CSoutput.n61 gnd 0.035023f
C1734 CSoutput.n62 gnd 0.148383f
C1735 CSoutput.n63 gnd 0.034547f
C1736 CSoutput.t201 gnd 0.324994f
C1737 CSoutput.n64 gnd 0.145152f
C1738 CSoutput.n65 gnd 0.04069f
C1739 CSoutput.n66 gnd 0.049132f
C1740 CSoutput.n67 gnd 0.049132f
C1741 CSoutput.n68 gnd 0.049132f
C1742 CSoutput.n69 gnd 0.039528f
C1743 CSoutput.n70 gnd 0.145152f
C1744 CSoutput.n71 gnd 0.041006f
C1745 CSoutput.n72 gnd 0.035864f
C1746 CSoutput.n73 gnd 0.049132f
C1747 CSoutput.n74 gnd 0.049132f
C1748 CSoutput.n75 gnd 0.037193f
C1749 CSoutput.n76 gnd 0.022089f
C1750 CSoutput.t204 gnd 0.365154f
C1751 CSoutput.n77 gnd 0.181394f
C1752 CSoutput.n78 gnd 0.742185f
C1753 CSoutput.t65 gnd 0.061285f
C1754 CSoutput.t123 gnd 0.061285f
C1755 CSoutput.n79 gnd 0.474486f
C1756 CSoutput.t72 gnd 0.061285f
C1757 CSoutput.t98 gnd 0.061285f
C1758 CSoutput.n80 gnd 0.47364f
C1759 CSoutput.n81 gnd 0.480744f
C1760 CSoutput.t177 gnd 0.061285f
C1761 CSoutput.t116 gnd 0.061285f
C1762 CSoutput.n82 gnd 0.47364f
C1763 CSoutput.n83 gnd 0.23689f
C1764 CSoutput.t74 gnd 0.061285f
C1765 CSoutput.t156 gnd 0.061285f
C1766 CSoutput.n84 gnd 0.47364f
C1767 CSoutput.n85 gnd 0.23689f
C1768 CSoutput.t81 gnd 0.061285f
C1769 CSoutput.t138 gnd 0.061285f
C1770 CSoutput.n86 gnd 0.47364f
C1771 CSoutput.n87 gnd 0.23689f
C1772 CSoutput.t103 gnd 0.061285f
C1773 CSoutput.t124 gnd 0.061285f
C1774 CSoutput.n88 gnd 0.47364f
C1775 CSoutput.n89 gnd 0.23689f
C1776 CSoutput.t119 gnd 0.061285f
C1777 CSoutput.t165 gnd 0.061285f
C1778 CSoutput.n90 gnd 0.47364f
C1779 CSoutput.n91 gnd 0.23689f
C1780 CSoutput.t91 gnd 0.061285f
C1781 CSoutput.t143 gnd 0.061285f
C1782 CSoutput.n92 gnd 0.47364f
C1783 CSoutput.n93 gnd 0.23689f
C1784 CSoutput.t112 gnd 0.061285f
C1785 CSoutput.t158 gnd 0.061285f
C1786 CSoutput.n94 gnd 0.47364f
C1787 CSoutput.n95 gnd 0.23689f
C1788 CSoutput.t128 gnd 0.061285f
C1789 CSoutput.t173 gnd 0.061285f
C1790 CSoutput.n96 gnd 0.47364f
C1791 CSoutput.n97 gnd 0.434402f
C1792 CSoutput.t86 gnd 0.061285f
C1793 CSoutput.t166 gnd 0.061285f
C1794 CSoutput.n98 gnd 0.474486f
C1795 CSoutput.t136 gnd 0.061285f
C1796 CSoutput.t134 gnd 0.061285f
C1797 CSoutput.n99 gnd 0.47364f
C1798 CSoutput.n100 gnd 0.480744f
C1799 CSoutput.t120 gnd 0.061285f
C1800 CSoutput.t83 gnd 0.061285f
C1801 CSoutput.n101 gnd 0.47364f
C1802 CSoutput.n102 gnd 0.23689f
C1803 CSoutput.t64 gnd 0.061285f
C1804 CSoutput.t122 gnd 0.061285f
C1805 CSoutput.n103 gnd 0.47364f
C1806 CSoutput.n104 gnd 0.23689f
C1807 CSoutput.t117 gnd 0.061285f
C1808 CSoutput.t80 gnd 0.061285f
C1809 CSoutput.n105 gnd 0.47364f
C1810 CSoutput.n106 gnd 0.23689f
C1811 CSoutput.t62 gnd 0.061285f
C1812 CSoutput.t60 gnd 0.061285f
C1813 CSoutput.n107 gnd 0.47364f
C1814 CSoutput.n108 gnd 0.23689f
C1815 CSoutput.t139 gnd 0.061285f
C1816 CSoutput.t99 gnd 0.061285f
C1817 CSoutput.n109 gnd 0.47364f
C1818 CSoutput.n110 gnd 0.23689f
C1819 CSoutput.t93 gnd 0.061285f
C1820 CSoutput.t59 gnd 0.061285f
C1821 CSoutput.n111 gnd 0.47364f
C1822 CSoutput.n112 gnd 0.23689f
C1823 CSoutput.t162 gnd 0.061285f
C1824 CSoutput.t135 gnd 0.061285f
C1825 CSoutput.n113 gnd 0.47364f
C1826 CSoutput.n114 gnd 0.23689f
C1827 CSoutput.t121 gnd 0.061285f
C1828 CSoutput.t84 gnd 0.061285f
C1829 CSoutput.n115 gnd 0.47364f
C1830 CSoutput.n116 gnd 0.353263f
C1831 CSoutput.n117 gnd 0.445463f
C1832 CSoutput.t104 gnd 0.061285f
C1833 CSoutput.t178 gnd 0.061285f
C1834 CSoutput.n118 gnd 0.474486f
C1835 CSoutput.t147 gnd 0.061285f
C1836 CSoutput.t145 gnd 0.061285f
C1837 CSoutput.n119 gnd 0.47364f
C1838 CSoutput.n120 gnd 0.480744f
C1839 CSoutput.t130 gnd 0.061285f
C1840 CSoutput.t100 gnd 0.061285f
C1841 CSoutput.n121 gnd 0.47364f
C1842 CSoutput.n122 gnd 0.23689f
C1843 CSoutput.t77 gnd 0.061285f
C1844 CSoutput.t132 gnd 0.061285f
C1845 CSoutput.n123 gnd 0.47364f
C1846 CSoutput.n124 gnd 0.23689f
C1847 CSoutput.t129 gnd 0.061285f
C1848 CSoutput.t97 gnd 0.061285f
C1849 CSoutput.n125 gnd 0.47364f
C1850 CSoutput.n126 gnd 0.23689f
C1851 CSoutput.t76 gnd 0.061285f
C1852 CSoutput.t75 gnd 0.061285f
C1853 CSoutput.n127 gnd 0.47364f
C1854 CSoutput.n128 gnd 0.23689f
C1855 CSoutput.t148 gnd 0.061285f
C1856 CSoutput.t113 gnd 0.061285f
C1857 CSoutput.n129 gnd 0.47364f
C1858 CSoutput.n130 gnd 0.23689f
C1859 CSoutput.t108 gnd 0.061285f
C1860 CSoutput.t71 gnd 0.061285f
C1861 CSoutput.n131 gnd 0.47364f
C1862 CSoutput.n132 gnd 0.23689f
C1863 CSoutput.t174 gnd 0.061285f
C1864 CSoutput.t146 gnd 0.061285f
C1865 CSoutput.n133 gnd 0.47364f
C1866 CSoutput.n134 gnd 0.23689f
C1867 CSoutput.t131 gnd 0.061285f
C1868 CSoutput.t101 gnd 0.061285f
C1869 CSoutput.n135 gnd 0.47364f
C1870 CSoutput.n136 gnd 0.353263f
C1871 CSoutput.n137 gnd 0.497913f
C1872 CSoutput.n138 gnd 9.07579f
C1873 CSoutput.n140 gnd 0.869128f
C1874 CSoutput.n141 gnd 0.651846f
C1875 CSoutput.n142 gnd 0.869128f
C1876 CSoutput.n143 gnd 0.869128f
C1877 CSoutput.n144 gnd 2.33996f
C1878 CSoutput.n145 gnd 0.869128f
C1879 CSoutput.n146 gnd 0.869128f
C1880 CSoutput.t199 gnd 1.08641f
C1881 CSoutput.n147 gnd 0.869128f
C1882 CSoutput.n148 gnd 0.869128f
C1883 CSoutput.n152 gnd 0.869128f
C1884 CSoutput.n156 gnd 0.869128f
C1885 CSoutput.n157 gnd 0.869128f
C1886 CSoutput.n159 gnd 0.869128f
C1887 CSoutput.n164 gnd 0.869128f
C1888 CSoutput.n166 gnd 0.869128f
C1889 CSoutput.n167 gnd 0.869128f
C1890 CSoutput.n169 gnd 0.869128f
C1891 CSoutput.n170 gnd 0.869128f
C1892 CSoutput.n172 gnd 0.869128f
C1893 CSoutput.t194 gnd 14.523f
C1894 CSoutput.n174 gnd 0.869128f
C1895 CSoutput.n175 gnd 0.651846f
C1896 CSoutput.n176 gnd 0.869128f
C1897 CSoutput.n177 gnd 0.869128f
C1898 CSoutput.n178 gnd 2.33996f
C1899 CSoutput.n179 gnd 0.869128f
C1900 CSoutput.n180 gnd 0.869128f
C1901 CSoutput.t206 gnd 1.08641f
C1902 CSoutput.n181 gnd 0.869128f
C1903 CSoutput.n182 gnd 0.869128f
C1904 CSoutput.n186 gnd 0.869128f
C1905 CSoutput.n190 gnd 0.869128f
C1906 CSoutput.n191 gnd 0.869128f
C1907 CSoutput.n193 gnd 0.869128f
C1908 CSoutput.n198 gnd 0.869128f
C1909 CSoutput.n200 gnd 0.869128f
C1910 CSoutput.n201 gnd 0.869128f
C1911 CSoutput.n203 gnd 0.869128f
C1912 CSoutput.n204 gnd 0.869128f
C1913 CSoutput.n206 gnd 0.869128f
C1914 CSoutput.n207 gnd 0.651846f
C1915 CSoutput.n209 gnd 0.869128f
C1916 CSoutput.n210 gnd 0.651846f
C1917 CSoutput.n211 gnd 0.869128f
C1918 CSoutput.n212 gnd 0.869128f
C1919 CSoutput.n213 gnd 2.33996f
C1920 CSoutput.n214 gnd 0.869128f
C1921 CSoutput.n215 gnd 0.869128f
C1922 CSoutput.t196 gnd 1.08641f
C1923 CSoutput.n216 gnd 0.869128f
C1924 CSoutput.n217 gnd 2.33996f
C1925 CSoutput.n219 gnd 0.869128f
C1926 CSoutput.n220 gnd 0.869128f
C1927 CSoutput.n222 gnd 0.869128f
C1928 CSoutput.n223 gnd 0.869128f
C1929 CSoutput.t207 gnd 14.2863f
C1930 CSoutput.t213 gnd 14.523f
C1931 CSoutput.n229 gnd 2.72658f
C1932 CSoutput.n230 gnd 11.1071f
C1933 CSoutput.n231 gnd 11.5719f
C1934 CSoutput.n236 gnd 2.95362f
C1935 CSoutput.n242 gnd 0.869128f
C1936 CSoutput.n244 gnd 0.869128f
C1937 CSoutput.n246 gnd 0.869128f
C1938 CSoutput.n248 gnd 0.869128f
C1939 CSoutput.n250 gnd 0.869128f
C1940 CSoutput.n256 gnd 0.869128f
C1941 CSoutput.n263 gnd 1.59452f
C1942 CSoutput.n264 gnd 1.59452f
C1943 CSoutput.n265 gnd 0.869128f
C1944 CSoutput.n266 gnd 0.869128f
C1945 CSoutput.n268 gnd 0.651846f
C1946 CSoutput.n269 gnd 0.558247f
C1947 CSoutput.n271 gnd 0.651846f
C1948 CSoutput.n272 gnd 0.558247f
C1949 CSoutput.n273 gnd 0.651846f
C1950 CSoutput.n275 gnd 0.869128f
C1951 CSoutput.n277 gnd 2.33996f
C1952 CSoutput.n278 gnd 2.72658f
C1953 CSoutput.n279 gnd 10.2157f
C1954 CSoutput.n281 gnd 0.651846f
C1955 CSoutput.n282 gnd 1.67724f
C1956 CSoutput.n283 gnd 0.651846f
C1957 CSoutput.n285 gnd 0.869128f
C1958 CSoutput.n287 gnd 2.33996f
C1959 CSoutput.n288 gnd 5.09735f
C1960 CSoutput.t149 gnd 0.061285f
C1961 CSoutput.t63 gnd 0.061285f
C1962 CSoutput.n289 gnd 0.474486f
C1963 CSoutput.t96 gnd 0.061285f
C1964 CSoutput.t70 gnd 0.061285f
C1965 CSoutput.n290 gnd 0.47364f
C1966 CSoutput.n291 gnd 0.480744f
C1967 CSoutput.t115 gnd 0.061285f
C1968 CSoutput.t90 gnd 0.061285f
C1969 CSoutput.n292 gnd 0.47364f
C1970 CSoutput.n293 gnd 0.23689f
C1971 CSoutput.t155 gnd 0.061285f
C1972 CSoutput.t73 gnd 0.061285f
C1973 CSoutput.n294 gnd 0.47364f
C1974 CSoutput.n295 gnd 0.23689f
C1975 CSoutput.t137 gnd 0.061285f
C1976 CSoutput.t78 gnd 0.061285f
C1977 CSoutput.n296 gnd 0.47364f
C1978 CSoutput.n297 gnd 0.23689f
C1979 CSoutput.t151 gnd 0.061285f
C1980 CSoutput.t102 gnd 0.061285f
C1981 CSoutput.n298 gnd 0.47364f
C1982 CSoutput.n299 gnd 0.23689f
C1983 CSoutput.t164 gnd 0.061285f
C1984 CSoutput.t118 gnd 0.061285f
C1985 CSoutput.n300 gnd 0.47364f
C1986 CSoutput.n301 gnd 0.23689f
C1987 CSoutput.t142 gnd 0.061285f
C1988 CSoutput.t92 gnd 0.061285f
C1989 CSoutput.n302 gnd 0.47364f
C1990 CSoutput.n303 gnd 0.23689f
C1991 CSoutput.t157 gnd 0.061285f
C1992 CSoutput.t110 gnd 0.061285f
C1993 CSoutput.n304 gnd 0.47364f
C1994 CSoutput.n305 gnd 0.23689f
C1995 CSoutput.t172 gnd 0.061285f
C1996 CSoutput.t126 gnd 0.061285f
C1997 CSoutput.n306 gnd 0.47364f
C1998 CSoutput.n307 gnd 0.434402f
C1999 CSoutput.t95 gnd 0.061285f
C2000 CSoutput.t163 gnd 0.061285f
C2001 CSoutput.n308 gnd 0.474486f
C2002 CSoutput.t87 gnd 0.061285f
C2003 CSoutput.t89 gnd 0.061285f
C2004 CSoutput.n309 gnd 0.47364f
C2005 CSoutput.n310 gnd 0.480744f
C2006 CSoutput.t160 gnd 0.061285f
C2007 CSoutput.t161 gnd 0.061285f
C2008 CSoutput.n311 gnd 0.47364f
C2009 CSoutput.n312 gnd 0.23689f
C2010 CSoutput.t69 gnd 0.061285f
C2011 CSoutput.t144 gnd 0.061285f
C2012 CSoutput.n313 gnd 0.47364f
C2013 CSoutput.n314 gnd 0.23689f
C2014 CSoutput.t154 gnd 0.061285f
C2015 CSoutput.t66 gnd 0.061285f
C2016 CSoutput.n315 gnd 0.47364f
C2017 CSoutput.n316 gnd 0.23689f
C2018 CSoutput.t114 gnd 0.061285f
C2019 CSoutput.t141 gnd 0.061285f
C2020 CSoutput.n317 gnd 0.47364f
C2021 CSoutput.n318 gnd 0.23689f
C2022 CSoutput.t168 gnd 0.061285f
C2023 CSoutput.t94 gnd 0.061285f
C2024 CSoutput.n319 gnd 0.47364f
C2025 CSoutput.n320 gnd 0.23689f
C2026 CSoutput.t140 gnd 0.061285f
C2027 CSoutput.t176 gnd 0.061285f
C2028 CSoutput.n321 gnd 0.47364f
C2029 CSoutput.n322 gnd 0.23689f
C2030 CSoutput.t88 gnd 0.061285f
C2031 CSoutput.t125 gnd 0.061285f
C2032 CSoutput.n323 gnd 0.47364f
C2033 CSoutput.n324 gnd 0.23689f
C2034 CSoutput.t159 gnd 0.061285f
C2035 CSoutput.t68 gnd 0.061285f
C2036 CSoutput.n325 gnd 0.47364f
C2037 CSoutput.n326 gnd 0.353263f
C2038 CSoutput.n327 gnd 0.445463f
C2039 CSoutput.t111 gnd 0.061285f
C2040 CSoutput.t175 gnd 0.061285f
C2041 CSoutput.n328 gnd 0.474486f
C2042 CSoutput.t105 gnd 0.061285f
C2043 CSoutput.t107 gnd 0.061285f
C2044 CSoutput.n329 gnd 0.47364f
C2045 CSoutput.n330 gnd 0.480744f
C2046 CSoutput.t169 gnd 0.061285f
C2047 CSoutput.t171 gnd 0.061285f
C2048 CSoutput.n331 gnd 0.47364f
C2049 CSoutput.n332 gnd 0.23689f
C2050 CSoutput.t85 gnd 0.061285f
C2051 CSoutput.t153 gnd 0.061285f
C2052 CSoutput.n333 gnd 0.47364f
C2053 CSoutput.n334 gnd 0.23689f
C2054 CSoutput.t167 gnd 0.061285f
C2055 CSoutput.t79 gnd 0.061285f
C2056 CSoutput.n335 gnd 0.47364f
C2057 CSoutput.n336 gnd 0.23689f
C2058 CSoutput.t127 gnd 0.061285f
C2059 CSoutput.t152 gnd 0.061285f
C2060 CSoutput.n337 gnd 0.47364f
C2061 CSoutput.n338 gnd 0.23689f
C2062 CSoutput.t61 gnd 0.061285f
C2063 CSoutput.t109 gnd 0.061285f
C2064 CSoutput.n339 gnd 0.47364f
C2065 CSoutput.n340 gnd 0.23689f
C2066 CSoutput.t150 gnd 0.061285f
C2067 CSoutput.t67 gnd 0.061285f
C2068 CSoutput.n341 gnd 0.47364f
C2069 CSoutput.n342 gnd 0.23689f
C2070 CSoutput.t106 gnd 0.061285f
C2071 CSoutput.t133 gnd 0.061285f
C2072 CSoutput.n343 gnd 0.47364f
C2073 CSoutput.n344 gnd 0.23689f
C2074 CSoutput.t170 gnd 0.061285f
C2075 CSoutput.t82 gnd 0.061285f
C2076 CSoutput.n345 gnd 0.473638f
C2077 CSoutput.n346 gnd 0.353265f
C2078 CSoutput.n347 gnd 0.497913f
C2079 CSoutput.n348 gnd 13.1652f
C2080 CSoutput.t38 gnd 0.053624f
C2081 CSoutput.t10 gnd 0.053624f
C2082 CSoutput.n349 gnd 0.475427f
C2083 CSoutput.t53 gnd 0.053624f
C2084 CSoutput.t39 gnd 0.053624f
C2085 CSoutput.n350 gnd 0.473841f
C2086 CSoutput.n351 gnd 0.441531f
C2087 CSoutput.t25 gnd 0.053624f
C2088 CSoutput.t34 gnd 0.053624f
C2089 CSoutput.n352 gnd 0.473841f
C2090 CSoutput.n353 gnd 0.217654f
C2091 CSoutput.t1 gnd 0.053624f
C2092 CSoutput.t52 gnd 0.053624f
C2093 CSoutput.n354 gnd 0.473841f
C2094 CSoutput.n355 gnd 0.217654f
C2095 CSoutput.t35 gnd 0.053624f
C2096 CSoutput.t36 gnd 0.053624f
C2097 CSoutput.n356 gnd 0.473841f
C2098 CSoutput.n357 gnd 0.217654f
C2099 CSoutput.t57 gnd 0.053624f
C2100 CSoutput.t12 gnd 0.053624f
C2101 CSoutput.n358 gnd 0.473841f
C2102 CSoutput.n359 gnd 0.401451f
C2103 CSoutput.t6 gnd 0.053624f
C2104 CSoutput.t47 gnd 0.053624f
C2105 CSoutput.n360 gnd 0.475427f
C2106 CSoutput.t14 gnd 0.053624f
C2107 CSoutput.t29 gnd 0.053624f
C2108 CSoutput.n361 gnd 0.473841f
C2109 CSoutput.n362 gnd 0.441531f
C2110 CSoutput.t187 gnd 0.053624f
C2111 CSoutput.t23 gnd 0.053624f
C2112 CSoutput.n363 gnd 0.473841f
C2113 CSoutput.n364 gnd 0.217654f
C2114 CSoutput.t183 gnd 0.053624f
C2115 CSoutput.t5 gnd 0.053624f
C2116 CSoutput.n365 gnd 0.473841f
C2117 CSoutput.n366 gnd 0.217654f
C2118 CSoutput.t22 gnd 0.053624f
C2119 CSoutput.t56 gnd 0.053624f
C2120 CSoutput.n367 gnd 0.473841f
C2121 CSoutput.n368 gnd 0.217654f
C2122 CSoutput.t189 gnd 0.053624f
C2123 CSoutput.t2 gnd 0.053624f
C2124 CSoutput.n369 gnd 0.473841f
C2125 CSoutput.n370 gnd 0.330446f
C2126 CSoutput.n371 gnd 0.416795f
C2127 CSoutput.t185 gnd 0.053624f
C2128 CSoutput.t0 gnd 0.053624f
C2129 CSoutput.n372 gnd 0.475427f
C2130 CSoutput.t9 gnd 0.053624f
C2131 CSoutput.t44 gnd 0.053624f
C2132 CSoutput.n373 gnd 0.473841f
C2133 CSoutput.n374 gnd 0.441531f
C2134 CSoutput.t188 gnd 0.053624f
C2135 CSoutput.t7 gnd 0.053624f
C2136 CSoutput.n375 gnd 0.473841f
C2137 CSoutput.n376 gnd 0.217654f
C2138 CSoutput.t37 gnd 0.053624f
C2139 CSoutput.t3 gnd 0.053624f
C2140 CSoutput.n377 gnd 0.473841f
C2141 CSoutput.n378 gnd 0.217654f
C2142 CSoutput.t26 gnd 0.053624f
C2143 CSoutput.t41 gnd 0.053624f
C2144 CSoutput.n379 gnd 0.473841f
C2145 CSoutput.n380 gnd 0.217654f
C2146 CSoutput.t28 gnd 0.053624f
C2147 CSoutput.t27 gnd 0.053624f
C2148 CSoutput.n381 gnd 0.473841f
C2149 CSoutput.n382 gnd 0.330446f
C2150 CSoutput.n383 gnd 0.447572f
C2151 CSoutput.n384 gnd 12.937201f
C2152 CSoutput.t49 gnd 0.053624f
C2153 CSoutput.t181 gnd 0.053624f
C2154 CSoutput.n385 gnd 0.475427f
C2155 CSoutput.t191 gnd 0.053624f
C2156 CSoutput.t32 gnd 0.053624f
C2157 CSoutput.n386 gnd 0.473841f
C2158 CSoutput.n387 gnd 0.441531f
C2159 CSoutput.t8 gnd 0.053624f
C2160 CSoutput.t43 gnd 0.053624f
C2161 CSoutput.n388 gnd 0.473841f
C2162 CSoutput.n389 gnd 0.217654f
C2163 CSoutput.t54 gnd 0.053624f
C2164 CSoutput.t184 gnd 0.053624f
C2165 CSoutput.n390 gnd 0.473841f
C2166 CSoutput.n391 gnd 0.217654f
C2167 CSoutput.t179 gnd 0.053624f
C2168 CSoutput.t48 gnd 0.053624f
C2169 CSoutput.n392 gnd 0.473841f
C2170 CSoutput.n393 gnd 0.217654f
C2171 CSoutput.t4 gnd 0.053624f
C2172 CSoutput.t11 gnd 0.053624f
C2173 CSoutput.n394 gnd 0.473841f
C2174 CSoutput.n395 gnd 0.401451f
C2175 CSoutput.t20 gnd 0.053624f
C2176 CSoutput.t186 gnd 0.053624f
C2177 CSoutput.n396 gnd 0.475427f
C2178 CSoutput.t30 gnd 0.053624f
C2179 CSoutput.t50 gnd 0.053624f
C2180 CSoutput.n397 gnd 0.473841f
C2181 CSoutput.n398 gnd 0.441531f
C2182 CSoutput.t51 gnd 0.053624f
C2183 CSoutput.t17 gnd 0.053624f
C2184 CSoutput.n399 gnd 0.473841f
C2185 CSoutput.n400 gnd 0.217654f
C2186 CSoutput.t180 gnd 0.053624f
C2187 CSoutput.t19 gnd 0.053624f
C2188 CSoutput.n401 gnd 0.473841f
C2189 CSoutput.n402 gnd 0.217654f
C2190 CSoutput.t190 gnd 0.053624f
C2191 CSoutput.t21 gnd 0.053624f
C2192 CSoutput.n403 gnd 0.473841f
C2193 CSoutput.n404 gnd 0.217654f
C2194 CSoutput.t182 gnd 0.053624f
C2195 CSoutput.t15 gnd 0.053624f
C2196 CSoutput.n405 gnd 0.473841f
C2197 CSoutput.n406 gnd 0.330446f
C2198 CSoutput.n407 gnd 0.416795f
C2199 CSoutput.t58 gnd 0.053624f
C2200 CSoutput.t31 gnd 0.053624f
C2201 CSoutput.n408 gnd 0.475427f
C2202 CSoutput.t24 gnd 0.053624f
C2203 CSoutput.t40 gnd 0.053624f
C2204 CSoutput.n409 gnd 0.473841f
C2205 CSoutput.n410 gnd 0.441531f
C2206 CSoutput.t33 gnd 0.053624f
C2207 CSoutput.t13 gnd 0.053624f
C2208 CSoutput.n411 gnd 0.473841f
C2209 CSoutput.n412 gnd 0.217654f
C2210 CSoutput.t42 gnd 0.053624f
C2211 CSoutput.t55 gnd 0.053624f
C2212 CSoutput.n413 gnd 0.473841f
C2213 CSoutput.n414 gnd 0.217654f
C2214 CSoutput.t16 gnd 0.053624f
C2215 CSoutput.t18 gnd 0.053624f
C2216 CSoutput.n415 gnd 0.473841f
C2217 CSoutput.n416 gnd 0.217654f
C2218 CSoutput.t46 gnd 0.053624f
C2219 CSoutput.t45 gnd 0.053624f
C2220 CSoutput.n417 gnd 0.473841f
C2221 CSoutput.n418 gnd 0.330446f
C2222 CSoutput.n419 gnd 0.447572f
C2223 CSoutput.n420 gnd 7.49367f
C2224 CSoutput.n421 gnd 14.7889f
C2225 vdd.t36 gnd 0.038214f
C2226 vdd.t23 gnd 0.038214f
C2227 vdd.n0 gnd 0.301396f
C2228 vdd.t48 gnd 0.038214f
C2229 vdd.t15 gnd 0.038214f
C2230 vdd.n1 gnd 0.300898f
C2231 vdd.n2 gnd 0.277486f
C2232 vdd.t4 gnd 0.038214f
C2233 vdd.t38 gnd 0.038214f
C2234 vdd.n3 gnd 0.300898f
C2235 vdd.n4 gnd 0.140335f
C2236 vdd.t40 gnd 0.038214f
C2237 vdd.t11 gnd 0.038214f
C2238 vdd.n5 gnd 0.300898f
C2239 vdd.n6 gnd 0.131678f
C2240 vdd.t50 gnd 0.038214f
C2241 vdd.t6 gnd 0.038214f
C2242 vdd.n7 gnd 0.301396f
C2243 vdd.t21 gnd 0.038214f
C2244 vdd.t34 gnd 0.038214f
C2245 vdd.n8 gnd 0.300898f
C2246 vdd.n9 gnd 0.277486f
C2247 vdd.t30 gnd 0.038214f
C2248 vdd.t303 gnd 0.038214f
C2249 vdd.n10 gnd 0.300898f
C2250 vdd.n11 gnd 0.140335f
C2251 vdd.t1 gnd 0.038214f
C2252 vdd.t32 gnd 0.038214f
C2253 vdd.n12 gnd 0.300898f
C2254 vdd.n13 gnd 0.131678f
C2255 vdd.n14 gnd 0.093094f
C2256 vdd.t51 gnd 0.02123f
C2257 vdd.t56 gnd 0.02123f
C2258 vdd.n15 gnd 0.19541f
C2259 vdd.t62 gnd 0.02123f
C2260 vdd.t27 gnd 0.02123f
C2261 vdd.n16 gnd 0.194839f
C2262 vdd.n17 gnd 0.33908f
C2263 vdd.t53 gnd 0.02123f
C2264 vdd.t300 gnd 0.02123f
C2265 vdd.n18 gnd 0.194839f
C2266 vdd.n19 gnd 0.140282f
C2267 vdd.t54 gnd 0.02123f
C2268 vdd.t28 gnd 0.02123f
C2269 vdd.n20 gnd 0.19541f
C2270 vdd.t58 gnd 0.02123f
C2271 vdd.t57 gnd 0.02123f
C2272 vdd.n21 gnd 0.194839f
C2273 vdd.n22 gnd 0.33908f
C2274 vdd.t60 gnd 0.02123f
C2275 vdd.t61 gnd 0.02123f
C2276 vdd.n23 gnd 0.194839f
C2277 vdd.n24 gnd 0.140282f
C2278 vdd.t301 gnd 0.02123f
C2279 vdd.t52 gnd 0.02123f
C2280 vdd.n25 gnd 0.194839f
C2281 vdd.t55 gnd 0.02123f
C2282 vdd.t59 gnd 0.02123f
C2283 vdd.n26 gnd 0.194839f
C2284 vdd.n27 gnd 21.2722f
C2285 vdd.n28 gnd 8.36097f
C2286 vdd.n29 gnd 0.00579f
C2287 vdd.n30 gnd 0.005373f
C2288 vdd.n31 gnd 0.002972f
C2289 vdd.n32 gnd 0.006824f
C2290 vdd.n33 gnd 0.002887f
C2291 vdd.n34 gnd 0.003057f
C2292 vdd.n35 gnd 0.005373f
C2293 vdd.n36 gnd 0.002887f
C2294 vdd.n37 gnd 0.006824f
C2295 vdd.n38 gnd 0.003057f
C2296 vdd.n39 gnd 0.005373f
C2297 vdd.n40 gnd 0.002887f
C2298 vdd.n41 gnd 0.005118f
C2299 vdd.n42 gnd 0.005134f
C2300 vdd.t268 gnd 0.014662f
C2301 vdd.n43 gnd 0.032622f
C2302 vdd.n44 gnd 0.169772f
C2303 vdd.n45 gnd 0.002887f
C2304 vdd.n46 gnd 0.003057f
C2305 vdd.n47 gnd 0.006824f
C2306 vdd.n48 gnd 0.006824f
C2307 vdd.n49 gnd 0.003057f
C2308 vdd.n50 gnd 0.002887f
C2309 vdd.n51 gnd 0.005373f
C2310 vdd.n52 gnd 0.005373f
C2311 vdd.n53 gnd 0.002887f
C2312 vdd.n54 gnd 0.003057f
C2313 vdd.n55 gnd 0.006824f
C2314 vdd.n56 gnd 0.006824f
C2315 vdd.n57 gnd 0.003057f
C2316 vdd.n58 gnd 0.002887f
C2317 vdd.n59 gnd 0.005373f
C2318 vdd.n60 gnd 0.005373f
C2319 vdd.n61 gnd 0.002887f
C2320 vdd.n62 gnd 0.003057f
C2321 vdd.n63 gnd 0.006824f
C2322 vdd.n64 gnd 0.006824f
C2323 vdd.n65 gnd 0.016134f
C2324 vdd.n66 gnd 0.002972f
C2325 vdd.n67 gnd 0.002887f
C2326 vdd.n68 gnd 0.013888f
C2327 vdd.n69 gnd 0.009696f
C2328 vdd.t153 gnd 0.033967f
C2329 vdd.t200 gnd 0.033967f
C2330 vdd.n70 gnd 0.233448f
C2331 vdd.n71 gnd 0.183571f
C2332 vdd.t164 gnd 0.033967f
C2333 vdd.t226 gnd 0.033967f
C2334 vdd.n72 gnd 0.233448f
C2335 vdd.n73 gnd 0.148141f
C2336 vdd.t191 gnd 0.033967f
C2337 vdd.t274 gnd 0.033967f
C2338 vdd.n74 gnd 0.233448f
C2339 vdd.n75 gnd 0.148141f
C2340 vdd.t169 gnd 0.033967f
C2341 vdd.t255 gnd 0.033967f
C2342 vdd.n76 gnd 0.233448f
C2343 vdd.n77 gnd 0.148141f
C2344 vdd.t173 gnd 0.033967f
C2345 vdd.t270 gnd 0.033967f
C2346 vdd.n78 gnd 0.233448f
C2347 vdd.n79 gnd 0.148141f
C2348 vdd.t209 gnd 0.033967f
C2349 vdd.t285 gnd 0.033967f
C2350 vdd.n80 gnd 0.233448f
C2351 vdd.n81 gnd 0.148141f
C2352 vdd.t229 gnd 0.033967f
C2353 vdd.t261 gnd 0.033967f
C2354 vdd.n82 gnd 0.233448f
C2355 vdd.n83 gnd 0.148141f
C2356 vdd.t194 gnd 0.033967f
C2357 vdd.t276 gnd 0.033967f
C2358 vdd.n84 gnd 0.233448f
C2359 vdd.n85 gnd 0.148141f
C2360 vdd.t218 gnd 0.033967f
C2361 vdd.t292 gnd 0.033967f
C2362 vdd.n86 gnd 0.233448f
C2363 vdd.n87 gnd 0.148141f
C2364 vdd.n88 gnd 0.00579f
C2365 vdd.n89 gnd 0.005373f
C2366 vdd.n90 gnd 0.002972f
C2367 vdd.n91 gnd 0.006824f
C2368 vdd.n92 gnd 0.002887f
C2369 vdd.n93 gnd 0.003057f
C2370 vdd.n94 gnd 0.005373f
C2371 vdd.n95 gnd 0.002887f
C2372 vdd.n96 gnd 0.006824f
C2373 vdd.n97 gnd 0.003057f
C2374 vdd.n98 gnd 0.005373f
C2375 vdd.n99 gnd 0.002887f
C2376 vdd.n100 gnd 0.005118f
C2377 vdd.n101 gnd 0.005134f
C2378 vdd.t244 gnd 0.014662f
C2379 vdd.n102 gnd 0.032622f
C2380 vdd.n103 gnd 0.169772f
C2381 vdd.n104 gnd 0.002887f
C2382 vdd.n105 gnd 0.003057f
C2383 vdd.n106 gnd 0.006824f
C2384 vdd.n107 gnd 0.006824f
C2385 vdd.n108 gnd 0.003057f
C2386 vdd.n109 gnd 0.002887f
C2387 vdd.n110 gnd 0.005373f
C2388 vdd.n111 gnd 0.005373f
C2389 vdd.n112 gnd 0.002887f
C2390 vdd.n113 gnd 0.003057f
C2391 vdd.n114 gnd 0.006824f
C2392 vdd.n115 gnd 0.006824f
C2393 vdd.n116 gnd 0.003057f
C2394 vdd.n117 gnd 0.002887f
C2395 vdd.n118 gnd 0.005373f
C2396 vdd.n119 gnd 0.005373f
C2397 vdd.n120 gnd 0.002887f
C2398 vdd.n121 gnd 0.003057f
C2399 vdd.n122 gnd 0.006824f
C2400 vdd.n123 gnd 0.006824f
C2401 vdd.n124 gnd 0.016134f
C2402 vdd.n125 gnd 0.002972f
C2403 vdd.n126 gnd 0.002887f
C2404 vdd.n127 gnd 0.013888f
C2405 vdd.n128 gnd 0.009391f
C2406 vdd.n129 gnd 0.110218f
C2407 vdd.n130 gnd 0.00579f
C2408 vdd.n131 gnd 0.005373f
C2409 vdd.n132 gnd 0.002972f
C2410 vdd.n133 gnd 0.006824f
C2411 vdd.n134 gnd 0.002887f
C2412 vdd.n135 gnd 0.003057f
C2413 vdd.n136 gnd 0.005373f
C2414 vdd.n137 gnd 0.002887f
C2415 vdd.n138 gnd 0.006824f
C2416 vdd.n139 gnd 0.003057f
C2417 vdd.n140 gnd 0.005373f
C2418 vdd.n141 gnd 0.002887f
C2419 vdd.n142 gnd 0.005118f
C2420 vdd.n143 gnd 0.005134f
C2421 vdd.t199 gnd 0.014662f
C2422 vdd.n144 gnd 0.032622f
C2423 vdd.n145 gnd 0.169772f
C2424 vdd.n146 gnd 0.002887f
C2425 vdd.n147 gnd 0.003057f
C2426 vdd.n148 gnd 0.006824f
C2427 vdd.n149 gnd 0.006824f
C2428 vdd.n150 gnd 0.003057f
C2429 vdd.n151 gnd 0.002887f
C2430 vdd.n152 gnd 0.005373f
C2431 vdd.n153 gnd 0.005373f
C2432 vdd.n154 gnd 0.002887f
C2433 vdd.n155 gnd 0.003057f
C2434 vdd.n156 gnd 0.006824f
C2435 vdd.n157 gnd 0.006824f
C2436 vdd.n158 gnd 0.003057f
C2437 vdd.n159 gnd 0.002887f
C2438 vdd.n160 gnd 0.005373f
C2439 vdd.n161 gnd 0.005373f
C2440 vdd.n162 gnd 0.002887f
C2441 vdd.n163 gnd 0.003057f
C2442 vdd.n164 gnd 0.006824f
C2443 vdd.n165 gnd 0.006824f
C2444 vdd.n166 gnd 0.016134f
C2445 vdd.n167 gnd 0.002972f
C2446 vdd.n168 gnd 0.002887f
C2447 vdd.n169 gnd 0.013888f
C2448 vdd.n170 gnd 0.009696f
C2449 vdd.t284 gnd 0.033967f
C2450 vdd.t186 gnd 0.033967f
C2451 vdd.n171 gnd 0.233448f
C2452 vdd.n172 gnd 0.183571f
C2453 vdd.t189 gnd 0.033967f
C2454 vdd.t280 gnd 0.033967f
C2455 vdd.n173 gnd 0.233448f
C2456 vdd.n174 gnd 0.148141f
C2457 vdd.t281 gnd 0.033967f
C2458 vdd.t162 gnd 0.033967f
C2459 vdd.n175 gnd 0.233448f
C2460 vdd.n176 gnd 0.148141f
C2461 vdd.t263 gnd 0.033967f
C2462 vdd.t273 gnd 0.033967f
C2463 vdd.n177 gnd 0.233448f
C2464 vdd.n178 gnd 0.148141f
C2465 vdd.t158 gnd 0.033967f
C2466 vdd.t224 gnd 0.033967f
C2467 vdd.n179 gnd 0.233448f
C2468 vdd.n180 gnd 0.148141f
C2469 vdd.t260 gnd 0.033967f
C2470 vdd.t288 gnd 0.033967f
C2471 vdd.n181 gnd 0.233448f
C2472 vdd.n182 gnd 0.148141f
C2473 vdd.t197 gnd 0.033967f
C2474 vdd.t259 gnd 0.033967f
C2475 vdd.n183 gnd 0.233448f
C2476 vdd.n184 gnd 0.148141f
C2477 vdd.t296 gnd 0.033967f
C2478 vdd.t188 gnd 0.033967f
C2479 vdd.n185 gnd 0.233448f
C2480 vdd.n186 gnd 0.148141f
C2481 vdd.t243 gnd 0.033967f
C2482 vdd.t279 gnd 0.033967f
C2483 vdd.n187 gnd 0.233448f
C2484 vdd.n188 gnd 0.148141f
C2485 vdd.n189 gnd 0.00579f
C2486 vdd.n190 gnd 0.005373f
C2487 vdd.n191 gnd 0.002972f
C2488 vdd.n192 gnd 0.006824f
C2489 vdd.n193 gnd 0.002887f
C2490 vdd.n194 gnd 0.003057f
C2491 vdd.n195 gnd 0.005373f
C2492 vdd.n196 gnd 0.002887f
C2493 vdd.n197 gnd 0.006824f
C2494 vdd.n198 gnd 0.003057f
C2495 vdd.n199 gnd 0.005373f
C2496 vdd.n200 gnd 0.002887f
C2497 vdd.n201 gnd 0.005118f
C2498 vdd.n202 gnd 0.005134f
C2499 vdd.t145 gnd 0.014662f
C2500 vdd.n203 gnd 0.032622f
C2501 vdd.n204 gnd 0.169772f
C2502 vdd.n205 gnd 0.002887f
C2503 vdd.n206 gnd 0.003057f
C2504 vdd.n207 gnd 0.006824f
C2505 vdd.n208 gnd 0.006824f
C2506 vdd.n209 gnd 0.003057f
C2507 vdd.n210 gnd 0.002887f
C2508 vdd.n211 gnd 0.005373f
C2509 vdd.n212 gnd 0.005373f
C2510 vdd.n213 gnd 0.002887f
C2511 vdd.n214 gnd 0.003057f
C2512 vdd.n215 gnd 0.006824f
C2513 vdd.n216 gnd 0.006824f
C2514 vdd.n217 gnd 0.003057f
C2515 vdd.n218 gnd 0.002887f
C2516 vdd.n219 gnd 0.005373f
C2517 vdd.n220 gnd 0.005373f
C2518 vdd.n221 gnd 0.002887f
C2519 vdd.n222 gnd 0.003057f
C2520 vdd.n223 gnd 0.006824f
C2521 vdd.n224 gnd 0.006824f
C2522 vdd.n225 gnd 0.016134f
C2523 vdd.n226 gnd 0.002972f
C2524 vdd.n227 gnd 0.002887f
C2525 vdd.n228 gnd 0.013888f
C2526 vdd.n229 gnd 0.009391f
C2527 vdd.n230 gnd 0.065568f
C2528 vdd.n231 gnd 0.23626f
C2529 vdd.n232 gnd 0.00579f
C2530 vdd.n233 gnd 0.005373f
C2531 vdd.n234 gnd 0.002972f
C2532 vdd.n235 gnd 0.006824f
C2533 vdd.n236 gnd 0.002887f
C2534 vdd.n237 gnd 0.003057f
C2535 vdd.n238 gnd 0.005373f
C2536 vdd.n239 gnd 0.002887f
C2537 vdd.n240 gnd 0.006824f
C2538 vdd.n241 gnd 0.003057f
C2539 vdd.n242 gnd 0.005373f
C2540 vdd.n243 gnd 0.002887f
C2541 vdd.n244 gnd 0.005118f
C2542 vdd.n245 gnd 0.005134f
C2543 vdd.t219 gnd 0.014662f
C2544 vdd.n246 gnd 0.032622f
C2545 vdd.n247 gnd 0.169772f
C2546 vdd.n248 gnd 0.002887f
C2547 vdd.n249 gnd 0.003057f
C2548 vdd.n250 gnd 0.006824f
C2549 vdd.n251 gnd 0.006824f
C2550 vdd.n252 gnd 0.003057f
C2551 vdd.n253 gnd 0.002887f
C2552 vdd.n254 gnd 0.005373f
C2553 vdd.n255 gnd 0.005373f
C2554 vdd.n256 gnd 0.002887f
C2555 vdd.n257 gnd 0.003057f
C2556 vdd.n258 gnd 0.006824f
C2557 vdd.n259 gnd 0.006824f
C2558 vdd.n260 gnd 0.003057f
C2559 vdd.n261 gnd 0.002887f
C2560 vdd.n262 gnd 0.005373f
C2561 vdd.n263 gnd 0.005373f
C2562 vdd.n264 gnd 0.002887f
C2563 vdd.n265 gnd 0.003057f
C2564 vdd.n266 gnd 0.006824f
C2565 vdd.n267 gnd 0.006824f
C2566 vdd.n268 gnd 0.016134f
C2567 vdd.n269 gnd 0.002972f
C2568 vdd.n270 gnd 0.002887f
C2569 vdd.n271 gnd 0.013888f
C2570 vdd.n272 gnd 0.009696f
C2571 vdd.t295 gnd 0.033967f
C2572 vdd.t212 gnd 0.033967f
C2573 vdd.n273 gnd 0.233448f
C2574 vdd.n274 gnd 0.183571f
C2575 vdd.t214 gnd 0.033967f
C2576 vdd.t289 gnd 0.033967f
C2577 vdd.n275 gnd 0.233448f
C2578 vdd.n276 gnd 0.148141f
C2579 vdd.t290 gnd 0.033967f
C2580 vdd.t183 gnd 0.033967f
C2581 vdd.n277 gnd 0.233448f
C2582 vdd.n278 gnd 0.148141f
C2583 vdd.t272 gnd 0.033967f
C2584 vdd.t287 gnd 0.033967f
C2585 vdd.n279 gnd 0.233448f
C2586 vdd.n280 gnd 0.148141f
C2587 vdd.t174 gnd 0.033967f
C2588 vdd.t245 gnd 0.033967f
C2589 vdd.n281 gnd 0.233448f
C2590 vdd.n282 gnd 0.148141f
C2591 vdd.t271 gnd 0.033967f
C2592 vdd.t151 gnd 0.033967f
C2593 vdd.n283 gnd 0.233448f
C2594 vdd.n284 gnd 0.148141f
C2595 vdd.t216 gnd 0.033967f
C2596 vdd.t269 gnd 0.033967f
C2597 vdd.n285 gnd 0.233448f
C2598 vdd.n286 gnd 0.148141f
C2599 vdd.t160 gnd 0.033967f
C2600 vdd.t213 gnd 0.033967f
C2601 vdd.n287 gnd 0.233448f
C2602 vdd.n288 gnd 0.148141f
C2603 vdd.t251 gnd 0.033967f
C2604 vdd.t291 gnd 0.033967f
C2605 vdd.n289 gnd 0.233448f
C2606 vdd.n290 gnd 0.148141f
C2607 vdd.n291 gnd 0.00579f
C2608 vdd.n292 gnd 0.005373f
C2609 vdd.n293 gnd 0.002972f
C2610 vdd.n294 gnd 0.006824f
C2611 vdd.n295 gnd 0.002887f
C2612 vdd.n296 gnd 0.003057f
C2613 vdd.n297 gnd 0.005373f
C2614 vdd.n298 gnd 0.002887f
C2615 vdd.n299 gnd 0.006824f
C2616 vdd.n300 gnd 0.003057f
C2617 vdd.n301 gnd 0.005373f
C2618 vdd.n302 gnd 0.002887f
C2619 vdd.n303 gnd 0.005118f
C2620 vdd.n304 gnd 0.005134f
C2621 vdd.t142 gnd 0.014662f
C2622 vdd.n305 gnd 0.032622f
C2623 vdd.n306 gnd 0.169772f
C2624 vdd.n307 gnd 0.002887f
C2625 vdd.n308 gnd 0.003057f
C2626 vdd.n309 gnd 0.006824f
C2627 vdd.n310 gnd 0.006824f
C2628 vdd.n311 gnd 0.003057f
C2629 vdd.n312 gnd 0.002887f
C2630 vdd.n313 gnd 0.005373f
C2631 vdd.n314 gnd 0.005373f
C2632 vdd.n315 gnd 0.002887f
C2633 vdd.n316 gnd 0.003057f
C2634 vdd.n317 gnd 0.006824f
C2635 vdd.n318 gnd 0.006824f
C2636 vdd.n319 gnd 0.003057f
C2637 vdd.n320 gnd 0.002887f
C2638 vdd.n321 gnd 0.005373f
C2639 vdd.n322 gnd 0.005373f
C2640 vdd.n323 gnd 0.002887f
C2641 vdd.n324 gnd 0.003057f
C2642 vdd.n325 gnd 0.006824f
C2643 vdd.n326 gnd 0.006824f
C2644 vdd.n327 gnd 0.016134f
C2645 vdd.n328 gnd 0.002972f
C2646 vdd.n329 gnd 0.002887f
C2647 vdd.n330 gnd 0.013888f
C2648 vdd.n331 gnd 0.009391f
C2649 vdd.n332 gnd 0.065568f
C2650 vdd.n333 gnd 0.270467f
C2651 vdd.n334 gnd 0.008109f
C2652 vdd.n335 gnd 0.01055f
C2653 vdd.n336 gnd 0.008492f
C2654 vdd.n337 gnd 0.008492f
C2655 vdd.n338 gnd 0.01055f
C2656 vdd.n339 gnd 0.01055f
C2657 vdd.n340 gnd 0.770922f
C2658 vdd.n341 gnd 0.01055f
C2659 vdd.n342 gnd 0.01055f
C2660 vdd.n343 gnd 0.01055f
C2661 vdd.n344 gnd 0.835614f
C2662 vdd.n345 gnd 0.01055f
C2663 vdd.n346 gnd 0.01055f
C2664 vdd.n347 gnd 0.01055f
C2665 vdd.n348 gnd 0.01055f
C2666 vdd.n349 gnd 0.008492f
C2667 vdd.n350 gnd 0.01055f
C2668 vdd.t150 gnd 0.539106f
C2669 vdd.n351 gnd 0.01055f
C2670 vdd.n352 gnd 0.01055f
C2671 vdd.n353 gnd 0.01055f
C2672 vdd.t258 gnd 0.539106f
C2673 vdd.n354 gnd 0.01055f
C2674 vdd.n355 gnd 0.01055f
C2675 vdd.n356 gnd 0.01055f
C2676 vdd.n357 gnd 0.01055f
C2677 vdd.n358 gnd 0.01055f
C2678 vdd.n359 gnd 0.008492f
C2679 vdd.n360 gnd 0.01055f
C2680 vdd.n361 gnd 0.60919f
C2681 vdd.n362 gnd 0.01055f
C2682 vdd.n363 gnd 0.01055f
C2683 vdd.n364 gnd 0.01055f
C2684 vdd.t187 gnd 0.539106f
C2685 vdd.n365 gnd 0.01055f
C2686 vdd.n366 gnd 0.01055f
C2687 vdd.n367 gnd 0.01055f
C2688 vdd.n368 gnd 0.01055f
C2689 vdd.n369 gnd 0.01055f
C2690 vdd.n370 gnd 0.008492f
C2691 vdd.n371 gnd 0.01055f
C2692 vdd.t217 gnd 0.539106f
C2693 vdd.n372 gnd 0.01055f
C2694 vdd.n373 gnd 0.01055f
C2695 vdd.n374 gnd 0.01055f
C2696 vdd.n375 gnd 0.630754f
C2697 vdd.n376 gnd 0.01055f
C2698 vdd.n377 gnd 0.01055f
C2699 vdd.n378 gnd 0.01055f
C2700 vdd.n379 gnd 0.01055f
C2701 vdd.n380 gnd 0.01055f
C2702 vdd.n381 gnd 0.008492f
C2703 vdd.n382 gnd 0.01055f
C2704 vdd.t141 gnd 0.539106f
C2705 vdd.n383 gnd 0.01055f
C2706 vdd.n384 gnd 0.01055f
C2707 vdd.n385 gnd 0.01055f
C2708 vdd.n386 gnd 0.544497f
C2709 vdd.n387 gnd 0.01055f
C2710 vdd.n388 gnd 0.01055f
C2711 vdd.n389 gnd 0.01055f
C2712 vdd.n390 gnd 0.01055f
C2713 vdd.n391 gnd 0.025523f
C2714 vdd.n392 gnd 0.026069f
C2715 vdd.t76 gnd 0.539106f
C2716 vdd.n393 gnd 0.025523f
C2717 vdd.n425 gnd 0.01055f
C2718 vdd.t104 gnd 0.129799f
C2719 vdd.t103 gnd 0.138719f
C2720 vdd.t102 gnd 0.169516f
C2721 vdd.n426 gnd 0.217295f
C2722 vdd.n427 gnd 0.183417f
C2723 vdd.n428 gnd 0.013927f
C2724 vdd.n429 gnd 0.01055f
C2725 vdd.n430 gnd 0.008492f
C2726 vdd.n431 gnd 0.01055f
C2727 vdd.n432 gnd 0.008492f
C2728 vdd.n433 gnd 0.01055f
C2729 vdd.n434 gnd 0.008492f
C2730 vdd.n435 gnd 0.01055f
C2731 vdd.n436 gnd 0.008492f
C2732 vdd.n437 gnd 0.01055f
C2733 vdd.n438 gnd 0.008492f
C2734 vdd.n439 gnd 0.01055f
C2735 vdd.t78 gnd 0.129799f
C2736 vdd.t77 gnd 0.138719f
C2737 vdd.t75 gnd 0.169516f
C2738 vdd.n440 gnd 0.217295f
C2739 vdd.n441 gnd 0.183417f
C2740 vdd.n442 gnd 0.008492f
C2741 vdd.n443 gnd 0.01055f
C2742 vdd.n444 gnd 0.008492f
C2743 vdd.n445 gnd 0.01055f
C2744 vdd.n446 gnd 0.008492f
C2745 vdd.n447 gnd 0.01055f
C2746 vdd.n448 gnd 0.008492f
C2747 vdd.n449 gnd 0.01055f
C2748 vdd.n450 gnd 0.008492f
C2749 vdd.n451 gnd 0.01055f
C2750 vdd.t95 gnd 0.129799f
C2751 vdd.t94 gnd 0.138719f
C2752 vdd.t93 gnd 0.169516f
C2753 vdd.n452 gnd 0.217295f
C2754 vdd.n453 gnd 0.183417f
C2755 vdd.n454 gnd 0.018173f
C2756 vdd.n455 gnd 0.01055f
C2757 vdd.n456 gnd 0.008492f
C2758 vdd.n457 gnd 0.01055f
C2759 vdd.n458 gnd 0.008492f
C2760 vdd.n459 gnd 0.01055f
C2761 vdd.n460 gnd 0.008492f
C2762 vdd.n461 gnd 0.01055f
C2763 vdd.n462 gnd 0.008492f
C2764 vdd.n463 gnd 0.01055f
C2765 vdd.n464 gnd 0.026069f
C2766 vdd.n465 gnd 0.007048f
C2767 vdd.n466 gnd 0.008492f
C2768 vdd.n467 gnd 0.01055f
C2769 vdd.n468 gnd 0.01055f
C2770 vdd.n469 gnd 0.008492f
C2771 vdd.n470 gnd 0.01055f
C2772 vdd.n471 gnd 0.01055f
C2773 vdd.n472 gnd 0.01055f
C2774 vdd.n473 gnd 0.01055f
C2775 vdd.n474 gnd 0.01055f
C2776 vdd.n475 gnd 0.008492f
C2777 vdd.n476 gnd 0.008492f
C2778 vdd.n477 gnd 0.01055f
C2779 vdd.n478 gnd 0.01055f
C2780 vdd.n479 gnd 0.008492f
C2781 vdd.n480 gnd 0.01055f
C2782 vdd.n481 gnd 0.01055f
C2783 vdd.n482 gnd 0.01055f
C2784 vdd.n483 gnd 0.01055f
C2785 vdd.n484 gnd 0.01055f
C2786 vdd.n485 gnd 0.008492f
C2787 vdd.n486 gnd 0.008492f
C2788 vdd.n487 gnd 0.01055f
C2789 vdd.n488 gnd 0.01055f
C2790 vdd.n489 gnd 0.008492f
C2791 vdd.n490 gnd 0.01055f
C2792 vdd.n491 gnd 0.01055f
C2793 vdd.n492 gnd 0.01055f
C2794 vdd.n493 gnd 0.01055f
C2795 vdd.n494 gnd 0.01055f
C2796 vdd.n495 gnd 0.008492f
C2797 vdd.n496 gnd 0.008492f
C2798 vdd.n497 gnd 0.01055f
C2799 vdd.n498 gnd 0.01055f
C2800 vdd.n499 gnd 0.008492f
C2801 vdd.n500 gnd 0.01055f
C2802 vdd.n501 gnd 0.01055f
C2803 vdd.n502 gnd 0.01055f
C2804 vdd.n503 gnd 0.01055f
C2805 vdd.n504 gnd 0.01055f
C2806 vdd.n505 gnd 0.008492f
C2807 vdd.n506 gnd 0.008492f
C2808 vdd.n507 gnd 0.01055f
C2809 vdd.n508 gnd 0.01055f
C2810 vdd.n509 gnd 0.007091f
C2811 vdd.n510 gnd 0.01055f
C2812 vdd.n511 gnd 0.01055f
C2813 vdd.n512 gnd 0.01055f
C2814 vdd.n513 gnd 0.01055f
C2815 vdd.n514 gnd 0.01055f
C2816 vdd.n515 gnd 0.007091f
C2817 vdd.n516 gnd 0.008492f
C2818 vdd.n517 gnd 0.01055f
C2819 vdd.n518 gnd 0.01055f
C2820 vdd.n519 gnd 0.008492f
C2821 vdd.n520 gnd 0.01055f
C2822 vdd.n521 gnd 0.01055f
C2823 vdd.n522 gnd 0.01055f
C2824 vdd.n523 gnd 0.01055f
C2825 vdd.n524 gnd 0.01055f
C2826 vdd.n525 gnd 0.008492f
C2827 vdd.n526 gnd 0.008492f
C2828 vdd.n527 gnd 0.01055f
C2829 vdd.n528 gnd 0.01055f
C2830 vdd.n529 gnd 0.008492f
C2831 vdd.n530 gnd 0.01055f
C2832 vdd.n531 gnd 0.01055f
C2833 vdd.n532 gnd 0.01055f
C2834 vdd.n533 gnd 0.01055f
C2835 vdd.n534 gnd 0.01055f
C2836 vdd.n535 gnd 0.008492f
C2837 vdd.n536 gnd 0.008492f
C2838 vdd.n537 gnd 0.01055f
C2839 vdd.n538 gnd 0.01055f
C2840 vdd.n539 gnd 0.008492f
C2841 vdd.n540 gnd 0.01055f
C2842 vdd.n541 gnd 0.01055f
C2843 vdd.n542 gnd 0.01055f
C2844 vdd.n543 gnd 0.01055f
C2845 vdd.n544 gnd 0.01055f
C2846 vdd.n545 gnd 0.008492f
C2847 vdd.n546 gnd 0.008492f
C2848 vdd.n547 gnd 0.01055f
C2849 vdd.n548 gnd 0.01055f
C2850 vdd.n549 gnd 0.008492f
C2851 vdd.n550 gnd 0.01055f
C2852 vdd.n551 gnd 0.01055f
C2853 vdd.n552 gnd 0.01055f
C2854 vdd.n553 gnd 0.01055f
C2855 vdd.n554 gnd 0.01055f
C2856 vdd.n555 gnd 0.008492f
C2857 vdd.n556 gnd 0.008492f
C2858 vdd.n557 gnd 0.01055f
C2859 vdd.n558 gnd 0.01055f
C2860 vdd.n559 gnd 0.008492f
C2861 vdd.n560 gnd 0.01055f
C2862 vdd.n561 gnd 0.01055f
C2863 vdd.n562 gnd 0.01055f
C2864 vdd.n563 gnd 0.01055f
C2865 vdd.n564 gnd 0.01055f
C2866 vdd.n565 gnd 0.005774f
C2867 vdd.n566 gnd 0.018173f
C2868 vdd.n567 gnd 0.01055f
C2869 vdd.n568 gnd 0.01055f
C2870 vdd.n569 gnd 0.008407f
C2871 vdd.n570 gnd 0.01055f
C2872 vdd.n571 gnd 0.01055f
C2873 vdd.n572 gnd 0.01055f
C2874 vdd.n573 gnd 0.01055f
C2875 vdd.n574 gnd 0.01055f
C2876 vdd.n575 gnd 0.008492f
C2877 vdd.n576 gnd 0.008492f
C2878 vdd.n577 gnd 0.01055f
C2879 vdd.n578 gnd 0.01055f
C2880 vdd.n579 gnd 0.008492f
C2881 vdd.n580 gnd 0.01055f
C2882 vdd.n581 gnd 0.01055f
C2883 vdd.n582 gnd 0.01055f
C2884 vdd.n583 gnd 0.01055f
C2885 vdd.n584 gnd 0.01055f
C2886 vdd.n585 gnd 0.008492f
C2887 vdd.n586 gnd 0.008492f
C2888 vdd.n587 gnd 0.01055f
C2889 vdd.n588 gnd 0.01055f
C2890 vdd.n589 gnd 0.008492f
C2891 vdd.n590 gnd 0.01055f
C2892 vdd.n591 gnd 0.01055f
C2893 vdd.n592 gnd 0.01055f
C2894 vdd.n593 gnd 0.01055f
C2895 vdd.n594 gnd 0.01055f
C2896 vdd.n595 gnd 0.008492f
C2897 vdd.n596 gnd 0.008492f
C2898 vdd.n597 gnd 0.01055f
C2899 vdd.n598 gnd 0.01055f
C2900 vdd.n599 gnd 0.008492f
C2901 vdd.n600 gnd 0.01055f
C2902 vdd.n601 gnd 0.01055f
C2903 vdd.n602 gnd 0.01055f
C2904 vdd.n603 gnd 0.01055f
C2905 vdd.n604 gnd 0.01055f
C2906 vdd.n605 gnd 0.008492f
C2907 vdd.n606 gnd 0.008492f
C2908 vdd.n607 gnd 0.01055f
C2909 vdd.n608 gnd 0.01055f
C2910 vdd.n609 gnd 0.008492f
C2911 vdd.n610 gnd 0.01055f
C2912 vdd.n611 gnd 0.01055f
C2913 vdd.n612 gnd 0.01055f
C2914 vdd.n613 gnd 0.01055f
C2915 vdd.n614 gnd 0.01055f
C2916 vdd.n615 gnd 0.008492f
C2917 vdd.n616 gnd 0.01055f
C2918 vdd.n617 gnd 0.008492f
C2919 vdd.n618 gnd 0.004458f
C2920 vdd.n619 gnd 0.01055f
C2921 vdd.n620 gnd 0.01055f
C2922 vdd.n621 gnd 0.008492f
C2923 vdd.n622 gnd 0.01055f
C2924 vdd.n623 gnd 0.008492f
C2925 vdd.n624 gnd 0.01055f
C2926 vdd.n625 gnd 0.008492f
C2927 vdd.n626 gnd 0.01055f
C2928 vdd.n627 gnd 0.008492f
C2929 vdd.n628 gnd 0.01055f
C2930 vdd.n629 gnd 0.008492f
C2931 vdd.n630 gnd 0.01055f
C2932 vdd.n631 gnd 0.008492f
C2933 vdd.n632 gnd 0.01055f
C2934 vdd.n633 gnd 0.587625f
C2935 vdd.t157 gnd 0.539106f
C2936 vdd.n634 gnd 0.01055f
C2937 vdd.n635 gnd 0.008492f
C2938 vdd.n636 gnd 0.01055f
C2939 vdd.n637 gnd 0.008492f
C2940 vdd.n638 gnd 0.01055f
C2941 vdd.t168 gnd 0.539106f
C2942 vdd.n639 gnd 0.01055f
C2943 vdd.n640 gnd 0.008492f
C2944 vdd.n641 gnd 0.01055f
C2945 vdd.n642 gnd 0.008492f
C2946 vdd.n643 gnd 0.01055f
C2947 vdd.t161 gnd 0.539106f
C2948 vdd.n644 gnd 0.673882f
C2949 vdd.n645 gnd 0.01055f
C2950 vdd.n646 gnd 0.008492f
C2951 vdd.n647 gnd 0.01055f
C2952 vdd.n648 gnd 0.008492f
C2953 vdd.n649 gnd 0.01055f
C2954 vdd.t190 gnd 0.539106f
C2955 vdd.n650 gnd 0.01055f
C2956 vdd.n651 gnd 0.008492f
C2957 vdd.n652 gnd 0.01055f
C2958 vdd.n653 gnd 0.008492f
C2959 vdd.n654 gnd 0.01055f
C2960 vdd.n655 gnd 0.749357f
C2961 vdd.n656 gnd 0.894916f
C2962 vdd.t225 gnd 0.539106f
C2963 vdd.n657 gnd 0.01055f
C2964 vdd.n658 gnd 0.008492f
C2965 vdd.n659 gnd 0.01055f
C2966 vdd.n660 gnd 0.008492f
C2967 vdd.n661 gnd 0.01055f
C2968 vdd.n662 gnd 0.566061f
C2969 vdd.n663 gnd 0.01055f
C2970 vdd.n664 gnd 0.008492f
C2971 vdd.n665 gnd 0.01055f
C2972 vdd.n666 gnd 0.008492f
C2973 vdd.n667 gnd 0.01055f
C2974 vdd.t152 gnd 0.539106f
C2975 vdd.t185 gnd 0.539106f
C2976 vdd.n668 gnd 0.01055f
C2977 vdd.n669 gnd 0.008492f
C2978 vdd.n670 gnd 0.01055f
C2979 vdd.n671 gnd 0.008492f
C2980 vdd.n672 gnd 0.01055f
C2981 vdd.t198 gnd 0.539106f
C2982 vdd.n673 gnd 0.01055f
C2983 vdd.n674 gnd 0.008492f
C2984 vdd.n675 gnd 0.01055f
C2985 vdd.n676 gnd 0.008492f
C2986 vdd.n677 gnd 0.01055f
C2987 vdd.n678 gnd 1.07821f
C2988 vdd.n679 gnd 0.878743f
C2989 vdd.n680 gnd 0.01055f
C2990 vdd.n681 gnd 0.008492f
C2991 vdd.n682 gnd 0.025523f
C2992 vdd.n683 gnd 0.007048f
C2993 vdd.n684 gnd 0.025523f
C2994 vdd.t64 gnd 0.539106f
C2995 vdd.n685 gnd 0.025523f
C2996 vdd.n686 gnd 0.007048f
C2997 vdd.n687 gnd 0.009073f
C2998 vdd.t87 gnd 0.129799f
C2999 vdd.t88 gnd 0.138719f
C3000 vdd.t86 gnd 0.169516f
C3001 vdd.n688 gnd 0.217295f
C3002 vdd.n689 gnd 0.182567f
C3003 vdd.n690 gnd 0.013078f
C3004 vdd.n691 gnd 0.01055f
C3005 vdd.n692 gnd 10.965401f
C3006 vdd.n723 gnd 1.48254f
C3007 vdd.n724 gnd 0.01055f
C3008 vdd.n725 gnd 0.01055f
C3009 vdd.n726 gnd 0.026069f
C3010 vdd.n727 gnd 0.009073f
C3011 vdd.n728 gnd 0.01055f
C3012 vdd.n729 gnd 0.008492f
C3013 vdd.n730 gnd 0.006752f
C3014 vdd.n731 gnd 0.033676f
C3015 vdd.n732 gnd 0.008492f
C3016 vdd.n733 gnd 0.01055f
C3017 vdd.n734 gnd 0.01055f
C3018 vdd.n735 gnd 0.01055f
C3019 vdd.n736 gnd 0.01055f
C3020 vdd.n737 gnd 0.01055f
C3021 vdd.n738 gnd 0.01055f
C3022 vdd.n739 gnd 0.01055f
C3023 vdd.n740 gnd 0.01055f
C3024 vdd.n741 gnd 0.01055f
C3025 vdd.n742 gnd 0.01055f
C3026 vdd.n743 gnd 0.01055f
C3027 vdd.n744 gnd 0.01055f
C3028 vdd.n745 gnd 0.01055f
C3029 vdd.n746 gnd 0.01055f
C3030 vdd.n747 gnd 0.007091f
C3031 vdd.n748 gnd 0.01055f
C3032 vdd.n749 gnd 0.01055f
C3033 vdd.n750 gnd 0.01055f
C3034 vdd.n751 gnd 0.01055f
C3035 vdd.n752 gnd 0.01055f
C3036 vdd.n753 gnd 0.01055f
C3037 vdd.n754 gnd 0.01055f
C3038 vdd.n755 gnd 0.01055f
C3039 vdd.n756 gnd 0.01055f
C3040 vdd.n757 gnd 0.01055f
C3041 vdd.n758 gnd 0.01055f
C3042 vdd.n759 gnd 0.01055f
C3043 vdd.n760 gnd 0.01055f
C3044 vdd.n761 gnd 0.01055f
C3045 vdd.n762 gnd 0.01055f
C3046 vdd.n763 gnd 0.01055f
C3047 vdd.n764 gnd 0.01055f
C3048 vdd.n765 gnd 0.01055f
C3049 vdd.n766 gnd 0.01055f
C3050 vdd.n767 gnd 0.008407f
C3051 vdd.t65 gnd 0.129799f
C3052 vdd.t66 gnd 0.138719f
C3053 vdd.t63 gnd 0.169516f
C3054 vdd.n768 gnd 0.217295f
C3055 vdd.n769 gnd 0.182567f
C3056 vdd.n770 gnd 0.01055f
C3057 vdd.n771 gnd 0.01055f
C3058 vdd.n772 gnd 0.01055f
C3059 vdd.n773 gnd 0.01055f
C3060 vdd.n774 gnd 0.01055f
C3061 vdd.n775 gnd 0.01055f
C3062 vdd.n776 gnd 0.01055f
C3063 vdd.n777 gnd 0.01055f
C3064 vdd.n778 gnd 0.01055f
C3065 vdd.n779 gnd 0.01055f
C3066 vdd.n780 gnd 0.01055f
C3067 vdd.n781 gnd 0.01055f
C3068 vdd.n782 gnd 0.01055f
C3069 vdd.n783 gnd 0.006752f
C3070 vdd.n785 gnd 0.007174f
C3071 vdd.n786 gnd 0.007174f
C3072 vdd.n787 gnd 0.007174f
C3073 vdd.n788 gnd 0.007174f
C3074 vdd.n789 gnd 0.007174f
C3075 vdd.n790 gnd 0.007174f
C3076 vdd.n792 gnd 0.007174f
C3077 vdd.n793 gnd 0.007174f
C3078 vdd.n795 gnd 0.007174f
C3079 vdd.n796 gnd 0.005223f
C3080 vdd.n798 gnd 0.007174f
C3081 vdd.t70 gnd 0.289914f
C3082 vdd.t69 gnd 0.296763f
C3083 vdd.t67 gnd 0.189267f
C3084 vdd.n799 gnd 0.102288f
C3085 vdd.n800 gnd 0.058021f
C3086 vdd.n801 gnd 0.010253f
C3087 vdd.n802 gnd 0.016447f
C3088 vdd.n804 gnd 0.007174f
C3089 vdd.n805 gnd 0.733184f
C3090 vdd.n806 gnd 0.015538f
C3091 vdd.n807 gnd 0.015538f
C3092 vdd.n808 gnd 0.007174f
C3093 vdd.n809 gnd 0.016536f
C3094 vdd.n810 gnd 0.007174f
C3095 vdd.n811 gnd 0.007174f
C3096 vdd.n812 gnd 0.007174f
C3097 vdd.n813 gnd 0.007174f
C3098 vdd.n814 gnd 0.007174f
C3099 vdd.n816 gnd 0.007174f
C3100 vdd.n817 gnd 0.007174f
C3101 vdd.n819 gnd 0.007174f
C3102 vdd.n820 gnd 0.007174f
C3103 vdd.n822 gnd 0.007174f
C3104 vdd.n823 gnd 0.007174f
C3105 vdd.n825 gnd 0.007174f
C3106 vdd.n826 gnd 0.007174f
C3107 vdd.n828 gnd 0.007174f
C3108 vdd.n829 gnd 0.007174f
C3109 vdd.n831 gnd 0.007174f
C3110 vdd.t98 gnd 0.289914f
C3111 vdd.t97 gnd 0.296763f
C3112 vdd.t96 gnd 0.189267f
C3113 vdd.n832 gnd 0.102288f
C3114 vdd.n833 gnd 0.058021f
C3115 vdd.n834 gnd 0.007174f
C3116 vdd.n836 gnd 0.007174f
C3117 vdd.n837 gnd 0.007174f
C3118 vdd.t68 gnd 0.366592f
C3119 vdd.n838 gnd 0.007174f
C3120 vdd.n839 gnd 0.007174f
C3121 vdd.n840 gnd 0.007174f
C3122 vdd.n841 gnd 0.007174f
C3123 vdd.n842 gnd 0.007174f
C3124 vdd.n843 gnd 0.733184f
C3125 vdd.n844 gnd 0.007174f
C3126 vdd.n845 gnd 0.007174f
C3127 vdd.n846 gnd 0.598408f
C3128 vdd.n847 gnd 0.007174f
C3129 vdd.n848 gnd 0.007174f
C3130 vdd.n849 gnd 0.007174f
C3131 vdd.n850 gnd 0.007174f
C3132 vdd.n851 gnd 0.733184f
C3133 vdd.n852 gnd 0.007174f
C3134 vdd.n853 gnd 0.007174f
C3135 vdd.n854 gnd 0.007174f
C3136 vdd.n855 gnd 0.007174f
C3137 vdd.n856 gnd 0.007174f
C3138 vdd.t19 gnd 0.366592f
C3139 vdd.n857 gnd 0.007174f
C3140 vdd.n858 gnd 0.007174f
C3141 vdd.n859 gnd 0.007174f
C3142 vdd.n860 gnd 0.007174f
C3143 vdd.n861 gnd 0.007174f
C3144 vdd.t16 gnd 0.366592f
C3145 vdd.n862 gnd 0.007174f
C3146 vdd.n863 gnd 0.007174f
C3147 vdd.n864 gnd 0.727793f
C3148 vdd.n865 gnd 0.007174f
C3149 vdd.n866 gnd 0.007174f
C3150 vdd.n867 gnd 0.007174f
C3151 vdd.t43 gnd 0.366592f
C3152 vdd.n868 gnd 0.007174f
C3153 vdd.n869 gnd 0.007174f
C3154 vdd.n870 gnd 0.566061f
C3155 vdd.n871 gnd 0.007174f
C3156 vdd.n872 gnd 0.007174f
C3157 vdd.n873 gnd 0.007174f
C3158 vdd.n874 gnd 0.490586f
C3159 vdd.n875 gnd 0.007174f
C3160 vdd.n876 gnd 0.007174f
C3161 vdd.n877 gnd 0.404329f
C3162 vdd.n878 gnd 0.007174f
C3163 vdd.n879 gnd 0.007174f
C3164 vdd.n880 gnd 0.007174f
C3165 vdd.n881 gnd 0.603799f
C3166 vdd.n882 gnd 0.007174f
C3167 vdd.n883 gnd 0.007174f
C3168 vdd.t299 gnd 0.366592f
C3169 vdd.n884 gnd 0.007174f
C3170 vdd.t84 gnd 0.296763f
C3171 vdd.t82 gnd 0.189267f
C3172 vdd.t85 gnd 0.296763f
C3173 vdd.n885 gnd 0.166793f
C3174 vdd.n886 gnd 0.007174f
C3175 vdd.n887 gnd 0.007174f
C3176 vdd.n888 gnd 0.733184f
C3177 vdd.n889 gnd 0.007174f
C3178 vdd.n890 gnd 0.007174f
C3179 vdd.t83 gnd 0.285726f
C3180 vdd.t25 gnd 0.129385f
C3181 vdd.n891 gnd 0.007174f
C3182 vdd.n892 gnd 0.007174f
C3183 vdd.n893 gnd 0.007174f
C3184 vdd.t13 gnd 0.366592f
C3185 vdd.n894 gnd 0.007174f
C3186 vdd.n895 gnd 0.007174f
C3187 vdd.n896 gnd 0.007174f
C3188 vdd.n897 gnd 0.007174f
C3189 vdd.n898 gnd 0.007174f
C3190 vdd.t18 gnd 0.366592f
C3191 vdd.n899 gnd 0.007174f
C3192 vdd.n900 gnd 0.007174f
C3193 vdd.n901 gnd 0.652318f
C3194 vdd.n902 gnd 0.007174f
C3195 vdd.n903 gnd 0.007174f
C3196 vdd.n904 gnd 0.007174f
C3197 vdd.n905 gnd 0.404329f
C3198 vdd.n906 gnd 0.007174f
C3199 vdd.n907 gnd 0.007174f
C3200 vdd.t5 gnd 0.366592f
C3201 vdd.n908 gnd 0.007174f
C3202 vdd.n909 gnd 0.007174f
C3203 vdd.n910 gnd 0.007174f
C3204 vdd.n911 gnd 0.566061f
C3205 vdd.n912 gnd 0.007174f
C3206 vdd.n913 gnd 0.007174f
C3207 vdd.t9 gnd 0.269553f
C3208 vdd.t49 gnd 0.328855f
C3209 vdd.n914 gnd 0.007174f
C3210 vdd.n915 gnd 0.007174f
C3211 vdd.n916 gnd 0.007174f
C3212 vdd.t33 gnd 0.366592f
C3213 vdd.n917 gnd 0.007174f
C3214 vdd.n918 gnd 0.007174f
C3215 vdd.t8 gnd 0.366592f
C3216 vdd.n919 gnd 0.007174f
C3217 vdd.n920 gnd 0.007174f
C3218 vdd.n921 gnd 0.007174f
C3219 vdd.t20 gnd 0.366592f
C3220 vdd.n922 gnd 0.007174f
C3221 vdd.n923 gnd 0.007174f
C3222 vdd.t46 gnd 0.366592f
C3223 vdd.n924 gnd 0.007174f
C3224 vdd.n925 gnd 0.007174f
C3225 vdd.n926 gnd 0.007174f
C3226 vdd.n927 gnd 0.733184f
C3227 vdd.n928 gnd 0.007174f
C3228 vdd.n929 gnd 0.007174f
C3229 vdd.n930 gnd 0.50676f
C3230 vdd.n931 gnd 0.007174f
C3231 vdd.n932 gnd 0.007174f
C3232 vdd.n933 gnd 0.007174f
C3233 vdd.t302 gnd 0.366592f
C3234 vdd.n934 gnd 0.007174f
C3235 vdd.n935 gnd 0.007174f
C3236 vdd.n936 gnd 0.007174f
C3237 vdd.n937 gnd 0.007174f
C3238 vdd.n938 gnd 0.007174f
C3239 vdd.t29 gnd 0.366592f
C3240 vdd.n939 gnd 0.007174f
C3241 vdd.n940 gnd 0.007174f
C3242 vdd.t114 gnd 0.366592f
C3243 vdd.n941 gnd 0.007174f
C3244 vdd.n942 gnd 0.016536f
C3245 vdd.n943 gnd 0.016536f
C3246 vdd.t31 gnd 0.646927f
C3247 vdd.n944 gnd 0.015538f
C3248 vdd.n945 gnd 0.015538f
C3249 vdd.n946 gnd 0.409721f
C3250 vdd.n947 gnd 0.016536f
C3251 vdd.n948 gnd 0.007174f
C3252 vdd.n949 gnd 0.007174f
C3253 vdd.t39 gnd 0.646927f
C3254 vdd.n967 gnd 0.016536f
C3255 vdd.n985 gnd 0.015538f
C3256 vdd.n986 gnd 0.007174f
C3257 vdd.n987 gnd 0.015538f
C3258 vdd.t135 gnd 0.289914f
C3259 vdd.t134 gnd 0.296763f
C3260 vdd.t133 gnd 0.189267f
C3261 vdd.n988 gnd 0.102288f
C3262 vdd.n989 gnd 0.058021f
C3263 vdd.n990 gnd 0.016447f
C3264 vdd.n991 gnd 0.007174f
C3265 vdd.n992 gnd 0.409721f
C3266 vdd.n993 gnd 0.015538f
C3267 vdd.n994 gnd 0.007174f
C3268 vdd.n995 gnd 0.016536f
C3269 vdd.n996 gnd 0.007174f
C3270 vdd.t112 gnd 0.289914f
C3271 vdd.t111 gnd 0.296763f
C3272 vdd.t109 gnd 0.189267f
C3273 vdd.n997 gnd 0.102288f
C3274 vdd.n998 gnd 0.058021f
C3275 vdd.n999 gnd 0.010253f
C3276 vdd.n1000 gnd 0.007174f
C3277 vdd.n1001 gnd 0.007174f
C3278 vdd.t110 gnd 0.366592f
C3279 vdd.n1002 gnd 0.007174f
C3280 vdd.t37 gnd 0.366592f
C3281 vdd.n1003 gnd 0.007174f
C3282 vdd.n1004 gnd 0.007174f
C3283 vdd.n1005 gnd 0.007174f
C3284 vdd.n1006 gnd 0.007174f
C3285 vdd.n1007 gnd 0.007174f
C3286 vdd.n1008 gnd 0.733184f
C3287 vdd.n1009 gnd 0.007174f
C3288 vdd.n1010 gnd 0.007174f
C3289 vdd.t3 gnd 0.366592f
C3290 vdd.n1011 gnd 0.007174f
C3291 vdd.n1012 gnd 0.007174f
C3292 vdd.n1013 gnd 0.007174f
C3293 vdd.n1014 gnd 0.007174f
C3294 vdd.n1015 gnd 0.50676f
C3295 vdd.n1016 gnd 0.007174f
C3296 vdd.n1017 gnd 0.007174f
C3297 vdd.n1018 gnd 0.007174f
C3298 vdd.n1019 gnd 0.007174f
C3299 vdd.n1020 gnd 0.007174f
C3300 vdd.t44 gnd 0.366592f
C3301 vdd.n1021 gnd 0.007174f
C3302 vdd.n1022 gnd 0.007174f
C3303 vdd.t14 gnd 0.366592f
C3304 vdd.n1023 gnd 0.007174f
C3305 vdd.n1024 gnd 0.007174f
C3306 vdd.n1025 gnd 0.007174f
C3307 vdd.t12 gnd 0.366592f
C3308 vdd.n1026 gnd 0.007174f
C3309 vdd.n1027 gnd 0.007174f
C3310 vdd.t47 gnd 0.366592f
C3311 vdd.n1028 gnd 0.007174f
C3312 vdd.n1029 gnd 0.007174f
C3313 vdd.n1030 gnd 0.007174f
C3314 vdd.t22 gnd 0.328855f
C3315 vdd.n1031 gnd 0.007174f
C3316 vdd.n1032 gnd 0.007174f
C3317 vdd.n1033 gnd 0.566061f
C3318 vdd.n1034 gnd 0.007174f
C3319 vdd.n1035 gnd 0.007174f
C3320 vdd.n1036 gnd 0.007174f
C3321 vdd.t35 gnd 0.366592f
C3322 vdd.n1037 gnd 0.007174f
C3323 vdd.n1038 gnd 0.007174f
C3324 vdd.t7 gnd 0.269553f
C3325 vdd.n1039 gnd 0.404329f
C3326 vdd.n1040 gnd 0.007174f
C3327 vdd.n1041 gnd 0.007174f
C3328 vdd.n1042 gnd 0.007174f
C3329 vdd.n1043 gnd 0.652318f
C3330 vdd.n1044 gnd 0.007174f
C3331 vdd.n1045 gnd 0.007174f
C3332 vdd.t42 gnd 0.366592f
C3333 vdd.n1046 gnd 0.007174f
C3334 vdd.n1047 gnd 0.007174f
C3335 vdd.n1048 gnd 0.007174f
C3336 vdd.n1049 gnd 0.733184f
C3337 vdd.n1050 gnd 0.007174f
C3338 vdd.n1051 gnd 0.007174f
C3339 vdd.t24 gnd 0.366592f
C3340 vdd.n1052 gnd 0.007174f
C3341 vdd.n1053 gnd 0.007174f
C3342 vdd.n1054 gnd 0.007174f
C3343 vdd.t26 gnd 0.129385f
C3344 vdd.n1055 gnd 0.007174f
C3345 vdd.n1056 gnd 0.007174f
C3346 vdd.n1057 gnd 0.007174f
C3347 vdd.t125 gnd 0.296763f
C3348 vdd.t123 gnd 0.189267f
C3349 vdd.t126 gnd 0.296763f
C3350 vdd.n1058 gnd 0.166793f
C3351 vdd.n1059 gnd 0.007174f
C3352 vdd.n1060 gnd 0.007174f
C3353 vdd.t41 gnd 0.366592f
C3354 vdd.n1061 gnd 0.007174f
C3355 vdd.n1062 gnd 0.007174f
C3356 vdd.t124 gnd 0.285726f
C3357 vdd.n1063 gnd 0.603799f
C3358 vdd.n1064 gnd 0.007174f
C3359 vdd.n1065 gnd 0.007174f
C3360 vdd.n1066 gnd 0.007174f
C3361 vdd.n1067 gnd 0.404329f
C3362 vdd.n1068 gnd 0.007174f
C3363 vdd.n1069 gnd 0.007174f
C3364 vdd.n1070 gnd 0.490586f
C3365 vdd.n1071 gnd 0.007174f
C3366 vdd.n1072 gnd 0.007174f
C3367 vdd.n1073 gnd 0.007174f
C3368 vdd.n1074 gnd 0.566061f
C3369 vdd.n1075 gnd 0.007174f
C3370 vdd.n1076 gnd 0.007174f
C3371 vdd.t45 gnd 0.366592f
C3372 vdd.n1077 gnd 0.007174f
C3373 vdd.n1078 gnd 0.007174f
C3374 vdd.n1079 gnd 0.007174f
C3375 vdd.n1080 gnd 0.727793f
C3376 vdd.n1081 gnd 0.007174f
C3377 vdd.n1082 gnd 0.007174f
C3378 vdd.t2 gnd 0.366592f
C3379 vdd.n1083 gnd 0.007174f
C3380 vdd.n1084 gnd 0.007174f
C3381 vdd.n1085 gnd 0.007174f
C3382 vdd.n1086 gnd 0.733184f
C3383 vdd.n1087 gnd 0.007174f
C3384 vdd.n1088 gnd 0.007174f
C3385 vdd.t17 gnd 0.366592f
C3386 vdd.n1089 gnd 0.007174f
C3387 vdd.n1090 gnd 0.007174f
C3388 vdd.n1091 gnd 0.007174f
C3389 vdd.n1092 gnd 0.733184f
C3390 vdd.n1093 gnd 0.007174f
C3391 vdd.n1094 gnd 0.007174f
C3392 vdd.n1095 gnd 0.007174f
C3393 vdd.n1096 gnd 0.007174f
C3394 vdd.n1097 gnd 0.007174f
C3395 vdd.n1098 gnd 0.598408f
C3396 vdd.n1099 gnd 0.007174f
C3397 vdd.n1100 gnd 0.007174f
C3398 vdd.n1101 gnd 0.007174f
C3399 vdd.n1102 gnd 0.007174f
C3400 vdd.n1103 gnd 0.007174f
C3401 vdd.n1104 gnd 0.733184f
C3402 vdd.n1105 gnd 0.007174f
C3403 vdd.n1106 gnd 0.007174f
C3404 vdd.t72 gnd 0.366592f
C3405 vdd.n1107 gnd 0.007174f
C3406 vdd.n1108 gnd 0.016536f
C3407 vdd.n1109 gnd 0.016536f
C3408 vdd.n1110 gnd 10.965401f
C3409 vdd.n1111 gnd 0.015538f
C3410 vdd.n1112 gnd 0.015538f
C3411 vdd.n1113 gnd 0.016536f
C3412 vdd.n1114 gnd 0.007174f
C3413 vdd.n1116 gnd 0.007174f
C3414 vdd.n1117 gnd 0.007174f
C3415 vdd.n1118 gnd 0.007174f
C3416 vdd.n1119 gnd 0.007174f
C3417 vdd.n1120 gnd 0.007174f
C3418 vdd.n1121 gnd 0.007174f
C3419 vdd.n1122 gnd 0.037749f
C3420 vdd.n1123 gnd 0.007174f
C3421 vdd.n1124 gnd 0.007174f
C3422 vdd.n1125 gnd 0.007174f
C3423 vdd.n1126 gnd 0.007174f
C3424 vdd.n1127 gnd 0.007174f
C3425 vdd.n1128 gnd 0.007174f
C3426 vdd.n1129 gnd 0.007174f
C3427 vdd.t137 gnd 0.289914f
C3428 vdd.t138 gnd 0.296763f
C3429 vdd.t136 gnd 0.189267f
C3430 vdd.n1130 gnd 0.102288f
C3431 vdd.n1131 gnd 0.058021f
C3432 vdd.n1132 gnd 0.007174f
C3433 vdd.n1133 gnd 0.007174f
C3434 vdd.n1134 gnd 0.007174f
C3435 vdd.n1135 gnd 0.007174f
C3436 vdd.t73 gnd 0.289914f
C3437 vdd.t74 gnd 0.296763f
C3438 vdd.t71 gnd 0.189267f
C3439 vdd.n1136 gnd 0.102288f
C3440 vdd.n1137 gnd 0.058021f
C3441 vdd.n1138 gnd 0.007174f
C3442 vdd.n1139 gnd 0.007174f
C3443 vdd.n1140 gnd 0.007174f
C3444 vdd.n1141 gnd 0.007174f
C3445 vdd.n1142 gnd 0.007174f
C3446 vdd.n1143 gnd 0.007174f
C3447 vdd.n1144 gnd 0.006752f
C3448 vdd.n1147 gnd 0.026069f
C3449 vdd.n1148 gnd 0.008492f
C3450 vdd.n1149 gnd 0.01055f
C3451 vdd.n1151 gnd 0.01055f
C3452 vdd.n1152 gnd 0.007048f
C3453 vdd.t90 gnd 0.539106f
C3454 vdd.n1153 gnd 11.375099f
C3455 vdd.n1154 gnd 0.01055f
C3456 vdd.n1155 gnd 0.026069f
C3457 vdd.n1156 gnd 0.008492f
C3458 vdd.n1157 gnd 0.01055f
C3459 vdd.n1158 gnd 0.008492f
C3460 vdd.n1159 gnd 0.01055f
C3461 vdd.n1160 gnd 1.07821f
C3462 vdd.n1161 gnd 0.01055f
C3463 vdd.n1162 gnd 0.008492f
C3464 vdd.n1163 gnd 0.008492f
C3465 vdd.n1164 gnd 0.01055f
C3466 vdd.n1165 gnd 0.008492f
C3467 vdd.n1166 gnd 0.01055f
C3468 vdd.t238 gnd 0.539106f
C3469 vdd.n1167 gnd 0.01055f
C3470 vdd.n1168 gnd 0.008492f
C3471 vdd.n1169 gnd 0.01055f
C3472 vdd.n1170 gnd 0.008492f
C3473 vdd.n1171 gnd 0.01055f
C3474 vdd.t155 gnd 0.539106f
C3475 vdd.n1172 gnd 0.01055f
C3476 vdd.n1173 gnd 0.008492f
C3477 vdd.n1174 gnd 0.01055f
C3478 vdd.n1175 gnd 0.008492f
C3479 vdd.n1176 gnd 0.01055f
C3480 vdd.n1177 gnd 0.867961f
C3481 vdd.n1178 gnd 0.894916f
C3482 vdd.t202 gnd 0.539106f
C3483 vdd.n1179 gnd 0.01055f
C3484 vdd.n1180 gnd 0.008492f
C3485 vdd.n1181 gnd 0.01055f
C3486 vdd.n1182 gnd 0.008492f
C3487 vdd.n1183 gnd 0.01055f
C3488 vdd.n1184 gnd 0.684665f
C3489 vdd.n1185 gnd 0.01055f
C3490 vdd.n1186 gnd 0.008492f
C3491 vdd.n1187 gnd 0.01055f
C3492 vdd.n1188 gnd 0.008492f
C3493 vdd.n1189 gnd 0.01055f
C3494 vdd.t232 gnd 0.539106f
C3495 vdd.t179 gnd 0.539106f
C3496 vdd.n1190 gnd 0.01055f
C3497 vdd.n1191 gnd 0.008492f
C3498 vdd.n1192 gnd 0.01055f
C3499 vdd.n1193 gnd 0.008492f
C3500 vdd.n1194 gnd 0.01055f
C3501 vdd.t236 gnd 0.539106f
C3502 vdd.n1195 gnd 0.01055f
C3503 vdd.n1196 gnd 0.008492f
C3504 vdd.n1197 gnd 0.01055f
C3505 vdd.n1198 gnd 0.008492f
C3506 vdd.n1199 gnd 0.01055f
C3507 vdd.t143 gnd 0.539106f
C3508 vdd.n1200 gnd 0.760139f
C3509 vdd.n1201 gnd 0.01055f
C3510 vdd.n1202 gnd 0.008492f
C3511 vdd.n1203 gnd 0.01055f
C3512 vdd.n1204 gnd 0.008492f
C3513 vdd.n1205 gnd 0.01055f
C3514 vdd.n1206 gnd 0.846396f
C3515 vdd.n1207 gnd 0.01055f
C3516 vdd.n1208 gnd 0.008492f
C3517 vdd.n1209 gnd 0.01055f
C3518 vdd.n1210 gnd 0.008492f
C3519 vdd.n1211 gnd 0.01055f
C3520 vdd.n1212 gnd 0.6631f
C3521 vdd.t177 gnd 0.539106f
C3522 vdd.n1213 gnd 0.01055f
C3523 vdd.n1214 gnd 0.008492f
C3524 vdd.n1215 gnd 0.01055f
C3525 vdd.n1216 gnd 0.008492f
C3526 vdd.n1217 gnd 0.01055f
C3527 vdd.t148 gnd 0.539106f
C3528 vdd.n1218 gnd 0.01055f
C3529 vdd.n1219 gnd 0.008492f
C3530 vdd.n1220 gnd 0.01055f
C3531 vdd.n1221 gnd 0.008492f
C3532 vdd.n1222 gnd 0.01055f
C3533 vdd.t204 gnd 0.539106f
C3534 vdd.n1223 gnd 0.598408f
C3535 vdd.n1224 gnd 0.01055f
C3536 vdd.n1225 gnd 0.008492f
C3537 vdd.n1226 gnd 0.01055f
C3538 vdd.n1227 gnd 0.008492f
C3539 vdd.n1228 gnd 0.01055f
C3540 vdd.t230 gnd 0.539106f
C3541 vdd.n1229 gnd 0.01055f
C3542 vdd.n1230 gnd 0.008492f
C3543 vdd.n1231 gnd 0.01055f
C3544 vdd.n1232 gnd 0.008492f
C3545 vdd.n1233 gnd 0.01055f
C3546 vdd.n1234 gnd 0.824832f
C3547 vdd.n1235 gnd 0.894916f
C3548 vdd.t139 gnd 0.539106f
C3549 vdd.n1236 gnd 0.01055f
C3550 vdd.n1237 gnd 0.008492f
C3551 vdd.n1238 gnd 0.01055f
C3552 vdd.n1239 gnd 0.008492f
C3553 vdd.n1240 gnd 0.01055f
C3554 vdd.n1241 gnd 0.641536f
C3555 vdd.n1242 gnd 0.01055f
C3556 vdd.n1243 gnd 0.008492f
C3557 vdd.n1244 gnd 0.01055f
C3558 vdd.n1245 gnd 0.008492f
C3559 vdd.n1246 gnd 0.01055f
C3560 vdd.t220 gnd 0.539106f
C3561 vdd.t240 gnd 0.539106f
C3562 vdd.n1247 gnd 0.01055f
C3563 vdd.n1248 gnd 0.008492f
C3564 vdd.n1249 gnd 0.01055f
C3565 vdd.n1250 gnd 0.008492f
C3566 vdd.n1251 gnd 0.01055f
C3567 vdd.t181 gnd 0.539106f
C3568 vdd.n1252 gnd 0.01055f
C3569 vdd.n1253 gnd 0.008492f
C3570 vdd.n1254 gnd 0.01055f
C3571 vdd.n1255 gnd 0.008492f
C3572 vdd.n1256 gnd 0.01055f
C3573 vdd.t234 gnd 0.539106f
C3574 vdd.n1257 gnd 0.803268f
C3575 vdd.n1258 gnd 0.01055f
C3576 vdd.n1259 gnd 0.008492f
C3577 vdd.n1260 gnd 0.01055f
C3578 vdd.n1261 gnd 0.008492f
C3579 vdd.n1262 gnd 0.01055f
C3580 vdd.n1263 gnd 1.07821f
C3581 vdd.n1264 gnd 0.01055f
C3582 vdd.n1265 gnd 0.008492f
C3583 vdd.n1266 gnd 0.025523f
C3584 vdd.n1267 gnd 0.007048f
C3585 vdd.n1268 gnd 0.025523f
C3586 vdd.t106 gnd 0.539106f
C3587 vdd.n1269 gnd 0.025523f
C3588 vdd.n1270 gnd 0.007048f
C3589 vdd.n1271 gnd 0.01055f
C3590 vdd.n1272 gnd 0.008492f
C3591 vdd.n1273 gnd 0.01055f
C3592 vdd.n1304 gnd 0.026069f
C3593 vdd.n1305 gnd 1.59036f
C3594 vdd.n1306 gnd 0.01055f
C3595 vdd.n1307 gnd 0.008492f
C3596 vdd.n1308 gnd 0.01055f
C3597 vdd.n1309 gnd 0.01055f
C3598 vdd.n1310 gnd 0.01055f
C3599 vdd.n1311 gnd 0.01055f
C3600 vdd.n1312 gnd 0.01055f
C3601 vdd.n1313 gnd 0.008492f
C3602 vdd.n1314 gnd 0.01055f
C3603 vdd.n1315 gnd 0.01055f
C3604 vdd.n1316 gnd 0.01055f
C3605 vdd.n1317 gnd 0.01055f
C3606 vdd.n1318 gnd 0.01055f
C3607 vdd.n1319 gnd 0.008492f
C3608 vdd.n1320 gnd 0.01055f
C3609 vdd.n1321 gnd 0.01055f
C3610 vdd.n1322 gnd 0.01055f
C3611 vdd.n1323 gnd 0.01055f
C3612 vdd.n1324 gnd 0.01055f
C3613 vdd.n1325 gnd 0.008492f
C3614 vdd.n1326 gnd 0.01055f
C3615 vdd.n1327 gnd 0.01055f
C3616 vdd.n1328 gnd 0.01055f
C3617 vdd.n1329 gnd 0.01055f
C3618 vdd.n1330 gnd 0.01055f
C3619 vdd.t131 gnd 0.129799f
C3620 vdd.t132 gnd 0.138719f
C3621 vdd.t130 gnd 0.169516f
C3622 vdd.n1331 gnd 0.217295f
C3623 vdd.n1332 gnd 0.183417f
C3624 vdd.n1333 gnd 0.018173f
C3625 vdd.n1334 gnd 0.01055f
C3626 vdd.n1335 gnd 0.01055f
C3627 vdd.n1336 gnd 0.01055f
C3628 vdd.n1337 gnd 0.01055f
C3629 vdd.n1338 gnd 0.01055f
C3630 vdd.n1339 gnd 0.008492f
C3631 vdd.n1340 gnd 0.01055f
C3632 vdd.n1341 gnd 0.01055f
C3633 vdd.n1342 gnd 0.01055f
C3634 vdd.n1343 gnd 0.01055f
C3635 vdd.n1344 gnd 0.01055f
C3636 vdd.n1345 gnd 0.008492f
C3637 vdd.n1346 gnd 0.01055f
C3638 vdd.n1347 gnd 0.01055f
C3639 vdd.n1348 gnd 0.01055f
C3640 vdd.n1349 gnd 0.01055f
C3641 vdd.n1350 gnd 0.01055f
C3642 vdd.n1351 gnd 0.008492f
C3643 vdd.n1352 gnd 0.01055f
C3644 vdd.n1353 gnd 0.01055f
C3645 vdd.n1354 gnd 0.01055f
C3646 vdd.n1355 gnd 0.01055f
C3647 vdd.n1356 gnd 0.01055f
C3648 vdd.n1357 gnd 0.008492f
C3649 vdd.n1358 gnd 0.01055f
C3650 vdd.n1359 gnd 0.01055f
C3651 vdd.n1360 gnd 0.01055f
C3652 vdd.n1361 gnd 0.01055f
C3653 vdd.n1362 gnd 0.01055f
C3654 vdd.n1363 gnd 0.008492f
C3655 vdd.n1364 gnd 0.01055f
C3656 vdd.n1365 gnd 0.01055f
C3657 vdd.n1366 gnd 0.01055f
C3658 vdd.n1367 gnd 0.01055f
C3659 vdd.n1368 gnd 0.008492f
C3660 vdd.n1369 gnd 0.01055f
C3661 vdd.n1370 gnd 0.01055f
C3662 vdd.n1371 gnd 0.01055f
C3663 vdd.n1372 gnd 0.01055f
C3664 vdd.n1373 gnd 0.01055f
C3665 vdd.n1374 gnd 0.008492f
C3666 vdd.n1375 gnd 0.01055f
C3667 vdd.n1376 gnd 0.01055f
C3668 vdd.n1377 gnd 0.01055f
C3669 vdd.n1378 gnd 0.01055f
C3670 vdd.n1379 gnd 0.01055f
C3671 vdd.n1380 gnd 0.008492f
C3672 vdd.n1381 gnd 0.01055f
C3673 vdd.n1382 gnd 0.01055f
C3674 vdd.n1383 gnd 0.01055f
C3675 vdd.n1384 gnd 0.01055f
C3676 vdd.n1385 gnd 0.01055f
C3677 vdd.n1386 gnd 0.008492f
C3678 vdd.n1387 gnd 0.01055f
C3679 vdd.n1388 gnd 0.01055f
C3680 vdd.n1389 gnd 0.01055f
C3681 vdd.n1390 gnd 0.01055f
C3682 vdd.n1391 gnd 0.01055f
C3683 vdd.n1392 gnd 0.008492f
C3684 vdd.n1393 gnd 0.01055f
C3685 vdd.n1394 gnd 0.01055f
C3686 vdd.n1395 gnd 0.01055f
C3687 vdd.n1396 gnd 0.01055f
C3688 vdd.t107 gnd 0.129799f
C3689 vdd.t108 gnd 0.138719f
C3690 vdd.t105 gnd 0.169516f
C3691 vdd.n1397 gnd 0.217295f
C3692 vdd.n1398 gnd 0.183417f
C3693 vdd.n1399 gnd 0.013927f
C3694 vdd.n1400 gnd 0.004034f
C3695 vdd.n1401 gnd 0.026069f
C3696 vdd.n1402 gnd 0.01055f
C3697 vdd.n1403 gnd 0.004458f
C3698 vdd.n1404 gnd 0.008492f
C3699 vdd.n1405 gnd 0.008492f
C3700 vdd.n1406 gnd 0.01055f
C3701 vdd.n1407 gnd 0.01055f
C3702 vdd.n1408 gnd 0.01055f
C3703 vdd.n1409 gnd 0.008492f
C3704 vdd.n1410 gnd 0.008492f
C3705 vdd.n1411 gnd 0.008492f
C3706 vdd.n1412 gnd 0.01055f
C3707 vdd.n1413 gnd 0.01055f
C3708 vdd.n1414 gnd 0.01055f
C3709 vdd.n1415 gnd 0.008492f
C3710 vdd.n1416 gnd 0.008492f
C3711 vdd.n1417 gnd 0.008492f
C3712 vdd.n1418 gnd 0.01055f
C3713 vdd.n1419 gnd 0.01055f
C3714 vdd.n1420 gnd 0.01055f
C3715 vdd.n1421 gnd 0.008492f
C3716 vdd.n1422 gnd 0.008492f
C3717 vdd.n1423 gnd 0.008492f
C3718 vdd.n1424 gnd 0.01055f
C3719 vdd.n1425 gnd 0.01055f
C3720 vdd.n1426 gnd 0.01055f
C3721 vdd.n1427 gnd 0.008492f
C3722 vdd.n1428 gnd 0.008492f
C3723 vdd.n1429 gnd 0.008492f
C3724 vdd.n1430 gnd 0.01055f
C3725 vdd.n1431 gnd 0.01055f
C3726 vdd.n1432 gnd 0.01055f
C3727 vdd.n1433 gnd 0.008407f
C3728 vdd.n1434 gnd 0.01055f
C3729 vdd.t118 gnd 0.129799f
C3730 vdd.t119 gnd 0.138719f
C3731 vdd.t117 gnd 0.169516f
C3732 vdd.n1435 gnd 0.217295f
C3733 vdd.n1436 gnd 0.183417f
C3734 vdd.n1437 gnd 0.018173f
C3735 vdd.n1438 gnd 0.005774f
C3736 vdd.n1439 gnd 0.01055f
C3737 vdd.n1440 gnd 0.01055f
C3738 vdd.n1441 gnd 0.01055f
C3739 vdd.n1442 gnd 0.008492f
C3740 vdd.n1443 gnd 0.008492f
C3741 vdd.n1444 gnd 0.008492f
C3742 vdd.n1445 gnd 0.01055f
C3743 vdd.n1446 gnd 0.01055f
C3744 vdd.n1447 gnd 0.01055f
C3745 vdd.n1448 gnd 0.008492f
C3746 vdd.n1449 gnd 0.008492f
C3747 vdd.n1450 gnd 0.008492f
C3748 vdd.n1451 gnd 0.01055f
C3749 vdd.n1452 gnd 0.01055f
C3750 vdd.n1453 gnd 0.01055f
C3751 vdd.n1454 gnd 0.008492f
C3752 vdd.n1455 gnd 0.008492f
C3753 vdd.n1456 gnd 0.008492f
C3754 vdd.n1457 gnd 0.01055f
C3755 vdd.n1458 gnd 0.01055f
C3756 vdd.n1459 gnd 0.01055f
C3757 vdd.n1460 gnd 0.008492f
C3758 vdd.n1461 gnd 0.008492f
C3759 vdd.n1462 gnd 0.008492f
C3760 vdd.n1463 gnd 0.01055f
C3761 vdd.n1464 gnd 0.01055f
C3762 vdd.n1465 gnd 0.01055f
C3763 vdd.n1466 gnd 0.008492f
C3764 vdd.n1467 gnd 0.008492f
C3765 vdd.n1468 gnd 0.007091f
C3766 vdd.n1469 gnd 0.01055f
C3767 vdd.n1470 gnd 0.01055f
C3768 vdd.n1471 gnd 0.01055f
C3769 vdd.n1472 gnd 0.007091f
C3770 vdd.n1473 gnd 0.008492f
C3771 vdd.n1474 gnd 0.008492f
C3772 vdd.n1475 gnd 0.01055f
C3773 vdd.n1476 gnd 0.01055f
C3774 vdd.n1477 gnd 0.01055f
C3775 vdd.n1478 gnd 0.008492f
C3776 vdd.n1479 gnd 0.008492f
C3777 vdd.n1480 gnd 0.008492f
C3778 vdd.n1481 gnd 0.01055f
C3779 vdd.n1482 gnd 0.01055f
C3780 vdd.n1483 gnd 0.01055f
C3781 vdd.n1484 gnd 0.008492f
C3782 vdd.n1485 gnd 0.008492f
C3783 vdd.n1486 gnd 0.008492f
C3784 vdd.n1487 gnd 0.01055f
C3785 vdd.n1488 gnd 0.01055f
C3786 vdd.n1489 gnd 0.01055f
C3787 vdd.n1490 gnd 0.008492f
C3788 vdd.n1491 gnd 0.008492f
C3789 vdd.n1492 gnd 0.008492f
C3790 vdd.n1493 gnd 0.01055f
C3791 vdd.n1494 gnd 0.01055f
C3792 vdd.n1495 gnd 0.01055f
C3793 vdd.n1496 gnd 0.008492f
C3794 vdd.n1497 gnd 0.01055f
C3795 vdd.n1498 gnd 2.55536f
C3796 vdd.n1500 gnd 0.026069f
C3797 vdd.n1501 gnd 0.007048f
C3798 vdd.n1502 gnd 0.026069f
C3799 vdd.n1503 gnd 0.025523f
C3800 vdd.n1504 gnd 0.01055f
C3801 vdd.n1505 gnd 0.008492f
C3802 vdd.n1506 gnd 0.01055f
C3803 vdd.n1507 gnd 0.544497f
C3804 vdd.n1508 gnd 0.01055f
C3805 vdd.n1509 gnd 0.008492f
C3806 vdd.n1510 gnd 0.01055f
C3807 vdd.n1511 gnd 0.01055f
C3808 vdd.n1512 gnd 0.01055f
C3809 vdd.n1513 gnd 0.008492f
C3810 vdd.n1514 gnd 0.01055f
C3811 vdd.n1515 gnd 0.986564f
C3812 vdd.n1516 gnd 1.07821f
C3813 vdd.n1517 gnd 0.01055f
C3814 vdd.n1518 gnd 0.008492f
C3815 vdd.n1519 gnd 0.01055f
C3816 vdd.n1520 gnd 0.01055f
C3817 vdd.n1521 gnd 0.01055f
C3818 vdd.n1522 gnd 0.008492f
C3819 vdd.n1523 gnd 0.01055f
C3820 vdd.n1524 gnd 0.630754f
C3821 vdd.n1525 gnd 0.01055f
C3822 vdd.n1526 gnd 0.008492f
C3823 vdd.n1527 gnd 0.01055f
C3824 vdd.n1528 gnd 0.01055f
C3825 vdd.n1529 gnd 0.01055f
C3826 vdd.n1530 gnd 0.008492f
C3827 vdd.n1531 gnd 0.01055f
C3828 vdd.n1532 gnd 0.619972f
C3829 vdd.n1533 gnd 0.81405f
C3830 vdd.n1534 gnd 0.01055f
C3831 vdd.n1535 gnd 0.008492f
C3832 vdd.n1536 gnd 0.01055f
C3833 vdd.n1537 gnd 0.01055f
C3834 vdd.n1538 gnd 0.01055f
C3835 vdd.n1539 gnd 0.008492f
C3836 vdd.n1540 gnd 0.01055f
C3837 vdd.n1541 gnd 0.894916f
C3838 vdd.n1542 gnd 0.01055f
C3839 vdd.n1543 gnd 0.008492f
C3840 vdd.n1544 gnd 0.01055f
C3841 vdd.n1545 gnd 0.01055f
C3842 vdd.n1546 gnd 0.01055f
C3843 vdd.n1547 gnd 0.008492f
C3844 vdd.n1548 gnd 0.01055f
C3845 vdd.t192 gnd 0.539106f
C3846 vdd.n1549 gnd 0.792486f
C3847 vdd.n1550 gnd 0.01055f
C3848 vdd.n1551 gnd 0.008492f
C3849 vdd.n1552 gnd 0.01055f
C3850 vdd.n1553 gnd 0.01055f
C3851 vdd.n1554 gnd 0.01055f
C3852 vdd.n1555 gnd 0.008492f
C3853 vdd.n1556 gnd 0.01055f
C3854 vdd.n1557 gnd 0.60919f
C3855 vdd.n1558 gnd 0.01055f
C3856 vdd.n1559 gnd 0.008492f
C3857 vdd.n1560 gnd 0.01055f
C3858 vdd.n1561 gnd 0.01055f
C3859 vdd.n1562 gnd 0.01055f
C3860 vdd.n1563 gnd 0.008492f
C3861 vdd.n1564 gnd 0.01055f
C3862 vdd.n1565 gnd 0.781704f
C3863 vdd.n1566 gnd 0.652318f
C3864 vdd.n1567 gnd 0.01055f
C3865 vdd.n1568 gnd 0.008492f
C3866 vdd.n1569 gnd 0.01055f
C3867 vdd.n1570 gnd 0.01055f
C3868 vdd.n1571 gnd 0.01055f
C3869 vdd.n1572 gnd 0.008492f
C3870 vdd.n1573 gnd 0.01055f
C3871 vdd.n1574 gnd 0.835614f
C3872 vdd.n1575 gnd 0.01055f
C3873 vdd.n1576 gnd 0.008492f
C3874 vdd.n1577 gnd 0.01055f
C3875 vdd.n1578 gnd 0.01055f
C3876 vdd.n1579 gnd 0.01055f
C3877 vdd.n1580 gnd 0.008492f
C3878 vdd.n1581 gnd 0.01055f
C3879 vdd.t146 gnd 0.539106f
C3880 vdd.n1582 gnd 0.894916f
C3881 vdd.n1583 gnd 0.01055f
C3882 vdd.n1584 gnd 0.008492f
C3883 vdd.n1585 gnd 0.01055f
C3884 vdd.n1586 gnd 0.008109f
C3885 vdd.n1587 gnd 0.00579f
C3886 vdd.n1588 gnd 0.005373f
C3887 vdd.n1589 gnd 0.002972f
C3888 vdd.n1590 gnd 0.006824f
C3889 vdd.n1591 gnd 0.002887f
C3890 vdd.n1592 gnd 0.003057f
C3891 vdd.n1593 gnd 0.005373f
C3892 vdd.n1594 gnd 0.002887f
C3893 vdd.n1595 gnd 0.006824f
C3894 vdd.n1596 gnd 0.003057f
C3895 vdd.n1597 gnd 0.005373f
C3896 vdd.n1598 gnd 0.002887f
C3897 vdd.n1599 gnd 0.005118f
C3898 vdd.n1600 gnd 0.005134f
C3899 vdd.t239 gnd 0.014662f
C3900 vdd.n1601 gnd 0.032622f
C3901 vdd.n1602 gnd 0.169772f
C3902 vdd.n1603 gnd 0.002887f
C3903 vdd.n1604 gnd 0.003057f
C3904 vdd.n1605 gnd 0.006824f
C3905 vdd.n1606 gnd 0.006824f
C3906 vdd.n1607 gnd 0.003057f
C3907 vdd.n1608 gnd 0.002887f
C3908 vdd.n1609 gnd 0.005373f
C3909 vdd.n1610 gnd 0.005373f
C3910 vdd.n1611 gnd 0.002887f
C3911 vdd.n1612 gnd 0.003057f
C3912 vdd.n1613 gnd 0.006824f
C3913 vdd.n1614 gnd 0.006824f
C3914 vdd.n1615 gnd 0.003057f
C3915 vdd.n1616 gnd 0.002887f
C3916 vdd.n1617 gnd 0.005373f
C3917 vdd.n1618 gnd 0.005373f
C3918 vdd.n1619 gnd 0.002887f
C3919 vdd.n1620 gnd 0.003057f
C3920 vdd.n1621 gnd 0.006824f
C3921 vdd.n1622 gnd 0.006824f
C3922 vdd.n1623 gnd 0.016134f
C3923 vdd.n1624 gnd 0.002972f
C3924 vdd.n1625 gnd 0.002887f
C3925 vdd.n1626 gnd 0.013888f
C3926 vdd.n1627 gnd 0.009696f
C3927 vdd.t203 gnd 0.033967f
C3928 vdd.t156 gnd 0.033967f
C3929 vdd.n1628 gnd 0.233448f
C3930 vdd.n1629 gnd 0.183571f
C3931 vdd.t227 gnd 0.033967f
C3932 vdd.t167 gnd 0.033967f
C3933 vdd.n1630 gnd 0.233448f
C3934 vdd.n1631 gnd 0.148141f
C3935 vdd.t275 gnd 0.033967f
C3936 vdd.t297 gnd 0.033967f
C3937 vdd.n1632 gnd 0.233448f
C3938 vdd.n1633 gnd 0.148141f
C3939 vdd.t256 gnd 0.033967f
C3940 vdd.t144 gnd 0.033967f
C3941 vdd.n1634 gnd 0.233448f
C3942 vdd.n1635 gnd 0.148141f
C3943 vdd.t242 gnd 0.033967f
C3944 vdd.t178 gnd 0.033967f
C3945 vdd.n1636 gnd 0.233448f
C3946 vdd.n1637 gnd 0.148141f
C3947 vdd.t286 gnd 0.033967f
C3948 vdd.t210 gnd 0.033967f
C3949 vdd.n1638 gnd 0.233448f
C3950 vdd.n1639 gnd 0.148141f
C3951 vdd.t262 gnd 0.033967f
C3952 vdd.t231 gnd 0.033967f
C3953 vdd.n1640 gnd 0.233448f
C3954 vdd.n1641 gnd 0.148141f
C3955 vdd.t277 gnd 0.033967f
C3956 vdd.t193 gnd 0.033967f
C3957 vdd.n1642 gnd 0.233448f
C3958 vdd.n1643 gnd 0.148141f
C3959 vdd.t293 gnd 0.033967f
C3960 vdd.t221 gnd 0.033967f
C3961 vdd.n1644 gnd 0.233448f
C3962 vdd.n1645 gnd 0.148141f
C3963 vdd.n1646 gnd 0.00579f
C3964 vdd.n1647 gnd 0.005373f
C3965 vdd.n1648 gnd 0.002972f
C3966 vdd.n1649 gnd 0.006824f
C3967 vdd.n1650 gnd 0.002887f
C3968 vdd.n1651 gnd 0.003057f
C3969 vdd.n1652 gnd 0.005373f
C3970 vdd.n1653 gnd 0.002887f
C3971 vdd.n1654 gnd 0.006824f
C3972 vdd.n1655 gnd 0.003057f
C3973 vdd.n1656 gnd 0.005373f
C3974 vdd.n1657 gnd 0.002887f
C3975 vdd.n1658 gnd 0.005118f
C3976 vdd.n1659 gnd 0.005134f
C3977 vdd.t246 gnd 0.014662f
C3978 vdd.n1660 gnd 0.032622f
C3979 vdd.n1661 gnd 0.169772f
C3980 vdd.n1662 gnd 0.002887f
C3981 vdd.n1663 gnd 0.003057f
C3982 vdd.n1664 gnd 0.006824f
C3983 vdd.n1665 gnd 0.006824f
C3984 vdd.n1666 gnd 0.003057f
C3985 vdd.n1667 gnd 0.002887f
C3986 vdd.n1668 gnd 0.005373f
C3987 vdd.n1669 gnd 0.005373f
C3988 vdd.n1670 gnd 0.002887f
C3989 vdd.n1671 gnd 0.003057f
C3990 vdd.n1672 gnd 0.006824f
C3991 vdd.n1673 gnd 0.006824f
C3992 vdd.n1674 gnd 0.003057f
C3993 vdd.n1675 gnd 0.002887f
C3994 vdd.n1676 gnd 0.005373f
C3995 vdd.n1677 gnd 0.005373f
C3996 vdd.n1678 gnd 0.002887f
C3997 vdd.n1679 gnd 0.003057f
C3998 vdd.n1680 gnd 0.006824f
C3999 vdd.n1681 gnd 0.006824f
C4000 vdd.n1682 gnd 0.016134f
C4001 vdd.n1683 gnd 0.002972f
C4002 vdd.n1684 gnd 0.002887f
C4003 vdd.n1685 gnd 0.013888f
C4004 vdd.n1686 gnd 0.009391f
C4005 vdd.n1687 gnd 0.110218f
C4006 vdd.n1688 gnd 0.00579f
C4007 vdd.n1689 gnd 0.005373f
C4008 vdd.n1690 gnd 0.002972f
C4009 vdd.n1691 gnd 0.006824f
C4010 vdd.n1692 gnd 0.002887f
C4011 vdd.n1693 gnd 0.003057f
C4012 vdd.n1694 gnd 0.005373f
C4013 vdd.n1695 gnd 0.002887f
C4014 vdd.n1696 gnd 0.006824f
C4015 vdd.n1697 gnd 0.003057f
C4016 vdd.n1698 gnd 0.005373f
C4017 vdd.n1699 gnd 0.002887f
C4018 vdd.n1700 gnd 0.005118f
C4019 vdd.n1701 gnd 0.005134f
C4020 vdd.t282 gnd 0.014662f
C4021 vdd.n1702 gnd 0.032622f
C4022 vdd.n1703 gnd 0.169772f
C4023 vdd.n1704 gnd 0.002887f
C4024 vdd.n1705 gnd 0.003057f
C4025 vdd.n1706 gnd 0.006824f
C4026 vdd.n1707 gnd 0.006824f
C4027 vdd.n1708 gnd 0.003057f
C4028 vdd.n1709 gnd 0.002887f
C4029 vdd.n1710 gnd 0.005373f
C4030 vdd.n1711 gnd 0.005373f
C4031 vdd.n1712 gnd 0.002887f
C4032 vdd.n1713 gnd 0.003057f
C4033 vdd.n1714 gnd 0.006824f
C4034 vdd.n1715 gnd 0.006824f
C4035 vdd.n1716 gnd 0.003057f
C4036 vdd.n1717 gnd 0.002887f
C4037 vdd.n1718 gnd 0.005373f
C4038 vdd.n1719 gnd 0.005373f
C4039 vdd.n1720 gnd 0.002887f
C4040 vdd.n1721 gnd 0.003057f
C4041 vdd.n1722 gnd 0.006824f
C4042 vdd.n1723 gnd 0.006824f
C4043 vdd.n1724 gnd 0.016134f
C4044 vdd.n1725 gnd 0.002972f
C4045 vdd.n1726 gnd 0.002887f
C4046 vdd.n1727 gnd 0.013888f
C4047 vdd.n1728 gnd 0.009696f
C4048 vdd.t252 gnd 0.033967f
C4049 vdd.t184 gnd 0.033967f
C4050 vdd.n1729 gnd 0.233448f
C4051 vdd.n1730 gnd 0.183571f
C4052 vdd.t180 gnd 0.033967f
C4053 vdd.t253 gnd 0.033967f
C4054 vdd.n1731 gnd 0.233448f
C4055 vdd.n1732 gnd 0.148141f
C4056 vdd.t237 gnd 0.033967f
C4057 vdd.t233 gnd 0.033967f
C4058 vdd.n1733 gnd 0.233448f
C4059 vdd.n1734 gnd 0.148141f
C4060 vdd.t176 gnd 0.033967f
C4061 vdd.t154 gnd 0.033967f
C4062 vdd.n1735 gnd 0.233448f
C4063 vdd.n1736 gnd 0.148141f
C4064 vdd.t147 gnd 0.033967f
C4065 vdd.t228 gnd 0.033967f
C4066 vdd.n1737 gnd 0.233448f
C4067 vdd.n1738 gnd 0.148141f
C4068 vdd.t205 gnd 0.033967f
C4069 vdd.t149 gnd 0.033967f
C4070 vdd.n1739 gnd 0.233448f
C4071 vdd.n1740 gnd 0.148141f
C4072 vdd.t140 gnd 0.033967f
C4073 vdd.t257 gnd 0.033967f
C4074 vdd.n1741 gnd 0.233448f
C4075 vdd.n1742 gnd 0.148141f
C4076 vdd.t241 gnd 0.033967f
C4077 vdd.t195 gnd 0.033967f
C4078 vdd.n1743 gnd 0.233448f
C4079 vdd.n1744 gnd 0.148141f
C4080 vdd.t182 gnd 0.033967f
C4081 vdd.t283 gnd 0.033967f
C4082 vdd.n1745 gnd 0.233448f
C4083 vdd.n1746 gnd 0.148141f
C4084 vdd.n1747 gnd 0.00579f
C4085 vdd.n1748 gnd 0.005373f
C4086 vdd.n1749 gnd 0.002972f
C4087 vdd.n1750 gnd 0.006824f
C4088 vdd.n1751 gnd 0.002887f
C4089 vdd.n1752 gnd 0.003057f
C4090 vdd.n1753 gnd 0.005373f
C4091 vdd.n1754 gnd 0.002887f
C4092 vdd.n1755 gnd 0.006824f
C4093 vdd.n1756 gnd 0.003057f
C4094 vdd.n1757 gnd 0.005373f
C4095 vdd.n1758 gnd 0.002887f
C4096 vdd.n1759 gnd 0.005118f
C4097 vdd.n1760 gnd 0.005134f
C4098 vdd.t235 gnd 0.014662f
C4099 vdd.n1761 gnd 0.032622f
C4100 vdd.n1762 gnd 0.169772f
C4101 vdd.n1763 gnd 0.002887f
C4102 vdd.n1764 gnd 0.003057f
C4103 vdd.n1765 gnd 0.006824f
C4104 vdd.n1766 gnd 0.006824f
C4105 vdd.n1767 gnd 0.003057f
C4106 vdd.n1768 gnd 0.002887f
C4107 vdd.n1769 gnd 0.005373f
C4108 vdd.n1770 gnd 0.005373f
C4109 vdd.n1771 gnd 0.002887f
C4110 vdd.n1772 gnd 0.003057f
C4111 vdd.n1773 gnd 0.006824f
C4112 vdd.n1774 gnd 0.006824f
C4113 vdd.n1775 gnd 0.003057f
C4114 vdd.n1776 gnd 0.002887f
C4115 vdd.n1777 gnd 0.005373f
C4116 vdd.n1778 gnd 0.005373f
C4117 vdd.n1779 gnd 0.002887f
C4118 vdd.n1780 gnd 0.003057f
C4119 vdd.n1781 gnd 0.006824f
C4120 vdd.n1782 gnd 0.006824f
C4121 vdd.n1783 gnd 0.016134f
C4122 vdd.n1784 gnd 0.002972f
C4123 vdd.n1785 gnd 0.002887f
C4124 vdd.n1786 gnd 0.013888f
C4125 vdd.n1787 gnd 0.009391f
C4126 vdd.n1788 gnd 0.065568f
C4127 vdd.n1789 gnd 0.23626f
C4128 vdd.n1790 gnd 0.00579f
C4129 vdd.n1791 gnd 0.005373f
C4130 vdd.n1792 gnd 0.002972f
C4131 vdd.n1793 gnd 0.006824f
C4132 vdd.n1794 gnd 0.002887f
C4133 vdd.n1795 gnd 0.003057f
C4134 vdd.n1796 gnd 0.005373f
C4135 vdd.n1797 gnd 0.002887f
C4136 vdd.n1798 gnd 0.006824f
C4137 vdd.n1799 gnd 0.003057f
C4138 vdd.n1800 gnd 0.005373f
C4139 vdd.n1801 gnd 0.002887f
C4140 vdd.n1802 gnd 0.005118f
C4141 vdd.n1803 gnd 0.005134f
C4142 vdd.t298 gnd 0.014662f
C4143 vdd.n1804 gnd 0.032622f
C4144 vdd.n1805 gnd 0.169772f
C4145 vdd.n1806 gnd 0.002887f
C4146 vdd.n1807 gnd 0.003057f
C4147 vdd.n1808 gnd 0.006824f
C4148 vdd.n1809 gnd 0.006824f
C4149 vdd.n1810 gnd 0.003057f
C4150 vdd.n1811 gnd 0.002887f
C4151 vdd.n1812 gnd 0.005373f
C4152 vdd.n1813 gnd 0.005373f
C4153 vdd.n1814 gnd 0.002887f
C4154 vdd.n1815 gnd 0.003057f
C4155 vdd.n1816 gnd 0.006824f
C4156 vdd.n1817 gnd 0.006824f
C4157 vdd.n1818 gnd 0.003057f
C4158 vdd.n1819 gnd 0.002887f
C4159 vdd.n1820 gnd 0.005373f
C4160 vdd.n1821 gnd 0.005373f
C4161 vdd.n1822 gnd 0.002887f
C4162 vdd.n1823 gnd 0.003057f
C4163 vdd.n1824 gnd 0.006824f
C4164 vdd.n1825 gnd 0.006824f
C4165 vdd.n1826 gnd 0.016134f
C4166 vdd.n1827 gnd 0.002972f
C4167 vdd.n1828 gnd 0.002887f
C4168 vdd.n1829 gnd 0.013888f
C4169 vdd.n1830 gnd 0.009696f
C4170 vdd.t264 gnd 0.033967f
C4171 vdd.t211 gnd 0.033967f
C4172 vdd.n1831 gnd 0.233448f
C4173 vdd.n1832 gnd 0.183571f
C4174 vdd.t206 gnd 0.033967f
C4175 vdd.t266 gnd 0.033967f
C4176 vdd.n1833 gnd 0.233448f
C4177 vdd.n1834 gnd 0.148141f
C4178 vdd.t250 gnd 0.033967f
C4179 vdd.t248 gnd 0.033967f
C4180 vdd.n1835 gnd 0.233448f
C4181 vdd.n1836 gnd 0.148141f
C4182 vdd.t201 gnd 0.033967f
C4183 vdd.t172 gnd 0.033967f
C4184 vdd.n1837 gnd 0.233448f
C4185 vdd.n1838 gnd 0.148141f
C4186 vdd.t170 gnd 0.033967f
C4187 vdd.t247 gnd 0.033967f
C4188 vdd.n1839 gnd 0.233448f
C4189 vdd.n1840 gnd 0.148141f
C4190 vdd.t222 gnd 0.033967f
C4191 vdd.t171 gnd 0.033967f
C4192 vdd.n1841 gnd 0.233448f
C4193 vdd.n1842 gnd 0.148141f
C4194 vdd.t165 gnd 0.033967f
C4195 vdd.t267 gnd 0.033967f
C4196 vdd.n1843 gnd 0.233448f
C4197 vdd.n1844 gnd 0.148141f
C4198 vdd.t265 gnd 0.033967f
C4199 vdd.t215 gnd 0.033967f
C4200 vdd.n1845 gnd 0.233448f
C4201 vdd.n1846 gnd 0.148141f
C4202 vdd.t207 gnd 0.033967f
C4203 vdd.t294 gnd 0.033967f
C4204 vdd.n1847 gnd 0.233448f
C4205 vdd.n1848 gnd 0.148141f
C4206 vdd.n1849 gnd 0.00579f
C4207 vdd.n1850 gnd 0.005373f
C4208 vdd.n1851 gnd 0.002972f
C4209 vdd.n1852 gnd 0.006824f
C4210 vdd.n1853 gnd 0.002887f
C4211 vdd.n1854 gnd 0.003057f
C4212 vdd.n1855 gnd 0.005373f
C4213 vdd.n1856 gnd 0.002887f
C4214 vdd.n1857 gnd 0.006824f
C4215 vdd.n1858 gnd 0.003057f
C4216 vdd.n1859 gnd 0.005373f
C4217 vdd.n1860 gnd 0.002887f
C4218 vdd.n1861 gnd 0.005118f
C4219 vdd.n1862 gnd 0.005134f
C4220 vdd.t249 gnd 0.014662f
C4221 vdd.n1863 gnd 0.032622f
C4222 vdd.n1864 gnd 0.169772f
C4223 vdd.n1865 gnd 0.002887f
C4224 vdd.n1866 gnd 0.003057f
C4225 vdd.n1867 gnd 0.006824f
C4226 vdd.n1868 gnd 0.006824f
C4227 vdd.n1869 gnd 0.003057f
C4228 vdd.n1870 gnd 0.002887f
C4229 vdd.n1871 gnd 0.005373f
C4230 vdd.n1872 gnd 0.005373f
C4231 vdd.n1873 gnd 0.002887f
C4232 vdd.n1874 gnd 0.003057f
C4233 vdd.n1875 gnd 0.006824f
C4234 vdd.n1876 gnd 0.006824f
C4235 vdd.n1877 gnd 0.003057f
C4236 vdd.n1878 gnd 0.002887f
C4237 vdd.n1879 gnd 0.005373f
C4238 vdd.n1880 gnd 0.005373f
C4239 vdd.n1881 gnd 0.002887f
C4240 vdd.n1882 gnd 0.003057f
C4241 vdd.n1883 gnd 0.006824f
C4242 vdd.n1884 gnd 0.006824f
C4243 vdd.n1885 gnd 0.016134f
C4244 vdd.n1886 gnd 0.002972f
C4245 vdd.n1887 gnd 0.002887f
C4246 vdd.n1888 gnd 0.013888f
C4247 vdd.n1889 gnd 0.009391f
C4248 vdd.n1890 gnd 0.065568f
C4249 vdd.n1891 gnd 0.270467f
C4250 vdd.n1892 gnd 2.96492f
C4251 vdd.n1893 gnd 0.622309f
C4252 vdd.n1894 gnd 0.008109f
C4253 vdd.n1895 gnd 0.008492f
C4254 vdd.n1896 gnd 0.01055f
C4255 vdd.n1897 gnd 0.770922f
C4256 vdd.n1898 gnd 0.01055f
C4257 vdd.n1899 gnd 0.008492f
C4258 vdd.n1900 gnd 0.01055f
C4259 vdd.n1901 gnd 0.01055f
C4260 vdd.n1902 gnd 0.01055f
C4261 vdd.n1903 gnd 0.008492f
C4262 vdd.n1904 gnd 0.01055f
C4263 vdd.n1905 gnd 0.894916f
C4264 vdd.t175 gnd 0.539106f
C4265 vdd.n1906 gnd 0.587625f
C4266 vdd.n1907 gnd 0.01055f
C4267 vdd.n1908 gnd 0.008492f
C4268 vdd.n1909 gnd 0.01055f
C4269 vdd.n1910 gnd 0.01055f
C4270 vdd.n1911 gnd 0.01055f
C4271 vdd.n1912 gnd 0.008492f
C4272 vdd.n1913 gnd 0.01055f
C4273 vdd.n1914 gnd 0.673882f
C4274 vdd.n1915 gnd 0.01055f
C4275 vdd.n1916 gnd 0.008492f
C4276 vdd.n1917 gnd 0.01055f
C4277 vdd.n1918 gnd 0.01055f
C4278 vdd.n1919 gnd 0.01055f
C4279 vdd.n1920 gnd 0.008492f
C4280 vdd.n1921 gnd 0.01055f
C4281 vdd.n1922 gnd 0.576843f
C4282 vdd.n1923 gnd 0.857178f
C4283 vdd.n1924 gnd 0.01055f
C4284 vdd.n1925 gnd 0.008492f
C4285 vdd.n1926 gnd 0.01055f
C4286 vdd.n1927 gnd 0.01055f
C4287 vdd.n1928 gnd 0.01055f
C4288 vdd.n1929 gnd 0.008492f
C4289 vdd.n1930 gnd 0.01055f
C4290 vdd.n1931 gnd 0.894916f
C4291 vdd.n1932 gnd 0.01055f
C4292 vdd.n1933 gnd 0.008492f
C4293 vdd.n1934 gnd 0.01055f
C4294 vdd.n1935 gnd 0.01055f
C4295 vdd.n1936 gnd 0.01055f
C4296 vdd.n1937 gnd 0.008492f
C4297 vdd.n1938 gnd 0.01055f
C4298 vdd.t166 gnd 0.539106f
C4299 vdd.n1939 gnd 0.749357f
C4300 vdd.n1940 gnd 0.01055f
C4301 vdd.n1941 gnd 0.008492f
C4302 vdd.n1942 gnd 0.01055f
C4303 vdd.n1943 gnd 0.01055f
C4304 vdd.n1944 gnd 0.01055f
C4305 vdd.n1945 gnd 0.008492f
C4306 vdd.n1946 gnd 0.01055f
C4307 vdd.n1947 gnd 0.566061f
C4308 vdd.n1948 gnd 0.01055f
C4309 vdd.n1949 gnd 0.008492f
C4310 vdd.n1950 gnd 0.01055f
C4311 vdd.n1951 gnd 0.01055f
C4312 vdd.n1952 gnd 0.01055f
C4313 vdd.n1953 gnd 0.008492f
C4314 vdd.n1954 gnd 0.01055f
C4315 vdd.n1955 gnd 0.738575f
C4316 vdd.n1956 gnd 0.695447f
C4317 vdd.n1957 gnd 0.01055f
C4318 vdd.n1958 gnd 0.008492f
C4319 vdd.n1959 gnd 0.01055f
C4320 vdd.n1960 gnd 0.01055f
C4321 vdd.n1961 gnd 0.01055f
C4322 vdd.n1962 gnd 0.008492f
C4323 vdd.n1963 gnd 0.01055f
C4324 vdd.n1964 gnd 0.878743f
C4325 vdd.n1965 gnd 0.01055f
C4326 vdd.n1966 gnd 0.008492f
C4327 vdd.n1967 gnd 0.01055f
C4328 vdd.n1968 gnd 0.01055f
C4329 vdd.n1969 gnd 0.025523f
C4330 vdd.n1970 gnd 0.01055f
C4331 vdd.n1971 gnd 0.01055f
C4332 vdd.n1972 gnd 0.008492f
C4333 vdd.n1973 gnd 0.01055f
C4334 vdd.n1974 gnd 0.652318f
C4335 vdd.n1975 gnd 1.07821f
C4336 vdd.n1976 gnd 0.01055f
C4337 vdd.n1977 gnd 0.008492f
C4338 vdd.n1978 gnd 0.01055f
C4339 vdd.n1979 gnd 0.01055f
C4340 vdd.n1980 gnd 0.009073f
C4341 vdd.n1981 gnd 0.008492f
C4342 vdd.n1983 gnd 0.01055f
C4343 vdd.n1985 gnd 0.008492f
C4344 vdd.n1986 gnd 0.01055f
C4345 vdd.n1987 gnd 0.008492f
C4346 vdd.n1989 gnd 0.01055f
C4347 vdd.n1990 gnd 0.008492f
C4348 vdd.n1991 gnd 0.01055f
C4349 vdd.n1992 gnd 0.01055f
C4350 vdd.n1993 gnd 0.01055f
C4351 vdd.n1994 gnd 0.01055f
C4352 vdd.n1995 gnd 0.01055f
C4353 vdd.n1996 gnd 0.008492f
C4354 vdd.n1998 gnd 0.01055f
C4355 vdd.n1999 gnd 0.01055f
C4356 vdd.n2000 gnd 0.01055f
C4357 vdd.n2001 gnd 0.01055f
C4358 vdd.n2002 gnd 0.01055f
C4359 vdd.n2003 gnd 0.008492f
C4360 vdd.n2005 gnd 0.01055f
C4361 vdd.n2006 gnd 0.01055f
C4362 vdd.n2007 gnd 0.01055f
C4363 vdd.n2008 gnd 0.01055f
C4364 vdd.n2009 gnd 0.007091f
C4365 vdd.t122 gnd 0.129799f
C4366 vdd.t121 gnd 0.138719f
C4367 vdd.t120 gnd 0.169516f
C4368 vdd.n2010 gnd 0.217295f
C4369 vdd.n2011 gnd 0.182567f
C4370 vdd.n2013 gnd 0.01055f
C4371 vdd.n2014 gnd 0.01055f
C4372 vdd.n2015 gnd 0.008492f
C4373 vdd.n2016 gnd 0.01055f
C4374 vdd.n2018 gnd 0.01055f
C4375 vdd.n2019 gnd 0.01055f
C4376 vdd.n2020 gnd 0.01055f
C4377 vdd.n2021 gnd 0.01055f
C4378 vdd.n2022 gnd 0.008492f
C4379 vdd.n2024 gnd 0.01055f
C4380 vdd.n2025 gnd 0.01055f
C4381 vdd.n2026 gnd 0.01055f
C4382 vdd.n2027 gnd 0.01055f
C4383 vdd.n2028 gnd 0.01055f
C4384 vdd.n2029 gnd 0.008492f
C4385 vdd.n2031 gnd 0.01055f
C4386 vdd.n2032 gnd 0.01055f
C4387 vdd.n2033 gnd 0.01055f
C4388 vdd.n2034 gnd 0.01055f
C4389 vdd.n2035 gnd 0.01055f
C4390 vdd.n2036 gnd 0.008492f
C4391 vdd.n2038 gnd 0.01055f
C4392 vdd.n2039 gnd 0.01055f
C4393 vdd.n2040 gnd 0.01055f
C4394 vdd.n2041 gnd 0.01055f
C4395 vdd.n2042 gnd 0.01055f
C4396 vdd.n2043 gnd 0.008492f
C4397 vdd.n2045 gnd 0.01055f
C4398 vdd.n2046 gnd 0.01055f
C4399 vdd.n2047 gnd 0.01055f
C4400 vdd.n2048 gnd 0.01055f
C4401 vdd.n2049 gnd 0.008407f
C4402 vdd.t101 gnd 0.129799f
C4403 vdd.t100 gnd 0.138719f
C4404 vdd.t99 gnd 0.169516f
C4405 vdd.n2050 gnd 0.217295f
C4406 vdd.n2051 gnd 0.182567f
C4407 vdd.n2053 gnd 0.01055f
C4408 vdd.n2054 gnd 0.01055f
C4409 vdd.n2055 gnd 0.008492f
C4410 vdd.n2056 gnd 0.01055f
C4411 vdd.n2058 gnd 0.01055f
C4412 vdd.n2059 gnd 0.01055f
C4413 vdd.n2060 gnd 0.01055f
C4414 vdd.n2061 gnd 0.01055f
C4415 vdd.n2062 gnd 0.008492f
C4416 vdd.n2064 gnd 0.01055f
C4417 vdd.n2065 gnd 0.01055f
C4418 vdd.n2066 gnd 0.01055f
C4419 vdd.n2067 gnd 0.01055f
C4420 vdd.n2068 gnd 0.01055f
C4421 vdd.n2069 gnd 0.008492f
C4422 vdd.n2071 gnd 0.01055f
C4423 vdd.n2072 gnd 0.01055f
C4424 vdd.n2073 gnd 0.01055f
C4425 vdd.n2074 gnd 0.01055f
C4426 vdd.n2075 gnd 0.01055f
C4427 vdd.n2076 gnd 0.01055f
C4428 vdd.n2077 gnd 0.008492f
C4429 vdd.n2079 gnd 0.01055f
C4430 vdd.n2081 gnd 0.01055f
C4431 vdd.n2082 gnd 0.008492f
C4432 vdd.n2083 gnd 0.008492f
C4433 vdd.n2084 gnd 0.01055f
C4434 vdd.n2086 gnd 0.01055f
C4435 vdd.n2087 gnd 0.008492f
C4436 vdd.n2088 gnd 0.008492f
C4437 vdd.n2089 gnd 0.01055f
C4438 vdd.n2091 gnd 0.01055f
C4439 vdd.n2092 gnd 0.01055f
C4440 vdd.n2093 gnd 0.008492f
C4441 vdd.n2094 gnd 0.008492f
C4442 vdd.n2095 gnd 0.008492f
C4443 vdd.n2096 gnd 0.01055f
C4444 vdd.n2098 gnd 0.01055f
C4445 vdd.n2099 gnd 0.01055f
C4446 vdd.n2100 gnd 0.008492f
C4447 vdd.n2101 gnd 0.008492f
C4448 vdd.n2102 gnd 0.008492f
C4449 vdd.n2103 gnd 0.01055f
C4450 vdd.n2105 gnd 0.01055f
C4451 vdd.n2106 gnd 0.01055f
C4452 vdd.n2107 gnd 0.008492f
C4453 vdd.n2108 gnd 0.008492f
C4454 vdd.n2109 gnd 0.008492f
C4455 vdd.n2110 gnd 0.01055f
C4456 vdd.n2112 gnd 0.01055f
C4457 vdd.n2113 gnd 0.01055f
C4458 vdd.n2114 gnd 0.008492f
C4459 vdd.n2115 gnd 0.01055f
C4460 vdd.n2116 gnd 0.01055f
C4461 vdd.n2117 gnd 0.01055f
C4462 vdd.n2118 gnd 0.017323f
C4463 vdd.n2119 gnd 0.005774f
C4464 vdd.n2120 gnd 0.008492f
C4465 vdd.n2121 gnd 0.01055f
C4466 vdd.n2123 gnd 0.01055f
C4467 vdd.n2124 gnd 0.01055f
C4468 vdd.n2125 gnd 0.008492f
C4469 vdd.n2126 gnd 0.008492f
C4470 vdd.n2127 gnd 0.008492f
C4471 vdd.n2128 gnd 0.01055f
C4472 vdd.n2130 gnd 0.01055f
C4473 vdd.n2131 gnd 0.01055f
C4474 vdd.n2132 gnd 0.008492f
C4475 vdd.n2133 gnd 0.008492f
C4476 vdd.n2134 gnd 0.008492f
C4477 vdd.n2135 gnd 0.01055f
C4478 vdd.n2137 gnd 0.01055f
C4479 vdd.n2138 gnd 0.01055f
C4480 vdd.n2139 gnd 0.008492f
C4481 vdd.n2140 gnd 0.008492f
C4482 vdd.n2141 gnd 0.008492f
C4483 vdd.n2142 gnd 0.01055f
C4484 vdd.n2144 gnd 0.01055f
C4485 vdd.n2145 gnd 0.01055f
C4486 vdd.n2146 gnd 0.008492f
C4487 vdd.n2147 gnd 0.008492f
C4488 vdd.n2148 gnd 0.008492f
C4489 vdd.n2149 gnd 0.01055f
C4490 vdd.n2151 gnd 0.01055f
C4491 vdd.n2152 gnd 0.01055f
C4492 vdd.n2153 gnd 0.008492f
C4493 vdd.n2154 gnd 0.01055f
C4494 vdd.n2155 gnd 0.01055f
C4495 vdd.n2156 gnd 0.01055f
C4496 vdd.n2157 gnd 0.017323f
C4497 vdd.n2158 gnd 0.007091f
C4498 vdd.n2159 gnd 0.008492f
C4499 vdd.n2160 gnd 0.01055f
C4500 vdd.n2162 gnd 0.01055f
C4501 vdd.n2163 gnd 0.01055f
C4502 vdd.n2164 gnd 0.008492f
C4503 vdd.n2165 gnd 0.008492f
C4504 vdd.n2166 gnd 0.008492f
C4505 vdd.n2167 gnd 0.01055f
C4506 vdd.n2169 gnd 0.01055f
C4507 vdd.n2170 gnd 0.01055f
C4508 vdd.n2171 gnd 0.008492f
C4509 vdd.n2172 gnd 0.008492f
C4510 vdd.n2173 gnd 0.008492f
C4511 vdd.n2174 gnd 0.01055f
C4512 vdd.n2176 gnd 0.01055f
C4513 vdd.n2177 gnd 0.01055f
C4514 vdd.n2179 gnd 0.01055f
C4515 vdd.n2180 gnd 0.008492f
C4516 vdd.n2181 gnd 0.006752f
C4517 vdd.n2182 gnd 0.95976f
C4518 vdd.n2184 gnd 0.008492f
C4519 vdd.n2185 gnd 0.008492f
C4520 vdd.n2186 gnd 0.01055f
C4521 vdd.n2188 gnd 0.01055f
C4522 vdd.n2189 gnd 0.01055f
C4523 vdd.n2190 gnd 0.008492f
C4524 vdd.n2191 gnd 0.007048f
C4525 vdd.n2192 gnd 0.026069f
C4526 vdd.n2193 gnd 0.025523f
C4527 vdd.n2194 gnd 0.007048f
C4528 vdd.n2195 gnd 0.025523f
C4529 vdd.n2196 gnd 1.48254f
C4530 vdd.n2197 gnd 0.025523f
C4531 vdd.n2198 gnd 0.026069f
C4532 vdd.n2199 gnd 0.004034f
C4533 vdd.t92 gnd 0.129799f
C4534 vdd.t91 gnd 0.138719f
C4535 vdd.t89 gnd 0.169516f
C4536 vdd.n2200 gnd 0.217295f
C4537 vdd.n2201 gnd 0.182567f
C4538 vdd.n2202 gnd 0.013078f
C4539 vdd.n2203 gnd 0.004458f
C4540 vdd.n2204 gnd 0.009073f
C4541 vdd.n2205 gnd 0.95976f
C4542 vdd.n2206 gnd 0.037749f
C4543 vdd.n2207 gnd 0.007174f
C4544 vdd.n2208 gnd 0.007174f
C4545 vdd.n2209 gnd 0.007174f
C4546 vdd.n2210 gnd 0.007174f
C4547 vdd.n2211 gnd 0.007174f
C4548 vdd.n2212 gnd 0.007174f
C4549 vdd.n2213 gnd 0.007174f
C4550 vdd.n2214 gnd 0.007174f
C4551 vdd.n2216 gnd 0.007174f
C4552 vdd.n2218 gnd 0.007174f
C4553 vdd.n2219 gnd 0.007174f
C4554 vdd.n2220 gnd 0.007174f
C4555 vdd.n2221 gnd 0.007174f
C4556 vdd.n2222 gnd 0.007174f
C4557 vdd.n2224 gnd 0.007174f
C4558 vdd.n2226 gnd 0.007174f
C4559 vdd.n2227 gnd 0.007174f
C4560 vdd.n2228 gnd 0.007174f
C4561 vdd.n2229 gnd 0.007174f
C4562 vdd.n2230 gnd 0.007174f
C4563 vdd.n2232 gnd 0.007174f
C4564 vdd.n2234 gnd 0.007174f
C4565 vdd.n2235 gnd 0.007174f
C4566 vdd.n2236 gnd 0.007174f
C4567 vdd.n2237 gnd 0.007174f
C4568 vdd.n2238 gnd 0.007174f
C4569 vdd.n2240 gnd 0.007174f
C4570 vdd.n2242 gnd 0.007174f
C4571 vdd.n2243 gnd 0.007174f
C4572 vdd.n2244 gnd 0.007174f
C4573 vdd.n2245 gnd 0.007174f
C4574 vdd.n2246 gnd 0.007174f
C4575 vdd.n2248 gnd 0.007174f
C4576 vdd.n2250 gnd 0.007174f
C4577 vdd.n2251 gnd 0.007174f
C4578 vdd.n2252 gnd 0.007174f
C4579 vdd.n2253 gnd 0.007174f
C4580 vdd.n2254 gnd 0.007174f
C4581 vdd.n2256 gnd 0.007174f
C4582 vdd.n2258 gnd 0.007174f
C4583 vdd.n2259 gnd 0.007174f
C4584 vdd.n2260 gnd 0.007174f
C4585 vdd.n2261 gnd 0.007174f
C4586 vdd.n2262 gnd 0.007174f
C4587 vdd.n2264 gnd 0.007174f
C4588 vdd.n2266 gnd 0.007174f
C4589 vdd.n2267 gnd 0.007174f
C4590 vdd.n2268 gnd 0.007174f
C4591 vdd.n2269 gnd 0.007174f
C4592 vdd.n2270 gnd 0.007174f
C4593 vdd.n2272 gnd 0.007174f
C4594 vdd.n2274 gnd 0.007174f
C4595 vdd.n2275 gnd 0.007174f
C4596 vdd.n2276 gnd 0.005223f
C4597 vdd.n2277 gnd 0.010253f
C4598 vdd.n2278 gnd 0.005539f
C4599 vdd.n2279 gnd 0.007174f
C4600 vdd.n2281 gnd 0.007174f
C4601 vdd.n2282 gnd 0.016536f
C4602 vdd.n2283 gnd 0.016536f
C4603 vdd.n2284 gnd 0.015538f
C4604 vdd.n2285 gnd 0.007174f
C4605 vdd.n2286 gnd 0.007174f
C4606 vdd.n2287 gnd 0.007174f
C4607 vdd.n2288 gnd 0.007174f
C4608 vdd.n2289 gnd 0.007174f
C4609 vdd.n2290 gnd 0.007174f
C4610 vdd.n2291 gnd 0.007174f
C4611 vdd.n2292 gnd 0.007174f
C4612 vdd.n2293 gnd 0.007174f
C4613 vdd.n2294 gnd 0.007174f
C4614 vdd.n2295 gnd 0.007174f
C4615 vdd.n2296 gnd 0.007174f
C4616 vdd.n2297 gnd 0.007174f
C4617 vdd.n2298 gnd 0.007174f
C4618 vdd.n2299 gnd 0.007174f
C4619 vdd.n2300 gnd 0.007174f
C4620 vdd.n2301 gnd 0.007174f
C4621 vdd.n2302 gnd 0.007174f
C4622 vdd.n2303 gnd 0.007174f
C4623 vdd.n2304 gnd 0.007174f
C4624 vdd.n2305 gnd 0.007174f
C4625 vdd.n2306 gnd 0.007174f
C4626 vdd.n2307 gnd 0.007174f
C4627 vdd.n2308 gnd 0.007174f
C4628 vdd.n2309 gnd 0.007174f
C4629 vdd.n2310 gnd 0.007174f
C4630 vdd.n2311 gnd 0.007174f
C4631 vdd.n2312 gnd 0.007174f
C4632 vdd.n2313 gnd 0.007174f
C4633 vdd.n2314 gnd 0.007174f
C4634 vdd.n2315 gnd 0.007174f
C4635 vdd.n2316 gnd 0.007174f
C4636 vdd.n2317 gnd 0.007174f
C4637 vdd.n2318 gnd 0.007174f
C4638 vdd.n2319 gnd 0.007174f
C4639 vdd.n2320 gnd 0.007174f
C4640 vdd.n2321 gnd 0.007174f
C4641 vdd.n2322 gnd 0.007174f
C4642 vdd.n2323 gnd 0.007174f
C4643 vdd.n2324 gnd 0.007174f
C4644 vdd.n2325 gnd 0.007174f
C4645 vdd.n2326 gnd 0.007174f
C4646 vdd.n2327 gnd 0.007174f
C4647 vdd.n2328 gnd 0.007174f
C4648 vdd.n2329 gnd 0.007174f
C4649 vdd.n2330 gnd 0.007174f
C4650 vdd.n2331 gnd 0.007174f
C4651 vdd.n2332 gnd 0.007174f
C4652 vdd.n2333 gnd 0.007174f
C4653 vdd.n2334 gnd 0.436676f
C4654 vdd.n2335 gnd 0.007174f
C4655 vdd.n2336 gnd 0.007174f
C4656 vdd.n2337 gnd 0.007174f
C4657 vdd.n2338 gnd 0.007174f
C4658 vdd.n2339 gnd 0.007174f
C4659 vdd.n2340 gnd 0.007174f
C4660 vdd.n2341 gnd 0.007174f
C4661 vdd.n2342 gnd 0.007174f
C4662 vdd.n2343 gnd 0.007174f
C4663 vdd.n2344 gnd 0.007174f
C4664 vdd.n2345 gnd 0.007174f
C4665 vdd.n2346 gnd 0.6631f
C4666 vdd.n2347 gnd 0.007174f
C4667 vdd.n2348 gnd 0.007174f
C4668 vdd.n2349 gnd 0.007174f
C4669 vdd.n2350 gnd 0.007174f
C4670 vdd.n2351 gnd 0.007174f
C4671 vdd.n2352 gnd 0.007174f
C4672 vdd.n2353 gnd 0.007174f
C4673 vdd.n2354 gnd 0.007174f
C4674 vdd.n2355 gnd 0.007174f
C4675 vdd.n2356 gnd 0.007174f
C4676 vdd.n2357 gnd 0.007174f
C4677 vdd.n2358 gnd 0.231816f
C4678 vdd.n2359 gnd 0.007174f
C4679 vdd.n2360 gnd 0.007174f
C4680 vdd.n2361 gnd 0.007174f
C4681 vdd.n2362 gnd 0.007174f
C4682 vdd.n2363 gnd 0.007174f
C4683 vdd.n2364 gnd 0.007174f
C4684 vdd.n2365 gnd 0.007174f
C4685 vdd.n2366 gnd 0.007174f
C4686 vdd.n2367 gnd 0.007174f
C4687 vdd.n2368 gnd 0.007174f
C4688 vdd.n2369 gnd 0.007174f
C4689 vdd.n2370 gnd 0.007174f
C4690 vdd.n2371 gnd 0.007174f
C4691 vdd.n2372 gnd 0.007174f
C4692 vdd.n2373 gnd 0.007174f
C4693 vdd.n2374 gnd 0.007174f
C4694 vdd.n2375 gnd 0.007174f
C4695 vdd.n2376 gnd 0.007174f
C4696 vdd.n2377 gnd 0.007174f
C4697 vdd.n2378 gnd 0.007174f
C4698 vdd.n2379 gnd 0.007174f
C4699 vdd.n2380 gnd 0.007174f
C4700 vdd.n2381 gnd 0.007174f
C4701 vdd.n2382 gnd 0.007174f
C4702 vdd.n2383 gnd 0.007174f
C4703 vdd.n2384 gnd 0.007174f
C4704 vdd.n2385 gnd 0.007174f
C4705 vdd.n2386 gnd 0.007174f
C4706 vdd.n2387 gnd 0.007174f
C4707 vdd.n2388 gnd 0.007174f
C4708 vdd.n2389 gnd 0.007174f
C4709 vdd.n2390 gnd 0.007174f
C4710 vdd.n2391 gnd 0.007174f
C4711 vdd.n2392 gnd 0.007174f
C4712 vdd.n2393 gnd 0.007174f
C4713 vdd.n2394 gnd 0.015538f
C4714 vdd.n2395 gnd 0.016536f
C4715 vdd.n2396 gnd 0.016536f
C4716 vdd.n2398 gnd 0.007174f
C4717 vdd.n2400 gnd 0.007174f
C4718 vdd.n2401 gnd 0.005539f
C4719 vdd.n2402 gnd 0.010253f
C4720 vdd.n2403 gnd 0.005223f
C4721 vdd.n2404 gnd 0.007174f
C4722 vdd.n2405 gnd 0.007174f
C4723 vdd.n2407 gnd 0.007174f
C4724 vdd.n2409 gnd 0.007174f
C4725 vdd.n2410 gnd 0.007174f
C4726 vdd.n2411 gnd 0.007174f
C4727 vdd.n2412 gnd 0.007174f
C4728 vdd.n2413 gnd 0.007174f
C4729 vdd.n2415 gnd 0.007174f
C4730 vdd.n2417 gnd 0.007174f
C4731 vdd.n2418 gnd 0.007174f
C4732 vdd.n2419 gnd 0.007174f
C4733 vdd.n2420 gnd 0.007174f
C4734 vdd.n2421 gnd 0.007174f
C4735 vdd.n2423 gnd 0.007174f
C4736 vdd.n2425 gnd 0.007174f
C4737 vdd.n2426 gnd 0.007174f
C4738 vdd.n2427 gnd 0.007174f
C4739 vdd.n2428 gnd 0.007174f
C4740 vdd.n2429 gnd 0.007174f
C4741 vdd.n2431 gnd 0.007174f
C4742 vdd.n2433 gnd 0.007174f
C4743 vdd.n2434 gnd 0.007174f
C4744 vdd.n2435 gnd 0.007174f
C4745 vdd.n2436 gnd 0.007174f
C4746 vdd.n2437 gnd 0.007174f
C4747 vdd.n2439 gnd 0.007174f
C4748 vdd.n2441 gnd 0.007174f
C4749 vdd.n2442 gnd 0.007174f
C4750 vdd.n2443 gnd 0.007174f
C4751 vdd.n2444 gnd 0.007174f
C4752 vdd.n2445 gnd 0.007174f
C4753 vdd.n2447 gnd 0.007174f
C4754 vdd.n2449 gnd 0.007174f
C4755 vdd.n2450 gnd 0.007174f
C4756 vdd.n2451 gnd 0.007174f
C4757 vdd.n2452 gnd 0.007174f
C4758 vdd.n2453 gnd 0.007174f
C4759 vdd.n2455 gnd 0.007174f
C4760 vdd.n2456 gnd 0.007174f
C4761 vdd.n2457 gnd 0.007174f
C4762 vdd.n2458 gnd 0.007174f
C4763 vdd.n2459 gnd 0.007174f
C4764 vdd.n2460 gnd 0.007174f
C4765 vdd.n2462 gnd 0.007174f
C4766 vdd.n2463 gnd 0.007174f
C4767 vdd.n2464 gnd 0.016536f
C4768 vdd.n2465 gnd 0.015538f
C4769 vdd.n2466 gnd 0.015538f
C4770 vdd.n2467 gnd 1.01352f
C4771 vdd.n2468 gnd 0.015538f
C4772 vdd.n2469 gnd 0.015538f
C4773 vdd.n2470 gnd 0.007174f
C4774 vdd.n2471 gnd 0.007174f
C4775 vdd.n2472 gnd 0.007174f
C4776 vdd.n2473 gnd 0.501369f
C4777 vdd.n2474 gnd 0.007174f
C4778 vdd.n2475 gnd 0.007174f
C4779 vdd.n2476 gnd 0.007174f
C4780 vdd.n2477 gnd 0.007174f
C4781 vdd.n2478 gnd 0.007174f
C4782 vdd.n2479 gnd 0.733184f
C4783 vdd.n2480 gnd 0.007174f
C4784 vdd.n2481 gnd 0.007174f
C4785 vdd.n2482 gnd 0.007174f
C4786 vdd.n2483 gnd 0.007174f
C4787 vdd.n2484 gnd 0.007174f
C4788 vdd.n2485 gnd 0.733184f
C4789 vdd.n2486 gnd 0.007174f
C4790 vdd.n2487 gnd 0.007174f
C4791 vdd.n2488 gnd 0.007174f
C4792 vdd.n2489 gnd 0.007174f
C4793 vdd.n2490 gnd 0.007174f
C4794 vdd.n2491 gnd 0.371983f
C4795 vdd.n2492 gnd 0.007174f
C4796 vdd.n2493 gnd 0.007174f
C4797 vdd.n2494 gnd 0.007174f
C4798 vdd.n2495 gnd 0.007174f
C4799 vdd.n2496 gnd 0.007174f
C4800 vdd.n2497 gnd 0.533715f
C4801 vdd.n2498 gnd 0.007174f
C4802 vdd.n2499 gnd 0.007174f
C4803 vdd.n2500 gnd 0.007174f
C4804 vdd.n2501 gnd 0.007174f
C4805 vdd.n2502 gnd 0.007174f
C4806 vdd.n2503 gnd 0.695447f
C4807 vdd.n2504 gnd 0.007174f
C4808 vdd.n2505 gnd 0.007174f
C4809 vdd.n2506 gnd 0.007174f
C4810 vdd.n2507 gnd 0.007174f
C4811 vdd.n2508 gnd 0.007174f
C4812 vdd.n2509 gnd 0.733184f
C4813 vdd.n2510 gnd 0.007174f
C4814 vdd.n2511 gnd 0.007174f
C4815 vdd.n2512 gnd 0.007174f
C4816 vdd.n2513 gnd 0.007174f
C4817 vdd.n2514 gnd 0.007174f
C4818 vdd.n2515 gnd 0.60919f
C4819 vdd.n2516 gnd 0.007174f
C4820 vdd.n2517 gnd 0.007174f
C4821 vdd.n2518 gnd 0.005908f
C4822 vdd.n2519 gnd 0.020783f
C4823 vdd.n2520 gnd 0.004853f
C4824 vdd.n2521 gnd 0.007174f
C4825 vdd.n2522 gnd 0.447458f
C4826 vdd.n2523 gnd 0.007174f
C4827 vdd.n2524 gnd 0.007174f
C4828 vdd.n2525 gnd 0.007174f
C4829 vdd.n2526 gnd 0.007174f
C4830 vdd.n2527 gnd 0.007174f
C4831 vdd.n2528 gnd 0.447458f
C4832 vdd.n2529 gnd 0.007174f
C4833 vdd.n2530 gnd 0.007174f
C4834 vdd.n2531 gnd 0.007174f
C4835 vdd.n2532 gnd 0.007174f
C4836 vdd.n2533 gnd 0.007174f
C4837 vdd.n2534 gnd 0.60919f
C4838 vdd.n2535 gnd 0.007174f
C4839 vdd.n2536 gnd 0.007174f
C4840 vdd.n2537 gnd 0.007174f
C4841 vdd.n2538 gnd 0.007174f
C4842 vdd.n2539 gnd 0.007174f
C4843 vdd.n2540 gnd 0.625363f
C4844 vdd.n2541 gnd 0.007174f
C4845 vdd.n2542 gnd 0.007174f
C4846 vdd.n2543 gnd 0.007174f
C4847 vdd.n2544 gnd 0.007174f
C4848 vdd.n2545 gnd 0.007174f
C4849 vdd.n2546 gnd 0.463631f
C4850 vdd.n2547 gnd 0.007174f
C4851 vdd.n2548 gnd 0.007174f
C4852 vdd.n2549 gnd 0.007174f
C4853 vdd.n2550 gnd 0.007174f
C4854 vdd.n2551 gnd 0.007174f
C4855 vdd.n2552 gnd 0.231816f
C4856 vdd.n2553 gnd 0.007174f
C4857 vdd.n2554 gnd 0.007174f
C4858 vdd.n2555 gnd 0.007174f
C4859 vdd.n2556 gnd 0.007174f
C4860 vdd.n2557 gnd 0.007174f
C4861 vdd.n2558 gnd 0.231816f
C4862 vdd.n2559 gnd 0.007174f
C4863 vdd.n2560 gnd 0.007174f
C4864 vdd.n2561 gnd 0.007174f
C4865 vdd.n2562 gnd 0.007174f
C4866 vdd.n2563 gnd 0.007174f
C4867 vdd.n2564 gnd 0.733184f
C4868 vdd.n2565 gnd 0.007174f
C4869 vdd.n2566 gnd 0.007174f
C4870 vdd.n2567 gnd 0.007174f
C4871 vdd.n2568 gnd 0.007174f
C4872 vdd.n2569 gnd 0.007174f
C4873 vdd.n2570 gnd 0.007174f
C4874 vdd.n2571 gnd 0.007174f
C4875 vdd.n2572 gnd 0.528324f
C4876 vdd.n2573 gnd 0.007174f
C4877 vdd.n2574 gnd 0.007174f
C4878 vdd.n2575 gnd 0.007174f
C4879 vdd.n2576 gnd 0.007174f
C4880 vdd.n2577 gnd 0.007174f
C4881 vdd.n2578 gnd 0.007174f
C4882 vdd.n2579 gnd 0.45824f
C4883 vdd.n2580 gnd 0.007174f
C4884 vdd.n2581 gnd 0.007174f
C4885 vdd.n2582 gnd 0.007174f
C4886 vdd.n2583 gnd 0.016447f
C4887 vdd.n2584 gnd 0.015626f
C4888 vdd.n2585 gnd 0.007174f
C4889 vdd.n2586 gnd 0.007174f
C4890 vdd.n2587 gnd 0.005539f
C4891 vdd.n2588 gnd 0.007174f
C4892 vdd.n2589 gnd 0.007174f
C4893 vdd.n2590 gnd 0.005223f
C4894 vdd.n2591 gnd 0.007174f
C4895 vdd.n2592 gnd 0.007174f
C4896 vdd.n2593 gnd 0.007174f
C4897 vdd.n2594 gnd 0.007174f
C4898 vdd.n2595 gnd 0.007174f
C4899 vdd.n2596 gnd 0.007174f
C4900 vdd.n2597 gnd 0.007174f
C4901 vdd.n2598 gnd 0.007174f
C4902 vdd.n2599 gnd 0.007174f
C4903 vdd.n2600 gnd 0.007174f
C4904 vdd.n2601 gnd 0.007174f
C4905 vdd.n2602 gnd 0.007174f
C4906 vdd.n2603 gnd 0.007174f
C4907 vdd.n2604 gnd 0.007174f
C4908 vdd.n2605 gnd 0.007174f
C4909 vdd.n2606 gnd 0.007174f
C4910 vdd.n2607 gnd 0.007174f
C4911 vdd.n2608 gnd 0.007174f
C4912 vdd.n2609 gnd 0.007174f
C4913 vdd.n2610 gnd 0.007174f
C4914 vdd.n2611 gnd 0.007174f
C4915 vdd.n2612 gnd 0.007174f
C4916 vdd.n2613 gnd 0.007174f
C4917 vdd.n2614 gnd 0.007174f
C4918 vdd.n2615 gnd 0.007174f
C4919 vdd.n2616 gnd 0.007174f
C4920 vdd.n2617 gnd 0.007174f
C4921 vdd.n2618 gnd 0.007174f
C4922 vdd.n2619 gnd 0.007174f
C4923 vdd.n2620 gnd 0.007174f
C4924 vdd.n2621 gnd 0.007174f
C4925 vdd.n2622 gnd 0.007174f
C4926 vdd.n2623 gnd 0.007174f
C4927 vdd.n2624 gnd 0.007174f
C4928 vdd.n2625 gnd 0.007174f
C4929 vdd.n2626 gnd 0.007174f
C4930 vdd.n2627 gnd 0.007174f
C4931 vdd.n2628 gnd 0.007174f
C4932 vdd.n2629 gnd 0.007174f
C4933 vdd.n2630 gnd 0.007174f
C4934 vdd.n2631 gnd 0.007174f
C4935 vdd.n2632 gnd 0.007174f
C4936 vdd.n2633 gnd 0.007174f
C4937 vdd.n2634 gnd 0.007174f
C4938 vdd.n2635 gnd 0.007174f
C4939 vdd.n2636 gnd 0.007174f
C4940 vdd.n2637 gnd 0.007174f
C4941 vdd.n2638 gnd 0.007174f
C4942 vdd.n2639 gnd 0.007174f
C4943 vdd.n2640 gnd 0.007174f
C4944 vdd.n2641 gnd 0.007174f
C4945 vdd.n2642 gnd 0.007174f
C4946 vdd.n2643 gnd 0.007174f
C4947 vdd.n2644 gnd 0.007174f
C4948 vdd.n2645 gnd 0.007174f
C4949 vdd.n2646 gnd 0.007174f
C4950 vdd.n2647 gnd 0.007174f
C4951 vdd.n2648 gnd 0.007174f
C4952 vdd.n2649 gnd 0.007174f
C4953 vdd.n2650 gnd 0.007174f
C4954 vdd.n2651 gnd 0.016536f
C4955 vdd.n2652 gnd 0.015538f
C4956 vdd.n2653 gnd 0.015538f
C4957 vdd.n2654 gnd 0.851787f
C4958 vdd.n2655 gnd 0.015538f
C4959 vdd.n2656 gnd 0.016536f
C4960 vdd.n2657 gnd 0.015626f
C4961 vdd.n2658 gnd 0.007174f
C4962 vdd.n2659 gnd 0.007174f
C4963 vdd.n2660 gnd 0.007174f
C4964 vdd.n2661 gnd 0.005539f
C4965 vdd.n2662 gnd 0.010253f
C4966 vdd.n2663 gnd 0.005223f
C4967 vdd.n2664 gnd 0.007174f
C4968 vdd.n2665 gnd 0.007174f
C4969 vdd.n2666 gnd 0.007174f
C4970 vdd.n2667 gnd 0.007174f
C4971 vdd.n2668 gnd 0.007174f
C4972 vdd.n2669 gnd 0.007174f
C4973 vdd.n2670 gnd 0.007174f
C4974 vdd.n2671 gnd 0.007174f
C4975 vdd.n2672 gnd 0.007174f
C4976 vdd.n2673 gnd 0.007174f
C4977 vdd.n2674 gnd 0.007174f
C4978 vdd.n2675 gnd 0.007174f
C4979 vdd.n2676 gnd 0.007174f
C4980 vdd.n2677 gnd 0.007174f
C4981 vdd.n2678 gnd 0.007174f
C4982 vdd.n2679 gnd 0.007174f
C4983 vdd.n2680 gnd 0.007174f
C4984 vdd.n2681 gnd 0.007174f
C4985 vdd.n2682 gnd 0.007174f
C4986 vdd.n2683 gnd 0.007174f
C4987 vdd.n2684 gnd 0.007174f
C4988 vdd.n2685 gnd 0.007174f
C4989 vdd.n2686 gnd 0.007174f
C4990 vdd.n2687 gnd 0.007174f
C4991 vdd.n2688 gnd 0.007174f
C4992 vdd.n2689 gnd 0.007174f
C4993 vdd.n2690 gnd 0.007174f
C4994 vdd.n2691 gnd 0.007174f
C4995 vdd.n2692 gnd 0.007174f
C4996 vdd.n2693 gnd 0.007174f
C4997 vdd.n2694 gnd 0.007174f
C4998 vdd.n2695 gnd 0.007174f
C4999 vdd.n2696 gnd 0.007174f
C5000 vdd.n2697 gnd 0.007174f
C5001 vdd.n2698 gnd 0.007174f
C5002 vdd.n2699 gnd 0.007174f
C5003 vdd.n2700 gnd 0.007174f
C5004 vdd.n2701 gnd 0.007174f
C5005 vdd.n2702 gnd 0.007174f
C5006 vdd.n2703 gnd 0.007174f
C5007 vdd.n2704 gnd 0.007174f
C5008 vdd.n2705 gnd 0.007174f
C5009 vdd.n2706 gnd 0.007174f
C5010 vdd.n2707 gnd 0.007174f
C5011 vdd.n2708 gnd 0.007174f
C5012 vdd.n2709 gnd 0.007174f
C5013 vdd.n2710 gnd 0.007174f
C5014 vdd.n2711 gnd 0.007174f
C5015 vdd.n2712 gnd 0.007174f
C5016 vdd.n2713 gnd 0.007174f
C5017 vdd.n2714 gnd 0.007174f
C5018 vdd.n2715 gnd 0.007174f
C5019 vdd.n2716 gnd 0.007174f
C5020 vdd.n2717 gnd 0.007174f
C5021 vdd.n2718 gnd 0.007174f
C5022 vdd.n2719 gnd 0.007174f
C5023 vdd.n2720 gnd 0.007174f
C5024 vdd.n2721 gnd 0.007174f
C5025 vdd.n2722 gnd 0.007174f
C5026 vdd.n2723 gnd 0.007174f
C5027 vdd.n2724 gnd 0.016536f
C5028 vdd.n2725 gnd 0.016536f
C5029 vdd.n2726 gnd 0.894916f
C5030 vdd.t10 gnd 3.18073f
C5031 vdd.t0 gnd 3.18073f
C5032 vdd.n2760 gnd 0.007174f
C5033 vdd.t128 gnd 0.289914f
C5034 vdd.t129 gnd 0.296763f
C5035 vdd.t127 gnd 0.189267f
C5036 vdd.n2761 gnd 0.102288f
C5037 vdd.n2762 gnd 0.058021f
C5038 vdd.n2763 gnd 0.010253f
C5039 vdd.n2764 gnd 0.007174f
C5040 vdd.n2765 gnd 0.007174f
C5041 vdd.n2766 gnd 0.007174f
C5042 vdd.n2767 gnd 0.007174f
C5043 vdd.n2768 gnd 0.007174f
C5044 vdd.n2769 gnd 0.007174f
C5045 vdd.n2770 gnd 0.007174f
C5046 vdd.n2771 gnd 0.007174f
C5047 vdd.n2772 gnd 0.007174f
C5048 vdd.n2773 gnd 0.007174f
C5049 vdd.n2774 gnd 0.007174f
C5050 vdd.n2775 gnd 0.007174f
C5051 vdd.n2776 gnd 0.007174f
C5052 vdd.n2777 gnd 0.007174f
C5053 vdd.n2778 gnd 0.007174f
C5054 vdd.n2779 gnd 0.007174f
C5055 vdd.n2780 gnd 0.007174f
C5056 vdd.n2781 gnd 0.007174f
C5057 vdd.n2782 gnd 0.007174f
C5058 vdd.n2783 gnd 0.007174f
C5059 vdd.n2784 gnd 0.007174f
C5060 vdd.n2785 gnd 0.007174f
C5061 vdd.n2786 gnd 0.007174f
C5062 vdd.n2787 gnd 0.007174f
C5063 vdd.n2788 gnd 0.007174f
C5064 vdd.n2789 gnd 0.007174f
C5065 vdd.n2790 gnd 0.007174f
C5066 vdd.n2791 gnd 0.007174f
C5067 vdd.n2792 gnd 0.007174f
C5068 vdd.n2793 gnd 0.007174f
C5069 vdd.n2794 gnd 0.007174f
C5070 vdd.n2795 gnd 0.007174f
C5071 vdd.n2796 gnd 0.007174f
C5072 vdd.n2797 gnd 0.007174f
C5073 vdd.n2798 gnd 0.007174f
C5074 vdd.n2799 gnd 0.007174f
C5075 vdd.n2800 gnd 0.007174f
C5076 vdd.n2801 gnd 0.007174f
C5077 vdd.n2802 gnd 0.007174f
C5078 vdd.n2803 gnd 0.007174f
C5079 vdd.n2804 gnd 0.007174f
C5080 vdd.n2805 gnd 0.007174f
C5081 vdd.n2806 gnd 0.007174f
C5082 vdd.n2807 gnd 0.007174f
C5083 vdd.n2808 gnd 0.007174f
C5084 vdd.n2809 gnd 0.007174f
C5085 vdd.n2810 gnd 0.007174f
C5086 vdd.n2811 gnd 0.007174f
C5087 vdd.n2812 gnd 0.007174f
C5088 vdd.n2813 gnd 0.007174f
C5089 vdd.n2814 gnd 0.007174f
C5090 vdd.n2815 gnd 0.007174f
C5091 vdd.n2816 gnd 0.007174f
C5092 vdd.n2817 gnd 0.007174f
C5093 vdd.n2818 gnd 0.007174f
C5094 vdd.n2819 gnd 0.007174f
C5095 vdd.n2820 gnd 0.007174f
C5096 vdd.n2821 gnd 0.007174f
C5097 vdd.n2822 gnd 0.007174f
C5098 vdd.n2823 gnd 0.007174f
C5099 vdd.n2824 gnd 0.005223f
C5100 vdd.n2825 gnd 0.007174f
C5101 vdd.n2826 gnd 0.007174f
C5102 vdd.n2827 gnd 0.005539f
C5103 vdd.n2828 gnd 0.007174f
C5104 vdd.n2829 gnd 0.007174f
C5105 vdd.t115 gnd 0.289914f
C5106 vdd.t116 gnd 0.296763f
C5107 vdd.t113 gnd 0.189267f
C5108 vdd.n2830 gnd 0.102288f
C5109 vdd.n2831 gnd 0.058021f
C5110 vdd.n2832 gnd 0.007174f
C5111 vdd.n2833 gnd 0.007174f
C5112 vdd.n2834 gnd 0.007174f
C5113 vdd.n2835 gnd 0.007174f
C5114 vdd.n2836 gnd 0.007174f
C5115 vdd.n2837 gnd 0.007174f
C5116 vdd.n2838 gnd 0.007174f
C5117 vdd.n2839 gnd 0.007174f
C5118 vdd.n2840 gnd 0.007174f
C5119 vdd.n2841 gnd 0.007174f
C5120 vdd.n2842 gnd 0.007174f
C5121 vdd.n2843 gnd 0.007174f
C5122 vdd.n2844 gnd 0.007174f
C5123 vdd.n2845 gnd 0.007174f
C5124 vdd.n2846 gnd 0.007174f
C5125 vdd.n2847 gnd 0.007174f
C5126 vdd.n2848 gnd 0.007174f
C5127 vdd.n2849 gnd 0.007174f
C5128 vdd.n2850 gnd 0.007174f
C5129 vdd.n2851 gnd 0.007174f
C5130 vdd.n2852 gnd 0.007174f
C5131 vdd.n2853 gnd 0.007174f
C5132 vdd.n2854 gnd 0.007174f
C5133 vdd.n2855 gnd 0.007174f
C5134 vdd.n2856 gnd 0.007174f
C5135 vdd.n2857 gnd 0.007174f
C5136 vdd.n2858 gnd 0.007174f
C5137 vdd.n2859 gnd 0.007174f
C5138 vdd.n2860 gnd 0.007174f
C5139 vdd.n2861 gnd 0.007174f
C5140 vdd.n2862 gnd 0.007174f
C5141 vdd.n2863 gnd 0.007174f
C5142 vdd.n2864 gnd 0.007174f
C5143 vdd.n2865 gnd 0.007174f
C5144 vdd.n2866 gnd 0.007174f
C5145 vdd.n2867 gnd 0.007174f
C5146 vdd.n2868 gnd 0.007174f
C5147 vdd.n2869 gnd 0.007174f
C5148 vdd.n2870 gnd 0.007174f
C5149 vdd.n2871 gnd 0.007174f
C5150 vdd.n2872 gnd 0.007174f
C5151 vdd.n2873 gnd 0.007174f
C5152 vdd.n2874 gnd 0.007174f
C5153 vdd.n2875 gnd 0.007174f
C5154 vdd.n2876 gnd 0.007174f
C5155 vdd.n2877 gnd 0.007174f
C5156 vdd.n2878 gnd 0.007174f
C5157 vdd.n2879 gnd 0.007174f
C5158 vdd.n2880 gnd 0.007174f
C5159 vdd.n2881 gnd 0.007174f
C5160 vdd.n2882 gnd 0.007174f
C5161 vdd.n2883 gnd 0.007174f
C5162 vdd.n2884 gnd 0.007174f
C5163 vdd.n2885 gnd 0.007174f
C5164 vdd.n2886 gnd 0.007174f
C5165 vdd.n2887 gnd 0.007174f
C5166 vdd.n2888 gnd 0.007174f
C5167 vdd.n2889 gnd 0.005223f
C5168 vdd.n2890 gnd 0.010253f
C5169 vdd.n2891 gnd 0.005539f
C5170 vdd.n2892 gnd 0.007174f
C5171 vdd.n2893 gnd 0.007174f
C5172 vdd.n2894 gnd 0.007174f
C5173 vdd.n2895 gnd 0.016536f
C5174 vdd.n2896 gnd 0.016536f
C5175 vdd.n2897 gnd 0.015538f
C5176 vdd.n2898 gnd 0.007174f
C5177 vdd.n2899 gnd 0.007174f
C5178 vdd.n2900 gnd 0.007174f
C5179 vdd.n2901 gnd 0.007174f
C5180 vdd.n2902 gnd 0.007174f
C5181 vdd.n2903 gnd 0.007174f
C5182 vdd.n2904 gnd 0.007174f
C5183 vdd.n2905 gnd 0.007174f
C5184 vdd.n2906 gnd 0.007174f
C5185 vdd.n2907 gnd 0.007174f
C5186 vdd.n2908 gnd 0.007174f
C5187 vdd.n2909 gnd 0.007174f
C5188 vdd.n2910 gnd 0.007174f
C5189 vdd.n2911 gnd 0.007174f
C5190 vdd.n2912 gnd 0.007174f
C5191 vdd.n2913 gnd 0.007174f
C5192 vdd.n2914 gnd 0.007174f
C5193 vdd.n2915 gnd 0.007174f
C5194 vdd.n2916 gnd 0.007174f
C5195 vdd.n2917 gnd 0.007174f
C5196 vdd.n2918 gnd 0.007174f
C5197 vdd.n2919 gnd 0.007174f
C5198 vdd.n2920 gnd 0.007174f
C5199 vdd.n2921 gnd 0.007174f
C5200 vdd.n2922 gnd 0.007174f
C5201 vdd.n2923 gnd 0.007174f
C5202 vdd.n2924 gnd 0.007174f
C5203 vdd.n2925 gnd 0.007174f
C5204 vdd.n2926 gnd 0.007174f
C5205 vdd.n2927 gnd 0.007174f
C5206 vdd.n2928 gnd 0.007174f
C5207 vdd.n2929 gnd 0.007174f
C5208 vdd.n2930 gnd 0.007174f
C5209 vdd.n2931 gnd 0.007174f
C5210 vdd.n2932 gnd 0.007174f
C5211 vdd.n2933 gnd 0.007174f
C5212 vdd.n2934 gnd 0.007174f
C5213 vdd.n2935 gnd 0.007174f
C5214 vdd.n2936 gnd 0.007174f
C5215 vdd.n2937 gnd 0.007174f
C5216 vdd.n2938 gnd 0.007174f
C5217 vdd.n2939 gnd 0.007174f
C5218 vdd.n2940 gnd 0.007174f
C5219 vdd.n2941 gnd 0.007174f
C5220 vdd.n2942 gnd 0.007174f
C5221 vdd.n2943 gnd 0.007174f
C5222 vdd.n2944 gnd 0.007174f
C5223 vdd.n2945 gnd 0.007174f
C5224 vdd.n2946 gnd 0.007174f
C5225 vdd.n2947 gnd 0.007174f
C5226 vdd.n2948 gnd 0.007174f
C5227 vdd.n2949 gnd 0.007174f
C5228 vdd.n2950 gnd 0.007174f
C5229 vdd.n2951 gnd 0.007174f
C5230 vdd.n2952 gnd 0.007174f
C5231 vdd.n2953 gnd 0.007174f
C5232 vdd.n2954 gnd 0.007174f
C5233 vdd.n2955 gnd 0.007174f
C5234 vdd.n2956 gnd 0.007174f
C5235 vdd.n2957 gnd 0.007174f
C5236 vdd.n2958 gnd 0.007174f
C5237 vdd.n2959 gnd 0.007174f
C5238 vdd.n2960 gnd 0.007174f
C5239 vdd.n2961 gnd 0.007174f
C5240 vdd.n2962 gnd 0.007174f
C5241 vdd.n2963 gnd 0.007174f
C5242 vdd.n2964 gnd 0.007174f
C5243 vdd.n2965 gnd 0.007174f
C5244 vdd.n2966 gnd 0.007174f
C5245 vdd.n2967 gnd 0.007174f
C5246 vdd.n2968 gnd 0.007174f
C5247 vdd.n2969 gnd 0.007174f
C5248 vdd.n2970 gnd 0.007174f
C5249 vdd.n2971 gnd 0.007174f
C5250 vdd.n2972 gnd 0.007174f
C5251 vdd.n2973 gnd 0.007174f
C5252 vdd.n2974 gnd 0.007174f
C5253 vdd.n2975 gnd 0.007174f
C5254 vdd.n2976 gnd 0.007174f
C5255 vdd.n2977 gnd 0.231816f
C5256 vdd.n2978 gnd 0.007174f
C5257 vdd.n2979 gnd 0.007174f
C5258 vdd.n2980 gnd 0.007174f
C5259 vdd.n2981 gnd 0.007174f
C5260 vdd.n2982 gnd 0.007174f
C5261 vdd.n2983 gnd 0.007174f
C5262 vdd.n2984 gnd 0.007174f
C5263 vdd.n2985 gnd 0.007174f
C5264 vdd.n2986 gnd 0.007174f
C5265 vdd.n2987 gnd 0.007174f
C5266 vdd.n2988 gnd 0.007174f
C5267 vdd.n2989 gnd 0.6631f
C5268 vdd.n2990 gnd 0.007174f
C5269 vdd.n2991 gnd 0.007174f
C5270 vdd.n2992 gnd 0.007174f
C5271 vdd.n2993 gnd 0.007174f
C5272 vdd.n2994 gnd 0.007174f
C5273 vdd.n2995 gnd 0.007174f
C5274 vdd.n2996 gnd 0.007174f
C5275 vdd.n2997 gnd 0.007174f
C5276 vdd.n2998 gnd 0.007174f
C5277 vdd.n2999 gnd 0.007174f
C5278 vdd.n3000 gnd 0.007174f
C5279 vdd.n3001 gnd 0.436676f
C5280 vdd.n3002 gnd 0.007174f
C5281 vdd.n3003 gnd 0.007174f
C5282 vdd.n3004 gnd 0.007174f
C5283 vdd.n3005 gnd 0.007174f
C5284 vdd.n3006 gnd 0.007174f
C5285 vdd.n3007 gnd 0.015538f
C5286 vdd.n3008 gnd 0.016536f
C5287 vdd.n3009 gnd 0.016536f
C5288 vdd.n3010 gnd 0.894916f
C5289 vdd.n3012 gnd 0.007174f
C5290 vdd.n3013 gnd 0.007174f
C5291 vdd.n3014 gnd 0.016536f
C5292 vdd.n3015 gnd 0.015538f
C5293 vdd.n3016 gnd 0.015538f
C5294 vdd.n3017 gnd 0.851787f
C5295 vdd.n3018 gnd 0.015538f
C5296 vdd.n3019 gnd 0.015538f
C5297 vdd.n3020 gnd 0.007174f
C5298 vdd.n3021 gnd 0.007174f
C5299 vdd.n3022 gnd 0.007174f
C5300 vdd.n3023 gnd 0.45824f
C5301 vdd.n3024 gnd 0.007174f
C5302 vdd.n3025 gnd 0.007174f
C5303 vdd.n3026 gnd 0.007174f
C5304 vdd.n3027 gnd 0.007174f
C5305 vdd.n3028 gnd 0.007174f
C5306 vdd.n3029 gnd 0.528324f
C5307 vdd.n3030 gnd 0.007174f
C5308 vdd.n3031 gnd 0.007174f
C5309 vdd.n3032 gnd 0.007174f
C5310 vdd.n3033 gnd 0.007174f
C5311 vdd.n3034 gnd 0.007174f
C5312 vdd.n3035 gnd 0.733184f
C5313 vdd.n3036 gnd 0.007174f
C5314 vdd.n3037 gnd 0.007174f
C5315 vdd.n3038 gnd 0.007174f
C5316 vdd.n3039 gnd 0.007174f
C5317 vdd.n3040 gnd 0.007174f
C5318 vdd.n3041 gnd 0.231816f
C5319 vdd.n3042 gnd 0.007174f
C5320 vdd.n3043 gnd 0.007174f
C5321 vdd.n3044 gnd 0.007174f
C5322 vdd.n3045 gnd 0.007174f
C5323 vdd.n3046 gnd 0.007174f
C5324 vdd.n3047 gnd 0.231816f
C5325 vdd.n3048 gnd 0.007174f
C5326 vdd.n3049 gnd 0.007174f
C5327 vdd.n3050 gnd 0.007174f
C5328 vdd.n3051 gnd 0.007174f
C5329 vdd.n3052 gnd 0.007174f
C5330 vdd.n3053 gnd 0.463631f
C5331 vdd.n3054 gnd 0.007174f
C5332 vdd.n3055 gnd 0.007174f
C5333 vdd.n3056 gnd 0.007174f
C5334 vdd.n3057 gnd 0.007174f
C5335 vdd.n3058 gnd 0.007174f
C5336 vdd.n3059 gnd 0.625363f
C5337 vdd.n3060 gnd 0.007174f
C5338 vdd.n3061 gnd 0.007174f
C5339 vdd.n3062 gnd 0.007174f
C5340 vdd.n3063 gnd 0.007174f
C5341 vdd.n3064 gnd 0.007174f
C5342 vdd.n3065 gnd 0.60919f
C5343 vdd.n3066 gnd 0.007174f
C5344 vdd.n3067 gnd 0.007174f
C5345 vdd.n3068 gnd 0.007174f
C5346 vdd.n3069 gnd 0.007174f
C5347 vdd.n3070 gnd 0.007174f
C5348 vdd.n3071 gnd 0.447458f
C5349 vdd.n3072 gnd 0.007174f
C5350 vdd.n3073 gnd 0.007174f
C5351 vdd.n3074 gnd 0.007174f
C5352 vdd.n3075 gnd 0.007174f
C5353 vdd.n3076 gnd 0.007174f
C5354 vdd.n3077 gnd 0.447458f
C5355 vdd.n3078 gnd 0.007174f
C5356 vdd.n3079 gnd 0.004853f
C5357 vdd.n3080 gnd 0.020783f
C5358 vdd.n3081 gnd 0.005908f
C5359 vdd.n3082 gnd 0.007174f
C5360 vdd.n3083 gnd 0.007174f
C5361 vdd.n3084 gnd 0.60919f
C5362 vdd.n3085 gnd 0.007174f
C5363 vdd.n3086 gnd 0.007174f
C5364 vdd.n3087 gnd 0.007174f
C5365 vdd.n3088 gnd 0.007174f
C5366 vdd.n3089 gnd 0.007174f
C5367 vdd.n3090 gnd 0.733184f
C5368 vdd.n3091 gnd 0.007174f
C5369 vdd.n3092 gnd 0.007174f
C5370 vdd.n3093 gnd 0.007174f
C5371 vdd.n3094 gnd 0.007174f
C5372 vdd.n3095 gnd 0.007174f
C5373 vdd.n3096 gnd 0.695447f
C5374 vdd.n3097 gnd 0.007174f
C5375 vdd.n3098 gnd 0.007174f
C5376 vdd.n3099 gnd 0.007174f
C5377 vdd.n3100 gnd 0.007174f
C5378 vdd.n3101 gnd 0.007174f
C5379 vdd.n3102 gnd 0.533715f
C5380 vdd.n3103 gnd 0.007174f
C5381 vdd.n3104 gnd 0.007174f
C5382 vdd.n3105 gnd 0.007174f
C5383 vdd.n3106 gnd 0.007174f
C5384 vdd.n3107 gnd 0.007174f
C5385 vdd.n3108 gnd 0.371983f
C5386 vdd.n3109 gnd 0.007174f
C5387 vdd.n3110 gnd 0.007174f
C5388 vdd.n3111 gnd 0.007174f
C5389 vdd.n3112 gnd 0.007174f
C5390 vdd.n3113 gnd 0.007174f
C5391 vdd.n3114 gnd 0.733184f
C5392 vdd.n3115 gnd 0.007174f
C5393 vdd.n3116 gnd 0.007174f
C5394 vdd.n3117 gnd 0.007174f
C5395 vdd.n3118 gnd 0.007174f
C5396 vdd.n3119 gnd 0.007174f
C5397 vdd.n3120 gnd 0.007174f
C5398 vdd.n3122 gnd 0.007174f
C5399 vdd.n3123 gnd 0.007174f
C5400 vdd.n3125 gnd 0.007174f
C5401 vdd.n3126 gnd 0.007174f
C5402 vdd.n3129 gnd 0.007174f
C5403 vdd.n3130 gnd 0.007174f
C5404 vdd.n3131 gnd 0.007174f
C5405 vdd.n3132 gnd 0.007174f
C5406 vdd.n3134 gnd 0.007174f
C5407 vdd.n3135 gnd 0.007174f
C5408 vdd.n3136 gnd 0.007174f
C5409 vdd.n3137 gnd 0.007174f
C5410 vdd.n3138 gnd 0.007174f
C5411 vdd.n3139 gnd 0.007174f
C5412 vdd.n3141 gnd 0.007174f
C5413 vdd.n3142 gnd 0.007174f
C5414 vdd.n3143 gnd 0.007174f
C5415 vdd.n3144 gnd 0.007174f
C5416 vdd.n3145 gnd 0.007174f
C5417 vdd.n3146 gnd 0.007174f
C5418 vdd.n3148 gnd 0.007174f
C5419 vdd.n3149 gnd 0.007174f
C5420 vdd.n3150 gnd 0.007174f
C5421 vdd.n3151 gnd 0.007174f
C5422 vdd.n3152 gnd 0.007174f
C5423 vdd.n3153 gnd 0.007174f
C5424 vdd.n3155 gnd 0.007174f
C5425 vdd.n3156 gnd 0.016536f
C5426 vdd.n3157 gnd 0.016536f
C5427 vdd.n3158 gnd 0.015538f
C5428 vdd.n3159 gnd 0.007174f
C5429 vdd.n3160 gnd 0.007174f
C5430 vdd.n3161 gnd 0.007174f
C5431 vdd.n3162 gnd 0.007174f
C5432 vdd.n3163 gnd 0.007174f
C5433 vdd.n3164 gnd 0.007174f
C5434 vdd.n3165 gnd 0.733184f
C5435 vdd.n3166 gnd 0.007174f
C5436 vdd.n3167 gnd 0.007174f
C5437 vdd.n3168 gnd 0.007174f
C5438 vdd.n3169 gnd 0.007174f
C5439 vdd.n3170 gnd 0.007174f
C5440 vdd.n3171 gnd 0.501369f
C5441 vdd.n3172 gnd 0.007174f
C5442 vdd.n3173 gnd 0.007174f
C5443 vdd.n3174 gnd 0.007174f
C5444 vdd.n3175 gnd 0.016447f
C5445 vdd.n3176 gnd 0.015626f
C5446 vdd.n3177 gnd 0.016536f
C5447 vdd.n3179 gnd 0.007174f
C5448 vdd.n3180 gnd 0.007174f
C5449 vdd.n3181 gnd 0.005539f
C5450 vdd.n3182 gnd 0.010253f
C5451 vdd.n3183 gnd 0.005223f
C5452 vdd.n3184 gnd 0.007174f
C5453 vdd.n3185 gnd 0.007174f
C5454 vdd.n3187 gnd 0.007174f
C5455 vdd.n3188 gnd 0.007174f
C5456 vdd.n3189 gnd 0.007174f
C5457 vdd.n3190 gnd 0.007174f
C5458 vdd.n3191 gnd 0.007174f
C5459 vdd.n3192 gnd 0.007174f
C5460 vdd.n3194 gnd 0.007174f
C5461 vdd.n3195 gnd 0.007174f
C5462 vdd.n3196 gnd 0.007174f
C5463 vdd.n3197 gnd 0.007174f
C5464 vdd.n3198 gnd 0.007174f
C5465 vdd.n3199 gnd 0.007174f
C5466 vdd.n3201 gnd 0.007174f
C5467 vdd.n3202 gnd 0.007174f
C5468 vdd.n3203 gnd 0.007174f
C5469 vdd.n3204 gnd 0.007174f
C5470 vdd.n3205 gnd 0.007174f
C5471 vdd.n3206 gnd 0.007174f
C5472 vdd.n3208 gnd 0.007174f
C5473 vdd.n3209 gnd 0.007174f
C5474 vdd.n3210 gnd 0.007174f
C5475 vdd.n3212 gnd 0.007174f
C5476 vdd.n3213 gnd 0.007174f
C5477 vdd.n3214 gnd 0.007174f
C5478 vdd.n3215 gnd 0.007174f
C5479 vdd.n3216 gnd 0.007174f
C5480 vdd.n3217 gnd 0.007174f
C5481 vdd.n3219 gnd 0.007174f
C5482 vdd.n3220 gnd 0.007174f
C5483 vdd.n3221 gnd 0.007174f
C5484 vdd.n3222 gnd 0.007174f
C5485 vdd.n3223 gnd 0.007174f
C5486 vdd.n3224 gnd 0.007174f
C5487 vdd.n3226 gnd 0.007174f
C5488 vdd.n3227 gnd 0.007174f
C5489 vdd.n3228 gnd 0.007174f
C5490 vdd.n3229 gnd 0.007174f
C5491 vdd.n3230 gnd 0.007174f
C5492 vdd.n3231 gnd 0.007174f
C5493 vdd.n3233 gnd 0.007174f
C5494 vdd.n3234 gnd 0.007174f
C5495 vdd.n3236 gnd 0.007174f
C5496 vdd.n3237 gnd 0.007174f
C5497 vdd.n3238 gnd 0.016536f
C5498 vdd.n3239 gnd 0.015538f
C5499 vdd.n3240 gnd 0.015538f
C5500 vdd.n3241 gnd 1.01352f
C5501 vdd.n3242 gnd 0.015538f
C5502 vdd.n3243 gnd 0.016536f
C5503 vdd.n3244 gnd 0.015626f
C5504 vdd.n3245 gnd 0.007174f
C5505 vdd.n3246 gnd 0.005539f
C5506 vdd.n3247 gnd 0.007174f
C5507 vdd.n3249 gnd 0.007174f
C5508 vdd.n3250 gnd 0.007174f
C5509 vdd.n3251 gnd 0.007174f
C5510 vdd.n3252 gnd 0.007174f
C5511 vdd.n3253 gnd 0.007174f
C5512 vdd.n3254 gnd 0.007174f
C5513 vdd.n3256 gnd 0.007174f
C5514 vdd.n3257 gnd 0.007174f
C5515 vdd.n3258 gnd 0.007174f
C5516 vdd.n3259 gnd 0.007174f
C5517 vdd.n3260 gnd 0.007174f
C5518 vdd.n3261 gnd 0.007174f
C5519 vdd.n3263 gnd 0.007174f
C5520 vdd.n3264 gnd 0.007174f
C5521 vdd.n3265 gnd 0.007174f
C5522 vdd.n3266 gnd 0.007174f
C5523 vdd.n3267 gnd 0.007174f
C5524 vdd.n3268 gnd 0.007174f
C5525 vdd.n3270 gnd 0.007174f
C5526 vdd.n3271 gnd 0.007174f
C5527 vdd.n3273 gnd 0.007174f
C5528 vdd.n3274 gnd 0.033676f
C5529 vdd.n3275 gnd 0.963832f
C5530 vdd.n3277 gnd 0.004458f
C5531 vdd.n3278 gnd 0.008492f
C5532 vdd.n3279 gnd 0.01055f
C5533 vdd.n3280 gnd 0.01055f
C5534 vdd.n3281 gnd 0.008492f
C5535 vdd.n3282 gnd 0.008492f
C5536 vdd.n3283 gnd 0.01055f
C5537 vdd.n3284 gnd 0.01055f
C5538 vdd.n3285 gnd 0.008492f
C5539 vdd.n3286 gnd 0.008492f
C5540 vdd.n3287 gnd 0.01055f
C5541 vdd.n3288 gnd 0.01055f
C5542 vdd.n3289 gnd 0.008492f
C5543 vdd.n3290 gnd 0.008492f
C5544 vdd.n3291 gnd 0.01055f
C5545 vdd.n3292 gnd 0.01055f
C5546 vdd.n3293 gnd 0.008492f
C5547 vdd.n3294 gnd 0.008492f
C5548 vdd.n3295 gnd 0.01055f
C5549 vdd.n3296 gnd 0.01055f
C5550 vdd.n3297 gnd 0.008492f
C5551 vdd.n3298 gnd 0.008492f
C5552 vdd.n3299 gnd 0.01055f
C5553 vdd.n3300 gnd 0.01055f
C5554 vdd.n3301 gnd 0.008492f
C5555 vdd.n3302 gnd 0.008492f
C5556 vdd.n3303 gnd 0.01055f
C5557 vdd.n3304 gnd 0.01055f
C5558 vdd.n3305 gnd 0.008492f
C5559 vdd.n3306 gnd 0.008492f
C5560 vdd.n3307 gnd 0.01055f
C5561 vdd.n3308 gnd 0.01055f
C5562 vdd.n3309 gnd 0.008492f
C5563 vdd.n3310 gnd 0.008492f
C5564 vdd.n3311 gnd 0.01055f
C5565 vdd.n3312 gnd 0.01055f
C5566 vdd.n3313 gnd 0.008492f
C5567 vdd.n3314 gnd 0.01055f
C5568 vdd.n3315 gnd 0.01055f
C5569 vdd.n3316 gnd 0.008492f
C5570 vdd.n3317 gnd 0.01055f
C5571 vdd.n3318 gnd 0.01055f
C5572 vdd.n3319 gnd 0.01055f
C5573 vdd.n3320 gnd 0.017323f
C5574 vdd.n3321 gnd 0.01055f
C5575 vdd.n3322 gnd 0.01055f
C5576 vdd.n3323 gnd 0.005774f
C5577 vdd.n3324 gnd 0.008492f
C5578 vdd.n3325 gnd 0.01055f
C5579 vdd.n3326 gnd 0.01055f
C5580 vdd.n3327 gnd 0.008492f
C5581 vdd.n3328 gnd 0.008492f
C5582 vdd.n3329 gnd 0.01055f
C5583 vdd.n3330 gnd 0.01055f
C5584 vdd.n3331 gnd 0.008492f
C5585 vdd.n3332 gnd 0.008492f
C5586 vdd.n3333 gnd 0.01055f
C5587 vdd.n3334 gnd 0.01055f
C5588 vdd.n3335 gnd 0.008492f
C5589 vdd.n3336 gnd 0.008492f
C5590 vdd.n3337 gnd 0.01055f
C5591 vdd.n3338 gnd 0.01055f
C5592 vdd.n3339 gnd 0.008492f
C5593 vdd.n3340 gnd 0.008492f
C5594 vdd.n3341 gnd 0.01055f
C5595 vdd.n3342 gnd 0.01055f
C5596 vdd.n3343 gnd 0.008492f
C5597 vdd.n3344 gnd 0.008492f
C5598 vdd.n3345 gnd 0.01055f
C5599 vdd.n3346 gnd 0.01055f
C5600 vdd.n3347 gnd 0.008492f
C5601 vdd.n3348 gnd 0.008492f
C5602 vdd.n3349 gnd 0.01055f
C5603 vdd.n3350 gnd 0.01055f
C5604 vdd.n3351 gnd 0.008492f
C5605 vdd.n3352 gnd 0.008492f
C5606 vdd.n3353 gnd 0.01055f
C5607 vdd.n3354 gnd 0.01055f
C5608 vdd.n3355 gnd 0.008492f
C5609 vdd.n3356 gnd 0.008492f
C5610 vdd.n3357 gnd 0.01055f
C5611 vdd.n3358 gnd 0.01055f
C5612 vdd.n3359 gnd 0.008492f
C5613 vdd.n3360 gnd 0.01055f
C5614 vdd.n3361 gnd 0.01055f
C5615 vdd.n3362 gnd 0.008492f
C5616 vdd.n3363 gnd 0.01055f
C5617 vdd.n3364 gnd 0.01055f
C5618 vdd.n3365 gnd 0.01055f
C5619 vdd.t80 gnd 0.129799f
C5620 vdd.t81 gnd 0.138719f
C5621 vdd.t79 gnd 0.169516f
C5622 vdd.n3366 gnd 0.217295f
C5623 vdd.n3367 gnd 0.182567f
C5624 vdd.n3368 gnd 0.017323f
C5625 vdd.n3369 gnd 0.01055f
C5626 vdd.n3370 gnd 0.01055f
C5627 vdd.n3371 gnd 0.007091f
C5628 vdd.n3372 gnd 0.008492f
C5629 vdd.n3373 gnd 0.01055f
C5630 vdd.n3374 gnd 0.01055f
C5631 vdd.n3375 gnd 0.008492f
C5632 vdd.n3376 gnd 0.008492f
C5633 vdd.n3377 gnd 0.01055f
C5634 vdd.n3378 gnd 0.01055f
C5635 vdd.n3379 gnd 0.008492f
C5636 vdd.n3380 gnd 0.008492f
C5637 vdd.n3381 gnd 0.01055f
C5638 vdd.n3382 gnd 0.01055f
C5639 vdd.n3383 gnd 0.008492f
C5640 vdd.n3384 gnd 0.008492f
C5641 vdd.n3385 gnd 0.01055f
C5642 vdd.n3386 gnd 0.01055f
C5643 vdd.n3387 gnd 0.008492f
C5644 vdd.n3388 gnd 0.008492f
C5645 vdd.n3389 gnd 0.01055f
C5646 vdd.n3390 gnd 0.01055f
C5647 vdd.n3391 gnd 0.008492f
C5648 vdd.n3392 gnd 0.008492f
C5649 vdd.n3393 gnd 0.01055f
C5650 vdd.n3394 gnd 0.01055f
C5651 vdd.n3395 gnd 0.008492f
C5652 vdd.n3396 gnd 0.008492f
C5653 vdd.n3398 gnd 0.963832f
C5654 vdd.n3400 gnd 0.008492f
C5655 vdd.n3401 gnd 0.008492f
C5656 vdd.n3402 gnd 0.007048f
C5657 vdd.n3403 gnd 0.026069f
C5658 vdd.n3405 gnd 11.375099f
C5659 vdd.n3406 gnd 0.026069f
C5660 vdd.n3407 gnd 0.004034f
C5661 vdd.n3408 gnd 0.026069f
C5662 vdd.n3409 gnd 0.025523f
C5663 vdd.n3410 gnd 0.01055f
C5664 vdd.n3411 gnd 0.008492f
C5665 vdd.n3412 gnd 0.01055f
C5666 vdd.n3413 gnd 0.652318f
C5667 vdd.n3414 gnd 0.01055f
C5668 vdd.n3415 gnd 0.008492f
C5669 vdd.n3416 gnd 0.01055f
C5670 vdd.n3417 gnd 0.01055f
C5671 vdd.n3418 gnd 0.01055f
C5672 vdd.n3419 gnd 0.008492f
C5673 vdd.n3420 gnd 0.01055f
C5674 vdd.n3421 gnd 1.07821f
C5675 vdd.n3422 gnd 0.01055f
C5676 vdd.n3423 gnd 0.008492f
C5677 vdd.n3424 gnd 0.01055f
C5678 vdd.n3425 gnd 0.01055f
C5679 vdd.n3426 gnd 0.01055f
C5680 vdd.n3427 gnd 0.008492f
C5681 vdd.n3428 gnd 0.01055f
C5682 vdd.n3429 gnd 0.695447f
C5683 vdd.n3430 gnd 0.738575f
C5684 vdd.n3431 gnd 0.01055f
C5685 vdd.n3432 gnd 0.008492f
C5686 vdd.n3433 gnd 0.01055f
C5687 vdd.n3434 gnd 0.01055f
C5688 vdd.n3435 gnd 0.01055f
C5689 vdd.n3436 gnd 0.008492f
C5690 vdd.n3437 gnd 0.01055f
C5691 vdd.n3438 gnd 0.894916f
C5692 vdd.n3439 gnd 0.01055f
C5693 vdd.n3440 gnd 0.008492f
C5694 vdd.n3441 gnd 0.01055f
C5695 vdd.n3442 gnd 0.01055f
C5696 vdd.n3443 gnd 0.01055f
C5697 vdd.n3444 gnd 0.008492f
C5698 vdd.n3445 gnd 0.01055f
C5699 vdd.t163 gnd 0.539106f
C5700 vdd.n3446 gnd 0.867961f
C5701 vdd.n3447 gnd 0.01055f
C5702 vdd.n3448 gnd 0.008492f
C5703 vdd.n3449 gnd 0.01055f
C5704 vdd.n3450 gnd 0.01055f
C5705 vdd.n3451 gnd 0.01055f
C5706 vdd.n3452 gnd 0.008492f
C5707 vdd.n3453 gnd 0.01055f
C5708 vdd.n3454 gnd 0.684665f
C5709 vdd.n3455 gnd 0.01055f
C5710 vdd.n3456 gnd 0.008492f
C5711 vdd.n3457 gnd 0.01055f
C5712 vdd.n3458 gnd 0.01055f
C5713 vdd.n3459 gnd 0.01055f
C5714 vdd.n3460 gnd 0.008492f
C5715 vdd.n3461 gnd 0.01055f
C5716 vdd.n3462 gnd 0.857178f
C5717 vdd.n3463 gnd 0.576843f
C5718 vdd.n3464 gnd 0.01055f
C5719 vdd.n3465 gnd 0.008492f
C5720 vdd.n3466 gnd 0.01055f
C5721 vdd.n3467 gnd 0.01055f
C5722 vdd.n3468 gnd 0.01055f
C5723 vdd.n3469 gnd 0.008492f
C5724 vdd.n3470 gnd 0.01055f
C5725 vdd.n3471 gnd 0.760139f
C5726 vdd.n3472 gnd 0.01055f
C5727 vdd.n3473 gnd 0.008492f
C5728 vdd.n3474 gnd 0.01055f
C5729 vdd.n3475 gnd 0.01055f
C5730 vdd.n3476 gnd 0.01055f
C5731 vdd.n3477 gnd 0.01055f
C5732 vdd.n3478 gnd 0.01055f
C5733 vdd.n3479 gnd 0.008492f
C5734 vdd.n3480 gnd 0.008492f
C5735 vdd.n3481 gnd 0.01055f
C5736 vdd.t254 gnd 0.539106f
C5737 vdd.n3482 gnd 0.894916f
C5738 vdd.n3483 gnd 0.01055f
C5739 vdd.n3484 gnd 0.008492f
C5740 vdd.n3485 gnd 0.01055f
C5741 vdd.n3486 gnd 0.01055f
C5742 vdd.n3487 gnd 0.01055f
C5743 vdd.n3488 gnd 0.008492f
C5744 vdd.n3489 gnd 0.01055f
C5745 vdd.n3490 gnd 0.846396f
C5746 vdd.n3491 gnd 0.01055f
C5747 vdd.n3492 gnd 0.01055f
C5748 vdd.n3493 gnd 0.008492f
C5749 vdd.n3494 gnd 0.008492f
C5750 vdd.n3495 gnd 0.01055f
C5751 vdd.n3496 gnd 0.01055f
C5752 vdd.n3497 gnd 0.01055f
C5753 vdd.n3498 gnd 0.008492f
C5754 vdd.n3499 gnd 0.01055f
C5755 vdd.n3500 gnd 0.008492f
C5756 vdd.n3501 gnd 0.008492f
C5757 vdd.n3502 gnd 0.01055f
C5758 vdd.n3503 gnd 0.01055f
C5759 vdd.n3504 gnd 0.01055f
C5760 vdd.n3505 gnd 0.008492f
C5761 vdd.n3506 gnd 0.01055f
C5762 vdd.n3507 gnd 0.008492f
C5763 vdd.n3508 gnd 0.008492f
C5764 vdd.n3509 gnd 0.01055f
C5765 vdd.n3510 gnd 0.01055f
C5766 vdd.n3511 gnd 0.01055f
C5767 vdd.n3512 gnd 0.008492f
C5768 vdd.n3513 gnd 0.894916f
C5769 vdd.n3514 gnd 0.01055f
C5770 vdd.n3515 gnd 0.008492f
C5771 vdd.n3516 gnd 0.008492f
C5772 vdd.n3517 gnd 0.01055f
C5773 vdd.n3518 gnd 0.01055f
C5774 vdd.n3519 gnd 0.01055f
C5775 vdd.n3520 gnd 0.008492f
C5776 vdd.n3521 gnd 0.01055f
C5777 vdd.n3522 gnd 0.008492f
C5778 vdd.n3523 gnd 0.008492f
C5779 vdd.n3524 gnd 0.01055f
C5780 vdd.n3525 gnd 0.01055f
C5781 vdd.n3526 gnd 0.01055f
C5782 vdd.n3527 gnd 0.008492f
C5783 vdd.n3528 gnd 0.01055f
C5784 vdd.n3529 gnd 0.008492f
C5785 vdd.n3530 gnd 0.007048f
C5786 vdd.n3531 gnd 0.025523f
C5787 vdd.n3532 gnd 0.026069f
C5788 vdd.n3533 gnd 0.004034f
C5789 vdd.n3534 gnd 0.026069f
C5790 vdd.n3536 gnd 2.55536f
C5791 vdd.n3537 gnd 1.59036f
C5792 vdd.n3538 gnd 0.025523f
C5793 vdd.n3539 gnd 0.007048f
C5794 vdd.n3540 gnd 0.008492f
C5795 vdd.n3541 gnd 0.008492f
C5796 vdd.n3542 gnd 0.01055f
C5797 vdd.n3543 gnd 1.07821f
C5798 vdd.n3544 gnd 1.07821f
C5799 vdd.n3545 gnd 0.986564f
C5800 vdd.n3546 gnd 0.01055f
C5801 vdd.n3547 gnd 0.008492f
C5802 vdd.n3548 gnd 0.008492f
C5803 vdd.n3549 gnd 0.008492f
C5804 vdd.n3550 gnd 0.01055f
C5805 vdd.n3551 gnd 0.803268f
C5806 vdd.t278 gnd 0.539106f
C5807 vdd.n3552 gnd 0.81405f
C5808 vdd.n3553 gnd 0.619972f
C5809 vdd.n3554 gnd 0.01055f
C5810 vdd.n3555 gnd 0.008492f
C5811 vdd.n3556 gnd 0.008492f
C5812 vdd.n3557 gnd 0.008492f
C5813 vdd.n3558 gnd 0.01055f
C5814 vdd.n3559 gnd 0.641536f
C5815 vdd.n3560 gnd 0.792486f
C5816 vdd.t159 gnd 0.539106f
C5817 vdd.n3561 gnd 0.824832f
C5818 vdd.n3562 gnd 0.01055f
C5819 vdd.n3563 gnd 0.008492f
C5820 vdd.n3564 gnd 0.008492f
C5821 vdd.n3565 gnd 0.008492f
C5822 vdd.n3566 gnd 0.01055f
C5823 vdd.n3567 gnd 0.894916f
C5824 vdd.t196 gnd 0.539106f
C5825 vdd.n3568 gnd 0.652318f
C5826 vdd.n3569 gnd 0.781704f
C5827 vdd.n3570 gnd 0.01055f
C5828 vdd.n3571 gnd 0.008492f
C5829 vdd.n3572 gnd 0.008492f
C5830 vdd.n3573 gnd 0.008492f
C5831 vdd.n3574 gnd 0.01055f
C5832 vdd.n3575 gnd 0.598408f
C5833 vdd.t208 gnd 0.539106f
C5834 vdd.n3576 gnd 0.894916f
C5835 vdd.t223 gnd 0.539106f
C5836 vdd.n3577 gnd 0.6631f
C5837 vdd.n3578 gnd 0.01055f
C5838 vdd.n3579 gnd 0.008492f
C5839 vdd.n3580 gnd 0.008109f
C5840 vdd.n3581 gnd 0.622309f
C5841 vdd.n3582 gnd 2.95346f
C5842 a_n8964_8799.n0 gnd 2.72898f
C5843 a_n8964_8799.n1 gnd 1.65342f
C5844 a_n8964_8799.n2 gnd 3.78285f
C5845 a_n8964_8799.n3 gnd 0.206316f
C5846 a_n8964_8799.n4 gnd 0.283299f
C5847 a_n8964_8799.n5 gnd 0.206316f
C5848 a_n8964_8799.n6 gnd 0.206316f
C5849 a_n8964_8799.n7 gnd 0.206316f
C5850 a_n8964_8799.n8 gnd 0.206316f
C5851 a_n8964_8799.n9 gnd 0.206316f
C5852 a_n8964_8799.n10 gnd 0.214532f
C5853 a_n8964_8799.n11 gnd 0.206316f
C5854 a_n8964_8799.n12 gnd 0.283299f
C5855 a_n8964_8799.n13 gnd 0.206316f
C5856 a_n8964_8799.n14 gnd 0.206316f
C5857 a_n8964_8799.n15 gnd 0.206316f
C5858 a_n8964_8799.n16 gnd 0.206316f
C5859 a_n8964_8799.n17 gnd 0.206316f
C5860 a_n8964_8799.n18 gnd 0.214532f
C5861 a_n8964_8799.n19 gnd 0.206316f
C5862 a_n8964_8799.n20 gnd 0.447177f
C5863 a_n8964_8799.n21 gnd 0.206316f
C5864 a_n8964_8799.n22 gnd 0.206316f
C5865 a_n8964_8799.n23 gnd 0.206316f
C5866 a_n8964_8799.n24 gnd 0.206316f
C5867 a_n8964_8799.n25 gnd 0.206316f
C5868 a_n8964_8799.n26 gnd 0.214532f
C5869 a_n8964_8799.n27 gnd 0.206316f
C5870 a_n8964_8799.n28 gnd 0.31769f
C5871 a_n8964_8799.n29 gnd 0.206316f
C5872 a_n8964_8799.n30 gnd 0.206316f
C5873 a_n8964_8799.n31 gnd 0.206316f
C5874 a_n8964_8799.n32 gnd 0.206316f
C5875 a_n8964_8799.n33 gnd 0.206316f
C5876 a_n8964_8799.n34 gnd 0.180141f
C5877 a_n8964_8799.n35 gnd 0.206316f
C5878 a_n8964_8799.n36 gnd 0.31769f
C5879 a_n8964_8799.n37 gnd 0.206316f
C5880 a_n8964_8799.n38 gnd 0.206316f
C5881 a_n8964_8799.n39 gnd 0.206316f
C5882 a_n8964_8799.n40 gnd 0.206316f
C5883 a_n8964_8799.n41 gnd 0.206316f
C5884 a_n8964_8799.n42 gnd 0.180141f
C5885 a_n8964_8799.n43 gnd 0.206316f
C5886 a_n8964_8799.n44 gnd 0.31769f
C5887 a_n8964_8799.n45 gnd 0.206316f
C5888 a_n8964_8799.n46 gnd 0.206316f
C5889 a_n8964_8799.n47 gnd 0.206316f
C5890 a_n8964_8799.n48 gnd 0.206316f
C5891 a_n8964_8799.n49 gnd 0.206316f
C5892 a_n8964_8799.n50 gnd 0.344019f
C5893 a_n8964_8799.n51 gnd 1.51213f
C5894 a_n8964_8799.n52 gnd 2.76027f
C5895 a_n8964_8799.n53 gnd 1.51214f
C5896 a_n8964_8799.n54 gnd 3.9057f
C5897 a_n8964_8799.n55 gnd 0.248385f
C5898 a_n8964_8799.n56 gnd 0.003631f
C5899 a_n8964_8799.n57 gnd 0.009572f
C5900 a_n8964_8799.n58 gnd 0.010458f
C5901 a_n8964_8799.n59 gnd 0.005526f
C5902 a_n8964_8799.n61 gnd 0.004637f
C5903 a_n8964_8799.n62 gnd 0.010029f
C5904 a_n8964_8799.n63 gnd 0.010029f
C5905 a_n8964_8799.n64 gnd 0.004637f
C5906 a_n8964_8799.n66 gnd 0.005526f
C5907 a_n8964_8799.n67 gnd 0.010458f
C5908 a_n8964_8799.n68 gnd 0.009572f
C5909 a_n8964_8799.n69 gnd 0.003631f
C5910 a_n8964_8799.n70 gnd 0.248385f
C5911 a_n8964_8799.n71 gnd 0.003631f
C5912 a_n8964_8799.n72 gnd 0.009572f
C5913 a_n8964_8799.n73 gnd 0.010458f
C5914 a_n8964_8799.n74 gnd 0.005526f
C5915 a_n8964_8799.n76 gnd 0.004637f
C5916 a_n8964_8799.n77 gnd 0.010029f
C5917 a_n8964_8799.n78 gnd 0.010029f
C5918 a_n8964_8799.n79 gnd 0.004637f
C5919 a_n8964_8799.n81 gnd 0.005526f
C5920 a_n8964_8799.n82 gnd 0.010458f
C5921 a_n8964_8799.n83 gnd 0.009572f
C5922 a_n8964_8799.n84 gnd 0.003631f
C5923 a_n8964_8799.n85 gnd 0.248385f
C5924 a_n8964_8799.n86 gnd 0.003631f
C5925 a_n8964_8799.n87 gnd 0.009572f
C5926 a_n8964_8799.n88 gnd 0.010458f
C5927 a_n8964_8799.n89 gnd 0.005526f
C5928 a_n8964_8799.n91 gnd 0.004637f
C5929 a_n8964_8799.n92 gnd 0.010029f
C5930 a_n8964_8799.n93 gnd 0.010029f
C5931 a_n8964_8799.n94 gnd 0.004637f
C5932 a_n8964_8799.n96 gnd 0.005526f
C5933 a_n8964_8799.n97 gnd 0.010458f
C5934 a_n8964_8799.n98 gnd 0.009572f
C5935 a_n8964_8799.n99 gnd 0.003631f
C5936 a_n8964_8799.n100 gnd 0.003631f
C5937 a_n8964_8799.n101 gnd 0.009572f
C5938 a_n8964_8799.n102 gnd 0.010458f
C5939 a_n8964_8799.n103 gnd 0.005526f
C5940 a_n8964_8799.n105 gnd 0.004637f
C5941 a_n8964_8799.n106 gnd 0.010029f
C5942 a_n8964_8799.n107 gnd 0.010029f
C5943 a_n8964_8799.n108 gnd 0.004637f
C5944 a_n8964_8799.n110 gnd 0.005526f
C5945 a_n8964_8799.n111 gnd 0.010458f
C5946 a_n8964_8799.n112 gnd 0.009572f
C5947 a_n8964_8799.n113 gnd 0.003631f
C5948 a_n8964_8799.n114 gnd 0.248385f
C5949 a_n8964_8799.n115 gnd 0.003631f
C5950 a_n8964_8799.n116 gnd 0.009572f
C5951 a_n8964_8799.n117 gnd 0.010458f
C5952 a_n8964_8799.n118 gnd 0.005526f
C5953 a_n8964_8799.n120 gnd 0.004637f
C5954 a_n8964_8799.n121 gnd 0.010029f
C5955 a_n8964_8799.n122 gnd 0.010029f
C5956 a_n8964_8799.n123 gnd 0.004637f
C5957 a_n8964_8799.n125 gnd 0.005526f
C5958 a_n8964_8799.n126 gnd 0.010458f
C5959 a_n8964_8799.n127 gnd 0.009572f
C5960 a_n8964_8799.n128 gnd 0.003631f
C5961 a_n8964_8799.n129 gnd 0.248385f
C5962 a_n8964_8799.n130 gnd 0.003631f
C5963 a_n8964_8799.n131 gnd 0.009572f
C5964 a_n8964_8799.n132 gnd 0.010458f
C5965 a_n8964_8799.n133 gnd 0.005526f
C5966 a_n8964_8799.n135 gnd 0.004637f
C5967 a_n8964_8799.n136 gnd 0.010029f
C5968 a_n8964_8799.n137 gnd 0.010029f
C5969 a_n8964_8799.n138 gnd 0.004637f
C5970 a_n8964_8799.n140 gnd 0.005526f
C5971 a_n8964_8799.n141 gnd 0.010458f
C5972 a_n8964_8799.n142 gnd 0.009572f
C5973 a_n8964_8799.n143 gnd 0.003631f
C5974 a_n8964_8799.n144 gnd 0.248385f
C5975 a_n8964_8799.t10 gnd 0.143103f
C5976 a_n8964_8799.t26 gnd 0.143103f
C5977 a_n8964_8799.t4 gnd 0.143103f
C5978 a_n8964_8799.n145 gnd 1.12868f
C5979 a_n8964_8799.t5 gnd 0.143103f
C5980 a_n8964_8799.t11 gnd 0.143103f
C5981 a_n8964_8799.n146 gnd 1.12682f
C5982 a_n8964_8799.t8 gnd 0.143103f
C5983 a_n8964_8799.t32 gnd 0.143103f
C5984 a_n8964_8799.n147 gnd 1.12682f
C5985 a_n8964_8799.t33 gnd 0.143103f
C5986 a_n8964_8799.t24 gnd 0.143103f
C5987 a_n8964_8799.n148 gnd 1.12682f
C5988 a_n8964_8799.t9 gnd 0.143103f
C5989 a_n8964_8799.t18 gnd 0.143103f
C5990 a_n8964_8799.n149 gnd 1.12682f
C5991 a_n8964_8799.t34 gnd 0.111303f
C5992 a_n8964_8799.t6 gnd 0.111303f
C5993 a_n8964_8799.n150 gnd 0.986409f
C5994 a_n8964_8799.t20 gnd 0.111303f
C5995 a_n8964_8799.t35 gnd 0.111303f
C5996 a_n8964_8799.n151 gnd 0.983508f
C5997 a_n8964_8799.t21 gnd 0.111303f
C5998 a_n8964_8799.t2 gnd 0.111303f
C5999 a_n8964_8799.n152 gnd 0.986408f
C6000 a_n8964_8799.t12 gnd 0.111303f
C6001 a_n8964_8799.t30 gnd 0.111303f
C6002 a_n8964_8799.n153 gnd 0.983508f
C6003 a_n8964_8799.t23 gnd 0.111303f
C6004 a_n8964_8799.t16 gnd 0.111303f
C6005 a_n8964_8799.n154 gnd 0.986408f
C6006 a_n8964_8799.t28 gnd 0.111303f
C6007 a_n8964_8799.t29 gnd 0.111303f
C6008 a_n8964_8799.n155 gnd 0.983508f
C6009 a_n8964_8799.t1 gnd 0.111303f
C6010 a_n8964_8799.t19 gnd 0.111303f
C6011 a_n8964_8799.n156 gnd 0.983508f
C6012 a_n8964_8799.t22 gnd 0.111303f
C6013 a_n8964_8799.t15 gnd 0.111303f
C6014 a_n8964_8799.n157 gnd 0.983508f
C6015 a_n8964_8799.t69 gnd 0.593373f
C6016 a_n8964_8799.n158 gnd 0.267144f
C6017 a_n8964_8799.t114 gnd 0.593373f
C6018 a_n8964_8799.t137 gnd 0.593373f
C6019 a_n8964_8799.n159 gnd 0.269058f
C6020 a_n8964_8799.t82 gnd 0.593373f
C6021 a_n8964_8799.t85 gnd 0.593373f
C6022 a_n8964_8799.n160 gnd 0.262309f
C6023 a_n8964_8799.t138 gnd 0.593373f
C6024 a_n8964_8799.t143 gnd 0.593373f
C6025 a_n8964_8799.n161 gnd 0.266258f
C6026 a_n8964_8799.t68 gnd 0.593373f
C6027 a_n8964_8799.t113 gnd 0.593373f
C6028 a_n8964_8799.t83 gnd 0.604603f
C6029 a_n8964_8799.n162 gnd 0.248746f
C6030 a_n8964_8799.n163 gnd 0.269428f
C6031 a_n8964_8799.t40 gnd 0.593373f
C6032 a_n8964_8799.n164 gnd 0.267144f
C6033 a_n8964_8799.n165 gnd 0.262945f
C6034 a_n8964_8799.t106 gnd 0.593373f
C6035 a_n8964_8799.n166 gnd 0.261673f
C6036 a_n8964_8799.t66 gnd 0.593373f
C6037 a_n8964_8799.n167 gnd 0.268805f
C6038 a_n8964_8799.t101 gnd 0.593373f
C6039 a_n8964_8799.n168 gnd 0.269058f
C6040 a_n8964_8799.n169 gnd 0.266687f
C6041 a_n8964_8799.t139 gnd 0.593373f
C6042 a_n8964_8799.n170 gnd 0.262309f
C6043 a_n8964_8799.t117 gnd 0.593373f
C6044 a_n8964_8799.n171 gnd 0.266687f
C6045 a_n8964_8799.n172 gnd 0.268805f
C6046 a_n8964_8799.t84 gnd 0.593373f
C6047 a_n8964_8799.n173 gnd 0.266258f
C6048 a_n8964_8799.n174 gnd 0.261673f
C6049 a_n8964_8799.t67 gnd 0.593373f
C6050 a_n8964_8799.n175 gnd 0.262945f
C6051 a_n8964_8799.t110 gnd 0.593373f
C6052 a_n8964_8799.n176 gnd 0.269428f
C6053 a_n8964_8799.t36 gnd 0.604593f
C6054 a_n8964_8799.t80 gnd 0.593373f
C6055 a_n8964_8799.n177 gnd 0.267144f
C6056 a_n8964_8799.t131 gnd 0.593373f
C6057 a_n8964_8799.t150 gnd 0.593373f
C6058 a_n8964_8799.n178 gnd 0.269058f
C6059 a_n8964_8799.t92 gnd 0.593373f
C6060 a_n8964_8799.t97 gnd 0.593373f
C6061 a_n8964_8799.n179 gnd 0.262309f
C6062 a_n8964_8799.t152 gnd 0.593373f
C6063 a_n8964_8799.t155 gnd 0.593373f
C6064 a_n8964_8799.n180 gnd 0.266258f
C6065 a_n8964_8799.t79 gnd 0.593373f
C6066 a_n8964_8799.t130 gnd 0.593373f
C6067 a_n8964_8799.t93 gnd 0.604603f
C6068 a_n8964_8799.n181 gnd 0.248746f
C6069 a_n8964_8799.n182 gnd 0.269428f
C6070 a_n8964_8799.t52 gnd 0.593373f
C6071 a_n8964_8799.n183 gnd 0.267144f
C6072 a_n8964_8799.n184 gnd 0.262945f
C6073 a_n8964_8799.t121 gnd 0.593373f
C6074 a_n8964_8799.n185 gnd 0.261673f
C6075 a_n8964_8799.t75 gnd 0.593373f
C6076 a_n8964_8799.n186 gnd 0.268805f
C6077 a_n8964_8799.t115 gnd 0.593373f
C6078 a_n8964_8799.n187 gnd 0.269058f
C6079 a_n8964_8799.n188 gnd 0.266687f
C6080 a_n8964_8799.t154 gnd 0.593373f
C6081 a_n8964_8799.n189 gnd 0.262309f
C6082 a_n8964_8799.t134 gnd 0.593373f
C6083 a_n8964_8799.n190 gnd 0.266687f
C6084 a_n8964_8799.n191 gnd 0.268805f
C6085 a_n8964_8799.t94 gnd 0.593373f
C6086 a_n8964_8799.n192 gnd 0.266258f
C6087 a_n8964_8799.n193 gnd 0.261673f
C6088 a_n8964_8799.t78 gnd 0.593373f
C6089 a_n8964_8799.n194 gnd 0.262945f
C6090 a_n8964_8799.t128 gnd 0.593373f
C6091 a_n8964_8799.n195 gnd 0.269428f
C6092 a_n8964_8799.t48 gnd 0.604593f
C6093 a_n8964_8799.n196 gnd 0.892053f
C6094 a_n8964_8799.t116 gnd 0.593373f
C6095 a_n8964_8799.n197 gnd 0.267144f
C6096 a_n8964_8799.t98 gnd 0.593373f
C6097 a_n8964_8799.t140 gnd 0.593373f
C6098 a_n8964_8799.n198 gnd 0.269058f
C6099 a_n8964_8799.t58 gnd 0.593373f
C6100 a_n8964_8799.t133 gnd 0.593373f
C6101 a_n8964_8799.n199 gnd 0.262309f
C6102 a_n8964_8799.t111 gnd 0.593373f
C6103 a_n8964_8799.t71 gnd 0.593373f
C6104 a_n8964_8799.n200 gnd 0.266258f
C6105 a_n8964_8799.t56 gnd 0.593373f
C6106 a_n8964_8799.t41 gnd 0.593373f
C6107 a_n8964_8799.t86 gnd 0.604603f
C6108 a_n8964_8799.n201 gnd 0.248746f
C6109 a_n8964_8799.n202 gnd 0.269428f
C6110 a_n8964_8799.t102 gnd 0.593373f
C6111 a_n8964_8799.n203 gnd 0.267144f
C6112 a_n8964_8799.n204 gnd 0.262945f
C6113 a_n8964_8799.t123 gnd 0.593373f
C6114 a_n8964_8799.n205 gnd 0.261673f
C6115 a_n8964_8799.t95 gnd 0.593373f
C6116 a_n8964_8799.n206 gnd 0.268805f
C6117 a_n8964_8799.t49 gnd 0.593373f
C6118 a_n8964_8799.n207 gnd 0.269058f
C6119 a_n8964_8799.n208 gnd 0.266687f
C6120 a_n8964_8799.t90 gnd 0.593373f
C6121 a_n8964_8799.n209 gnd 0.262309f
C6122 a_n8964_8799.t76 gnd 0.593373f
C6123 a_n8964_8799.n210 gnd 0.266687f
C6124 a_n8964_8799.n211 gnd 0.268805f
C6125 a_n8964_8799.t37 gnd 0.593373f
C6126 a_n8964_8799.n212 gnd 0.266258f
C6127 a_n8964_8799.n213 gnd 0.261673f
C6128 a_n8964_8799.t142 gnd 0.593373f
C6129 a_n8964_8799.n214 gnd 0.262945f
C6130 a_n8964_8799.t149 gnd 0.593373f
C6131 a_n8964_8799.n215 gnd 0.269428f
C6132 a_n8964_8799.t91 gnd 0.604593f
C6133 a_n8964_8799.n216 gnd 1.68955f
C6134 a_n8964_8799.t103 gnd 0.604593f
C6135 a_n8964_8799.t39 gnd 0.593373f
C6136 a_n8964_8799.t109 gnd 0.593373f
C6137 a_n8964_8799.n217 gnd 0.267144f
C6138 a_n8964_8799.t107 gnd 0.593373f
C6139 a_n8964_8799.t45 gnd 0.593373f
C6140 a_n8964_8799.t43 gnd 0.593373f
C6141 a_n8964_8799.n218 gnd 0.266258f
C6142 a_n8964_8799.t129 gnd 0.593373f
C6143 a_n8964_8799.t61 gnd 0.593373f
C6144 a_n8964_8799.t47 gnd 0.593373f
C6145 a_n8964_8799.n219 gnd 0.266687f
C6146 a_n8964_8799.t135 gnd 0.593373f
C6147 a_n8964_8799.t87 gnd 0.593373f
C6148 a_n8964_8799.t62 gnd 0.593373f
C6149 a_n8964_8799.n220 gnd 0.266687f
C6150 a_n8964_8799.t153 gnd 0.593373f
C6151 a_n8964_8799.t105 gnd 0.593373f
C6152 a_n8964_8799.t64 gnd 0.593373f
C6153 a_n8964_8799.n221 gnd 0.266258f
C6154 a_n8964_8799.t147 gnd 0.593373f
C6155 a_n8964_8799.t108 gnd 0.593373f
C6156 a_n8964_8799.t81 gnd 0.593373f
C6157 a_n8964_8799.n222 gnd 0.267144f
C6158 a_n8964_8799.t132 gnd 0.604603f
C6159 a_n8964_8799.n223 gnd 0.248746f
C6160 a_n8964_8799.t44 gnd 0.593373f
C6161 a_n8964_8799.n224 gnd 0.269428f
C6162 a_n8964_8799.n225 gnd 0.262945f
C6163 a_n8964_8799.n226 gnd 0.261673f
C6164 a_n8964_8799.n227 gnd 0.268805f
C6165 a_n8964_8799.n228 gnd 0.269058f
C6166 a_n8964_8799.n229 gnd 0.262309f
C6167 a_n8964_8799.n230 gnd 0.262309f
C6168 a_n8964_8799.n231 gnd 0.269058f
C6169 a_n8964_8799.n232 gnd 0.268805f
C6170 a_n8964_8799.n233 gnd 0.261673f
C6171 a_n8964_8799.n234 gnd 0.262945f
C6172 a_n8964_8799.n235 gnd 0.269428f
C6173 a_n8964_8799.t119 gnd 0.604593f
C6174 a_n8964_8799.t51 gnd 0.593373f
C6175 a_n8964_8799.t127 gnd 0.593373f
C6176 a_n8964_8799.n236 gnd 0.267144f
C6177 a_n8964_8799.t125 gnd 0.593373f
C6178 a_n8964_8799.t54 gnd 0.593373f
C6179 a_n8964_8799.t53 gnd 0.593373f
C6180 a_n8964_8799.n237 gnd 0.266258f
C6181 a_n8964_8799.t145 gnd 0.593373f
C6182 a_n8964_8799.t70 gnd 0.593373f
C6183 a_n8964_8799.t60 gnd 0.593373f
C6184 a_n8964_8799.n238 gnd 0.266687f
C6185 a_n8964_8799.t148 gnd 0.593373f
C6186 a_n8964_8799.t100 gnd 0.593373f
C6187 a_n8964_8799.t73 gnd 0.593373f
C6188 a_n8964_8799.n239 gnd 0.266687f
C6189 a_n8964_8799.t46 gnd 0.593373f
C6190 a_n8964_8799.t120 gnd 0.593373f
C6191 a_n8964_8799.t74 gnd 0.593373f
C6192 a_n8964_8799.n240 gnd 0.266258f
C6193 a_n8964_8799.t38 gnd 0.593373f
C6194 a_n8964_8799.t126 gnd 0.593373f
C6195 a_n8964_8799.t89 gnd 0.593373f
C6196 a_n8964_8799.n241 gnd 0.267144f
C6197 a_n8964_8799.t146 gnd 0.604603f
C6198 a_n8964_8799.n242 gnd 0.248746f
C6199 a_n8964_8799.t55 gnd 0.593373f
C6200 a_n8964_8799.n243 gnd 0.269428f
C6201 a_n8964_8799.n244 gnd 0.262945f
C6202 a_n8964_8799.n245 gnd 0.261673f
C6203 a_n8964_8799.n246 gnd 0.268805f
C6204 a_n8964_8799.n247 gnd 0.269058f
C6205 a_n8964_8799.n248 gnd 0.262309f
C6206 a_n8964_8799.n249 gnd 0.262309f
C6207 a_n8964_8799.n250 gnd 0.269058f
C6208 a_n8964_8799.n251 gnd 0.268805f
C6209 a_n8964_8799.n252 gnd 0.261673f
C6210 a_n8964_8799.n253 gnd 0.262945f
C6211 a_n8964_8799.n254 gnd 0.269428f
C6212 a_n8964_8799.n255 gnd 0.892053f
C6213 a_n8964_8799.t65 gnd 0.604593f
C6214 a_n8964_8799.t151 gnd 0.593373f
C6215 a_n8964_8799.t118 gnd 0.593373f
C6216 a_n8964_8799.n256 gnd 0.267144f
C6217 a_n8964_8799.t144 gnd 0.593373f
C6218 a_n8964_8799.t99 gnd 0.593373f
C6219 a_n8964_8799.t124 gnd 0.593373f
C6220 a_n8964_8799.n257 gnd 0.266258f
C6221 a_n8964_8799.t59 gnd 0.593373f
C6222 a_n8964_8799.t141 gnd 0.593373f
C6223 a_n8964_8799.t77 gnd 0.593373f
C6224 a_n8964_8799.n258 gnd 0.266687f
C6225 a_n8964_8799.t136 gnd 0.593373f
C6226 a_n8964_8799.t63 gnd 0.593373f
C6227 a_n8964_8799.t112 gnd 0.593373f
C6228 a_n8964_8799.n259 gnd 0.266687f
C6229 a_n8964_8799.t50 gnd 0.593373f
C6230 a_n8964_8799.t96 gnd 0.593373f
C6231 a_n8964_8799.t72 gnd 0.593373f
C6232 a_n8964_8799.n260 gnd 0.266258f
C6233 a_n8964_8799.t122 gnd 0.593373f
C6234 a_n8964_8799.t57 gnd 0.593373f
C6235 a_n8964_8799.t104 gnd 0.593373f
C6236 a_n8964_8799.n261 gnd 0.267144f
C6237 a_n8964_8799.t88 gnd 0.604603f
C6238 a_n8964_8799.n262 gnd 0.248746f
C6239 a_n8964_8799.t42 gnd 0.593373f
C6240 a_n8964_8799.n263 gnd 0.269428f
C6241 a_n8964_8799.n264 gnd 0.262945f
C6242 a_n8964_8799.n265 gnd 0.261673f
C6243 a_n8964_8799.n266 gnd 0.268805f
C6244 a_n8964_8799.n267 gnd 0.269058f
C6245 a_n8964_8799.n268 gnd 0.262309f
C6246 a_n8964_8799.n269 gnd 0.262309f
C6247 a_n8964_8799.n270 gnd 0.269058f
C6248 a_n8964_8799.n271 gnd 0.268805f
C6249 a_n8964_8799.n272 gnd 0.261673f
C6250 a_n8964_8799.n273 gnd 0.262945f
C6251 a_n8964_8799.n274 gnd 0.269428f
C6252 a_n8964_8799.n275 gnd 1.30305f
C6253 a_n8964_8799.n276 gnd 15.571901f
C6254 a_n8964_8799.n277 gnd 4.34263f
C6255 a_n8964_8799.n278 gnd 6.93963f
C6256 a_n8964_8799.t7 gnd 0.143103f
C6257 a_n8964_8799.t25 gnd 0.143103f
C6258 a_n8964_8799.n279 gnd 1.12867f
C6259 a_n8964_8799.t27 gnd 0.143103f
C6260 a_n8964_8799.t3 gnd 0.143103f
C6261 a_n8964_8799.n280 gnd 1.12682f
C6262 a_n8964_8799.t13 gnd 0.143103f
C6263 a_n8964_8799.t14 gnd 0.143103f
C6264 a_n8964_8799.n281 gnd 1.12682f
C6265 a_n8964_8799.t31 gnd 0.143103f
C6266 a_n8964_8799.t17 gnd 0.143103f
C6267 a_n8964_8799.n282 gnd 1.12682f
C6268 a_n8964_8799.n283 gnd 1.12682f
C6269 a_n8964_8799.t0 gnd 0.143103f
.ends

