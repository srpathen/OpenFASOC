* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 gnd.t221 gnd.t218 gnd.t220 gnd.t219 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X1 commonsourceibias.t47 commonsourceibias.t46 gnd.t269 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X2 gnd.t235 commonsourceibias.t48 CSoutput.t127 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X3 gnd.t217 gnd.t215 gnd.t216 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X4 vdd.t138 a_n6972_8799.t36 CSoutput.t63 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X5 a_n1986_8322.t19 a_n2848_n452.t48 vdd.t154 vdd.t153 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X6 a_n1808_13878.t11 a_n2848_n452.t45 a_n2848_n452.t46 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X7 a_n6972_8799.t20 plus.t5 a_n3106_n452.t27 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X8 output.t3 outputibias.t8 gnd.t101 gnd.t100 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X9 gnd.t92 commonsourceibias.t49 CSoutput.t126 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X10 a_n3106_n452.t26 plus.t6 a_n6972_8799.t11 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X11 vdd.t164 CSoutput.t144 output.t19 gnd.t93 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X12 a_n2848_n452.t40 a_n2848_n452.t39 a_n1808_13878.t10 vdd.t142 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 a_n1808_13878.t9 a_n2848_n452.t43 a_n2848_n452.t44 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X14 vdd.t255 vdd.t253 vdd.t254 vdd.t231 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X15 CSoutput.t76 a_n6972_8799.t37 vdd.t137 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X16 a_n1808_13878.t19 a_n2848_n452.t49 vdd.t156 vdd.t155 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 gnd.t53 commonsourceibias.t44 commonsourceibias.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 vdd.t176 CSoutput.t145 output.t18 gnd.t94 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X19 vdd.t252 vdd.t250 vdd.t251 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X20 CSoutput.t56 a_n6972_8799.t38 vdd.t136 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 vdd.t135 a_n6972_8799.t39 CSoutput.t44 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 gnd.t63 commonsourceibias.t50 CSoutput.t125 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 outputibias.t7 outputibias.t6 gnd.t262 gnd.t261 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X24 CSoutput.t20 a_n6972_8799.t40 vdd.t134 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X25 a_n1986_8322.t11 a_n2848_n452.t50 a_n6972_8799.t12 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X26 a_n2848_n452.t17 minus.t5 a_n3106_n452.t49 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 a_n6972_8799.t5 plus.t7 a_n3106_n452.t25 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X28 gnd.t90 commonsourceibias.t42 commonsourceibias.t43 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X29 CSoutput.t69 a_n6972_8799.t41 vdd.t133 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 plus.t4 gnd.t212 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X31 a_n2848_n452.t16 minus.t6 a_n3106_n452.t48 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X32 vdd.t132 a_n6972_8799.t42 CSoutput.t134 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X33 CSoutput.t124 commonsourceibias.t51 gnd.t43 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 CSoutput.t146 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X35 gnd.t227 commonsourceibias.t40 commonsourceibias.t41 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X36 CSoutput.t74 a_n6972_8799.t43 vdd.t131 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 vdd.t130 a_n6972_8799.t44 CSoutput.t0 vdd.t96 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 a_n3106_n452.t24 plus.t8 a_n6972_8799.t32 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X39 a_n6972_8799.t13 a_n2848_n452.t51 a_n1986_8322.t10 vdd.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X40 CSoutput.t67 a_n6972_8799.t45 vdd.t129 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X41 vdd.t128 a_n6972_8799.t46 CSoutput.t42 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X42 a_n3106_n452.t47 minus.t7 a_n2848_n452.t15 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X43 CSoutput.t123 commonsourceibias.t52 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 a_n3106_n452.t0 diffpairibias.t16 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X45 output.t17 CSoutput.t147 vdd.t172 gnd.t283 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X46 vdd.t170 CSoutput.t148 output.t16 gnd.t284 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X47 CSoutput.t122 commonsourceibias.t53 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 CSoutput.t24 a_n6972_8799.t47 vdd.t127 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X49 CSoutput.t128 a_n6972_8799.t48 vdd.t126 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X50 vdd.t249 vdd.t247 vdd.t248 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X51 vdd.t246 vdd.t244 vdd.t245 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X52 CSoutput.t121 commonsourceibias.t54 gnd.t291 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X53 gnd.t211 gnd.t209 gnd.t210 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X54 CSoutput.t4 a_n6972_8799.t49 vdd.t125 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 a_n3106_n452.t23 plus.t9 a_n6972_8799.t17 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X56 a_n1808_13878.t8 a_n2848_n452.t33 a_n2848_n452.t34 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X57 vdd.t124 a_n6972_8799.t50 CSoutput.t2 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X58 a_n3106_n452.t22 plus.t10 a_n6972_8799.t26 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X59 a_n3106_n452.t46 minus.t8 a_n2848_n452.t14 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X60 diffpairibias.t15 diffpairibias.t14 gnd.t229 gnd.t228 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 a_n2848_n452.t36 a_n2848_n452.t35 a_n1808_13878.t7 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X62 CSoutput.t78 a_n6972_8799.t51 vdd.t123 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X63 gnd.t208 gnd.t206 gnd.t207 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X64 vdd.t243 vdd.t241 vdd.t242 vdd.t216 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X65 CSoutput.t71 a_n6972_8799.t52 vdd.t122 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 vdd.t121 a_n6972_8799.t53 CSoutput.t129 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X67 gnd.t12 commonsourceibias.t55 CSoutput.t120 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X68 gnd.t106 commonsourceibias.t56 CSoutput.t119 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 diffpairibias.t13 diffpairibias.t12 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X70 CSoutput.t130 a_n6972_8799.t54 vdd.t120 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 gnd.t287 commonsourceibias.t57 CSoutput.t118 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X72 commonsourceibias.t39 commonsourceibias.t38 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X73 vdd.t119 a_n6972_8799.t55 CSoutput.t22 vdd.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 vdd.t117 a_n6972_8799.t56 CSoutput.t131 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X75 vdd.t178 CSoutput.t149 output.t15 gnd.t285 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X76 CSoutput.t135 a_n6972_8799.t57 vdd.t116 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X77 vdd.t115 a_n6972_8799.t58 CSoutput.t10 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X78 CSoutput.t23 a_n6972_8799.t59 vdd.t114 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X79 a_n3106_n452.t45 minus.t9 a_n2848_n452.t13 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X80 a_n3106_n452.t21 plus.t11 a_n6972_8799.t15 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X81 vdd.t113 a_n6972_8799.t60 CSoutput.t34 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 gnd.t248 commonsourceibias.t58 CSoutput.t117 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X83 a_n6972_8799.t16 plus.t12 a_n3106_n452.t20 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X84 commonsourceibias.t37 commonsourceibias.t36 gnd.t257 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 CSoutput.t133 a_n6972_8799.t61 vdd.t112 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 CSoutput.t50 a_n6972_8799.t62 vdd.t111 vdd.t100 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 a_n3106_n452.t43 diffpairibias.t17 gnd.t253 gnd.t252 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X88 gnd.t282 commonsourceibias.t34 commonsourceibias.t35 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X89 CSoutput.t39 a_n6972_8799.t63 vdd.t110 vdd.t100 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X90 a_n3106_n452.t19 plus.t13 a_n6972_8799.t31 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X91 vdd.t109 a_n6972_8799.t64 CSoutput.t29 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X92 gnd.t36 commonsourceibias.t32 commonsourceibias.t33 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X93 commonsourceibias.t31 commonsourceibias.t30 gnd.t73 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n2848_n452.t24 a_n2848_n452.t23 a_n1808_13878.t6 vdd.t147 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X95 outputibias.t5 outputibias.t4 gnd.t274 gnd.t273 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X96 a_n2848_n452.t26 a_n2848_n452.t25 a_n1808_13878.t5 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X97 vdd.t108 a_n6972_8799.t65 CSoutput.t141 vdd.t96 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X98 vdd.t107 a_n6972_8799.t66 CSoutput.t51 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n6972_8799.t2 a_n2848_n452.t52 a_n1986_8322.t9 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 CSoutput.t116 commonsourceibias.t59 gnd.t104 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X101 vdd.t106 a_n6972_8799.t67 CSoutput.t40 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n2848_n452.t18 minus.t10 a_n3106_n452.t50 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X103 CSoutput.t115 commonsourceibias.t60 gnd.t87 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 vdd.t105 a_n6972_8799.t68 CSoutput.t54 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 gnd.t78 commonsourceibias.t61 CSoutput.t114 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X106 gnd.t205 gnd.t202 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X107 commonsourceibias.t29 commonsourceibias.t28 gnd.t279 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 CSoutput.t58 a_n6972_8799.t69 vdd.t104 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X109 CSoutput.t113 commonsourceibias.t62 gnd.t264 gnd.t263 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X110 CSoutput.t150 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X111 outputibias.t3 outputibias.t2 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X112 vdd.t103 a_n6972_8799.t70 CSoutput.t45 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X113 vdd.t240 vdd.t238 vdd.t239 vdd.t224 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X114 CSoutput.t77 a_n6972_8799.t71 vdd.t102 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X115 vdd.t237 vdd.t234 vdd.t236 vdd.t235 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X116 a_n3106_n452.t31 diffpairibias.t18 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X117 vdd.t233 vdd.t230 vdd.t232 vdd.t231 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X118 gnd.t201 gnd.t199 minus.t4 gnd.t200 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X119 gnd.t198 gnd.t196 gnd.t197 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X120 commonsourceibias.t27 commonsourceibias.t26 gnd.t89 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X121 vdd.t2 a_n2848_n452.t53 a_n1986_8322.t18 vdd.t1 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X122 vdd.t229 vdd.t227 vdd.t228 vdd.t220 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X123 CSoutput.t79 a_n6972_8799.t72 vdd.t101 vdd.t100 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X124 a_n1986_8322.t17 a_n2848_n452.t54 vdd.t261 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X125 vdd.t99 a_n6972_8799.t73 CSoutput.t28 vdd.t98 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 gnd.t266 commonsourceibias.t24 commonsourceibias.t25 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t281 commonsourceibias.t63 CSoutput.t112 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 vdd.t263 a_n2848_n452.t55 a_n1808_13878.t18 vdd.t262 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X129 gnd.t195 gnd.t193 plus.t3 gnd.t194 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X130 gnd.t26 commonsourceibias.t64 CSoutput.t111 gnd.t25 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X131 a_n2848_n452.t22 minus.t11 a_n3106_n452.t54 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X132 a_n6972_8799.t33 plus.t14 a_n3106_n452.t18 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X133 gnd.t265 commonsourceibias.t65 CSoutput.t110 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X134 vdd.t226 vdd.t223 vdd.t225 vdd.t224 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X135 a_n6972_8799.t23 plus.t15 a_n3106_n452.t17 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X136 a_n2848_n452.t21 minus.t12 a_n3106_n452.t53 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X137 diffpairibias.t11 diffpairibias.t10 gnd.t40 gnd.t39 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X138 vdd.t175 CSoutput.t151 output.t14 gnd.t68 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X139 vdd.t222 vdd.t219 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 vdd.t97 a_n6972_8799.t74 CSoutput.t143 vdd.t96 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 gnd.t267 commonsourceibias.t66 CSoutput.t109 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 outputibias.t1 outputibias.t0 gnd.t278 gnd.t277 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X143 a_n6972_8799.t22 a_n2848_n452.t56 a_n1986_8322.t8 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 a_n1986_8322.t16 a_n2848_n452.t57 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X145 vdd.t218 vdd.t215 vdd.t217 vdd.t216 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X146 gnd.t247 commonsourceibias.t67 CSoutput.t108 gnd.t246 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 vdd.t95 a_n6972_8799.t75 CSoutput.t49 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 a_n2848_n452.t42 a_n2848_n452.t41 a_n1808_13878.t4 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X149 a_n3106_n452.t52 minus.t13 a_n2848_n452.t20 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X150 CSoutput.t152 a_n1986_8322.t23 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X151 CSoutput.t30 a_n6972_8799.t76 vdd.t94 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X152 a_n6972_8799.t9 a_n2848_n452.t58 a_n1986_8322.t7 vdd.t10 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 CSoutput.t107 commonsourceibias.t68 gnd.t237 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 CSoutput.t153 a_n1986_8322.t22 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X155 a_n1808_13878.t3 a_n2848_n452.t27 a_n2848_n452.t28 vdd.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X156 a_n3106_n452.t16 plus.t16 a_n6972_8799.t35 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X157 a_n2848_n452.t19 minus.t14 a_n3106_n452.t51 gnd.t99 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X158 vdd.t93 a_n6972_8799.t77 CSoutput.t138 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 CSoutput.t32 a_n6972_8799.t78 vdd.t92 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X160 vdd.t141 a_n2848_n452.t59 a_n1986_8322.t15 vdd.t140 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X161 gnd.t192 gnd.t189 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X162 a_n3106_n452.t28 diffpairibias.t19 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X163 CSoutput.t46 a_n6972_8799.t79 vdd.t91 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X164 CSoutput.t106 commonsourceibias.t69 gnd.t98 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 a_n6972_8799.t0 plus.t17 a_n3106_n452.t15 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X166 CSoutput.t105 commonsourceibias.t70 gnd.t14 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X167 a_n3106_n452.t32 diffpairibias.t20 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X168 vdd.t90 a_n6972_8799.t80 CSoutput.t137 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X169 gnd.t6 commonsourceibias.t71 CSoutput.t104 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X170 CSoutput.t103 commonsourceibias.t72 gnd.t62 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 a_n6972_8799.t27 plus.t18 a_n3106_n452.t14 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X172 vdd.t89 a_n6972_8799.t81 CSoutput.t27 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 minus.t3 gnd.t186 gnd.t188 gnd.t187 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X174 gnd.t185 gnd.t183 gnd.t184 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X175 diffpairibias.t9 diffpairibias.t8 gnd.t271 gnd.t270 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X176 a_n2848_n452.t12 minus.t15 a_n3106_n452.t44 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X177 CSoutput.t35 a_n6972_8799.t82 vdd.t88 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X178 a_n3106_n452.t13 plus.t19 a_n6972_8799.t24 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X179 CSoutput.t142 a_n6972_8799.t83 vdd.t86 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X180 CSoutput.t102 commonsourceibias.t73 gnd.t236 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X181 gnd.t56 commonsourceibias.t74 CSoutput.t101 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 vdd.t214 vdd.t212 vdd.t213 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X183 a_n1808_13878.t17 a_n2848_n452.t60 vdd.t257 vdd.t256 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X184 vdd.t259 a_n2848_n452.t61 a_n1808_13878.t16 vdd.t258 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X185 gnd.t88 commonsourceibias.t22 commonsourceibias.t23 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 gnd.t241 commonsourceibias.t75 CSoutput.t100 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X187 output.t13 CSoutput.t154 vdd.t167 gnd.t27 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X188 CSoutput.t59 a_n6972_8799.t84 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 vdd.t83 a_n6972_8799.t85 CSoutput.t36 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 gnd.t8 commonsourceibias.t76 CSoutput.t99 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 a_n3106_n452.t2 minus.t16 a_n2848_n452.t1 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X192 diffpairibias.t7 diffpairibias.t6 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X193 CSoutput.t37 a_n6972_8799.t86 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X194 gnd.t46 commonsourceibias.t20 commonsourceibias.t21 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 output.t12 CSoutput.t155 vdd.t168 gnd.t28 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X196 vdd.t79 a_n6972_8799.t87 CSoutput.t41 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X197 CSoutput.t98 commonsourceibias.t77 gnd.t111 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 a_n3106_n452.t42 minus.t17 a_n2848_n452.t11 gnd.t232 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X199 a_n3106_n452.t12 plus.t20 a_n6972_8799.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X200 gnd.t182 gnd.t180 gnd.t181 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X201 gnd.t179 gnd.t177 gnd.t178 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X202 a_n1986_8322.t6 a_n2848_n452.t62 a_n6972_8799.t18 vdd.t142 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X203 CSoutput.t17 a_n6972_8799.t88 vdd.t78 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X204 CSoutput.t97 commonsourceibias.t78 gnd.t24 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X205 a_n3106_n452.t1 minus.t18 a_n2848_n452.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X206 vdd.t77 a_n6972_8799.t89 CSoutput.t43 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 vdd.t75 a_n6972_8799.t90 CSoutput.t8 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 CSoutput.t55 a_n6972_8799.t91 vdd.t73 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X209 vdd.t72 a_n6972_8799.t92 CSoutput.t11 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X210 vdd.t158 a_n2848_n452.t63 a_n1986_8322.t14 vdd.t157 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X211 gnd.t33 commonsourceibias.t18 commonsourceibias.t19 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 a_n1808_13878.t15 a_n2848_n452.t64 vdd.t8 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X213 gnd.t176 gnd.t173 gnd.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X214 minus.t2 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X215 CSoutput.t96 commonsourceibias.t79 gnd.t75 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X216 a_n3106_n452.t41 diffpairibias.t21 gnd.t245 gnd.t244 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X217 vdd.t71 a_n6972_8799.t93 CSoutput.t70 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X218 CSoutput.t73 a_n6972_8799.t94 vdd.t70 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X219 a_n6972_8799.t30 plus.t21 a_n3106_n452.t11 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X220 a_n2848_n452.t4 minus.t19 a_n3106_n452.t30 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X221 CSoutput.t95 commonsourceibias.t80 gnd.t48 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 output.t11 CSoutput.t156 vdd.t166 gnd.t81 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X223 CSoutput.t19 a_n6972_8799.t95 vdd.t69 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X224 a_n3106_n452.t29 minus.t20 a_n2848_n452.t3 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X225 CSoutput.t157 a_n1986_8322.t21 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X226 vdd.t211 vdd.t209 vdd.t210 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X227 CSoutput.t94 commonsourceibias.t81 gnd.t95 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 gnd.t169 gnd.t166 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X229 a_n1986_8322.t5 a_n2848_n452.t65 a_n6972_8799.t4 vdd.t9 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X230 vdd.t208 vdd.t206 vdd.t207 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X231 vdd.t151 a_n2848_n452.t66 a_n1986_8322.t13 vdd.t150 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 vdd.t68 a_n6972_8799.t96 CSoutput.t38 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 CSoutput.t57 a_n6972_8799.t97 vdd.t67 vdd.t66 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 gnd.t91 commonsourceibias.t82 CSoutput.t93 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 output.t2 outputibias.t9 gnd.t18 gnd.t17 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X236 CSoutput.t140 a_n6972_8799.t98 vdd.t65 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 a_n3106_n452.t36 minus.t21 a_n2848_n452.t8 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X238 gnd.t165 gnd.t163 gnd.t164 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X239 vdd.t165 CSoutput.t158 output.t10 gnd.t82 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X240 vdd.t64 a_n6972_8799.t99 CSoutput.t53 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X241 vdd.t63 a_n6972_8799.t100 CSoutput.t72 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 a_n3106_n452.t38 minus.t22 a_n2848_n452.t10 gnd.t110 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X243 gnd.t162 gnd.t160 gnd.t161 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X244 output.t1 outputibias.t10 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X245 diffpairibias.t5 diffpairibias.t4 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X246 vdd.t205 vdd.t202 vdd.t204 vdd.t203 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X247 CSoutput.t9 a_n6972_8799.t101 vdd.t62 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 a_n1808_13878.t2 a_n2848_n452.t37 a_n2848_n452.t38 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X249 gnd.t268 commonsourceibias.t83 CSoutput.t92 gnd.t55 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 CSoutput.t91 commonsourceibias.t84 gnd.t57 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X251 a_n1986_8322.t4 a_n2848_n452.t67 a_n6972_8799.t14 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X252 gnd.t159 gnd.t156 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X253 gnd.t290 commonsourceibias.t85 CSoutput.t90 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X254 gnd.t260 commonsourceibias.t16 commonsourceibias.t17 gnd.t240 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X255 vdd.t61 a_n6972_8799.t102 CSoutput.t1 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 CSoutput.t3 a_n6972_8799.t103 vdd.t60 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 a_n3106_n452.t34 minus.t23 a_n2848_n452.t6 gnd.t80 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X258 gnd.t155 gnd.t152 gnd.t154 gnd.t153 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X259 vdd.t177 CSoutput.t159 output.t9 gnd.t83 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X260 output.t8 CSoutput.t160 vdd.t173 gnd.t84 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X261 vdd.t58 a_n6972_8799.t104 CSoutput.t132 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 CSoutput.t75 a_n6972_8799.t105 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 a_n1986_8322.t12 a_n2848_n452.t68 vdd.t144 vdd.t143 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X264 gnd.t151 gnd.t149 plus.t2 gnd.t150 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X265 gnd.t148 gnd.t146 gnd.t147 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X266 CSoutput.t89 commonsourceibias.t86 gnd.t52 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X267 gnd.t145 gnd.t142 gnd.t144 gnd.t143 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X268 CSoutput.t88 commonsourceibias.t87 gnd.t112 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X269 gnd.t141 gnd.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X270 output.t7 CSoutput.t161 vdd.t171 gnd.t85 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X271 vdd.t146 a_n2848_n452.t69 a_n1808_13878.t14 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X272 vdd.t201 vdd.t199 vdd.t200 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X273 CSoutput.t31 a_n6972_8799.t106 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X274 CSoutput.t21 a_n6972_8799.t107 vdd.t52 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 vdd.t51 a_n6972_8799.t108 CSoutput.t6 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 vdd.t49 a_n6972_8799.t109 CSoutput.t7 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X277 vdd.t198 vdd.t195 vdd.t197 vdd.t196 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X278 a_n1986_8322.t3 a_n2848_n452.t70 a_n6972_8799.t7 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X279 a_n3106_n452.t10 plus.t22 a_n6972_8799.t28 gnd.t234 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X280 output.t0 outputibias.t11 gnd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X281 vdd.t194 vdd.t192 vdd.t193 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X282 a_n6972_8799.t8 a_n2848_n452.t71 a_n1986_8322.t2 vdd.t139 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X283 a_n1808_13878.t13 a_n2848_n452.t72 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X284 vdd.t48 a_n6972_8799.t110 CSoutput.t14 vdd.t47 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 CSoutput.t33 a_n6972_8799.t111 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 gnd.t137 gnd.t135 minus.t1 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X287 a_n2848_n452.t5 minus.t24 a_n3106_n452.t33 gnd.t74 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X288 a_n6972_8799.t29 plus.t23 a_n3106_n452.t9 gnd.t254 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X289 CSoutput.t87 commonsourceibias.t88 gnd.t42 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X290 vdd.t44 a_n6972_8799.t112 CSoutput.t47 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 a_n2848_n452.t7 minus.t25 a_n3106_n452.t35 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X292 CSoutput.t15 a_n6972_8799.t113 vdd.t43 vdd.t42 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 commonsourceibias.t15 commonsourceibias.t14 gnd.t256 gnd.t61 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 gnd.t72 commonsourceibias.t89 CSoutput.t86 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 vdd.t179 CSoutput.t162 output.t6 gnd.t250 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X296 vdd.t191 vdd.t188 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X297 vdd.t187 vdd.t184 vdd.t186 vdd.t185 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X298 gnd.t113 commonsourceibias.t90 CSoutput.t85 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 CSoutput.t139 a_n6972_8799.t114 vdd.t41 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X300 vdd.t40 a_n6972_8799.t115 CSoutput.t61 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X301 a_n1808_13878.t1 a_n2848_n452.t31 a_n2848_n452.t32 vdd.t149 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X302 gnd.t134 gnd.t131 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X303 a_n3106_n452.t55 minus.t26 a_n2848_n452.t47 gnd.t286 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X304 a_n3106_n452.t40 diffpairibias.t22 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X305 gnd.t45 commonsourceibias.t91 CSoutput.t84 gnd.t44 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X306 commonsourceibias.t13 commonsourceibias.t12 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X307 a_n6972_8799.t10 plus.t24 a_n3106_n452.t8 gnd.t47 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X308 CSoutput.t52 a_n6972_8799.t116 vdd.t39 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X309 vdd.t38 a_n6972_8799.t117 CSoutput.t5 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X310 diffpairibias.t3 diffpairibias.t2 gnd.t109 gnd.t108 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X311 a_n6972_8799.t21 a_n2848_n452.t73 a_n1986_8322.t1 vdd.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X312 a_n2848_n452.t30 a_n2848_n452.t29 a_n1808_13878.t0 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X313 vdd.t37 a_n6972_8799.t118 CSoutput.t64 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X314 gnd.t130 gnd.t128 plus.t1 gnd.t129 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X315 a_n2848_n452.t2 minus.t27 a_n3106_n452.t3 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X316 vdd.t36 a_n6972_8799.t119 CSoutput.t68 vdd.t35 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X317 CSoutput.t65 a_n6972_8799.t120 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X318 commonsourceibias.t11 commonsourceibias.t10 gnd.t69 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 gnd.t77 commonsourceibias.t92 CSoutput.t83 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X320 vdd.t183 vdd.t180 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X321 vdd.t32 a_n6972_8799.t121 CSoutput.t12 vdd.t31 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X322 CSoutput.t163 a_n1986_8322.t20 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X323 diffpairibias.t1 diffpairibias.t0 gnd.t231 gnd.t230 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X324 CSoutput.t66 a_n6972_8799.t122 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 CSoutput.t82 commonsourceibias.t93 gnd.t223 gnd.t9 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X327 vdd.t28 a_n6972_8799.t123 CSoutput.t25 vdd.t27 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X328 output.t5 CSoutput.t164 vdd.t169 gnd.t251 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X329 plus.t0 gnd.t121 gnd.t123 gnd.t122 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X330 gnd.t120 gnd.t117 gnd.t119 gnd.t118 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X331 CSoutput.t81 commonsourceibias.t94 gnd.t280 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 commonsourceibias.t9 commonsourceibias.t8 gnd.t259 gnd.t58 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 gnd.t116 gnd.t114 minus.t0 gnd.t115 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X334 a_n6972_8799.t6 plus.t25 a_n3106_n452.t7 gnd.t35 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X335 vdd.t5 a_n2848_n452.t74 a_n1808_13878.t12 vdd.t4 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X336 CSoutput.t136 a_n6972_8799.t124 vdd.t26 vdd.t25 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 CSoutput.t80 commonsourceibias.t95 gnd.t60 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X338 a_n6972_8799.t25 plus.t26 a_n3106_n452.t6 gnd.t226 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X339 a_n2848_n452.t9 minus.t28 a_n3106_n452.t37 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X340 output.t4 CSoutput.t165 vdd.t174 gnd.t249 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X341 vdd.t24 a_n6972_8799.t125 CSoutput.t60 vdd.t23 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X342 CSoutput.t16 a_n6972_8799.t126 vdd.t22 vdd.t21 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X343 vdd.t20 a_n6972_8799.t127 CSoutput.t62 vdd.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X344 gnd.t71 commonsourceibias.t6 commonsourceibias.t7 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X345 commonsourceibias.t5 commonsourceibias.t4 gnd.t272 gnd.t13 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 CSoutput.t48 a_n6972_8799.t128 vdd.t18 vdd.t17 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 vdd.t16 a_n6972_8799.t129 CSoutput.t18 vdd.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 a_n1986_8322.t0 a_n2848_n452.t75 a_n6972_8799.t3 vdd.t6 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X349 a_n3106_n452.t5 plus.t27 a_n6972_8799.t34 gnd.t31 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X350 commonsourceibias.t3 commonsourceibias.t2 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X351 vdd.t14 a_n6972_8799.t130 CSoutput.t26 vdd.t13 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X352 CSoutput.t13 a_n6972_8799.t131 vdd.t12 vdd.t11 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X353 a_n3106_n452.t4 plus.t28 a_n6972_8799.t19 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X354 gnd.t258 commonsourceibias.t0 commonsourceibias.t1 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X355 a_n3106_n452.t39 diffpairibias.t23 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 gnd.n6510 gnd.n404 1655.14
R1 gnd.n5914 gnd.n4574 939.716
R2 gnd.n6800 gnd.n84 838.452
R3 gnd.n6963 gnd.n80 838.452
R4 gnd.n1363 gnd.n1310 838.452
R5 gnd.n4152 gnd.n1365 838.452
R6 gnd.n4368 gnd.n1163 838.452
R7 gnd.n2864 gnd.n1161 838.452
R8 gnd.n2356 gnd.n905 838.452
R9 gnd.n2418 gnd.n2357 838.452
R10 gnd.n6961 gnd.n86 819.232
R11 gnd.n155 gnd.n82 819.232
R12 gnd.n4155 gnd.n4154 819.232
R13 gnd.n4227 gnd.n1314 819.232
R14 gnd.n4370 gnd.n1158 819.232
R15 gnd.n2178 gnd.n1160 819.232
R16 gnd.n4496 gnd.n4495 819.232
R17 gnd.n4572 gnd.n909 819.232
R18 gnd.n2057 gnd.n1168 771.183
R19 gnd.n4239 gnd.n1271 771.183
R20 gnd.n2909 gnd.n1977 771.183
R21 gnd.n3893 gnd.n1274 771.183
R22 gnd.n864 gnd.n850 766.379
R23 gnd.n5830 gnd.n5829 766.379
R24 gnd.n5045 gnd.n4944 766.379
R25 gnd.n5043 gnd.n4946 766.379
R26 gnd.n5915 gnd.n855 756.769
R27 gnd.n5816 gnd.n5815 756.769
R28 gnd.n5177 gnd.n4906 756.769
R29 gnd.n5163 gnd.n4895 756.769
R30 gnd.n6118 gnd.n636 723.135
R31 gnd.n6509 gnd.n405 723.135
R32 gnd.n6722 gnd.n6721 723.135
R33 gnd.n2315 gnd.n2309 723.135
R34 gnd.n6118 gnd.n6117 585
R35 gnd.n6119 gnd.n6118 585
R36 gnd.n6116 gnd.n638 585
R37 gnd.n638 gnd.n637 585
R38 gnd.n6115 gnd.n6114 585
R39 gnd.n6114 gnd.n6113 585
R40 gnd.n643 gnd.n642 585
R41 gnd.n6112 gnd.n643 585
R42 gnd.n6110 gnd.n6109 585
R43 gnd.n6111 gnd.n6110 585
R44 gnd.n6108 gnd.n645 585
R45 gnd.n645 gnd.n644 585
R46 gnd.n6107 gnd.n6106 585
R47 gnd.n6106 gnd.n6105 585
R48 gnd.n651 gnd.n650 585
R49 gnd.n6104 gnd.n651 585
R50 gnd.n6102 gnd.n6101 585
R51 gnd.n6103 gnd.n6102 585
R52 gnd.n6100 gnd.n653 585
R53 gnd.n653 gnd.n652 585
R54 gnd.n6099 gnd.n6098 585
R55 gnd.n6098 gnd.n6097 585
R56 gnd.n659 gnd.n658 585
R57 gnd.n6096 gnd.n659 585
R58 gnd.n6094 gnd.n6093 585
R59 gnd.n6095 gnd.n6094 585
R60 gnd.n6092 gnd.n661 585
R61 gnd.n661 gnd.n660 585
R62 gnd.n6091 gnd.n6090 585
R63 gnd.n6090 gnd.n6089 585
R64 gnd.n667 gnd.n666 585
R65 gnd.n6088 gnd.n667 585
R66 gnd.n6086 gnd.n6085 585
R67 gnd.n6087 gnd.n6086 585
R68 gnd.n6084 gnd.n669 585
R69 gnd.n669 gnd.n668 585
R70 gnd.n6083 gnd.n6082 585
R71 gnd.n6082 gnd.n6081 585
R72 gnd.n675 gnd.n674 585
R73 gnd.n6080 gnd.n675 585
R74 gnd.n6078 gnd.n6077 585
R75 gnd.n6079 gnd.n6078 585
R76 gnd.n6076 gnd.n677 585
R77 gnd.n677 gnd.n676 585
R78 gnd.n6075 gnd.n6074 585
R79 gnd.n6074 gnd.n6073 585
R80 gnd.n683 gnd.n682 585
R81 gnd.n6072 gnd.n683 585
R82 gnd.n6070 gnd.n6069 585
R83 gnd.n6071 gnd.n6070 585
R84 gnd.n6068 gnd.n685 585
R85 gnd.n685 gnd.n684 585
R86 gnd.n6067 gnd.n6066 585
R87 gnd.n6066 gnd.n6065 585
R88 gnd.n691 gnd.n690 585
R89 gnd.n6064 gnd.n691 585
R90 gnd.n6062 gnd.n6061 585
R91 gnd.n6063 gnd.n6062 585
R92 gnd.n6060 gnd.n693 585
R93 gnd.n693 gnd.n692 585
R94 gnd.n6059 gnd.n6058 585
R95 gnd.n6058 gnd.n6057 585
R96 gnd.n699 gnd.n698 585
R97 gnd.n6056 gnd.n699 585
R98 gnd.n6054 gnd.n6053 585
R99 gnd.n6055 gnd.n6054 585
R100 gnd.n6052 gnd.n701 585
R101 gnd.n701 gnd.n700 585
R102 gnd.n6051 gnd.n6050 585
R103 gnd.n6050 gnd.n6049 585
R104 gnd.n707 gnd.n706 585
R105 gnd.n6048 gnd.n707 585
R106 gnd.n6046 gnd.n6045 585
R107 gnd.n6047 gnd.n6046 585
R108 gnd.n6044 gnd.n709 585
R109 gnd.n709 gnd.n708 585
R110 gnd.n6043 gnd.n6042 585
R111 gnd.n6042 gnd.n6041 585
R112 gnd.n715 gnd.n714 585
R113 gnd.n6040 gnd.n715 585
R114 gnd.n6038 gnd.n6037 585
R115 gnd.n6039 gnd.n6038 585
R116 gnd.n6036 gnd.n717 585
R117 gnd.n717 gnd.n716 585
R118 gnd.n6035 gnd.n6034 585
R119 gnd.n6034 gnd.n6033 585
R120 gnd.n723 gnd.n722 585
R121 gnd.n6032 gnd.n723 585
R122 gnd.n6030 gnd.n6029 585
R123 gnd.n6031 gnd.n6030 585
R124 gnd.n6028 gnd.n725 585
R125 gnd.n725 gnd.n724 585
R126 gnd.n6027 gnd.n6026 585
R127 gnd.n6026 gnd.n6025 585
R128 gnd.n731 gnd.n730 585
R129 gnd.n6024 gnd.n731 585
R130 gnd.n6022 gnd.n6021 585
R131 gnd.n6023 gnd.n6022 585
R132 gnd.n6020 gnd.n733 585
R133 gnd.n733 gnd.n732 585
R134 gnd.n6019 gnd.n6018 585
R135 gnd.n6018 gnd.n6017 585
R136 gnd.n739 gnd.n738 585
R137 gnd.n6016 gnd.n739 585
R138 gnd.n6014 gnd.n6013 585
R139 gnd.n6015 gnd.n6014 585
R140 gnd.n6012 gnd.n741 585
R141 gnd.n741 gnd.n740 585
R142 gnd.n6011 gnd.n6010 585
R143 gnd.n6010 gnd.n6009 585
R144 gnd.n747 gnd.n746 585
R145 gnd.n6008 gnd.n747 585
R146 gnd.n6006 gnd.n6005 585
R147 gnd.n6007 gnd.n6006 585
R148 gnd.n6004 gnd.n749 585
R149 gnd.n749 gnd.n748 585
R150 gnd.n6003 gnd.n6002 585
R151 gnd.n6002 gnd.n6001 585
R152 gnd.n755 gnd.n754 585
R153 gnd.n6000 gnd.n755 585
R154 gnd.n5998 gnd.n5997 585
R155 gnd.n5999 gnd.n5998 585
R156 gnd.n5996 gnd.n757 585
R157 gnd.n757 gnd.n756 585
R158 gnd.n5995 gnd.n5994 585
R159 gnd.n5994 gnd.n5993 585
R160 gnd.n763 gnd.n762 585
R161 gnd.n5992 gnd.n763 585
R162 gnd.n5990 gnd.n5989 585
R163 gnd.n5991 gnd.n5990 585
R164 gnd.n5988 gnd.n765 585
R165 gnd.n765 gnd.n764 585
R166 gnd.n5987 gnd.n5986 585
R167 gnd.n5986 gnd.n5985 585
R168 gnd.n771 gnd.n770 585
R169 gnd.n5984 gnd.n771 585
R170 gnd.n5982 gnd.n5981 585
R171 gnd.n5983 gnd.n5982 585
R172 gnd.n5980 gnd.n773 585
R173 gnd.n773 gnd.n772 585
R174 gnd.n5979 gnd.n5978 585
R175 gnd.n5978 gnd.n5977 585
R176 gnd.n779 gnd.n778 585
R177 gnd.n5976 gnd.n779 585
R178 gnd.n5974 gnd.n5973 585
R179 gnd.n5975 gnd.n5974 585
R180 gnd.n5972 gnd.n781 585
R181 gnd.n781 gnd.n780 585
R182 gnd.n5971 gnd.n5970 585
R183 gnd.n5970 gnd.n5969 585
R184 gnd.n787 gnd.n786 585
R185 gnd.n5968 gnd.n787 585
R186 gnd.n5966 gnd.n5965 585
R187 gnd.n5967 gnd.n5966 585
R188 gnd.n5964 gnd.n789 585
R189 gnd.n789 gnd.n788 585
R190 gnd.n5963 gnd.n5962 585
R191 gnd.n5962 gnd.n5961 585
R192 gnd.n795 gnd.n794 585
R193 gnd.n5960 gnd.n795 585
R194 gnd.n5958 gnd.n5957 585
R195 gnd.n5959 gnd.n5958 585
R196 gnd.n5956 gnd.n797 585
R197 gnd.n797 gnd.n796 585
R198 gnd.n5955 gnd.n5954 585
R199 gnd.n5954 gnd.n5953 585
R200 gnd.n803 gnd.n802 585
R201 gnd.n5952 gnd.n803 585
R202 gnd.n636 gnd.n635 585
R203 gnd.n6120 gnd.n636 585
R204 gnd.n6123 gnd.n6122 585
R205 gnd.n6122 gnd.n6121 585
R206 gnd.n633 gnd.n632 585
R207 gnd.n632 gnd.n631 585
R208 gnd.n6128 gnd.n6127 585
R209 gnd.n6129 gnd.n6128 585
R210 gnd.n630 gnd.n629 585
R211 gnd.n6130 gnd.n630 585
R212 gnd.n6133 gnd.n6132 585
R213 gnd.n6132 gnd.n6131 585
R214 gnd.n627 gnd.n626 585
R215 gnd.n626 gnd.n625 585
R216 gnd.n6138 gnd.n6137 585
R217 gnd.n6139 gnd.n6138 585
R218 gnd.n624 gnd.n623 585
R219 gnd.n6140 gnd.n624 585
R220 gnd.n6143 gnd.n6142 585
R221 gnd.n6142 gnd.n6141 585
R222 gnd.n621 gnd.n620 585
R223 gnd.n620 gnd.n619 585
R224 gnd.n6148 gnd.n6147 585
R225 gnd.n6149 gnd.n6148 585
R226 gnd.n618 gnd.n617 585
R227 gnd.n6150 gnd.n618 585
R228 gnd.n6153 gnd.n6152 585
R229 gnd.n6152 gnd.n6151 585
R230 gnd.n615 gnd.n614 585
R231 gnd.n614 gnd.n613 585
R232 gnd.n6158 gnd.n6157 585
R233 gnd.n6159 gnd.n6158 585
R234 gnd.n612 gnd.n611 585
R235 gnd.n6160 gnd.n612 585
R236 gnd.n6163 gnd.n6162 585
R237 gnd.n6162 gnd.n6161 585
R238 gnd.n609 gnd.n608 585
R239 gnd.n608 gnd.n607 585
R240 gnd.n6168 gnd.n6167 585
R241 gnd.n6169 gnd.n6168 585
R242 gnd.n606 gnd.n605 585
R243 gnd.n6170 gnd.n606 585
R244 gnd.n6173 gnd.n6172 585
R245 gnd.n6172 gnd.n6171 585
R246 gnd.n603 gnd.n602 585
R247 gnd.n602 gnd.n601 585
R248 gnd.n6178 gnd.n6177 585
R249 gnd.n6179 gnd.n6178 585
R250 gnd.n600 gnd.n599 585
R251 gnd.n6180 gnd.n600 585
R252 gnd.n6183 gnd.n6182 585
R253 gnd.n6182 gnd.n6181 585
R254 gnd.n597 gnd.n596 585
R255 gnd.n596 gnd.n595 585
R256 gnd.n6188 gnd.n6187 585
R257 gnd.n6189 gnd.n6188 585
R258 gnd.n594 gnd.n593 585
R259 gnd.n6190 gnd.n594 585
R260 gnd.n6193 gnd.n6192 585
R261 gnd.n6192 gnd.n6191 585
R262 gnd.n591 gnd.n590 585
R263 gnd.n590 gnd.n589 585
R264 gnd.n6198 gnd.n6197 585
R265 gnd.n6199 gnd.n6198 585
R266 gnd.n588 gnd.n587 585
R267 gnd.n6200 gnd.n588 585
R268 gnd.n6203 gnd.n6202 585
R269 gnd.n6202 gnd.n6201 585
R270 gnd.n585 gnd.n584 585
R271 gnd.n584 gnd.n583 585
R272 gnd.n6208 gnd.n6207 585
R273 gnd.n6209 gnd.n6208 585
R274 gnd.n582 gnd.n581 585
R275 gnd.n6210 gnd.n582 585
R276 gnd.n6213 gnd.n6212 585
R277 gnd.n6212 gnd.n6211 585
R278 gnd.n579 gnd.n578 585
R279 gnd.n578 gnd.n577 585
R280 gnd.n6218 gnd.n6217 585
R281 gnd.n6219 gnd.n6218 585
R282 gnd.n576 gnd.n575 585
R283 gnd.n6220 gnd.n576 585
R284 gnd.n6223 gnd.n6222 585
R285 gnd.n6222 gnd.n6221 585
R286 gnd.n573 gnd.n572 585
R287 gnd.n572 gnd.n571 585
R288 gnd.n6228 gnd.n6227 585
R289 gnd.n6229 gnd.n6228 585
R290 gnd.n570 gnd.n569 585
R291 gnd.n6230 gnd.n570 585
R292 gnd.n6233 gnd.n6232 585
R293 gnd.n6232 gnd.n6231 585
R294 gnd.n567 gnd.n566 585
R295 gnd.n566 gnd.n565 585
R296 gnd.n6238 gnd.n6237 585
R297 gnd.n6239 gnd.n6238 585
R298 gnd.n564 gnd.n563 585
R299 gnd.n6240 gnd.n564 585
R300 gnd.n6243 gnd.n6242 585
R301 gnd.n6242 gnd.n6241 585
R302 gnd.n561 gnd.n560 585
R303 gnd.n560 gnd.n559 585
R304 gnd.n6248 gnd.n6247 585
R305 gnd.n6249 gnd.n6248 585
R306 gnd.n558 gnd.n557 585
R307 gnd.n6250 gnd.n558 585
R308 gnd.n6253 gnd.n6252 585
R309 gnd.n6252 gnd.n6251 585
R310 gnd.n555 gnd.n554 585
R311 gnd.n554 gnd.n553 585
R312 gnd.n6258 gnd.n6257 585
R313 gnd.n6259 gnd.n6258 585
R314 gnd.n552 gnd.n551 585
R315 gnd.n6260 gnd.n552 585
R316 gnd.n6263 gnd.n6262 585
R317 gnd.n6262 gnd.n6261 585
R318 gnd.n549 gnd.n548 585
R319 gnd.n548 gnd.n547 585
R320 gnd.n6268 gnd.n6267 585
R321 gnd.n6269 gnd.n6268 585
R322 gnd.n546 gnd.n545 585
R323 gnd.n6270 gnd.n546 585
R324 gnd.n6273 gnd.n6272 585
R325 gnd.n6272 gnd.n6271 585
R326 gnd.n543 gnd.n542 585
R327 gnd.n542 gnd.n541 585
R328 gnd.n6278 gnd.n6277 585
R329 gnd.n6279 gnd.n6278 585
R330 gnd.n540 gnd.n539 585
R331 gnd.n6280 gnd.n540 585
R332 gnd.n6283 gnd.n6282 585
R333 gnd.n6282 gnd.n6281 585
R334 gnd.n537 gnd.n536 585
R335 gnd.n536 gnd.n535 585
R336 gnd.n6288 gnd.n6287 585
R337 gnd.n6289 gnd.n6288 585
R338 gnd.n534 gnd.n533 585
R339 gnd.n6290 gnd.n534 585
R340 gnd.n6293 gnd.n6292 585
R341 gnd.n6292 gnd.n6291 585
R342 gnd.n531 gnd.n530 585
R343 gnd.n530 gnd.n529 585
R344 gnd.n6298 gnd.n6297 585
R345 gnd.n6299 gnd.n6298 585
R346 gnd.n528 gnd.n527 585
R347 gnd.n6300 gnd.n528 585
R348 gnd.n6303 gnd.n6302 585
R349 gnd.n6302 gnd.n6301 585
R350 gnd.n525 gnd.n524 585
R351 gnd.n524 gnd.n523 585
R352 gnd.n6308 gnd.n6307 585
R353 gnd.n6309 gnd.n6308 585
R354 gnd.n522 gnd.n521 585
R355 gnd.n6310 gnd.n522 585
R356 gnd.n6313 gnd.n6312 585
R357 gnd.n6312 gnd.n6311 585
R358 gnd.n519 gnd.n518 585
R359 gnd.n518 gnd.n517 585
R360 gnd.n6318 gnd.n6317 585
R361 gnd.n6319 gnd.n6318 585
R362 gnd.n516 gnd.n515 585
R363 gnd.n6320 gnd.n516 585
R364 gnd.n6323 gnd.n6322 585
R365 gnd.n6322 gnd.n6321 585
R366 gnd.n513 gnd.n512 585
R367 gnd.n512 gnd.n511 585
R368 gnd.n6328 gnd.n6327 585
R369 gnd.n6329 gnd.n6328 585
R370 gnd.n510 gnd.n509 585
R371 gnd.n6330 gnd.n510 585
R372 gnd.n6333 gnd.n6332 585
R373 gnd.n6332 gnd.n6331 585
R374 gnd.n507 gnd.n506 585
R375 gnd.n506 gnd.n505 585
R376 gnd.n6338 gnd.n6337 585
R377 gnd.n6339 gnd.n6338 585
R378 gnd.n504 gnd.n503 585
R379 gnd.n6340 gnd.n504 585
R380 gnd.n6343 gnd.n6342 585
R381 gnd.n6342 gnd.n6341 585
R382 gnd.n501 gnd.n500 585
R383 gnd.n500 gnd.n499 585
R384 gnd.n6348 gnd.n6347 585
R385 gnd.n6349 gnd.n6348 585
R386 gnd.n498 gnd.n497 585
R387 gnd.n6350 gnd.n498 585
R388 gnd.n6353 gnd.n6352 585
R389 gnd.n6352 gnd.n6351 585
R390 gnd.n495 gnd.n494 585
R391 gnd.n494 gnd.n493 585
R392 gnd.n6358 gnd.n6357 585
R393 gnd.n6359 gnd.n6358 585
R394 gnd.n492 gnd.n491 585
R395 gnd.n6360 gnd.n492 585
R396 gnd.n6363 gnd.n6362 585
R397 gnd.n6362 gnd.n6361 585
R398 gnd.n489 gnd.n488 585
R399 gnd.n488 gnd.n487 585
R400 gnd.n6368 gnd.n6367 585
R401 gnd.n6369 gnd.n6368 585
R402 gnd.n486 gnd.n485 585
R403 gnd.n6370 gnd.n486 585
R404 gnd.n6373 gnd.n6372 585
R405 gnd.n6372 gnd.n6371 585
R406 gnd.n483 gnd.n482 585
R407 gnd.n482 gnd.n481 585
R408 gnd.n6378 gnd.n6377 585
R409 gnd.n6379 gnd.n6378 585
R410 gnd.n480 gnd.n479 585
R411 gnd.n6380 gnd.n480 585
R412 gnd.n6383 gnd.n6382 585
R413 gnd.n6382 gnd.n6381 585
R414 gnd.n477 gnd.n476 585
R415 gnd.n476 gnd.n475 585
R416 gnd.n6388 gnd.n6387 585
R417 gnd.n6389 gnd.n6388 585
R418 gnd.n474 gnd.n473 585
R419 gnd.n6390 gnd.n474 585
R420 gnd.n6393 gnd.n6392 585
R421 gnd.n6392 gnd.n6391 585
R422 gnd.n471 gnd.n470 585
R423 gnd.n470 gnd.n469 585
R424 gnd.n6398 gnd.n6397 585
R425 gnd.n6399 gnd.n6398 585
R426 gnd.n468 gnd.n467 585
R427 gnd.n6400 gnd.n468 585
R428 gnd.n6403 gnd.n6402 585
R429 gnd.n6402 gnd.n6401 585
R430 gnd.n465 gnd.n464 585
R431 gnd.n464 gnd.n463 585
R432 gnd.n6408 gnd.n6407 585
R433 gnd.n6409 gnd.n6408 585
R434 gnd.n462 gnd.n461 585
R435 gnd.n6410 gnd.n462 585
R436 gnd.n6413 gnd.n6412 585
R437 gnd.n6412 gnd.n6411 585
R438 gnd.n459 gnd.n458 585
R439 gnd.n458 gnd.n457 585
R440 gnd.n6418 gnd.n6417 585
R441 gnd.n6419 gnd.n6418 585
R442 gnd.n456 gnd.n455 585
R443 gnd.n6420 gnd.n456 585
R444 gnd.n6423 gnd.n6422 585
R445 gnd.n6422 gnd.n6421 585
R446 gnd.n453 gnd.n452 585
R447 gnd.n452 gnd.n451 585
R448 gnd.n6428 gnd.n6427 585
R449 gnd.n6429 gnd.n6428 585
R450 gnd.n450 gnd.n449 585
R451 gnd.n6430 gnd.n450 585
R452 gnd.n6433 gnd.n6432 585
R453 gnd.n6432 gnd.n6431 585
R454 gnd.n447 gnd.n446 585
R455 gnd.n446 gnd.n445 585
R456 gnd.n6438 gnd.n6437 585
R457 gnd.n6439 gnd.n6438 585
R458 gnd.n444 gnd.n443 585
R459 gnd.n6440 gnd.n444 585
R460 gnd.n6443 gnd.n6442 585
R461 gnd.n6442 gnd.n6441 585
R462 gnd.n441 gnd.n440 585
R463 gnd.n440 gnd.n439 585
R464 gnd.n6448 gnd.n6447 585
R465 gnd.n6449 gnd.n6448 585
R466 gnd.n438 gnd.n437 585
R467 gnd.n6450 gnd.n438 585
R468 gnd.n6453 gnd.n6452 585
R469 gnd.n6452 gnd.n6451 585
R470 gnd.n435 gnd.n434 585
R471 gnd.n434 gnd.n433 585
R472 gnd.n6458 gnd.n6457 585
R473 gnd.n6459 gnd.n6458 585
R474 gnd.n432 gnd.n431 585
R475 gnd.n6460 gnd.n432 585
R476 gnd.n6463 gnd.n6462 585
R477 gnd.n6462 gnd.n6461 585
R478 gnd.n429 gnd.n428 585
R479 gnd.n428 gnd.n427 585
R480 gnd.n6468 gnd.n6467 585
R481 gnd.n6469 gnd.n6468 585
R482 gnd.n426 gnd.n425 585
R483 gnd.n6470 gnd.n426 585
R484 gnd.n6473 gnd.n6472 585
R485 gnd.n6472 gnd.n6471 585
R486 gnd.n423 gnd.n422 585
R487 gnd.n422 gnd.n421 585
R488 gnd.n6478 gnd.n6477 585
R489 gnd.n6479 gnd.n6478 585
R490 gnd.n420 gnd.n419 585
R491 gnd.n6480 gnd.n420 585
R492 gnd.n6483 gnd.n6482 585
R493 gnd.n6482 gnd.n6481 585
R494 gnd.n417 gnd.n416 585
R495 gnd.n416 gnd.n415 585
R496 gnd.n6488 gnd.n6487 585
R497 gnd.n6489 gnd.n6488 585
R498 gnd.n414 gnd.n413 585
R499 gnd.n6490 gnd.n414 585
R500 gnd.n6493 gnd.n6492 585
R501 gnd.n6492 gnd.n6491 585
R502 gnd.n411 gnd.n410 585
R503 gnd.n410 gnd.n409 585
R504 gnd.n6499 gnd.n6498 585
R505 gnd.n6500 gnd.n6499 585
R506 gnd.n408 gnd.n407 585
R507 gnd.n6501 gnd.n408 585
R508 gnd.n6504 gnd.n6503 585
R509 gnd.n6503 gnd.n6502 585
R510 gnd.n6505 gnd.n405 585
R511 gnd.n405 gnd.n404 585
R512 gnd.n280 gnd.n279 585
R513 gnd.n6712 gnd.n279 585
R514 gnd.n6715 gnd.n6714 585
R515 gnd.n6714 gnd.n6713 585
R516 gnd.n283 gnd.n282 585
R517 gnd.n6711 gnd.n283 585
R518 gnd.n6709 gnd.n6708 585
R519 gnd.n6710 gnd.n6709 585
R520 gnd.n286 gnd.n285 585
R521 gnd.n285 gnd.n284 585
R522 gnd.n6704 gnd.n6703 585
R523 gnd.n6703 gnd.n6702 585
R524 gnd.n289 gnd.n288 585
R525 gnd.n6701 gnd.n289 585
R526 gnd.n6699 gnd.n6698 585
R527 gnd.n6700 gnd.n6699 585
R528 gnd.n292 gnd.n291 585
R529 gnd.n291 gnd.n290 585
R530 gnd.n6694 gnd.n6693 585
R531 gnd.n6693 gnd.n6692 585
R532 gnd.n295 gnd.n294 585
R533 gnd.n6691 gnd.n295 585
R534 gnd.n6689 gnd.n6688 585
R535 gnd.n6690 gnd.n6689 585
R536 gnd.n298 gnd.n297 585
R537 gnd.n297 gnd.n296 585
R538 gnd.n6684 gnd.n6683 585
R539 gnd.n6683 gnd.n6682 585
R540 gnd.n301 gnd.n300 585
R541 gnd.n6681 gnd.n301 585
R542 gnd.n6679 gnd.n6678 585
R543 gnd.n6680 gnd.n6679 585
R544 gnd.n304 gnd.n303 585
R545 gnd.n303 gnd.n302 585
R546 gnd.n6674 gnd.n6673 585
R547 gnd.n6673 gnd.n6672 585
R548 gnd.n307 gnd.n306 585
R549 gnd.n6671 gnd.n307 585
R550 gnd.n6669 gnd.n6668 585
R551 gnd.n6670 gnd.n6669 585
R552 gnd.n310 gnd.n309 585
R553 gnd.n309 gnd.n308 585
R554 gnd.n6664 gnd.n6663 585
R555 gnd.n6663 gnd.n6662 585
R556 gnd.n313 gnd.n312 585
R557 gnd.n6661 gnd.n313 585
R558 gnd.n6659 gnd.n6658 585
R559 gnd.n6660 gnd.n6659 585
R560 gnd.n316 gnd.n315 585
R561 gnd.n315 gnd.n314 585
R562 gnd.n6654 gnd.n6653 585
R563 gnd.n6653 gnd.n6652 585
R564 gnd.n319 gnd.n318 585
R565 gnd.n6651 gnd.n319 585
R566 gnd.n6649 gnd.n6648 585
R567 gnd.n6650 gnd.n6649 585
R568 gnd.n322 gnd.n321 585
R569 gnd.n321 gnd.n320 585
R570 gnd.n6644 gnd.n6643 585
R571 gnd.n6643 gnd.n6642 585
R572 gnd.n325 gnd.n324 585
R573 gnd.n6641 gnd.n325 585
R574 gnd.n6639 gnd.n6638 585
R575 gnd.n6640 gnd.n6639 585
R576 gnd.n328 gnd.n327 585
R577 gnd.n327 gnd.n326 585
R578 gnd.n6634 gnd.n6633 585
R579 gnd.n6633 gnd.n6632 585
R580 gnd.n331 gnd.n330 585
R581 gnd.n6631 gnd.n331 585
R582 gnd.n6629 gnd.n6628 585
R583 gnd.n6630 gnd.n6629 585
R584 gnd.n334 gnd.n333 585
R585 gnd.n333 gnd.n332 585
R586 gnd.n6624 gnd.n6623 585
R587 gnd.n6623 gnd.n6622 585
R588 gnd.n337 gnd.n336 585
R589 gnd.n6621 gnd.n337 585
R590 gnd.n6619 gnd.n6618 585
R591 gnd.n6620 gnd.n6619 585
R592 gnd.n340 gnd.n339 585
R593 gnd.n339 gnd.n338 585
R594 gnd.n6614 gnd.n6613 585
R595 gnd.n6613 gnd.n6612 585
R596 gnd.n343 gnd.n342 585
R597 gnd.n6611 gnd.n343 585
R598 gnd.n6609 gnd.n6608 585
R599 gnd.n6610 gnd.n6609 585
R600 gnd.n346 gnd.n345 585
R601 gnd.n345 gnd.n344 585
R602 gnd.n6604 gnd.n6603 585
R603 gnd.n6603 gnd.n6602 585
R604 gnd.n349 gnd.n348 585
R605 gnd.n6601 gnd.n349 585
R606 gnd.n6599 gnd.n6598 585
R607 gnd.n6600 gnd.n6599 585
R608 gnd.n352 gnd.n351 585
R609 gnd.n351 gnd.n350 585
R610 gnd.n6594 gnd.n6593 585
R611 gnd.n6593 gnd.n6592 585
R612 gnd.n355 gnd.n354 585
R613 gnd.n6591 gnd.n355 585
R614 gnd.n6589 gnd.n6588 585
R615 gnd.n6590 gnd.n6589 585
R616 gnd.n358 gnd.n357 585
R617 gnd.n357 gnd.n356 585
R618 gnd.n6584 gnd.n6583 585
R619 gnd.n6583 gnd.n6582 585
R620 gnd.n361 gnd.n360 585
R621 gnd.n6581 gnd.n361 585
R622 gnd.n6579 gnd.n6578 585
R623 gnd.n6580 gnd.n6579 585
R624 gnd.n364 gnd.n363 585
R625 gnd.n363 gnd.n362 585
R626 gnd.n6574 gnd.n6573 585
R627 gnd.n6573 gnd.n6572 585
R628 gnd.n367 gnd.n366 585
R629 gnd.n6571 gnd.n367 585
R630 gnd.n6569 gnd.n6568 585
R631 gnd.n6570 gnd.n6569 585
R632 gnd.n370 gnd.n369 585
R633 gnd.n369 gnd.n368 585
R634 gnd.n6564 gnd.n6563 585
R635 gnd.n6563 gnd.n6562 585
R636 gnd.n373 gnd.n372 585
R637 gnd.n6561 gnd.n373 585
R638 gnd.n6559 gnd.n6558 585
R639 gnd.n6560 gnd.n6559 585
R640 gnd.n376 gnd.n375 585
R641 gnd.n375 gnd.n374 585
R642 gnd.n6554 gnd.n6553 585
R643 gnd.n6553 gnd.n6552 585
R644 gnd.n379 gnd.n378 585
R645 gnd.n6551 gnd.n379 585
R646 gnd.n6549 gnd.n6548 585
R647 gnd.n6550 gnd.n6549 585
R648 gnd.n382 gnd.n381 585
R649 gnd.n381 gnd.n380 585
R650 gnd.n6544 gnd.n6543 585
R651 gnd.n6543 gnd.n6542 585
R652 gnd.n385 gnd.n384 585
R653 gnd.n6541 gnd.n385 585
R654 gnd.n6539 gnd.n6538 585
R655 gnd.n6540 gnd.n6539 585
R656 gnd.n388 gnd.n387 585
R657 gnd.n387 gnd.n386 585
R658 gnd.n6534 gnd.n6533 585
R659 gnd.n6533 gnd.n6532 585
R660 gnd.n391 gnd.n390 585
R661 gnd.n6531 gnd.n391 585
R662 gnd.n6529 gnd.n6528 585
R663 gnd.n6530 gnd.n6529 585
R664 gnd.n394 gnd.n393 585
R665 gnd.n393 gnd.n392 585
R666 gnd.n6524 gnd.n6523 585
R667 gnd.n6523 gnd.n6522 585
R668 gnd.n397 gnd.n396 585
R669 gnd.n6521 gnd.n397 585
R670 gnd.n6519 gnd.n6518 585
R671 gnd.n6520 gnd.n6519 585
R672 gnd.n400 gnd.n399 585
R673 gnd.n399 gnd.n398 585
R674 gnd.n6514 gnd.n6513 585
R675 gnd.n6513 gnd.n6512 585
R676 gnd.n403 gnd.n402 585
R677 gnd.n6511 gnd.n403 585
R678 gnd.n6509 gnd.n6508 585
R679 gnd.n6510 gnd.n6509 585
R680 gnd.n4368 gnd.n4367 585
R681 gnd.n4369 gnd.n4368 585
R682 gnd.n1149 gnd.n1148 585
R683 gnd.n2577 gnd.n1149 585
R684 gnd.n4377 gnd.n4376 585
R685 gnd.n4376 gnd.n4375 585
R686 gnd.n4378 gnd.n1143 585
R687 gnd.n2569 gnd.n1143 585
R688 gnd.n4380 gnd.n4379 585
R689 gnd.n4381 gnd.n4380 585
R690 gnd.n1127 gnd.n1126 585
R691 gnd.n2560 gnd.n1127 585
R692 gnd.n4389 gnd.n4388 585
R693 gnd.n4388 gnd.n4387 585
R694 gnd.n4390 gnd.n1121 585
R695 gnd.n2552 gnd.n1121 585
R696 gnd.n4392 gnd.n4391 585
R697 gnd.n4393 gnd.n4392 585
R698 gnd.n1105 gnd.n1104 585
R699 gnd.n2544 gnd.n1105 585
R700 gnd.n4401 gnd.n4400 585
R701 gnd.n4400 gnd.n4399 585
R702 gnd.n4402 gnd.n1099 585
R703 gnd.n2536 gnd.n1099 585
R704 gnd.n4404 gnd.n4403 585
R705 gnd.n4405 gnd.n4404 585
R706 gnd.n1084 gnd.n1083 585
R707 gnd.n2528 gnd.n1084 585
R708 gnd.n4413 gnd.n4412 585
R709 gnd.n4412 gnd.n4411 585
R710 gnd.n4414 gnd.n1078 585
R711 gnd.n2520 gnd.n1078 585
R712 gnd.n4416 gnd.n4415 585
R713 gnd.n4417 gnd.n4416 585
R714 gnd.n1065 gnd.n1064 585
R715 gnd.n2512 gnd.n1065 585
R716 gnd.n4426 gnd.n4425 585
R717 gnd.n4425 gnd.n4424 585
R718 gnd.n4427 gnd.n1060 585
R719 gnd.n2504 gnd.n1060 585
R720 gnd.n4429 gnd.n4428 585
R721 gnd.n4430 gnd.n4429 585
R722 gnd.n1048 gnd.n1047 585
R723 gnd.n2496 gnd.n1048 585
R724 gnd.n4439 gnd.n4438 585
R725 gnd.n4438 gnd.n4437 585
R726 gnd.n4440 gnd.n1040 585
R727 gnd.n2488 gnd.n1040 585
R728 gnd.n4442 gnd.n4441 585
R729 gnd.n4443 gnd.n4442 585
R730 gnd.n1041 gnd.n1039 585
R731 gnd.n2480 gnd.n1039 585
R732 gnd.n1023 gnd.n1022 585
R733 gnd.n2326 gnd.n1023 585
R734 gnd.n4453 gnd.n4452 585
R735 gnd.n4452 gnd.n4451 585
R736 gnd.n4454 gnd.n1017 585
R737 gnd.n2471 gnd.n1017 585
R738 gnd.n4456 gnd.n4455 585
R739 gnd.n4457 gnd.n4456 585
R740 gnd.n1001 gnd.n1000 585
R741 gnd.n2461 gnd.n1001 585
R742 gnd.n4465 gnd.n4464 585
R743 gnd.n4464 gnd.n4463 585
R744 gnd.n4466 gnd.n995 585
R745 gnd.n1002 gnd.n995 585
R746 gnd.n4468 gnd.n4467 585
R747 gnd.n4469 gnd.n4468 585
R748 gnd.n982 gnd.n981 585
R749 gnd.n985 gnd.n982 585
R750 gnd.n4477 gnd.n4476 585
R751 gnd.n4476 gnd.n4475 585
R752 gnd.n4478 gnd.n976 585
R753 gnd.n976 gnd.n974 585
R754 gnd.n4480 gnd.n4479 585
R755 gnd.n4481 gnd.n4480 585
R756 gnd.n977 gnd.n975 585
R757 gnd.n975 gnd.n962 585
R758 gnd.n2423 gnd.n963 585
R759 gnd.n4487 gnd.n963 585
R760 gnd.n2360 gnd.n2358 585
R761 gnd.n2358 gnd.n960 585
R762 gnd.n2428 gnd.n2427 585
R763 gnd.n2435 gnd.n2428 585
R764 gnd.n2359 gnd.n2357 585
R765 gnd.n2357 gnd.n906 585
R766 gnd.n2419 gnd.n2418 585
R767 gnd.n2417 gnd.n2416 585
R768 gnd.n2415 gnd.n2414 585
R769 gnd.n2413 gnd.n2412 585
R770 gnd.n2411 gnd.n2410 585
R771 gnd.n2409 gnd.n2408 585
R772 gnd.n2407 gnd.n2406 585
R773 gnd.n2405 gnd.n2404 585
R774 gnd.n2403 gnd.n2402 585
R775 gnd.n2401 gnd.n2400 585
R776 gnd.n2399 gnd.n2398 585
R777 gnd.n2397 gnd.n2396 585
R778 gnd.n2395 gnd.n2394 585
R779 gnd.n2393 gnd.n2392 585
R780 gnd.n2391 gnd.n2390 585
R781 gnd.n2389 gnd.n2388 585
R782 gnd.n2387 gnd.n2386 585
R783 gnd.n2379 gnd.n2376 585
R784 gnd.n2382 gnd.n905 585
R785 gnd.n4574 gnd.n905 585
R786 gnd.n2865 gnd.n2864 585
R787 gnd.n2866 gnd.n2017 585
R788 gnd.n2116 gnd.n2014 585
R789 gnd.n2115 gnd.n2114 585
R790 gnd.n2027 gnd.n2026 585
R791 gnd.n2103 gnd.n2102 585
R792 gnd.n2101 gnd.n2100 585
R793 gnd.n2089 gnd.n2034 585
R794 gnd.n2091 gnd.n2090 585
R795 gnd.n2088 gnd.n2040 585
R796 gnd.n2039 gnd.n2038 585
R797 gnd.n2079 gnd.n2078 585
R798 gnd.n2077 gnd.n2076 585
R799 gnd.n2065 gnd.n2046 585
R800 gnd.n2067 gnd.n2066 585
R801 gnd.n2064 gnd.n2054 585
R802 gnd.n2053 gnd.n2052 585
R803 gnd.n2051 gnd.n2050 585
R804 gnd.n1165 gnd.n1163 585
R805 gnd.n2862 gnd.n1163 585
R806 gnd.n2186 gnd.n1161 585
R807 gnd.n4369 gnd.n1161 585
R808 gnd.n2576 gnd.n2575 585
R809 gnd.n2577 gnd.n2576 585
R810 gnd.n2185 gnd.n1152 585
R811 gnd.n4375 gnd.n1152 585
R812 gnd.n2571 gnd.n2570 585
R813 gnd.n2570 gnd.n2569 585
R814 gnd.n2188 gnd.n1141 585
R815 gnd.n4381 gnd.n1141 585
R816 gnd.n2559 gnd.n2558 585
R817 gnd.n2560 gnd.n2559 585
R818 gnd.n2192 gnd.n1130 585
R819 gnd.n4387 gnd.n1130 585
R820 gnd.n2554 gnd.n2553 585
R821 gnd.n2553 gnd.n2552 585
R822 gnd.n2194 gnd.n1119 585
R823 gnd.n4393 gnd.n1119 585
R824 gnd.n2543 gnd.n2542 585
R825 gnd.n2544 gnd.n2543 585
R826 gnd.n2198 gnd.n1108 585
R827 gnd.n4399 gnd.n1108 585
R828 gnd.n2538 gnd.n2537 585
R829 gnd.n2537 gnd.n2536 585
R830 gnd.n2200 gnd.n1098 585
R831 gnd.n4405 gnd.n1098 585
R832 gnd.n2527 gnd.n2526 585
R833 gnd.n2528 gnd.n2527 585
R834 gnd.n2205 gnd.n1087 585
R835 gnd.n4411 gnd.n1087 585
R836 gnd.n2522 gnd.n2521 585
R837 gnd.n2521 gnd.n2520 585
R838 gnd.n2207 gnd.n1076 585
R839 gnd.n4417 gnd.n1076 585
R840 gnd.n2511 gnd.n2510 585
R841 gnd.n2512 gnd.n2511 585
R842 gnd.n2211 gnd.n1068 585
R843 gnd.n4424 gnd.n1068 585
R844 gnd.n2506 gnd.n2505 585
R845 gnd.n2505 gnd.n2504 585
R846 gnd.n2213 gnd.n1059 585
R847 gnd.n4430 gnd.n1059 585
R848 gnd.n2495 gnd.n2494 585
R849 gnd.n2496 gnd.n2495 585
R850 gnd.n2219 gnd.n1051 585
R851 gnd.n4437 gnd.n1051 585
R852 gnd.n2490 gnd.n2489 585
R853 gnd.n2489 gnd.n2488 585
R854 gnd.n2221 gnd.n1037 585
R855 gnd.n4443 gnd.n1037 585
R856 gnd.n2479 gnd.n2478 585
R857 gnd.n2480 gnd.n2479 585
R858 gnd.n2328 gnd.n2327 585
R859 gnd.n2327 gnd.n2326 585
R860 gnd.n2474 gnd.n1026 585
R861 gnd.n4451 gnd.n1026 585
R862 gnd.n2473 gnd.n2472 585
R863 gnd.n2472 gnd.n2471 585
R864 gnd.n2330 gnd.n1015 585
R865 gnd.n4457 gnd.n1015 585
R866 gnd.n2460 gnd.n2459 585
R867 gnd.n2461 gnd.n2460 585
R868 gnd.n2349 gnd.n1004 585
R869 gnd.n4463 gnd.n1004 585
R870 gnd.n2454 gnd.n2453 585
R871 gnd.n2453 gnd.n1002 585
R872 gnd.n2452 gnd.n994 585
R873 gnd.n4469 gnd.n994 585
R874 gnd.n2451 gnd.n2450 585
R875 gnd.n2450 gnd.n985 585
R876 gnd.n2351 gnd.n984 585
R877 gnd.n4475 gnd.n984 585
R878 gnd.n2446 gnd.n2445 585
R879 gnd.n2445 gnd.n974 585
R880 gnd.n2444 gnd.n973 585
R881 gnd.n4481 gnd.n973 585
R882 gnd.n2443 gnd.n2442 585
R883 gnd.n2442 gnd.n962 585
R884 gnd.n2353 gnd.n961 585
R885 gnd.n4487 gnd.n961 585
R886 gnd.n2438 gnd.n2437 585
R887 gnd.n2437 gnd.n960 585
R888 gnd.n2436 gnd.n2355 585
R889 gnd.n2436 gnd.n2435 585
R890 gnd.n2380 gnd.n2356 585
R891 gnd.n2356 gnd.n906 585
R892 gnd.n6866 gnd.n84 585
R893 gnd.n6962 gnd.n84 585
R894 gnd.n6867 gnd.n6798 585
R895 gnd.n6798 gnd.n81 585
R896 gnd.n6868 gnd.n163 585
R897 gnd.n6882 gnd.n163 585
R898 gnd.n175 gnd.n173 585
R899 gnd.n173 gnd.n162 585
R900 gnd.n6873 gnd.n6872 585
R901 gnd.n6874 gnd.n6873 585
R902 gnd.n174 gnd.n172 585
R903 gnd.n172 gnd.n170 585
R904 gnd.n6794 gnd.n6793 585
R905 gnd.n6793 gnd.n6792 585
R906 gnd.n178 gnd.n177 585
R907 gnd.n188 gnd.n178 585
R908 gnd.n6783 gnd.n6782 585
R909 gnd.n6784 gnd.n6783 585
R910 gnd.n190 gnd.n189 585
R911 gnd.n189 gnd.n186 585
R912 gnd.n6778 gnd.n6777 585
R913 gnd.n6777 gnd.n6776 585
R914 gnd.n193 gnd.n192 585
R915 gnd.n194 gnd.n193 585
R916 gnd.n6767 gnd.n6766 585
R917 gnd.n6768 gnd.n6767 585
R918 gnd.n204 gnd.n203 585
R919 gnd.n268 gnd.n203 585
R920 gnd.n6762 gnd.n6761 585
R921 gnd.n6761 gnd.n6760 585
R922 gnd.n207 gnd.n206 585
R923 gnd.n6728 gnd.n207 585
R924 gnd.n6751 gnd.n6750 585
R925 gnd.n6752 gnd.n6751 585
R926 gnd.n225 gnd.n224 585
R927 gnd.n6733 gnd.n224 585
R928 gnd.n6746 gnd.n6745 585
R929 gnd.n6745 gnd.n6744 585
R930 gnd.n228 gnd.n227 585
R931 gnd.n6739 gnd.n228 585
R932 gnd.n4117 gnd.n4116 585
R933 gnd.n4116 gnd.n4115 585
R934 gnd.n1396 gnd.n1393 585
R935 gnd.n4099 gnd.n1396 585
R936 gnd.n4121 gnd.n1392 585
R937 gnd.n1402 gnd.n1392 585
R938 gnd.n4122 gnd.n1391 585
R939 gnd.n4091 gnd.n1391 585
R940 gnd.n4123 gnd.n1390 585
R941 gnd.n4071 gnd.n1390 585
R942 gnd.n1417 gnd.n1388 585
R943 gnd.n4082 gnd.n1417 585
R944 gnd.n4127 gnd.n1387 585
R945 gnd.n4077 gnd.n1387 585
R946 gnd.n4128 gnd.n1386 585
R947 gnd.n4059 gnd.n1386 585
R948 gnd.n4129 gnd.n1385 585
R949 gnd.n1437 gnd.n1385 585
R950 gnd.n1446 gnd.n1383 585
R951 gnd.n4051 gnd.n1446 585
R952 gnd.n4133 gnd.n1382 585
R953 gnd.n3936 gnd.n1382 585
R954 gnd.n4134 gnd.n1381 585
R955 gnd.n4040 gnd.n1381 585
R956 gnd.n4135 gnd.n1380 585
R957 gnd.n4025 gnd.n1380 585
R958 gnd.n3941 gnd.n1378 585
R959 gnd.n3942 gnd.n3941 585
R960 gnd.n4139 gnd.n1377 585
R961 gnd.n4016 gnd.n1377 585
R962 gnd.n4140 gnd.n1376 585
R963 gnd.n3946 gnd.n1376 585
R964 gnd.n4141 gnd.n1375 585
R965 gnd.n4006 gnd.n1375 585
R966 gnd.n3993 gnd.n1373 585
R967 gnd.n3994 gnd.n3993 585
R968 gnd.n4145 gnd.n1372 585
R969 gnd.n1487 gnd.n1372 585
R970 gnd.n4146 gnd.n1371 585
R971 gnd.n3984 gnd.n1371 585
R972 gnd.n4147 gnd.n1370 585
R973 gnd.n3956 gnd.n1370 585
R974 gnd.n1367 gnd.n1366 585
R975 gnd.n3974 gnd.n1366 585
R976 gnd.n4152 gnd.n4151 585
R977 gnd.n4153 gnd.n4152 585
R978 gnd.n1548 gnd.n1365 585
R979 gnd.n1552 gnd.n1551 585
R980 gnd.n1554 gnd.n1553 585
R981 gnd.n1543 gnd.n1542 585
R982 gnd.n1566 gnd.n1544 585
R983 gnd.n1568 gnd.n1567 585
R984 gnd.n1570 gnd.n1569 585
R985 gnd.n1534 gnd.n1533 585
R986 gnd.n1583 gnd.n1535 585
R987 gnd.n1585 gnd.n1584 585
R988 gnd.n1587 gnd.n1586 585
R989 gnd.n1525 gnd.n1524 585
R990 gnd.n1600 gnd.n1526 585
R991 gnd.n1602 gnd.n1601 585
R992 gnd.n1604 gnd.n1603 585
R993 gnd.n1516 gnd.n1515 585
R994 gnd.n1617 gnd.n1517 585
R995 gnd.n1618 gnd.n1512 585
R996 gnd.n1619 gnd.n1310 585
R997 gnd.n4229 gnd.n1310 585
R998 gnd.n6837 gnd.n80 585
R999 gnd.n6838 gnd.n6836 585
R1000 gnd.n6839 gnd.n6832 585
R1001 gnd.n6830 gnd.n6828 585
R1002 gnd.n6843 gnd.n6827 585
R1003 gnd.n6844 gnd.n6825 585
R1004 gnd.n6845 gnd.n6824 585
R1005 gnd.n6822 gnd.n6820 585
R1006 gnd.n6849 gnd.n6819 585
R1007 gnd.n6850 gnd.n6817 585
R1008 gnd.n6851 gnd.n6816 585
R1009 gnd.n6814 gnd.n6812 585
R1010 gnd.n6855 gnd.n6811 585
R1011 gnd.n6856 gnd.n6809 585
R1012 gnd.n6857 gnd.n6808 585
R1013 gnd.n6806 gnd.n6804 585
R1014 gnd.n6861 gnd.n6803 585
R1015 gnd.n6862 gnd.n6801 585
R1016 gnd.n6863 gnd.n6800 585
R1017 gnd.n6800 gnd.n94 585
R1018 gnd.n6964 gnd.n6963 585
R1019 gnd.n6963 gnd.n6962 585
R1020 gnd.n79 gnd.n77 585
R1021 gnd.n81 gnd.n79 585
R1022 gnd.n6968 gnd.n76 585
R1023 gnd.n6882 gnd.n76 585
R1024 gnd.n6969 gnd.n75 585
R1025 gnd.n162 gnd.n75 585
R1026 gnd.n6970 gnd.n74 585
R1027 gnd.n6874 gnd.n74 585
R1028 gnd.n169 gnd.n72 585
R1029 gnd.n170 gnd.n169 585
R1030 gnd.n6974 gnd.n71 585
R1031 gnd.n6792 gnd.n71 585
R1032 gnd.n6975 gnd.n70 585
R1033 gnd.n188 gnd.n70 585
R1034 gnd.n6976 gnd.n69 585
R1035 gnd.n6784 gnd.n69 585
R1036 gnd.n185 gnd.n67 585
R1037 gnd.n186 gnd.n185 585
R1038 gnd.n6980 gnd.n66 585
R1039 gnd.n6776 gnd.n66 585
R1040 gnd.n6981 gnd.n65 585
R1041 gnd.n194 gnd.n65 585
R1042 gnd.n6982 gnd.n64 585
R1043 gnd.n6768 gnd.n64 585
R1044 gnd.n267 gnd.n62 585
R1045 gnd.n268 gnd.n267 585
R1046 gnd.n6986 gnd.n61 585
R1047 gnd.n6760 gnd.n61 585
R1048 gnd.n6987 gnd.n60 585
R1049 gnd.n6728 gnd.n60 585
R1050 gnd.n6988 gnd.n59 585
R1051 gnd.n6752 gnd.n59 585
R1052 gnd.n6732 gnd.n57 585
R1053 gnd.n6733 gnd.n6732 585
R1054 gnd.n6992 gnd.n56 585
R1055 gnd.n6744 gnd.n56 585
R1056 gnd.n6993 gnd.n55 585
R1057 gnd.n6739 gnd.n55 585
R1058 gnd.n6994 gnd.n54 585
R1059 gnd.n4115 gnd.n54 585
R1060 gnd.n1404 gnd.n52 585
R1061 gnd.n4099 gnd.n1404 585
R1062 gnd.n1411 gnd.n1409 585
R1063 gnd.n1409 gnd.n1402 585
R1064 gnd.n4089 gnd.n4088 585
R1065 gnd.n4091 gnd.n4089 585
R1066 gnd.n1410 gnd.n1408 585
R1067 gnd.n4071 gnd.n1408 585
R1068 gnd.n4084 gnd.n4083 585
R1069 gnd.n4083 gnd.n4082 585
R1070 gnd.n1414 gnd.n1413 585
R1071 gnd.n4077 gnd.n1414 585
R1072 gnd.n4058 gnd.n4057 585
R1073 gnd.n4059 gnd.n4058 585
R1074 gnd.n1439 gnd.n1438 585
R1075 gnd.n1438 gnd.n1437 585
R1076 gnd.n4053 gnd.n4052 585
R1077 gnd.n4052 gnd.n4051 585
R1078 gnd.n1442 gnd.n1441 585
R1079 gnd.n3936 gnd.n1442 585
R1080 gnd.n1465 gnd.n1455 585
R1081 gnd.n4040 gnd.n1455 585
R1082 gnd.n4024 gnd.n4023 585
R1083 gnd.n4025 gnd.n4024 585
R1084 gnd.n1464 gnd.n1463 585
R1085 gnd.n3942 gnd.n1463 585
R1086 gnd.n4018 gnd.n4017 585
R1087 gnd.n4017 gnd.n4016 585
R1088 gnd.n1468 gnd.n1467 585
R1089 gnd.n3946 gnd.n1468 585
R1090 gnd.n1491 gnd.n1480 585
R1091 gnd.n4006 gnd.n1480 585
R1092 gnd.n3992 gnd.n3991 585
R1093 gnd.n3994 gnd.n3992 585
R1094 gnd.n1490 gnd.n1489 585
R1095 gnd.n1489 gnd.n1487 585
R1096 gnd.n3986 gnd.n3985 585
R1097 gnd.n3985 gnd.n3984 585
R1098 gnd.n1494 gnd.n1493 585
R1099 gnd.n3956 gnd.n1494 585
R1100 gnd.n3916 gnd.n3915 585
R1101 gnd.n3974 gnd.n3916 585
R1102 gnd.n1503 gnd.n1363 585
R1103 gnd.n4153 gnd.n1363 585
R1104 gnd.n850 gnd.n849 585
R1105 gnd.n853 gnd.n850 585
R1106 gnd.n5925 gnd.n5924 585
R1107 gnd.n5924 gnd.n5923 585
R1108 gnd.n5926 gnd.n844 585
R1109 gnd.n5822 gnd.n844 585
R1110 gnd.n5928 gnd.n5927 585
R1111 gnd.n5929 gnd.n5928 585
R1112 gnd.n845 gnd.n843 585
R1113 gnd.n843 gnd.n839 585
R1114 gnd.n825 gnd.n824 585
R1115 gnd.n828 gnd.n825 585
R1116 gnd.n5939 gnd.n5938 585
R1117 gnd.n5938 gnd.n5937 585
R1118 gnd.n5940 gnd.n819 585
R1119 gnd.n5543 gnd.n819 585
R1120 gnd.n5942 gnd.n5941 585
R1121 gnd.n5943 gnd.n5942 585
R1122 gnd.n820 gnd.n818 585
R1123 gnd.n5527 gnd.n818 585
R1124 gnd.n5518 gnd.n5517 585
R1125 gnd.n5517 gnd.n806 585
R1126 gnd.n5516 gnd.n4647 585
R1127 gnd.n5516 gnd.n804 585
R1128 gnd.n5515 gnd.n4649 585
R1129 gnd.n5515 gnd.n5514 585
R1130 gnd.n5505 gnd.n4648 585
R1131 gnd.n4660 gnd.n4648 585
R1132 gnd.n5504 gnd.n5503 585
R1133 gnd.n5503 gnd.n5502 585
R1134 gnd.n4657 gnd.n4655 585
R1135 gnd.n5489 gnd.n4657 585
R1136 gnd.n5480 gnd.n5479 585
R1137 gnd.n5479 gnd.n5478 585
R1138 gnd.n4672 gnd.n4671 585
R1139 gnd.n4680 gnd.n4672 585
R1140 gnd.n5457 gnd.n5456 585
R1141 gnd.n5458 gnd.n5457 585
R1142 gnd.n4683 gnd.n4682 585
R1143 gnd.n4691 gnd.n4682 585
R1144 gnd.n5431 gnd.n4703 585
R1145 gnd.n4703 gnd.n4690 585
R1146 gnd.n5433 gnd.n5432 585
R1147 gnd.n5434 gnd.n5433 585
R1148 gnd.n4704 gnd.n4702 585
R1149 gnd.n4702 gnd.n4698 585
R1150 gnd.n5420 gnd.n5419 585
R1151 gnd.n5419 gnd.n5418 585
R1152 gnd.n4709 gnd.n4708 585
R1153 gnd.n4719 gnd.n4709 585
R1154 gnd.n5409 gnd.n5408 585
R1155 gnd.n5408 gnd.n5407 585
R1156 gnd.n4716 gnd.n4715 585
R1157 gnd.n5395 gnd.n4716 585
R1158 gnd.n5369 gnd.n4773 585
R1159 gnd.n4773 gnd.n4726 585
R1160 gnd.n5371 gnd.n5370 585
R1161 gnd.n5372 gnd.n5371 585
R1162 gnd.n4774 gnd.n4772 585
R1163 gnd.n4782 gnd.n4772 585
R1164 gnd.n5347 gnd.n4794 585
R1165 gnd.n4794 gnd.n4781 585
R1166 gnd.n5349 gnd.n5348 585
R1167 gnd.n5350 gnd.n5349 585
R1168 gnd.n4795 gnd.n4793 585
R1169 gnd.n4793 gnd.n4789 585
R1170 gnd.n5335 gnd.n5334 585
R1171 gnd.n5334 gnd.n5333 585
R1172 gnd.n4800 gnd.n4799 585
R1173 gnd.n4809 gnd.n4800 585
R1174 gnd.n5324 gnd.n5323 585
R1175 gnd.n5323 gnd.n5322 585
R1176 gnd.n4807 gnd.n4806 585
R1177 gnd.n5310 gnd.n4807 585
R1178 gnd.n5282 gnd.n5281 585
R1179 gnd.n5281 gnd.n4816 585
R1180 gnd.n5283 gnd.n4827 585
R1181 gnd.n5274 gnd.n4827 585
R1182 gnd.n5285 gnd.n5284 585
R1183 gnd.n5286 gnd.n5285 585
R1184 gnd.n4828 gnd.n4826 585
R1185 gnd.n4842 gnd.n4826 585
R1186 gnd.n5266 gnd.n5265 585
R1187 gnd.n5265 gnd.n5264 585
R1188 gnd.n4839 gnd.n4838 585
R1189 gnd.n5249 gnd.n4839 585
R1190 gnd.n5236 gnd.n4859 585
R1191 gnd.n4859 gnd.n4849 585
R1192 gnd.n5238 gnd.n5237 585
R1193 gnd.n5239 gnd.n5238 585
R1194 gnd.n4860 gnd.n4858 585
R1195 gnd.n4868 gnd.n4858 585
R1196 gnd.n5212 gnd.n4880 585
R1197 gnd.n4880 gnd.n4867 585
R1198 gnd.n5214 gnd.n5213 585
R1199 gnd.n5215 gnd.n5214 585
R1200 gnd.n4881 gnd.n4879 585
R1201 gnd.n4879 gnd.n4875 585
R1202 gnd.n5200 gnd.n5199 585
R1203 gnd.n5199 gnd.n5198 585
R1204 gnd.n4886 gnd.n4885 585
R1205 gnd.n4890 gnd.n4886 585
R1206 gnd.n5184 gnd.n5183 585
R1207 gnd.n5185 gnd.n5184 585
R1208 gnd.n4901 gnd.n4900 585
R1209 gnd.n4900 gnd.n4896 585
R1210 gnd.n5174 gnd.n5173 585
R1211 gnd.n5175 gnd.n5174 585
R1212 gnd.n4910 gnd.n4909 585
R1213 gnd.n4909 gnd.n4907 585
R1214 gnd.n5168 gnd.n5167 585
R1215 gnd.n5167 gnd.n5166 585
R1216 gnd.n4914 gnd.n4913 585
R1217 gnd.n4922 gnd.n4914 585
R1218 gnd.n5075 gnd.n5074 585
R1219 gnd.n5076 gnd.n5075 585
R1220 gnd.n4924 gnd.n4923 585
R1221 gnd.n4923 gnd.n4921 585
R1222 gnd.n5070 gnd.n5069 585
R1223 gnd.n5069 gnd.n5068 585
R1224 gnd.n4927 gnd.n4926 585
R1225 gnd.n4928 gnd.n4927 585
R1226 gnd.n5059 gnd.n5058 585
R1227 gnd.n5060 gnd.n5059 585
R1228 gnd.n4936 gnd.n4935 585
R1229 gnd.n4935 gnd.n4934 585
R1230 gnd.n5054 gnd.n5053 585
R1231 gnd.n5053 gnd.n5052 585
R1232 gnd.n4939 gnd.n4938 585
R1233 gnd.n4940 gnd.n4939 585
R1234 gnd.n5043 gnd.n5042 585
R1235 gnd.n5044 gnd.n5043 585
R1236 gnd.n5039 gnd.n4946 585
R1237 gnd.n5038 gnd.n5037 585
R1238 gnd.n5035 gnd.n4948 585
R1239 gnd.n5035 gnd.n4945 585
R1240 gnd.n5034 gnd.n5033 585
R1241 gnd.n5032 gnd.n5031 585
R1242 gnd.n5030 gnd.n4953 585
R1243 gnd.n5028 gnd.n5027 585
R1244 gnd.n5026 gnd.n4954 585
R1245 gnd.n5025 gnd.n5024 585
R1246 gnd.n5022 gnd.n4959 585
R1247 gnd.n5020 gnd.n5019 585
R1248 gnd.n5018 gnd.n4960 585
R1249 gnd.n5017 gnd.n5016 585
R1250 gnd.n5014 gnd.n4965 585
R1251 gnd.n5012 gnd.n5011 585
R1252 gnd.n5010 gnd.n4966 585
R1253 gnd.n5009 gnd.n5008 585
R1254 gnd.n5006 gnd.n4971 585
R1255 gnd.n5004 gnd.n5003 585
R1256 gnd.n5002 gnd.n4972 585
R1257 gnd.n5001 gnd.n5000 585
R1258 gnd.n4998 gnd.n4977 585
R1259 gnd.n4996 gnd.n4995 585
R1260 gnd.n4993 gnd.n4978 585
R1261 gnd.n4992 gnd.n4991 585
R1262 gnd.n4989 gnd.n4987 585
R1263 gnd.n4985 gnd.n4944 585
R1264 gnd.n5831 gnd.n5830 585
R1265 gnd.n5833 gnd.n5832 585
R1266 gnd.n5835 gnd.n5834 585
R1267 gnd.n5837 gnd.n5836 585
R1268 gnd.n5839 gnd.n5838 585
R1269 gnd.n5841 gnd.n5840 585
R1270 gnd.n5843 gnd.n5842 585
R1271 gnd.n5845 gnd.n5844 585
R1272 gnd.n5847 gnd.n5846 585
R1273 gnd.n5849 gnd.n5848 585
R1274 gnd.n5851 gnd.n5850 585
R1275 gnd.n5853 gnd.n5852 585
R1276 gnd.n5855 gnd.n5854 585
R1277 gnd.n5857 gnd.n5856 585
R1278 gnd.n5859 gnd.n5858 585
R1279 gnd.n5861 gnd.n5860 585
R1280 gnd.n5863 gnd.n5862 585
R1281 gnd.n5865 gnd.n5864 585
R1282 gnd.n5867 gnd.n5866 585
R1283 gnd.n5869 gnd.n5868 585
R1284 gnd.n5871 gnd.n5870 585
R1285 gnd.n5873 gnd.n5872 585
R1286 gnd.n5875 gnd.n5874 585
R1287 gnd.n5877 gnd.n5876 585
R1288 gnd.n5879 gnd.n5878 585
R1289 gnd.n5880 gnd.n4601 585
R1290 gnd.n5881 gnd.n864 585
R1291 gnd.n5914 gnd.n864 585
R1292 gnd.n5829 gnd.n5828 585
R1293 gnd.n5829 gnd.n853 585
R1294 gnd.n4630 gnd.n851 585
R1295 gnd.n5923 gnd.n851 585
R1296 gnd.n5824 gnd.n5823 585
R1297 gnd.n5823 gnd.n5822 585
R1298 gnd.n4632 gnd.n841 585
R1299 gnd.n5929 gnd.n841 585
R1300 gnd.n5537 gnd.n5536 585
R1301 gnd.n5537 gnd.n839 585
R1302 gnd.n5539 gnd.n5538 585
R1303 gnd.n5538 gnd.n828 585
R1304 gnd.n5540 gnd.n826 585
R1305 gnd.n5937 gnd.n826 585
R1306 gnd.n5542 gnd.n5541 585
R1307 gnd.n5543 gnd.n5542 585
R1308 gnd.n4641 gnd.n816 585
R1309 gnd.n5943 gnd.n816 585
R1310 gnd.n5529 gnd.n5528 585
R1311 gnd.n5528 gnd.n5527 585
R1312 gnd.n4644 gnd.n4643 585
R1313 gnd.n4644 gnd.n806 585
R1314 gnd.n5470 gnd.n5469 585
R1315 gnd.n5469 gnd.n804 585
R1316 gnd.n5471 gnd.n4651 585
R1317 gnd.n5514 gnd.n4651 585
R1318 gnd.n5473 gnd.n5472 585
R1319 gnd.n5472 gnd.n4660 585
R1320 gnd.n5474 gnd.n4658 585
R1321 gnd.n5502 gnd.n4658 585
R1322 gnd.n5475 gnd.n4668 585
R1323 gnd.n5489 gnd.n4668 585
R1324 gnd.n5477 gnd.n5476 585
R1325 gnd.n5478 gnd.n5477 585
R1326 gnd.n4675 gnd.n4674 585
R1327 gnd.n4680 gnd.n4674 585
R1328 gnd.n5460 gnd.n5459 585
R1329 gnd.n5459 gnd.n5458 585
R1330 gnd.n4678 gnd.n4677 585
R1331 gnd.n4691 gnd.n4678 585
R1332 gnd.n5385 gnd.n5384 585
R1333 gnd.n5384 gnd.n4690 585
R1334 gnd.n5386 gnd.n4700 585
R1335 gnd.n5434 gnd.n4700 585
R1336 gnd.n5388 gnd.n5387 585
R1337 gnd.n5387 gnd.n4698 585
R1338 gnd.n5389 gnd.n4711 585
R1339 gnd.n5418 gnd.n4711 585
R1340 gnd.n5391 gnd.n5390 585
R1341 gnd.n5390 gnd.n4719 585
R1342 gnd.n5392 gnd.n4718 585
R1343 gnd.n5407 gnd.n4718 585
R1344 gnd.n5394 gnd.n5393 585
R1345 gnd.n5395 gnd.n5394 585
R1346 gnd.n4730 gnd.n4729 585
R1347 gnd.n4729 gnd.n4726 585
R1348 gnd.n5374 gnd.n5373 585
R1349 gnd.n5373 gnd.n5372 585
R1350 gnd.n4769 gnd.n4768 585
R1351 gnd.n4782 gnd.n4769 585
R1352 gnd.n5295 gnd.n5294 585
R1353 gnd.n5294 gnd.n4781 585
R1354 gnd.n5296 gnd.n4791 585
R1355 gnd.n5350 gnd.n4791 585
R1356 gnd.n5299 gnd.n5298 585
R1357 gnd.n5298 gnd.n4789 585
R1358 gnd.n5300 gnd.n4802 585
R1359 gnd.n5333 gnd.n4802 585
R1360 gnd.n5303 gnd.n5302 585
R1361 gnd.n5302 gnd.n4809 585
R1362 gnd.n5304 gnd.n4808 585
R1363 gnd.n5322 gnd.n4808 585
R1364 gnd.n5307 gnd.n5306 585
R1365 gnd.n5310 gnd.n5307 585
R1366 gnd.n5292 gnd.n4818 585
R1367 gnd.n4818 gnd.n4816 585
R1368 gnd.n4823 gnd.n4819 585
R1369 gnd.n5274 gnd.n4823 585
R1370 gnd.n5288 gnd.n5287 585
R1371 gnd.n5287 gnd.n5286 585
R1372 gnd.n4822 gnd.n4821 585
R1373 gnd.n4842 gnd.n4822 585
R1374 gnd.n5246 gnd.n4841 585
R1375 gnd.n5264 gnd.n4841 585
R1376 gnd.n5248 gnd.n5247 585
R1377 gnd.n5249 gnd.n5248 585
R1378 gnd.n4852 gnd.n4851 585
R1379 gnd.n4851 gnd.n4849 585
R1380 gnd.n5241 gnd.n5240 585
R1381 gnd.n5240 gnd.n5239 585
R1382 gnd.n4855 gnd.n4854 585
R1383 gnd.n4868 gnd.n4855 585
R1384 gnd.n5092 gnd.n5091 585
R1385 gnd.n5091 gnd.n4867 585
R1386 gnd.n5093 gnd.n4877 585
R1387 gnd.n5215 gnd.n4877 585
R1388 gnd.n5095 gnd.n5094 585
R1389 gnd.n5094 gnd.n4875 585
R1390 gnd.n5096 gnd.n4887 585
R1391 gnd.n5198 gnd.n4887 585
R1392 gnd.n5098 gnd.n5097 585
R1393 gnd.n5097 gnd.n4890 585
R1394 gnd.n5099 gnd.n4898 585
R1395 gnd.n5185 gnd.n4898 585
R1396 gnd.n5101 gnd.n5100 585
R1397 gnd.n5100 gnd.n4896 585
R1398 gnd.n5102 gnd.n4908 585
R1399 gnd.n5175 gnd.n4908 585
R1400 gnd.n5103 gnd.n4916 585
R1401 gnd.n4916 gnd.n4907 585
R1402 gnd.n5105 gnd.n5104 585
R1403 gnd.n5166 gnd.n5105 585
R1404 gnd.n4917 gnd.n4915 585
R1405 gnd.n4922 gnd.n4915 585
R1406 gnd.n5078 gnd.n5077 585
R1407 gnd.n5077 gnd.n5076 585
R1408 gnd.n4920 gnd.n4919 585
R1409 gnd.n4921 gnd.n4920 585
R1410 gnd.n5067 gnd.n5066 585
R1411 gnd.n5068 gnd.n5067 585
R1412 gnd.n4930 gnd.n4929 585
R1413 gnd.n4929 gnd.n4928 585
R1414 gnd.n5062 gnd.n5061 585
R1415 gnd.n5061 gnd.n5060 585
R1416 gnd.n4933 gnd.n4932 585
R1417 gnd.n4934 gnd.n4933 585
R1418 gnd.n5051 gnd.n5050 585
R1419 gnd.n5052 gnd.n5051 585
R1420 gnd.n4942 gnd.n4941 585
R1421 gnd.n4941 gnd.n4940 585
R1422 gnd.n5046 gnd.n5045 585
R1423 gnd.n5045 gnd.n5044 585
R1424 gnd.n5919 gnd.n855 585
R1425 gnd.n863 gnd.n855 585
R1426 gnd.n5921 gnd.n5920 585
R1427 gnd.n5922 gnd.n5921 585
R1428 gnd.n856 gnd.n854 585
R1429 gnd.n5821 gnd.n854 585
R1430 gnd.n838 gnd.n837 585
R1431 gnd.n842 gnd.n838 585
R1432 gnd.n5932 gnd.n5931 585
R1433 gnd.n5931 gnd.n5930 585
R1434 gnd.n5933 gnd.n830 585
R1435 gnd.n4634 gnd.n830 585
R1436 gnd.n5935 gnd.n5934 585
R1437 gnd.n5936 gnd.n5935 585
R1438 gnd.n831 gnd.n829 585
R1439 gnd.n5544 gnd.n829 585
R1440 gnd.n814 gnd.n813 585
R1441 gnd.n817 gnd.n814 585
R1442 gnd.n5946 gnd.n5945 585
R1443 gnd.n5945 gnd.n5944 585
R1444 gnd.n5947 gnd.n808 585
R1445 gnd.n5526 gnd.n808 585
R1446 gnd.n5949 gnd.n5948 585
R1447 gnd.n5950 gnd.n5949 585
R1448 gnd.n809 gnd.n807 585
R1449 gnd.n5513 gnd.n807 585
R1450 gnd.n5498 gnd.n4662 585
R1451 gnd.n4662 gnd.n4650 585
R1452 gnd.n5500 gnd.n5499 585
R1453 gnd.n5501 gnd.n5500 585
R1454 gnd.n4663 gnd.n4661 585
R1455 gnd.n5488 gnd.n4661 585
R1456 gnd.n5492 gnd.n5491 585
R1457 gnd.n5491 gnd.n5490 585
R1458 gnd.n4666 gnd.n4665 585
R1459 gnd.n4673 gnd.n4666 585
R1460 gnd.n5444 gnd.n5443 585
R1461 gnd.n5443 gnd.n4681 585
R1462 gnd.n5445 gnd.n4693 585
R1463 gnd.n4693 gnd.n4679 585
R1464 gnd.n5447 gnd.n5446 585
R1465 gnd.n5448 gnd.n5447 585
R1466 gnd.n4694 gnd.n4692 585
R1467 gnd.n4701 gnd.n4692 585
R1468 gnd.n5437 gnd.n5436 585
R1469 gnd.n5436 gnd.n5435 585
R1470 gnd.n4697 gnd.n4696 585
R1471 gnd.n5417 gnd.n4697 585
R1472 gnd.n5403 gnd.n4721 585
R1473 gnd.n4721 gnd.n4710 585
R1474 gnd.n5405 gnd.n5404 585
R1475 gnd.n5406 gnd.n5405 585
R1476 gnd.n4722 gnd.n4720 585
R1477 gnd.n4720 gnd.n4717 585
R1478 gnd.n5398 gnd.n5397 585
R1479 gnd.n5397 gnd.n5396 585
R1480 gnd.n4725 gnd.n4724 585
R1481 gnd.n4771 gnd.n4725 585
R1482 gnd.n5358 gnd.n4784 585
R1483 gnd.n4784 gnd.n4770 585
R1484 gnd.n5360 gnd.n5359 585
R1485 gnd.n5361 gnd.n5360 585
R1486 gnd.n4785 gnd.n4783 585
R1487 gnd.n4792 gnd.n4783 585
R1488 gnd.n5353 gnd.n5352 585
R1489 gnd.n5352 gnd.n5351 585
R1490 gnd.n4788 gnd.n4787 585
R1491 gnd.n5332 gnd.n4788 585
R1492 gnd.n5318 gnd.n4811 585
R1493 gnd.n4811 gnd.n4801 585
R1494 gnd.n5320 gnd.n5319 585
R1495 gnd.n5321 gnd.n5320 585
R1496 gnd.n4812 gnd.n4810 585
R1497 gnd.n5309 gnd.n4810 585
R1498 gnd.n5313 gnd.n5312 585
R1499 gnd.n5312 gnd.n5311 585
R1500 gnd.n4815 gnd.n4814 585
R1501 gnd.n5275 gnd.n4815 585
R1502 gnd.n5259 gnd.n5258 585
R1503 gnd.n5258 gnd.n4825 585
R1504 gnd.n5260 gnd.n4844 585
R1505 gnd.n4844 gnd.n4824 585
R1506 gnd.n5262 gnd.n5261 585
R1507 gnd.n5263 gnd.n5262 585
R1508 gnd.n4845 gnd.n4843 585
R1509 gnd.n4843 gnd.n4840 585
R1510 gnd.n5252 gnd.n5251 585
R1511 gnd.n5251 gnd.n5250 585
R1512 gnd.n4848 gnd.n4847 585
R1513 gnd.n4857 gnd.n4848 585
R1514 gnd.n5223 gnd.n4870 585
R1515 gnd.n4870 gnd.n4856 585
R1516 gnd.n5225 gnd.n5224 585
R1517 gnd.n5226 gnd.n5225 585
R1518 gnd.n4871 gnd.n4869 585
R1519 gnd.n4878 gnd.n4869 585
R1520 gnd.n5218 gnd.n5217 585
R1521 gnd.n5217 gnd.n5216 585
R1522 gnd.n4874 gnd.n4873 585
R1523 gnd.n5197 gnd.n4874 585
R1524 gnd.n5193 gnd.n5192 585
R1525 gnd.n5194 gnd.n5193 585
R1526 gnd.n4892 gnd.n4891 585
R1527 gnd.n4899 gnd.n4891 585
R1528 gnd.n5188 gnd.n5187 585
R1529 gnd.n5187 gnd.n5186 585
R1530 gnd.n4895 gnd.n4894 585
R1531 gnd.n5176 gnd.n4895 585
R1532 gnd.n5163 gnd.n5162 585
R1533 gnd.n5161 gnd.n5114 585
R1534 gnd.n5160 gnd.n5113 585
R1535 gnd.n5165 gnd.n5113 585
R1536 gnd.n5159 gnd.n5158 585
R1537 gnd.n5157 gnd.n5156 585
R1538 gnd.n5155 gnd.n5154 585
R1539 gnd.n5153 gnd.n5152 585
R1540 gnd.n5151 gnd.n5150 585
R1541 gnd.n5149 gnd.n5148 585
R1542 gnd.n5147 gnd.n5146 585
R1543 gnd.n5145 gnd.n5144 585
R1544 gnd.n5143 gnd.n5142 585
R1545 gnd.n5141 gnd.n5140 585
R1546 gnd.n5139 gnd.n5138 585
R1547 gnd.n5137 gnd.n5136 585
R1548 gnd.n5135 gnd.n5134 585
R1549 gnd.n5130 gnd.n4906 585
R1550 gnd.n5815 gnd.n4596 585
R1551 gnd.n5887 gnd.n5886 585
R1552 gnd.n5889 gnd.n5888 585
R1553 gnd.n5891 gnd.n5890 585
R1554 gnd.n5893 gnd.n5892 585
R1555 gnd.n5895 gnd.n5894 585
R1556 gnd.n5897 gnd.n5896 585
R1557 gnd.n5899 gnd.n5898 585
R1558 gnd.n5901 gnd.n5900 585
R1559 gnd.n5903 gnd.n5902 585
R1560 gnd.n5905 gnd.n5904 585
R1561 gnd.n5907 gnd.n5906 585
R1562 gnd.n5909 gnd.n5908 585
R1563 gnd.n5910 gnd.n4582 585
R1564 gnd.n5912 gnd.n5911 585
R1565 gnd.n862 gnd.n861 585
R1566 gnd.n5916 gnd.n5915 585
R1567 gnd.n5915 gnd.n5914 585
R1568 gnd.n5817 gnd.n5816 585
R1569 gnd.n5816 gnd.n863 585
R1570 gnd.n5818 gnd.n852 585
R1571 gnd.n5922 gnd.n852 585
R1572 gnd.n5820 gnd.n5819 585
R1573 gnd.n5821 gnd.n5820 585
R1574 gnd.n5811 gnd.n4633 585
R1575 gnd.n4633 gnd.n842 585
R1576 gnd.n5809 gnd.n840 585
R1577 gnd.n5930 gnd.n840 585
R1578 gnd.n4636 gnd.n4635 585
R1579 gnd.n4635 gnd.n4634 585
R1580 gnd.n5547 gnd.n827 585
R1581 gnd.n5936 gnd.n827 585
R1582 gnd.n5546 gnd.n5545 585
R1583 gnd.n5545 gnd.n5544 585
R1584 gnd.n4640 gnd.n4638 585
R1585 gnd.n4640 gnd.n817 585
R1586 gnd.n5523 gnd.n815 585
R1587 gnd.n5944 gnd.n815 585
R1588 gnd.n5525 gnd.n5524 585
R1589 gnd.n5526 gnd.n5525 585
R1590 gnd.n4645 gnd.n805 585
R1591 gnd.n5950 gnd.n805 585
R1592 gnd.n5512 gnd.n5511 585
R1593 gnd.n5513 gnd.n5512 585
R1594 gnd.n4653 gnd.n4652 585
R1595 gnd.n4652 gnd.n4650 585
R1596 gnd.n5485 gnd.n4659 585
R1597 gnd.n5501 gnd.n4659 585
R1598 gnd.n5487 gnd.n5486 585
R1599 gnd.n5488 gnd.n5487 585
R1600 gnd.n4669 gnd.n4667 585
R1601 gnd.n5490 gnd.n4667 585
R1602 gnd.n5451 gnd.n4687 585
R1603 gnd.n5451 gnd.n4673 585
R1604 gnd.n5453 gnd.n5452 585
R1605 gnd.n5452 gnd.n4681 585
R1606 gnd.n5450 gnd.n4686 585
R1607 gnd.n5450 gnd.n4679 585
R1608 gnd.n5449 gnd.n4689 585
R1609 gnd.n5449 gnd.n5448 585
R1610 gnd.n5426 gnd.n4688 585
R1611 gnd.n4701 gnd.n4688 585
R1612 gnd.n5425 gnd.n4699 585
R1613 gnd.n5435 gnd.n4699 585
R1614 gnd.n5416 gnd.n4706 585
R1615 gnd.n5417 gnd.n5416 585
R1616 gnd.n5415 gnd.n5414 585
R1617 gnd.n5415 gnd.n4710 585
R1618 gnd.n5413 gnd.n4712 585
R1619 gnd.n5406 gnd.n4712 585
R1620 gnd.n4727 gnd.n4713 585
R1621 gnd.n4727 gnd.n4717 585
R1622 gnd.n5366 gnd.n4728 585
R1623 gnd.n5396 gnd.n4728 585
R1624 gnd.n5365 gnd.n5364 585
R1625 gnd.n5364 gnd.n4771 585
R1626 gnd.n5363 gnd.n4778 585
R1627 gnd.n5363 gnd.n4770 585
R1628 gnd.n5362 gnd.n4780 585
R1629 gnd.n5362 gnd.n5361 585
R1630 gnd.n5341 gnd.n4779 585
R1631 gnd.n4792 gnd.n4779 585
R1632 gnd.n5340 gnd.n4790 585
R1633 gnd.n5351 gnd.n4790 585
R1634 gnd.n5331 gnd.n4797 585
R1635 gnd.n5332 gnd.n5331 585
R1636 gnd.n5330 gnd.n5329 585
R1637 gnd.n5330 gnd.n4801 585
R1638 gnd.n5328 gnd.n4803 585
R1639 gnd.n5321 gnd.n4803 585
R1640 gnd.n5308 gnd.n4804 585
R1641 gnd.n5309 gnd.n5308 585
R1642 gnd.n5278 gnd.n4817 585
R1643 gnd.n5311 gnd.n4817 585
R1644 gnd.n5277 gnd.n5276 585
R1645 gnd.n5276 gnd.n5275 585
R1646 gnd.n5273 gnd.n4834 585
R1647 gnd.n5273 gnd.n4825 585
R1648 gnd.n5272 gnd.n5271 585
R1649 gnd.n5272 gnd.n4824 585
R1650 gnd.n4836 gnd.n4835 585
R1651 gnd.n5263 gnd.n4835 585
R1652 gnd.n5232 gnd.n5231 585
R1653 gnd.n5231 gnd.n4840 585
R1654 gnd.n5233 gnd.n4850 585
R1655 gnd.n5250 gnd.n4850 585
R1656 gnd.n5230 gnd.n5229 585
R1657 gnd.n5229 gnd.n4857 585
R1658 gnd.n5228 gnd.n4864 585
R1659 gnd.n5228 gnd.n4856 585
R1660 gnd.n5227 gnd.n4866 585
R1661 gnd.n5227 gnd.n5226 585
R1662 gnd.n5206 gnd.n4865 585
R1663 gnd.n4878 gnd.n4865 585
R1664 gnd.n5205 gnd.n4876 585
R1665 gnd.n5216 gnd.n4876 585
R1666 gnd.n5196 gnd.n4883 585
R1667 gnd.n5197 gnd.n5196 585
R1668 gnd.n5195 gnd.n4889 585
R1669 gnd.n5195 gnd.n5194 585
R1670 gnd.n5180 gnd.n4888 585
R1671 gnd.n4899 gnd.n4888 585
R1672 gnd.n5179 gnd.n4897 585
R1673 gnd.n5186 gnd.n4897 585
R1674 gnd.n5178 gnd.n5177 585
R1675 gnd.n5177 gnd.n5176 585
R1676 gnd.n4371 gnd.n4370 585
R1677 gnd.n4370 gnd.n4369 585
R1678 gnd.n4372 gnd.n1153 585
R1679 gnd.n2577 gnd.n1153 585
R1680 gnd.n4374 gnd.n4373 585
R1681 gnd.n4375 gnd.n4374 585
R1682 gnd.n1138 gnd.n1137 585
R1683 gnd.n2569 gnd.n1138 585
R1684 gnd.n4383 gnd.n4382 585
R1685 gnd.n4382 gnd.n4381 585
R1686 gnd.n4384 gnd.n1132 585
R1687 gnd.n2560 gnd.n1132 585
R1688 gnd.n4386 gnd.n4385 585
R1689 gnd.n4387 gnd.n4386 585
R1690 gnd.n1116 gnd.n1115 585
R1691 gnd.n2552 gnd.n1116 585
R1692 gnd.n4395 gnd.n4394 585
R1693 gnd.n4394 gnd.n4393 585
R1694 gnd.n4396 gnd.n1110 585
R1695 gnd.n2544 gnd.n1110 585
R1696 gnd.n4398 gnd.n4397 585
R1697 gnd.n4399 gnd.n4398 585
R1698 gnd.n1095 gnd.n1094 585
R1699 gnd.n2536 gnd.n1095 585
R1700 gnd.n4407 gnd.n4406 585
R1701 gnd.n4406 gnd.n4405 585
R1702 gnd.n4408 gnd.n1089 585
R1703 gnd.n2528 gnd.n1089 585
R1704 gnd.n4410 gnd.n4409 585
R1705 gnd.n4411 gnd.n4410 585
R1706 gnd.n1073 gnd.n1072 585
R1707 gnd.n2520 gnd.n1073 585
R1708 gnd.n4419 gnd.n4418 585
R1709 gnd.n4418 gnd.n4417 585
R1710 gnd.n4420 gnd.n1070 585
R1711 gnd.n2512 gnd.n1070 585
R1712 gnd.n4423 gnd.n4422 585
R1713 gnd.n4424 gnd.n4423 585
R1714 gnd.n1071 gnd.n1056 585
R1715 gnd.n2504 gnd.n1056 585
R1716 gnd.n4432 gnd.n4431 585
R1717 gnd.n4431 gnd.n4430 585
R1718 gnd.n4433 gnd.n1053 585
R1719 gnd.n2496 gnd.n1053 585
R1720 gnd.n4436 gnd.n4435 585
R1721 gnd.n4437 gnd.n4436 585
R1722 gnd.n1054 gnd.n1034 585
R1723 gnd.n2488 gnd.n1034 585
R1724 gnd.n4445 gnd.n4444 585
R1725 gnd.n4444 gnd.n4443 585
R1726 gnd.n4446 gnd.n1032 585
R1727 gnd.n2480 gnd.n1032 585
R1728 gnd.n4448 gnd.n1028 585
R1729 gnd.n2326 gnd.n1028 585
R1730 gnd.n4450 gnd.n4449 585
R1731 gnd.n4451 gnd.n4450 585
R1732 gnd.n1012 gnd.n1011 585
R1733 gnd.n2471 gnd.n1012 585
R1734 gnd.n4459 gnd.n4458 585
R1735 gnd.n4458 gnd.n4457 585
R1736 gnd.n4460 gnd.n1006 585
R1737 gnd.n2461 gnd.n1006 585
R1738 gnd.n4462 gnd.n4461 585
R1739 gnd.n4463 gnd.n4462 585
R1740 gnd.n992 gnd.n991 585
R1741 gnd.n1002 gnd.n992 585
R1742 gnd.n4471 gnd.n4470 585
R1743 gnd.n4470 gnd.n4469 585
R1744 gnd.n4472 gnd.n986 585
R1745 gnd.n986 gnd.n985 585
R1746 gnd.n4474 gnd.n4473 585
R1747 gnd.n4475 gnd.n4474 585
R1748 gnd.n971 gnd.n970 585
R1749 gnd.n974 gnd.n971 585
R1750 gnd.n4483 gnd.n4482 585
R1751 gnd.n4482 gnd.n4481 585
R1752 gnd.n4484 gnd.n965 585
R1753 gnd.n965 gnd.n962 585
R1754 gnd.n4486 gnd.n4485 585
R1755 gnd.n4487 gnd.n4486 585
R1756 gnd.n966 gnd.n964 585
R1757 gnd.n964 gnd.n960 585
R1758 gnd.n2434 gnd.n2433 585
R1759 gnd.n2435 gnd.n2434 585
R1760 gnd.n2429 gnd.n909 585
R1761 gnd.n909 gnd.n906 585
R1762 gnd.n4572 gnd.n4571 585
R1763 gnd.n4570 gnd.n908 585
R1764 gnd.n4569 gnd.n907 585
R1765 gnd.n4574 gnd.n907 585
R1766 gnd.n4568 gnd.n4567 585
R1767 gnd.n4566 gnd.n4565 585
R1768 gnd.n4564 gnd.n4563 585
R1769 gnd.n4562 gnd.n4561 585
R1770 gnd.n4560 gnd.n4559 585
R1771 gnd.n4558 gnd.n4557 585
R1772 gnd.n4556 gnd.n4555 585
R1773 gnd.n4554 gnd.n4553 585
R1774 gnd.n4552 gnd.n4551 585
R1775 gnd.n4550 gnd.n4549 585
R1776 gnd.n4548 gnd.n4547 585
R1777 gnd.n4546 gnd.n4545 585
R1778 gnd.n4544 gnd.n4543 585
R1779 gnd.n4542 gnd.n4541 585
R1780 gnd.n4540 gnd.n4539 585
R1781 gnd.n4537 gnd.n4536 585
R1782 gnd.n4535 gnd.n4534 585
R1783 gnd.n4533 gnd.n4532 585
R1784 gnd.n4531 gnd.n4530 585
R1785 gnd.n4529 gnd.n4528 585
R1786 gnd.n4527 gnd.n4526 585
R1787 gnd.n4525 gnd.n4524 585
R1788 gnd.n4523 gnd.n4522 585
R1789 gnd.n4521 gnd.n4520 585
R1790 gnd.n4519 gnd.n4518 585
R1791 gnd.n4517 gnd.n4516 585
R1792 gnd.n4515 gnd.n4514 585
R1793 gnd.n4513 gnd.n4512 585
R1794 gnd.n4511 gnd.n4510 585
R1795 gnd.n4509 gnd.n4508 585
R1796 gnd.n4507 gnd.n4506 585
R1797 gnd.n4505 gnd.n4504 585
R1798 gnd.n4503 gnd.n4502 585
R1799 gnd.n4501 gnd.n948 585
R1800 gnd.n952 gnd.n949 585
R1801 gnd.n4497 gnd.n4496 585
R1802 gnd.n2179 gnd.n2178 585
R1803 gnd.n2585 gnd.n2584 585
R1804 gnd.n2587 gnd.n2586 585
R1805 gnd.n2589 gnd.n2588 585
R1806 gnd.n2591 gnd.n2590 585
R1807 gnd.n2593 gnd.n2592 585
R1808 gnd.n2595 gnd.n2594 585
R1809 gnd.n2597 gnd.n2596 585
R1810 gnd.n2599 gnd.n2598 585
R1811 gnd.n2601 gnd.n2600 585
R1812 gnd.n2603 gnd.n2602 585
R1813 gnd.n2605 gnd.n2604 585
R1814 gnd.n2607 gnd.n2606 585
R1815 gnd.n2609 gnd.n2608 585
R1816 gnd.n2611 gnd.n2610 585
R1817 gnd.n2613 gnd.n2612 585
R1818 gnd.n2615 gnd.n2614 585
R1819 gnd.n2617 gnd.n2616 585
R1820 gnd.n2619 gnd.n2618 585
R1821 gnd.n2622 gnd.n2621 585
R1822 gnd.n2620 gnd.n2157 585
R1823 gnd.n2835 gnd.n2834 585
R1824 gnd.n2837 gnd.n2836 585
R1825 gnd.n2839 gnd.n2838 585
R1826 gnd.n2841 gnd.n2840 585
R1827 gnd.n2843 gnd.n2842 585
R1828 gnd.n2845 gnd.n2844 585
R1829 gnd.n2847 gnd.n2846 585
R1830 gnd.n2849 gnd.n2848 585
R1831 gnd.n2851 gnd.n2850 585
R1832 gnd.n2853 gnd.n2852 585
R1833 gnd.n2855 gnd.n2854 585
R1834 gnd.n2857 gnd.n2856 585
R1835 gnd.n2858 gnd.n2138 585
R1836 gnd.n2860 gnd.n2859 585
R1837 gnd.n2139 gnd.n2137 585
R1838 gnd.n2140 gnd.n1158 585
R1839 gnd.n2862 gnd.n1158 585
R1840 gnd.n2580 gnd.n1160 585
R1841 gnd.n4369 gnd.n1160 585
R1842 gnd.n2579 gnd.n2578 585
R1843 gnd.n2578 gnd.n2577 585
R1844 gnd.n2183 gnd.n1151 585
R1845 gnd.n4375 gnd.n1151 585
R1846 gnd.n2568 gnd.n2567 585
R1847 gnd.n2569 gnd.n2568 585
R1848 gnd.n2189 gnd.n1140 585
R1849 gnd.n4381 gnd.n1140 585
R1850 gnd.n2562 gnd.n2561 585
R1851 gnd.n2561 gnd.n2560 585
R1852 gnd.n2191 gnd.n1129 585
R1853 gnd.n4387 gnd.n1129 585
R1854 gnd.n2551 gnd.n2550 585
R1855 gnd.n2552 gnd.n2551 585
R1856 gnd.n2195 gnd.n1118 585
R1857 gnd.n4393 gnd.n1118 585
R1858 gnd.n2546 gnd.n2545 585
R1859 gnd.n2545 gnd.n2544 585
R1860 gnd.n2197 gnd.n1107 585
R1861 gnd.n4399 gnd.n1107 585
R1862 gnd.n2535 gnd.n2534 585
R1863 gnd.n2536 gnd.n2535 585
R1864 gnd.n2202 gnd.n1097 585
R1865 gnd.n4405 gnd.n1097 585
R1866 gnd.n2530 gnd.n2529 585
R1867 gnd.n2529 gnd.n2528 585
R1868 gnd.n2204 gnd.n1086 585
R1869 gnd.n4411 gnd.n1086 585
R1870 gnd.n2519 gnd.n2518 585
R1871 gnd.n2520 gnd.n2519 585
R1872 gnd.n2208 gnd.n1075 585
R1873 gnd.n4417 gnd.n1075 585
R1874 gnd.n2514 gnd.n2513 585
R1875 gnd.n2513 gnd.n2512 585
R1876 gnd.n2210 gnd.n1067 585
R1877 gnd.n4424 gnd.n1067 585
R1878 gnd.n2503 gnd.n2502 585
R1879 gnd.n2504 gnd.n2503 585
R1880 gnd.n2215 gnd.n1058 585
R1881 gnd.n4430 gnd.n1058 585
R1882 gnd.n2498 gnd.n2497 585
R1883 gnd.n2497 gnd.n2496 585
R1884 gnd.n2218 gnd.n1050 585
R1885 gnd.n4437 gnd.n1050 585
R1886 gnd.n2487 gnd.n2486 585
R1887 gnd.n2488 gnd.n2487 585
R1888 gnd.n2222 gnd.n1036 585
R1889 gnd.n4443 gnd.n1036 585
R1890 gnd.n2482 gnd.n2481 585
R1891 gnd.n2481 gnd.n2480 585
R1892 gnd.n2225 gnd.n2224 585
R1893 gnd.n2326 gnd.n2225 585
R1894 gnd.n2468 gnd.n1025 585
R1895 gnd.n4451 gnd.n1025 585
R1896 gnd.n2470 gnd.n2469 585
R1897 gnd.n2471 gnd.n2470 585
R1898 gnd.n2331 gnd.n1014 585
R1899 gnd.n4457 gnd.n1014 585
R1900 gnd.n2463 gnd.n2462 585
R1901 gnd.n2462 gnd.n2461 585
R1902 gnd.n2348 gnd.n1003 585
R1903 gnd.n4463 gnd.n1003 585
R1904 gnd.n2347 gnd.n2346 585
R1905 gnd.n2346 gnd.n1002 585
R1906 gnd.n2333 gnd.n993 585
R1907 gnd.n4469 gnd.n993 585
R1908 gnd.n2342 gnd.n2341 585
R1909 gnd.n2341 gnd.n985 585
R1910 gnd.n2340 gnd.n983 585
R1911 gnd.n4475 gnd.n983 585
R1912 gnd.n2339 gnd.n2338 585
R1913 gnd.n2338 gnd.n974 585
R1914 gnd.n2335 gnd.n972 585
R1915 gnd.n4481 gnd.n972 585
R1916 gnd.n959 gnd.n957 585
R1917 gnd.n962 gnd.n959 585
R1918 gnd.n4489 gnd.n4488 585
R1919 gnd.n4488 gnd.n4487 585
R1920 gnd.n958 gnd.n955 585
R1921 gnd.n960 gnd.n958 585
R1922 gnd.n4493 gnd.n954 585
R1923 gnd.n2435 gnd.n954 585
R1924 gnd.n4495 gnd.n4494 585
R1925 gnd.n4495 gnd.n906 585
R1926 gnd.n6961 gnd.n6960 585
R1927 gnd.n6962 gnd.n6961 585
R1928 gnd.n87 gnd.n85 585
R1929 gnd.n85 gnd.n81 585
R1930 gnd.n6881 gnd.n6880 585
R1931 gnd.n6882 gnd.n6881 585
R1932 gnd.n165 gnd.n164 585
R1933 gnd.n164 gnd.n162 585
R1934 gnd.n6876 gnd.n6875 585
R1935 gnd.n6875 gnd.n6874 585
R1936 gnd.n168 gnd.n167 585
R1937 gnd.n170 gnd.n168 585
R1938 gnd.n6791 gnd.n6790 585
R1939 gnd.n6792 gnd.n6791 585
R1940 gnd.n181 gnd.n180 585
R1941 gnd.n188 gnd.n180 585
R1942 gnd.n6786 gnd.n6785 585
R1943 gnd.n6785 gnd.n6784 585
R1944 gnd.n184 gnd.n183 585
R1945 gnd.n186 gnd.n184 585
R1946 gnd.n6775 gnd.n6774 585
R1947 gnd.n6776 gnd.n6775 585
R1948 gnd.n197 gnd.n196 585
R1949 gnd.n196 gnd.n194 585
R1950 gnd.n6770 gnd.n6769 585
R1951 gnd.n6769 gnd.n6768 585
R1952 gnd.n200 gnd.n199 585
R1953 gnd.n268 gnd.n200 585
R1954 gnd.n6759 gnd.n6758 585
R1955 gnd.n6760 gnd.n6759 585
R1956 gnd.n211 gnd.n210 585
R1957 gnd.n6728 gnd.n210 585
R1958 gnd.n6754 gnd.n6753 585
R1959 gnd.n6753 gnd.n6752 585
R1960 gnd.n220 gnd.n219 585
R1961 gnd.n6733 gnd.n220 585
R1962 gnd.n6743 gnd.n6742 585
R1963 gnd.n6744 gnd.n6743 585
R1964 gnd.n6741 gnd.n6740 585
R1965 gnd.n6740 gnd.n6739 585
R1966 gnd.n4096 gnd.n232 585
R1967 gnd.n4115 gnd.n232 585
R1968 gnd.n4098 gnd.n4097 585
R1969 gnd.n4099 gnd.n4098 585
R1970 gnd.n4095 gnd.n4094 585
R1971 gnd.n4095 gnd.n1402 585
R1972 gnd.n4093 gnd.n4092 585
R1973 gnd.n4092 gnd.n4091 585
R1974 gnd.n4079 gnd.n1405 585
R1975 gnd.n4071 gnd.n1405 585
R1976 gnd.n4081 gnd.n4080 585
R1977 gnd.n4082 gnd.n4081 585
R1978 gnd.n4078 gnd.n1419 585
R1979 gnd.n4078 gnd.n4077 585
R1980 gnd.n4047 gnd.n1418 585
R1981 gnd.n4059 gnd.n1418 585
R1982 gnd.n4048 gnd.n1448 585
R1983 gnd.n1448 gnd.n1437 585
R1984 gnd.n4050 gnd.n4049 585
R1985 gnd.n4051 gnd.n4050 585
R1986 gnd.n1449 gnd.n1447 585
R1987 gnd.n3936 gnd.n1447 585
R1988 gnd.n4042 gnd.n4041 585
R1989 gnd.n4041 gnd.n4040 585
R1990 gnd.n1452 gnd.n1451 585
R1991 gnd.n4025 gnd.n1452 585
R1992 gnd.n4013 gnd.n1473 585
R1993 gnd.n3942 gnd.n1473 585
R1994 gnd.n4015 gnd.n4014 585
R1995 gnd.n4016 gnd.n4015 585
R1996 gnd.n1474 gnd.n1472 585
R1997 gnd.n3946 gnd.n1472 585
R1998 gnd.n4008 gnd.n4007 585
R1999 gnd.n4007 gnd.n4006 585
R2000 gnd.n1477 gnd.n1476 585
R2001 gnd.n3994 gnd.n1477 585
R2002 gnd.n3981 gnd.n1499 585
R2003 gnd.n1499 gnd.n1487 585
R2004 gnd.n3983 gnd.n3982 585
R2005 gnd.n3984 gnd.n3983 585
R2006 gnd.n1500 gnd.n1498 585
R2007 gnd.n3956 gnd.n1498 585
R2008 gnd.n3976 gnd.n3975 585
R2009 gnd.n3975 gnd.n3974 585
R2010 gnd.n1502 gnd.n1314 585
R2011 gnd.n4153 gnd.n1314 585
R2012 gnd.n4227 gnd.n4226 585
R2013 gnd.n4225 gnd.n1313 585
R2014 gnd.n4224 gnd.n1312 585
R2015 gnd.n4229 gnd.n1312 585
R2016 gnd.n4223 gnd.n4222 585
R2017 gnd.n4221 gnd.n4220 585
R2018 gnd.n4219 gnd.n4218 585
R2019 gnd.n4217 gnd.n4216 585
R2020 gnd.n4215 gnd.n4214 585
R2021 gnd.n4213 gnd.n4212 585
R2022 gnd.n4211 gnd.n4210 585
R2023 gnd.n4209 gnd.n4208 585
R2024 gnd.n4207 gnd.n4206 585
R2025 gnd.n4205 gnd.n4204 585
R2026 gnd.n4203 gnd.n4202 585
R2027 gnd.n4201 gnd.n4200 585
R2028 gnd.n4199 gnd.n4198 585
R2029 gnd.n4196 gnd.n4195 585
R2030 gnd.n4194 gnd.n4193 585
R2031 gnd.n4192 gnd.n4191 585
R2032 gnd.n4190 gnd.n4189 585
R2033 gnd.n4188 gnd.n4187 585
R2034 gnd.n4186 gnd.n4185 585
R2035 gnd.n4184 gnd.n4183 585
R2036 gnd.n4182 gnd.n4181 585
R2037 gnd.n4180 gnd.n4179 585
R2038 gnd.n4178 gnd.n4177 585
R2039 gnd.n4176 gnd.n4175 585
R2040 gnd.n4174 gnd.n4173 585
R2041 gnd.n4172 gnd.n4171 585
R2042 gnd.n4170 gnd.n4169 585
R2043 gnd.n4168 gnd.n4167 585
R2044 gnd.n4166 gnd.n4165 585
R2045 gnd.n4164 gnd.n4163 585
R2046 gnd.n4162 gnd.n4161 585
R2047 gnd.n4160 gnd.n1354 585
R2048 gnd.n1358 gnd.n1355 585
R2049 gnd.n4156 gnd.n4155 585
R2050 gnd.n156 gnd.n155 585
R2051 gnd.n6890 gnd.n151 585
R2052 gnd.n6892 gnd.n6891 585
R2053 gnd.n6894 gnd.n149 585
R2054 gnd.n6896 gnd.n6895 585
R2055 gnd.n6897 gnd.n144 585
R2056 gnd.n6899 gnd.n6898 585
R2057 gnd.n6901 gnd.n142 585
R2058 gnd.n6903 gnd.n6902 585
R2059 gnd.n6904 gnd.n137 585
R2060 gnd.n6906 gnd.n6905 585
R2061 gnd.n6908 gnd.n135 585
R2062 gnd.n6910 gnd.n6909 585
R2063 gnd.n6911 gnd.n130 585
R2064 gnd.n6913 gnd.n6912 585
R2065 gnd.n6915 gnd.n128 585
R2066 gnd.n6917 gnd.n6916 585
R2067 gnd.n6918 gnd.n123 585
R2068 gnd.n6920 gnd.n6919 585
R2069 gnd.n6922 gnd.n121 585
R2070 gnd.n6924 gnd.n6923 585
R2071 gnd.n6928 gnd.n116 585
R2072 gnd.n6930 gnd.n6929 585
R2073 gnd.n6932 gnd.n114 585
R2074 gnd.n6934 gnd.n6933 585
R2075 gnd.n6935 gnd.n109 585
R2076 gnd.n6937 gnd.n6936 585
R2077 gnd.n6939 gnd.n107 585
R2078 gnd.n6941 gnd.n6940 585
R2079 gnd.n6942 gnd.n102 585
R2080 gnd.n6944 gnd.n6943 585
R2081 gnd.n6946 gnd.n100 585
R2082 gnd.n6948 gnd.n6947 585
R2083 gnd.n6949 gnd.n95 585
R2084 gnd.n6951 gnd.n6950 585
R2085 gnd.n6953 gnd.n92 585
R2086 gnd.n6955 gnd.n6954 585
R2087 gnd.n6956 gnd.n90 585
R2088 gnd.n6957 gnd.n86 585
R2089 gnd.n94 gnd.n86 585
R2090 gnd.n6886 gnd.n82 585
R2091 gnd.n6962 gnd.n82 585
R2092 gnd.n6885 gnd.n6884 585
R2093 gnd.n6884 gnd.n81 585
R2094 gnd.n6883 gnd.n160 585
R2095 gnd.n6883 gnd.n6882 585
R2096 gnd.n253 gnd.n161 585
R2097 gnd.n162 gnd.n161 585
R2098 gnd.n254 gnd.n171 585
R2099 gnd.n6874 gnd.n171 585
R2100 gnd.n256 gnd.n255 585
R2101 gnd.n255 gnd.n170 585
R2102 gnd.n257 gnd.n179 585
R2103 gnd.n6792 gnd.n179 585
R2104 gnd.n259 gnd.n258 585
R2105 gnd.n258 gnd.n188 585
R2106 gnd.n260 gnd.n187 585
R2107 gnd.n6784 gnd.n187 585
R2108 gnd.n262 gnd.n261 585
R2109 gnd.n261 gnd.n186 585
R2110 gnd.n263 gnd.n195 585
R2111 gnd.n6776 gnd.n195 585
R2112 gnd.n265 gnd.n264 585
R2113 gnd.n264 gnd.n194 585
R2114 gnd.n266 gnd.n202 585
R2115 gnd.n6768 gnd.n202 585
R2116 gnd.n270 gnd.n269 585
R2117 gnd.n269 gnd.n268 585
R2118 gnd.n271 gnd.n208 585
R2119 gnd.n6760 gnd.n208 585
R2120 gnd.n6730 gnd.n6729 585
R2121 gnd.n6729 gnd.n6728 585
R2122 gnd.n6731 gnd.n222 585
R2123 gnd.n6752 gnd.n222 585
R2124 gnd.n6735 gnd.n6734 585
R2125 gnd.n6734 gnd.n6733 585
R2126 gnd.n6736 gnd.n230 585
R2127 gnd.n6744 gnd.n230 585
R2128 gnd.n6738 gnd.n6737 585
R2129 gnd.n6739 gnd.n6738 585
R2130 gnd.n234 gnd.n233 585
R2131 gnd.n4115 gnd.n233 585
R2132 gnd.n1428 gnd.n1403 585
R2133 gnd.n4099 gnd.n1403 585
R2134 gnd.n1430 gnd.n1429 585
R2135 gnd.n1429 gnd.n1402 585
R2136 gnd.n1431 gnd.n1407 585
R2137 gnd.n4091 gnd.n1407 585
R2138 gnd.n4073 gnd.n4072 585
R2139 gnd.n4072 gnd.n4071 585
R2140 gnd.n4074 gnd.n1416 585
R2141 gnd.n4082 gnd.n1416 585
R2142 gnd.n4076 gnd.n4075 585
R2143 gnd.n4077 gnd.n4076 585
R2144 gnd.n1422 gnd.n1421 585
R2145 gnd.n4059 gnd.n1421 585
R2146 gnd.n3934 gnd.n3933 585
R2147 gnd.n3933 gnd.n1437 585
R2148 gnd.n3935 gnd.n1444 585
R2149 gnd.n4051 gnd.n1444 585
R2150 gnd.n3938 gnd.n3937 585
R2151 gnd.n3937 gnd.n3936 585
R2152 gnd.n3939 gnd.n1454 585
R2153 gnd.n4040 gnd.n1454 585
R2154 gnd.n3940 gnd.n1462 585
R2155 gnd.n4025 gnd.n1462 585
R2156 gnd.n3944 gnd.n3943 585
R2157 gnd.n3943 gnd.n3942 585
R2158 gnd.n3945 gnd.n1470 585
R2159 gnd.n4016 gnd.n1470 585
R2160 gnd.n3948 gnd.n3947 585
R2161 gnd.n3947 gnd.n3946 585
R2162 gnd.n3949 gnd.n1479 585
R2163 gnd.n4006 gnd.n1479 585
R2164 gnd.n3950 gnd.n1488 585
R2165 gnd.n3994 gnd.n1488 585
R2166 gnd.n3952 gnd.n3951 585
R2167 gnd.n3951 gnd.n1487 585
R2168 gnd.n3953 gnd.n1496 585
R2169 gnd.n3984 gnd.n1496 585
R2170 gnd.n3955 gnd.n3954 585
R2171 gnd.n3956 gnd.n3955 585
R2172 gnd.n3917 gnd.n1360 585
R2173 gnd.n3974 gnd.n1360 585
R2174 gnd.n4154 gnd.n1361 585
R2175 gnd.n4154 gnd.n4153 585
R2176 gnd.n3718 gnd.n3717 585
R2177 gnd.n3717 gnd.n3716 585
R2178 gnd.n3719 gnd.n3517 585
R2179 gnd.n3517 gnd.n1650 585
R2180 gnd.n3721 gnd.n3720 585
R2181 gnd.n3722 gnd.n3721 585
R2182 gnd.n3519 gnd.n3516 585
R2183 gnd.n3516 gnd.n1658 585
R2184 gnd.n3518 gnd.n3507 585
R2185 gnd.n3507 gnd.n1657 585
R2186 gnd.n3730 gnd.n3506 585
R2187 gnd.n3730 gnd.n3729 585
R2188 gnd.n3732 gnd.n3731 585
R2189 gnd.n3731 gnd.n1665 585
R2190 gnd.n3733 gnd.n3503 585
R2191 gnd.n3503 gnd.n1664 585
R2192 gnd.n3735 gnd.n3734 585
R2193 gnd.n3736 gnd.n3735 585
R2194 gnd.n3505 gnd.n3502 585
R2195 gnd.n3502 gnd.n1672 585
R2196 gnd.n3504 gnd.n3495 585
R2197 gnd.n3495 gnd.n1671 585
R2198 gnd.n3746 gnd.n3494 585
R2199 gnd.n3746 gnd.n3745 585
R2200 gnd.n3748 gnd.n3747 585
R2201 gnd.n3747 gnd.n1679 585
R2202 gnd.n3749 gnd.n3491 585
R2203 gnd.n3491 gnd.n1678 585
R2204 gnd.n3751 gnd.n3750 585
R2205 gnd.n3752 gnd.n3751 585
R2206 gnd.n3493 gnd.n3490 585
R2207 gnd.n3490 gnd.n1685 585
R2208 gnd.n3492 gnd.n3479 585
R2209 gnd.n3758 gnd.n3479 585
R2210 gnd.n3761 gnd.n3478 585
R2211 gnd.n3761 gnd.n3760 585
R2212 gnd.n3763 gnd.n3762 585
R2213 gnd.n3762 gnd.n1692 585
R2214 gnd.n3764 gnd.n3475 585
R2215 gnd.n3475 gnd.n1691 585
R2216 gnd.n3766 gnd.n3765 585
R2217 gnd.n3767 gnd.n3766 585
R2218 gnd.n3477 gnd.n3474 585
R2219 gnd.n3474 gnd.n1699 585
R2220 gnd.n3476 gnd.n3466 585
R2221 gnd.n3466 gnd.n1698 585
R2222 gnd.n3776 gnd.n3465 585
R2223 gnd.n3776 gnd.n3775 585
R2224 gnd.n3778 gnd.n3777 585
R2225 gnd.n3777 gnd.n1705 585
R2226 gnd.n3779 gnd.n1730 585
R2227 gnd.n1730 gnd.n1729 585
R2228 gnd.n3781 gnd.n3780 585
R2229 gnd.n3782 gnd.n3781 585
R2230 gnd.n3464 gnd.n1728 585
R2231 gnd.n1728 gnd.n1712 585
R2232 gnd.n3463 gnd.n3462 585
R2233 gnd.n3462 gnd.n1711 585
R2234 gnd.n3461 gnd.n3457 585
R2235 gnd.n3461 gnd.n3460 585
R2236 gnd.n3456 gnd.n1719 585
R2237 gnd.n3790 gnd.n1719 585
R2238 gnd.n3455 gnd.n3454 585
R2239 gnd.n3454 gnd.n1718 585
R2240 gnd.n3453 gnd.n1731 585
R2241 gnd.n3453 gnd.n3452 585
R2242 gnd.n3321 gnd.n1732 585
R2243 gnd.n3331 gnd.n1732 585
R2244 gnd.n3322 gnd.n3320 585
R2245 gnd.n3320 gnd.n1743 585
R2246 gnd.n3324 gnd.n3323 585
R2247 gnd.n3324 gnd.n1741 585
R2248 gnd.n3325 gnd.n3319 585
R2249 gnd.n3339 gnd.n3325 585
R2250 gnd.n3342 gnd.n3341 585
R2251 gnd.n3341 gnd.n3340 585
R2252 gnd.n3343 gnd.n3316 585
R2253 gnd.n3316 gnd.n1750 585
R2254 gnd.n3345 gnd.n3344 585
R2255 gnd.n3346 gnd.n3345 585
R2256 gnd.n3318 gnd.n3315 585
R2257 gnd.n3315 gnd.n1757 585
R2258 gnd.n3317 gnd.n3305 585
R2259 gnd.n3352 gnd.n3305 585
R2260 gnd.n3355 gnd.n3304 585
R2261 gnd.n3355 gnd.n3354 585
R2262 gnd.n3357 gnd.n3356 585
R2263 gnd.n3356 gnd.n1764 585
R2264 gnd.n3358 gnd.n3301 585
R2265 gnd.n3301 gnd.n1763 585
R2266 gnd.n3360 gnd.n3359 585
R2267 gnd.n3361 gnd.n3360 585
R2268 gnd.n3303 gnd.n3300 585
R2269 gnd.n3300 gnd.n1772 585
R2270 gnd.n3302 gnd.n3292 585
R2271 gnd.n3292 gnd.n1770 585
R2272 gnd.n3370 gnd.n3291 585
R2273 gnd.n3370 gnd.n3369 585
R2274 gnd.n3372 gnd.n3371 585
R2275 gnd.n3371 gnd.n1779 585
R2276 gnd.n3373 gnd.n1806 585
R2277 gnd.n1806 gnd.n1778 585
R2278 gnd.n3375 gnd.n3374 585
R2279 gnd.n3376 gnd.n3375 585
R2280 gnd.n3290 gnd.n1805 585
R2281 gnd.n1805 gnd.n1787 585
R2282 gnd.n3289 gnd.n3288 585
R2283 gnd.n3288 gnd.n1785 585
R2284 gnd.n3287 gnd.n3286 585
R2285 gnd.n3287 gnd.n1796 585
R2286 gnd.n3285 gnd.n1794 585
R2287 gnd.n3384 gnd.n1794 585
R2288 gnd.n3284 gnd.n3283 585
R2289 gnd.n3283 gnd.n1793 585
R2290 gnd.n3282 gnd.n1807 585
R2291 gnd.n3282 gnd.n3281 585
R2292 gnd.n3150 gnd.n1808 585
R2293 gnd.n3160 gnd.n1808 585
R2294 gnd.n3151 gnd.n3149 585
R2295 gnd.n3149 gnd.n1819 585
R2296 gnd.n3153 gnd.n3152 585
R2297 gnd.n3153 gnd.n1818 585
R2298 gnd.n3154 gnd.n3148 585
R2299 gnd.n3168 gnd.n3154 585
R2300 gnd.n3171 gnd.n3170 585
R2301 gnd.n3170 gnd.n3169 585
R2302 gnd.n3172 gnd.n3145 585
R2303 gnd.n3145 gnd.n1826 585
R2304 gnd.n3174 gnd.n3173 585
R2305 gnd.n3175 gnd.n3174 585
R2306 gnd.n3147 gnd.n3144 585
R2307 gnd.n3144 gnd.n3141 585
R2308 gnd.n3146 gnd.n3133 585
R2309 gnd.n3181 gnd.n3133 585
R2310 gnd.n3184 gnd.n3132 585
R2311 gnd.n3184 gnd.n3183 585
R2312 gnd.n3186 gnd.n3185 585
R2313 gnd.n3185 gnd.n1838 585
R2314 gnd.n3187 gnd.n3129 585
R2315 gnd.n3129 gnd.n1837 585
R2316 gnd.n3189 gnd.n3188 585
R2317 gnd.n3190 gnd.n3189 585
R2318 gnd.n3131 gnd.n3128 585
R2319 gnd.n3128 gnd.n1844 585
R2320 gnd.n3130 gnd.n3117 585
R2321 gnd.n3196 gnd.n3117 585
R2322 gnd.n3199 gnd.n3116 585
R2323 gnd.n3199 gnd.n3198 585
R2324 gnd.n3201 gnd.n3200 585
R2325 gnd.n3200 gnd.n1851 585
R2326 gnd.n3202 gnd.n1877 585
R2327 gnd.n1877 gnd.n1850 585
R2328 gnd.n3204 gnd.n3203 585
R2329 gnd.n3205 gnd.n3204 585
R2330 gnd.n3115 gnd.n1876 585
R2331 gnd.n1876 gnd.n1858 585
R2332 gnd.n3114 gnd.n3113 585
R2333 gnd.n3113 gnd.n1857 585
R2334 gnd.n3112 gnd.n3111 585
R2335 gnd.n3112 gnd.n1866 585
R2336 gnd.n3110 gnd.n1864 585
R2337 gnd.n3213 gnd.n1864 585
R2338 gnd.n3109 gnd.n3108 585
R2339 gnd.n3108 gnd.n3107 585
R2340 gnd.n1879 gnd.n1878 585
R2341 gnd.n1880 gnd.n1879 585
R2342 gnd.n2986 gnd.n2985 585
R2343 gnd.n2987 gnd.n2986 585
R2344 gnd.n2984 gnd.n2982 585
R2345 gnd.n2982 gnd.n1889 585
R2346 gnd.n2983 gnd.n2974 585
R2347 gnd.n2974 gnd.n1888 585
R2348 gnd.n2996 gnd.n2973 585
R2349 gnd.n2996 gnd.n2995 585
R2350 gnd.n2998 gnd.n2997 585
R2351 gnd.n2997 gnd.n1898 585
R2352 gnd.n2999 gnd.n2970 585
R2353 gnd.n2970 gnd.n1896 585
R2354 gnd.n3001 gnd.n3000 585
R2355 gnd.n3002 gnd.n3001 585
R2356 gnd.n2972 gnd.n2969 585
R2357 gnd.n2969 gnd.n1904 585
R2358 gnd.n2971 gnd.n2959 585
R2359 gnd.n3008 gnd.n2959 585
R2360 gnd.n3011 gnd.n2958 585
R2361 gnd.n3011 gnd.n3010 585
R2362 gnd.n3013 gnd.n3012 585
R2363 gnd.n3012 gnd.n1912 585
R2364 gnd.n3014 gnd.n2955 585
R2365 gnd.n2955 gnd.n1910 585
R2366 gnd.n3016 gnd.n3015 585
R2367 gnd.n3017 gnd.n3016 585
R2368 gnd.n2957 gnd.n2954 585
R2369 gnd.n2954 gnd.n1919 585
R2370 gnd.n2956 gnd.n2946 585
R2371 gnd.n2946 gnd.n1918 585
R2372 gnd.n3026 gnd.n2945 585
R2373 gnd.n3026 gnd.n3025 585
R2374 gnd.n3028 gnd.n3027 585
R2375 gnd.n3027 gnd.n1926 585
R2376 gnd.n3029 gnd.n1953 585
R2377 gnd.n1953 gnd.n1952 585
R2378 gnd.n3031 gnd.n3030 585
R2379 gnd.n3032 gnd.n3031 585
R2380 gnd.n2944 gnd.n1950 585
R2381 gnd.n1950 gnd.n1933 585
R2382 gnd.n2943 gnd.n2942 585
R2383 gnd.n2942 gnd.n1932 585
R2384 gnd.n2941 gnd.n2940 585
R2385 gnd.n2941 gnd.n1942 585
R2386 gnd.n2939 gnd.n1939 585
R2387 gnd.n3040 gnd.n1939 585
R2388 gnd.n2938 gnd.n2937 585
R2389 gnd.n2937 gnd.n2936 585
R2390 gnd.n1955 gnd.n1954 585
R2391 gnd.n1956 gnd.n1955 585
R2392 gnd.n2756 gnd.n2755 585
R2393 gnd.n2757 gnd.n2756 585
R2394 gnd.n2754 gnd.n2648 585
R2395 gnd.n2648 gnd.n1964 585
R2396 gnd.n2753 gnd.n2752 585
R2397 gnd.n2752 gnd.n1963 585
R2398 gnd.n2751 gnd.n2750 585
R2399 gnd.n2749 gnd.n2748 585
R2400 gnd.n2747 gnd.n2671 585
R2401 gnd.n2747 gnd.n1973 585
R2402 gnd.n2746 gnd.n2745 585
R2403 gnd.n2744 gnd.n2743 585
R2404 gnd.n2742 gnd.n2673 585
R2405 gnd.n2740 gnd.n2739 585
R2406 gnd.n2738 gnd.n2674 585
R2407 gnd.n2737 gnd.n2736 585
R2408 gnd.n2734 gnd.n2675 585
R2409 gnd.n2732 gnd.n2731 585
R2410 gnd.n2730 gnd.n2676 585
R2411 gnd.n2729 gnd.n2728 585
R2412 gnd.n2726 gnd.n2677 585
R2413 gnd.n2724 gnd.n2723 585
R2414 gnd.n2722 gnd.n2678 585
R2415 gnd.n2721 gnd.n2720 585
R2416 gnd.n2718 gnd.n2679 585
R2417 gnd.n2716 gnd.n2715 585
R2418 gnd.n2714 gnd.n2680 585
R2419 gnd.n2713 gnd.n2712 585
R2420 gnd.n2710 gnd.n2681 585
R2421 gnd.n2708 gnd.n2707 585
R2422 gnd.n2706 gnd.n2682 585
R2423 gnd.n2705 gnd.n2704 585
R2424 gnd.n2702 gnd.n2683 585
R2425 gnd.n2700 gnd.n2699 585
R2426 gnd.n2698 gnd.n2684 585
R2427 gnd.n2697 gnd.n2696 585
R2428 gnd.n2694 gnd.n2693 585
R2429 gnd.n2692 gnd.n2691 585
R2430 gnd.n2690 gnd.n2627 585
R2431 gnd.n2832 gnd.n2831 585
R2432 gnd.n2829 gnd.n2626 585
R2433 gnd.n2827 gnd.n2826 585
R2434 gnd.n2825 gnd.n2629 585
R2435 gnd.n2823 gnd.n2822 585
R2436 gnd.n2820 gnd.n2632 585
R2437 gnd.n2818 gnd.n2817 585
R2438 gnd.n2816 gnd.n2633 585
R2439 gnd.n2815 gnd.n2814 585
R2440 gnd.n2812 gnd.n2634 585
R2441 gnd.n2810 gnd.n2809 585
R2442 gnd.n2808 gnd.n2635 585
R2443 gnd.n2807 gnd.n2806 585
R2444 gnd.n2804 gnd.n2636 585
R2445 gnd.n2802 gnd.n2801 585
R2446 gnd.n2800 gnd.n2637 585
R2447 gnd.n2799 gnd.n2798 585
R2448 gnd.n2796 gnd.n2638 585
R2449 gnd.n2794 gnd.n2793 585
R2450 gnd.n2792 gnd.n2639 585
R2451 gnd.n2791 gnd.n2790 585
R2452 gnd.n2788 gnd.n2640 585
R2453 gnd.n2786 gnd.n2785 585
R2454 gnd.n2784 gnd.n2641 585
R2455 gnd.n2783 gnd.n2782 585
R2456 gnd.n2780 gnd.n2642 585
R2457 gnd.n2778 gnd.n2777 585
R2458 gnd.n2776 gnd.n2643 585
R2459 gnd.n2775 gnd.n2774 585
R2460 gnd.n2772 gnd.n2644 585
R2461 gnd.n2770 gnd.n2769 585
R2462 gnd.n2768 gnd.n2645 585
R2463 gnd.n2767 gnd.n2766 585
R2464 gnd.n3649 gnd.n3648 585
R2465 gnd.n3651 gnd.n3650 585
R2466 gnd.n3653 gnd.n3652 585
R2467 gnd.n3655 gnd.n3654 585
R2468 gnd.n3657 gnd.n3656 585
R2469 gnd.n3659 gnd.n3658 585
R2470 gnd.n3661 gnd.n3660 585
R2471 gnd.n3663 gnd.n3662 585
R2472 gnd.n3665 gnd.n3664 585
R2473 gnd.n3667 gnd.n3666 585
R2474 gnd.n3669 gnd.n3668 585
R2475 gnd.n3671 gnd.n3670 585
R2476 gnd.n3673 gnd.n3672 585
R2477 gnd.n3675 gnd.n3674 585
R2478 gnd.n3677 gnd.n3676 585
R2479 gnd.n3679 gnd.n3678 585
R2480 gnd.n3681 gnd.n3680 585
R2481 gnd.n3683 gnd.n3682 585
R2482 gnd.n3685 gnd.n3684 585
R2483 gnd.n3687 gnd.n3686 585
R2484 gnd.n3689 gnd.n3688 585
R2485 gnd.n3691 gnd.n3690 585
R2486 gnd.n3693 gnd.n3692 585
R2487 gnd.n3695 gnd.n3694 585
R2488 gnd.n3697 gnd.n3696 585
R2489 gnd.n3699 gnd.n3698 585
R2490 gnd.n3701 gnd.n3700 585
R2491 gnd.n3703 gnd.n3702 585
R2492 gnd.n3705 gnd.n3704 585
R2493 gnd.n3708 gnd.n3707 585
R2494 gnd.n3710 gnd.n3709 585
R2495 gnd.n3712 gnd.n3711 585
R2496 gnd.n3714 gnd.n3713 585
R2497 gnd.n3625 gnd.n1331 585
R2498 gnd.n3624 gnd.n3623 585
R2499 gnd.n3622 gnd.n3621 585
R2500 gnd.n3620 gnd.n3619 585
R2501 gnd.n3617 gnd.n3616 585
R2502 gnd.n3615 gnd.n3614 585
R2503 gnd.n3613 gnd.n3612 585
R2504 gnd.n3611 gnd.n3610 585
R2505 gnd.n3609 gnd.n3608 585
R2506 gnd.n3607 gnd.n3606 585
R2507 gnd.n3605 gnd.n3604 585
R2508 gnd.n3603 gnd.n3602 585
R2509 gnd.n3601 gnd.n3600 585
R2510 gnd.n3599 gnd.n3598 585
R2511 gnd.n3597 gnd.n3596 585
R2512 gnd.n3595 gnd.n3594 585
R2513 gnd.n3593 gnd.n3592 585
R2514 gnd.n3591 gnd.n3590 585
R2515 gnd.n3589 gnd.n3588 585
R2516 gnd.n3587 gnd.n3586 585
R2517 gnd.n3585 gnd.n3584 585
R2518 gnd.n3583 gnd.n3582 585
R2519 gnd.n3581 gnd.n3580 585
R2520 gnd.n3579 gnd.n3578 585
R2521 gnd.n3577 gnd.n3576 585
R2522 gnd.n3575 gnd.n3574 585
R2523 gnd.n3573 gnd.n3572 585
R2524 gnd.n3571 gnd.n3570 585
R2525 gnd.n3569 gnd.n3568 585
R2526 gnd.n3567 gnd.n3566 585
R2527 gnd.n3565 gnd.n3564 585
R2528 gnd.n3563 gnd.n3562 585
R2529 gnd.n3561 gnd.n3540 585
R2530 gnd.n3647 gnd.n3541 585
R2531 gnd.n3716 gnd.n3541 585
R2532 gnd.n3646 gnd.n3514 585
R2533 gnd.n3514 gnd.n1650 585
R2534 gnd.n3723 gnd.n3513 585
R2535 gnd.n3723 gnd.n3722 585
R2536 gnd.n3725 gnd.n3724 585
R2537 gnd.n3724 gnd.n1658 585
R2538 gnd.n3726 gnd.n3510 585
R2539 gnd.n3510 gnd.n1657 585
R2540 gnd.n3728 gnd.n3727 585
R2541 gnd.n3729 gnd.n3728 585
R2542 gnd.n3512 gnd.n3509 585
R2543 gnd.n3509 gnd.n1665 585
R2544 gnd.n3511 gnd.n3500 585
R2545 gnd.n3500 gnd.n1664 585
R2546 gnd.n3737 gnd.n3499 585
R2547 gnd.n3737 gnd.n3736 585
R2548 gnd.n3739 gnd.n3738 585
R2549 gnd.n3738 gnd.n1672 585
R2550 gnd.n3740 gnd.n3497 585
R2551 gnd.n3497 gnd.n1671 585
R2552 gnd.n3742 gnd.n3741 585
R2553 gnd.n3745 gnd.n3742 585
R2554 gnd.n3498 gnd.n3496 585
R2555 gnd.n3496 gnd.n1679 585
R2556 gnd.n3488 gnd.n3487 585
R2557 gnd.n3488 gnd.n1678 585
R2558 gnd.n3754 gnd.n3753 585
R2559 gnd.n3753 gnd.n3752 585
R2560 gnd.n3755 gnd.n3482 585
R2561 gnd.n3482 gnd.n1685 585
R2562 gnd.n3757 gnd.n3756 585
R2563 gnd.n3758 gnd.n3757 585
R2564 gnd.n3486 gnd.n3480 585
R2565 gnd.n3760 gnd.n3480 585
R2566 gnd.n3485 gnd.n3484 585
R2567 gnd.n3484 gnd.n1692 585
R2568 gnd.n3483 gnd.n3472 585
R2569 gnd.n3472 gnd.n1691 585
R2570 gnd.n3768 gnd.n3471 585
R2571 gnd.n3768 gnd.n3767 585
R2572 gnd.n3770 gnd.n3769 585
R2573 gnd.n3769 gnd.n1699 585
R2574 gnd.n3771 gnd.n3468 585
R2575 gnd.n3468 gnd.n1698 585
R2576 gnd.n3773 gnd.n3772 585
R2577 gnd.n3775 gnd.n3773 585
R2578 gnd.n3470 gnd.n3467 585
R2579 gnd.n3467 gnd.n1705 585
R2580 gnd.n3469 gnd.n1725 585
R2581 gnd.n1729 gnd.n1725 585
R2582 gnd.n3783 gnd.n1726 585
R2583 gnd.n3783 gnd.n3782 585
R2584 gnd.n3784 gnd.n1724 585
R2585 gnd.n3784 gnd.n1712 585
R2586 gnd.n3786 gnd.n3785 585
R2587 gnd.n3785 gnd.n1711 585
R2588 gnd.n3787 gnd.n1722 585
R2589 gnd.n3460 gnd.n1722 585
R2590 gnd.n3789 gnd.n3788 585
R2591 gnd.n3790 gnd.n3789 585
R2592 gnd.n1723 gnd.n1721 585
R2593 gnd.n1721 gnd.n1718 585
R2594 gnd.n3329 gnd.n1734 585
R2595 gnd.n3452 gnd.n1734 585
R2596 gnd.n3332 gnd.n3330 585
R2597 gnd.n3332 gnd.n3331 585
R2598 gnd.n3334 gnd.n3333 585
R2599 gnd.n3333 gnd.n1743 585
R2600 gnd.n3335 gnd.n3327 585
R2601 gnd.n3327 gnd.n1741 585
R2602 gnd.n3337 gnd.n3336 585
R2603 gnd.n3339 gnd.n3337 585
R2604 gnd.n3328 gnd.n3326 585
R2605 gnd.n3340 gnd.n3326 585
R2606 gnd.n3313 gnd.n3312 585
R2607 gnd.n3313 gnd.n1750 585
R2608 gnd.n3348 gnd.n3347 585
R2609 gnd.n3347 gnd.n3346 585
R2610 gnd.n3349 gnd.n3307 585
R2611 gnd.n3307 gnd.n1757 585
R2612 gnd.n3351 gnd.n3350 585
R2613 gnd.n3352 gnd.n3351 585
R2614 gnd.n3311 gnd.n3306 585
R2615 gnd.n3354 gnd.n3306 585
R2616 gnd.n3310 gnd.n3309 585
R2617 gnd.n3309 gnd.n1764 585
R2618 gnd.n3308 gnd.n3298 585
R2619 gnd.n3298 gnd.n1763 585
R2620 gnd.n3362 gnd.n3297 585
R2621 gnd.n3362 gnd.n3361 585
R2622 gnd.n3364 gnd.n3363 585
R2623 gnd.n3363 gnd.n1772 585
R2624 gnd.n3365 gnd.n3294 585
R2625 gnd.n3294 gnd.n1770 585
R2626 gnd.n3367 gnd.n3366 585
R2627 gnd.n3369 gnd.n3367 585
R2628 gnd.n3296 gnd.n3293 585
R2629 gnd.n3293 gnd.n1779 585
R2630 gnd.n3295 gnd.n1802 585
R2631 gnd.n1802 gnd.n1778 585
R2632 gnd.n3377 gnd.n1803 585
R2633 gnd.n3377 gnd.n3376 585
R2634 gnd.n3378 gnd.n1801 585
R2635 gnd.n3378 gnd.n1787 585
R2636 gnd.n3380 gnd.n3379 585
R2637 gnd.n3379 gnd.n1785 585
R2638 gnd.n3381 gnd.n1799 585
R2639 gnd.n1799 gnd.n1796 585
R2640 gnd.n3383 gnd.n3382 585
R2641 gnd.n3384 gnd.n3383 585
R2642 gnd.n1800 gnd.n1798 585
R2643 gnd.n1798 gnd.n1793 585
R2644 gnd.n3158 gnd.n1811 585
R2645 gnd.n3281 gnd.n1811 585
R2646 gnd.n3161 gnd.n3159 585
R2647 gnd.n3161 gnd.n3160 585
R2648 gnd.n3163 gnd.n3162 585
R2649 gnd.n3162 gnd.n1819 585
R2650 gnd.n3164 gnd.n3156 585
R2651 gnd.n3156 gnd.n1818 585
R2652 gnd.n3166 gnd.n3165 585
R2653 gnd.n3168 gnd.n3166 585
R2654 gnd.n3157 gnd.n3155 585
R2655 gnd.n3169 gnd.n3155 585
R2656 gnd.n3140 gnd.n3139 585
R2657 gnd.n3140 gnd.n1826 585
R2658 gnd.n3177 gnd.n3176 585
R2659 gnd.n3176 gnd.n3175 585
R2660 gnd.n3178 gnd.n3135 585
R2661 gnd.n3141 gnd.n3135 585
R2662 gnd.n3180 gnd.n3179 585
R2663 gnd.n3181 gnd.n3180 585
R2664 gnd.n3138 gnd.n3134 585
R2665 gnd.n3183 gnd.n3134 585
R2666 gnd.n3137 gnd.n3136 585
R2667 gnd.n3136 gnd.n1838 585
R2668 gnd.n3125 gnd.n3124 585
R2669 gnd.n3125 gnd.n1837 585
R2670 gnd.n3192 gnd.n3191 585
R2671 gnd.n3191 gnd.n3190 585
R2672 gnd.n3193 gnd.n3119 585
R2673 gnd.n3119 gnd.n1844 585
R2674 gnd.n3195 gnd.n3194 585
R2675 gnd.n3196 gnd.n3195 585
R2676 gnd.n3123 gnd.n3118 585
R2677 gnd.n3198 gnd.n3118 585
R2678 gnd.n3122 gnd.n3121 585
R2679 gnd.n3121 gnd.n1851 585
R2680 gnd.n3120 gnd.n1872 585
R2681 gnd.n1872 gnd.n1850 585
R2682 gnd.n3206 gnd.n1873 585
R2683 gnd.n3206 gnd.n3205 585
R2684 gnd.n3207 gnd.n1871 585
R2685 gnd.n3207 gnd.n1858 585
R2686 gnd.n3209 gnd.n3208 585
R2687 gnd.n3208 gnd.n1857 585
R2688 gnd.n3210 gnd.n1869 585
R2689 gnd.n1869 gnd.n1866 585
R2690 gnd.n3212 gnd.n3211 585
R2691 gnd.n3213 gnd.n3212 585
R2692 gnd.n1870 gnd.n1868 585
R2693 gnd.n3107 gnd.n1868 585
R2694 gnd.n2980 gnd.n2979 585
R2695 gnd.n2980 gnd.n1880 585
R2696 gnd.n2988 gnd.n2978 585
R2697 gnd.n2988 gnd.n2987 585
R2698 gnd.n2990 gnd.n2989 585
R2699 gnd.n2989 gnd.n1889 585
R2700 gnd.n2991 gnd.n2976 585
R2701 gnd.n2976 gnd.n1888 585
R2702 gnd.n2993 gnd.n2992 585
R2703 gnd.n2995 gnd.n2993 585
R2704 gnd.n2977 gnd.n2975 585
R2705 gnd.n2975 gnd.n1898 585
R2706 gnd.n2967 gnd.n2966 585
R2707 gnd.n2967 gnd.n1896 585
R2708 gnd.n3004 gnd.n3003 585
R2709 gnd.n3003 gnd.n3002 585
R2710 gnd.n3005 gnd.n2961 585
R2711 gnd.n2961 gnd.n1904 585
R2712 gnd.n3007 gnd.n3006 585
R2713 gnd.n3008 gnd.n3007 585
R2714 gnd.n2965 gnd.n2960 585
R2715 gnd.n3010 gnd.n2960 585
R2716 gnd.n2964 gnd.n2963 585
R2717 gnd.n2963 gnd.n1912 585
R2718 gnd.n2962 gnd.n2952 585
R2719 gnd.n2952 gnd.n1910 585
R2720 gnd.n3018 gnd.n2951 585
R2721 gnd.n3018 gnd.n3017 585
R2722 gnd.n3020 gnd.n3019 585
R2723 gnd.n3019 gnd.n1919 585
R2724 gnd.n3021 gnd.n2948 585
R2725 gnd.n2948 gnd.n1918 585
R2726 gnd.n3023 gnd.n3022 585
R2727 gnd.n3025 gnd.n3023 585
R2728 gnd.n2950 gnd.n2947 585
R2729 gnd.n2947 gnd.n1926 585
R2730 gnd.n2949 gnd.n1948 585
R2731 gnd.n1952 gnd.n1948 585
R2732 gnd.n3033 gnd.n1949 585
R2733 gnd.n3033 gnd.n3032 585
R2734 gnd.n3034 gnd.n1947 585
R2735 gnd.n3034 gnd.n1933 585
R2736 gnd.n3036 gnd.n3035 585
R2737 gnd.n3035 gnd.n1932 585
R2738 gnd.n3037 gnd.n1945 585
R2739 gnd.n1945 gnd.n1942 585
R2740 gnd.n3039 gnd.n3038 585
R2741 gnd.n3040 gnd.n3039 585
R2742 gnd.n1946 gnd.n1944 585
R2743 gnd.n2936 gnd.n1944 585
R2744 gnd.n2760 gnd.n2759 585
R2745 gnd.n2759 gnd.n1956 585
R2746 gnd.n2761 gnd.n2758 585
R2747 gnd.n2758 gnd.n2757 585
R2748 gnd.n2763 gnd.n2762 585
R2749 gnd.n2763 gnd.n1964 585
R2750 gnd.n2764 gnd.n2646 585
R2751 gnd.n2764 gnd.n1963 585
R2752 gnd.n2311 gnd.n2309 585
R2753 gnd.n2309 gnd.n1005 585
R2754 gnd.n6721 gnd.n6719 585
R2755 gnd.n6721 gnd.n6720 585
R2756 gnd.n6723 gnd.n6722 585
R2757 gnd.n6722 gnd.n201 585
R2758 gnd.n6724 gnd.n273 585
R2759 gnd.n273 gnd.n209 585
R2760 gnd.n6726 gnd.n6725 585
R2761 gnd.n6727 gnd.n6726 585
R2762 gnd.n274 gnd.n272 585
R2763 gnd.n272 gnd.n223 585
R2764 gnd.n4107 gnd.n4106 585
R2765 gnd.n4107 gnd.n221 585
R2766 gnd.n4109 gnd.n4108 585
R2767 gnd.n4108 gnd.n231 585
R2768 gnd.n4110 gnd.n1399 585
R2769 gnd.n1399 gnd.n229 585
R2770 gnd.n4113 gnd.n4112 585
R2771 gnd.n4114 gnd.n4113 585
R2772 gnd.n4104 gnd.n1398 585
R2773 gnd.n1398 gnd.n1397 585
R2774 gnd.n4102 gnd.n4101 585
R2775 gnd.n4101 gnd.n4100 585
R2776 gnd.n1401 gnd.n1400 585
R2777 gnd.n4090 gnd.n1401 585
R2778 gnd.n4067 gnd.n1433 585
R2779 gnd.n1433 gnd.n1406 585
R2780 gnd.n4069 gnd.n4068 585
R2781 gnd.n4070 gnd.n4069 585
R2782 gnd.n4064 gnd.n1432 585
R2783 gnd.n1432 gnd.n1415 585
R2784 gnd.n4063 gnd.n4062 585
R2785 gnd.n4062 gnd.n1420 585
R2786 gnd.n4061 gnd.n1434 585
R2787 gnd.n4061 gnd.n4060 585
R2788 gnd.n4035 gnd.n1436 585
R2789 gnd.n1445 gnd.n1436 585
R2790 gnd.n4036 gnd.n1457 585
R2791 gnd.n1457 gnd.n1443 585
R2792 gnd.n4038 gnd.n4037 585
R2793 gnd.n4039 gnd.n4038 585
R2794 gnd.n1458 gnd.n1456 585
R2795 gnd.n1456 gnd.n1453 585
R2796 gnd.n4028 gnd.n4027 585
R2797 gnd.n4027 gnd.n4026 585
R2798 gnd.n1461 gnd.n1460 585
R2799 gnd.n1471 gnd.n1461 585
R2800 gnd.n4002 gnd.n1482 585
R2801 gnd.n1482 gnd.n1469 585
R2802 gnd.n4004 gnd.n4003 585
R2803 gnd.n4005 gnd.n4004 585
R2804 gnd.n1483 gnd.n1481 585
R2805 gnd.n1481 gnd.n1478 585
R2806 gnd.n3997 gnd.n3996 585
R2807 gnd.n3996 gnd.n3995 585
R2808 gnd.n1486 gnd.n1485 585
R2809 gnd.n1497 gnd.n1486 585
R2810 gnd.n3970 gnd.n3958 585
R2811 gnd.n3958 gnd.n1495 585
R2812 gnd.n3972 gnd.n3971 585
R2813 gnd.n3973 gnd.n3972 585
R2814 gnd.n3959 gnd.n3957 585
R2815 gnd.n3957 gnd.n1364 585
R2816 gnd.n3965 gnd.n3964 585
R2817 gnd.n3964 gnd.n1362 585
R2818 gnd.n3963 gnd.n3962 585
R2819 gnd.n3963 gnd.n1311 585
R2820 gnd.n1282 gnd.n1281 585
R2821 gnd.n4230 gnd.n1282 585
R2822 gnd.n4233 gnd.n4232 585
R2823 gnd.n4232 gnd.n4231 585
R2824 gnd.n4234 gnd.n1276 585
R2825 gnd.n1276 gnd.n1275 585
R2826 gnd.n4236 gnd.n4235 585
R2827 gnd.n4237 gnd.n4236 585
R2828 gnd.n1277 gnd.n1273 585
R2829 gnd.n4238 gnd.n1273 585
R2830 gnd.n3880 gnd.n1645 585
R2831 gnd.n1645 gnd.n1272 585
R2832 gnd.n3882 gnd.n3881 585
R2833 gnd.n3883 gnd.n3882 585
R2834 gnd.n1646 gnd.n1644 585
R2835 gnd.n3715 gnd.n1644 585
R2836 gnd.n3874 gnd.n3873 585
R2837 gnd.n3873 gnd.n3872 585
R2838 gnd.n1649 gnd.n1648 585
R2839 gnd.n3515 gnd.n1649 585
R2840 gnd.n3861 gnd.n3860 585
R2841 gnd.n3862 gnd.n3861 585
R2842 gnd.n1660 gnd.n1659 585
R2843 gnd.n3729 gnd.n1659 585
R2844 gnd.n3856 gnd.n3855 585
R2845 gnd.n3855 gnd.n3854 585
R2846 gnd.n1663 gnd.n1662 585
R2847 gnd.n3501 gnd.n1663 585
R2848 gnd.n3845 gnd.n3844 585
R2849 gnd.n3846 gnd.n3845 585
R2850 gnd.n1674 gnd.n1673 585
R2851 gnd.n3744 gnd.n1673 585
R2852 gnd.n3840 gnd.n3839 585
R2853 gnd.n3839 gnd.n3838 585
R2854 gnd.n1677 gnd.n1676 585
R2855 gnd.n3489 gnd.n1677 585
R2856 gnd.n3829 gnd.n3828 585
R2857 gnd.n3830 gnd.n3829 585
R2858 gnd.n1687 gnd.n1686 585
R2859 gnd.n3759 gnd.n1686 585
R2860 gnd.n3824 gnd.n3823 585
R2861 gnd.n3823 gnd.n3822 585
R2862 gnd.n1690 gnd.n1689 585
R2863 gnd.n3473 gnd.n1690 585
R2864 gnd.n3813 gnd.n3812 585
R2865 gnd.n3814 gnd.n3813 585
R2866 gnd.n1701 gnd.n1700 585
R2867 gnd.t232 gnd.n1700 585
R2868 gnd.n3808 gnd.n3807 585
R2869 gnd.n3807 gnd.n3806 585
R2870 gnd.n1704 gnd.n1703 585
R2871 gnd.n1727 gnd.n1704 585
R2872 gnd.n3797 gnd.n3796 585
R2873 gnd.n3798 gnd.n3797 585
R2874 gnd.n1714 gnd.n1713 585
R2875 gnd.n3459 gnd.n1713 585
R2876 gnd.n3792 gnd.n3791 585
R2877 gnd.n3791 gnd.n3790 585
R2878 gnd.n1717 gnd.n1716 585
R2879 gnd.n3451 gnd.n1717 585
R2880 gnd.n3439 gnd.n1745 585
R2881 gnd.n1745 gnd.n1733 585
R2882 gnd.n3441 gnd.n3440 585
R2883 gnd.n3442 gnd.n3441 585
R2884 gnd.n1746 gnd.n1744 585
R2885 gnd.n3338 gnd.n1744 585
R2886 gnd.n3434 gnd.n3433 585
R2887 gnd.n3433 gnd.n3432 585
R2888 gnd.n1749 gnd.n1748 585
R2889 gnd.n3314 gnd.n1749 585
R2890 gnd.n3423 gnd.n3422 585
R2891 gnd.n3424 gnd.n3423 585
R2892 gnd.n1759 gnd.n1758 585
R2893 gnd.n3353 gnd.n1758 585
R2894 gnd.n3418 gnd.n3417 585
R2895 gnd.n3417 gnd.n3416 585
R2896 gnd.n1762 gnd.n1761 585
R2897 gnd.n3299 gnd.n1762 585
R2898 gnd.n3407 gnd.n3406 585
R2899 gnd.n3408 gnd.n3407 585
R2900 gnd.n1774 gnd.n1773 585
R2901 gnd.n3368 gnd.n1773 585
R2902 gnd.n3402 gnd.n3401 585
R2903 gnd.n3401 gnd.n3400 585
R2904 gnd.n1777 gnd.n1776 585
R2905 gnd.n1804 gnd.n1777 585
R2906 gnd.n3391 gnd.n3390 585
R2907 gnd.n3392 gnd.n3391 585
R2908 gnd.n1789 gnd.n1788 585
R2909 gnd.n1795 gnd.n1788 585
R2910 gnd.n3386 gnd.n3385 585
R2911 gnd.n3385 gnd.n3384 585
R2912 gnd.n1792 gnd.n1791 585
R2913 gnd.n3280 gnd.n1792 585
R2914 gnd.n3268 gnd.n1821 585
R2915 gnd.n1821 gnd.n1810 585
R2916 gnd.n3270 gnd.n3269 585
R2917 gnd.n3271 gnd.n3270 585
R2918 gnd.n1822 gnd.n1820 585
R2919 gnd.n3167 gnd.n1820 585
R2920 gnd.n3263 gnd.n3262 585
R2921 gnd.n3262 gnd.n3261 585
R2922 gnd.n1825 gnd.n1824 585
R2923 gnd.n3143 gnd.n1825 585
R2924 gnd.n3252 gnd.n3251 585
R2925 gnd.n3253 gnd.n3252 585
R2926 gnd.n1833 gnd.n1832 585
R2927 gnd.n3182 gnd.n1832 585
R2928 gnd.n3247 gnd.n3246 585
R2929 gnd.n3246 gnd.n3245 585
R2930 gnd.n1836 gnd.n1835 585
R2931 gnd.n3127 gnd.n1836 585
R2932 gnd.n3236 gnd.n3235 585
R2933 gnd.n3237 gnd.n3236 585
R2934 gnd.n1846 gnd.n1845 585
R2935 gnd.n3197 gnd.n1845 585
R2936 gnd.n3231 gnd.n3230 585
R2937 gnd.n3230 gnd.n3229 585
R2938 gnd.n1849 gnd.n1848 585
R2939 gnd.n1875 gnd.n1849 585
R2940 gnd.n3220 gnd.n3219 585
R2941 gnd.n3221 gnd.n3220 585
R2942 gnd.n1860 gnd.n1859 585
R2943 gnd.n1865 gnd.n1859 585
R2944 gnd.n3215 gnd.n3214 585
R2945 gnd.n3214 gnd.n3213 585
R2946 gnd.n1863 gnd.n1862 585
R2947 gnd.n3106 gnd.n1863 585
R2948 gnd.n3094 gnd.n1891 585
R2949 gnd.n2981 gnd.n1891 585
R2950 gnd.n3096 gnd.n3095 585
R2951 gnd.n3097 gnd.n3096 585
R2952 gnd.n1892 gnd.n1890 585
R2953 gnd.n2994 gnd.n1890 585
R2954 gnd.n3089 gnd.n3088 585
R2955 gnd.n3088 gnd.t79 585
R2956 gnd.n1895 gnd.n1894 585
R2957 gnd.n2968 gnd.n1895 585
R2958 gnd.n3079 gnd.n3078 585
R2959 gnd.n3080 gnd.n3079 585
R2960 gnd.n1906 gnd.n1905 585
R2961 gnd.n3009 gnd.n1905 585
R2962 gnd.n3074 gnd.n3073 585
R2963 gnd.n3073 gnd.n3072 585
R2964 gnd.n1909 gnd.n1908 585
R2965 gnd.n2953 gnd.n1909 585
R2966 gnd.n3063 gnd.n3062 585
R2967 gnd.n3064 gnd.n3063 585
R2968 gnd.n1921 gnd.n1920 585
R2969 gnd.n3024 gnd.n1920 585
R2970 gnd.n3058 gnd.n3057 585
R2971 gnd.n3057 gnd.n3056 585
R2972 gnd.n1924 gnd.n1923 585
R2973 gnd.n1951 gnd.n1924 585
R2974 gnd.n3047 gnd.n3046 585
R2975 gnd.n3048 gnd.n3047 585
R2976 gnd.n1935 gnd.n1934 585
R2977 gnd.n1941 gnd.n1934 585
R2978 gnd.n3042 gnd.n3041 585
R2979 gnd.n3041 gnd.n3040 585
R2980 gnd.n1938 gnd.n1937 585
R2981 gnd.n2935 gnd.n1938 585
R2982 gnd.n2923 gnd.n1966 585
R2983 gnd.n2647 gnd.n1966 585
R2984 gnd.n2925 gnd.n2924 585
R2985 gnd.n2926 gnd.n2925 585
R2986 gnd.n1967 gnd.n1965 585
R2987 gnd.n1972 gnd.n1965 585
R2988 gnd.n2918 gnd.n2917 585
R2989 gnd.n2917 gnd.n2916 585
R2990 gnd.n1970 gnd.n1969 585
R2991 gnd.n1979 gnd.n1970 585
R2992 gnd.n2907 gnd.n2906 585
R2993 gnd.n2908 gnd.n2907 585
R2994 gnd.n1981 gnd.n1980 585
R2995 gnd.n1980 gnd.n1978 585
R2996 gnd.n2902 gnd.n2901 585
R2997 gnd.n2901 gnd.n2900 585
R2998 gnd.n1984 gnd.n1983 585
R2999 gnd.n1985 gnd.n1984 585
R3000 gnd.n2263 gnd.n2262 585
R3001 gnd.n2263 gnd.n2118 585
R3002 gnd.n2265 gnd.n2264 585
R3003 gnd.n2264 gnd.n2018 585
R3004 gnd.n2266 gnd.n2256 585
R3005 gnd.n2256 gnd.n1162 585
R3006 gnd.n2268 gnd.n2267 585
R3007 gnd.n2268 gnd.n1159 585
R3008 gnd.n2269 gnd.n2255 585
R3009 gnd.n2269 gnd.n2184 585
R3010 gnd.n2271 gnd.n2270 585
R3011 gnd.n2270 gnd.n1150 585
R3012 gnd.n2272 gnd.n2250 585
R3013 gnd.n2250 gnd.n1142 585
R3014 gnd.n2274 gnd.n2273 585
R3015 gnd.n2274 gnd.n1139 585
R3016 gnd.n2275 gnd.n2249 585
R3017 gnd.n2275 gnd.n1131 585
R3018 gnd.n2277 gnd.n2276 585
R3019 gnd.n2276 gnd.n1128 585
R3020 gnd.n2278 gnd.n2244 585
R3021 gnd.n2244 gnd.n1120 585
R3022 gnd.n2280 gnd.n2279 585
R3023 gnd.n2280 gnd.n1117 585
R3024 gnd.n2281 gnd.n2243 585
R3025 gnd.n2281 gnd.n1109 585
R3026 gnd.n2283 gnd.n2282 585
R3027 gnd.n2282 gnd.n1106 585
R3028 gnd.n2284 gnd.n2238 585
R3029 gnd.n2238 gnd.n2201 585
R3030 gnd.n2286 gnd.n2285 585
R3031 gnd.n2286 gnd.n1096 585
R3032 gnd.n2287 gnd.n2237 585
R3033 gnd.n2287 gnd.n1088 585
R3034 gnd.n2289 gnd.n2288 585
R3035 gnd.n2288 gnd.n1085 585
R3036 gnd.n2290 gnd.n2235 585
R3037 gnd.n2235 gnd.n1077 585
R3038 gnd.n2292 gnd.n2291 585
R3039 gnd.n2292 gnd.n1074 585
R3040 gnd.n2294 gnd.n2293 585
R3041 gnd.n2293 gnd.n1069 585
R3042 gnd.n2296 gnd.n2295 585
R3043 gnd.n2296 gnd.n1066 585
R3044 gnd.n2298 gnd.n2297 585
R3045 gnd.n2297 gnd.n2214 585
R3046 gnd.n2300 gnd.n2299 585
R3047 gnd.n2300 gnd.n1057 585
R3048 gnd.n2302 gnd.n2301 585
R3049 gnd.n2302 gnd.n1052 585
R3050 gnd.n2303 gnd.n2234 585
R3051 gnd.n2303 gnd.n1049 585
R3052 gnd.n2305 gnd.n2304 585
R3053 gnd.n2304 gnd.n1038 585
R3054 gnd.n2229 gnd.n2227 585
R3055 gnd.n2227 gnd.n1035 585
R3056 gnd.n2324 gnd.n2323 585
R3057 gnd.n2325 gnd.n2324 585
R3058 gnd.n2228 gnd.n2226 585
R3059 gnd.n2226 gnd.n1027 585
R3060 gnd.n2318 gnd.n2317 585
R3061 gnd.n2317 gnd.n1024 585
R3062 gnd.n2316 gnd.n2308 585
R3063 gnd.n2316 gnd.n1016 585
R3064 gnd.n2315 gnd.n2314 585
R3065 gnd.n2315 gnd.n1013 585
R3066 gnd.n4240 gnd.n4239 585
R3067 gnd.n4239 gnd.n4238 585
R3068 gnd.n4241 gnd.n1269 585
R3069 gnd.n1272 gnd.n1269 585
R3070 gnd.n4242 gnd.n1268 585
R3071 gnd.n3883 gnd.n1268 585
R3072 gnd.n3542 gnd.n1266 585
R3073 gnd.n3715 gnd.n3542 585
R3074 gnd.n4246 gnd.n1265 585
R3075 gnd.n3872 gnd.n1265 585
R3076 gnd.n4247 gnd.n1264 585
R3077 gnd.n3515 gnd.n1264 585
R3078 gnd.n4248 gnd.n1263 585
R3079 gnd.n3862 gnd.n1263 585
R3080 gnd.n3508 gnd.n1261 585
R3081 gnd.n3729 gnd.n3508 585
R3082 gnd.n4252 gnd.n1260 585
R3083 gnd.n3854 gnd.n1260 585
R3084 gnd.n4253 gnd.n1259 585
R3085 gnd.n3501 gnd.n1259 585
R3086 gnd.n4254 gnd.n1258 585
R3087 gnd.n3846 gnd.n1258 585
R3088 gnd.n3743 gnd.n1256 585
R3089 gnd.n3744 gnd.n3743 585
R3090 gnd.n4258 gnd.n1255 585
R3091 gnd.n3838 gnd.n1255 585
R3092 gnd.n4259 gnd.n1254 585
R3093 gnd.n3489 gnd.n1254 585
R3094 gnd.n4260 gnd.n1253 585
R3095 gnd.n3830 gnd.n1253 585
R3096 gnd.n3481 gnd.n1251 585
R3097 gnd.n3759 gnd.n3481 585
R3098 gnd.n4264 gnd.n1250 585
R3099 gnd.n3822 gnd.n1250 585
R3100 gnd.n4265 gnd.n1249 585
R3101 gnd.n3473 gnd.n1249 585
R3102 gnd.n4266 gnd.n1248 585
R3103 gnd.n3814 gnd.n1248 585
R3104 gnd.n3774 gnd.n1246 585
R3105 gnd.t232 gnd.n3774 585
R3106 gnd.n4270 gnd.n1245 585
R3107 gnd.n3806 gnd.n1245 585
R3108 gnd.n4271 gnd.n1244 585
R3109 gnd.n1727 gnd.n1244 585
R3110 gnd.n4272 gnd.n1243 585
R3111 gnd.n3798 gnd.n1243 585
R3112 gnd.n3458 gnd.n1241 585
R3113 gnd.n3459 gnd.n3458 585
R3114 gnd.n4276 gnd.n1240 585
R3115 gnd.n3790 gnd.n1240 585
R3116 gnd.n4277 gnd.n1239 585
R3117 gnd.n3451 gnd.n1239 585
R3118 gnd.n4278 gnd.n1238 585
R3119 gnd.n1733 gnd.n1238 585
R3120 gnd.n1742 gnd.n1236 585
R3121 gnd.n3442 gnd.n1742 585
R3122 gnd.n4282 gnd.n1235 585
R3123 gnd.n3338 gnd.n1235 585
R3124 gnd.n4283 gnd.n1234 585
R3125 gnd.n3432 gnd.n1234 585
R3126 gnd.n4284 gnd.n1233 585
R3127 gnd.n3314 gnd.n1233 585
R3128 gnd.n1756 gnd.n1231 585
R3129 gnd.n3424 gnd.n1756 585
R3130 gnd.n4288 gnd.n1230 585
R3131 gnd.n3353 gnd.n1230 585
R3132 gnd.n4289 gnd.n1229 585
R3133 gnd.n3416 gnd.n1229 585
R3134 gnd.n4290 gnd.n1228 585
R3135 gnd.n3299 gnd.n1228 585
R3136 gnd.n1771 gnd.n1226 585
R3137 gnd.n3408 gnd.n1771 585
R3138 gnd.n4294 gnd.n1225 585
R3139 gnd.n3368 gnd.n1225 585
R3140 gnd.n4295 gnd.n1224 585
R3141 gnd.n3400 gnd.n1224 585
R3142 gnd.n4296 gnd.n1223 585
R3143 gnd.n1804 gnd.n1223 585
R3144 gnd.n1786 gnd.n1221 585
R3145 gnd.n3392 gnd.n1786 585
R3146 gnd.n4300 gnd.n1220 585
R3147 gnd.n1795 gnd.n1220 585
R3148 gnd.n4301 gnd.n1219 585
R3149 gnd.n3384 gnd.n1219 585
R3150 gnd.n4302 gnd.n1218 585
R3151 gnd.n3280 gnd.n1218 585
R3152 gnd.n1809 gnd.n1216 585
R3153 gnd.n1810 gnd.n1809 585
R3154 gnd.n4306 gnd.n1215 585
R3155 gnd.n3271 gnd.n1215 585
R3156 gnd.n4307 gnd.n1214 585
R3157 gnd.n3167 gnd.n1214 585
R3158 gnd.n4308 gnd.n1213 585
R3159 gnd.n3261 gnd.n1213 585
R3160 gnd.n3142 gnd.n1211 585
R3161 gnd.n3143 gnd.n3142 585
R3162 gnd.n4312 gnd.n1210 585
R3163 gnd.n3253 gnd.n1210 585
R3164 gnd.n4313 gnd.n1209 585
R3165 gnd.n3182 gnd.n1209 585
R3166 gnd.n4314 gnd.n1208 585
R3167 gnd.n3245 gnd.n1208 585
R3168 gnd.n3126 gnd.n1206 585
R3169 gnd.n3127 gnd.n3126 585
R3170 gnd.n4318 gnd.n1205 585
R3171 gnd.n3237 gnd.n1205 585
R3172 gnd.n4319 gnd.n1204 585
R3173 gnd.n3197 gnd.n1204 585
R3174 gnd.n4320 gnd.n1203 585
R3175 gnd.n3229 gnd.n1203 585
R3176 gnd.n1874 gnd.n1201 585
R3177 gnd.n1875 gnd.n1874 585
R3178 gnd.n4324 gnd.n1200 585
R3179 gnd.n3221 gnd.n1200 585
R3180 gnd.n4325 gnd.n1199 585
R3181 gnd.n1865 gnd.n1199 585
R3182 gnd.n4326 gnd.n1198 585
R3183 gnd.n3213 gnd.n1198 585
R3184 gnd.n1881 gnd.n1196 585
R3185 gnd.n3106 gnd.n1881 585
R3186 gnd.n4330 gnd.n1195 585
R3187 gnd.n2981 gnd.n1195 585
R3188 gnd.n4331 gnd.n1194 585
R3189 gnd.n3097 gnd.n1194 585
R3190 gnd.n4332 gnd.n1193 585
R3191 gnd.n2994 gnd.n1193 585
R3192 gnd.n1897 gnd.n1191 585
R3193 gnd.t79 gnd.n1897 585
R3194 gnd.n4336 gnd.n1190 585
R3195 gnd.n2968 gnd.n1190 585
R3196 gnd.n4337 gnd.n1189 585
R3197 gnd.n3080 gnd.n1189 585
R3198 gnd.n4338 gnd.n1188 585
R3199 gnd.n3009 gnd.n1188 585
R3200 gnd.n1911 gnd.n1186 585
R3201 gnd.n3072 gnd.n1911 585
R3202 gnd.n4342 gnd.n1185 585
R3203 gnd.n2953 gnd.n1185 585
R3204 gnd.n4343 gnd.n1184 585
R3205 gnd.n3064 gnd.n1184 585
R3206 gnd.n4344 gnd.n1183 585
R3207 gnd.n3024 gnd.n1183 585
R3208 gnd.n1925 gnd.n1181 585
R3209 gnd.n3056 gnd.n1925 585
R3210 gnd.n4348 gnd.n1180 585
R3211 gnd.n1951 gnd.n1180 585
R3212 gnd.n4349 gnd.n1179 585
R3213 gnd.n3048 gnd.n1179 585
R3214 gnd.n4350 gnd.n1178 585
R3215 gnd.n1941 gnd.n1178 585
R3216 gnd.n1940 gnd.n1176 585
R3217 gnd.n3040 gnd.n1940 585
R3218 gnd.n4354 gnd.n1175 585
R3219 gnd.n2935 gnd.n1175 585
R3220 gnd.n4355 gnd.n1174 585
R3221 gnd.n2647 gnd.n1174 585
R3222 gnd.n4356 gnd.n1173 585
R3223 gnd.n2926 gnd.n1173 585
R3224 gnd.n1971 gnd.n1171 585
R3225 gnd.n1972 gnd.n1971 585
R3226 gnd.n4360 gnd.n1170 585
R3227 gnd.n2916 gnd.n1170 585
R3228 gnd.n4361 gnd.n1169 585
R3229 gnd.n1979 gnd.n1169 585
R3230 gnd.n4362 gnd.n1168 585
R3231 gnd.n2908 gnd.n1168 585
R3232 gnd.n2058 gnd.n2057 585
R3233 gnd.n2061 gnd.n2060 585
R3234 gnd.n2059 gnd.n2048 585
R3235 gnd.n2071 gnd.n2070 585
R3236 gnd.n2073 gnd.n2072 585
R3237 gnd.n2043 gnd.n2042 585
R3238 gnd.n2082 gnd.n2044 585
R3239 gnd.n2085 gnd.n2084 585
R3240 gnd.n2083 gnd.n2036 585
R3241 gnd.n2095 gnd.n2094 585
R3242 gnd.n2097 gnd.n2096 585
R3243 gnd.n2031 gnd.n2030 585
R3244 gnd.n2107 gnd.n2032 585
R3245 gnd.n2109 gnd.n2108 585
R3246 gnd.n2111 gnd.n2110 585
R3247 gnd.n2011 gnd.n2010 585
R3248 gnd.n2869 gnd.n2012 585
R3249 gnd.n2872 gnd.n2871 585
R3250 gnd.n2870 gnd.n2007 585
R3251 gnd.n2878 gnd.n2877 585
R3252 gnd.n2880 gnd.n2879 585
R3253 gnd.n2883 gnd.n2882 585
R3254 gnd.n2881 gnd.n2005 585
R3255 gnd.n2888 gnd.n2887 585
R3256 gnd.n2890 gnd.n2889 585
R3257 gnd.n2893 gnd.n2892 585
R3258 gnd.n2000 gnd.n1999 585
R3259 gnd.n2898 gnd.n2897 585
R3260 gnd.n2001 gnd.n1977 585
R3261 gnd.n2900 gnd.n1977 585
R3262 gnd.n3887 gnd.n1274 585
R3263 gnd.n4238 gnd.n1274 585
R3264 gnd.n3886 gnd.n3885 585
R3265 gnd.n3885 gnd.n1272 585
R3266 gnd.n3884 gnd.n1642 585
R3267 gnd.n3884 gnd.n3883 585
R3268 gnd.n1653 gnd.n1643 585
R3269 gnd.n3715 gnd.n1643 585
R3270 gnd.n3871 gnd.n3870 585
R3271 gnd.n3872 gnd.n3871 585
R3272 gnd.n1652 gnd.n1651 585
R3273 gnd.n3515 gnd.n1651 585
R3274 gnd.n3864 gnd.n3863 585
R3275 gnd.n3863 gnd.n3862 585
R3276 gnd.n1656 gnd.n1655 585
R3277 gnd.n3729 gnd.n1656 585
R3278 gnd.n3853 gnd.n3852 585
R3279 gnd.n3854 gnd.n3853 585
R3280 gnd.n1667 gnd.n1666 585
R3281 gnd.n3501 gnd.n1666 585
R3282 gnd.n3848 gnd.n3847 585
R3283 gnd.n3847 gnd.n3846 585
R3284 gnd.n1670 gnd.n1669 585
R3285 gnd.n3744 gnd.n1670 585
R3286 gnd.n3837 gnd.n3836 585
R3287 gnd.n3838 gnd.n3837 585
R3288 gnd.n1681 gnd.n1680 585
R3289 gnd.n3489 gnd.n1680 585
R3290 gnd.n3832 gnd.n3831 585
R3291 gnd.n3831 gnd.n3830 585
R3292 gnd.n1684 gnd.n1683 585
R3293 gnd.n3759 gnd.n1684 585
R3294 gnd.n3821 gnd.n3820 585
R3295 gnd.n3822 gnd.n3821 585
R3296 gnd.n1694 gnd.n1693 585
R3297 gnd.n3473 gnd.n1693 585
R3298 gnd.n3816 gnd.n3815 585
R3299 gnd.n3815 gnd.n3814 585
R3300 gnd.n1697 gnd.n1696 585
R3301 gnd.t232 gnd.n1697 585
R3302 gnd.n3805 gnd.n3804 585
R3303 gnd.n3806 gnd.n3805 585
R3304 gnd.n1707 gnd.n1706 585
R3305 gnd.n1727 gnd.n1706 585
R3306 gnd.n3800 gnd.n3799 585
R3307 gnd.n3799 gnd.n3798 585
R3308 gnd.n1710 gnd.n1709 585
R3309 gnd.n3459 gnd.n1710 585
R3310 gnd.n1737 gnd.n1720 585
R3311 gnd.n3790 gnd.n1720 585
R3312 gnd.n3450 gnd.n3449 585
R3313 gnd.n3451 gnd.n3450 585
R3314 gnd.n1736 gnd.n1735 585
R3315 gnd.n1735 gnd.n1733 585
R3316 gnd.n3444 gnd.n3443 585
R3317 gnd.n3443 gnd.n3442 585
R3318 gnd.n1740 gnd.n1739 585
R3319 gnd.n3338 gnd.n1740 585
R3320 gnd.n3431 gnd.n3430 585
R3321 gnd.n3432 gnd.n3431 585
R3322 gnd.n1752 gnd.n1751 585
R3323 gnd.n3314 gnd.n1751 585
R3324 gnd.n3426 gnd.n3425 585
R3325 gnd.n3425 gnd.n3424 585
R3326 gnd.n1755 gnd.n1754 585
R3327 gnd.n3353 gnd.n1755 585
R3328 gnd.n3415 gnd.n3414 585
R3329 gnd.n3416 gnd.n3415 585
R3330 gnd.n1766 gnd.n1765 585
R3331 gnd.n3299 gnd.n1765 585
R3332 gnd.n3410 gnd.n3409 585
R3333 gnd.n3409 gnd.n3408 585
R3334 gnd.n1769 gnd.n1768 585
R3335 gnd.n3368 gnd.n1769 585
R3336 gnd.n3399 gnd.n3398 585
R3337 gnd.n3400 gnd.n3399 585
R3338 gnd.n1781 gnd.n1780 585
R3339 gnd.n1804 gnd.n1780 585
R3340 gnd.n3394 gnd.n3393 585
R3341 gnd.n3393 gnd.n3392 585
R3342 gnd.n1784 gnd.n1783 585
R3343 gnd.n1795 gnd.n1784 585
R3344 gnd.n1814 gnd.n1797 585
R3345 gnd.n3384 gnd.n1797 585
R3346 gnd.n3279 gnd.n3278 585
R3347 gnd.n3280 gnd.n3279 585
R3348 gnd.n1813 gnd.n1812 585
R3349 gnd.n1812 gnd.n1810 585
R3350 gnd.n3273 gnd.n3272 585
R3351 gnd.n3272 gnd.n3271 585
R3352 gnd.n1817 gnd.n1816 585
R3353 gnd.n3167 gnd.n1817 585
R3354 gnd.n3260 gnd.n3259 585
R3355 gnd.n3261 gnd.n3260 585
R3356 gnd.n1828 gnd.n1827 585
R3357 gnd.n3143 gnd.n1827 585
R3358 gnd.n3255 gnd.n3254 585
R3359 gnd.n3254 gnd.n3253 585
R3360 gnd.n1831 gnd.n1830 585
R3361 gnd.n3182 gnd.n1831 585
R3362 gnd.n3244 gnd.n3243 585
R3363 gnd.n3245 gnd.n3244 585
R3364 gnd.n1840 gnd.n1839 585
R3365 gnd.n3127 gnd.n1839 585
R3366 gnd.n3239 gnd.n3238 585
R3367 gnd.n3238 gnd.n3237 585
R3368 gnd.n1843 gnd.n1842 585
R3369 gnd.n3197 gnd.n1843 585
R3370 gnd.n3228 gnd.n3227 585
R3371 gnd.n3229 gnd.n3228 585
R3372 gnd.n1853 gnd.n1852 585
R3373 gnd.n1875 gnd.n1852 585
R3374 gnd.n3223 gnd.n3222 585
R3375 gnd.n3222 gnd.n3221 585
R3376 gnd.n1856 gnd.n1855 585
R3377 gnd.n1865 gnd.n1856 585
R3378 gnd.n1884 gnd.n1867 585
R3379 gnd.n3213 gnd.n1867 585
R3380 gnd.n3105 gnd.n3104 585
R3381 gnd.n3106 gnd.n3105 585
R3382 gnd.n1883 gnd.n1882 585
R3383 gnd.n2981 gnd.n1882 585
R3384 gnd.n3099 gnd.n3098 585
R3385 gnd.n3098 gnd.n3097 585
R3386 gnd.n1887 gnd.n1886 585
R3387 gnd.n2994 gnd.n1887 585
R3388 gnd.n3087 gnd.n3086 585
R3389 gnd.t79 gnd.n3087 585
R3390 gnd.n1900 gnd.n1899 585
R3391 gnd.n2968 gnd.n1899 585
R3392 gnd.n3082 gnd.n3081 585
R3393 gnd.n3081 gnd.n3080 585
R3394 gnd.n1903 gnd.n1902 585
R3395 gnd.n3009 gnd.n1903 585
R3396 gnd.n3071 gnd.n3070 585
R3397 gnd.n3072 gnd.n3071 585
R3398 gnd.n1914 gnd.n1913 585
R3399 gnd.n2953 gnd.n1913 585
R3400 gnd.n3066 gnd.n3065 585
R3401 gnd.n3065 gnd.n3064 585
R3402 gnd.n1917 gnd.n1916 585
R3403 gnd.n3024 gnd.n1917 585
R3404 gnd.n3055 gnd.n3054 585
R3405 gnd.n3056 gnd.n3055 585
R3406 gnd.n1928 gnd.n1927 585
R3407 gnd.n1951 gnd.n1927 585
R3408 gnd.n3050 gnd.n3049 585
R3409 gnd.n3049 gnd.n3048 585
R3410 gnd.n1931 gnd.n1930 585
R3411 gnd.n1941 gnd.n1931 585
R3412 gnd.n1959 gnd.n1943 585
R3413 gnd.n3040 gnd.n1943 585
R3414 gnd.n2934 gnd.n2933 585
R3415 gnd.n2935 gnd.n2934 585
R3416 gnd.n1958 gnd.n1957 585
R3417 gnd.n2647 gnd.n1957 585
R3418 gnd.n2928 gnd.n2927 585
R3419 gnd.n2927 gnd.n2926 585
R3420 gnd.n1962 gnd.n1961 585
R3421 gnd.n1972 gnd.n1962 585
R3422 gnd.n2915 gnd.n2914 585
R3423 gnd.n2916 gnd.n2915 585
R3424 gnd.n1975 gnd.n1974 585
R3425 gnd.n1979 gnd.n1974 585
R3426 gnd.n2910 gnd.n2909 585
R3427 gnd.n2909 gnd.n2908 585
R3428 gnd.n3894 gnd.n3893 585
R3429 gnd.n3893 gnd.n1275 585
R3430 gnd.n3895 gnd.n3892 585
R3431 gnd.n3890 gnd.n1640 585
R3432 gnd.n3899 gnd.n1639 585
R3433 gnd.n3903 gnd.n1637 585
R3434 gnd.n3904 gnd.n1636 585
R3435 gnd.n1634 gnd.n1632 585
R3436 gnd.n3908 gnd.n1631 585
R3437 gnd.n3909 gnd.n1629 585
R3438 gnd.n3910 gnd.n1628 585
R3439 gnd.n1626 gnd.n1506 585
R3440 gnd.n1625 gnd.n1507 585
R3441 gnd.n1623 gnd.n1622 585
R3442 gnd.n1509 gnd.n1508 585
R3443 gnd.n1613 gnd.n1612 585
R3444 gnd.n1610 gnd.n1519 585
R3445 gnd.n1608 gnd.n1607 585
R3446 gnd.n1521 gnd.n1520 585
R3447 gnd.n1596 gnd.n1595 585
R3448 gnd.n1593 gnd.n1528 585
R3449 gnd.n1591 gnd.n1590 585
R3450 gnd.n1530 gnd.n1529 585
R3451 gnd.n1579 gnd.n1578 585
R3452 gnd.n1576 gnd.n1537 585
R3453 gnd.n1574 gnd.n1573 585
R3454 gnd.n1539 gnd.n1538 585
R3455 gnd.n1562 gnd.n1561 585
R3456 gnd.n1559 gnd.n1557 585
R3457 gnd.n1546 gnd.n1271 585
R3458 gnd.n3717 gnd.n3540 506.916
R3459 gnd.n3648 gnd.n3541 506.916
R3460 gnd.n2766 gnd.n2764 506.916
R3461 gnd.n2752 gnd.n2751 506.916
R3462 gnd.n6120 gnd.n6119 475.281
R3463 gnd.n2630 gnd.t209 389.64
R3464 gnd.n3644 gnd.t142 389.64
R3465 gnd.n2685 gnd.t156 389.64
R3466 gnd.n3559 gnd.t196 389.64
R3467 gnd.n2003 gnd.t189 371.625
R3468 gnd.n6833 gnd.t177 371.625
R3469 gnd.n1513 gnd.t163 371.625
R3470 gnd.n2015 gnd.t183 371.625
R3471 gnd.n1334 gnd.t160 371.625
R3472 gnd.n1356 gnd.t131 371.625
R3473 gnd.n157 gnd.t117 371.625
R3474 gnd.n6925 gnd.t146 371.625
R3475 gnd.n928 gnd.t215 371.625
R3476 gnd.n950 gnd.t206 371.625
R3477 gnd.n2377 gnd.t202 371.625
R3478 gnd.n2180 gnd.t138 371.625
R3479 gnd.n2158 gnd.t180 371.625
R3480 gnd.n3900 gnd.t173 371.625
R3481 gnd.n5131 gnd.t124 323.425
R3482 gnd.n4597 gnd.t166 323.425
R3483 gnd.n5799 gnd.n5773 289.615
R3484 gnd.n5767 gnd.n5741 289.615
R3485 gnd.n5735 gnd.n5709 289.615
R3486 gnd.n5704 gnd.n5678 289.615
R3487 gnd.n5672 gnd.n5646 289.615
R3488 gnd.n5640 gnd.n5614 289.615
R3489 gnd.n5608 gnd.n5582 289.615
R3490 gnd.n5577 gnd.n5551 289.615
R3491 gnd.n4981 gnd.t218 279.217
R3492 gnd.n4623 gnd.t152 279.217
R3493 gnd.n2655 gnd.t195 260.649
R3494 gnd.n3531 gnd.t201 260.649
R3495 gnd.n2670 gnd.n1973 256.663
R3496 gnd.n2672 gnd.n1973 256.663
R3497 gnd.n2741 gnd.n1973 256.663
R3498 gnd.n2735 gnd.n1973 256.663
R3499 gnd.n2733 gnd.n1973 256.663
R3500 gnd.n2727 gnd.n1973 256.663
R3501 gnd.n2725 gnd.n1973 256.663
R3502 gnd.n2719 gnd.n1973 256.663
R3503 gnd.n2717 gnd.n1973 256.663
R3504 gnd.n2711 gnd.n1973 256.663
R3505 gnd.n2709 gnd.n1973 256.663
R3506 gnd.n2703 gnd.n1973 256.663
R3507 gnd.n2701 gnd.n1973 256.663
R3508 gnd.n2695 gnd.n1973 256.663
R3509 gnd.n2688 gnd.n1973 256.663
R3510 gnd.n2689 gnd.n1973 256.663
R3511 gnd.n2832 gnd.n2628 256.663
R3512 gnd.n2830 gnd.n1973 256.663
R3513 gnd.n2828 gnd.n1973 256.663
R3514 gnd.n2821 gnd.n1973 256.663
R3515 gnd.n2819 gnd.n1973 256.663
R3516 gnd.n2813 gnd.n1973 256.663
R3517 gnd.n2811 gnd.n1973 256.663
R3518 gnd.n2805 gnd.n1973 256.663
R3519 gnd.n2803 gnd.n1973 256.663
R3520 gnd.n2797 gnd.n1973 256.663
R3521 gnd.n2795 gnd.n1973 256.663
R3522 gnd.n2789 gnd.n1973 256.663
R3523 gnd.n2787 gnd.n1973 256.663
R3524 gnd.n2781 gnd.n1973 256.663
R3525 gnd.n2779 gnd.n1973 256.663
R3526 gnd.n2773 gnd.n1973 256.663
R3527 gnd.n2771 gnd.n1973 256.663
R3528 gnd.n2765 gnd.n1973 256.663
R3529 gnd.n3714 gnd.n3627 256.663
R3530 gnd.n3714 gnd.n3628 256.663
R3531 gnd.n3714 gnd.n3629 256.663
R3532 gnd.n3714 gnd.n3630 256.663
R3533 gnd.n3714 gnd.n3631 256.663
R3534 gnd.n3714 gnd.n3632 256.663
R3535 gnd.n3714 gnd.n3633 256.663
R3536 gnd.n3714 gnd.n3634 256.663
R3537 gnd.n3714 gnd.n3635 256.663
R3538 gnd.n3714 gnd.n3636 256.663
R3539 gnd.n3714 gnd.n3637 256.663
R3540 gnd.n3714 gnd.n3638 256.663
R3541 gnd.n3714 gnd.n3639 256.663
R3542 gnd.n3714 gnd.n3640 256.663
R3543 gnd.n3714 gnd.n3641 256.663
R3544 gnd.n3714 gnd.n3642 256.663
R3545 gnd.n3643 gnd.n1331 256.663
R3546 gnd.n3714 gnd.n3626 256.663
R3547 gnd.n3714 gnd.n3558 256.663
R3548 gnd.n3714 gnd.n3557 256.663
R3549 gnd.n3714 gnd.n3556 256.663
R3550 gnd.n3714 gnd.n3555 256.663
R3551 gnd.n3714 gnd.n3554 256.663
R3552 gnd.n3714 gnd.n3553 256.663
R3553 gnd.n3714 gnd.n3552 256.663
R3554 gnd.n3714 gnd.n3551 256.663
R3555 gnd.n3714 gnd.n3550 256.663
R3556 gnd.n3714 gnd.n3549 256.663
R3557 gnd.n3714 gnd.n3548 256.663
R3558 gnd.n3714 gnd.n3547 256.663
R3559 gnd.n3714 gnd.n3546 256.663
R3560 gnd.n3714 gnd.n3545 256.663
R3561 gnd.n3714 gnd.n3544 256.663
R3562 gnd.n3714 gnd.n3543 256.663
R3563 gnd.n4574 gnd.n896 242.672
R3564 gnd.n4574 gnd.n897 242.672
R3565 gnd.n4574 gnd.n898 242.672
R3566 gnd.n4574 gnd.n899 242.672
R3567 gnd.n4574 gnd.n900 242.672
R3568 gnd.n4574 gnd.n901 242.672
R3569 gnd.n4574 gnd.n902 242.672
R3570 gnd.n4574 gnd.n903 242.672
R3571 gnd.n4574 gnd.n904 242.672
R3572 gnd.n2863 gnd.n2862 242.672
R3573 gnd.n2862 gnd.n2117 242.672
R3574 gnd.n2862 gnd.n2025 242.672
R3575 gnd.n2862 gnd.n2024 242.672
R3576 gnd.n2862 gnd.n2023 242.672
R3577 gnd.n2862 gnd.n2022 242.672
R3578 gnd.n2862 gnd.n2021 242.672
R3579 gnd.n2862 gnd.n2020 242.672
R3580 gnd.n2862 gnd.n2019 242.672
R3581 gnd.n4229 gnd.n1301 242.672
R3582 gnd.n4229 gnd.n1302 242.672
R3583 gnd.n4229 gnd.n1303 242.672
R3584 gnd.n4229 gnd.n1304 242.672
R3585 gnd.n4229 gnd.n1305 242.672
R3586 gnd.n4229 gnd.n1306 242.672
R3587 gnd.n4229 gnd.n1307 242.672
R3588 gnd.n4229 gnd.n1308 242.672
R3589 gnd.n4229 gnd.n1309 242.672
R3590 gnd.n6835 gnd.n94 242.672
R3591 gnd.n6831 gnd.n94 242.672
R3592 gnd.n6826 gnd.n94 242.672
R3593 gnd.n6823 gnd.n94 242.672
R3594 gnd.n6818 gnd.n94 242.672
R3595 gnd.n6815 gnd.n94 242.672
R3596 gnd.n6810 gnd.n94 242.672
R3597 gnd.n6807 gnd.n94 242.672
R3598 gnd.n6802 gnd.n94 242.672
R3599 gnd.n5036 gnd.n4945 242.672
R3600 gnd.n4949 gnd.n4945 242.672
R3601 gnd.n5029 gnd.n4945 242.672
R3602 gnd.n5023 gnd.n4945 242.672
R3603 gnd.n5021 gnd.n4945 242.672
R3604 gnd.n5015 gnd.n4945 242.672
R3605 gnd.n5013 gnd.n4945 242.672
R3606 gnd.n5007 gnd.n4945 242.672
R3607 gnd.n5005 gnd.n4945 242.672
R3608 gnd.n4999 gnd.n4945 242.672
R3609 gnd.n4997 gnd.n4945 242.672
R3610 gnd.n4990 gnd.n4945 242.672
R3611 gnd.n4988 gnd.n4945 242.672
R3612 gnd.n5914 gnd.n877 242.672
R3613 gnd.n5914 gnd.n876 242.672
R3614 gnd.n5914 gnd.n875 242.672
R3615 gnd.n5914 gnd.n874 242.672
R3616 gnd.n5914 gnd.n873 242.672
R3617 gnd.n5914 gnd.n872 242.672
R3618 gnd.n5914 gnd.n871 242.672
R3619 gnd.n5914 gnd.n870 242.672
R3620 gnd.n5914 gnd.n869 242.672
R3621 gnd.n5914 gnd.n868 242.672
R3622 gnd.n5914 gnd.n867 242.672
R3623 gnd.n5914 gnd.n866 242.672
R3624 gnd.n5914 gnd.n865 242.672
R3625 gnd.n5165 gnd.n5164 242.672
R3626 gnd.n5165 gnd.n5106 242.672
R3627 gnd.n5165 gnd.n5107 242.672
R3628 gnd.n5165 gnd.n5108 242.672
R3629 gnd.n5165 gnd.n5109 242.672
R3630 gnd.n5165 gnd.n5110 242.672
R3631 gnd.n5165 gnd.n5111 242.672
R3632 gnd.n5165 gnd.n5112 242.672
R3633 gnd.n5914 gnd.n4575 242.672
R3634 gnd.n5914 gnd.n4576 242.672
R3635 gnd.n5914 gnd.n4577 242.672
R3636 gnd.n5914 gnd.n4578 242.672
R3637 gnd.n5914 gnd.n4579 242.672
R3638 gnd.n5914 gnd.n4580 242.672
R3639 gnd.n5914 gnd.n4581 242.672
R3640 gnd.n5914 gnd.n5913 242.672
R3641 gnd.n4574 gnd.n4573 242.672
R3642 gnd.n4574 gnd.n878 242.672
R3643 gnd.n4574 gnd.n879 242.672
R3644 gnd.n4574 gnd.n880 242.672
R3645 gnd.n4574 gnd.n881 242.672
R3646 gnd.n4574 gnd.n882 242.672
R3647 gnd.n4574 gnd.n883 242.672
R3648 gnd.n4574 gnd.n884 242.672
R3649 gnd.n4574 gnd.n885 242.672
R3650 gnd.n4574 gnd.n886 242.672
R3651 gnd.n4574 gnd.n887 242.672
R3652 gnd.n4574 gnd.n888 242.672
R3653 gnd.n4574 gnd.n889 242.672
R3654 gnd.n4574 gnd.n890 242.672
R3655 gnd.n4574 gnd.n891 242.672
R3656 gnd.n4574 gnd.n892 242.672
R3657 gnd.n4574 gnd.n893 242.672
R3658 gnd.n4574 gnd.n894 242.672
R3659 gnd.n4574 gnd.n895 242.672
R3660 gnd.n2862 gnd.n2119 242.672
R3661 gnd.n2862 gnd.n2120 242.672
R3662 gnd.n2862 gnd.n2121 242.672
R3663 gnd.n2862 gnd.n2122 242.672
R3664 gnd.n2862 gnd.n2123 242.672
R3665 gnd.n2862 gnd.n2124 242.672
R3666 gnd.n2862 gnd.n2125 242.672
R3667 gnd.n2862 gnd.n2126 242.672
R3668 gnd.n2862 gnd.n2127 242.672
R3669 gnd.n2862 gnd.n2128 242.672
R3670 gnd.n2862 gnd.n2129 242.672
R3671 gnd.n2833 gnd.n2160 242.672
R3672 gnd.n2862 gnd.n2130 242.672
R3673 gnd.n2862 gnd.n2131 242.672
R3674 gnd.n2862 gnd.n2132 242.672
R3675 gnd.n2862 gnd.n2133 242.672
R3676 gnd.n2862 gnd.n2134 242.672
R3677 gnd.n2862 gnd.n2135 242.672
R3678 gnd.n2862 gnd.n2136 242.672
R3679 gnd.n2862 gnd.n2861 242.672
R3680 gnd.n4229 gnd.n4228 242.672
R3681 gnd.n4229 gnd.n1283 242.672
R3682 gnd.n4229 gnd.n1284 242.672
R3683 gnd.n4229 gnd.n1285 242.672
R3684 gnd.n4229 gnd.n1286 242.672
R3685 gnd.n4229 gnd.n1287 242.672
R3686 gnd.n4229 gnd.n1288 242.672
R3687 gnd.n4229 gnd.n1289 242.672
R3688 gnd.n4197 gnd.n1332 242.672
R3689 gnd.n4229 gnd.n1290 242.672
R3690 gnd.n4229 gnd.n1291 242.672
R3691 gnd.n4229 gnd.n1292 242.672
R3692 gnd.n4229 gnd.n1293 242.672
R3693 gnd.n4229 gnd.n1294 242.672
R3694 gnd.n4229 gnd.n1295 242.672
R3695 gnd.n4229 gnd.n1296 242.672
R3696 gnd.n4229 gnd.n1297 242.672
R3697 gnd.n4229 gnd.n1298 242.672
R3698 gnd.n4229 gnd.n1299 242.672
R3699 gnd.n4229 gnd.n1300 242.672
R3700 gnd.n154 gnd.n94 242.672
R3701 gnd.n6893 gnd.n94 242.672
R3702 gnd.n150 gnd.n94 242.672
R3703 gnd.n6900 gnd.n94 242.672
R3704 gnd.n143 gnd.n94 242.672
R3705 gnd.n6907 gnd.n94 242.672
R3706 gnd.n136 gnd.n94 242.672
R3707 gnd.n6914 gnd.n94 242.672
R3708 gnd.n129 gnd.n94 242.672
R3709 gnd.n6921 gnd.n94 242.672
R3710 gnd.n122 gnd.n94 242.672
R3711 gnd.n6931 gnd.n94 242.672
R3712 gnd.n115 gnd.n94 242.672
R3713 gnd.n6938 gnd.n94 242.672
R3714 gnd.n108 gnd.n94 242.672
R3715 gnd.n6945 gnd.n94 242.672
R3716 gnd.n101 gnd.n94 242.672
R3717 gnd.n6952 gnd.n94 242.672
R3718 gnd.n94 gnd.n93 242.672
R3719 gnd.n2900 gnd.n1986 242.672
R3720 gnd.n2900 gnd.n1987 242.672
R3721 gnd.n2900 gnd.n1988 242.672
R3722 gnd.n2900 gnd.n1989 242.672
R3723 gnd.n2900 gnd.n1990 242.672
R3724 gnd.n2900 gnd.n1991 242.672
R3725 gnd.n2900 gnd.n1992 242.672
R3726 gnd.n2900 gnd.n1993 242.672
R3727 gnd.n2900 gnd.n1994 242.672
R3728 gnd.n2900 gnd.n1995 242.672
R3729 gnd.n2900 gnd.n1996 242.672
R3730 gnd.n2900 gnd.n1997 242.672
R3731 gnd.n2900 gnd.n1998 242.672
R3732 gnd.n2900 gnd.n2899 242.672
R3733 gnd.n3891 gnd.n1275 242.672
R3734 gnd.n1638 gnd.n1275 242.672
R3735 gnd.n1635 gnd.n1275 242.672
R3736 gnd.n1630 gnd.n1275 242.672
R3737 gnd.n1627 gnd.n1275 242.672
R3738 gnd.n1624 gnd.n1275 242.672
R3739 gnd.n1611 gnd.n1275 242.672
R3740 gnd.n1609 gnd.n1275 242.672
R3741 gnd.n1594 gnd.n1275 242.672
R3742 gnd.n1592 gnd.n1275 242.672
R3743 gnd.n1577 gnd.n1275 242.672
R3744 gnd.n1575 gnd.n1275 242.672
R3745 gnd.n1560 gnd.n1275 242.672
R3746 gnd.n1558 gnd.n1275 242.672
R3747 gnd.n90 gnd.n86 240.244
R3748 gnd.n6954 gnd.n6953 240.244
R3749 gnd.n6951 gnd.n95 240.244
R3750 gnd.n6947 gnd.n6946 240.244
R3751 gnd.n6944 gnd.n102 240.244
R3752 gnd.n6940 gnd.n6939 240.244
R3753 gnd.n6937 gnd.n109 240.244
R3754 gnd.n6933 gnd.n6932 240.244
R3755 gnd.n6930 gnd.n116 240.244
R3756 gnd.n6923 gnd.n6922 240.244
R3757 gnd.n6920 gnd.n123 240.244
R3758 gnd.n6916 gnd.n6915 240.244
R3759 gnd.n6913 gnd.n130 240.244
R3760 gnd.n6909 gnd.n6908 240.244
R3761 gnd.n6906 gnd.n137 240.244
R3762 gnd.n6902 gnd.n6901 240.244
R3763 gnd.n6899 gnd.n144 240.244
R3764 gnd.n6895 gnd.n6894 240.244
R3765 gnd.n6892 gnd.n151 240.244
R3766 gnd.n4154 gnd.n1360 240.244
R3767 gnd.n3955 gnd.n1360 240.244
R3768 gnd.n3955 gnd.n1496 240.244
R3769 gnd.n3951 gnd.n1496 240.244
R3770 gnd.n3951 gnd.n1488 240.244
R3771 gnd.n1488 gnd.n1479 240.244
R3772 gnd.n3947 gnd.n1479 240.244
R3773 gnd.n3947 gnd.n1470 240.244
R3774 gnd.n3943 gnd.n1470 240.244
R3775 gnd.n3943 gnd.n1462 240.244
R3776 gnd.n1462 gnd.n1454 240.244
R3777 gnd.n3937 gnd.n1454 240.244
R3778 gnd.n3937 gnd.n1444 240.244
R3779 gnd.n3933 gnd.n1444 240.244
R3780 gnd.n3933 gnd.n1421 240.244
R3781 gnd.n4076 gnd.n1421 240.244
R3782 gnd.n4076 gnd.n1416 240.244
R3783 gnd.n4072 gnd.n1416 240.244
R3784 gnd.n4072 gnd.n1407 240.244
R3785 gnd.n1429 gnd.n1407 240.244
R3786 gnd.n1429 gnd.n1403 240.244
R3787 gnd.n1403 gnd.n233 240.244
R3788 gnd.n6738 gnd.n233 240.244
R3789 gnd.n6738 gnd.n230 240.244
R3790 gnd.n6734 gnd.n230 240.244
R3791 gnd.n6734 gnd.n222 240.244
R3792 gnd.n6729 gnd.n222 240.244
R3793 gnd.n6729 gnd.n208 240.244
R3794 gnd.n269 gnd.n208 240.244
R3795 gnd.n269 gnd.n202 240.244
R3796 gnd.n264 gnd.n202 240.244
R3797 gnd.n264 gnd.n195 240.244
R3798 gnd.n261 gnd.n195 240.244
R3799 gnd.n261 gnd.n187 240.244
R3800 gnd.n258 gnd.n187 240.244
R3801 gnd.n258 gnd.n179 240.244
R3802 gnd.n255 gnd.n179 240.244
R3803 gnd.n255 gnd.n171 240.244
R3804 gnd.n171 gnd.n161 240.244
R3805 gnd.n6883 gnd.n161 240.244
R3806 gnd.n6884 gnd.n6883 240.244
R3807 gnd.n6884 gnd.n82 240.244
R3808 gnd.n1313 gnd.n1312 240.244
R3809 gnd.n4222 gnd.n1312 240.244
R3810 gnd.n4220 gnd.n4219 240.244
R3811 gnd.n4216 gnd.n4215 240.244
R3812 gnd.n4212 gnd.n4211 240.244
R3813 gnd.n4208 gnd.n4207 240.244
R3814 gnd.n4204 gnd.n4203 240.244
R3815 gnd.n4200 gnd.n4199 240.244
R3816 gnd.n4195 gnd.n4194 240.244
R3817 gnd.n4191 gnd.n4190 240.244
R3818 gnd.n4187 gnd.n4186 240.244
R3819 gnd.n4183 gnd.n4182 240.244
R3820 gnd.n4179 gnd.n4178 240.244
R3821 gnd.n4175 gnd.n4174 240.244
R3822 gnd.n4171 gnd.n4170 240.244
R3823 gnd.n4167 gnd.n4166 240.244
R3824 gnd.n4163 gnd.n4162 240.244
R3825 gnd.n1355 gnd.n1354 240.244
R3826 gnd.n3975 gnd.n1314 240.244
R3827 gnd.n3975 gnd.n1498 240.244
R3828 gnd.n3983 gnd.n1498 240.244
R3829 gnd.n3983 gnd.n1499 240.244
R3830 gnd.n1499 gnd.n1477 240.244
R3831 gnd.n4007 gnd.n1477 240.244
R3832 gnd.n4007 gnd.n1472 240.244
R3833 gnd.n4015 gnd.n1472 240.244
R3834 gnd.n4015 gnd.n1473 240.244
R3835 gnd.n1473 gnd.n1452 240.244
R3836 gnd.n4041 gnd.n1452 240.244
R3837 gnd.n4041 gnd.n1447 240.244
R3838 gnd.n4050 gnd.n1447 240.244
R3839 gnd.n4050 gnd.n1448 240.244
R3840 gnd.n1448 gnd.n1418 240.244
R3841 gnd.n4078 gnd.n1418 240.244
R3842 gnd.n4081 gnd.n4078 240.244
R3843 gnd.n4081 gnd.n1405 240.244
R3844 gnd.n4092 gnd.n1405 240.244
R3845 gnd.n4095 gnd.n4092 240.244
R3846 gnd.n4098 gnd.n4095 240.244
R3847 gnd.n4098 gnd.n232 240.244
R3848 gnd.n6740 gnd.n232 240.244
R3849 gnd.n6743 gnd.n6740 240.244
R3850 gnd.n6743 gnd.n220 240.244
R3851 gnd.n6753 gnd.n220 240.244
R3852 gnd.n6753 gnd.n210 240.244
R3853 gnd.n6759 gnd.n210 240.244
R3854 gnd.n6759 gnd.n200 240.244
R3855 gnd.n6769 gnd.n200 240.244
R3856 gnd.n6769 gnd.n196 240.244
R3857 gnd.n6775 gnd.n196 240.244
R3858 gnd.n6775 gnd.n184 240.244
R3859 gnd.n6785 gnd.n184 240.244
R3860 gnd.n6785 gnd.n180 240.244
R3861 gnd.n6791 gnd.n180 240.244
R3862 gnd.n6791 gnd.n168 240.244
R3863 gnd.n6875 gnd.n168 240.244
R3864 gnd.n6875 gnd.n164 240.244
R3865 gnd.n6881 gnd.n164 240.244
R3866 gnd.n6881 gnd.n85 240.244
R3867 gnd.n6961 gnd.n85 240.244
R3868 gnd.n2137 gnd.n1158 240.244
R3869 gnd.n2860 gnd.n2138 240.244
R3870 gnd.n2856 gnd.n2855 240.244
R3871 gnd.n2852 gnd.n2851 240.244
R3872 gnd.n2848 gnd.n2847 240.244
R3873 gnd.n2844 gnd.n2843 240.244
R3874 gnd.n2840 gnd.n2839 240.244
R3875 gnd.n2836 gnd.n2835 240.244
R3876 gnd.n2621 gnd.n2620 240.244
R3877 gnd.n2618 gnd.n2617 240.244
R3878 gnd.n2614 gnd.n2613 240.244
R3879 gnd.n2610 gnd.n2609 240.244
R3880 gnd.n2606 gnd.n2605 240.244
R3881 gnd.n2602 gnd.n2601 240.244
R3882 gnd.n2598 gnd.n2597 240.244
R3883 gnd.n2594 gnd.n2593 240.244
R3884 gnd.n2590 gnd.n2589 240.244
R3885 gnd.n2586 gnd.n2585 240.244
R3886 gnd.n4495 gnd.n954 240.244
R3887 gnd.n958 gnd.n954 240.244
R3888 gnd.n4488 gnd.n958 240.244
R3889 gnd.n4488 gnd.n959 240.244
R3890 gnd.n972 gnd.n959 240.244
R3891 gnd.n2338 gnd.n972 240.244
R3892 gnd.n2338 gnd.n983 240.244
R3893 gnd.n2341 gnd.n983 240.244
R3894 gnd.n2341 gnd.n993 240.244
R3895 gnd.n2346 gnd.n993 240.244
R3896 gnd.n2346 gnd.n1003 240.244
R3897 gnd.n2462 gnd.n1003 240.244
R3898 gnd.n2462 gnd.n1014 240.244
R3899 gnd.n2470 gnd.n1014 240.244
R3900 gnd.n2470 gnd.n1025 240.244
R3901 gnd.n2225 gnd.n1025 240.244
R3902 gnd.n2481 gnd.n2225 240.244
R3903 gnd.n2481 gnd.n1036 240.244
R3904 gnd.n2487 gnd.n1036 240.244
R3905 gnd.n2487 gnd.n1050 240.244
R3906 gnd.n2497 gnd.n1050 240.244
R3907 gnd.n2497 gnd.n1058 240.244
R3908 gnd.n2503 gnd.n1058 240.244
R3909 gnd.n2503 gnd.n1067 240.244
R3910 gnd.n2513 gnd.n1067 240.244
R3911 gnd.n2513 gnd.n1075 240.244
R3912 gnd.n2519 gnd.n1075 240.244
R3913 gnd.n2519 gnd.n1086 240.244
R3914 gnd.n2529 gnd.n1086 240.244
R3915 gnd.n2529 gnd.n1097 240.244
R3916 gnd.n2535 gnd.n1097 240.244
R3917 gnd.n2535 gnd.n1107 240.244
R3918 gnd.n2545 gnd.n1107 240.244
R3919 gnd.n2545 gnd.n1118 240.244
R3920 gnd.n2551 gnd.n1118 240.244
R3921 gnd.n2551 gnd.n1129 240.244
R3922 gnd.n2561 gnd.n1129 240.244
R3923 gnd.n2561 gnd.n1140 240.244
R3924 gnd.n2568 gnd.n1140 240.244
R3925 gnd.n2568 gnd.n1151 240.244
R3926 gnd.n2578 gnd.n1151 240.244
R3927 gnd.n2578 gnd.n1160 240.244
R3928 gnd.n908 gnd.n907 240.244
R3929 gnd.n4567 gnd.n907 240.244
R3930 gnd.n4565 gnd.n4564 240.244
R3931 gnd.n4561 gnd.n4560 240.244
R3932 gnd.n4557 gnd.n4556 240.244
R3933 gnd.n4553 gnd.n4552 240.244
R3934 gnd.n4549 gnd.n4548 240.244
R3935 gnd.n4545 gnd.n4544 240.244
R3936 gnd.n4541 gnd.n4540 240.244
R3937 gnd.n4536 gnd.n4535 240.244
R3938 gnd.n4532 gnd.n4531 240.244
R3939 gnd.n4528 gnd.n4527 240.244
R3940 gnd.n4524 gnd.n4523 240.244
R3941 gnd.n4520 gnd.n4519 240.244
R3942 gnd.n4516 gnd.n4515 240.244
R3943 gnd.n4512 gnd.n4511 240.244
R3944 gnd.n4508 gnd.n4507 240.244
R3945 gnd.n4504 gnd.n4503 240.244
R3946 gnd.n949 gnd.n948 240.244
R3947 gnd.n2434 gnd.n909 240.244
R3948 gnd.n2434 gnd.n964 240.244
R3949 gnd.n4486 gnd.n964 240.244
R3950 gnd.n4486 gnd.n965 240.244
R3951 gnd.n4482 gnd.n965 240.244
R3952 gnd.n4482 gnd.n971 240.244
R3953 gnd.n4474 gnd.n971 240.244
R3954 gnd.n4474 gnd.n986 240.244
R3955 gnd.n4470 gnd.n986 240.244
R3956 gnd.n4470 gnd.n992 240.244
R3957 gnd.n4462 gnd.n992 240.244
R3958 gnd.n4462 gnd.n1006 240.244
R3959 gnd.n4458 gnd.n1006 240.244
R3960 gnd.n4458 gnd.n1012 240.244
R3961 gnd.n4450 gnd.n1012 240.244
R3962 gnd.n4450 gnd.n1028 240.244
R3963 gnd.n1032 gnd.n1028 240.244
R3964 gnd.n4444 gnd.n1032 240.244
R3965 gnd.n4444 gnd.n1034 240.244
R3966 gnd.n4436 gnd.n1034 240.244
R3967 gnd.n4436 gnd.n1053 240.244
R3968 gnd.n4431 gnd.n1053 240.244
R3969 gnd.n4431 gnd.n1056 240.244
R3970 gnd.n4423 gnd.n1056 240.244
R3971 gnd.n4423 gnd.n1070 240.244
R3972 gnd.n4418 gnd.n1070 240.244
R3973 gnd.n4418 gnd.n1073 240.244
R3974 gnd.n4410 gnd.n1073 240.244
R3975 gnd.n4410 gnd.n1089 240.244
R3976 gnd.n4406 gnd.n1089 240.244
R3977 gnd.n4406 gnd.n1095 240.244
R3978 gnd.n4398 gnd.n1095 240.244
R3979 gnd.n4398 gnd.n1110 240.244
R3980 gnd.n4394 gnd.n1110 240.244
R3981 gnd.n4394 gnd.n1116 240.244
R3982 gnd.n4386 gnd.n1116 240.244
R3983 gnd.n4386 gnd.n1132 240.244
R3984 gnd.n4382 gnd.n1132 240.244
R3985 gnd.n4382 gnd.n1138 240.244
R3986 gnd.n4374 gnd.n1138 240.244
R3987 gnd.n4374 gnd.n1153 240.244
R3988 gnd.n4370 gnd.n1153 240.244
R3989 gnd.n5915 gnd.n862 240.244
R3990 gnd.n5912 gnd.n4582 240.244
R3991 gnd.n5908 gnd.n5907 240.244
R3992 gnd.n5904 gnd.n5903 240.244
R3993 gnd.n5900 gnd.n5899 240.244
R3994 gnd.n5896 gnd.n5895 240.244
R3995 gnd.n5892 gnd.n5891 240.244
R3996 gnd.n5888 gnd.n5887 240.244
R3997 gnd.n5177 gnd.n4897 240.244
R3998 gnd.n4897 gnd.n4888 240.244
R3999 gnd.n5195 gnd.n4888 240.244
R4000 gnd.n5196 gnd.n5195 240.244
R4001 gnd.n5196 gnd.n4876 240.244
R4002 gnd.n4876 gnd.n4865 240.244
R4003 gnd.n5227 gnd.n4865 240.244
R4004 gnd.n5228 gnd.n5227 240.244
R4005 gnd.n5229 gnd.n5228 240.244
R4006 gnd.n5229 gnd.n4850 240.244
R4007 gnd.n5231 gnd.n4850 240.244
R4008 gnd.n5231 gnd.n4835 240.244
R4009 gnd.n5272 gnd.n4835 240.244
R4010 gnd.n5273 gnd.n5272 240.244
R4011 gnd.n5276 gnd.n5273 240.244
R4012 gnd.n5276 gnd.n4817 240.244
R4013 gnd.n5308 gnd.n4817 240.244
R4014 gnd.n5308 gnd.n4803 240.244
R4015 gnd.n5330 gnd.n4803 240.244
R4016 gnd.n5331 gnd.n5330 240.244
R4017 gnd.n5331 gnd.n4790 240.244
R4018 gnd.n4790 gnd.n4779 240.244
R4019 gnd.n5362 gnd.n4779 240.244
R4020 gnd.n5363 gnd.n5362 240.244
R4021 gnd.n5364 gnd.n5363 240.244
R4022 gnd.n5364 gnd.n4728 240.244
R4023 gnd.n4728 gnd.n4727 240.244
R4024 gnd.n4727 gnd.n4712 240.244
R4025 gnd.n5415 gnd.n4712 240.244
R4026 gnd.n5416 gnd.n5415 240.244
R4027 gnd.n5416 gnd.n4699 240.244
R4028 gnd.n4699 gnd.n4688 240.244
R4029 gnd.n5449 gnd.n4688 240.244
R4030 gnd.n5450 gnd.n5449 240.244
R4031 gnd.n5452 gnd.n5450 240.244
R4032 gnd.n5452 gnd.n5451 240.244
R4033 gnd.n5451 gnd.n4667 240.244
R4034 gnd.n5487 gnd.n4667 240.244
R4035 gnd.n5487 gnd.n4659 240.244
R4036 gnd.n4659 gnd.n4652 240.244
R4037 gnd.n5512 gnd.n4652 240.244
R4038 gnd.n5512 gnd.n805 240.244
R4039 gnd.n5525 gnd.n805 240.244
R4040 gnd.n5525 gnd.n815 240.244
R4041 gnd.n4640 gnd.n815 240.244
R4042 gnd.n5545 gnd.n4640 240.244
R4043 gnd.n5545 gnd.n827 240.244
R4044 gnd.n4635 gnd.n827 240.244
R4045 gnd.n4635 gnd.n840 240.244
R4046 gnd.n4633 gnd.n840 240.244
R4047 gnd.n5820 gnd.n4633 240.244
R4048 gnd.n5820 gnd.n852 240.244
R4049 gnd.n5816 gnd.n852 240.244
R4050 gnd.n5114 gnd.n5113 240.244
R4051 gnd.n5158 gnd.n5113 240.244
R4052 gnd.n5156 gnd.n5155 240.244
R4053 gnd.n5152 gnd.n5151 240.244
R4054 gnd.n5148 gnd.n5147 240.244
R4055 gnd.n5144 gnd.n5143 240.244
R4056 gnd.n5140 gnd.n5139 240.244
R4057 gnd.n5136 gnd.n5135 240.244
R4058 gnd.n5187 gnd.n4895 240.244
R4059 gnd.n5187 gnd.n4891 240.244
R4060 gnd.n5193 gnd.n4891 240.244
R4061 gnd.n5193 gnd.n4874 240.244
R4062 gnd.n5217 gnd.n4874 240.244
R4063 gnd.n5217 gnd.n4869 240.244
R4064 gnd.n5225 gnd.n4869 240.244
R4065 gnd.n5225 gnd.n4870 240.244
R4066 gnd.n4870 gnd.n4848 240.244
R4067 gnd.n5251 gnd.n4848 240.244
R4068 gnd.n5251 gnd.n4843 240.244
R4069 gnd.n5262 gnd.n4843 240.244
R4070 gnd.n5262 gnd.n4844 240.244
R4071 gnd.n5258 gnd.n4844 240.244
R4072 gnd.n5258 gnd.n4815 240.244
R4073 gnd.n5312 gnd.n4815 240.244
R4074 gnd.n5312 gnd.n4810 240.244
R4075 gnd.n5320 gnd.n4810 240.244
R4076 gnd.n5320 gnd.n4811 240.244
R4077 gnd.n4811 gnd.n4788 240.244
R4078 gnd.n5352 gnd.n4788 240.244
R4079 gnd.n5352 gnd.n4783 240.244
R4080 gnd.n5360 gnd.n4783 240.244
R4081 gnd.n5360 gnd.n4784 240.244
R4082 gnd.n4784 gnd.n4725 240.244
R4083 gnd.n5397 gnd.n4725 240.244
R4084 gnd.n5397 gnd.n4720 240.244
R4085 gnd.n5405 gnd.n4720 240.244
R4086 gnd.n5405 gnd.n4721 240.244
R4087 gnd.n4721 gnd.n4697 240.244
R4088 gnd.n5436 gnd.n4697 240.244
R4089 gnd.n5436 gnd.n4692 240.244
R4090 gnd.n5447 gnd.n4692 240.244
R4091 gnd.n5447 gnd.n4693 240.244
R4092 gnd.n5443 gnd.n4693 240.244
R4093 gnd.n5443 gnd.n4666 240.244
R4094 gnd.n5491 gnd.n4666 240.244
R4095 gnd.n5491 gnd.n4661 240.244
R4096 gnd.n5500 gnd.n4661 240.244
R4097 gnd.n5500 gnd.n4662 240.244
R4098 gnd.n4662 gnd.n807 240.244
R4099 gnd.n5949 gnd.n807 240.244
R4100 gnd.n5949 gnd.n808 240.244
R4101 gnd.n5945 gnd.n808 240.244
R4102 gnd.n5945 gnd.n814 240.244
R4103 gnd.n829 gnd.n814 240.244
R4104 gnd.n5935 gnd.n829 240.244
R4105 gnd.n5935 gnd.n830 240.244
R4106 gnd.n5931 gnd.n830 240.244
R4107 gnd.n5931 gnd.n838 240.244
R4108 gnd.n854 gnd.n838 240.244
R4109 gnd.n5921 gnd.n854 240.244
R4110 gnd.n5921 gnd.n855 240.244
R4111 gnd.n4601 gnd.n864 240.244
R4112 gnd.n5878 gnd.n5877 240.244
R4113 gnd.n5874 gnd.n5873 240.244
R4114 gnd.n5870 gnd.n5869 240.244
R4115 gnd.n5866 gnd.n5865 240.244
R4116 gnd.n5862 gnd.n5861 240.244
R4117 gnd.n5858 gnd.n5857 240.244
R4118 gnd.n5854 gnd.n5853 240.244
R4119 gnd.n5850 gnd.n5849 240.244
R4120 gnd.n5846 gnd.n5845 240.244
R4121 gnd.n5842 gnd.n5841 240.244
R4122 gnd.n5838 gnd.n5837 240.244
R4123 gnd.n5834 gnd.n5833 240.244
R4124 gnd.n5045 gnd.n4941 240.244
R4125 gnd.n5051 gnd.n4941 240.244
R4126 gnd.n5051 gnd.n4933 240.244
R4127 gnd.n5061 gnd.n4933 240.244
R4128 gnd.n5061 gnd.n4929 240.244
R4129 gnd.n5067 gnd.n4929 240.244
R4130 gnd.n5067 gnd.n4920 240.244
R4131 gnd.n5077 gnd.n4920 240.244
R4132 gnd.n5077 gnd.n4915 240.244
R4133 gnd.n5105 gnd.n4915 240.244
R4134 gnd.n5105 gnd.n4916 240.244
R4135 gnd.n4916 gnd.n4908 240.244
R4136 gnd.n5100 gnd.n4908 240.244
R4137 gnd.n5100 gnd.n4898 240.244
R4138 gnd.n5097 gnd.n4898 240.244
R4139 gnd.n5097 gnd.n4887 240.244
R4140 gnd.n5094 gnd.n4887 240.244
R4141 gnd.n5094 gnd.n4877 240.244
R4142 gnd.n5091 gnd.n4877 240.244
R4143 gnd.n5091 gnd.n4855 240.244
R4144 gnd.n5240 gnd.n4855 240.244
R4145 gnd.n5240 gnd.n4851 240.244
R4146 gnd.n5248 gnd.n4851 240.244
R4147 gnd.n5248 gnd.n4841 240.244
R4148 gnd.n4841 gnd.n4822 240.244
R4149 gnd.n5287 gnd.n4822 240.244
R4150 gnd.n5287 gnd.n4823 240.244
R4151 gnd.n4823 gnd.n4818 240.244
R4152 gnd.n5307 gnd.n4818 240.244
R4153 gnd.n5307 gnd.n4808 240.244
R4154 gnd.n5302 gnd.n4808 240.244
R4155 gnd.n5302 gnd.n4802 240.244
R4156 gnd.n5298 gnd.n4802 240.244
R4157 gnd.n5298 gnd.n4791 240.244
R4158 gnd.n5294 gnd.n4791 240.244
R4159 gnd.n5294 gnd.n4769 240.244
R4160 gnd.n5373 gnd.n4769 240.244
R4161 gnd.n5373 gnd.n4729 240.244
R4162 gnd.n5394 gnd.n4729 240.244
R4163 gnd.n5394 gnd.n4718 240.244
R4164 gnd.n5390 gnd.n4718 240.244
R4165 gnd.n5390 gnd.n4711 240.244
R4166 gnd.n5387 gnd.n4711 240.244
R4167 gnd.n5387 gnd.n4700 240.244
R4168 gnd.n5384 gnd.n4700 240.244
R4169 gnd.n5384 gnd.n4678 240.244
R4170 gnd.n5459 gnd.n4678 240.244
R4171 gnd.n5459 gnd.n4674 240.244
R4172 gnd.n5477 gnd.n4674 240.244
R4173 gnd.n5477 gnd.n4668 240.244
R4174 gnd.n4668 gnd.n4658 240.244
R4175 gnd.n5472 gnd.n4658 240.244
R4176 gnd.n5472 gnd.n4651 240.244
R4177 gnd.n5469 gnd.n4651 240.244
R4178 gnd.n5469 gnd.n4644 240.244
R4179 gnd.n5528 gnd.n4644 240.244
R4180 gnd.n5528 gnd.n816 240.244
R4181 gnd.n5542 gnd.n816 240.244
R4182 gnd.n5542 gnd.n826 240.244
R4183 gnd.n5538 gnd.n826 240.244
R4184 gnd.n5538 gnd.n5537 240.244
R4185 gnd.n5537 gnd.n841 240.244
R4186 gnd.n5823 gnd.n841 240.244
R4187 gnd.n5823 gnd.n851 240.244
R4188 gnd.n5829 gnd.n851 240.244
R4189 gnd.n5037 gnd.n5035 240.244
R4190 gnd.n5035 gnd.n5034 240.244
R4191 gnd.n5031 gnd.n5030 240.244
R4192 gnd.n5028 gnd.n4954 240.244
R4193 gnd.n5024 gnd.n5022 240.244
R4194 gnd.n5020 gnd.n4960 240.244
R4195 gnd.n5016 gnd.n5014 240.244
R4196 gnd.n5012 gnd.n4966 240.244
R4197 gnd.n5008 gnd.n5006 240.244
R4198 gnd.n5004 gnd.n4972 240.244
R4199 gnd.n5000 gnd.n4998 240.244
R4200 gnd.n4996 gnd.n4978 240.244
R4201 gnd.n4991 gnd.n4989 240.244
R4202 gnd.n5043 gnd.n4939 240.244
R4203 gnd.n5053 gnd.n4939 240.244
R4204 gnd.n5053 gnd.n4935 240.244
R4205 gnd.n5059 gnd.n4935 240.244
R4206 gnd.n5059 gnd.n4927 240.244
R4207 gnd.n5069 gnd.n4927 240.244
R4208 gnd.n5069 gnd.n4923 240.244
R4209 gnd.n5075 gnd.n4923 240.244
R4210 gnd.n5075 gnd.n4914 240.244
R4211 gnd.n5167 gnd.n4914 240.244
R4212 gnd.n5167 gnd.n4909 240.244
R4213 gnd.n5174 gnd.n4909 240.244
R4214 gnd.n5174 gnd.n4900 240.244
R4215 gnd.n5184 gnd.n4900 240.244
R4216 gnd.n5184 gnd.n4886 240.244
R4217 gnd.n5199 gnd.n4886 240.244
R4218 gnd.n5199 gnd.n4879 240.244
R4219 gnd.n5214 gnd.n4879 240.244
R4220 gnd.n5214 gnd.n4880 240.244
R4221 gnd.n4880 gnd.n4858 240.244
R4222 gnd.n5238 gnd.n4858 240.244
R4223 gnd.n5238 gnd.n4859 240.244
R4224 gnd.n4859 gnd.n4839 240.244
R4225 gnd.n5265 gnd.n4839 240.244
R4226 gnd.n5265 gnd.n4826 240.244
R4227 gnd.n5285 gnd.n4826 240.244
R4228 gnd.n5285 gnd.n4827 240.244
R4229 gnd.n5281 gnd.n4827 240.244
R4230 gnd.n5281 gnd.n4807 240.244
R4231 gnd.n5323 gnd.n4807 240.244
R4232 gnd.n5323 gnd.n4800 240.244
R4233 gnd.n5334 gnd.n4800 240.244
R4234 gnd.n5334 gnd.n4793 240.244
R4235 gnd.n5349 gnd.n4793 240.244
R4236 gnd.n5349 gnd.n4794 240.244
R4237 gnd.n4794 gnd.n4772 240.244
R4238 gnd.n5371 gnd.n4772 240.244
R4239 gnd.n5371 gnd.n4773 240.244
R4240 gnd.n4773 gnd.n4716 240.244
R4241 gnd.n5408 gnd.n4716 240.244
R4242 gnd.n5408 gnd.n4709 240.244
R4243 gnd.n5419 gnd.n4709 240.244
R4244 gnd.n5419 gnd.n4702 240.244
R4245 gnd.n5433 gnd.n4702 240.244
R4246 gnd.n5433 gnd.n4703 240.244
R4247 gnd.n4703 gnd.n4682 240.244
R4248 gnd.n5457 gnd.n4682 240.244
R4249 gnd.n5457 gnd.n4672 240.244
R4250 gnd.n5479 gnd.n4672 240.244
R4251 gnd.n5479 gnd.n4657 240.244
R4252 gnd.n5503 gnd.n4657 240.244
R4253 gnd.n5503 gnd.n4648 240.244
R4254 gnd.n5515 gnd.n4648 240.244
R4255 gnd.n5516 gnd.n5515 240.244
R4256 gnd.n5517 gnd.n5516 240.244
R4257 gnd.n5517 gnd.n818 240.244
R4258 gnd.n5942 gnd.n818 240.244
R4259 gnd.n5942 gnd.n819 240.244
R4260 gnd.n5938 gnd.n819 240.244
R4261 gnd.n5938 gnd.n825 240.244
R4262 gnd.n843 gnd.n825 240.244
R4263 gnd.n5928 gnd.n843 240.244
R4264 gnd.n5928 gnd.n844 240.244
R4265 gnd.n5924 gnd.n844 240.244
R4266 gnd.n5924 gnd.n850 240.244
R4267 gnd.n6801 gnd.n6800 240.244
R4268 gnd.n6806 gnd.n6803 240.244
R4269 gnd.n6809 gnd.n6808 240.244
R4270 gnd.n6814 gnd.n6811 240.244
R4271 gnd.n6817 gnd.n6816 240.244
R4272 gnd.n6822 gnd.n6819 240.244
R4273 gnd.n6825 gnd.n6824 240.244
R4274 gnd.n6830 gnd.n6827 240.244
R4275 gnd.n6836 gnd.n6832 240.244
R4276 gnd.n3916 gnd.n1363 240.244
R4277 gnd.n3916 gnd.n1494 240.244
R4278 gnd.n3985 gnd.n1494 240.244
R4279 gnd.n3985 gnd.n1489 240.244
R4280 gnd.n3992 gnd.n1489 240.244
R4281 gnd.n3992 gnd.n1480 240.244
R4282 gnd.n1480 gnd.n1468 240.244
R4283 gnd.n4017 gnd.n1468 240.244
R4284 gnd.n4017 gnd.n1463 240.244
R4285 gnd.n4024 gnd.n1463 240.244
R4286 gnd.n4024 gnd.n1455 240.244
R4287 gnd.n1455 gnd.n1442 240.244
R4288 gnd.n4052 gnd.n1442 240.244
R4289 gnd.n4052 gnd.n1438 240.244
R4290 gnd.n4058 gnd.n1438 240.244
R4291 gnd.n4058 gnd.n1414 240.244
R4292 gnd.n4083 gnd.n1414 240.244
R4293 gnd.n4083 gnd.n1408 240.244
R4294 gnd.n4089 gnd.n1408 240.244
R4295 gnd.n4089 gnd.n1409 240.244
R4296 gnd.n1409 gnd.n1404 240.244
R4297 gnd.n1404 gnd.n54 240.244
R4298 gnd.n55 gnd.n54 240.244
R4299 gnd.n56 gnd.n55 240.244
R4300 gnd.n6732 gnd.n56 240.244
R4301 gnd.n6732 gnd.n59 240.244
R4302 gnd.n60 gnd.n59 240.244
R4303 gnd.n61 gnd.n60 240.244
R4304 gnd.n267 gnd.n61 240.244
R4305 gnd.n267 gnd.n64 240.244
R4306 gnd.n65 gnd.n64 240.244
R4307 gnd.n66 gnd.n65 240.244
R4308 gnd.n185 gnd.n66 240.244
R4309 gnd.n185 gnd.n69 240.244
R4310 gnd.n70 gnd.n69 240.244
R4311 gnd.n71 gnd.n70 240.244
R4312 gnd.n169 gnd.n71 240.244
R4313 gnd.n169 gnd.n74 240.244
R4314 gnd.n75 gnd.n74 240.244
R4315 gnd.n76 gnd.n75 240.244
R4316 gnd.n79 gnd.n76 240.244
R4317 gnd.n6963 gnd.n79 240.244
R4318 gnd.n1553 gnd.n1552 240.244
R4319 gnd.n1544 gnd.n1543 240.244
R4320 gnd.n1569 gnd.n1568 240.244
R4321 gnd.n1535 gnd.n1534 240.244
R4322 gnd.n1586 gnd.n1585 240.244
R4323 gnd.n1526 gnd.n1525 240.244
R4324 gnd.n1603 gnd.n1602 240.244
R4325 gnd.n1517 gnd.n1516 240.244
R4326 gnd.n1512 gnd.n1310 240.244
R4327 gnd.n4152 gnd.n1366 240.244
R4328 gnd.n1370 gnd.n1366 240.244
R4329 gnd.n1371 gnd.n1370 240.244
R4330 gnd.n1372 gnd.n1371 240.244
R4331 gnd.n3993 gnd.n1372 240.244
R4332 gnd.n3993 gnd.n1375 240.244
R4333 gnd.n1376 gnd.n1375 240.244
R4334 gnd.n1377 gnd.n1376 240.244
R4335 gnd.n3941 gnd.n1377 240.244
R4336 gnd.n3941 gnd.n1380 240.244
R4337 gnd.n1381 gnd.n1380 240.244
R4338 gnd.n1382 gnd.n1381 240.244
R4339 gnd.n1446 gnd.n1382 240.244
R4340 gnd.n1446 gnd.n1385 240.244
R4341 gnd.n1386 gnd.n1385 240.244
R4342 gnd.n1387 gnd.n1386 240.244
R4343 gnd.n1417 gnd.n1387 240.244
R4344 gnd.n1417 gnd.n1390 240.244
R4345 gnd.n1391 gnd.n1390 240.244
R4346 gnd.n1392 gnd.n1391 240.244
R4347 gnd.n1396 gnd.n1392 240.244
R4348 gnd.n4116 gnd.n1396 240.244
R4349 gnd.n4116 gnd.n228 240.244
R4350 gnd.n6745 gnd.n228 240.244
R4351 gnd.n6745 gnd.n224 240.244
R4352 gnd.n6751 gnd.n224 240.244
R4353 gnd.n6751 gnd.n207 240.244
R4354 gnd.n6761 gnd.n207 240.244
R4355 gnd.n6761 gnd.n203 240.244
R4356 gnd.n6767 gnd.n203 240.244
R4357 gnd.n6767 gnd.n193 240.244
R4358 gnd.n6777 gnd.n193 240.244
R4359 gnd.n6777 gnd.n189 240.244
R4360 gnd.n6783 gnd.n189 240.244
R4361 gnd.n6783 gnd.n178 240.244
R4362 gnd.n6793 gnd.n178 240.244
R4363 gnd.n6793 gnd.n172 240.244
R4364 gnd.n6873 gnd.n172 240.244
R4365 gnd.n6873 gnd.n173 240.244
R4366 gnd.n173 gnd.n163 240.244
R4367 gnd.n6798 gnd.n163 240.244
R4368 gnd.n6798 gnd.n84 240.244
R4369 gnd.n2050 gnd.n1163 240.244
R4370 gnd.n2054 gnd.n2053 240.244
R4371 gnd.n2066 gnd.n2065 240.244
R4372 gnd.n2078 gnd.n2077 240.244
R4373 gnd.n2040 gnd.n2039 240.244
R4374 gnd.n2090 gnd.n2089 240.244
R4375 gnd.n2102 gnd.n2101 240.244
R4376 gnd.n2115 gnd.n2026 240.244
R4377 gnd.n2116 gnd.n2017 240.244
R4378 gnd.n2436 gnd.n2356 240.244
R4379 gnd.n2437 gnd.n2436 240.244
R4380 gnd.n2437 gnd.n961 240.244
R4381 gnd.n2442 gnd.n961 240.244
R4382 gnd.n2442 gnd.n973 240.244
R4383 gnd.n2445 gnd.n973 240.244
R4384 gnd.n2445 gnd.n984 240.244
R4385 gnd.n2450 gnd.n984 240.244
R4386 gnd.n2450 gnd.n994 240.244
R4387 gnd.n2453 gnd.n994 240.244
R4388 gnd.n2453 gnd.n1004 240.244
R4389 gnd.n2460 gnd.n1004 240.244
R4390 gnd.n2460 gnd.n1015 240.244
R4391 gnd.n2472 gnd.n1015 240.244
R4392 gnd.n2472 gnd.n1026 240.244
R4393 gnd.n2327 gnd.n1026 240.244
R4394 gnd.n2479 gnd.n2327 240.244
R4395 gnd.n2479 gnd.n1037 240.244
R4396 gnd.n2489 gnd.n1037 240.244
R4397 gnd.n2489 gnd.n1051 240.244
R4398 gnd.n2495 gnd.n1051 240.244
R4399 gnd.n2495 gnd.n1059 240.244
R4400 gnd.n2505 gnd.n1059 240.244
R4401 gnd.n2505 gnd.n1068 240.244
R4402 gnd.n2511 gnd.n1068 240.244
R4403 gnd.n2511 gnd.n1076 240.244
R4404 gnd.n2521 gnd.n1076 240.244
R4405 gnd.n2521 gnd.n1087 240.244
R4406 gnd.n2527 gnd.n1087 240.244
R4407 gnd.n2527 gnd.n1098 240.244
R4408 gnd.n2537 gnd.n1098 240.244
R4409 gnd.n2537 gnd.n1108 240.244
R4410 gnd.n2543 gnd.n1108 240.244
R4411 gnd.n2543 gnd.n1119 240.244
R4412 gnd.n2553 gnd.n1119 240.244
R4413 gnd.n2553 gnd.n1130 240.244
R4414 gnd.n2559 gnd.n1130 240.244
R4415 gnd.n2559 gnd.n1141 240.244
R4416 gnd.n2570 gnd.n1141 240.244
R4417 gnd.n2570 gnd.n1152 240.244
R4418 gnd.n2576 gnd.n1152 240.244
R4419 gnd.n2576 gnd.n1161 240.244
R4420 gnd.n2416 gnd.n2415 240.244
R4421 gnd.n2412 gnd.n2411 240.244
R4422 gnd.n2408 gnd.n2407 240.244
R4423 gnd.n2404 gnd.n2403 240.244
R4424 gnd.n2400 gnd.n2399 240.244
R4425 gnd.n2396 gnd.n2395 240.244
R4426 gnd.n2392 gnd.n2391 240.244
R4427 gnd.n2388 gnd.n2387 240.244
R4428 gnd.n2376 gnd.n905 240.244
R4429 gnd.n2428 gnd.n2357 240.244
R4430 gnd.n2428 gnd.n2358 240.244
R4431 gnd.n2358 gnd.n963 240.244
R4432 gnd.n975 gnd.n963 240.244
R4433 gnd.n4480 gnd.n975 240.244
R4434 gnd.n4480 gnd.n976 240.244
R4435 gnd.n4476 gnd.n976 240.244
R4436 gnd.n4476 gnd.n982 240.244
R4437 gnd.n4468 gnd.n982 240.244
R4438 gnd.n4468 gnd.n995 240.244
R4439 gnd.n4464 gnd.n995 240.244
R4440 gnd.n4464 gnd.n1001 240.244
R4441 gnd.n4456 gnd.n1001 240.244
R4442 gnd.n4456 gnd.n1017 240.244
R4443 gnd.n4452 gnd.n1017 240.244
R4444 gnd.n4452 gnd.n1023 240.244
R4445 gnd.n1039 gnd.n1023 240.244
R4446 gnd.n4442 gnd.n1039 240.244
R4447 gnd.n4442 gnd.n1040 240.244
R4448 gnd.n4438 gnd.n1040 240.244
R4449 gnd.n4438 gnd.n1048 240.244
R4450 gnd.n4429 gnd.n1048 240.244
R4451 gnd.n4429 gnd.n1060 240.244
R4452 gnd.n4425 gnd.n1060 240.244
R4453 gnd.n4425 gnd.n1065 240.244
R4454 gnd.n4416 gnd.n1065 240.244
R4455 gnd.n4416 gnd.n1078 240.244
R4456 gnd.n4412 gnd.n1078 240.244
R4457 gnd.n4412 gnd.n1084 240.244
R4458 gnd.n4404 gnd.n1084 240.244
R4459 gnd.n4404 gnd.n1099 240.244
R4460 gnd.n4400 gnd.n1099 240.244
R4461 gnd.n4400 gnd.n1105 240.244
R4462 gnd.n4392 gnd.n1105 240.244
R4463 gnd.n4392 gnd.n1121 240.244
R4464 gnd.n4388 gnd.n1121 240.244
R4465 gnd.n4388 gnd.n1127 240.244
R4466 gnd.n4380 gnd.n1127 240.244
R4467 gnd.n4380 gnd.n1143 240.244
R4468 gnd.n4376 gnd.n1143 240.244
R4469 gnd.n4376 gnd.n1149 240.244
R4470 gnd.n4368 gnd.n1149 240.244
R4471 gnd.n6122 gnd.n636 240.244
R4472 gnd.n6122 gnd.n632 240.244
R4473 gnd.n6128 gnd.n632 240.244
R4474 gnd.n6128 gnd.n630 240.244
R4475 gnd.n6132 gnd.n630 240.244
R4476 gnd.n6132 gnd.n626 240.244
R4477 gnd.n6138 gnd.n626 240.244
R4478 gnd.n6138 gnd.n624 240.244
R4479 gnd.n6142 gnd.n624 240.244
R4480 gnd.n6142 gnd.n620 240.244
R4481 gnd.n6148 gnd.n620 240.244
R4482 gnd.n6148 gnd.n618 240.244
R4483 gnd.n6152 gnd.n618 240.244
R4484 gnd.n6152 gnd.n614 240.244
R4485 gnd.n6158 gnd.n614 240.244
R4486 gnd.n6158 gnd.n612 240.244
R4487 gnd.n6162 gnd.n612 240.244
R4488 gnd.n6162 gnd.n608 240.244
R4489 gnd.n6168 gnd.n608 240.244
R4490 gnd.n6168 gnd.n606 240.244
R4491 gnd.n6172 gnd.n606 240.244
R4492 gnd.n6172 gnd.n602 240.244
R4493 gnd.n6178 gnd.n602 240.244
R4494 gnd.n6178 gnd.n600 240.244
R4495 gnd.n6182 gnd.n600 240.244
R4496 gnd.n6182 gnd.n596 240.244
R4497 gnd.n6188 gnd.n596 240.244
R4498 gnd.n6188 gnd.n594 240.244
R4499 gnd.n6192 gnd.n594 240.244
R4500 gnd.n6192 gnd.n590 240.244
R4501 gnd.n6198 gnd.n590 240.244
R4502 gnd.n6198 gnd.n588 240.244
R4503 gnd.n6202 gnd.n588 240.244
R4504 gnd.n6202 gnd.n584 240.244
R4505 gnd.n6208 gnd.n584 240.244
R4506 gnd.n6208 gnd.n582 240.244
R4507 gnd.n6212 gnd.n582 240.244
R4508 gnd.n6212 gnd.n578 240.244
R4509 gnd.n6218 gnd.n578 240.244
R4510 gnd.n6218 gnd.n576 240.244
R4511 gnd.n6222 gnd.n576 240.244
R4512 gnd.n6222 gnd.n572 240.244
R4513 gnd.n6228 gnd.n572 240.244
R4514 gnd.n6228 gnd.n570 240.244
R4515 gnd.n6232 gnd.n570 240.244
R4516 gnd.n6232 gnd.n566 240.244
R4517 gnd.n6238 gnd.n566 240.244
R4518 gnd.n6238 gnd.n564 240.244
R4519 gnd.n6242 gnd.n564 240.244
R4520 gnd.n6242 gnd.n560 240.244
R4521 gnd.n6248 gnd.n560 240.244
R4522 gnd.n6248 gnd.n558 240.244
R4523 gnd.n6252 gnd.n558 240.244
R4524 gnd.n6252 gnd.n554 240.244
R4525 gnd.n6258 gnd.n554 240.244
R4526 gnd.n6258 gnd.n552 240.244
R4527 gnd.n6262 gnd.n552 240.244
R4528 gnd.n6262 gnd.n548 240.244
R4529 gnd.n6268 gnd.n548 240.244
R4530 gnd.n6268 gnd.n546 240.244
R4531 gnd.n6272 gnd.n546 240.244
R4532 gnd.n6272 gnd.n542 240.244
R4533 gnd.n6278 gnd.n542 240.244
R4534 gnd.n6278 gnd.n540 240.244
R4535 gnd.n6282 gnd.n540 240.244
R4536 gnd.n6282 gnd.n536 240.244
R4537 gnd.n6288 gnd.n536 240.244
R4538 gnd.n6288 gnd.n534 240.244
R4539 gnd.n6292 gnd.n534 240.244
R4540 gnd.n6292 gnd.n530 240.244
R4541 gnd.n6298 gnd.n530 240.244
R4542 gnd.n6298 gnd.n528 240.244
R4543 gnd.n6302 gnd.n528 240.244
R4544 gnd.n6302 gnd.n524 240.244
R4545 gnd.n6308 gnd.n524 240.244
R4546 gnd.n6308 gnd.n522 240.244
R4547 gnd.n6312 gnd.n522 240.244
R4548 gnd.n6312 gnd.n518 240.244
R4549 gnd.n6318 gnd.n518 240.244
R4550 gnd.n6318 gnd.n516 240.244
R4551 gnd.n6322 gnd.n516 240.244
R4552 gnd.n6322 gnd.n512 240.244
R4553 gnd.n6328 gnd.n512 240.244
R4554 gnd.n6328 gnd.n510 240.244
R4555 gnd.n6332 gnd.n510 240.244
R4556 gnd.n6332 gnd.n506 240.244
R4557 gnd.n6338 gnd.n506 240.244
R4558 gnd.n6338 gnd.n504 240.244
R4559 gnd.n6342 gnd.n504 240.244
R4560 gnd.n6342 gnd.n500 240.244
R4561 gnd.n6348 gnd.n500 240.244
R4562 gnd.n6348 gnd.n498 240.244
R4563 gnd.n6352 gnd.n498 240.244
R4564 gnd.n6352 gnd.n494 240.244
R4565 gnd.n6358 gnd.n494 240.244
R4566 gnd.n6358 gnd.n492 240.244
R4567 gnd.n6362 gnd.n492 240.244
R4568 gnd.n6362 gnd.n488 240.244
R4569 gnd.n6368 gnd.n488 240.244
R4570 gnd.n6368 gnd.n486 240.244
R4571 gnd.n6372 gnd.n486 240.244
R4572 gnd.n6372 gnd.n482 240.244
R4573 gnd.n6378 gnd.n482 240.244
R4574 gnd.n6378 gnd.n480 240.244
R4575 gnd.n6382 gnd.n480 240.244
R4576 gnd.n6382 gnd.n476 240.244
R4577 gnd.n6388 gnd.n476 240.244
R4578 gnd.n6388 gnd.n474 240.244
R4579 gnd.n6392 gnd.n474 240.244
R4580 gnd.n6392 gnd.n470 240.244
R4581 gnd.n6398 gnd.n470 240.244
R4582 gnd.n6398 gnd.n468 240.244
R4583 gnd.n6402 gnd.n468 240.244
R4584 gnd.n6402 gnd.n464 240.244
R4585 gnd.n6408 gnd.n464 240.244
R4586 gnd.n6408 gnd.n462 240.244
R4587 gnd.n6412 gnd.n462 240.244
R4588 gnd.n6412 gnd.n458 240.244
R4589 gnd.n6418 gnd.n458 240.244
R4590 gnd.n6418 gnd.n456 240.244
R4591 gnd.n6422 gnd.n456 240.244
R4592 gnd.n6422 gnd.n452 240.244
R4593 gnd.n6428 gnd.n452 240.244
R4594 gnd.n6428 gnd.n450 240.244
R4595 gnd.n6432 gnd.n450 240.244
R4596 gnd.n6432 gnd.n446 240.244
R4597 gnd.n6438 gnd.n446 240.244
R4598 gnd.n6438 gnd.n444 240.244
R4599 gnd.n6442 gnd.n444 240.244
R4600 gnd.n6442 gnd.n440 240.244
R4601 gnd.n6448 gnd.n440 240.244
R4602 gnd.n6448 gnd.n438 240.244
R4603 gnd.n6452 gnd.n438 240.244
R4604 gnd.n6452 gnd.n434 240.244
R4605 gnd.n6458 gnd.n434 240.244
R4606 gnd.n6458 gnd.n432 240.244
R4607 gnd.n6462 gnd.n432 240.244
R4608 gnd.n6462 gnd.n428 240.244
R4609 gnd.n6468 gnd.n428 240.244
R4610 gnd.n6468 gnd.n426 240.244
R4611 gnd.n6472 gnd.n426 240.244
R4612 gnd.n6472 gnd.n422 240.244
R4613 gnd.n6478 gnd.n422 240.244
R4614 gnd.n6478 gnd.n420 240.244
R4615 gnd.n6482 gnd.n420 240.244
R4616 gnd.n6482 gnd.n416 240.244
R4617 gnd.n6488 gnd.n416 240.244
R4618 gnd.n6488 gnd.n414 240.244
R4619 gnd.n6492 gnd.n414 240.244
R4620 gnd.n6492 gnd.n410 240.244
R4621 gnd.n6499 gnd.n410 240.244
R4622 gnd.n6499 gnd.n408 240.244
R4623 gnd.n6503 gnd.n408 240.244
R4624 gnd.n6503 gnd.n405 240.244
R4625 gnd.n6509 gnd.n403 240.244
R4626 gnd.n6513 gnd.n403 240.244
R4627 gnd.n6513 gnd.n399 240.244
R4628 gnd.n6519 gnd.n399 240.244
R4629 gnd.n6519 gnd.n397 240.244
R4630 gnd.n6523 gnd.n397 240.244
R4631 gnd.n6523 gnd.n393 240.244
R4632 gnd.n6529 gnd.n393 240.244
R4633 gnd.n6529 gnd.n391 240.244
R4634 gnd.n6533 gnd.n391 240.244
R4635 gnd.n6533 gnd.n387 240.244
R4636 gnd.n6539 gnd.n387 240.244
R4637 gnd.n6539 gnd.n385 240.244
R4638 gnd.n6543 gnd.n385 240.244
R4639 gnd.n6543 gnd.n381 240.244
R4640 gnd.n6549 gnd.n381 240.244
R4641 gnd.n6549 gnd.n379 240.244
R4642 gnd.n6553 gnd.n379 240.244
R4643 gnd.n6553 gnd.n375 240.244
R4644 gnd.n6559 gnd.n375 240.244
R4645 gnd.n6559 gnd.n373 240.244
R4646 gnd.n6563 gnd.n373 240.244
R4647 gnd.n6563 gnd.n369 240.244
R4648 gnd.n6569 gnd.n369 240.244
R4649 gnd.n6569 gnd.n367 240.244
R4650 gnd.n6573 gnd.n367 240.244
R4651 gnd.n6573 gnd.n363 240.244
R4652 gnd.n6579 gnd.n363 240.244
R4653 gnd.n6579 gnd.n361 240.244
R4654 gnd.n6583 gnd.n361 240.244
R4655 gnd.n6583 gnd.n357 240.244
R4656 gnd.n6589 gnd.n357 240.244
R4657 gnd.n6589 gnd.n355 240.244
R4658 gnd.n6593 gnd.n355 240.244
R4659 gnd.n6593 gnd.n351 240.244
R4660 gnd.n6599 gnd.n351 240.244
R4661 gnd.n6599 gnd.n349 240.244
R4662 gnd.n6603 gnd.n349 240.244
R4663 gnd.n6603 gnd.n345 240.244
R4664 gnd.n6609 gnd.n345 240.244
R4665 gnd.n6609 gnd.n343 240.244
R4666 gnd.n6613 gnd.n343 240.244
R4667 gnd.n6613 gnd.n339 240.244
R4668 gnd.n6619 gnd.n339 240.244
R4669 gnd.n6619 gnd.n337 240.244
R4670 gnd.n6623 gnd.n337 240.244
R4671 gnd.n6623 gnd.n333 240.244
R4672 gnd.n6629 gnd.n333 240.244
R4673 gnd.n6629 gnd.n331 240.244
R4674 gnd.n6633 gnd.n331 240.244
R4675 gnd.n6633 gnd.n327 240.244
R4676 gnd.n6639 gnd.n327 240.244
R4677 gnd.n6639 gnd.n325 240.244
R4678 gnd.n6643 gnd.n325 240.244
R4679 gnd.n6643 gnd.n321 240.244
R4680 gnd.n6649 gnd.n321 240.244
R4681 gnd.n6649 gnd.n319 240.244
R4682 gnd.n6653 gnd.n319 240.244
R4683 gnd.n6653 gnd.n315 240.244
R4684 gnd.n6659 gnd.n315 240.244
R4685 gnd.n6659 gnd.n313 240.244
R4686 gnd.n6663 gnd.n313 240.244
R4687 gnd.n6663 gnd.n309 240.244
R4688 gnd.n6669 gnd.n309 240.244
R4689 gnd.n6669 gnd.n307 240.244
R4690 gnd.n6673 gnd.n307 240.244
R4691 gnd.n6673 gnd.n303 240.244
R4692 gnd.n6679 gnd.n303 240.244
R4693 gnd.n6679 gnd.n301 240.244
R4694 gnd.n6683 gnd.n301 240.244
R4695 gnd.n6683 gnd.n297 240.244
R4696 gnd.n6689 gnd.n297 240.244
R4697 gnd.n6689 gnd.n295 240.244
R4698 gnd.n6693 gnd.n295 240.244
R4699 gnd.n6693 gnd.n291 240.244
R4700 gnd.n6699 gnd.n291 240.244
R4701 gnd.n6699 gnd.n289 240.244
R4702 gnd.n6703 gnd.n289 240.244
R4703 gnd.n6703 gnd.n285 240.244
R4704 gnd.n6709 gnd.n285 240.244
R4705 gnd.n6709 gnd.n283 240.244
R4706 gnd.n6714 gnd.n283 240.244
R4707 gnd.n6714 gnd.n279 240.244
R4708 gnd.n6721 gnd.n279 240.244
R4709 gnd.n2316 gnd.n2315 240.244
R4710 gnd.n2317 gnd.n2316 240.244
R4711 gnd.n2317 gnd.n2226 240.244
R4712 gnd.n2324 gnd.n2226 240.244
R4713 gnd.n2324 gnd.n2227 240.244
R4714 gnd.n2304 gnd.n2227 240.244
R4715 gnd.n2304 gnd.n2303 240.244
R4716 gnd.n2303 gnd.n2302 240.244
R4717 gnd.n2302 gnd.n2300 240.244
R4718 gnd.n2300 gnd.n2297 240.244
R4719 gnd.n2297 gnd.n2296 240.244
R4720 gnd.n2296 gnd.n2293 240.244
R4721 gnd.n2293 gnd.n2292 240.244
R4722 gnd.n2292 gnd.n2235 240.244
R4723 gnd.n2288 gnd.n2235 240.244
R4724 gnd.n2288 gnd.n2287 240.244
R4725 gnd.n2287 gnd.n2286 240.244
R4726 gnd.n2286 gnd.n2238 240.244
R4727 gnd.n2282 gnd.n2238 240.244
R4728 gnd.n2282 gnd.n2281 240.244
R4729 gnd.n2281 gnd.n2280 240.244
R4730 gnd.n2280 gnd.n2244 240.244
R4731 gnd.n2276 gnd.n2244 240.244
R4732 gnd.n2276 gnd.n2275 240.244
R4733 gnd.n2275 gnd.n2274 240.244
R4734 gnd.n2274 gnd.n2250 240.244
R4735 gnd.n2270 gnd.n2250 240.244
R4736 gnd.n2270 gnd.n2269 240.244
R4737 gnd.n2269 gnd.n2268 240.244
R4738 gnd.n2268 gnd.n2256 240.244
R4739 gnd.n2264 gnd.n2256 240.244
R4740 gnd.n2264 gnd.n2263 240.244
R4741 gnd.n2263 gnd.n1984 240.244
R4742 gnd.n2901 gnd.n1984 240.244
R4743 gnd.n2901 gnd.n1980 240.244
R4744 gnd.n2907 gnd.n1980 240.244
R4745 gnd.n2907 gnd.n1970 240.244
R4746 gnd.n2917 gnd.n1970 240.244
R4747 gnd.n2917 gnd.n1965 240.244
R4748 gnd.n2925 gnd.n1965 240.244
R4749 gnd.n2925 gnd.n1966 240.244
R4750 gnd.n1966 gnd.n1938 240.244
R4751 gnd.n3041 gnd.n1938 240.244
R4752 gnd.n3041 gnd.n1934 240.244
R4753 gnd.n3047 gnd.n1934 240.244
R4754 gnd.n3047 gnd.n1924 240.244
R4755 gnd.n3057 gnd.n1924 240.244
R4756 gnd.n3057 gnd.n1920 240.244
R4757 gnd.n3063 gnd.n1920 240.244
R4758 gnd.n3063 gnd.n1909 240.244
R4759 gnd.n3073 gnd.n1909 240.244
R4760 gnd.n3073 gnd.n1905 240.244
R4761 gnd.n3079 gnd.n1905 240.244
R4762 gnd.n3079 gnd.n1895 240.244
R4763 gnd.n3088 gnd.n1895 240.244
R4764 gnd.n3088 gnd.n1890 240.244
R4765 gnd.n3096 gnd.n1890 240.244
R4766 gnd.n3096 gnd.n1891 240.244
R4767 gnd.n1891 gnd.n1863 240.244
R4768 gnd.n3214 gnd.n1863 240.244
R4769 gnd.n3214 gnd.n1859 240.244
R4770 gnd.n3220 gnd.n1859 240.244
R4771 gnd.n3220 gnd.n1849 240.244
R4772 gnd.n3230 gnd.n1849 240.244
R4773 gnd.n3230 gnd.n1845 240.244
R4774 gnd.n3236 gnd.n1845 240.244
R4775 gnd.n3236 gnd.n1836 240.244
R4776 gnd.n3246 gnd.n1836 240.244
R4777 gnd.n3246 gnd.n1832 240.244
R4778 gnd.n3252 gnd.n1832 240.244
R4779 gnd.n3252 gnd.n1825 240.244
R4780 gnd.n3262 gnd.n1825 240.244
R4781 gnd.n3262 gnd.n1820 240.244
R4782 gnd.n3270 gnd.n1820 240.244
R4783 gnd.n3270 gnd.n1821 240.244
R4784 gnd.n1821 gnd.n1792 240.244
R4785 gnd.n3385 gnd.n1792 240.244
R4786 gnd.n3385 gnd.n1788 240.244
R4787 gnd.n3391 gnd.n1788 240.244
R4788 gnd.n3391 gnd.n1777 240.244
R4789 gnd.n3401 gnd.n1777 240.244
R4790 gnd.n3401 gnd.n1773 240.244
R4791 gnd.n3407 gnd.n1773 240.244
R4792 gnd.n3407 gnd.n1762 240.244
R4793 gnd.n3417 gnd.n1762 240.244
R4794 gnd.n3417 gnd.n1758 240.244
R4795 gnd.n3423 gnd.n1758 240.244
R4796 gnd.n3423 gnd.n1749 240.244
R4797 gnd.n3433 gnd.n1749 240.244
R4798 gnd.n3433 gnd.n1744 240.244
R4799 gnd.n3441 gnd.n1744 240.244
R4800 gnd.n3441 gnd.n1745 240.244
R4801 gnd.n1745 gnd.n1717 240.244
R4802 gnd.n3791 gnd.n1717 240.244
R4803 gnd.n3791 gnd.n1713 240.244
R4804 gnd.n3797 gnd.n1713 240.244
R4805 gnd.n3797 gnd.n1704 240.244
R4806 gnd.n3807 gnd.n1704 240.244
R4807 gnd.n3807 gnd.n1700 240.244
R4808 gnd.n3813 gnd.n1700 240.244
R4809 gnd.n3813 gnd.n1690 240.244
R4810 gnd.n3823 gnd.n1690 240.244
R4811 gnd.n3823 gnd.n1686 240.244
R4812 gnd.n3829 gnd.n1686 240.244
R4813 gnd.n3829 gnd.n1677 240.244
R4814 gnd.n3839 gnd.n1677 240.244
R4815 gnd.n3839 gnd.n1673 240.244
R4816 gnd.n3845 gnd.n1673 240.244
R4817 gnd.n3845 gnd.n1663 240.244
R4818 gnd.n3855 gnd.n1663 240.244
R4819 gnd.n3855 gnd.n1659 240.244
R4820 gnd.n3861 gnd.n1659 240.244
R4821 gnd.n3861 gnd.n1649 240.244
R4822 gnd.n3873 gnd.n1649 240.244
R4823 gnd.n3873 gnd.n1644 240.244
R4824 gnd.n3882 gnd.n1644 240.244
R4825 gnd.n3882 gnd.n1645 240.244
R4826 gnd.n1645 gnd.n1273 240.244
R4827 gnd.n4236 gnd.n1273 240.244
R4828 gnd.n4236 gnd.n1276 240.244
R4829 gnd.n4232 gnd.n1276 240.244
R4830 gnd.n4232 gnd.n1282 240.244
R4831 gnd.n3963 gnd.n1282 240.244
R4832 gnd.n3964 gnd.n3963 240.244
R4833 gnd.n3964 gnd.n3957 240.244
R4834 gnd.n3972 gnd.n3957 240.244
R4835 gnd.n3972 gnd.n3958 240.244
R4836 gnd.n3958 gnd.n1486 240.244
R4837 gnd.n3996 gnd.n1486 240.244
R4838 gnd.n3996 gnd.n1481 240.244
R4839 gnd.n4004 gnd.n1481 240.244
R4840 gnd.n4004 gnd.n1482 240.244
R4841 gnd.n1482 gnd.n1461 240.244
R4842 gnd.n4027 gnd.n1461 240.244
R4843 gnd.n4027 gnd.n1456 240.244
R4844 gnd.n4038 gnd.n1456 240.244
R4845 gnd.n4038 gnd.n1457 240.244
R4846 gnd.n1457 gnd.n1436 240.244
R4847 gnd.n4061 gnd.n1436 240.244
R4848 gnd.n4062 gnd.n4061 240.244
R4849 gnd.n4062 gnd.n1432 240.244
R4850 gnd.n4069 gnd.n1432 240.244
R4851 gnd.n4069 gnd.n1433 240.244
R4852 gnd.n1433 gnd.n1401 240.244
R4853 gnd.n4101 gnd.n1401 240.244
R4854 gnd.n4101 gnd.n1398 240.244
R4855 gnd.n4113 gnd.n1398 240.244
R4856 gnd.n4113 gnd.n1399 240.244
R4857 gnd.n4108 gnd.n1399 240.244
R4858 gnd.n4108 gnd.n4107 240.244
R4859 gnd.n4107 gnd.n272 240.244
R4860 gnd.n6726 gnd.n272 240.244
R4861 gnd.n6726 gnd.n273 240.244
R4862 gnd.n6722 gnd.n273 240.244
R4863 gnd.n6118 gnd.n638 240.244
R4864 gnd.n6114 gnd.n638 240.244
R4865 gnd.n6114 gnd.n643 240.244
R4866 gnd.n6110 gnd.n643 240.244
R4867 gnd.n6110 gnd.n645 240.244
R4868 gnd.n6106 gnd.n645 240.244
R4869 gnd.n6106 gnd.n651 240.244
R4870 gnd.n6102 gnd.n651 240.244
R4871 gnd.n6102 gnd.n653 240.244
R4872 gnd.n6098 gnd.n653 240.244
R4873 gnd.n6098 gnd.n659 240.244
R4874 gnd.n6094 gnd.n659 240.244
R4875 gnd.n6094 gnd.n661 240.244
R4876 gnd.n6090 gnd.n661 240.244
R4877 gnd.n6090 gnd.n667 240.244
R4878 gnd.n6086 gnd.n667 240.244
R4879 gnd.n6086 gnd.n669 240.244
R4880 gnd.n6082 gnd.n669 240.244
R4881 gnd.n6082 gnd.n675 240.244
R4882 gnd.n6078 gnd.n675 240.244
R4883 gnd.n6078 gnd.n677 240.244
R4884 gnd.n6074 gnd.n677 240.244
R4885 gnd.n6074 gnd.n683 240.244
R4886 gnd.n6070 gnd.n683 240.244
R4887 gnd.n6070 gnd.n685 240.244
R4888 gnd.n6066 gnd.n685 240.244
R4889 gnd.n6066 gnd.n691 240.244
R4890 gnd.n6062 gnd.n691 240.244
R4891 gnd.n6062 gnd.n693 240.244
R4892 gnd.n6058 gnd.n693 240.244
R4893 gnd.n6058 gnd.n699 240.244
R4894 gnd.n6054 gnd.n699 240.244
R4895 gnd.n6054 gnd.n701 240.244
R4896 gnd.n6050 gnd.n701 240.244
R4897 gnd.n6050 gnd.n707 240.244
R4898 gnd.n6046 gnd.n707 240.244
R4899 gnd.n6046 gnd.n709 240.244
R4900 gnd.n6042 gnd.n709 240.244
R4901 gnd.n6042 gnd.n715 240.244
R4902 gnd.n6038 gnd.n715 240.244
R4903 gnd.n6038 gnd.n717 240.244
R4904 gnd.n6034 gnd.n717 240.244
R4905 gnd.n6034 gnd.n723 240.244
R4906 gnd.n6030 gnd.n723 240.244
R4907 gnd.n6030 gnd.n725 240.244
R4908 gnd.n6026 gnd.n725 240.244
R4909 gnd.n6026 gnd.n731 240.244
R4910 gnd.n6022 gnd.n731 240.244
R4911 gnd.n6022 gnd.n733 240.244
R4912 gnd.n6018 gnd.n733 240.244
R4913 gnd.n6018 gnd.n739 240.244
R4914 gnd.n6014 gnd.n739 240.244
R4915 gnd.n6014 gnd.n741 240.244
R4916 gnd.n6010 gnd.n741 240.244
R4917 gnd.n6010 gnd.n747 240.244
R4918 gnd.n6006 gnd.n747 240.244
R4919 gnd.n6006 gnd.n749 240.244
R4920 gnd.n6002 gnd.n749 240.244
R4921 gnd.n6002 gnd.n755 240.244
R4922 gnd.n5998 gnd.n755 240.244
R4923 gnd.n5998 gnd.n757 240.244
R4924 gnd.n5994 gnd.n757 240.244
R4925 gnd.n5994 gnd.n763 240.244
R4926 gnd.n5990 gnd.n763 240.244
R4927 gnd.n5990 gnd.n765 240.244
R4928 gnd.n5986 gnd.n765 240.244
R4929 gnd.n5986 gnd.n771 240.244
R4930 gnd.n5982 gnd.n771 240.244
R4931 gnd.n5982 gnd.n773 240.244
R4932 gnd.n5978 gnd.n773 240.244
R4933 gnd.n5978 gnd.n779 240.244
R4934 gnd.n5974 gnd.n779 240.244
R4935 gnd.n5974 gnd.n781 240.244
R4936 gnd.n5970 gnd.n781 240.244
R4937 gnd.n5970 gnd.n787 240.244
R4938 gnd.n5966 gnd.n787 240.244
R4939 gnd.n5966 gnd.n789 240.244
R4940 gnd.n5962 gnd.n789 240.244
R4941 gnd.n5962 gnd.n795 240.244
R4942 gnd.n5958 gnd.n795 240.244
R4943 gnd.n5958 gnd.n797 240.244
R4944 gnd.n5954 gnd.n797 240.244
R4945 gnd.n5954 gnd.n803 240.244
R4946 gnd.n2309 gnd.n803 240.244
R4947 gnd.n1169 gnd.n1168 240.244
R4948 gnd.n1170 gnd.n1169 240.244
R4949 gnd.n1971 gnd.n1170 240.244
R4950 gnd.n1971 gnd.n1173 240.244
R4951 gnd.n1174 gnd.n1173 240.244
R4952 gnd.n1175 gnd.n1174 240.244
R4953 gnd.n1940 gnd.n1175 240.244
R4954 gnd.n1940 gnd.n1178 240.244
R4955 gnd.n1179 gnd.n1178 240.244
R4956 gnd.n1180 gnd.n1179 240.244
R4957 gnd.n1925 gnd.n1180 240.244
R4958 gnd.n1925 gnd.n1183 240.244
R4959 gnd.n1184 gnd.n1183 240.244
R4960 gnd.n1185 gnd.n1184 240.244
R4961 gnd.n1911 gnd.n1185 240.244
R4962 gnd.n1911 gnd.n1188 240.244
R4963 gnd.n1189 gnd.n1188 240.244
R4964 gnd.n1190 gnd.n1189 240.244
R4965 gnd.n1897 gnd.n1190 240.244
R4966 gnd.n1897 gnd.n1193 240.244
R4967 gnd.n1194 gnd.n1193 240.244
R4968 gnd.n1195 gnd.n1194 240.244
R4969 gnd.n1881 gnd.n1195 240.244
R4970 gnd.n1881 gnd.n1198 240.244
R4971 gnd.n1199 gnd.n1198 240.244
R4972 gnd.n1200 gnd.n1199 240.244
R4973 gnd.n1874 gnd.n1200 240.244
R4974 gnd.n1874 gnd.n1203 240.244
R4975 gnd.n1204 gnd.n1203 240.244
R4976 gnd.n1205 gnd.n1204 240.244
R4977 gnd.n3126 gnd.n1205 240.244
R4978 gnd.n3126 gnd.n1208 240.244
R4979 gnd.n1209 gnd.n1208 240.244
R4980 gnd.n1210 gnd.n1209 240.244
R4981 gnd.n3142 gnd.n1210 240.244
R4982 gnd.n3142 gnd.n1213 240.244
R4983 gnd.n1214 gnd.n1213 240.244
R4984 gnd.n1215 gnd.n1214 240.244
R4985 gnd.n1809 gnd.n1215 240.244
R4986 gnd.n1809 gnd.n1218 240.244
R4987 gnd.n1219 gnd.n1218 240.244
R4988 gnd.n1220 gnd.n1219 240.244
R4989 gnd.n1786 gnd.n1220 240.244
R4990 gnd.n1786 gnd.n1223 240.244
R4991 gnd.n1224 gnd.n1223 240.244
R4992 gnd.n1225 gnd.n1224 240.244
R4993 gnd.n1771 gnd.n1225 240.244
R4994 gnd.n1771 gnd.n1228 240.244
R4995 gnd.n1229 gnd.n1228 240.244
R4996 gnd.n1230 gnd.n1229 240.244
R4997 gnd.n1756 gnd.n1230 240.244
R4998 gnd.n1756 gnd.n1233 240.244
R4999 gnd.n1234 gnd.n1233 240.244
R5000 gnd.n1235 gnd.n1234 240.244
R5001 gnd.n1742 gnd.n1235 240.244
R5002 gnd.n1742 gnd.n1238 240.244
R5003 gnd.n1239 gnd.n1238 240.244
R5004 gnd.n1240 gnd.n1239 240.244
R5005 gnd.n3458 gnd.n1240 240.244
R5006 gnd.n3458 gnd.n1243 240.244
R5007 gnd.n1244 gnd.n1243 240.244
R5008 gnd.n1245 gnd.n1244 240.244
R5009 gnd.n3774 gnd.n1245 240.244
R5010 gnd.n3774 gnd.n1248 240.244
R5011 gnd.n1249 gnd.n1248 240.244
R5012 gnd.n1250 gnd.n1249 240.244
R5013 gnd.n3481 gnd.n1250 240.244
R5014 gnd.n3481 gnd.n1253 240.244
R5015 gnd.n1254 gnd.n1253 240.244
R5016 gnd.n1255 gnd.n1254 240.244
R5017 gnd.n3743 gnd.n1255 240.244
R5018 gnd.n3743 gnd.n1258 240.244
R5019 gnd.n1259 gnd.n1258 240.244
R5020 gnd.n1260 gnd.n1259 240.244
R5021 gnd.n3508 gnd.n1260 240.244
R5022 gnd.n3508 gnd.n1263 240.244
R5023 gnd.n1264 gnd.n1263 240.244
R5024 gnd.n1265 gnd.n1264 240.244
R5025 gnd.n3542 gnd.n1265 240.244
R5026 gnd.n3542 gnd.n1268 240.244
R5027 gnd.n1269 gnd.n1268 240.244
R5028 gnd.n4239 gnd.n1269 240.244
R5029 gnd.n2060 gnd.n2059 240.244
R5030 gnd.n2072 gnd.n2071 240.244
R5031 gnd.n2044 gnd.n2043 240.244
R5032 gnd.n2084 gnd.n2083 240.244
R5033 gnd.n2096 gnd.n2095 240.244
R5034 gnd.n2032 gnd.n2031 240.244
R5035 gnd.n2110 gnd.n2109 240.244
R5036 gnd.n2012 gnd.n2011 240.244
R5037 gnd.n2871 gnd.n2870 240.244
R5038 gnd.n2879 gnd.n2878 240.244
R5039 gnd.n2882 gnd.n2881 240.244
R5040 gnd.n2889 gnd.n2888 240.244
R5041 gnd.n2892 gnd.n1999 240.244
R5042 gnd.n2898 gnd.n1977 240.244
R5043 gnd.n2909 gnd.n1974 240.244
R5044 gnd.n2915 gnd.n1974 240.244
R5045 gnd.n2915 gnd.n1962 240.244
R5046 gnd.n2927 gnd.n1962 240.244
R5047 gnd.n2927 gnd.n1957 240.244
R5048 gnd.n2934 gnd.n1957 240.244
R5049 gnd.n2934 gnd.n1943 240.244
R5050 gnd.n1943 gnd.n1931 240.244
R5051 gnd.n3049 gnd.n1931 240.244
R5052 gnd.n3049 gnd.n1927 240.244
R5053 gnd.n3055 gnd.n1927 240.244
R5054 gnd.n3055 gnd.n1917 240.244
R5055 gnd.n3065 gnd.n1917 240.244
R5056 gnd.n3065 gnd.n1913 240.244
R5057 gnd.n3071 gnd.n1913 240.244
R5058 gnd.n3071 gnd.n1903 240.244
R5059 gnd.n3081 gnd.n1903 240.244
R5060 gnd.n3081 gnd.n1899 240.244
R5061 gnd.n3087 gnd.n1899 240.244
R5062 gnd.n3087 gnd.n1887 240.244
R5063 gnd.n3098 gnd.n1887 240.244
R5064 gnd.n3098 gnd.n1882 240.244
R5065 gnd.n3105 gnd.n1882 240.244
R5066 gnd.n3105 gnd.n1867 240.244
R5067 gnd.n1867 gnd.n1856 240.244
R5068 gnd.n3222 gnd.n1856 240.244
R5069 gnd.n3222 gnd.n1852 240.244
R5070 gnd.n3228 gnd.n1852 240.244
R5071 gnd.n3228 gnd.n1843 240.244
R5072 gnd.n3238 gnd.n1843 240.244
R5073 gnd.n3238 gnd.n1839 240.244
R5074 gnd.n3244 gnd.n1839 240.244
R5075 gnd.n3244 gnd.n1831 240.244
R5076 gnd.n3254 gnd.n1831 240.244
R5077 gnd.n3254 gnd.n1827 240.244
R5078 gnd.n3260 gnd.n1827 240.244
R5079 gnd.n3260 gnd.n1817 240.244
R5080 gnd.n3272 gnd.n1817 240.244
R5081 gnd.n3272 gnd.n1812 240.244
R5082 gnd.n3279 gnd.n1812 240.244
R5083 gnd.n3279 gnd.n1797 240.244
R5084 gnd.n1797 gnd.n1784 240.244
R5085 gnd.n3393 gnd.n1784 240.244
R5086 gnd.n3393 gnd.n1780 240.244
R5087 gnd.n3399 gnd.n1780 240.244
R5088 gnd.n3399 gnd.n1769 240.244
R5089 gnd.n3409 gnd.n1769 240.244
R5090 gnd.n3409 gnd.n1765 240.244
R5091 gnd.n3415 gnd.n1765 240.244
R5092 gnd.n3415 gnd.n1755 240.244
R5093 gnd.n3425 gnd.n1755 240.244
R5094 gnd.n3425 gnd.n1751 240.244
R5095 gnd.n3431 gnd.n1751 240.244
R5096 gnd.n3431 gnd.n1740 240.244
R5097 gnd.n3443 gnd.n1740 240.244
R5098 gnd.n3443 gnd.n1735 240.244
R5099 gnd.n3450 gnd.n1735 240.244
R5100 gnd.n3450 gnd.n1720 240.244
R5101 gnd.n1720 gnd.n1710 240.244
R5102 gnd.n3799 gnd.n1710 240.244
R5103 gnd.n3799 gnd.n1706 240.244
R5104 gnd.n3805 gnd.n1706 240.244
R5105 gnd.n3805 gnd.n1697 240.244
R5106 gnd.n3815 gnd.n1697 240.244
R5107 gnd.n3815 gnd.n1693 240.244
R5108 gnd.n3821 gnd.n1693 240.244
R5109 gnd.n3821 gnd.n1684 240.244
R5110 gnd.n3831 gnd.n1684 240.244
R5111 gnd.n3831 gnd.n1680 240.244
R5112 gnd.n3837 gnd.n1680 240.244
R5113 gnd.n3837 gnd.n1670 240.244
R5114 gnd.n3847 gnd.n1670 240.244
R5115 gnd.n3847 gnd.n1666 240.244
R5116 gnd.n3853 gnd.n1666 240.244
R5117 gnd.n3853 gnd.n1656 240.244
R5118 gnd.n3863 gnd.n1656 240.244
R5119 gnd.n3863 gnd.n1651 240.244
R5120 gnd.n3871 gnd.n1651 240.244
R5121 gnd.n3871 gnd.n1643 240.244
R5122 gnd.n3884 gnd.n1643 240.244
R5123 gnd.n3885 gnd.n3884 240.244
R5124 gnd.n3885 gnd.n1274 240.244
R5125 gnd.n1561 gnd.n1559 240.244
R5126 gnd.n1574 gnd.n1538 240.244
R5127 gnd.n1578 gnd.n1576 240.244
R5128 gnd.n1591 gnd.n1529 240.244
R5129 gnd.n1595 gnd.n1593 240.244
R5130 gnd.n1608 gnd.n1520 240.244
R5131 gnd.n1612 gnd.n1610 240.244
R5132 gnd.n1623 gnd.n1508 240.244
R5133 gnd.n1626 gnd.n1625 240.244
R5134 gnd.n1629 gnd.n1628 240.244
R5135 gnd.n1634 gnd.n1631 240.244
R5136 gnd.n1637 gnd.n1636 240.244
R5137 gnd.n3890 gnd.n1639 240.244
R5138 gnd.n3893 gnd.n3892 240.244
R5139 gnd.n2655 gnd.n2654 240.132
R5140 gnd.n3531 gnd.n3530 240.132
R5141 gnd.n6121 gnd.n6120 225.874
R5142 gnd.n6121 gnd.n631 225.874
R5143 gnd.n6129 gnd.n631 225.874
R5144 gnd.n6130 gnd.n6129 225.874
R5145 gnd.n6131 gnd.n6130 225.874
R5146 gnd.n6131 gnd.n625 225.874
R5147 gnd.n6139 gnd.n625 225.874
R5148 gnd.n6140 gnd.n6139 225.874
R5149 gnd.n6141 gnd.n6140 225.874
R5150 gnd.n6141 gnd.n619 225.874
R5151 gnd.n6149 gnd.n619 225.874
R5152 gnd.n6150 gnd.n6149 225.874
R5153 gnd.n6151 gnd.n6150 225.874
R5154 gnd.n6151 gnd.n613 225.874
R5155 gnd.n6159 gnd.n613 225.874
R5156 gnd.n6160 gnd.n6159 225.874
R5157 gnd.n6161 gnd.n6160 225.874
R5158 gnd.n6161 gnd.n607 225.874
R5159 gnd.n6169 gnd.n607 225.874
R5160 gnd.n6170 gnd.n6169 225.874
R5161 gnd.n6171 gnd.n6170 225.874
R5162 gnd.n6171 gnd.n601 225.874
R5163 gnd.n6179 gnd.n601 225.874
R5164 gnd.n6180 gnd.n6179 225.874
R5165 gnd.n6181 gnd.n6180 225.874
R5166 gnd.n6181 gnd.n595 225.874
R5167 gnd.n6189 gnd.n595 225.874
R5168 gnd.n6190 gnd.n6189 225.874
R5169 gnd.n6191 gnd.n6190 225.874
R5170 gnd.n6191 gnd.n589 225.874
R5171 gnd.n6199 gnd.n589 225.874
R5172 gnd.n6200 gnd.n6199 225.874
R5173 gnd.n6201 gnd.n6200 225.874
R5174 gnd.n6201 gnd.n583 225.874
R5175 gnd.n6209 gnd.n583 225.874
R5176 gnd.n6210 gnd.n6209 225.874
R5177 gnd.n6211 gnd.n6210 225.874
R5178 gnd.n6211 gnd.n577 225.874
R5179 gnd.n6219 gnd.n577 225.874
R5180 gnd.n6220 gnd.n6219 225.874
R5181 gnd.n6221 gnd.n6220 225.874
R5182 gnd.n6221 gnd.n571 225.874
R5183 gnd.n6229 gnd.n571 225.874
R5184 gnd.n6230 gnd.n6229 225.874
R5185 gnd.n6231 gnd.n6230 225.874
R5186 gnd.n6231 gnd.n565 225.874
R5187 gnd.n6239 gnd.n565 225.874
R5188 gnd.n6240 gnd.n6239 225.874
R5189 gnd.n6241 gnd.n6240 225.874
R5190 gnd.n6241 gnd.n559 225.874
R5191 gnd.n6249 gnd.n559 225.874
R5192 gnd.n6250 gnd.n6249 225.874
R5193 gnd.n6251 gnd.n6250 225.874
R5194 gnd.n6251 gnd.n553 225.874
R5195 gnd.n6259 gnd.n553 225.874
R5196 gnd.n6260 gnd.n6259 225.874
R5197 gnd.n6261 gnd.n6260 225.874
R5198 gnd.n6261 gnd.n547 225.874
R5199 gnd.n6269 gnd.n547 225.874
R5200 gnd.n6270 gnd.n6269 225.874
R5201 gnd.n6271 gnd.n6270 225.874
R5202 gnd.n6271 gnd.n541 225.874
R5203 gnd.n6279 gnd.n541 225.874
R5204 gnd.n6280 gnd.n6279 225.874
R5205 gnd.n6281 gnd.n6280 225.874
R5206 gnd.n6281 gnd.n535 225.874
R5207 gnd.n6289 gnd.n535 225.874
R5208 gnd.n6290 gnd.n6289 225.874
R5209 gnd.n6291 gnd.n6290 225.874
R5210 gnd.n6291 gnd.n529 225.874
R5211 gnd.n6299 gnd.n529 225.874
R5212 gnd.n6300 gnd.n6299 225.874
R5213 gnd.n6301 gnd.n6300 225.874
R5214 gnd.n6301 gnd.n523 225.874
R5215 gnd.n6309 gnd.n523 225.874
R5216 gnd.n6310 gnd.n6309 225.874
R5217 gnd.n6311 gnd.n6310 225.874
R5218 gnd.n6311 gnd.n517 225.874
R5219 gnd.n6319 gnd.n517 225.874
R5220 gnd.n6320 gnd.n6319 225.874
R5221 gnd.n6321 gnd.n6320 225.874
R5222 gnd.n6321 gnd.n511 225.874
R5223 gnd.n6329 gnd.n511 225.874
R5224 gnd.n6330 gnd.n6329 225.874
R5225 gnd.n6331 gnd.n6330 225.874
R5226 gnd.n6331 gnd.n505 225.874
R5227 gnd.n6339 gnd.n505 225.874
R5228 gnd.n6340 gnd.n6339 225.874
R5229 gnd.n6341 gnd.n6340 225.874
R5230 gnd.n6341 gnd.n499 225.874
R5231 gnd.n6349 gnd.n499 225.874
R5232 gnd.n6350 gnd.n6349 225.874
R5233 gnd.n6351 gnd.n6350 225.874
R5234 gnd.n6351 gnd.n493 225.874
R5235 gnd.n6359 gnd.n493 225.874
R5236 gnd.n6360 gnd.n6359 225.874
R5237 gnd.n6361 gnd.n6360 225.874
R5238 gnd.n6361 gnd.n487 225.874
R5239 gnd.n6369 gnd.n487 225.874
R5240 gnd.n6370 gnd.n6369 225.874
R5241 gnd.n6371 gnd.n6370 225.874
R5242 gnd.n6371 gnd.n481 225.874
R5243 gnd.n6379 gnd.n481 225.874
R5244 gnd.n6380 gnd.n6379 225.874
R5245 gnd.n6381 gnd.n6380 225.874
R5246 gnd.n6381 gnd.n475 225.874
R5247 gnd.n6389 gnd.n475 225.874
R5248 gnd.n6390 gnd.n6389 225.874
R5249 gnd.n6391 gnd.n6390 225.874
R5250 gnd.n6391 gnd.n469 225.874
R5251 gnd.n6399 gnd.n469 225.874
R5252 gnd.n6400 gnd.n6399 225.874
R5253 gnd.n6401 gnd.n6400 225.874
R5254 gnd.n6401 gnd.n463 225.874
R5255 gnd.n6409 gnd.n463 225.874
R5256 gnd.n6410 gnd.n6409 225.874
R5257 gnd.n6411 gnd.n6410 225.874
R5258 gnd.n6411 gnd.n457 225.874
R5259 gnd.n6419 gnd.n457 225.874
R5260 gnd.n6420 gnd.n6419 225.874
R5261 gnd.n6421 gnd.n6420 225.874
R5262 gnd.n6421 gnd.n451 225.874
R5263 gnd.n6429 gnd.n451 225.874
R5264 gnd.n6430 gnd.n6429 225.874
R5265 gnd.n6431 gnd.n6430 225.874
R5266 gnd.n6431 gnd.n445 225.874
R5267 gnd.n6439 gnd.n445 225.874
R5268 gnd.n6440 gnd.n6439 225.874
R5269 gnd.n6441 gnd.n6440 225.874
R5270 gnd.n6441 gnd.n439 225.874
R5271 gnd.n6449 gnd.n439 225.874
R5272 gnd.n6450 gnd.n6449 225.874
R5273 gnd.n6451 gnd.n6450 225.874
R5274 gnd.n6451 gnd.n433 225.874
R5275 gnd.n6459 gnd.n433 225.874
R5276 gnd.n6460 gnd.n6459 225.874
R5277 gnd.n6461 gnd.n6460 225.874
R5278 gnd.n6461 gnd.n427 225.874
R5279 gnd.n6469 gnd.n427 225.874
R5280 gnd.n6470 gnd.n6469 225.874
R5281 gnd.n6471 gnd.n6470 225.874
R5282 gnd.n6471 gnd.n421 225.874
R5283 gnd.n6479 gnd.n421 225.874
R5284 gnd.n6480 gnd.n6479 225.874
R5285 gnd.n6481 gnd.n6480 225.874
R5286 gnd.n6481 gnd.n415 225.874
R5287 gnd.n6489 gnd.n415 225.874
R5288 gnd.n6490 gnd.n6489 225.874
R5289 gnd.n6491 gnd.n6490 225.874
R5290 gnd.n6491 gnd.n409 225.874
R5291 gnd.n6500 gnd.n409 225.874
R5292 gnd.n6501 gnd.n6500 225.874
R5293 gnd.n6502 gnd.n6501 225.874
R5294 gnd.n6502 gnd.n404 225.874
R5295 gnd.n4981 gnd.t221 224.174
R5296 gnd.n4623 gnd.t154 224.174
R5297 gnd.n1332 gnd.n1289 199.319
R5298 gnd.n1332 gnd.n1290 199.319
R5299 gnd.n2160 gnd.n2130 199.319
R5300 gnd.n2160 gnd.n2129 199.319
R5301 gnd.n2656 gnd.n2653 186.49
R5302 gnd.n3532 gnd.n3529 186.49
R5303 gnd.n5800 gnd.n5799 185
R5304 gnd.n5798 gnd.n5797 185
R5305 gnd.n5777 gnd.n5776 185
R5306 gnd.n5792 gnd.n5791 185
R5307 gnd.n5790 gnd.n5789 185
R5308 gnd.n5781 gnd.n5780 185
R5309 gnd.n5784 gnd.n5783 185
R5310 gnd.n5768 gnd.n5767 185
R5311 gnd.n5766 gnd.n5765 185
R5312 gnd.n5745 gnd.n5744 185
R5313 gnd.n5760 gnd.n5759 185
R5314 gnd.n5758 gnd.n5757 185
R5315 gnd.n5749 gnd.n5748 185
R5316 gnd.n5752 gnd.n5751 185
R5317 gnd.n5736 gnd.n5735 185
R5318 gnd.n5734 gnd.n5733 185
R5319 gnd.n5713 gnd.n5712 185
R5320 gnd.n5728 gnd.n5727 185
R5321 gnd.n5726 gnd.n5725 185
R5322 gnd.n5717 gnd.n5716 185
R5323 gnd.n5720 gnd.n5719 185
R5324 gnd.n5705 gnd.n5704 185
R5325 gnd.n5703 gnd.n5702 185
R5326 gnd.n5682 gnd.n5681 185
R5327 gnd.n5697 gnd.n5696 185
R5328 gnd.n5695 gnd.n5694 185
R5329 gnd.n5686 gnd.n5685 185
R5330 gnd.n5689 gnd.n5688 185
R5331 gnd.n5673 gnd.n5672 185
R5332 gnd.n5671 gnd.n5670 185
R5333 gnd.n5650 gnd.n5649 185
R5334 gnd.n5665 gnd.n5664 185
R5335 gnd.n5663 gnd.n5662 185
R5336 gnd.n5654 gnd.n5653 185
R5337 gnd.n5657 gnd.n5656 185
R5338 gnd.n5641 gnd.n5640 185
R5339 gnd.n5639 gnd.n5638 185
R5340 gnd.n5618 gnd.n5617 185
R5341 gnd.n5633 gnd.n5632 185
R5342 gnd.n5631 gnd.n5630 185
R5343 gnd.n5622 gnd.n5621 185
R5344 gnd.n5625 gnd.n5624 185
R5345 gnd.n5609 gnd.n5608 185
R5346 gnd.n5607 gnd.n5606 185
R5347 gnd.n5586 gnd.n5585 185
R5348 gnd.n5601 gnd.n5600 185
R5349 gnd.n5599 gnd.n5598 185
R5350 gnd.n5590 gnd.n5589 185
R5351 gnd.n5593 gnd.n5592 185
R5352 gnd.n5578 gnd.n5577 185
R5353 gnd.n5576 gnd.n5575 185
R5354 gnd.n5555 gnd.n5554 185
R5355 gnd.n5570 gnd.n5569 185
R5356 gnd.n5568 gnd.n5567 185
R5357 gnd.n5559 gnd.n5558 185
R5358 gnd.n5562 gnd.n5561 185
R5359 gnd.n4982 gnd.t220 178.987
R5360 gnd.n4624 gnd.t155 178.987
R5361 gnd.n1 gnd.t245 170.774
R5362 gnd.n7 gnd.t65 170.103
R5363 gnd.n6 gnd.t243 170.103
R5364 gnd.n5 gnd.t67 170.103
R5365 gnd.n4 gnd.t239 170.103
R5366 gnd.n3 gnd.t50 170.103
R5367 gnd.n2 gnd.t3 170.103
R5368 gnd.n1 gnd.t253 170.103
R5369 gnd.n3564 gnd.n3563 163.367
R5370 gnd.n3568 gnd.n3567 163.367
R5371 gnd.n3572 gnd.n3571 163.367
R5372 gnd.n3576 gnd.n3575 163.367
R5373 gnd.n3580 gnd.n3579 163.367
R5374 gnd.n3584 gnd.n3583 163.367
R5375 gnd.n3588 gnd.n3587 163.367
R5376 gnd.n3592 gnd.n3591 163.367
R5377 gnd.n3596 gnd.n3595 163.367
R5378 gnd.n3600 gnd.n3599 163.367
R5379 gnd.n3604 gnd.n3603 163.367
R5380 gnd.n3608 gnd.n3607 163.367
R5381 gnd.n3612 gnd.n3611 163.367
R5382 gnd.n3616 gnd.n3615 163.367
R5383 gnd.n3621 gnd.n3620 163.367
R5384 gnd.n3625 gnd.n3624 163.367
R5385 gnd.n3713 gnd.n3712 163.367
R5386 gnd.n3709 gnd.n3708 163.367
R5387 gnd.n3704 gnd.n3703 163.367
R5388 gnd.n3700 gnd.n3699 163.367
R5389 gnd.n3696 gnd.n3695 163.367
R5390 gnd.n3692 gnd.n3691 163.367
R5391 gnd.n3688 gnd.n3687 163.367
R5392 gnd.n3684 gnd.n3683 163.367
R5393 gnd.n3680 gnd.n3679 163.367
R5394 gnd.n3676 gnd.n3675 163.367
R5395 gnd.n3672 gnd.n3671 163.367
R5396 gnd.n3668 gnd.n3667 163.367
R5397 gnd.n3664 gnd.n3663 163.367
R5398 gnd.n3660 gnd.n3659 163.367
R5399 gnd.n3656 gnd.n3655 163.367
R5400 gnd.n3652 gnd.n3651 163.367
R5401 gnd.n2764 gnd.n2763 163.367
R5402 gnd.n2763 gnd.n2758 163.367
R5403 gnd.n2759 gnd.n2758 163.367
R5404 gnd.n2759 gnd.n1944 163.367
R5405 gnd.n3039 gnd.n1944 163.367
R5406 gnd.n3039 gnd.n1945 163.367
R5407 gnd.n3035 gnd.n1945 163.367
R5408 gnd.n3035 gnd.n3034 163.367
R5409 gnd.n3034 gnd.n3033 163.367
R5410 gnd.n3033 gnd.n1948 163.367
R5411 gnd.n2947 gnd.n1948 163.367
R5412 gnd.n3023 gnd.n2947 163.367
R5413 gnd.n3023 gnd.n2948 163.367
R5414 gnd.n3019 gnd.n2948 163.367
R5415 gnd.n3019 gnd.n3018 163.367
R5416 gnd.n3018 gnd.n2952 163.367
R5417 gnd.n2963 gnd.n2952 163.367
R5418 gnd.n2963 gnd.n2960 163.367
R5419 gnd.n3007 gnd.n2960 163.367
R5420 gnd.n3007 gnd.n2961 163.367
R5421 gnd.n3003 gnd.n2961 163.367
R5422 gnd.n3003 gnd.n2967 163.367
R5423 gnd.n2975 gnd.n2967 163.367
R5424 gnd.n2993 gnd.n2975 163.367
R5425 gnd.n2993 gnd.n2976 163.367
R5426 gnd.n2989 gnd.n2976 163.367
R5427 gnd.n2989 gnd.n2988 163.367
R5428 gnd.n2988 gnd.n2980 163.367
R5429 gnd.n2980 gnd.n1868 163.367
R5430 gnd.n3212 gnd.n1868 163.367
R5431 gnd.n3212 gnd.n1869 163.367
R5432 gnd.n3208 gnd.n1869 163.367
R5433 gnd.n3208 gnd.n3207 163.367
R5434 gnd.n3207 gnd.n3206 163.367
R5435 gnd.n3206 gnd.n1872 163.367
R5436 gnd.n3121 gnd.n1872 163.367
R5437 gnd.n3121 gnd.n3118 163.367
R5438 gnd.n3195 gnd.n3118 163.367
R5439 gnd.n3195 gnd.n3119 163.367
R5440 gnd.n3191 gnd.n3119 163.367
R5441 gnd.n3191 gnd.n3125 163.367
R5442 gnd.n3136 gnd.n3125 163.367
R5443 gnd.n3136 gnd.n3134 163.367
R5444 gnd.n3180 gnd.n3134 163.367
R5445 gnd.n3180 gnd.n3135 163.367
R5446 gnd.n3176 gnd.n3135 163.367
R5447 gnd.n3176 gnd.n3140 163.367
R5448 gnd.n3155 gnd.n3140 163.367
R5449 gnd.n3166 gnd.n3155 163.367
R5450 gnd.n3166 gnd.n3156 163.367
R5451 gnd.n3162 gnd.n3156 163.367
R5452 gnd.n3162 gnd.n3161 163.367
R5453 gnd.n3161 gnd.n1811 163.367
R5454 gnd.n1811 gnd.n1798 163.367
R5455 gnd.n3383 gnd.n1798 163.367
R5456 gnd.n3383 gnd.n1799 163.367
R5457 gnd.n3379 gnd.n1799 163.367
R5458 gnd.n3379 gnd.n3378 163.367
R5459 gnd.n3378 gnd.n3377 163.367
R5460 gnd.n3377 gnd.n1802 163.367
R5461 gnd.n3293 gnd.n1802 163.367
R5462 gnd.n3367 gnd.n3293 163.367
R5463 gnd.n3367 gnd.n3294 163.367
R5464 gnd.n3363 gnd.n3294 163.367
R5465 gnd.n3363 gnd.n3362 163.367
R5466 gnd.n3362 gnd.n3298 163.367
R5467 gnd.n3309 gnd.n3298 163.367
R5468 gnd.n3309 gnd.n3306 163.367
R5469 gnd.n3351 gnd.n3306 163.367
R5470 gnd.n3351 gnd.n3307 163.367
R5471 gnd.n3347 gnd.n3307 163.367
R5472 gnd.n3347 gnd.n3313 163.367
R5473 gnd.n3326 gnd.n3313 163.367
R5474 gnd.n3337 gnd.n3326 163.367
R5475 gnd.n3337 gnd.n3327 163.367
R5476 gnd.n3333 gnd.n3327 163.367
R5477 gnd.n3333 gnd.n3332 163.367
R5478 gnd.n3332 gnd.n1734 163.367
R5479 gnd.n1734 gnd.n1721 163.367
R5480 gnd.n3789 gnd.n1721 163.367
R5481 gnd.n3789 gnd.n1722 163.367
R5482 gnd.n3785 gnd.n1722 163.367
R5483 gnd.n3785 gnd.n3784 163.367
R5484 gnd.n3784 gnd.n3783 163.367
R5485 gnd.n3783 gnd.n1725 163.367
R5486 gnd.n3467 gnd.n1725 163.367
R5487 gnd.n3773 gnd.n3467 163.367
R5488 gnd.n3773 gnd.n3468 163.367
R5489 gnd.n3769 gnd.n3468 163.367
R5490 gnd.n3769 gnd.n3768 163.367
R5491 gnd.n3768 gnd.n3472 163.367
R5492 gnd.n3484 gnd.n3472 163.367
R5493 gnd.n3484 gnd.n3480 163.367
R5494 gnd.n3757 gnd.n3480 163.367
R5495 gnd.n3757 gnd.n3482 163.367
R5496 gnd.n3753 gnd.n3482 163.367
R5497 gnd.n3753 gnd.n3488 163.367
R5498 gnd.n3496 gnd.n3488 163.367
R5499 gnd.n3742 gnd.n3496 163.367
R5500 gnd.n3742 gnd.n3497 163.367
R5501 gnd.n3738 gnd.n3497 163.367
R5502 gnd.n3738 gnd.n3737 163.367
R5503 gnd.n3737 gnd.n3500 163.367
R5504 gnd.n3509 gnd.n3500 163.367
R5505 gnd.n3728 gnd.n3509 163.367
R5506 gnd.n3728 gnd.n3510 163.367
R5507 gnd.n3724 gnd.n3510 163.367
R5508 gnd.n3724 gnd.n3723 163.367
R5509 gnd.n3723 gnd.n3514 163.367
R5510 gnd.n3541 gnd.n3514 163.367
R5511 gnd.n2748 gnd.n2747 163.367
R5512 gnd.n2747 gnd.n2746 163.367
R5513 gnd.n2743 gnd.n2742 163.367
R5514 gnd.n2740 gnd.n2674 163.367
R5515 gnd.n2736 gnd.n2734 163.367
R5516 gnd.n2732 gnd.n2676 163.367
R5517 gnd.n2728 gnd.n2726 163.367
R5518 gnd.n2724 gnd.n2678 163.367
R5519 gnd.n2720 gnd.n2718 163.367
R5520 gnd.n2716 gnd.n2680 163.367
R5521 gnd.n2712 gnd.n2710 163.367
R5522 gnd.n2708 gnd.n2682 163.367
R5523 gnd.n2704 gnd.n2702 163.367
R5524 gnd.n2700 gnd.n2684 163.367
R5525 gnd.n2696 gnd.n2694 163.367
R5526 gnd.n2691 gnd.n2690 163.367
R5527 gnd.n2831 gnd.n2829 163.367
R5528 gnd.n2827 gnd.n2629 163.367
R5529 gnd.n2822 gnd.n2820 163.367
R5530 gnd.n2818 gnd.n2633 163.367
R5531 gnd.n2814 gnd.n2812 163.367
R5532 gnd.n2810 gnd.n2635 163.367
R5533 gnd.n2806 gnd.n2804 163.367
R5534 gnd.n2802 gnd.n2637 163.367
R5535 gnd.n2798 gnd.n2796 163.367
R5536 gnd.n2794 gnd.n2639 163.367
R5537 gnd.n2790 gnd.n2788 163.367
R5538 gnd.n2786 gnd.n2641 163.367
R5539 gnd.n2782 gnd.n2780 163.367
R5540 gnd.n2778 gnd.n2643 163.367
R5541 gnd.n2774 gnd.n2772 163.367
R5542 gnd.n2770 gnd.n2645 163.367
R5543 gnd.n2752 gnd.n2648 163.367
R5544 gnd.n2756 gnd.n2648 163.367
R5545 gnd.n2756 gnd.n1955 163.367
R5546 gnd.n2937 gnd.n1955 163.367
R5547 gnd.n2937 gnd.n1939 163.367
R5548 gnd.n2941 gnd.n1939 163.367
R5549 gnd.n2942 gnd.n2941 163.367
R5550 gnd.n2942 gnd.n1950 163.367
R5551 gnd.n3031 gnd.n1950 163.367
R5552 gnd.n3031 gnd.n1953 163.367
R5553 gnd.n3027 gnd.n1953 163.367
R5554 gnd.n3027 gnd.n3026 163.367
R5555 gnd.n3026 gnd.n2946 163.367
R5556 gnd.n2954 gnd.n2946 163.367
R5557 gnd.n3016 gnd.n2954 163.367
R5558 gnd.n3016 gnd.n2955 163.367
R5559 gnd.n3012 gnd.n2955 163.367
R5560 gnd.n3012 gnd.n3011 163.367
R5561 gnd.n3011 gnd.n2959 163.367
R5562 gnd.n2969 gnd.n2959 163.367
R5563 gnd.n3001 gnd.n2969 163.367
R5564 gnd.n3001 gnd.n2970 163.367
R5565 gnd.n2997 gnd.n2970 163.367
R5566 gnd.n2997 gnd.n2996 163.367
R5567 gnd.n2996 gnd.n2974 163.367
R5568 gnd.n2982 gnd.n2974 163.367
R5569 gnd.n2986 gnd.n2982 163.367
R5570 gnd.n2986 gnd.n1879 163.367
R5571 gnd.n3108 gnd.n1879 163.367
R5572 gnd.n3108 gnd.n1864 163.367
R5573 gnd.n3112 gnd.n1864 163.367
R5574 gnd.n3113 gnd.n3112 163.367
R5575 gnd.n3113 gnd.n1876 163.367
R5576 gnd.n3204 gnd.n1876 163.367
R5577 gnd.n3204 gnd.n1877 163.367
R5578 gnd.n3200 gnd.n1877 163.367
R5579 gnd.n3200 gnd.n3199 163.367
R5580 gnd.n3199 gnd.n3117 163.367
R5581 gnd.n3128 gnd.n3117 163.367
R5582 gnd.n3189 gnd.n3128 163.367
R5583 gnd.n3189 gnd.n3129 163.367
R5584 gnd.n3185 gnd.n3129 163.367
R5585 gnd.n3185 gnd.n3184 163.367
R5586 gnd.n3184 gnd.n3133 163.367
R5587 gnd.n3144 gnd.n3133 163.367
R5588 gnd.n3174 gnd.n3144 163.367
R5589 gnd.n3174 gnd.n3145 163.367
R5590 gnd.n3170 gnd.n3145 163.367
R5591 gnd.n3170 gnd.n3154 163.367
R5592 gnd.n3154 gnd.n3153 163.367
R5593 gnd.n3153 gnd.n3149 163.367
R5594 gnd.n3149 gnd.n1808 163.367
R5595 gnd.n3282 gnd.n1808 163.367
R5596 gnd.n3283 gnd.n3282 163.367
R5597 gnd.n3283 gnd.n1794 163.367
R5598 gnd.n3287 gnd.n1794 163.367
R5599 gnd.n3288 gnd.n3287 163.367
R5600 gnd.n3288 gnd.n1805 163.367
R5601 gnd.n3375 gnd.n1805 163.367
R5602 gnd.n3375 gnd.n1806 163.367
R5603 gnd.n3371 gnd.n1806 163.367
R5604 gnd.n3371 gnd.n3370 163.367
R5605 gnd.n3370 gnd.n3292 163.367
R5606 gnd.n3300 gnd.n3292 163.367
R5607 gnd.n3360 gnd.n3300 163.367
R5608 gnd.n3360 gnd.n3301 163.367
R5609 gnd.n3356 gnd.n3301 163.367
R5610 gnd.n3356 gnd.n3355 163.367
R5611 gnd.n3355 gnd.n3305 163.367
R5612 gnd.n3315 gnd.n3305 163.367
R5613 gnd.n3345 gnd.n3315 163.367
R5614 gnd.n3345 gnd.n3316 163.367
R5615 gnd.n3341 gnd.n3316 163.367
R5616 gnd.n3341 gnd.n3325 163.367
R5617 gnd.n3325 gnd.n3324 163.367
R5618 gnd.n3324 gnd.n3320 163.367
R5619 gnd.n3320 gnd.n1732 163.367
R5620 gnd.n3453 gnd.n1732 163.367
R5621 gnd.n3454 gnd.n3453 163.367
R5622 gnd.n3454 gnd.n1719 163.367
R5623 gnd.n3461 gnd.n1719 163.367
R5624 gnd.n3462 gnd.n3461 163.367
R5625 gnd.n3462 gnd.n1728 163.367
R5626 gnd.n3781 gnd.n1728 163.367
R5627 gnd.n3781 gnd.n1730 163.367
R5628 gnd.n3777 gnd.n1730 163.367
R5629 gnd.n3777 gnd.n3776 163.367
R5630 gnd.n3776 gnd.n3466 163.367
R5631 gnd.n3474 gnd.n3466 163.367
R5632 gnd.n3766 gnd.n3474 163.367
R5633 gnd.n3766 gnd.n3475 163.367
R5634 gnd.n3762 gnd.n3475 163.367
R5635 gnd.n3762 gnd.n3761 163.367
R5636 gnd.n3761 gnd.n3479 163.367
R5637 gnd.n3490 gnd.n3479 163.367
R5638 gnd.n3751 gnd.n3490 163.367
R5639 gnd.n3751 gnd.n3491 163.367
R5640 gnd.n3747 gnd.n3491 163.367
R5641 gnd.n3747 gnd.n3746 163.367
R5642 gnd.n3746 gnd.n3495 163.367
R5643 gnd.n3502 gnd.n3495 163.367
R5644 gnd.n3735 gnd.n3502 163.367
R5645 gnd.n3735 gnd.n3503 163.367
R5646 gnd.n3731 gnd.n3503 163.367
R5647 gnd.n3731 gnd.n3730 163.367
R5648 gnd.n3730 gnd.n3507 163.367
R5649 gnd.n3516 gnd.n3507 163.367
R5650 gnd.n3721 gnd.n3516 163.367
R5651 gnd.n3721 gnd.n3517 163.367
R5652 gnd.n3717 gnd.n3517 163.367
R5653 gnd.n6511 gnd.n6510 157.424
R5654 gnd.n6512 gnd.n6511 157.424
R5655 gnd.n6512 gnd.n398 157.424
R5656 gnd.n6520 gnd.n398 157.424
R5657 gnd.n6521 gnd.n6520 157.424
R5658 gnd.n6522 gnd.n6521 157.424
R5659 gnd.n6522 gnd.n392 157.424
R5660 gnd.n6530 gnd.n392 157.424
R5661 gnd.n6531 gnd.n6530 157.424
R5662 gnd.n6532 gnd.n6531 157.424
R5663 gnd.n6532 gnd.n386 157.424
R5664 gnd.n6540 gnd.n386 157.424
R5665 gnd.n6541 gnd.n6540 157.424
R5666 gnd.n6542 gnd.n6541 157.424
R5667 gnd.n6542 gnd.n380 157.424
R5668 gnd.n6550 gnd.n380 157.424
R5669 gnd.n6551 gnd.n6550 157.424
R5670 gnd.n6552 gnd.n6551 157.424
R5671 gnd.n6552 gnd.n374 157.424
R5672 gnd.n6560 gnd.n374 157.424
R5673 gnd.n6561 gnd.n6560 157.424
R5674 gnd.n6562 gnd.n6561 157.424
R5675 gnd.n6562 gnd.n368 157.424
R5676 gnd.n6570 gnd.n368 157.424
R5677 gnd.n6571 gnd.n6570 157.424
R5678 gnd.n6572 gnd.n6571 157.424
R5679 gnd.n6572 gnd.n362 157.424
R5680 gnd.n6580 gnd.n362 157.424
R5681 gnd.n6581 gnd.n6580 157.424
R5682 gnd.n6582 gnd.n6581 157.424
R5683 gnd.n6582 gnd.n356 157.424
R5684 gnd.n6590 gnd.n356 157.424
R5685 gnd.n6591 gnd.n6590 157.424
R5686 gnd.n6592 gnd.n6591 157.424
R5687 gnd.n6592 gnd.n350 157.424
R5688 gnd.n6600 gnd.n350 157.424
R5689 gnd.n6601 gnd.n6600 157.424
R5690 gnd.n6602 gnd.n6601 157.424
R5691 gnd.n6602 gnd.n344 157.424
R5692 gnd.n6610 gnd.n344 157.424
R5693 gnd.n6611 gnd.n6610 157.424
R5694 gnd.n6612 gnd.n6611 157.424
R5695 gnd.n6612 gnd.n338 157.424
R5696 gnd.n6620 gnd.n338 157.424
R5697 gnd.n6621 gnd.n6620 157.424
R5698 gnd.n6622 gnd.n6621 157.424
R5699 gnd.n6622 gnd.n332 157.424
R5700 gnd.n6630 gnd.n332 157.424
R5701 gnd.n6631 gnd.n6630 157.424
R5702 gnd.n6632 gnd.n6631 157.424
R5703 gnd.n6632 gnd.n326 157.424
R5704 gnd.n6640 gnd.n326 157.424
R5705 gnd.n6641 gnd.n6640 157.424
R5706 gnd.n6642 gnd.n6641 157.424
R5707 gnd.n6642 gnd.n320 157.424
R5708 gnd.n6650 gnd.n320 157.424
R5709 gnd.n6651 gnd.n6650 157.424
R5710 gnd.n6652 gnd.n6651 157.424
R5711 gnd.n6652 gnd.n314 157.424
R5712 gnd.n6660 gnd.n314 157.424
R5713 gnd.n6661 gnd.n6660 157.424
R5714 gnd.n6662 gnd.n6661 157.424
R5715 gnd.n6662 gnd.n308 157.424
R5716 gnd.n6670 gnd.n308 157.424
R5717 gnd.n6671 gnd.n6670 157.424
R5718 gnd.n6672 gnd.n6671 157.424
R5719 gnd.n6672 gnd.n302 157.424
R5720 gnd.n6680 gnd.n302 157.424
R5721 gnd.n6681 gnd.n6680 157.424
R5722 gnd.n6682 gnd.n6681 157.424
R5723 gnd.n6682 gnd.n296 157.424
R5724 gnd.n6690 gnd.n296 157.424
R5725 gnd.n6691 gnd.n6690 157.424
R5726 gnd.n6692 gnd.n6691 157.424
R5727 gnd.n6692 gnd.n290 157.424
R5728 gnd.n6700 gnd.n290 157.424
R5729 gnd.n6701 gnd.n6700 157.424
R5730 gnd.n6702 gnd.n6701 157.424
R5731 gnd.n6702 gnd.n284 157.424
R5732 gnd.n6710 gnd.n284 157.424
R5733 gnd.n6711 gnd.n6710 157.424
R5734 gnd.n6713 gnd.n6711 157.424
R5735 gnd.n6713 gnd.n6712 157.424
R5736 gnd.n3538 gnd.n3537 156.462
R5737 gnd.n5740 gnd.n5708 153.042
R5738 gnd.n5804 gnd.n5803 152.079
R5739 gnd.n5772 gnd.n5771 152.079
R5740 gnd.n5740 gnd.n5739 152.079
R5741 gnd.n2661 gnd.n2660 152
R5742 gnd.n2662 gnd.n2651 152
R5743 gnd.n2664 gnd.n2663 152
R5744 gnd.n2666 gnd.n2649 152
R5745 gnd.n2668 gnd.n2667 152
R5746 gnd.n3536 gnd.n3520 152
R5747 gnd.n3528 gnd.n3521 152
R5748 gnd.n3527 gnd.n3526 152
R5749 gnd.n3525 gnd.n3522 152
R5750 gnd.n3523 gnd.t199 150.546
R5751 gnd.t101 gnd.n5782 147.661
R5752 gnd.t18 gnd.n5750 147.661
R5753 gnd.t22 gnd.n5718 147.661
R5754 gnd.t16 gnd.n5687 147.661
R5755 gnd.t274 gnd.n5655 147.661
R5756 gnd.t262 gnd.n5623 147.661
R5757 gnd.t278 gnd.n5591 147.661
R5758 gnd.t38 gnd.n5560 147.661
R5759 gnd.n3643 gnd.n3626 143.351
R5760 gnd.n2689 gnd.n2628 143.351
R5761 gnd.n2830 gnd.n2628 143.351
R5762 gnd.n2658 gnd.t128 130.484
R5763 gnd.n2667 gnd.t193 126.766
R5764 gnd.n2665 gnd.t121 126.766
R5765 gnd.n2651 gnd.t149 126.766
R5766 gnd.n2659 gnd.t212 126.766
R5767 gnd.n3524 gnd.t186 126.766
R5768 gnd.n3526 gnd.t114 126.766
R5769 gnd.n3535 gnd.t170 126.766
R5770 gnd.n3537 gnd.t135 126.766
R5771 gnd.n5799 gnd.n5798 104.615
R5772 gnd.n5798 gnd.n5776 104.615
R5773 gnd.n5791 gnd.n5776 104.615
R5774 gnd.n5791 gnd.n5790 104.615
R5775 gnd.n5790 gnd.n5780 104.615
R5776 gnd.n5783 gnd.n5780 104.615
R5777 gnd.n5767 gnd.n5766 104.615
R5778 gnd.n5766 gnd.n5744 104.615
R5779 gnd.n5759 gnd.n5744 104.615
R5780 gnd.n5759 gnd.n5758 104.615
R5781 gnd.n5758 gnd.n5748 104.615
R5782 gnd.n5751 gnd.n5748 104.615
R5783 gnd.n5735 gnd.n5734 104.615
R5784 gnd.n5734 gnd.n5712 104.615
R5785 gnd.n5727 gnd.n5712 104.615
R5786 gnd.n5727 gnd.n5726 104.615
R5787 gnd.n5726 gnd.n5716 104.615
R5788 gnd.n5719 gnd.n5716 104.615
R5789 gnd.n5704 gnd.n5703 104.615
R5790 gnd.n5703 gnd.n5681 104.615
R5791 gnd.n5696 gnd.n5681 104.615
R5792 gnd.n5696 gnd.n5695 104.615
R5793 gnd.n5695 gnd.n5685 104.615
R5794 gnd.n5688 gnd.n5685 104.615
R5795 gnd.n5672 gnd.n5671 104.615
R5796 gnd.n5671 gnd.n5649 104.615
R5797 gnd.n5664 gnd.n5649 104.615
R5798 gnd.n5664 gnd.n5663 104.615
R5799 gnd.n5663 gnd.n5653 104.615
R5800 gnd.n5656 gnd.n5653 104.615
R5801 gnd.n5640 gnd.n5639 104.615
R5802 gnd.n5639 gnd.n5617 104.615
R5803 gnd.n5632 gnd.n5617 104.615
R5804 gnd.n5632 gnd.n5631 104.615
R5805 gnd.n5631 gnd.n5621 104.615
R5806 gnd.n5624 gnd.n5621 104.615
R5807 gnd.n5608 gnd.n5607 104.615
R5808 gnd.n5607 gnd.n5585 104.615
R5809 gnd.n5600 gnd.n5585 104.615
R5810 gnd.n5600 gnd.n5599 104.615
R5811 gnd.n5599 gnd.n5589 104.615
R5812 gnd.n5592 gnd.n5589 104.615
R5813 gnd.n5577 gnd.n5576 104.615
R5814 gnd.n5576 gnd.n5554 104.615
R5815 gnd.n5569 gnd.n5554 104.615
R5816 gnd.n5569 gnd.n5568 104.615
R5817 gnd.n5568 gnd.n5558 104.615
R5818 gnd.n5561 gnd.n5558 104.615
R5819 gnd.n5131 gnd.t127 100.632
R5820 gnd.n4597 gnd.t168 100.632
R5821 gnd.n6954 gnd.n93 99.6594
R5822 gnd.n6952 gnd.n6951 99.6594
R5823 gnd.n6947 gnd.n101 99.6594
R5824 gnd.n6945 gnd.n6944 99.6594
R5825 gnd.n6940 gnd.n108 99.6594
R5826 gnd.n6938 gnd.n6937 99.6594
R5827 gnd.n6933 gnd.n115 99.6594
R5828 gnd.n6931 gnd.n6930 99.6594
R5829 gnd.n6923 gnd.n122 99.6594
R5830 gnd.n6921 gnd.n6920 99.6594
R5831 gnd.n6916 gnd.n129 99.6594
R5832 gnd.n6914 gnd.n6913 99.6594
R5833 gnd.n6909 gnd.n136 99.6594
R5834 gnd.n6907 gnd.n6906 99.6594
R5835 gnd.n6902 gnd.n143 99.6594
R5836 gnd.n6900 gnd.n6899 99.6594
R5837 gnd.n6895 gnd.n150 99.6594
R5838 gnd.n6893 gnd.n6892 99.6594
R5839 gnd.n155 gnd.n154 99.6594
R5840 gnd.n4228 gnd.n4227 99.6594
R5841 gnd.n4222 gnd.n1283 99.6594
R5842 gnd.n4219 gnd.n1284 99.6594
R5843 gnd.n4215 gnd.n1285 99.6594
R5844 gnd.n4211 gnd.n1286 99.6594
R5845 gnd.n4207 gnd.n1287 99.6594
R5846 gnd.n4203 gnd.n1288 99.6594
R5847 gnd.n4199 gnd.n1289 99.6594
R5848 gnd.n4194 gnd.n1291 99.6594
R5849 gnd.n4190 gnd.n1292 99.6594
R5850 gnd.n4186 gnd.n1293 99.6594
R5851 gnd.n4182 gnd.n1294 99.6594
R5852 gnd.n4178 gnd.n1295 99.6594
R5853 gnd.n4174 gnd.n1296 99.6594
R5854 gnd.n4170 gnd.n1297 99.6594
R5855 gnd.n4166 gnd.n1298 99.6594
R5856 gnd.n4162 gnd.n1299 99.6594
R5857 gnd.n1355 gnd.n1300 99.6594
R5858 gnd.n2861 gnd.n2860 99.6594
R5859 gnd.n2856 gnd.n2136 99.6594
R5860 gnd.n2852 gnd.n2135 99.6594
R5861 gnd.n2848 gnd.n2134 99.6594
R5862 gnd.n2844 gnd.n2133 99.6594
R5863 gnd.n2840 gnd.n2132 99.6594
R5864 gnd.n2836 gnd.n2131 99.6594
R5865 gnd.n2620 gnd.n2129 99.6594
R5866 gnd.n2618 gnd.n2128 99.6594
R5867 gnd.n2614 gnd.n2127 99.6594
R5868 gnd.n2610 gnd.n2126 99.6594
R5869 gnd.n2606 gnd.n2125 99.6594
R5870 gnd.n2602 gnd.n2124 99.6594
R5871 gnd.n2598 gnd.n2123 99.6594
R5872 gnd.n2594 gnd.n2122 99.6594
R5873 gnd.n2590 gnd.n2121 99.6594
R5874 gnd.n2586 gnd.n2120 99.6594
R5875 gnd.n2178 gnd.n2119 99.6594
R5876 gnd.n4573 gnd.n4572 99.6594
R5877 gnd.n4567 gnd.n878 99.6594
R5878 gnd.n4564 gnd.n879 99.6594
R5879 gnd.n4560 gnd.n880 99.6594
R5880 gnd.n4556 gnd.n881 99.6594
R5881 gnd.n4552 gnd.n882 99.6594
R5882 gnd.n4548 gnd.n883 99.6594
R5883 gnd.n4544 gnd.n884 99.6594
R5884 gnd.n4540 gnd.n885 99.6594
R5885 gnd.n4535 gnd.n886 99.6594
R5886 gnd.n4531 gnd.n887 99.6594
R5887 gnd.n4527 gnd.n888 99.6594
R5888 gnd.n4523 gnd.n889 99.6594
R5889 gnd.n4519 gnd.n890 99.6594
R5890 gnd.n4515 gnd.n891 99.6594
R5891 gnd.n4511 gnd.n892 99.6594
R5892 gnd.n4507 gnd.n893 99.6594
R5893 gnd.n4503 gnd.n894 99.6594
R5894 gnd.n949 gnd.n895 99.6594
R5895 gnd.n5913 gnd.n5912 99.6594
R5896 gnd.n5908 gnd.n4581 99.6594
R5897 gnd.n5904 gnd.n4580 99.6594
R5898 gnd.n5900 gnd.n4579 99.6594
R5899 gnd.n5896 gnd.n4578 99.6594
R5900 gnd.n5892 gnd.n4577 99.6594
R5901 gnd.n5888 gnd.n4576 99.6594
R5902 gnd.n5815 gnd.n4575 99.6594
R5903 gnd.n5164 gnd.n5163 99.6594
R5904 gnd.n5158 gnd.n5106 99.6594
R5905 gnd.n5155 gnd.n5107 99.6594
R5906 gnd.n5151 gnd.n5108 99.6594
R5907 gnd.n5147 gnd.n5109 99.6594
R5908 gnd.n5143 gnd.n5110 99.6594
R5909 gnd.n5139 gnd.n5111 99.6594
R5910 gnd.n5135 gnd.n5112 99.6594
R5911 gnd.n5878 gnd.n865 99.6594
R5912 gnd.n5874 gnd.n866 99.6594
R5913 gnd.n5870 gnd.n867 99.6594
R5914 gnd.n5866 gnd.n868 99.6594
R5915 gnd.n5862 gnd.n869 99.6594
R5916 gnd.n5858 gnd.n870 99.6594
R5917 gnd.n5854 gnd.n871 99.6594
R5918 gnd.n5850 gnd.n872 99.6594
R5919 gnd.n5846 gnd.n873 99.6594
R5920 gnd.n5842 gnd.n874 99.6594
R5921 gnd.n5838 gnd.n875 99.6594
R5922 gnd.n5834 gnd.n876 99.6594
R5923 gnd.n5830 gnd.n877 99.6594
R5924 gnd.n5036 gnd.n4946 99.6594
R5925 gnd.n5034 gnd.n4949 99.6594
R5926 gnd.n5030 gnd.n5029 99.6594
R5927 gnd.n5023 gnd.n4954 99.6594
R5928 gnd.n5022 gnd.n5021 99.6594
R5929 gnd.n5015 gnd.n4960 99.6594
R5930 gnd.n5014 gnd.n5013 99.6594
R5931 gnd.n5007 gnd.n4966 99.6594
R5932 gnd.n5006 gnd.n5005 99.6594
R5933 gnd.n4999 gnd.n4972 99.6594
R5934 gnd.n4998 gnd.n4997 99.6594
R5935 gnd.n4990 gnd.n4978 99.6594
R5936 gnd.n4989 gnd.n4988 99.6594
R5937 gnd.n6803 gnd.n6802 99.6594
R5938 gnd.n6808 gnd.n6807 99.6594
R5939 gnd.n6811 gnd.n6810 99.6594
R5940 gnd.n6816 gnd.n6815 99.6594
R5941 gnd.n6819 gnd.n6818 99.6594
R5942 gnd.n6824 gnd.n6823 99.6594
R5943 gnd.n6827 gnd.n6826 99.6594
R5944 gnd.n6832 gnd.n6831 99.6594
R5945 gnd.n6835 gnd.n80 99.6594
R5946 gnd.n1365 gnd.n1301 99.6594
R5947 gnd.n1553 gnd.n1302 99.6594
R5948 gnd.n1544 gnd.n1303 99.6594
R5949 gnd.n1569 gnd.n1304 99.6594
R5950 gnd.n1535 gnd.n1305 99.6594
R5951 gnd.n1586 gnd.n1306 99.6594
R5952 gnd.n1526 gnd.n1307 99.6594
R5953 gnd.n1603 gnd.n1308 99.6594
R5954 gnd.n1517 gnd.n1309 99.6594
R5955 gnd.n2053 gnd.n2019 99.6594
R5956 gnd.n2066 gnd.n2020 99.6594
R5957 gnd.n2077 gnd.n2021 99.6594
R5958 gnd.n2039 gnd.n2022 99.6594
R5959 gnd.n2090 gnd.n2023 99.6594
R5960 gnd.n2101 gnd.n2024 99.6594
R5961 gnd.n2026 gnd.n2025 99.6594
R5962 gnd.n2117 gnd.n2116 99.6594
R5963 gnd.n2864 gnd.n2863 99.6594
R5964 gnd.n2418 gnd.n896 99.6594
R5965 gnd.n2415 gnd.n897 99.6594
R5966 gnd.n2411 gnd.n898 99.6594
R5967 gnd.n2407 gnd.n899 99.6594
R5968 gnd.n2403 gnd.n900 99.6594
R5969 gnd.n2399 gnd.n901 99.6594
R5970 gnd.n2395 gnd.n902 99.6594
R5971 gnd.n2391 gnd.n903 99.6594
R5972 gnd.n2387 gnd.n904 99.6594
R5973 gnd.n2416 gnd.n896 99.6594
R5974 gnd.n2412 gnd.n897 99.6594
R5975 gnd.n2408 gnd.n898 99.6594
R5976 gnd.n2404 gnd.n899 99.6594
R5977 gnd.n2400 gnd.n900 99.6594
R5978 gnd.n2396 gnd.n901 99.6594
R5979 gnd.n2392 gnd.n902 99.6594
R5980 gnd.n2388 gnd.n903 99.6594
R5981 gnd.n2376 gnd.n904 99.6594
R5982 gnd.n2863 gnd.n2017 99.6594
R5983 gnd.n2117 gnd.n2115 99.6594
R5984 gnd.n2102 gnd.n2025 99.6594
R5985 gnd.n2089 gnd.n2024 99.6594
R5986 gnd.n2040 gnd.n2023 99.6594
R5987 gnd.n2078 gnd.n2022 99.6594
R5988 gnd.n2065 gnd.n2021 99.6594
R5989 gnd.n2054 gnd.n2020 99.6594
R5990 gnd.n2050 gnd.n2019 99.6594
R5991 gnd.n1552 gnd.n1301 99.6594
R5992 gnd.n1543 gnd.n1302 99.6594
R5993 gnd.n1568 gnd.n1303 99.6594
R5994 gnd.n1534 gnd.n1304 99.6594
R5995 gnd.n1585 gnd.n1305 99.6594
R5996 gnd.n1525 gnd.n1306 99.6594
R5997 gnd.n1602 gnd.n1307 99.6594
R5998 gnd.n1516 gnd.n1308 99.6594
R5999 gnd.n1512 gnd.n1309 99.6594
R6000 gnd.n6836 gnd.n6835 99.6594
R6001 gnd.n6831 gnd.n6830 99.6594
R6002 gnd.n6826 gnd.n6825 99.6594
R6003 gnd.n6823 gnd.n6822 99.6594
R6004 gnd.n6818 gnd.n6817 99.6594
R6005 gnd.n6815 gnd.n6814 99.6594
R6006 gnd.n6810 gnd.n6809 99.6594
R6007 gnd.n6807 gnd.n6806 99.6594
R6008 gnd.n6802 gnd.n6801 99.6594
R6009 gnd.n5037 gnd.n5036 99.6594
R6010 gnd.n5031 gnd.n4949 99.6594
R6011 gnd.n5029 gnd.n5028 99.6594
R6012 gnd.n5024 gnd.n5023 99.6594
R6013 gnd.n5021 gnd.n5020 99.6594
R6014 gnd.n5016 gnd.n5015 99.6594
R6015 gnd.n5013 gnd.n5012 99.6594
R6016 gnd.n5008 gnd.n5007 99.6594
R6017 gnd.n5005 gnd.n5004 99.6594
R6018 gnd.n5000 gnd.n4999 99.6594
R6019 gnd.n4997 gnd.n4996 99.6594
R6020 gnd.n4991 gnd.n4990 99.6594
R6021 gnd.n4988 gnd.n4944 99.6594
R6022 gnd.n5833 gnd.n877 99.6594
R6023 gnd.n5837 gnd.n876 99.6594
R6024 gnd.n5841 gnd.n875 99.6594
R6025 gnd.n5845 gnd.n874 99.6594
R6026 gnd.n5849 gnd.n873 99.6594
R6027 gnd.n5853 gnd.n872 99.6594
R6028 gnd.n5857 gnd.n871 99.6594
R6029 gnd.n5861 gnd.n870 99.6594
R6030 gnd.n5865 gnd.n869 99.6594
R6031 gnd.n5869 gnd.n868 99.6594
R6032 gnd.n5873 gnd.n867 99.6594
R6033 gnd.n5877 gnd.n866 99.6594
R6034 gnd.n4601 gnd.n865 99.6594
R6035 gnd.n5164 gnd.n5114 99.6594
R6036 gnd.n5156 gnd.n5106 99.6594
R6037 gnd.n5152 gnd.n5107 99.6594
R6038 gnd.n5148 gnd.n5108 99.6594
R6039 gnd.n5144 gnd.n5109 99.6594
R6040 gnd.n5140 gnd.n5110 99.6594
R6041 gnd.n5136 gnd.n5111 99.6594
R6042 gnd.n5112 gnd.n4906 99.6594
R6043 gnd.n5887 gnd.n4575 99.6594
R6044 gnd.n5891 gnd.n4576 99.6594
R6045 gnd.n5895 gnd.n4577 99.6594
R6046 gnd.n5899 gnd.n4578 99.6594
R6047 gnd.n5903 gnd.n4579 99.6594
R6048 gnd.n5907 gnd.n4580 99.6594
R6049 gnd.n4582 gnd.n4581 99.6594
R6050 gnd.n5913 gnd.n862 99.6594
R6051 gnd.n4573 gnd.n908 99.6594
R6052 gnd.n4565 gnd.n878 99.6594
R6053 gnd.n4561 gnd.n879 99.6594
R6054 gnd.n4557 gnd.n880 99.6594
R6055 gnd.n4553 gnd.n881 99.6594
R6056 gnd.n4549 gnd.n882 99.6594
R6057 gnd.n4545 gnd.n883 99.6594
R6058 gnd.n4541 gnd.n884 99.6594
R6059 gnd.n4536 gnd.n885 99.6594
R6060 gnd.n4532 gnd.n886 99.6594
R6061 gnd.n4528 gnd.n887 99.6594
R6062 gnd.n4524 gnd.n888 99.6594
R6063 gnd.n4520 gnd.n889 99.6594
R6064 gnd.n4516 gnd.n890 99.6594
R6065 gnd.n4512 gnd.n891 99.6594
R6066 gnd.n4508 gnd.n892 99.6594
R6067 gnd.n4504 gnd.n893 99.6594
R6068 gnd.n948 gnd.n894 99.6594
R6069 gnd.n4496 gnd.n895 99.6594
R6070 gnd.n2585 gnd.n2119 99.6594
R6071 gnd.n2589 gnd.n2120 99.6594
R6072 gnd.n2593 gnd.n2121 99.6594
R6073 gnd.n2597 gnd.n2122 99.6594
R6074 gnd.n2601 gnd.n2123 99.6594
R6075 gnd.n2605 gnd.n2124 99.6594
R6076 gnd.n2609 gnd.n2125 99.6594
R6077 gnd.n2613 gnd.n2126 99.6594
R6078 gnd.n2617 gnd.n2127 99.6594
R6079 gnd.n2621 gnd.n2128 99.6594
R6080 gnd.n2835 gnd.n2130 99.6594
R6081 gnd.n2839 gnd.n2131 99.6594
R6082 gnd.n2843 gnd.n2132 99.6594
R6083 gnd.n2847 gnd.n2133 99.6594
R6084 gnd.n2851 gnd.n2134 99.6594
R6085 gnd.n2855 gnd.n2135 99.6594
R6086 gnd.n2138 gnd.n2136 99.6594
R6087 gnd.n2861 gnd.n2137 99.6594
R6088 gnd.n4228 gnd.n1313 99.6594
R6089 gnd.n4220 gnd.n1283 99.6594
R6090 gnd.n4216 gnd.n1284 99.6594
R6091 gnd.n4212 gnd.n1285 99.6594
R6092 gnd.n4208 gnd.n1286 99.6594
R6093 gnd.n4204 gnd.n1287 99.6594
R6094 gnd.n4200 gnd.n1288 99.6594
R6095 gnd.n4195 gnd.n1290 99.6594
R6096 gnd.n4191 gnd.n1291 99.6594
R6097 gnd.n4187 gnd.n1292 99.6594
R6098 gnd.n4183 gnd.n1293 99.6594
R6099 gnd.n4179 gnd.n1294 99.6594
R6100 gnd.n4175 gnd.n1295 99.6594
R6101 gnd.n4171 gnd.n1296 99.6594
R6102 gnd.n4167 gnd.n1297 99.6594
R6103 gnd.n4163 gnd.n1298 99.6594
R6104 gnd.n1354 gnd.n1299 99.6594
R6105 gnd.n4155 gnd.n1300 99.6594
R6106 gnd.n154 gnd.n151 99.6594
R6107 gnd.n6894 gnd.n6893 99.6594
R6108 gnd.n150 gnd.n144 99.6594
R6109 gnd.n6901 gnd.n6900 99.6594
R6110 gnd.n143 gnd.n137 99.6594
R6111 gnd.n6908 gnd.n6907 99.6594
R6112 gnd.n136 gnd.n130 99.6594
R6113 gnd.n6915 gnd.n6914 99.6594
R6114 gnd.n129 gnd.n123 99.6594
R6115 gnd.n6922 gnd.n6921 99.6594
R6116 gnd.n122 gnd.n116 99.6594
R6117 gnd.n6932 gnd.n6931 99.6594
R6118 gnd.n115 gnd.n109 99.6594
R6119 gnd.n6939 gnd.n6938 99.6594
R6120 gnd.n108 gnd.n102 99.6594
R6121 gnd.n6946 gnd.n6945 99.6594
R6122 gnd.n101 gnd.n95 99.6594
R6123 gnd.n6953 gnd.n6952 99.6594
R6124 gnd.n93 gnd.n90 99.6594
R6125 gnd.n2057 gnd.n1986 99.6594
R6126 gnd.n2059 gnd.n1987 99.6594
R6127 gnd.n2072 gnd.n1988 99.6594
R6128 gnd.n2044 gnd.n1989 99.6594
R6129 gnd.n2083 gnd.n1990 99.6594
R6130 gnd.n2096 gnd.n1991 99.6594
R6131 gnd.n2032 gnd.n1992 99.6594
R6132 gnd.n2110 gnd.n1993 99.6594
R6133 gnd.n2012 gnd.n1994 99.6594
R6134 gnd.n2870 gnd.n1995 99.6594
R6135 gnd.n2879 gnd.n1996 99.6594
R6136 gnd.n2881 gnd.n1997 99.6594
R6137 gnd.n2889 gnd.n1998 99.6594
R6138 gnd.n2899 gnd.n1999 99.6594
R6139 gnd.n2060 gnd.n1986 99.6594
R6140 gnd.n2071 gnd.n1987 99.6594
R6141 gnd.n2043 gnd.n1988 99.6594
R6142 gnd.n2084 gnd.n1989 99.6594
R6143 gnd.n2095 gnd.n1990 99.6594
R6144 gnd.n2031 gnd.n1991 99.6594
R6145 gnd.n2109 gnd.n1992 99.6594
R6146 gnd.n2011 gnd.n1993 99.6594
R6147 gnd.n2871 gnd.n1994 99.6594
R6148 gnd.n2878 gnd.n1995 99.6594
R6149 gnd.n2882 gnd.n1996 99.6594
R6150 gnd.n2888 gnd.n1997 99.6594
R6151 gnd.n2892 gnd.n1998 99.6594
R6152 gnd.n2899 gnd.n2898 99.6594
R6153 gnd.n1558 gnd.n1271 99.6594
R6154 gnd.n1561 gnd.n1560 99.6594
R6155 gnd.n1575 gnd.n1574 99.6594
R6156 gnd.n1578 gnd.n1577 99.6594
R6157 gnd.n1592 gnd.n1591 99.6594
R6158 gnd.n1595 gnd.n1594 99.6594
R6159 gnd.n1609 gnd.n1608 99.6594
R6160 gnd.n1612 gnd.n1611 99.6594
R6161 gnd.n1624 gnd.n1623 99.6594
R6162 gnd.n1627 gnd.n1626 99.6594
R6163 gnd.n1630 gnd.n1629 99.6594
R6164 gnd.n1635 gnd.n1634 99.6594
R6165 gnd.n1638 gnd.n1637 99.6594
R6166 gnd.n3891 gnd.n3890 99.6594
R6167 gnd.n3892 gnd.n3891 99.6594
R6168 gnd.n1639 gnd.n1638 99.6594
R6169 gnd.n1636 gnd.n1635 99.6594
R6170 gnd.n1631 gnd.n1630 99.6594
R6171 gnd.n1628 gnd.n1627 99.6594
R6172 gnd.n1625 gnd.n1624 99.6594
R6173 gnd.n1611 gnd.n1508 99.6594
R6174 gnd.n1610 gnd.n1609 99.6594
R6175 gnd.n1594 gnd.n1520 99.6594
R6176 gnd.n1593 gnd.n1592 99.6594
R6177 gnd.n1577 gnd.n1529 99.6594
R6178 gnd.n1576 gnd.n1575 99.6594
R6179 gnd.n1560 gnd.n1538 99.6594
R6180 gnd.n1559 gnd.n1558 99.6594
R6181 gnd.n2003 gnd.t192 98.63
R6182 gnd.n6833 gnd.t178 98.63
R6183 gnd.n1513 gnd.t165 98.63
R6184 gnd.n2015 gnd.t184 98.63
R6185 gnd.n1334 gnd.t162 98.63
R6186 gnd.n1356 gnd.t134 98.63
R6187 gnd.n157 gnd.t119 98.63
R6188 gnd.n6925 gnd.t147 98.63
R6189 gnd.n928 gnd.t217 98.63
R6190 gnd.n950 gnd.t208 98.63
R6191 gnd.n2377 gnd.t205 98.63
R6192 gnd.n2180 gnd.t140 98.63
R6193 gnd.n2158 gnd.t181 98.63
R6194 gnd.n3900 gnd.t175 98.63
R6195 gnd.n2630 gnd.t211 96.6984
R6196 gnd.n3644 gnd.t144 96.6984
R6197 gnd.n2685 gnd.t159 96.6906
R6198 gnd.n3559 gnd.t197 96.6906
R6199 gnd.n6712 gnd.n83 94.4549
R6200 gnd.n2658 gnd.n2657 81.8399
R6201 gnd.n5132 gnd.t126 74.8376
R6202 gnd.n4598 gnd.t169 74.8376
R6203 gnd.n2631 gnd.t210 72.8438
R6204 gnd.n3645 gnd.t145 72.8438
R6205 gnd.n2659 gnd.n2652 72.8411
R6206 gnd.n2665 gnd.n2650 72.8411
R6207 gnd.n3535 gnd.n3534 72.8411
R6208 gnd.n2004 gnd.t191 72.836
R6209 gnd.n2686 gnd.t158 72.836
R6210 gnd.n3560 gnd.t198 72.836
R6211 gnd.n6834 gnd.t179 72.836
R6212 gnd.n1514 gnd.t164 72.836
R6213 gnd.n2016 gnd.t185 72.836
R6214 gnd.n1335 gnd.t161 72.836
R6215 gnd.n1357 gnd.t133 72.836
R6216 gnd.n158 gnd.t120 72.836
R6217 gnd.n6926 gnd.t148 72.836
R6218 gnd.n929 gnd.t216 72.836
R6219 gnd.n951 gnd.t207 72.836
R6220 gnd.n2378 gnd.t204 72.836
R6221 gnd.n2181 gnd.t141 72.836
R6222 gnd.n2159 gnd.t182 72.836
R6223 gnd.n3901 gnd.t176 72.836
R6224 gnd.n3563 gnd.n3543 71.676
R6225 gnd.n3567 gnd.n3544 71.676
R6226 gnd.n3571 gnd.n3545 71.676
R6227 gnd.n3575 gnd.n3546 71.676
R6228 gnd.n3579 gnd.n3547 71.676
R6229 gnd.n3583 gnd.n3548 71.676
R6230 gnd.n3587 gnd.n3549 71.676
R6231 gnd.n3591 gnd.n3550 71.676
R6232 gnd.n3595 gnd.n3551 71.676
R6233 gnd.n3599 gnd.n3552 71.676
R6234 gnd.n3603 gnd.n3553 71.676
R6235 gnd.n3607 gnd.n3554 71.676
R6236 gnd.n3611 gnd.n3555 71.676
R6237 gnd.n3615 gnd.n3556 71.676
R6238 gnd.n3620 gnd.n3557 71.676
R6239 gnd.n3624 gnd.n3558 71.676
R6240 gnd.n3713 gnd.n3643 71.676
R6241 gnd.n3709 gnd.n3642 71.676
R6242 gnd.n3704 gnd.n3641 71.676
R6243 gnd.n3700 gnd.n3640 71.676
R6244 gnd.n3696 gnd.n3639 71.676
R6245 gnd.n3692 gnd.n3638 71.676
R6246 gnd.n3688 gnd.n3637 71.676
R6247 gnd.n3684 gnd.n3636 71.676
R6248 gnd.n3680 gnd.n3635 71.676
R6249 gnd.n3676 gnd.n3634 71.676
R6250 gnd.n3672 gnd.n3633 71.676
R6251 gnd.n3668 gnd.n3632 71.676
R6252 gnd.n3664 gnd.n3631 71.676
R6253 gnd.n3660 gnd.n3630 71.676
R6254 gnd.n3656 gnd.n3629 71.676
R6255 gnd.n3652 gnd.n3628 71.676
R6256 gnd.n3648 gnd.n3627 71.676
R6257 gnd.n2751 gnd.n2670 71.676
R6258 gnd.n2746 gnd.n2672 71.676
R6259 gnd.n2742 gnd.n2741 71.676
R6260 gnd.n2735 gnd.n2674 71.676
R6261 gnd.n2734 gnd.n2733 71.676
R6262 gnd.n2727 gnd.n2676 71.676
R6263 gnd.n2726 gnd.n2725 71.676
R6264 gnd.n2719 gnd.n2678 71.676
R6265 gnd.n2718 gnd.n2717 71.676
R6266 gnd.n2711 gnd.n2680 71.676
R6267 gnd.n2710 gnd.n2709 71.676
R6268 gnd.n2703 gnd.n2682 71.676
R6269 gnd.n2702 gnd.n2701 71.676
R6270 gnd.n2695 gnd.n2684 71.676
R6271 gnd.n2694 gnd.n2688 71.676
R6272 gnd.n2690 gnd.n2689 71.676
R6273 gnd.n2829 gnd.n2828 71.676
R6274 gnd.n2821 gnd.n2629 71.676
R6275 gnd.n2820 gnd.n2819 71.676
R6276 gnd.n2813 gnd.n2633 71.676
R6277 gnd.n2812 gnd.n2811 71.676
R6278 gnd.n2805 gnd.n2635 71.676
R6279 gnd.n2804 gnd.n2803 71.676
R6280 gnd.n2797 gnd.n2637 71.676
R6281 gnd.n2796 gnd.n2795 71.676
R6282 gnd.n2789 gnd.n2639 71.676
R6283 gnd.n2788 gnd.n2787 71.676
R6284 gnd.n2781 gnd.n2641 71.676
R6285 gnd.n2780 gnd.n2779 71.676
R6286 gnd.n2773 gnd.n2643 71.676
R6287 gnd.n2772 gnd.n2771 71.676
R6288 gnd.n2765 gnd.n2645 71.676
R6289 gnd.n2748 gnd.n2670 71.676
R6290 gnd.n2743 gnd.n2672 71.676
R6291 gnd.n2741 gnd.n2740 71.676
R6292 gnd.n2736 gnd.n2735 71.676
R6293 gnd.n2733 gnd.n2732 71.676
R6294 gnd.n2728 gnd.n2727 71.676
R6295 gnd.n2725 gnd.n2724 71.676
R6296 gnd.n2720 gnd.n2719 71.676
R6297 gnd.n2717 gnd.n2716 71.676
R6298 gnd.n2712 gnd.n2711 71.676
R6299 gnd.n2709 gnd.n2708 71.676
R6300 gnd.n2704 gnd.n2703 71.676
R6301 gnd.n2701 gnd.n2700 71.676
R6302 gnd.n2696 gnd.n2695 71.676
R6303 gnd.n2691 gnd.n2688 71.676
R6304 gnd.n2831 gnd.n2830 71.676
R6305 gnd.n2828 gnd.n2827 71.676
R6306 gnd.n2822 gnd.n2821 71.676
R6307 gnd.n2819 gnd.n2818 71.676
R6308 gnd.n2814 gnd.n2813 71.676
R6309 gnd.n2811 gnd.n2810 71.676
R6310 gnd.n2806 gnd.n2805 71.676
R6311 gnd.n2803 gnd.n2802 71.676
R6312 gnd.n2798 gnd.n2797 71.676
R6313 gnd.n2795 gnd.n2794 71.676
R6314 gnd.n2790 gnd.n2789 71.676
R6315 gnd.n2787 gnd.n2786 71.676
R6316 gnd.n2782 gnd.n2781 71.676
R6317 gnd.n2779 gnd.n2778 71.676
R6318 gnd.n2774 gnd.n2773 71.676
R6319 gnd.n2771 gnd.n2770 71.676
R6320 gnd.n2766 gnd.n2765 71.676
R6321 gnd.n3651 gnd.n3627 71.676
R6322 gnd.n3655 gnd.n3628 71.676
R6323 gnd.n3659 gnd.n3629 71.676
R6324 gnd.n3663 gnd.n3630 71.676
R6325 gnd.n3667 gnd.n3631 71.676
R6326 gnd.n3671 gnd.n3632 71.676
R6327 gnd.n3675 gnd.n3633 71.676
R6328 gnd.n3679 gnd.n3634 71.676
R6329 gnd.n3683 gnd.n3635 71.676
R6330 gnd.n3687 gnd.n3636 71.676
R6331 gnd.n3691 gnd.n3637 71.676
R6332 gnd.n3695 gnd.n3638 71.676
R6333 gnd.n3699 gnd.n3639 71.676
R6334 gnd.n3703 gnd.n3640 71.676
R6335 gnd.n3708 gnd.n3641 71.676
R6336 gnd.n3712 gnd.n3642 71.676
R6337 gnd.n3626 gnd.n3625 71.676
R6338 gnd.n3621 gnd.n3558 71.676
R6339 gnd.n3616 gnd.n3557 71.676
R6340 gnd.n3612 gnd.n3556 71.676
R6341 gnd.n3608 gnd.n3555 71.676
R6342 gnd.n3604 gnd.n3554 71.676
R6343 gnd.n3600 gnd.n3553 71.676
R6344 gnd.n3596 gnd.n3552 71.676
R6345 gnd.n3592 gnd.n3551 71.676
R6346 gnd.n3588 gnd.n3550 71.676
R6347 gnd.n3584 gnd.n3549 71.676
R6348 gnd.n3580 gnd.n3548 71.676
R6349 gnd.n3576 gnd.n3547 71.676
R6350 gnd.n3572 gnd.n3546 71.676
R6351 gnd.n3568 gnd.n3545 71.676
R6352 gnd.n3564 gnd.n3544 71.676
R6353 gnd.n3543 gnd.n3540 71.676
R6354 gnd.n8 gnd.t229 69.1507
R6355 gnd.n14 gnd.t231 68.4792
R6356 gnd.n13 gnd.t271 68.4792
R6357 gnd.n12 gnd.t40 68.4792
R6358 gnd.n11 gnd.t289 68.4792
R6359 gnd.n10 gnd.t109 68.4792
R6360 gnd.n9 gnd.t225 68.4792
R6361 gnd.n8 gnd.t276 68.4792
R6362 gnd.n5044 gnd.n4945 64.369
R6363 gnd.n4574 gnd.n906 63.0944
R6364 gnd.n2824 gnd.n2631 59.5399
R6365 gnd.n3706 gnd.n3645 59.5399
R6366 gnd.n2687 gnd.n2686 59.5399
R6367 gnd.n3618 gnd.n3560 59.5399
R6368 gnd.n2669 gnd.n2668 59.1804
R6369 gnd.n5914 gnd.n863 57.3586
R6370 gnd.n4755 gnd.t20 56.607
R6371 gnd.n40 gnd.t36 56.607
R6372 gnd.n4732 gnd.t236 56.407
R6373 gnd.n4743 gnd.t57 56.407
R6374 gnd.n17 gnd.t78 56.407
R6375 gnd.n28 gnd.t6 56.407
R6376 gnd.n4764 gnd.t260 55.8337
R6377 gnd.n4741 gnd.t265 55.8337
R6378 gnd.n4752 gnd.t241 55.8337
R6379 gnd.n49 gnd.t269 55.8337
R6380 gnd.n26 gnd.t291 55.8337
R6381 gnd.n37 gnd.t264 55.8337
R6382 gnd.n2656 gnd.n2655 54.358
R6383 gnd.n3532 gnd.n3531 54.358
R6384 gnd.n4755 gnd.n4754 53.0052
R6385 gnd.n4757 gnd.n4756 53.0052
R6386 gnd.n4759 gnd.n4758 53.0052
R6387 gnd.n4761 gnd.n4760 53.0052
R6388 gnd.n4763 gnd.n4762 53.0052
R6389 gnd.n4732 gnd.n4731 53.0052
R6390 gnd.n4734 gnd.n4733 53.0052
R6391 gnd.n4736 gnd.n4735 53.0052
R6392 gnd.n4738 gnd.n4737 53.0052
R6393 gnd.n4740 gnd.n4739 53.0052
R6394 gnd.n4743 gnd.n4742 53.0052
R6395 gnd.n4745 gnd.n4744 53.0052
R6396 gnd.n4747 gnd.n4746 53.0052
R6397 gnd.n4749 gnd.n4748 53.0052
R6398 gnd.n4751 gnd.n4750 53.0052
R6399 gnd.n48 gnd.n47 53.0052
R6400 gnd.n46 gnd.n45 53.0052
R6401 gnd.n44 gnd.n43 53.0052
R6402 gnd.n42 gnd.n41 53.0052
R6403 gnd.n40 gnd.n39 53.0052
R6404 gnd.n25 gnd.n24 53.0052
R6405 gnd.n23 gnd.n22 53.0052
R6406 gnd.n21 gnd.n20 53.0052
R6407 gnd.n19 gnd.n18 53.0052
R6408 gnd.n17 gnd.n16 53.0052
R6409 gnd.n36 gnd.n35 53.0052
R6410 gnd.n34 gnd.n33 53.0052
R6411 gnd.n32 gnd.n31 53.0052
R6412 gnd.n30 gnd.n29 53.0052
R6413 gnd.n28 gnd.n27 53.0052
R6414 gnd.n3523 gnd.n3522 52.4801
R6415 gnd.n5783 gnd.t101 52.3082
R6416 gnd.n5751 gnd.t18 52.3082
R6417 gnd.n5719 gnd.t22 52.3082
R6418 gnd.n5688 gnd.t16 52.3082
R6419 gnd.n5656 gnd.t274 52.3082
R6420 gnd.n5624 gnd.t262 52.3082
R6421 gnd.n5592 gnd.t278 52.3082
R6422 gnd.n5561 gnd.t38 52.3082
R6423 gnd.n5613 gnd.n5581 51.4173
R6424 gnd.n5677 gnd.n5676 50.455
R6425 gnd.n5645 gnd.n5644 50.455
R6426 gnd.n5613 gnd.n5612 50.455
R6427 gnd.n6962 gnd.n83 49.0735
R6428 gnd.n4197 gnd.n1331 45.6325
R6429 gnd.n2833 gnd.n2832 45.6325
R6430 gnd.n4982 gnd.n4981 45.1884
R6431 gnd.n4624 gnd.n4623 45.1884
R6432 gnd.n3539 gnd.n3538 44.3322
R6433 gnd.n2659 gnd.n2658 44.3189
R6434 gnd.n2891 gnd.n2004 42.2793
R6435 gnd.n4994 gnd.n4982 42.2793
R6436 gnd.n4625 gnd.n4624 42.2793
R6437 gnd.n5134 gnd.n5132 42.2793
R6438 gnd.n5886 gnd.n4598 42.2793
R6439 gnd.n6838 gnd.n6834 42.2793
R6440 gnd.n1618 gnd.n1514 42.2793
R6441 gnd.n2866 gnd.n2016 42.2793
R6442 gnd.n1358 gnd.n1357 42.2793
R6443 gnd.n6890 gnd.n158 42.2793
R6444 gnd.n6927 gnd.n6926 42.2793
R6445 gnd.n4538 gnd.n929 42.2793
R6446 gnd.n952 gnd.n951 42.2793
R6447 gnd.n2379 gnd.n2378 42.2793
R6448 gnd.n2584 gnd.n2181 42.2793
R6449 gnd.n3902 gnd.n3901 42.2793
R6450 gnd.n2657 gnd.n2656 41.6274
R6451 gnd.n3533 gnd.n3532 41.6274
R6452 gnd.n2666 gnd.n2665 40.8975
R6453 gnd.n3536 gnd.n3535 40.8975
R6454 gnd.n6119 gnd.n637 38.7261
R6455 gnd.n6113 gnd.n637 38.7261
R6456 gnd.n6113 gnd.n6112 38.7261
R6457 gnd.n6112 gnd.n6111 38.7261
R6458 gnd.n6111 gnd.n644 38.7261
R6459 gnd.n6105 gnd.n644 38.7261
R6460 gnd.n6105 gnd.n6104 38.7261
R6461 gnd.n6104 gnd.n6103 38.7261
R6462 gnd.n6103 gnd.n652 38.7261
R6463 gnd.n6097 gnd.n652 38.7261
R6464 gnd.n6097 gnd.n6096 38.7261
R6465 gnd.n6096 gnd.n6095 38.7261
R6466 gnd.n6095 gnd.n660 38.7261
R6467 gnd.n6089 gnd.n660 38.7261
R6468 gnd.n6089 gnd.n6088 38.7261
R6469 gnd.n6088 gnd.n6087 38.7261
R6470 gnd.n6087 gnd.n668 38.7261
R6471 gnd.n6081 gnd.n668 38.7261
R6472 gnd.n6081 gnd.n6080 38.7261
R6473 gnd.n6080 gnd.n6079 38.7261
R6474 gnd.n6079 gnd.n676 38.7261
R6475 gnd.n6073 gnd.n676 38.7261
R6476 gnd.n6073 gnd.n6072 38.7261
R6477 gnd.n6072 gnd.n6071 38.7261
R6478 gnd.n6071 gnd.n684 38.7261
R6479 gnd.n6065 gnd.n684 38.7261
R6480 gnd.n6065 gnd.n6064 38.7261
R6481 gnd.n6064 gnd.n6063 38.7261
R6482 gnd.n6063 gnd.n692 38.7261
R6483 gnd.n6057 gnd.n692 38.7261
R6484 gnd.n6057 gnd.n6056 38.7261
R6485 gnd.n6056 gnd.n6055 38.7261
R6486 gnd.n6055 gnd.n700 38.7261
R6487 gnd.n6049 gnd.n700 38.7261
R6488 gnd.n6049 gnd.n6048 38.7261
R6489 gnd.n6048 gnd.n6047 38.7261
R6490 gnd.n6047 gnd.n708 38.7261
R6491 gnd.n6041 gnd.n708 38.7261
R6492 gnd.n6041 gnd.n6040 38.7261
R6493 gnd.n6040 gnd.n6039 38.7261
R6494 gnd.n6039 gnd.n716 38.7261
R6495 gnd.n6033 gnd.n716 38.7261
R6496 gnd.n6033 gnd.n6032 38.7261
R6497 gnd.n6032 gnd.n6031 38.7261
R6498 gnd.n6031 gnd.n724 38.7261
R6499 gnd.n6025 gnd.n724 38.7261
R6500 gnd.n6025 gnd.n6024 38.7261
R6501 gnd.n6024 gnd.n6023 38.7261
R6502 gnd.n6023 gnd.n732 38.7261
R6503 gnd.n6017 gnd.n732 38.7261
R6504 gnd.n6017 gnd.n6016 38.7261
R6505 gnd.n6016 gnd.n6015 38.7261
R6506 gnd.n6015 gnd.n740 38.7261
R6507 gnd.n6009 gnd.n740 38.7261
R6508 gnd.n6009 gnd.n6008 38.7261
R6509 gnd.n6008 gnd.n6007 38.7261
R6510 gnd.n6007 gnd.n748 38.7261
R6511 gnd.n6001 gnd.n748 38.7261
R6512 gnd.n6001 gnd.n6000 38.7261
R6513 gnd.n6000 gnd.n5999 38.7261
R6514 gnd.n5999 gnd.n756 38.7261
R6515 gnd.n5993 gnd.n756 38.7261
R6516 gnd.n5993 gnd.n5992 38.7261
R6517 gnd.n5992 gnd.n5991 38.7261
R6518 gnd.n5991 gnd.n764 38.7261
R6519 gnd.n5985 gnd.n764 38.7261
R6520 gnd.n5985 gnd.n5984 38.7261
R6521 gnd.n5984 gnd.n5983 38.7261
R6522 gnd.n5983 gnd.n772 38.7261
R6523 gnd.n5977 gnd.n772 38.7261
R6524 gnd.n5977 gnd.n5976 38.7261
R6525 gnd.n5976 gnd.n5975 38.7261
R6526 gnd.n5975 gnd.n780 38.7261
R6527 gnd.n5969 gnd.n780 38.7261
R6528 gnd.n5969 gnd.n5968 38.7261
R6529 gnd.n5968 gnd.n5967 38.7261
R6530 gnd.n5967 gnd.n788 38.7261
R6531 gnd.n5961 gnd.n788 38.7261
R6532 gnd.n5961 gnd.n5960 38.7261
R6533 gnd.n5960 gnd.n5959 38.7261
R6534 gnd.n5959 gnd.n796 38.7261
R6535 gnd.n5953 gnd.n796 38.7261
R6536 gnd.n5953 gnd.n5952 38.7261
R6537 gnd.n4197 gnd.n1335 36.9518
R6538 gnd.n2833 gnd.n2159 36.9518
R6539 gnd.n2665 gnd.n2664 35.055
R6540 gnd.n2660 gnd.n2659 35.055
R6541 gnd.n3525 gnd.n3524 35.055
R6542 gnd.n3535 gnd.n3521 35.055
R6543 gnd.n3649 gnd.n3647 32.9371
R6544 gnd.n2767 gnd.n2646 32.9371
R6545 gnd.n5044 gnd.n4940 31.8661
R6546 gnd.n5052 gnd.n4940 31.8661
R6547 gnd.n5060 gnd.n4934 31.8661
R6548 gnd.n5060 gnd.n4928 31.8661
R6549 gnd.n5068 gnd.n4928 31.8661
R6550 gnd.n5068 gnd.n4921 31.8661
R6551 gnd.n5076 gnd.n4921 31.8661
R6552 gnd.n5076 gnd.n4922 31.8661
R6553 gnd.n5175 gnd.n4907 31.8661
R6554 gnd.n2435 gnd.n906 31.8661
R6555 gnd.n4487 gnd.n960 31.8661
R6556 gnd.n4487 gnd.n962 31.8661
R6557 gnd.n4481 gnd.n962 31.8661
R6558 gnd.n4481 gnd.n974 31.8661
R6559 gnd.n4475 gnd.n985 31.8661
R6560 gnd.n4469 gnd.n985 31.8661
R6561 gnd.n4463 gnd.n1002 31.8661
R6562 gnd.n2018 gnd.n1162 31.8661
R6563 gnd.n2118 gnd.n1985 31.8661
R6564 gnd.n2900 gnd.n1985 31.8661
R6565 gnd.n2900 gnd.n1978 31.8661
R6566 gnd.n2908 gnd.n1978 31.8661
R6567 gnd.n2908 gnd.n1979 31.8661
R6568 gnd.n4238 gnd.n1272 31.8661
R6569 gnd.n4238 gnd.n4237 31.8661
R6570 gnd.n4237 gnd.n1275 31.8661
R6571 gnd.n4231 gnd.n1275 31.8661
R6572 gnd.n4231 gnd.n4230 31.8661
R6573 gnd.n1362 gnd.n1311 31.8661
R6574 gnd.n6776 gnd.n194 31.8661
R6575 gnd.n6784 gnd.n186 31.8661
R6576 gnd.n6784 gnd.n188 31.8661
R6577 gnd.n6792 gnd.n170 31.8661
R6578 gnd.n6874 gnd.n170 31.8661
R6579 gnd.n6874 gnd.n162 31.8661
R6580 gnd.n6882 gnd.n162 31.8661
R6581 gnd.n6962 gnd.n81 31.8661
R6582 gnd.n1002 gnd.t58 30.9101
R6583 gnd.n6776 gnd.t25 30.9101
R6584 gnd.n2862 gnd.n2118 27.4049
R6585 gnd.n4230 gnd.n4229 27.4049
R6586 gnd.n2461 gnd.n1013 26.7676
R6587 gnd.n4457 gnd.n1016 26.7676
R6588 gnd.n4451 gnd.n1027 26.7676
R6589 gnd.n2326 gnd.n2325 26.7676
R6590 gnd.n4443 gnd.n1038 26.7676
R6591 gnd.n4437 gnd.n1052 26.7676
R6592 gnd.n2496 gnd.n1057 26.7676
R6593 gnd.n2504 gnd.n1066 26.7676
R6594 gnd.n4424 gnd.n1069 26.7676
R6595 gnd.n2512 gnd.n1074 26.7676
R6596 gnd.n4417 gnd.n1077 26.7676
R6597 gnd.n4411 gnd.n1088 26.7676
R6598 gnd.n2528 gnd.n1096 26.7676
R6599 gnd.n2536 gnd.n1106 26.7676
R6600 gnd.n4399 gnd.n1109 26.7676
R6601 gnd.n2544 gnd.n1117 26.7676
R6602 gnd.n4393 gnd.n1120 26.7676
R6603 gnd.n4387 gnd.n1131 26.7676
R6604 gnd.n2560 gnd.n1139 26.7676
R6605 gnd.n4381 gnd.n1142 26.7676
R6606 gnd.n2569 gnd.n1150 26.7676
R6607 gnd.n2577 gnd.n1159 26.7676
R6608 gnd.n4369 gnd.n1162 26.7676
R6609 gnd.n4153 gnd.n1362 26.7676
R6610 gnd.n3974 gnd.n1364 26.7676
R6611 gnd.n3984 gnd.n1495 26.7676
R6612 gnd.n1497 gnd.n1487 26.7676
R6613 gnd.n3995 gnd.n3994 26.7676
R6614 gnd.n4006 gnd.n1478 26.7676
R6615 gnd.n4016 gnd.n1469 26.7676
R6616 gnd.n3942 gnd.n1471 26.7676
R6617 gnd.n4026 gnd.n4025 26.7676
R6618 gnd.n4040 gnd.n1453 26.7676
R6619 gnd.n4051 gnd.n1443 26.7676
R6620 gnd.n1445 gnd.n1437 26.7676
R6621 gnd.n4077 gnd.n1420 26.7676
R6622 gnd.n4082 gnd.n1415 26.7676
R6623 gnd.n4071 gnd.n4070 26.7676
R6624 gnd.n4091 gnd.n1406 26.7676
R6625 gnd.n4100 gnd.n4099 26.7676
R6626 gnd.n4115 gnd.n1397 26.7676
R6627 gnd.n6744 gnd.n229 26.7676
R6628 gnd.n6752 gnd.n221 26.7676
R6629 gnd.n6728 gnd.n223 26.7676
R6630 gnd.n268 gnd.n209 26.7676
R6631 gnd.n6768 gnd.n201 26.7676
R6632 gnd.t55 gnd.n1035 26.4489
R6633 gnd.t86 gnd.n231 26.4489
R6634 gnd.n2004 gnd.n2003 25.7944
R6635 gnd.n5132 gnd.n5131 25.7944
R6636 gnd.n4598 gnd.n4597 25.7944
R6637 gnd.n6834 gnd.n6833 25.7944
R6638 gnd.n1514 gnd.n1513 25.7944
R6639 gnd.n2016 gnd.n2015 25.7944
R6640 gnd.n1335 gnd.n1334 25.7944
R6641 gnd.n1357 gnd.n1356 25.7944
R6642 gnd.n158 gnd.n157 25.7944
R6643 gnd.n6926 gnd.n6925 25.7944
R6644 gnd.n929 gnd.n928 25.7944
R6645 gnd.n951 gnd.n950 25.7944
R6646 gnd.n2378 gnd.n2377 25.7944
R6647 gnd.n2181 gnd.n2180 25.7944
R6648 gnd.n2159 gnd.n2158 25.7944
R6649 gnd.n3901 gnd.n3900 25.7944
R6650 gnd.n5176 gnd.n4896 24.8557
R6651 gnd.n4899 gnd.n4890 24.8557
R6652 gnd.n5197 gnd.n4875 24.8557
R6653 gnd.n5216 gnd.n5215 24.8557
R6654 gnd.n5226 gnd.n4868 24.8557
R6655 gnd.n5239 gnd.n4856 24.8557
R6656 gnd.n5264 gnd.n4840 24.8557
R6657 gnd.n5263 gnd.n4842 24.8557
R6658 gnd.n5286 gnd.n4824 24.8557
R6659 gnd.n5275 gnd.n4816 24.8557
R6660 gnd.n5311 gnd.n5310 24.8557
R6661 gnd.n5321 gnd.n4809 24.8557
R6662 gnd.n5333 gnd.n4801 24.8557
R6663 gnd.n5332 gnd.n4789 24.8557
R6664 gnd.n5351 gnd.n5350 24.8557
R6665 gnd.n5372 gnd.n4770 24.8557
R6666 gnd.n5396 gnd.n5395 24.8557
R6667 gnd.n5407 gnd.n4717 24.8557
R6668 gnd.n5406 gnd.n4719 24.8557
R6669 gnd.n5418 gnd.n4710 24.8557
R6670 gnd.n5435 gnd.n5434 24.8557
R6671 gnd.n4701 gnd.n4690 24.8557
R6672 gnd.n5458 gnd.n4679 24.8557
R6673 gnd.n4681 gnd.n4680 24.8557
R6674 gnd.n5478 gnd.n4673 24.8557
R6675 gnd.n5490 gnd.n5489 24.8557
R6676 gnd.n5501 gnd.n4660 24.8557
R6677 gnd.n5514 gnd.n4650 24.8557
R6678 gnd.n5950 gnd.n806 24.8557
R6679 gnd.n5944 gnd.n5943 24.8557
R6680 gnd.n5543 gnd.n817 24.8557
R6681 gnd.n5936 gnd.n828 24.8557
R6682 gnd.n4634 gnd.n839 24.8557
R6683 gnd.n5930 gnd.n5929 24.8557
R6684 gnd.n5922 gnd.n853 24.8557
R6685 gnd.n2631 gnd.n2630 23.855
R6686 gnd.n3645 gnd.n3644 23.855
R6687 gnd.n2686 gnd.n2685 23.855
R6688 gnd.n3560 gnd.n3559 23.855
R6689 gnd.n5194 gnd.t37 23.2624
R6690 gnd.n1973 gnd.n1972 23.2624
R6691 gnd.n3715 gnd.n3714 23.2624
R6692 gnd.n5952 gnd.n5951 23.2358
R6693 gnd.n5186 gnd.t125 22.6251
R6694 gnd.n3040 gnd.n1942 21.6691
R6695 gnd.n3032 gnd.n1933 21.6691
R6696 gnd.n3017 gnd.n1919 21.6691
R6697 gnd.n3002 gnd.n1904 21.6691
R6698 gnd.n2995 gnd.n1898 21.6691
R6699 gnd.n3213 gnd.n1866 21.6691
R6700 gnd.n3198 gnd.n1851 21.6691
R6701 gnd.n3190 gnd.n1844 21.6691
R6702 gnd.n3183 gnd.n1838 21.6691
R6703 gnd.n3175 gnd.n3141 21.6691
R6704 gnd.n3169 gnd.n3168 21.6691
R6705 gnd.n3384 gnd.n1793 21.6691
R6706 gnd.n3384 gnd.n1796 21.6691
R6707 gnd.n3369 gnd.n1779 21.6691
R6708 gnd.n3361 gnd.n1772 21.6691
R6709 gnd.n3354 gnd.n1764 21.6691
R6710 gnd.n3346 gnd.n1757 21.6691
R6711 gnd.n3340 gnd.n3339 21.6691
R6712 gnd.n3790 gnd.n1718 21.6691
R6713 gnd.n3775 gnd.n1705 21.6691
R6714 gnd.n3767 gnd.n1699 21.6691
R6715 gnd.n3752 gnd.n1685 21.6691
R6716 gnd.n3736 gnd.n1672 21.6691
R6717 gnd.n3722 gnd.n1650 21.6691
R6718 gnd.n5166 gnd.t15 21.3504
R6719 gnd.n2488 gnd.t102 21.3504
R6720 gnd.n6739 gnd.t44 21.3504
R6721 gnd.t32 gnd.n1005 21.0318
R6722 gnd.n6720 gnd.t23 21.0318
R6723 gnd.n2753 gnd.n2669 20.7615
R6724 gnd.n3718 gnd.n3539 20.7615
R6725 gnd.t83 gnd.n804 20.7131
R6726 gnd.n2520 gnd.t105 20.7131
R6727 gnd.t29 gnd.n4059 20.7131
R6728 gnd.t122 gnd.n1964 20.3945
R6729 gnd.n2647 gnd.n1956 20.3945
R6730 gnd.n3048 gnd.n1932 20.3945
R6731 gnd.n2981 gnd.n1880 20.3945
R6732 gnd.n3221 gnd.n1857 20.3945
R6733 gnd.n3281 gnd.n1810 20.3945
R6734 gnd.n3392 gnd.n1785 20.3945
R6735 gnd.n3452 gnd.n1733 20.3945
R6736 gnd.n3798 gnd.n1711 20.3945
R6737 gnd.t81 gnd.n4691 20.0758
R6738 gnd.n4475 gnd.t240 20.0758
R6739 gnd.n2552 gnd.t19 20.0758
R6740 gnd.t143 gnd.t230 20.0758
R6741 gnd.n3946 gnd.t5 20.0758
R6742 gnd.n188 gnd.t263 20.0758
R6743 gnd.n2653 gnd.t214 19.8005
R6744 gnd.n2653 gnd.t130 19.8005
R6745 gnd.n2654 gnd.t123 19.8005
R6746 gnd.n2654 gnd.t151 19.8005
R6747 gnd.n3529 gnd.t172 19.8005
R6748 gnd.n3529 gnd.t137 19.8005
R6749 gnd.n3530 gnd.t188 19.8005
R6750 gnd.n3530 gnd.t116 19.8005
R6751 gnd.n2650 gnd.n2649 19.5087
R6752 gnd.n2663 gnd.n2650 19.5087
R6753 gnd.n2661 gnd.n2652 19.5087
R6754 gnd.n3534 gnd.n3528 19.5087
R6755 gnd.t285 gnd.n4726 19.4385
R6756 gnd.n2910 gnd.n1975 19.3944
R6757 gnd.n2914 gnd.n1975 19.3944
R6758 gnd.n2914 gnd.n1961 19.3944
R6759 gnd.n2928 gnd.n1961 19.3944
R6760 gnd.n2928 gnd.n1958 19.3944
R6761 gnd.n2933 gnd.n1958 19.3944
R6762 gnd.n2933 gnd.n1959 19.3944
R6763 gnd.n1959 gnd.n1930 19.3944
R6764 gnd.n3050 gnd.n1930 19.3944
R6765 gnd.n3050 gnd.n1928 19.3944
R6766 gnd.n3054 gnd.n1928 19.3944
R6767 gnd.n3054 gnd.n1916 19.3944
R6768 gnd.n3066 gnd.n1916 19.3944
R6769 gnd.n3066 gnd.n1914 19.3944
R6770 gnd.n3070 gnd.n1914 19.3944
R6771 gnd.n3070 gnd.n1902 19.3944
R6772 gnd.n3082 gnd.n1902 19.3944
R6773 gnd.n3082 gnd.n1900 19.3944
R6774 gnd.n3086 gnd.n1900 19.3944
R6775 gnd.n3086 gnd.n1886 19.3944
R6776 gnd.n3099 gnd.n1886 19.3944
R6777 gnd.n3099 gnd.n1883 19.3944
R6778 gnd.n3104 gnd.n1883 19.3944
R6779 gnd.n3104 gnd.n1884 19.3944
R6780 gnd.n1884 gnd.n1855 19.3944
R6781 gnd.n3223 gnd.n1855 19.3944
R6782 gnd.n3223 gnd.n1853 19.3944
R6783 gnd.n3227 gnd.n1853 19.3944
R6784 gnd.n3227 gnd.n1842 19.3944
R6785 gnd.n3239 gnd.n1842 19.3944
R6786 gnd.n3239 gnd.n1840 19.3944
R6787 gnd.n3243 gnd.n1840 19.3944
R6788 gnd.n3243 gnd.n1830 19.3944
R6789 gnd.n3255 gnd.n1830 19.3944
R6790 gnd.n3255 gnd.n1828 19.3944
R6791 gnd.n3259 gnd.n1828 19.3944
R6792 gnd.n3259 gnd.n1816 19.3944
R6793 gnd.n3273 gnd.n1816 19.3944
R6794 gnd.n3273 gnd.n1813 19.3944
R6795 gnd.n3278 gnd.n1813 19.3944
R6796 gnd.n3278 gnd.n1814 19.3944
R6797 gnd.n1814 gnd.n1783 19.3944
R6798 gnd.n3394 gnd.n1783 19.3944
R6799 gnd.n3394 gnd.n1781 19.3944
R6800 gnd.n3398 gnd.n1781 19.3944
R6801 gnd.n3398 gnd.n1768 19.3944
R6802 gnd.n3410 gnd.n1768 19.3944
R6803 gnd.n3410 gnd.n1766 19.3944
R6804 gnd.n3414 gnd.n1766 19.3944
R6805 gnd.n3414 gnd.n1754 19.3944
R6806 gnd.n3426 gnd.n1754 19.3944
R6807 gnd.n3426 gnd.n1752 19.3944
R6808 gnd.n3430 gnd.n1752 19.3944
R6809 gnd.n3430 gnd.n1739 19.3944
R6810 gnd.n3444 gnd.n1739 19.3944
R6811 gnd.n3444 gnd.n1736 19.3944
R6812 gnd.n3449 gnd.n1736 19.3944
R6813 gnd.n3449 gnd.n1737 19.3944
R6814 gnd.n1737 gnd.n1709 19.3944
R6815 gnd.n3800 gnd.n1709 19.3944
R6816 gnd.n3800 gnd.n1707 19.3944
R6817 gnd.n3804 gnd.n1707 19.3944
R6818 gnd.n3804 gnd.n1696 19.3944
R6819 gnd.n3816 gnd.n1696 19.3944
R6820 gnd.n3816 gnd.n1694 19.3944
R6821 gnd.n3820 gnd.n1694 19.3944
R6822 gnd.n3820 gnd.n1683 19.3944
R6823 gnd.n3832 gnd.n1683 19.3944
R6824 gnd.n3832 gnd.n1681 19.3944
R6825 gnd.n3836 gnd.n1681 19.3944
R6826 gnd.n3836 gnd.n1669 19.3944
R6827 gnd.n3848 gnd.n1669 19.3944
R6828 gnd.n3848 gnd.n1667 19.3944
R6829 gnd.n3852 gnd.n1667 19.3944
R6830 gnd.n3852 gnd.n1655 19.3944
R6831 gnd.n3864 gnd.n1655 19.3944
R6832 gnd.n3864 gnd.n1652 19.3944
R6833 gnd.n3870 gnd.n1652 19.3944
R6834 gnd.n3870 gnd.n1653 19.3944
R6835 gnd.n1653 gnd.n1642 19.3944
R6836 gnd.n3886 gnd.n1642 19.3944
R6837 gnd.n3887 gnd.n3886 19.3944
R6838 gnd.n2893 gnd.n2000 19.3944
R6839 gnd.n2897 gnd.n2000 19.3944
R6840 gnd.n2897 gnd.n2001 19.3944
R6841 gnd.n2061 gnd.n2058 19.3944
R6842 gnd.n2061 gnd.n2048 19.3944
R6843 gnd.n2070 gnd.n2048 19.3944
R6844 gnd.n2073 gnd.n2070 19.3944
R6845 gnd.n2073 gnd.n2042 19.3944
R6846 gnd.n2082 gnd.n2042 19.3944
R6847 gnd.n2085 gnd.n2082 19.3944
R6848 gnd.n2085 gnd.n2036 19.3944
R6849 gnd.n2094 gnd.n2036 19.3944
R6850 gnd.n2097 gnd.n2094 19.3944
R6851 gnd.n2097 gnd.n2030 19.3944
R6852 gnd.n2107 gnd.n2030 19.3944
R6853 gnd.n2108 gnd.n2107 19.3944
R6854 gnd.n2111 gnd.n2108 19.3944
R6855 gnd.n2111 gnd.n2010 19.3944
R6856 gnd.n2869 gnd.n2010 19.3944
R6857 gnd.n2872 gnd.n2869 19.3944
R6858 gnd.n2872 gnd.n2007 19.3944
R6859 gnd.n2877 gnd.n2007 19.3944
R6860 gnd.n2880 gnd.n2877 19.3944
R6861 gnd.n2883 gnd.n2880 19.3944
R6862 gnd.n2883 gnd.n2005 19.3944
R6863 gnd.n2887 gnd.n2005 19.3944
R6864 gnd.n2890 gnd.n2887 19.3944
R6865 gnd.n5039 gnd.n5038 19.3944
R6866 gnd.n5038 gnd.n4948 19.3944
R6867 gnd.n5033 gnd.n4948 19.3944
R6868 gnd.n5033 gnd.n5032 19.3944
R6869 gnd.n5032 gnd.n4953 19.3944
R6870 gnd.n5027 gnd.n4953 19.3944
R6871 gnd.n5027 gnd.n5026 19.3944
R6872 gnd.n5026 gnd.n5025 19.3944
R6873 gnd.n5025 gnd.n4959 19.3944
R6874 gnd.n5019 gnd.n4959 19.3944
R6875 gnd.n5019 gnd.n5018 19.3944
R6876 gnd.n5018 gnd.n5017 19.3944
R6877 gnd.n5017 gnd.n4965 19.3944
R6878 gnd.n5011 gnd.n4965 19.3944
R6879 gnd.n5011 gnd.n5010 19.3944
R6880 gnd.n5010 gnd.n5009 19.3944
R6881 gnd.n5009 gnd.n4971 19.3944
R6882 gnd.n5003 gnd.n4971 19.3944
R6883 gnd.n5003 gnd.n5002 19.3944
R6884 gnd.n5002 gnd.n5001 19.3944
R6885 gnd.n5001 gnd.n4977 19.3944
R6886 gnd.n4995 gnd.n4977 19.3944
R6887 gnd.n4993 gnd.n4992 19.3944
R6888 gnd.n4992 gnd.n4987 19.3944
R6889 gnd.n4987 gnd.n4985 19.3944
R6890 gnd.n5836 gnd.n5835 19.3944
R6891 gnd.n5835 gnd.n5832 19.3944
R6892 gnd.n5832 gnd.n5831 19.3944
R6893 gnd.n5881 gnd.n5880 19.3944
R6894 gnd.n5880 gnd.n5879 19.3944
R6895 gnd.n5879 gnd.n5876 19.3944
R6896 gnd.n5876 gnd.n5875 19.3944
R6897 gnd.n5875 gnd.n5872 19.3944
R6898 gnd.n5872 gnd.n5871 19.3944
R6899 gnd.n5871 gnd.n5868 19.3944
R6900 gnd.n5868 gnd.n5867 19.3944
R6901 gnd.n5867 gnd.n5864 19.3944
R6902 gnd.n5864 gnd.n5863 19.3944
R6903 gnd.n5863 gnd.n5860 19.3944
R6904 gnd.n5860 gnd.n5859 19.3944
R6905 gnd.n5859 gnd.n5856 19.3944
R6906 gnd.n5856 gnd.n5855 19.3944
R6907 gnd.n5855 gnd.n5852 19.3944
R6908 gnd.n5852 gnd.n5851 19.3944
R6909 gnd.n5851 gnd.n5848 19.3944
R6910 gnd.n5848 gnd.n5847 19.3944
R6911 gnd.n5847 gnd.n5844 19.3944
R6912 gnd.n5844 gnd.n5843 19.3944
R6913 gnd.n5843 gnd.n5840 19.3944
R6914 gnd.n5840 gnd.n5839 19.3944
R6915 gnd.n5179 gnd.n5178 19.3944
R6916 gnd.n5180 gnd.n5179 19.3944
R6917 gnd.n5180 gnd.n4889 19.3944
R6918 gnd.n4889 gnd.n4883 19.3944
R6919 gnd.n5205 gnd.n4883 19.3944
R6920 gnd.n5206 gnd.n5205 19.3944
R6921 gnd.n5206 gnd.n4866 19.3944
R6922 gnd.n4866 gnd.n4864 19.3944
R6923 gnd.n5230 gnd.n4864 19.3944
R6924 gnd.n5233 gnd.n5230 19.3944
R6925 gnd.n5233 gnd.n5232 19.3944
R6926 gnd.n5232 gnd.n4836 19.3944
R6927 gnd.n5271 gnd.n4836 19.3944
R6928 gnd.n5271 gnd.n4834 19.3944
R6929 gnd.n5277 gnd.n4834 19.3944
R6930 gnd.n5278 gnd.n5277 19.3944
R6931 gnd.n5278 gnd.n4804 19.3944
R6932 gnd.n5328 gnd.n4804 19.3944
R6933 gnd.n5329 gnd.n5328 19.3944
R6934 gnd.n5329 gnd.n4797 19.3944
R6935 gnd.n5340 gnd.n4797 19.3944
R6936 gnd.n5341 gnd.n5340 19.3944
R6937 gnd.n5341 gnd.n4780 19.3944
R6938 gnd.n4780 gnd.n4778 19.3944
R6939 gnd.n5365 gnd.n4778 19.3944
R6940 gnd.n5366 gnd.n5365 19.3944
R6941 gnd.n5366 gnd.n4713 19.3944
R6942 gnd.n5413 gnd.n4713 19.3944
R6943 gnd.n5414 gnd.n5413 19.3944
R6944 gnd.n5414 gnd.n4706 19.3944
R6945 gnd.n5425 gnd.n4706 19.3944
R6946 gnd.n5426 gnd.n5425 19.3944
R6947 gnd.n5426 gnd.n4689 19.3944
R6948 gnd.n4689 gnd.n4686 19.3944
R6949 gnd.n5453 gnd.n4686 19.3944
R6950 gnd.n5453 gnd.n4687 19.3944
R6951 gnd.n4687 gnd.n4669 19.3944
R6952 gnd.n5486 gnd.n4669 19.3944
R6953 gnd.n5486 gnd.n5485 19.3944
R6954 gnd.n5485 gnd.n4653 19.3944
R6955 gnd.n5511 gnd.n4653 19.3944
R6956 gnd.n5511 gnd.n4645 19.3944
R6957 gnd.n5524 gnd.n4645 19.3944
R6958 gnd.n5524 gnd.n5523 19.3944
R6959 gnd.n5523 gnd.n4638 19.3944
R6960 gnd.n5546 gnd.n4638 19.3944
R6961 gnd.n5547 gnd.n5546 19.3944
R6962 gnd.n5547 gnd.n4636 19.3944
R6963 gnd.n5809 gnd.n4636 19.3944
R6964 gnd.n5811 gnd.n5809 19.3944
R6965 gnd.n5819 gnd.n5811 19.3944
R6966 gnd.n5819 gnd.n5818 19.3944
R6967 gnd.n5818 gnd.n5817 19.3944
R6968 gnd.n5162 gnd.n5161 19.3944
R6969 gnd.n5161 gnd.n5160 19.3944
R6970 gnd.n5160 gnd.n5159 19.3944
R6971 gnd.n5159 gnd.n5157 19.3944
R6972 gnd.n5157 gnd.n5154 19.3944
R6973 gnd.n5154 gnd.n5153 19.3944
R6974 gnd.n5153 gnd.n5150 19.3944
R6975 gnd.n5150 gnd.n5149 19.3944
R6976 gnd.n5149 gnd.n5146 19.3944
R6977 gnd.n5146 gnd.n5145 19.3944
R6978 gnd.n5145 gnd.n5142 19.3944
R6979 gnd.n5142 gnd.n5141 19.3944
R6980 gnd.n5141 gnd.n5138 19.3944
R6981 gnd.n5138 gnd.n5137 19.3944
R6982 gnd.n5188 gnd.n4894 19.3944
R6983 gnd.n5188 gnd.n4892 19.3944
R6984 gnd.n5192 gnd.n4892 19.3944
R6985 gnd.n5192 gnd.n4873 19.3944
R6986 gnd.n5218 gnd.n4873 19.3944
R6987 gnd.n5218 gnd.n4871 19.3944
R6988 gnd.n5224 gnd.n4871 19.3944
R6989 gnd.n5224 gnd.n5223 19.3944
R6990 gnd.n5223 gnd.n4847 19.3944
R6991 gnd.n5252 gnd.n4847 19.3944
R6992 gnd.n5252 gnd.n4845 19.3944
R6993 gnd.n5261 gnd.n4845 19.3944
R6994 gnd.n5261 gnd.n5260 19.3944
R6995 gnd.n5260 gnd.n5259 19.3944
R6996 gnd.n5259 gnd.n4814 19.3944
R6997 gnd.n5313 gnd.n4814 19.3944
R6998 gnd.n5313 gnd.n4812 19.3944
R6999 gnd.n5319 gnd.n4812 19.3944
R7000 gnd.n5319 gnd.n5318 19.3944
R7001 gnd.n5318 gnd.n4787 19.3944
R7002 gnd.n5353 gnd.n4787 19.3944
R7003 gnd.n5353 gnd.n4785 19.3944
R7004 gnd.n5359 gnd.n4785 19.3944
R7005 gnd.n5359 gnd.n5358 19.3944
R7006 gnd.n5358 gnd.n4724 19.3944
R7007 gnd.n5398 gnd.n4724 19.3944
R7008 gnd.n5398 gnd.n4722 19.3944
R7009 gnd.n5404 gnd.n4722 19.3944
R7010 gnd.n5404 gnd.n5403 19.3944
R7011 gnd.n5403 gnd.n4696 19.3944
R7012 gnd.n5437 gnd.n4696 19.3944
R7013 gnd.n5437 gnd.n4694 19.3944
R7014 gnd.n5446 gnd.n4694 19.3944
R7015 gnd.n5446 gnd.n5445 19.3944
R7016 gnd.n5445 gnd.n5444 19.3944
R7017 gnd.n5444 gnd.n4665 19.3944
R7018 gnd.n5492 gnd.n4665 19.3944
R7019 gnd.n5492 gnd.n4663 19.3944
R7020 gnd.n5499 gnd.n4663 19.3944
R7021 gnd.n5499 gnd.n5498 19.3944
R7022 gnd.n5498 gnd.n809 19.3944
R7023 gnd.n5948 gnd.n809 19.3944
R7024 gnd.n5948 gnd.n5947 19.3944
R7025 gnd.n5947 gnd.n5946 19.3944
R7026 gnd.n5946 gnd.n813 19.3944
R7027 gnd.n831 gnd.n813 19.3944
R7028 gnd.n5934 gnd.n831 19.3944
R7029 gnd.n5934 gnd.n5933 19.3944
R7030 gnd.n5933 gnd.n5932 19.3944
R7031 gnd.n5932 gnd.n837 19.3944
R7032 gnd.n856 gnd.n837 19.3944
R7033 gnd.n5920 gnd.n856 19.3944
R7034 gnd.n5920 gnd.n5919 19.3944
R7035 gnd.n5916 gnd.n861 19.3944
R7036 gnd.n5911 gnd.n861 19.3944
R7037 gnd.n5911 gnd.n5910 19.3944
R7038 gnd.n5910 gnd.n5909 19.3944
R7039 gnd.n5909 gnd.n5906 19.3944
R7040 gnd.n5906 gnd.n5905 19.3944
R7041 gnd.n5905 gnd.n5902 19.3944
R7042 gnd.n5902 gnd.n5901 19.3944
R7043 gnd.n5901 gnd.n5898 19.3944
R7044 gnd.n5898 gnd.n5897 19.3944
R7045 gnd.n5897 gnd.n5894 19.3944
R7046 gnd.n5894 gnd.n5893 19.3944
R7047 gnd.n5893 gnd.n5890 19.3944
R7048 gnd.n5890 gnd.n5889 19.3944
R7049 gnd.n5046 gnd.n4942 19.3944
R7050 gnd.n5050 gnd.n4942 19.3944
R7051 gnd.n5050 gnd.n4932 19.3944
R7052 gnd.n5062 gnd.n4932 19.3944
R7053 gnd.n5062 gnd.n4930 19.3944
R7054 gnd.n5066 gnd.n4930 19.3944
R7055 gnd.n5066 gnd.n4919 19.3944
R7056 gnd.n5078 gnd.n4919 19.3944
R7057 gnd.n5078 gnd.n4917 19.3944
R7058 gnd.n5104 gnd.n4917 19.3944
R7059 gnd.n5104 gnd.n5103 19.3944
R7060 gnd.n5103 gnd.n5102 19.3944
R7061 gnd.n5102 gnd.n5101 19.3944
R7062 gnd.n5101 gnd.n5099 19.3944
R7063 gnd.n5099 gnd.n5098 19.3944
R7064 gnd.n5098 gnd.n5096 19.3944
R7065 gnd.n5096 gnd.n5095 19.3944
R7066 gnd.n5095 gnd.n5093 19.3944
R7067 gnd.n5093 gnd.n5092 19.3944
R7068 gnd.n5092 gnd.n4854 19.3944
R7069 gnd.n5241 gnd.n4854 19.3944
R7070 gnd.n5241 gnd.n4852 19.3944
R7071 gnd.n5247 gnd.n4852 19.3944
R7072 gnd.n5247 gnd.n5246 19.3944
R7073 gnd.n5246 gnd.n4821 19.3944
R7074 gnd.n5288 gnd.n4821 19.3944
R7075 gnd.n5288 gnd.n4819 19.3944
R7076 gnd.n5292 gnd.n4819 19.3944
R7077 gnd.n5306 gnd.n5292 19.3944
R7078 gnd.n5304 gnd.n5303 19.3944
R7079 gnd.n5300 gnd.n5299 19.3944
R7080 gnd.n5296 gnd.n5295 19.3944
R7081 gnd.n5374 gnd.n4768 19.3944
R7082 gnd.n5374 gnd.n4730 19.3944
R7083 gnd.n5393 gnd.n4730 19.3944
R7084 gnd.n5393 gnd.n5392 19.3944
R7085 gnd.n5392 gnd.n5391 19.3944
R7086 gnd.n5391 gnd.n5389 19.3944
R7087 gnd.n5389 gnd.n5388 19.3944
R7088 gnd.n5388 gnd.n5386 19.3944
R7089 gnd.n5386 gnd.n5385 19.3944
R7090 gnd.n5385 gnd.n4677 19.3944
R7091 gnd.n5460 gnd.n4677 19.3944
R7092 gnd.n5460 gnd.n4675 19.3944
R7093 gnd.n5476 gnd.n4675 19.3944
R7094 gnd.n5476 gnd.n5475 19.3944
R7095 gnd.n5475 gnd.n5474 19.3944
R7096 gnd.n5474 gnd.n5473 19.3944
R7097 gnd.n5473 gnd.n5471 19.3944
R7098 gnd.n5471 gnd.n5470 19.3944
R7099 gnd.n5470 gnd.n4643 19.3944
R7100 gnd.n5529 gnd.n4643 19.3944
R7101 gnd.n5529 gnd.n4641 19.3944
R7102 gnd.n5541 gnd.n4641 19.3944
R7103 gnd.n5541 gnd.n5540 19.3944
R7104 gnd.n5540 gnd.n5539 19.3944
R7105 gnd.n5539 gnd.n5536 19.3944
R7106 gnd.n5536 gnd.n4632 19.3944
R7107 gnd.n5824 gnd.n4632 19.3944
R7108 gnd.n5824 gnd.n4630 19.3944
R7109 gnd.n5828 gnd.n4630 19.3944
R7110 gnd.n5042 gnd.n4938 19.3944
R7111 gnd.n5054 gnd.n4938 19.3944
R7112 gnd.n5054 gnd.n4936 19.3944
R7113 gnd.n5058 gnd.n4936 19.3944
R7114 gnd.n5058 gnd.n4926 19.3944
R7115 gnd.n5070 gnd.n4926 19.3944
R7116 gnd.n5070 gnd.n4924 19.3944
R7117 gnd.n5074 gnd.n4924 19.3944
R7118 gnd.n5074 gnd.n4913 19.3944
R7119 gnd.n5168 gnd.n4913 19.3944
R7120 gnd.n5168 gnd.n4910 19.3944
R7121 gnd.n5173 gnd.n4910 19.3944
R7122 gnd.n5173 gnd.n4901 19.3944
R7123 gnd.n5183 gnd.n4901 19.3944
R7124 gnd.n5183 gnd.n4885 19.3944
R7125 gnd.n5200 gnd.n4885 19.3944
R7126 gnd.n5200 gnd.n4881 19.3944
R7127 gnd.n5213 gnd.n4881 19.3944
R7128 gnd.n5213 gnd.n5212 19.3944
R7129 gnd.n5212 gnd.n4860 19.3944
R7130 gnd.n5237 gnd.n4860 19.3944
R7131 gnd.n5237 gnd.n5236 19.3944
R7132 gnd.n5236 gnd.n4838 19.3944
R7133 gnd.n5266 gnd.n4838 19.3944
R7134 gnd.n5266 gnd.n4828 19.3944
R7135 gnd.n5284 gnd.n4828 19.3944
R7136 gnd.n5284 gnd.n5283 19.3944
R7137 gnd.n5283 gnd.n5282 19.3944
R7138 gnd.n5282 gnd.n4806 19.3944
R7139 gnd.n5324 gnd.n4806 19.3944
R7140 gnd.n5324 gnd.n4799 19.3944
R7141 gnd.n5335 gnd.n4799 19.3944
R7142 gnd.n5335 gnd.n4795 19.3944
R7143 gnd.n5348 gnd.n4795 19.3944
R7144 gnd.n5348 gnd.n5347 19.3944
R7145 gnd.n5347 gnd.n4774 19.3944
R7146 gnd.n5370 gnd.n4774 19.3944
R7147 gnd.n5370 gnd.n5369 19.3944
R7148 gnd.n5369 gnd.n4715 19.3944
R7149 gnd.n5409 gnd.n4715 19.3944
R7150 gnd.n5409 gnd.n4708 19.3944
R7151 gnd.n5420 gnd.n4708 19.3944
R7152 gnd.n5420 gnd.n4704 19.3944
R7153 gnd.n5432 gnd.n4704 19.3944
R7154 gnd.n5432 gnd.n5431 19.3944
R7155 gnd.n5431 gnd.n4683 19.3944
R7156 gnd.n5456 gnd.n4683 19.3944
R7157 gnd.n5456 gnd.n4671 19.3944
R7158 gnd.n5480 gnd.n4671 19.3944
R7159 gnd.n5480 gnd.n4655 19.3944
R7160 gnd.n5504 gnd.n4655 19.3944
R7161 gnd.n5505 gnd.n5504 19.3944
R7162 gnd.n5505 gnd.n4649 19.3944
R7163 gnd.n4649 gnd.n4647 19.3944
R7164 gnd.n5518 gnd.n4647 19.3944
R7165 gnd.n5518 gnd.n820 19.3944
R7166 gnd.n5941 gnd.n820 19.3944
R7167 gnd.n5941 gnd.n5940 19.3944
R7168 gnd.n5940 gnd.n5939 19.3944
R7169 gnd.n5939 gnd.n824 19.3944
R7170 gnd.n845 gnd.n824 19.3944
R7171 gnd.n5927 gnd.n845 19.3944
R7172 gnd.n5927 gnd.n5926 19.3944
R7173 gnd.n5926 gnd.n5925 19.3944
R7174 gnd.n5925 gnd.n849 19.3944
R7175 gnd.n3915 gnd.n1503 19.3944
R7176 gnd.n3915 gnd.n1493 19.3944
R7177 gnd.n3986 gnd.n1493 19.3944
R7178 gnd.n3986 gnd.n1490 19.3944
R7179 gnd.n3991 gnd.n1490 19.3944
R7180 gnd.n3991 gnd.n1491 19.3944
R7181 gnd.n1491 gnd.n1467 19.3944
R7182 gnd.n4018 gnd.n1467 19.3944
R7183 gnd.n4018 gnd.n1464 19.3944
R7184 gnd.n4023 gnd.n1464 19.3944
R7185 gnd.n4023 gnd.n1465 19.3944
R7186 gnd.n1465 gnd.n1441 19.3944
R7187 gnd.n4053 gnd.n1441 19.3944
R7188 gnd.n4053 gnd.n1439 19.3944
R7189 gnd.n4057 gnd.n1439 19.3944
R7190 gnd.n4057 gnd.n1413 19.3944
R7191 gnd.n4084 gnd.n1413 19.3944
R7192 gnd.n4084 gnd.n1410 19.3944
R7193 gnd.n4088 gnd.n1410 19.3944
R7194 gnd.n4088 gnd.n1411 19.3944
R7195 gnd.n1411 gnd.n52 19.3944
R7196 gnd.n6994 gnd.n52 19.3944
R7197 gnd.n6994 gnd.n6993 19.3944
R7198 gnd.n6993 gnd.n6992 19.3944
R7199 gnd.n6992 gnd.n57 19.3944
R7200 gnd.n6988 gnd.n57 19.3944
R7201 gnd.n6988 gnd.n6987 19.3944
R7202 gnd.n6987 gnd.n6986 19.3944
R7203 gnd.n6986 gnd.n62 19.3944
R7204 gnd.n6982 gnd.n62 19.3944
R7205 gnd.n6982 gnd.n6981 19.3944
R7206 gnd.n6981 gnd.n6980 19.3944
R7207 gnd.n6980 gnd.n67 19.3944
R7208 gnd.n6976 gnd.n67 19.3944
R7209 gnd.n6976 gnd.n6975 19.3944
R7210 gnd.n6975 gnd.n6974 19.3944
R7211 gnd.n6974 gnd.n72 19.3944
R7212 gnd.n6970 gnd.n72 19.3944
R7213 gnd.n6970 gnd.n6969 19.3944
R7214 gnd.n6969 gnd.n6968 19.3944
R7215 gnd.n6968 gnd.n77 19.3944
R7216 gnd.n6964 gnd.n77 19.3944
R7217 gnd.n6863 gnd.n6862 19.3944
R7218 gnd.n6862 gnd.n6861 19.3944
R7219 gnd.n6861 gnd.n6804 19.3944
R7220 gnd.n6857 gnd.n6804 19.3944
R7221 gnd.n6857 gnd.n6856 19.3944
R7222 gnd.n6856 gnd.n6855 19.3944
R7223 gnd.n6855 gnd.n6812 19.3944
R7224 gnd.n6851 gnd.n6812 19.3944
R7225 gnd.n6851 gnd.n6850 19.3944
R7226 gnd.n6850 gnd.n6849 19.3944
R7227 gnd.n6849 gnd.n6820 19.3944
R7228 gnd.n6845 gnd.n6820 19.3944
R7229 gnd.n6845 gnd.n6844 19.3944
R7230 gnd.n6844 gnd.n6843 19.3944
R7231 gnd.n6843 gnd.n6828 19.3944
R7232 gnd.n6839 gnd.n6828 19.3944
R7233 gnd.n1551 gnd.n1548 19.3944
R7234 gnd.n1554 gnd.n1551 19.3944
R7235 gnd.n1554 gnd.n1542 19.3944
R7236 gnd.n1566 gnd.n1542 19.3944
R7237 gnd.n1567 gnd.n1566 19.3944
R7238 gnd.n1570 gnd.n1567 19.3944
R7239 gnd.n1570 gnd.n1533 19.3944
R7240 gnd.n1583 gnd.n1533 19.3944
R7241 gnd.n1584 gnd.n1583 19.3944
R7242 gnd.n1587 gnd.n1584 19.3944
R7243 gnd.n1587 gnd.n1524 19.3944
R7244 gnd.n1600 gnd.n1524 19.3944
R7245 gnd.n1601 gnd.n1600 19.3944
R7246 gnd.n1604 gnd.n1601 19.3944
R7247 gnd.n1604 gnd.n1515 19.3944
R7248 gnd.n1617 gnd.n1515 19.3944
R7249 gnd.n4151 gnd.n1367 19.3944
R7250 gnd.n4147 gnd.n1367 19.3944
R7251 gnd.n4147 gnd.n4146 19.3944
R7252 gnd.n4146 gnd.n4145 19.3944
R7253 gnd.n4145 gnd.n1373 19.3944
R7254 gnd.n4141 gnd.n1373 19.3944
R7255 gnd.n4141 gnd.n4140 19.3944
R7256 gnd.n4140 gnd.n4139 19.3944
R7257 gnd.n4139 gnd.n1378 19.3944
R7258 gnd.n4135 gnd.n1378 19.3944
R7259 gnd.n4135 gnd.n4134 19.3944
R7260 gnd.n4134 gnd.n4133 19.3944
R7261 gnd.n4133 gnd.n1383 19.3944
R7262 gnd.n4129 gnd.n1383 19.3944
R7263 gnd.n4129 gnd.n4128 19.3944
R7264 gnd.n4128 gnd.n4127 19.3944
R7265 gnd.n4127 gnd.n1388 19.3944
R7266 gnd.n4123 gnd.n1388 19.3944
R7267 gnd.n4123 gnd.n4122 19.3944
R7268 gnd.n4122 gnd.n4121 19.3944
R7269 gnd.n4121 gnd.n1393 19.3944
R7270 gnd.n4117 gnd.n1393 19.3944
R7271 gnd.n4117 gnd.n227 19.3944
R7272 gnd.n6746 gnd.n227 19.3944
R7273 gnd.n6746 gnd.n225 19.3944
R7274 gnd.n6750 gnd.n225 19.3944
R7275 gnd.n6750 gnd.n206 19.3944
R7276 gnd.n6762 gnd.n206 19.3944
R7277 gnd.n6762 gnd.n204 19.3944
R7278 gnd.n6766 gnd.n204 19.3944
R7279 gnd.n6766 gnd.n192 19.3944
R7280 gnd.n6778 gnd.n192 19.3944
R7281 gnd.n6778 gnd.n190 19.3944
R7282 gnd.n6782 gnd.n190 19.3944
R7283 gnd.n6782 gnd.n177 19.3944
R7284 gnd.n6794 gnd.n177 19.3944
R7285 gnd.n6794 gnd.n174 19.3944
R7286 gnd.n6872 gnd.n174 19.3944
R7287 gnd.n6872 gnd.n175 19.3944
R7288 gnd.n6868 gnd.n175 19.3944
R7289 gnd.n6868 gnd.n6867 19.3944
R7290 gnd.n6867 gnd.n6866 19.3944
R7291 gnd.n2051 gnd.n1165 19.3944
R7292 gnd.n2052 gnd.n2051 19.3944
R7293 gnd.n2064 gnd.n2052 19.3944
R7294 gnd.n2067 gnd.n2064 19.3944
R7295 gnd.n2067 gnd.n2046 19.3944
R7296 gnd.n2076 gnd.n2046 19.3944
R7297 gnd.n2079 gnd.n2076 19.3944
R7298 gnd.n2079 gnd.n2038 19.3944
R7299 gnd.n2088 gnd.n2038 19.3944
R7300 gnd.n2091 gnd.n2088 19.3944
R7301 gnd.n2091 gnd.n2034 19.3944
R7302 gnd.n2100 gnd.n2034 19.3944
R7303 gnd.n2103 gnd.n2100 19.3944
R7304 gnd.n2103 gnd.n2027 19.3944
R7305 gnd.n2114 gnd.n2027 19.3944
R7306 gnd.n2114 gnd.n2014 19.3944
R7307 gnd.n6508 gnd.n402 19.3944
R7308 gnd.n6514 gnd.n402 19.3944
R7309 gnd.n6514 gnd.n400 19.3944
R7310 gnd.n6518 gnd.n400 19.3944
R7311 gnd.n6518 gnd.n396 19.3944
R7312 gnd.n6524 gnd.n396 19.3944
R7313 gnd.n6524 gnd.n394 19.3944
R7314 gnd.n6528 gnd.n394 19.3944
R7315 gnd.n6528 gnd.n390 19.3944
R7316 gnd.n6534 gnd.n390 19.3944
R7317 gnd.n6534 gnd.n388 19.3944
R7318 gnd.n6538 gnd.n388 19.3944
R7319 gnd.n6538 gnd.n384 19.3944
R7320 gnd.n6544 gnd.n384 19.3944
R7321 gnd.n6544 gnd.n382 19.3944
R7322 gnd.n6548 gnd.n382 19.3944
R7323 gnd.n6548 gnd.n378 19.3944
R7324 gnd.n6554 gnd.n378 19.3944
R7325 gnd.n6554 gnd.n376 19.3944
R7326 gnd.n6558 gnd.n376 19.3944
R7327 gnd.n6558 gnd.n372 19.3944
R7328 gnd.n6564 gnd.n372 19.3944
R7329 gnd.n6564 gnd.n370 19.3944
R7330 gnd.n6568 gnd.n370 19.3944
R7331 gnd.n6568 gnd.n366 19.3944
R7332 gnd.n6574 gnd.n366 19.3944
R7333 gnd.n6574 gnd.n364 19.3944
R7334 gnd.n6578 gnd.n364 19.3944
R7335 gnd.n6578 gnd.n360 19.3944
R7336 gnd.n6584 gnd.n360 19.3944
R7337 gnd.n6584 gnd.n358 19.3944
R7338 gnd.n6588 gnd.n358 19.3944
R7339 gnd.n6588 gnd.n354 19.3944
R7340 gnd.n6594 gnd.n354 19.3944
R7341 gnd.n6594 gnd.n352 19.3944
R7342 gnd.n6598 gnd.n352 19.3944
R7343 gnd.n6598 gnd.n348 19.3944
R7344 gnd.n6604 gnd.n348 19.3944
R7345 gnd.n6604 gnd.n346 19.3944
R7346 gnd.n6608 gnd.n346 19.3944
R7347 gnd.n6608 gnd.n342 19.3944
R7348 gnd.n6614 gnd.n342 19.3944
R7349 gnd.n6614 gnd.n340 19.3944
R7350 gnd.n6618 gnd.n340 19.3944
R7351 gnd.n6618 gnd.n336 19.3944
R7352 gnd.n6624 gnd.n336 19.3944
R7353 gnd.n6624 gnd.n334 19.3944
R7354 gnd.n6628 gnd.n334 19.3944
R7355 gnd.n6628 gnd.n330 19.3944
R7356 gnd.n6634 gnd.n330 19.3944
R7357 gnd.n6634 gnd.n328 19.3944
R7358 gnd.n6638 gnd.n328 19.3944
R7359 gnd.n6638 gnd.n324 19.3944
R7360 gnd.n6644 gnd.n324 19.3944
R7361 gnd.n6644 gnd.n322 19.3944
R7362 gnd.n6648 gnd.n322 19.3944
R7363 gnd.n6648 gnd.n318 19.3944
R7364 gnd.n6654 gnd.n318 19.3944
R7365 gnd.n6654 gnd.n316 19.3944
R7366 gnd.n6658 gnd.n316 19.3944
R7367 gnd.n6658 gnd.n312 19.3944
R7368 gnd.n6664 gnd.n312 19.3944
R7369 gnd.n6664 gnd.n310 19.3944
R7370 gnd.n6668 gnd.n310 19.3944
R7371 gnd.n6668 gnd.n306 19.3944
R7372 gnd.n6674 gnd.n306 19.3944
R7373 gnd.n6674 gnd.n304 19.3944
R7374 gnd.n6678 gnd.n304 19.3944
R7375 gnd.n6678 gnd.n300 19.3944
R7376 gnd.n6684 gnd.n300 19.3944
R7377 gnd.n6684 gnd.n298 19.3944
R7378 gnd.n6688 gnd.n298 19.3944
R7379 gnd.n6688 gnd.n294 19.3944
R7380 gnd.n6694 gnd.n294 19.3944
R7381 gnd.n6694 gnd.n292 19.3944
R7382 gnd.n6698 gnd.n292 19.3944
R7383 gnd.n6698 gnd.n288 19.3944
R7384 gnd.n6704 gnd.n288 19.3944
R7385 gnd.n6704 gnd.n286 19.3944
R7386 gnd.n6708 gnd.n286 19.3944
R7387 gnd.n6708 gnd.n282 19.3944
R7388 gnd.n6715 gnd.n282 19.3944
R7389 gnd.n6715 gnd.n280 19.3944
R7390 gnd.n6719 gnd.n280 19.3944
R7391 gnd.n6123 gnd.n635 19.3944
R7392 gnd.n6123 gnd.n633 19.3944
R7393 gnd.n6127 gnd.n633 19.3944
R7394 gnd.n6127 gnd.n629 19.3944
R7395 gnd.n6133 gnd.n629 19.3944
R7396 gnd.n6133 gnd.n627 19.3944
R7397 gnd.n6137 gnd.n627 19.3944
R7398 gnd.n6137 gnd.n623 19.3944
R7399 gnd.n6143 gnd.n623 19.3944
R7400 gnd.n6143 gnd.n621 19.3944
R7401 gnd.n6147 gnd.n621 19.3944
R7402 gnd.n6147 gnd.n617 19.3944
R7403 gnd.n6153 gnd.n617 19.3944
R7404 gnd.n6153 gnd.n615 19.3944
R7405 gnd.n6157 gnd.n615 19.3944
R7406 gnd.n6157 gnd.n611 19.3944
R7407 gnd.n6163 gnd.n611 19.3944
R7408 gnd.n6163 gnd.n609 19.3944
R7409 gnd.n6167 gnd.n609 19.3944
R7410 gnd.n6167 gnd.n605 19.3944
R7411 gnd.n6173 gnd.n605 19.3944
R7412 gnd.n6173 gnd.n603 19.3944
R7413 gnd.n6177 gnd.n603 19.3944
R7414 gnd.n6177 gnd.n599 19.3944
R7415 gnd.n6183 gnd.n599 19.3944
R7416 gnd.n6183 gnd.n597 19.3944
R7417 gnd.n6187 gnd.n597 19.3944
R7418 gnd.n6187 gnd.n593 19.3944
R7419 gnd.n6193 gnd.n593 19.3944
R7420 gnd.n6193 gnd.n591 19.3944
R7421 gnd.n6197 gnd.n591 19.3944
R7422 gnd.n6197 gnd.n587 19.3944
R7423 gnd.n6203 gnd.n587 19.3944
R7424 gnd.n6203 gnd.n585 19.3944
R7425 gnd.n6207 gnd.n585 19.3944
R7426 gnd.n6207 gnd.n581 19.3944
R7427 gnd.n6213 gnd.n581 19.3944
R7428 gnd.n6213 gnd.n579 19.3944
R7429 gnd.n6217 gnd.n579 19.3944
R7430 gnd.n6217 gnd.n575 19.3944
R7431 gnd.n6223 gnd.n575 19.3944
R7432 gnd.n6223 gnd.n573 19.3944
R7433 gnd.n6227 gnd.n573 19.3944
R7434 gnd.n6227 gnd.n569 19.3944
R7435 gnd.n6233 gnd.n569 19.3944
R7436 gnd.n6233 gnd.n567 19.3944
R7437 gnd.n6237 gnd.n567 19.3944
R7438 gnd.n6237 gnd.n563 19.3944
R7439 gnd.n6243 gnd.n563 19.3944
R7440 gnd.n6243 gnd.n561 19.3944
R7441 gnd.n6247 gnd.n561 19.3944
R7442 gnd.n6247 gnd.n557 19.3944
R7443 gnd.n6253 gnd.n557 19.3944
R7444 gnd.n6253 gnd.n555 19.3944
R7445 gnd.n6257 gnd.n555 19.3944
R7446 gnd.n6257 gnd.n551 19.3944
R7447 gnd.n6263 gnd.n551 19.3944
R7448 gnd.n6263 gnd.n549 19.3944
R7449 gnd.n6267 gnd.n549 19.3944
R7450 gnd.n6267 gnd.n545 19.3944
R7451 gnd.n6273 gnd.n545 19.3944
R7452 gnd.n6273 gnd.n543 19.3944
R7453 gnd.n6277 gnd.n543 19.3944
R7454 gnd.n6277 gnd.n539 19.3944
R7455 gnd.n6283 gnd.n539 19.3944
R7456 gnd.n6283 gnd.n537 19.3944
R7457 gnd.n6287 gnd.n537 19.3944
R7458 gnd.n6287 gnd.n533 19.3944
R7459 gnd.n6293 gnd.n533 19.3944
R7460 gnd.n6293 gnd.n531 19.3944
R7461 gnd.n6297 gnd.n531 19.3944
R7462 gnd.n6297 gnd.n527 19.3944
R7463 gnd.n6303 gnd.n527 19.3944
R7464 gnd.n6303 gnd.n525 19.3944
R7465 gnd.n6307 gnd.n525 19.3944
R7466 gnd.n6307 gnd.n521 19.3944
R7467 gnd.n6313 gnd.n521 19.3944
R7468 gnd.n6313 gnd.n519 19.3944
R7469 gnd.n6317 gnd.n519 19.3944
R7470 gnd.n6317 gnd.n515 19.3944
R7471 gnd.n6323 gnd.n515 19.3944
R7472 gnd.n6323 gnd.n513 19.3944
R7473 gnd.n6327 gnd.n513 19.3944
R7474 gnd.n6327 gnd.n509 19.3944
R7475 gnd.n6333 gnd.n509 19.3944
R7476 gnd.n6333 gnd.n507 19.3944
R7477 gnd.n6337 gnd.n507 19.3944
R7478 gnd.n6337 gnd.n503 19.3944
R7479 gnd.n6343 gnd.n503 19.3944
R7480 gnd.n6343 gnd.n501 19.3944
R7481 gnd.n6347 gnd.n501 19.3944
R7482 gnd.n6347 gnd.n497 19.3944
R7483 gnd.n6353 gnd.n497 19.3944
R7484 gnd.n6353 gnd.n495 19.3944
R7485 gnd.n6357 gnd.n495 19.3944
R7486 gnd.n6357 gnd.n491 19.3944
R7487 gnd.n6363 gnd.n491 19.3944
R7488 gnd.n6363 gnd.n489 19.3944
R7489 gnd.n6367 gnd.n489 19.3944
R7490 gnd.n6367 gnd.n485 19.3944
R7491 gnd.n6373 gnd.n485 19.3944
R7492 gnd.n6373 gnd.n483 19.3944
R7493 gnd.n6377 gnd.n483 19.3944
R7494 gnd.n6377 gnd.n479 19.3944
R7495 gnd.n6383 gnd.n479 19.3944
R7496 gnd.n6383 gnd.n477 19.3944
R7497 gnd.n6387 gnd.n477 19.3944
R7498 gnd.n6387 gnd.n473 19.3944
R7499 gnd.n6393 gnd.n473 19.3944
R7500 gnd.n6393 gnd.n471 19.3944
R7501 gnd.n6397 gnd.n471 19.3944
R7502 gnd.n6397 gnd.n467 19.3944
R7503 gnd.n6403 gnd.n467 19.3944
R7504 gnd.n6403 gnd.n465 19.3944
R7505 gnd.n6407 gnd.n465 19.3944
R7506 gnd.n6407 gnd.n461 19.3944
R7507 gnd.n6413 gnd.n461 19.3944
R7508 gnd.n6413 gnd.n459 19.3944
R7509 gnd.n6417 gnd.n459 19.3944
R7510 gnd.n6417 gnd.n455 19.3944
R7511 gnd.n6423 gnd.n455 19.3944
R7512 gnd.n6423 gnd.n453 19.3944
R7513 gnd.n6427 gnd.n453 19.3944
R7514 gnd.n6427 gnd.n449 19.3944
R7515 gnd.n6433 gnd.n449 19.3944
R7516 gnd.n6433 gnd.n447 19.3944
R7517 gnd.n6437 gnd.n447 19.3944
R7518 gnd.n6437 gnd.n443 19.3944
R7519 gnd.n6443 gnd.n443 19.3944
R7520 gnd.n6443 gnd.n441 19.3944
R7521 gnd.n6447 gnd.n441 19.3944
R7522 gnd.n6447 gnd.n437 19.3944
R7523 gnd.n6453 gnd.n437 19.3944
R7524 gnd.n6453 gnd.n435 19.3944
R7525 gnd.n6457 gnd.n435 19.3944
R7526 gnd.n6457 gnd.n431 19.3944
R7527 gnd.n6463 gnd.n431 19.3944
R7528 gnd.n6463 gnd.n429 19.3944
R7529 gnd.n6467 gnd.n429 19.3944
R7530 gnd.n6467 gnd.n425 19.3944
R7531 gnd.n6473 gnd.n425 19.3944
R7532 gnd.n6473 gnd.n423 19.3944
R7533 gnd.n6477 gnd.n423 19.3944
R7534 gnd.n6477 gnd.n419 19.3944
R7535 gnd.n6483 gnd.n419 19.3944
R7536 gnd.n6483 gnd.n417 19.3944
R7537 gnd.n6487 gnd.n417 19.3944
R7538 gnd.n6487 gnd.n413 19.3944
R7539 gnd.n6493 gnd.n413 19.3944
R7540 gnd.n6493 gnd.n411 19.3944
R7541 gnd.n6498 gnd.n411 19.3944
R7542 gnd.n6498 gnd.n407 19.3944
R7543 gnd.n6504 gnd.n407 19.3944
R7544 gnd.n6505 gnd.n6504 19.3944
R7545 gnd.n4226 gnd.n4225 19.3944
R7546 gnd.n4225 gnd.n4224 19.3944
R7547 gnd.n4224 gnd.n4223 19.3944
R7548 gnd.n4223 gnd.n4221 19.3944
R7549 gnd.n4221 gnd.n4218 19.3944
R7550 gnd.n4218 gnd.n4217 19.3944
R7551 gnd.n4217 gnd.n4214 19.3944
R7552 gnd.n4214 gnd.n4213 19.3944
R7553 gnd.n4213 gnd.n4210 19.3944
R7554 gnd.n4210 gnd.n4209 19.3944
R7555 gnd.n4209 gnd.n4206 19.3944
R7556 gnd.n4206 gnd.n4205 19.3944
R7557 gnd.n4205 gnd.n4202 19.3944
R7558 gnd.n4202 gnd.n4201 19.3944
R7559 gnd.n4201 gnd.n4198 19.3944
R7560 gnd.n4196 gnd.n4193 19.3944
R7561 gnd.n4193 gnd.n4192 19.3944
R7562 gnd.n4192 gnd.n4189 19.3944
R7563 gnd.n4189 gnd.n4188 19.3944
R7564 gnd.n4188 gnd.n4185 19.3944
R7565 gnd.n4185 gnd.n4184 19.3944
R7566 gnd.n4184 gnd.n4181 19.3944
R7567 gnd.n4181 gnd.n4180 19.3944
R7568 gnd.n4180 gnd.n4177 19.3944
R7569 gnd.n4177 gnd.n4176 19.3944
R7570 gnd.n4176 gnd.n4173 19.3944
R7571 gnd.n4173 gnd.n4172 19.3944
R7572 gnd.n4172 gnd.n4169 19.3944
R7573 gnd.n4169 gnd.n4168 19.3944
R7574 gnd.n4168 gnd.n4165 19.3944
R7575 gnd.n4165 gnd.n4164 19.3944
R7576 gnd.n4164 gnd.n4161 19.3944
R7577 gnd.n4161 gnd.n4160 19.3944
R7578 gnd.n3917 gnd.n1361 19.3944
R7579 gnd.n3954 gnd.n3917 19.3944
R7580 gnd.n3954 gnd.n3953 19.3944
R7581 gnd.n3953 gnd.n3952 19.3944
R7582 gnd.n3952 gnd.n3950 19.3944
R7583 gnd.n3950 gnd.n3949 19.3944
R7584 gnd.n3949 gnd.n3948 19.3944
R7585 gnd.n3948 gnd.n3945 19.3944
R7586 gnd.n3945 gnd.n3944 19.3944
R7587 gnd.n3944 gnd.n3940 19.3944
R7588 gnd.n3940 gnd.n3939 19.3944
R7589 gnd.n3939 gnd.n3938 19.3944
R7590 gnd.n3938 gnd.n3935 19.3944
R7591 gnd.n3935 gnd.n3934 19.3944
R7592 gnd.n3934 gnd.n1422 19.3944
R7593 gnd.n4075 gnd.n1422 19.3944
R7594 gnd.n4075 gnd.n4074 19.3944
R7595 gnd.n4074 gnd.n4073 19.3944
R7596 gnd.n4073 gnd.n1431 19.3944
R7597 gnd.n1431 gnd.n1430 19.3944
R7598 gnd.n1430 gnd.n1428 19.3944
R7599 gnd.n1428 gnd.n234 19.3944
R7600 gnd.n6737 gnd.n234 19.3944
R7601 gnd.n6737 gnd.n6736 19.3944
R7602 gnd.n6736 gnd.n6735 19.3944
R7603 gnd.n6735 gnd.n6731 19.3944
R7604 gnd.n6731 gnd.n6730 19.3944
R7605 gnd.n6730 gnd.n271 19.3944
R7606 gnd.n271 gnd.n270 19.3944
R7607 gnd.n270 gnd.n266 19.3944
R7608 gnd.n266 gnd.n265 19.3944
R7609 gnd.n265 gnd.n263 19.3944
R7610 gnd.n263 gnd.n262 19.3944
R7611 gnd.n262 gnd.n260 19.3944
R7612 gnd.n260 gnd.n259 19.3944
R7613 gnd.n259 gnd.n257 19.3944
R7614 gnd.n257 gnd.n256 19.3944
R7615 gnd.n256 gnd.n254 19.3944
R7616 gnd.n254 gnd.n253 19.3944
R7617 gnd.n253 gnd.n160 19.3944
R7618 gnd.n6885 gnd.n160 19.3944
R7619 gnd.n6886 gnd.n6885 19.3944
R7620 gnd.n6924 gnd.n121 19.3944
R7621 gnd.n6919 gnd.n121 19.3944
R7622 gnd.n6919 gnd.n6918 19.3944
R7623 gnd.n6918 gnd.n6917 19.3944
R7624 gnd.n6917 gnd.n128 19.3944
R7625 gnd.n6912 gnd.n128 19.3944
R7626 gnd.n6912 gnd.n6911 19.3944
R7627 gnd.n6911 gnd.n6910 19.3944
R7628 gnd.n6910 gnd.n135 19.3944
R7629 gnd.n6905 gnd.n135 19.3944
R7630 gnd.n6905 gnd.n6904 19.3944
R7631 gnd.n6904 gnd.n6903 19.3944
R7632 gnd.n6903 gnd.n142 19.3944
R7633 gnd.n6898 gnd.n142 19.3944
R7634 gnd.n6898 gnd.n6897 19.3944
R7635 gnd.n6897 gnd.n6896 19.3944
R7636 gnd.n6896 gnd.n149 19.3944
R7637 gnd.n6891 gnd.n149 19.3944
R7638 gnd.n6957 gnd.n6956 19.3944
R7639 gnd.n6956 gnd.n6955 19.3944
R7640 gnd.n6955 gnd.n92 19.3944
R7641 gnd.n6950 gnd.n92 19.3944
R7642 gnd.n6950 gnd.n6949 19.3944
R7643 gnd.n6949 gnd.n6948 19.3944
R7644 gnd.n6948 gnd.n100 19.3944
R7645 gnd.n6943 gnd.n100 19.3944
R7646 gnd.n6943 gnd.n6942 19.3944
R7647 gnd.n6942 gnd.n6941 19.3944
R7648 gnd.n6941 gnd.n107 19.3944
R7649 gnd.n6936 gnd.n107 19.3944
R7650 gnd.n6936 gnd.n6935 19.3944
R7651 gnd.n6935 gnd.n6934 19.3944
R7652 gnd.n6934 gnd.n114 19.3944
R7653 gnd.n6929 gnd.n114 19.3944
R7654 gnd.n6929 gnd.n6928 19.3944
R7655 gnd.n3976 gnd.n1502 19.3944
R7656 gnd.n3976 gnd.n1500 19.3944
R7657 gnd.n3982 gnd.n1500 19.3944
R7658 gnd.n3982 gnd.n3981 19.3944
R7659 gnd.n3981 gnd.n1476 19.3944
R7660 gnd.n4008 gnd.n1476 19.3944
R7661 gnd.n4008 gnd.n1474 19.3944
R7662 gnd.n4014 gnd.n1474 19.3944
R7663 gnd.n4014 gnd.n4013 19.3944
R7664 gnd.n4013 gnd.n1451 19.3944
R7665 gnd.n4042 gnd.n1451 19.3944
R7666 gnd.n4042 gnd.n1449 19.3944
R7667 gnd.n4049 gnd.n1449 19.3944
R7668 gnd.n4049 gnd.n4048 19.3944
R7669 gnd.n4048 gnd.n4047 19.3944
R7670 gnd.n4047 gnd.n1419 19.3944
R7671 gnd.n4080 gnd.n4079 19.3944
R7672 gnd.n4094 gnd.n4093 19.3944
R7673 gnd.n4097 gnd.n4096 19.3944
R7674 gnd.n6742 gnd.n6741 19.3944
R7675 gnd.n6754 gnd.n219 19.3944
R7676 gnd.n6754 gnd.n211 19.3944
R7677 gnd.n6758 gnd.n211 19.3944
R7678 gnd.n6758 gnd.n199 19.3944
R7679 gnd.n6770 gnd.n199 19.3944
R7680 gnd.n6770 gnd.n197 19.3944
R7681 gnd.n6774 gnd.n197 19.3944
R7682 gnd.n6774 gnd.n183 19.3944
R7683 gnd.n6786 gnd.n183 19.3944
R7684 gnd.n6786 gnd.n181 19.3944
R7685 gnd.n6790 gnd.n181 19.3944
R7686 gnd.n6790 gnd.n167 19.3944
R7687 gnd.n6876 gnd.n167 19.3944
R7688 gnd.n6876 gnd.n165 19.3944
R7689 gnd.n6880 gnd.n165 19.3944
R7690 gnd.n6880 gnd.n87 19.3944
R7691 gnd.n6960 gnd.n87 19.3944
R7692 gnd.n2314 gnd.n2308 19.3944
R7693 gnd.n2318 gnd.n2308 19.3944
R7694 gnd.n2318 gnd.n2228 19.3944
R7695 gnd.n2323 gnd.n2228 19.3944
R7696 gnd.n2305 gnd.n2229 19.3944
R7697 gnd.n2301 gnd.n2234 19.3944
R7698 gnd.n2299 gnd.n2298 19.3944
R7699 gnd.n2295 gnd.n2294 19.3944
R7700 gnd.n2291 gnd.n2290 19.3944
R7701 gnd.n2290 gnd.n2289 19.3944
R7702 gnd.n2289 gnd.n2237 19.3944
R7703 gnd.n2285 gnd.n2237 19.3944
R7704 gnd.n2285 gnd.n2284 19.3944
R7705 gnd.n2284 gnd.n2283 19.3944
R7706 gnd.n2283 gnd.n2243 19.3944
R7707 gnd.n2279 gnd.n2243 19.3944
R7708 gnd.n2279 gnd.n2278 19.3944
R7709 gnd.n2278 gnd.n2277 19.3944
R7710 gnd.n2277 gnd.n2249 19.3944
R7711 gnd.n2273 gnd.n2249 19.3944
R7712 gnd.n2273 gnd.n2272 19.3944
R7713 gnd.n2272 gnd.n2271 19.3944
R7714 gnd.n2271 gnd.n2255 19.3944
R7715 gnd.n2267 gnd.n2255 19.3944
R7716 gnd.n2267 gnd.n2266 19.3944
R7717 gnd.n2266 gnd.n2265 19.3944
R7718 gnd.n2265 gnd.n2262 19.3944
R7719 gnd.n2262 gnd.n1983 19.3944
R7720 gnd.n2902 gnd.n1983 19.3944
R7721 gnd.n2902 gnd.n1981 19.3944
R7722 gnd.n2906 gnd.n1981 19.3944
R7723 gnd.n2906 gnd.n1969 19.3944
R7724 gnd.n2918 gnd.n1969 19.3944
R7725 gnd.n2918 gnd.n1967 19.3944
R7726 gnd.n2924 gnd.n1967 19.3944
R7727 gnd.n2924 gnd.n2923 19.3944
R7728 gnd.n2923 gnd.n1937 19.3944
R7729 gnd.n3042 gnd.n1937 19.3944
R7730 gnd.n3042 gnd.n1935 19.3944
R7731 gnd.n3046 gnd.n1935 19.3944
R7732 gnd.n3046 gnd.n1923 19.3944
R7733 gnd.n3058 gnd.n1923 19.3944
R7734 gnd.n3058 gnd.n1921 19.3944
R7735 gnd.n3062 gnd.n1921 19.3944
R7736 gnd.n3062 gnd.n1908 19.3944
R7737 gnd.n3074 gnd.n1908 19.3944
R7738 gnd.n3074 gnd.n1906 19.3944
R7739 gnd.n3078 gnd.n1906 19.3944
R7740 gnd.n3078 gnd.n1894 19.3944
R7741 gnd.n3089 gnd.n1894 19.3944
R7742 gnd.n3089 gnd.n1892 19.3944
R7743 gnd.n3095 gnd.n1892 19.3944
R7744 gnd.n3095 gnd.n3094 19.3944
R7745 gnd.n3094 gnd.n1862 19.3944
R7746 gnd.n3215 gnd.n1862 19.3944
R7747 gnd.n3215 gnd.n1860 19.3944
R7748 gnd.n3219 gnd.n1860 19.3944
R7749 gnd.n3219 gnd.n1848 19.3944
R7750 gnd.n3231 gnd.n1848 19.3944
R7751 gnd.n3231 gnd.n1846 19.3944
R7752 gnd.n3235 gnd.n1846 19.3944
R7753 gnd.n3235 gnd.n1835 19.3944
R7754 gnd.n3247 gnd.n1835 19.3944
R7755 gnd.n3247 gnd.n1833 19.3944
R7756 gnd.n3251 gnd.n1833 19.3944
R7757 gnd.n3251 gnd.n1824 19.3944
R7758 gnd.n3263 gnd.n1824 19.3944
R7759 gnd.n3263 gnd.n1822 19.3944
R7760 gnd.n3269 gnd.n1822 19.3944
R7761 gnd.n3269 gnd.n3268 19.3944
R7762 gnd.n3268 gnd.n1791 19.3944
R7763 gnd.n3386 gnd.n1791 19.3944
R7764 gnd.n3386 gnd.n1789 19.3944
R7765 gnd.n3390 gnd.n1789 19.3944
R7766 gnd.n3390 gnd.n1776 19.3944
R7767 gnd.n3402 gnd.n1776 19.3944
R7768 gnd.n3402 gnd.n1774 19.3944
R7769 gnd.n3406 gnd.n1774 19.3944
R7770 gnd.n3406 gnd.n1761 19.3944
R7771 gnd.n3418 gnd.n1761 19.3944
R7772 gnd.n3418 gnd.n1759 19.3944
R7773 gnd.n3422 gnd.n1759 19.3944
R7774 gnd.n3422 gnd.n1748 19.3944
R7775 gnd.n3434 gnd.n1748 19.3944
R7776 gnd.n3434 gnd.n1746 19.3944
R7777 gnd.n3440 gnd.n1746 19.3944
R7778 gnd.n3440 gnd.n3439 19.3944
R7779 gnd.n3439 gnd.n1716 19.3944
R7780 gnd.n3792 gnd.n1716 19.3944
R7781 gnd.n3792 gnd.n1714 19.3944
R7782 gnd.n3796 gnd.n1714 19.3944
R7783 gnd.n3796 gnd.n1703 19.3944
R7784 gnd.n3808 gnd.n1703 19.3944
R7785 gnd.n3808 gnd.n1701 19.3944
R7786 gnd.n3812 gnd.n1701 19.3944
R7787 gnd.n3812 gnd.n1689 19.3944
R7788 gnd.n3824 gnd.n1689 19.3944
R7789 gnd.n3824 gnd.n1687 19.3944
R7790 gnd.n3828 gnd.n1687 19.3944
R7791 gnd.n3828 gnd.n1676 19.3944
R7792 gnd.n3840 gnd.n1676 19.3944
R7793 gnd.n3840 gnd.n1674 19.3944
R7794 gnd.n3844 gnd.n1674 19.3944
R7795 gnd.n3844 gnd.n1662 19.3944
R7796 gnd.n3856 gnd.n1662 19.3944
R7797 gnd.n3856 gnd.n1660 19.3944
R7798 gnd.n3860 gnd.n1660 19.3944
R7799 gnd.n3860 gnd.n1648 19.3944
R7800 gnd.n3874 gnd.n1648 19.3944
R7801 gnd.n3874 gnd.n1646 19.3944
R7802 gnd.n3881 gnd.n1646 19.3944
R7803 gnd.n3881 gnd.n3880 19.3944
R7804 gnd.n3880 gnd.n1277 19.3944
R7805 gnd.n4235 gnd.n1277 19.3944
R7806 gnd.n4235 gnd.n4234 19.3944
R7807 gnd.n4234 gnd.n4233 19.3944
R7808 gnd.n4233 gnd.n1281 19.3944
R7809 gnd.n3962 gnd.n1281 19.3944
R7810 gnd.n3965 gnd.n3962 19.3944
R7811 gnd.n3965 gnd.n3959 19.3944
R7812 gnd.n3971 gnd.n3959 19.3944
R7813 gnd.n3971 gnd.n3970 19.3944
R7814 gnd.n3970 gnd.n1485 19.3944
R7815 gnd.n3997 gnd.n1485 19.3944
R7816 gnd.n3997 gnd.n1483 19.3944
R7817 gnd.n4003 gnd.n1483 19.3944
R7818 gnd.n4003 gnd.n4002 19.3944
R7819 gnd.n4002 gnd.n1460 19.3944
R7820 gnd.n4028 gnd.n1460 19.3944
R7821 gnd.n4028 gnd.n1458 19.3944
R7822 gnd.n4037 gnd.n1458 19.3944
R7823 gnd.n4037 gnd.n4036 19.3944
R7824 gnd.n4036 gnd.n4035 19.3944
R7825 gnd.n4035 gnd.n1434 19.3944
R7826 gnd.n4063 gnd.n1434 19.3944
R7827 gnd.n4064 gnd.n4063 19.3944
R7828 gnd.n4068 gnd.n4067 19.3944
R7829 gnd.n4102 gnd.n1400 19.3944
R7830 gnd.n4112 gnd.n4104 19.3944
R7831 gnd.n4110 gnd.n4109 19.3944
R7832 gnd.n4106 gnd.n274 19.3944
R7833 gnd.n6725 gnd.n274 19.3944
R7834 gnd.n6725 gnd.n6724 19.3944
R7835 gnd.n6724 gnd.n6723 19.3944
R7836 gnd.n4571 gnd.n4570 19.3944
R7837 gnd.n4570 gnd.n4569 19.3944
R7838 gnd.n4569 gnd.n4568 19.3944
R7839 gnd.n4568 gnd.n4566 19.3944
R7840 gnd.n4566 gnd.n4563 19.3944
R7841 gnd.n4563 gnd.n4562 19.3944
R7842 gnd.n4562 gnd.n4559 19.3944
R7843 gnd.n4559 gnd.n4558 19.3944
R7844 gnd.n4558 gnd.n4555 19.3944
R7845 gnd.n4555 gnd.n4554 19.3944
R7846 gnd.n4554 gnd.n4551 19.3944
R7847 gnd.n4551 gnd.n4550 19.3944
R7848 gnd.n4550 gnd.n4547 19.3944
R7849 gnd.n4547 gnd.n4546 19.3944
R7850 gnd.n4546 gnd.n4543 19.3944
R7851 gnd.n4543 gnd.n4542 19.3944
R7852 gnd.n4542 gnd.n4539 19.3944
R7853 gnd.n4537 gnd.n4534 19.3944
R7854 gnd.n4534 gnd.n4533 19.3944
R7855 gnd.n4533 gnd.n4530 19.3944
R7856 gnd.n4530 gnd.n4529 19.3944
R7857 gnd.n4529 gnd.n4526 19.3944
R7858 gnd.n4526 gnd.n4525 19.3944
R7859 gnd.n4525 gnd.n4522 19.3944
R7860 gnd.n4522 gnd.n4521 19.3944
R7861 gnd.n4521 gnd.n4518 19.3944
R7862 gnd.n4518 gnd.n4517 19.3944
R7863 gnd.n4517 gnd.n4514 19.3944
R7864 gnd.n4514 gnd.n4513 19.3944
R7865 gnd.n4513 gnd.n4510 19.3944
R7866 gnd.n4510 gnd.n4509 19.3944
R7867 gnd.n4509 gnd.n4506 19.3944
R7868 gnd.n4506 gnd.n4505 19.3944
R7869 gnd.n4505 gnd.n4502 19.3944
R7870 gnd.n4502 gnd.n4501 19.3944
R7871 gnd.n2427 gnd.n2359 19.3944
R7872 gnd.n2427 gnd.n2360 19.3944
R7873 gnd.n2423 gnd.n2360 19.3944
R7874 gnd.n2423 gnd.n977 19.3944
R7875 gnd.n4479 gnd.n977 19.3944
R7876 gnd.n4479 gnd.n4478 19.3944
R7877 gnd.n4478 gnd.n4477 19.3944
R7878 gnd.n4477 gnd.n981 19.3944
R7879 gnd.n4467 gnd.n981 19.3944
R7880 gnd.n4467 gnd.n4466 19.3944
R7881 gnd.n4466 gnd.n4465 19.3944
R7882 gnd.n4465 gnd.n1000 19.3944
R7883 gnd.n4455 gnd.n1000 19.3944
R7884 gnd.n4455 gnd.n4454 19.3944
R7885 gnd.n4454 gnd.n4453 19.3944
R7886 gnd.n4453 gnd.n1022 19.3944
R7887 gnd.n1041 gnd.n1022 19.3944
R7888 gnd.n4441 gnd.n1041 19.3944
R7889 gnd.n4441 gnd.n4440 19.3944
R7890 gnd.n4440 gnd.n4439 19.3944
R7891 gnd.n4439 gnd.n1047 19.3944
R7892 gnd.n4428 gnd.n1047 19.3944
R7893 gnd.n4428 gnd.n4427 19.3944
R7894 gnd.n4427 gnd.n4426 19.3944
R7895 gnd.n4426 gnd.n1064 19.3944
R7896 gnd.n4415 gnd.n1064 19.3944
R7897 gnd.n4415 gnd.n4414 19.3944
R7898 gnd.n4414 gnd.n4413 19.3944
R7899 gnd.n4413 gnd.n1083 19.3944
R7900 gnd.n4403 gnd.n1083 19.3944
R7901 gnd.n4403 gnd.n4402 19.3944
R7902 gnd.n4402 gnd.n4401 19.3944
R7903 gnd.n4401 gnd.n1104 19.3944
R7904 gnd.n4391 gnd.n1104 19.3944
R7905 gnd.n4391 gnd.n4390 19.3944
R7906 gnd.n4390 gnd.n4389 19.3944
R7907 gnd.n4389 gnd.n1126 19.3944
R7908 gnd.n4379 gnd.n1126 19.3944
R7909 gnd.n4379 gnd.n4378 19.3944
R7910 gnd.n4378 gnd.n4377 19.3944
R7911 gnd.n4377 gnd.n1148 19.3944
R7912 gnd.n4367 gnd.n1148 19.3944
R7913 gnd.n2419 gnd.n2417 19.3944
R7914 gnd.n2417 gnd.n2414 19.3944
R7915 gnd.n2414 gnd.n2413 19.3944
R7916 gnd.n2413 gnd.n2410 19.3944
R7917 gnd.n2410 gnd.n2409 19.3944
R7918 gnd.n2409 gnd.n2406 19.3944
R7919 gnd.n2406 gnd.n2405 19.3944
R7920 gnd.n2405 gnd.n2402 19.3944
R7921 gnd.n2402 gnd.n2401 19.3944
R7922 gnd.n2401 gnd.n2398 19.3944
R7923 gnd.n2398 gnd.n2397 19.3944
R7924 gnd.n2397 gnd.n2394 19.3944
R7925 gnd.n2394 gnd.n2393 19.3944
R7926 gnd.n2393 gnd.n2390 19.3944
R7927 gnd.n2390 gnd.n2389 19.3944
R7928 gnd.n2389 gnd.n2386 19.3944
R7929 gnd.n2380 gnd.n2355 19.3944
R7930 gnd.n2438 gnd.n2355 19.3944
R7931 gnd.n2438 gnd.n2353 19.3944
R7932 gnd.n2443 gnd.n2353 19.3944
R7933 gnd.n2444 gnd.n2443 19.3944
R7934 gnd.n2446 gnd.n2444 19.3944
R7935 gnd.n2446 gnd.n2351 19.3944
R7936 gnd.n2451 gnd.n2351 19.3944
R7937 gnd.n2452 gnd.n2451 19.3944
R7938 gnd.n2454 gnd.n2452 19.3944
R7939 gnd.n2454 gnd.n2349 19.3944
R7940 gnd.n2459 gnd.n2349 19.3944
R7941 gnd.n2459 gnd.n2330 19.3944
R7942 gnd.n2473 gnd.n2330 19.3944
R7943 gnd.n2474 gnd.n2473 19.3944
R7944 gnd.n2474 gnd.n2328 19.3944
R7945 gnd.n2478 gnd.n2328 19.3944
R7946 gnd.n2478 gnd.n2221 19.3944
R7947 gnd.n2490 gnd.n2221 19.3944
R7948 gnd.n2490 gnd.n2219 19.3944
R7949 gnd.n2494 gnd.n2219 19.3944
R7950 gnd.n2494 gnd.n2213 19.3944
R7951 gnd.n2506 gnd.n2213 19.3944
R7952 gnd.n2506 gnd.n2211 19.3944
R7953 gnd.n2510 gnd.n2211 19.3944
R7954 gnd.n2510 gnd.n2207 19.3944
R7955 gnd.n2522 gnd.n2207 19.3944
R7956 gnd.n2522 gnd.n2205 19.3944
R7957 gnd.n2526 gnd.n2205 19.3944
R7958 gnd.n2526 gnd.n2200 19.3944
R7959 gnd.n2538 gnd.n2200 19.3944
R7960 gnd.n2538 gnd.n2198 19.3944
R7961 gnd.n2542 gnd.n2198 19.3944
R7962 gnd.n2542 gnd.n2194 19.3944
R7963 gnd.n2554 gnd.n2194 19.3944
R7964 gnd.n2554 gnd.n2192 19.3944
R7965 gnd.n2558 gnd.n2192 19.3944
R7966 gnd.n2558 gnd.n2188 19.3944
R7967 gnd.n2571 gnd.n2188 19.3944
R7968 gnd.n2571 gnd.n2185 19.3944
R7969 gnd.n2575 gnd.n2185 19.3944
R7970 gnd.n2575 gnd.n2186 19.3944
R7971 gnd.n4494 gnd.n4493 19.3944
R7972 gnd.n4493 gnd.n955 19.3944
R7973 gnd.n4489 gnd.n955 19.3944
R7974 gnd.n4489 gnd.n957 19.3944
R7975 gnd.n2335 gnd.n957 19.3944
R7976 gnd.n2339 gnd.n2335 19.3944
R7977 gnd.n2340 gnd.n2339 19.3944
R7978 gnd.n2342 gnd.n2340 19.3944
R7979 gnd.n2342 gnd.n2333 19.3944
R7980 gnd.n2347 gnd.n2333 19.3944
R7981 gnd.n2348 gnd.n2347 19.3944
R7982 gnd.n2463 gnd.n2348 19.3944
R7983 gnd.n2463 gnd.n2331 19.3944
R7984 gnd.n2469 gnd.n2331 19.3944
R7985 gnd.n2469 gnd.n2468 19.3944
R7986 gnd.n2468 gnd.n2224 19.3944
R7987 gnd.n2482 gnd.n2224 19.3944
R7988 gnd.n2482 gnd.n2222 19.3944
R7989 gnd.n2486 gnd.n2222 19.3944
R7990 gnd.n2486 gnd.n2218 19.3944
R7991 gnd.n2498 gnd.n2218 19.3944
R7992 gnd.n2498 gnd.n2215 19.3944
R7993 gnd.n2502 gnd.n2215 19.3944
R7994 gnd.n2502 gnd.n2210 19.3944
R7995 gnd.n2514 gnd.n2210 19.3944
R7996 gnd.n2514 gnd.n2208 19.3944
R7997 gnd.n2518 gnd.n2208 19.3944
R7998 gnd.n2518 gnd.n2204 19.3944
R7999 gnd.n2530 gnd.n2204 19.3944
R8000 gnd.n2530 gnd.n2202 19.3944
R8001 gnd.n2534 gnd.n2202 19.3944
R8002 gnd.n2534 gnd.n2197 19.3944
R8003 gnd.n2546 gnd.n2197 19.3944
R8004 gnd.n2546 gnd.n2195 19.3944
R8005 gnd.n2550 gnd.n2195 19.3944
R8006 gnd.n2550 gnd.n2191 19.3944
R8007 gnd.n2562 gnd.n2191 19.3944
R8008 gnd.n2562 gnd.n2189 19.3944
R8009 gnd.n2567 gnd.n2189 19.3944
R8010 gnd.n2567 gnd.n2183 19.3944
R8011 gnd.n2579 gnd.n2183 19.3944
R8012 gnd.n2580 gnd.n2579 19.3944
R8013 gnd.n2622 gnd.n2157 19.3944
R8014 gnd.n2622 gnd.n2619 19.3944
R8015 gnd.n2619 gnd.n2616 19.3944
R8016 gnd.n2616 gnd.n2615 19.3944
R8017 gnd.n2615 gnd.n2612 19.3944
R8018 gnd.n2612 gnd.n2611 19.3944
R8019 gnd.n2611 gnd.n2608 19.3944
R8020 gnd.n2608 gnd.n2607 19.3944
R8021 gnd.n2607 gnd.n2604 19.3944
R8022 gnd.n2604 gnd.n2603 19.3944
R8023 gnd.n2603 gnd.n2600 19.3944
R8024 gnd.n2600 gnd.n2599 19.3944
R8025 gnd.n2599 gnd.n2596 19.3944
R8026 gnd.n2596 gnd.n2595 19.3944
R8027 gnd.n2595 gnd.n2592 19.3944
R8028 gnd.n2592 gnd.n2591 19.3944
R8029 gnd.n2591 gnd.n2588 19.3944
R8030 gnd.n2588 gnd.n2587 19.3944
R8031 gnd.n2140 gnd.n2139 19.3944
R8032 gnd.n2859 gnd.n2139 19.3944
R8033 gnd.n2859 gnd.n2858 19.3944
R8034 gnd.n2858 gnd.n2857 19.3944
R8035 gnd.n2857 gnd.n2854 19.3944
R8036 gnd.n2854 gnd.n2853 19.3944
R8037 gnd.n2853 gnd.n2850 19.3944
R8038 gnd.n2850 gnd.n2849 19.3944
R8039 gnd.n2849 gnd.n2846 19.3944
R8040 gnd.n2846 gnd.n2845 19.3944
R8041 gnd.n2845 gnd.n2842 19.3944
R8042 gnd.n2842 gnd.n2841 19.3944
R8043 gnd.n2841 gnd.n2838 19.3944
R8044 gnd.n2838 gnd.n2837 19.3944
R8045 gnd.n2837 gnd.n2834 19.3944
R8046 gnd.n2433 gnd.n2429 19.3944
R8047 gnd.n2433 gnd.n966 19.3944
R8048 gnd.n4485 gnd.n966 19.3944
R8049 gnd.n4485 gnd.n4484 19.3944
R8050 gnd.n4484 gnd.n4483 19.3944
R8051 gnd.n4483 gnd.n970 19.3944
R8052 gnd.n4473 gnd.n970 19.3944
R8053 gnd.n4473 gnd.n4472 19.3944
R8054 gnd.n4472 gnd.n4471 19.3944
R8055 gnd.n4471 gnd.n991 19.3944
R8056 gnd.n4461 gnd.n991 19.3944
R8057 gnd.n4461 gnd.n4460 19.3944
R8058 gnd.n4460 gnd.n4459 19.3944
R8059 gnd.n4459 gnd.n1011 19.3944
R8060 gnd.n4449 gnd.n1011 19.3944
R8061 gnd.n4449 gnd.n4448 19.3944
R8062 gnd.n4446 gnd.n4445 19.3944
R8063 gnd.n4435 gnd.n1054 19.3944
R8064 gnd.n4433 gnd.n4432 19.3944
R8065 gnd.n4422 gnd.n1071 19.3944
R8066 gnd.n4420 gnd.n4419 19.3944
R8067 gnd.n4419 gnd.n1072 19.3944
R8068 gnd.n4409 gnd.n1072 19.3944
R8069 gnd.n4409 gnd.n4408 19.3944
R8070 gnd.n4408 gnd.n4407 19.3944
R8071 gnd.n4407 gnd.n1094 19.3944
R8072 gnd.n4397 gnd.n1094 19.3944
R8073 gnd.n4397 gnd.n4396 19.3944
R8074 gnd.n4396 gnd.n4395 19.3944
R8075 gnd.n4395 gnd.n1115 19.3944
R8076 gnd.n4385 gnd.n1115 19.3944
R8077 gnd.n4385 gnd.n4384 19.3944
R8078 gnd.n4384 gnd.n4383 19.3944
R8079 gnd.n4383 gnd.n1137 19.3944
R8080 gnd.n4373 gnd.n1137 19.3944
R8081 gnd.n4373 gnd.n4372 19.3944
R8082 gnd.n4372 gnd.n4371 19.3944
R8083 gnd.n6117 gnd.n6116 19.3944
R8084 gnd.n6116 gnd.n6115 19.3944
R8085 gnd.n6115 gnd.n642 19.3944
R8086 gnd.n6109 gnd.n642 19.3944
R8087 gnd.n6109 gnd.n6108 19.3944
R8088 gnd.n6108 gnd.n6107 19.3944
R8089 gnd.n6107 gnd.n650 19.3944
R8090 gnd.n6101 gnd.n650 19.3944
R8091 gnd.n6101 gnd.n6100 19.3944
R8092 gnd.n6100 gnd.n6099 19.3944
R8093 gnd.n6099 gnd.n658 19.3944
R8094 gnd.n6093 gnd.n658 19.3944
R8095 gnd.n6093 gnd.n6092 19.3944
R8096 gnd.n6092 gnd.n6091 19.3944
R8097 gnd.n6091 gnd.n666 19.3944
R8098 gnd.n6085 gnd.n666 19.3944
R8099 gnd.n6085 gnd.n6084 19.3944
R8100 gnd.n6084 gnd.n6083 19.3944
R8101 gnd.n6083 gnd.n674 19.3944
R8102 gnd.n6077 gnd.n674 19.3944
R8103 gnd.n6077 gnd.n6076 19.3944
R8104 gnd.n6076 gnd.n6075 19.3944
R8105 gnd.n6075 gnd.n682 19.3944
R8106 gnd.n6069 gnd.n682 19.3944
R8107 gnd.n6069 gnd.n6068 19.3944
R8108 gnd.n6068 gnd.n6067 19.3944
R8109 gnd.n6067 gnd.n690 19.3944
R8110 gnd.n6061 gnd.n690 19.3944
R8111 gnd.n6061 gnd.n6060 19.3944
R8112 gnd.n6060 gnd.n6059 19.3944
R8113 gnd.n6059 gnd.n698 19.3944
R8114 gnd.n6053 gnd.n698 19.3944
R8115 gnd.n6053 gnd.n6052 19.3944
R8116 gnd.n6052 gnd.n6051 19.3944
R8117 gnd.n6051 gnd.n706 19.3944
R8118 gnd.n6045 gnd.n706 19.3944
R8119 gnd.n6045 gnd.n6044 19.3944
R8120 gnd.n6044 gnd.n6043 19.3944
R8121 gnd.n6043 gnd.n714 19.3944
R8122 gnd.n6037 gnd.n714 19.3944
R8123 gnd.n6037 gnd.n6036 19.3944
R8124 gnd.n6036 gnd.n6035 19.3944
R8125 gnd.n6035 gnd.n722 19.3944
R8126 gnd.n6029 gnd.n722 19.3944
R8127 gnd.n6029 gnd.n6028 19.3944
R8128 gnd.n6028 gnd.n6027 19.3944
R8129 gnd.n6027 gnd.n730 19.3944
R8130 gnd.n6021 gnd.n730 19.3944
R8131 gnd.n6021 gnd.n6020 19.3944
R8132 gnd.n6020 gnd.n6019 19.3944
R8133 gnd.n6019 gnd.n738 19.3944
R8134 gnd.n6013 gnd.n738 19.3944
R8135 gnd.n6013 gnd.n6012 19.3944
R8136 gnd.n6012 gnd.n6011 19.3944
R8137 gnd.n6011 gnd.n746 19.3944
R8138 gnd.n6005 gnd.n746 19.3944
R8139 gnd.n6005 gnd.n6004 19.3944
R8140 gnd.n6004 gnd.n6003 19.3944
R8141 gnd.n6003 gnd.n754 19.3944
R8142 gnd.n5997 gnd.n754 19.3944
R8143 gnd.n5997 gnd.n5996 19.3944
R8144 gnd.n5996 gnd.n5995 19.3944
R8145 gnd.n5995 gnd.n762 19.3944
R8146 gnd.n5989 gnd.n762 19.3944
R8147 gnd.n5989 gnd.n5988 19.3944
R8148 gnd.n5988 gnd.n5987 19.3944
R8149 gnd.n5987 gnd.n770 19.3944
R8150 gnd.n5981 gnd.n770 19.3944
R8151 gnd.n5981 gnd.n5980 19.3944
R8152 gnd.n5980 gnd.n5979 19.3944
R8153 gnd.n5979 gnd.n778 19.3944
R8154 gnd.n5973 gnd.n778 19.3944
R8155 gnd.n5973 gnd.n5972 19.3944
R8156 gnd.n5972 gnd.n5971 19.3944
R8157 gnd.n5971 gnd.n786 19.3944
R8158 gnd.n5965 gnd.n786 19.3944
R8159 gnd.n5965 gnd.n5964 19.3944
R8160 gnd.n5964 gnd.n5963 19.3944
R8161 gnd.n5963 gnd.n794 19.3944
R8162 gnd.n5957 gnd.n794 19.3944
R8163 gnd.n5957 gnd.n5956 19.3944
R8164 gnd.n5956 gnd.n5955 19.3944
R8165 gnd.n5955 gnd.n802 19.3944
R8166 gnd.n2311 gnd.n802 19.3944
R8167 gnd.n4362 gnd.n4361 19.3944
R8168 gnd.n4361 gnd.n4360 19.3944
R8169 gnd.n4360 gnd.n1171 19.3944
R8170 gnd.n4356 gnd.n1171 19.3944
R8171 gnd.n4356 gnd.n4355 19.3944
R8172 gnd.n4355 gnd.n4354 19.3944
R8173 gnd.n4354 gnd.n1176 19.3944
R8174 gnd.n4350 gnd.n1176 19.3944
R8175 gnd.n4350 gnd.n4349 19.3944
R8176 gnd.n4349 gnd.n4348 19.3944
R8177 gnd.n4348 gnd.n1181 19.3944
R8178 gnd.n4344 gnd.n1181 19.3944
R8179 gnd.n4344 gnd.n4343 19.3944
R8180 gnd.n4343 gnd.n4342 19.3944
R8181 gnd.n4342 gnd.n1186 19.3944
R8182 gnd.n4338 gnd.n1186 19.3944
R8183 gnd.n4338 gnd.n4337 19.3944
R8184 gnd.n4337 gnd.n4336 19.3944
R8185 gnd.n4336 gnd.n1191 19.3944
R8186 gnd.n4332 gnd.n1191 19.3944
R8187 gnd.n4332 gnd.n4331 19.3944
R8188 gnd.n4331 gnd.n4330 19.3944
R8189 gnd.n4330 gnd.n1196 19.3944
R8190 gnd.n4326 gnd.n1196 19.3944
R8191 gnd.n4326 gnd.n4325 19.3944
R8192 gnd.n4325 gnd.n4324 19.3944
R8193 gnd.n4324 gnd.n1201 19.3944
R8194 gnd.n4320 gnd.n1201 19.3944
R8195 gnd.n4320 gnd.n4319 19.3944
R8196 gnd.n4319 gnd.n4318 19.3944
R8197 gnd.n4318 gnd.n1206 19.3944
R8198 gnd.n4314 gnd.n1206 19.3944
R8199 gnd.n4314 gnd.n4313 19.3944
R8200 gnd.n4313 gnd.n4312 19.3944
R8201 gnd.n4312 gnd.n1211 19.3944
R8202 gnd.n4308 gnd.n1211 19.3944
R8203 gnd.n4308 gnd.n4307 19.3944
R8204 gnd.n4307 gnd.n4306 19.3944
R8205 gnd.n4306 gnd.n1216 19.3944
R8206 gnd.n4302 gnd.n1216 19.3944
R8207 gnd.n4302 gnd.n4301 19.3944
R8208 gnd.n4301 gnd.n4300 19.3944
R8209 gnd.n4300 gnd.n1221 19.3944
R8210 gnd.n4296 gnd.n1221 19.3944
R8211 gnd.n4296 gnd.n4295 19.3944
R8212 gnd.n4295 gnd.n4294 19.3944
R8213 gnd.n4294 gnd.n1226 19.3944
R8214 gnd.n4290 gnd.n1226 19.3944
R8215 gnd.n4290 gnd.n4289 19.3944
R8216 gnd.n4289 gnd.n4288 19.3944
R8217 gnd.n4288 gnd.n1231 19.3944
R8218 gnd.n4284 gnd.n1231 19.3944
R8219 gnd.n4284 gnd.n4283 19.3944
R8220 gnd.n4283 gnd.n4282 19.3944
R8221 gnd.n4282 gnd.n1236 19.3944
R8222 gnd.n4278 gnd.n1236 19.3944
R8223 gnd.n4278 gnd.n4277 19.3944
R8224 gnd.n4277 gnd.n4276 19.3944
R8225 gnd.n4276 gnd.n1241 19.3944
R8226 gnd.n4272 gnd.n1241 19.3944
R8227 gnd.n4272 gnd.n4271 19.3944
R8228 gnd.n4271 gnd.n4270 19.3944
R8229 gnd.n4270 gnd.n1246 19.3944
R8230 gnd.n4266 gnd.n1246 19.3944
R8231 gnd.n4266 gnd.n4265 19.3944
R8232 gnd.n4265 gnd.n4264 19.3944
R8233 gnd.n4264 gnd.n1251 19.3944
R8234 gnd.n4260 gnd.n1251 19.3944
R8235 gnd.n4260 gnd.n4259 19.3944
R8236 gnd.n4259 gnd.n4258 19.3944
R8237 gnd.n4258 gnd.n1256 19.3944
R8238 gnd.n4254 gnd.n1256 19.3944
R8239 gnd.n4254 gnd.n4253 19.3944
R8240 gnd.n4253 gnd.n4252 19.3944
R8241 gnd.n4252 gnd.n1261 19.3944
R8242 gnd.n4248 gnd.n1261 19.3944
R8243 gnd.n4248 gnd.n4247 19.3944
R8244 gnd.n4247 gnd.n4246 19.3944
R8245 gnd.n4246 gnd.n1266 19.3944
R8246 gnd.n4242 gnd.n1266 19.3944
R8247 gnd.n4242 gnd.n4241 19.3944
R8248 gnd.n4241 gnd.n4240 19.3944
R8249 gnd.n3899 gnd.n1640 19.3944
R8250 gnd.n3895 gnd.n1640 19.3944
R8251 gnd.n3895 gnd.n3894 19.3944
R8252 gnd.n1557 gnd.n1546 19.3944
R8253 gnd.n1562 gnd.n1557 19.3944
R8254 gnd.n1562 gnd.n1539 19.3944
R8255 gnd.n1573 gnd.n1539 19.3944
R8256 gnd.n1573 gnd.n1537 19.3944
R8257 gnd.n1579 gnd.n1537 19.3944
R8258 gnd.n1579 gnd.n1530 19.3944
R8259 gnd.n1590 gnd.n1530 19.3944
R8260 gnd.n1590 gnd.n1528 19.3944
R8261 gnd.n1596 gnd.n1528 19.3944
R8262 gnd.n1596 gnd.n1521 19.3944
R8263 gnd.n1607 gnd.n1521 19.3944
R8264 gnd.n1607 gnd.n1519 19.3944
R8265 gnd.n1613 gnd.n1519 19.3944
R8266 gnd.n1613 gnd.n1509 19.3944
R8267 gnd.n1622 gnd.n1509 19.3944
R8268 gnd.n1622 gnd.n1507 19.3944
R8269 gnd.n1507 gnd.n1506 19.3944
R8270 gnd.n3910 gnd.n1506 19.3944
R8271 gnd.n3910 gnd.n3909 19.3944
R8272 gnd.n3909 gnd.n3908 19.3944
R8273 gnd.n3908 gnd.n1632 19.3944
R8274 gnd.n3904 gnd.n1632 19.3944
R8275 gnd.n3904 gnd.n3903 19.3944
R8276 gnd.n3107 gnd.t34 19.1199
R8277 gnd.n3229 gnd.n1850 19.1199
R8278 gnd.n3167 gnd.n1818 19.1199
R8279 gnd.n3400 gnd.n1778 19.1199
R8280 gnd.n3338 gnd.n1741 19.1199
R8281 gnd.n3460 gnd.t96 19.1199
R8282 gnd.n3716 gnd.n3715 19.1199
R8283 gnd.n5322 gnd.t283 18.8012
R8284 gnd.n5361 gnd.t17 18.8012
R8285 gnd.n5165 gnd.n4907 18.4825
R8286 gnd.t187 gnd.n1665 18.4825
R8287 gnd.n4198 gnd.n4197 18.4247
R8288 gnd.n2834 gnd.n2833 18.4247
R8289 gnd.n6839 gnd.n6838 18.2308
R8290 gnd.n1618 gnd.n1617 18.2308
R8291 gnd.n2866 gnd.n2014 18.2308
R8292 gnd.n2386 gnd.n2379 18.2308
R8293 gnd.t94 gnd.n4849 18.1639
R8294 gnd.n1952 gnd.t228 18.1639
R8295 gnd.t64 gnd.n1671 18.1639
R8296 gnd.n3064 gnd.n1918 17.8452
R8297 gnd.n2968 gnd.n1896 17.8452
R8298 gnd.n3143 gnd.n1826 17.8452
R8299 gnd.n3408 gnd.n1770 17.8452
R8300 gnd.n3814 gnd.n1698 17.8452
R8301 gnd.n3489 gnd.n1678 17.8452
R8302 gnd.n4878 gnd.t249 17.5266
R8303 gnd.n3237 gnd.t224 17.5266
R8304 gnd.n3314 gnd.t66 17.5266
R8305 gnd.t1 gnd.n1926 17.2079
R8306 gnd.n3745 gnd.t47 17.2079
R8307 gnd.t68 gnd.n4825 16.8893
R8308 gnd.n2435 gnd.t203 16.8893
R8309 gnd.n2201 gnd.t9 16.8893
R8310 gnd.n4039 gnd.t11 16.8893
R8311 gnd.t118 gnd.n81 16.8893
R8312 gnd.n3072 gnd.n1910 16.5706
R8313 gnd.n3009 gnd.n3008 16.5706
R8314 gnd.n3245 gnd.n1837 16.5706
R8315 gnd.n3182 gnd.n3181 16.5706
R8316 gnd.n3416 gnd.n1763 16.5706
R8317 gnd.n3353 gnd.n3352 16.5706
R8318 gnd.n3822 gnd.n1691 16.5706
R8319 gnd.n3759 gnd.n3758 16.5706
R8320 gnd.t219 gnd.n4934 16.2519
R8321 gnd.n4792 gnd.t84 16.2519
R8322 gnd.n2214 gnd.t70 16.2519
R8323 gnd.n1979 gnd.t190 16.2519
R8324 gnd.t174 gnd.n1272 16.2519
R8325 gnd.n4090 gnd.t51 16.2519
R8326 gnd.n2987 gnd.t110 15.9333
R8327 gnd.t74 gnd.n1712 15.9333
R8328 gnd.n5784 gnd.n5782 15.6674
R8329 gnd.n5752 gnd.n5750 15.6674
R8330 gnd.n5720 gnd.n5718 15.6674
R8331 gnd.n5689 gnd.n5687 15.6674
R8332 gnd.n5657 gnd.n5655 15.6674
R8333 gnd.n5625 gnd.n5623 15.6674
R8334 gnd.n5593 gnd.n5591 15.6674
R8335 gnd.n5562 gnd.n5560 15.6674
R8336 gnd.n5052 gnd.t219 15.6146
R8337 gnd.n5822 gnd.t153 15.6146
R8338 gnd.n5923 gnd.t167 15.6146
R8339 gnd.t13 gnd.n1024 15.6146
R8340 gnd.n2916 gnd.t190 15.6146
R8341 gnd.n3883 gnd.t174 15.6146
R8342 gnd.n6727 gnd.t246 15.6146
R8343 gnd.n3524 gnd.n3523 15.0827
R8344 gnd.n2657 gnd.n2652 15.0481
R8345 gnd.n3534 gnd.n3533 15.0481
R8346 gnd.n5488 gnd.t251 14.9773
R8347 gnd.t203 gnd.n960 14.9773
R8348 gnd.n4375 gnd.t139 14.9773
R8349 gnd.t132 gnd.n3956 14.9773
R8350 gnd.n6882 gnd.t118 14.9773
R8351 gnd.n3080 gnd.t4 14.6587
R8352 gnd.n3473 gnd.t226 14.6587
R8353 gnd.t273 gnd.n5526 14.34
R8354 gnd.n5544 gnd.t93 14.34
R8355 gnd.n3024 gnd.n1918 14.0214
R8356 gnd.t79 gnd.n1896 14.0214
R8357 gnd.n3197 gnd.n3196 14.0214
R8358 gnd.n3261 gnd.n1826 14.0214
R8359 gnd.n3368 gnd.n1770 14.0214
R8360 gnd.n3432 gnd.n1750 14.0214
R8361 gnd.t232 gnd.n1698 14.0214
R8362 gnd.n3838 gnd.n1678 14.0214
R8363 gnd.n3515 gnd.t115 14.0214
R8364 gnd.n94 gnd.n83 14.0214
R8365 gnd.t21 gnd.n5249 13.7027
R8366 gnd.t252 gnd.n1912 13.7027
R8367 gnd.n3760 gnd.t270 13.7027
R8368 gnd.n5134 gnd.n5130 13.5763
R8369 gnd.n5886 gnd.n4596 13.5763
R8370 gnd.n4160 gnd.n1358 13.5763
R8371 gnd.n6891 gnd.n6890 13.5763
R8372 gnd.n4501 gnd.n952 13.5763
R8373 gnd.n2587 gnd.n2584 13.5763
R8374 gnd.n5166 gnd.n5165 13.384
R8375 gnd.n2668 gnd.n2649 13.1884
R8376 gnd.n2663 gnd.n2662 13.1884
R8377 gnd.n2662 gnd.n2661 13.1884
R8378 gnd.n3527 gnd.n3522 13.1884
R8379 gnd.n3528 gnd.n3527 13.1884
R8380 gnd.n2664 gnd.n2651 13.146
R8381 gnd.n2660 gnd.n2651 13.146
R8382 gnd.n3526 gnd.n3525 13.146
R8383 gnd.n3526 gnd.n3521 13.146
R8384 gnd.n5785 gnd.n5781 12.8005
R8385 gnd.n5753 gnd.n5749 12.8005
R8386 gnd.n5721 gnd.n5717 12.8005
R8387 gnd.n5690 gnd.n5686 12.8005
R8388 gnd.n5658 gnd.n5654 12.8005
R8389 gnd.n5626 gnd.n5622 12.8005
R8390 gnd.n5594 gnd.n5590 12.8005
R8391 gnd.n5563 gnd.n5559 12.8005
R8392 gnd.n2926 gnd.n1963 12.7467
R8393 gnd.t150 gnd.t157 12.7467
R8394 gnd.n1952 gnd.n1951 12.7467
R8395 gnd.t254 gnd.n1910 12.7467
R8396 gnd.n3097 gnd.n1888 12.7467
R8397 gnd.n1875 gnd.n1850 12.7467
R8398 gnd.n3271 gnd.n1818 12.7467
R8399 gnd.t107 gnd.n1819 12.7467
R8400 gnd.n3376 gnd.t54 12.7467
R8401 gnd.n1804 gnd.n1778 12.7467
R8402 gnd.n3442 gnd.n1741 12.7467
R8403 gnd.n1729 gnd.n1727 12.7467
R8404 gnd.n3758 gnd.t97 12.7467
R8405 gnd.n3846 gnd.n1671 12.7467
R8406 gnd.t200 gnd.n1664 12.7467
R8407 gnd.t275 gnd.n1888 12.4281
R8408 gnd.n1729 gnd.t242 12.4281
R8409 gnd.n5137 gnd.n5134 12.4126
R8410 gnd.n5889 gnd.n5886 12.4126
R8411 gnd.n4156 gnd.n1358 12.4126
R8412 gnd.n6890 gnd.n156 12.4126
R8413 gnd.n4497 gnd.n952 12.4126
R8414 gnd.n2584 gnd.n2179 12.4126
R8415 gnd.n2750 gnd.n2669 12.1761
R8416 gnd.n3561 gnd.n3539 12.1761
R8417 gnd.n5789 gnd.n5788 12.0247
R8418 gnd.n5757 gnd.n5756 12.0247
R8419 gnd.n5725 gnd.n5724 12.0247
R8420 gnd.n5694 gnd.n5693 12.0247
R8421 gnd.n5662 gnd.n5661 12.0247
R8422 gnd.n5630 gnd.n5629 12.0247
R8423 gnd.n5598 gnd.n5597 12.0247
R8424 gnd.n5567 gnd.n5566 12.0247
R8425 gnd.t240 gnd.n974 11.7908
R8426 gnd.n2184 gnd.t139 11.7908
R8427 gnd.n3973 gnd.t132 11.7908
R8428 gnd.n6792 gnd.t263 11.7908
R8429 gnd.n2935 gnd.n1956 11.4721
R8430 gnd.n3106 gnd.n1880 11.4721
R8431 gnd.n1865 gnd.n1857 11.4721
R8432 gnd.n3281 gnd.n3280 11.4721
R8433 gnd.n1795 gnd.n1785 11.4721
R8434 gnd.n3452 gnd.n3451 11.4721
R8435 gnd.n3459 gnd.n1711 11.4721
R8436 gnd.n3854 gnd.n1664 11.4721
R8437 gnd.n3862 gnd.n1658 11.4721
R8438 gnd.n5792 gnd.n5779 11.249
R8439 gnd.n5760 gnd.n5747 11.249
R8440 gnd.n5728 gnd.n5715 11.249
R8441 gnd.n5697 gnd.n5684 11.249
R8442 gnd.n5665 gnd.n5652 11.249
R8443 gnd.n5633 gnd.n5620 11.249
R8444 gnd.n5601 gnd.n5588 11.249
R8445 gnd.n5570 gnd.n5557 11.249
R8446 gnd.n5250 gnd.t21 11.1535
R8447 gnd.n2471 gnd.t13 11.1535
R8448 gnd.n6760 gnd.t246 11.1535
R8449 gnd.t194 gnd.n1963 10.8348
R8450 gnd.t222 gnd.n1858 10.8348
R8451 gnd.n3205 gnd.t222 10.8348
R8452 gnd.t0 gnd.n1743 10.8348
R8453 gnd.n3331 gnd.t0 10.8348
R8454 gnd.n3711 gnd.n3710 10.6151
R8455 gnd.n3710 gnd.n3707 10.6151
R8456 gnd.n3705 gnd.n3702 10.6151
R8457 gnd.n3702 gnd.n3701 10.6151
R8458 gnd.n3701 gnd.n3698 10.6151
R8459 gnd.n3698 gnd.n3697 10.6151
R8460 gnd.n3697 gnd.n3694 10.6151
R8461 gnd.n3694 gnd.n3693 10.6151
R8462 gnd.n3693 gnd.n3690 10.6151
R8463 gnd.n3690 gnd.n3689 10.6151
R8464 gnd.n3689 gnd.n3686 10.6151
R8465 gnd.n3686 gnd.n3685 10.6151
R8466 gnd.n3685 gnd.n3682 10.6151
R8467 gnd.n3682 gnd.n3681 10.6151
R8468 gnd.n3681 gnd.n3678 10.6151
R8469 gnd.n3678 gnd.n3677 10.6151
R8470 gnd.n3677 gnd.n3674 10.6151
R8471 gnd.n3674 gnd.n3673 10.6151
R8472 gnd.n3673 gnd.n3670 10.6151
R8473 gnd.n3670 gnd.n3669 10.6151
R8474 gnd.n3669 gnd.n3666 10.6151
R8475 gnd.n3666 gnd.n3665 10.6151
R8476 gnd.n3665 gnd.n3662 10.6151
R8477 gnd.n3662 gnd.n3661 10.6151
R8478 gnd.n3661 gnd.n3658 10.6151
R8479 gnd.n3658 gnd.n3657 10.6151
R8480 gnd.n3657 gnd.n3654 10.6151
R8481 gnd.n3654 gnd.n3653 10.6151
R8482 gnd.n3653 gnd.n3650 10.6151
R8483 gnd.n3650 gnd.n3649 10.6151
R8484 gnd.n2762 gnd.n2646 10.6151
R8485 gnd.n2762 gnd.n2761 10.6151
R8486 gnd.n2761 gnd.n2760 10.6151
R8487 gnd.n2760 gnd.n1946 10.6151
R8488 gnd.n3038 gnd.n1946 10.6151
R8489 gnd.n3038 gnd.n3037 10.6151
R8490 gnd.n3037 gnd.n3036 10.6151
R8491 gnd.n3036 gnd.n1947 10.6151
R8492 gnd.n1949 gnd.n1947 10.6151
R8493 gnd.n2949 gnd.n1949 10.6151
R8494 gnd.n2950 gnd.n2949 10.6151
R8495 gnd.n3022 gnd.n2950 10.6151
R8496 gnd.n3022 gnd.n3021 10.6151
R8497 gnd.n3021 gnd.n3020 10.6151
R8498 gnd.n3020 gnd.n2951 10.6151
R8499 gnd.n2962 gnd.n2951 10.6151
R8500 gnd.n2964 gnd.n2962 10.6151
R8501 gnd.n2965 gnd.n2964 10.6151
R8502 gnd.n3006 gnd.n2965 10.6151
R8503 gnd.n3006 gnd.n3005 10.6151
R8504 gnd.n3005 gnd.n3004 10.6151
R8505 gnd.n3004 gnd.n2966 10.6151
R8506 gnd.n2977 gnd.n2966 10.6151
R8507 gnd.n2992 gnd.n2977 10.6151
R8508 gnd.n2992 gnd.n2991 10.6151
R8509 gnd.n2991 gnd.n2990 10.6151
R8510 gnd.n2990 gnd.n2978 10.6151
R8511 gnd.n2979 gnd.n2978 10.6151
R8512 gnd.n2979 gnd.n1870 10.6151
R8513 gnd.n3211 gnd.n1870 10.6151
R8514 gnd.n3211 gnd.n3210 10.6151
R8515 gnd.n3210 gnd.n3209 10.6151
R8516 gnd.n3209 gnd.n1871 10.6151
R8517 gnd.n1873 gnd.n1871 10.6151
R8518 gnd.n3120 gnd.n1873 10.6151
R8519 gnd.n3122 gnd.n3120 10.6151
R8520 gnd.n3123 gnd.n3122 10.6151
R8521 gnd.n3194 gnd.n3123 10.6151
R8522 gnd.n3194 gnd.n3193 10.6151
R8523 gnd.n3193 gnd.n3192 10.6151
R8524 gnd.n3192 gnd.n3124 10.6151
R8525 gnd.n3137 gnd.n3124 10.6151
R8526 gnd.n3138 gnd.n3137 10.6151
R8527 gnd.n3179 gnd.n3138 10.6151
R8528 gnd.n3179 gnd.n3178 10.6151
R8529 gnd.n3178 gnd.n3177 10.6151
R8530 gnd.n3177 gnd.n3139 10.6151
R8531 gnd.n3157 gnd.n3139 10.6151
R8532 gnd.n3165 gnd.n3157 10.6151
R8533 gnd.n3165 gnd.n3164 10.6151
R8534 gnd.n3164 gnd.n3163 10.6151
R8535 gnd.n3163 gnd.n3159 10.6151
R8536 gnd.n3159 gnd.n3158 10.6151
R8537 gnd.n3158 gnd.n1800 10.6151
R8538 gnd.n3382 gnd.n1800 10.6151
R8539 gnd.n3382 gnd.n3381 10.6151
R8540 gnd.n3381 gnd.n3380 10.6151
R8541 gnd.n3380 gnd.n1801 10.6151
R8542 gnd.n1803 gnd.n1801 10.6151
R8543 gnd.n3295 gnd.n1803 10.6151
R8544 gnd.n3296 gnd.n3295 10.6151
R8545 gnd.n3366 gnd.n3296 10.6151
R8546 gnd.n3366 gnd.n3365 10.6151
R8547 gnd.n3365 gnd.n3364 10.6151
R8548 gnd.n3364 gnd.n3297 10.6151
R8549 gnd.n3308 gnd.n3297 10.6151
R8550 gnd.n3310 gnd.n3308 10.6151
R8551 gnd.n3311 gnd.n3310 10.6151
R8552 gnd.n3350 gnd.n3311 10.6151
R8553 gnd.n3350 gnd.n3349 10.6151
R8554 gnd.n3349 gnd.n3348 10.6151
R8555 gnd.n3348 gnd.n3312 10.6151
R8556 gnd.n3328 gnd.n3312 10.6151
R8557 gnd.n3336 gnd.n3328 10.6151
R8558 gnd.n3336 gnd.n3335 10.6151
R8559 gnd.n3335 gnd.n3334 10.6151
R8560 gnd.n3334 gnd.n3330 10.6151
R8561 gnd.n3330 gnd.n3329 10.6151
R8562 gnd.n3329 gnd.n1723 10.6151
R8563 gnd.n3788 gnd.n1723 10.6151
R8564 gnd.n3788 gnd.n3787 10.6151
R8565 gnd.n3787 gnd.n3786 10.6151
R8566 gnd.n3786 gnd.n1724 10.6151
R8567 gnd.n1726 gnd.n1724 10.6151
R8568 gnd.n3469 gnd.n1726 10.6151
R8569 gnd.n3470 gnd.n3469 10.6151
R8570 gnd.n3772 gnd.n3470 10.6151
R8571 gnd.n3772 gnd.n3771 10.6151
R8572 gnd.n3771 gnd.n3770 10.6151
R8573 gnd.n3770 gnd.n3471 10.6151
R8574 gnd.n3483 gnd.n3471 10.6151
R8575 gnd.n3485 gnd.n3483 10.6151
R8576 gnd.n3486 gnd.n3485 10.6151
R8577 gnd.n3756 gnd.n3486 10.6151
R8578 gnd.n3756 gnd.n3755 10.6151
R8579 gnd.n3755 gnd.n3754 10.6151
R8580 gnd.n3754 gnd.n3487 10.6151
R8581 gnd.n3498 gnd.n3487 10.6151
R8582 gnd.n3741 gnd.n3498 10.6151
R8583 gnd.n3741 gnd.n3740 10.6151
R8584 gnd.n3740 gnd.n3739 10.6151
R8585 gnd.n3739 gnd.n3499 10.6151
R8586 gnd.n3511 gnd.n3499 10.6151
R8587 gnd.n3512 gnd.n3511 10.6151
R8588 gnd.n3727 gnd.n3512 10.6151
R8589 gnd.n3727 gnd.n3726 10.6151
R8590 gnd.n3726 gnd.n3725 10.6151
R8591 gnd.n3725 gnd.n3513 10.6151
R8592 gnd.n3646 gnd.n3513 10.6151
R8593 gnd.n3647 gnd.n3646 10.6151
R8594 gnd.n2826 gnd.n2626 10.6151
R8595 gnd.n2826 gnd.n2825 10.6151
R8596 gnd.n2823 gnd.n2632 10.6151
R8597 gnd.n2817 gnd.n2632 10.6151
R8598 gnd.n2817 gnd.n2816 10.6151
R8599 gnd.n2816 gnd.n2815 10.6151
R8600 gnd.n2815 gnd.n2634 10.6151
R8601 gnd.n2809 gnd.n2634 10.6151
R8602 gnd.n2809 gnd.n2808 10.6151
R8603 gnd.n2808 gnd.n2807 10.6151
R8604 gnd.n2807 gnd.n2636 10.6151
R8605 gnd.n2801 gnd.n2636 10.6151
R8606 gnd.n2801 gnd.n2800 10.6151
R8607 gnd.n2800 gnd.n2799 10.6151
R8608 gnd.n2799 gnd.n2638 10.6151
R8609 gnd.n2793 gnd.n2638 10.6151
R8610 gnd.n2793 gnd.n2792 10.6151
R8611 gnd.n2792 gnd.n2791 10.6151
R8612 gnd.n2791 gnd.n2640 10.6151
R8613 gnd.n2785 gnd.n2640 10.6151
R8614 gnd.n2785 gnd.n2784 10.6151
R8615 gnd.n2784 gnd.n2783 10.6151
R8616 gnd.n2783 gnd.n2642 10.6151
R8617 gnd.n2777 gnd.n2642 10.6151
R8618 gnd.n2777 gnd.n2776 10.6151
R8619 gnd.n2776 gnd.n2775 10.6151
R8620 gnd.n2775 gnd.n2644 10.6151
R8621 gnd.n2769 gnd.n2644 10.6151
R8622 gnd.n2769 gnd.n2768 10.6151
R8623 gnd.n2768 gnd.n2767 10.6151
R8624 gnd.n2750 gnd.n2749 10.6151
R8625 gnd.n2749 gnd.n2671 10.6151
R8626 gnd.n2745 gnd.n2671 10.6151
R8627 gnd.n2745 gnd.n2744 10.6151
R8628 gnd.n2744 gnd.n2673 10.6151
R8629 gnd.n2739 gnd.n2673 10.6151
R8630 gnd.n2739 gnd.n2738 10.6151
R8631 gnd.n2738 gnd.n2737 10.6151
R8632 gnd.n2737 gnd.n2675 10.6151
R8633 gnd.n2731 gnd.n2675 10.6151
R8634 gnd.n2731 gnd.n2730 10.6151
R8635 gnd.n2730 gnd.n2729 10.6151
R8636 gnd.n2729 gnd.n2677 10.6151
R8637 gnd.n2723 gnd.n2677 10.6151
R8638 gnd.n2723 gnd.n2722 10.6151
R8639 gnd.n2722 gnd.n2721 10.6151
R8640 gnd.n2721 gnd.n2679 10.6151
R8641 gnd.n2715 gnd.n2679 10.6151
R8642 gnd.n2715 gnd.n2714 10.6151
R8643 gnd.n2714 gnd.n2713 10.6151
R8644 gnd.n2713 gnd.n2681 10.6151
R8645 gnd.n2707 gnd.n2681 10.6151
R8646 gnd.n2707 gnd.n2706 10.6151
R8647 gnd.n2706 gnd.n2705 10.6151
R8648 gnd.n2705 gnd.n2683 10.6151
R8649 gnd.n2699 gnd.n2683 10.6151
R8650 gnd.n2699 gnd.n2698 10.6151
R8651 gnd.n2698 gnd.n2697 10.6151
R8652 gnd.n2693 gnd.n2692 10.6151
R8653 gnd.n2692 gnd.n2627 10.6151
R8654 gnd.n3562 gnd.n3561 10.6151
R8655 gnd.n3565 gnd.n3562 10.6151
R8656 gnd.n3566 gnd.n3565 10.6151
R8657 gnd.n3569 gnd.n3566 10.6151
R8658 gnd.n3570 gnd.n3569 10.6151
R8659 gnd.n3573 gnd.n3570 10.6151
R8660 gnd.n3574 gnd.n3573 10.6151
R8661 gnd.n3577 gnd.n3574 10.6151
R8662 gnd.n3578 gnd.n3577 10.6151
R8663 gnd.n3581 gnd.n3578 10.6151
R8664 gnd.n3582 gnd.n3581 10.6151
R8665 gnd.n3585 gnd.n3582 10.6151
R8666 gnd.n3586 gnd.n3585 10.6151
R8667 gnd.n3589 gnd.n3586 10.6151
R8668 gnd.n3590 gnd.n3589 10.6151
R8669 gnd.n3593 gnd.n3590 10.6151
R8670 gnd.n3594 gnd.n3593 10.6151
R8671 gnd.n3597 gnd.n3594 10.6151
R8672 gnd.n3598 gnd.n3597 10.6151
R8673 gnd.n3601 gnd.n3598 10.6151
R8674 gnd.n3602 gnd.n3601 10.6151
R8675 gnd.n3605 gnd.n3602 10.6151
R8676 gnd.n3606 gnd.n3605 10.6151
R8677 gnd.n3609 gnd.n3606 10.6151
R8678 gnd.n3610 gnd.n3609 10.6151
R8679 gnd.n3613 gnd.n3610 10.6151
R8680 gnd.n3614 gnd.n3613 10.6151
R8681 gnd.n3617 gnd.n3614 10.6151
R8682 gnd.n3622 gnd.n3619 10.6151
R8683 gnd.n3623 gnd.n3622 10.6151
R8684 gnd.n2754 gnd.n2753 10.6151
R8685 gnd.n2755 gnd.n2754 10.6151
R8686 gnd.n2755 gnd.n1954 10.6151
R8687 gnd.n2938 gnd.n1954 10.6151
R8688 gnd.n2939 gnd.n2938 10.6151
R8689 gnd.n2940 gnd.n2939 10.6151
R8690 gnd.n2943 gnd.n2940 10.6151
R8691 gnd.n2944 gnd.n2943 10.6151
R8692 gnd.n3030 gnd.n2944 10.6151
R8693 gnd.n3030 gnd.n3029 10.6151
R8694 gnd.n3029 gnd.n3028 10.6151
R8695 gnd.n3028 gnd.n2945 10.6151
R8696 gnd.n2956 gnd.n2945 10.6151
R8697 gnd.n2957 gnd.n2956 10.6151
R8698 gnd.n3015 gnd.n2957 10.6151
R8699 gnd.n3015 gnd.n3014 10.6151
R8700 gnd.n3014 gnd.n3013 10.6151
R8701 gnd.n3013 gnd.n2958 10.6151
R8702 gnd.n2971 gnd.n2958 10.6151
R8703 gnd.n2972 gnd.n2971 10.6151
R8704 gnd.n3000 gnd.n2972 10.6151
R8705 gnd.n3000 gnd.n2999 10.6151
R8706 gnd.n2999 gnd.n2998 10.6151
R8707 gnd.n2998 gnd.n2973 10.6151
R8708 gnd.n2983 gnd.n2973 10.6151
R8709 gnd.n2984 gnd.n2983 10.6151
R8710 gnd.n2985 gnd.n2984 10.6151
R8711 gnd.n2985 gnd.n1878 10.6151
R8712 gnd.n3109 gnd.n1878 10.6151
R8713 gnd.n3110 gnd.n3109 10.6151
R8714 gnd.n3111 gnd.n3110 10.6151
R8715 gnd.n3114 gnd.n3111 10.6151
R8716 gnd.n3115 gnd.n3114 10.6151
R8717 gnd.n3203 gnd.n3115 10.6151
R8718 gnd.n3203 gnd.n3202 10.6151
R8719 gnd.n3202 gnd.n3201 10.6151
R8720 gnd.n3201 gnd.n3116 10.6151
R8721 gnd.n3130 gnd.n3116 10.6151
R8722 gnd.n3131 gnd.n3130 10.6151
R8723 gnd.n3188 gnd.n3131 10.6151
R8724 gnd.n3188 gnd.n3187 10.6151
R8725 gnd.n3187 gnd.n3186 10.6151
R8726 gnd.n3186 gnd.n3132 10.6151
R8727 gnd.n3146 gnd.n3132 10.6151
R8728 gnd.n3147 gnd.n3146 10.6151
R8729 gnd.n3173 gnd.n3147 10.6151
R8730 gnd.n3173 gnd.n3172 10.6151
R8731 gnd.n3172 gnd.n3171 10.6151
R8732 gnd.n3171 gnd.n3148 10.6151
R8733 gnd.n3152 gnd.n3148 10.6151
R8734 gnd.n3152 gnd.n3151 10.6151
R8735 gnd.n3151 gnd.n3150 10.6151
R8736 gnd.n3150 gnd.n1807 10.6151
R8737 gnd.n3284 gnd.n1807 10.6151
R8738 gnd.n3285 gnd.n3284 10.6151
R8739 gnd.n3286 gnd.n3285 10.6151
R8740 gnd.n3289 gnd.n3286 10.6151
R8741 gnd.n3290 gnd.n3289 10.6151
R8742 gnd.n3374 gnd.n3290 10.6151
R8743 gnd.n3374 gnd.n3373 10.6151
R8744 gnd.n3373 gnd.n3372 10.6151
R8745 gnd.n3372 gnd.n3291 10.6151
R8746 gnd.n3302 gnd.n3291 10.6151
R8747 gnd.n3303 gnd.n3302 10.6151
R8748 gnd.n3359 gnd.n3303 10.6151
R8749 gnd.n3359 gnd.n3358 10.6151
R8750 gnd.n3358 gnd.n3357 10.6151
R8751 gnd.n3357 gnd.n3304 10.6151
R8752 gnd.n3317 gnd.n3304 10.6151
R8753 gnd.n3318 gnd.n3317 10.6151
R8754 gnd.n3344 gnd.n3318 10.6151
R8755 gnd.n3344 gnd.n3343 10.6151
R8756 gnd.n3343 gnd.n3342 10.6151
R8757 gnd.n3342 gnd.n3319 10.6151
R8758 gnd.n3323 gnd.n3319 10.6151
R8759 gnd.n3323 gnd.n3322 10.6151
R8760 gnd.n3322 gnd.n3321 10.6151
R8761 gnd.n3321 gnd.n1731 10.6151
R8762 gnd.n3455 gnd.n1731 10.6151
R8763 gnd.n3456 gnd.n3455 10.6151
R8764 gnd.n3457 gnd.n3456 10.6151
R8765 gnd.n3463 gnd.n3457 10.6151
R8766 gnd.n3464 gnd.n3463 10.6151
R8767 gnd.n3780 gnd.n3464 10.6151
R8768 gnd.n3780 gnd.n3779 10.6151
R8769 gnd.n3779 gnd.n3778 10.6151
R8770 gnd.n3778 gnd.n3465 10.6151
R8771 gnd.n3476 gnd.n3465 10.6151
R8772 gnd.n3477 gnd.n3476 10.6151
R8773 gnd.n3765 gnd.n3477 10.6151
R8774 gnd.n3765 gnd.n3764 10.6151
R8775 gnd.n3764 gnd.n3763 10.6151
R8776 gnd.n3763 gnd.n3478 10.6151
R8777 gnd.n3492 gnd.n3478 10.6151
R8778 gnd.n3493 gnd.n3492 10.6151
R8779 gnd.n3750 gnd.n3493 10.6151
R8780 gnd.n3750 gnd.n3749 10.6151
R8781 gnd.n3749 gnd.n3748 10.6151
R8782 gnd.n3748 gnd.n3494 10.6151
R8783 gnd.n3504 gnd.n3494 10.6151
R8784 gnd.n3505 gnd.n3504 10.6151
R8785 gnd.n3734 gnd.n3505 10.6151
R8786 gnd.n3734 gnd.n3733 10.6151
R8787 gnd.n3733 gnd.n3732 10.6151
R8788 gnd.n3732 gnd.n3506 10.6151
R8789 gnd.n3518 gnd.n3506 10.6151
R8790 gnd.n3519 gnd.n3518 10.6151
R8791 gnd.n3720 gnd.n3519 10.6151
R8792 gnd.n3720 gnd.n3719 10.6151
R8793 gnd.n3719 gnd.n3718 10.6151
R8794 gnd.n4922 gnd.t15 10.5161
R8795 gnd.n5527 gnd.t273 10.5161
R8796 gnd.n5937 gnd.t93 10.5161
R8797 gnd.n4430 gnd.t70 10.5161
R8798 gnd.t51 gnd.n1402 10.5161
R8799 gnd.n5793 gnd.n5777 10.4732
R8800 gnd.n5761 gnd.n5745 10.4732
R8801 gnd.n5729 gnd.n5713 10.4732
R8802 gnd.n5698 gnd.n5682 10.4732
R8803 gnd.n5666 gnd.n5650 10.4732
R8804 gnd.n5634 gnd.n5618 10.4732
R8805 gnd.n5602 gnd.n5586 10.4732
R8806 gnd.n5571 gnd.n5555 10.4732
R8807 gnd.n2936 gnd.n2935 10.1975
R8808 gnd.n1942 gnd.n1941 10.1975
R8809 gnd.n3107 gnd.n3106 10.1975
R8810 gnd.n3280 gnd.n1793 10.1975
R8811 gnd.n1796 gnd.n1795 10.1975
R8812 gnd.n3460 gnd.n3459 10.1975
R8813 gnd.n3854 gnd.n1665 10.1975
R8814 gnd.n3862 gnd.n1657 10.1975
R8815 gnd.n5502 gnd.t251 9.87883
R8816 gnd.n2461 gnd.t32 9.87883
R8817 gnd.n4405 gnd.t9 9.87883
R8818 gnd.n3936 gnd.t11 9.87883
R8819 gnd.n6768 gnd.t23 9.87883
R8820 gnd.n5797 gnd.n5796 9.69747
R8821 gnd.n5765 gnd.n5764 9.69747
R8822 gnd.n5733 gnd.n5732 9.69747
R8823 gnd.n5702 gnd.n5701 9.69747
R8824 gnd.n5670 gnd.n5669 9.69747
R8825 gnd.n5638 gnd.n5637 9.69747
R8826 gnd.n5606 gnd.n5605 9.69747
R8827 gnd.n5575 gnd.n5574 9.69747
R8828 gnd.n6997 gnd.n50 9.6512
R8829 gnd.n3127 gnd.t31 9.56018
R8830 gnd.n3424 gnd.t255 9.56018
R8831 gnd.n4365 gnd.n1165 9.45599
R8832 gnd.n1548 gnd.n1368 9.45599
R8833 gnd.n5803 gnd.n5802 9.45567
R8834 gnd.n5771 gnd.n5770 9.45567
R8835 gnd.n5739 gnd.n5738 9.45567
R8836 gnd.n5708 gnd.n5707 9.45567
R8837 gnd.n5676 gnd.n5675 9.45567
R8838 gnd.n5644 gnd.n5643 9.45567
R8839 gnd.n5612 gnd.n5611 9.45567
R8840 gnd.n5581 gnd.n5580 9.45567
R8841 gnd.n4766 gnd.n4765 9.39724
R8842 gnd.n5802 gnd.n5801 9.3005
R8843 gnd.n5775 gnd.n5774 9.3005
R8844 gnd.n5796 gnd.n5795 9.3005
R8845 gnd.n5794 gnd.n5793 9.3005
R8846 gnd.n5779 gnd.n5778 9.3005
R8847 gnd.n5788 gnd.n5787 9.3005
R8848 gnd.n5786 gnd.n5785 9.3005
R8849 gnd.n5770 gnd.n5769 9.3005
R8850 gnd.n5743 gnd.n5742 9.3005
R8851 gnd.n5764 gnd.n5763 9.3005
R8852 gnd.n5762 gnd.n5761 9.3005
R8853 gnd.n5747 gnd.n5746 9.3005
R8854 gnd.n5756 gnd.n5755 9.3005
R8855 gnd.n5754 gnd.n5753 9.3005
R8856 gnd.n5738 gnd.n5737 9.3005
R8857 gnd.n5711 gnd.n5710 9.3005
R8858 gnd.n5732 gnd.n5731 9.3005
R8859 gnd.n5730 gnd.n5729 9.3005
R8860 gnd.n5715 gnd.n5714 9.3005
R8861 gnd.n5724 gnd.n5723 9.3005
R8862 gnd.n5722 gnd.n5721 9.3005
R8863 gnd.n5707 gnd.n5706 9.3005
R8864 gnd.n5680 gnd.n5679 9.3005
R8865 gnd.n5701 gnd.n5700 9.3005
R8866 gnd.n5699 gnd.n5698 9.3005
R8867 gnd.n5684 gnd.n5683 9.3005
R8868 gnd.n5693 gnd.n5692 9.3005
R8869 gnd.n5691 gnd.n5690 9.3005
R8870 gnd.n5675 gnd.n5674 9.3005
R8871 gnd.n5648 gnd.n5647 9.3005
R8872 gnd.n5669 gnd.n5668 9.3005
R8873 gnd.n5667 gnd.n5666 9.3005
R8874 gnd.n5652 gnd.n5651 9.3005
R8875 gnd.n5661 gnd.n5660 9.3005
R8876 gnd.n5659 gnd.n5658 9.3005
R8877 gnd.n5643 gnd.n5642 9.3005
R8878 gnd.n5616 gnd.n5615 9.3005
R8879 gnd.n5637 gnd.n5636 9.3005
R8880 gnd.n5635 gnd.n5634 9.3005
R8881 gnd.n5620 gnd.n5619 9.3005
R8882 gnd.n5629 gnd.n5628 9.3005
R8883 gnd.n5627 gnd.n5626 9.3005
R8884 gnd.n5611 gnd.n5610 9.3005
R8885 gnd.n5584 gnd.n5583 9.3005
R8886 gnd.n5605 gnd.n5604 9.3005
R8887 gnd.n5603 gnd.n5602 9.3005
R8888 gnd.n5588 gnd.n5587 9.3005
R8889 gnd.n5597 gnd.n5596 9.3005
R8890 gnd.n5595 gnd.n5594 9.3005
R8891 gnd.n5580 gnd.n5579 9.3005
R8892 gnd.n5553 gnd.n5552 9.3005
R8893 gnd.n5574 gnd.n5573 9.3005
R8894 gnd.n5572 gnd.n5571 9.3005
R8895 gnd.n5557 gnd.n5556 9.3005
R8896 gnd.n5566 gnd.n5565 9.3005
R8897 gnd.n5564 gnd.n5563 9.3005
R8898 gnd.n861 gnd.n860 9.3005
R8899 gnd.n5911 gnd.n4583 9.3005
R8900 gnd.n5910 gnd.n4584 9.3005
R8901 gnd.n5909 gnd.n4585 9.3005
R8902 gnd.n5906 gnd.n4586 9.3005
R8903 gnd.n5905 gnd.n4587 9.3005
R8904 gnd.n5902 gnd.n4588 9.3005
R8905 gnd.n5901 gnd.n4589 9.3005
R8906 gnd.n5898 gnd.n4590 9.3005
R8907 gnd.n5897 gnd.n4591 9.3005
R8908 gnd.n5894 gnd.n4592 9.3005
R8909 gnd.n5893 gnd.n4593 9.3005
R8910 gnd.n5890 gnd.n4594 9.3005
R8911 gnd.n5889 gnd.n4595 9.3005
R8912 gnd.n5886 gnd.n5885 9.3005
R8913 gnd.n5884 gnd.n4596 9.3005
R8914 gnd.n5917 gnd.n5916 9.3005
R8915 gnd.n5189 gnd.n5188 9.3005
R8916 gnd.n5190 gnd.n4892 9.3005
R8917 gnd.n5192 gnd.n5191 9.3005
R8918 gnd.n4873 gnd.n4872 9.3005
R8919 gnd.n5219 gnd.n5218 9.3005
R8920 gnd.n5220 gnd.n4871 9.3005
R8921 gnd.n5224 gnd.n5221 9.3005
R8922 gnd.n5223 gnd.n5222 9.3005
R8923 gnd.n4847 gnd.n4846 9.3005
R8924 gnd.n5253 gnd.n5252 9.3005
R8925 gnd.n5254 gnd.n4845 9.3005
R8926 gnd.n5261 gnd.n5255 9.3005
R8927 gnd.n5260 gnd.n5256 9.3005
R8928 gnd.n5259 gnd.n5257 9.3005
R8929 gnd.n4814 gnd.n4813 9.3005
R8930 gnd.n5314 gnd.n5313 9.3005
R8931 gnd.n5315 gnd.n4812 9.3005
R8932 gnd.n5319 gnd.n5316 9.3005
R8933 gnd.n5318 gnd.n5317 9.3005
R8934 gnd.n4787 gnd.n4786 9.3005
R8935 gnd.n5354 gnd.n5353 9.3005
R8936 gnd.n5355 gnd.n4785 9.3005
R8937 gnd.n5359 gnd.n5356 9.3005
R8938 gnd.n5358 gnd.n5357 9.3005
R8939 gnd.n4724 gnd.n4723 9.3005
R8940 gnd.n5399 gnd.n5398 9.3005
R8941 gnd.n5400 gnd.n4722 9.3005
R8942 gnd.n5404 gnd.n5401 9.3005
R8943 gnd.n5403 gnd.n5402 9.3005
R8944 gnd.n4696 gnd.n4695 9.3005
R8945 gnd.n5438 gnd.n5437 9.3005
R8946 gnd.n5439 gnd.n4694 9.3005
R8947 gnd.n5446 gnd.n5440 9.3005
R8948 gnd.n5445 gnd.n5441 9.3005
R8949 gnd.n5444 gnd.n5442 9.3005
R8950 gnd.n4665 gnd.n4664 9.3005
R8951 gnd.n5493 gnd.n5492 9.3005
R8952 gnd.n5494 gnd.n4663 9.3005
R8953 gnd.n5499 gnd.n5495 9.3005
R8954 gnd.n5498 gnd.n5497 9.3005
R8955 gnd.n5496 gnd.n809 9.3005
R8956 gnd.n5948 gnd.n810 9.3005
R8957 gnd.n5947 gnd.n811 9.3005
R8958 gnd.n5946 gnd.n812 9.3005
R8959 gnd.n832 gnd.n813 9.3005
R8960 gnd.n833 gnd.n831 9.3005
R8961 gnd.n5934 gnd.n834 9.3005
R8962 gnd.n5933 gnd.n835 9.3005
R8963 gnd.n5932 gnd.n836 9.3005
R8964 gnd.n857 gnd.n837 9.3005
R8965 gnd.n858 gnd.n856 9.3005
R8966 gnd.n5920 gnd.n859 9.3005
R8967 gnd.n5919 gnd.n5918 9.3005
R8968 gnd.n4894 gnd.n4893 9.3005
R8969 gnd.n5134 gnd.n5133 9.3005
R8970 gnd.n5137 gnd.n5129 9.3005
R8971 gnd.n5138 gnd.n5128 9.3005
R8972 gnd.n5141 gnd.n5127 9.3005
R8973 gnd.n5142 gnd.n5126 9.3005
R8974 gnd.n5145 gnd.n5125 9.3005
R8975 gnd.n5146 gnd.n5124 9.3005
R8976 gnd.n5149 gnd.n5123 9.3005
R8977 gnd.n5150 gnd.n5122 9.3005
R8978 gnd.n5153 gnd.n5121 9.3005
R8979 gnd.n5154 gnd.n5120 9.3005
R8980 gnd.n5157 gnd.n5119 9.3005
R8981 gnd.n5159 gnd.n5118 9.3005
R8982 gnd.n5160 gnd.n5117 9.3005
R8983 gnd.n5161 gnd.n5116 9.3005
R8984 gnd.n5162 gnd.n5115 9.3005
R8985 gnd.n5130 gnd.n4911 9.3005
R8986 gnd.n5179 gnd.n4902 9.3005
R8987 gnd.n5181 gnd.n5180 9.3005
R8988 gnd.n4889 gnd.n4884 9.3005
R8989 gnd.n5202 gnd.n4883 9.3005
R8990 gnd.n5205 gnd.n5204 9.3005
R8991 gnd.n5207 gnd.n5206 9.3005
R8992 gnd.n5210 gnd.n4866 9.3005
R8993 gnd.n5208 gnd.n4864 9.3005
R8994 gnd.n5230 gnd.n4862 9.3005
R8995 gnd.n5234 gnd.n5233 9.3005
R8996 gnd.n5232 gnd.n4837 9.3005
R8997 gnd.n5268 gnd.n4836 9.3005
R8998 gnd.n5271 gnd.n5270 9.3005
R8999 gnd.n4834 gnd.n4833 9.3005
R9000 gnd.n5277 gnd.n4831 9.3005
R9001 gnd.n5279 gnd.n5278 9.3005
R9002 gnd.n4805 gnd.n4804 9.3005
R9003 gnd.n5328 gnd.n5327 9.3005
R9004 gnd.n5329 gnd.n4798 9.3005
R9005 gnd.n5337 gnd.n4797 9.3005
R9006 gnd.n5340 gnd.n5339 9.3005
R9007 gnd.n5342 gnd.n5341 9.3005
R9008 gnd.n5345 gnd.n4780 9.3005
R9009 gnd.n5343 gnd.n4778 9.3005
R9010 gnd.n5365 gnd.n4776 9.3005
R9011 gnd.n5367 gnd.n5366 9.3005
R9012 gnd.n4714 gnd.n4713 9.3005
R9013 gnd.n5413 gnd.n5412 9.3005
R9014 gnd.n5414 gnd.n4707 9.3005
R9015 gnd.n5422 gnd.n4706 9.3005
R9016 gnd.n5425 gnd.n5424 9.3005
R9017 gnd.n5427 gnd.n5426 9.3005
R9018 gnd.n5429 gnd.n4689 9.3005
R9019 gnd.n4686 gnd.n4684 9.3005
R9020 gnd.n5454 gnd.n5453 9.3005
R9021 gnd.n4687 gnd.n4670 9.3005
R9022 gnd.n5482 gnd.n4669 9.3005
R9023 gnd.n5486 gnd.n5484 9.3005
R9024 gnd.n5485 gnd.n4654 9.3005
R9025 gnd.n5507 gnd.n4653 9.3005
R9026 gnd.n5511 gnd.n5510 9.3005
R9027 gnd.n4646 gnd.n4645 9.3005
R9028 gnd.n5524 gnd.n5520 9.3005
R9029 gnd.n5523 gnd.n5522 9.3005
R9030 gnd.n4638 gnd.n4637 9.3005
R9031 gnd.n5546 gnd.n4639 9.3005
R9032 gnd.n5548 gnd.n5547 9.3005
R9033 gnd.n5550 gnd.n4636 9.3005
R9034 gnd.n5809 gnd.n5808 9.3005
R9035 gnd.n5811 gnd.n5810 9.3005
R9036 gnd.n5819 gnd.n5812 9.3005
R9037 gnd.n5818 gnd.n5814 9.3005
R9038 gnd.n5817 gnd.n4599 9.3005
R9039 gnd.n5178 gnd.n4905 9.3005
R9040 gnd.n5880 gnd.n4600 9.3005
R9041 gnd.n5879 gnd.n4602 9.3005
R9042 gnd.n5876 gnd.n4603 9.3005
R9043 gnd.n5875 gnd.n4604 9.3005
R9044 gnd.n5872 gnd.n4605 9.3005
R9045 gnd.n5871 gnd.n4606 9.3005
R9046 gnd.n5868 gnd.n4607 9.3005
R9047 gnd.n5867 gnd.n4608 9.3005
R9048 gnd.n5864 gnd.n4609 9.3005
R9049 gnd.n5863 gnd.n4610 9.3005
R9050 gnd.n5860 gnd.n4611 9.3005
R9051 gnd.n5859 gnd.n4612 9.3005
R9052 gnd.n5856 gnd.n4613 9.3005
R9053 gnd.n5855 gnd.n4614 9.3005
R9054 gnd.n5852 gnd.n4615 9.3005
R9055 gnd.n5851 gnd.n4616 9.3005
R9056 gnd.n5848 gnd.n4617 9.3005
R9057 gnd.n5847 gnd.n4618 9.3005
R9058 gnd.n5844 gnd.n4619 9.3005
R9059 gnd.n5843 gnd.n4620 9.3005
R9060 gnd.n5840 gnd.n4621 9.3005
R9061 gnd.n5839 gnd.n4622 9.3005
R9062 gnd.n5836 gnd.n4626 9.3005
R9063 gnd.n5835 gnd.n4627 9.3005
R9064 gnd.n5832 gnd.n4628 9.3005
R9065 gnd.n5831 gnd.n4629 9.3005
R9066 gnd.n5882 gnd.n5881 9.3005
R9067 gnd.n5375 gnd.n5374 9.3005
R9068 gnd.n5376 gnd.n4730 9.3005
R9069 gnd.n5393 gnd.n5377 9.3005
R9070 gnd.n5392 gnd.n5378 9.3005
R9071 gnd.n5391 gnd.n5379 9.3005
R9072 gnd.n5389 gnd.n5380 9.3005
R9073 gnd.n5388 gnd.n5381 9.3005
R9074 gnd.n5386 gnd.n5382 9.3005
R9075 gnd.n5385 gnd.n5383 9.3005
R9076 gnd.n4677 gnd.n4676 9.3005
R9077 gnd.n5461 gnd.n5460 9.3005
R9078 gnd.n5462 gnd.n4675 9.3005
R9079 gnd.n5476 gnd.n5463 9.3005
R9080 gnd.n5475 gnd.n5464 9.3005
R9081 gnd.n5474 gnd.n5465 9.3005
R9082 gnd.n5473 gnd.n5466 9.3005
R9083 gnd.n5471 gnd.n5467 9.3005
R9084 gnd.n5470 gnd.n5468 9.3005
R9085 gnd.n4643 gnd.n4642 9.3005
R9086 gnd.n5530 gnd.n5529 9.3005
R9087 gnd.n5531 gnd.n4641 9.3005
R9088 gnd.n5541 gnd.n5532 9.3005
R9089 gnd.n5540 gnd.n5533 9.3005
R9090 gnd.n5539 gnd.n5534 9.3005
R9091 gnd.n5536 gnd.n5535 9.3005
R9092 gnd.n4632 gnd.n4631 9.3005
R9093 gnd.n5825 gnd.n5824 9.3005
R9094 gnd.n5826 gnd.n4630 9.3005
R9095 gnd.n5828 gnd.n5827 9.3005
R9096 gnd.n5048 gnd.n4942 9.3005
R9097 gnd.n5050 gnd.n5049 9.3005
R9098 gnd.n4932 gnd.n4931 9.3005
R9099 gnd.n5063 gnd.n5062 9.3005
R9100 gnd.n5064 gnd.n4930 9.3005
R9101 gnd.n5066 gnd.n5065 9.3005
R9102 gnd.n4919 gnd.n4918 9.3005
R9103 gnd.n5079 gnd.n5078 9.3005
R9104 gnd.n5080 gnd.n4917 9.3005
R9105 gnd.n5104 gnd.n5081 9.3005
R9106 gnd.n5103 gnd.n5082 9.3005
R9107 gnd.n5102 gnd.n5083 9.3005
R9108 gnd.n5101 gnd.n5084 9.3005
R9109 gnd.n5099 gnd.n5085 9.3005
R9110 gnd.n5098 gnd.n5086 9.3005
R9111 gnd.n5096 gnd.n5087 9.3005
R9112 gnd.n5095 gnd.n5088 9.3005
R9113 gnd.n5093 gnd.n5089 9.3005
R9114 gnd.n5092 gnd.n5090 9.3005
R9115 gnd.n4854 gnd.n4853 9.3005
R9116 gnd.n5242 gnd.n5241 9.3005
R9117 gnd.n5243 gnd.n4852 9.3005
R9118 gnd.n5247 gnd.n5244 9.3005
R9119 gnd.n5246 gnd.n5245 9.3005
R9120 gnd.n4821 gnd.n4820 9.3005
R9121 gnd.n5289 gnd.n5288 9.3005
R9122 gnd.n5290 gnd.n4819 9.3005
R9123 gnd.n5292 gnd.n5291 9.3005
R9124 gnd.n5047 gnd.n5046 9.3005
R9125 gnd.n4987 gnd.n4986 9.3005
R9126 gnd.n4992 gnd.n4984 9.3005
R9127 gnd.n4993 gnd.n4983 9.3005
R9128 gnd.n4995 gnd.n4980 9.3005
R9129 gnd.n4979 gnd.n4977 9.3005
R9130 gnd.n5001 gnd.n4976 9.3005
R9131 gnd.n5002 gnd.n4975 9.3005
R9132 gnd.n5003 gnd.n4974 9.3005
R9133 gnd.n4973 gnd.n4971 9.3005
R9134 gnd.n5009 gnd.n4970 9.3005
R9135 gnd.n5010 gnd.n4969 9.3005
R9136 gnd.n5011 gnd.n4968 9.3005
R9137 gnd.n4967 gnd.n4965 9.3005
R9138 gnd.n5017 gnd.n4964 9.3005
R9139 gnd.n5018 gnd.n4963 9.3005
R9140 gnd.n5019 gnd.n4962 9.3005
R9141 gnd.n4961 gnd.n4959 9.3005
R9142 gnd.n5025 gnd.n4958 9.3005
R9143 gnd.n5026 gnd.n4957 9.3005
R9144 gnd.n5027 gnd.n4956 9.3005
R9145 gnd.n4955 gnd.n4953 9.3005
R9146 gnd.n5032 gnd.n4952 9.3005
R9147 gnd.n5033 gnd.n4951 9.3005
R9148 gnd.n4950 gnd.n4948 9.3005
R9149 gnd.n5038 gnd.n4947 9.3005
R9150 gnd.n5040 gnd.n5039 9.3005
R9151 gnd.n4985 gnd.n4943 9.3005
R9152 gnd.n4938 gnd.n4937 9.3005
R9153 gnd.n5055 gnd.n5054 9.3005
R9154 gnd.n5056 gnd.n4936 9.3005
R9155 gnd.n5058 gnd.n5057 9.3005
R9156 gnd.n4926 gnd.n4925 9.3005
R9157 gnd.n5071 gnd.n5070 9.3005
R9158 gnd.n5072 gnd.n4924 9.3005
R9159 gnd.n5074 gnd.n5073 9.3005
R9160 gnd.n4913 gnd.n4912 9.3005
R9161 gnd.n5169 gnd.n5168 9.3005
R9162 gnd.n5171 gnd.n4910 9.3005
R9163 gnd.n5173 gnd.n5172 9.3005
R9164 gnd.n4904 gnd.n4901 9.3005
R9165 gnd.n5183 gnd.n5182 9.3005
R9166 gnd.n4903 gnd.n4885 9.3005
R9167 gnd.n5201 gnd.n5200 9.3005
R9168 gnd.n5203 gnd.n4881 9.3005
R9169 gnd.n5213 gnd.n4882 9.3005
R9170 gnd.n5212 gnd.n5211 9.3005
R9171 gnd.n5209 gnd.n4860 9.3005
R9172 gnd.n5237 gnd.n4861 9.3005
R9173 gnd.n5236 gnd.n5235 9.3005
R9174 gnd.n4863 gnd.n4838 9.3005
R9175 gnd.n5267 gnd.n5266 9.3005
R9176 gnd.n5269 gnd.n4828 9.3005
R9177 gnd.n5284 gnd.n4829 9.3005
R9178 gnd.n5283 gnd.n4830 9.3005
R9179 gnd.n5282 gnd.n5280 9.3005
R9180 gnd.n4832 gnd.n4806 9.3005
R9181 gnd.n5325 gnd.n5324 9.3005
R9182 gnd.n5326 gnd.n4799 9.3005
R9183 gnd.n5336 gnd.n5335 9.3005
R9184 gnd.n5338 gnd.n4795 9.3005
R9185 gnd.n5348 gnd.n4796 9.3005
R9186 gnd.n5347 gnd.n5346 9.3005
R9187 gnd.n5344 gnd.n4774 9.3005
R9188 gnd.n5370 gnd.n4775 9.3005
R9189 gnd.n5369 gnd.n5368 9.3005
R9190 gnd.n4777 gnd.n4715 9.3005
R9191 gnd.n5410 gnd.n5409 9.3005
R9192 gnd.n5411 gnd.n4708 9.3005
R9193 gnd.n5421 gnd.n5420 9.3005
R9194 gnd.n5423 gnd.n4704 9.3005
R9195 gnd.n5432 gnd.n4705 9.3005
R9196 gnd.n5431 gnd.n5430 9.3005
R9197 gnd.n5428 gnd.n4683 9.3005
R9198 gnd.n5456 gnd.n5455 9.3005
R9199 gnd.n4685 gnd.n4671 9.3005
R9200 gnd.n5481 gnd.n5480 9.3005
R9201 gnd.n5483 gnd.n4655 9.3005
R9202 gnd.n5504 gnd.n4656 9.3005
R9203 gnd.n5506 gnd.n5505 9.3005
R9204 gnd.n5508 gnd.n4649 9.3005
R9205 gnd.n5509 gnd.n4647 9.3005
R9206 gnd.n5519 gnd.n5518 9.3005
R9207 gnd.n5521 gnd.n820 9.3005
R9208 gnd.n5941 gnd.n821 9.3005
R9209 gnd.n5940 gnd.n822 9.3005
R9210 gnd.n5939 gnd.n823 9.3005
R9211 gnd.n5549 gnd.n824 9.3005
R9212 gnd.n5807 gnd.n845 9.3005
R9213 gnd.n5927 gnd.n846 9.3005
R9214 gnd.n5926 gnd.n847 9.3005
R9215 gnd.n5925 gnd.n848 9.3005
R9216 gnd.n5813 gnd.n849 9.3005
R9217 gnd.n5042 gnd.n5041 9.3005
R9218 gnd.n635 gnd.n634 9.3005
R9219 gnd.n6124 gnd.n6123 9.3005
R9220 gnd.n6125 gnd.n633 9.3005
R9221 gnd.n6127 gnd.n6126 9.3005
R9222 gnd.n629 gnd.n628 9.3005
R9223 gnd.n6134 gnd.n6133 9.3005
R9224 gnd.n6135 gnd.n627 9.3005
R9225 gnd.n6137 gnd.n6136 9.3005
R9226 gnd.n623 gnd.n622 9.3005
R9227 gnd.n6144 gnd.n6143 9.3005
R9228 gnd.n6145 gnd.n621 9.3005
R9229 gnd.n6147 gnd.n6146 9.3005
R9230 gnd.n617 gnd.n616 9.3005
R9231 gnd.n6154 gnd.n6153 9.3005
R9232 gnd.n6155 gnd.n615 9.3005
R9233 gnd.n6157 gnd.n6156 9.3005
R9234 gnd.n611 gnd.n610 9.3005
R9235 gnd.n6164 gnd.n6163 9.3005
R9236 gnd.n6165 gnd.n609 9.3005
R9237 gnd.n6167 gnd.n6166 9.3005
R9238 gnd.n605 gnd.n604 9.3005
R9239 gnd.n6174 gnd.n6173 9.3005
R9240 gnd.n6175 gnd.n603 9.3005
R9241 gnd.n6177 gnd.n6176 9.3005
R9242 gnd.n599 gnd.n598 9.3005
R9243 gnd.n6184 gnd.n6183 9.3005
R9244 gnd.n6185 gnd.n597 9.3005
R9245 gnd.n6187 gnd.n6186 9.3005
R9246 gnd.n593 gnd.n592 9.3005
R9247 gnd.n6194 gnd.n6193 9.3005
R9248 gnd.n6195 gnd.n591 9.3005
R9249 gnd.n6197 gnd.n6196 9.3005
R9250 gnd.n587 gnd.n586 9.3005
R9251 gnd.n6204 gnd.n6203 9.3005
R9252 gnd.n6205 gnd.n585 9.3005
R9253 gnd.n6207 gnd.n6206 9.3005
R9254 gnd.n581 gnd.n580 9.3005
R9255 gnd.n6214 gnd.n6213 9.3005
R9256 gnd.n6215 gnd.n579 9.3005
R9257 gnd.n6217 gnd.n6216 9.3005
R9258 gnd.n575 gnd.n574 9.3005
R9259 gnd.n6224 gnd.n6223 9.3005
R9260 gnd.n6225 gnd.n573 9.3005
R9261 gnd.n6227 gnd.n6226 9.3005
R9262 gnd.n569 gnd.n568 9.3005
R9263 gnd.n6234 gnd.n6233 9.3005
R9264 gnd.n6235 gnd.n567 9.3005
R9265 gnd.n6237 gnd.n6236 9.3005
R9266 gnd.n563 gnd.n562 9.3005
R9267 gnd.n6244 gnd.n6243 9.3005
R9268 gnd.n6245 gnd.n561 9.3005
R9269 gnd.n6247 gnd.n6246 9.3005
R9270 gnd.n557 gnd.n556 9.3005
R9271 gnd.n6254 gnd.n6253 9.3005
R9272 gnd.n6255 gnd.n555 9.3005
R9273 gnd.n6257 gnd.n6256 9.3005
R9274 gnd.n551 gnd.n550 9.3005
R9275 gnd.n6264 gnd.n6263 9.3005
R9276 gnd.n6265 gnd.n549 9.3005
R9277 gnd.n6267 gnd.n6266 9.3005
R9278 gnd.n545 gnd.n544 9.3005
R9279 gnd.n6274 gnd.n6273 9.3005
R9280 gnd.n6275 gnd.n543 9.3005
R9281 gnd.n6277 gnd.n6276 9.3005
R9282 gnd.n539 gnd.n538 9.3005
R9283 gnd.n6284 gnd.n6283 9.3005
R9284 gnd.n6285 gnd.n537 9.3005
R9285 gnd.n6287 gnd.n6286 9.3005
R9286 gnd.n533 gnd.n532 9.3005
R9287 gnd.n6294 gnd.n6293 9.3005
R9288 gnd.n6295 gnd.n531 9.3005
R9289 gnd.n6297 gnd.n6296 9.3005
R9290 gnd.n527 gnd.n526 9.3005
R9291 gnd.n6304 gnd.n6303 9.3005
R9292 gnd.n6305 gnd.n525 9.3005
R9293 gnd.n6307 gnd.n6306 9.3005
R9294 gnd.n521 gnd.n520 9.3005
R9295 gnd.n6314 gnd.n6313 9.3005
R9296 gnd.n6315 gnd.n519 9.3005
R9297 gnd.n6317 gnd.n6316 9.3005
R9298 gnd.n515 gnd.n514 9.3005
R9299 gnd.n6324 gnd.n6323 9.3005
R9300 gnd.n6325 gnd.n513 9.3005
R9301 gnd.n6327 gnd.n6326 9.3005
R9302 gnd.n509 gnd.n508 9.3005
R9303 gnd.n6334 gnd.n6333 9.3005
R9304 gnd.n6335 gnd.n507 9.3005
R9305 gnd.n6337 gnd.n6336 9.3005
R9306 gnd.n503 gnd.n502 9.3005
R9307 gnd.n6344 gnd.n6343 9.3005
R9308 gnd.n6345 gnd.n501 9.3005
R9309 gnd.n6347 gnd.n6346 9.3005
R9310 gnd.n497 gnd.n496 9.3005
R9311 gnd.n6354 gnd.n6353 9.3005
R9312 gnd.n6355 gnd.n495 9.3005
R9313 gnd.n6357 gnd.n6356 9.3005
R9314 gnd.n491 gnd.n490 9.3005
R9315 gnd.n6364 gnd.n6363 9.3005
R9316 gnd.n6365 gnd.n489 9.3005
R9317 gnd.n6367 gnd.n6366 9.3005
R9318 gnd.n485 gnd.n484 9.3005
R9319 gnd.n6374 gnd.n6373 9.3005
R9320 gnd.n6375 gnd.n483 9.3005
R9321 gnd.n6377 gnd.n6376 9.3005
R9322 gnd.n479 gnd.n478 9.3005
R9323 gnd.n6384 gnd.n6383 9.3005
R9324 gnd.n6385 gnd.n477 9.3005
R9325 gnd.n6387 gnd.n6386 9.3005
R9326 gnd.n473 gnd.n472 9.3005
R9327 gnd.n6394 gnd.n6393 9.3005
R9328 gnd.n6395 gnd.n471 9.3005
R9329 gnd.n6397 gnd.n6396 9.3005
R9330 gnd.n467 gnd.n466 9.3005
R9331 gnd.n6404 gnd.n6403 9.3005
R9332 gnd.n6405 gnd.n465 9.3005
R9333 gnd.n6407 gnd.n6406 9.3005
R9334 gnd.n461 gnd.n460 9.3005
R9335 gnd.n6414 gnd.n6413 9.3005
R9336 gnd.n6415 gnd.n459 9.3005
R9337 gnd.n6417 gnd.n6416 9.3005
R9338 gnd.n455 gnd.n454 9.3005
R9339 gnd.n6424 gnd.n6423 9.3005
R9340 gnd.n6425 gnd.n453 9.3005
R9341 gnd.n6427 gnd.n6426 9.3005
R9342 gnd.n449 gnd.n448 9.3005
R9343 gnd.n6434 gnd.n6433 9.3005
R9344 gnd.n6435 gnd.n447 9.3005
R9345 gnd.n6437 gnd.n6436 9.3005
R9346 gnd.n443 gnd.n442 9.3005
R9347 gnd.n6444 gnd.n6443 9.3005
R9348 gnd.n6445 gnd.n441 9.3005
R9349 gnd.n6447 gnd.n6446 9.3005
R9350 gnd.n437 gnd.n436 9.3005
R9351 gnd.n6454 gnd.n6453 9.3005
R9352 gnd.n6455 gnd.n435 9.3005
R9353 gnd.n6457 gnd.n6456 9.3005
R9354 gnd.n431 gnd.n430 9.3005
R9355 gnd.n6464 gnd.n6463 9.3005
R9356 gnd.n6465 gnd.n429 9.3005
R9357 gnd.n6467 gnd.n6466 9.3005
R9358 gnd.n425 gnd.n424 9.3005
R9359 gnd.n6474 gnd.n6473 9.3005
R9360 gnd.n6475 gnd.n423 9.3005
R9361 gnd.n6477 gnd.n6476 9.3005
R9362 gnd.n419 gnd.n418 9.3005
R9363 gnd.n6484 gnd.n6483 9.3005
R9364 gnd.n6485 gnd.n417 9.3005
R9365 gnd.n6487 gnd.n6486 9.3005
R9366 gnd.n413 gnd.n412 9.3005
R9367 gnd.n6494 gnd.n6493 9.3005
R9368 gnd.n6495 gnd.n411 9.3005
R9369 gnd.n6498 gnd.n6497 9.3005
R9370 gnd.n6496 gnd.n407 9.3005
R9371 gnd.n6504 gnd.n406 9.3005
R9372 gnd.n6506 gnd.n6505 9.3005
R9373 gnd.n402 gnd.n401 9.3005
R9374 gnd.n6515 gnd.n6514 9.3005
R9375 gnd.n6516 gnd.n400 9.3005
R9376 gnd.n6518 gnd.n6517 9.3005
R9377 gnd.n396 gnd.n395 9.3005
R9378 gnd.n6525 gnd.n6524 9.3005
R9379 gnd.n6526 gnd.n394 9.3005
R9380 gnd.n6528 gnd.n6527 9.3005
R9381 gnd.n390 gnd.n389 9.3005
R9382 gnd.n6535 gnd.n6534 9.3005
R9383 gnd.n6536 gnd.n388 9.3005
R9384 gnd.n6538 gnd.n6537 9.3005
R9385 gnd.n384 gnd.n383 9.3005
R9386 gnd.n6545 gnd.n6544 9.3005
R9387 gnd.n6546 gnd.n382 9.3005
R9388 gnd.n6548 gnd.n6547 9.3005
R9389 gnd.n378 gnd.n377 9.3005
R9390 gnd.n6555 gnd.n6554 9.3005
R9391 gnd.n6556 gnd.n376 9.3005
R9392 gnd.n6558 gnd.n6557 9.3005
R9393 gnd.n372 gnd.n371 9.3005
R9394 gnd.n6565 gnd.n6564 9.3005
R9395 gnd.n6566 gnd.n370 9.3005
R9396 gnd.n6568 gnd.n6567 9.3005
R9397 gnd.n366 gnd.n365 9.3005
R9398 gnd.n6575 gnd.n6574 9.3005
R9399 gnd.n6576 gnd.n364 9.3005
R9400 gnd.n6578 gnd.n6577 9.3005
R9401 gnd.n360 gnd.n359 9.3005
R9402 gnd.n6585 gnd.n6584 9.3005
R9403 gnd.n6586 gnd.n358 9.3005
R9404 gnd.n6588 gnd.n6587 9.3005
R9405 gnd.n354 gnd.n353 9.3005
R9406 gnd.n6595 gnd.n6594 9.3005
R9407 gnd.n6596 gnd.n352 9.3005
R9408 gnd.n6598 gnd.n6597 9.3005
R9409 gnd.n348 gnd.n347 9.3005
R9410 gnd.n6605 gnd.n6604 9.3005
R9411 gnd.n6606 gnd.n346 9.3005
R9412 gnd.n6608 gnd.n6607 9.3005
R9413 gnd.n342 gnd.n341 9.3005
R9414 gnd.n6615 gnd.n6614 9.3005
R9415 gnd.n6616 gnd.n340 9.3005
R9416 gnd.n6618 gnd.n6617 9.3005
R9417 gnd.n336 gnd.n335 9.3005
R9418 gnd.n6625 gnd.n6624 9.3005
R9419 gnd.n6626 gnd.n334 9.3005
R9420 gnd.n6628 gnd.n6627 9.3005
R9421 gnd.n330 gnd.n329 9.3005
R9422 gnd.n6635 gnd.n6634 9.3005
R9423 gnd.n6636 gnd.n328 9.3005
R9424 gnd.n6638 gnd.n6637 9.3005
R9425 gnd.n324 gnd.n323 9.3005
R9426 gnd.n6645 gnd.n6644 9.3005
R9427 gnd.n6646 gnd.n322 9.3005
R9428 gnd.n6648 gnd.n6647 9.3005
R9429 gnd.n318 gnd.n317 9.3005
R9430 gnd.n6655 gnd.n6654 9.3005
R9431 gnd.n6656 gnd.n316 9.3005
R9432 gnd.n6658 gnd.n6657 9.3005
R9433 gnd.n312 gnd.n311 9.3005
R9434 gnd.n6665 gnd.n6664 9.3005
R9435 gnd.n6666 gnd.n310 9.3005
R9436 gnd.n6668 gnd.n6667 9.3005
R9437 gnd.n306 gnd.n305 9.3005
R9438 gnd.n6675 gnd.n6674 9.3005
R9439 gnd.n6676 gnd.n304 9.3005
R9440 gnd.n6678 gnd.n6677 9.3005
R9441 gnd.n300 gnd.n299 9.3005
R9442 gnd.n6685 gnd.n6684 9.3005
R9443 gnd.n6686 gnd.n298 9.3005
R9444 gnd.n6688 gnd.n6687 9.3005
R9445 gnd.n294 gnd.n293 9.3005
R9446 gnd.n6695 gnd.n6694 9.3005
R9447 gnd.n6696 gnd.n292 9.3005
R9448 gnd.n6698 gnd.n6697 9.3005
R9449 gnd.n288 gnd.n287 9.3005
R9450 gnd.n6705 gnd.n6704 9.3005
R9451 gnd.n6706 gnd.n286 9.3005
R9452 gnd.n6708 gnd.n6707 9.3005
R9453 gnd.n282 gnd.n281 9.3005
R9454 gnd.n6716 gnd.n6715 9.3005
R9455 gnd.n6717 gnd.n280 9.3005
R9456 gnd.n6719 gnd.n6718 9.3005
R9457 gnd.n6508 gnd.n6507 9.3005
R9458 gnd.n6956 gnd.n89 9.3005
R9459 gnd.n6955 gnd.n91 9.3005
R9460 gnd.n96 gnd.n92 9.3005
R9461 gnd.n6950 gnd.n97 9.3005
R9462 gnd.n6949 gnd.n98 9.3005
R9463 gnd.n6948 gnd.n99 9.3005
R9464 gnd.n103 gnd.n100 9.3005
R9465 gnd.n6943 gnd.n104 9.3005
R9466 gnd.n6942 gnd.n105 9.3005
R9467 gnd.n6941 gnd.n106 9.3005
R9468 gnd.n110 gnd.n107 9.3005
R9469 gnd.n6936 gnd.n111 9.3005
R9470 gnd.n6935 gnd.n112 9.3005
R9471 gnd.n6934 gnd.n113 9.3005
R9472 gnd.n117 gnd.n114 9.3005
R9473 gnd.n6929 gnd.n118 9.3005
R9474 gnd.n6928 gnd.n119 9.3005
R9475 gnd.n6924 gnd.n120 9.3005
R9476 gnd.n124 gnd.n121 9.3005
R9477 gnd.n6919 gnd.n125 9.3005
R9478 gnd.n6918 gnd.n126 9.3005
R9479 gnd.n6917 gnd.n127 9.3005
R9480 gnd.n131 gnd.n128 9.3005
R9481 gnd.n6912 gnd.n132 9.3005
R9482 gnd.n6911 gnd.n133 9.3005
R9483 gnd.n6910 gnd.n134 9.3005
R9484 gnd.n138 gnd.n135 9.3005
R9485 gnd.n6905 gnd.n139 9.3005
R9486 gnd.n6904 gnd.n140 9.3005
R9487 gnd.n6903 gnd.n141 9.3005
R9488 gnd.n145 gnd.n142 9.3005
R9489 gnd.n6898 gnd.n146 9.3005
R9490 gnd.n6897 gnd.n147 9.3005
R9491 gnd.n6896 gnd.n148 9.3005
R9492 gnd.n152 gnd.n149 9.3005
R9493 gnd.n6891 gnd.n153 9.3005
R9494 gnd.n6890 gnd.n6889 9.3005
R9495 gnd.n6888 gnd.n156 9.3005
R9496 gnd.n6958 gnd.n6957 9.3005
R9497 gnd.n3918 gnd.n3917 9.3005
R9498 gnd.n3954 gnd.n3919 9.3005
R9499 gnd.n3953 gnd.n3920 9.3005
R9500 gnd.n3952 gnd.n3921 9.3005
R9501 gnd.n3950 gnd.n3922 9.3005
R9502 gnd.n3949 gnd.n3923 9.3005
R9503 gnd.n3948 gnd.n3924 9.3005
R9504 gnd.n3945 gnd.n3925 9.3005
R9505 gnd.n3944 gnd.n3926 9.3005
R9506 gnd.n3940 gnd.n3927 9.3005
R9507 gnd.n3939 gnd.n3928 9.3005
R9508 gnd.n3938 gnd.n3929 9.3005
R9509 gnd.n3935 gnd.n3930 9.3005
R9510 gnd.n3934 gnd.n3932 9.3005
R9511 gnd.n3931 gnd.n1422 9.3005
R9512 gnd.n4075 gnd.n1423 9.3005
R9513 gnd.n4074 gnd.n1424 9.3005
R9514 gnd.n4073 gnd.n1425 9.3005
R9515 gnd.n1431 gnd.n1426 9.3005
R9516 gnd.n1430 gnd.n1427 9.3005
R9517 gnd.n1428 gnd.n1395 9.3005
R9518 gnd.n1394 gnd.n234 9.3005
R9519 gnd.n6737 gnd.n235 9.3005
R9520 gnd.n6736 gnd.n236 9.3005
R9521 gnd.n6735 gnd.n237 9.3005
R9522 gnd.n6731 gnd.n238 9.3005
R9523 gnd.n6730 gnd.n239 9.3005
R9524 gnd.n271 gnd.n240 9.3005
R9525 gnd.n270 gnd.n241 9.3005
R9526 gnd.n266 gnd.n242 9.3005
R9527 gnd.n265 gnd.n243 9.3005
R9528 gnd.n263 gnd.n244 9.3005
R9529 gnd.n262 gnd.n245 9.3005
R9530 gnd.n260 gnd.n246 9.3005
R9531 gnd.n259 gnd.n247 9.3005
R9532 gnd.n257 gnd.n248 9.3005
R9533 gnd.n256 gnd.n249 9.3005
R9534 gnd.n254 gnd.n250 9.3005
R9535 gnd.n253 gnd.n252 9.3005
R9536 gnd.n251 gnd.n160 9.3005
R9537 gnd.n6885 gnd.n159 9.3005
R9538 gnd.n6887 gnd.n6886 9.3005
R9539 gnd.n1361 gnd.n1359 9.3005
R9540 gnd.n4160 gnd.n4159 9.3005
R9541 gnd.n4161 gnd.n1353 9.3005
R9542 gnd.n4164 gnd.n1352 9.3005
R9543 gnd.n4165 gnd.n1351 9.3005
R9544 gnd.n4168 gnd.n1350 9.3005
R9545 gnd.n4169 gnd.n1349 9.3005
R9546 gnd.n4172 gnd.n1348 9.3005
R9547 gnd.n4173 gnd.n1347 9.3005
R9548 gnd.n4176 gnd.n1346 9.3005
R9549 gnd.n4177 gnd.n1345 9.3005
R9550 gnd.n4180 gnd.n1344 9.3005
R9551 gnd.n4181 gnd.n1343 9.3005
R9552 gnd.n4184 gnd.n1342 9.3005
R9553 gnd.n4185 gnd.n1341 9.3005
R9554 gnd.n4188 gnd.n1340 9.3005
R9555 gnd.n4189 gnd.n1339 9.3005
R9556 gnd.n4192 gnd.n1338 9.3005
R9557 gnd.n4193 gnd.n1337 9.3005
R9558 gnd.n4196 gnd.n1336 9.3005
R9559 gnd.n4198 gnd.n1330 9.3005
R9560 gnd.n4201 gnd.n1329 9.3005
R9561 gnd.n4202 gnd.n1328 9.3005
R9562 gnd.n4205 gnd.n1327 9.3005
R9563 gnd.n4206 gnd.n1326 9.3005
R9564 gnd.n4209 gnd.n1325 9.3005
R9565 gnd.n4210 gnd.n1324 9.3005
R9566 gnd.n4213 gnd.n1323 9.3005
R9567 gnd.n4214 gnd.n1322 9.3005
R9568 gnd.n4217 gnd.n1321 9.3005
R9569 gnd.n4218 gnd.n1320 9.3005
R9570 gnd.n4221 gnd.n1319 9.3005
R9571 gnd.n4223 gnd.n1318 9.3005
R9572 gnd.n4224 gnd.n1317 9.3005
R9573 gnd.n4225 gnd.n1316 9.3005
R9574 gnd.n4226 gnd.n1315 9.3005
R9575 gnd.n4158 gnd.n1358 9.3005
R9576 gnd.n4157 gnd.n4156 9.3005
R9577 gnd.n3977 gnd.n3976 9.3005
R9578 gnd.n3978 gnd.n1500 9.3005
R9579 gnd.n3982 gnd.n3979 9.3005
R9580 gnd.n3981 gnd.n3980 9.3005
R9581 gnd.n1476 gnd.n1475 9.3005
R9582 gnd.n4009 gnd.n4008 9.3005
R9583 gnd.n4010 gnd.n1474 9.3005
R9584 gnd.n4014 gnd.n4011 9.3005
R9585 gnd.n4013 gnd.n4012 9.3005
R9586 gnd.n1451 gnd.n1450 9.3005
R9587 gnd.n4043 gnd.n4042 9.3005
R9588 gnd.n4044 gnd.n1449 9.3005
R9589 gnd.n4049 gnd.n4045 9.3005
R9590 gnd.n4048 gnd.n4046 9.3005
R9591 gnd.n4047 gnd.n212 9.3005
R9592 gnd.n6756 gnd.n211 9.3005
R9593 gnd.n6758 gnd.n6757 9.3005
R9594 gnd.n199 gnd.n198 9.3005
R9595 gnd.n6771 gnd.n6770 9.3005
R9596 gnd.n6772 gnd.n197 9.3005
R9597 gnd.n6774 gnd.n6773 9.3005
R9598 gnd.n183 gnd.n182 9.3005
R9599 gnd.n6787 gnd.n6786 9.3005
R9600 gnd.n6788 gnd.n181 9.3005
R9601 gnd.n6790 gnd.n6789 9.3005
R9602 gnd.n167 gnd.n166 9.3005
R9603 gnd.n6877 gnd.n6876 9.3005
R9604 gnd.n6878 gnd.n165 9.3005
R9605 gnd.n6880 gnd.n6879 9.3005
R9606 gnd.n88 gnd.n87 9.3005
R9607 gnd.n6960 gnd.n6959 9.3005
R9608 gnd.n1502 gnd.n1501 9.3005
R9609 gnd.n6755 gnd.n6754 9.3005
R9610 gnd.n2290 gnd.n2230 9.3005
R9611 gnd.n2289 gnd.n2236 9.3005
R9612 gnd.n2239 gnd.n2237 9.3005
R9613 gnd.n2285 gnd.n2240 9.3005
R9614 gnd.n2284 gnd.n2241 9.3005
R9615 gnd.n2283 gnd.n2242 9.3005
R9616 gnd.n2245 gnd.n2243 9.3005
R9617 gnd.n2279 gnd.n2246 9.3005
R9618 gnd.n2278 gnd.n2247 9.3005
R9619 gnd.n2277 gnd.n2248 9.3005
R9620 gnd.n2251 gnd.n2249 9.3005
R9621 gnd.n2273 gnd.n2252 9.3005
R9622 gnd.n2272 gnd.n2253 9.3005
R9623 gnd.n2271 gnd.n2254 9.3005
R9624 gnd.n2257 gnd.n2255 9.3005
R9625 gnd.n2267 gnd.n2258 9.3005
R9626 gnd.n2266 gnd.n2259 9.3005
R9627 gnd.n2265 gnd.n2260 9.3005
R9628 gnd.n2262 gnd.n2261 9.3005
R9629 gnd.n1983 gnd.n1982 9.3005
R9630 gnd.n2903 gnd.n2902 9.3005
R9631 gnd.n2904 gnd.n1981 9.3005
R9632 gnd.n2906 gnd.n2905 9.3005
R9633 gnd.n1969 gnd.n1968 9.3005
R9634 gnd.n2919 gnd.n2918 9.3005
R9635 gnd.n2920 gnd.n1967 9.3005
R9636 gnd.n2924 gnd.n2921 9.3005
R9637 gnd.n2923 gnd.n2922 9.3005
R9638 gnd.n1937 gnd.n1936 9.3005
R9639 gnd.n3043 gnd.n3042 9.3005
R9640 gnd.n3044 gnd.n1935 9.3005
R9641 gnd.n3046 gnd.n3045 9.3005
R9642 gnd.n1923 gnd.n1922 9.3005
R9643 gnd.n3059 gnd.n3058 9.3005
R9644 gnd.n3060 gnd.n1921 9.3005
R9645 gnd.n3062 gnd.n3061 9.3005
R9646 gnd.n1908 gnd.n1907 9.3005
R9647 gnd.n3075 gnd.n3074 9.3005
R9648 gnd.n3076 gnd.n1906 9.3005
R9649 gnd.n3078 gnd.n3077 9.3005
R9650 gnd.n1894 gnd.n1893 9.3005
R9651 gnd.n3090 gnd.n3089 9.3005
R9652 gnd.n3091 gnd.n1892 9.3005
R9653 gnd.n3095 gnd.n3092 9.3005
R9654 gnd.n3094 gnd.n3093 9.3005
R9655 gnd.n1862 gnd.n1861 9.3005
R9656 gnd.n3216 gnd.n3215 9.3005
R9657 gnd.n3217 gnd.n1860 9.3005
R9658 gnd.n3219 gnd.n3218 9.3005
R9659 gnd.n1848 gnd.n1847 9.3005
R9660 gnd.n3232 gnd.n3231 9.3005
R9661 gnd.n3233 gnd.n1846 9.3005
R9662 gnd.n3235 gnd.n3234 9.3005
R9663 gnd.n1835 gnd.n1834 9.3005
R9664 gnd.n3248 gnd.n3247 9.3005
R9665 gnd.n3249 gnd.n1833 9.3005
R9666 gnd.n3251 gnd.n3250 9.3005
R9667 gnd.n1824 gnd.n1823 9.3005
R9668 gnd.n3264 gnd.n3263 9.3005
R9669 gnd.n3265 gnd.n1822 9.3005
R9670 gnd.n3269 gnd.n3266 9.3005
R9671 gnd.n3268 gnd.n3267 9.3005
R9672 gnd.n1791 gnd.n1790 9.3005
R9673 gnd.n3387 gnd.n3386 9.3005
R9674 gnd.n3388 gnd.n1789 9.3005
R9675 gnd.n3390 gnd.n3389 9.3005
R9676 gnd.n1776 gnd.n1775 9.3005
R9677 gnd.n3403 gnd.n3402 9.3005
R9678 gnd.n3404 gnd.n1774 9.3005
R9679 gnd.n3406 gnd.n3405 9.3005
R9680 gnd.n1761 gnd.n1760 9.3005
R9681 gnd.n3419 gnd.n3418 9.3005
R9682 gnd.n3420 gnd.n1759 9.3005
R9683 gnd.n3422 gnd.n3421 9.3005
R9684 gnd.n1748 gnd.n1747 9.3005
R9685 gnd.n3435 gnd.n3434 9.3005
R9686 gnd.n3436 gnd.n1746 9.3005
R9687 gnd.n3440 gnd.n3437 9.3005
R9688 gnd.n3439 gnd.n3438 9.3005
R9689 gnd.n1716 gnd.n1715 9.3005
R9690 gnd.n3793 gnd.n3792 9.3005
R9691 gnd.n3794 gnd.n1714 9.3005
R9692 gnd.n3796 gnd.n3795 9.3005
R9693 gnd.n1703 gnd.n1702 9.3005
R9694 gnd.n3809 gnd.n3808 9.3005
R9695 gnd.n3810 gnd.n1701 9.3005
R9696 gnd.n3812 gnd.n3811 9.3005
R9697 gnd.n1689 gnd.n1688 9.3005
R9698 gnd.n3825 gnd.n3824 9.3005
R9699 gnd.n3826 gnd.n1687 9.3005
R9700 gnd.n3828 gnd.n3827 9.3005
R9701 gnd.n1676 gnd.n1675 9.3005
R9702 gnd.n3841 gnd.n3840 9.3005
R9703 gnd.n3842 gnd.n1674 9.3005
R9704 gnd.n3844 gnd.n3843 9.3005
R9705 gnd.n1662 gnd.n1661 9.3005
R9706 gnd.n3857 gnd.n3856 9.3005
R9707 gnd.n3858 gnd.n1660 9.3005
R9708 gnd.n3860 gnd.n3859 9.3005
R9709 gnd.n1648 gnd.n1647 9.3005
R9710 gnd.n3875 gnd.n3874 9.3005
R9711 gnd.n3876 gnd.n1646 9.3005
R9712 gnd.n3881 gnd.n3877 9.3005
R9713 gnd.n3880 gnd.n3879 9.3005
R9714 gnd.n3878 gnd.n1277 9.3005
R9715 gnd.n4235 gnd.n1278 9.3005
R9716 gnd.n4234 gnd.n1279 9.3005
R9717 gnd.n4233 gnd.n1280 9.3005
R9718 gnd.n3960 gnd.n1281 9.3005
R9719 gnd.n3962 gnd.n3961 9.3005
R9720 gnd.n3966 gnd.n3965 9.3005
R9721 gnd.n3967 gnd.n3959 9.3005
R9722 gnd.n3971 gnd.n3968 9.3005
R9723 gnd.n3970 gnd.n3969 9.3005
R9724 gnd.n1485 gnd.n1484 9.3005
R9725 gnd.n3998 gnd.n3997 9.3005
R9726 gnd.n3999 gnd.n1483 9.3005
R9727 gnd.n4003 gnd.n4000 9.3005
R9728 gnd.n4002 gnd.n4001 9.3005
R9729 gnd.n1460 gnd.n1459 9.3005
R9730 gnd.n4029 gnd.n4028 9.3005
R9731 gnd.n4030 gnd.n1458 9.3005
R9732 gnd.n4037 gnd.n4031 9.3005
R9733 gnd.n4036 gnd.n4032 9.3005
R9734 gnd.n4035 gnd.n4034 9.3005
R9735 gnd.n4033 gnd.n1434 9.3005
R9736 gnd.n4063 gnd.n1435 9.3005
R9737 gnd.n275 gnd.n274 9.3005
R9738 gnd.n6725 gnd.n276 9.3005
R9739 gnd.n6724 gnd.n277 9.3005
R9740 gnd.n6723 gnd.n278 9.3005
R9741 gnd.n2494 gnd.n2493 9.3005
R9742 gnd.n2355 gnd.n2354 9.3005
R9743 gnd.n2439 gnd.n2438 9.3005
R9744 gnd.n2440 gnd.n2353 9.3005
R9745 gnd.n2443 gnd.n2441 9.3005
R9746 gnd.n2444 gnd.n2352 9.3005
R9747 gnd.n2447 gnd.n2446 9.3005
R9748 gnd.n2448 gnd.n2351 9.3005
R9749 gnd.n2451 gnd.n2449 9.3005
R9750 gnd.n2452 gnd.n2350 9.3005
R9751 gnd.n2455 gnd.n2454 9.3005
R9752 gnd.n2456 gnd.n2349 9.3005
R9753 gnd.n2459 gnd.n2458 9.3005
R9754 gnd.n2457 gnd.n2330 9.3005
R9755 gnd.n2473 gnd.n2329 9.3005
R9756 gnd.n2475 gnd.n2474 9.3005
R9757 gnd.n2476 gnd.n2328 9.3005
R9758 gnd.n2478 gnd.n2477 9.3005
R9759 gnd.n2221 gnd.n2220 9.3005
R9760 gnd.n2491 gnd.n2490 9.3005
R9761 gnd.n2492 gnd.n2219 9.3005
R9762 gnd.n2381 gnd.n2380 9.3005
R9763 gnd.n2386 gnd.n2385 9.3005
R9764 gnd.n2389 gnd.n2375 9.3005
R9765 gnd.n2390 gnd.n2374 9.3005
R9766 gnd.n2393 gnd.n2373 9.3005
R9767 gnd.n2394 gnd.n2372 9.3005
R9768 gnd.n2397 gnd.n2371 9.3005
R9769 gnd.n2398 gnd.n2370 9.3005
R9770 gnd.n2401 gnd.n2369 9.3005
R9771 gnd.n2402 gnd.n2368 9.3005
R9772 gnd.n2405 gnd.n2367 9.3005
R9773 gnd.n2406 gnd.n2366 9.3005
R9774 gnd.n2409 gnd.n2365 9.3005
R9775 gnd.n2410 gnd.n2364 9.3005
R9776 gnd.n2413 gnd.n2363 9.3005
R9777 gnd.n2414 gnd.n2362 9.3005
R9778 gnd.n2417 gnd.n2361 9.3005
R9779 gnd.n2420 gnd.n2419 9.3005
R9780 gnd.n2384 gnd.n2379 9.3005
R9781 gnd.n2383 gnd.n2382 9.3005
R9782 gnd.n2427 gnd.n2426 9.3005
R9783 gnd.n2425 gnd.n2360 9.3005
R9784 gnd.n2424 gnd.n2423 9.3005
R9785 gnd.n2422 gnd.n977 9.3005
R9786 gnd.n4479 gnd.n978 9.3005
R9787 gnd.n4478 gnd.n979 9.3005
R9788 gnd.n4477 gnd.n980 9.3005
R9789 gnd.n996 gnd.n981 9.3005
R9790 gnd.n4467 gnd.n997 9.3005
R9791 gnd.n4466 gnd.n998 9.3005
R9792 gnd.n4465 gnd.n999 9.3005
R9793 gnd.n1018 gnd.n1000 9.3005
R9794 gnd.n4455 gnd.n1019 9.3005
R9795 gnd.n4454 gnd.n1020 9.3005
R9796 gnd.n4453 gnd.n1021 9.3005
R9797 gnd.n1042 gnd.n1022 9.3005
R9798 gnd.n1043 gnd.n1041 9.3005
R9799 gnd.n4441 gnd.n1044 9.3005
R9800 gnd.n4440 gnd.n1045 9.3005
R9801 gnd.n4439 gnd.n1046 9.3005
R9802 gnd.n2216 gnd.n1047 9.3005
R9803 gnd.n4428 gnd.n1061 9.3005
R9804 gnd.n4427 gnd.n1062 9.3005
R9805 gnd.n4426 gnd.n1063 9.3005
R9806 gnd.n1079 gnd.n1064 9.3005
R9807 gnd.n4415 gnd.n1080 9.3005
R9808 gnd.n4414 gnd.n1081 9.3005
R9809 gnd.n4413 gnd.n1082 9.3005
R9810 gnd.n1100 gnd.n1083 9.3005
R9811 gnd.n4403 gnd.n1101 9.3005
R9812 gnd.n4402 gnd.n1102 9.3005
R9813 gnd.n4401 gnd.n1103 9.3005
R9814 gnd.n1122 gnd.n1104 9.3005
R9815 gnd.n4391 gnd.n1123 9.3005
R9816 gnd.n4390 gnd.n1124 9.3005
R9817 gnd.n4389 gnd.n1125 9.3005
R9818 gnd.n1144 gnd.n1126 9.3005
R9819 gnd.n4379 gnd.n1145 9.3005
R9820 gnd.n4378 gnd.n1146 9.3005
R9821 gnd.n4377 gnd.n1147 9.3005
R9822 gnd.n1164 gnd.n1148 9.3005
R9823 gnd.n4367 gnd.n4366 9.3005
R9824 gnd.n2421 gnd.n2359 9.3005
R9825 gnd.n2834 gnd.n2156 9.3005
R9826 gnd.n2837 gnd.n2155 9.3005
R9827 gnd.n2838 gnd.n2154 9.3005
R9828 gnd.n2841 gnd.n2153 9.3005
R9829 gnd.n2842 gnd.n2152 9.3005
R9830 gnd.n2845 gnd.n2151 9.3005
R9831 gnd.n2846 gnd.n2150 9.3005
R9832 gnd.n2849 gnd.n2149 9.3005
R9833 gnd.n2850 gnd.n2148 9.3005
R9834 gnd.n2853 gnd.n2147 9.3005
R9835 gnd.n2854 gnd.n2146 9.3005
R9836 gnd.n2857 gnd.n2145 9.3005
R9837 gnd.n2858 gnd.n2144 9.3005
R9838 gnd.n2859 gnd.n2143 9.3005
R9839 gnd.n2142 gnd.n2139 9.3005
R9840 gnd.n2141 gnd.n2140 9.3005
R9841 gnd.n2623 gnd.n2622 9.3005
R9842 gnd.n2619 gnd.n2161 9.3005
R9843 gnd.n2616 gnd.n2162 9.3005
R9844 gnd.n2615 gnd.n2163 9.3005
R9845 gnd.n2612 gnd.n2164 9.3005
R9846 gnd.n2611 gnd.n2165 9.3005
R9847 gnd.n2608 gnd.n2166 9.3005
R9848 gnd.n2607 gnd.n2167 9.3005
R9849 gnd.n2604 gnd.n2168 9.3005
R9850 gnd.n2603 gnd.n2169 9.3005
R9851 gnd.n2600 gnd.n2170 9.3005
R9852 gnd.n2599 gnd.n2171 9.3005
R9853 gnd.n2596 gnd.n2172 9.3005
R9854 gnd.n2595 gnd.n2173 9.3005
R9855 gnd.n2592 gnd.n2174 9.3005
R9856 gnd.n2591 gnd.n2175 9.3005
R9857 gnd.n2588 gnd.n2176 9.3005
R9858 gnd.n2587 gnd.n2177 9.3005
R9859 gnd.n2584 gnd.n2583 9.3005
R9860 gnd.n2582 gnd.n2179 9.3005
R9861 gnd.n2624 gnd.n2157 9.3005
R9862 gnd.n4493 gnd.n4492 9.3005
R9863 gnd.n4491 gnd.n955 9.3005
R9864 gnd.n4490 gnd.n4489 9.3005
R9865 gnd.n957 gnd.n956 9.3005
R9866 gnd.n2336 gnd.n2335 9.3005
R9867 gnd.n2339 gnd.n2337 9.3005
R9868 gnd.n2340 gnd.n2334 9.3005
R9869 gnd.n2343 gnd.n2342 9.3005
R9870 gnd.n2344 gnd.n2333 9.3005
R9871 gnd.n2347 gnd.n2345 9.3005
R9872 gnd.n2348 gnd.n2332 9.3005
R9873 gnd.n2464 gnd.n2463 9.3005
R9874 gnd.n2465 gnd.n2331 9.3005
R9875 gnd.n2469 gnd.n2466 9.3005
R9876 gnd.n2468 gnd.n2467 9.3005
R9877 gnd.n2224 gnd.n2223 9.3005
R9878 gnd.n2483 gnd.n2482 9.3005
R9879 gnd.n2484 gnd.n2222 9.3005
R9880 gnd.n2486 gnd.n2485 9.3005
R9881 gnd.n2218 gnd.n2217 9.3005
R9882 gnd.n2499 gnd.n2498 9.3005
R9883 gnd.n2500 gnd.n2215 9.3005
R9884 gnd.n2502 gnd.n2501 9.3005
R9885 gnd.n2210 gnd.n2209 9.3005
R9886 gnd.n2515 gnd.n2514 9.3005
R9887 gnd.n2516 gnd.n2208 9.3005
R9888 gnd.n2518 gnd.n2517 9.3005
R9889 gnd.n2204 gnd.n2203 9.3005
R9890 gnd.n2531 gnd.n2530 9.3005
R9891 gnd.n2532 gnd.n2202 9.3005
R9892 gnd.n2534 gnd.n2533 9.3005
R9893 gnd.n2197 gnd.n2196 9.3005
R9894 gnd.n2547 gnd.n2546 9.3005
R9895 gnd.n2548 gnd.n2195 9.3005
R9896 gnd.n2550 gnd.n2549 9.3005
R9897 gnd.n2191 gnd.n2190 9.3005
R9898 gnd.n2563 gnd.n2562 9.3005
R9899 gnd.n2564 gnd.n2189 9.3005
R9900 gnd.n2567 gnd.n2566 9.3005
R9901 gnd.n2565 gnd.n2183 9.3005
R9902 gnd.n2579 gnd.n2182 9.3005
R9903 gnd.n2581 gnd.n2580 9.3005
R9904 gnd.n4494 gnd.n953 9.3005
R9905 gnd.n4501 gnd.n4500 9.3005
R9906 gnd.n4502 gnd.n947 9.3005
R9907 gnd.n4505 gnd.n946 9.3005
R9908 gnd.n4506 gnd.n945 9.3005
R9909 gnd.n4509 gnd.n944 9.3005
R9910 gnd.n4510 gnd.n943 9.3005
R9911 gnd.n4513 gnd.n942 9.3005
R9912 gnd.n4514 gnd.n941 9.3005
R9913 gnd.n4517 gnd.n940 9.3005
R9914 gnd.n4518 gnd.n939 9.3005
R9915 gnd.n4521 gnd.n938 9.3005
R9916 gnd.n4522 gnd.n937 9.3005
R9917 gnd.n4525 gnd.n936 9.3005
R9918 gnd.n4526 gnd.n935 9.3005
R9919 gnd.n4529 gnd.n934 9.3005
R9920 gnd.n4530 gnd.n933 9.3005
R9921 gnd.n4533 gnd.n932 9.3005
R9922 gnd.n4534 gnd.n931 9.3005
R9923 gnd.n4537 gnd.n930 9.3005
R9924 gnd.n4539 gnd.n927 9.3005
R9925 gnd.n4542 gnd.n926 9.3005
R9926 gnd.n4543 gnd.n925 9.3005
R9927 gnd.n4546 gnd.n924 9.3005
R9928 gnd.n4547 gnd.n923 9.3005
R9929 gnd.n4550 gnd.n922 9.3005
R9930 gnd.n4551 gnd.n921 9.3005
R9931 gnd.n4554 gnd.n920 9.3005
R9932 gnd.n4555 gnd.n919 9.3005
R9933 gnd.n4558 gnd.n918 9.3005
R9934 gnd.n4559 gnd.n917 9.3005
R9935 gnd.n4562 gnd.n916 9.3005
R9936 gnd.n4563 gnd.n915 9.3005
R9937 gnd.n4566 gnd.n914 9.3005
R9938 gnd.n4568 gnd.n913 9.3005
R9939 gnd.n4569 gnd.n912 9.3005
R9940 gnd.n4570 gnd.n911 9.3005
R9941 gnd.n4571 gnd.n910 9.3005
R9942 gnd.n4499 gnd.n952 9.3005
R9943 gnd.n4498 gnd.n4497 9.3005
R9944 gnd.n2433 gnd.n2432 9.3005
R9945 gnd.n2431 gnd.n966 9.3005
R9946 gnd.n4485 gnd.n967 9.3005
R9947 gnd.n4484 gnd.n968 9.3005
R9948 gnd.n4483 gnd.n969 9.3005
R9949 gnd.n987 gnd.n970 9.3005
R9950 gnd.n4473 gnd.n988 9.3005
R9951 gnd.n4472 gnd.n989 9.3005
R9952 gnd.n4471 gnd.n990 9.3005
R9953 gnd.n1007 gnd.n991 9.3005
R9954 gnd.n4461 gnd.n1008 9.3005
R9955 gnd.n4460 gnd.n1009 9.3005
R9956 gnd.n4459 gnd.n1010 9.3005
R9957 gnd.n1029 gnd.n1011 9.3005
R9958 gnd.n4449 gnd.n1030 9.3005
R9959 gnd.n1090 gnd.n1072 9.3005
R9960 gnd.n4409 gnd.n1091 9.3005
R9961 gnd.n4408 gnd.n1092 9.3005
R9962 gnd.n4407 gnd.n1093 9.3005
R9963 gnd.n1111 gnd.n1094 9.3005
R9964 gnd.n4397 gnd.n1112 9.3005
R9965 gnd.n4396 gnd.n1113 9.3005
R9966 gnd.n4395 gnd.n1114 9.3005
R9967 gnd.n1133 gnd.n1115 9.3005
R9968 gnd.n4385 gnd.n1134 9.3005
R9969 gnd.n4384 gnd.n1135 9.3005
R9970 gnd.n4383 gnd.n1136 9.3005
R9971 gnd.n1154 gnd.n1137 9.3005
R9972 gnd.n4373 gnd.n1155 9.3005
R9973 gnd.n4372 gnd.n1156 9.3005
R9974 gnd.n4371 gnd.n1157 9.3005
R9975 gnd.n2430 gnd.n2429 9.3005
R9976 gnd.n4419 gnd.n1031 9.3005
R9977 gnd.n2308 gnd.n2307 9.3005
R9978 gnd.n2319 gnd.n2318 9.3005
R9979 gnd.n2320 gnd.n2228 9.3005
R9980 gnd.n2314 gnd.n2313 9.3005
R9981 gnd.n2310 gnd.n802 9.3005
R9982 gnd.n5955 gnd.n801 9.3005
R9983 gnd.n5956 gnd.n800 9.3005
R9984 gnd.n5957 gnd.n799 9.3005
R9985 gnd.n798 gnd.n794 9.3005
R9986 gnd.n5963 gnd.n793 9.3005
R9987 gnd.n5964 gnd.n792 9.3005
R9988 gnd.n5965 gnd.n791 9.3005
R9989 gnd.n790 gnd.n786 9.3005
R9990 gnd.n5971 gnd.n785 9.3005
R9991 gnd.n5972 gnd.n784 9.3005
R9992 gnd.n5973 gnd.n783 9.3005
R9993 gnd.n782 gnd.n778 9.3005
R9994 gnd.n5979 gnd.n777 9.3005
R9995 gnd.n5980 gnd.n776 9.3005
R9996 gnd.n5981 gnd.n775 9.3005
R9997 gnd.n774 gnd.n770 9.3005
R9998 gnd.n5987 gnd.n769 9.3005
R9999 gnd.n5988 gnd.n768 9.3005
R10000 gnd.n5989 gnd.n767 9.3005
R10001 gnd.n766 gnd.n762 9.3005
R10002 gnd.n5995 gnd.n761 9.3005
R10003 gnd.n5996 gnd.n760 9.3005
R10004 gnd.n5997 gnd.n759 9.3005
R10005 gnd.n758 gnd.n754 9.3005
R10006 gnd.n6003 gnd.n753 9.3005
R10007 gnd.n6004 gnd.n752 9.3005
R10008 gnd.n6005 gnd.n751 9.3005
R10009 gnd.n750 gnd.n746 9.3005
R10010 gnd.n6011 gnd.n745 9.3005
R10011 gnd.n6012 gnd.n744 9.3005
R10012 gnd.n6013 gnd.n743 9.3005
R10013 gnd.n742 gnd.n738 9.3005
R10014 gnd.n6019 gnd.n737 9.3005
R10015 gnd.n6020 gnd.n736 9.3005
R10016 gnd.n6021 gnd.n735 9.3005
R10017 gnd.n734 gnd.n730 9.3005
R10018 gnd.n6027 gnd.n729 9.3005
R10019 gnd.n6028 gnd.n728 9.3005
R10020 gnd.n6029 gnd.n727 9.3005
R10021 gnd.n726 gnd.n722 9.3005
R10022 gnd.n6035 gnd.n721 9.3005
R10023 gnd.n6036 gnd.n720 9.3005
R10024 gnd.n6037 gnd.n719 9.3005
R10025 gnd.n718 gnd.n714 9.3005
R10026 gnd.n6043 gnd.n713 9.3005
R10027 gnd.n6044 gnd.n712 9.3005
R10028 gnd.n6045 gnd.n711 9.3005
R10029 gnd.n710 gnd.n706 9.3005
R10030 gnd.n6051 gnd.n705 9.3005
R10031 gnd.n6052 gnd.n704 9.3005
R10032 gnd.n6053 gnd.n703 9.3005
R10033 gnd.n702 gnd.n698 9.3005
R10034 gnd.n6059 gnd.n697 9.3005
R10035 gnd.n6060 gnd.n696 9.3005
R10036 gnd.n6061 gnd.n695 9.3005
R10037 gnd.n694 gnd.n690 9.3005
R10038 gnd.n6067 gnd.n689 9.3005
R10039 gnd.n6068 gnd.n688 9.3005
R10040 gnd.n6069 gnd.n687 9.3005
R10041 gnd.n686 gnd.n682 9.3005
R10042 gnd.n6075 gnd.n681 9.3005
R10043 gnd.n6076 gnd.n680 9.3005
R10044 gnd.n6077 gnd.n679 9.3005
R10045 gnd.n678 gnd.n674 9.3005
R10046 gnd.n6083 gnd.n673 9.3005
R10047 gnd.n6084 gnd.n672 9.3005
R10048 gnd.n6085 gnd.n671 9.3005
R10049 gnd.n670 gnd.n666 9.3005
R10050 gnd.n6091 gnd.n665 9.3005
R10051 gnd.n6092 gnd.n664 9.3005
R10052 gnd.n6093 gnd.n663 9.3005
R10053 gnd.n662 gnd.n658 9.3005
R10054 gnd.n6099 gnd.n657 9.3005
R10055 gnd.n6100 gnd.n656 9.3005
R10056 gnd.n6101 gnd.n655 9.3005
R10057 gnd.n654 gnd.n650 9.3005
R10058 gnd.n6107 gnd.n649 9.3005
R10059 gnd.n6108 gnd.n648 9.3005
R10060 gnd.n6109 gnd.n647 9.3005
R10061 gnd.n646 gnd.n642 9.3005
R10062 gnd.n6115 gnd.n641 9.3005
R10063 gnd.n6116 gnd.n640 9.3005
R10064 gnd.n6117 gnd.n639 9.3005
R10065 gnd.n2312 gnd.n2311 9.3005
R10066 gnd.n1557 gnd.n1556 9.3005
R10067 gnd.n1563 gnd.n1562 9.3005
R10068 gnd.n1564 gnd.n1539 9.3005
R10069 gnd.n1573 gnd.n1572 9.3005
R10070 gnd.n1541 gnd.n1537 9.3005
R10071 gnd.n1580 gnd.n1579 9.3005
R10072 gnd.n1581 gnd.n1530 9.3005
R10073 gnd.n1590 gnd.n1589 9.3005
R10074 gnd.n1532 gnd.n1528 9.3005
R10075 gnd.n1597 gnd.n1596 9.3005
R10076 gnd.n1598 gnd.n1521 9.3005
R10077 gnd.n1607 gnd.n1606 9.3005
R10078 gnd.n1523 gnd.n1519 9.3005
R10079 gnd.n1614 gnd.n1613 9.3005
R10080 gnd.n1615 gnd.n1509 9.3005
R10081 gnd.n1622 gnd.n1621 9.3005
R10082 gnd.n1511 gnd.n1507 9.3005
R10083 gnd.n1506 gnd.n1504 9.3005
R10084 gnd.n1547 gnd.n1546 9.3005
R10085 gnd.n1617 gnd.n1616 9.3005
R10086 gnd.n1518 gnd.n1515 9.3005
R10087 gnd.n1605 gnd.n1604 9.3005
R10088 gnd.n1601 gnd.n1522 9.3005
R10089 gnd.n1600 gnd.n1599 9.3005
R10090 gnd.n1527 gnd.n1524 9.3005
R10091 gnd.n1588 gnd.n1587 9.3005
R10092 gnd.n1584 gnd.n1531 9.3005
R10093 gnd.n1583 gnd.n1582 9.3005
R10094 gnd.n1536 gnd.n1533 9.3005
R10095 gnd.n1571 gnd.n1570 9.3005
R10096 gnd.n1567 gnd.n1540 9.3005
R10097 gnd.n1566 gnd.n1565 9.3005
R10098 gnd.n1545 gnd.n1542 9.3005
R10099 gnd.n1555 gnd.n1554 9.3005
R10100 gnd.n1551 gnd.n1550 9.3005
R10101 gnd.n1618 gnd.n1510 9.3005
R10102 gnd.n1620 gnd.n1619 9.3005
R10103 gnd.n3911 gnd.n3910 9.3005
R10104 gnd.n3909 gnd.n1505 9.3005
R10105 gnd.n3908 gnd.n3907 9.3005
R10106 gnd.n3906 gnd.n1632 9.3005
R10107 gnd.n3905 gnd.n3904 9.3005
R10108 gnd.n3903 gnd.n1633 9.3005
R10109 gnd.n3899 gnd.n3898 9.3005
R10110 gnd.n3897 gnd.n1640 9.3005
R10111 gnd.n3896 gnd.n3895 9.3005
R10112 gnd.n3894 gnd.n3889 9.3005
R10113 gnd.n2912 gnd.n1975 9.3005
R10114 gnd.n2914 gnd.n2913 9.3005
R10115 gnd.n1961 gnd.n1960 9.3005
R10116 gnd.n2929 gnd.n2928 9.3005
R10117 gnd.n2930 gnd.n1958 9.3005
R10118 gnd.n2933 gnd.n2932 9.3005
R10119 gnd.n2931 gnd.n1959 9.3005
R10120 gnd.n1930 gnd.n1929 9.3005
R10121 gnd.n3051 gnd.n3050 9.3005
R10122 gnd.n3052 gnd.n1928 9.3005
R10123 gnd.n3054 gnd.n3053 9.3005
R10124 gnd.n1916 gnd.n1915 9.3005
R10125 gnd.n3067 gnd.n3066 9.3005
R10126 gnd.n3068 gnd.n1914 9.3005
R10127 gnd.n3070 gnd.n3069 9.3005
R10128 gnd.n1902 gnd.n1901 9.3005
R10129 gnd.n3083 gnd.n3082 9.3005
R10130 gnd.n3084 gnd.n1900 9.3005
R10131 gnd.n3086 gnd.n3085 9.3005
R10132 gnd.n1886 gnd.n1885 9.3005
R10133 gnd.n3100 gnd.n3099 9.3005
R10134 gnd.n3101 gnd.n1883 9.3005
R10135 gnd.n3104 gnd.n3103 9.3005
R10136 gnd.n3102 gnd.n1884 9.3005
R10137 gnd.n1855 gnd.n1854 9.3005
R10138 gnd.n3224 gnd.n3223 9.3005
R10139 gnd.n3225 gnd.n1853 9.3005
R10140 gnd.n3227 gnd.n3226 9.3005
R10141 gnd.n1842 gnd.n1841 9.3005
R10142 gnd.n3240 gnd.n3239 9.3005
R10143 gnd.n3241 gnd.n1840 9.3005
R10144 gnd.n3243 gnd.n3242 9.3005
R10145 gnd.n1830 gnd.n1829 9.3005
R10146 gnd.n3256 gnd.n3255 9.3005
R10147 gnd.n3257 gnd.n1828 9.3005
R10148 gnd.n3259 gnd.n3258 9.3005
R10149 gnd.n1816 gnd.n1815 9.3005
R10150 gnd.n3274 gnd.n3273 9.3005
R10151 gnd.n3275 gnd.n1813 9.3005
R10152 gnd.n3278 gnd.n3277 9.3005
R10153 gnd.n3276 gnd.n1814 9.3005
R10154 gnd.n1783 gnd.n1782 9.3005
R10155 gnd.n3395 gnd.n3394 9.3005
R10156 gnd.n3396 gnd.n1781 9.3005
R10157 gnd.n3398 gnd.n3397 9.3005
R10158 gnd.n1768 gnd.n1767 9.3005
R10159 gnd.n3411 gnd.n3410 9.3005
R10160 gnd.n3412 gnd.n1766 9.3005
R10161 gnd.n3414 gnd.n3413 9.3005
R10162 gnd.n1754 gnd.n1753 9.3005
R10163 gnd.n3427 gnd.n3426 9.3005
R10164 gnd.n3428 gnd.n1752 9.3005
R10165 gnd.n3430 gnd.n3429 9.3005
R10166 gnd.n1739 gnd.n1738 9.3005
R10167 gnd.n3445 gnd.n3444 9.3005
R10168 gnd.n3446 gnd.n1736 9.3005
R10169 gnd.n3449 gnd.n3448 9.3005
R10170 gnd.n3447 gnd.n1737 9.3005
R10171 gnd.n1709 gnd.n1708 9.3005
R10172 gnd.n3801 gnd.n3800 9.3005
R10173 gnd.n3802 gnd.n1707 9.3005
R10174 gnd.n3804 gnd.n3803 9.3005
R10175 gnd.n1696 gnd.n1695 9.3005
R10176 gnd.n3817 gnd.n3816 9.3005
R10177 gnd.n3818 gnd.n1694 9.3005
R10178 gnd.n3820 gnd.n3819 9.3005
R10179 gnd.n1683 gnd.n1682 9.3005
R10180 gnd.n3833 gnd.n3832 9.3005
R10181 gnd.n3834 gnd.n1681 9.3005
R10182 gnd.n3836 gnd.n3835 9.3005
R10183 gnd.n1669 gnd.n1668 9.3005
R10184 gnd.n3849 gnd.n3848 9.3005
R10185 gnd.n3850 gnd.n1667 9.3005
R10186 gnd.n3852 gnd.n3851 9.3005
R10187 gnd.n1655 gnd.n1654 9.3005
R10188 gnd.n3865 gnd.n3864 9.3005
R10189 gnd.n3866 gnd.n1652 9.3005
R10190 gnd.n3870 gnd.n3869 9.3005
R10191 gnd.n3868 gnd.n1653 9.3005
R10192 gnd.n3867 gnd.n1642 9.3005
R10193 gnd.n3886 gnd.n1641 9.3005
R10194 gnd.n3888 gnd.n3887 9.3005
R10195 gnd.n2911 gnd.n2910 9.3005
R10196 gnd.n2897 gnd.n2896 9.3005
R10197 gnd.n2895 gnd.n2000 9.3005
R10198 gnd.n2894 gnd.n2893 9.3005
R10199 gnd.n2890 gnd.n2002 9.3005
R10200 gnd.n2887 gnd.n2886 9.3005
R10201 gnd.n2885 gnd.n2005 9.3005
R10202 gnd.n2884 gnd.n2883 9.3005
R10203 gnd.n2880 gnd.n2006 9.3005
R10204 gnd.n2877 gnd.n2876 9.3005
R10205 gnd.n2001 gnd.n1976 9.3005
R10206 gnd.n2213 gnd.n2212 9.3005
R10207 gnd.n2507 gnd.n2506 9.3005
R10208 gnd.n2508 gnd.n2211 9.3005
R10209 gnd.n2510 gnd.n2509 9.3005
R10210 gnd.n2207 gnd.n2206 9.3005
R10211 gnd.n2523 gnd.n2522 9.3005
R10212 gnd.n2524 gnd.n2205 9.3005
R10213 gnd.n2526 gnd.n2525 9.3005
R10214 gnd.n2200 gnd.n2199 9.3005
R10215 gnd.n2539 gnd.n2538 9.3005
R10216 gnd.n2540 gnd.n2198 9.3005
R10217 gnd.n2542 gnd.n2541 9.3005
R10218 gnd.n2194 gnd.n2193 9.3005
R10219 gnd.n2555 gnd.n2554 9.3005
R10220 gnd.n2556 gnd.n2192 9.3005
R10221 gnd.n2558 gnd.n2557 9.3005
R10222 gnd.n2188 gnd.n2187 9.3005
R10223 gnd.n2572 gnd.n2571 9.3005
R10224 gnd.n2573 gnd.n2185 9.3005
R10225 gnd.n2575 gnd.n2574 9.3005
R10226 gnd.n2186 gnd.n2008 9.3005
R10227 gnd.n2874 gnd.n2007 9.3005
R10228 gnd.n2873 gnd.n2872 9.3005
R10229 gnd.n2869 gnd.n2868 9.3005
R10230 gnd.n2013 gnd.n2010 9.3005
R10231 gnd.n2112 gnd.n2111 9.3005
R10232 gnd.n2108 gnd.n2028 9.3005
R10233 gnd.n2107 gnd.n2106 9.3005
R10234 gnd.n2033 gnd.n2030 9.3005
R10235 gnd.n2098 gnd.n2097 9.3005
R10236 gnd.n2094 gnd.n2093 9.3005
R10237 gnd.n2037 gnd.n2036 9.3005
R10238 gnd.n2086 gnd.n2085 9.3005
R10239 gnd.n2082 gnd.n2081 9.3005
R10240 gnd.n2045 gnd.n2042 9.3005
R10241 gnd.n2074 gnd.n2073 9.3005
R10242 gnd.n2070 gnd.n2069 9.3005
R10243 gnd.n2049 gnd.n2048 9.3005
R10244 gnd.n2062 gnd.n2061 9.3005
R10245 gnd.n2058 gnd.n2056 9.3005
R10246 gnd.n2051 gnd.n1166 9.3005
R10247 gnd.n2055 gnd.n2052 9.3005
R10248 gnd.n2064 gnd.n2063 9.3005
R10249 gnd.n2068 gnd.n2067 9.3005
R10250 gnd.n2047 gnd.n2046 9.3005
R10251 gnd.n2076 gnd.n2075 9.3005
R10252 gnd.n2080 gnd.n2079 9.3005
R10253 gnd.n2041 gnd.n2038 9.3005
R10254 gnd.n2088 gnd.n2087 9.3005
R10255 gnd.n2092 gnd.n2091 9.3005
R10256 gnd.n2035 gnd.n2034 9.3005
R10257 gnd.n2100 gnd.n2099 9.3005
R10258 gnd.n2104 gnd.n2103 9.3005
R10259 gnd.n2105 gnd.n2027 9.3005
R10260 gnd.n2114 gnd.n2113 9.3005
R10261 gnd.n2029 gnd.n2014 9.3005
R10262 gnd.n2867 gnd.n2866 9.3005
R10263 gnd.n2865 gnd.n2009 9.3005
R10264 gnd.n4361 gnd.n1167 9.3005
R10265 gnd.n4360 gnd.n4359 9.3005
R10266 gnd.n4358 gnd.n1171 9.3005
R10267 gnd.n4357 gnd.n4356 9.3005
R10268 gnd.n4355 gnd.n1172 9.3005
R10269 gnd.n4354 gnd.n4353 9.3005
R10270 gnd.n4352 gnd.n1176 9.3005
R10271 gnd.n4351 gnd.n4350 9.3005
R10272 gnd.n4349 gnd.n1177 9.3005
R10273 gnd.n4348 gnd.n4347 9.3005
R10274 gnd.n4346 gnd.n1181 9.3005
R10275 gnd.n4345 gnd.n4344 9.3005
R10276 gnd.n4343 gnd.n1182 9.3005
R10277 gnd.n4342 gnd.n4341 9.3005
R10278 gnd.n4340 gnd.n1186 9.3005
R10279 gnd.n4339 gnd.n4338 9.3005
R10280 gnd.n4337 gnd.n1187 9.3005
R10281 gnd.n4336 gnd.n4335 9.3005
R10282 gnd.n4334 gnd.n1191 9.3005
R10283 gnd.n4333 gnd.n4332 9.3005
R10284 gnd.n4331 gnd.n1192 9.3005
R10285 gnd.n4330 gnd.n4329 9.3005
R10286 gnd.n4328 gnd.n1196 9.3005
R10287 gnd.n4327 gnd.n4326 9.3005
R10288 gnd.n4325 gnd.n1197 9.3005
R10289 gnd.n4324 gnd.n4323 9.3005
R10290 gnd.n4322 gnd.n1201 9.3005
R10291 gnd.n4321 gnd.n4320 9.3005
R10292 gnd.n4319 gnd.n1202 9.3005
R10293 gnd.n4318 gnd.n4317 9.3005
R10294 gnd.n4316 gnd.n1206 9.3005
R10295 gnd.n4315 gnd.n4314 9.3005
R10296 gnd.n4313 gnd.n1207 9.3005
R10297 gnd.n4312 gnd.n4311 9.3005
R10298 gnd.n4310 gnd.n1211 9.3005
R10299 gnd.n4309 gnd.n4308 9.3005
R10300 gnd.n4307 gnd.n1212 9.3005
R10301 gnd.n4306 gnd.n4305 9.3005
R10302 gnd.n4304 gnd.n1216 9.3005
R10303 gnd.n4303 gnd.n4302 9.3005
R10304 gnd.n4301 gnd.n1217 9.3005
R10305 gnd.n4300 gnd.n4299 9.3005
R10306 gnd.n4298 gnd.n1221 9.3005
R10307 gnd.n4297 gnd.n4296 9.3005
R10308 gnd.n4295 gnd.n1222 9.3005
R10309 gnd.n4294 gnd.n4293 9.3005
R10310 gnd.n4292 gnd.n1226 9.3005
R10311 gnd.n4291 gnd.n4290 9.3005
R10312 gnd.n4289 gnd.n1227 9.3005
R10313 gnd.n4288 gnd.n4287 9.3005
R10314 gnd.n4286 gnd.n1231 9.3005
R10315 gnd.n4285 gnd.n4284 9.3005
R10316 gnd.n4283 gnd.n1232 9.3005
R10317 gnd.n4282 gnd.n4281 9.3005
R10318 gnd.n4280 gnd.n1236 9.3005
R10319 gnd.n4279 gnd.n4278 9.3005
R10320 gnd.n4277 gnd.n1237 9.3005
R10321 gnd.n4276 gnd.n4275 9.3005
R10322 gnd.n4274 gnd.n1241 9.3005
R10323 gnd.n4273 gnd.n4272 9.3005
R10324 gnd.n4271 gnd.n1242 9.3005
R10325 gnd.n4270 gnd.n4269 9.3005
R10326 gnd.n4268 gnd.n1246 9.3005
R10327 gnd.n4267 gnd.n4266 9.3005
R10328 gnd.n4265 gnd.n1247 9.3005
R10329 gnd.n4264 gnd.n4263 9.3005
R10330 gnd.n4262 gnd.n1251 9.3005
R10331 gnd.n4261 gnd.n4260 9.3005
R10332 gnd.n4259 gnd.n1252 9.3005
R10333 gnd.n4258 gnd.n4257 9.3005
R10334 gnd.n4256 gnd.n1256 9.3005
R10335 gnd.n4255 gnd.n4254 9.3005
R10336 gnd.n4253 gnd.n1257 9.3005
R10337 gnd.n4252 gnd.n4251 9.3005
R10338 gnd.n4250 gnd.n1261 9.3005
R10339 gnd.n4249 gnd.n4248 9.3005
R10340 gnd.n4247 gnd.n1262 9.3005
R10341 gnd.n4246 gnd.n4245 9.3005
R10342 gnd.n4244 gnd.n1266 9.3005
R10343 gnd.n4243 gnd.n4242 9.3005
R10344 gnd.n4241 gnd.n1267 9.3005
R10345 gnd.n4240 gnd.n1270 9.3005
R10346 gnd.n4363 gnd.n4362 9.3005
R10347 gnd.n4149 gnd.n1367 9.3005
R10348 gnd.n4148 gnd.n4147 9.3005
R10349 gnd.n4146 gnd.n1369 9.3005
R10350 gnd.n4145 gnd.n4144 9.3005
R10351 gnd.n4143 gnd.n1373 9.3005
R10352 gnd.n4142 gnd.n4141 9.3005
R10353 gnd.n4140 gnd.n1374 9.3005
R10354 gnd.n4139 gnd.n4138 9.3005
R10355 gnd.n4137 gnd.n1378 9.3005
R10356 gnd.n4136 gnd.n4135 9.3005
R10357 gnd.n4134 gnd.n1379 9.3005
R10358 gnd.n4133 gnd.n4132 9.3005
R10359 gnd.n4131 gnd.n1383 9.3005
R10360 gnd.n4130 gnd.n4129 9.3005
R10361 gnd.n4128 gnd.n1384 9.3005
R10362 gnd.n4127 gnd.n4126 9.3005
R10363 gnd.n4125 gnd.n1388 9.3005
R10364 gnd.n4124 gnd.n4123 9.3005
R10365 gnd.n4122 gnd.n1389 9.3005
R10366 gnd.n4121 gnd.n4120 9.3005
R10367 gnd.n4119 gnd.n1393 9.3005
R10368 gnd.n4118 gnd.n4117 9.3005
R10369 gnd.n227 gnd.n226 9.3005
R10370 gnd.n6747 gnd.n6746 9.3005
R10371 gnd.n6748 gnd.n225 9.3005
R10372 gnd.n6750 gnd.n6749 9.3005
R10373 gnd.n206 gnd.n205 9.3005
R10374 gnd.n6763 gnd.n6762 9.3005
R10375 gnd.n6764 gnd.n204 9.3005
R10376 gnd.n6766 gnd.n6765 9.3005
R10377 gnd.n192 gnd.n191 9.3005
R10378 gnd.n6779 gnd.n6778 9.3005
R10379 gnd.n6780 gnd.n190 9.3005
R10380 gnd.n6782 gnd.n6781 9.3005
R10381 gnd.n177 gnd.n176 9.3005
R10382 gnd.n6795 gnd.n6794 9.3005
R10383 gnd.n6796 gnd.n174 9.3005
R10384 gnd.n6872 gnd.n6871 9.3005
R10385 gnd.n6870 gnd.n175 9.3005
R10386 gnd.n6869 gnd.n6868 9.3005
R10387 gnd.n6867 gnd.n6797 9.3005
R10388 gnd.n6866 gnd.n6865 9.3005
R10389 gnd.n4151 gnd.n4150 9.3005
R10390 gnd.n6862 gnd.n6799 9.3005
R10391 gnd.n6861 gnd.n6860 9.3005
R10392 gnd.n6859 gnd.n6804 9.3005
R10393 gnd.n6858 gnd.n6857 9.3005
R10394 gnd.n6856 gnd.n6805 9.3005
R10395 gnd.n6855 gnd.n6854 9.3005
R10396 gnd.n6853 gnd.n6812 9.3005
R10397 gnd.n6852 gnd.n6851 9.3005
R10398 gnd.n6850 gnd.n6813 9.3005
R10399 gnd.n6849 gnd.n6848 9.3005
R10400 gnd.n6847 gnd.n6820 9.3005
R10401 gnd.n6846 gnd.n6845 9.3005
R10402 gnd.n6844 gnd.n6821 9.3005
R10403 gnd.n6843 gnd.n6842 9.3005
R10404 gnd.n6841 gnd.n6828 9.3005
R10405 gnd.n6840 gnd.n6839 9.3005
R10406 gnd.n6838 gnd.n6829 9.3005
R10407 gnd.n6837 gnd.n78 9.3005
R10408 gnd.n6864 gnd.n6863 9.3005
R10409 gnd.n3915 gnd.n3914 9.3005
R10410 gnd.n1493 gnd.n1492 9.3005
R10411 gnd.n3987 gnd.n3986 9.3005
R10412 gnd.n3988 gnd.n1490 9.3005
R10413 gnd.n3991 gnd.n3990 9.3005
R10414 gnd.n3989 gnd.n1491 9.3005
R10415 gnd.n1467 gnd.n1466 9.3005
R10416 gnd.n4019 gnd.n4018 9.3005
R10417 gnd.n4020 gnd.n1464 9.3005
R10418 gnd.n4023 gnd.n4022 9.3005
R10419 gnd.n4021 gnd.n1465 9.3005
R10420 gnd.n1441 gnd.n1440 9.3005
R10421 gnd.n4054 gnd.n4053 9.3005
R10422 gnd.n4055 gnd.n1439 9.3005
R10423 gnd.n4057 gnd.n4056 9.3005
R10424 gnd.n1413 gnd.n1412 9.3005
R10425 gnd.n4085 gnd.n4084 9.3005
R10426 gnd.n4086 gnd.n1410 9.3005
R10427 gnd.n4088 gnd.n4087 9.3005
R10428 gnd.n1411 gnd.n51 9.3005
R10429 gnd.n6996 gnd.n52 9.3005
R10430 gnd.n6995 gnd.n6994 9.3005
R10431 gnd.n6993 gnd.n53 9.3005
R10432 gnd.n6992 gnd.n6991 9.3005
R10433 gnd.n6990 gnd.n57 9.3005
R10434 gnd.n6989 gnd.n6988 9.3005
R10435 gnd.n6987 gnd.n58 9.3005
R10436 gnd.n6986 gnd.n6985 9.3005
R10437 gnd.n6984 gnd.n62 9.3005
R10438 gnd.n6983 gnd.n6982 9.3005
R10439 gnd.n6981 gnd.n63 9.3005
R10440 gnd.n6980 gnd.n6979 9.3005
R10441 gnd.n6978 gnd.n67 9.3005
R10442 gnd.n6977 gnd.n6976 9.3005
R10443 gnd.n6975 gnd.n68 9.3005
R10444 gnd.n6974 gnd.n6973 9.3005
R10445 gnd.n6972 gnd.n72 9.3005
R10446 gnd.n6971 gnd.n6970 9.3005
R10447 gnd.n6969 gnd.n73 9.3005
R10448 gnd.n6968 gnd.n6967 9.3005
R10449 gnd.n6966 gnd.n77 9.3005
R10450 gnd.n6965 gnd.n6964 9.3005
R10451 gnd.n3913 gnd.n1503 9.3005
R10452 gnd.t250 gnd.n4698 9.24152
R10453 gnd.t153 gnd.n842 9.24152
R10454 gnd.n5821 gnd.t167 9.24152
R10455 gnd.t261 gnd.t250 8.92286
R10456 gnd.n2926 gnd.n1964 8.92286
R10457 gnd.n3097 gnd.n1889 8.92286
R10458 gnd.n3205 gnd.n1875 8.92286
R10459 gnd.n3271 gnd.n1819 8.92286
R10460 gnd.n3376 gnd.n1804 8.92286
R10461 gnd.n3442 gnd.n1743 8.92286
R10462 gnd.n3782 gnd.n1727 8.92286
R10463 gnd.n3846 gnd.n1672 8.92286
R10464 gnd.n3872 gnd.n1650 8.92286
R10465 gnd.n5800 gnd.n5775 8.92171
R10466 gnd.n5768 gnd.n5743 8.92171
R10467 gnd.n5736 gnd.n5711 8.92171
R10468 gnd.n5705 gnd.n5680 8.92171
R10469 gnd.n5673 gnd.n5648 8.92171
R10470 gnd.n5641 gnd.n5616 8.92171
R10471 gnd.n5609 gnd.n5584 8.92171
R10472 gnd.n5578 gnd.n5553 8.92171
R10473 gnd.n3538 gnd.n3520 8.72777
R10474 gnd.t84 gnd.n4781 8.60421
R10475 gnd.n2916 gnd.n1973 8.60421
R10476 gnd.n3160 gnd.t108 8.60421
R10477 gnd.t238 gnd.n1787 8.60421
R10478 gnd.n4753 gnd.n4741 8.43467
R10479 gnd.n38 gnd.n26 8.43467
R10480 gnd.n2493 gnd.n0 8.41456
R10481 gnd.n6997 gnd.n6996 8.41456
R10482 gnd.n1972 gnd.t194 8.28555
R10483 gnd.n5801 gnd.n5773 8.14595
R10484 gnd.n5769 gnd.n5741 8.14595
R10485 gnd.n5737 gnd.n5709 8.14595
R10486 gnd.n5706 gnd.n5678 8.14595
R10487 gnd.n5674 gnd.n5646 8.14595
R10488 gnd.n5642 gnd.n5614 8.14595
R10489 gnd.n5610 gnd.n5582 8.14595
R10490 gnd.n5579 gnd.n5551 8.14595
R10491 gnd.n5806 gnd.n5805 7.97301
R10492 gnd.n5274 gnd.t68 7.9669
R10493 gnd.n3010 gnd.t252 7.9669
R10494 gnd.t270 gnd.n1692 7.9669
R10495 gnd.n6838 gnd.n6837 7.75808
R10496 gnd.n1619 gnd.n1618 7.75808
R10497 gnd.n2866 gnd.n2865 7.75808
R10498 gnd.n2382 gnd.n2379 7.75808
R10499 gnd.n1941 gnd.t213 7.64824
R10500 gnd.n3025 gnd.n3024 7.64824
R10501 gnd.t79 gnd.n1898 7.64824
R10502 gnd.n3181 gnd.t35 7.64824
R10503 gnd.n3253 gnd.t35 7.64824
R10504 gnd.n3299 gnd.t234 7.64824
R10505 gnd.t234 gnd.n1763 7.64824
R10506 gnd.n3775 gnd.t232 7.64824
R10507 gnd.n3838 gnd.n1679 7.64824
R10508 gnd.n3501 gnd.t200 7.64824
R10509 gnd.t249 gnd.n4867 7.32958
R10510 gnd.t244 gnd.t150 7.32958
R10511 gnd.n2667 gnd.n2666 7.30353
R10512 gnd.n3537 gnd.n3536 7.30353
R10513 gnd.n5176 gnd.n5175 7.01093
R10514 gnd.n5186 gnd.n4896 7.01093
R10515 gnd.n5185 gnd.n4899 7.01093
R10516 gnd.n5194 gnd.n4890 7.01093
R10517 gnd.n5198 gnd.n5197 7.01093
R10518 gnd.n5216 gnd.n4875 7.01093
R10519 gnd.n5215 gnd.n4878 7.01093
R10520 gnd.n5226 gnd.n4867 7.01093
R10521 gnd.n4868 gnd.n4856 7.01093
R10522 gnd.n5239 gnd.n4857 7.01093
R10523 gnd.n5250 gnd.n4849 7.01093
R10524 gnd.n5249 gnd.n4840 7.01093
R10525 gnd.n4842 gnd.n4824 7.01093
R10526 gnd.n5286 gnd.n4825 7.01093
R10527 gnd.n5275 gnd.n5274 7.01093
R10528 gnd.n5311 gnd.n4816 7.01093
R10529 gnd.n5322 gnd.n5321 7.01093
R10530 gnd.n4809 gnd.n4801 7.01093
R10531 gnd.n5351 gnd.n4789 7.01093
R10532 gnd.n5350 gnd.n4792 7.01093
R10533 gnd.n5361 gnd.n4781 7.01093
R10534 gnd.n4782 gnd.n4770 7.01093
R10535 gnd.n5372 gnd.n4771 7.01093
R10536 gnd.n5396 gnd.n4726 7.01093
R10537 gnd.n5395 gnd.n4717 7.01093
R10538 gnd.n4719 gnd.n4710 7.01093
R10539 gnd.n5418 gnd.n5417 7.01093
R10540 gnd.n5435 gnd.n4698 7.01093
R10541 gnd.n5434 gnd.n4701 7.01093
R10542 gnd.n5448 gnd.n4690 7.01093
R10543 gnd.n4691 gnd.n4679 7.01093
R10544 gnd.n5458 gnd.n4681 7.01093
R10545 gnd.n5489 gnd.n5488 7.01093
R10546 gnd.n5502 gnd.n5501 7.01093
R10547 gnd.n4660 gnd.n4650 7.01093
R10548 gnd.n5514 gnd.n5513 7.01093
R10549 gnd.n5526 gnd.n806 7.01093
R10550 gnd.n5943 gnd.n817 7.01093
R10551 gnd.n5544 gnd.n5543 7.01093
R10552 gnd.n5937 gnd.n5936 7.01093
R10553 gnd.n4634 gnd.n828 7.01093
R10554 gnd.n5930 gnd.n839 7.01093
R10555 gnd.n5929 gnd.n842 7.01093
R10556 gnd.n5822 gnd.n5821 7.01093
R10557 gnd.n5923 gnd.n5922 7.01093
R10558 gnd.n863 gnd.n853 7.01093
R10559 gnd.n3261 gnd.t80 7.01093
R10560 gnd.t99 gnd.n3368 7.01093
R10561 gnd.n3872 gnd.t171 7.01093
R10562 gnd.n4857 gnd.t94 6.69227
R10563 gnd.n5417 gnd.t261 6.69227
R10564 gnd.n5944 gnd.t27 6.69227
R10565 gnd.t19 gnd.n1128 6.69227
R10566 gnd.n2994 gnd.t275 6.69227
R10567 gnd.n3806 gnd.t242 6.69227
R10568 gnd.n4005 gnd.t5 6.69227
R10569 gnd.n3707 gnd.n3706 6.5566
R10570 gnd.n2825 gnd.n2824 6.5566
R10571 gnd.n2693 gnd.n2687 6.5566
R10572 gnd.n3619 gnd.n3618 6.5566
R10573 gnd.n3017 gnd.n2953 6.37362
R10574 gnd.n3080 gnd.n1904 6.37362
R10575 gnd.n3190 gnd.n3127 6.37362
R10576 gnd.n3424 gnd.n1757 6.37362
R10577 gnd.n3767 gnd.n3473 6.37362
R10578 gnd.n3830 gnd.n1685 6.37362
R10579 gnd.t115 gnd.n1658 6.37362
R10580 gnd.n2893 gnd.n2891 6.20656
R10581 gnd.n6927 gnd.n6924 6.20656
R10582 gnd.n4538 gnd.n4537 6.20656
R10583 gnd.n3902 gnd.n3899 6.20656
R10584 gnd.n5310 gnd.t277 6.05496
R10585 gnd.n5309 gnd.t283 6.05496
R10586 gnd.t17 gnd.n4782 6.05496
R10587 gnd.t284 gnd.n4673 6.05496
R10588 gnd.t105 gnd.n1085 6.05496
R10589 gnd.n4060 gnd.t29 6.05496
R10590 gnd.n5803 gnd.n5773 5.81868
R10591 gnd.n5771 gnd.n5741 5.81868
R10592 gnd.n5739 gnd.n5709 5.81868
R10593 gnd.n5708 gnd.n5678 5.81868
R10594 gnd.n5676 gnd.n5646 5.81868
R10595 gnd.n5644 gnd.n5614 5.81868
R10596 gnd.n5612 gnd.n5582 5.81868
R10597 gnd.n5581 gnd.n5551 5.81868
R10598 gnd.n3032 gnd.t129 5.73631
R10599 gnd.t110 gnd.n1889 5.73631
R10600 gnd.t31 gnd.n1837 5.73631
R10601 gnd.n3352 gnd.t255 5.73631
R10602 gnd.n3782 gnd.t74 5.73631
R10603 gnd.n3716 gnd.t171 5.73631
R10604 gnd.n3711 gnd.n1331 5.62001
R10605 gnd.n2832 gnd.n2626 5.62001
R10606 gnd.n2832 gnd.n2627 5.62001
R10607 gnd.n3623 gnd.n1331 5.62001
R10608 gnd.n4994 gnd.n4993 5.4308
R10609 gnd.n5836 gnd.n4625 5.4308
R10610 gnd.n4771 gnd.t285 5.41765
R10611 gnd.t85 gnd.n5406 5.41765
R10612 gnd.n5490 gnd.t100 5.41765
R10613 gnd.t102 gnd.n1049 5.41765
R10614 gnd.t2 gnd.n1865 5.41765
R10615 gnd.n3451 gnd.t39 5.41765
R10616 gnd.n4114 gnd.t44 5.41765
R10617 gnd.n4457 gnd.n1013 5.09899
R10618 gnd.n2471 gnd.n1016 5.09899
R10619 gnd.n4451 gnd.n1024 5.09899
R10620 gnd.n2326 gnd.n1027 5.09899
R10621 gnd.n2480 gnd.n2325 5.09899
R10622 gnd.n4443 gnd.n1035 5.09899
R10623 gnd.n2488 gnd.n1038 5.09899
R10624 gnd.n4437 gnd.n1049 5.09899
R10625 gnd.n2496 gnd.n1052 5.09899
R10626 gnd.n4430 gnd.n1057 5.09899
R10627 gnd.n2504 gnd.n2214 5.09899
R10628 gnd.n4424 gnd.n1066 5.09899
R10629 gnd.n4417 gnd.n1074 5.09899
R10630 gnd.n2520 gnd.n1077 5.09899
R10631 gnd.n4411 gnd.n1085 5.09899
R10632 gnd.n2528 gnd.n1088 5.09899
R10633 gnd.n4405 gnd.n1096 5.09899
R10634 gnd.n2536 gnd.n2201 5.09899
R10635 gnd.n4399 gnd.n1106 5.09899
R10636 gnd.n4393 gnd.n1117 5.09899
R10637 gnd.n2552 gnd.n1120 5.09899
R10638 gnd.n4387 gnd.n1128 5.09899
R10639 gnd.n2560 gnd.n1131 5.09899
R10640 gnd.n4381 gnd.n1139 5.09899
R10641 gnd.n2569 gnd.n1142 5.09899
R10642 gnd.n4375 gnd.n1150 5.09899
R10643 gnd.n2577 gnd.n2184 5.09899
R10644 gnd.n4369 gnd.n1159 5.09899
R10645 gnd.n3072 gnd.n1912 5.09899
R10646 gnd.n3010 gnd.n3009 5.09899
R10647 gnd.t233 gnd.n3197 5.09899
R10648 gnd.n3245 gnd.n1838 5.09899
R10649 gnd.n3183 gnd.n3182 5.09899
R10650 gnd.n3416 gnd.n1764 5.09899
R10651 gnd.n3354 gnd.n3353 5.09899
R10652 gnd.n3432 gnd.t286 5.09899
R10653 gnd.n3822 gnd.n1692 5.09899
R10654 gnd.n3760 gnd.n3759 5.09899
R10655 gnd.n4153 gnd.n1364 5.09899
R10656 gnd.n3974 gnd.n3973 5.09899
R10657 gnd.n3956 gnd.n1495 5.09899
R10658 gnd.n3984 gnd.n1497 5.09899
R10659 gnd.n3995 gnd.n1487 5.09899
R10660 gnd.n3994 gnd.n1478 5.09899
R10661 gnd.n4006 gnd.n4005 5.09899
R10662 gnd.n3946 gnd.n1469 5.09899
R10663 gnd.n4016 gnd.n1471 5.09899
R10664 gnd.n4025 gnd.n1453 5.09899
R10665 gnd.n4040 gnd.n4039 5.09899
R10666 gnd.n3936 gnd.n1443 5.09899
R10667 gnd.n4051 gnd.n1445 5.09899
R10668 gnd.n4060 gnd.n1437 5.09899
R10669 gnd.n4059 gnd.n1420 5.09899
R10670 gnd.n4077 gnd.n1415 5.09899
R10671 gnd.n4071 gnd.n1406 5.09899
R10672 gnd.n4091 gnd.n4090 5.09899
R10673 gnd.n4100 gnd.n1402 5.09899
R10674 gnd.n4099 gnd.n1397 5.09899
R10675 gnd.n4115 gnd.n4114 5.09899
R10676 gnd.n6739 gnd.n229 5.09899
R10677 gnd.n6744 gnd.n231 5.09899
R10678 gnd.n6733 gnd.n221 5.09899
R10679 gnd.n6752 gnd.n223 5.09899
R10680 gnd.n6728 gnd.n6727 5.09899
R10681 gnd.n6760 gnd.n209 5.09899
R10682 gnd.n268 gnd.n201 5.09899
R10683 gnd.n5801 gnd.n5800 5.04292
R10684 gnd.n5769 gnd.n5768 5.04292
R10685 gnd.n5737 gnd.n5736 5.04292
R10686 gnd.n5706 gnd.n5705 5.04292
R10687 gnd.n5674 gnd.n5673 5.04292
R10688 gnd.n5642 gnd.n5641 5.04292
R10689 gnd.n5610 gnd.n5609 5.04292
R10690 gnd.n5579 gnd.n5578 5.04292
R10691 gnd.n4765 gnd.n4764 4.82753
R10692 gnd.n50 gnd.n49 4.82753
R10693 gnd.t82 gnd.n5332 4.78034
R10694 gnd.n5448 gnd.t81 4.78034
R10695 gnd.t41 gnd.n1069 4.78034
R10696 gnd.n1866 gnd.t2 4.78034
R10697 gnd.t39 gnd.n1718 4.78034
R10698 gnd.n3714 gnd.t136 4.78034
R10699 gnd.n4070 gnd.t7 4.78034
R10700 gnd.n5306 gnd.n5305 4.74817
R10701 gnd.n5301 gnd.n5300 4.74817
R10702 gnd.n5297 gnd.n5296 4.74817
R10703 gnd.n5293 gnd.n4768 4.74817
R10704 gnd.n5305 gnd.n5304 4.74817
R10705 gnd.n5303 gnd.n5301 4.74817
R10706 gnd.n5299 gnd.n5297 4.74817
R10707 gnd.n5295 gnd.n5293 4.74817
R10708 gnd.n4080 gnd.n218 4.74817
R10709 gnd.n4093 gnd.n217 4.74817
R10710 gnd.n4097 gnd.n216 4.74817
R10711 gnd.n6741 gnd.n215 4.74817
R10712 gnd.n219 gnd.n214 4.74817
R10713 gnd.n1419 gnd.n218 4.74817
R10714 gnd.n4079 gnd.n217 4.74817
R10715 gnd.n4094 gnd.n216 4.74817
R10716 gnd.n4096 gnd.n215 4.74817
R10717 gnd.n6742 gnd.n214 4.74817
R10718 gnd.n2323 gnd.n2322 4.74817
R10719 gnd.n2306 gnd.n2234 4.74817
R10720 gnd.n2299 gnd.n2233 4.74817
R10721 gnd.n2295 gnd.n2232 4.74817
R10722 gnd.n2291 gnd.n2231 4.74817
R10723 gnd.n4068 gnd.n4065 4.74817
R10724 gnd.n4066 gnd.n1400 4.74817
R10725 gnd.n4104 gnd.n4103 4.74817
R10726 gnd.n4111 gnd.n4110 4.74817
R10727 gnd.n4106 gnd.n4105 4.74817
R10728 gnd.n4065 gnd.n4064 4.74817
R10729 gnd.n4067 gnd.n4066 4.74817
R10730 gnd.n4103 gnd.n4102 4.74817
R10731 gnd.n4112 gnd.n4111 4.74817
R10732 gnd.n4109 gnd.n4105 4.74817
R10733 gnd.n4447 gnd.n4446 4.74817
R10734 gnd.n1054 gnd.n1033 4.74817
R10735 gnd.n4434 gnd.n4433 4.74817
R10736 gnd.n1071 gnd.n1055 4.74817
R10737 gnd.n4421 gnd.n4420 4.74817
R10738 gnd.n4448 gnd.n4447 4.74817
R10739 gnd.n4445 gnd.n1033 4.74817
R10740 gnd.n4435 gnd.n4434 4.74817
R10741 gnd.n4432 gnd.n1055 4.74817
R10742 gnd.n4422 gnd.n4421 4.74817
R10743 gnd.n2322 gnd.n2229 4.74817
R10744 gnd.n2306 gnd.n2305 4.74817
R10745 gnd.n2301 gnd.n2233 4.74817
R10746 gnd.n2298 gnd.n2232 4.74817
R10747 gnd.n2294 gnd.n2231 4.74817
R10748 gnd.n4753 gnd.n4752 4.7074
R10749 gnd.n38 gnd.n37 4.7074
R10750 gnd.n4765 gnd.n4753 4.65959
R10751 gnd.n50 gnd.n38 4.65959
R10752 gnd.n4197 gnd.n1333 4.6132
R10753 gnd.n2833 gnd.n2625 4.6132
R10754 gnd.n2862 gnd.n2018 4.46168
R10755 gnd.n3025 gnd.t1 4.46168
R10756 gnd.t47 gnd.n1679 4.46168
R10757 gnd.n4229 gnd.n1311 4.46168
R10758 gnd.n3533 gnd.n3520 4.46111
R10759 gnd.n5786 gnd.n5782 4.38594
R10760 gnd.n5754 gnd.n5750 4.38594
R10761 gnd.n5722 gnd.n5718 4.38594
R10762 gnd.n5691 gnd.n5687 4.38594
R10763 gnd.n5659 gnd.n5655 4.38594
R10764 gnd.n5627 gnd.n5623 4.38594
R10765 gnd.n5595 gnd.n5591 4.38594
R10766 gnd.n5564 gnd.n5560 4.38594
R10767 gnd.n5797 gnd.n5775 4.26717
R10768 gnd.n5765 gnd.n5743 4.26717
R10769 gnd.n5733 gnd.n5711 4.26717
R10770 gnd.n5702 gnd.n5680 4.26717
R10771 gnd.n5670 gnd.n5648 4.26717
R10772 gnd.n5638 gnd.n5616 4.26717
R10773 gnd.n5606 gnd.n5584 4.26717
R10774 gnd.n5575 gnd.n5553 4.26717
R10775 gnd.t28 gnd.n5263 4.14303
R10776 gnd.n5513 gnd.t83 4.14303
R10777 gnd.t76 gnd.n1109 4.14303
R10778 gnd.n3141 gnd.t49 4.14303
R10779 gnd.n3361 gnd.t288 4.14303
R10780 gnd.n4026 gnd.t61 4.14303
R10781 gnd.n5805 gnd.n5804 4.08274
R10782 gnd.n3706 gnd.n3705 4.05904
R10783 gnd.n2824 gnd.n2823 4.05904
R10784 gnd.n2697 gnd.n2687 4.05904
R10785 gnd.n3618 gnd.n3617 4.05904
R10786 gnd.n15 gnd.n7 3.99943
R10787 gnd.n5951 gnd.n804 3.82437
R10788 gnd.t213 gnd.n1932 3.82437
R10789 gnd.n3064 gnd.n1919 3.82437
R10790 gnd.n3002 gnd.n2968 3.82437
R10791 gnd.n3237 gnd.n1844 3.82437
R10792 gnd.n3175 gnd.n3143 3.82437
R10793 gnd.n3408 gnd.n1772 3.82437
R10794 gnd.n3346 gnd.n3314 3.82437
R10795 gnd.n3814 gnd.n1699 3.82437
R10796 gnd.n3752 gnd.n3489 3.82437
R10797 gnd.n3883 gnd.t136 3.82437
R10798 gnd.n5805 gnd.n5677 3.70378
R10799 gnd.n4767 gnd.n4766 3.65935
R10800 gnd.n15 gnd.n14 3.60163
R10801 gnd.n5796 gnd.n5777 3.49141
R10802 gnd.n5764 gnd.n5745 3.49141
R10803 gnd.n5732 gnd.n5713 3.49141
R10804 gnd.n5701 gnd.n5682 3.49141
R10805 gnd.n5669 gnd.n5650 3.49141
R10806 gnd.n5637 gnd.n5618 3.49141
R10807 gnd.n5605 gnd.n5586 3.49141
R10808 gnd.n5574 gnd.n5555 3.49141
R10809 gnd.n5951 gnd.n5950 3.18706
R10810 gnd.n1951 gnd.t129 3.18706
R10811 gnd.n3729 gnd.t187 3.18706
R10812 gnd.n5264 gnd.t28 2.8684
R10813 gnd.n4754 gnd.t10 2.82907
R10814 gnd.n4754 gnd.t88 2.82907
R10815 gnd.n4756 gnd.t279 2.82907
R10816 gnd.n4756 gnd.t258 2.82907
R10817 gnd.n4758 gnd.t103 2.82907
R10818 gnd.n4758 gnd.t71 2.82907
R10819 gnd.n4760 gnd.t272 2.82907
R10820 gnd.n4760 gnd.t90 2.82907
R10821 gnd.n4762 gnd.t259 2.82907
R10822 gnd.n4762 gnd.t33 2.82907
R10823 gnd.n4731 gnd.t223 2.82907
R10824 gnd.n4731 gnd.t290 2.82907
R10825 gnd.n4733 gnd.t75 2.82907
R10826 gnd.n4733 gnd.t106 2.82907
R10827 gnd.n4735 gnd.t112 2.82907
R10828 gnd.n4735 gnd.t72 2.82907
R10829 gnd.n4737 gnd.t14 2.82907
R10830 gnd.n4737 gnd.t56 2.82907
R10831 gnd.n4739 gnd.t59 2.82907
R10832 gnd.n4739 gnd.t91 2.82907
R10833 gnd.n4742 gnd.t43 2.82907
R10834 gnd.n4742 gnd.t77 2.82907
R10835 gnd.n4744 gnd.t42 2.82907
R10836 gnd.n4744 gnd.t281 2.82907
R10837 gnd.n4746 gnd.t280 2.82907
R10838 gnd.n4746 gnd.t235 2.82907
R10839 gnd.n4748 gnd.t48 2.82907
R10840 gnd.n4748 gnd.t268 2.82907
R10841 gnd.n4750 gnd.t104 2.82907
R10842 gnd.n4750 gnd.t113 2.82907
R10843 gnd.n47 gnd.t69 2.82907
R10844 gnd.n47 gnd.t227 2.82907
R10845 gnd.n45 gnd.t89 2.82907
R10846 gnd.n45 gnd.t282 2.82907
R10847 gnd.n43 gnd.t257 2.82907
R10848 gnd.n43 gnd.t53 2.82907
R10849 gnd.n41 gnd.t73 2.82907
R10850 gnd.n41 gnd.t46 2.82907
R10851 gnd.n39 gnd.t256 2.82907
R10852 gnd.n39 gnd.t266 2.82907
R10853 gnd.n24 gnd.t237 2.82907
R10854 gnd.n24 gnd.t287 2.82907
R10855 gnd.n22 gnd.t87 2.82907
R10856 gnd.n22 gnd.t248 2.82907
R10857 gnd.n20 gnd.t111 2.82907
R10858 gnd.n20 gnd.t45 2.82907
R10859 gnd.n18 gnd.t60 2.82907
R10860 gnd.n18 gnd.t267 2.82907
R10861 gnd.n16 gnd.t62 2.82907
R10862 gnd.n16 gnd.t92 2.82907
R10863 gnd.n35 gnd.t24 2.82907
R10864 gnd.n35 gnd.t26 2.82907
R10865 gnd.n33 gnd.t98 2.82907
R10866 gnd.n33 gnd.t247 2.82907
R10867 gnd.n31 gnd.t52 2.82907
R10868 gnd.n31 gnd.t63 2.82907
R10869 gnd.n29 gnd.t30 2.82907
R10870 gnd.n29 gnd.t8 2.82907
R10871 gnd.n27 gnd.t95 2.82907
R10872 gnd.n27 gnd.t12 2.82907
R10873 gnd.n5793 gnd.n5792 2.71565
R10874 gnd.n5761 gnd.n5760 2.71565
R10875 gnd.n5729 gnd.n5728 2.71565
R10876 gnd.n5698 gnd.n5697 2.71565
R10877 gnd.n5666 gnd.n5665 2.71565
R10878 gnd.n5634 gnd.n5633 2.71565
R10879 gnd.n5602 gnd.n5601 2.71565
R10880 gnd.n5571 gnd.n5570 2.71565
R10881 gnd.n3056 gnd.n1926 2.54975
R10882 gnd.n2953 gnd.t254 2.54975
R10883 gnd.n2995 gnd.n2994 2.54975
R10884 gnd.n3213 gnd.t34 2.54975
R10885 gnd.n3229 gnd.n1851 2.54975
R10886 gnd.n3198 gnd.t233 2.54975
R10887 gnd.n3168 gnd.n3167 2.54975
R10888 gnd.n3400 gnd.n1779 2.54975
R10889 gnd.n3340 gnd.t286 2.54975
R10890 gnd.n3339 gnd.n3338 2.54975
R10891 gnd.n3790 gnd.t96 2.54975
R10892 gnd.n3806 gnd.n1705 2.54975
R10893 gnd.n3830 gnd.t97 2.54975
R10894 gnd.n3745 gnd.n3744 2.54975
R10895 gnd.n5305 gnd.n4767 2.27742
R10896 gnd.n5301 gnd.n4767 2.27742
R10897 gnd.n5297 gnd.n4767 2.27742
R10898 gnd.n5293 gnd.n4767 2.27742
R10899 gnd.n6755 gnd.n218 2.27742
R10900 gnd.n6755 gnd.n217 2.27742
R10901 gnd.n6755 gnd.n216 2.27742
R10902 gnd.n6755 gnd.n215 2.27742
R10903 gnd.n6755 gnd.n214 2.27742
R10904 gnd.n4065 gnd.n213 2.27742
R10905 gnd.n4066 gnd.n213 2.27742
R10906 gnd.n4103 gnd.n213 2.27742
R10907 gnd.n4111 gnd.n213 2.27742
R10908 gnd.n4105 gnd.n213 2.27742
R10909 gnd.n4447 gnd.n1031 2.27742
R10910 gnd.n1033 gnd.n1031 2.27742
R10911 gnd.n4434 gnd.n1031 2.27742
R10912 gnd.n1055 gnd.n1031 2.27742
R10913 gnd.n4421 gnd.n1031 2.27742
R10914 gnd.n2322 gnd.n2321 2.27742
R10915 gnd.n2321 gnd.n2306 2.27742
R10916 gnd.n2321 gnd.n2233 2.27742
R10917 gnd.n2321 gnd.n2232 2.27742
R10918 gnd.n2321 gnd.n2231 2.27742
R10919 gnd.t125 gnd.n5185 2.23109
R10920 gnd.n5333 gnd.t82 2.23109
R10921 gnd.n3253 gnd.t49 2.23109
R10922 gnd.t288 gnd.n3299 2.23109
R10923 gnd.n5789 gnd.n5779 1.93989
R10924 gnd.n5757 gnd.n5747 1.93989
R10925 gnd.n5725 gnd.n5715 1.93989
R10926 gnd.n5694 gnd.n5684 1.93989
R10927 gnd.n5662 gnd.n5652 1.93989
R10928 gnd.n5630 gnd.n5620 1.93989
R10929 gnd.n5598 gnd.n5588 1.93989
R10930 gnd.n5567 gnd.n5557 1.93989
R10931 gnd.n5198 gnd.t37 1.59378
R10932 gnd.n5407 gnd.t85 1.59378
R10933 gnd.n5478 gnd.t100 1.59378
R10934 gnd.n2757 gnd.t122 1.27512
R10935 gnd.n2757 gnd.n2647 1.27512
R10936 gnd.n3048 gnd.n1933 1.27512
R10937 gnd.n2987 gnd.n2981 1.27512
R10938 gnd.n3221 gnd.n1858 1.27512
R10939 gnd.n3160 gnd.n1810 1.27512
R10940 gnd.n3392 gnd.n1787 1.27512
R10941 gnd.n3331 gnd.n1733 1.27512
R10942 gnd.n3798 gnd.n1712 1.27512
R10943 gnd.n3736 gnd.n3501 1.27512
R10944 gnd.n3722 gnd.n3515 1.27512
R10945 gnd.n4995 gnd.n4994 1.16414
R10946 gnd.n5839 gnd.n4625 1.16414
R10947 gnd.n5788 gnd.n5781 1.16414
R10948 gnd.n5756 gnd.n5749 1.16414
R10949 gnd.n5724 gnd.n5717 1.16414
R10950 gnd.n5693 gnd.n5686 1.16414
R10951 gnd.n5661 gnd.n5654 1.16414
R10952 gnd.n5629 gnd.n5622 1.16414
R10953 gnd.n5597 gnd.n5590 1.16414
R10954 gnd.n5566 gnd.n5559 1.16414
R10955 gnd.n4197 gnd.n4196 0.970197
R10956 gnd.n2833 gnd.n2157 0.970197
R10957 gnd.n5772 gnd.n5740 0.962709
R10958 gnd.n5804 gnd.n5772 0.962709
R10959 gnd.n5645 gnd.n5613 0.962709
R10960 gnd.n5677 gnd.n5645 0.962709
R10961 gnd.t277 gnd.n5309 0.956468
R10962 gnd.n4680 gnd.t284 0.956468
R10963 gnd.n4469 gnd.t58 0.956468
R10964 gnd.n4463 gnd.n1005 0.956468
R10965 gnd.n2544 gnd.t76 0.956468
R10966 gnd.n2936 gnd.t244 0.956468
R10967 gnd.n3056 gnd.t228 0.956468
R10968 gnd.n3744 gnd.t64 0.956468
R10969 gnd.t230 gnd.n1657 0.956468
R10970 gnd.n3942 gnd.t61 0.956468
R10971 gnd.n6720 gnd.n194 0.956468
R10972 gnd.t25 gnd.n186 0.956468
R10973 gnd.n4761 gnd.n4759 0.773756
R10974 gnd.n46 gnd.n44 0.773756
R10975 gnd.n4764 gnd.n4763 0.773756
R10976 gnd.n4763 gnd.n4761 0.773756
R10977 gnd.n4759 gnd.n4757 0.773756
R10978 gnd.n4757 gnd.n4755 0.773756
R10979 gnd.n42 gnd.n40 0.773756
R10980 gnd.n44 gnd.n42 0.773756
R10981 gnd.n48 gnd.n46 0.773756
R10982 gnd.n49 gnd.n48 0.773756
R10983 gnd.n2 gnd.n1 0.672012
R10984 gnd.n3 gnd.n2 0.672012
R10985 gnd.n4 gnd.n3 0.672012
R10986 gnd.n5 gnd.n4 0.672012
R10987 gnd.n6 gnd.n5 0.672012
R10988 gnd.n7 gnd.n6 0.672012
R10989 gnd.n9 gnd.n8 0.672012
R10990 gnd.n10 gnd.n9 0.672012
R10991 gnd.n11 gnd.n10 0.672012
R10992 gnd.n12 gnd.n11 0.672012
R10993 gnd.n13 gnd.n12 0.672012
R10994 gnd.n14 gnd.n13 0.672012
R10995 gnd.n3040 gnd.t157 0.637812
R10996 gnd.n3008 gnd.t4 0.637812
R10997 gnd.n3169 gnd.t80 0.637812
R10998 gnd.n3369 gnd.t99 0.637812
R10999 gnd.t226 gnd.n1691 0.637812
R11000 gnd.n3729 gnd.t143 0.637812
R11001 gnd.n4741 gnd.n4740 0.573776
R11002 gnd.n4740 gnd.n4738 0.573776
R11003 gnd.n4738 gnd.n4736 0.573776
R11004 gnd.n4736 gnd.n4734 0.573776
R11005 gnd.n4734 gnd.n4732 0.573776
R11006 gnd.n4752 gnd.n4751 0.573776
R11007 gnd.n4751 gnd.n4749 0.573776
R11008 gnd.n4749 gnd.n4747 0.573776
R11009 gnd.n4747 gnd.n4745 0.573776
R11010 gnd.n4745 gnd.n4743 0.573776
R11011 gnd.n19 gnd.n17 0.573776
R11012 gnd.n21 gnd.n19 0.573776
R11013 gnd.n23 gnd.n21 0.573776
R11014 gnd.n25 gnd.n23 0.573776
R11015 gnd.n26 gnd.n25 0.573776
R11016 gnd.n30 gnd.n28 0.573776
R11017 gnd.n32 gnd.n30 0.573776
R11018 gnd.n34 gnd.n32 0.573776
R11019 gnd.n36 gnd.n34 0.573776
R11020 gnd.n37 gnd.n36 0.573776
R11021 gnd gnd.n0 0.551497
R11022 gnd.n6755 gnd.n213 0.548625
R11023 gnd.n2321 gnd.n1031 0.548625
R11024 gnd.n2383 gnd.n2381 0.532512
R11025 gnd.n2421 gnd.n2420 0.532512
R11026 gnd.n6865 gnd.n6864 0.532512
R11027 gnd.n6965 gnd.n78 0.532512
R11028 gnd.n4364 gnd.n4363 0.523366
R11029 gnd.n1549 gnd.n1270 0.523366
R11030 gnd.n6959 gnd.n6958 0.520317
R11031 gnd.n6888 gnd.n6887 0.520317
R11032 gnd.n4157 gnd.n1359 0.520317
R11033 gnd.n1501 gnd.n1315 0.520317
R11034 gnd.n2141 gnd.n1157 0.520317
R11035 gnd.n2582 gnd.n2581 0.520317
R11036 gnd.n4498 gnd.n953 0.520317
R11037 gnd.n2430 gnd.n910 0.520317
R11038 gnd.n3889 gnd.n3888 0.489829
R11039 gnd.n2911 gnd.n1976 0.489829
R11040 gnd.n5827 gnd.n4629 0.486781
R11041 gnd.n5047 gnd.n4943 0.48678
R11042 gnd.n5918 gnd.n5917 0.480683
R11043 gnd.n5115 gnd.n4893 0.480683
R11044 gnd.n6998 gnd.n6997 0.470187
R11045 gnd.n639 gnd.n634 0.459342
R11046 gnd.n6507 gnd.n6506 0.459342
R11047 gnd.n6718 gnd.n278 0.459342
R11048 gnd.n2313 gnd.n2312 0.459342
R11049 gnd.n4366 gnd.n4365 0.432431
R11050 gnd.n4150 gnd.n1368 0.432431
R11051 gnd.n2891 gnd.n2890 0.388379
R11052 gnd.n5785 gnd.n5784 0.388379
R11053 gnd.n5753 gnd.n5752 0.388379
R11054 gnd.n5721 gnd.n5720 0.388379
R11055 gnd.n5690 gnd.n5689 0.388379
R11056 gnd.n5658 gnd.n5657 0.388379
R11057 gnd.n5626 gnd.n5625 0.388379
R11058 gnd.n5594 gnd.n5593 0.388379
R11059 gnd.n5563 gnd.n5562 0.388379
R11060 gnd.n6928 gnd.n6927 0.388379
R11061 gnd.n4539 gnd.n4538 0.388379
R11062 gnd.n3903 gnd.n3902 0.388379
R11063 gnd.n6998 gnd.n15 0.374463
R11064 gnd.n5527 gnd.t27 0.319156
R11065 gnd.n2480 gnd.t55 0.319156
R11066 gnd.n2512 gnd.t41 0.319156
R11067 gnd.n3196 gnd.t224 0.319156
R11068 gnd.t108 gnd.t107 0.319156
R11069 gnd.t54 gnd.t238 0.319156
R11070 gnd.t66 gnd.n1750 0.319156
R11071 gnd.n4082 gnd.t7 0.319156
R11072 gnd.n6733 gnd.t86 0.319156
R11073 gnd.n5041 gnd.n5040 0.311721
R11074 gnd.n2875 gnd.n2008 0.302329
R11075 gnd.n3913 gnd.n3912 0.302329
R11076 gnd gnd.n6998 0.295112
R11077 gnd.n5884 gnd.n5883 0.268793
R11078 gnd.n5883 gnd.n5882 0.241354
R11079 gnd.n1333 gnd.n1330 0.229039
R11080 gnd.n1336 gnd.n1333 0.229039
R11081 gnd.n2625 gnd.n2156 0.229039
R11082 gnd.n2625 gnd.n2624 0.229039
R11083 gnd.n5170 gnd.n4911 0.206293
R11084 gnd.n5802 gnd.n5774 0.155672
R11085 gnd.n5795 gnd.n5774 0.155672
R11086 gnd.n5795 gnd.n5794 0.155672
R11087 gnd.n5794 gnd.n5778 0.155672
R11088 gnd.n5787 gnd.n5778 0.155672
R11089 gnd.n5787 gnd.n5786 0.155672
R11090 gnd.n5770 gnd.n5742 0.155672
R11091 gnd.n5763 gnd.n5742 0.155672
R11092 gnd.n5763 gnd.n5762 0.155672
R11093 gnd.n5762 gnd.n5746 0.155672
R11094 gnd.n5755 gnd.n5746 0.155672
R11095 gnd.n5755 gnd.n5754 0.155672
R11096 gnd.n5738 gnd.n5710 0.155672
R11097 gnd.n5731 gnd.n5710 0.155672
R11098 gnd.n5731 gnd.n5730 0.155672
R11099 gnd.n5730 gnd.n5714 0.155672
R11100 gnd.n5723 gnd.n5714 0.155672
R11101 gnd.n5723 gnd.n5722 0.155672
R11102 gnd.n5707 gnd.n5679 0.155672
R11103 gnd.n5700 gnd.n5679 0.155672
R11104 gnd.n5700 gnd.n5699 0.155672
R11105 gnd.n5699 gnd.n5683 0.155672
R11106 gnd.n5692 gnd.n5683 0.155672
R11107 gnd.n5692 gnd.n5691 0.155672
R11108 gnd.n5675 gnd.n5647 0.155672
R11109 gnd.n5668 gnd.n5647 0.155672
R11110 gnd.n5668 gnd.n5667 0.155672
R11111 gnd.n5667 gnd.n5651 0.155672
R11112 gnd.n5660 gnd.n5651 0.155672
R11113 gnd.n5660 gnd.n5659 0.155672
R11114 gnd.n5643 gnd.n5615 0.155672
R11115 gnd.n5636 gnd.n5615 0.155672
R11116 gnd.n5636 gnd.n5635 0.155672
R11117 gnd.n5635 gnd.n5619 0.155672
R11118 gnd.n5628 gnd.n5619 0.155672
R11119 gnd.n5628 gnd.n5627 0.155672
R11120 gnd.n5611 gnd.n5583 0.155672
R11121 gnd.n5604 gnd.n5583 0.155672
R11122 gnd.n5604 gnd.n5603 0.155672
R11123 gnd.n5603 gnd.n5587 0.155672
R11124 gnd.n5596 gnd.n5587 0.155672
R11125 gnd.n5596 gnd.n5595 0.155672
R11126 gnd.n5580 gnd.n5552 0.155672
R11127 gnd.n5573 gnd.n5552 0.155672
R11128 gnd.n5573 gnd.n5572 0.155672
R11129 gnd.n5572 gnd.n5556 0.155672
R11130 gnd.n5565 gnd.n5556 0.155672
R11131 gnd.n5565 gnd.n5564 0.155672
R11132 gnd.n5917 gnd.n860 0.152939
R11133 gnd.n4583 gnd.n860 0.152939
R11134 gnd.n4584 gnd.n4583 0.152939
R11135 gnd.n4585 gnd.n4584 0.152939
R11136 gnd.n4586 gnd.n4585 0.152939
R11137 gnd.n4587 gnd.n4586 0.152939
R11138 gnd.n4588 gnd.n4587 0.152939
R11139 gnd.n4589 gnd.n4588 0.152939
R11140 gnd.n4590 gnd.n4589 0.152939
R11141 gnd.n4591 gnd.n4590 0.152939
R11142 gnd.n4592 gnd.n4591 0.152939
R11143 gnd.n4593 gnd.n4592 0.152939
R11144 gnd.n4594 gnd.n4593 0.152939
R11145 gnd.n4595 gnd.n4594 0.152939
R11146 gnd.n5885 gnd.n4595 0.152939
R11147 gnd.n5885 gnd.n5884 0.152939
R11148 gnd.n5189 gnd.n4893 0.152939
R11149 gnd.n5190 gnd.n5189 0.152939
R11150 gnd.n5191 gnd.n5190 0.152939
R11151 gnd.n5191 gnd.n4872 0.152939
R11152 gnd.n5219 gnd.n4872 0.152939
R11153 gnd.n5220 gnd.n5219 0.152939
R11154 gnd.n5221 gnd.n5220 0.152939
R11155 gnd.n5222 gnd.n5221 0.152939
R11156 gnd.n5222 gnd.n4846 0.152939
R11157 gnd.n5253 gnd.n4846 0.152939
R11158 gnd.n5254 gnd.n5253 0.152939
R11159 gnd.n5255 gnd.n5254 0.152939
R11160 gnd.n5256 gnd.n5255 0.152939
R11161 gnd.n5257 gnd.n5256 0.152939
R11162 gnd.n5257 gnd.n4813 0.152939
R11163 gnd.n5314 gnd.n4813 0.152939
R11164 gnd.n5315 gnd.n5314 0.152939
R11165 gnd.n5316 gnd.n5315 0.152939
R11166 gnd.n5317 gnd.n5316 0.152939
R11167 gnd.n5317 gnd.n4786 0.152939
R11168 gnd.n5354 gnd.n4786 0.152939
R11169 gnd.n5355 gnd.n5354 0.152939
R11170 gnd.n5356 gnd.n5355 0.152939
R11171 gnd.n5357 gnd.n5356 0.152939
R11172 gnd.n5357 gnd.n4723 0.152939
R11173 gnd.n5399 gnd.n4723 0.152939
R11174 gnd.n5400 gnd.n5399 0.152939
R11175 gnd.n5401 gnd.n5400 0.152939
R11176 gnd.n5402 gnd.n5401 0.152939
R11177 gnd.n5402 gnd.n4695 0.152939
R11178 gnd.n5438 gnd.n4695 0.152939
R11179 gnd.n5439 gnd.n5438 0.152939
R11180 gnd.n5440 gnd.n5439 0.152939
R11181 gnd.n5441 gnd.n5440 0.152939
R11182 gnd.n5442 gnd.n5441 0.152939
R11183 gnd.n5442 gnd.n4664 0.152939
R11184 gnd.n5493 gnd.n4664 0.152939
R11185 gnd.n5494 gnd.n5493 0.152939
R11186 gnd.n5495 gnd.n5494 0.152939
R11187 gnd.n5497 gnd.n5495 0.152939
R11188 gnd.n5497 gnd.n5496 0.152939
R11189 gnd.n5496 gnd.n810 0.152939
R11190 gnd.n811 gnd.n810 0.152939
R11191 gnd.n812 gnd.n811 0.152939
R11192 gnd.n832 gnd.n812 0.152939
R11193 gnd.n833 gnd.n832 0.152939
R11194 gnd.n834 gnd.n833 0.152939
R11195 gnd.n835 gnd.n834 0.152939
R11196 gnd.n836 gnd.n835 0.152939
R11197 gnd.n857 gnd.n836 0.152939
R11198 gnd.n858 gnd.n857 0.152939
R11199 gnd.n859 gnd.n858 0.152939
R11200 gnd.n5918 gnd.n859 0.152939
R11201 gnd.n5116 gnd.n5115 0.152939
R11202 gnd.n5117 gnd.n5116 0.152939
R11203 gnd.n5118 gnd.n5117 0.152939
R11204 gnd.n5119 gnd.n5118 0.152939
R11205 gnd.n5120 gnd.n5119 0.152939
R11206 gnd.n5121 gnd.n5120 0.152939
R11207 gnd.n5122 gnd.n5121 0.152939
R11208 gnd.n5123 gnd.n5122 0.152939
R11209 gnd.n5124 gnd.n5123 0.152939
R11210 gnd.n5125 gnd.n5124 0.152939
R11211 gnd.n5126 gnd.n5125 0.152939
R11212 gnd.n5127 gnd.n5126 0.152939
R11213 gnd.n5128 gnd.n5127 0.152939
R11214 gnd.n5129 gnd.n5128 0.152939
R11215 gnd.n5133 gnd.n5129 0.152939
R11216 gnd.n5133 gnd.n4911 0.152939
R11217 gnd.n5882 gnd.n4600 0.152939
R11218 gnd.n4602 gnd.n4600 0.152939
R11219 gnd.n4603 gnd.n4602 0.152939
R11220 gnd.n4604 gnd.n4603 0.152939
R11221 gnd.n4605 gnd.n4604 0.152939
R11222 gnd.n4606 gnd.n4605 0.152939
R11223 gnd.n4607 gnd.n4606 0.152939
R11224 gnd.n4608 gnd.n4607 0.152939
R11225 gnd.n4609 gnd.n4608 0.152939
R11226 gnd.n4610 gnd.n4609 0.152939
R11227 gnd.n4611 gnd.n4610 0.152939
R11228 gnd.n4612 gnd.n4611 0.152939
R11229 gnd.n4613 gnd.n4612 0.152939
R11230 gnd.n4614 gnd.n4613 0.152939
R11231 gnd.n4615 gnd.n4614 0.152939
R11232 gnd.n4616 gnd.n4615 0.152939
R11233 gnd.n4617 gnd.n4616 0.152939
R11234 gnd.n4618 gnd.n4617 0.152939
R11235 gnd.n4619 gnd.n4618 0.152939
R11236 gnd.n4620 gnd.n4619 0.152939
R11237 gnd.n4621 gnd.n4620 0.152939
R11238 gnd.n4622 gnd.n4621 0.152939
R11239 gnd.n4626 gnd.n4622 0.152939
R11240 gnd.n4627 gnd.n4626 0.152939
R11241 gnd.n4628 gnd.n4627 0.152939
R11242 gnd.n4629 gnd.n4628 0.152939
R11243 gnd.n5376 gnd.n5375 0.152939
R11244 gnd.n5377 gnd.n5376 0.152939
R11245 gnd.n5378 gnd.n5377 0.152939
R11246 gnd.n5379 gnd.n5378 0.152939
R11247 gnd.n5380 gnd.n5379 0.152939
R11248 gnd.n5381 gnd.n5380 0.152939
R11249 gnd.n5382 gnd.n5381 0.152939
R11250 gnd.n5383 gnd.n5382 0.152939
R11251 gnd.n5383 gnd.n4676 0.152939
R11252 gnd.n5461 gnd.n4676 0.152939
R11253 gnd.n5462 gnd.n5461 0.152939
R11254 gnd.n5463 gnd.n5462 0.152939
R11255 gnd.n5464 gnd.n5463 0.152939
R11256 gnd.n5465 gnd.n5464 0.152939
R11257 gnd.n5466 gnd.n5465 0.152939
R11258 gnd.n5467 gnd.n5466 0.152939
R11259 gnd.n5468 gnd.n5467 0.152939
R11260 gnd.n5468 gnd.n4642 0.152939
R11261 gnd.n5530 gnd.n4642 0.152939
R11262 gnd.n5531 gnd.n5530 0.152939
R11263 gnd.n5532 gnd.n5531 0.152939
R11264 gnd.n5533 gnd.n5532 0.152939
R11265 gnd.n5534 gnd.n5533 0.152939
R11266 gnd.n5535 gnd.n5534 0.152939
R11267 gnd.n5535 gnd.n4631 0.152939
R11268 gnd.n5825 gnd.n4631 0.152939
R11269 gnd.n5826 gnd.n5825 0.152939
R11270 gnd.n5827 gnd.n5826 0.152939
R11271 gnd.n5048 gnd.n5047 0.152939
R11272 gnd.n5049 gnd.n5048 0.152939
R11273 gnd.n5049 gnd.n4931 0.152939
R11274 gnd.n5063 gnd.n4931 0.152939
R11275 gnd.n5064 gnd.n5063 0.152939
R11276 gnd.n5065 gnd.n5064 0.152939
R11277 gnd.n5065 gnd.n4918 0.152939
R11278 gnd.n5079 gnd.n4918 0.152939
R11279 gnd.n5080 gnd.n5079 0.152939
R11280 gnd.n5081 gnd.n5080 0.152939
R11281 gnd.n5082 gnd.n5081 0.152939
R11282 gnd.n5083 gnd.n5082 0.152939
R11283 gnd.n5084 gnd.n5083 0.152939
R11284 gnd.n5085 gnd.n5084 0.152939
R11285 gnd.n5086 gnd.n5085 0.152939
R11286 gnd.n5087 gnd.n5086 0.152939
R11287 gnd.n5088 gnd.n5087 0.152939
R11288 gnd.n5089 gnd.n5088 0.152939
R11289 gnd.n5090 gnd.n5089 0.152939
R11290 gnd.n5090 gnd.n4853 0.152939
R11291 gnd.n5242 gnd.n4853 0.152939
R11292 gnd.n5243 gnd.n5242 0.152939
R11293 gnd.n5244 gnd.n5243 0.152939
R11294 gnd.n5245 gnd.n5244 0.152939
R11295 gnd.n5245 gnd.n4820 0.152939
R11296 gnd.n5289 gnd.n4820 0.152939
R11297 gnd.n5290 gnd.n5289 0.152939
R11298 gnd.n5291 gnd.n5290 0.152939
R11299 gnd.n5040 gnd.n4947 0.152939
R11300 gnd.n4950 gnd.n4947 0.152939
R11301 gnd.n4951 gnd.n4950 0.152939
R11302 gnd.n4952 gnd.n4951 0.152939
R11303 gnd.n4955 gnd.n4952 0.152939
R11304 gnd.n4956 gnd.n4955 0.152939
R11305 gnd.n4957 gnd.n4956 0.152939
R11306 gnd.n4958 gnd.n4957 0.152939
R11307 gnd.n4961 gnd.n4958 0.152939
R11308 gnd.n4962 gnd.n4961 0.152939
R11309 gnd.n4963 gnd.n4962 0.152939
R11310 gnd.n4964 gnd.n4963 0.152939
R11311 gnd.n4967 gnd.n4964 0.152939
R11312 gnd.n4968 gnd.n4967 0.152939
R11313 gnd.n4969 gnd.n4968 0.152939
R11314 gnd.n4970 gnd.n4969 0.152939
R11315 gnd.n4973 gnd.n4970 0.152939
R11316 gnd.n4974 gnd.n4973 0.152939
R11317 gnd.n4975 gnd.n4974 0.152939
R11318 gnd.n4976 gnd.n4975 0.152939
R11319 gnd.n4979 gnd.n4976 0.152939
R11320 gnd.n4980 gnd.n4979 0.152939
R11321 gnd.n4983 gnd.n4980 0.152939
R11322 gnd.n4984 gnd.n4983 0.152939
R11323 gnd.n4986 gnd.n4984 0.152939
R11324 gnd.n4986 gnd.n4943 0.152939
R11325 gnd.n6124 gnd.n634 0.152939
R11326 gnd.n6125 gnd.n6124 0.152939
R11327 gnd.n6126 gnd.n6125 0.152939
R11328 gnd.n6126 gnd.n628 0.152939
R11329 gnd.n6134 gnd.n628 0.152939
R11330 gnd.n6135 gnd.n6134 0.152939
R11331 gnd.n6136 gnd.n6135 0.152939
R11332 gnd.n6136 gnd.n622 0.152939
R11333 gnd.n6144 gnd.n622 0.152939
R11334 gnd.n6145 gnd.n6144 0.152939
R11335 gnd.n6146 gnd.n6145 0.152939
R11336 gnd.n6146 gnd.n616 0.152939
R11337 gnd.n6154 gnd.n616 0.152939
R11338 gnd.n6155 gnd.n6154 0.152939
R11339 gnd.n6156 gnd.n6155 0.152939
R11340 gnd.n6156 gnd.n610 0.152939
R11341 gnd.n6164 gnd.n610 0.152939
R11342 gnd.n6165 gnd.n6164 0.152939
R11343 gnd.n6166 gnd.n6165 0.152939
R11344 gnd.n6166 gnd.n604 0.152939
R11345 gnd.n6174 gnd.n604 0.152939
R11346 gnd.n6175 gnd.n6174 0.152939
R11347 gnd.n6176 gnd.n6175 0.152939
R11348 gnd.n6176 gnd.n598 0.152939
R11349 gnd.n6184 gnd.n598 0.152939
R11350 gnd.n6185 gnd.n6184 0.152939
R11351 gnd.n6186 gnd.n6185 0.152939
R11352 gnd.n6186 gnd.n592 0.152939
R11353 gnd.n6194 gnd.n592 0.152939
R11354 gnd.n6195 gnd.n6194 0.152939
R11355 gnd.n6196 gnd.n6195 0.152939
R11356 gnd.n6196 gnd.n586 0.152939
R11357 gnd.n6204 gnd.n586 0.152939
R11358 gnd.n6205 gnd.n6204 0.152939
R11359 gnd.n6206 gnd.n6205 0.152939
R11360 gnd.n6206 gnd.n580 0.152939
R11361 gnd.n6214 gnd.n580 0.152939
R11362 gnd.n6215 gnd.n6214 0.152939
R11363 gnd.n6216 gnd.n6215 0.152939
R11364 gnd.n6216 gnd.n574 0.152939
R11365 gnd.n6224 gnd.n574 0.152939
R11366 gnd.n6225 gnd.n6224 0.152939
R11367 gnd.n6226 gnd.n6225 0.152939
R11368 gnd.n6226 gnd.n568 0.152939
R11369 gnd.n6234 gnd.n568 0.152939
R11370 gnd.n6235 gnd.n6234 0.152939
R11371 gnd.n6236 gnd.n6235 0.152939
R11372 gnd.n6236 gnd.n562 0.152939
R11373 gnd.n6244 gnd.n562 0.152939
R11374 gnd.n6245 gnd.n6244 0.152939
R11375 gnd.n6246 gnd.n6245 0.152939
R11376 gnd.n6246 gnd.n556 0.152939
R11377 gnd.n6254 gnd.n556 0.152939
R11378 gnd.n6255 gnd.n6254 0.152939
R11379 gnd.n6256 gnd.n6255 0.152939
R11380 gnd.n6256 gnd.n550 0.152939
R11381 gnd.n6264 gnd.n550 0.152939
R11382 gnd.n6265 gnd.n6264 0.152939
R11383 gnd.n6266 gnd.n6265 0.152939
R11384 gnd.n6266 gnd.n544 0.152939
R11385 gnd.n6274 gnd.n544 0.152939
R11386 gnd.n6275 gnd.n6274 0.152939
R11387 gnd.n6276 gnd.n6275 0.152939
R11388 gnd.n6276 gnd.n538 0.152939
R11389 gnd.n6284 gnd.n538 0.152939
R11390 gnd.n6285 gnd.n6284 0.152939
R11391 gnd.n6286 gnd.n6285 0.152939
R11392 gnd.n6286 gnd.n532 0.152939
R11393 gnd.n6294 gnd.n532 0.152939
R11394 gnd.n6295 gnd.n6294 0.152939
R11395 gnd.n6296 gnd.n6295 0.152939
R11396 gnd.n6296 gnd.n526 0.152939
R11397 gnd.n6304 gnd.n526 0.152939
R11398 gnd.n6305 gnd.n6304 0.152939
R11399 gnd.n6306 gnd.n6305 0.152939
R11400 gnd.n6306 gnd.n520 0.152939
R11401 gnd.n6314 gnd.n520 0.152939
R11402 gnd.n6315 gnd.n6314 0.152939
R11403 gnd.n6316 gnd.n6315 0.152939
R11404 gnd.n6316 gnd.n514 0.152939
R11405 gnd.n6324 gnd.n514 0.152939
R11406 gnd.n6325 gnd.n6324 0.152939
R11407 gnd.n6326 gnd.n6325 0.152939
R11408 gnd.n6326 gnd.n508 0.152939
R11409 gnd.n6334 gnd.n508 0.152939
R11410 gnd.n6335 gnd.n6334 0.152939
R11411 gnd.n6336 gnd.n6335 0.152939
R11412 gnd.n6336 gnd.n502 0.152939
R11413 gnd.n6344 gnd.n502 0.152939
R11414 gnd.n6345 gnd.n6344 0.152939
R11415 gnd.n6346 gnd.n6345 0.152939
R11416 gnd.n6346 gnd.n496 0.152939
R11417 gnd.n6354 gnd.n496 0.152939
R11418 gnd.n6355 gnd.n6354 0.152939
R11419 gnd.n6356 gnd.n6355 0.152939
R11420 gnd.n6356 gnd.n490 0.152939
R11421 gnd.n6364 gnd.n490 0.152939
R11422 gnd.n6365 gnd.n6364 0.152939
R11423 gnd.n6366 gnd.n6365 0.152939
R11424 gnd.n6366 gnd.n484 0.152939
R11425 gnd.n6374 gnd.n484 0.152939
R11426 gnd.n6375 gnd.n6374 0.152939
R11427 gnd.n6376 gnd.n6375 0.152939
R11428 gnd.n6376 gnd.n478 0.152939
R11429 gnd.n6384 gnd.n478 0.152939
R11430 gnd.n6385 gnd.n6384 0.152939
R11431 gnd.n6386 gnd.n6385 0.152939
R11432 gnd.n6386 gnd.n472 0.152939
R11433 gnd.n6394 gnd.n472 0.152939
R11434 gnd.n6395 gnd.n6394 0.152939
R11435 gnd.n6396 gnd.n6395 0.152939
R11436 gnd.n6396 gnd.n466 0.152939
R11437 gnd.n6404 gnd.n466 0.152939
R11438 gnd.n6405 gnd.n6404 0.152939
R11439 gnd.n6406 gnd.n6405 0.152939
R11440 gnd.n6406 gnd.n460 0.152939
R11441 gnd.n6414 gnd.n460 0.152939
R11442 gnd.n6415 gnd.n6414 0.152939
R11443 gnd.n6416 gnd.n6415 0.152939
R11444 gnd.n6416 gnd.n454 0.152939
R11445 gnd.n6424 gnd.n454 0.152939
R11446 gnd.n6425 gnd.n6424 0.152939
R11447 gnd.n6426 gnd.n6425 0.152939
R11448 gnd.n6426 gnd.n448 0.152939
R11449 gnd.n6434 gnd.n448 0.152939
R11450 gnd.n6435 gnd.n6434 0.152939
R11451 gnd.n6436 gnd.n6435 0.152939
R11452 gnd.n6436 gnd.n442 0.152939
R11453 gnd.n6444 gnd.n442 0.152939
R11454 gnd.n6445 gnd.n6444 0.152939
R11455 gnd.n6446 gnd.n6445 0.152939
R11456 gnd.n6446 gnd.n436 0.152939
R11457 gnd.n6454 gnd.n436 0.152939
R11458 gnd.n6455 gnd.n6454 0.152939
R11459 gnd.n6456 gnd.n6455 0.152939
R11460 gnd.n6456 gnd.n430 0.152939
R11461 gnd.n6464 gnd.n430 0.152939
R11462 gnd.n6465 gnd.n6464 0.152939
R11463 gnd.n6466 gnd.n6465 0.152939
R11464 gnd.n6466 gnd.n424 0.152939
R11465 gnd.n6474 gnd.n424 0.152939
R11466 gnd.n6475 gnd.n6474 0.152939
R11467 gnd.n6476 gnd.n6475 0.152939
R11468 gnd.n6476 gnd.n418 0.152939
R11469 gnd.n6484 gnd.n418 0.152939
R11470 gnd.n6485 gnd.n6484 0.152939
R11471 gnd.n6486 gnd.n6485 0.152939
R11472 gnd.n6486 gnd.n412 0.152939
R11473 gnd.n6494 gnd.n412 0.152939
R11474 gnd.n6495 gnd.n6494 0.152939
R11475 gnd.n6497 gnd.n6495 0.152939
R11476 gnd.n6497 gnd.n6496 0.152939
R11477 gnd.n6496 gnd.n406 0.152939
R11478 gnd.n6506 gnd.n406 0.152939
R11479 gnd.n6507 gnd.n401 0.152939
R11480 gnd.n6515 gnd.n401 0.152939
R11481 gnd.n6516 gnd.n6515 0.152939
R11482 gnd.n6517 gnd.n6516 0.152939
R11483 gnd.n6517 gnd.n395 0.152939
R11484 gnd.n6525 gnd.n395 0.152939
R11485 gnd.n6526 gnd.n6525 0.152939
R11486 gnd.n6527 gnd.n6526 0.152939
R11487 gnd.n6527 gnd.n389 0.152939
R11488 gnd.n6535 gnd.n389 0.152939
R11489 gnd.n6536 gnd.n6535 0.152939
R11490 gnd.n6537 gnd.n6536 0.152939
R11491 gnd.n6537 gnd.n383 0.152939
R11492 gnd.n6545 gnd.n383 0.152939
R11493 gnd.n6546 gnd.n6545 0.152939
R11494 gnd.n6547 gnd.n6546 0.152939
R11495 gnd.n6547 gnd.n377 0.152939
R11496 gnd.n6555 gnd.n377 0.152939
R11497 gnd.n6556 gnd.n6555 0.152939
R11498 gnd.n6557 gnd.n6556 0.152939
R11499 gnd.n6557 gnd.n371 0.152939
R11500 gnd.n6565 gnd.n371 0.152939
R11501 gnd.n6566 gnd.n6565 0.152939
R11502 gnd.n6567 gnd.n6566 0.152939
R11503 gnd.n6567 gnd.n365 0.152939
R11504 gnd.n6575 gnd.n365 0.152939
R11505 gnd.n6576 gnd.n6575 0.152939
R11506 gnd.n6577 gnd.n6576 0.152939
R11507 gnd.n6577 gnd.n359 0.152939
R11508 gnd.n6585 gnd.n359 0.152939
R11509 gnd.n6586 gnd.n6585 0.152939
R11510 gnd.n6587 gnd.n6586 0.152939
R11511 gnd.n6587 gnd.n353 0.152939
R11512 gnd.n6595 gnd.n353 0.152939
R11513 gnd.n6596 gnd.n6595 0.152939
R11514 gnd.n6597 gnd.n6596 0.152939
R11515 gnd.n6597 gnd.n347 0.152939
R11516 gnd.n6605 gnd.n347 0.152939
R11517 gnd.n6606 gnd.n6605 0.152939
R11518 gnd.n6607 gnd.n6606 0.152939
R11519 gnd.n6607 gnd.n341 0.152939
R11520 gnd.n6615 gnd.n341 0.152939
R11521 gnd.n6616 gnd.n6615 0.152939
R11522 gnd.n6617 gnd.n6616 0.152939
R11523 gnd.n6617 gnd.n335 0.152939
R11524 gnd.n6625 gnd.n335 0.152939
R11525 gnd.n6626 gnd.n6625 0.152939
R11526 gnd.n6627 gnd.n6626 0.152939
R11527 gnd.n6627 gnd.n329 0.152939
R11528 gnd.n6635 gnd.n329 0.152939
R11529 gnd.n6636 gnd.n6635 0.152939
R11530 gnd.n6637 gnd.n6636 0.152939
R11531 gnd.n6637 gnd.n323 0.152939
R11532 gnd.n6645 gnd.n323 0.152939
R11533 gnd.n6646 gnd.n6645 0.152939
R11534 gnd.n6647 gnd.n6646 0.152939
R11535 gnd.n6647 gnd.n317 0.152939
R11536 gnd.n6655 gnd.n317 0.152939
R11537 gnd.n6656 gnd.n6655 0.152939
R11538 gnd.n6657 gnd.n6656 0.152939
R11539 gnd.n6657 gnd.n311 0.152939
R11540 gnd.n6665 gnd.n311 0.152939
R11541 gnd.n6666 gnd.n6665 0.152939
R11542 gnd.n6667 gnd.n6666 0.152939
R11543 gnd.n6667 gnd.n305 0.152939
R11544 gnd.n6675 gnd.n305 0.152939
R11545 gnd.n6676 gnd.n6675 0.152939
R11546 gnd.n6677 gnd.n6676 0.152939
R11547 gnd.n6677 gnd.n299 0.152939
R11548 gnd.n6685 gnd.n299 0.152939
R11549 gnd.n6686 gnd.n6685 0.152939
R11550 gnd.n6687 gnd.n6686 0.152939
R11551 gnd.n6687 gnd.n293 0.152939
R11552 gnd.n6695 gnd.n293 0.152939
R11553 gnd.n6696 gnd.n6695 0.152939
R11554 gnd.n6697 gnd.n6696 0.152939
R11555 gnd.n6697 gnd.n287 0.152939
R11556 gnd.n6705 gnd.n287 0.152939
R11557 gnd.n6706 gnd.n6705 0.152939
R11558 gnd.n6707 gnd.n6706 0.152939
R11559 gnd.n6707 gnd.n281 0.152939
R11560 gnd.n6716 gnd.n281 0.152939
R11561 gnd.n6717 gnd.n6716 0.152939
R11562 gnd.n6718 gnd.n6717 0.152939
R11563 gnd.n276 gnd.n275 0.152939
R11564 gnd.n277 gnd.n276 0.152939
R11565 gnd.n278 gnd.n277 0.152939
R11566 gnd.n6756 gnd.n6755 0.152939
R11567 gnd.n6757 gnd.n6756 0.152939
R11568 gnd.n6757 gnd.n198 0.152939
R11569 gnd.n6771 gnd.n198 0.152939
R11570 gnd.n6772 gnd.n6771 0.152939
R11571 gnd.n6773 gnd.n6772 0.152939
R11572 gnd.n6773 gnd.n182 0.152939
R11573 gnd.n6787 gnd.n182 0.152939
R11574 gnd.n6788 gnd.n6787 0.152939
R11575 gnd.n6789 gnd.n6788 0.152939
R11576 gnd.n6789 gnd.n166 0.152939
R11577 gnd.n6877 gnd.n166 0.152939
R11578 gnd.n6878 gnd.n6877 0.152939
R11579 gnd.n6879 gnd.n6878 0.152939
R11580 gnd.n6879 gnd.n88 0.152939
R11581 gnd.n6959 gnd.n88 0.152939
R11582 gnd.n6958 gnd.n89 0.152939
R11583 gnd.n91 gnd.n89 0.152939
R11584 gnd.n96 gnd.n91 0.152939
R11585 gnd.n97 gnd.n96 0.152939
R11586 gnd.n98 gnd.n97 0.152939
R11587 gnd.n99 gnd.n98 0.152939
R11588 gnd.n103 gnd.n99 0.152939
R11589 gnd.n104 gnd.n103 0.152939
R11590 gnd.n105 gnd.n104 0.152939
R11591 gnd.n106 gnd.n105 0.152939
R11592 gnd.n110 gnd.n106 0.152939
R11593 gnd.n111 gnd.n110 0.152939
R11594 gnd.n112 gnd.n111 0.152939
R11595 gnd.n113 gnd.n112 0.152939
R11596 gnd.n117 gnd.n113 0.152939
R11597 gnd.n118 gnd.n117 0.152939
R11598 gnd.n119 gnd.n118 0.152939
R11599 gnd.n120 gnd.n119 0.152939
R11600 gnd.n124 gnd.n120 0.152939
R11601 gnd.n125 gnd.n124 0.152939
R11602 gnd.n126 gnd.n125 0.152939
R11603 gnd.n127 gnd.n126 0.152939
R11604 gnd.n131 gnd.n127 0.152939
R11605 gnd.n132 gnd.n131 0.152939
R11606 gnd.n133 gnd.n132 0.152939
R11607 gnd.n134 gnd.n133 0.152939
R11608 gnd.n138 gnd.n134 0.152939
R11609 gnd.n139 gnd.n138 0.152939
R11610 gnd.n140 gnd.n139 0.152939
R11611 gnd.n141 gnd.n140 0.152939
R11612 gnd.n145 gnd.n141 0.152939
R11613 gnd.n146 gnd.n145 0.152939
R11614 gnd.n147 gnd.n146 0.152939
R11615 gnd.n148 gnd.n147 0.152939
R11616 gnd.n152 gnd.n148 0.152939
R11617 gnd.n153 gnd.n152 0.152939
R11618 gnd.n6889 gnd.n153 0.152939
R11619 gnd.n6889 gnd.n6888 0.152939
R11620 gnd.n3918 gnd.n1359 0.152939
R11621 gnd.n3919 gnd.n3918 0.152939
R11622 gnd.n3920 gnd.n3919 0.152939
R11623 gnd.n3921 gnd.n3920 0.152939
R11624 gnd.n3922 gnd.n3921 0.152939
R11625 gnd.n3923 gnd.n3922 0.152939
R11626 gnd.n3924 gnd.n3923 0.152939
R11627 gnd.n3925 gnd.n3924 0.152939
R11628 gnd.n3926 gnd.n3925 0.152939
R11629 gnd.n3927 gnd.n3926 0.152939
R11630 gnd.n3928 gnd.n3927 0.152939
R11631 gnd.n3929 gnd.n3928 0.152939
R11632 gnd.n3930 gnd.n3929 0.152939
R11633 gnd.n3932 gnd.n3930 0.152939
R11634 gnd.n3932 gnd.n3931 0.152939
R11635 gnd.n3931 gnd.n1423 0.152939
R11636 gnd.n1424 gnd.n1423 0.152939
R11637 gnd.n1425 gnd.n1424 0.152939
R11638 gnd.n1426 gnd.n1425 0.152939
R11639 gnd.n1427 gnd.n1426 0.152939
R11640 gnd.n1427 gnd.n1395 0.152939
R11641 gnd.n1395 gnd.n1394 0.152939
R11642 gnd.n1394 gnd.n235 0.152939
R11643 gnd.n236 gnd.n235 0.152939
R11644 gnd.n237 gnd.n236 0.152939
R11645 gnd.n238 gnd.n237 0.152939
R11646 gnd.n239 gnd.n238 0.152939
R11647 gnd.n240 gnd.n239 0.152939
R11648 gnd.n241 gnd.n240 0.152939
R11649 gnd.n242 gnd.n241 0.152939
R11650 gnd.n243 gnd.n242 0.152939
R11651 gnd.n244 gnd.n243 0.152939
R11652 gnd.n245 gnd.n244 0.152939
R11653 gnd.n246 gnd.n245 0.152939
R11654 gnd.n247 gnd.n246 0.152939
R11655 gnd.n248 gnd.n247 0.152939
R11656 gnd.n249 gnd.n248 0.152939
R11657 gnd.n250 gnd.n249 0.152939
R11658 gnd.n252 gnd.n250 0.152939
R11659 gnd.n252 gnd.n251 0.152939
R11660 gnd.n251 gnd.n159 0.152939
R11661 gnd.n6887 gnd.n159 0.152939
R11662 gnd.n1316 gnd.n1315 0.152939
R11663 gnd.n1317 gnd.n1316 0.152939
R11664 gnd.n1318 gnd.n1317 0.152939
R11665 gnd.n1319 gnd.n1318 0.152939
R11666 gnd.n1320 gnd.n1319 0.152939
R11667 gnd.n1321 gnd.n1320 0.152939
R11668 gnd.n1322 gnd.n1321 0.152939
R11669 gnd.n1323 gnd.n1322 0.152939
R11670 gnd.n1324 gnd.n1323 0.152939
R11671 gnd.n1325 gnd.n1324 0.152939
R11672 gnd.n1326 gnd.n1325 0.152939
R11673 gnd.n1327 gnd.n1326 0.152939
R11674 gnd.n1328 gnd.n1327 0.152939
R11675 gnd.n1329 gnd.n1328 0.152939
R11676 gnd.n1330 gnd.n1329 0.152939
R11677 gnd.n1337 gnd.n1336 0.152939
R11678 gnd.n1338 gnd.n1337 0.152939
R11679 gnd.n1339 gnd.n1338 0.152939
R11680 gnd.n1340 gnd.n1339 0.152939
R11681 gnd.n1341 gnd.n1340 0.152939
R11682 gnd.n1342 gnd.n1341 0.152939
R11683 gnd.n1343 gnd.n1342 0.152939
R11684 gnd.n1344 gnd.n1343 0.152939
R11685 gnd.n1345 gnd.n1344 0.152939
R11686 gnd.n1346 gnd.n1345 0.152939
R11687 gnd.n1347 gnd.n1346 0.152939
R11688 gnd.n1348 gnd.n1347 0.152939
R11689 gnd.n1349 gnd.n1348 0.152939
R11690 gnd.n1350 gnd.n1349 0.152939
R11691 gnd.n1351 gnd.n1350 0.152939
R11692 gnd.n1352 gnd.n1351 0.152939
R11693 gnd.n1353 gnd.n1352 0.152939
R11694 gnd.n4159 gnd.n1353 0.152939
R11695 gnd.n4159 gnd.n4158 0.152939
R11696 gnd.n4158 gnd.n4157 0.152939
R11697 gnd.n3977 gnd.n1501 0.152939
R11698 gnd.n3978 gnd.n3977 0.152939
R11699 gnd.n3979 gnd.n3978 0.152939
R11700 gnd.n3980 gnd.n3979 0.152939
R11701 gnd.n3980 gnd.n1475 0.152939
R11702 gnd.n4009 gnd.n1475 0.152939
R11703 gnd.n4010 gnd.n4009 0.152939
R11704 gnd.n4011 gnd.n4010 0.152939
R11705 gnd.n4012 gnd.n4011 0.152939
R11706 gnd.n4012 gnd.n1450 0.152939
R11707 gnd.n4043 gnd.n1450 0.152939
R11708 gnd.n4044 gnd.n4043 0.152939
R11709 gnd.n4045 gnd.n4044 0.152939
R11710 gnd.n4046 gnd.n4045 0.152939
R11711 gnd.n4046 gnd.n212 0.152939
R11712 gnd.n6755 gnd.n212 0.152939
R11713 gnd.n2236 gnd.n2230 0.152939
R11714 gnd.n2239 gnd.n2236 0.152939
R11715 gnd.n2240 gnd.n2239 0.152939
R11716 gnd.n2241 gnd.n2240 0.152939
R11717 gnd.n2242 gnd.n2241 0.152939
R11718 gnd.n2245 gnd.n2242 0.152939
R11719 gnd.n2246 gnd.n2245 0.152939
R11720 gnd.n2247 gnd.n2246 0.152939
R11721 gnd.n2248 gnd.n2247 0.152939
R11722 gnd.n2251 gnd.n2248 0.152939
R11723 gnd.n2252 gnd.n2251 0.152939
R11724 gnd.n2253 gnd.n2252 0.152939
R11725 gnd.n2254 gnd.n2253 0.152939
R11726 gnd.n2257 gnd.n2254 0.152939
R11727 gnd.n2258 gnd.n2257 0.152939
R11728 gnd.n2259 gnd.n2258 0.152939
R11729 gnd.n2260 gnd.n2259 0.152939
R11730 gnd.n2261 gnd.n2260 0.152939
R11731 gnd.n2261 gnd.n1982 0.152939
R11732 gnd.n2903 gnd.n1982 0.152939
R11733 gnd.n2904 gnd.n2903 0.152939
R11734 gnd.n2905 gnd.n2904 0.152939
R11735 gnd.n2905 gnd.n1968 0.152939
R11736 gnd.n2919 gnd.n1968 0.152939
R11737 gnd.n2920 gnd.n2919 0.152939
R11738 gnd.n2921 gnd.n2920 0.152939
R11739 gnd.n2922 gnd.n2921 0.152939
R11740 gnd.n2922 gnd.n1936 0.152939
R11741 gnd.n3043 gnd.n1936 0.152939
R11742 gnd.n3044 gnd.n3043 0.152939
R11743 gnd.n3045 gnd.n3044 0.152939
R11744 gnd.n3045 gnd.n1922 0.152939
R11745 gnd.n3059 gnd.n1922 0.152939
R11746 gnd.n3060 gnd.n3059 0.152939
R11747 gnd.n3061 gnd.n3060 0.152939
R11748 gnd.n3061 gnd.n1907 0.152939
R11749 gnd.n3075 gnd.n1907 0.152939
R11750 gnd.n3076 gnd.n3075 0.152939
R11751 gnd.n3077 gnd.n3076 0.152939
R11752 gnd.n3077 gnd.n1893 0.152939
R11753 gnd.n3090 gnd.n1893 0.152939
R11754 gnd.n3091 gnd.n3090 0.152939
R11755 gnd.n3092 gnd.n3091 0.152939
R11756 gnd.n3093 gnd.n3092 0.152939
R11757 gnd.n3093 gnd.n1861 0.152939
R11758 gnd.n3216 gnd.n1861 0.152939
R11759 gnd.n3217 gnd.n3216 0.152939
R11760 gnd.n3218 gnd.n3217 0.152939
R11761 gnd.n3218 gnd.n1847 0.152939
R11762 gnd.n3232 gnd.n1847 0.152939
R11763 gnd.n3233 gnd.n3232 0.152939
R11764 gnd.n3234 gnd.n3233 0.152939
R11765 gnd.n3234 gnd.n1834 0.152939
R11766 gnd.n3248 gnd.n1834 0.152939
R11767 gnd.n3249 gnd.n3248 0.152939
R11768 gnd.n3250 gnd.n3249 0.152939
R11769 gnd.n3250 gnd.n1823 0.152939
R11770 gnd.n3264 gnd.n1823 0.152939
R11771 gnd.n3265 gnd.n3264 0.152939
R11772 gnd.n3266 gnd.n3265 0.152939
R11773 gnd.n3267 gnd.n3266 0.152939
R11774 gnd.n3267 gnd.n1790 0.152939
R11775 gnd.n3387 gnd.n1790 0.152939
R11776 gnd.n3388 gnd.n3387 0.152939
R11777 gnd.n3389 gnd.n3388 0.152939
R11778 gnd.n3389 gnd.n1775 0.152939
R11779 gnd.n3403 gnd.n1775 0.152939
R11780 gnd.n3404 gnd.n3403 0.152939
R11781 gnd.n3405 gnd.n3404 0.152939
R11782 gnd.n3405 gnd.n1760 0.152939
R11783 gnd.n3419 gnd.n1760 0.152939
R11784 gnd.n3420 gnd.n3419 0.152939
R11785 gnd.n3421 gnd.n3420 0.152939
R11786 gnd.n3421 gnd.n1747 0.152939
R11787 gnd.n3435 gnd.n1747 0.152939
R11788 gnd.n3436 gnd.n3435 0.152939
R11789 gnd.n3437 gnd.n3436 0.152939
R11790 gnd.n3438 gnd.n3437 0.152939
R11791 gnd.n3438 gnd.n1715 0.152939
R11792 gnd.n3793 gnd.n1715 0.152939
R11793 gnd.n3794 gnd.n3793 0.152939
R11794 gnd.n3795 gnd.n3794 0.152939
R11795 gnd.n3795 gnd.n1702 0.152939
R11796 gnd.n3809 gnd.n1702 0.152939
R11797 gnd.n3810 gnd.n3809 0.152939
R11798 gnd.n3811 gnd.n3810 0.152939
R11799 gnd.n3811 gnd.n1688 0.152939
R11800 gnd.n3825 gnd.n1688 0.152939
R11801 gnd.n3826 gnd.n3825 0.152939
R11802 gnd.n3827 gnd.n3826 0.152939
R11803 gnd.n3827 gnd.n1675 0.152939
R11804 gnd.n3841 gnd.n1675 0.152939
R11805 gnd.n3842 gnd.n3841 0.152939
R11806 gnd.n3843 gnd.n3842 0.152939
R11807 gnd.n3843 gnd.n1661 0.152939
R11808 gnd.n3857 gnd.n1661 0.152939
R11809 gnd.n3858 gnd.n3857 0.152939
R11810 gnd.n3859 gnd.n3858 0.152939
R11811 gnd.n3859 gnd.n1647 0.152939
R11812 gnd.n3875 gnd.n1647 0.152939
R11813 gnd.n3876 gnd.n3875 0.152939
R11814 gnd.n3877 gnd.n3876 0.152939
R11815 gnd.n3879 gnd.n3877 0.152939
R11816 gnd.n3879 gnd.n3878 0.152939
R11817 gnd.n3878 gnd.n1278 0.152939
R11818 gnd.n1279 gnd.n1278 0.152939
R11819 gnd.n1280 gnd.n1279 0.152939
R11820 gnd.n3960 gnd.n1280 0.152939
R11821 gnd.n3961 gnd.n3960 0.152939
R11822 gnd.n3966 gnd.n3961 0.152939
R11823 gnd.n3967 gnd.n3966 0.152939
R11824 gnd.n3968 gnd.n3967 0.152939
R11825 gnd.n3969 gnd.n3968 0.152939
R11826 gnd.n3969 gnd.n1484 0.152939
R11827 gnd.n3998 gnd.n1484 0.152939
R11828 gnd.n3999 gnd.n3998 0.152939
R11829 gnd.n4000 gnd.n3999 0.152939
R11830 gnd.n4001 gnd.n4000 0.152939
R11831 gnd.n4001 gnd.n1459 0.152939
R11832 gnd.n4029 gnd.n1459 0.152939
R11833 gnd.n4030 gnd.n4029 0.152939
R11834 gnd.n4031 gnd.n4030 0.152939
R11835 gnd.n4032 gnd.n4031 0.152939
R11836 gnd.n4034 gnd.n4032 0.152939
R11837 gnd.n4034 gnd.n4033 0.152939
R11838 gnd.n4033 gnd.n1435 0.152939
R11839 gnd.n2381 gnd.n2354 0.152939
R11840 gnd.n2439 gnd.n2354 0.152939
R11841 gnd.n2440 gnd.n2439 0.152939
R11842 gnd.n2441 gnd.n2440 0.152939
R11843 gnd.n2441 gnd.n2352 0.152939
R11844 gnd.n2447 gnd.n2352 0.152939
R11845 gnd.n2448 gnd.n2447 0.152939
R11846 gnd.n2449 gnd.n2448 0.152939
R11847 gnd.n2449 gnd.n2350 0.152939
R11848 gnd.n2455 gnd.n2350 0.152939
R11849 gnd.n2456 gnd.n2455 0.152939
R11850 gnd.n2458 gnd.n2456 0.152939
R11851 gnd.n2458 gnd.n2457 0.152939
R11852 gnd.n2457 gnd.n2329 0.152939
R11853 gnd.n2475 gnd.n2329 0.152939
R11854 gnd.n2476 gnd.n2475 0.152939
R11855 gnd.n2477 gnd.n2476 0.152939
R11856 gnd.n2477 gnd.n2220 0.152939
R11857 gnd.n2491 gnd.n2220 0.152939
R11858 gnd.n2492 gnd.n2491 0.152939
R11859 gnd.n2420 gnd.n2361 0.152939
R11860 gnd.n2362 gnd.n2361 0.152939
R11861 gnd.n2363 gnd.n2362 0.152939
R11862 gnd.n2364 gnd.n2363 0.152939
R11863 gnd.n2365 gnd.n2364 0.152939
R11864 gnd.n2366 gnd.n2365 0.152939
R11865 gnd.n2367 gnd.n2366 0.152939
R11866 gnd.n2368 gnd.n2367 0.152939
R11867 gnd.n2369 gnd.n2368 0.152939
R11868 gnd.n2370 gnd.n2369 0.152939
R11869 gnd.n2371 gnd.n2370 0.152939
R11870 gnd.n2372 gnd.n2371 0.152939
R11871 gnd.n2373 gnd.n2372 0.152939
R11872 gnd.n2374 gnd.n2373 0.152939
R11873 gnd.n2375 gnd.n2374 0.152939
R11874 gnd.n2385 gnd.n2375 0.152939
R11875 gnd.n2385 gnd.n2384 0.152939
R11876 gnd.n2384 gnd.n2383 0.152939
R11877 gnd.n2426 gnd.n2421 0.152939
R11878 gnd.n2426 gnd.n2425 0.152939
R11879 gnd.n2425 gnd.n2424 0.152939
R11880 gnd.n2424 gnd.n2422 0.152939
R11881 gnd.n2422 gnd.n978 0.152939
R11882 gnd.n979 gnd.n978 0.152939
R11883 gnd.n980 gnd.n979 0.152939
R11884 gnd.n996 gnd.n980 0.152939
R11885 gnd.n997 gnd.n996 0.152939
R11886 gnd.n998 gnd.n997 0.152939
R11887 gnd.n999 gnd.n998 0.152939
R11888 gnd.n1018 gnd.n999 0.152939
R11889 gnd.n1019 gnd.n1018 0.152939
R11890 gnd.n1020 gnd.n1019 0.152939
R11891 gnd.n1021 gnd.n1020 0.152939
R11892 gnd.n1042 gnd.n1021 0.152939
R11893 gnd.n1043 gnd.n1042 0.152939
R11894 gnd.n1044 gnd.n1043 0.152939
R11895 gnd.n1045 gnd.n1044 0.152939
R11896 gnd.n1046 gnd.n1045 0.152939
R11897 gnd.n2216 gnd.n1046 0.152939
R11898 gnd.n2216 gnd.n1061 0.152939
R11899 gnd.n1062 gnd.n1061 0.152939
R11900 gnd.n1063 gnd.n1062 0.152939
R11901 gnd.n1079 gnd.n1063 0.152939
R11902 gnd.n1080 gnd.n1079 0.152939
R11903 gnd.n1081 gnd.n1080 0.152939
R11904 gnd.n1082 gnd.n1081 0.152939
R11905 gnd.n1100 gnd.n1082 0.152939
R11906 gnd.n1101 gnd.n1100 0.152939
R11907 gnd.n1102 gnd.n1101 0.152939
R11908 gnd.n1103 gnd.n1102 0.152939
R11909 gnd.n1122 gnd.n1103 0.152939
R11910 gnd.n1123 gnd.n1122 0.152939
R11911 gnd.n1124 gnd.n1123 0.152939
R11912 gnd.n1125 gnd.n1124 0.152939
R11913 gnd.n1144 gnd.n1125 0.152939
R11914 gnd.n1145 gnd.n1144 0.152939
R11915 gnd.n1146 gnd.n1145 0.152939
R11916 gnd.n1147 gnd.n1146 0.152939
R11917 gnd.n1164 gnd.n1147 0.152939
R11918 gnd.n4366 gnd.n1164 0.152939
R11919 gnd.n1090 gnd.n1031 0.152939
R11920 gnd.n1091 gnd.n1090 0.152939
R11921 gnd.n1092 gnd.n1091 0.152939
R11922 gnd.n1093 gnd.n1092 0.152939
R11923 gnd.n1111 gnd.n1093 0.152939
R11924 gnd.n1112 gnd.n1111 0.152939
R11925 gnd.n1113 gnd.n1112 0.152939
R11926 gnd.n1114 gnd.n1113 0.152939
R11927 gnd.n1133 gnd.n1114 0.152939
R11928 gnd.n1134 gnd.n1133 0.152939
R11929 gnd.n1135 gnd.n1134 0.152939
R11930 gnd.n1136 gnd.n1135 0.152939
R11931 gnd.n1154 gnd.n1136 0.152939
R11932 gnd.n1155 gnd.n1154 0.152939
R11933 gnd.n1156 gnd.n1155 0.152939
R11934 gnd.n1157 gnd.n1156 0.152939
R11935 gnd.n2142 gnd.n2141 0.152939
R11936 gnd.n2143 gnd.n2142 0.152939
R11937 gnd.n2144 gnd.n2143 0.152939
R11938 gnd.n2145 gnd.n2144 0.152939
R11939 gnd.n2146 gnd.n2145 0.152939
R11940 gnd.n2147 gnd.n2146 0.152939
R11941 gnd.n2148 gnd.n2147 0.152939
R11942 gnd.n2149 gnd.n2148 0.152939
R11943 gnd.n2150 gnd.n2149 0.152939
R11944 gnd.n2151 gnd.n2150 0.152939
R11945 gnd.n2152 gnd.n2151 0.152939
R11946 gnd.n2153 gnd.n2152 0.152939
R11947 gnd.n2154 gnd.n2153 0.152939
R11948 gnd.n2155 gnd.n2154 0.152939
R11949 gnd.n2156 gnd.n2155 0.152939
R11950 gnd.n2624 gnd.n2623 0.152939
R11951 gnd.n2623 gnd.n2161 0.152939
R11952 gnd.n2162 gnd.n2161 0.152939
R11953 gnd.n2163 gnd.n2162 0.152939
R11954 gnd.n2164 gnd.n2163 0.152939
R11955 gnd.n2165 gnd.n2164 0.152939
R11956 gnd.n2166 gnd.n2165 0.152939
R11957 gnd.n2167 gnd.n2166 0.152939
R11958 gnd.n2168 gnd.n2167 0.152939
R11959 gnd.n2169 gnd.n2168 0.152939
R11960 gnd.n2170 gnd.n2169 0.152939
R11961 gnd.n2171 gnd.n2170 0.152939
R11962 gnd.n2172 gnd.n2171 0.152939
R11963 gnd.n2173 gnd.n2172 0.152939
R11964 gnd.n2174 gnd.n2173 0.152939
R11965 gnd.n2175 gnd.n2174 0.152939
R11966 gnd.n2176 gnd.n2175 0.152939
R11967 gnd.n2177 gnd.n2176 0.152939
R11968 gnd.n2583 gnd.n2177 0.152939
R11969 gnd.n2583 gnd.n2582 0.152939
R11970 gnd.n4492 gnd.n953 0.152939
R11971 gnd.n4492 gnd.n4491 0.152939
R11972 gnd.n4491 gnd.n4490 0.152939
R11973 gnd.n4490 gnd.n956 0.152939
R11974 gnd.n2336 gnd.n956 0.152939
R11975 gnd.n2337 gnd.n2336 0.152939
R11976 gnd.n2337 gnd.n2334 0.152939
R11977 gnd.n2343 gnd.n2334 0.152939
R11978 gnd.n2344 gnd.n2343 0.152939
R11979 gnd.n2345 gnd.n2344 0.152939
R11980 gnd.n2345 gnd.n2332 0.152939
R11981 gnd.n2464 gnd.n2332 0.152939
R11982 gnd.n2465 gnd.n2464 0.152939
R11983 gnd.n2466 gnd.n2465 0.152939
R11984 gnd.n2467 gnd.n2466 0.152939
R11985 gnd.n2467 gnd.n2223 0.152939
R11986 gnd.n2483 gnd.n2223 0.152939
R11987 gnd.n2484 gnd.n2483 0.152939
R11988 gnd.n2485 gnd.n2484 0.152939
R11989 gnd.n2485 gnd.n2217 0.152939
R11990 gnd.n2499 gnd.n2217 0.152939
R11991 gnd.n2500 gnd.n2499 0.152939
R11992 gnd.n2501 gnd.n2500 0.152939
R11993 gnd.n2501 gnd.n2209 0.152939
R11994 gnd.n2515 gnd.n2209 0.152939
R11995 gnd.n2516 gnd.n2515 0.152939
R11996 gnd.n2517 gnd.n2516 0.152939
R11997 gnd.n2517 gnd.n2203 0.152939
R11998 gnd.n2531 gnd.n2203 0.152939
R11999 gnd.n2532 gnd.n2531 0.152939
R12000 gnd.n2533 gnd.n2532 0.152939
R12001 gnd.n2533 gnd.n2196 0.152939
R12002 gnd.n2547 gnd.n2196 0.152939
R12003 gnd.n2548 gnd.n2547 0.152939
R12004 gnd.n2549 gnd.n2548 0.152939
R12005 gnd.n2549 gnd.n2190 0.152939
R12006 gnd.n2563 gnd.n2190 0.152939
R12007 gnd.n2564 gnd.n2563 0.152939
R12008 gnd.n2566 gnd.n2564 0.152939
R12009 gnd.n2566 gnd.n2565 0.152939
R12010 gnd.n2565 gnd.n2182 0.152939
R12011 gnd.n2581 gnd.n2182 0.152939
R12012 gnd.n911 gnd.n910 0.152939
R12013 gnd.n912 gnd.n911 0.152939
R12014 gnd.n913 gnd.n912 0.152939
R12015 gnd.n914 gnd.n913 0.152939
R12016 gnd.n915 gnd.n914 0.152939
R12017 gnd.n916 gnd.n915 0.152939
R12018 gnd.n917 gnd.n916 0.152939
R12019 gnd.n918 gnd.n917 0.152939
R12020 gnd.n919 gnd.n918 0.152939
R12021 gnd.n920 gnd.n919 0.152939
R12022 gnd.n921 gnd.n920 0.152939
R12023 gnd.n922 gnd.n921 0.152939
R12024 gnd.n923 gnd.n922 0.152939
R12025 gnd.n924 gnd.n923 0.152939
R12026 gnd.n925 gnd.n924 0.152939
R12027 gnd.n926 gnd.n925 0.152939
R12028 gnd.n927 gnd.n926 0.152939
R12029 gnd.n930 gnd.n927 0.152939
R12030 gnd.n931 gnd.n930 0.152939
R12031 gnd.n932 gnd.n931 0.152939
R12032 gnd.n933 gnd.n932 0.152939
R12033 gnd.n934 gnd.n933 0.152939
R12034 gnd.n935 gnd.n934 0.152939
R12035 gnd.n936 gnd.n935 0.152939
R12036 gnd.n937 gnd.n936 0.152939
R12037 gnd.n938 gnd.n937 0.152939
R12038 gnd.n939 gnd.n938 0.152939
R12039 gnd.n940 gnd.n939 0.152939
R12040 gnd.n941 gnd.n940 0.152939
R12041 gnd.n942 gnd.n941 0.152939
R12042 gnd.n943 gnd.n942 0.152939
R12043 gnd.n944 gnd.n943 0.152939
R12044 gnd.n945 gnd.n944 0.152939
R12045 gnd.n946 gnd.n945 0.152939
R12046 gnd.n947 gnd.n946 0.152939
R12047 gnd.n4500 gnd.n947 0.152939
R12048 gnd.n4500 gnd.n4499 0.152939
R12049 gnd.n4499 gnd.n4498 0.152939
R12050 gnd.n2432 gnd.n2430 0.152939
R12051 gnd.n2432 gnd.n2431 0.152939
R12052 gnd.n2431 gnd.n967 0.152939
R12053 gnd.n968 gnd.n967 0.152939
R12054 gnd.n969 gnd.n968 0.152939
R12055 gnd.n987 gnd.n969 0.152939
R12056 gnd.n988 gnd.n987 0.152939
R12057 gnd.n989 gnd.n988 0.152939
R12058 gnd.n990 gnd.n989 0.152939
R12059 gnd.n1007 gnd.n990 0.152939
R12060 gnd.n1008 gnd.n1007 0.152939
R12061 gnd.n1009 gnd.n1008 0.152939
R12062 gnd.n1010 gnd.n1009 0.152939
R12063 gnd.n1029 gnd.n1010 0.152939
R12064 gnd.n1030 gnd.n1029 0.152939
R12065 gnd.n1031 gnd.n1030 0.152939
R12066 gnd.n2313 gnd.n2307 0.152939
R12067 gnd.n2319 gnd.n2307 0.152939
R12068 gnd.n2320 gnd.n2319 0.152939
R12069 gnd.n640 gnd.n639 0.152939
R12070 gnd.n641 gnd.n640 0.152939
R12071 gnd.n646 gnd.n641 0.152939
R12072 gnd.n647 gnd.n646 0.152939
R12073 gnd.n648 gnd.n647 0.152939
R12074 gnd.n649 gnd.n648 0.152939
R12075 gnd.n654 gnd.n649 0.152939
R12076 gnd.n655 gnd.n654 0.152939
R12077 gnd.n656 gnd.n655 0.152939
R12078 gnd.n657 gnd.n656 0.152939
R12079 gnd.n662 gnd.n657 0.152939
R12080 gnd.n663 gnd.n662 0.152939
R12081 gnd.n664 gnd.n663 0.152939
R12082 gnd.n665 gnd.n664 0.152939
R12083 gnd.n670 gnd.n665 0.152939
R12084 gnd.n671 gnd.n670 0.152939
R12085 gnd.n672 gnd.n671 0.152939
R12086 gnd.n673 gnd.n672 0.152939
R12087 gnd.n678 gnd.n673 0.152939
R12088 gnd.n679 gnd.n678 0.152939
R12089 gnd.n680 gnd.n679 0.152939
R12090 gnd.n681 gnd.n680 0.152939
R12091 gnd.n686 gnd.n681 0.152939
R12092 gnd.n687 gnd.n686 0.152939
R12093 gnd.n688 gnd.n687 0.152939
R12094 gnd.n689 gnd.n688 0.152939
R12095 gnd.n694 gnd.n689 0.152939
R12096 gnd.n695 gnd.n694 0.152939
R12097 gnd.n696 gnd.n695 0.152939
R12098 gnd.n697 gnd.n696 0.152939
R12099 gnd.n702 gnd.n697 0.152939
R12100 gnd.n703 gnd.n702 0.152939
R12101 gnd.n704 gnd.n703 0.152939
R12102 gnd.n705 gnd.n704 0.152939
R12103 gnd.n710 gnd.n705 0.152939
R12104 gnd.n711 gnd.n710 0.152939
R12105 gnd.n712 gnd.n711 0.152939
R12106 gnd.n713 gnd.n712 0.152939
R12107 gnd.n718 gnd.n713 0.152939
R12108 gnd.n719 gnd.n718 0.152939
R12109 gnd.n720 gnd.n719 0.152939
R12110 gnd.n721 gnd.n720 0.152939
R12111 gnd.n726 gnd.n721 0.152939
R12112 gnd.n727 gnd.n726 0.152939
R12113 gnd.n728 gnd.n727 0.152939
R12114 gnd.n729 gnd.n728 0.152939
R12115 gnd.n734 gnd.n729 0.152939
R12116 gnd.n735 gnd.n734 0.152939
R12117 gnd.n736 gnd.n735 0.152939
R12118 gnd.n737 gnd.n736 0.152939
R12119 gnd.n742 gnd.n737 0.152939
R12120 gnd.n743 gnd.n742 0.152939
R12121 gnd.n744 gnd.n743 0.152939
R12122 gnd.n745 gnd.n744 0.152939
R12123 gnd.n750 gnd.n745 0.152939
R12124 gnd.n751 gnd.n750 0.152939
R12125 gnd.n752 gnd.n751 0.152939
R12126 gnd.n753 gnd.n752 0.152939
R12127 gnd.n758 gnd.n753 0.152939
R12128 gnd.n759 gnd.n758 0.152939
R12129 gnd.n760 gnd.n759 0.152939
R12130 gnd.n761 gnd.n760 0.152939
R12131 gnd.n766 gnd.n761 0.152939
R12132 gnd.n767 gnd.n766 0.152939
R12133 gnd.n768 gnd.n767 0.152939
R12134 gnd.n769 gnd.n768 0.152939
R12135 gnd.n774 gnd.n769 0.152939
R12136 gnd.n775 gnd.n774 0.152939
R12137 gnd.n776 gnd.n775 0.152939
R12138 gnd.n777 gnd.n776 0.152939
R12139 gnd.n782 gnd.n777 0.152939
R12140 gnd.n783 gnd.n782 0.152939
R12141 gnd.n784 gnd.n783 0.152939
R12142 gnd.n785 gnd.n784 0.152939
R12143 gnd.n790 gnd.n785 0.152939
R12144 gnd.n791 gnd.n790 0.152939
R12145 gnd.n792 gnd.n791 0.152939
R12146 gnd.n793 gnd.n792 0.152939
R12147 gnd.n798 gnd.n793 0.152939
R12148 gnd.n799 gnd.n798 0.152939
R12149 gnd.n800 gnd.n799 0.152939
R12150 gnd.n801 gnd.n800 0.152939
R12151 gnd.n2310 gnd.n801 0.152939
R12152 gnd.n2312 gnd.n2310 0.152939
R12153 gnd.n3911 gnd.n1505 0.152939
R12154 gnd.n3907 gnd.n1505 0.152939
R12155 gnd.n3907 gnd.n3906 0.152939
R12156 gnd.n3906 gnd.n3905 0.152939
R12157 gnd.n3905 gnd.n1633 0.152939
R12158 gnd.n3898 gnd.n1633 0.152939
R12159 gnd.n3898 gnd.n3897 0.152939
R12160 gnd.n3897 gnd.n3896 0.152939
R12161 gnd.n3896 gnd.n3889 0.152939
R12162 gnd.n2912 gnd.n2911 0.152939
R12163 gnd.n2913 gnd.n2912 0.152939
R12164 gnd.n2913 gnd.n1960 0.152939
R12165 gnd.n2929 gnd.n1960 0.152939
R12166 gnd.n2930 gnd.n2929 0.152939
R12167 gnd.n2932 gnd.n2930 0.152939
R12168 gnd.n2932 gnd.n2931 0.152939
R12169 gnd.n2931 gnd.n1929 0.152939
R12170 gnd.n3051 gnd.n1929 0.152939
R12171 gnd.n3052 gnd.n3051 0.152939
R12172 gnd.n3053 gnd.n3052 0.152939
R12173 gnd.n3053 gnd.n1915 0.152939
R12174 gnd.n3067 gnd.n1915 0.152939
R12175 gnd.n3068 gnd.n3067 0.152939
R12176 gnd.n3069 gnd.n3068 0.152939
R12177 gnd.n3069 gnd.n1901 0.152939
R12178 gnd.n3083 gnd.n1901 0.152939
R12179 gnd.n3084 gnd.n3083 0.152939
R12180 gnd.n3085 gnd.n3084 0.152939
R12181 gnd.n3085 gnd.n1885 0.152939
R12182 gnd.n3100 gnd.n1885 0.152939
R12183 gnd.n3101 gnd.n3100 0.152939
R12184 gnd.n3103 gnd.n3101 0.152939
R12185 gnd.n3103 gnd.n3102 0.152939
R12186 gnd.n3102 gnd.n1854 0.152939
R12187 gnd.n3224 gnd.n1854 0.152939
R12188 gnd.n3225 gnd.n3224 0.152939
R12189 gnd.n3226 gnd.n3225 0.152939
R12190 gnd.n3226 gnd.n1841 0.152939
R12191 gnd.n3240 gnd.n1841 0.152939
R12192 gnd.n3241 gnd.n3240 0.152939
R12193 gnd.n3242 gnd.n3241 0.152939
R12194 gnd.n3242 gnd.n1829 0.152939
R12195 gnd.n3256 gnd.n1829 0.152939
R12196 gnd.n3257 gnd.n3256 0.152939
R12197 gnd.n3258 gnd.n3257 0.152939
R12198 gnd.n3258 gnd.n1815 0.152939
R12199 gnd.n3274 gnd.n1815 0.152939
R12200 gnd.n3275 gnd.n3274 0.152939
R12201 gnd.n3277 gnd.n3275 0.152939
R12202 gnd.n3277 gnd.n3276 0.152939
R12203 gnd.n3276 gnd.n1782 0.152939
R12204 gnd.n3395 gnd.n1782 0.152939
R12205 gnd.n3396 gnd.n3395 0.152939
R12206 gnd.n3397 gnd.n3396 0.152939
R12207 gnd.n3397 gnd.n1767 0.152939
R12208 gnd.n3411 gnd.n1767 0.152939
R12209 gnd.n3412 gnd.n3411 0.152939
R12210 gnd.n3413 gnd.n3412 0.152939
R12211 gnd.n3413 gnd.n1753 0.152939
R12212 gnd.n3427 gnd.n1753 0.152939
R12213 gnd.n3428 gnd.n3427 0.152939
R12214 gnd.n3429 gnd.n3428 0.152939
R12215 gnd.n3429 gnd.n1738 0.152939
R12216 gnd.n3445 gnd.n1738 0.152939
R12217 gnd.n3446 gnd.n3445 0.152939
R12218 gnd.n3448 gnd.n3446 0.152939
R12219 gnd.n3448 gnd.n3447 0.152939
R12220 gnd.n3447 gnd.n1708 0.152939
R12221 gnd.n3801 gnd.n1708 0.152939
R12222 gnd.n3802 gnd.n3801 0.152939
R12223 gnd.n3803 gnd.n3802 0.152939
R12224 gnd.n3803 gnd.n1695 0.152939
R12225 gnd.n3817 gnd.n1695 0.152939
R12226 gnd.n3818 gnd.n3817 0.152939
R12227 gnd.n3819 gnd.n3818 0.152939
R12228 gnd.n3819 gnd.n1682 0.152939
R12229 gnd.n3833 gnd.n1682 0.152939
R12230 gnd.n3834 gnd.n3833 0.152939
R12231 gnd.n3835 gnd.n3834 0.152939
R12232 gnd.n3835 gnd.n1668 0.152939
R12233 gnd.n3849 gnd.n1668 0.152939
R12234 gnd.n3850 gnd.n3849 0.152939
R12235 gnd.n3851 gnd.n3850 0.152939
R12236 gnd.n3851 gnd.n1654 0.152939
R12237 gnd.n3865 gnd.n1654 0.152939
R12238 gnd.n3866 gnd.n3865 0.152939
R12239 gnd.n3869 gnd.n3866 0.152939
R12240 gnd.n3869 gnd.n3868 0.152939
R12241 gnd.n3868 gnd.n3867 0.152939
R12242 gnd.n3867 gnd.n1641 0.152939
R12243 gnd.n3888 gnd.n1641 0.152939
R12244 gnd.n2876 gnd.n2006 0.152939
R12245 gnd.n2884 gnd.n2006 0.152939
R12246 gnd.n2885 gnd.n2884 0.152939
R12247 gnd.n2886 gnd.n2885 0.152939
R12248 gnd.n2886 gnd.n2002 0.152939
R12249 gnd.n2894 gnd.n2002 0.152939
R12250 gnd.n2895 gnd.n2894 0.152939
R12251 gnd.n2896 gnd.n2895 0.152939
R12252 gnd.n2896 gnd.n1976 0.152939
R12253 gnd.n2507 gnd.n2212 0.152939
R12254 gnd.n2508 gnd.n2507 0.152939
R12255 gnd.n2509 gnd.n2508 0.152939
R12256 gnd.n2509 gnd.n2206 0.152939
R12257 gnd.n2523 gnd.n2206 0.152939
R12258 gnd.n2524 gnd.n2523 0.152939
R12259 gnd.n2525 gnd.n2524 0.152939
R12260 gnd.n2525 gnd.n2199 0.152939
R12261 gnd.n2539 gnd.n2199 0.152939
R12262 gnd.n2540 gnd.n2539 0.152939
R12263 gnd.n2541 gnd.n2540 0.152939
R12264 gnd.n2541 gnd.n2193 0.152939
R12265 gnd.n2555 gnd.n2193 0.152939
R12266 gnd.n2556 gnd.n2555 0.152939
R12267 gnd.n2557 gnd.n2556 0.152939
R12268 gnd.n2557 gnd.n2187 0.152939
R12269 gnd.n2572 gnd.n2187 0.152939
R12270 gnd.n2573 gnd.n2572 0.152939
R12271 gnd.n2574 gnd.n2573 0.152939
R12272 gnd.n2574 gnd.n2008 0.152939
R12273 gnd.n4363 gnd.n1167 0.152939
R12274 gnd.n4359 gnd.n1167 0.152939
R12275 gnd.n4359 gnd.n4358 0.152939
R12276 gnd.n4358 gnd.n4357 0.152939
R12277 gnd.n4357 gnd.n1172 0.152939
R12278 gnd.n4353 gnd.n1172 0.152939
R12279 gnd.n4353 gnd.n4352 0.152939
R12280 gnd.n4352 gnd.n4351 0.152939
R12281 gnd.n4351 gnd.n1177 0.152939
R12282 gnd.n4347 gnd.n1177 0.152939
R12283 gnd.n4347 gnd.n4346 0.152939
R12284 gnd.n4346 gnd.n4345 0.152939
R12285 gnd.n4345 gnd.n1182 0.152939
R12286 gnd.n4341 gnd.n1182 0.152939
R12287 gnd.n4341 gnd.n4340 0.152939
R12288 gnd.n4340 gnd.n4339 0.152939
R12289 gnd.n4339 gnd.n1187 0.152939
R12290 gnd.n4335 gnd.n1187 0.152939
R12291 gnd.n4335 gnd.n4334 0.152939
R12292 gnd.n4334 gnd.n4333 0.152939
R12293 gnd.n4333 gnd.n1192 0.152939
R12294 gnd.n4329 gnd.n1192 0.152939
R12295 gnd.n4329 gnd.n4328 0.152939
R12296 gnd.n4328 gnd.n4327 0.152939
R12297 gnd.n4327 gnd.n1197 0.152939
R12298 gnd.n4323 gnd.n1197 0.152939
R12299 gnd.n4323 gnd.n4322 0.152939
R12300 gnd.n4322 gnd.n4321 0.152939
R12301 gnd.n4321 gnd.n1202 0.152939
R12302 gnd.n4317 gnd.n1202 0.152939
R12303 gnd.n4317 gnd.n4316 0.152939
R12304 gnd.n4316 gnd.n4315 0.152939
R12305 gnd.n4315 gnd.n1207 0.152939
R12306 gnd.n4311 gnd.n1207 0.152939
R12307 gnd.n4311 gnd.n4310 0.152939
R12308 gnd.n4310 gnd.n4309 0.152939
R12309 gnd.n4309 gnd.n1212 0.152939
R12310 gnd.n4305 gnd.n1212 0.152939
R12311 gnd.n4305 gnd.n4304 0.152939
R12312 gnd.n4304 gnd.n4303 0.152939
R12313 gnd.n4303 gnd.n1217 0.152939
R12314 gnd.n4299 gnd.n1217 0.152939
R12315 gnd.n4299 gnd.n4298 0.152939
R12316 gnd.n4298 gnd.n4297 0.152939
R12317 gnd.n4297 gnd.n1222 0.152939
R12318 gnd.n4293 gnd.n1222 0.152939
R12319 gnd.n4293 gnd.n4292 0.152939
R12320 gnd.n4292 gnd.n4291 0.152939
R12321 gnd.n4291 gnd.n1227 0.152939
R12322 gnd.n4287 gnd.n1227 0.152939
R12323 gnd.n4287 gnd.n4286 0.152939
R12324 gnd.n4286 gnd.n4285 0.152939
R12325 gnd.n4285 gnd.n1232 0.152939
R12326 gnd.n4281 gnd.n1232 0.152939
R12327 gnd.n4281 gnd.n4280 0.152939
R12328 gnd.n4280 gnd.n4279 0.152939
R12329 gnd.n4279 gnd.n1237 0.152939
R12330 gnd.n4275 gnd.n1237 0.152939
R12331 gnd.n4275 gnd.n4274 0.152939
R12332 gnd.n4274 gnd.n4273 0.152939
R12333 gnd.n4273 gnd.n1242 0.152939
R12334 gnd.n4269 gnd.n1242 0.152939
R12335 gnd.n4269 gnd.n4268 0.152939
R12336 gnd.n4268 gnd.n4267 0.152939
R12337 gnd.n4267 gnd.n1247 0.152939
R12338 gnd.n4263 gnd.n1247 0.152939
R12339 gnd.n4263 gnd.n4262 0.152939
R12340 gnd.n4262 gnd.n4261 0.152939
R12341 gnd.n4261 gnd.n1252 0.152939
R12342 gnd.n4257 gnd.n1252 0.152939
R12343 gnd.n4257 gnd.n4256 0.152939
R12344 gnd.n4256 gnd.n4255 0.152939
R12345 gnd.n4255 gnd.n1257 0.152939
R12346 gnd.n4251 gnd.n1257 0.152939
R12347 gnd.n4251 gnd.n4250 0.152939
R12348 gnd.n4250 gnd.n4249 0.152939
R12349 gnd.n4249 gnd.n1262 0.152939
R12350 gnd.n4245 gnd.n1262 0.152939
R12351 gnd.n4245 gnd.n4244 0.152939
R12352 gnd.n4244 gnd.n4243 0.152939
R12353 gnd.n4243 gnd.n1267 0.152939
R12354 gnd.n1270 gnd.n1267 0.152939
R12355 gnd.n4150 gnd.n4149 0.152939
R12356 gnd.n4149 gnd.n4148 0.152939
R12357 gnd.n4148 gnd.n1369 0.152939
R12358 gnd.n4144 gnd.n1369 0.152939
R12359 gnd.n4144 gnd.n4143 0.152939
R12360 gnd.n4143 gnd.n4142 0.152939
R12361 gnd.n4142 gnd.n1374 0.152939
R12362 gnd.n4138 gnd.n1374 0.152939
R12363 gnd.n4138 gnd.n4137 0.152939
R12364 gnd.n4137 gnd.n4136 0.152939
R12365 gnd.n4136 gnd.n1379 0.152939
R12366 gnd.n4132 gnd.n1379 0.152939
R12367 gnd.n4132 gnd.n4131 0.152939
R12368 gnd.n4131 gnd.n4130 0.152939
R12369 gnd.n4130 gnd.n1384 0.152939
R12370 gnd.n4126 gnd.n1384 0.152939
R12371 gnd.n4126 gnd.n4125 0.152939
R12372 gnd.n4125 gnd.n4124 0.152939
R12373 gnd.n4124 gnd.n1389 0.152939
R12374 gnd.n4120 gnd.n1389 0.152939
R12375 gnd.n4120 gnd.n4119 0.152939
R12376 gnd.n4119 gnd.n4118 0.152939
R12377 gnd.n4118 gnd.n226 0.152939
R12378 gnd.n6747 gnd.n226 0.152939
R12379 gnd.n6748 gnd.n6747 0.152939
R12380 gnd.n6749 gnd.n6748 0.152939
R12381 gnd.n6749 gnd.n205 0.152939
R12382 gnd.n6763 gnd.n205 0.152939
R12383 gnd.n6764 gnd.n6763 0.152939
R12384 gnd.n6765 gnd.n6764 0.152939
R12385 gnd.n6765 gnd.n191 0.152939
R12386 gnd.n6779 gnd.n191 0.152939
R12387 gnd.n6780 gnd.n6779 0.152939
R12388 gnd.n6781 gnd.n6780 0.152939
R12389 gnd.n6781 gnd.n176 0.152939
R12390 gnd.n6795 gnd.n176 0.152939
R12391 gnd.n6796 gnd.n6795 0.152939
R12392 gnd.n6871 gnd.n6796 0.152939
R12393 gnd.n6871 gnd.n6870 0.152939
R12394 gnd.n6870 gnd.n6869 0.152939
R12395 gnd.n6869 gnd.n6797 0.152939
R12396 gnd.n6865 gnd.n6797 0.152939
R12397 gnd.n6864 gnd.n6799 0.152939
R12398 gnd.n6860 gnd.n6799 0.152939
R12399 gnd.n6860 gnd.n6859 0.152939
R12400 gnd.n6859 gnd.n6858 0.152939
R12401 gnd.n6858 gnd.n6805 0.152939
R12402 gnd.n6854 gnd.n6805 0.152939
R12403 gnd.n6854 gnd.n6853 0.152939
R12404 gnd.n6853 gnd.n6852 0.152939
R12405 gnd.n6852 gnd.n6813 0.152939
R12406 gnd.n6848 gnd.n6813 0.152939
R12407 gnd.n6848 gnd.n6847 0.152939
R12408 gnd.n6847 gnd.n6846 0.152939
R12409 gnd.n6846 gnd.n6821 0.152939
R12410 gnd.n6842 gnd.n6821 0.152939
R12411 gnd.n6842 gnd.n6841 0.152939
R12412 gnd.n6841 gnd.n6840 0.152939
R12413 gnd.n6840 gnd.n6829 0.152939
R12414 gnd.n6829 gnd.n78 0.152939
R12415 gnd.n3914 gnd.n3913 0.152939
R12416 gnd.n3914 gnd.n1492 0.152939
R12417 gnd.n3987 gnd.n1492 0.152939
R12418 gnd.n3988 gnd.n3987 0.152939
R12419 gnd.n3990 gnd.n3988 0.152939
R12420 gnd.n3990 gnd.n3989 0.152939
R12421 gnd.n3989 gnd.n1466 0.152939
R12422 gnd.n4019 gnd.n1466 0.152939
R12423 gnd.n4020 gnd.n4019 0.152939
R12424 gnd.n4022 gnd.n4020 0.152939
R12425 gnd.n4022 gnd.n4021 0.152939
R12426 gnd.n4021 gnd.n1440 0.152939
R12427 gnd.n4054 gnd.n1440 0.152939
R12428 gnd.n4055 gnd.n4054 0.152939
R12429 gnd.n4056 gnd.n4055 0.152939
R12430 gnd.n4056 gnd.n1412 0.152939
R12431 gnd.n4085 gnd.n1412 0.152939
R12432 gnd.n4086 gnd.n4085 0.152939
R12433 gnd.n4087 gnd.n4086 0.152939
R12434 gnd.n4087 gnd.n51 0.152939
R12435 gnd.n6996 gnd.n51 0.152939
R12436 gnd.n6996 gnd.n6995 0.152939
R12437 gnd.n6995 gnd.n53 0.152939
R12438 gnd.n6991 gnd.n53 0.152939
R12439 gnd.n6991 gnd.n6990 0.152939
R12440 gnd.n6990 gnd.n6989 0.152939
R12441 gnd.n6989 gnd.n58 0.152939
R12442 gnd.n6985 gnd.n58 0.152939
R12443 gnd.n6985 gnd.n6984 0.152939
R12444 gnd.n6984 gnd.n6983 0.152939
R12445 gnd.n6983 gnd.n63 0.152939
R12446 gnd.n6979 gnd.n63 0.152939
R12447 gnd.n6979 gnd.n6978 0.152939
R12448 gnd.n6978 gnd.n6977 0.152939
R12449 gnd.n6977 gnd.n68 0.152939
R12450 gnd.n6973 gnd.n68 0.152939
R12451 gnd.n6973 gnd.n6972 0.152939
R12452 gnd.n6972 gnd.n6971 0.152939
R12453 gnd.n6971 gnd.n73 0.152939
R12454 gnd.n6967 gnd.n73 0.152939
R12455 gnd.n6967 gnd.n6966 0.152939
R12456 gnd.n6966 gnd.n6965 0.152939
R12457 gnd.n3912 gnd.n3911 0.151415
R12458 gnd.n2876 gnd.n2875 0.151415
R12459 gnd.n2493 gnd.n2492 0.145814
R12460 gnd.n2493 gnd.n2212 0.145814
R12461 gnd.n2321 gnd.n2230 0.128549
R12462 gnd.n1435 gnd.n213 0.128549
R12463 gnd.n4766 gnd.n0 0.127478
R12464 gnd.n5375 gnd.n4767 0.0767195
R12465 gnd.n5291 gnd.n4767 0.0767195
R12466 gnd.n4365 gnd.n4364 0.063
R12467 gnd.n1549 gnd.n1368 0.063
R12468 gnd.n5883 gnd.n4599 0.0477147
R12469 gnd.n5041 gnd.n4937 0.0442063
R12470 gnd.n5055 gnd.n4937 0.0442063
R12471 gnd.n5056 gnd.n5055 0.0442063
R12472 gnd.n5057 gnd.n5056 0.0442063
R12473 gnd.n5057 gnd.n4925 0.0442063
R12474 gnd.n5071 gnd.n4925 0.0442063
R12475 gnd.n5072 gnd.n5071 0.0442063
R12476 gnd.n5073 gnd.n5072 0.0442063
R12477 gnd.n5073 gnd.n4912 0.0442063
R12478 gnd.n5169 gnd.n4912 0.0442063
R12479 gnd.n5172 gnd.n5171 0.0344674
R12480 gnd.n1511 gnd.n1504 0.0344674
R12481 gnd.n2874 gnd.n2873 0.0344674
R12482 gnd.n4905 gnd.n4904 0.0269946
R12483 gnd.n5182 gnd.n4902 0.0269946
R12484 gnd.n5181 gnd.n4903 0.0269946
R12485 gnd.n5201 gnd.n4884 0.0269946
R12486 gnd.n5203 gnd.n5202 0.0269946
R12487 gnd.n5204 gnd.n4882 0.0269946
R12488 gnd.n5211 gnd.n5207 0.0269946
R12489 gnd.n5210 gnd.n5209 0.0269946
R12490 gnd.n5208 gnd.n4861 0.0269946
R12491 gnd.n5235 gnd.n4862 0.0269946
R12492 gnd.n5234 gnd.n4863 0.0269946
R12493 gnd.n5267 gnd.n4837 0.0269946
R12494 gnd.n5269 gnd.n5268 0.0269946
R12495 gnd.n5270 gnd.n4829 0.0269946
R12496 gnd.n4833 gnd.n4830 0.0269946
R12497 gnd.n5280 gnd.n4831 0.0269946
R12498 gnd.n5279 gnd.n4832 0.0269946
R12499 gnd.n5325 gnd.n4805 0.0269946
R12500 gnd.n5327 gnd.n5326 0.0269946
R12501 gnd.n5336 gnd.n4798 0.0269946
R12502 gnd.n5338 gnd.n5337 0.0269946
R12503 gnd.n5339 gnd.n4796 0.0269946
R12504 gnd.n5346 gnd.n5342 0.0269946
R12505 gnd.n5345 gnd.n5344 0.0269946
R12506 gnd.n5343 gnd.n4775 0.0269946
R12507 gnd.n5368 gnd.n4776 0.0269946
R12508 gnd.n5367 gnd.n4777 0.0269946
R12509 gnd.n5410 gnd.n4714 0.0269946
R12510 gnd.n5412 gnd.n5411 0.0269946
R12511 gnd.n5421 gnd.n4707 0.0269946
R12512 gnd.n5423 gnd.n5422 0.0269946
R12513 gnd.n5424 gnd.n4705 0.0269946
R12514 gnd.n5430 gnd.n5427 0.0269946
R12515 gnd.n5429 gnd.n5428 0.0269946
R12516 gnd.n5455 gnd.n4684 0.0269946
R12517 gnd.n5454 gnd.n4685 0.0269946
R12518 gnd.n5481 gnd.n4670 0.0269946
R12519 gnd.n5483 gnd.n5482 0.0269946
R12520 gnd.n5484 gnd.n4656 0.0269946
R12521 gnd.n5506 gnd.n4654 0.0269946
R12522 gnd.n5508 gnd.n5507 0.0269946
R12523 gnd.n5510 gnd.n5509 0.0269946
R12524 gnd.n5519 gnd.n4646 0.0269946
R12525 gnd.n5521 gnd.n5520 0.0269946
R12526 gnd.n5522 gnd.n821 0.0269946
R12527 gnd.n4637 gnd.n822 0.0269946
R12528 gnd.n4639 gnd.n823 0.0269946
R12529 gnd.n5549 gnd.n5548 0.0269946
R12530 gnd.n5808 gnd.n846 0.0269946
R12531 gnd.n5810 gnd.n847 0.0269946
R12532 gnd.n5812 gnd.n848 0.0269946
R12533 gnd.n5814 gnd.n5813 0.0269946
R12534 gnd.n275 gnd.n213 0.0248902
R12535 gnd.n2321 gnd.n2320 0.0248902
R12536 gnd.n1550 gnd.n1549 0.0246168
R12537 gnd.n4364 gnd.n1166 0.0246168
R12538 gnd.n5171 gnd.n5170 0.0202011
R12539 gnd.n1550 gnd.n1547 0.0174837
R12540 gnd.n1555 gnd.n1547 0.0174837
R12541 gnd.n1556 gnd.n1555 0.0174837
R12542 gnd.n1556 gnd.n1545 0.0174837
R12543 gnd.n1563 gnd.n1545 0.0174837
R12544 gnd.n1565 gnd.n1563 0.0174837
R12545 gnd.n1565 gnd.n1564 0.0174837
R12546 gnd.n1564 gnd.n1540 0.0174837
R12547 gnd.n1572 gnd.n1540 0.0174837
R12548 gnd.n1572 gnd.n1571 0.0174837
R12549 gnd.n1571 gnd.n1541 0.0174837
R12550 gnd.n1541 gnd.n1536 0.0174837
R12551 gnd.n1580 gnd.n1536 0.0174837
R12552 gnd.n1582 gnd.n1580 0.0174837
R12553 gnd.n1582 gnd.n1581 0.0174837
R12554 gnd.n1581 gnd.n1531 0.0174837
R12555 gnd.n1589 gnd.n1531 0.0174837
R12556 gnd.n1589 gnd.n1588 0.0174837
R12557 gnd.n1588 gnd.n1532 0.0174837
R12558 gnd.n1532 gnd.n1527 0.0174837
R12559 gnd.n1597 gnd.n1527 0.0174837
R12560 gnd.n1599 gnd.n1597 0.0174837
R12561 gnd.n1599 gnd.n1598 0.0174837
R12562 gnd.n1598 gnd.n1522 0.0174837
R12563 gnd.n1606 gnd.n1522 0.0174837
R12564 gnd.n1606 gnd.n1605 0.0174837
R12565 gnd.n1605 gnd.n1523 0.0174837
R12566 gnd.n1523 gnd.n1518 0.0174837
R12567 gnd.n1614 gnd.n1518 0.0174837
R12568 gnd.n1616 gnd.n1614 0.0174837
R12569 gnd.n1616 gnd.n1615 0.0174837
R12570 gnd.n1615 gnd.n1510 0.0174837
R12571 gnd.n1621 gnd.n1510 0.0174837
R12572 gnd.n1621 gnd.n1620 0.0174837
R12573 gnd.n1620 gnd.n1511 0.0174837
R12574 gnd.n2056 gnd.n1166 0.0174837
R12575 gnd.n2056 gnd.n2055 0.0174837
R12576 gnd.n2062 gnd.n2055 0.0174837
R12577 gnd.n2063 gnd.n2062 0.0174837
R12578 gnd.n2063 gnd.n2049 0.0174837
R12579 gnd.n2068 gnd.n2049 0.0174837
R12580 gnd.n2069 gnd.n2068 0.0174837
R12581 gnd.n2069 gnd.n2047 0.0174837
R12582 gnd.n2074 gnd.n2047 0.0174837
R12583 gnd.n2075 gnd.n2074 0.0174837
R12584 gnd.n2075 gnd.n2045 0.0174837
R12585 gnd.n2080 gnd.n2045 0.0174837
R12586 gnd.n2081 gnd.n2080 0.0174837
R12587 gnd.n2081 gnd.n2041 0.0174837
R12588 gnd.n2086 gnd.n2041 0.0174837
R12589 gnd.n2087 gnd.n2086 0.0174837
R12590 gnd.n2087 gnd.n2037 0.0174837
R12591 gnd.n2092 gnd.n2037 0.0174837
R12592 gnd.n2093 gnd.n2092 0.0174837
R12593 gnd.n2093 gnd.n2035 0.0174837
R12594 gnd.n2098 gnd.n2035 0.0174837
R12595 gnd.n2099 gnd.n2098 0.0174837
R12596 gnd.n2099 gnd.n2033 0.0174837
R12597 gnd.n2104 gnd.n2033 0.0174837
R12598 gnd.n2106 gnd.n2104 0.0174837
R12599 gnd.n2106 gnd.n2105 0.0174837
R12600 gnd.n2105 gnd.n2028 0.0174837
R12601 gnd.n2113 gnd.n2028 0.0174837
R12602 gnd.n2113 gnd.n2112 0.0174837
R12603 gnd.n2112 gnd.n2029 0.0174837
R12604 gnd.n2029 gnd.n2013 0.0174837
R12605 gnd.n2867 gnd.n2013 0.0174837
R12606 gnd.n2868 gnd.n2867 0.0174837
R12607 gnd.n2868 gnd.n2009 0.0174837
R12608 gnd.n2873 gnd.n2009 0.0174837
R12609 gnd.n5170 gnd.n5169 0.0148637
R12610 gnd.n5806 gnd.n5550 0.0144266
R12611 gnd.n5807 gnd.n5806 0.0130679
R12612 gnd.n5172 gnd.n4905 0.00797283
R12613 gnd.n4904 gnd.n4902 0.00797283
R12614 gnd.n5182 gnd.n5181 0.00797283
R12615 gnd.n4903 gnd.n4884 0.00797283
R12616 gnd.n5202 gnd.n5201 0.00797283
R12617 gnd.n5204 gnd.n5203 0.00797283
R12618 gnd.n5207 gnd.n4882 0.00797283
R12619 gnd.n5211 gnd.n5210 0.00797283
R12620 gnd.n5209 gnd.n5208 0.00797283
R12621 gnd.n4862 gnd.n4861 0.00797283
R12622 gnd.n5235 gnd.n5234 0.00797283
R12623 gnd.n4863 gnd.n4837 0.00797283
R12624 gnd.n5268 gnd.n5267 0.00797283
R12625 gnd.n5270 gnd.n5269 0.00797283
R12626 gnd.n4833 gnd.n4829 0.00797283
R12627 gnd.n4831 gnd.n4830 0.00797283
R12628 gnd.n5280 gnd.n5279 0.00797283
R12629 gnd.n4832 gnd.n4805 0.00797283
R12630 gnd.n5327 gnd.n5325 0.00797283
R12631 gnd.n5326 gnd.n4798 0.00797283
R12632 gnd.n5337 gnd.n5336 0.00797283
R12633 gnd.n5339 gnd.n5338 0.00797283
R12634 gnd.n5342 gnd.n4796 0.00797283
R12635 gnd.n5346 gnd.n5345 0.00797283
R12636 gnd.n5344 gnd.n5343 0.00797283
R12637 gnd.n4776 gnd.n4775 0.00797283
R12638 gnd.n5368 gnd.n5367 0.00797283
R12639 gnd.n4777 gnd.n4714 0.00797283
R12640 gnd.n5412 gnd.n5410 0.00797283
R12641 gnd.n5411 gnd.n4707 0.00797283
R12642 gnd.n5422 gnd.n5421 0.00797283
R12643 gnd.n5424 gnd.n5423 0.00797283
R12644 gnd.n5427 gnd.n4705 0.00797283
R12645 gnd.n5430 gnd.n5429 0.00797283
R12646 gnd.n5428 gnd.n4684 0.00797283
R12647 gnd.n5455 gnd.n5454 0.00797283
R12648 gnd.n4685 gnd.n4670 0.00797283
R12649 gnd.n5482 gnd.n5481 0.00797283
R12650 gnd.n5484 gnd.n5483 0.00797283
R12651 gnd.n4656 gnd.n4654 0.00797283
R12652 gnd.n5507 gnd.n5506 0.00797283
R12653 gnd.n5510 gnd.n5508 0.00797283
R12654 gnd.n5509 gnd.n4646 0.00797283
R12655 gnd.n5520 gnd.n5519 0.00797283
R12656 gnd.n5522 gnd.n5521 0.00797283
R12657 gnd.n4637 gnd.n821 0.00797283
R12658 gnd.n4639 gnd.n822 0.00797283
R12659 gnd.n5548 gnd.n823 0.00797283
R12660 gnd.n5550 gnd.n5549 0.00797283
R12661 gnd.n5808 gnd.n5807 0.00797283
R12662 gnd.n5810 gnd.n846 0.00797283
R12663 gnd.n5812 gnd.n847 0.00797283
R12664 gnd.n5814 gnd.n848 0.00797283
R12665 gnd.n5813 gnd.n4599 0.00797283
R12666 gnd.n4119 gnd.n1395 0.00614909
R12667 gnd.n2499 gnd.n2216 0.00614909
R12668 gnd.n3912 gnd.n1504 0.000839674
R12669 gnd.n2875 gnd.n2874 0.000839674
R12670 commonsourceibias.n25 commonsourceibias.t46 230.006
R12671 commonsourceibias.n91 commonsourceibias.t62 230.006
R12672 commonsourceibias.n154 commonsourceibias.t54 230.006
R12673 commonsourceibias.n258 commonsourceibias.t16 230.006
R12674 commonsourceibias.n217 commonsourceibias.t75 230.006
R12675 commonsourceibias.n355 commonsourceibias.t65 230.006
R12676 commonsourceibias.n70 commonsourceibias.t32 207.983
R12677 commonsourceibias.n136 commonsourceibias.t71 207.983
R12678 commonsourceibias.n199 commonsourceibias.t61 207.983
R12679 commonsourceibias.n304 commonsourceibias.t2 207.983
R12680 commonsourceibias.n338 commonsourceibias.t84 207.983
R12681 commonsourceibias.n401 commonsourceibias.t73 207.983
R12682 commonsourceibias.n10 commonsourceibias.t14 168.701
R12683 commonsourceibias.n63 commonsourceibias.t24 168.701
R12684 commonsourceibias.n57 commonsourceibias.t30 168.701
R12685 commonsourceibias.n16 commonsourceibias.t20 168.701
R12686 commonsourceibias.n49 commonsourceibias.t36 168.701
R12687 commonsourceibias.n43 commonsourceibias.t44 168.701
R12688 commonsourceibias.n19 commonsourceibias.t26 168.701
R12689 commonsourceibias.n21 commonsourceibias.t34 168.701
R12690 commonsourceibias.n23 commonsourceibias.t10 168.701
R12691 commonsourceibias.n26 commonsourceibias.t40 168.701
R12692 commonsourceibias.n1 commonsourceibias.t81 168.701
R12693 commonsourceibias.n129 commonsourceibias.t55 168.701
R12694 commonsourceibias.n123 commonsourceibias.t53 168.701
R12695 commonsourceibias.n7 commonsourceibias.t76 168.701
R12696 commonsourceibias.n115 commonsourceibias.t86 168.701
R12697 commonsourceibias.n109 commonsourceibias.t50 168.701
R12698 commonsourceibias.n85 commonsourceibias.t69 168.701
R12699 commonsourceibias.n87 commonsourceibias.t67 168.701
R12700 commonsourceibias.n89 commonsourceibias.t78 168.701
R12701 commonsourceibias.n92 commonsourceibias.t64 168.701
R12702 commonsourceibias.n155 commonsourceibias.t57 168.701
R12703 commonsourceibias.n152 commonsourceibias.t68 168.701
R12704 commonsourceibias.n150 commonsourceibias.t58 168.701
R12705 commonsourceibias.n148 commonsourceibias.t60 168.701
R12706 commonsourceibias.n172 commonsourceibias.t91 168.701
R12707 commonsourceibias.n178 commonsourceibias.t77 168.701
R12708 commonsourceibias.n145 commonsourceibias.t66 168.701
R12709 commonsourceibias.n186 commonsourceibias.t95 168.701
R12710 commonsourceibias.n192 commonsourceibias.t49 168.701
R12711 commonsourceibias.n139 commonsourceibias.t72 168.701
R12712 commonsourceibias.n259 commonsourceibias.t8 168.701
R12713 commonsourceibias.n256 commonsourceibias.t18 168.701
R12714 commonsourceibias.n254 commonsourceibias.t4 168.701
R12715 commonsourceibias.n252 commonsourceibias.t42 168.701
R12716 commonsourceibias.n276 commonsourceibias.t12 168.701
R12717 commonsourceibias.n282 commonsourceibias.t6 168.701
R12718 commonsourceibias.n284 commonsourceibias.t28 168.701
R12719 commonsourceibias.n291 commonsourceibias.t0 168.701
R12720 commonsourceibias.n297 commonsourceibias.t38 168.701
R12721 commonsourceibias.n244 commonsourceibias.t22 168.701
R12722 commonsourceibias.n203 commonsourceibias.t92 168.701
R12723 commonsourceibias.n331 commonsourceibias.t51 168.701
R12724 commonsourceibias.n325 commonsourceibias.t63 168.701
R12725 commonsourceibias.n318 commonsourceibias.t88 168.701
R12726 commonsourceibias.n316 commonsourceibias.t48 168.701
R12727 commonsourceibias.n218 commonsourceibias.t59 168.701
R12728 commonsourceibias.n215 commonsourceibias.t90 168.701
R12729 commonsourceibias.n213 commonsourceibias.t80 168.701
R12730 commonsourceibias.n211 commonsourceibias.t83 168.701
R12731 commonsourceibias.n235 commonsourceibias.t94 168.701
R12732 commonsourceibias.n356 commonsourceibias.t52 168.701
R12733 commonsourceibias.n353 commonsourceibias.t82 168.701
R12734 commonsourceibias.n351 commonsourceibias.t70 168.701
R12735 commonsourceibias.n349 commonsourceibias.t74 168.701
R12736 commonsourceibias.n373 commonsourceibias.t87 168.701
R12737 commonsourceibias.n379 commonsourceibias.t89 168.701
R12738 commonsourceibias.n381 commonsourceibias.t79 168.701
R12739 commonsourceibias.n388 commonsourceibias.t56 168.701
R12740 commonsourceibias.n394 commonsourceibias.t93 168.701
R12741 commonsourceibias.n341 commonsourceibias.t85 168.701
R12742 commonsourceibias.n27 commonsourceibias.n24 161.3
R12743 commonsourceibias.n29 commonsourceibias.n28 161.3
R12744 commonsourceibias.n31 commonsourceibias.n30 161.3
R12745 commonsourceibias.n32 commonsourceibias.n22 161.3
R12746 commonsourceibias.n34 commonsourceibias.n33 161.3
R12747 commonsourceibias.n36 commonsourceibias.n35 161.3
R12748 commonsourceibias.n37 commonsourceibias.n20 161.3
R12749 commonsourceibias.n39 commonsourceibias.n38 161.3
R12750 commonsourceibias.n41 commonsourceibias.n40 161.3
R12751 commonsourceibias.n42 commonsourceibias.n18 161.3
R12752 commonsourceibias.n45 commonsourceibias.n44 161.3
R12753 commonsourceibias.n46 commonsourceibias.n17 161.3
R12754 commonsourceibias.n48 commonsourceibias.n47 161.3
R12755 commonsourceibias.n50 commonsourceibias.n15 161.3
R12756 commonsourceibias.n52 commonsourceibias.n51 161.3
R12757 commonsourceibias.n53 commonsourceibias.n14 161.3
R12758 commonsourceibias.n55 commonsourceibias.n54 161.3
R12759 commonsourceibias.n56 commonsourceibias.n13 161.3
R12760 commonsourceibias.n59 commonsourceibias.n58 161.3
R12761 commonsourceibias.n60 commonsourceibias.n12 161.3
R12762 commonsourceibias.n62 commonsourceibias.n61 161.3
R12763 commonsourceibias.n64 commonsourceibias.n11 161.3
R12764 commonsourceibias.n66 commonsourceibias.n65 161.3
R12765 commonsourceibias.n68 commonsourceibias.n67 161.3
R12766 commonsourceibias.n69 commonsourceibias.n9 161.3
R12767 commonsourceibias.n93 commonsourceibias.n90 161.3
R12768 commonsourceibias.n95 commonsourceibias.n94 161.3
R12769 commonsourceibias.n97 commonsourceibias.n96 161.3
R12770 commonsourceibias.n98 commonsourceibias.n88 161.3
R12771 commonsourceibias.n100 commonsourceibias.n99 161.3
R12772 commonsourceibias.n102 commonsourceibias.n101 161.3
R12773 commonsourceibias.n103 commonsourceibias.n86 161.3
R12774 commonsourceibias.n105 commonsourceibias.n104 161.3
R12775 commonsourceibias.n107 commonsourceibias.n106 161.3
R12776 commonsourceibias.n108 commonsourceibias.n84 161.3
R12777 commonsourceibias.n111 commonsourceibias.n110 161.3
R12778 commonsourceibias.n112 commonsourceibias.n8 161.3
R12779 commonsourceibias.n114 commonsourceibias.n113 161.3
R12780 commonsourceibias.n116 commonsourceibias.n6 161.3
R12781 commonsourceibias.n118 commonsourceibias.n117 161.3
R12782 commonsourceibias.n119 commonsourceibias.n5 161.3
R12783 commonsourceibias.n121 commonsourceibias.n120 161.3
R12784 commonsourceibias.n122 commonsourceibias.n4 161.3
R12785 commonsourceibias.n125 commonsourceibias.n124 161.3
R12786 commonsourceibias.n126 commonsourceibias.n3 161.3
R12787 commonsourceibias.n128 commonsourceibias.n127 161.3
R12788 commonsourceibias.n130 commonsourceibias.n2 161.3
R12789 commonsourceibias.n132 commonsourceibias.n131 161.3
R12790 commonsourceibias.n134 commonsourceibias.n133 161.3
R12791 commonsourceibias.n135 commonsourceibias.n0 161.3
R12792 commonsourceibias.n198 commonsourceibias.n138 161.3
R12793 commonsourceibias.n197 commonsourceibias.n196 161.3
R12794 commonsourceibias.n195 commonsourceibias.n194 161.3
R12795 commonsourceibias.n193 commonsourceibias.n140 161.3
R12796 commonsourceibias.n191 commonsourceibias.n190 161.3
R12797 commonsourceibias.n189 commonsourceibias.n141 161.3
R12798 commonsourceibias.n188 commonsourceibias.n187 161.3
R12799 commonsourceibias.n185 commonsourceibias.n142 161.3
R12800 commonsourceibias.n184 commonsourceibias.n183 161.3
R12801 commonsourceibias.n182 commonsourceibias.n143 161.3
R12802 commonsourceibias.n181 commonsourceibias.n180 161.3
R12803 commonsourceibias.n179 commonsourceibias.n144 161.3
R12804 commonsourceibias.n177 commonsourceibias.n176 161.3
R12805 commonsourceibias.n175 commonsourceibias.n146 161.3
R12806 commonsourceibias.n174 commonsourceibias.n173 161.3
R12807 commonsourceibias.n171 commonsourceibias.n147 161.3
R12808 commonsourceibias.n170 commonsourceibias.n169 161.3
R12809 commonsourceibias.n168 commonsourceibias.n167 161.3
R12810 commonsourceibias.n166 commonsourceibias.n149 161.3
R12811 commonsourceibias.n165 commonsourceibias.n164 161.3
R12812 commonsourceibias.n163 commonsourceibias.n162 161.3
R12813 commonsourceibias.n161 commonsourceibias.n151 161.3
R12814 commonsourceibias.n160 commonsourceibias.n159 161.3
R12815 commonsourceibias.n158 commonsourceibias.n157 161.3
R12816 commonsourceibias.n156 commonsourceibias.n153 161.3
R12817 commonsourceibias.n303 commonsourceibias.n243 161.3
R12818 commonsourceibias.n302 commonsourceibias.n301 161.3
R12819 commonsourceibias.n300 commonsourceibias.n299 161.3
R12820 commonsourceibias.n298 commonsourceibias.n245 161.3
R12821 commonsourceibias.n296 commonsourceibias.n295 161.3
R12822 commonsourceibias.n294 commonsourceibias.n246 161.3
R12823 commonsourceibias.n293 commonsourceibias.n292 161.3
R12824 commonsourceibias.n290 commonsourceibias.n247 161.3
R12825 commonsourceibias.n289 commonsourceibias.n288 161.3
R12826 commonsourceibias.n287 commonsourceibias.n248 161.3
R12827 commonsourceibias.n286 commonsourceibias.n285 161.3
R12828 commonsourceibias.n283 commonsourceibias.n249 161.3
R12829 commonsourceibias.n281 commonsourceibias.n280 161.3
R12830 commonsourceibias.n279 commonsourceibias.n250 161.3
R12831 commonsourceibias.n278 commonsourceibias.n277 161.3
R12832 commonsourceibias.n275 commonsourceibias.n251 161.3
R12833 commonsourceibias.n274 commonsourceibias.n273 161.3
R12834 commonsourceibias.n272 commonsourceibias.n271 161.3
R12835 commonsourceibias.n270 commonsourceibias.n253 161.3
R12836 commonsourceibias.n269 commonsourceibias.n268 161.3
R12837 commonsourceibias.n267 commonsourceibias.n266 161.3
R12838 commonsourceibias.n265 commonsourceibias.n255 161.3
R12839 commonsourceibias.n264 commonsourceibias.n263 161.3
R12840 commonsourceibias.n262 commonsourceibias.n261 161.3
R12841 commonsourceibias.n260 commonsourceibias.n257 161.3
R12842 commonsourceibias.n237 commonsourceibias.n236 161.3
R12843 commonsourceibias.n234 commonsourceibias.n210 161.3
R12844 commonsourceibias.n233 commonsourceibias.n232 161.3
R12845 commonsourceibias.n231 commonsourceibias.n230 161.3
R12846 commonsourceibias.n229 commonsourceibias.n212 161.3
R12847 commonsourceibias.n228 commonsourceibias.n227 161.3
R12848 commonsourceibias.n226 commonsourceibias.n225 161.3
R12849 commonsourceibias.n224 commonsourceibias.n214 161.3
R12850 commonsourceibias.n223 commonsourceibias.n222 161.3
R12851 commonsourceibias.n221 commonsourceibias.n220 161.3
R12852 commonsourceibias.n219 commonsourceibias.n216 161.3
R12853 commonsourceibias.n313 commonsourceibias.n209 161.3
R12854 commonsourceibias.n337 commonsourceibias.n202 161.3
R12855 commonsourceibias.n336 commonsourceibias.n335 161.3
R12856 commonsourceibias.n334 commonsourceibias.n333 161.3
R12857 commonsourceibias.n332 commonsourceibias.n204 161.3
R12858 commonsourceibias.n330 commonsourceibias.n329 161.3
R12859 commonsourceibias.n328 commonsourceibias.n205 161.3
R12860 commonsourceibias.n327 commonsourceibias.n326 161.3
R12861 commonsourceibias.n324 commonsourceibias.n206 161.3
R12862 commonsourceibias.n323 commonsourceibias.n322 161.3
R12863 commonsourceibias.n321 commonsourceibias.n207 161.3
R12864 commonsourceibias.n320 commonsourceibias.n319 161.3
R12865 commonsourceibias.n317 commonsourceibias.n208 161.3
R12866 commonsourceibias.n315 commonsourceibias.n314 161.3
R12867 commonsourceibias.n400 commonsourceibias.n340 161.3
R12868 commonsourceibias.n399 commonsourceibias.n398 161.3
R12869 commonsourceibias.n397 commonsourceibias.n396 161.3
R12870 commonsourceibias.n395 commonsourceibias.n342 161.3
R12871 commonsourceibias.n393 commonsourceibias.n392 161.3
R12872 commonsourceibias.n391 commonsourceibias.n343 161.3
R12873 commonsourceibias.n390 commonsourceibias.n389 161.3
R12874 commonsourceibias.n387 commonsourceibias.n344 161.3
R12875 commonsourceibias.n386 commonsourceibias.n385 161.3
R12876 commonsourceibias.n384 commonsourceibias.n345 161.3
R12877 commonsourceibias.n383 commonsourceibias.n382 161.3
R12878 commonsourceibias.n380 commonsourceibias.n346 161.3
R12879 commonsourceibias.n378 commonsourceibias.n377 161.3
R12880 commonsourceibias.n376 commonsourceibias.n347 161.3
R12881 commonsourceibias.n375 commonsourceibias.n374 161.3
R12882 commonsourceibias.n372 commonsourceibias.n348 161.3
R12883 commonsourceibias.n371 commonsourceibias.n370 161.3
R12884 commonsourceibias.n369 commonsourceibias.n368 161.3
R12885 commonsourceibias.n367 commonsourceibias.n350 161.3
R12886 commonsourceibias.n366 commonsourceibias.n365 161.3
R12887 commonsourceibias.n364 commonsourceibias.n363 161.3
R12888 commonsourceibias.n362 commonsourceibias.n352 161.3
R12889 commonsourceibias.n361 commonsourceibias.n360 161.3
R12890 commonsourceibias.n359 commonsourceibias.n358 161.3
R12891 commonsourceibias.n357 commonsourceibias.n354 161.3
R12892 commonsourceibias.n80 commonsourceibias.n78 81.5057
R12893 commonsourceibias.n240 commonsourceibias.n238 81.5057
R12894 commonsourceibias.n80 commonsourceibias.n79 80.9324
R12895 commonsourceibias.n82 commonsourceibias.n81 80.9324
R12896 commonsourceibias.n77 commonsourceibias.n76 80.9324
R12897 commonsourceibias.n75 commonsourceibias.n74 80.9324
R12898 commonsourceibias.n73 commonsourceibias.n72 80.9324
R12899 commonsourceibias.n307 commonsourceibias.n306 80.9324
R12900 commonsourceibias.n309 commonsourceibias.n308 80.9324
R12901 commonsourceibias.n311 commonsourceibias.n310 80.9324
R12902 commonsourceibias.n242 commonsourceibias.n241 80.9324
R12903 commonsourceibias.n240 commonsourceibias.n239 80.9324
R12904 commonsourceibias.n71 commonsourceibias.n70 80.6037
R12905 commonsourceibias.n137 commonsourceibias.n136 80.6037
R12906 commonsourceibias.n200 commonsourceibias.n199 80.6037
R12907 commonsourceibias.n305 commonsourceibias.n304 80.6037
R12908 commonsourceibias.n339 commonsourceibias.n338 80.6037
R12909 commonsourceibias.n402 commonsourceibias.n401 80.6037
R12910 commonsourceibias.n65 commonsourceibias.n64 56.5617
R12911 commonsourceibias.n51 commonsourceibias.n50 56.5617
R12912 commonsourceibias.n42 commonsourceibias.n41 56.5617
R12913 commonsourceibias.n28 commonsourceibias.n27 56.5617
R12914 commonsourceibias.n131 commonsourceibias.n130 56.5617
R12915 commonsourceibias.n117 commonsourceibias.n116 56.5617
R12916 commonsourceibias.n108 commonsourceibias.n107 56.5617
R12917 commonsourceibias.n94 commonsourceibias.n93 56.5617
R12918 commonsourceibias.n157 commonsourceibias.n156 56.5617
R12919 commonsourceibias.n171 commonsourceibias.n170 56.5617
R12920 commonsourceibias.n180 commonsourceibias.n179 56.5617
R12921 commonsourceibias.n194 commonsourceibias.n193 56.5617
R12922 commonsourceibias.n261 commonsourceibias.n260 56.5617
R12923 commonsourceibias.n275 commonsourceibias.n274 56.5617
R12924 commonsourceibias.n285 commonsourceibias.n283 56.5617
R12925 commonsourceibias.n299 commonsourceibias.n298 56.5617
R12926 commonsourceibias.n333 commonsourceibias.n332 56.5617
R12927 commonsourceibias.n319 commonsourceibias.n317 56.5617
R12928 commonsourceibias.n220 commonsourceibias.n219 56.5617
R12929 commonsourceibias.n234 commonsourceibias.n233 56.5617
R12930 commonsourceibias.n358 commonsourceibias.n357 56.5617
R12931 commonsourceibias.n372 commonsourceibias.n371 56.5617
R12932 commonsourceibias.n382 commonsourceibias.n380 56.5617
R12933 commonsourceibias.n396 commonsourceibias.n395 56.5617
R12934 commonsourceibias.n56 commonsourceibias.n55 56.0773
R12935 commonsourceibias.n37 commonsourceibias.n36 56.0773
R12936 commonsourceibias.n122 commonsourceibias.n121 56.0773
R12937 commonsourceibias.n103 commonsourceibias.n102 56.0773
R12938 commonsourceibias.n166 commonsourceibias.n165 56.0773
R12939 commonsourceibias.n185 commonsourceibias.n184 56.0773
R12940 commonsourceibias.n270 commonsourceibias.n269 56.0773
R12941 commonsourceibias.n290 commonsourceibias.n289 56.0773
R12942 commonsourceibias.n324 commonsourceibias.n323 56.0773
R12943 commonsourceibias.n229 commonsourceibias.n228 56.0773
R12944 commonsourceibias.n367 commonsourceibias.n366 56.0773
R12945 commonsourceibias.n387 commonsourceibias.n386 56.0773
R12946 commonsourceibias.n70 commonsourceibias.n69 46.0096
R12947 commonsourceibias.n136 commonsourceibias.n135 46.0096
R12948 commonsourceibias.n199 commonsourceibias.n198 46.0096
R12949 commonsourceibias.n304 commonsourceibias.n303 46.0096
R12950 commonsourceibias.n338 commonsourceibias.n337 46.0096
R12951 commonsourceibias.n401 commonsourceibias.n400 46.0096
R12952 commonsourceibias.n58 commonsourceibias.n12 41.5458
R12953 commonsourceibias.n33 commonsourceibias.n32 41.5458
R12954 commonsourceibias.n124 commonsourceibias.n3 41.5458
R12955 commonsourceibias.n99 commonsourceibias.n98 41.5458
R12956 commonsourceibias.n162 commonsourceibias.n161 41.5458
R12957 commonsourceibias.n187 commonsourceibias.n141 41.5458
R12958 commonsourceibias.n266 commonsourceibias.n265 41.5458
R12959 commonsourceibias.n292 commonsourceibias.n246 41.5458
R12960 commonsourceibias.n326 commonsourceibias.n205 41.5458
R12961 commonsourceibias.n225 commonsourceibias.n224 41.5458
R12962 commonsourceibias.n363 commonsourceibias.n362 41.5458
R12963 commonsourceibias.n389 commonsourceibias.n343 41.5458
R12964 commonsourceibias.n48 commonsourceibias.n17 40.577
R12965 commonsourceibias.n44 commonsourceibias.n17 40.577
R12966 commonsourceibias.n114 commonsourceibias.n8 40.577
R12967 commonsourceibias.n110 commonsourceibias.n8 40.577
R12968 commonsourceibias.n173 commonsourceibias.n146 40.577
R12969 commonsourceibias.n177 commonsourceibias.n146 40.577
R12970 commonsourceibias.n277 commonsourceibias.n250 40.577
R12971 commonsourceibias.n281 commonsourceibias.n250 40.577
R12972 commonsourceibias.n315 commonsourceibias.n209 40.577
R12973 commonsourceibias.n236 commonsourceibias.n209 40.577
R12974 commonsourceibias.n374 commonsourceibias.n347 40.577
R12975 commonsourceibias.n378 commonsourceibias.n347 40.577
R12976 commonsourceibias.n62 commonsourceibias.n12 39.6083
R12977 commonsourceibias.n32 commonsourceibias.n31 39.6083
R12978 commonsourceibias.n128 commonsourceibias.n3 39.6083
R12979 commonsourceibias.n98 commonsourceibias.n97 39.6083
R12980 commonsourceibias.n161 commonsourceibias.n160 39.6083
R12981 commonsourceibias.n191 commonsourceibias.n141 39.6083
R12982 commonsourceibias.n265 commonsourceibias.n264 39.6083
R12983 commonsourceibias.n296 commonsourceibias.n246 39.6083
R12984 commonsourceibias.n330 commonsourceibias.n205 39.6083
R12985 commonsourceibias.n224 commonsourceibias.n223 39.6083
R12986 commonsourceibias.n362 commonsourceibias.n361 39.6083
R12987 commonsourceibias.n393 commonsourceibias.n343 39.6083
R12988 commonsourceibias.n26 commonsourceibias.n25 33.0515
R12989 commonsourceibias.n92 commonsourceibias.n91 33.0515
R12990 commonsourceibias.n155 commonsourceibias.n154 33.0515
R12991 commonsourceibias.n259 commonsourceibias.n258 33.0515
R12992 commonsourceibias.n218 commonsourceibias.n217 33.0515
R12993 commonsourceibias.n356 commonsourceibias.n355 33.0515
R12994 commonsourceibias.n25 commonsourceibias.n24 28.5514
R12995 commonsourceibias.n91 commonsourceibias.n90 28.5514
R12996 commonsourceibias.n154 commonsourceibias.n153 28.5514
R12997 commonsourceibias.n258 commonsourceibias.n257 28.5514
R12998 commonsourceibias.n217 commonsourceibias.n216 28.5514
R12999 commonsourceibias.n355 commonsourceibias.n354 28.5514
R13000 commonsourceibias.n69 commonsourceibias.n68 26.0455
R13001 commonsourceibias.n135 commonsourceibias.n134 26.0455
R13002 commonsourceibias.n198 commonsourceibias.n197 26.0455
R13003 commonsourceibias.n303 commonsourceibias.n302 26.0455
R13004 commonsourceibias.n337 commonsourceibias.n336 26.0455
R13005 commonsourceibias.n400 commonsourceibias.n399 26.0455
R13006 commonsourceibias.n55 commonsourceibias.n14 25.0767
R13007 commonsourceibias.n38 commonsourceibias.n37 25.0767
R13008 commonsourceibias.n121 commonsourceibias.n5 25.0767
R13009 commonsourceibias.n104 commonsourceibias.n103 25.0767
R13010 commonsourceibias.n167 commonsourceibias.n166 25.0767
R13011 commonsourceibias.n184 commonsourceibias.n143 25.0767
R13012 commonsourceibias.n271 commonsourceibias.n270 25.0767
R13013 commonsourceibias.n289 commonsourceibias.n248 25.0767
R13014 commonsourceibias.n323 commonsourceibias.n207 25.0767
R13015 commonsourceibias.n230 commonsourceibias.n229 25.0767
R13016 commonsourceibias.n368 commonsourceibias.n367 25.0767
R13017 commonsourceibias.n386 commonsourceibias.n345 25.0767
R13018 commonsourceibias.n51 commonsourceibias.n16 24.3464
R13019 commonsourceibias.n41 commonsourceibias.n19 24.3464
R13020 commonsourceibias.n117 commonsourceibias.n7 24.3464
R13021 commonsourceibias.n107 commonsourceibias.n85 24.3464
R13022 commonsourceibias.n170 commonsourceibias.n148 24.3464
R13023 commonsourceibias.n180 commonsourceibias.n145 24.3464
R13024 commonsourceibias.n274 commonsourceibias.n252 24.3464
R13025 commonsourceibias.n285 commonsourceibias.n284 24.3464
R13026 commonsourceibias.n319 commonsourceibias.n318 24.3464
R13027 commonsourceibias.n233 commonsourceibias.n211 24.3464
R13028 commonsourceibias.n371 commonsourceibias.n349 24.3464
R13029 commonsourceibias.n382 commonsourceibias.n381 24.3464
R13030 commonsourceibias.n65 commonsourceibias.n10 23.8546
R13031 commonsourceibias.n27 commonsourceibias.n26 23.8546
R13032 commonsourceibias.n131 commonsourceibias.n1 23.8546
R13033 commonsourceibias.n93 commonsourceibias.n92 23.8546
R13034 commonsourceibias.n156 commonsourceibias.n155 23.8546
R13035 commonsourceibias.n194 commonsourceibias.n139 23.8546
R13036 commonsourceibias.n260 commonsourceibias.n259 23.8546
R13037 commonsourceibias.n299 commonsourceibias.n244 23.8546
R13038 commonsourceibias.n333 commonsourceibias.n203 23.8546
R13039 commonsourceibias.n219 commonsourceibias.n218 23.8546
R13040 commonsourceibias.n357 commonsourceibias.n356 23.8546
R13041 commonsourceibias.n396 commonsourceibias.n341 23.8546
R13042 commonsourceibias.n64 commonsourceibias.n63 16.9689
R13043 commonsourceibias.n28 commonsourceibias.n23 16.9689
R13044 commonsourceibias.n130 commonsourceibias.n129 16.9689
R13045 commonsourceibias.n94 commonsourceibias.n89 16.9689
R13046 commonsourceibias.n157 commonsourceibias.n152 16.9689
R13047 commonsourceibias.n193 commonsourceibias.n192 16.9689
R13048 commonsourceibias.n261 commonsourceibias.n256 16.9689
R13049 commonsourceibias.n298 commonsourceibias.n297 16.9689
R13050 commonsourceibias.n332 commonsourceibias.n331 16.9689
R13051 commonsourceibias.n220 commonsourceibias.n215 16.9689
R13052 commonsourceibias.n358 commonsourceibias.n353 16.9689
R13053 commonsourceibias.n395 commonsourceibias.n394 16.9689
R13054 commonsourceibias.n50 commonsourceibias.n49 16.477
R13055 commonsourceibias.n43 commonsourceibias.n42 16.477
R13056 commonsourceibias.n116 commonsourceibias.n115 16.477
R13057 commonsourceibias.n109 commonsourceibias.n108 16.477
R13058 commonsourceibias.n172 commonsourceibias.n171 16.477
R13059 commonsourceibias.n179 commonsourceibias.n178 16.477
R13060 commonsourceibias.n276 commonsourceibias.n275 16.477
R13061 commonsourceibias.n283 commonsourceibias.n282 16.477
R13062 commonsourceibias.n317 commonsourceibias.n316 16.477
R13063 commonsourceibias.n235 commonsourceibias.n234 16.477
R13064 commonsourceibias.n373 commonsourceibias.n372 16.477
R13065 commonsourceibias.n380 commonsourceibias.n379 16.477
R13066 commonsourceibias.n57 commonsourceibias.n56 15.9852
R13067 commonsourceibias.n36 commonsourceibias.n21 15.9852
R13068 commonsourceibias.n123 commonsourceibias.n122 15.9852
R13069 commonsourceibias.n102 commonsourceibias.n87 15.9852
R13070 commonsourceibias.n165 commonsourceibias.n150 15.9852
R13071 commonsourceibias.n186 commonsourceibias.n185 15.9852
R13072 commonsourceibias.n269 commonsourceibias.n254 15.9852
R13073 commonsourceibias.n291 commonsourceibias.n290 15.9852
R13074 commonsourceibias.n325 commonsourceibias.n324 15.9852
R13075 commonsourceibias.n228 commonsourceibias.n213 15.9852
R13076 commonsourceibias.n366 commonsourceibias.n351 15.9852
R13077 commonsourceibias.n388 commonsourceibias.n387 15.9852
R13078 commonsourceibias.n73 commonsourceibias.n71 13.2057
R13079 commonsourceibias.n307 commonsourceibias.n305 13.2057
R13080 commonsourceibias.n404 commonsourceibias.n201 11.9876
R13081 commonsourceibias.n404 commonsourceibias.n403 10.3347
R13082 commonsourceibias.n112 commonsourceibias.n83 9.50363
R13083 commonsourceibias.n313 commonsourceibias.n312 9.50363
R13084 commonsourceibias.n201 commonsourceibias.n137 8.732
R13085 commonsourceibias.n403 commonsourceibias.n339 8.732
R13086 commonsourceibias.n58 commonsourceibias.n57 8.60764
R13087 commonsourceibias.n33 commonsourceibias.n21 8.60764
R13088 commonsourceibias.n124 commonsourceibias.n123 8.60764
R13089 commonsourceibias.n99 commonsourceibias.n87 8.60764
R13090 commonsourceibias.n162 commonsourceibias.n150 8.60764
R13091 commonsourceibias.n187 commonsourceibias.n186 8.60764
R13092 commonsourceibias.n266 commonsourceibias.n254 8.60764
R13093 commonsourceibias.n292 commonsourceibias.n291 8.60764
R13094 commonsourceibias.n326 commonsourceibias.n325 8.60764
R13095 commonsourceibias.n225 commonsourceibias.n213 8.60764
R13096 commonsourceibias.n363 commonsourceibias.n351 8.60764
R13097 commonsourceibias.n389 commonsourceibias.n388 8.60764
R13098 commonsourceibias.n49 commonsourceibias.n48 8.11581
R13099 commonsourceibias.n44 commonsourceibias.n43 8.11581
R13100 commonsourceibias.n115 commonsourceibias.n114 8.11581
R13101 commonsourceibias.n110 commonsourceibias.n109 8.11581
R13102 commonsourceibias.n173 commonsourceibias.n172 8.11581
R13103 commonsourceibias.n178 commonsourceibias.n177 8.11581
R13104 commonsourceibias.n277 commonsourceibias.n276 8.11581
R13105 commonsourceibias.n282 commonsourceibias.n281 8.11581
R13106 commonsourceibias.n316 commonsourceibias.n315 8.11581
R13107 commonsourceibias.n236 commonsourceibias.n235 8.11581
R13108 commonsourceibias.n374 commonsourceibias.n373 8.11581
R13109 commonsourceibias.n379 commonsourceibias.n378 8.11581
R13110 commonsourceibias.n63 commonsourceibias.n62 7.62397
R13111 commonsourceibias.n31 commonsourceibias.n23 7.62397
R13112 commonsourceibias.n129 commonsourceibias.n128 7.62397
R13113 commonsourceibias.n97 commonsourceibias.n89 7.62397
R13114 commonsourceibias.n160 commonsourceibias.n152 7.62397
R13115 commonsourceibias.n192 commonsourceibias.n191 7.62397
R13116 commonsourceibias.n264 commonsourceibias.n256 7.62397
R13117 commonsourceibias.n297 commonsourceibias.n296 7.62397
R13118 commonsourceibias.n331 commonsourceibias.n330 7.62397
R13119 commonsourceibias.n223 commonsourceibias.n215 7.62397
R13120 commonsourceibias.n361 commonsourceibias.n353 7.62397
R13121 commonsourceibias.n394 commonsourceibias.n393 7.62397
R13122 commonsourceibias.n201 commonsourceibias.n200 5.00473
R13123 commonsourceibias.n403 commonsourceibias.n402 5.00473
R13124 commonsourceibias commonsourceibias.n404 3.87639
R13125 commonsourceibias.n78 commonsourceibias.t41 2.82907
R13126 commonsourceibias.n78 commonsourceibias.t47 2.82907
R13127 commonsourceibias.n79 commonsourceibias.t35 2.82907
R13128 commonsourceibias.n79 commonsourceibias.t11 2.82907
R13129 commonsourceibias.n81 commonsourceibias.t45 2.82907
R13130 commonsourceibias.n81 commonsourceibias.t27 2.82907
R13131 commonsourceibias.n76 commonsourceibias.t21 2.82907
R13132 commonsourceibias.n76 commonsourceibias.t37 2.82907
R13133 commonsourceibias.n74 commonsourceibias.t25 2.82907
R13134 commonsourceibias.n74 commonsourceibias.t31 2.82907
R13135 commonsourceibias.n72 commonsourceibias.t33 2.82907
R13136 commonsourceibias.n72 commonsourceibias.t15 2.82907
R13137 commonsourceibias.n306 commonsourceibias.t23 2.82907
R13138 commonsourceibias.n306 commonsourceibias.t3 2.82907
R13139 commonsourceibias.n308 commonsourceibias.t1 2.82907
R13140 commonsourceibias.n308 commonsourceibias.t39 2.82907
R13141 commonsourceibias.n310 commonsourceibias.t7 2.82907
R13142 commonsourceibias.n310 commonsourceibias.t29 2.82907
R13143 commonsourceibias.n241 commonsourceibias.t43 2.82907
R13144 commonsourceibias.n241 commonsourceibias.t13 2.82907
R13145 commonsourceibias.n239 commonsourceibias.t19 2.82907
R13146 commonsourceibias.n239 commonsourceibias.t5 2.82907
R13147 commonsourceibias.n238 commonsourceibias.t17 2.82907
R13148 commonsourceibias.n238 commonsourceibias.t9 2.82907
R13149 commonsourceibias.n68 commonsourceibias.n10 0.738255
R13150 commonsourceibias.n134 commonsourceibias.n1 0.738255
R13151 commonsourceibias.n197 commonsourceibias.n139 0.738255
R13152 commonsourceibias.n302 commonsourceibias.n244 0.738255
R13153 commonsourceibias.n336 commonsourceibias.n203 0.738255
R13154 commonsourceibias.n399 commonsourceibias.n341 0.738255
R13155 commonsourceibias.n75 commonsourceibias.n73 0.573776
R13156 commonsourceibias.n77 commonsourceibias.n75 0.573776
R13157 commonsourceibias.n82 commonsourceibias.n80 0.573776
R13158 commonsourceibias.n242 commonsourceibias.n240 0.573776
R13159 commonsourceibias.n311 commonsourceibias.n309 0.573776
R13160 commonsourceibias.n309 commonsourceibias.n307 0.573776
R13161 commonsourceibias.n83 commonsourceibias.n77 0.287138
R13162 commonsourceibias.n83 commonsourceibias.n82 0.287138
R13163 commonsourceibias.n312 commonsourceibias.n242 0.287138
R13164 commonsourceibias.n312 commonsourceibias.n311 0.287138
R13165 commonsourceibias.n71 commonsourceibias.n9 0.285035
R13166 commonsourceibias.n137 commonsourceibias.n0 0.285035
R13167 commonsourceibias.n200 commonsourceibias.n138 0.285035
R13168 commonsourceibias.n305 commonsourceibias.n243 0.285035
R13169 commonsourceibias.n339 commonsourceibias.n202 0.285035
R13170 commonsourceibias.n402 commonsourceibias.n340 0.285035
R13171 commonsourceibias.n16 commonsourceibias.n14 0.246418
R13172 commonsourceibias.n38 commonsourceibias.n19 0.246418
R13173 commonsourceibias.n7 commonsourceibias.n5 0.246418
R13174 commonsourceibias.n104 commonsourceibias.n85 0.246418
R13175 commonsourceibias.n167 commonsourceibias.n148 0.246418
R13176 commonsourceibias.n145 commonsourceibias.n143 0.246418
R13177 commonsourceibias.n271 commonsourceibias.n252 0.246418
R13178 commonsourceibias.n284 commonsourceibias.n248 0.246418
R13179 commonsourceibias.n318 commonsourceibias.n207 0.246418
R13180 commonsourceibias.n230 commonsourceibias.n211 0.246418
R13181 commonsourceibias.n368 commonsourceibias.n349 0.246418
R13182 commonsourceibias.n381 commonsourceibias.n345 0.246418
R13183 commonsourceibias.n67 commonsourceibias.n9 0.189894
R13184 commonsourceibias.n67 commonsourceibias.n66 0.189894
R13185 commonsourceibias.n66 commonsourceibias.n11 0.189894
R13186 commonsourceibias.n61 commonsourceibias.n11 0.189894
R13187 commonsourceibias.n61 commonsourceibias.n60 0.189894
R13188 commonsourceibias.n60 commonsourceibias.n59 0.189894
R13189 commonsourceibias.n59 commonsourceibias.n13 0.189894
R13190 commonsourceibias.n54 commonsourceibias.n13 0.189894
R13191 commonsourceibias.n54 commonsourceibias.n53 0.189894
R13192 commonsourceibias.n53 commonsourceibias.n52 0.189894
R13193 commonsourceibias.n52 commonsourceibias.n15 0.189894
R13194 commonsourceibias.n47 commonsourceibias.n15 0.189894
R13195 commonsourceibias.n47 commonsourceibias.n46 0.189894
R13196 commonsourceibias.n46 commonsourceibias.n45 0.189894
R13197 commonsourceibias.n45 commonsourceibias.n18 0.189894
R13198 commonsourceibias.n40 commonsourceibias.n18 0.189894
R13199 commonsourceibias.n40 commonsourceibias.n39 0.189894
R13200 commonsourceibias.n39 commonsourceibias.n20 0.189894
R13201 commonsourceibias.n35 commonsourceibias.n20 0.189894
R13202 commonsourceibias.n35 commonsourceibias.n34 0.189894
R13203 commonsourceibias.n34 commonsourceibias.n22 0.189894
R13204 commonsourceibias.n30 commonsourceibias.n22 0.189894
R13205 commonsourceibias.n30 commonsourceibias.n29 0.189894
R13206 commonsourceibias.n29 commonsourceibias.n24 0.189894
R13207 commonsourceibias.n111 commonsourceibias.n84 0.189894
R13208 commonsourceibias.n106 commonsourceibias.n84 0.189894
R13209 commonsourceibias.n106 commonsourceibias.n105 0.189894
R13210 commonsourceibias.n105 commonsourceibias.n86 0.189894
R13211 commonsourceibias.n101 commonsourceibias.n86 0.189894
R13212 commonsourceibias.n101 commonsourceibias.n100 0.189894
R13213 commonsourceibias.n100 commonsourceibias.n88 0.189894
R13214 commonsourceibias.n96 commonsourceibias.n88 0.189894
R13215 commonsourceibias.n96 commonsourceibias.n95 0.189894
R13216 commonsourceibias.n95 commonsourceibias.n90 0.189894
R13217 commonsourceibias.n133 commonsourceibias.n0 0.189894
R13218 commonsourceibias.n133 commonsourceibias.n132 0.189894
R13219 commonsourceibias.n132 commonsourceibias.n2 0.189894
R13220 commonsourceibias.n127 commonsourceibias.n2 0.189894
R13221 commonsourceibias.n127 commonsourceibias.n126 0.189894
R13222 commonsourceibias.n126 commonsourceibias.n125 0.189894
R13223 commonsourceibias.n125 commonsourceibias.n4 0.189894
R13224 commonsourceibias.n120 commonsourceibias.n4 0.189894
R13225 commonsourceibias.n120 commonsourceibias.n119 0.189894
R13226 commonsourceibias.n119 commonsourceibias.n118 0.189894
R13227 commonsourceibias.n118 commonsourceibias.n6 0.189894
R13228 commonsourceibias.n113 commonsourceibias.n6 0.189894
R13229 commonsourceibias.n196 commonsourceibias.n138 0.189894
R13230 commonsourceibias.n196 commonsourceibias.n195 0.189894
R13231 commonsourceibias.n195 commonsourceibias.n140 0.189894
R13232 commonsourceibias.n190 commonsourceibias.n140 0.189894
R13233 commonsourceibias.n190 commonsourceibias.n189 0.189894
R13234 commonsourceibias.n189 commonsourceibias.n188 0.189894
R13235 commonsourceibias.n188 commonsourceibias.n142 0.189894
R13236 commonsourceibias.n183 commonsourceibias.n142 0.189894
R13237 commonsourceibias.n183 commonsourceibias.n182 0.189894
R13238 commonsourceibias.n182 commonsourceibias.n181 0.189894
R13239 commonsourceibias.n181 commonsourceibias.n144 0.189894
R13240 commonsourceibias.n176 commonsourceibias.n144 0.189894
R13241 commonsourceibias.n176 commonsourceibias.n175 0.189894
R13242 commonsourceibias.n175 commonsourceibias.n174 0.189894
R13243 commonsourceibias.n174 commonsourceibias.n147 0.189894
R13244 commonsourceibias.n169 commonsourceibias.n147 0.189894
R13245 commonsourceibias.n169 commonsourceibias.n168 0.189894
R13246 commonsourceibias.n168 commonsourceibias.n149 0.189894
R13247 commonsourceibias.n164 commonsourceibias.n149 0.189894
R13248 commonsourceibias.n164 commonsourceibias.n163 0.189894
R13249 commonsourceibias.n163 commonsourceibias.n151 0.189894
R13250 commonsourceibias.n159 commonsourceibias.n151 0.189894
R13251 commonsourceibias.n159 commonsourceibias.n158 0.189894
R13252 commonsourceibias.n158 commonsourceibias.n153 0.189894
R13253 commonsourceibias.n262 commonsourceibias.n257 0.189894
R13254 commonsourceibias.n263 commonsourceibias.n262 0.189894
R13255 commonsourceibias.n263 commonsourceibias.n255 0.189894
R13256 commonsourceibias.n267 commonsourceibias.n255 0.189894
R13257 commonsourceibias.n268 commonsourceibias.n267 0.189894
R13258 commonsourceibias.n268 commonsourceibias.n253 0.189894
R13259 commonsourceibias.n272 commonsourceibias.n253 0.189894
R13260 commonsourceibias.n273 commonsourceibias.n272 0.189894
R13261 commonsourceibias.n273 commonsourceibias.n251 0.189894
R13262 commonsourceibias.n278 commonsourceibias.n251 0.189894
R13263 commonsourceibias.n279 commonsourceibias.n278 0.189894
R13264 commonsourceibias.n280 commonsourceibias.n279 0.189894
R13265 commonsourceibias.n280 commonsourceibias.n249 0.189894
R13266 commonsourceibias.n286 commonsourceibias.n249 0.189894
R13267 commonsourceibias.n287 commonsourceibias.n286 0.189894
R13268 commonsourceibias.n288 commonsourceibias.n287 0.189894
R13269 commonsourceibias.n288 commonsourceibias.n247 0.189894
R13270 commonsourceibias.n293 commonsourceibias.n247 0.189894
R13271 commonsourceibias.n294 commonsourceibias.n293 0.189894
R13272 commonsourceibias.n295 commonsourceibias.n294 0.189894
R13273 commonsourceibias.n295 commonsourceibias.n245 0.189894
R13274 commonsourceibias.n300 commonsourceibias.n245 0.189894
R13275 commonsourceibias.n301 commonsourceibias.n300 0.189894
R13276 commonsourceibias.n301 commonsourceibias.n243 0.189894
R13277 commonsourceibias.n221 commonsourceibias.n216 0.189894
R13278 commonsourceibias.n222 commonsourceibias.n221 0.189894
R13279 commonsourceibias.n222 commonsourceibias.n214 0.189894
R13280 commonsourceibias.n226 commonsourceibias.n214 0.189894
R13281 commonsourceibias.n227 commonsourceibias.n226 0.189894
R13282 commonsourceibias.n227 commonsourceibias.n212 0.189894
R13283 commonsourceibias.n231 commonsourceibias.n212 0.189894
R13284 commonsourceibias.n232 commonsourceibias.n231 0.189894
R13285 commonsourceibias.n232 commonsourceibias.n210 0.189894
R13286 commonsourceibias.n237 commonsourceibias.n210 0.189894
R13287 commonsourceibias.n314 commonsourceibias.n208 0.189894
R13288 commonsourceibias.n320 commonsourceibias.n208 0.189894
R13289 commonsourceibias.n321 commonsourceibias.n320 0.189894
R13290 commonsourceibias.n322 commonsourceibias.n321 0.189894
R13291 commonsourceibias.n322 commonsourceibias.n206 0.189894
R13292 commonsourceibias.n327 commonsourceibias.n206 0.189894
R13293 commonsourceibias.n328 commonsourceibias.n327 0.189894
R13294 commonsourceibias.n329 commonsourceibias.n328 0.189894
R13295 commonsourceibias.n329 commonsourceibias.n204 0.189894
R13296 commonsourceibias.n334 commonsourceibias.n204 0.189894
R13297 commonsourceibias.n335 commonsourceibias.n334 0.189894
R13298 commonsourceibias.n335 commonsourceibias.n202 0.189894
R13299 commonsourceibias.n359 commonsourceibias.n354 0.189894
R13300 commonsourceibias.n360 commonsourceibias.n359 0.189894
R13301 commonsourceibias.n360 commonsourceibias.n352 0.189894
R13302 commonsourceibias.n364 commonsourceibias.n352 0.189894
R13303 commonsourceibias.n365 commonsourceibias.n364 0.189894
R13304 commonsourceibias.n365 commonsourceibias.n350 0.189894
R13305 commonsourceibias.n369 commonsourceibias.n350 0.189894
R13306 commonsourceibias.n370 commonsourceibias.n369 0.189894
R13307 commonsourceibias.n370 commonsourceibias.n348 0.189894
R13308 commonsourceibias.n375 commonsourceibias.n348 0.189894
R13309 commonsourceibias.n376 commonsourceibias.n375 0.189894
R13310 commonsourceibias.n377 commonsourceibias.n376 0.189894
R13311 commonsourceibias.n377 commonsourceibias.n346 0.189894
R13312 commonsourceibias.n383 commonsourceibias.n346 0.189894
R13313 commonsourceibias.n384 commonsourceibias.n383 0.189894
R13314 commonsourceibias.n385 commonsourceibias.n384 0.189894
R13315 commonsourceibias.n385 commonsourceibias.n344 0.189894
R13316 commonsourceibias.n390 commonsourceibias.n344 0.189894
R13317 commonsourceibias.n391 commonsourceibias.n390 0.189894
R13318 commonsourceibias.n392 commonsourceibias.n391 0.189894
R13319 commonsourceibias.n392 commonsourceibias.n342 0.189894
R13320 commonsourceibias.n397 commonsourceibias.n342 0.189894
R13321 commonsourceibias.n398 commonsourceibias.n397 0.189894
R13322 commonsourceibias.n398 commonsourceibias.n340 0.189894
R13323 commonsourceibias.n112 commonsourceibias.n111 0.170955
R13324 commonsourceibias.n113 commonsourceibias.n112 0.170955
R13325 commonsourceibias.n313 commonsourceibias.n237 0.170955
R13326 commonsourceibias.n314 commonsourceibias.n313 0.170955
R13327 CSoutput.n19 CSoutput.t165 184.661
R13328 CSoutput.n78 CSoutput.n77 165.8
R13329 CSoutput.n76 CSoutput.n0 165.8
R13330 CSoutput.n75 CSoutput.n74 165.8
R13331 CSoutput.n73 CSoutput.n72 165.8
R13332 CSoutput.n71 CSoutput.n2 165.8
R13333 CSoutput.n69 CSoutput.n68 165.8
R13334 CSoutput.n67 CSoutput.n3 165.8
R13335 CSoutput.n66 CSoutput.n65 165.8
R13336 CSoutput.n63 CSoutput.n4 165.8
R13337 CSoutput.n61 CSoutput.n60 165.8
R13338 CSoutput.n59 CSoutput.n5 165.8
R13339 CSoutput.n58 CSoutput.n57 165.8
R13340 CSoutput.n55 CSoutput.n6 165.8
R13341 CSoutput.n54 CSoutput.n53 165.8
R13342 CSoutput.n52 CSoutput.n51 165.8
R13343 CSoutput.n50 CSoutput.n8 165.8
R13344 CSoutput.n48 CSoutput.n47 165.8
R13345 CSoutput.n46 CSoutput.n9 165.8
R13346 CSoutput.n45 CSoutput.n44 165.8
R13347 CSoutput.n42 CSoutput.n10 165.8
R13348 CSoutput.n41 CSoutput.n40 165.8
R13349 CSoutput.n39 CSoutput.n38 165.8
R13350 CSoutput.n37 CSoutput.n12 165.8
R13351 CSoutput.n35 CSoutput.n34 165.8
R13352 CSoutput.n33 CSoutput.n13 165.8
R13353 CSoutput.n32 CSoutput.n31 165.8
R13354 CSoutput.n29 CSoutput.n14 165.8
R13355 CSoutput.n28 CSoutput.n27 165.8
R13356 CSoutput.n26 CSoutput.n25 165.8
R13357 CSoutput.n24 CSoutput.n16 165.8
R13358 CSoutput.n22 CSoutput.n21 165.8
R13359 CSoutput.n20 CSoutput.n17 165.8
R13360 CSoutput.n77 CSoutput.t144 162.194
R13361 CSoutput.n18 CSoutput.t145 120.501
R13362 CSoutput.n23 CSoutput.t155 120.501
R13363 CSoutput.n15 CSoutput.t151 120.501
R13364 CSoutput.n30 CSoutput.t147 120.501
R13365 CSoutput.n36 CSoutput.t158 120.501
R13366 CSoutput.n11 CSoutput.t160 120.501
R13367 CSoutput.n43 CSoutput.t149 120.501
R13368 CSoutput.n49 CSoutput.t161 120.501
R13369 CSoutput.n7 CSoutput.t162 120.501
R13370 CSoutput.n56 CSoutput.t156 120.501
R13371 CSoutput.n62 CSoutput.t148 120.501
R13372 CSoutput.n64 CSoutput.t164 120.501
R13373 CSoutput.n70 CSoutput.t159 120.501
R13374 CSoutput.n1 CSoutput.t154 120.501
R13375 CSoutput.n310 CSoutput.n308 103.469
R13376 CSoutput.n294 CSoutput.n292 103.469
R13377 CSoutput.n279 CSoutput.n277 103.469
R13378 CSoutput.n112 CSoutput.n110 103.469
R13379 CSoutput.n96 CSoutput.n94 103.469
R13380 CSoutput.n81 CSoutput.n79 103.469
R13381 CSoutput.n320 CSoutput.n319 103.111
R13382 CSoutput.n318 CSoutput.n317 103.111
R13383 CSoutput.n316 CSoutput.n315 103.111
R13384 CSoutput.n314 CSoutput.n313 103.111
R13385 CSoutput.n312 CSoutput.n311 103.111
R13386 CSoutput.n310 CSoutput.n309 103.111
R13387 CSoutput.n306 CSoutput.n305 103.111
R13388 CSoutput.n304 CSoutput.n303 103.111
R13389 CSoutput.n302 CSoutput.n301 103.111
R13390 CSoutput.n300 CSoutput.n299 103.111
R13391 CSoutput.n298 CSoutput.n297 103.111
R13392 CSoutput.n296 CSoutput.n295 103.111
R13393 CSoutput.n294 CSoutput.n293 103.111
R13394 CSoutput.n291 CSoutput.n290 103.111
R13395 CSoutput.n289 CSoutput.n288 103.111
R13396 CSoutput.n287 CSoutput.n286 103.111
R13397 CSoutput.n285 CSoutput.n284 103.111
R13398 CSoutput.n283 CSoutput.n282 103.111
R13399 CSoutput.n281 CSoutput.n280 103.111
R13400 CSoutput.n279 CSoutput.n278 103.111
R13401 CSoutput.n112 CSoutput.n111 103.111
R13402 CSoutput.n114 CSoutput.n113 103.111
R13403 CSoutput.n116 CSoutput.n115 103.111
R13404 CSoutput.n118 CSoutput.n117 103.111
R13405 CSoutput.n120 CSoutput.n119 103.111
R13406 CSoutput.n122 CSoutput.n121 103.111
R13407 CSoutput.n124 CSoutput.n123 103.111
R13408 CSoutput.n96 CSoutput.n95 103.111
R13409 CSoutput.n98 CSoutput.n97 103.111
R13410 CSoutput.n100 CSoutput.n99 103.111
R13411 CSoutput.n102 CSoutput.n101 103.111
R13412 CSoutput.n104 CSoutput.n103 103.111
R13413 CSoutput.n106 CSoutput.n105 103.111
R13414 CSoutput.n108 CSoutput.n107 103.111
R13415 CSoutput.n81 CSoutput.n80 103.111
R13416 CSoutput.n83 CSoutput.n82 103.111
R13417 CSoutput.n85 CSoutput.n84 103.111
R13418 CSoutput.n87 CSoutput.n86 103.111
R13419 CSoutput.n89 CSoutput.n88 103.111
R13420 CSoutput.n91 CSoutput.n90 103.111
R13421 CSoutput.n93 CSoutput.n92 103.111
R13422 CSoutput.n322 CSoutput.n321 103.111
R13423 CSoutput.n338 CSoutput.n336 81.5057
R13424 CSoutput.n327 CSoutput.n325 81.5057
R13425 CSoutput.n362 CSoutput.n360 81.5057
R13426 CSoutput.n351 CSoutput.n349 81.5057
R13427 CSoutput.n346 CSoutput.n345 80.9324
R13428 CSoutput.n344 CSoutput.n343 80.9324
R13429 CSoutput.n342 CSoutput.n341 80.9324
R13430 CSoutput.n340 CSoutput.n339 80.9324
R13431 CSoutput.n338 CSoutput.n337 80.9324
R13432 CSoutput.n335 CSoutput.n334 80.9324
R13433 CSoutput.n333 CSoutput.n332 80.9324
R13434 CSoutput.n331 CSoutput.n330 80.9324
R13435 CSoutput.n329 CSoutput.n328 80.9324
R13436 CSoutput.n327 CSoutput.n326 80.9324
R13437 CSoutput.n362 CSoutput.n361 80.9324
R13438 CSoutput.n364 CSoutput.n363 80.9324
R13439 CSoutput.n366 CSoutput.n365 80.9324
R13440 CSoutput.n368 CSoutput.n367 80.9324
R13441 CSoutput.n370 CSoutput.n369 80.9324
R13442 CSoutput.n351 CSoutput.n350 80.9324
R13443 CSoutput.n353 CSoutput.n352 80.9324
R13444 CSoutput.n355 CSoutput.n354 80.9324
R13445 CSoutput.n357 CSoutput.n356 80.9324
R13446 CSoutput.n359 CSoutput.n358 80.9324
R13447 CSoutput.n25 CSoutput.n24 48.1486
R13448 CSoutput.n69 CSoutput.n3 48.1486
R13449 CSoutput.n38 CSoutput.n37 48.1486
R13450 CSoutput.n42 CSoutput.n41 48.1486
R13451 CSoutput.n51 CSoutput.n50 48.1486
R13452 CSoutput.n55 CSoutput.n54 48.1486
R13453 CSoutput.n22 CSoutput.n17 46.462
R13454 CSoutput.n72 CSoutput.n71 46.462
R13455 CSoutput.n20 CSoutput.n19 44.9055
R13456 CSoutput.n29 CSoutput.n28 43.7635
R13457 CSoutput.n65 CSoutput.n63 43.7635
R13458 CSoutput.n35 CSoutput.n13 41.7396
R13459 CSoutput.n57 CSoutput.n5 41.7396
R13460 CSoutput.n44 CSoutput.n9 37.0171
R13461 CSoutput.n48 CSoutput.n9 37.0171
R13462 CSoutput.n76 CSoutput.n75 34.9932
R13463 CSoutput.n31 CSoutput.n13 32.2947
R13464 CSoutput.n61 CSoutput.n5 32.2947
R13465 CSoutput.n30 CSoutput.n29 29.6014
R13466 CSoutput.n63 CSoutput.n62 29.6014
R13467 CSoutput.n19 CSoutput.n18 28.4085
R13468 CSoutput.n18 CSoutput.n17 25.1176
R13469 CSoutput.n72 CSoutput.n1 25.1176
R13470 CSoutput.n43 CSoutput.n42 22.0922
R13471 CSoutput.n50 CSoutput.n49 22.0922
R13472 CSoutput.n77 CSoutput.n76 21.8586
R13473 CSoutput.n37 CSoutput.n36 18.9681
R13474 CSoutput.n56 CSoutput.n55 18.9681
R13475 CSoutput.n25 CSoutput.n15 17.6292
R13476 CSoutput.n64 CSoutput.n3 17.6292
R13477 CSoutput.n24 CSoutput.n23 15.844
R13478 CSoutput.n70 CSoutput.n69 15.844
R13479 CSoutput.n38 CSoutput.n11 14.5051
R13480 CSoutput.n54 CSoutput.n7 14.5051
R13481 CSoutput.n373 CSoutput.n78 11.6139
R13482 CSoutput.n41 CSoutput.n11 11.3811
R13483 CSoutput.n51 CSoutput.n7 11.3811
R13484 CSoutput.n23 CSoutput.n22 10.0422
R13485 CSoutput.n71 CSoutput.n70 10.0422
R13486 CSoutput.n307 CSoutput.n291 9.25285
R13487 CSoutput.n109 CSoutput.n93 9.25285
R13488 CSoutput.n347 CSoutput.n335 8.97993
R13489 CSoutput.n371 CSoutput.n359 8.97993
R13490 CSoutput.n348 CSoutput.n324 8.72024
R13491 CSoutput.n28 CSoutput.n15 8.25698
R13492 CSoutput.n65 CSoutput.n64 8.25698
R13493 CSoutput.n348 CSoutput.n347 7.89345
R13494 CSoutput.n372 CSoutput.n371 7.89345
R13495 CSoutput.n324 CSoutput.n323 7.12641
R13496 CSoutput.n126 CSoutput.n125 7.12641
R13497 CSoutput.n36 CSoutput.n35 6.91809
R13498 CSoutput.n57 CSoutput.n56 6.91809
R13499 CSoutput.n347 CSoutput.n346 5.25266
R13500 CSoutput.n371 CSoutput.n370 5.25266
R13501 CSoutput.n323 CSoutput.n322 5.1449
R13502 CSoutput.n307 CSoutput.n306 5.1449
R13503 CSoutput.n125 CSoutput.n124 5.1449
R13504 CSoutput.n109 CSoutput.n108 5.1449
R13505 CSoutput.n373 CSoutput.n126 5.1278
R13506 CSoutput.n217 CSoutput.n170 4.5005
R13507 CSoutput.n186 CSoutput.n170 4.5005
R13508 CSoutput.n181 CSoutput.n165 4.5005
R13509 CSoutput.n181 CSoutput.n167 4.5005
R13510 CSoutput.n181 CSoutput.n164 4.5005
R13511 CSoutput.n181 CSoutput.n168 4.5005
R13512 CSoutput.n181 CSoutput.n163 4.5005
R13513 CSoutput.n181 CSoutput.t150 4.5005
R13514 CSoutput.n181 CSoutput.n162 4.5005
R13515 CSoutput.n181 CSoutput.n169 4.5005
R13516 CSoutput.n181 CSoutput.n170 4.5005
R13517 CSoutput.n179 CSoutput.n165 4.5005
R13518 CSoutput.n179 CSoutput.n167 4.5005
R13519 CSoutput.n179 CSoutput.n164 4.5005
R13520 CSoutput.n179 CSoutput.n168 4.5005
R13521 CSoutput.n179 CSoutput.n163 4.5005
R13522 CSoutput.n179 CSoutput.t150 4.5005
R13523 CSoutput.n179 CSoutput.n162 4.5005
R13524 CSoutput.n179 CSoutput.n169 4.5005
R13525 CSoutput.n179 CSoutput.n170 4.5005
R13526 CSoutput.n178 CSoutput.n165 4.5005
R13527 CSoutput.n178 CSoutput.n167 4.5005
R13528 CSoutput.n178 CSoutput.n164 4.5005
R13529 CSoutput.n178 CSoutput.n168 4.5005
R13530 CSoutput.n178 CSoutput.n163 4.5005
R13531 CSoutput.n178 CSoutput.t150 4.5005
R13532 CSoutput.n178 CSoutput.n162 4.5005
R13533 CSoutput.n178 CSoutput.n169 4.5005
R13534 CSoutput.n178 CSoutput.n170 4.5005
R13535 CSoutput.n263 CSoutput.n165 4.5005
R13536 CSoutput.n263 CSoutput.n167 4.5005
R13537 CSoutput.n263 CSoutput.n164 4.5005
R13538 CSoutput.n263 CSoutput.n168 4.5005
R13539 CSoutput.n263 CSoutput.n163 4.5005
R13540 CSoutput.n263 CSoutput.t150 4.5005
R13541 CSoutput.n263 CSoutput.n162 4.5005
R13542 CSoutput.n263 CSoutput.n169 4.5005
R13543 CSoutput.n263 CSoutput.n170 4.5005
R13544 CSoutput.n261 CSoutput.n165 4.5005
R13545 CSoutput.n261 CSoutput.n167 4.5005
R13546 CSoutput.n261 CSoutput.n164 4.5005
R13547 CSoutput.n261 CSoutput.n168 4.5005
R13548 CSoutput.n261 CSoutput.n163 4.5005
R13549 CSoutput.n261 CSoutput.t150 4.5005
R13550 CSoutput.n261 CSoutput.n162 4.5005
R13551 CSoutput.n261 CSoutput.n169 4.5005
R13552 CSoutput.n259 CSoutput.n165 4.5005
R13553 CSoutput.n259 CSoutput.n167 4.5005
R13554 CSoutput.n259 CSoutput.n164 4.5005
R13555 CSoutput.n259 CSoutput.n168 4.5005
R13556 CSoutput.n259 CSoutput.n163 4.5005
R13557 CSoutput.n259 CSoutput.t150 4.5005
R13558 CSoutput.n259 CSoutput.n162 4.5005
R13559 CSoutput.n259 CSoutput.n169 4.5005
R13560 CSoutput.n189 CSoutput.n165 4.5005
R13561 CSoutput.n189 CSoutput.n167 4.5005
R13562 CSoutput.n189 CSoutput.n164 4.5005
R13563 CSoutput.n189 CSoutput.n168 4.5005
R13564 CSoutput.n189 CSoutput.n163 4.5005
R13565 CSoutput.n189 CSoutput.t150 4.5005
R13566 CSoutput.n189 CSoutput.n162 4.5005
R13567 CSoutput.n189 CSoutput.n169 4.5005
R13568 CSoutput.n189 CSoutput.n170 4.5005
R13569 CSoutput.n188 CSoutput.n165 4.5005
R13570 CSoutput.n188 CSoutput.n167 4.5005
R13571 CSoutput.n188 CSoutput.n164 4.5005
R13572 CSoutput.n188 CSoutput.n168 4.5005
R13573 CSoutput.n188 CSoutput.n163 4.5005
R13574 CSoutput.n188 CSoutput.t150 4.5005
R13575 CSoutput.n188 CSoutput.n162 4.5005
R13576 CSoutput.n188 CSoutput.n169 4.5005
R13577 CSoutput.n188 CSoutput.n170 4.5005
R13578 CSoutput.n192 CSoutput.n165 4.5005
R13579 CSoutput.n192 CSoutput.n167 4.5005
R13580 CSoutput.n192 CSoutput.n164 4.5005
R13581 CSoutput.n192 CSoutput.n168 4.5005
R13582 CSoutput.n192 CSoutput.n163 4.5005
R13583 CSoutput.n192 CSoutput.t150 4.5005
R13584 CSoutput.n192 CSoutput.n162 4.5005
R13585 CSoutput.n192 CSoutput.n169 4.5005
R13586 CSoutput.n192 CSoutput.n170 4.5005
R13587 CSoutput.n191 CSoutput.n165 4.5005
R13588 CSoutput.n191 CSoutput.n167 4.5005
R13589 CSoutput.n191 CSoutput.n164 4.5005
R13590 CSoutput.n191 CSoutput.n168 4.5005
R13591 CSoutput.n191 CSoutput.n163 4.5005
R13592 CSoutput.n191 CSoutput.t150 4.5005
R13593 CSoutput.n191 CSoutput.n162 4.5005
R13594 CSoutput.n191 CSoutput.n169 4.5005
R13595 CSoutput.n191 CSoutput.n170 4.5005
R13596 CSoutput.n174 CSoutput.n165 4.5005
R13597 CSoutput.n174 CSoutput.n167 4.5005
R13598 CSoutput.n174 CSoutput.n164 4.5005
R13599 CSoutput.n174 CSoutput.n168 4.5005
R13600 CSoutput.n174 CSoutput.n163 4.5005
R13601 CSoutput.n174 CSoutput.t150 4.5005
R13602 CSoutput.n174 CSoutput.n162 4.5005
R13603 CSoutput.n174 CSoutput.n169 4.5005
R13604 CSoutput.n174 CSoutput.n170 4.5005
R13605 CSoutput.n266 CSoutput.n165 4.5005
R13606 CSoutput.n266 CSoutput.n167 4.5005
R13607 CSoutput.n266 CSoutput.n164 4.5005
R13608 CSoutput.n266 CSoutput.n168 4.5005
R13609 CSoutput.n266 CSoutput.n163 4.5005
R13610 CSoutput.n266 CSoutput.t150 4.5005
R13611 CSoutput.n266 CSoutput.n162 4.5005
R13612 CSoutput.n266 CSoutput.n169 4.5005
R13613 CSoutput.n266 CSoutput.n170 4.5005
R13614 CSoutput.n253 CSoutput.n224 4.5005
R13615 CSoutput.n253 CSoutput.n230 4.5005
R13616 CSoutput.n211 CSoutput.n200 4.5005
R13617 CSoutput.n211 CSoutput.n202 4.5005
R13618 CSoutput.n211 CSoutput.n199 4.5005
R13619 CSoutput.n211 CSoutput.n203 4.5005
R13620 CSoutput.n211 CSoutput.n198 4.5005
R13621 CSoutput.n211 CSoutput.t146 4.5005
R13622 CSoutput.n211 CSoutput.n197 4.5005
R13623 CSoutput.n211 CSoutput.n204 4.5005
R13624 CSoutput.n253 CSoutput.n211 4.5005
R13625 CSoutput.n232 CSoutput.n200 4.5005
R13626 CSoutput.n232 CSoutput.n202 4.5005
R13627 CSoutput.n232 CSoutput.n199 4.5005
R13628 CSoutput.n232 CSoutput.n203 4.5005
R13629 CSoutput.n232 CSoutput.n198 4.5005
R13630 CSoutput.n232 CSoutput.t146 4.5005
R13631 CSoutput.n232 CSoutput.n197 4.5005
R13632 CSoutput.n232 CSoutput.n204 4.5005
R13633 CSoutput.n253 CSoutput.n232 4.5005
R13634 CSoutput.n210 CSoutput.n200 4.5005
R13635 CSoutput.n210 CSoutput.n202 4.5005
R13636 CSoutput.n210 CSoutput.n199 4.5005
R13637 CSoutput.n210 CSoutput.n203 4.5005
R13638 CSoutput.n210 CSoutput.n198 4.5005
R13639 CSoutput.n210 CSoutput.t146 4.5005
R13640 CSoutput.n210 CSoutput.n197 4.5005
R13641 CSoutput.n210 CSoutput.n204 4.5005
R13642 CSoutput.n253 CSoutput.n210 4.5005
R13643 CSoutput.n234 CSoutput.n200 4.5005
R13644 CSoutput.n234 CSoutput.n202 4.5005
R13645 CSoutput.n234 CSoutput.n199 4.5005
R13646 CSoutput.n234 CSoutput.n203 4.5005
R13647 CSoutput.n234 CSoutput.n198 4.5005
R13648 CSoutput.n234 CSoutput.t146 4.5005
R13649 CSoutput.n234 CSoutput.n197 4.5005
R13650 CSoutput.n234 CSoutput.n204 4.5005
R13651 CSoutput.n253 CSoutput.n234 4.5005
R13652 CSoutput.n200 CSoutput.n195 4.5005
R13653 CSoutput.n202 CSoutput.n195 4.5005
R13654 CSoutput.n199 CSoutput.n195 4.5005
R13655 CSoutput.n203 CSoutput.n195 4.5005
R13656 CSoutput.n198 CSoutput.n195 4.5005
R13657 CSoutput.t146 CSoutput.n195 4.5005
R13658 CSoutput.n197 CSoutput.n195 4.5005
R13659 CSoutput.n204 CSoutput.n195 4.5005
R13660 CSoutput.n256 CSoutput.n200 4.5005
R13661 CSoutput.n256 CSoutput.n202 4.5005
R13662 CSoutput.n256 CSoutput.n199 4.5005
R13663 CSoutput.n256 CSoutput.n203 4.5005
R13664 CSoutput.n256 CSoutput.n198 4.5005
R13665 CSoutput.n256 CSoutput.t146 4.5005
R13666 CSoutput.n256 CSoutput.n197 4.5005
R13667 CSoutput.n256 CSoutput.n204 4.5005
R13668 CSoutput.n254 CSoutput.n200 4.5005
R13669 CSoutput.n254 CSoutput.n202 4.5005
R13670 CSoutput.n254 CSoutput.n199 4.5005
R13671 CSoutput.n254 CSoutput.n203 4.5005
R13672 CSoutput.n254 CSoutput.n198 4.5005
R13673 CSoutput.n254 CSoutput.t146 4.5005
R13674 CSoutput.n254 CSoutput.n197 4.5005
R13675 CSoutput.n254 CSoutput.n204 4.5005
R13676 CSoutput.n254 CSoutput.n253 4.5005
R13677 CSoutput.n236 CSoutput.n200 4.5005
R13678 CSoutput.n236 CSoutput.n202 4.5005
R13679 CSoutput.n236 CSoutput.n199 4.5005
R13680 CSoutput.n236 CSoutput.n203 4.5005
R13681 CSoutput.n236 CSoutput.n198 4.5005
R13682 CSoutput.n236 CSoutput.t146 4.5005
R13683 CSoutput.n236 CSoutput.n197 4.5005
R13684 CSoutput.n236 CSoutput.n204 4.5005
R13685 CSoutput.n253 CSoutput.n236 4.5005
R13686 CSoutput.n208 CSoutput.n200 4.5005
R13687 CSoutput.n208 CSoutput.n202 4.5005
R13688 CSoutput.n208 CSoutput.n199 4.5005
R13689 CSoutput.n208 CSoutput.n203 4.5005
R13690 CSoutput.n208 CSoutput.n198 4.5005
R13691 CSoutput.n208 CSoutput.t146 4.5005
R13692 CSoutput.n208 CSoutput.n197 4.5005
R13693 CSoutput.n208 CSoutput.n204 4.5005
R13694 CSoutput.n253 CSoutput.n208 4.5005
R13695 CSoutput.n238 CSoutput.n200 4.5005
R13696 CSoutput.n238 CSoutput.n202 4.5005
R13697 CSoutput.n238 CSoutput.n199 4.5005
R13698 CSoutput.n238 CSoutput.n203 4.5005
R13699 CSoutput.n238 CSoutput.n198 4.5005
R13700 CSoutput.n238 CSoutput.t146 4.5005
R13701 CSoutput.n238 CSoutput.n197 4.5005
R13702 CSoutput.n238 CSoutput.n204 4.5005
R13703 CSoutput.n253 CSoutput.n238 4.5005
R13704 CSoutput.n207 CSoutput.n200 4.5005
R13705 CSoutput.n207 CSoutput.n202 4.5005
R13706 CSoutput.n207 CSoutput.n199 4.5005
R13707 CSoutput.n207 CSoutput.n203 4.5005
R13708 CSoutput.n207 CSoutput.n198 4.5005
R13709 CSoutput.n207 CSoutput.t146 4.5005
R13710 CSoutput.n207 CSoutput.n197 4.5005
R13711 CSoutput.n207 CSoutput.n204 4.5005
R13712 CSoutput.n253 CSoutput.n207 4.5005
R13713 CSoutput.n252 CSoutput.n200 4.5005
R13714 CSoutput.n252 CSoutput.n202 4.5005
R13715 CSoutput.n252 CSoutput.n199 4.5005
R13716 CSoutput.n252 CSoutput.n203 4.5005
R13717 CSoutput.n252 CSoutput.n198 4.5005
R13718 CSoutput.n252 CSoutput.t146 4.5005
R13719 CSoutput.n252 CSoutput.n197 4.5005
R13720 CSoutput.n252 CSoutput.n204 4.5005
R13721 CSoutput.n253 CSoutput.n252 4.5005
R13722 CSoutput.n251 CSoutput.n136 4.5005
R13723 CSoutput.n152 CSoutput.n136 4.5005
R13724 CSoutput.n147 CSoutput.n131 4.5005
R13725 CSoutput.n147 CSoutput.n133 4.5005
R13726 CSoutput.n147 CSoutput.n130 4.5005
R13727 CSoutput.n147 CSoutput.n134 4.5005
R13728 CSoutput.n147 CSoutput.n129 4.5005
R13729 CSoutput.n147 CSoutput.t163 4.5005
R13730 CSoutput.n147 CSoutput.n128 4.5005
R13731 CSoutput.n147 CSoutput.n135 4.5005
R13732 CSoutput.n147 CSoutput.n136 4.5005
R13733 CSoutput.n145 CSoutput.n131 4.5005
R13734 CSoutput.n145 CSoutput.n133 4.5005
R13735 CSoutput.n145 CSoutput.n130 4.5005
R13736 CSoutput.n145 CSoutput.n134 4.5005
R13737 CSoutput.n145 CSoutput.n129 4.5005
R13738 CSoutput.n145 CSoutput.t163 4.5005
R13739 CSoutput.n145 CSoutput.n128 4.5005
R13740 CSoutput.n145 CSoutput.n135 4.5005
R13741 CSoutput.n145 CSoutput.n136 4.5005
R13742 CSoutput.n144 CSoutput.n131 4.5005
R13743 CSoutput.n144 CSoutput.n133 4.5005
R13744 CSoutput.n144 CSoutput.n130 4.5005
R13745 CSoutput.n144 CSoutput.n134 4.5005
R13746 CSoutput.n144 CSoutput.n129 4.5005
R13747 CSoutput.n144 CSoutput.t163 4.5005
R13748 CSoutput.n144 CSoutput.n128 4.5005
R13749 CSoutput.n144 CSoutput.n135 4.5005
R13750 CSoutput.n144 CSoutput.n136 4.5005
R13751 CSoutput.n273 CSoutput.n131 4.5005
R13752 CSoutput.n273 CSoutput.n133 4.5005
R13753 CSoutput.n273 CSoutput.n130 4.5005
R13754 CSoutput.n273 CSoutput.n134 4.5005
R13755 CSoutput.n273 CSoutput.n129 4.5005
R13756 CSoutput.n273 CSoutput.t163 4.5005
R13757 CSoutput.n273 CSoutput.n128 4.5005
R13758 CSoutput.n273 CSoutput.n135 4.5005
R13759 CSoutput.n273 CSoutput.n136 4.5005
R13760 CSoutput.n271 CSoutput.n131 4.5005
R13761 CSoutput.n271 CSoutput.n133 4.5005
R13762 CSoutput.n271 CSoutput.n130 4.5005
R13763 CSoutput.n271 CSoutput.n134 4.5005
R13764 CSoutput.n271 CSoutput.n129 4.5005
R13765 CSoutput.n271 CSoutput.t163 4.5005
R13766 CSoutput.n271 CSoutput.n128 4.5005
R13767 CSoutput.n271 CSoutput.n135 4.5005
R13768 CSoutput.n269 CSoutput.n131 4.5005
R13769 CSoutput.n269 CSoutput.n133 4.5005
R13770 CSoutput.n269 CSoutput.n130 4.5005
R13771 CSoutput.n269 CSoutput.n134 4.5005
R13772 CSoutput.n269 CSoutput.n129 4.5005
R13773 CSoutput.n269 CSoutput.t163 4.5005
R13774 CSoutput.n269 CSoutput.n128 4.5005
R13775 CSoutput.n269 CSoutput.n135 4.5005
R13776 CSoutput.n155 CSoutput.n131 4.5005
R13777 CSoutput.n155 CSoutput.n133 4.5005
R13778 CSoutput.n155 CSoutput.n130 4.5005
R13779 CSoutput.n155 CSoutput.n134 4.5005
R13780 CSoutput.n155 CSoutput.n129 4.5005
R13781 CSoutput.n155 CSoutput.t163 4.5005
R13782 CSoutput.n155 CSoutput.n128 4.5005
R13783 CSoutput.n155 CSoutput.n135 4.5005
R13784 CSoutput.n155 CSoutput.n136 4.5005
R13785 CSoutput.n154 CSoutput.n131 4.5005
R13786 CSoutput.n154 CSoutput.n133 4.5005
R13787 CSoutput.n154 CSoutput.n130 4.5005
R13788 CSoutput.n154 CSoutput.n134 4.5005
R13789 CSoutput.n154 CSoutput.n129 4.5005
R13790 CSoutput.n154 CSoutput.t163 4.5005
R13791 CSoutput.n154 CSoutput.n128 4.5005
R13792 CSoutput.n154 CSoutput.n135 4.5005
R13793 CSoutput.n154 CSoutput.n136 4.5005
R13794 CSoutput.n158 CSoutput.n131 4.5005
R13795 CSoutput.n158 CSoutput.n133 4.5005
R13796 CSoutput.n158 CSoutput.n130 4.5005
R13797 CSoutput.n158 CSoutput.n134 4.5005
R13798 CSoutput.n158 CSoutput.n129 4.5005
R13799 CSoutput.n158 CSoutput.t163 4.5005
R13800 CSoutput.n158 CSoutput.n128 4.5005
R13801 CSoutput.n158 CSoutput.n135 4.5005
R13802 CSoutput.n158 CSoutput.n136 4.5005
R13803 CSoutput.n157 CSoutput.n131 4.5005
R13804 CSoutput.n157 CSoutput.n133 4.5005
R13805 CSoutput.n157 CSoutput.n130 4.5005
R13806 CSoutput.n157 CSoutput.n134 4.5005
R13807 CSoutput.n157 CSoutput.n129 4.5005
R13808 CSoutput.n157 CSoutput.t163 4.5005
R13809 CSoutput.n157 CSoutput.n128 4.5005
R13810 CSoutput.n157 CSoutput.n135 4.5005
R13811 CSoutput.n157 CSoutput.n136 4.5005
R13812 CSoutput.n140 CSoutput.n131 4.5005
R13813 CSoutput.n140 CSoutput.n133 4.5005
R13814 CSoutput.n140 CSoutput.n130 4.5005
R13815 CSoutput.n140 CSoutput.n134 4.5005
R13816 CSoutput.n140 CSoutput.n129 4.5005
R13817 CSoutput.n140 CSoutput.t163 4.5005
R13818 CSoutput.n140 CSoutput.n128 4.5005
R13819 CSoutput.n140 CSoutput.n135 4.5005
R13820 CSoutput.n140 CSoutput.n136 4.5005
R13821 CSoutput.n276 CSoutput.n131 4.5005
R13822 CSoutput.n276 CSoutput.n133 4.5005
R13823 CSoutput.n276 CSoutput.n130 4.5005
R13824 CSoutput.n276 CSoutput.n134 4.5005
R13825 CSoutput.n276 CSoutput.n129 4.5005
R13826 CSoutput.n276 CSoutput.t163 4.5005
R13827 CSoutput.n276 CSoutput.n128 4.5005
R13828 CSoutput.n276 CSoutput.n135 4.5005
R13829 CSoutput.n276 CSoutput.n136 4.5005
R13830 CSoutput.n323 CSoutput.n307 4.10845
R13831 CSoutput.n125 CSoutput.n109 4.10845
R13832 CSoutput.n321 CSoutput.t47 4.06363
R13833 CSoutput.n321 CSoutput.t135 4.06363
R13834 CSoutput.n319 CSoutput.t134 4.06363
R13835 CSoutput.n319 CSoutput.t69 4.06363
R13836 CSoutput.n317 CSoutput.t53 4.06363
R13837 CSoutput.n317 CSoutput.t140 4.06363
R13838 CSoutput.n315 CSoutput.t70 4.06363
R13839 CSoutput.n315 CSoutput.t20 4.06363
R13840 CSoutput.n313 CSoutput.t68 4.06363
R13841 CSoutput.n313 CSoutput.t19 4.06363
R13842 CSoutput.n311 CSoutput.t27 4.06363
R13843 CSoutput.n311 CSoutput.t39 4.06363
R13844 CSoutput.n309 CSoutput.t10 4.06363
R13845 CSoutput.n309 CSoutput.t52 4.06363
R13846 CSoutput.n308 CSoutput.t137 4.06363
R13847 CSoutput.n308 CSoutput.t46 4.06363
R13848 CSoutput.n305 CSoutput.t25 4.06363
R13849 CSoutput.n305 CSoutput.t77 4.06363
R13850 CSoutput.n303 CSoutput.t129 4.06363
R13851 CSoutput.n303 CSoutput.t71 4.06363
R13852 CSoutput.n301 CSoutput.t6 4.06363
R13853 CSoutput.n301 CSoutput.t21 4.06363
R13854 CSoutput.n299 CSoutput.t132 4.06363
R13855 CSoutput.n299 CSoutput.t4 4.06363
R13856 CSoutput.n297 CSoutput.t63 4.06363
R13857 CSoutput.n297 CSoutput.t75 4.06363
R13858 CSoutput.n295 CSoutput.t11 4.06363
R13859 CSoutput.n295 CSoutput.t79 4.06363
R13860 CSoutput.n293 CSoutput.t45 4.06363
R13861 CSoutput.n293 CSoutput.t48 4.06363
R13862 CSoutput.n292 CSoutput.t41 4.06363
R13863 CSoutput.n292 CSoutput.t37 4.06363
R13864 CSoutput.n290 CSoutput.t131 4.06363
R13865 CSoutput.n290 CSoutput.t65 4.06363
R13866 CSoutput.n288 CSoutput.t43 4.06363
R13867 CSoutput.n288 CSoutput.t31 4.06363
R13868 CSoutput.n286 CSoutput.t1 4.06363
R13869 CSoutput.n286 CSoutput.t66 4.06363
R13870 CSoutput.n284 CSoutput.t51 4.06363
R13871 CSoutput.n284 CSoutput.t16 4.06363
R13872 CSoutput.n282 CSoutput.t38 4.06363
R13873 CSoutput.n282 CSoutput.t74 4.06363
R13874 CSoutput.n280 CSoutput.t14 4.06363
R13875 CSoutput.n280 CSoutput.t50 4.06363
R13876 CSoutput.n278 CSoutput.t8 4.06363
R13877 CSoutput.n278 CSoutput.t56 4.06363
R13878 CSoutput.n277 CSoutput.t26 4.06363
R13879 CSoutput.n277 CSoutput.t78 4.06363
R13880 CSoutput.n110 CSoutput.t42 4.06363
R13881 CSoutput.n110 CSoutput.t67 4.06363
R13882 CSoutput.n111 CSoutput.t29 4.06363
R13883 CSoutput.n111 CSoutput.t139 4.06363
R13884 CSoutput.n113 CSoutput.t5 4.06363
R13885 CSoutput.n113 CSoutput.t24 4.06363
R13886 CSoutput.n115 CSoutput.t141 4.06363
R13887 CSoutput.n115 CSoutput.t142 4.06363
R13888 CSoutput.n117 CSoutput.t72 4.06363
R13889 CSoutput.n117 CSoutput.t76 4.06363
R13890 CSoutput.n119 CSoutput.t54 4.06363
R13891 CSoutput.n119 CSoutput.t58 4.06363
R13892 CSoutput.n121 CSoutput.t138 4.06363
R13893 CSoutput.n121 CSoutput.t9 4.06363
R13894 CSoutput.n123 CSoutput.t61 4.06363
R13895 CSoutput.n123 CSoutput.t32 4.06363
R13896 CSoutput.n94 CSoutput.t22 4.06363
R13897 CSoutput.n94 CSoutput.t23 4.06363
R13898 CSoutput.n95 CSoutput.t28 4.06363
R13899 CSoutput.n95 CSoutput.t136 4.06363
R13900 CSoutput.n97 CSoutput.t18 4.06363
R13901 CSoutput.n97 CSoutput.t133 4.06363
R13902 CSoutput.n99 CSoutput.t143 4.06363
R13903 CSoutput.n99 CSoutput.t73 4.06363
R13904 CSoutput.n101 CSoutput.t7 4.06363
R13905 CSoutput.n101 CSoutput.t128 4.06363
R13906 CSoutput.n103 CSoutput.t49 4.06363
R13907 CSoutput.n103 CSoutput.t30 4.06363
R13908 CSoutput.n105 CSoutput.t36 4.06363
R13909 CSoutput.n105 CSoutput.t15 4.06363
R13910 CSoutput.n107 CSoutput.t60 4.06363
R13911 CSoutput.n107 CSoutput.t59 4.06363
R13912 CSoutput.n79 CSoutput.t2 4.06363
R13913 CSoutput.n79 CSoutput.t13 4.06363
R13914 CSoutput.n80 CSoutput.t40 4.06363
R13915 CSoutput.n80 CSoutput.t55 4.06363
R13916 CSoutput.n82 CSoutput.t34 4.06363
R13917 CSoutput.n82 CSoutput.t33 4.06363
R13918 CSoutput.n84 CSoutput.t0 4.06363
R13919 CSoutput.n84 CSoutput.t57 4.06363
R13920 CSoutput.n86 CSoutput.t62 4.06363
R13921 CSoutput.n86 CSoutput.t35 4.06363
R13922 CSoutput.n88 CSoutput.t12 4.06363
R13923 CSoutput.n88 CSoutput.t3 4.06363
R13924 CSoutput.n90 CSoutput.t44 4.06363
R13925 CSoutput.n90 CSoutput.t17 4.06363
R13926 CSoutput.n92 CSoutput.t64 4.06363
R13927 CSoutput.n92 CSoutput.t130 4.06363
R13928 CSoutput.n44 CSoutput.n43 3.79402
R13929 CSoutput.n49 CSoutput.n48 3.79402
R13930 CSoutput.n373 CSoutput.n372 3.57343
R13931 CSoutput.n345 CSoutput.t118 2.82907
R13932 CSoutput.n345 CSoutput.t121 2.82907
R13933 CSoutput.n343 CSoutput.t117 2.82907
R13934 CSoutput.n343 CSoutput.t107 2.82907
R13935 CSoutput.n341 CSoutput.t84 2.82907
R13936 CSoutput.n341 CSoutput.t115 2.82907
R13937 CSoutput.n339 CSoutput.t109 2.82907
R13938 CSoutput.n339 CSoutput.t98 2.82907
R13939 CSoutput.n337 CSoutput.t126 2.82907
R13940 CSoutput.n337 CSoutput.t80 2.82907
R13941 CSoutput.n336 CSoutput.t114 2.82907
R13942 CSoutput.n336 CSoutput.t103 2.82907
R13943 CSoutput.n334 CSoutput.t111 2.82907
R13944 CSoutput.n334 CSoutput.t113 2.82907
R13945 CSoutput.n332 CSoutput.t108 2.82907
R13946 CSoutput.n332 CSoutput.t97 2.82907
R13947 CSoutput.n330 CSoutput.t125 2.82907
R13948 CSoutput.n330 CSoutput.t106 2.82907
R13949 CSoutput.n328 CSoutput.t99 2.82907
R13950 CSoutput.n328 CSoutput.t89 2.82907
R13951 CSoutput.n326 CSoutput.t120 2.82907
R13952 CSoutput.n326 CSoutput.t122 2.82907
R13953 CSoutput.n325 CSoutput.t104 2.82907
R13954 CSoutput.n325 CSoutput.t94 2.82907
R13955 CSoutput.n360 CSoutput.t90 2.82907
R13956 CSoutput.n360 CSoutput.t102 2.82907
R13957 CSoutput.n361 CSoutput.t119 2.82907
R13958 CSoutput.n361 CSoutput.t82 2.82907
R13959 CSoutput.n363 CSoutput.t86 2.82907
R13960 CSoutput.n363 CSoutput.t96 2.82907
R13961 CSoutput.n365 CSoutput.t101 2.82907
R13962 CSoutput.n365 CSoutput.t88 2.82907
R13963 CSoutput.n367 CSoutput.t93 2.82907
R13964 CSoutput.n367 CSoutput.t105 2.82907
R13965 CSoutput.n369 CSoutput.t110 2.82907
R13966 CSoutput.n369 CSoutput.t123 2.82907
R13967 CSoutput.n349 CSoutput.t83 2.82907
R13968 CSoutput.n349 CSoutput.t91 2.82907
R13969 CSoutput.n350 CSoutput.t112 2.82907
R13970 CSoutput.n350 CSoutput.t124 2.82907
R13971 CSoutput.n352 CSoutput.t127 2.82907
R13972 CSoutput.n352 CSoutput.t87 2.82907
R13973 CSoutput.n354 CSoutput.t92 2.82907
R13974 CSoutput.n354 CSoutput.t81 2.82907
R13975 CSoutput.n356 CSoutput.t85 2.82907
R13976 CSoutput.n356 CSoutput.t95 2.82907
R13977 CSoutput.n358 CSoutput.t100 2.82907
R13978 CSoutput.n358 CSoutput.t116 2.82907
R13979 CSoutput.n372 CSoutput.n348 2.75627
R13980 CSoutput.n75 CSoutput.n1 2.45513
R13981 CSoutput.n324 CSoutput.n126 2.36742
R13982 CSoutput.n217 CSoutput.n215 2.251
R13983 CSoutput.n217 CSoutput.n214 2.251
R13984 CSoutput.n217 CSoutput.n213 2.251
R13985 CSoutput.n217 CSoutput.n212 2.251
R13986 CSoutput.n186 CSoutput.n185 2.251
R13987 CSoutput.n186 CSoutput.n184 2.251
R13988 CSoutput.n186 CSoutput.n183 2.251
R13989 CSoutput.n186 CSoutput.n182 2.251
R13990 CSoutput.n259 CSoutput.n258 2.251
R13991 CSoutput.n224 CSoutput.n222 2.251
R13992 CSoutput.n224 CSoutput.n221 2.251
R13993 CSoutput.n224 CSoutput.n220 2.251
R13994 CSoutput.n242 CSoutput.n224 2.251
R13995 CSoutput.n230 CSoutput.n229 2.251
R13996 CSoutput.n230 CSoutput.n228 2.251
R13997 CSoutput.n230 CSoutput.n227 2.251
R13998 CSoutput.n230 CSoutput.n226 2.251
R13999 CSoutput.n256 CSoutput.n196 2.251
R14000 CSoutput.n251 CSoutput.n249 2.251
R14001 CSoutput.n251 CSoutput.n248 2.251
R14002 CSoutput.n251 CSoutput.n247 2.251
R14003 CSoutput.n251 CSoutput.n246 2.251
R14004 CSoutput.n152 CSoutput.n151 2.251
R14005 CSoutput.n152 CSoutput.n150 2.251
R14006 CSoutput.n152 CSoutput.n149 2.251
R14007 CSoutput.n152 CSoutput.n148 2.251
R14008 CSoutput.n269 CSoutput.n268 2.251
R14009 CSoutput.n186 CSoutput.n166 2.2505
R14010 CSoutput.n181 CSoutput.n166 2.2505
R14011 CSoutput.n179 CSoutput.n166 2.2505
R14012 CSoutput.n178 CSoutput.n166 2.2505
R14013 CSoutput.n263 CSoutput.n166 2.2505
R14014 CSoutput.n261 CSoutput.n166 2.2505
R14015 CSoutput.n259 CSoutput.n166 2.2505
R14016 CSoutput.n189 CSoutput.n166 2.2505
R14017 CSoutput.n188 CSoutput.n166 2.2505
R14018 CSoutput.n192 CSoutput.n166 2.2505
R14019 CSoutput.n191 CSoutput.n166 2.2505
R14020 CSoutput.n174 CSoutput.n166 2.2505
R14021 CSoutput.n266 CSoutput.n166 2.2505
R14022 CSoutput.n266 CSoutput.n265 2.2505
R14023 CSoutput.n230 CSoutput.n201 2.2505
R14024 CSoutput.n211 CSoutput.n201 2.2505
R14025 CSoutput.n232 CSoutput.n201 2.2505
R14026 CSoutput.n210 CSoutput.n201 2.2505
R14027 CSoutput.n234 CSoutput.n201 2.2505
R14028 CSoutput.n201 CSoutput.n195 2.2505
R14029 CSoutput.n256 CSoutput.n201 2.2505
R14030 CSoutput.n254 CSoutput.n201 2.2505
R14031 CSoutput.n236 CSoutput.n201 2.2505
R14032 CSoutput.n208 CSoutput.n201 2.2505
R14033 CSoutput.n238 CSoutput.n201 2.2505
R14034 CSoutput.n207 CSoutput.n201 2.2505
R14035 CSoutput.n252 CSoutput.n201 2.2505
R14036 CSoutput.n252 CSoutput.n205 2.2505
R14037 CSoutput.n152 CSoutput.n132 2.2505
R14038 CSoutput.n147 CSoutput.n132 2.2505
R14039 CSoutput.n145 CSoutput.n132 2.2505
R14040 CSoutput.n144 CSoutput.n132 2.2505
R14041 CSoutput.n273 CSoutput.n132 2.2505
R14042 CSoutput.n271 CSoutput.n132 2.2505
R14043 CSoutput.n269 CSoutput.n132 2.2505
R14044 CSoutput.n155 CSoutput.n132 2.2505
R14045 CSoutput.n154 CSoutput.n132 2.2505
R14046 CSoutput.n158 CSoutput.n132 2.2505
R14047 CSoutput.n157 CSoutput.n132 2.2505
R14048 CSoutput.n140 CSoutput.n132 2.2505
R14049 CSoutput.n276 CSoutput.n132 2.2505
R14050 CSoutput.n276 CSoutput.n275 2.2505
R14051 CSoutput.n194 CSoutput.n187 2.25024
R14052 CSoutput.n194 CSoutput.n180 2.25024
R14053 CSoutput.n262 CSoutput.n194 2.25024
R14054 CSoutput.n194 CSoutput.n190 2.25024
R14055 CSoutput.n194 CSoutput.n193 2.25024
R14056 CSoutput.n194 CSoutput.n161 2.25024
R14057 CSoutput.n244 CSoutput.n241 2.25024
R14058 CSoutput.n244 CSoutput.n240 2.25024
R14059 CSoutput.n244 CSoutput.n239 2.25024
R14060 CSoutput.n244 CSoutput.n206 2.25024
R14061 CSoutput.n244 CSoutput.n243 2.25024
R14062 CSoutput.n245 CSoutput.n244 2.25024
R14063 CSoutput.n160 CSoutput.n153 2.25024
R14064 CSoutput.n160 CSoutput.n146 2.25024
R14065 CSoutput.n272 CSoutput.n160 2.25024
R14066 CSoutput.n160 CSoutput.n156 2.25024
R14067 CSoutput.n160 CSoutput.n159 2.25024
R14068 CSoutput.n160 CSoutput.n127 2.25024
R14069 CSoutput.n261 CSoutput.n171 1.50111
R14070 CSoutput.n209 CSoutput.n195 1.50111
R14071 CSoutput.n271 CSoutput.n137 1.50111
R14072 CSoutput.n217 CSoutput.n216 1.501
R14073 CSoutput.n224 CSoutput.n223 1.501
R14074 CSoutput.n251 CSoutput.n250 1.501
R14075 CSoutput.n265 CSoutput.n176 1.12536
R14076 CSoutput.n265 CSoutput.n177 1.12536
R14077 CSoutput.n265 CSoutput.n264 1.12536
R14078 CSoutput.n225 CSoutput.n205 1.12536
R14079 CSoutput.n231 CSoutput.n205 1.12536
R14080 CSoutput.n233 CSoutput.n205 1.12536
R14081 CSoutput.n275 CSoutput.n142 1.12536
R14082 CSoutput.n275 CSoutput.n143 1.12536
R14083 CSoutput.n275 CSoutput.n274 1.12536
R14084 CSoutput.n265 CSoutput.n172 1.12536
R14085 CSoutput.n265 CSoutput.n173 1.12536
R14086 CSoutput.n265 CSoutput.n175 1.12536
R14087 CSoutput.n255 CSoutput.n205 1.12536
R14088 CSoutput.n235 CSoutput.n205 1.12536
R14089 CSoutput.n237 CSoutput.n205 1.12536
R14090 CSoutput.n275 CSoutput.n138 1.12536
R14091 CSoutput.n275 CSoutput.n139 1.12536
R14092 CSoutput.n275 CSoutput.n141 1.12536
R14093 CSoutput.n31 CSoutput.n30 0.669944
R14094 CSoutput.n62 CSoutput.n61 0.669944
R14095 CSoutput.n340 CSoutput.n338 0.573776
R14096 CSoutput.n342 CSoutput.n340 0.573776
R14097 CSoutput.n344 CSoutput.n342 0.573776
R14098 CSoutput.n346 CSoutput.n344 0.573776
R14099 CSoutput.n329 CSoutput.n327 0.573776
R14100 CSoutput.n331 CSoutput.n329 0.573776
R14101 CSoutput.n333 CSoutput.n331 0.573776
R14102 CSoutput.n335 CSoutput.n333 0.573776
R14103 CSoutput.n370 CSoutput.n368 0.573776
R14104 CSoutput.n368 CSoutput.n366 0.573776
R14105 CSoutput.n366 CSoutput.n364 0.573776
R14106 CSoutput.n364 CSoutput.n362 0.573776
R14107 CSoutput.n359 CSoutput.n357 0.573776
R14108 CSoutput.n357 CSoutput.n355 0.573776
R14109 CSoutput.n355 CSoutput.n353 0.573776
R14110 CSoutput.n353 CSoutput.n351 0.573776
R14111 CSoutput.n373 CSoutput.n276 0.53442
R14112 CSoutput.n312 CSoutput.n310 0.358259
R14113 CSoutput.n314 CSoutput.n312 0.358259
R14114 CSoutput.n316 CSoutput.n314 0.358259
R14115 CSoutput.n318 CSoutput.n316 0.358259
R14116 CSoutput.n320 CSoutput.n318 0.358259
R14117 CSoutput.n322 CSoutput.n320 0.358259
R14118 CSoutput.n296 CSoutput.n294 0.358259
R14119 CSoutput.n298 CSoutput.n296 0.358259
R14120 CSoutput.n300 CSoutput.n298 0.358259
R14121 CSoutput.n302 CSoutput.n300 0.358259
R14122 CSoutput.n304 CSoutput.n302 0.358259
R14123 CSoutput.n306 CSoutput.n304 0.358259
R14124 CSoutput.n281 CSoutput.n279 0.358259
R14125 CSoutput.n283 CSoutput.n281 0.358259
R14126 CSoutput.n285 CSoutput.n283 0.358259
R14127 CSoutput.n287 CSoutput.n285 0.358259
R14128 CSoutput.n289 CSoutput.n287 0.358259
R14129 CSoutput.n291 CSoutput.n289 0.358259
R14130 CSoutput.n124 CSoutput.n122 0.358259
R14131 CSoutput.n122 CSoutput.n120 0.358259
R14132 CSoutput.n120 CSoutput.n118 0.358259
R14133 CSoutput.n118 CSoutput.n116 0.358259
R14134 CSoutput.n116 CSoutput.n114 0.358259
R14135 CSoutput.n114 CSoutput.n112 0.358259
R14136 CSoutput.n108 CSoutput.n106 0.358259
R14137 CSoutput.n106 CSoutput.n104 0.358259
R14138 CSoutput.n104 CSoutput.n102 0.358259
R14139 CSoutput.n102 CSoutput.n100 0.358259
R14140 CSoutput.n100 CSoutput.n98 0.358259
R14141 CSoutput.n98 CSoutput.n96 0.358259
R14142 CSoutput.n93 CSoutput.n91 0.358259
R14143 CSoutput.n91 CSoutput.n89 0.358259
R14144 CSoutput.n89 CSoutput.n87 0.358259
R14145 CSoutput.n87 CSoutput.n85 0.358259
R14146 CSoutput.n85 CSoutput.n83 0.358259
R14147 CSoutput.n83 CSoutput.n81 0.358259
R14148 CSoutput.n21 CSoutput.n20 0.169105
R14149 CSoutput.n21 CSoutput.n16 0.169105
R14150 CSoutput.n26 CSoutput.n16 0.169105
R14151 CSoutput.n27 CSoutput.n26 0.169105
R14152 CSoutput.n27 CSoutput.n14 0.169105
R14153 CSoutput.n32 CSoutput.n14 0.169105
R14154 CSoutput.n33 CSoutput.n32 0.169105
R14155 CSoutput.n34 CSoutput.n33 0.169105
R14156 CSoutput.n34 CSoutput.n12 0.169105
R14157 CSoutput.n39 CSoutput.n12 0.169105
R14158 CSoutput.n40 CSoutput.n39 0.169105
R14159 CSoutput.n40 CSoutput.n10 0.169105
R14160 CSoutput.n45 CSoutput.n10 0.169105
R14161 CSoutput.n46 CSoutput.n45 0.169105
R14162 CSoutput.n47 CSoutput.n46 0.169105
R14163 CSoutput.n47 CSoutput.n8 0.169105
R14164 CSoutput.n52 CSoutput.n8 0.169105
R14165 CSoutput.n53 CSoutput.n52 0.169105
R14166 CSoutput.n53 CSoutput.n6 0.169105
R14167 CSoutput.n58 CSoutput.n6 0.169105
R14168 CSoutput.n59 CSoutput.n58 0.169105
R14169 CSoutput.n60 CSoutput.n59 0.169105
R14170 CSoutput.n60 CSoutput.n4 0.169105
R14171 CSoutput.n66 CSoutput.n4 0.169105
R14172 CSoutput.n67 CSoutput.n66 0.169105
R14173 CSoutput.n68 CSoutput.n67 0.169105
R14174 CSoutput.n68 CSoutput.n2 0.169105
R14175 CSoutput.n73 CSoutput.n2 0.169105
R14176 CSoutput.n74 CSoutput.n73 0.169105
R14177 CSoutput.n74 CSoutput.n0 0.169105
R14178 CSoutput.n78 CSoutput.n0 0.169105
R14179 CSoutput.n219 CSoutput.n218 0.0910737
R14180 CSoutput.n270 CSoutput.n267 0.0723685
R14181 CSoutput.n224 CSoutput.n219 0.0522944
R14182 CSoutput.n267 CSoutput.n266 0.0499135
R14183 CSoutput.n218 CSoutput.n217 0.0499135
R14184 CSoutput.n252 CSoutput.n251 0.0464294
R14185 CSoutput.n260 CSoutput.n257 0.0391444
R14186 CSoutput.n219 CSoutput.t153 0.023435
R14187 CSoutput.n267 CSoutput.t152 0.02262
R14188 CSoutput.n218 CSoutput.t157 0.02262
R14189 CSoutput CSoutput.n373 0.0052
R14190 CSoutput.n189 CSoutput.n172 0.00365111
R14191 CSoutput.n192 CSoutput.n173 0.00365111
R14192 CSoutput.n175 CSoutput.n174 0.00365111
R14193 CSoutput.n217 CSoutput.n176 0.00365111
R14194 CSoutput.n181 CSoutput.n177 0.00365111
R14195 CSoutput.n264 CSoutput.n178 0.00365111
R14196 CSoutput.n255 CSoutput.n254 0.00365111
R14197 CSoutput.n235 CSoutput.n208 0.00365111
R14198 CSoutput.n237 CSoutput.n207 0.00365111
R14199 CSoutput.n225 CSoutput.n224 0.00365111
R14200 CSoutput.n231 CSoutput.n211 0.00365111
R14201 CSoutput.n233 CSoutput.n210 0.00365111
R14202 CSoutput.n155 CSoutput.n138 0.00365111
R14203 CSoutput.n158 CSoutput.n139 0.00365111
R14204 CSoutput.n141 CSoutput.n140 0.00365111
R14205 CSoutput.n251 CSoutput.n142 0.00365111
R14206 CSoutput.n147 CSoutput.n143 0.00365111
R14207 CSoutput.n274 CSoutput.n144 0.00365111
R14208 CSoutput.n186 CSoutput.n176 0.00340054
R14209 CSoutput.n179 CSoutput.n177 0.00340054
R14210 CSoutput.n264 CSoutput.n263 0.00340054
R14211 CSoutput.n259 CSoutput.n172 0.00340054
R14212 CSoutput.n188 CSoutput.n173 0.00340054
R14213 CSoutput.n191 CSoutput.n175 0.00340054
R14214 CSoutput.n230 CSoutput.n225 0.00340054
R14215 CSoutput.n232 CSoutput.n231 0.00340054
R14216 CSoutput.n234 CSoutput.n233 0.00340054
R14217 CSoutput.n256 CSoutput.n255 0.00340054
R14218 CSoutput.n236 CSoutput.n235 0.00340054
R14219 CSoutput.n238 CSoutput.n237 0.00340054
R14220 CSoutput.n152 CSoutput.n142 0.00340054
R14221 CSoutput.n145 CSoutput.n143 0.00340054
R14222 CSoutput.n274 CSoutput.n273 0.00340054
R14223 CSoutput.n269 CSoutput.n138 0.00340054
R14224 CSoutput.n154 CSoutput.n139 0.00340054
R14225 CSoutput.n157 CSoutput.n141 0.00340054
R14226 CSoutput.n187 CSoutput.n181 0.00252698
R14227 CSoutput.n180 CSoutput.n178 0.00252698
R14228 CSoutput.n262 CSoutput.n261 0.00252698
R14229 CSoutput.n190 CSoutput.n188 0.00252698
R14230 CSoutput.n193 CSoutput.n191 0.00252698
R14231 CSoutput.n266 CSoutput.n161 0.00252698
R14232 CSoutput.n187 CSoutput.n186 0.00252698
R14233 CSoutput.n180 CSoutput.n179 0.00252698
R14234 CSoutput.n263 CSoutput.n262 0.00252698
R14235 CSoutput.n190 CSoutput.n189 0.00252698
R14236 CSoutput.n193 CSoutput.n192 0.00252698
R14237 CSoutput.n174 CSoutput.n161 0.00252698
R14238 CSoutput.n241 CSoutput.n211 0.00252698
R14239 CSoutput.n240 CSoutput.n210 0.00252698
R14240 CSoutput.n239 CSoutput.n195 0.00252698
R14241 CSoutput.n236 CSoutput.n206 0.00252698
R14242 CSoutput.n243 CSoutput.n238 0.00252698
R14243 CSoutput.n252 CSoutput.n245 0.00252698
R14244 CSoutput.n241 CSoutput.n230 0.00252698
R14245 CSoutput.n240 CSoutput.n232 0.00252698
R14246 CSoutput.n239 CSoutput.n234 0.00252698
R14247 CSoutput.n254 CSoutput.n206 0.00252698
R14248 CSoutput.n243 CSoutput.n208 0.00252698
R14249 CSoutput.n245 CSoutput.n207 0.00252698
R14250 CSoutput.n153 CSoutput.n147 0.00252698
R14251 CSoutput.n146 CSoutput.n144 0.00252698
R14252 CSoutput.n272 CSoutput.n271 0.00252698
R14253 CSoutput.n156 CSoutput.n154 0.00252698
R14254 CSoutput.n159 CSoutput.n157 0.00252698
R14255 CSoutput.n276 CSoutput.n127 0.00252698
R14256 CSoutput.n153 CSoutput.n152 0.00252698
R14257 CSoutput.n146 CSoutput.n145 0.00252698
R14258 CSoutput.n273 CSoutput.n272 0.00252698
R14259 CSoutput.n156 CSoutput.n155 0.00252698
R14260 CSoutput.n159 CSoutput.n158 0.00252698
R14261 CSoutput.n140 CSoutput.n127 0.00252698
R14262 CSoutput.n261 CSoutput.n260 0.0020275
R14263 CSoutput.n260 CSoutput.n259 0.0020275
R14264 CSoutput.n257 CSoutput.n195 0.0020275
R14265 CSoutput.n257 CSoutput.n256 0.0020275
R14266 CSoutput.n271 CSoutput.n270 0.0020275
R14267 CSoutput.n270 CSoutput.n269 0.0020275
R14268 CSoutput.n171 CSoutput.n170 0.00166668
R14269 CSoutput.n253 CSoutput.n209 0.00166668
R14270 CSoutput.n137 CSoutput.n136 0.00166668
R14271 CSoutput.n275 CSoutput.n137 0.00133328
R14272 CSoutput.n209 CSoutput.n205 0.00133328
R14273 CSoutput.n265 CSoutput.n171 0.00133328
R14274 CSoutput.n268 CSoutput.n160 0.001
R14275 CSoutput.n246 CSoutput.n160 0.001
R14276 CSoutput.n148 CSoutput.n128 0.001
R14277 CSoutput.n247 CSoutput.n128 0.001
R14278 CSoutput.n149 CSoutput.n129 0.001
R14279 CSoutput.n248 CSoutput.n129 0.001
R14280 CSoutput.n150 CSoutput.n130 0.001
R14281 CSoutput.n249 CSoutput.n130 0.001
R14282 CSoutput.n151 CSoutput.n131 0.001
R14283 CSoutput.n250 CSoutput.n131 0.001
R14284 CSoutput.n244 CSoutput.n196 0.001
R14285 CSoutput.n244 CSoutput.n242 0.001
R14286 CSoutput.n226 CSoutput.n197 0.001
R14287 CSoutput.n220 CSoutput.n197 0.001
R14288 CSoutput.n227 CSoutput.n198 0.001
R14289 CSoutput.n221 CSoutput.n198 0.001
R14290 CSoutput.n228 CSoutput.n199 0.001
R14291 CSoutput.n222 CSoutput.n199 0.001
R14292 CSoutput.n229 CSoutput.n200 0.001
R14293 CSoutput.n223 CSoutput.n200 0.001
R14294 CSoutput.n258 CSoutput.n194 0.001
R14295 CSoutput.n212 CSoutput.n194 0.001
R14296 CSoutput.n182 CSoutput.n162 0.001
R14297 CSoutput.n213 CSoutput.n162 0.001
R14298 CSoutput.n183 CSoutput.n163 0.001
R14299 CSoutput.n214 CSoutput.n163 0.001
R14300 CSoutput.n184 CSoutput.n164 0.001
R14301 CSoutput.n215 CSoutput.n164 0.001
R14302 CSoutput.n185 CSoutput.n165 0.001
R14303 CSoutput.n216 CSoutput.n165 0.001
R14304 CSoutput.n216 CSoutput.n166 0.001
R14305 CSoutput.n215 CSoutput.n167 0.001
R14306 CSoutput.n214 CSoutput.n168 0.001
R14307 CSoutput.n213 CSoutput.t150 0.001
R14308 CSoutput.n212 CSoutput.n169 0.001
R14309 CSoutput.n185 CSoutput.n167 0.001
R14310 CSoutput.n184 CSoutput.n168 0.001
R14311 CSoutput.n183 CSoutput.t150 0.001
R14312 CSoutput.n182 CSoutput.n169 0.001
R14313 CSoutput.n258 CSoutput.n170 0.001
R14314 CSoutput.n223 CSoutput.n201 0.001
R14315 CSoutput.n222 CSoutput.n202 0.001
R14316 CSoutput.n221 CSoutput.n203 0.001
R14317 CSoutput.n220 CSoutput.t146 0.001
R14318 CSoutput.n242 CSoutput.n204 0.001
R14319 CSoutput.n229 CSoutput.n202 0.001
R14320 CSoutput.n228 CSoutput.n203 0.001
R14321 CSoutput.n227 CSoutput.t146 0.001
R14322 CSoutput.n226 CSoutput.n204 0.001
R14323 CSoutput.n253 CSoutput.n196 0.001
R14324 CSoutput.n250 CSoutput.n132 0.001
R14325 CSoutput.n249 CSoutput.n133 0.001
R14326 CSoutput.n248 CSoutput.n134 0.001
R14327 CSoutput.n247 CSoutput.t163 0.001
R14328 CSoutput.n246 CSoutput.n135 0.001
R14329 CSoutput.n151 CSoutput.n133 0.001
R14330 CSoutput.n150 CSoutput.n134 0.001
R14331 CSoutput.n149 CSoutput.t163 0.001
R14332 CSoutput.n148 CSoutput.n135 0.001
R14333 CSoutput.n268 CSoutput.n136 0.001
R14334 a_n6972_8799.n184 a_n6972_8799.t57 485.149
R14335 a_n6972_8799.n200 a_n6972_8799.t71 485.149
R14336 a_n6972_8799.n217 a_n6972_8799.t120 485.149
R14337 a_n6972_8799.n133 a_n6972_8799.t115 485.149
R14338 a_n6972_8799.n149 a_n6972_8799.t125 485.149
R14339 a_n6972_8799.n166 a_n6972_8799.t118 485.149
R14340 a_n6972_8799.n194 a_n6972_8799.t80 464.166
R14341 a_n6972_8799.n193 a_n6972_8799.t79 464.166
R14342 a_n6972_8799.n179 a_n6972_8799.t58 464.166
R14343 a_n6972_8799.n192 a_n6972_8799.t116 464.166
R14344 a_n6972_8799.n191 a_n6972_8799.t81 464.166
R14345 a_n6972_8799.n180 a_n6972_8799.t63 464.166
R14346 a_n6972_8799.n190 a_n6972_8799.t119 464.166
R14347 a_n6972_8799.n189 a_n6972_8799.t95 464.166
R14348 a_n6972_8799.n181 a_n6972_8799.t93 464.166
R14349 a_n6972_8799.n188 a_n6972_8799.t40 464.166
R14350 a_n6972_8799.n187 a_n6972_8799.t99 464.166
R14351 a_n6972_8799.n182 a_n6972_8799.t98 464.166
R14352 a_n6972_8799.n186 a_n6972_8799.t42 464.166
R14353 a_n6972_8799.n185 a_n6972_8799.t41 464.166
R14354 a_n6972_8799.n183 a_n6972_8799.t112 464.166
R14355 a_n6972_8799.n210 a_n6972_8799.t87 464.166
R14356 a_n6972_8799.n209 a_n6972_8799.t86 464.166
R14357 a_n6972_8799.n195 a_n6972_8799.t70 464.166
R14358 a_n6972_8799.n208 a_n6972_8799.t128 464.166
R14359 a_n6972_8799.n207 a_n6972_8799.t92 464.166
R14360 a_n6972_8799.n196 a_n6972_8799.t72 464.166
R14361 a_n6972_8799.n206 a_n6972_8799.t36 464.166
R14362 a_n6972_8799.n205 a_n6972_8799.t105 464.166
R14363 a_n6972_8799.n197 a_n6972_8799.t104 464.166
R14364 a_n6972_8799.n204 a_n6972_8799.t49 464.166
R14365 a_n6972_8799.n203 a_n6972_8799.t108 464.166
R14366 a_n6972_8799.n198 a_n6972_8799.t107 464.166
R14367 a_n6972_8799.n202 a_n6972_8799.t53 464.166
R14368 a_n6972_8799.n201 a_n6972_8799.t52 464.166
R14369 a_n6972_8799.n199 a_n6972_8799.t123 464.166
R14370 a_n6972_8799.n227 a_n6972_8799.t130 464.166
R14371 a_n6972_8799.n226 a_n6972_8799.t51 464.166
R14372 a_n6972_8799.n212 a_n6972_8799.t90 464.166
R14373 a_n6972_8799.n225 a_n6972_8799.t38 464.166
R14374 a_n6972_8799.n224 a_n6972_8799.t110 464.166
R14375 a_n6972_8799.n213 a_n6972_8799.t62 464.166
R14376 a_n6972_8799.n223 a_n6972_8799.t96 464.166
R14377 a_n6972_8799.n222 a_n6972_8799.t43 464.166
R14378 a_n6972_8799.n214 a_n6972_8799.t66 464.166
R14379 a_n6972_8799.n221 a_n6972_8799.t126 464.166
R14380 a_n6972_8799.n220 a_n6972_8799.t102 464.166
R14381 a_n6972_8799.n215 a_n6972_8799.t122 464.166
R14382 a_n6972_8799.n219 a_n6972_8799.t89 464.166
R14383 a_n6972_8799.n218 a_n6972_8799.t106 464.166
R14384 a_n6972_8799.n216 a_n6972_8799.t56 464.166
R14385 a_n6972_8799.n132 a_n6972_8799.t78 464.166
R14386 a_n6972_8799.n135 a_n6972_8799.t77 464.166
R14387 a_n6972_8799.n131 a_n6972_8799.t101 464.166
R14388 a_n6972_8799.n136 a_n6972_8799.t68 464.166
R14389 a_n6972_8799.n137 a_n6972_8799.t69 464.166
R14390 a_n6972_8799.n138 a_n6972_8799.t100 464.166
R14391 a_n6972_8799.n139 a_n6972_8799.t37 464.166
R14392 a_n6972_8799.n130 a_n6972_8799.t65 464.166
R14393 a_n6972_8799.n140 a_n6972_8799.t83 464.166
R14394 a_n6972_8799.n141 a_n6972_8799.t117 464.166
R14395 a_n6972_8799.n142 a_n6972_8799.t47 464.166
R14396 a_n6972_8799.n143 a_n6972_8799.t64 464.166
R14397 a_n6972_8799.n129 a_n6972_8799.t114 464.166
R14398 a_n6972_8799.n144 a_n6972_8799.t46 464.166
R14399 a_n6972_8799.n148 a_n6972_8799.t84 464.166
R14400 a_n6972_8799.n151 a_n6972_8799.t85 464.166
R14401 a_n6972_8799.n147 a_n6972_8799.t113 464.166
R14402 a_n6972_8799.n152 a_n6972_8799.t75 464.166
R14403 a_n6972_8799.n153 a_n6972_8799.t76 464.166
R14404 a_n6972_8799.n154 a_n6972_8799.t109 464.166
R14405 a_n6972_8799.n155 a_n6972_8799.t48 464.166
R14406 a_n6972_8799.n146 a_n6972_8799.t74 464.166
R14407 a_n6972_8799.n156 a_n6972_8799.t94 464.166
R14408 a_n6972_8799.n157 a_n6972_8799.t129 464.166
R14409 a_n6972_8799.n158 a_n6972_8799.t61 464.166
R14410 a_n6972_8799.n159 a_n6972_8799.t73 464.166
R14411 a_n6972_8799.n145 a_n6972_8799.t124 464.166
R14412 a_n6972_8799.n160 a_n6972_8799.t55 464.166
R14413 a_n6972_8799.n165 a_n6972_8799.t54 464.166
R14414 a_n6972_8799.n168 a_n6972_8799.t39 464.166
R14415 a_n6972_8799.n164 a_n6972_8799.t88 464.166
R14416 a_n6972_8799.n169 a_n6972_8799.t121 464.166
R14417 a_n6972_8799.n170 a_n6972_8799.t103 464.166
R14418 a_n6972_8799.n171 a_n6972_8799.t127 464.166
R14419 a_n6972_8799.n172 a_n6972_8799.t82 464.166
R14420 a_n6972_8799.n163 a_n6972_8799.t44 464.166
R14421 a_n6972_8799.n173 a_n6972_8799.t97 464.166
R14422 a_n6972_8799.n174 a_n6972_8799.t60 464.166
R14423 a_n6972_8799.n175 a_n6972_8799.t111 464.166
R14424 a_n6972_8799.n176 a_n6972_8799.t67 464.166
R14425 a_n6972_8799.n162 a_n6972_8799.t91 464.166
R14426 a_n6972_8799.n177 a_n6972_8799.t50 464.166
R14427 a_n6972_8799.n52 a_n6972_8799.n30 74.4178
R14428 a_n6972_8799.n185 a_n6972_8799.n52 12.4674
R14429 a_n6972_8799.n51 a_n6972_8799.n30 80.107
R14430 a_n6972_8799.n51 a_n6972_8799.n186 1.08907
R14431 a_n6972_8799.n31 a_n6972_8799.n50 75.3623
R14432 a_n6972_8799.n49 a_n6972_8799.n31 70.3058
R14433 a_n6972_8799.n33 a_n6972_8799.n48 70.1674
R14434 a_n6972_8799.n48 a_n6972_8799.n181 20.9683
R14435 a_n6972_8799.n47 a_n6972_8799.n33 75.0448
R14436 a_n6972_8799.n189 a_n6972_8799.n47 11.2134
R14437 a_n6972_8799.n46 a_n6972_8799.n32 80.4688
R14438 a_n6972_8799.n32 a_n6972_8799.n45 74.73
R14439 a_n6972_8799.n44 a_n6972_8799.n34 70.1674
R14440 a_n6972_8799.n192 a_n6972_8799.n44 20.9683
R14441 a_n6972_8799.n34 a_n6972_8799.n43 70.5844
R14442 a_n6972_8799.n43 a_n6972_8799.n179 20.1342
R14443 a_n6972_8799.n42 a_n6972_8799.n35 75.6825
R14444 a_n6972_8799.n193 a_n6972_8799.n42 9.93802
R14445 a_n6972_8799.n35 a_n6972_8799.n194 161.3
R14446 a_n6972_8799.n63 a_n6972_8799.n24 74.4178
R14447 a_n6972_8799.n201 a_n6972_8799.n63 12.4674
R14448 a_n6972_8799.n62 a_n6972_8799.n24 80.107
R14449 a_n6972_8799.n62 a_n6972_8799.n202 1.08907
R14450 a_n6972_8799.n25 a_n6972_8799.n61 75.3623
R14451 a_n6972_8799.n60 a_n6972_8799.n25 70.3058
R14452 a_n6972_8799.n27 a_n6972_8799.n59 70.1674
R14453 a_n6972_8799.n59 a_n6972_8799.n197 20.9683
R14454 a_n6972_8799.n58 a_n6972_8799.n27 75.0448
R14455 a_n6972_8799.n205 a_n6972_8799.n58 11.2134
R14456 a_n6972_8799.n57 a_n6972_8799.n26 80.4688
R14457 a_n6972_8799.n26 a_n6972_8799.n56 74.73
R14458 a_n6972_8799.n55 a_n6972_8799.n28 70.1674
R14459 a_n6972_8799.n208 a_n6972_8799.n55 20.9683
R14460 a_n6972_8799.n28 a_n6972_8799.n54 70.5844
R14461 a_n6972_8799.n54 a_n6972_8799.n195 20.1342
R14462 a_n6972_8799.n53 a_n6972_8799.n29 75.6825
R14463 a_n6972_8799.n209 a_n6972_8799.n53 9.93802
R14464 a_n6972_8799.n29 a_n6972_8799.n210 161.3
R14465 a_n6972_8799.n74 a_n6972_8799.n18 74.4178
R14466 a_n6972_8799.n218 a_n6972_8799.n74 12.4674
R14467 a_n6972_8799.n73 a_n6972_8799.n18 80.107
R14468 a_n6972_8799.n73 a_n6972_8799.n219 1.08907
R14469 a_n6972_8799.n19 a_n6972_8799.n72 75.3623
R14470 a_n6972_8799.n71 a_n6972_8799.n19 70.3058
R14471 a_n6972_8799.n21 a_n6972_8799.n70 70.1674
R14472 a_n6972_8799.n70 a_n6972_8799.n214 20.9683
R14473 a_n6972_8799.n69 a_n6972_8799.n21 75.0448
R14474 a_n6972_8799.n222 a_n6972_8799.n69 11.2134
R14475 a_n6972_8799.n68 a_n6972_8799.n20 80.4688
R14476 a_n6972_8799.n20 a_n6972_8799.n67 74.73
R14477 a_n6972_8799.n66 a_n6972_8799.n22 70.1674
R14478 a_n6972_8799.n225 a_n6972_8799.n66 20.9683
R14479 a_n6972_8799.n22 a_n6972_8799.n65 70.5844
R14480 a_n6972_8799.n65 a_n6972_8799.n212 20.1342
R14481 a_n6972_8799.n64 a_n6972_8799.n23 75.6825
R14482 a_n6972_8799.n226 a_n6972_8799.n64 9.93802
R14483 a_n6972_8799.n23 a_n6972_8799.n227 161.3
R14484 a_n6972_8799.n13 a_n6972_8799.n85 70.1674
R14485 a_n6972_8799.n144 a_n6972_8799.n85 20.9683
R14486 a_n6972_8799.n84 a_n6972_8799.n13 74.4178
R14487 a_n6972_8799.n84 a_n6972_8799.n129 12.4674
R14488 a_n6972_8799.n12 a_n6972_8799.n83 80.107
R14489 a_n6972_8799.n143 a_n6972_8799.n83 1.08907
R14490 a_n6972_8799.n82 a_n6972_8799.n12 75.3623
R14491 a_n6972_8799.n14 a_n6972_8799.n81 70.3058
R14492 a_n6972_8799.n80 a_n6972_8799.n14 70.1674
R14493 a_n6972_8799.n80 a_n6972_8799.n130 20.9683
R14494 a_n6972_8799.n15 a_n6972_8799.n79 75.0448
R14495 a_n6972_8799.n139 a_n6972_8799.n79 11.2134
R14496 a_n6972_8799.n78 a_n6972_8799.n15 80.4688
R14497 a_n6972_8799.n16 a_n6972_8799.n77 74.73
R14498 a_n6972_8799.n76 a_n6972_8799.n16 70.1674
R14499 a_n6972_8799.n76 a_n6972_8799.n131 20.9683
R14500 a_n6972_8799.n17 a_n6972_8799.n75 70.5844
R14501 a_n6972_8799.n135 a_n6972_8799.n75 20.1342
R14502 a_n6972_8799.n134 a_n6972_8799.n17 161.3
R14503 a_n6972_8799.n7 a_n6972_8799.n96 70.1674
R14504 a_n6972_8799.n160 a_n6972_8799.n96 20.9683
R14505 a_n6972_8799.n95 a_n6972_8799.n7 74.4178
R14506 a_n6972_8799.n95 a_n6972_8799.n145 12.4674
R14507 a_n6972_8799.n6 a_n6972_8799.n94 80.107
R14508 a_n6972_8799.n159 a_n6972_8799.n94 1.08907
R14509 a_n6972_8799.n93 a_n6972_8799.n6 75.3623
R14510 a_n6972_8799.n8 a_n6972_8799.n92 70.3058
R14511 a_n6972_8799.n91 a_n6972_8799.n8 70.1674
R14512 a_n6972_8799.n91 a_n6972_8799.n146 20.9683
R14513 a_n6972_8799.n9 a_n6972_8799.n90 75.0448
R14514 a_n6972_8799.n155 a_n6972_8799.n90 11.2134
R14515 a_n6972_8799.n89 a_n6972_8799.n9 80.4688
R14516 a_n6972_8799.n10 a_n6972_8799.n88 74.73
R14517 a_n6972_8799.n87 a_n6972_8799.n10 70.1674
R14518 a_n6972_8799.n87 a_n6972_8799.n147 20.9683
R14519 a_n6972_8799.n11 a_n6972_8799.n86 70.5844
R14520 a_n6972_8799.n151 a_n6972_8799.n86 20.1342
R14521 a_n6972_8799.n150 a_n6972_8799.n11 161.3
R14522 a_n6972_8799.n1 a_n6972_8799.n107 70.1674
R14523 a_n6972_8799.n177 a_n6972_8799.n107 20.9683
R14524 a_n6972_8799.n106 a_n6972_8799.n1 74.4178
R14525 a_n6972_8799.n106 a_n6972_8799.n162 12.4674
R14526 a_n6972_8799.n0 a_n6972_8799.n105 80.107
R14527 a_n6972_8799.n176 a_n6972_8799.n105 1.08907
R14528 a_n6972_8799.n104 a_n6972_8799.n0 75.3623
R14529 a_n6972_8799.n2 a_n6972_8799.n103 70.3058
R14530 a_n6972_8799.n102 a_n6972_8799.n2 70.1674
R14531 a_n6972_8799.n102 a_n6972_8799.n163 20.9683
R14532 a_n6972_8799.n3 a_n6972_8799.n101 75.0448
R14533 a_n6972_8799.n172 a_n6972_8799.n101 11.2134
R14534 a_n6972_8799.n100 a_n6972_8799.n3 80.4688
R14535 a_n6972_8799.n4 a_n6972_8799.n99 74.73
R14536 a_n6972_8799.n98 a_n6972_8799.n4 70.1674
R14537 a_n6972_8799.n98 a_n6972_8799.n164 20.9683
R14538 a_n6972_8799.n5 a_n6972_8799.n97 70.5844
R14539 a_n6972_8799.n168 a_n6972_8799.n97 20.1342
R14540 a_n6972_8799.n167 a_n6972_8799.n5 161.3
R14541 a_n6972_8799.n37 a_n6972_8799.n108 98.9633
R14542 a_n6972_8799.n36 a_n6972_8799.n109 98.9631
R14543 a_n6972_8799.n37 a_n6972_8799.n232 98.6055
R14544 a_n6972_8799.n36 a_n6972_8799.n110 98.6055
R14545 a_n6972_8799.n36 a_n6972_8799.n111 98.6055
R14546 a_n6972_8799.n233 a_n6972_8799.n37 98.6054
R14547 a_n6972_8799.n114 a_n6972_8799.n112 81.4626
R14548 a_n6972_8799.n122 a_n6972_8799.n120 81.4626
R14549 a_n6972_8799.n118 a_n6972_8799.n116 81.4626
R14550 a_n6972_8799.n125 a_n6972_8799.n124 80.9324
R14551 a_n6972_8799.n127 a_n6972_8799.n126 80.9324
R14552 a_n6972_8799.n41 a_n6972_8799.n128 80.9324
R14553 a_n6972_8799.n40 a_n6972_8799.n115 80.9324
R14554 a_n6972_8799.n114 a_n6972_8799.n113 80.9324
R14555 a_n6972_8799.n122 a_n6972_8799.n121 80.9324
R14556 a_n6972_8799.n39 a_n6972_8799.n123 80.9324
R14557 a_n6972_8799.n38 a_n6972_8799.n119 80.9324
R14558 a_n6972_8799.n118 a_n6972_8799.n117 80.9324
R14559 a_n6972_8799.n30 a_n6972_8799.n184 70.4033
R14560 a_n6972_8799.n24 a_n6972_8799.n200 70.4033
R14561 a_n6972_8799.n18 a_n6972_8799.n217 70.4033
R14562 a_n6972_8799.n17 a_n6972_8799.n133 70.4033
R14563 a_n6972_8799.n11 a_n6972_8799.n149 70.4033
R14564 a_n6972_8799.n5 a_n6972_8799.n166 70.4033
R14565 a_n6972_8799.n194 a_n6972_8799.n193 48.2005
R14566 a_n6972_8799.n44 a_n6972_8799.n191 20.9683
R14567 a_n6972_8799.n190 a_n6972_8799.n189 48.2005
R14568 a_n6972_8799.n188 a_n6972_8799.n48 20.9683
R14569 a_n6972_8799.n186 a_n6972_8799.n182 48.2005
R14570 a_n6972_8799.n210 a_n6972_8799.n209 48.2005
R14571 a_n6972_8799.n55 a_n6972_8799.n207 20.9683
R14572 a_n6972_8799.n206 a_n6972_8799.n205 48.2005
R14573 a_n6972_8799.n204 a_n6972_8799.n59 20.9683
R14574 a_n6972_8799.n202 a_n6972_8799.n198 48.2005
R14575 a_n6972_8799.n227 a_n6972_8799.n226 48.2005
R14576 a_n6972_8799.n66 a_n6972_8799.n224 20.9683
R14577 a_n6972_8799.n223 a_n6972_8799.n222 48.2005
R14578 a_n6972_8799.n221 a_n6972_8799.n70 20.9683
R14579 a_n6972_8799.n219 a_n6972_8799.n215 48.2005
R14580 a_n6972_8799.n136 a_n6972_8799.n76 20.9683
R14581 a_n6972_8799.n139 a_n6972_8799.n138 48.2005
R14582 a_n6972_8799.n140 a_n6972_8799.n80 20.9683
R14583 a_n6972_8799.n143 a_n6972_8799.n142 48.2005
R14584 a_n6972_8799.t45 a_n6972_8799.n85 485.135
R14585 a_n6972_8799.n152 a_n6972_8799.n87 20.9683
R14586 a_n6972_8799.n155 a_n6972_8799.n154 48.2005
R14587 a_n6972_8799.n156 a_n6972_8799.n91 20.9683
R14588 a_n6972_8799.n159 a_n6972_8799.n158 48.2005
R14589 a_n6972_8799.t59 a_n6972_8799.n96 485.135
R14590 a_n6972_8799.n169 a_n6972_8799.n98 20.9683
R14591 a_n6972_8799.n172 a_n6972_8799.n171 48.2005
R14592 a_n6972_8799.n173 a_n6972_8799.n102 20.9683
R14593 a_n6972_8799.n176 a_n6972_8799.n175 48.2005
R14594 a_n6972_8799.t131 a_n6972_8799.n107 485.135
R14595 a_n6972_8799.n46 a_n6972_8799.n180 47.835
R14596 a_n6972_8799.n49 a_n6972_8799.n187 20.6913
R14597 a_n6972_8799.n57 a_n6972_8799.n196 47.835
R14598 a_n6972_8799.n60 a_n6972_8799.n203 20.6913
R14599 a_n6972_8799.n68 a_n6972_8799.n213 47.835
R14600 a_n6972_8799.n71 a_n6972_8799.n220 20.6913
R14601 a_n6972_8799.n137 a_n6972_8799.n78 47.835
R14602 a_n6972_8799.n141 a_n6972_8799.n81 20.6913
R14603 a_n6972_8799.n153 a_n6972_8799.n89 47.835
R14604 a_n6972_8799.n157 a_n6972_8799.n92 20.6913
R14605 a_n6972_8799.n170 a_n6972_8799.n100 47.835
R14606 a_n6972_8799.n174 a_n6972_8799.n103 20.6913
R14607 a_n6972_8799.n192 a_n6972_8799.n43 22.3251
R14608 a_n6972_8799.n208 a_n6972_8799.n54 22.3251
R14609 a_n6972_8799.n225 a_n6972_8799.n65 22.3251
R14610 a_n6972_8799.n131 a_n6972_8799.n75 22.3251
R14611 a_n6972_8799.n147 a_n6972_8799.n86 22.3251
R14612 a_n6972_8799.n164 a_n6972_8799.n97 22.3251
R14613 a_n6972_8799.n125 a_n6972_8799.n39 34.3237
R14614 a_n6972_8799.n52 a_n6972_8799.n183 33.6462
R14615 a_n6972_8799.n63 a_n6972_8799.n199 33.6462
R14616 a_n6972_8799.n74 a_n6972_8799.n216 33.6462
R14617 a_n6972_8799.n135 a_n6972_8799.n134 27.0217
R14618 a_n6972_8799.n144 a_n6972_8799.n84 33.6462
R14619 a_n6972_8799.n151 a_n6972_8799.n150 27.0217
R14620 a_n6972_8799.n160 a_n6972_8799.n95 33.6462
R14621 a_n6972_8799.n168 a_n6972_8799.n167 27.0217
R14622 a_n6972_8799.n177 a_n6972_8799.n106 33.6462
R14623 a_n6972_8799.n45 a_n6972_8799.n180 11.843
R14624 a_n6972_8799.n187 a_n6972_8799.n50 36.139
R14625 a_n6972_8799.n56 a_n6972_8799.n196 11.843
R14626 a_n6972_8799.n203 a_n6972_8799.n61 36.139
R14627 a_n6972_8799.n67 a_n6972_8799.n213 11.843
R14628 a_n6972_8799.n220 a_n6972_8799.n72 36.139
R14629 a_n6972_8799.n137 a_n6972_8799.n77 11.843
R14630 a_n6972_8799.n141 a_n6972_8799.n82 36.139
R14631 a_n6972_8799.n153 a_n6972_8799.n88 11.843
R14632 a_n6972_8799.n157 a_n6972_8799.n93 36.139
R14633 a_n6972_8799.n170 a_n6972_8799.n99 11.843
R14634 a_n6972_8799.n174 a_n6972_8799.n104 36.139
R14635 a_n6972_8799.n47 a_n6972_8799.n181 35.3134
R14636 a_n6972_8799.n58 a_n6972_8799.n197 35.3134
R14637 a_n6972_8799.n69 a_n6972_8799.n214 35.3134
R14638 a_n6972_8799.n130 a_n6972_8799.n79 35.3134
R14639 a_n6972_8799.n146 a_n6972_8799.n90 35.3134
R14640 a_n6972_8799.n163 a_n6972_8799.n101 35.3134
R14641 a_n6972_8799.n191 a_n6972_8799.n45 34.4824
R14642 a_n6972_8799.n50 a_n6972_8799.n182 10.5784
R14643 a_n6972_8799.n207 a_n6972_8799.n56 34.4824
R14644 a_n6972_8799.n61 a_n6972_8799.n198 10.5784
R14645 a_n6972_8799.n224 a_n6972_8799.n67 34.4824
R14646 a_n6972_8799.n72 a_n6972_8799.n215 10.5784
R14647 a_n6972_8799.n77 a_n6972_8799.n136 34.4824
R14648 a_n6972_8799.n142 a_n6972_8799.n82 10.5784
R14649 a_n6972_8799.n88 a_n6972_8799.n152 34.4824
R14650 a_n6972_8799.n158 a_n6972_8799.n93 10.5784
R14651 a_n6972_8799.n99 a_n6972_8799.n169 34.4824
R14652 a_n6972_8799.n175 a_n6972_8799.n104 10.5784
R14653 a_n6972_8799.n42 a_n6972_8799.n179 36.9592
R14654 a_n6972_8799.n53 a_n6972_8799.n195 36.9592
R14655 a_n6972_8799.n64 a_n6972_8799.n212 36.9592
R14656 a_n6972_8799.n134 a_n6972_8799.n132 21.1793
R14657 a_n6972_8799.n150 a_n6972_8799.n148 21.1793
R14658 a_n6972_8799.n167 a_n6972_8799.n165 21.1793
R14659 a_n6972_8799.n184 a_n6972_8799.n183 20.9576
R14660 a_n6972_8799.n200 a_n6972_8799.n199 20.9576
R14661 a_n6972_8799.n217 a_n6972_8799.n216 20.9576
R14662 a_n6972_8799.n133 a_n6972_8799.n132 20.9576
R14663 a_n6972_8799.n149 a_n6972_8799.n148 20.9576
R14664 a_n6972_8799.n166 a_n6972_8799.n165 20.9576
R14665 a_n6972_8799.n230 a_n6972_8799.n41 12.3339
R14666 a_n6972_8799.n231 a_n6972_8799.n230 11.4887
R14667 a_n6972_8799.n211 a_n6972_8799.n35 9.07815
R14668 a_n6972_8799.n161 a_n6972_8799.n13 9.07815
R14669 a_n6972_8799.n229 a_n6972_8799.n178 6.93972
R14670 a_n6972_8799.n229 a_n6972_8799.n228 6.44309
R14671 a_n6972_8799.n211 a_n6972_8799.n29 4.9702
R14672 a_n6972_8799.n228 a_n6972_8799.n23 4.9702
R14673 a_n6972_8799.n161 a_n6972_8799.n7 4.9702
R14674 a_n6972_8799.n178 a_n6972_8799.n1 4.9702
R14675 a_n6972_8799.n228 a_n6972_8799.n211 4.10845
R14676 a_n6972_8799.n178 a_n6972_8799.n161 4.10845
R14677 a_n6972_8799.n232 a_n6972_8799.t14 3.61217
R14678 a_n6972_8799.n232 a_n6972_8799.t21 3.61217
R14679 a_n6972_8799.n108 a_n6972_8799.t3 3.61217
R14680 a_n6972_8799.n108 a_n6972_8799.t9 3.61217
R14681 a_n6972_8799.n109 a_n6972_8799.t4 3.61217
R14682 a_n6972_8799.n109 a_n6972_8799.t13 3.61217
R14683 a_n6972_8799.n110 a_n6972_8799.t12 3.61217
R14684 a_n6972_8799.n110 a_n6972_8799.t22 3.61217
R14685 a_n6972_8799.n111 a_n6972_8799.t7 3.61217
R14686 a_n6972_8799.n111 a_n6972_8799.t8 3.61217
R14687 a_n6972_8799.n233 a_n6972_8799.t18 3.61217
R14688 a_n6972_8799.t2 a_n6972_8799.n233 3.61217
R14689 a_n6972_8799.n230 a_n6972_8799.n229 3.4105
R14690 a_n6972_8799.n124 a_n6972_8799.t19 2.82907
R14691 a_n6972_8799.n124 a_n6972_8799.t10 2.82907
R14692 a_n6972_8799.n126 a_n6972_8799.t26 2.82907
R14693 a_n6972_8799.n126 a_n6972_8799.t25 2.82907
R14694 a_n6972_8799.n128 a_n6972_8799.t31 2.82907
R14695 a_n6972_8799.n128 a_n6972_8799.t23 2.82907
R14696 a_n6972_8799.n115 a_n6972_8799.t35 2.82907
R14697 a_n6972_8799.n115 a_n6972_8799.t0 2.82907
R14698 a_n6972_8799.n113 a_n6972_8799.t28 2.82907
R14699 a_n6972_8799.n113 a_n6972_8799.t30 2.82907
R14700 a_n6972_8799.n112 a_n6972_8799.t15 2.82907
R14701 a_n6972_8799.n112 a_n6972_8799.t20 2.82907
R14702 a_n6972_8799.n120 a_n6972_8799.t17 2.82907
R14703 a_n6972_8799.n120 a_n6972_8799.t33 2.82907
R14704 a_n6972_8799.n121 a_n6972_8799.t34 2.82907
R14705 a_n6972_8799.n121 a_n6972_8799.t6 2.82907
R14706 a_n6972_8799.n123 a_n6972_8799.t24 2.82907
R14707 a_n6972_8799.n123 a_n6972_8799.t27 2.82907
R14708 a_n6972_8799.n119 a_n6972_8799.t32 2.82907
R14709 a_n6972_8799.n119 a_n6972_8799.t5 2.82907
R14710 a_n6972_8799.n117 a_n6972_8799.t11 2.82907
R14711 a_n6972_8799.n117 a_n6972_8799.t16 2.82907
R14712 a_n6972_8799.n116 a_n6972_8799.t1 2.82907
R14713 a_n6972_8799.n116 a_n6972_8799.t29 2.82907
R14714 a_n6972_8799.n51 a_n6972_8799.n185 47.0982
R14715 a_n6972_8799.n62 a_n6972_8799.n201 47.0982
R14716 a_n6972_8799.n73 a_n6972_8799.n218 47.0982
R14717 a_n6972_8799.n129 a_n6972_8799.n83 47.0982
R14718 a_n6972_8799.n145 a_n6972_8799.n94 47.0982
R14719 a_n6972_8799.n162 a_n6972_8799.n105 47.0982
R14720 a_n6972_8799.n231 a_n6972_8799.n36 31.5519
R14721 a_n6972_8799.n46 a_n6972_8799.n190 0.365327
R14722 a_n6972_8799.n188 a_n6972_8799.n49 21.4216
R14723 a_n6972_8799.n57 a_n6972_8799.n206 0.365327
R14724 a_n6972_8799.n204 a_n6972_8799.n60 21.4216
R14725 a_n6972_8799.n68 a_n6972_8799.n223 0.365327
R14726 a_n6972_8799.n221 a_n6972_8799.n71 21.4216
R14727 a_n6972_8799.n138 a_n6972_8799.n78 0.365327
R14728 a_n6972_8799.n81 a_n6972_8799.n140 21.4216
R14729 a_n6972_8799.n154 a_n6972_8799.n89 0.365327
R14730 a_n6972_8799.n92 a_n6972_8799.n156 21.4216
R14731 a_n6972_8799.n171 a_n6972_8799.n100 0.365327
R14732 a_n6972_8799.n103 a_n6972_8799.n173 21.4216
R14733 a_n6972_8799.n37 a_n6972_8799.n231 17.6132
R14734 a_n6972_8799.n31 a_n6972_8799.n30 1.13686
R14735 a_n6972_8799.n25 a_n6972_8799.n24 1.13686
R14736 a_n6972_8799.n19 a_n6972_8799.n18 1.13686
R14737 a_n6972_8799.n13 a_n6972_8799.n12 1.13686
R14738 a_n6972_8799.n7 a_n6972_8799.n6 1.13686
R14739 a_n6972_8799.n1 a_n6972_8799.n0 1.13686
R14740 a_n6972_8799.n35 a_n6972_8799.n34 0.758076
R14741 a_n6972_8799.n32 a_n6972_8799.n34 0.758076
R14742 a_n6972_8799.n33 a_n6972_8799.n32 0.758076
R14743 a_n6972_8799.n33 a_n6972_8799.n31 0.758076
R14744 a_n6972_8799.n29 a_n6972_8799.n28 0.758076
R14745 a_n6972_8799.n26 a_n6972_8799.n28 0.758076
R14746 a_n6972_8799.n27 a_n6972_8799.n26 0.758076
R14747 a_n6972_8799.n27 a_n6972_8799.n25 0.758076
R14748 a_n6972_8799.n23 a_n6972_8799.n22 0.758076
R14749 a_n6972_8799.n20 a_n6972_8799.n22 0.758076
R14750 a_n6972_8799.n21 a_n6972_8799.n20 0.758076
R14751 a_n6972_8799.n21 a_n6972_8799.n19 0.758076
R14752 a_n6972_8799.n16 a_n6972_8799.n17 0.758076
R14753 a_n6972_8799.n15 a_n6972_8799.n16 0.758076
R14754 a_n6972_8799.n14 a_n6972_8799.n15 0.758076
R14755 a_n6972_8799.n12 a_n6972_8799.n14 0.758076
R14756 a_n6972_8799.n10 a_n6972_8799.n11 0.758076
R14757 a_n6972_8799.n9 a_n6972_8799.n10 0.758076
R14758 a_n6972_8799.n8 a_n6972_8799.n9 0.758076
R14759 a_n6972_8799.n6 a_n6972_8799.n8 0.758076
R14760 a_n6972_8799.n4 a_n6972_8799.n5 0.758076
R14761 a_n6972_8799.n3 a_n6972_8799.n4 0.758076
R14762 a_n6972_8799.n2 a_n6972_8799.n3 0.758076
R14763 a_n6972_8799.n0 a_n6972_8799.n2 0.758076
R14764 a_n6972_8799.n38 a_n6972_8799.n118 0.530672
R14765 a_n6972_8799.n39 a_n6972_8799.n122 0.530672
R14766 a_n6972_8799.n40 a_n6972_8799.n114 0.530672
R14767 a_n6972_8799.n41 a_n6972_8799.n127 0.530672
R14768 a_n6972_8799.n127 a_n6972_8799.n125 0.530672
R14769 a_n6972_8799.n41 a_n6972_8799.n40 0.530672
R14770 a_n6972_8799.n39 a_n6972_8799.n38 0.530672
R14771 vdd.n315 vdd.n279 756.745
R14772 vdd.n260 vdd.n224 756.745
R14773 vdd.n217 vdd.n181 756.745
R14774 vdd.n162 vdd.n126 756.745
R14775 vdd.n120 vdd.n84 756.745
R14776 vdd.n65 vdd.n29 756.745
R14777 vdd.n1684 vdd.n1648 756.745
R14778 vdd.n1739 vdd.n1703 756.745
R14779 vdd.n1586 vdd.n1550 756.745
R14780 vdd.n1641 vdd.n1605 756.745
R14781 vdd.n1489 vdd.n1453 756.745
R14782 vdd.n1544 vdd.n1508 756.745
R14783 vdd.n2094 vdd.t230 640.208
R14784 vdd.n936 vdd.t215 640.208
R14785 vdd.n2068 vdd.t253 640.208
R14786 vdd.n928 vdd.t241 640.208
R14787 vdd.n2839 vdd.t202 640.208
R14788 vdd.n2559 vdd.t238 640.208
R14789 vdd.n804 vdd.t219 640.208
R14790 vdd.n2556 vdd.t223 640.208
R14791 vdd.n768 vdd.t227 640.208
R14792 vdd.n998 vdd.t234 640.208
R14793 vdd.n1148 vdd.t184 592.009
R14794 vdd.n1304 vdd.t199 592.009
R14795 vdd.n1340 vdd.t206 592.009
R14796 vdd.n2250 vdd.t195 592.009
R14797 vdd.n1887 vdd.t209 592.009
R14798 vdd.n1847 vdd.t212 592.009
R14799 vdd.n405 vdd.t188 592.009
R14800 vdd.n419 vdd.t244 592.009
R14801 vdd.n431 vdd.t250 592.009
R14802 vdd.n723 vdd.t180 592.009
R14803 vdd.n686 vdd.t192 592.009
R14804 vdd.n3013 vdd.t247 592.009
R14805 vdd.n316 vdd.n315 585
R14806 vdd.n314 vdd.n281 585
R14807 vdd.n313 vdd.n312 585
R14808 vdd.n284 vdd.n282 585
R14809 vdd.n307 vdd.n306 585
R14810 vdd.n305 vdd.n304 585
R14811 vdd.n288 vdd.n287 585
R14812 vdd.n299 vdd.n298 585
R14813 vdd.n297 vdd.n296 585
R14814 vdd.n292 vdd.n291 585
R14815 vdd.n261 vdd.n260 585
R14816 vdd.n259 vdd.n226 585
R14817 vdd.n258 vdd.n257 585
R14818 vdd.n229 vdd.n227 585
R14819 vdd.n252 vdd.n251 585
R14820 vdd.n250 vdd.n249 585
R14821 vdd.n233 vdd.n232 585
R14822 vdd.n244 vdd.n243 585
R14823 vdd.n242 vdd.n241 585
R14824 vdd.n237 vdd.n236 585
R14825 vdd.n218 vdd.n217 585
R14826 vdd.n216 vdd.n183 585
R14827 vdd.n215 vdd.n214 585
R14828 vdd.n186 vdd.n184 585
R14829 vdd.n209 vdd.n208 585
R14830 vdd.n207 vdd.n206 585
R14831 vdd.n190 vdd.n189 585
R14832 vdd.n201 vdd.n200 585
R14833 vdd.n199 vdd.n198 585
R14834 vdd.n194 vdd.n193 585
R14835 vdd.n163 vdd.n162 585
R14836 vdd.n161 vdd.n128 585
R14837 vdd.n160 vdd.n159 585
R14838 vdd.n131 vdd.n129 585
R14839 vdd.n154 vdd.n153 585
R14840 vdd.n152 vdd.n151 585
R14841 vdd.n135 vdd.n134 585
R14842 vdd.n146 vdd.n145 585
R14843 vdd.n144 vdd.n143 585
R14844 vdd.n139 vdd.n138 585
R14845 vdd.n121 vdd.n120 585
R14846 vdd.n119 vdd.n86 585
R14847 vdd.n118 vdd.n117 585
R14848 vdd.n89 vdd.n87 585
R14849 vdd.n112 vdd.n111 585
R14850 vdd.n110 vdd.n109 585
R14851 vdd.n93 vdd.n92 585
R14852 vdd.n104 vdd.n103 585
R14853 vdd.n102 vdd.n101 585
R14854 vdd.n97 vdd.n96 585
R14855 vdd.n66 vdd.n65 585
R14856 vdd.n64 vdd.n31 585
R14857 vdd.n63 vdd.n62 585
R14858 vdd.n34 vdd.n32 585
R14859 vdd.n57 vdd.n56 585
R14860 vdd.n55 vdd.n54 585
R14861 vdd.n38 vdd.n37 585
R14862 vdd.n49 vdd.n48 585
R14863 vdd.n47 vdd.n46 585
R14864 vdd.n42 vdd.n41 585
R14865 vdd.n1685 vdd.n1684 585
R14866 vdd.n1683 vdd.n1650 585
R14867 vdd.n1682 vdd.n1681 585
R14868 vdd.n1653 vdd.n1651 585
R14869 vdd.n1676 vdd.n1675 585
R14870 vdd.n1674 vdd.n1673 585
R14871 vdd.n1657 vdd.n1656 585
R14872 vdd.n1668 vdd.n1667 585
R14873 vdd.n1666 vdd.n1665 585
R14874 vdd.n1661 vdd.n1660 585
R14875 vdd.n1740 vdd.n1739 585
R14876 vdd.n1738 vdd.n1705 585
R14877 vdd.n1737 vdd.n1736 585
R14878 vdd.n1708 vdd.n1706 585
R14879 vdd.n1731 vdd.n1730 585
R14880 vdd.n1729 vdd.n1728 585
R14881 vdd.n1712 vdd.n1711 585
R14882 vdd.n1723 vdd.n1722 585
R14883 vdd.n1721 vdd.n1720 585
R14884 vdd.n1716 vdd.n1715 585
R14885 vdd.n1587 vdd.n1586 585
R14886 vdd.n1585 vdd.n1552 585
R14887 vdd.n1584 vdd.n1583 585
R14888 vdd.n1555 vdd.n1553 585
R14889 vdd.n1578 vdd.n1577 585
R14890 vdd.n1576 vdd.n1575 585
R14891 vdd.n1559 vdd.n1558 585
R14892 vdd.n1570 vdd.n1569 585
R14893 vdd.n1568 vdd.n1567 585
R14894 vdd.n1563 vdd.n1562 585
R14895 vdd.n1642 vdd.n1641 585
R14896 vdd.n1640 vdd.n1607 585
R14897 vdd.n1639 vdd.n1638 585
R14898 vdd.n1610 vdd.n1608 585
R14899 vdd.n1633 vdd.n1632 585
R14900 vdd.n1631 vdd.n1630 585
R14901 vdd.n1614 vdd.n1613 585
R14902 vdd.n1625 vdd.n1624 585
R14903 vdd.n1623 vdd.n1622 585
R14904 vdd.n1618 vdd.n1617 585
R14905 vdd.n1490 vdd.n1489 585
R14906 vdd.n1488 vdd.n1455 585
R14907 vdd.n1487 vdd.n1486 585
R14908 vdd.n1458 vdd.n1456 585
R14909 vdd.n1481 vdd.n1480 585
R14910 vdd.n1479 vdd.n1478 585
R14911 vdd.n1462 vdd.n1461 585
R14912 vdd.n1473 vdd.n1472 585
R14913 vdd.n1471 vdd.n1470 585
R14914 vdd.n1466 vdd.n1465 585
R14915 vdd.n1545 vdd.n1544 585
R14916 vdd.n1543 vdd.n1510 585
R14917 vdd.n1542 vdd.n1541 585
R14918 vdd.n1513 vdd.n1511 585
R14919 vdd.n1536 vdd.n1535 585
R14920 vdd.n1534 vdd.n1533 585
R14921 vdd.n1517 vdd.n1516 585
R14922 vdd.n1528 vdd.n1527 585
R14923 vdd.n1526 vdd.n1525 585
R14924 vdd.n1521 vdd.n1520 585
R14925 vdd.n445 vdd.n370 462.44
R14926 vdd.n3251 vdd.n372 462.44
R14927 vdd.n3146 vdd.n657 462.44
R14928 vdd.n3144 vdd.n660 462.44
R14929 vdd.n2245 vdd.n1047 462.44
R14930 vdd.n2248 vdd.n2247 462.44
R14931 vdd.n1375 vdd.n1145 462.44
R14932 vdd.n1372 vdd.n1143 462.44
R14933 vdd.n293 vdd.t116 329.043
R14934 vdd.n238 vdd.t90 329.043
R14935 vdd.n195 vdd.t102 329.043
R14936 vdd.n140 vdd.t79 329.043
R14937 vdd.n98 vdd.t34 329.043
R14938 vdd.n43 vdd.t14 329.043
R14939 vdd.n1662 vdd.t129 329.043
R14940 vdd.n1717 vdd.t40 329.043
R14941 vdd.n1564 vdd.t114 329.043
R14942 vdd.n1619 vdd.t24 329.043
R14943 vdd.n1467 vdd.t12 329.043
R14944 vdd.n1522 vdd.t37 329.043
R14945 vdd.n1148 vdd.t187 319.788
R14946 vdd.n1304 vdd.t201 319.788
R14947 vdd.n1340 vdd.t208 319.788
R14948 vdd.n2250 vdd.t197 319.788
R14949 vdd.n1887 vdd.t210 319.788
R14950 vdd.n1847 vdd.t213 319.788
R14951 vdd.n405 vdd.t190 319.788
R14952 vdd.n419 vdd.t245 319.788
R14953 vdd.n431 vdd.t251 319.788
R14954 vdd.n723 vdd.t183 319.788
R14955 vdd.n686 vdd.t194 319.788
R14956 vdd.n3013 vdd.t249 319.788
R14957 vdd.n1149 vdd.t186 303.69
R14958 vdd.n1305 vdd.t200 303.69
R14959 vdd.n1341 vdd.t207 303.69
R14960 vdd.n2251 vdd.t198 303.69
R14961 vdd.n1888 vdd.t211 303.69
R14962 vdd.n1848 vdd.t214 303.69
R14963 vdd.n406 vdd.t191 303.69
R14964 vdd.n420 vdd.t246 303.69
R14965 vdd.n432 vdd.t252 303.69
R14966 vdd.n724 vdd.t182 303.69
R14967 vdd.n687 vdd.t193 303.69
R14968 vdd.n3014 vdd.t248 303.69
R14969 vdd.n2782 vdd.n884 297.074
R14970 vdd.n2975 vdd.n778 297.074
R14971 vdd.n2912 vdd.n775 297.074
R14972 vdd.n2705 vdd.n885 297.074
R14973 vdd.n2520 vdd.n925 297.074
R14974 vdd.n2451 vdd.n2450 297.074
R14975 vdd.n2197 vdd.n1021 297.074
R14976 vdd.n2293 vdd.n1019 297.074
R14977 vdd.n2891 vdd.n776 297.074
R14978 vdd.n2978 vdd.n2977 297.074
R14979 vdd.n2554 vdd.n886 297.074
R14980 vdd.n2780 vdd.n887 297.074
R14981 vdd.n2448 vdd.n934 297.074
R14982 vdd.n932 vdd.n907 297.074
R14983 vdd.n2134 vdd.n1022 297.074
R14984 vdd.n2291 vdd.n1023 297.074
R14985 vdd.n2893 vdd.n776 185
R14986 vdd.n2976 vdd.n776 185
R14987 vdd.n2895 vdd.n2894 185
R14988 vdd.n2894 vdd.n774 185
R14989 vdd.n2896 vdd.n810 185
R14990 vdd.n2906 vdd.n810 185
R14991 vdd.n2897 vdd.n819 185
R14992 vdd.n819 vdd.n817 185
R14993 vdd.n2899 vdd.n2898 185
R14994 vdd.n2900 vdd.n2899 185
R14995 vdd.n2852 vdd.n818 185
R14996 vdd.n818 vdd.n814 185
R14997 vdd.n2851 vdd.n2850 185
R14998 vdd.n2850 vdd.n2849 185
R14999 vdd.n821 vdd.n820 185
R15000 vdd.n822 vdd.n821 185
R15001 vdd.n2842 vdd.n2841 185
R15002 vdd.n2843 vdd.n2842 185
R15003 vdd.n2838 vdd.n831 185
R15004 vdd.n831 vdd.n828 185
R15005 vdd.n2837 vdd.n2836 185
R15006 vdd.n2836 vdd.n2835 185
R15007 vdd.n833 vdd.n832 185
R15008 vdd.n841 vdd.n833 185
R15009 vdd.n2828 vdd.n2827 185
R15010 vdd.n2829 vdd.n2828 185
R15011 vdd.n2826 vdd.n842 185
R15012 vdd.n2677 vdd.n842 185
R15013 vdd.n2825 vdd.n2824 185
R15014 vdd.n2824 vdd.n2823 185
R15015 vdd.n844 vdd.n843 185
R15016 vdd.n845 vdd.n844 185
R15017 vdd.n2816 vdd.n2815 185
R15018 vdd.n2817 vdd.n2816 185
R15019 vdd.n2814 vdd.n854 185
R15020 vdd.n854 vdd.n851 185
R15021 vdd.n2813 vdd.n2812 185
R15022 vdd.n2812 vdd.n2811 185
R15023 vdd.n856 vdd.n855 185
R15024 vdd.n864 vdd.n856 185
R15025 vdd.n2804 vdd.n2803 185
R15026 vdd.n2805 vdd.n2804 185
R15027 vdd.n2802 vdd.n865 185
R15028 vdd.n871 vdd.n865 185
R15029 vdd.n2801 vdd.n2800 185
R15030 vdd.n2800 vdd.n2799 185
R15031 vdd.n867 vdd.n866 185
R15032 vdd.n868 vdd.n867 185
R15033 vdd.n2792 vdd.n2791 185
R15034 vdd.n2793 vdd.n2792 185
R15035 vdd.n2790 vdd.n877 185
R15036 vdd.n2698 vdd.n877 185
R15037 vdd.n2789 vdd.n2788 185
R15038 vdd.n2788 vdd.n2787 185
R15039 vdd.n879 vdd.n878 185
R15040 vdd.t256 vdd.n879 185
R15041 vdd.n2780 vdd.n2779 185
R15042 vdd.n2781 vdd.n2780 185
R15043 vdd.n2778 vdd.n887 185
R15044 vdd.n2777 vdd.n2776 185
R15045 vdd.n889 vdd.n888 185
R15046 vdd.n2563 vdd.n2562 185
R15047 vdd.n2565 vdd.n2564 185
R15048 vdd.n2567 vdd.n2566 185
R15049 vdd.n2569 vdd.n2568 185
R15050 vdd.n2571 vdd.n2570 185
R15051 vdd.n2573 vdd.n2572 185
R15052 vdd.n2575 vdd.n2574 185
R15053 vdd.n2577 vdd.n2576 185
R15054 vdd.n2579 vdd.n2578 185
R15055 vdd.n2581 vdd.n2580 185
R15056 vdd.n2583 vdd.n2582 185
R15057 vdd.n2585 vdd.n2584 185
R15058 vdd.n2587 vdd.n2586 185
R15059 vdd.n2589 vdd.n2588 185
R15060 vdd.n2591 vdd.n2590 185
R15061 vdd.n2593 vdd.n2592 185
R15062 vdd.n2595 vdd.n2594 185
R15063 vdd.n2597 vdd.n2596 185
R15064 vdd.n2599 vdd.n2598 185
R15065 vdd.n2601 vdd.n2600 185
R15066 vdd.n2603 vdd.n2602 185
R15067 vdd.n2605 vdd.n2604 185
R15068 vdd.n2607 vdd.n2606 185
R15069 vdd.n2609 vdd.n2608 185
R15070 vdd.n2611 vdd.n2610 185
R15071 vdd.n2613 vdd.n2612 185
R15072 vdd.n2615 vdd.n2614 185
R15073 vdd.n2617 vdd.n2616 185
R15074 vdd.n2619 vdd.n2618 185
R15075 vdd.n2621 vdd.n2620 185
R15076 vdd.n2623 vdd.n2622 185
R15077 vdd.n2624 vdd.n2554 185
R15078 vdd.n2774 vdd.n2554 185
R15079 vdd.n2979 vdd.n2978 185
R15080 vdd.n2980 vdd.n767 185
R15081 vdd.n2982 vdd.n2981 185
R15082 vdd.n2984 vdd.n765 185
R15083 vdd.n2986 vdd.n2985 185
R15084 vdd.n2987 vdd.n764 185
R15085 vdd.n2989 vdd.n2988 185
R15086 vdd.n2991 vdd.n762 185
R15087 vdd.n2993 vdd.n2992 185
R15088 vdd.n2994 vdd.n761 185
R15089 vdd.n2996 vdd.n2995 185
R15090 vdd.n2998 vdd.n759 185
R15091 vdd.n3000 vdd.n2999 185
R15092 vdd.n3001 vdd.n758 185
R15093 vdd.n3003 vdd.n3002 185
R15094 vdd.n3005 vdd.n757 185
R15095 vdd.n3006 vdd.n754 185
R15096 vdd.n3009 vdd.n3008 185
R15097 vdd.n755 vdd.n753 185
R15098 vdd.n2865 vdd.n2864 185
R15099 vdd.n2867 vdd.n2866 185
R15100 vdd.n2869 vdd.n2861 185
R15101 vdd.n2871 vdd.n2870 185
R15102 vdd.n2872 vdd.n2860 185
R15103 vdd.n2874 vdd.n2873 185
R15104 vdd.n2876 vdd.n2858 185
R15105 vdd.n2878 vdd.n2877 185
R15106 vdd.n2879 vdd.n2857 185
R15107 vdd.n2881 vdd.n2880 185
R15108 vdd.n2883 vdd.n2855 185
R15109 vdd.n2885 vdd.n2884 185
R15110 vdd.n2886 vdd.n2854 185
R15111 vdd.n2888 vdd.n2887 185
R15112 vdd.n2890 vdd.n2853 185
R15113 vdd.n2892 vdd.n2891 185
R15114 vdd.n2891 vdd.n756 185
R15115 vdd.n2977 vdd.n771 185
R15116 vdd.n2977 vdd.n2976 185
R15117 vdd.n2629 vdd.n773 185
R15118 vdd.n774 vdd.n773 185
R15119 vdd.n2630 vdd.n809 185
R15120 vdd.n2906 vdd.n809 185
R15121 vdd.n2632 vdd.n2631 185
R15122 vdd.n2631 vdd.n817 185
R15123 vdd.n2633 vdd.n816 185
R15124 vdd.n2900 vdd.n816 185
R15125 vdd.n2635 vdd.n2634 185
R15126 vdd.n2634 vdd.n814 185
R15127 vdd.n2636 vdd.n824 185
R15128 vdd.n2849 vdd.n824 185
R15129 vdd.n2638 vdd.n2637 185
R15130 vdd.n2637 vdd.n822 185
R15131 vdd.n2639 vdd.n830 185
R15132 vdd.n2843 vdd.n830 185
R15133 vdd.n2641 vdd.n2640 185
R15134 vdd.n2640 vdd.n828 185
R15135 vdd.n2642 vdd.n835 185
R15136 vdd.n2835 vdd.n835 185
R15137 vdd.n2644 vdd.n2643 185
R15138 vdd.n2643 vdd.n841 185
R15139 vdd.n2645 vdd.n840 185
R15140 vdd.n2829 vdd.n840 185
R15141 vdd.n2679 vdd.n2678 185
R15142 vdd.n2678 vdd.n2677 185
R15143 vdd.n2680 vdd.n847 185
R15144 vdd.n2823 vdd.n847 185
R15145 vdd.n2682 vdd.n2681 185
R15146 vdd.n2681 vdd.n845 185
R15147 vdd.n2683 vdd.n853 185
R15148 vdd.n2817 vdd.n853 185
R15149 vdd.n2685 vdd.n2684 185
R15150 vdd.n2684 vdd.n851 185
R15151 vdd.n2686 vdd.n858 185
R15152 vdd.n2811 vdd.n858 185
R15153 vdd.n2688 vdd.n2687 185
R15154 vdd.n2687 vdd.n864 185
R15155 vdd.n2689 vdd.n863 185
R15156 vdd.n2805 vdd.n863 185
R15157 vdd.n2691 vdd.n2690 185
R15158 vdd.n2690 vdd.n871 185
R15159 vdd.n2692 vdd.n870 185
R15160 vdd.n2799 vdd.n870 185
R15161 vdd.n2694 vdd.n2693 185
R15162 vdd.n2693 vdd.n868 185
R15163 vdd.n2695 vdd.n876 185
R15164 vdd.n2793 vdd.n876 185
R15165 vdd.n2697 vdd.n2696 185
R15166 vdd.n2698 vdd.n2697 185
R15167 vdd.n2628 vdd.n881 185
R15168 vdd.n2787 vdd.n881 185
R15169 vdd.n2627 vdd.n2626 185
R15170 vdd.n2626 vdd.t256 185
R15171 vdd.n2625 vdd.n886 185
R15172 vdd.n2781 vdd.n886 185
R15173 vdd.n2245 vdd.n2244 185
R15174 vdd.n2246 vdd.n2245 185
R15175 vdd.n1048 vdd.n1046 185
R15176 vdd.n1046 vdd.n1044 185
R15177 vdd.n1814 vdd.n1813 185
R15178 vdd.n1813 vdd.n1812 185
R15179 vdd.n1051 vdd.n1050 185
R15180 vdd.n1052 vdd.n1051 185
R15181 vdd.n1801 vdd.n1800 185
R15182 vdd.n1802 vdd.n1801 185
R15183 vdd.n1060 vdd.n1059 185
R15184 vdd.n1793 vdd.n1059 185
R15185 vdd.n1796 vdd.n1795 185
R15186 vdd.n1795 vdd.n1794 185
R15187 vdd.n1063 vdd.n1062 185
R15188 vdd.n1069 vdd.n1063 185
R15189 vdd.n1784 vdd.n1783 185
R15190 vdd.n1785 vdd.n1784 185
R15191 vdd.n1071 vdd.n1070 185
R15192 vdd.n1776 vdd.n1070 185
R15193 vdd.n1779 vdd.n1778 185
R15194 vdd.n1778 vdd.n1777 185
R15195 vdd.n1074 vdd.n1073 185
R15196 vdd.n1075 vdd.n1074 185
R15197 vdd.n1767 vdd.n1766 185
R15198 vdd.n1768 vdd.n1767 185
R15199 vdd.n1083 vdd.n1082 185
R15200 vdd.n1082 vdd.n1081 185
R15201 vdd.n1762 vdd.n1761 185
R15202 vdd.n1761 vdd.n1760 185
R15203 vdd.n1086 vdd.n1085 185
R15204 vdd.n1092 vdd.n1086 185
R15205 vdd.n1751 vdd.n1750 185
R15206 vdd.n1752 vdd.n1751 185
R15207 vdd.n1094 vdd.n1093 185
R15208 vdd.n1448 vdd.n1093 185
R15209 vdd.n1451 vdd.n1450 185
R15210 vdd.n1450 vdd.n1449 185
R15211 vdd.n1097 vdd.n1096 185
R15212 vdd.n1104 vdd.n1097 185
R15213 vdd.n1439 vdd.n1438 185
R15214 vdd.n1440 vdd.n1439 185
R15215 vdd.n1106 vdd.n1105 185
R15216 vdd.n1105 vdd.n1103 185
R15217 vdd.n1434 vdd.n1433 185
R15218 vdd.n1433 vdd.n1432 185
R15219 vdd.n1109 vdd.n1108 185
R15220 vdd.n1110 vdd.n1109 185
R15221 vdd.n1423 vdd.n1422 185
R15222 vdd.n1424 vdd.n1423 185
R15223 vdd.n1117 vdd.n1116 185
R15224 vdd.n1415 vdd.n1116 185
R15225 vdd.n1418 vdd.n1417 185
R15226 vdd.n1417 vdd.n1416 185
R15227 vdd.n1120 vdd.n1119 185
R15228 vdd.n1126 vdd.n1120 185
R15229 vdd.n1406 vdd.n1405 185
R15230 vdd.n1407 vdd.n1406 185
R15231 vdd.n1128 vdd.n1127 185
R15232 vdd.n1398 vdd.n1127 185
R15233 vdd.n1401 vdd.n1400 185
R15234 vdd.n1400 vdd.n1399 185
R15235 vdd.n1131 vdd.n1130 185
R15236 vdd.n1132 vdd.n1131 185
R15237 vdd.n1389 vdd.n1388 185
R15238 vdd.n1390 vdd.n1389 185
R15239 vdd.n1140 vdd.n1139 185
R15240 vdd.n1139 vdd.n1138 185
R15241 vdd.n1384 vdd.n1383 185
R15242 vdd.n1383 vdd.n1382 185
R15243 vdd.n1143 vdd.n1142 185
R15244 vdd.n1144 vdd.n1143 185
R15245 vdd.n1372 vdd.n1371 185
R15246 vdd.n1370 vdd.n1183 185
R15247 vdd.n1185 vdd.n1182 185
R15248 vdd.n1374 vdd.n1182 185
R15249 vdd.n1366 vdd.n1187 185
R15250 vdd.n1365 vdd.n1188 185
R15251 vdd.n1364 vdd.n1189 185
R15252 vdd.n1192 vdd.n1190 185
R15253 vdd.n1360 vdd.n1193 185
R15254 vdd.n1359 vdd.n1194 185
R15255 vdd.n1358 vdd.n1195 185
R15256 vdd.n1198 vdd.n1196 185
R15257 vdd.n1354 vdd.n1199 185
R15258 vdd.n1353 vdd.n1200 185
R15259 vdd.n1352 vdd.n1201 185
R15260 vdd.n1204 vdd.n1202 185
R15261 vdd.n1348 vdd.n1205 185
R15262 vdd.n1347 vdd.n1206 185
R15263 vdd.n1346 vdd.n1207 185
R15264 vdd.n1338 vdd.n1208 185
R15265 vdd.n1342 vdd.n1339 185
R15266 vdd.n1337 vdd.n1210 185
R15267 vdd.n1336 vdd.n1211 185
R15268 vdd.n1214 vdd.n1212 185
R15269 vdd.n1332 vdd.n1215 185
R15270 vdd.n1331 vdd.n1216 185
R15271 vdd.n1330 vdd.n1217 185
R15272 vdd.n1220 vdd.n1218 185
R15273 vdd.n1326 vdd.n1221 185
R15274 vdd.n1325 vdd.n1222 185
R15275 vdd.n1324 vdd.n1223 185
R15276 vdd.n1226 vdd.n1224 185
R15277 vdd.n1320 vdd.n1227 185
R15278 vdd.n1319 vdd.n1228 185
R15279 vdd.n1318 vdd.n1229 185
R15280 vdd.n1232 vdd.n1230 185
R15281 vdd.n1314 vdd.n1233 185
R15282 vdd.n1313 vdd.n1234 185
R15283 vdd.n1312 vdd.n1235 185
R15284 vdd.n1238 vdd.n1236 185
R15285 vdd.n1308 vdd.n1239 185
R15286 vdd.n1307 vdd.n1240 185
R15287 vdd.n1306 vdd.n1303 185
R15288 vdd.n1243 vdd.n1241 185
R15289 vdd.n1299 vdd.n1244 185
R15290 vdd.n1298 vdd.n1245 185
R15291 vdd.n1297 vdd.n1246 185
R15292 vdd.n1249 vdd.n1247 185
R15293 vdd.n1293 vdd.n1250 185
R15294 vdd.n1292 vdd.n1251 185
R15295 vdd.n1291 vdd.n1252 185
R15296 vdd.n1255 vdd.n1253 185
R15297 vdd.n1287 vdd.n1256 185
R15298 vdd.n1286 vdd.n1257 185
R15299 vdd.n1285 vdd.n1258 185
R15300 vdd.n1261 vdd.n1259 185
R15301 vdd.n1281 vdd.n1262 185
R15302 vdd.n1280 vdd.n1263 185
R15303 vdd.n1279 vdd.n1264 185
R15304 vdd.n1267 vdd.n1265 185
R15305 vdd.n1275 vdd.n1268 185
R15306 vdd.n1274 vdd.n1269 185
R15307 vdd.n1273 vdd.n1270 185
R15308 vdd.n1271 vdd.n1151 185
R15309 vdd.n1376 vdd.n1375 185
R15310 vdd.n1375 vdd.n1374 185
R15311 vdd.n2249 vdd.n2248 185
R15312 vdd.n2253 vdd.n1040 185
R15313 vdd.n1916 vdd.n1039 185
R15314 vdd.n1919 vdd.n1918 185
R15315 vdd.n1921 vdd.n1920 185
R15316 vdd.n1924 vdd.n1923 185
R15317 vdd.n1926 vdd.n1925 185
R15318 vdd.n1928 vdd.n1914 185
R15319 vdd.n1930 vdd.n1929 185
R15320 vdd.n1931 vdd.n1908 185
R15321 vdd.n1933 vdd.n1932 185
R15322 vdd.n1935 vdd.n1906 185
R15323 vdd.n1937 vdd.n1936 185
R15324 vdd.n1938 vdd.n1901 185
R15325 vdd.n1940 vdd.n1939 185
R15326 vdd.n1942 vdd.n1899 185
R15327 vdd.n1944 vdd.n1943 185
R15328 vdd.n1945 vdd.n1895 185
R15329 vdd.n1947 vdd.n1946 185
R15330 vdd.n1949 vdd.n1892 185
R15331 vdd.n1951 vdd.n1950 185
R15332 vdd.n1893 vdd.n1886 185
R15333 vdd.n1955 vdd.n1890 185
R15334 vdd.n1956 vdd.n1882 185
R15335 vdd.n1958 vdd.n1957 185
R15336 vdd.n1960 vdd.n1880 185
R15337 vdd.n1962 vdd.n1961 185
R15338 vdd.n1963 vdd.n1875 185
R15339 vdd.n1965 vdd.n1964 185
R15340 vdd.n1967 vdd.n1873 185
R15341 vdd.n1969 vdd.n1968 185
R15342 vdd.n1970 vdd.n1868 185
R15343 vdd.n1972 vdd.n1971 185
R15344 vdd.n1974 vdd.n1866 185
R15345 vdd.n1976 vdd.n1975 185
R15346 vdd.n1977 vdd.n1861 185
R15347 vdd.n1979 vdd.n1978 185
R15348 vdd.n1981 vdd.n1859 185
R15349 vdd.n1983 vdd.n1982 185
R15350 vdd.n1984 vdd.n1855 185
R15351 vdd.n1986 vdd.n1985 185
R15352 vdd.n1988 vdd.n1852 185
R15353 vdd.n1990 vdd.n1989 185
R15354 vdd.n1853 vdd.n1846 185
R15355 vdd.n1994 vdd.n1850 185
R15356 vdd.n1995 vdd.n1842 185
R15357 vdd.n1997 vdd.n1996 185
R15358 vdd.n1999 vdd.n1840 185
R15359 vdd.n2001 vdd.n2000 185
R15360 vdd.n2002 vdd.n1835 185
R15361 vdd.n2004 vdd.n2003 185
R15362 vdd.n2006 vdd.n1833 185
R15363 vdd.n2008 vdd.n2007 185
R15364 vdd.n2009 vdd.n1828 185
R15365 vdd.n2011 vdd.n2010 185
R15366 vdd.n2013 vdd.n1827 185
R15367 vdd.n2014 vdd.n1824 185
R15368 vdd.n2017 vdd.n2016 185
R15369 vdd.n1826 vdd.n1822 185
R15370 vdd.n2234 vdd.n1820 185
R15371 vdd.n2236 vdd.n2235 185
R15372 vdd.n2238 vdd.n1818 185
R15373 vdd.n2240 vdd.n2239 185
R15374 vdd.n2241 vdd.n1047 185
R15375 vdd.n2247 vdd.n1043 185
R15376 vdd.n2247 vdd.n2246 185
R15377 vdd.n1055 vdd.n1042 185
R15378 vdd.n1044 vdd.n1042 185
R15379 vdd.n1811 vdd.n1810 185
R15380 vdd.n1812 vdd.n1811 185
R15381 vdd.n1054 vdd.n1053 185
R15382 vdd.n1053 vdd.n1052 185
R15383 vdd.n1804 vdd.n1803 185
R15384 vdd.n1803 vdd.n1802 185
R15385 vdd.n1058 vdd.n1057 185
R15386 vdd.n1793 vdd.n1058 185
R15387 vdd.n1792 vdd.n1791 185
R15388 vdd.n1794 vdd.n1792 185
R15389 vdd.n1065 vdd.n1064 185
R15390 vdd.n1069 vdd.n1064 185
R15391 vdd.n1787 vdd.n1786 185
R15392 vdd.n1786 vdd.n1785 185
R15393 vdd.n1068 vdd.n1067 185
R15394 vdd.n1776 vdd.n1068 185
R15395 vdd.n1775 vdd.n1774 185
R15396 vdd.n1777 vdd.n1775 185
R15397 vdd.n1077 vdd.n1076 185
R15398 vdd.n1076 vdd.n1075 185
R15399 vdd.n1770 vdd.n1769 185
R15400 vdd.n1769 vdd.n1768 185
R15401 vdd.n1080 vdd.n1079 185
R15402 vdd.n1081 vdd.n1080 185
R15403 vdd.n1759 vdd.n1758 185
R15404 vdd.n1760 vdd.n1759 185
R15405 vdd.n1088 vdd.n1087 185
R15406 vdd.n1092 vdd.n1087 185
R15407 vdd.n1754 vdd.n1753 185
R15408 vdd.n1753 vdd.n1752 185
R15409 vdd.n1091 vdd.n1090 185
R15410 vdd.n1448 vdd.n1091 185
R15411 vdd.n1447 vdd.n1446 185
R15412 vdd.n1449 vdd.n1447 185
R15413 vdd.n1099 vdd.n1098 185
R15414 vdd.n1104 vdd.n1098 185
R15415 vdd.n1442 vdd.n1441 185
R15416 vdd.n1441 vdd.n1440 185
R15417 vdd.n1102 vdd.n1101 185
R15418 vdd.n1103 vdd.n1102 185
R15419 vdd.n1431 vdd.n1430 185
R15420 vdd.n1432 vdd.n1431 185
R15421 vdd.n1112 vdd.n1111 185
R15422 vdd.n1111 vdd.n1110 185
R15423 vdd.n1426 vdd.n1425 185
R15424 vdd.n1425 vdd.n1424 185
R15425 vdd.n1115 vdd.n1114 185
R15426 vdd.n1415 vdd.n1115 185
R15427 vdd.n1414 vdd.n1413 185
R15428 vdd.n1416 vdd.n1414 185
R15429 vdd.n1122 vdd.n1121 185
R15430 vdd.n1126 vdd.n1121 185
R15431 vdd.n1409 vdd.n1408 185
R15432 vdd.n1408 vdd.n1407 185
R15433 vdd.n1125 vdd.n1124 185
R15434 vdd.n1398 vdd.n1125 185
R15435 vdd.n1397 vdd.n1396 185
R15436 vdd.n1399 vdd.n1397 185
R15437 vdd.n1134 vdd.n1133 185
R15438 vdd.n1133 vdd.n1132 185
R15439 vdd.n1392 vdd.n1391 185
R15440 vdd.n1391 vdd.n1390 185
R15441 vdd.n1137 vdd.n1136 185
R15442 vdd.n1138 vdd.n1137 185
R15443 vdd.n1381 vdd.n1380 185
R15444 vdd.n1382 vdd.n1381 185
R15445 vdd.n1146 vdd.n1145 185
R15446 vdd.n1145 vdd.n1144 185
R15447 vdd.n927 vdd.n925 185
R15448 vdd.n2449 vdd.n925 185
R15449 vdd.n2371 vdd.n944 185
R15450 vdd.n944 vdd.t1 185
R15451 vdd.n2373 vdd.n2372 185
R15452 vdd.n2374 vdd.n2373 185
R15453 vdd.n2370 vdd.n943 185
R15454 vdd.n2073 vdd.n943 185
R15455 vdd.n2369 vdd.n2368 185
R15456 vdd.n2368 vdd.n2367 185
R15457 vdd.n946 vdd.n945 185
R15458 vdd.n947 vdd.n946 185
R15459 vdd.n2358 vdd.n2357 185
R15460 vdd.n2359 vdd.n2358 185
R15461 vdd.n2356 vdd.n957 185
R15462 vdd.n957 vdd.n954 185
R15463 vdd.n2355 vdd.n2354 185
R15464 vdd.n2354 vdd.n2353 185
R15465 vdd.n959 vdd.n958 185
R15466 vdd.n960 vdd.n959 185
R15467 vdd.n2346 vdd.n2345 185
R15468 vdd.n2347 vdd.n2346 185
R15469 vdd.n2344 vdd.n968 185
R15470 vdd.n973 vdd.n968 185
R15471 vdd.n2343 vdd.n2342 185
R15472 vdd.n2342 vdd.n2341 185
R15473 vdd.n970 vdd.n969 185
R15474 vdd.n979 vdd.n970 185
R15475 vdd.n2334 vdd.n2333 185
R15476 vdd.n2335 vdd.n2334 185
R15477 vdd.n2332 vdd.n980 185
R15478 vdd.n2174 vdd.n980 185
R15479 vdd.n2331 vdd.n2330 185
R15480 vdd.n2330 vdd.n2329 185
R15481 vdd.n982 vdd.n981 185
R15482 vdd.n983 vdd.n982 185
R15483 vdd.n2322 vdd.n2321 185
R15484 vdd.n2323 vdd.n2322 185
R15485 vdd.n2320 vdd.n992 185
R15486 vdd.n992 vdd.n989 185
R15487 vdd.n2319 vdd.n2318 185
R15488 vdd.n2318 vdd.n2317 185
R15489 vdd.n994 vdd.n993 185
R15490 vdd.n1004 vdd.n994 185
R15491 vdd.n2309 vdd.n2308 185
R15492 vdd.n2310 vdd.n2309 185
R15493 vdd.n2307 vdd.n1005 185
R15494 vdd.n1005 vdd.n1001 185
R15495 vdd.n2306 vdd.n2305 185
R15496 vdd.n2305 vdd.n2304 185
R15497 vdd.n1007 vdd.n1006 185
R15498 vdd.n1008 vdd.n1007 185
R15499 vdd.n2297 vdd.n2296 185
R15500 vdd.n2298 vdd.n2297 185
R15501 vdd.n2295 vdd.n1017 185
R15502 vdd.n1017 vdd.n1014 185
R15503 vdd.n2294 vdd.n2293 185
R15504 vdd.n2293 vdd.n2292 185
R15505 vdd.n1019 vdd.n1018 185
R15506 vdd.n2029 vdd.n2028 185
R15507 vdd.n2030 vdd.n2026 185
R15508 vdd.n2026 vdd.n1020 185
R15509 vdd.n2032 vdd.n2031 185
R15510 vdd.n2034 vdd.n2025 185
R15511 vdd.n2037 vdd.n2036 185
R15512 vdd.n2038 vdd.n2024 185
R15513 vdd.n2040 vdd.n2039 185
R15514 vdd.n2042 vdd.n2023 185
R15515 vdd.n2045 vdd.n2044 185
R15516 vdd.n2046 vdd.n2022 185
R15517 vdd.n2048 vdd.n2047 185
R15518 vdd.n2050 vdd.n2021 185
R15519 vdd.n2053 vdd.n2052 185
R15520 vdd.n2054 vdd.n2020 185
R15521 vdd.n2056 vdd.n2055 185
R15522 vdd.n2058 vdd.n2019 185
R15523 vdd.n2231 vdd.n2059 185
R15524 vdd.n2230 vdd.n2229 185
R15525 vdd.n2227 vdd.n2060 185
R15526 vdd.n2225 vdd.n2224 185
R15527 vdd.n2223 vdd.n2061 185
R15528 vdd.n2222 vdd.n2221 185
R15529 vdd.n2219 vdd.n2062 185
R15530 vdd.n2217 vdd.n2216 185
R15531 vdd.n2215 vdd.n2063 185
R15532 vdd.n2214 vdd.n2213 185
R15533 vdd.n2211 vdd.n2064 185
R15534 vdd.n2209 vdd.n2208 185
R15535 vdd.n2207 vdd.n2065 185
R15536 vdd.n2206 vdd.n2205 185
R15537 vdd.n2203 vdd.n2066 185
R15538 vdd.n2201 vdd.n2200 185
R15539 vdd.n2199 vdd.n2067 185
R15540 vdd.n2198 vdd.n2197 185
R15541 vdd.n2452 vdd.n2451 185
R15542 vdd.n2454 vdd.n2453 185
R15543 vdd.n2456 vdd.n2455 185
R15544 vdd.n2459 vdd.n2458 185
R15545 vdd.n2461 vdd.n2460 185
R15546 vdd.n2463 vdd.n2462 185
R15547 vdd.n2465 vdd.n2464 185
R15548 vdd.n2467 vdd.n2466 185
R15549 vdd.n2469 vdd.n2468 185
R15550 vdd.n2471 vdd.n2470 185
R15551 vdd.n2473 vdd.n2472 185
R15552 vdd.n2475 vdd.n2474 185
R15553 vdd.n2477 vdd.n2476 185
R15554 vdd.n2479 vdd.n2478 185
R15555 vdd.n2481 vdd.n2480 185
R15556 vdd.n2483 vdd.n2482 185
R15557 vdd.n2485 vdd.n2484 185
R15558 vdd.n2487 vdd.n2486 185
R15559 vdd.n2489 vdd.n2488 185
R15560 vdd.n2491 vdd.n2490 185
R15561 vdd.n2493 vdd.n2492 185
R15562 vdd.n2495 vdd.n2494 185
R15563 vdd.n2497 vdd.n2496 185
R15564 vdd.n2499 vdd.n2498 185
R15565 vdd.n2501 vdd.n2500 185
R15566 vdd.n2503 vdd.n2502 185
R15567 vdd.n2505 vdd.n2504 185
R15568 vdd.n2507 vdd.n2506 185
R15569 vdd.n2509 vdd.n2508 185
R15570 vdd.n2511 vdd.n2510 185
R15571 vdd.n2513 vdd.n2512 185
R15572 vdd.n2515 vdd.n2514 185
R15573 vdd.n2517 vdd.n2516 185
R15574 vdd.n2518 vdd.n926 185
R15575 vdd.n2520 vdd.n2519 185
R15576 vdd.n2521 vdd.n2520 185
R15577 vdd.n2450 vdd.n930 185
R15578 vdd.n2450 vdd.n2449 185
R15579 vdd.n2071 vdd.n931 185
R15580 vdd.t1 vdd.n931 185
R15581 vdd.n2072 vdd.n941 185
R15582 vdd.n2374 vdd.n941 185
R15583 vdd.n2075 vdd.n2074 185
R15584 vdd.n2074 vdd.n2073 185
R15585 vdd.n2076 vdd.n948 185
R15586 vdd.n2367 vdd.n948 185
R15587 vdd.n2078 vdd.n2077 185
R15588 vdd.n2077 vdd.n947 185
R15589 vdd.n2079 vdd.n955 185
R15590 vdd.n2359 vdd.n955 185
R15591 vdd.n2081 vdd.n2080 185
R15592 vdd.n2080 vdd.n954 185
R15593 vdd.n2082 vdd.n961 185
R15594 vdd.n2353 vdd.n961 185
R15595 vdd.n2084 vdd.n2083 185
R15596 vdd.n2083 vdd.n960 185
R15597 vdd.n2085 vdd.n966 185
R15598 vdd.n2347 vdd.n966 185
R15599 vdd.n2087 vdd.n2086 185
R15600 vdd.n2086 vdd.n973 185
R15601 vdd.n2088 vdd.n971 185
R15602 vdd.n2341 vdd.n971 185
R15603 vdd.n2090 vdd.n2089 185
R15604 vdd.n2089 vdd.n979 185
R15605 vdd.n2091 vdd.n977 185
R15606 vdd.n2335 vdd.n977 185
R15607 vdd.n2176 vdd.n2175 185
R15608 vdd.n2175 vdd.n2174 185
R15609 vdd.n2177 vdd.n984 185
R15610 vdd.n2329 vdd.n984 185
R15611 vdd.n2179 vdd.n2178 185
R15612 vdd.n2178 vdd.n983 185
R15613 vdd.n2180 vdd.n990 185
R15614 vdd.n2323 vdd.n990 185
R15615 vdd.n2182 vdd.n2181 185
R15616 vdd.n2181 vdd.n989 185
R15617 vdd.n2183 vdd.n995 185
R15618 vdd.n2317 vdd.n995 185
R15619 vdd.n2185 vdd.n2184 185
R15620 vdd.n2184 vdd.n1004 185
R15621 vdd.n2186 vdd.n1002 185
R15622 vdd.n2310 vdd.n1002 185
R15623 vdd.n2188 vdd.n2187 185
R15624 vdd.n2187 vdd.n1001 185
R15625 vdd.n2189 vdd.n1009 185
R15626 vdd.n2304 vdd.n1009 185
R15627 vdd.n2191 vdd.n2190 185
R15628 vdd.n2190 vdd.n1008 185
R15629 vdd.n2192 vdd.n1015 185
R15630 vdd.n2298 vdd.n1015 185
R15631 vdd.n2194 vdd.n2193 185
R15632 vdd.n2193 vdd.n1014 185
R15633 vdd.n2195 vdd.n1021 185
R15634 vdd.n2292 vdd.n1021 185
R15635 vdd.n370 vdd.n369 185
R15636 vdd.n3254 vdd.n370 185
R15637 vdd.n3257 vdd.n3256 185
R15638 vdd.n3256 vdd.n3255 185
R15639 vdd.n3258 vdd.n364 185
R15640 vdd.n364 vdd.n363 185
R15641 vdd.n3260 vdd.n3259 185
R15642 vdd.n3261 vdd.n3260 185
R15643 vdd.n359 vdd.n358 185
R15644 vdd.n3262 vdd.n359 185
R15645 vdd.n3265 vdd.n3264 185
R15646 vdd.n3264 vdd.n3263 185
R15647 vdd.n3266 vdd.n353 185
R15648 vdd.n3236 vdd.n353 185
R15649 vdd.n3268 vdd.n3267 185
R15650 vdd.n3269 vdd.n3268 185
R15651 vdd.n348 vdd.n347 185
R15652 vdd.n3270 vdd.n348 185
R15653 vdd.n3273 vdd.n3272 185
R15654 vdd.n3272 vdd.n3271 185
R15655 vdd.n3274 vdd.n342 185
R15656 vdd.n349 vdd.n342 185
R15657 vdd.n3276 vdd.n3275 185
R15658 vdd.n3277 vdd.n3276 185
R15659 vdd.n338 vdd.n337 185
R15660 vdd.n3278 vdd.n338 185
R15661 vdd.n3281 vdd.n3280 185
R15662 vdd.n3280 vdd.n3279 185
R15663 vdd.n3282 vdd.n333 185
R15664 vdd.n333 vdd.n332 185
R15665 vdd.n3284 vdd.n3283 185
R15666 vdd.n3285 vdd.n3284 185
R15667 vdd.n327 vdd.n325 185
R15668 vdd.n3286 vdd.n327 185
R15669 vdd.n3289 vdd.n3288 185
R15670 vdd.n3288 vdd.n3287 185
R15671 vdd.n326 vdd.n324 185
R15672 vdd.n328 vdd.n326 185
R15673 vdd.n3212 vdd.n3211 185
R15674 vdd.n3213 vdd.n3212 185
R15675 vdd.n615 vdd.n614 185
R15676 vdd.n614 vdd.n613 185
R15677 vdd.n3207 vdd.n3206 185
R15678 vdd.n3206 vdd.n3205 185
R15679 vdd.n618 vdd.n617 185
R15680 vdd.n624 vdd.n618 185
R15681 vdd.n3193 vdd.n3192 185
R15682 vdd.n3194 vdd.n3193 185
R15683 vdd.n626 vdd.n625 185
R15684 vdd.n3185 vdd.n625 185
R15685 vdd.n3188 vdd.n3187 185
R15686 vdd.n3187 vdd.n3186 185
R15687 vdd.n629 vdd.n628 185
R15688 vdd.n636 vdd.n629 185
R15689 vdd.n3176 vdd.n3175 185
R15690 vdd.n3177 vdd.n3176 185
R15691 vdd.n638 vdd.n637 185
R15692 vdd.n637 vdd.n635 185
R15693 vdd.n3171 vdd.n3170 185
R15694 vdd.n3170 vdd.n3169 185
R15695 vdd.n641 vdd.n640 185
R15696 vdd.n642 vdd.n641 185
R15697 vdd.n3160 vdd.n3159 185
R15698 vdd.n3161 vdd.n3160 185
R15699 vdd.n650 vdd.n649 185
R15700 vdd.n649 vdd.n648 185
R15701 vdd.n3155 vdd.n3154 185
R15702 vdd.n3154 vdd.n3153 185
R15703 vdd.n653 vdd.n652 185
R15704 vdd.n659 vdd.n653 185
R15705 vdd.n3144 vdd.n3143 185
R15706 vdd.n3145 vdd.n3144 185
R15707 vdd.n3140 vdd.n660 185
R15708 vdd.n3139 vdd.n3138 185
R15709 vdd.n3136 vdd.n662 185
R15710 vdd.n3136 vdd.n658 185
R15711 vdd.n3135 vdd.n3134 185
R15712 vdd.n3133 vdd.n3132 185
R15713 vdd.n3131 vdd.n3130 185
R15714 vdd.n3129 vdd.n3128 185
R15715 vdd.n3127 vdd.n668 185
R15716 vdd.n3125 vdd.n3124 185
R15717 vdd.n3123 vdd.n669 185
R15718 vdd.n3122 vdd.n3121 185
R15719 vdd.n3119 vdd.n674 185
R15720 vdd.n3117 vdd.n3116 185
R15721 vdd.n3115 vdd.n675 185
R15722 vdd.n3114 vdd.n3113 185
R15723 vdd.n3111 vdd.n680 185
R15724 vdd.n3109 vdd.n3108 185
R15725 vdd.n3107 vdd.n681 185
R15726 vdd.n3106 vdd.n3105 185
R15727 vdd.n3103 vdd.n688 185
R15728 vdd.n3101 vdd.n3100 185
R15729 vdd.n3099 vdd.n689 185
R15730 vdd.n3098 vdd.n3097 185
R15731 vdd.n3095 vdd.n694 185
R15732 vdd.n3093 vdd.n3092 185
R15733 vdd.n3091 vdd.n695 185
R15734 vdd.n3090 vdd.n3089 185
R15735 vdd.n3087 vdd.n700 185
R15736 vdd.n3085 vdd.n3084 185
R15737 vdd.n3083 vdd.n701 185
R15738 vdd.n3082 vdd.n3081 185
R15739 vdd.n3079 vdd.n706 185
R15740 vdd.n3077 vdd.n3076 185
R15741 vdd.n3075 vdd.n707 185
R15742 vdd.n3074 vdd.n3073 185
R15743 vdd.n3071 vdd.n712 185
R15744 vdd.n3069 vdd.n3068 185
R15745 vdd.n3067 vdd.n713 185
R15746 vdd.n3066 vdd.n3065 185
R15747 vdd.n3063 vdd.n718 185
R15748 vdd.n3061 vdd.n3060 185
R15749 vdd.n3059 vdd.n719 185
R15750 vdd.n728 vdd.n722 185
R15751 vdd.n3055 vdd.n3054 185
R15752 vdd.n3052 vdd.n726 185
R15753 vdd.n3051 vdd.n3050 185
R15754 vdd.n3049 vdd.n3048 185
R15755 vdd.n3047 vdd.n732 185
R15756 vdd.n3045 vdd.n3044 185
R15757 vdd.n3043 vdd.n733 185
R15758 vdd.n3042 vdd.n3041 185
R15759 vdd.n3039 vdd.n738 185
R15760 vdd.n3037 vdd.n3036 185
R15761 vdd.n3035 vdd.n739 185
R15762 vdd.n3034 vdd.n3033 185
R15763 vdd.n3031 vdd.n744 185
R15764 vdd.n3029 vdd.n3028 185
R15765 vdd.n3027 vdd.n745 185
R15766 vdd.n3026 vdd.n3025 185
R15767 vdd.n3023 vdd.n3022 185
R15768 vdd.n3021 vdd.n3020 185
R15769 vdd.n3019 vdd.n3018 185
R15770 vdd.n3017 vdd.n3016 185
R15771 vdd.n3012 vdd.n657 185
R15772 vdd.n658 vdd.n657 185
R15773 vdd.n3251 vdd.n3250 185
R15774 vdd.n599 vdd.n404 185
R15775 vdd.n598 vdd.n597 185
R15776 vdd.n596 vdd.n595 185
R15777 vdd.n594 vdd.n409 185
R15778 vdd.n590 vdd.n589 185
R15779 vdd.n588 vdd.n587 185
R15780 vdd.n586 vdd.n585 185
R15781 vdd.n584 vdd.n411 185
R15782 vdd.n580 vdd.n579 185
R15783 vdd.n578 vdd.n577 185
R15784 vdd.n576 vdd.n575 185
R15785 vdd.n574 vdd.n413 185
R15786 vdd.n570 vdd.n569 185
R15787 vdd.n568 vdd.n567 185
R15788 vdd.n566 vdd.n565 185
R15789 vdd.n564 vdd.n415 185
R15790 vdd.n560 vdd.n559 185
R15791 vdd.n558 vdd.n557 185
R15792 vdd.n556 vdd.n555 185
R15793 vdd.n554 vdd.n417 185
R15794 vdd.n550 vdd.n549 185
R15795 vdd.n548 vdd.n547 185
R15796 vdd.n546 vdd.n545 185
R15797 vdd.n544 vdd.n421 185
R15798 vdd.n540 vdd.n539 185
R15799 vdd.n538 vdd.n537 185
R15800 vdd.n536 vdd.n535 185
R15801 vdd.n534 vdd.n423 185
R15802 vdd.n530 vdd.n529 185
R15803 vdd.n528 vdd.n527 185
R15804 vdd.n526 vdd.n525 185
R15805 vdd.n524 vdd.n425 185
R15806 vdd.n520 vdd.n519 185
R15807 vdd.n518 vdd.n517 185
R15808 vdd.n516 vdd.n515 185
R15809 vdd.n514 vdd.n427 185
R15810 vdd.n510 vdd.n509 185
R15811 vdd.n508 vdd.n507 185
R15812 vdd.n506 vdd.n505 185
R15813 vdd.n504 vdd.n429 185
R15814 vdd.n500 vdd.n499 185
R15815 vdd.n498 vdd.n497 185
R15816 vdd.n496 vdd.n495 185
R15817 vdd.n494 vdd.n433 185
R15818 vdd.n490 vdd.n489 185
R15819 vdd.n488 vdd.n487 185
R15820 vdd.n486 vdd.n485 185
R15821 vdd.n484 vdd.n435 185
R15822 vdd.n480 vdd.n479 185
R15823 vdd.n478 vdd.n477 185
R15824 vdd.n476 vdd.n475 185
R15825 vdd.n474 vdd.n437 185
R15826 vdd.n470 vdd.n469 185
R15827 vdd.n468 vdd.n467 185
R15828 vdd.n466 vdd.n465 185
R15829 vdd.n464 vdd.n439 185
R15830 vdd.n460 vdd.n459 185
R15831 vdd.n458 vdd.n457 185
R15832 vdd.n456 vdd.n455 185
R15833 vdd.n454 vdd.n441 185
R15834 vdd.n450 vdd.n449 185
R15835 vdd.n448 vdd.n447 185
R15836 vdd.n446 vdd.n445 185
R15837 vdd.n3247 vdd.n372 185
R15838 vdd.n3254 vdd.n372 185
R15839 vdd.n3246 vdd.n371 185
R15840 vdd.n3255 vdd.n371 185
R15841 vdd.n3245 vdd.n3244 185
R15842 vdd.n3244 vdd.n363 185
R15843 vdd.n602 vdd.n362 185
R15844 vdd.n3261 vdd.n362 185
R15845 vdd.n3240 vdd.n361 185
R15846 vdd.n3262 vdd.n361 185
R15847 vdd.n3239 vdd.n360 185
R15848 vdd.n3263 vdd.n360 185
R15849 vdd.n3238 vdd.n3237 185
R15850 vdd.n3237 vdd.n3236 185
R15851 vdd.n604 vdd.n352 185
R15852 vdd.n3269 vdd.n352 185
R15853 vdd.n3232 vdd.n351 185
R15854 vdd.n3270 vdd.n351 185
R15855 vdd.n3231 vdd.n350 185
R15856 vdd.n3271 vdd.n350 185
R15857 vdd.n3230 vdd.n3229 185
R15858 vdd.n3229 vdd.n349 185
R15859 vdd.n606 vdd.n341 185
R15860 vdd.n3277 vdd.n341 185
R15861 vdd.n3225 vdd.n340 185
R15862 vdd.n3278 vdd.n340 185
R15863 vdd.n3224 vdd.n339 185
R15864 vdd.n3279 vdd.n339 185
R15865 vdd.n3223 vdd.n3222 185
R15866 vdd.n3222 vdd.n332 185
R15867 vdd.n608 vdd.n331 185
R15868 vdd.n3285 vdd.n331 185
R15869 vdd.n3218 vdd.n330 185
R15870 vdd.n3286 vdd.n330 185
R15871 vdd.n3217 vdd.n329 185
R15872 vdd.n3287 vdd.n329 185
R15873 vdd.n3216 vdd.n3215 185
R15874 vdd.n3215 vdd.n328 185
R15875 vdd.n3214 vdd.n610 185
R15876 vdd.n3214 vdd.n3213 185
R15877 vdd.n3202 vdd.n612 185
R15878 vdd.n613 vdd.n612 185
R15879 vdd.n3204 vdd.n3203 185
R15880 vdd.n3205 vdd.n3204 185
R15881 vdd.n620 vdd.n619 185
R15882 vdd.n624 vdd.n619 185
R15883 vdd.n3196 vdd.n3195 185
R15884 vdd.n3195 vdd.n3194 185
R15885 vdd.n623 vdd.n622 185
R15886 vdd.n3185 vdd.n623 185
R15887 vdd.n3184 vdd.n3183 185
R15888 vdd.n3186 vdd.n3184 185
R15889 vdd.n631 vdd.n630 185
R15890 vdd.n636 vdd.n630 185
R15891 vdd.n3179 vdd.n3178 185
R15892 vdd.n3178 vdd.n3177 185
R15893 vdd.n634 vdd.n633 185
R15894 vdd.n635 vdd.n634 185
R15895 vdd.n3168 vdd.n3167 185
R15896 vdd.n3169 vdd.n3168 185
R15897 vdd.n644 vdd.n643 185
R15898 vdd.n643 vdd.n642 185
R15899 vdd.n3163 vdd.n3162 185
R15900 vdd.n3162 vdd.n3161 185
R15901 vdd.n647 vdd.n646 185
R15902 vdd.n648 vdd.n647 185
R15903 vdd.n3152 vdd.n3151 185
R15904 vdd.n3153 vdd.n3152 185
R15905 vdd.n655 vdd.n654 185
R15906 vdd.n659 vdd.n654 185
R15907 vdd.n3147 vdd.n3146 185
R15908 vdd.n3146 vdd.n3145 185
R15909 vdd.n884 vdd.n883 185
R15910 vdd.n2772 vdd.n2771 185
R15911 vdd.n2770 vdd.n2555 185
R15912 vdd.n2774 vdd.n2555 185
R15913 vdd.n2769 vdd.n2768 185
R15914 vdd.n2767 vdd.n2766 185
R15915 vdd.n2765 vdd.n2764 185
R15916 vdd.n2763 vdd.n2762 185
R15917 vdd.n2761 vdd.n2760 185
R15918 vdd.n2759 vdd.n2758 185
R15919 vdd.n2757 vdd.n2756 185
R15920 vdd.n2755 vdd.n2754 185
R15921 vdd.n2753 vdd.n2752 185
R15922 vdd.n2751 vdd.n2750 185
R15923 vdd.n2749 vdd.n2748 185
R15924 vdd.n2747 vdd.n2746 185
R15925 vdd.n2745 vdd.n2744 185
R15926 vdd.n2743 vdd.n2742 185
R15927 vdd.n2741 vdd.n2740 185
R15928 vdd.n2739 vdd.n2738 185
R15929 vdd.n2737 vdd.n2736 185
R15930 vdd.n2735 vdd.n2734 185
R15931 vdd.n2733 vdd.n2732 185
R15932 vdd.n2731 vdd.n2730 185
R15933 vdd.n2729 vdd.n2728 185
R15934 vdd.n2727 vdd.n2726 185
R15935 vdd.n2725 vdd.n2724 185
R15936 vdd.n2723 vdd.n2722 185
R15937 vdd.n2721 vdd.n2720 185
R15938 vdd.n2719 vdd.n2718 185
R15939 vdd.n2717 vdd.n2716 185
R15940 vdd.n2715 vdd.n2714 185
R15941 vdd.n2713 vdd.n2712 185
R15942 vdd.n2710 vdd.n2709 185
R15943 vdd.n2708 vdd.n2707 185
R15944 vdd.n2706 vdd.n2705 185
R15945 vdd.n2913 vdd.n2912 185
R15946 vdd.n2914 vdd.n803 185
R15947 vdd.n2916 vdd.n2915 185
R15948 vdd.n2918 vdd.n801 185
R15949 vdd.n2920 vdd.n2919 185
R15950 vdd.n2921 vdd.n800 185
R15951 vdd.n2923 vdd.n2922 185
R15952 vdd.n2925 vdd.n798 185
R15953 vdd.n2927 vdd.n2926 185
R15954 vdd.n2928 vdd.n797 185
R15955 vdd.n2930 vdd.n2929 185
R15956 vdd.n2932 vdd.n795 185
R15957 vdd.n2934 vdd.n2933 185
R15958 vdd.n2935 vdd.n794 185
R15959 vdd.n2937 vdd.n2936 185
R15960 vdd.n2939 vdd.n792 185
R15961 vdd.n2941 vdd.n2940 185
R15962 vdd.n2943 vdd.n791 185
R15963 vdd.n2945 vdd.n2944 185
R15964 vdd.n2947 vdd.n789 185
R15965 vdd.n2949 vdd.n2948 185
R15966 vdd.n2950 vdd.n788 185
R15967 vdd.n2952 vdd.n2951 185
R15968 vdd.n2954 vdd.n786 185
R15969 vdd.n2956 vdd.n2955 185
R15970 vdd.n2957 vdd.n785 185
R15971 vdd.n2959 vdd.n2958 185
R15972 vdd.n2961 vdd.n783 185
R15973 vdd.n2963 vdd.n2962 185
R15974 vdd.n2964 vdd.n782 185
R15975 vdd.n2966 vdd.n2965 185
R15976 vdd.n2968 vdd.n781 185
R15977 vdd.n2969 vdd.n780 185
R15978 vdd.n2972 vdd.n2971 185
R15979 vdd.n2973 vdd.n778 185
R15980 vdd.n778 vdd.n756 185
R15981 vdd.n2910 vdd.n775 185
R15982 vdd.n2976 vdd.n775 185
R15983 vdd.n2909 vdd.n2908 185
R15984 vdd.n2908 vdd.n774 185
R15985 vdd.n2907 vdd.n807 185
R15986 vdd.n2907 vdd.n2906 185
R15987 vdd.n2661 vdd.n808 185
R15988 vdd.n817 vdd.n808 185
R15989 vdd.n2662 vdd.n815 185
R15990 vdd.n2900 vdd.n815 185
R15991 vdd.n2664 vdd.n2663 185
R15992 vdd.n2663 vdd.n814 185
R15993 vdd.n2665 vdd.n823 185
R15994 vdd.n2849 vdd.n823 185
R15995 vdd.n2667 vdd.n2666 185
R15996 vdd.n2666 vdd.n822 185
R15997 vdd.n2668 vdd.n829 185
R15998 vdd.n2843 vdd.n829 185
R15999 vdd.n2670 vdd.n2669 185
R16000 vdd.n2669 vdd.n828 185
R16001 vdd.n2671 vdd.n834 185
R16002 vdd.n2835 vdd.n834 185
R16003 vdd.n2673 vdd.n2672 185
R16004 vdd.n2672 vdd.n841 185
R16005 vdd.n2674 vdd.n839 185
R16006 vdd.n2829 vdd.n839 185
R16007 vdd.n2676 vdd.n2675 185
R16008 vdd.n2677 vdd.n2676 185
R16009 vdd.n2660 vdd.n846 185
R16010 vdd.n2823 vdd.n846 185
R16011 vdd.n2659 vdd.n2658 185
R16012 vdd.n2658 vdd.n845 185
R16013 vdd.n2657 vdd.n852 185
R16014 vdd.n2817 vdd.n852 185
R16015 vdd.n2656 vdd.n2655 185
R16016 vdd.n2655 vdd.n851 185
R16017 vdd.n2654 vdd.n857 185
R16018 vdd.n2811 vdd.n857 185
R16019 vdd.n2653 vdd.n2652 185
R16020 vdd.n2652 vdd.n864 185
R16021 vdd.n2651 vdd.n862 185
R16022 vdd.n2805 vdd.n862 185
R16023 vdd.n2650 vdd.n2649 185
R16024 vdd.n2649 vdd.n871 185
R16025 vdd.n2648 vdd.n869 185
R16026 vdd.n2799 vdd.n869 185
R16027 vdd.n2647 vdd.n2646 185
R16028 vdd.n2646 vdd.n868 185
R16029 vdd.n2558 vdd.n875 185
R16030 vdd.n2793 vdd.n875 185
R16031 vdd.n2700 vdd.n2699 185
R16032 vdd.n2699 vdd.n2698 185
R16033 vdd.n2701 vdd.n880 185
R16034 vdd.n2787 vdd.n880 185
R16035 vdd.n2703 vdd.n2702 185
R16036 vdd.n2702 vdd.t256 185
R16037 vdd.n2704 vdd.n885 185
R16038 vdd.n2781 vdd.n885 185
R16039 vdd.n2783 vdd.n2782 185
R16040 vdd.n2782 vdd.n2781 185
R16041 vdd.n2784 vdd.n882 185
R16042 vdd.n882 vdd.t256 185
R16043 vdd.n2786 vdd.n2785 185
R16044 vdd.n2787 vdd.n2786 185
R16045 vdd.n874 vdd.n873 185
R16046 vdd.n2698 vdd.n874 185
R16047 vdd.n2795 vdd.n2794 185
R16048 vdd.n2794 vdd.n2793 185
R16049 vdd.n2796 vdd.n872 185
R16050 vdd.n872 vdd.n868 185
R16051 vdd.n2798 vdd.n2797 185
R16052 vdd.n2799 vdd.n2798 185
R16053 vdd.n861 vdd.n860 185
R16054 vdd.n871 vdd.n861 185
R16055 vdd.n2807 vdd.n2806 185
R16056 vdd.n2806 vdd.n2805 185
R16057 vdd.n2808 vdd.n859 185
R16058 vdd.n864 vdd.n859 185
R16059 vdd.n2810 vdd.n2809 185
R16060 vdd.n2811 vdd.n2810 185
R16061 vdd.n850 vdd.n849 185
R16062 vdd.n851 vdd.n850 185
R16063 vdd.n2819 vdd.n2818 185
R16064 vdd.n2818 vdd.n2817 185
R16065 vdd.n2820 vdd.n848 185
R16066 vdd.n848 vdd.n845 185
R16067 vdd.n2822 vdd.n2821 185
R16068 vdd.n2823 vdd.n2822 185
R16069 vdd.n838 vdd.n837 185
R16070 vdd.n2677 vdd.n838 185
R16071 vdd.n2831 vdd.n2830 185
R16072 vdd.n2830 vdd.n2829 185
R16073 vdd.n2832 vdd.n836 185
R16074 vdd.n841 vdd.n836 185
R16075 vdd.n2834 vdd.n2833 185
R16076 vdd.n2835 vdd.n2834 185
R16077 vdd.n827 vdd.n826 185
R16078 vdd.n828 vdd.n827 185
R16079 vdd.n2845 vdd.n2844 185
R16080 vdd.n2844 vdd.n2843 185
R16081 vdd.n2846 vdd.n825 185
R16082 vdd.n825 vdd.n822 185
R16083 vdd.n2848 vdd.n2847 185
R16084 vdd.n2849 vdd.n2848 185
R16085 vdd.n813 vdd.n812 185
R16086 vdd.n814 vdd.n813 185
R16087 vdd.n2902 vdd.n2901 185
R16088 vdd.n2901 vdd.n2900 185
R16089 vdd.n2903 vdd.n811 185
R16090 vdd.n817 vdd.n811 185
R16091 vdd.n2905 vdd.n2904 185
R16092 vdd.n2906 vdd.n2905 185
R16093 vdd.n779 vdd.n777 185
R16094 vdd.n777 vdd.n774 185
R16095 vdd.n2975 vdd.n2974 185
R16096 vdd.n2976 vdd.n2975 185
R16097 vdd.n2448 vdd.n2447 185
R16098 vdd.n2449 vdd.n2448 185
R16099 vdd.n935 vdd.n933 185
R16100 vdd.n933 vdd.t1 185
R16101 vdd.n2363 vdd.n942 185
R16102 vdd.n2374 vdd.n942 185
R16103 vdd.n2364 vdd.n951 185
R16104 vdd.n2073 vdd.n951 185
R16105 vdd.n2366 vdd.n2365 185
R16106 vdd.n2367 vdd.n2366 185
R16107 vdd.n2362 vdd.n950 185
R16108 vdd.n950 vdd.n947 185
R16109 vdd.n2361 vdd.n2360 185
R16110 vdd.n2360 vdd.n2359 185
R16111 vdd.n953 vdd.n952 185
R16112 vdd.n954 vdd.n953 185
R16113 vdd.n2352 vdd.n2351 185
R16114 vdd.n2353 vdd.n2352 185
R16115 vdd.n2350 vdd.n963 185
R16116 vdd.n963 vdd.n960 185
R16117 vdd.n2349 vdd.n2348 185
R16118 vdd.n2348 vdd.n2347 185
R16119 vdd.n965 vdd.n964 185
R16120 vdd.n973 vdd.n965 185
R16121 vdd.n2340 vdd.n2339 185
R16122 vdd.n2341 vdd.n2340 185
R16123 vdd.n2338 vdd.n974 185
R16124 vdd.n979 vdd.n974 185
R16125 vdd.n2337 vdd.n2336 185
R16126 vdd.n2336 vdd.n2335 185
R16127 vdd.n976 vdd.n975 185
R16128 vdd.n2174 vdd.n976 185
R16129 vdd.n2328 vdd.n2327 185
R16130 vdd.n2329 vdd.n2328 185
R16131 vdd.n2326 vdd.n986 185
R16132 vdd.n986 vdd.n983 185
R16133 vdd.n2325 vdd.n2324 185
R16134 vdd.n2324 vdd.n2323 185
R16135 vdd.n988 vdd.n987 185
R16136 vdd.n989 vdd.n988 185
R16137 vdd.n2316 vdd.n2315 185
R16138 vdd.n2317 vdd.n2316 185
R16139 vdd.n2313 vdd.n997 185
R16140 vdd.n1004 vdd.n997 185
R16141 vdd.n2312 vdd.n2311 185
R16142 vdd.n2311 vdd.n2310 185
R16143 vdd.n1000 vdd.n999 185
R16144 vdd.n1001 vdd.n1000 185
R16145 vdd.n2303 vdd.n2302 185
R16146 vdd.n2304 vdd.n2303 185
R16147 vdd.n2301 vdd.n1011 185
R16148 vdd.n1011 vdd.n1008 185
R16149 vdd.n2300 vdd.n2299 185
R16150 vdd.n2299 vdd.n2298 185
R16151 vdd.n1013 vdd.n1012 185
R16152 vdd.n1014 vdd.n1013 185
R16153 vdd.n2291 vdd.n2290 185
R16154 vdd.n2292 vdd.n2291 185
R16155 vdd.n2379 vdd.n907 185
R16156 vdd.n2521 vdd.n907 185
R16157 vdd.n2381 vdd.n2380 185
R16158 vdd.n2383 vdd.n2382 185
R16159 vdd.n2385 vdd.n2384 185
R16160 vdd.n2387 vdd.n2386 185
R16161 vdd.n2389 vdd.n2388 185
R16162 vdd.n2391 vdd.n2390 185
R16163 vdd.n2393 vdd.n2392 185
R16164 vdd.n2395 vdd.n2394 185
R16165 vdd.n2397 vdd.n2396 185
R16166 vdd.n2399 vdd.n2398 185
R16167 vdd.n2401 vdd.n2400 185
R16168 vdd.n2403 vdd.n2402 185
R16169 vdd.n2405 vdd.n2404 185
R16170 vdd.n2407 vdd.n2406 185
R16171 vdd.n2409 vdd.n2408 185
R16172 vdd.n2411 vdd.n2410 185
R16173 vdd.n2413 vdd.n2412 185
R16174 vdd.n2415 vdd.n2414 185
R16175 vdd.n2417 vdd.n2416 185
R16176 vdd.n2419 vdd.n2418 185
R16177 vdd.n2421 vdd.n2420 185
R16178 vdd.n2423 vdd.n2422 185
R16179 vdd.n2425 vdd.n2424 185
R16180 vdd.n2427 vdd.n2426 185
R16181 vdd.n2429 vdd.n2428 185
R16182 vdd.n2431 vdd.n2430 185
R16183 vdd.n2433 vdd.n2432 185
R16184 vdd.n2435 vdd.n2434 185
R16185 vdd.n2437 vdd.n2436 185
R16186 vdd.n2439 vdd.n2438 185
R16187 vdd.n2441 vdd.n2440 185
R16188 vdd.n2443 vdd.n2442 185
R16189 vdd.n2445 vdd.n2444 185
R16190 vdd.n2446 vdd.n934 185
R16191 vdd.n2378 vdd.n932 185
R16192 vdd.n2449 vdd.n932 185
R16193 vdd.n2377 vdd.n2376 185
R16194 vdd.n2376 vdd.t1 185
R16195 vdd.n2375 vdd.n939 185
R16196 vdd.n2375 vdd.n2374 185
R16197 vdd.n2155 vdd.n940 185
R16198 vdd.n2073 vdd.n940 185
R16199 vdd.n2156 vdd.n949 185
R16200 vdd.n2367 vdd.n949 185
R16201 vdd.n2158 vdd.n2157 185
R16202 vdd.n2157 vdd.n947 185
R16203 vdd.n2159 vdd.n956 185
R16204 vdd.n2359 vdd.n956 185
R16205 vdd.n2161 vdd.n2160 185
R16206 vdd.n2160 vdd.n954 185
R16207 vdd.n2162 vdd.n962 185
R16208 vdd.n2353 vdd.n962 185
R16209 vdd.n2164 vdd.n2163 185
R16210 vdd.n2163 vdd.n960 185
R16211 vdd.n2165 vdd.n967 185
R16212 vdd.n2347 vdd.n967 185
R16213 vdd.n2167 vdd.n2166 185
R16214 vdd.n2166 vdd.n973 185
R16215 vdd.n2168 vdd.n972 185
R16216 vdd.n2341 vdd.n972 185
R16217 vdd.n2170 vdd.n2169 185
R16218 vdd.n2169 vdd.n979 185
R16219 vdd.n2171 vdd.n978 185
R16220 vdd.n2335 vdd.n978 185
R16221 vdd.n2173 vdd.n2172 185
R16222 vdd.n2174 vdd.n2173 185
R16223 vdd.n2154 vdd.n985 185
R16224 vdd.n2329 vdd.n985 185
R16225 vdd.n2153 vdd.n2152 185
R16226 vdd.n2152 vdd.n983 185
R16227 vdd.n2151 vdd.n991 185
R16228 vdd.n2323 vdd.n991 185
R16229 vdd.n2150 vdd.n2149 185
R16230 vdd.n2149 vdd.n989 185
R16231 vdd.n2148 vdd.n996 185
R16232 vdd.n2317 vdd.n996 185
R16233 vdd.n2147 vdd.n2146 185
R16234 vdd.n2146 vdd.n1004 185
R16235 vdd.n2145 vdd.n1003 185
R16236 vdd.n2310 vdd.n1003 185
R16237 vdd.n2144 vdd.n2143 185
R16238 vdd.n2143 vdd.n1001 185
R16239 vdd.n2142 vdd.n1010 185
R16240 vdd.n2304 vdd.n1010 185
R16241 vdd.n2141 vdd.n2140 185
R16242 vdd.n2140 vdd.n1008 185
R16243 vdd.n2139 vdd.n1016 185
R16244 vdd.n2298 vdd.n1016 185
R16245 vdd.n2138 vdd.n2137 185
R16246 vdd.n2137 vdd.n1014 185
R16247 vdd.n2136 vdd.n1022 185
R16248 vdd.n2292 vdd.n1022 185
R16249 vdd.n2289 vdd.n1023 185
R16250 vdd.n2288 vdd.n2287 185
R16251 vdd.n2285 vdd.n1024 185
R16252 vdd.n2283 vdd.n2282 185
R16253 vdd.n2281 vdd.n1025 185
R16254 vdd.n2280 vdd.n2279 185
R16255 vdd.n2277 vdd.n1026 185
R16256 vdd.n2275 vdd.n2274 185
R16257 vdd.n2273 vdd.n1027 185
R16258 vdd.n2272 vdd.n2271 185
R16259 vdd.n2269 vdd.n1028 185
R16260 vdd.n2267 vdd.n2266 185
R16261 vdd.n2265 vdd.n1029 185
R16262 vdd.n2264 vdd.n2263 185
R16263 vdd.n2261 vdd.n1030 185
R16264 vdd.n2259 vdd.n2258 185
R16265 vdd.n2257 vdd.n1031 185
R16266 vdd.n2256 vdd.n1033 185
R16267 vdd.n2101 vdd.n1034 185
R16268 vdd.n2104 vdd.n2103 185
R16269 vdd.n2106 vdd.n2105 185
R16270 vdd.n2108 vdd.n2100 185
R16271 vdd.n2111 vdd.n2110 185
R16272 vdd.n2112 vdd.n2099 185
R16273 vdd.n2114 vdd.n2113 185
R16274 vdd.n2116 vdd.n2098 185
R16275 vdd.n2119 vdd.n2118 185
R16276 vdd.n2120 vdd.n2097 185
R16277 vdd.n2122 vdd.n2121 185
R16278 vdd.n2124 vdd.n2096 185
R16279 vdd.n2127 vdd.n2126 185
R16280 vdd.n2128 vdd.n2093 185
R16281 vdd.n2131 vdd.n2130 185
R16282 vdd.n2133 vdd.n2092 185
R16283 vdd.n2135 vdd.n2134 185
R16284 vdd.n2134 vdd.n1020 185
R16285 vdd.n315 vdd.n314 171.744
R16286 vdd.n314 vdd.n313 171.744
R16287 vdd.n313 vdd.n282 171.744
R16288 vdd.n306 vdd.n282 171.744
R16289 vdd.n306 vdd.n305 171.744
R16290 vdd.n305 vdd.n287 171.744
R16291 vdd.n298 vdd.n287 171.744
R16292 vdd.n298 vdd.n297 171.744
R16293 vdd.n297 vdd.n291 171.744
R16294 vdd.n260 vdd.n259 171.744
R16295 vdd.n259 vdd.n258 171.744
R16296 vdd.n258 vdd.n227 171.744
R16297 vdd.n251 vdd.n227 171.744
R16298 vdd.n251 vdd.n250 171.744
R16299 vdd.n250 vdd.n232 171.744
R16300 vdd.n243 vdd.n232 171.744
R16301 vdd.n243 vdd.n242 171.744
R16302 vdd.n242 vdd.n236 171.744
R16303 vdd.n217 vdd.n216 171.744
R16304 vdd.n216 vdd.n215 171.744
R16305 vdd.n215 vdd.n184 171.744
R16306 vdd.n208 vdd.n184 171.744
R16307 vdd.n208 vdd.n207 171.744
R16308 vdd.n207 vdd.n189 171.744
R16309 vdd.n200 vdd.n189 171.744
R16310 vdd.n200 vdd.n199 171.744
R16311 vdd.n199 vdd.n193 171.744
R16312 vdd.n162 vdd.n161 171.744
R16313 vdd.n161 vdd.n160 171.744
R16314 vdd.n160 vdd.n129 171.744
R16315 vdd.n153 vdd.n129 171.744
R16316 vdd.n153 vdd.n152 171.744
R16317 vdd.n152 vdd.n134 171.744
R16318 vdd.n145 vdd.n134 171.744
R16319 vdd.n145 vdd.n144 171.744
R16320 vdd.n144 vdd.n138 171.744
R16321 vdd.n120 vdd.n119 171.744
R16322 vdd.n119 vdd.n118 171.744
R16323 vdd.n118 vdd.n87 171.744
R16324 vdd.n111 vdd.n87 171.744
R16325 vdd.n111 vdd.n110 171.744
R16326 vdd.n110 vdd.n92 171.744
R16327 vdd.n103 vdd.n92 171.744
R16328 vdd.n103 vdd.n102 171.744
R16329 vdd.n102 vdd.n96 171.744
R16330 vdd.n65 vdd.n64 171.744
R16331 vdd.n64 vdd.n63 171.744
R16332 vdd.n63 vdd.n32 171.744
R16333 vdd.n56 vdd.n32 171.744
R16334 vdd.n56 vdd.n55 171.744
R16335 vdd.n55 vdd.n37 171.744
R16336 vdd.n48 vdd.n37 171.744
R16337 vdd.n48 vdd.n47 171.744
R16338 vdd.n47 vdd.n41 171.744
R16339 vdd.n1684 vdd.n1683 171.744
R16340 vdd.n1683 vdd.n1682 171.744
R16341 vdd.n1682 vdd.n1651 171.744
R16342 vdd.n1675 vdd.n1651 171.744
R16343 vdd.n1675 vdd.n1674 171.744
R16344 vdd.n1674 vdd.n1656 171.744
R16345 vdd.n1667 vdd.n1656 171.744
R16346 vdd.n1667 vdd.n1666 171.744
R16347 vdd.n1666 vdd.n1660 171.744
R16348 vdd.n1739 vdd.n1738 171.744
R16349 vdd.n1738 vdd.n1737 171.744
R16350 vdd.n1737 vdd.n1706 171.744
R16351 vdd.n1730 vdd.n1706 171.744
R16352 vdd.n1730 vdd.n1729 171.744
R16353 vdd.n1729 vdd.n1711 171.744
R16354 vdd.n1722 vdd.n1711 171.744
R16355 vdd.n1722 vdd.n1721 171.744
R16356 vdd.n1721 vdd.n1715 171.744
R16357 vdd.n1586 vdd.n1585 171.744
R16358 vdd.n1585 vdd.n1584 171.744
R16359 vdd.n1584 vdd.n1553 171.744
R16360 vdd.n1577 vdd.n1553 171.744
R16361 vdd.n1577 vdd.n1576 171.744
R16362 vdd.n1576 vdd.n1558 171.744
R16363 vdd.n1569 vdd.n1558 171.744
R16364 vdd.n1569 vdd.n1568 171.744
R16365 vdd.n1568 vdd.n1562 171.744
R16366 vdd.n1641 vdd.n1640 171.744
R16367 vdd.n1640 vdd.n1639 171.744
R16368 vdd.n1639 vdd.n1608 171.744
R16369 vdd.n1632 vdd.n1608 171.744
R16370 vdd.n1632 vdd.n1631 171.744
R16371 vdd.n1631 vdd.n1613 171.744
R16372 vdd.n1624 vdd.n1613 171.744
R16373 vdd.n1624 vdd.n1623 171.744
R16374 vdd.n1623 vdd.n1617 171.744
R16375 vdd.n1489 vdd.n1488 171.744
R16376 vdd.n1488 vdd.n1487 171.744
R16377 vdd.n1487 vdd.n1456 171.744
R16378 vdd.n1480 vdd.n1456 171.744
R16379 vdd.n1480 vdd.n1479 171.744
R16380 vdd.n1479 vdd.n1461 171.744
R16381 vdd.n1472 vdd.n1461 171.744
R16382 vdd.n1472 vdd.n1471 171.744
R16383 vdd.n1471 vdd.n1465 171.744
R16384 vdd.n1544 vdd.n1543 171.744
R16385 vdd.n1543 vdd.n1542 171.744
R16386 vdd.n1542 vdd.n1511 171.744
R16387 vdd.n1535 vdd.n1511 171.744
R16388 vdd.n1535 vdd.n1534 171.744
R16389 vdd.n1534 vdd.n1516 171.744
R16390 vdd.n1527 vdd.n1516 171.744
R16391 vdd.n1527 vdd.n1526 171.744
R16392 vdd.n1526 vdd.n1520 171.744
R16393 vdd.n449 vdd.n448 146.341
R16394 vdd.n455 vdd.n454 146.341
R16395 vdd.n459 vdd.n458 146.341
R16396 vdd.n465 vdd.n464 146.341
R16397 vdd.n469 vdd.n468 146.341
R16398 vdd.n475 vdd.n474 146.341
R16399 vdd.n479 vdd.n478 146.341
R16400 vdd.n485 vdd.n484 146.341
R16401 vdd.n489 vdd.n488 146.341
R16402 vdd.n495 vdd.n494 146.341
R16403 vdd.n499 vdd.n498 146.341
R16404 vdd.n505 vdd.n504 146.341
R16405 vdd.n509 vdd.n508 146.341
R16406 vdd.n515 vdd.n514 146.341
R16407 vdd.n519 vdd.n518 146.341
R16408 vdd.n525 vdd.n524 146.341
R16409 vdd.n529 vdd.n528 146.341
R16410 vdd.n535 vdd.n534 146.341
R16411 vdd.n539 vdd.n538 146.341
R16412 vdd.n545 vdd.n544 146.341
R16413 vdd.n549 vdd.n548 146.341
R16414 vdd.n555 vdd.n554 146.341
R16415 vdd.n559 vdd.n558 146.341
R16416 vdd.n565 vdd.n564 146.341
R16417 vdd.n569 vdd.n568 146.341
R16418 vdd.n575 vdd.n574 146.341
R16419 vdd.n579 vdd.n578 146.341
R16420 vdd.n585 vdd.n584 146.341
R16421 vdd.n589 vdd.n588 146.341
R16422 vdd.n595 vdd.n594 146.341
R16423 vdd.n597 vdd.n404 146.341
R16424 vdd.n3146 vdd.n654 146.341
R16425 vdd.n3152 vdd.n654 146.341
R16426 vdd.n3152 vdd.n647 146.341
R16427 vdd.n3162 vdd.n647 146.341
R16428 vdd.n3162 vdd.n643 146.341
R16429 vdd.n3168 vdd.n643 146.341
R16430 vdd.n3168 vdd.n634 146.341
R16431 vdd.n3178 vdd.n634 146.341
R16432 vdd.n3178 vdd.n630 146.341
R16433 vdd.n3184 vdd.n630 146.341
R16434 vdd.n3184 vdd.n623 146.341
R16435 vdd.n3195 vdd.n623 146.341
R16436 vdd.n3195 vdd.n619 146.341
R16437 vdd.n3204 vdd.n619 146.341
R16438 vdd.n3204 vdd.n612 146.341
R16439 vdd.n3214 vdd.n612 146.341
R16440 vdd.n3215 vdd.n3214 146.341
R16441 vdd.n3215 vdd.n329 146.341
R16442 vdd.n330 vdd.n329 146.341
R16443 vdd.n331 vdd.n330 146.341
R16444 vdd.n3222 vdd.n331 146.341
R16445 vdd.n3222 vdd.n339 146.341
R16446 vdd.n340 vdd.n339 146.341
R16447 vdd.n341 vdd.n340 146.341
R16448 vdd.n3229 vdd.n341 146.341
R16449 vdd.n3229 vdd.n350 146.341
R16450 vdd.n351 vdd.n350 146.341
R16451 vdd.n352 vdd.n351 146.341
R16452 vdd.n3237 vdd.n352 146.341
R16453 vdd.n3237 vdd.n360 146.341
R16454 vdd.n361 vdd.n360 146.341
R16455 vdd.n362 vdd.n361 146.341
R16456 vdd.n3244 vdd.n362 146.341
R16457 vdd.n3244 vdd.n371 146.341
R16458 vdd.n372 vdd.n371 146.341
R16459 vdd.n3138 vdd.n3136 146.341
R16460 vdd.n3136 vdd.n3135 146.341
R16461 vdd.n3132 vdd.n3131 146.341
R16462 vdd.n3128 vdd.n3127 146.341
R16463 vdd.n3125 vdd.n669 146.341
R16464 vdd.n3121 vdd.n3119 146.341
R16465 vdd.n3117 vdd.n675 146.341
R16466 vdd.n3113 vdd.n3111 146.341
R16467 vdd.n3109 vdd.n681 146.341
R16468 vdd.n3105 vdd.n3103 146.341
R16469 vdd.n3101 vdd.n689 146.341
R16470 vdd.n3097 vdd.n3095 146.341
R16471 vdd.n3093 vdd.n695 146.341
R16472 vdd.n3089 vdd.n3087 146.341
R16473 vdd.n3085 vdd.n701 146.341
R16474 vdd.n3081 vdd.n3079 146.341
R16475 vdd.n3077 vdd.n707 146.341
R16476 vdd.n3073 vdd.n3071 146.341
R16477 vdd.n3069 vdd.n713 146.341
R16478 vdd.n3065 vdd.n3063 146.341
R16479 vdd.n3061 vdd.n719 146.341
R16480 vdd.n3054 vdd.n728 146.341
R16481 vdd.n3052 vdd.n3051 146.341
R16482 vdd.n3048 vdd.n3047 146.341
R16483 vdd.n3045 vdd.n733 146.341
R16484 vdd.n3041 vdd.n3039 146.341
R16485 vdd.n3037 vdd.n739 146.341
R16486 vdd.n3033 vdd.n3031 146.341
R16487 vdd.n3029 vdd.n745 146.341
R16488 vdd.n3025 vdd.n3023 146.341
R16489 vdd.n3020 vdd.n3019 146.341
R16490 vdd.n3016 vdd.n657 146.341
R16491 vdd.n3144 vdd.n653 146.341
R16492 vdd.n3154 vdd.n653 146.341
R16493 vdd.n3154 vdd.n649 146.341
R16494 vdd.n3160 vdd.n649 146.341
R16495 vdd.n3160 vdd.n641 146.341
R16496 vdd.n3170 vdd.n641 146.341
R16497 vdd.n3170 vdd.n637 146.341
R16498 vdd.n3176 vdd.n637 146.341
R16499 vdd.n3176 vdd.n629 146.341
R16500 vdd.n3187 vdd.n629 146.341
R16501 vdd.n3187 vdd.n625 146.341
R16502 vdd.n3193 vdd.n625 146.341
R16503 vdd.n3193 vdd.n618 146.341
R16504 vdd.n3206 vdd.n618 146.341
R16505 vdd.n3206 vdd.n614 146.341
R16506 vdd.n3212 vdd.n614 146.341
R16507 vdd.n3212 vdd.n326 146.341
R16508 vdd.n3288 vdd.n326 146.341
R16509 vdd.n3288 vdd.n327 146.341
R16510 vdd.n3284 vdd.n327 146.341
R16511 vdd.n3284 vdd.n333 146.341
R16512 vdd.n3280 vdd.n333 146.341
R16513 vdd.n3280 vdd.n338 146.341
R16514 vdd.n3276 vdd.n338 146.341
R16515 vdd.n3276 vdd.n342 146.341
R16516 vdd.n3272 vdd.n342 146.341
R16517 vdd.n3272 vdd.n348 146.341
R16518 vdd.n3268 vdd.n348 146.341
R16519 vdd.n3268 vdd.n353 146.341
R16520 vdd.n3264 vdd.n353 146.341
R16521 vdd.n3264 vdd.n359 146.341
R16522 vdd.n3260 vdd.n359 146.341
R16523 vdd.n3260 vdd.n364 146.341
R16524 vdd.n3256 vdd.n364 146.341
R16525 vdd.n3256 vdd.n370 146.341
R16526 vdd.n2239 vdd.n2238 146.341
R16527 vdd.n2236 vdd.n1820 146.341
R16528 vdd.n2016 vdd.n1826 146.341
R16529 vdd.n2014 vdd.n2013 146.341
R16530 vdd.n2011 vdd.n1828 146.341
R16531 vdd.n2007 vdd.n2006 146.341
R16532 vdd.n2004 vdd.n1835 146.341
R16533 vdd.n2000 vdd.n1999 146.341
R16534 vdd.n1997 vdd.n1842 146.341
R16535 vdd.n1853 vdd.n1850 146.341
R16536 vdd.n1989 vdd.n1988 146.341
R16537 vdd.n1986 vdd.n1855 146.341
R16538 vdd.n1982 vdd.n1981 146.341
R16539 vdd.n1979 vdd.n1861 146.341
R16540 vdd.n1975 vdd.n1974 146.341
R16541 vdd.n1972 vdd.n1868 146.341
R16542 vdd.n1968 vdd.n1967 146.341
R16543 vdd.n1965 vdd.n1875 146.341
R16544 vdd.n1961 vdd.n1960 146.341
R16545 vdd.n1958 vdd.n1882 146.341
R16546 vdd.n1893 vdd.n1890 146.341
R16547 vdd.n1950 vdd.n1949 146.341
R16548 vdd.n1947 vdd.n1895 146.341
R16549 vdd.n1943 vdd.n1942 146.341
R16550 vdd.n1940 vdd.n1901 146.341
R16551 vdd.n1936 vdd.n1935 146.341
R16552 vdd.n1933 vdd.n1908 146.341
R16553 vdd.n1929 vdd.n1928 146.341
R16554 vdd.n1926 vdd.n1923 146.341
R16555 vdd.n1921 vdd.n1918 146.341
R16556 vdd.n1916 vdd.n1040 146.341
R16557 vdd.n1381 vdd.n1145 146.341
R16558 vdd.n1381 vdd.n1137 146.341
R16559 vdd.n1391 vdd.n1137 146.341
R16560 vdd.n1391 vdd.n1133 146.341
R16561 vdd.n1397 vdd.n1133 146.341
R16562 vdd.n1397 vdd.n1125 146.341
R16563 vdd.n1408 vdd.n1125 146.341
R16564 vdd.n1408 vdd.n1121 146.341
R16565 vdd.n1414 vdd.n1121 146.341
R16566 vdd.n1414 vdd.n1115 146.341
R16567 vdd.n1425 vdd.n1115 146.341
R16568 vdd.n1425 vdd.n1111 146.341
R16569 vdd.n1431 vdd.n1111 146.341
R16570 vdd.n1431 vdd.n1102 146.341
R16571 vdd.n1441 vdd.n1102 146.341
R16572 vdd.n1441 vdd.n1098 146.341
R16573 vdd.n1447 vdd.n1098 146.341
R16574 vdd.n1447 vdd.n1091 146.341
R16575 vdd.n1753 vdd.n1091 146.341
R16576 vdd.n1753 vdd.n1087 146.341
R16577 vdd.n1759 vdd.n1087 146.341
R16578 vdd.n1759 vdd.n1080 146.341
R16579 vdd.n1769 vdd.n1080 146.341
R16580 vdd.n1769 vdd.n1076 146.341
R16581 vdd.n1775 vdd.n1076 146.341
R16582 vdd.n1775 vdd.n1068 146.341
R16583 vdd.n1786 vdd.n1068 146.341
R16584 vdd.n1786 vdd.n1064 146.341
R16585 vdd.n1792 vdd.n1064 146.341
R16586 vdd.n1792 vdd.n1058 146.341
R16587 vdd.n1803 vdd.n1058 146.341
R16588 vdd.n1803 vdd.n1053 146.341
R16589 vdd.n1811 vdd.n1053 146.341
R16590 vdd.n1811 vdd.n1042 146.341
R16591 vdd.n2247 vdd.n1042 146.341
R16592 vdd.n1183 vdd.n1182 146.341
R16593 vdd.n1187 vdd.n1182 146.341
R16594 vdd.n1189 vdd.n1188 146.341
R16595 vdd.n1193 vdd.n1192 146.341
R16596 vdd.n1195 vdd.n1194 146.341
R16597 vdd.n1199 vdd.n1198 146.341
R16598 vdd.n1201 vdd.n1200 146.341
R16599 vdd.n1205 vdd.n1204 146.341
R16600 vdd.n1207 vdd.n1206 146.341
R16601 vdd.n1339 vdd.n1338 146.341
R16602 vdd.n1211 vdd.n1210 146.341
R16603 vdd.n1215 vdd.n1214 146.341
R16604 vdd.n1217 vdd.n1216 146.341
R16605 vdd.n1221 vdd.n1220 146.341
R16606 vdd.n1223 vdd.n1222 146.341
R16607 vdd.n1227 vdd.n1226 146.341
R16608 vdd.n1229 vdd.n1228 146.341
R16609 vdd.n1233 vdd.n1232 146.341
R16610 vdd.n1235 vdd.n1234 146.341
R16611 vdd.n1239 vdd.n1238 146.341
R16612 vdd.n1303 vdd.n1240 146.341
R16613 vdd.n1244 vdd.n1243 146.341
R16614 vdd.n1246 vdd.n1245 146.341
R16615 vdd.n1250 vdd.n1249 146.341
R16616 vdd.n1252 vdd.n1251 146.341
R16617 vdd.n1256 vdd.n1255 146.341
R16618 vdd.n1258 vdd.n1257 146.341
R16619 vdd.n1262 vdd.n1261 146.341
R16620 vdd.n1264 vdd.n1263 146.341
R16621 vdd.n1268 vdd.n1267 146.341
R16622 vdd.n1270 vdd.n1269 146.341
R16623 vdd.n1375 vdd.n1151 146.341
R16624 vdd.n1383 vdd.n1143 146.341
R16625 vdd.n1383 vdd.n1139 146.341
R16626 vdd.n1389 vdd.n1139 146.341
R16627 vdd.n1389 vdd.n1131 146.341
R16628 vdd.n1400 vdd.n1131 146.341
R16629 vdd.n1400 vdd.n1127 146.341
R16630 vdd.n1406 vdd.n1127 146.341
R16631 vdd.n1406 vdd.n1120 146.341
R16632 vdd.n1417 vdd.n1120 146.341
R16633 vdd.n1417 vdd.n1116 146.341
R16634 vdd.n1423 vdd.n1116 146.341
R16635 vdd.n1423 vdd.n1109 146.341
R16636 vdd.n1433 vdd.n1109 146.341
R16637 vdd.n1433 vdd.n1105 146.341
R16638 vdd.n1439 vdd.n1105 146.341
R16639 vdd.n1439 vdd.n1097 146.341
R16640 vdd.n1450 vdd.n1097 146.341
R16641 vdd.n1450 vdd.n1093 146.341
R16642 vdd.n1751 vdd.n1093 146.341
R16643 vdd.n1751 vdd.n1086 146.341
R16644 vdd.n1761 vdd.n1086 146.341
R16645 vdd.n1761 vdd.n1082 146.341
R16646 vdd.n1767 vdd.n1082 146.341
R16647 vdd.n1767 vdd.n1074 146.341
R16648 vdd.n1778 vdd.n1074 146.341
R16649 vdd.n1778 vdd.n1070 146.341
R16650 vdd.n1784 vdd.n1070 146.341
R16651 vdd.n1784 vdd.n1063 146.341
R16652 vdd.n1795 vdd.n1063 146.341
R16653 vdd.n1795 vdd.n1059 146.341
R16654 vdd.n1801 vdd.n1059 146.341
R16655 vdd.n1801 vdd.n1051 146.341
R16656 vdd.n1813 vdd.n1051 146.341
R16657 vdd.n1813 vdd.n1046 146.341
R16658 vdd.n2245 vdd.n1046 146.341
R16659 vdd.n1045 vdd.n1020 141.707
R16660 vdd.n756 vdd.n658 141.707
R16661 vdd.n2094 vdd.t233 127.284
R16662 vdd.n936 vdd.t217 127.284
R16663 vdd.n2068 vdd.t255 127.284
R16664 vdd.n928 vdd.t242 127.284
R16665 vdd.n2839 vdd.t204 127.284
R16666 vdd.n2839 vdd.t205 127.284
R16667 vdd.n2559 vdd.t240 127.284
R16668 vdd.n804 vdd.t221 127.284
R16669 vdd.n2556 vdd.t226 127.284
R16670 vdd.n768 vdd.t228 127.284
R16671 vdd.n998 vdd.t236 127.284
R16672 vdd.n998 vdd.t237 127.284
R16673 vdd.n22 vdd.n20 117.314
R16674 vdd.n17 vdd.n15 117.314
R16675 vdd.n27 vdd.n26 116.927
R16676 vdd.n24 vdd.n23 116.927
R16677 vdd.n22 vdd.n21 116.927
R16678 vdd.n17 vdd.n16 116.927
R16679 vdd.n19 vdd.n18 116.927
R16680 vdd.n27 vdd.n25 116.927
R16681 vdd.n2095 vdd.t232 111.188
R16682 vdd.n937 vdd.t218 111.188
R16683 vdd.n2069 vdd.t254 111.188
R16684 vdd.n929 vdd.t243 111.188
R16685 vdd.n2560 vdd.t239 111.188
R16686 vdd.n805 vdd.t222 111.188
R16687 vdd.n2557 vdd.t225 111.188
R16688 vdd.n769 vdd.t229 111.188
R16689 vdd.n2782 vdd.n882 99.5127
R16690 vdd.n2786 vdd.n882 99.5127
R16691 vdd.n2786 vdd.n874 99.5127
R16692 vdd.n2794 vdd.n874 99.5127
R16693 vdd.n2794 vdd.n872 99.5127
R16694 vdd.n2798 vdd.n872 99.5127
R16695 vdd.n2798 vdd.n861 99.5127
R16696 vdd.n2806 vdd.n861 99.5127
R16697 vdd.n2806 vdd.n859 99.5127
R16698 vdd.n2810 vdd.n859 99.5127
R16699 vdd.n2810 vdd.n850 99.5127
R16700 vdd.n2818 vdd.n850 99.5127
R16701 vdd.n2818 vdd.n848 99.5127
R16702 vdd.n2822 vdd.n848 99.5127
R16703 vdd.n2822 vdd.n838 99.5127
R16704 vdd.n2830 vdd.n838 99.5127
R16705 vdd.n2830 vdd.n836 99.5127
R16706 vdd.n2834 vdd.n836 99.5127
R16707 vdd.n2834 vdd.n827 99.5127
R16708 vdd.n2844 vdd.n827 99.5127
R16709 vdd.n2844 vdd.n825 99.5127
R16710 vdd.n2848 vdd.n825 99.5127
R16711 vdd.n2848 vdd.n813 99.5127
R16712 vdd.n2901 vdd.n813 99.5127
R16713 vdd.n2901 vdd.n811 99.5127
R16714 vdd.n2905 vdd.n811 99.5127
R16715 vdd.n2905 vdd.n777 99.5127
R16716 vdd.n2975 vdd.n777 99.5127
R16717 vdd.n2971 vdd.n778 99.5127
R16718 vdd.n2969 vdd.n2968 99.5127
R16719 vdd.n2966 vdd.n782 99.5127
R16720 vdd.n2962 vdd.n2961 99.5127
R16721 vdd.n2959 vdd.n785 99.5127
R16722 vdd.n2955 vdd.n2954 99.5127
R16723 vdd.n2952 vdd.n788 99.5127
R16724 vdd.n2948 vdd.n2947 99.5127
R16725 vdd.n2945 vdd.n791 99.5127
R16726 vdd.n2940 vdd.n2939 99.5127
R16727 vdd.n2937 vdd.n794 99.5127
R16728 vdd.n2933 vdd.n2932 99.5127
R16729 vdd.n2930 vdd.n797 99.5127
R16730 vdd.n2926 vdd.n2925 99.5127
R16731 vdd.n2923 vdd.n800 99.5127
R16732 vdd.n2919 vdd.n2918 99.5127
R16733 vdd.n2916 vdd.n803 99.5127
R16734 vdd.n2702 vdd.n885 99.5127
R16735 vdd.n2702 vdd.n880 99.5127
R16736 vdd.n2699 vdd.n880 99.5127
R16737 vdd.n2699 vdd.n875 99.5127
R16738 vdd.n2646 vdd.n875 99.5127
R16739 vdd.n2646 vdd.n869 99.5127
R16740 vdd.n2649 vdd.n869 99.5127
R16741 vdd.n2649 vdd.n862 99.5127
R16742 vdd.n2652 vdd.n862 99.5127
R16743 vdd.n2652 vdd.n857 99.5127
R16744 vdd.n2655 vdd.n857 99.5127
R16745 vdd.n2655 vdd.n852 99.5127
R16746 vdd.n2658 vdd.n852 99.5127
R16747 vdd.n2658 vdd.n846 99.5127
R16748 vdd.n2676 vdd.n846 99.5127
R16749 vdd.n2676 vdd.n839 99.5127
R16750 vdd.n2672 vdd.n839 99.5127
R16751 vdd.n2672 vdd.n834 99.5127
R16752 vdd.n2669 vdd.n834 99.5127
R16753 vdd.n2669 vdd.n829 99.5127
R16754 vdd.n2666 vdd.n829 99.5127
R16755 vdd.n2666 vdd.n823 99.5127
R16756 vdd.n2663 vdd.n823 99.5127
R16757 vdd.n2663 vdd.n815 99.5127
R16758 vdd.n815 vdd.n808 99.5127
R16759 vdd.n2907 vdd.n808 99.5127
R16760 vdd.n2908 vdd.n2907 99.5127
R16761 vdd.n2908 vdd.n775 99.5127
R16762 vdd.n2772 vdd.n2555 99.5127
R16763 vdd.n2768 vdd.n2555 99.5127
R16764 vdd.n2766 vdd.n2765 99.5127
R16765 vdd.n2762 vdd.n2761 99.5127
R16766 vdd.n2758 vdd.n2757 99.5127
R16767 vdd.n2754 vdd.n2753 99.5127
R16768 vdd.n2750 vdd.n2749 99.5127
R16769 vdd.n2746 vdd.n2745 99.5127
R16770 vdd.n2742 vdd.n2741 99.5127
R16771 vdd.n2738 vdd.n2737 99.5127
R16772 vdd.n2734 vdd.n2733 99.5127
R16773 vdd.n2730 vdd.n2729 99.5127
R16774 vdd.n2726 vdd.n2725 99.5127
R16775 vdd.n2722 vdd.n2721 99.5127
R16776 vdd.n2718 vdd.n2717 99.5127
R16777 vdd.n2714 vdd.n2713 99.5127
R16778 vdd.n2709 vdd.n2708 99.5127
R16779 vdd.n2520 vdd.n926 99.5127
R16780 vdd.n2516 vdd.n2515 99.5127
R16781 vdd.n2512 vdd.n2511 99.5127
R16782 vdd.n2508 vdd.n2507 99.5127
R16783 vdd.n2504 vdd.n2503 99.5127
R16784 vdd.n2500 vdd.n2499 99.5127
R16785 vdd.n2496 vdd.n2495 99.5127
R16786 vdd.n2492 vdd.n2491 99.5127
R16787 vdd.n2488 vdd.n2487 99.5127
R16788 vdd.n2484 vdd.n2483 99.5127
R16789 vdd.n2480 vdd.n2479 99.5127
R16790 vdd.n2476 vdd.n2475 99.5127
R16791 vdd.n2472 vdd.n2471 99.5127
R16792 vdd.n2468 vdd.n2467 99.5127
R16793 vdd.n2464 vdd.n2463 99.5127
R16794 vdd.n2460 vdd.n2459 99.5127
R16795 vdd.n2455 vdd.n2454 99.5127
R16796 vdd.n2193 vdd.n1021 99.5127
R16797 vdd.n2193 vdd.n1015 99.5127
R16798 vdd.n2190 vdd.n1015 99.5127
R16799 vdd.n2190 vdd.n1009 99.5127
R16800 vdd.n2187 vdd.n1009 99.5127
R16801 vdd.n2187 vdd.n1002 99.5127
R16802 vdd.n2184 vdd.n1002 99.5127
R16803 vdd.n2184 vdd.n995 99.5127
R16804 vdd.n2181 vdd.n995 99.5127
R16805 vdd.n2181 vdd.n990 99.5127
R16806 vdd.n2178 vdd.n990 99.5127
R16807 vdd.n2178 vdd.n984 99.5127
R16808 vdd.n2175 vdd.n984 99.5127
R16809 vdd.n2175 vdd.n977 99.5127
R16810 vdd.n2089 vdd.n977 99.5127
R16811 vdd.n2089 vdd.n971 99.5127
R16812 vdd.n2086 vdd.n971 99.5127
R16813 vdd.n2086 vdd.n966 99.5127
R16814 vdd.n2083 vdd.n966 99.5127
R16815 vdd.n2083 vdd.n961 99.5127
R16816 vdd.n2080 vdd.n961 99.5127
R16817 vdd.n2080 vdd.n955 99.5127
R16818 vdd.n2077 vdd.n955 99.5127
R16819 vdd.n2077 vdd.n948 99.5127
R16820 vdd.n2074 vdd.n948 99.5127
R16821 vdd.n2074 vdd.n941 99.5127
R16822 vdd.n941 vdd.n931 99.5127
R16823 vdd.n2450 vdd.n931 99.5127
R16824 vdd.n2028 vdd.n2026 99.5127
R16825 vdd.n2032 vdd.n2026 99.5127
R16826 vdd.n2036 vdd.n2034 99.5127
R16827 vdd.n2040 vdd.n2024 99.5127
R16828 vdd.n2044 vdd.n2042 99.5127
R16829 vdd.n2048 vdd.n2022 99.5127
R16830 vdd.n2052 vdd.n2050 99.5127
R16831 vdd.n2056 vdd.n2020 99.5127
R16832 vdd.n2059 vdd.n2058 99.5127
R16833 vdd.n2229 vdd.n2227 99.5127
R16834 vdd.n2225 vdd.n2061 99.5127
R16835 vdd.n2221 vdd.n2219 99.5127
R16836 vdd.n2217 vdd.n2063 99.5127
R16837 vdd.n2213 vdd.n2211 99.5127
R16838 vdd.n2209 vdd.n2065 99.5127
R16839 vdd.n2205 vdd.n2203 99.5127
R16840 vdd.n2201 vdd.n2067 99.5127
R16841 vdd.n2293 vdd.n1017 99.5127
R16842 vdd.n2297 vdd.n1017 99.5127
R16843 vdd.n2297 vdd.n1007 99.5127
R16844 vdd.n2305 vdd.n1007 99.5127
R16845 vdd.n2305 vdd.n1005 99.5127
R16846 vdd.n2309 vdd.n1005 99.5127
R16847 vdd.n2309 vdd.n994 99.5127
R16848 vdd.n2318 vdd.n994 99.5127
R16849 vdd.n2318 vdd.n992 99.5127
R16850 vdd.n2322 vdd.n992 99.5127
R16851 vdd.n2322 vdd.n982 99.5127
R16852 vdd.n2330 vdd.n982 99.5127
R16853 vdd.n2330 vdd.n980 99.5127
R16854 vdd.n2334 vdd.n980 99.5127
R16855 vdd.n2334 vdd.n970 99.5127
R16856 vdd.n2342 vdd.n970 99.5127
R16857 vdd.n2342 vdd.n968 99.5127
R16858 vdd.n2346 vdd.n968 99.5127
R16859 vdd.n2346 vdd.n959 99.5127
R16860 vdd.n2354 vdd.n959 99.5127
R16861 vdd.n2354 vdd.n957 99.5127
R16862 vdd.n2358 vdd.n957 99.5127
R16863 vdd.n2358 vdd.n946 99.5127
R16864 vdd.n2368 vdd.n946 99.5127
R16865 vdd.n2368 vdd.n943 99.5127
R16866 vdd.n2373 vdd.n943 99.5127
R16867 vdd.n2373 vdd.n944 99.5127
R16868 vdd.n944 vdd.n925 99.5127
R16869 vdd.n2891 vdd.n2890 99.5127
R16870 vdd.n2888 vdd.n2854 99.5127
R16871 vdd.n2884 vdd.n2883 99.5127
R16872 vdd.n2881 vdd.n2857 99.5127
R16873 vdd.n2877 vdd.n2876 99.5127
R16874 vdd.n2874 vdd.n2860 99.5127
R16875 vdd.n2870 vdd.n2869 99.5127
R16876 vdd.n2867 vdd.n2864 99.5127
R16877 vdd.n3008 vdd.n755 99.5127
R16878 vdd.n3006 vdd.n3005 99.5127
R16879 vdd.n3003 vdd.n758 99.5127
R16880 vdd.n2999 vdd.n2998 99.5127
R16881 vdd.n2996 vdd.n761 99.5127
R16882 vdd.n2992 vdd.n2991 99.5127
R16883 vdd.n2989 vdd.n764 99.5127
R16884 vdd.n2985 vdd.n2984 99.5127
R16885 vdd.n2982 vdd.n767 99.5127
R16886 vdd.n2626 vdd.n886 99.5127
R16887 vdd.n2626 vdd.n881 99.5127
R16888 vdd.n2697 vdd.n881 99.5127
R16889 vdd.n2697 vdd.n876 99.5127
R16890 vdd.n2693 vdd.n876 99.5127
R16891 vdd.n2693 vdd.n870 99.5127
R16892 vdd.n2690 vdd.n870 99.5127
R16893 vdd.n2690 vdd.n863 99.5127
R16894 vdd.n2687 vdd.n863 99.5127
R16895 vdd.n2687 vdd.n858 99.5127
R16896 vdd.n2684 vdd.n858 99.5127
R16897 vdd.n2684 vdd.n853 99.5127
R16898 vdd.n2681 vdd.n853 99.5127
R16899 vdd.n2681 vdd.n847 99.5127
R16900 vdd.n2678 vdd.n847 99.5127
R16901 vdd.n2678 vdd.n840 99.5127
R16902 vdd.n2643 vdd.n840 99.5127
R16903 vdd.n2643 vdd.n835 99.5127
R16904 vdd.n2640 vdd.n835 99.5127
R16905 vdd.n2640 vdd.n830 99.5127
R16906 vdd.n2637 vdd.n830 99.5127
R16907 vdd.n2637 vdd.n824 99.5127
R16908 vdd.n2634 vdd.n824 99.5127
R16909 vdd.n2634 vdd.n816 99.5127
R16910 vdd.n2631 vdd.n816 99.5127
R16911 vdd.n2631 vdd.n809 99.5127
R16912 vdd.n809 vdd.n773 99.5127
R16913 vdd.n2977 vdd.n773 99.5127
R16914 vdd.n2776 vdd.n889 99.5127
R16915 vdd.n2564 vdd.n2563 99.5127
R16916 vdd.n2568 vdd.n2567 99.5127
R16917 vdd.n2572 vdd.n2571 99.5127
R16918 vdd.n2576 vdd.n2575 99.5127
R16919 vdd.n2580 vdd.n2579 99.5127
R16920 vdd.n2584 vdd.n2583 99.5127
R16921 vdd.n2588 vdd.n2587 99.5127
R16922 vdd.n2592 vdd.n2591 99.5127
R16923 vdd.n2596 vdd.n2595 99.5127
R16924 vdd.n2600 vdd.n2599 99.5127
R16925 vdd.n2604 vdd.n2603 99.5127
R16926 vdd.n2608 vdd.n2607 99.5127
R16927 vdd.n2612 vdd.n2611 99.5127
R16928 vdd.n2616 vdd.n2615 99.5127
R16929 vdd.n2620 vdd.n2619 99.5127
R16930 vdd.n2622 vdd.n2554 99.5127
R16931 vdd.n2780 vdd.n879 99.5127
R16932 vdd.n2788 vdd.n879 99.5127
R16933 vdd.n2788 vdd.n877 99.5127
R16934 vdd.n2792 vdd.n877 99.5127
R16935 vdd.n2792 vdd.n867 99.5127
R16936 vdd.n2800 vdd.n867 99.5127
R16937 vdd.n2800 vdd.n865 99.5127
R16938 vdd.n2804 vdd.n865 99.5127
R16939 vdd.n2804 vdd.n856 99.5127
R16940 vdd.n2812 vdd.n856 99.5127
R16941 vdd.n2812 vdd.n854 99.5127
R16942 vdd.n2816 vdd.n854 99.5127
R16943 vdd.n2816 vdd.n844 99.5127
R16944 vdd.n2824 vdd.n844 99.5127
R16945 vdd.n2824 vdd.n842 99.5127
R16946 vdd.n2828 vdd.n842 99.5127
R16947 vdd.n2828 vdd.n833 99.5127
R16948 vdd.n2836 vdd.n833 99.5127
R16949 vdd.n2836 vdd.n831 99.5127
R16950 vdd.n2842 vdd.n831 99.5127
R16951 vdd.n2842 vdd.n821 99.5127
R16952 vdd.n2850 vdd.n821 99.5127
R16953 vdd.n2850 vdd.n818 99.5127
R16954 vdd.n2899 vdd.n818 99.5127
R16955 vdd.n2899 vdd.n819 99.5127
R16956 vdd.n819 vdd.n810 99.5127
R16957 vdd.n2894 vdd.n810 99.5127
R16958 vdd.n2894 vdd.n776 99.5127
R16959 vdd.n2444 vdd.n2443 99.5127
R16960 vdd.n2440 vdd.n2439 99.5127
R16961 vdd.n2436 vdd.n2435 99.5127
R16962 vdd.n2432 vdd.n2431 99.5127
R16963 vdd.n2428 vdd.n2427 99.5127
R16964 vdd.n2424 vdd.n2423 99.5127
R16965 vdd.n2420 vdd.n2419 99.5127
R16966 vdd.n2416 vdd.n2415 99.5127
R16967 vdd.n2412 vdd.n2411 99.5127
R16968 vdd.n2408 vdd.n2407 99.5127
R16969 vdd.n2404 vdd.n2403 99.5127
R16970 vdd.n2400 vdd.n2399 99.5127
R16971 vdd.n2396 vdd.n2395 99.5127
R16972 vdd.n2392 vdd.n2391 99.5127
R16973 vdd.n2388 vdd.n2387 99.5127
R16974 vdd.n2384 vdd.n2383 99.5127
R16975 vdd.n2380 vdd.n907 99.5127
R16976 vdd.n2137 vdd.n1022 99.5127
R16977 vdd.n2137 vdd.n1016 99.5127
R16978 vdd.n2140 vdd.n1016 99.5127
R16979 vdd.n2140 vdd.n1010 99.5127
R16980 vdd.n2143 vdd.n1010 99.5127
R16981 vdd.n2143 vdd.n1003 99.5127
R16982 vdd.n2146 vdd.n1003 99.5127
R16983 vdd.n2146 vdd.n996 99.5127
R16984 vdd.n2149 vdd.n996 99.5127
R16985 vdd.n2149 vdd.n991 99.5127
R16986 vdd.n2152 vdd.n991 99.5127
R16987 vdd.n2152 vdd.n985 99.5127
R16988 vdd.n2173 vdd.n985 99.5127
R16989 vdd.n2173 vdd.n978 99.5127
R16990 vdd.n2169 vdd.n978 99.5127
R16991 vdd.n2169 vdd.n972 99.5127
R16992 vdd.n2166 vdd.n972 99.5127
R16993 vdd.n2166 vdd.n967 99.5127
R16994 vdd.n2163 vdd.n967 99.5127
R16995 vdd.n2163 vdd.n962 99.5127
R16996 vdd.n2160 vdd.n962 99.5127
R16997 vdd.n2160 vdd.n956 99.5127
R16998 vdd.n2157 vdd.n956 99.5127
R16999 vdd.n2157 vdd.n949 99.5127
R17000 vdd.n949 vdd.n940 99.5127
R17001 vdd.n2375 vdd.n940 99.5127
R17002 vdd.n2376 vdd.n2375 99.5127
R17003 vdd.n2376 vdd.n932 99.5127
R17004 vdd.n2287 vdd.n2285 99.5127
R17005 vdd.n2283 vdd.n1025 99.5127
R17006 vdd.n2279 vdd.n2277 99.5127
R17007 vdd.n2275 vdd.n1027 99.5127
R17008 vdd.n2271 vdd.n2269 99.5127
R17009 vdd.n2267 vdd.n1029 99.5127
R17010 vdd.n2263 vdd.n2261 99.5127
R17011 vdd.n2259 vdd.n1031 99.5127
R17012 vdd.n2101 vdd.n1033 99.5127
R17013 vdd.n2106 vdd.n2103 99.5127
R17014 vdd.n2110 vdd.n2108 99.5127
R17015 vdd.n2114 vdd.n2099 99.5127
R17016 vdd.n2118 vdd.n2116 99.5127
R17017 vdd.n2122 vdd.n2097 99.5127
R17018 vdd.n2126 vdd.n2124 99.5127
R17019 vdd.n2131 vdd.n2093 99.5127
R17020 vdd.n2134 vdd.n2133 99.5127
R17021 vdd.n2291 vdd.n1013 99.5127
R17022 vdd.n2299 vdd.n1013 99.5127
R17023 vdd.n2299 vdd.n1011 99.5127
R17024 vdd.n2303 vdd.n1011 99.5127
R17025 vdd.n2303 vdd.n1000 99.5127
R17026 vdd.n2311 vdd.n1000 99.5127
R17027 vdd.n2311 vdd.n997 99.5127
R17028 vdd.n2316 vdd.n997 99.5127
R17029 vdd.n2316 vdd.n988 99.5127
R17030 vdd.n2324 vdd.n988 99.5127
R17031 vdd.n2324 vdd.n986 99.5127
R17032 vdd.n2328 vdd.n986 99.5127
R17033 vdd.n2328 vdd.n976 99.5127
R17034 vdd.n2336 vdd.n976 99.5127
R17035 vdd.n2336 vdd.n974 99.5127
R17036 vdd.n2340 vdd.n974 99.5127
R17037 vdd.n2340 vdd.n965 99.5127
R17038 vdd.n2348 vdd.n965 99.5127
R17039 vdd.n2348 vdd.n963 99.5127
R17040 vdd.n2352 vdd.n963 99.5127
R17041 vdd.n2352 vdd.n953 99.5127
R17042 vdd.n2360 vdd.n953 99.5127
R17043 vdd.n2360 vdd.n950 99.5127
R17044 vdd.n2366 vdd.n950 99.5127
R17045 vdd.n2366 vdd.n951 99.5127
R17046 vdd.n951 vdd.n942 99.5127
R17047 vdd.n942 vdd.n933 99.5127
R17048 vdd.n2448 vdd.n933 99.5127
R17049 vdd.n9 vdd.n7 98.9633
R17050 vdd.n2 vdd.n0 98.9633
R17051 vdd.n9 vdd.n8 98.6055
R17052 vdd.n11 vdd.n10 98.6055
R17053 vdd.n13 vdd.n12 98.6055
R17054 vdd.n6 vdd.n5 98.6055
R17055 vdd.n4 vdd.n3 98.6055
R17056 vdd.n2 vdd.n1 98.6055
R17057 vdd.t116 vdd.n291 85.8723
R17058 vdd.t90 vdd.n236 85.8723
R17059 vdd.t102 vdd.n193 85.8723
R17060 vdd.t79 vdd.n138 85.8723
R17061 vdd.t34 vdd.n96 85.8723
R17062 vdd.t14 vdd.n41 85.8723
R17063 vdd.t129 vdd.n1660 85.8723
R17064 vdd.t40 vdd.n1715 85.8723
R17065 vdd.t114 vdd.n1562 85.8723
R17066 vdd.t24 vdd.n1617 85.8723
R17067 vdd.t12 vdd.n1465 85.8723
R17068 vdd.t37 vdd.n1520 85.8723
R17069 vdd.n2840 vdd.n2839 78.546
R17070 vdd.n2314 vdd.n998 78.546
R17071 vdd.n278 vdd.n277 75.1835
R17072 vdd.n276 vdd.n275 75.1835
R17073 vdd.n274 vdd.n273 75.1835
R17074 vdd.n272 vdd.n271 75.1835
R17075 vdd.n270 vdd.n269 75.1835
R17076 vdd.n268 vdd.n267 75.1835
R17077 vdd.n266 vdd.n265 75.1835
R17078 vdd.n180 vdd.n179 75.1835
R17079 vdd.n178 vdd.n177 75.1835
R17080 vdd.n176 vdd.n175 75.1835
R17081 vdd.n174 vdd.n173 75.1835
R17082 vdd.n172 vdd.n171 75.1835
R17083 vdd.n170 vdd.n169 75.1835
R17084 vdd.n168 vdd.n167 75.1835
R17085 vdd.n83 vdd.n82 75.1835
R17086 vdd.n81 vdd.n80 75.1835
R17087 vdd.n79 vdd.n78 75.1835
R17088 vdd.n77 vdd.n76 75.1835
R17089 vdd.n75 vdd.n74 75.1835
R17090 vdd.n73 vdd.n72 75.1835
R17091 vdd.n71 vdd.n70 75.1835
R17092 vdd.n1690 vdd.n1689 75.1835
R17093 vdd.n1692 vdd.n1691 75.1835
R17094 vdd.n1694 vdd.n1693 75.1835
R17095 vdd.n1696 vdd.n1695 75.1835
R17096 vdd.n1698 vdd.n1697 75.1835
R17097 vdd.n1700 vdd.n1699 75.1835
R17098 vdd.n1702 vdd.n1701 75.1835
R17099 vdd.n1592 vdd.n1591 75.1835
R17100 vdd.n1594 vdd.n1593 75.1835
R17101 vdd.n1596 vdd.n1595 75.1835
R17102 vdd.n1598 vdd.n1597 75.1835
R17103 vdd.n1600 vdd.n1599 75.1835
R17104 vdd.n1602 vdd.n1601 75.1835
R17105 vdd.n1604 vdd.n1603 75.1835
R17106 vdd.n1495 vdd.n1494 75.1835
R17107 vdd.n1497 vdd.n1496 75.1835
R17108 vdd.n1499 vdd.n1498 75.1835
R17109 vdd.n1501 vdd.n1500 75.1835
R17110 vdd.n1503 vdd.n1502 75.1835
R17111 vdd.n1505 vdd.n1504 75.1835
R17112 vdd.n1507 vdd.n1506 75.1835
R17113 vdd.n2775 vdd.n2774 72.8958
R17114 vdd.n2774 vdd.n2538 72.8958
R17115 vdd.n2774 vdd.n2539 72.8958
R17116 vdd.n2774 vdd.n2540 72.8958
R17117 vdd.n2774 vdd.n2541 72.8958
R17118 vdd.n2774 vdd.n2542 72.8958
R17119 vdd.n2774 vdd.n2543 72.8958
R17120 vdd.n2774 vdd.n2544 72.8958
R17121 vdd.n2774 vdd.n2545 72.8958
R17122 vdd.n2774 vdd.n2546 72.8958
R17123 vdd.n2774 vdd.n2547 72.8958
R17124 vdd.n2774 vdd.n2548 72.8958
R17125 vdd.n2774 vdd.n2549 72.8958
R17126 vdd.n2774 vdd.n2550 72.8958
R17127 vdd.n2774 vdd.n2551 72.8958
R17128 vdd.n2774 vdd.n2552 72.8958
R17129 vdd.n2774 vdd.n2553 72.8958
R17130 vdd.n772 vdd.n756 72.8958
R17131 vdd.n2983 vdd.n756 72.8958
R17132 vdd.n766 vdd.n756 72.8958
R17133 vdd.n2990 vdd.n756 72.8958
R17134 vdd.n763 vdd.n756 72.8958
R17135 vdd.n2997 vdd.n756 72.8958
R17136 vdd.n760 vdd.n756 72.8958
R17137 vdd.n3004 vdd.n756 72.8958
R17138 vdd.n3007 vdd.n756 72.8958
R17139 vdd.n2863 vdd.n756 72.8958
R17140 vdd.n2868 vdd.n756 72.8958
R17141 vdd.n2862 vdd.n756 72.8958
R17142 vdd.n2875 vdd.n756 72.8958
R17143 vdd.n2859 vdd.n756 72.8958
R17144 vdd.n2882 vdd.n756 72.8958
R17145 vdd.n2856 vdd.n756 72.8958
R17146 vdd.n2889 vdd.n756 72.8958
R17147 vdd.n2027 vdd.n1020 72.8958
R17148 vdd.n2033 vdd.n1020 72.8958
R17149 vdd.n2035 vdd.n1020 72.8958
R17150 vdd.n2041 vdd.n1020 72.8958
R17151 vdd.n2043 vdd.n1020 72.8958
R17152 vdd.n2049 vdd.n1020 72.8958
R17153 vdd.n2051 vdd.n1020 72.8958
R17154 vdd.n2057 vdd.n1020 72.8958
R17155 vdd.n2228 vdd.n1020 72.8958
R17156 vdd.n2226 vdd.n1020 72.8958
R17157 vdd.n2220 vdd.n1020 72.8958
R17158 vdd.n2218 vdd.n1020 72.8958
R17159 vdd.n2212 vdd.n1020 72.8958
R17160 vdd.n2210 vdd.n1020 72.8958
R17161 vdd.n2204 vdd.n1020 72.8958
R17162 vdd.n2202 vdd.n1020 72.8958
R17163 vdd.n2196 vdd.n1020 72.8958
R17164 vdd.n2521 vdd.n908 72.8958
R17165 vdd.n2521 vdd.n909 72.8958
R17166 vdd.n2521 vdd.n910 72.8958
R17167 vdd.n2521 vdd.n911 72.8958
R17168 vdd.n2521 vdd.n912 72.8958
R17169 vdd.n2521 vdd.n913 72.8958
R17170 vdd.n2521 vdd.n914 72.8958
R17171 vdd.n2521 vdd.n915 72.8958
R17172 vdd.n2521 vdd.n916 72.8958
R17173 vdd.n2521 vdd.n917 72.8958
R17174 vdd.n2521 vdd.n918 72.8958
R17175 vdd.n2521 vdd.n919 72.8958
R17176 vdd.n2521 vdd.n920 72.8958
R17177 vdd.n2521 vdd.n921 72.8958
R17178 vdd.n2521 vdd.n922 72.8958
R17179 vdd.n2521 vdd.n923 72.8958
R17180 vdd.n2521 vdd.n924 72.8958
R17181 vdd.n2774 vdd.n2773 72.8958
R17182 vdd.n2774 vdd.n2522 72.8958
R17183 vdd.n2774 vdd.n2523 72.8958
R17184 vdd.n2774 vdd.n2524 72.8958
R17185 vdd.n2774 vdd.n2525 72.8958
R17186 vdd.n2774 vdd.n2526 72.8958
R17187 vdd.n2774 vdd.n2527 72.8958
R17188 vdd.n2774 vdd.n2528 72.8958
R17189 vdd.n2774 vdd.n2529 72.8958
R17190 vdd.n2774 vdd.n2530 72.8958
R17191 vdd.n2774 vdd.n2531 72.8958
R17192 vdd.n2774 vdd.n2532 72.8958
R17193 vdd.n2774 vdd.n2533 72.8958
R17194 vdd.n2774 vdd.n2534 72.8958
R17195 vdd.n2774 vdd.n2535 72.8958
R17196 vdd.n2774 vdd.n2536 72.8958
R17197 vdd.n2774 vdd.n2537 72.8958
R17198 vdd.n2911 vdd.n756 72.8958
R17199 vdd.n2917 vdd.n756 72.8958
R17200 vdd.n802 vdd.n756 72.8958
R17201 vdd.n2924 vdd.n756 72.8958
R17202 vdd.n799 vdd.n756 72.8958
R17203 vdd.n2931 vdd.n756 72.8958
R17204 vdd.n796 vdd.n756 72.8958
R17205 vdd.n2938 vdd.n756 72.8958
R17206 vdd.n793 vdd.n756 72.8958
R17207 vdd.n2946 vdd.n756 72.8958
R17208 vdd.n790 vdd.n756 72.8958
R17209 vdd.n2953 vdd.n756 72.8958
R17210 vdd.n787 vdd.n756 72.8958
R17211 vdd.n2960 vdd.n756 72.8958
R17212 vdd.n784 vdd.n756 72.8958
R17213 vdd.n2967 vdd.n756 72.8958
R17214 vdd.n2970 vdd.n756 72.8958
R17215 vdd.n2521 vdd.n906 72.8958
R17216 vdd.n2521 vdd.n905 72.8958
R17217 vdd.n2521 vdd.n904 72.8958
R17218 vdd.n2521 vdd.n903 72.8958
R17219 vdd.n2521 vdd.n902 72.8958
R17220 vdd.n2521 vdd.n901 72.8958
R17221 vdd.n2521 vdd.n900 72.8958
R17222 vdd.n2521 vdd.n899 72.8958
R17223 vdd.n2521 vdd.n898 72.8958
R17224 vdd.n2521 vdd.n897 72.8958
R17225 vdd.n2521 vdd.n896 72.8958
R17226 vdd.n2521 vdd.n895 72.8958
R17227 vdd.n2521 vdd.n894 72.8958
R17228 vdd.n2521 vdd.n893 72.8958
R17229 vdd.n2521 vdd.n892 72.8958
R17230 vdd.n2521 vdd.n891 72.8958
R17231 vdd.n2521 vdd.n890 72.8958
R17232 vdd.n2286 vdd.n1020 72.8958
R17233 vdd.n2284 vdd.n1020 72.8958
R17234 vdd.n2278 vdd.n1020 72.8958
R17235 vdd.n2276 vdd.n1020 72.8958
R17236 vdd.n2270 vdd.n1020 72.8958
R17237 vdd.n2268 vdd.n1020 72.8958
R17238 vdd.n2262 vdd.n1020 72.8958
R17239 vdd.n2260 vdd.n1020 72.8958
R17240 vdd.n1032 vdd.n1020 72.8958
R17241 vdd.n2102 vdd.n1020 72.8958
R17242 vdd.n2107 vdd.n1020 72.8958
R17243 vdd.n2109 vdd.n1020 72.8958
R17244 vdd.n2115 vdd.n1020 72.8958
R17245 vdd.n2117 vdd.n1020 72.8958
R17246 vdd.n2123 vdd.n1020 72.8958
R17247 vdd.n2125 vdd.n1020 72.8958
R17248 vdd.n2132 vdd.n1020 72.8958
R17249 vdd.n1374 vdd.n1373 66.2847
R17250 vdd.n1374 vdd.n1152 66.2847
R17251 vdd.n1374 vdd.n1153 66.2847
R17252 vdd.n1374 vdd.n1154 66.2847
R17253 vdd.n1374 vdd.n1155 66.2847
R17254 vdd.n1374 vdd.n1156 66.2847
R17255 vdd.n1374 vdd.n1157 66.2847
R17256 vdd.n1374 vdd.n1158 66.2847
R17257 vdd.n1374 vdd.n1159 66.2847
R17258 vdd.n1374 vdd.n1160 66.2847
R17259 vdd.n1374 vdd.n1161 66.2847
R17260 vdd.n1374 vdd.n1162 66.2847
R17261 vdd.n1374 vdd.n1163 66.2847
R17262 vdd.n1374 vdd.n1164 66.2847
R17263 vdd.n1374 vdd.n1165 66.2847
R17264 vdd.n1374 vdd.n1166 66.2847
R17265 vdd.n1374 vdd.n1167 66.2847
R17266 vdd.n1374 vdd.n1168 66.2847
R17267 vdd.n1374 vdd.n1169 66.2847
R17268 vdd.n1374 vdd.n1170 66.2847
R17269 vdd.n1374 vdd.n1171 66.2847
R17270 vdd.n1374 vdd.n1172 66.2847
R17271 vdd.n1374 vdd.n1173 66.2847
R17272 vdd.n1374 vdd.n1174 66.2847
R17273 vdd.n1374 vdd.n1175 66.2847
R17274 vdd.n1374 vdd.n1176 66.2847
R17275 vdd.n1374 vdd.n1177 66.2847
R17276 vdd.n1374 vdd.n1178 66.2847
R17277 vdd.n1374 vdd.n1179 66.2847
R17278 vdd.n1374 vdd.n1180 66.2847
R17279 vdd.n1374 vdd.n1181 66.2847
R17280 vdd.n1045 vdd.n1041 66.2847
R17281 vdd.n1917 vdd.n1045 66.2847
R17282 vdd.n1922 vdd.n1045 66.2847
R17283 vdd.n1927 vdd.n1045 66.2847
R17284 vdd.n1915 vdd.n1045 66.2847
R17285 vdd.n1934 vdd.n1045 66.2847
R17286 vdd.n1907 vdd.n1045 66.2847
R17287 vdd.n1941 vdd.n1045 66.2847
R17288 vdd.n1900 vdd.n1045 66.2847
R17289 vdd.n1948 vdd.n1045 66.2847
R17290 vdd.n1894 vdd.n1045 66.2847
R17291 vdd.n1889 vdd.n1045 66.2847
R17292 vdd.n1959 vdd.n1045 66.2847
R17293 vdd.n1881 vdd.n1045 66.2847
R17294 vdd.n1966 vdd.n1045 66.2847
R17295 vdd.n1874 vdd.n1045 66.2847
R17296 vdd.n1973 vdd.n1045 66.2847
R17297 vdd.n1867 vdd.n1045 66.2847
R17298 vdd.n1980 vdd.n1045 66.2847
R17299 vdd.n1860 vdd.n1045 66.2847
R17300 vdd.n1987 vdd.n1045 66.2847
R17301 vdd.n1854 vdd.n1045 66.2847
R17302 vdd.n1849 vdd.n1045 66.2847
R17303 vdd.n1998 vdd.n1045 66.2847
R17304 vdd.n1841 vdd.n1045 66.2847
R17305 vdd.n2005 vdd.n1045 66.2847
R17306 vdd.n1834 vdd.n1045 66.2847
R17307 vdd.n2012 vdd.n1045 66.2847
R17308 vdd.n2015 vdd.n1045 66.2847
R17309 vdd.n1825 vdd.n1045 66.2847
R17310 vdd.n2237 vdd.n1045 66.2847
R17311 vdd.n1819 vdd.n1045 66.2847
R17312 vdd.n3137 vdd.n658 66.2847
R17313 vdd.n663 vdd.n658 66.2847
R17314 vdd.n666 vdd.n658 66.2847
R17315 vdd.n3126 vdd.n658 66.2847
R17316 vdd.n3120 vdd.n658 66.2847
R17317 vdd.n3118 vdd.n658 66.2847
R17318 vdd.n3112 vdd.n658 66.2847
R17319 vdd.n3110 vdd.n658 66.2847
R17320 vdd.n3104 vdd.n658 66.2847
R17321 vdd.n3102 vdd.n658 66.2847
R17322 vdd.n3096 vdd.n658 66.2847
R17323 vdd.n3094 vdd.n658 66.2847
R17324 vdd.n3088 vdd.n658 66.2847
R17325 vdd.n3086 vdd.n658 66.2847
R17326 vdd.n3080 vdd.n658 66.2847
R17327 vdd.n3078 vdd.n658 66.2847
R17328 vdd.n3072 vdd.n658 66.2847
R17329 vdd.n3070 vdd.n658 66.2847
R17330 vdd.n3064 vdd.n658 66.2847
R17331 vdd.n3062 vdd.n658 66.2847
R17332 vdd.n727 vdd.n658 66.2847
R17333 vdd.n3053 vdd.n658 66.2847
R17334 vdd.n729 vdd.n658 66.2847
R17335 vdd.n3046 vdd.n658 66.2847
R17336 vdd.n3040 vdd.n658 66.2847
R17337 vdd.n3038 vdd.n658 66.2847
R17338 vdd.n3032 vdd.n658 66.2847
R17339 vdd.n3030 vdd.n658 66.2847
R17340 vdd.n3024 vdd.n658 66.2847
R17341 vdd.n750 vdd.n658 66.2847
R17342 vdd.n752 vdd.n658 66.2847
R17343 vdd.n3253 vdd.n3252 66.2847
R17344 vdd.n3253 vdd.n403 66.2847
R17345 vdd.n3253 vdd.n402 66.2847
R17346 vdd.n3253 vdd.n401 66.2847
R17347 vdd.n3253 vdd.n400 66.2847
R17348 vdd.n3253 vdd.n399 66.2847
R17349 vdd.n3253 vdd.n398 66.2847
R17350 vdd.n3253 vdd.n397 66.2847
R17351 vdd.n3253 vdd.n396 66.2847
R17352 vdd.n3253 vdd.n395 66.2847
R17353 vdd.n3253 vdd.n394 66.2847
R17354 vdd.n3253 vdd.n393 66.2847
R17355 vdd.n3253 vdd.n392 66.2847
R17356 vdd.n3253 vdd.n391 66.2847
R17357 vdd.n3253 vdd.n390 66.2847
R17358 vdd.n3253 vdd.n389 66.2847
R17359 vdd.n3253 vdd.n388 66.2847
R17360 vdd.n3253 vdd.n387 66.2847
R17361 vdd.n3253 vdd.n386 66.2847
R17362 vdd.n3253 vdd.n385 66.2847
R17363 vdd.n3253 vdd.n384 66.2847
R17364 vdd.n3253 vdd.n383 66.2847
R17365 vdd.n3253 vdd.n382 66.2847
R17366 vdd.n3253 vdd.n381 66.2847
R17367 vdd.n3253 vdd.n380 66.2847
R17368 vdd.n3253 vdd.n379 66.2847
R17369 vdd.n3253 vdd.n378 66.2847
R17370 vdd.n3253 vdd.n377 66.2847
R17371 vdd.n3253 vdd.n376 66.2847
R17372 vdd.n3253 vdd.n375 66.2847
R17373 vdd.n3253 vdd.n374 66.2847
R17374 vdd.n3253 vdd.n373 66.2847
R17375 vdd.n448 vdd.n373 52.4337
R17376 vdd.n454 vdd.n374 52.4337
R17377 vdd.n458 vdd.n375 52.4337
R17378 vdd.n464 vdd.n376 52.4337
R17379 vdd.n468 vdd.n377 52.4337
R17380 vdd.n474 vdd.n378 52.4337
R17381 vdd.n478 vdd.n379 52.4337
R17382 vdd.n484 vdd.n380 52.4337
R17383 vdd.n488 vdd.n381 52.4337
R17384 vdd.n494 vdd.n382 52.4337
R17385 vdd.n498 vdd.n383 52.4337
R17386 vdd.n504 vdd.n384 52.4337
R17387 vdd.n508 vdd.n385 52.4337
R17388 vdd.n514 vdd.n386 52.4337
R17389 vdd.n518 vdd.n387 52.4337
R17390 vdd.n524 vdd.n388 52.4337
R17391 vdd.n528 vdd.n389 52.4337
R17392 vdd.n534 vdd.n390 52.4337
R17393 vdd.n538 vdd.n391 52.4337
R17394 vdd.n544 vdd.n392 52.4337
R17395 vdd.n548 vdd.n393 52.4337
R17396 vdd.n554 vdd.n394 52.4337
R17397 vdd.n558 vdd.n395 52.4337
R17398 vdd.n564 vdd.n396 52.4337
R17399 vdd.n568 vdd.n397 52.4337
R17400 vdd.n574 vdd.n398 52.4337
R17401 vdd.n578 vdd.n399 52.4337
R17402 vdd.n584 vdd.n400 52.4337
R17403 vdd.n588 vdd.n401 52.4337
R17404 vdd.n594 vdd.n402 52.4337
R17405 vdd.n597 vdd.n403 52.4337
R17406 vdd.n3252 vdd.n3251 52.4337
R17407 vdd.n3137 vdd.n660 52.4337
R17408 vdd.n3135 vdd.n663 52.4337
R17409 vdd.n3131 vdd.n666 52.4337
R17410 vdd.n3127 vdd.n3126 52.4337
R17411 vdd.n3120 vdd.n669 52.4337
R17412 vdd.n3119 vdd.n3118 52.4337
R17413 vdd.n3112 vdd.n675 52.4337
R17414 vdd.n3111 vdd.n3110 52.4337
R17415 vdd.n3104 vdd.n681 52.4337
R17416 vdd.n3103 vdd.n3102 52.4337
R17417 vdd.n3096 vdd.n689 52.4337
R17418 vdd.n3095 vdd.n3094 52.4337
R17419 vdd.n3088 vdd.n695 52.4337
R17420 vdd.n3087 vdd.n3086 52.4337
R17421 vdd.n3080 vdd.n701 52.4337
R17422 vdd.n3079 vdd.n3078 52.4337
R17423 vdd.n3072 vdd.n707 52.4337
R17424 vdd.n3071 vdd.n3070 52.4337
R17425 vdd.n3064 vdd.n713 52.4337
R17426 vdd.n3063 vdd.n3062 52.4337
R17427 vdd.n727 vdd.n719 52.4337
R17428 vdd.n3054 vdd.n3053 52.4337
R17429 vdd.n3051 vdd.n729 52.4337
R17430 vdd.n3047 vdd.n3046 52.4337
R17431 vdd.n3040 vdd.n733 52.4337
R17432 vdd.n3039 vdd.n3038 52.4337
R17433 vdd.n3032 vdd.n739 52.4337
R17434 vdd.n3031 vdd.n3030 52.4337
R17435 vdd.n3024 vdd.n745 52.4337
R17436 vdd.n3023 vdd.n750 52.4337
R17437 vdd.n3019 vdd.n752 52.4337
R17438 vdd.n2239 vdd.n1819 52.4337
R17439 vdd.n2237 vdd.n2236 52.4337
R17440 vdd.n1826 vdd.n1825 52.4337
R17441 vdd.n2015 vdd.n2014 52.4337
R17442 vdd.n2012 vdd.n2011 52.4337
R17443 vdd.n2007 vdd.n1834 52.4337
R17444 vdd.n2005 vdd.n2004 52.4337
R17445 vdd.n2000 vdd.n1841 52.4337
R17446 vdd.n1998 vdd.n1997 52.4337
R17447 vdd.n1850 vdd.n1849 52.4337
R17448 vdd.n1989 vdd.n1854 52.4337
R17449 vdd.n1987 vdd.n1986 52.4337
R17450 vdd.n1982 vdd.n1860 52.4337
R17451 vdd.n1980 vdd.n1979 52.4337
R17452 vdd.n1975 vdd.n1867 52.4337
R17453 vdd.n1973 vdd.n1972 52.4337
R17454 vdd.n1968 vdd.n1874 52.4337
R17455 vdd.n1966 vdd.n1965 52.4337
R17456 vdd.n1961 vdd.n1881 52.4337
R17457 vdd.n1959 vdd.n1958 52.4337
R17458 vdd.n1890 vdd.n1889 52.4337
R17459 vdd.n1950 vdd.n1894 52.4337
R17460 vdd.n1948 vdd.n1947 52.4337
R17461 vdd.n1943 vdd.n1900 52.4337
R17462 vdd.n1941 vdd.n1940 52.4337
R17463 vdd.n1936 vdd.n1907 52.4337
R17464 vdd.n1934 vdd.n1933 52.4337
R17465 vdd.n1929 vdd.n1915 52.4337
R17466 vdd.n1927 vdd.n1926 52.4337
R17467 vdd.n1922 vdd.n1921 52.4337
R17468 vdd.n1917 vdd.n1916 52.4337
R17469 vdd.n2248 vdd.n1041 52.4337
R17470 vdd.n1373 vdd.n1372 52.4337
R17471 vdd.n1187 vdd.n1152 52.4337
R17472 vdd.n1189 vdd.n1153 52.4337
R17473 vdd.n1193 vdd.n1154 52.4337
R17474 vdd.n1195 vdd.n1155 52.4337
R17475 vdd.n1199 vdd.n1156 52.4337
R17476 vdd.n1201 vdd.n1157 52.4337
R17477 vdd.n1205 vdd.n1158 52.4337
R17478 vdd.n1207 vdd.n1159 52.4337
R17479 vdd.n1339 vdd.n1160 52.4337
R17480 vdd.n1211 vdd.n1161 52.4337
R17481 vdd.n1215 vdd.n1162 52.4337
R17482 vdd.n1217 vdd.n1163 52.4337
R17483 vdd.n1221 vdd.n1164 52.4337
R17484 vdd.n1223 vdd.n1165 52.4337
R17485 vdd.n1227 vdd.n1166 52.4337
R17486 vdd.n1229 vdd.n1167 52.4337
R17487 vdd.n1233 vdd.n1168 52.4337
R17488 vdd.n1235 vdd.n1169 52.4337
R17489 vdd.n1239 vdd.n1170 52.4337
R17490 vdd.n1303 vdd.n1171 52.4337
R17491 vdd.n1244 vdd.n1172 52.4337
R17492 vdd.n1246 vdd.n1173 52.4337
R17493 vdd.n1250 vdd.n1174 52.4337
R17494 vdd.n1252 vdd.n1175 52.4337
R17495 vdd.n1256 vdd.n1176 52.4337
R17496 vdd.n1258 vdd.n1177 52.4337
R17497 vdd.n1262 vdd.n1178 52.4337
R17498 vdd.n1264 vdd.n1179 52.4337
R17499 vdd.n1268 vdd.n1180 52.4337
R17500 vdd.n1270 vdd.n1181 52.4337
R17501 vdd.n1373 vdd.n1183 52.4337
R17502 vdd.n1188 vdd.n1152 52.4337
R17503 vdd.n1192 vdd.n1153 52.4337
R17504 vdd.n1194 vdd.n1154 52.4337
R17505 vdd.n1198 vdd.n1155 52.4337
R17506 vdd.n1200 vdd.n1156 52.4337
R17507 vdd.n1204 vdd.n1157 52.4337
R17508 vdd.n1206 vdd.n1158 52.4337
R17509 vdd.n1338 vdd.n1159 52.4337
R17510 vdd.n1210 vdd.n1160 52.4337
R17511 vdd.n1214 vdd.n1161 52.4337
R17512 vdd.n1216 vdd.n1162 52.4337
R17513 vdd.n1220 vdd.n1163 52.4337
R17514 vdd.n1222 vdd.n1164 52.4337
R17515 vdd.n1226 vdd.n1165 52.4337
R17516 vdd.n1228 vdd.n1166 52.4337
R17517 vdd.n1232 vdd.n1167 52.4337
R17518 vdd.n1234 vdd.n1168 52.4337
R17519 vdd.n1238 vdd.n1169 52.4337
R17520 vdd.n1240 vdd.n1170 52.4337
R17521 vdd.n1243 vdd.n1171 52.4337
R17522 vdd.n1245 vdd.n1172 52.4337
R17523 vdd.n1249 vdd.n1173 52.4337
R17524 vdd.n1251 vdd.n1174 52.4337
R17525 vdd.n1255 vdd.n1175 52.4337
R17526 vdd.n1257 vdd.n1176 52.4337
R17527 vdd.n1261 vdd.n1177 52.4337
R17528 vdd.n1263 vdd.n1178 52.4337
R17529 vdd.n1267 vdd.n1179 52.4337
R17530 vdd.n1269 vdd.n1180 52.4337
R17531 vdd.n1181 vdd.n1151 52.4337
R17532 vdd.n1041 vdd.n1040 52.4337
R17533 vdd.n1918 vdd.n1917 52.4337
R17534 vdd.n1923 vdd.n1922 52.4337
R17535 vdd.n1928 vdd.n1927 52.4337
R17536 vdd.n1915 vdd.n1908 52.4337
R17537 vdd.n1935 vdd.n1934 52.4337
R17538 vdd.n1907 vdd.n1901 52.4337
R17539 vdd.n1942 vdd.n1941 52.4337
R17540 vdd.n1900 vdd.n1895 52.4337
R17541 vdd.n1949 vdd.n1948 52.4337
R17542 vdd.n1894 vdd.n1893 52.4337
R17543 vdd.n1889 vdd.n1882 52.4337
R17544 vdd.n1960 vdd.n1959 52.4337
R17545 vdd.n1881 vdd.n1875 52.4337
R17546 vdd.n1967 vdd.n1966 52.4337
R17547 vdd.n1874 vdd.n1868 52.4337
R17548 vdd.n1974 vdd.n1973 52.4337
R17549 vdd.n1867 vdd.n1861 52.4337
R17550 vdd.n1981 vdd.n1980 52.4337
R17551 vdd.n1860 vdd.n1855 52.4337
R17552 vdd.n1988 vdd.n1987 52.4337
R17553 vdd.n1854 vdd.n1853 52.4337
R17554 vdd.n1849 vdd.n1842 52.4337
R17555 vdd.n1999 vdd.n1998 52.4337
R17556 vdd.n1841 vdd.n1835 52.4337
R17557 vdd.n2006 vdd.n2005 52.4337
R17558 vdd.n1834 vdd.n1828 52.4337
R17559 vdd.n2013 vdd.n2012 52.4337
R17560 vdd.n2016 vdd.n2015 52.4337
R17561 vdd.n1825 vdd.n1820 52.4337
R17562 vdd.n2238 vdd.n2237 52.4337
R17563 vdd.n1819 vdd.n1047 52.4337
R17564 vdd.n3138 vdd.n3137 52.4337
R17565 vdd.n3132 vdd.n663 52.4337
R17566 vdd.n3128 vdd.n666 52.4337
R17567 vdd.n3126 vdd.n3125 52.4337
R17568 vdd.n3121 vdd.n3120 52.4337
R17569 vdd.n3118 vdd.n3117 52.4337
R17570 vdd.n3113 vdd.n3112 52.4337
R17571 vdd.n3110 vdd.n3109 52.4337
R17572 vdd.n3105 vdd.n3104 52.4337
R17573 vdd.n3102 vdd.n3101 52.4337
R17574 vdd.n3097 vdd.n3096 52.4337
R17575 vdd.n3094 vdd.n3093 52.4337
R17576 vdd.n3089 vdd.n3088 52.4337
R17577 vdd.n3086 vdd.n3085 52.4337
R17578 vdd.n3081 vdd.n3080 52.4337
R17579 vdd.n3078 vdd.n3077 52.4337
R17580 vdd.n3073 vdd.n3072 52.4337
R17581 vdd.n3070 vdd.n3069 52.4337
R17582 vdd.n3065 vdd.n3064 52.4337
R17583 vdd.n3062 vdd.n3061 52.4337
R17584 vdd.n728 vdd.n727 52.4337
R17585 vdd.n3053 vdd.n3052 52.4337
R17586 vdd.n3048 vdd.n729 52.4337
R17587 vdd.n3046 vdd.n3045 52.4337
R17588 vdd.n3041 vdd.n3040 52.4337
R17589 vdd.n3038 vdd.n3037 52.4337
R17590 vdd.n3033 vdd.n3032 52.4337
R17591 vdd.n3030 vdd.n3029 52.4337
R17592 vdd.n3025 vdd.n3024 52.4337
R17593 vdd.n3020 vdd.n750 52.4337
R17594 vdd.n3016 vdd.n752 52.4337
R17595 vdd.n3252 vdd.n404 52.4337
R17596 vdd.n595 vdd.n403 52.4337
R17597 vdd.n589 vdd.n402 52.4337
R17598 vdd.n585 vdd.n401 52.4337
R17599 vdd.n579 vdd.n400 52.4337
R17600 vdd.n575 vdd.n399 52.4337
R17601 vdd.n569 vdd.n398 52.4337
R17602 vdd.n565 vdd.n397 52.4337
R17603 vdd.n559 vdd.n396 52.4337
R17604 vdd.n555 vdd.n395 52.4337
R17605 vdd.n549 vdd.n394 52.4337
R17606 vdd.n545 vdd.n393 52.4337
R17607 vdd.n539 vdd.n392 52.4337
R17608 vdd.n535 vdd.n391 52.4337
R17609 vdd.n529 vdd.n390 52.4337
R17610 vdd.n525 vdd.n389 52.4337
R17611 vdd.n519 vdd.n388 52.4337
R17612 vdd.n515 vdd.n387 52.4337
R17613 vdd.n509 vdd.n386 52.4337
R17614 vdd.n505 vdd.n385 52.4337
R17615 vdd.n499 vdd.n384 52.4337
R17616 vdd.n495 vdd.n383 52.4337
R17617 vdd.n489 vdd.n382 52.4337
R17618 vdd.n485 vdd.n381 52.4337
R17619 vdd.n479 vdd.n380 52.4337
R17620 vdd.n475 vdd.n379 52.4337
R17621 vdd.n469 vdd.n378 52.4337
R17622 vdd.n465 vdd.n377 52.4337
R17623 vdd.n459 vdd.n376 52.4337
R17624 vdd.n455 vdd.n375 52.4337
R17625 vdd.n449 vdd.n374 52.4337
R17626 vdd.n445 vdd.n373 52.4337
R17627 vdd.t160 vdd.t157 51.4683
R17628 vdd.n266 vdd.n264 42.0461
R17629 vdd.n168 vdd.n166 42.0461
R17630 vdd.n71 vdd.n69 42.0461
R17631 vdd.n1690 vdd.n1688 42.0461
R17632 vdd.n1592 vdd.n1590 42.0461
R17633 vdd.n1495 vdd.n1493 42.0461
R17634 vdd.n320 vdd.n319 41.6884
R17635 vdd.n222 vdd.n221 41.6884
R17636 vdd.n125 vdd.n124 41.6884
R17637 vdd.n1744 vdd.n1743 41.6884
R17638 vdd.n1646 vdd.n1645 41.6884
R17639 vdd.n1549 vdd.n1548 41.6884
R17640 vdd.n1150 vdd.n1149 41.1157
R17641 vdd.n1306 vdd.n1305 41.1157
R17642 vdd.n1342 vdd.n1341 41.1157
R17643 vdd.n407 vdd.n406 41.1157
R17644 vdd.n547 vdd.n420 41.1157
R17645 vdd.n433 vdd.n432 41.1157
R17646 vdd.n2970 vdd.n2969 39.2114
R17647 vdd.n2967 vdd.n2966 39.2114
R17648 vdd.n2962 vdd.n784 39.2114
R17649 vdd.n2960 vdd.n2959 39.2114
R17650 vdd.n2955 vdd.n787 39.2114
R17651 vdd.n2953 vdd.n2952 39.2114
R17652 vdd.n2948 vdd.n790 39.2114
R17653 vdd.n2946 vdd.n2945 39.2114
R17654 vdd.n2940 vdd.n793 39.2114
R17655 vdd.n2938 vdd.n2937 39.2114
R17656 vdd.n2933 vdd.n796 39.2114
R17657 vdd.n2931 vdd.n2930 39.2114
R17658 vdd.n2926 vdd.n799 39.2114
R17659 vdd.n2924 vdd.n2923 39.2114
R17660 vdd.n2919 vdd.n802 39.2114
R17661 vdd.n2917 vdd.n2916 39.2114
R17662 vdd.n2912 vdd.n2911 39.2114
R17663 vdd.n2773 vdd.n884 39.2114
R17664 vdd.n2768 vdd.n2522 39.2114
R17665 vdd.n2765 vdd.n2523 39.2114
R17666 vdd.n2761 vdd.n2524 39.2114
R17667 vdd.n2757 vdd.n2525 39.2114
R17668 vdd.n2753 vdd.n2526 39.2114
R17669 vdd.n2749 vdd.n2527 39.2114
R17670 vdd.n2745 vdd.n2528 39.2114
R17671 vdd.n2741 vdd.n2529 39.2114
R17672 vdd.n2737 vdd.n2530 39.2114
R17673 vdd.n2733 vdd.n2531 39.2114
R17674 vdd.n2729 vdd.n2532 39.2114
R17675 vdd.n2725 vdd.n2533 39.2114
R17676 vdd.n2721 vdd.n2534 39.2114
R17677 vdd.n2717 vdd.n2535 39.2114
R17678 vdd.n2713 vdd.n2536 39.2114
R17679 vdd.n2708 vdd.n2537 39.2114
R17680 vdd.n2516 vdd.n924 39.2114
R17681 vdd.n2512 vdd.n923 39.2114
R17682 vdd.n2508 vdd.n922 39.2114
R17683 vdd.n2504 vdd.n921 39.2114
R17684 vdd.n2500 vdd.n920 39.2114
R17685 vdd.n2496 vdd.n919 39.2114
R17686 vdd.n2492 vdd.n918 39.2114
R17687 vdd.n2488 vdd.n917 39.2114
R17688 vdd.n2484 vdd.n916 39.2114
R17689 vdd.n2480 vdd.n915 39.2114
R17690 vdd.n2476 vdd.n914 39.2114
R17691 vdd.n2472 vdd.n913 39.2114
R17692 vdd.n2468 vdd.n912 39.2114
R17693 vdd.n2464 vdd.n911 39.2114
R17694 vdd.n2460 vdd.n910 39.2114
R17695 vdd.n2455 vdd.n909 39.2114
R17696 vdd.n2451 vdd.n908 39.2114
R17697 vdd.n2027 vdd.n1019 39.2114
R17698 vdd.n2033 vdd.n2032 39.2114
R17699 vdd.n2036 vdd.n2035 39.2114
R17700 vdd.n2041 vdd.n2040 39.2114
R17701 vdd.n2044 vdd.n2043 39.2114
R17702 vdd.n2049 vdd.n2048 39.2114
R17703 vdd.n2052 vdd.n2051 39.2114
R17704 vdd.n2057 vdd.n2056 39.2114
R17705 vdd.n2228 vdd.n2059 39.2114
R17706 vdd.n2227 vdd.n2226 39.2114
R17707 vdd.n2220 vdd.n2061 39.2114
R17708 vdd.n2219 vdd.n2218 39.2114
R17709 vdd.n2212 vdd.n2063 39.2114
R17710 vdd.n2211 vdd.n2210 39.2114
R17711 vdd.n2204 vdd.n2065 39.2114
R17712 vdd.n2203 vdd.n2202 39.2114
R17713 vdd.n2196 vdd.n2067 39.2114
R17714 vdd.n2889 vdd.n2888 39.2114
R17715 vdd.n2884 vdd.n2856 39.2114
R17716 vdd.n2882 vdd.n2881 39.2114
R17717 vdd.n2877 vdd.n2859 39.2114
R17718 vdd.n2875 vdd.n2874 39.2114
R17719 vdd.n2870 vdd.n2862 39.2114
R17720 vdd.n2868 vdd.n2867 39.2114
R17721 vdd.n2863 vdd.n755 39.2114
R17722 vdd.n3007 vdd.n3006 39.2114
R17723 vdd.n3004 vdd.n3003 39.2114
R17724 vdd.n2999 vdd.n760 39.2114
R17725 vdd.n2997 vdd.n2996 39.2114
R17726 vdd.n2992 vdd.n763 39.2114
R17727 vdd.n2990 vdd.n2989 39.2114
R17728 vdd.n2985 vdd.n766 39.2114
R17729 vdd.n2983 vdd.n2982 39.2114
R17730 vdd.n2978 vdd.n772 39.2114
R17731 vdd.n2775 vdd.n887 39.2114
R17732 vdd.n2538 vdd.n889 39.2114
R17733 vdd.n2564 vdd.n2539 39.2114
R17734 vdd.n2568 vdd.n2540 39.2114
R17735 vdd.n2572 vdd.n2541 39.2114
R17736 vdd.n2576 vdd.n2542 39.2114
R17737 vdd.n2580 vdd.n2543 39.2114
R17738 vdd.n2584 vdd.n2544 39.2114
R17739 vdd.n2588 vdd.n2545 39.2114
R17740 vdd.n2592 vdd.n2546 39.2114
R17741 vdd.n2596 vdd.n2547 39.2114
R17742 vdd.n2600 vdd.n2548 39.2114
R17743 vdd.n2604 vdd.n2549 39.2114
R17744 vdd.n2608 vdd.n2550 39.2114
R17745 vdd.n2612 vdd.n2551 39.2114
R17746 vdd.n2616 vdd.n2552 39.2114
R17747 vdd.n2620 vdd.n2553 39.2114
R17748 vdd.n2776 vdd.n2775 39.2114
R17749 vdd.n2563 vdd.n2538 39.2114
R17750 vdd.n2567 vdd.n2539 39.2114
R17751 vdd.n2571 vdd.n2540 39.2114
R17752 vdd.n2575 vdd.n2541 39.2114
R17753 vdd.n2579 vdd.n2542 39.2114
R17754 vdd.n2583 vdd.n2543 39.2114
R17755 vdd.n2587 vdd.n2544 39.2114
R17756 vdd.n2591 vdd.n2545 39.2114
R17757 vdd.n2595 vdd.n2546 39.2114
R17758 vdd.n2599 vdd.n2547 39.2114
R17759 vdd.n2603 vdd.n2548 39.2114
R17760 vdd.n2607 vdd.n2549 39.2114
R17761 vdd.n2611 vdd.n2550 39.2114
R17762 vdd.n2615 vdd.n2551 39.2114
R17763 vdd.n2619 vdd.n2552 39.2114
R17764 vdd.n2622 vdd.n2553 39.2114
R17765 vdd.n772 vdd.n767 39.2114
R17766 vdd.n2984 vdd.n2983 39.2114
R17767 vdd.n766 vdd.n764 39.2114
R17768 vdd.n2991 vdd.n2990 39.2114
R17769 vdd.n763 vdd.n761 39.2114
R17770 vdd.n2998 vdd.n2997 39.2114
R17771 vdd.n760 vdd.n758 39.2114
R17772 vdd.n3005 vdd.n3004 39.2114
R17773 vdd.n3008 vdd.n3007 39.2114
R17774 vdd.n2864 vdd.n2863 39.2114
R17775 vdd.n2869 vdd.n2868 39.2114
R17776 vdd.n2862 vdd.n2860 39.2114
R17777 vdd.n2876 vdd.n2875 39.2114
R17778 vdd.n2859 vdd.n2857 39.2114
R17779 vdd.n2883 vdd.n2882 39.2114
R17780 vdd.n2856 vdd.n2854 39.2114
R17781 vdd.n2890 vdd.n2889 39.2114
R17782 vdd.n2028 vdd.n2027 39.2114
R17783 vdd.n2034 vdd.n2033 39.2114
R17784 vdd.n2035 vdd.n2024 39.2114
R17785 vdd.n2042 vdd.n2041 39.2114
R17786 vdd.n2043 vdd.n2022 39.2114
R17787 vdd.n2050 vdd.n2049 39.2114
R17788 vdd.n2051 vdd.n2020 39.2114
R17789 vdd.n2058 vdd.n2057 39.2114
R17790 vdd.n2229 vdd.n2228 39.2114
R17791 vdd.n2226 vdd.n2225 39.2114
R17792 vdd.n2221 vdd.n2220 39.2114
R17793 vdd.n2218 vdd.n2217 39.2114
R17794 vdd.n2213 vdd.n2212 39.2114
R17795 vdd.n2210 vdd.n2209 39.2114
R17796 vdd.n2205 vdd.n2204 39.2114
R17797 vdd.n2202 vdd.n2201 39.2114
R17798 vdd.n2197 vdd.n2196 39.2114
R17799 vdd.n2454 vdd.n908 39.2114
R17800 vdd.n2459 vdd.n909 39.2114
R17801 vdd.n2463 vdd.n910 39.2114
R17802 vdd.n2467 vdd.n911 39.2114
R17803 vdd.n2471 vdd.n912 39.2114
R17804 vdd.n2475 vdd.n913 39.2114
R17805 vdd.n2479 vdd.n914 39.2114
R17806 vdd.n2483 vdd.n915 39.2114
R17807 vdd.n2487 vdd.n916 39.2114
R17808 vdd.n2491 vdd.n917 39.2114
R17809 vdd.n2495 vdd.n918 39.2114
R17810 vdd.n2499 vdd.n919 39.2114
R17811 vdd.n2503 vdd.n920 39.2114
R17812 vdd.n2507 vdd.n921 39.2114
R17813 vdd.n2511 vdd.n922 39.2114
R17814 vdd.n2515 vdd.n923 39.2114
R17815 vdd.n926 vdd.n924 39.2114
R17816 vdd.n2773 vdd.n2772 39.2114
R17817 vdd.n2766 vdd.n2522 39.2114
R17818 vdd.n2762 vdd.n2523 39.2114
R17819 vdd.n2758 vdd.n2524 39.2114
R17820 vdd.n2754 vdd.n2525 39.2114
R17821 vdd.n2750 vdd.n2526 39.2114
R17822 vdd.n2746 vdd.n2527 39.2114
R17823 vdd.n2742 vdd.n2528 39.2114
R17824 vdd.n2738 vdd.n2529 39.2114
R17825 vdd.n2734 vdd.n2530 39.2114
R17826 vdd.n2730 vdd.n2531 39.2114
R17827 vdd.n2726 vdd.n2532 39.2114
R17828 vdd.n2722 vdd.n2533 39.2114
R17829 vdd.n2718 vdd.n2534 39.2114
R17830 vdd.n2714 vdd.n2535 39.2114
R17831 vdd.n2709 vdd.n2536 39.2114
R17832 vdd.n2705 vdd.n2537 39.2114
R17833 vdd.n2911 vdd.n803 39.2114
R17834 vdd.n2918 vdd.n2917 39.2114
R17835 vdd.n802 vdd.n800 39.2114
R17836 vdd.n2925 vdd.n2924 39.2114
R17837 vdd.n799 vdd.n797 39.2114
R17838 vdd.n2932 vdd.n2931 39.2114
R17839 vdd.n796 vdd.n794 39.2114
R17840 vdd.n2939 vdd.n2938 39.2114
R17841 vdd.n793 vdd.n791 39.2114
R17842 vdd.n2947 vdd.n2946 39.2114
R17843 vdd.n790 vdd.n788 39.2114
R17844 vdd.n2954 vdd.n2953 39.2114
R17845 vdd.n787 vdd.n785 39.2114
R17846 vdd.n2961 vdd.n2960 39.2114
R17847 vdd.n784 vdd.n782 39.2114
R17848 vdd.n2968 vdd.n2967 39.2114
R17849 vdd.n2971 vdd.n2970 39.2114
R17850 vdd.n934 vdd.n890 39.2114
R17851 vdd.n2443 vdd.n891 39.2114
R17852 vdd.n2439 vdd.n892 39.2114
R17853 vdd.n2435 vdd.n893 39.2114
R17854 vdd.n2431 vdd.n894 39.2114
R17855 vdd.n2427 vdd.n895 39.2114
R17856 vdd.n2423 vdd.n896 39.2114
R17857 vdd.n2419 vdd.n897 39.2114
R17858 vdd.n2415 vdd.n898 39.2114
R17859 vdd.n2411 vdd.n899 39.2114
R17860 vdd.n2407 vdd.n900 39.2114
R17861 vdd.n2403 vdd.n901 39.2114
R17862 vdd.n2399 vdd.n902 39.2114
R17863 vdd.n2395 vdd.n903 39.2114
R17864 vdd.n2391 vdd.n904 39.2114
R17865 vdd.n2387 vdd.n905 39.2114
R17866 vdd.n2383 vdd.n906 39.2114
R17867 vdd.n2286 vdd.n1023 39.2114
R17868 vdd.n2285 vdd.n2284 39.2114
R17869 vdd.n2278 vdd.n1025 39.2114
R17870 vdd.n2277 vdd.n2276 39.2114
R17871 vdd.n2270 vdd.n1027 39.2114
R17872 vdd.n2269 vdd.n2268 39.2114
R17873 vdd.n2262 vdd.n1029 39.2114
R17874 vdd.n2261 vdd.n2260 39.2114
R17875 vdd.n1032 vdd.n1031 39.2114
R17876 vdd.n2102 vdd.n2101 39.2114
R17877 vdd.n2107 vdd.n2106 39.2114
R17878 vdd.n2110 vdd.n2109 39.2114
R17879 vdd.n2115 vdd.n2114 39.2114
R17880 vdd.n2118 vdd.n2117 39.2114
R17881 vdd.n2123 vdd.n2122 39.2114
R17882 vdd.n2126 vdd.n2125 39.2114
R17883 vdd.n2132 vdd.n2131 39.2114
R17884 vdd.n2380 vdd.n906 39.2114
R17885 vdd.n2384 vdd.n905 39.2114
R17886 vdd.n2388 vdd.n904 39.2114
R17887 vdd.n2392 vdd.n903 39.2114
R17888 vdd.n2396 vdd.n902 39.2114
R17889 vdd.n2400 vdd.n901 39.2114
R17890 vdd.n2404 vdd.n900 39.2114
R17891 vdd.n2408 vdd.n899 39.2114
R17892 vdd.n2412 vdd.n898 39.2114
R17893 vdd.n2416 vdd.n897 39.2114
R17894 vdd.n2420 vdd.n896 39.2114
R17895 vdd.n2424 vdd.n895 39.2114
R17896 vdd.n2428 vdd.n894 39.2114
R17897 vdd.n2432 vdd.n893 39.2114
R17898 vdd.n2436 vdd.n892 39.2114
R17899 vdd.n2440 vdd.n891 39.2114
R17900 vdd.n2444 vdd.n890 39.2114
R17901 vdd.n2287 vdd.n2286 39.2114
R17902 vdd.n2284 vdd.n2283 39.2114
R17903 vdd.n2279 vdd.n2278 39.2114
R17904 vdd.n2276 vdd.n2275 39.2114
R17905 vdd.n2271 vdd.n2270 39.2114
R17906 vdd.n2268 vdd.n2267 39.2114
R17907 vdd.n2263 vdd.n2262 39.2114
R17908 vdd.n2260 vdd.n2259 39.2114
R17909 vdd.n1033 vdd.n1032 39.2114
R17910 vdd.n2103 vdd.n2102 39.2114
R17911 vdd.n2108 vdd.n2107 39.2114
R17912 vdd.n2109 vdd.n2099 39.2114
R17913 vdd.n2116 vdd.n2115 39.2114
R17914 vdd.n2117 vdd.n2097 39.2114
R17915 vdd.n2124 vdd.n2123 39.2114
R17916 vdd.n2125 vdd.n2093 39.2114
R17917 vdd.n2133 vdd.n2132 39.2114
R17918 vdd.n2252 vdd.n2251 37.2369
R17919 vdd.n1955 vdd.n1888 37.2369
R17920 vdd.n1994 vdd.n1848 37.2369
R17921 vdd.n3059 vdd.n724 37.2369
R17922 vdd.n688 vdd.n687 37.2369
R17923 vdd.n3015 vdd.n3014 37.2369
R17924 vdd.n2294 vdd.n1018 31.6883
R17925 vdd.n2519 vdd.n927 31.6883
R17926 vdd.n2452 vdd.n930 31.6883
R17927 vdd.n2198 vdd.n2195 31.6883
R17928 vdd.n2706 vdd.n2704 31.6883
R17929 vdd.n2913 vdd.n2910 31.6883
R17930 vdd.n2783 vdd.n883 31.6883
R17931 vdd.n2974 vdd.n2973 31.6883
R17932 vdd.n2893 vdd.n2892 31.6883
R17933 vdd.n2979 vdd.n771 31.6883
R17934 vdd.n2625 vdd.n2624 31.6883
R17935 vdd.n2779 vdd.n2778 31.6883
R17936 vdd.n2290 vdd.n2289 31.6883
R17937 vdd.n2447 vdd.n2446 31.6883
R17938 vdd.n2379 vdd.n2378 31.6883
R17939 vdd.n2136 vdd.n2135 31.6883
R17940 vdd.n2129 vdd.n2095 30.449
R17941 vdd.n938 vdd.n937 30.449
R17942 vdd.n2070 vdd.n2069 30.449
R17943 vdd.n2457 vdd.n929 30.449
R17944 vdd.n2561 vdd.n2560 30.449
R17945 vdd.n806 vdd.n805 30.449
R17946 vdd.n2711 vdd.n2557 30.449
R17947 vdd.n770 vdd.n769 30.449
R17948 vdd.n1380 vdd.n1146 19.3944
R17949 vdd.n1380 vdd.n1136 19.3944
R17950 vdd.n1392 vdd.n1136 19.3944
R17951 vdd.n1392 vdd.n1134 19.3944
R17952 vdd.n1396 vdd.n1134 19.3944
R17953 vdd.n1396 vdd.n1124 19.3944
R17954 vdd.n1409 vdd.n1124 19.3944
R17955 vdd.n1409 vdd.n1122 19.3944
R17956 vdd.n1413 vdd.n1122 19.3944
R17957 vdd.n1413 vdd.n1114 19.3944
R17958 vdd.n1426 vdd.n1114 19.3944
R17959 vdd.n1426 vdd.n1112 19.3944
R17960 vdd.n1430 vdd.n1112 19.3944
R17961 vdd.n1430 vdd.n1101 19.3944
R17962 vdd.n1442 vdd.n1101 19.3944
R17963 vdd.n1442 vdd.n1099 19.3944
R17964 vdd.n1446 vdd.n1099 19.3944
R17965 vdd.n1446 vdd.n1090 19.3944
R17966 vdd.n1754 vdd.n1090 19.3944
R17967 vdd.n1754 vdd.n1088 19.3944
R17968 vdd.n1758 vdd.n1088 19.3944
R17969 vdd.n1758 vdd.n1079 19.3944
R17970 vdd.n1770 vdd.n1079 19.3944
R17971 vdd.n1770 vdd.n1077 19.3944
R17972 vdd.n1774 vdd.n1077 19.3944
R17973 vdd.n1774 vdd.n1067 19.3944
R17974 vdd.n1787 vdd.n1067 19.3944
R17975 vdd.n1787 vdd.n1065 19.3944
R17976 vdd.n1791 vdd.n1065 19.3944
R17977 vdd.n1791 vdd.n1057 19.3944
R17978 vdd.n1804 vdd.n1057 19.3944
R17979 vdd.n1804 vdd.n1054 19.3944
R17980 vdd.n1810 vdd.n1054 19.3944
R17981 vdd.n1810 vdd.n1055 19.3944
R17982 vdd.n1055 vdd.n1043 19.3944
R17983 vdd.n1299 vdd.n1241 19.3944
R17984 vdd.n1299 vdd.n1298 19.3944
R17985 vdd.n1298 vdd.n1297 19.3944
R17986 vdd.n1297 vdd.n1247 19.3944
R17987 vdd.n1293 vdd.n1247 19.3944
R17988 vdd.n1293 vdd.n1292 19.3944
R17989 vdd.n1292 vdd.n1291 19.3944
R17990 vdd.n1291 vdd.n1253 19.3944
R17991 vdd.n1287 vdd.n1253 19.3944
R17992 vdd.n1287 vdd.n1286 19.3944
R17993 vdd.n1286 vdd.n1285 19.3944
R17994 vdd.n1285 vdd.n1259 19.3944
R17995 vdd.n1281 vdd.n1259 19.3944
R17996 vdd.n1281 vdd.n1280 19.3944
R17997 vdd.n1280 vdd.n1279 19.3944
R17998 vdd.n1279 vdd.n1265 19.3944
R17999 vdd.n1275 vdd.n1265 19.3944
R18000 vdd.n1275 vdd.n1274 19.3944
R18001 vdd.n1274 vdd.n1273 19.3944
R18002 vdd.n1273 vdd.n1271 19.3944
R18003 vdd.n1337 vdd.n1336 19.3944
R18004 vdd.n1336 vdd.n1212 19.3944
R18005 vdd.n1332 vdd.n1212 19.3944
R18006 vdd.n1332 vdd.n1331 19.3944
R18007 vdd.n1331 vdd.n1330 19.3944
R18008 vdd.n1330 vdd.n1218 19.3944
R18009 vdd.n1326 vdd.n1218 19.3944
R18010 vdd.n1326 vdd.n1325 19.3944
R18011 vdd.n1325 vdd.n1324 19.3944
R18012 vdd.n1324 vdd.n1224 19.3944
R18013 vdd.n1320 vdd.n1224 19.3944
R18014 vdd.n1320 vdd.n1319 19.3944
R18015 vdd.n1319 vdd.n1318 19.3944
R18016 vdd.n1318 vdd.n1230 19.3944
R18017 vdd.n1314 vdd.n1230 19.3944
R18018 vdd.n1314 vdd.n1313 19.3944
R18019 vdd.n1313 vdd.n1312 19.3944
R18020 vdd.n1312 vdd.n1236 19.3944
R18021 vdd.n1308 vdd.n1236 19.3944
R18022 vdd.n1308 vdd.n1307 19.3944
R18023 vdd.n1371 vdd.n1370 19.3944
R18024 vdd.n1370 vdd.n1185 19.3944
R18025 vdd.n1366 vdd.n1185 19.3944
R18026 vdd.n1366 vdd.n1365 19.3944
R18027 vdd.n1365 vdd.n1364 19.3944
R18028 vdd.n1364 vdd.n1190 19.3944
R18029 vdd.n1360 vdd.n1190 19.3944
R18030 vdd.n1360 vdd.n1359 19.3944
R18031 vdd.n1359 vdd.n1358 19.3944
R18032 vdd.n1358 vdd.n1196 19.3944
R18033 vdd.n1354 vdd.n1196 19.3944
R18034 vdd.n1354 vdd.n1353 19.3944
R18035 vdd.n1353 vdd.n1352 19.3944
R18036 vdd.n1352 vdd.n1202 19.3944
R18037 vdd.n1348 vdd.n1202 19.3944
R18038 vdd.n1348 vdd.n1347 19.3944
R18039 vdd.n1347 vdd.n1346 19.3944
R18040 vdd.n1346 vdd.n1208 19.3944
R18041 vdd.n1951 vdd.n1886 19.3944
R18042 vdd.n1951 vdd.n1892 19.3944
R18043 vdd.n1946 vdd.n1892 19.3944
R18044 vdd.n1946 vdd.n1945 19.3944
R18045 vdd.n1945 vdd.n1944 19.3944
R18046 vdd.n1944 vdd.n1899 19.3944
R18047 vdd.n1939 vdd.n1899 19.3944
R18048 vdd.n1939 vdd.n1938 19.3944
R18049 vdd.n1938 vdd.n1937 19.3944
R18050 vdd.n1937 vdd.n1906 19.3944
R18051 vdd.n1932 vdd.n1906 19.3944
R18052 vdd.n1932 vdd.n1931 19.3944
R18053 vdd.n1931 vdd.n1930 19.3944
R18054 vdd.n1930 vdd.n1914 19.3944
R18055 vdd.n1925 vdd.n1914 19.3944
R18056 vdd.n1925 vdd.n1924 19.3944
R18057 vdd.n1920 vdd.n1919 19.3944
R18058 vdd.n2253 vdd.n1039 19.3944
R18059 vdd.n1990 vdd.n1846 19.3944
R18060 vdd.n1990 vdd.n1852 19.3944
R18061 vdd.n1985 vdd.n1852 19.3944
R18062 vdd.n1985 vdd.n1984 19.3944
R18063 vdd.n1984 vdd.n1983 19.3944
R18064 vdd.n1983 vdd.n1859 19.3944
R18065 vdd.n1978 vdd.n1859 19.3944
R18066 vdd.n1978 vdd.n1977 19.3944
R18067 vdd.n1977 vdd.n1976 19.3944
R18068 vdd.n1976 vdd.n1866 19.3944
R18069 vdd.n1971 vdd.n1866 19.3944
R18070 vdd.n1971 vdd.n1970 19.3944
R18071 vdd.n1970 vdd.n1969 19.3944
R18072 vdd.n1969 vdd.n1873 19.3944
R18073 vdd.n1964 vdd.n1873 19.3944
R18074 vdd.n1964 vdd.n1963 19.3944
R18075 vdd.n1963 vdd.n1962 19.3944
R18076 vdd.n1962 vdd.n1880 19.3944
R18077 vdd.n1957 vdd.n1880 19.3944
R18078 vdd.n1957 vdd.n1956 19.3944
R18079 vdd.n2241 vdd.n2240 19.3944
R18080 vdd.n2240 vdd.n1818 19.3944
R18081 vdd.n2235 vdd.n2234 19.3944
R18082 vdd.n2017 vdd.n1822 19.3944
R18083 vdd.n2017 vdd.n1824 19.3944
R18084 vdd.n1827 vdd.n1824 19.3944
R18085 vdd.n2010 vdd.n1827 19.3944
R18086 vdd.n2010 vdd.n2009 19.3944
R18087 vdd.n2009 vdd.n2008 19.3944
R18088 vdd.n2008 vdd.n1833 19.3944
R18089 vdd.n2003 vdd.n1833 19.3944
R18090 vdd.n2003 vdd.n2002 19.3944
R18091 vdd.n2002 vdd.n2001 19.3944
R18092 vdd.n2001 vdd.n1840 19.3944
R18093 vdd.n1996 vdd.n1840 19.3944
R18094 vdd.n1996 vdd.n1995 19.3944
R18095 vdd.n1384 vdd.n1142 19.3944
R18096 vdd.n1384 vdd.n1140 19.3944
R18097 vdd.n1388 vdd.n1140 19.3944
R18098 vdd.n1388 vdd.n1130 19.3944
R18099 vdd.n1401 vdd.n1130 19.3944
R18100 vdd.n1401 vdd.n1128 19.3944
R18101 vdd.n1405 vdd.n1128 19.3944
R18102 vdd.n1405 vdd.n1119 19.3944
R18103 vdd.n1418 vdd.n1119 19.3944
R18104 vdd.n1418 vdd.n1117 19.3944
R18105 vdd.n1422 vdd.n1117 19.3944
R18106 vdd.n1422 vdd.n1108 19.3944
R18107 vdd.n1434 vdd.n1108 19.3944
R18108 vdd.n1434 vdd.n1106 19.3944
R18109 vdd.n1438 vdd.n1106 19.3944
R18110 vdd.n1438 vdd.n1096 19.3944
R18111 vdd.n1451 vdd.n1096 19.3944
R18112 vdd.n1451 vdd.n1094 19.3944
R18113 vdd.n1750 vdd.n1094 19.3944
R18114 vdd.n1750 vdd.n1085 19.3944
R18115 vdd.n1762 vdd.n1085 19.3944
R18116 vdd.n1762 vdd.n1083 19.3944
R18117 vdd.n1766 vdd.n1083 19.3944
R18118 vdd.n1766 vdd.n1073 19.3944
R18119 vdd.n1779 vdd.n1073 19.3944
R18120 vdd.n1779 vdd.n1071 19.3944
R18121 vdd.n1783 vdd.n1071 19.3944
R18122 vdd.n1783 vdd.n1062 19.3944
R18123 vdd.n1796 vdd.n1062 19.3944
R18124 vdd.n1796 vdd.n1060 19.3944
R18125 vdd.n1800 vdd.n1060 19.3944
R18126 vdd.n1800 vdd.n1050 19.3944
R18127 vdd.n1814 vdd.n1050 19.3944
R18128 vdd.n1814 vdd.n1048 19.3944
R18129 vdd.n2244 vdd.n1048 19.3944
R18130 vdd.n3147 vdd.n655 19.3944
R18131 vdd.n3151 vdd.n655 19.3944
R18132 vdd.n3151 vdd.n646 19.3944
R18133 vdd.n3163 vdd.n646 19.3944
R18134 vdd.n3163 vdd.n644 19.3944
R18135 vdd.n3167 vdd.n644 19.3944
R18136 vdd.n3167 vdd.n633 19.3944
R18137 vdd.n3179 vdd.n633 19.3944
R18138 vdd.n3179 vdd.n631 19.3944
R18139 vdd.n3183 vdd.n631 19.3944
R18140 vdd.n3183 vdd.n622 19.3944
R18141 vdd.n3196 vdd.n622 19.3944
R18142 vdd.n3196 vdd.n620 19.3944
R18143 vdd.n3203 vdd.n620 19.3944
R18144 vdd.n3203 vdd.n3202 19.3944
R18145 vdd.n3202 vdd.n610 19.3944
R18146 vdd.n3216 vdd.n610 19.3944
R18147 vdd.n3217 vdd.n3216 19.3944
R18148 vdd.n3218 vdd.n3217 19.3944
R18149 vdd.n3218 vdd.n608 19.3944
R18150 vdd.n3223 vdd.n608 19.3944
R18151 vdd.n3224 vdd.n3223 19.3944
R18152 vdd.n3225 vdd.n3224 19.3944
R18153 vdd.n3225 vdd.n606 19.3944
R18154 vdd.n3230 vdd.n606 19.3944
R18155 vdd.n3231 vdd.n3230 19.3944
R18156 vdd.n3232 vdd.n3231 19.3944
R18157 vdd.n3232 vdd.n604 19.3944
R18158 vdd.n3238 vdd.n604 19.3944
R18159 vdd.n3239 vdd.n3238 19.3944
R18160 vdd.n3240 vdd.n3239 19.3944
R18161 vdd.n3240 vdd.n602 19.3944
R18162 vdd.n3245 vdd.n602 19.3944
R18163 vdd.n3246 vdd.n3245 19.3944
R18164 vdd.n3247 vdd.n3246 19.3944
R18165 vdd.n550 vdd.n417 19.3944
R18166 vdd.n556 vdd.n417 19.3944
R18167 vdd.n557 vdd.n556 19.3944
R18168 vdd.n560 vdd.n557 19.3944
R18169 vdd.n560 vdd.n415 19.3944
R18170 vdd.n566 vdd.n415 19.3944
R18171 vdd.n567 vdd.n566 19.3944
R18172 vdd.n570 vdd.n567 19.3944
R18173 vdd.n570 vdd.n413 19.3944
R18174 vdd.n576 vdd.n413 19.3944
R18175 vdd.n577 vdd.n576 19.3944
R18176 vdd.n580 vdd.n577 19.3944
R18177 vdd.n580 vdd.n411 19.3944
R18178 vdd.n586 vdd.n411 19.3944
R18179 vdd.n587 vdd.n586 19.3944
R18180 vdd.n590 vdd.n587 19.3944
R18181 vdd.n590 vdd.n409 19.3944
R18182 vdd.n596 vdd.n409 19.3944
R18183 vdd.n598 vdd.n596 19.3944
R18184 vdd.n599 vdd.n598 19.3944
R18185 vdd.n497 vdd.n496 19.3944
R18186 vdd.n500 vdd.n497 19.3944
R18187 vdd.n500 vdd.n429 19.3944
R18188 vdd.n506 vdd.n429 19.3944
R18189 vdd.n507 vdd.n506 19.3944
R18190 vdd.n510 vdd.n507 19.3944
R18191 vdd.n510 vdd.n427 19.3944
R18192 vdd.n516 vdd.n427 19.3944
R18193 vdd.n517 vdd.n516 19.3944
R18194 vdd.n520 vdd.n517 19.3944
R18195 vdd.n520 vdd.n425 19.3944
R18196 vdd.n526 vdd.n425 19.3944
R18197 vdd.n527 vdd.n526 19.3944
R18198 vdd.n530 vdd.n527 19.3944
R18199 vdd.n530 vdd.n423 19.3944
R18200 vdd.n536 vdd.n423 19.3944
R18201 vdd.n537 vdd.n536 19.3944
R18202 vdd.n540 vdd.n537 19.3944
R18203 vdd.n540 vdd.n421 19.3944
R18204 vdd.n546 vdd.n421 19.3944
R18205 vdd.n447 vdd.n446 19.3944
R18206 vdd.n450 vdd.n447 19.3944
R18207 vdd.n450 vdd.n441 19.3944
R18208 vdd.n456 vdd.n441 19.3944
R18209 vdd.n457 vdd.n456 19.3944
R18210 vdd.n460 vdd.n457 19.3944
R18211 vdd.n460 vdd.n439 19.3944
R18212 vdd.n466 vdd.n439 19.3944
R18213 vdd.n467 vdd.n466 19.3944
R18214 vdd.n470 vdd.n467 19.3944
R18215 vdd.n470 vdd.n437 19.3944
R18216 vdd.n476 vdd.n437 19.3944
R18217 vdd.n477 vdd.n476 19.3944
R18218 vdd.n480 vdd.n477 19.3944
R18219 vdd.n480 vdd.n435 19.3944
R18220 vdd.n486 vdd.n435 19.3944
R18221 vdd.n487 vdd.n486 19.3944
R18222 vdd.n490 vdd.n487 19.3944
R18223 vdd.n3143 vdd.n652 19.3944
R18224 vdd.n3155 vdd.n652 19.3944
R18225 vdd.n3155 vdd.n650 19.3944
R18226 vdd.n3159 vdd.n650 19.3944
R18227 vdd.n3159 vdd.n640 19.3944
R18228 vdd.n3171 vdd.n640 19.3944
R18229 vdd.n3171 vdd.n638 19.3944
R18230 vdd.n3175 vdd.n638 19.3944
R18231 vdd.n3175 vdd.n628 19.3944
R18232 vdd.n3188 vdd.n628 19.3944
R18233 vdd.n3188 vdd.n626 19.3944
R18234 vdd.n3192 vdd.n626 19.3944
R18235 vdd.n3192 vdd.n617 19.3944
R18236 vdd.n3207 vdd.n617 19.3944
R18237 vdd.n3207 vdd.n615 19.3944
R18238 vdd.n3211 vdd.n615 19.3944
R18239 vdd.n3211 vdd.n324 19.3944
R18240 vdd.n3289 vdd.n324 19.3944
R18241 vdd.n3289 vdd.n325 19.3944
R18242 vdd.n3283 vdd.n325 19.3944
R18243 vdd.n3283 vdd.n3282 19.3944
R18244 vdd.n3282 vdd.n3281 19.3944
R18245 vdd.n3281 vdd.n337 19.3944
R18246 vdd.n3275 vdd.n337 19.3944
R18247 vdd.n3275 vdd.n3274 19.3944
R18248 vdd.n3274 vdd.n3273 19.3944
R18249 vdd.n3273 vdd.n347 19.3944
R18250 vdd.n3267 vdd.n347 19.3944
R18251 vdd.n3267 vdd.n3266 19.3944
R18252 vdd.n3266 vdd.n3265 19.3944
R18253 vdd.n3265 vdd.n358 19.3944
R18254 vdd.n3259 vdd.n358 19.3944
R18255 vdd.n3259 vdd.n3258 19.3944
R18256 vdd.n3258 vdd.n3257 19.3944
R18257 vdd.n3257 vdd.n369 19.3944
R18258 vdd.n3100 vdd.n3099 19.3944
R18259 vdd.n3099 vdd.n3098 19.3944
R18260 vdd.n3098 vdd.n694 19.3944
R18261 vdd.n3092 vdd.n694 19.3944
R18262 vdd.n3092 vdd.n3091 19.3944
R18263 vdd.n3091 vdd.n3090 19.3944
R18264 vdd.n3090 vdd.n700 19.3944
R18265 vdd.n3084 vdd.n700 19.3944
R18266 vdd.n3084 vdd.n3083 19.3944
R18267 vdd.n3083 vdd.n3082 19.3944
R18268 vdd.n3082 vdd.n706 19.3944
R18269 vdd.n3076 vdd.n706 19.3944
R18270 vdd.n3076 vdd.n3075 19.3944
R18271 vdd.n3075 vdd.n3074 19.3944
R18272 vdd.n3074 vdd.n712 19.3944
R18273 vdd.n3068 vdd.n712 19.3944
R18274 vdd.n3068 vdd.n3067 19.3944
R18275 vdd.n3067 vdd.n3066 19.3944
R18276 vdd.n3066 vdd.n718 19.3944
R18277 vdd.n3060 vdd.n718 19.3944
R18278 vdd.n3140 vdd.n3139 19.3944
R18279 vdd.n3139 vdd.n662 19.3944
R18280 vdd.n3134 vdd.n3133 19.3944
R18281 vdd.n3130 vdd.n3129 19.3944
R18282 vdd.n3129 vdd.n668 19.3944
R18283 vdd.n3124 vdd.n668 19.3944
R18284 vdd.n3124 vdd.n3123 19.3944
R18285 vdd.n3123 vdd.n3122 19.3944
R18286 vdd.n3122 vdd.n674 19.3944
R18287 vdd.n3116 vdd.n674 19.3944
R18288 vdd.n3116 vdd.n3115 19.3944
R18289 vdd.n3115 vdd.n3114 19.3944
R18290 vdd.n3114 vdd.n680 19.3944
R18291 vdd.n3108 vdd.n680 19.3944
R18292 vdd.n3108 vdd.n3107 19.3944
R18293 vdd.n3107 vdd.n3106 19.3944
R18294 vdd.n3055 vdd.n722 19.3944
R18295 vdd.n3055 vdd.n726 19.3944
R18296 vdd.n3050 vdd.n726 19.3944
R18297 vdd.n3050 vdd.n3049 19.3944
R18298 vdd.n3049 vdd.n732 19.3944
R18299 vdd.n3044 vdd.n732 19.3944
R18300 vdd.n3044 vdd.n3043 19.3944
R18301 vdd.n3043 vdd.n3042 19.3944
R18302 vdd.n3042 vdd.n738 19.3944
R18303 vdd.n3036 vdd.n738 19.3944
R18304 vdd.n3036 vdd.n3035 19.3944
R18305 vdd.n3035 vdd.n3034 19.3944
R18306 vdd.n3034 vdd.n744 19.3944
R18307 vdd.n3028 vdd.n744 19.3944
R18308 vdd.n3028 vdd.n3027 19.3944
R18309 vdd.n3027 vdd.n3026 19.3944
R18310 vdd.n3022 vdd.n3021 19.3944
R18311 vdd.n3018 vdd.n3017 19.3944
R18312 vdd.n1306 vdd.n1241 19.0066
R18313 vdd.n1955 vdd.n1886 19.0066
R18314 vdd.n550 vdd.n547 19.0066
R18315 vdd.n3059 vdd.n722 19.0066
R18316 vdd.n1374 vdd.n1144 18.5924
R18317 vdd.n2246 vdd.n1045 18.5924
R18318 vdd.n3145 vdd.n658 18.5924
R18319 vdd.n3254 vdd.n3253 18.5924
R18320 vdd.n2095 vdd.n2094 16.0975
R18321 vdd.n937 vdd.n936 16.0975
R18322 vdd.n1149 vdd.n1148 16.0975
R18323 vdd.n1305 vdd.n1304 16.0975
R18324 vdd.n1341 vdd.n1340 16.0975
R18325 vdd.n2251 vdd.n2250 16.0975
R18326 vdd.n1888 vdd.n1887 16.0975
R18327 vdd.n1848 vdd.n1847 16.0975
R18328 vdd.n2069 vdd.n2068 16.0975
R18329 vdd.n929 vdd.n928 16.0975
R18330 vdd.n2560 vdd.n2559 16.0975
R18331 vdd.n406 vdd.n405 16.0975
R18332 vdd.n420 vdd.n419 16.0975
R18333 vdd.n432 vdd.n431 16.0975
R18334 vdd.n724 vdd.n723 16.0975
R18335 vdd.n687 vdd.n686 16.0975
R18336 vdd.n805 vdd.n804 16.0975
R18337 vdd.n2557 vdd.n2556 16.0975
R18338 vdd.n3014 vdd.n3013 16.0975
R18339 vdd.n769 vdd.n768 16.0975
R18340 vdd.t157 vdd.n2521 15.4182
R18341 vdd.n2774 vdd.t160 15.4182
R18342 vdd.n28 vdd.n27 14.5238
R18343 vdd.n2292 vdd.n1020 14.5112
R18344 vdd.n2976 vdd.n756 14.5112
R18345 vdd.n316 vdd.n281 13.1884
R18346 vdd.n261 vdd.n226 13.1884
R18347 vdd.n218 vdd.n183 13.1884
R18348 vdd.n163 vdd.n128 13.1884
R18349 vdd.n121 vdd.n86 13.1884
R18350 vdd.n66 vdd.n31 13.1884
R18351 vdd.n1685 vdd.n1650 13.1884
R18352 vdd.n1740 vdd.n1705 13.1884
R18353 vdd.n1587 vdd.n1552 13.1884
R18354 vdd.n1642 vdd.n1607 13.1884
R18355 vdd.n1490 vdd.n1455 13.1884
R18356 vdd.n1545 vdd.n1510 13.1884
R18357 vdd.n1342 vdd.n1337 12.9944
R18358 vdd.n1342 vdd.n1208 12.9944
R18359 vdd.n1994 vdd.n1846 12.9944
R18360 vdd.n1995 vdd.n1994 12.9944
R18361 vdd.n496 vdd.n433 12.9944
R18362 vdd.n490 vdd.n433 12.9944
R18363 vdd.n3100 vdd.n688 12.9944
R18364 vdd.n3106 vdd.n688 12.9944
R18365 vdd.n317 vdd.n279 12.8005
R18366 vdd.n312 vdd.n283 12.8005
R18367 vdd.n262 vdd.n224 12.8005
R18368 vdd.n257 vdd.n228 12.8005
R18369 vdd.n219 vdd.n181 12.8005
R18370 vdd.n214 vdd.n185 12.8005
R18371 vdd.n164 vdd.n126 12.8005
R18372 vdd.n159 vdd.n130 12.8005
R18373 vdd.n122 vdd.n84 12.8005
R18374 vdd.n117 vdd.n88 12.8005
R18375 vdd.n67 vdd.n29 12.8005
R18376 vdd.n62 vdd.n33 12.8005
R18377 vdd.n1686 vdd.n1648 12.8005
R18378 vdd.n1681 vdd.n1652 12.8005
R18379 vdd.n1741 vdd.n1703 12.8005
R18380 vdd.n1736 vdd.n1707 12.8005
R18381 vdd.n1588 vdd.n1550 12.8005
R18382 vdd.n1583 vdd.n1554 12.8005
R18383 vdd.n1643 vdd.n1605 12.8005
R18384 vdd.n1638 vdd.n1609 12.8005
R18385 vdd.n1491 vdd.n1453 12.8005
R18386 vdd.n1486 vdd.n1457 12.8005
R18387 vdd.n1546 vdd.n1508 12.8005
R18388 vdd.n1541 vdd.n1512 12.8005
R18389 vdd.n311 vdd.n284 12.0247
R18390 vdd.n256 vdd.n229 12.0247
R18391 vdd.n213 vdd.n186 12.0247
R18392 vdd.n158 vdd.n131 12.0247
R18393 vdd.n116 vdd.n89 12.0247
R18394 vdd.n61 vdd.n34 12.0247
R18395 vdd.n1680 vdd.n1653 12.0247
R18396 vdd.n1735 vdd.n1708 12.0247
R18397 vdd.n1582 vdd.n1555 12.0247
R18398 vdd.n1637 vdd.n1610 12.0247
R18399 vdd.n1485 vdd.n1458 12.0247
R18400 vdd.n1540 vdd.n1513 12.0247
R18401 vdd.n1382 vdd.n1144 11.337
R18402 vdd.n1390 vdd.n1138 11.337
R18403 vdd.n1390 vdd.n1132 11.337
R18404 vdd.n1399 vdd.n1132 11.337
R18405 vdd.n1407 vdd.n1126 11.337
R18406 vdd.n1416 vdd.n1415 11.337
R18407 vdd.n1432 vdd.n1110 11.337
R18408 vdd.n1440 vdd.n1103 11.337
R18409 vdd.n1449 vdd.n1448 11.337
R18410 vdd.n1752 vdd.n1092 11.337
R18411 vdd.n1768 vdd.n1081 11.337
R18412 vdd.n1777 vdd.n1075 11.337
R18413 vdd.n1785 vdd.n1069 11.337
R18414 vdd.n1794 vdd.n1793 11.337
R18415 vdd.n1802 vdd.n1052 11.337
R18416 vdd.n1812 vdd.n1052 11.337
R18417 vdd.n2246 vdd.n1044 11.337
R18418 vdd.n3145 vdd.n659 11.337
R18419 vdd.n3153 vdd.n648 11.337
R18420 vdd.n3161 vdd.n648 11.337
R18421 vdd.n3169 vdd.n642 11.337
R18422 vdd.n3177 vdd.n635 11.337
R18423 vdd.n3186 vdd.n3185 11.337
R18424 vdd.n3194 vdd.n624 11.337
R18425 vdd.n3213 vdd.n613 11.337
R18426 vdd.n3287 vdd.n328 11.337
R18427 vdd.n3285 vdd.n332 11.337
R18428 vdd.n3279 vdd.n3278 11.337
R18429 vdd.n3271 vdd.n349 11.337
R18430 vdd.n3270 vdd.n3269 11.337
R18431 vdd.n3263 vdd.n3262 11.337
R18432 vdd.n3262 vdd.n3261 11.337
R18433 vdd.n3261 vdd.n363 11.337
R18434 vdd.n3255 vdd.n3254 11.337
R18435 vdd.n308 vdd.n307 11.249
R18436 vdd.n253 vdd.n252 11.249
R18437 vdd.n210 vdd.n209 11.249
R18438 vdd.n155 vdd.n154 11.249
R18439 vdd.n113 vdd.n112 11.249
R18440 vdd.n58 vdd.n57 11.249
R18441 vdd.n1677 vdd.n1676 11.249
R18442 vdd.n1732 vdd.n1731 11.249
R18443 vdd.n1579 vdd.n1578 11.249
R18444 vdd.n1634 vdd.n1633 11.249
R18445 vdd.n1482 vdd.n1481 11.249
R18446 vdd.n1537 vdd.n1536 11.249
R18447 vdd.n2449 vdd.t260 11.1103
R18448 vdd.n2781 vdd.t258 11.1103
R18449 vdd.n1802 vdd.t11 10.7702
R18450 vdd.n3161 vdd.t13 10.7702
R18451 vdd.n293 vdd.n292 10.7238
R18452 vdd.n238 vdd.n237 10.7238
R18453 vdd.n195 vdd.n194 10.7238
R18454 vdd.n140 vdd.n139 10.7238
R18455 vdd.n98 vdd.n97 10.7238
R18456 vdd.n43 vdd.n42 10.7238
R18457 vdd.n1662 vdd.n1661 10.7238
R18458 vdd.n1717 vdd.n1716 10.7238
R18459 vdd.n1564 vdd.n1563 10.7238
R18460 vdd.n1619 vdd.n1618 10.7238
R18461 vdd.n1467 vdd.n1466 10.7238
R18462 vdd.n1522 vdd.n1521 10.7238
R18463 vdd.n2295 vdd.n2294 10.6151
R18464 vdd.n2296 vdd.n2295 10.6151
R18465 vdd.n2296 vdd.n1006 10.6151
R18466 vdd.n2306 vdd.n1006 10.6151
R18467 vdd.n2307 vdd.n2306 10.6151
R18468 vdd.n2308 vdd.n2307 10.6151
R18469 vdd.n2308 vdd.n993 10.6151
R18470 vdd.n2319 vdd.n993 10.6151
R18471 vdd.n2320 vdd.n2319 10.6151
R18472 vdd.n2321 vdd.n2320 10.6151
R18473 vdd.n2321 vdd.n981 10.6151
R18474 vdd.n2331 vdd.n981 10.6151
R18475 vdd.n2332 vdd.n2331 10.6151
R18476 vdd.n2333 vdd.n2332 10.6151
R18477 vdd.n2333 vdd.n969 10.6151
R18478 vdd.n2343 vdd.n969 10.6151
R18479 vdd.n2344 vdd.n2343 10.6151
R18480 vdd.n2345 vdd.n2344 10.6151
R18481 vdd.n2345 vdd.n958 10.6151
R18482 vdd.n2355 vdd.n958 10.6151
R18483 vdd.n2356 vdd.n2355 10.6151
R18484 vdd.n2357 vdd.n2356 10.6151
R18485 vdd.n2357 vdd.n945 10.6151
R18486 vdd.n2369 vdd.n945 10.6151
R18487 vdd.n2370 vdd.n2369 10.6151
R18488 vdd.n2372 vdd.n2370 10.6151
R18489 vdd.n2372 vdd.n2371 10.6151
R18490 vdd.n2371 vdd.n927 10.6151
R18491 vdd.n2519 vdd.n2518 10.6151
R18492 vdd.n2518 vdd.n2517 10.6151
R18493 vdd.n2517 vdd.n2514 10.6151
R18494 vdd.n2514 vdd.n2513 10.6151
R18495 vdd.n2513 vdd.n2510 10.6151
R18496 vdd.n2510 vdd.n2509 10.6151
R18497 vdd.n2509 vdd.n2506 10.6151
R18498 vdd.n2506 vdd.n2505 10.6151
R18499 vdd.n2505 vdd.n2502 10.6151
R18500 vdd.n2502 vdd.n2501 10.6151
R18501 vdd.n2501 vdd.n2498 10.6151
R18502 vdd.n2498 vdd.n2497 10.6151
R18503 vdd.n2497 vdd.n2494 10.6151
R18504 vdd.n2494 vdd.n2493 10.6151
R18505 vdd.n2493 vdd.n2490 10.6151
R18506 vdd.n2490 vdd.n2489 10.6151
R18507 vdd.n2489 vdd.n2486 10.6151
R18508 vdd.n2486 vdd.n2485 10.6151
R18509 vdd.n2485 vdd.n2482 10.6151
R18510 vdd.n2482 vdd.n2481 10.6151
R18511 vdd.n2481 vdd.n2478 10.6151
R18512 vdd.n2478 vdd.n2477 10.6151
R18513 vdd.n2477 vdd.n2474 10.6151
R18514 vdd.n2474 vdd.n2473 10.6151
R18515 vdd.n2473 vdd.n2470 10.6151
R18516 vdd.n2470 vdd.n2469 10.6151
R18517 vdd.n2469 vdd.n2466 10.6151
R18518 vdd.n2466 vdd.n2465 10.6151
R18519 vdd.n2465 vdd.n2462 10.6151
R18520 vdd.n2462 vdd.n2461 10.6151
R18521 vdd.n2461 vdd.n2458 10.6151
R18522 vdd.n2456 vdd.n2453 10.6151
R18523 vdd.n2453 vdd.n2452 10.6151
R18524 vdd.n2195 vdd.n2194 10.6151
R18525 vdd.n2194 vdd.n2192 10.6151
R18526 vdd.n2192 vdd.n2191 10.6151
R18527 vdd.n2191 vdd.n2189 10.6151
R18528 vdd.n2189 vdd.n2188 10.6151
R18529 vdd.n2188 vdd.n2186 10.6151
R18530 vdd.n2186 vdd.n2185 10.6151
R18531 vdd.n2185 vdd.n2183 10.6151
R18532 vdd.n2183 vdd.n2182 10.6151
R18533 vdd.n2182 vdd.n2180 10.6151
R18534 vdd.n2180 vdd.n2179 10.6151
R18535 vdd.n2179 vdd.n2177 10.6151
R18536 vdd.n2177 vdd.n2176 10.6151
R18537 vdd.n2176 vdd.n2091 10.6151
R18538 vdd.n2091 vdd.n2090 10.6151
R18539 vdd.n2090 vdd.n2088 10.6151
R18540 vdd.n2088 vdd.n2087 10.6151
R18541 vdd.n2087 vdd.n2085 10.6151
R18542 vdd.n2085 vdd.n2084 10.6151
R18543 vdd.n2084 vdd.n2082 10.6151
R18544 vdd.n2082 vdd.n2081 10.6151
R18545 vdd.n2081 vdd.n2079 10.6151
R18546 vdd.n2079 vdd.n2078 10.6151
R18547 vdd.n2078 vdd.n2076 10.6151
R18548 vdd.n2076 vdd.n2075 10.6151
R18549 vdd.n2075 vdd.n2072 10.6151
R18550 vdd.n2072 vdd.n2071 10.6151
R18551 vdd.n2071 vdd.n930 10.6151
R18552 vdd.n2029 vdd.n1018 10.6151
R18553 vdd.n2030 vdd.n2029 10.6151
R18554 vdd.n2031 vdd.n2030 10.6151
R18555 vdd.n2031 vdd.n2025 10.6151
R18556 vdd.n2037 vdd.n2025 10.6151
R18557 vdd.n2038 vdd.n2037 10.6151
R18558 vdd.n2039 vdd.n2038 10.6151
R18559 vdd.n2039 vdd.n2023 10.6151
R18560 vdd.n2045 vdd.n2023 10.6151
R18561 vdd.n2046 vdd.n2045 10.6151
R18562 vdd.n2047 vdd.n2046 10.6151
R18563 vdd.n2047 vdd.n2021 10.6151
R18564 vdd.n2053 vdd.n2021 10.6151
R18565 vdd.n2054 vdd.n2053 10.6151
R18566 vdd.n2055 vdd.n2054 10.6151
R18567 vdd.n2055 vdd.n2019 10.6151
R18568 vdd.n2231 vdd.n2019 10.6151
R18569 vdd.n2231 vdd.n2230 10.6151
R18570 vdd.n2230 vdd.n2060 10.6151
R18571 vdd.n2224 vdd.n2060 10.6151
R18572 vdd.n2224 vdd.n2223 10.6151
R18573 vdd.n2223 vdd.n2222 10.6151
R18574 vdd.n2222 vdd.n2062 10.6151
R18575 vdd.n2216 vdd.n2062 10.6151
R18576 vdd.n2216 vdd.n2215 10.6151
R18577 vdd.n2215 vdd.n2214 10.6151
R18578 vdd.n2214 vdd.n2064 10.6151
R18579 vdd.n2208 vdd.n2064 10.6151
R18580 vdd.n2208 vdd.n2207 10.6151
R18581 vdd.n2207 vdd.n2206 10.6151
R18582 vdd.n2206 vdd.n2066 10.6151
R18583 vdd.n2200 vdd.n2199 10.6151
R18584 vdd.n2199 vdd.n2198 10.6151
R18585 vdd.n2704 vdd.n2703 10.6151
R18586 vdd.n2703 vdd.n2701 10.6151
R18587 vdd.n2701 vdd.n2700 10.6151
R18588 vdd.n2700 vdd.n2558 10.6151
R18589 vdd.n2647 vdd.n2558 10.6151
R18590 vdd.n2648 vdd.n2647 10.6151
R18591 vdd.n2650 vdd.n2648 10.6151
R18592 vdd.n2651 vdd.n2650 10.6151
R18593 vdd.n2653 vdd.n2651 10.6151
R18594 vdd.n2654 vdd.n2653 10.6151
R18595 vdd.n2656 vdd.n2654 10.6151
R18596 vdd.n2657 vdd.n2656 10.6151
R18597 vdd.n2659 vdd.n2657 10.6151
R18598 vdd.n2660 vdd.n2659 10.6151
R18599 vdd.n2675 vdd.n2660 10.6151
R18600 vdd.n2675 vdd.n2674 10.6151
R18601 vdd.n2674 vdd.n2673 10.6151
R18602 vdd.n2673 vdd.n2671 10.6151
R18603 vdd.n2671 vdd.n2670 10.6151
R18604 vdd.n2670 vdd.n2668 10.6151
R18605 vdd.n2668 vdd.n2667 10.6151
R18606 vdd.n2667 vdd.n2665 10.6151
R18607 vdd.n2665 vdd.n2664 10.6151
R18608 vdd.n2664 vdd.n2662 10.6151
R18609 vdd.n2662 vdd.n2661 10.6151
R18610 vdd.n2661 vdd.n807 10.6151
R18611 vdd.n2909 vdd.n807 10.6151
R18612 vdd.n2910 vdd.n2909 10.6151
R18613 vdd.n2771 vdd.n883 10.6151
R18614 vdd.n2771 vdd.n2770 10.6151
R18615 vdd.n2770 vdd.n2769 10.6151
R18616 vdd.n2769 vdd.n2767 10.6151
R18617 vdd.n2767 vdd.n2764 10.6151
R18618 vdd.n2764 vdd.n2763 10.6151
R18619 vdd.n2763 vdd.n2760 10.6151
R18620 vdd.n2760 vdd.n2759 10.6151
R18621 vdd.n2759 vdd.n2756 10.6151
R18622 vdd.n2756 vdd.n2755 10.6151
R18623 vdd.n2755 vdd.n2752 10.6151
R18624 vdd.n2752 vdd.n2751 10.6151
R18625 vdd.n2751 vdd.n2748 10.6151
R18626 vdd.n2748 vdd.n2747 10.6151
R18627 vdd.n2747 vdd.n2744 10.6151
R18628 vdd.n2744 vdd.n2743 10.6151
R18629 vdd.n2743 vdd.n2740 10.6151
R18630 vdd.n2740 vdd.n2739 10.6151
R18631 vdd.n2739 vdd.n2736 10.6151
R18632 vdd.n2736 vdd.n2735 10.6151
R18633 vdd.n2735 vdd.n2732 10.6151
R18634 vdd.n2732 vdd.n2731 10.6151
R18635 vdd.n2731 vdd.n2728 10.6151
R18636 vdd.n2728 vdd.n2727 10.6151
R18637 vdd.n2727 vdd.n2724 10.6151
R18638 vdd.n2724 vdd.n2723 10.6151
R18639 vdd.n2723 vdd.n2720 10.6151
R18640 vdd.n2720 vdd.n2719 10.6151
R18641 vdd.n2719 vdd.n2716 10.6151
R18642 vdd.n2716 vdd.n2715 10.6151
R18643 vdd.n2715 vdd.n2712 10.6151
R18644 vdd.n2710 vdd.n2707 10.6151
R18645 vdd.n2707 vdd.n2706 10.6151
R18646 vdd.n2784 vdd.n2783 10.6151
R18647 vdd.n2785 vdd.n2784 10.6151
R18648 vdd.n2785 vdd.n873 10.6151
R18649 vdd.n2795 vdd.n873 10.6151
R18650 vdd.n2796 vdd.n2795 10.6151
R18651 vdd.n2797 vdd.n2796 10.6151
R18652 vdd.n2797 vdd.n860 10.6151
R18653 vdd.n2807 vdd.n860 10.6151
R18654 vdd.n2808 vdd.n2807 10.6151
R18655 vdd.n2809 vdd.n2808 10.6151
R18656 vdd.n2809 vdd.n849 10.6151
R18657 vdd.n2819 vdd.n849 10.6151
R18658 vdd.n2820 vdd.n2819 10.6151
R18659 vdd.n2821 vdd.n2820 10.6151
R18660 vdd.n2821 vdd.n837 10.6151
R18661 vdd.n2831 vdd.n837 10.6151
R18662 vdd.n2832 vdd.n2831 10.6151
R18663 vdd.n2833 vdd.n2832 10.6151
R18664 vdd.n2833 vdd.n826 10.6151
R18665 vdd.n2845 vdd.n826 10.6151
R18666 vdd.n2846 vdd.n2845 10.6151
R18667 vdd.n2847 vdd.n2846 10.6151
R18668 vdd.n2847 vdd.n812 10.6151
R18669 vdd.n2902 vdd.n812 10.6151
R18670 vdd.n2903 vdd.n2902 10.6151
R18671 vdd.n2904 vdd.n2903 10.6151
R18672 vdd.n2904 vdd.n779 10.6151
R18673 vdd.n2974 vdd.n779 10.6151
R18674 vdd.n2973 vdd.n2972 10.6151
R18675 vdd.n2972 vdd.n780 10.6151
R18676 vdd.n781 vdd.n780 10.6151
R18677 vdd.n2965 vdd.n781 10.6151
R18678 vdd.n2965 vdd.n2964 10.6151
R18679 vdd.n2964 vdd.n2963 10.6151
R18680 vdd.n2963 vdd.n783 10.6151
R18681 vdd.n2958 vdd.n783 10.6151
R18682 vdd.n2958 vdd.n2957 10.6151
R18683 vdd.n2957 vdd.n2956 10.6151
R18684 vdd.n2956 vdd.n786 10.6151
R18685 vdd.n2951 vdd.n786 10.6151
R18686 vdd.n2951 vdd.n2950 10.6151
R18687 vdd.n2950 vdd.n2949 10.6151
R18688 vdd.n2949 vdd.n789 10.6151
R18689 vdd.n2944 vdd.n789 10.6151
R18690 vdd.n2944 vdd.n2943 10.6151
R18691 vdd.n2943 vdd.n2941 10.6151
R18692 vdd.n2941 vdd.n792 10.6151
R18693 vdd.n2936 vdd.n792 10.6151
R18694 vdd.n2936 vdd.n2935 10.6151
R18695 vdd.n2935 vdd.n2934 10.6151
R18696 vdd.n2934 vdd.n795 10.6151
R18697 vdd.n2929 vdd.n795 10.6151
R18698 vdd.n2929 vdd.n2928 10.6151
R18699 vdd.n2928 vdd.n2927 10.6151
R18700 vdd.n2927 vdd.n798 10.6151
R18701 vdd.n2922 vdd.n798 10.6151
R18702 vdd.n2922 vdd.n2921 10.6151
R18703 vdd.n2921 vdd.n2920 10.6151
R18704 vdd.n2920 vdd.n801 10.6151
R18705 vdd.n2915 vdd.n2914 10.6151
R18706 vdd.n2914 vdd.n2913 10.6151
R18707 vdd.n2892 vdd.n2853 10.6151
R18708 vdd.n2887 vdd.n2853 10.6151
R18709 vdd.n2887 vdd.n2886 10.6151
R18710 vdd.n2886 vdd.n2885 10.6151
R18711 vdd.n2885 vdd.n2855 10.6151
R18712 vdd.n2880 vdd.n2855 10.6151
R18713 vdd.n2880 vdd.n2879 10.6151
R18714 vdd.n2879 vdd.n2878 10.6151
R18715 vdd.n2878 vdd.n2858 10.6151
R18716 vdd.n2873 vdd.n2858 10.6151
R18717 vdd.n2873 vdd.n2872 10.6151
R18718 vdd.n2872 vdd.n2871 10.6151
R18719 vdd.n2871 vdd.n2861 10.6151
R18720 vdd.n2866 vdd.n2861 10.6151
R18721 vdd.n2866 vdd.n2865 10.6151
R18722 vdd.n2865 vdd.n753 10.6151
R18723 vdd.n3009 vdd.n753 10.6151
R18724 vdd.n3009 vdd.n754 10.6151
R18725 vdd.n757 vdd.n754 10.6151
R18726 vdd.n3002 vdd.n757 10.6151
R18727 vdd.n3002 vdd.n3001 10.6151
R18728 vdd.n3001 vdd.n3000 10.6151
R18729 vdd.n3000 vdd.n759 10.6151
R18730 vdd.n2995 vdd.n759 10.6151
R18731 vdd.n2995 vdd.n2994 10.6151
R18732 vdd.n2994 vdd.n2993 10.6151
R18733 vdd.n2993 vdd.n762 10.6151
R18734 vdd.n2988 vdd.n762 10.6151
R18735 vdd.n2988 vdd.n2987 10.6151
R18736 vdd.n2987 vdd.n2986 10.6151
R18737 vdd.n2986 vdd.n765 10.6151
R18738 vdd.n2981 vdd.n2980 10.6151
R18739 vdd.n2980 vdd.n2979 10.6151
R18740 vdd.n2627 vdd.n2625 10.6151
R18741 vdd.n2628 vdd.n2627 10.6151
R18742 vdd.n2696 vdd.n2628 10.6151
R18743 vdd.n2696 vdd.n2695 10.6151
R18744 vdd.n2695 vdd.n2694 10.6151
R18745 vdd.n2694 vdd.n2692 10.6151
R18746 vdd.n2692 vdd.n2691 10.6151
R18747 vdd.n2691 vdd.n2689 10.6151
R18748 vdd.n2689 vdd.n2688 10.6151
R18749 vdd.n2688 vdd.n2686 10.6151
R18750 vdd.n2686 vdd.n2685 10.6151
R18751 vdd.n2685 vdd.n2683 10.6151
R18752 vdd.n2683 vdd.n2682 10.6151
R18753 vdd.n2682 vdd.n2680 10.6151
R18754 vdd.n2680 vdd.n2679 10.6151
R18755 vdd.n2679 vdd.n2645 10.6151
R18756 vdd.n2645 vdd.n2644 10.6151
R18757 vdd.n2644 vdd.n2642 10.6151
R18758 vdd.n2642 vdd.n2641 10.6151
R18759 vdd.n2641 vdd.n2639 10.6151
R18760 vdd.n2639 vdd.n2638 10.6151
R18761 vdd.n2638 vdd.n2636 10.6151
R18762 vdd.n2636 vdd.n2635 10.6151
R18763 vdd.n2635 vdd.n2633 10.6151
R18764 vdd.n2633 vdd.n2632 10.6151
R18765 vdd.n2632 vdd.n2630 10.6151
R18766 vdd.n2630 vdd.n2629 10.6151
R18767 vdd.n2629 vdd.n771 10.6151
R18768 vdd.n2778 vdd.n2777 10.6151
R18769 vdd.n2777 vdd.n888 10.6151
R18770 vdd.n2562 vdd.n888 10.6151
R18771 vdd.n2565 vdd.n2562 10.6151
R18772 vdd.n2566 vdd.n2565 10.6151
R18773 vdd.n2569 vdd.n2566 10.6151
R18774 vdd.n2570 vdd.n2569 10.6151
R18775 vdd.n2573 vdd.n2570 10.6151
R18776 vdd.n2574 vdd.n2573 10.6151
R18777 vdd.n2577 vdd.n2574 10.6151
R18778 vdd.n2578 vdd.n2577 10.6151
R18779 vdd.n2581 vdd.n2578 10.6151
R18780 vdd.n2582 vdd.n2581 10.6151
R18781 vdd.n2585 vdd.n2582 10.6151
R18782 vdd.n2586 vdd.n2585 10.6151
R18783 vdd.n2589 vdd.n2586 10.6151
R18784 vdd.n2590 vdd.n2589 10.6151
R18785 vdd.n2593 vdd.n2590 10.6151
R18786 vdd.n2594 vdd.n2593 10.6151
R18787 vdd.n2597 vdd.n2594 10.6151
R18788 vdd.n2598 vdd.n2597 10.6151
R18789 vdd.n2601 vdd.n2598 10.6151
R18790 vdd.n2602 vdd.n2601 10.6151
R18791 vdd.n2605 vdd.n2602 10.6151
R18792 vdd.n2606 vdd.n2605 10.6151
R18793 vdd.n2609 vdd.n2606 10.6151
R18794 vdd.n2610 vdd.n2609 10.6151
R18795 vdd.n2613 vdd.n2610 10.6151
R18796 vdd.n2614 vdd.n2613 10.6151
R18797 vdd.n2617 vdd.n2614 10.6151
R18798 vdd.n2618 vdd.n2617 10.6151
R18799 vdd.n2623 vdd.n2621 10.6151
R18800 vdd.n2624 vdd.n2623 10.6151
R18801 vdd.n2779 vdd.n878 10.6151
R18802 vdd.n2789 vdd.n878 10.6151
R18803 vdd.n2790 vdd.n2789 10.6151
R18804 vdd.n2791 vdd.n2790 10.6151
R18805 vdd.n2791 vdd.n866 10.6151
R18806 vdd.n2801 vdd.n866 10.6151
R18807 vdd.n2802 vdd.n2801 10.6151
R18808 vdd.n2803 vdd.n2802 10.6151
R18809 vdd.n2803 vdd.n855 10.6151
R18810 vdd.n2813 vdd.n855 10.6151
R18811 vdd.n2814 vdd.n2813 10.6151
R18812 vdd.n2815 vdd.n2814 10.6151
R18813 vdd.n2815 vdd.n843 10.6151
R18814 vdd.n2825 vdd.n843 10.6151
R18815 vdd.n2826 vdd.n2825 10.6151
R18816 vdd.n2827 vdd.n2826 10.6151
R18817 vdd.n2827 vdd.n832 10.6151
R18818 vdd.n2837 vdd.n832 10.6151
R18819 vdd.n2838 vdd.n2837 10.6151
R18820 vdd.n2841 vdd.n2838 10.6151
R18821 vdd.n2851 vdd.n820 10.6151
R18822 vdd.n2852 vdd.n2851 10.6151
R18823 vdd.n2898 vdd.n2852 10.6151
R18824 vdd.n2898 vdd.n2897 10.6151
R18825 vdd.n2897 vdd.n2896 10.6151
R18826 vdd.n2896 vdd.n2895 10.6151
R18827 vdd.n2895 vdd.n2893 10.6151
R18828 vdd.n2290 vdd.n1012 10.6151
R18829 vdd.n2300 vdd.n1012 10.6151
R18830 vdd.n2301 vdd.n2300 10.6151
R18831 vdd.n2302 vdd.n2301 10.6151
R18832 vdd.n2302 vdd.n999 10.6151
R18833 vdd.n2312 vdd.n999 10.6151
R18834 vdd.n2313 vdd.n2312 10.6151
R18835 vdd.n2315 vdd.n987 10.6151
R18836 vdd.n2325 vdd.n987 10.6151
R18837 vdd.n2326 vdd.n2325 10.6151
R18838 vdd.n2327 vdd.n2326 10.6151
R18839 vdd.n2327 vdd.n975 10.6151
R18840 vdd.n2337 vdd.n975 10.6151
R18841 vdd.n2338 vdd.n2337 10.6151
R18842 vdd.n2339 vdd.n2338 10.6151
R18843 vdd.n2339 vdd.n964 10.6151
R18844 vdd.n2349 vdd.n964 10.6151
R18845 vdd.n2350 vdd.n2349 10.6151
R18846 vdd.n2351 vdd.n2350 10.6151
R18847 vdd.n2351 vdd.n952 10.6151
R18848 vdd.n2361 vdd.n952 10.6151
R18849 vdd.n2362 vdd.n2361 10.6151
R18850 vdd.n2365 vdd.n2362 10.6151
R18851 vdd.n2365 vdd.n2364 10.6151
R18852 vdd.n2364 vdd.n2363 10.6151
R18853 vdd.n2363 vdd.n935 10.6151
R18854 vdd.n2447 vdd.n935 10.6151
R18855 vdd.n2446 vdd.n2445 10.6151
R18856 vdd.n2445 vdd.n2442 10.6151
R18857 vdd.n2442 vdd.n2441 10.6151
R18858 vdd.n2441 vdd.n2438 10.6151
R18859 vdd.n2438 vdd.n2437 10.6151
R18860 vdd.n2437 vdd.n2434 10.6151
R18861 vdd.n2434 vdd.n2433 10.6151
R18862 vdd.n2433 vdd.n2430 10.6151
R18863 vdd.n2430 vdd.n2429 10.6151
R18864 vdd.n2429 vdd.n2426 10.6151
R18865 vdd.n2426 vdd.n2425 10.6151
R18866 vdd.n2425 vdd.n2422 10.6151
R18867 vdd.n2422 vdd.n2421 10.6151
R18868 vdd.n2421 vdd.n2418 10.6151
R18869 vdd.n2418 vdd.n2417 10.6151
R18870 vdd.n2417 vdd.n2414 10.6151
R18871 vdd.n2414 vdd.n2413 10.6151
R18872 vdd.n2413 vdd.n2410 10.6151
R18873 vdd.n2410 vdd.n2409 10.6151
R18874 vdd.n2409 vdd.n2406 10.6151
R18875 vdd.n2406 vdd.n2405 10.6151
R18876 vdd.n2405 vdd.n2402 10.6151
R18877 vdd.n2402 vdd.n2401 10.6151
R18878 vdd.n2401 vdd.n2398 10.6151
R18879 vdd.n2398 vdd.n2397 10.6151
R18880 vdd.n2397 vdd.n2394 10.6151
R18881 vdd.n2394 vdd.n2393 10.6151
R18882 vdd.n2393 vdd.n2390 10.6151
R18883 vdd.n2390 vdd.n2389 10.6151
R18884 vdd.n2389 vdd.n2386 10.6151
R18885 vdd.n2386 vdd.n2385 10.6151
R18886 vdd.n2382 vdd.n2381 10.6151
R18887 vdd.n2381 vdd.n2379 10.6151
R18888 vdd.n2138 vdd.n2136 10.6151
R18889 vdd.n2139 vdd.n2138 10.6151
R18890 vdd.n2141 vdd.n2139 10.6151
R18891 vdd.n2142 vdd.n2141 10.6151
R18892 vdd.n2144 vdd.n2142 10.6151
R18893 vdd.n2145 vdd.n2144 10.6151
R18894 vdd.n2147 vdd.n2145 10.6151
R18895 vdd.n2148 vdd.n2147 10.6151
R18896 vdd.n2150 vdd.n2148 10.6151
R18897 vdd.n2151 vdd.n2150 10.6151
R18898 vdd.n2153 vdd.n2151 10.6151
R18899 vdd.n2154 vdd.n2153 10.6151
R18900 vdd.n2172 vdd.n2154 10.6151
R18901 vdd.n2172 vdd.n2171 10.6151
R18902 vdd.n2171 vdd.n2170 10.6151
R18903 vdd.n2170 vdd.n2168 10.6151
R18904 vdd.n2168 vdd.n2167 10.6151
R18905 vdd.n2167 vdd.n2165 10.6151
R18906 vdd.n2165 vdd.n2164 10.6151
R18907 vdd.n2164 vdd.n2162 10.6151
R18908 vdd.n2162 vdd.n2161 10.6151
R18909 vdd.n2161 vdd.n2159 10.6151
R18910 vdd.n2159 vdd.n2158 10.6151
R18911 vdd.n2158 vdd.n2156 10.6151
R18912 vdd.n2156 vdd.n2155 10.6151
R18913 vdd.n2155 vdd.n939 10.6151
R18914 vdd.n2377 vdd.n939 10.6151
R18915 vdd.n2378 vdd.n2377 10.6151
R18916 vdd.n2289 vdd.n2288 10.6151
R18917 vdd.n2288 vdd.n1024 10.6151
R18918 vdd.n2282 vdd.n1024 10.6151
R18919 vdd.n2282 vdd.n2281 10.6151
R18920 vdd.n2281 vdd.n2280 10.6151
R18921 vdd.n2280 vdd.n1026 10.6151
R18922 vdd.n2274 vdd.n1026 10.6151
R18923 vdd.n2274 vdd.n2273 10.6151
R18924 vdd.n2273 vdd.n2272 10.6151
R18925 vdd.n2272 vdd.n1028 10.6151
R18926 vdd.n2266 vdd.n1028 10.6151
R18927 vdd.n2266 vdd.n2265 10.6151
R18928 vdd.n2265 vdd.n2264 10.6151
R18929 vdd.n2264 vdd.n1030 10.6151
R18930 vdd.n2258 vdd.n1030 10.6151
R18931 vdd.n2258 vdd.n2257 10.6151
R18932 vdd.n2257 vdd.n2256 10.6151
R18933 vdd.n2256 vdd.n1034 10.6151
R18934 vdd.n2104 vdd.n1034 10.6151
R18935 vdd.n2105 vdd.n2104 10.6151
R18936 vdd.n2105 vdd.n2100 10.6151
R18937 vdd.n2111 vdd.n2100 10.6151
R18938 vdd.n2112 vdd.n2111 10.6151
R18939 vdd.n2113 vdd.n2112 10.6151
R18940 vdd.n2113 vdd.n2098 10.6151
R18941 vdd.n2119 vdd.n2098 10.6151
R18942 vdd.n2120 vdd.n2119 10.6151
R18943 vdd.n2121 vdd.n2120 10.6151
R18944 vdd.n2121 vdd.n2096 10.6151
R18945 vdd.n2127 vdd.n2096 10.6151
R18946 vdd.n2128 vdd.n2127 10.6151
R18947 vdd.n2130 vdd.n2092 10.6151
R18948 vdd.n2135 vdd.n2092 10.6151
R18949 vdd.t98 vdd.n1776 10.5435
R18950 vdd.n636 vdd.t17 10.5435
R18951 vdd.n304 vdd.n286 10.4732
R18952 vdd.n249 vdd.n231 10.4732
R18953 vdd.n206 vdd.n188 10.4732
R18954 vdd.n151 vdd.n133 10.4732
R18955 vdd.n109 vdd.n91 10.4732
R18956 vdd.n54 vdd.n36 10.4732
R18957 vdd.n1673 vdd.n1655 10.4732
R18958 vdd.n1728 vdd.n1710 10.4732
R18959 vdd.n1575 vdd.n1557 10.4732
R18960 vdd.n1630 vdd.n1612 10.4732
R18961 vdd.n1478 vdd.n1460 10.4732
R18962 vdd.n1533 vdd.n1515 10.4732
R18963 vdd.n1760 vdd.t66 10.3167
R18964 vdd.n3205 vdd.t35 10.3167
R18965 vdd.t19 vdd.n1104 10.09
R18966 vdd.n1812 vdd.t196 10.09
R18967 vdd.n3153 vdd.t181 10.09
R18968 vdd.n3286 vdd.t21 10.09
R18969 vdd.n1424 vdd.t42 9.86327
R18970 vdd.n3277 vdd.t76 9.86327
R18971 vdd.n303 vdd.n288 9.69747
R18972 vdd.n248 vdd.n233 9.69747
R18973 vdd.n205 vdd.n190 9.69747
R18974 vdd.n150 vdd.n135 9.69747
R18975 vdd.n108 vdd.n93 9.69747
R18976 vdd.n53 vdd.n38 9.69747
R18977 vdd.n1672 vdd.n1657 9.69747
R18978 vdd.n1727 vdd.n1712 9.69747
R18979 vdd.n1574 vdd.n1559 9.69747
R18980 vdd.n1629 vdd.n1614 9.69747
R18981 vdd.n1477 vdd.n1462 9.69747
R18982 vdd.n1532 vdd.n1517 9.69747
R18983 vdd.n2232 vdd.n2231 9.67831
R18984 vdd.n2943 vdd.n2942 9.67831
R18985 vdd.n3010 vdd.n3009 9.67831
R18986 vdd.n2256 vdd.n2255 9.67831
R18987 vdd.t23 vdd.n1398 9.63654
R18988 vdd.n3236 vdd.t33 9.63654
R18989 vdd.n319 vdd.n318 9.45567
R18990 vdd.n264 vdd.n263 9.45567
R18991 vdd.n221 vdd.n220 9.45567
R18992 vdd.n166 vdd.n165 9.45567
R18993 vdd.n124 vdd.n123 9.45567
R18994 vdd.n69 vdd.n68 9.45567
R18995 vdd.n1688 vdd.n1687 9.45567
R18996 vdd.n1743 vdd.n1742 9.45567
R18997 vdd.n1590 vdd.n1589 9.45567
R18998 vdd.n1645 vdd.n1644 9.45567
R18999 vdd.n1493 vdd.n1492 9.45567
R19000 vdd.n1548 vdd.n1547 9.45567
R19001 vdd.n1992 vdd.n1846 9.3005
R19002 vdd.n1991 vdd.n1990 9.3005
R19003 vdd.n1852 vdd.n1851 9.3005
R19004 vdd.n1985 vdd.n1856 9.3005
R19005 vdd.n1984 vdd.n1857 9.3005
R19006 vdd.n1983 vdd.n1858 9.3005
R19007 vdd.n1862 vdd.n1859 9.3005
R19008 vdd.n1978 vdd.n1863 9.3005
R19009 vdd.n1977 vdd.n1864 9.3005
R19010 vdd.n1976 vdd.n1865 9.3005
R19011 vdd.n1869 vdd.n1866 9.3005
R19012 vdd.n1971 vdd.n1870 9.3005
R19013 vdd.n1970 vdd.n1871 9.3005
R19014 vdd.n1969 vdd.n1872 9.3005
R19015 vdd.n1876 vdd.n1873 9.3005
R19016 vdd.n1964 vdd.n1877 9.3005
R19017 vdd.n1963 vdd.n1878 9.3005
R19018 vdd.n1962 vdd.n1879 9.3005
R19019 vdd.n1883 vdd.n1880 9.3005
R19020 vdd.n1957 vdd.n1884 9.3005
R19021 vdd.n1956 vdd.n1885 9.3005
R19022 vdd.n1955 vdd.n1954 9.3005
R19023 vdd.n1953 vdd.n1886 9.3005
R19024 vdd.n1952 vdd.n1951 9.3005
R19025 vdd.n1892 vdd.n1891 9.3005
R19026 vdd.n1946 vdd.n1896 9.3005
R19027 vdd.n1945 vdd.n1897 9.3005
R19028 vdd.n1944 vdd.n1898 9.3005
R19029 vdd.n1902 vdd.n1899 9.3005
R19030 vdd.n1939 vdd.n1903 9.3005
R19031 vdd.n1938 vdd.n1904 9.3005
R19032 vdd.n1937 vdd.n1905 9.3005
R19033 vdd.n1909 vdd.n1906 9.3005
R19034 vdd.n1932 vdd.n1910 9.3005
R19035 vdd.n1931 vdd.n1911 9.3005
R19036 vdd.n1930 vdd.n1912 9.3005
R19037 vdd.n1914 vdd.n1913 9.3005
R19038 vdd.n1925 vdd.n1035 9.3005
R19039 vdd.n1994 vdd.n1993 9.3005
R19040 vdd.n2018 vdd.n2017 9.3005
R19041 vdd.n1824 vdd.n1823 9.3005
R19042 vdd.n1829 vdd.n1827 9.3005
R19043 vdd.n2010 vdd.n1830 9.3005
R19044 vdd.n2009 vdd.n1831 9.3005
R19045 vdd.n2008 vdd.n1832 9.3005
R19046 vdd.n1836 vdd.n1833 9.3005
R19047 vdd.n2003 vdd.n1837 9.3005
R19048 vdd.n2002 vdd.n1838 9.3005
R19049 vdd.n2001 vdd.n1839 9.3005
R19050 vdd.n1843 vdd.n1840 9.3005
R19051 vdd.n1996 vdd.n1844 9.3005
R19052 vdd.n1995 vdd.n1845 9.3005
R19053 vdd.n2240 vdd.n1817 9.3005
R19054 vdd.n2242 vdd.n2241 9.3005
R19055 vdd.n1748 vdd.n1094 9.3005
R19056 vdd.n1750 vdd.n1749 9.3005
R19057 vdd.n1085 vdd.n1084 9.3005
R19058 vdd.n1763 vdd.n1762 9.3005
R19059 vdd.n1764 vdd.n1083 9.3005
R19060 vdd.n1766 vdd.n1765 9.3005
R19061 vdd.n1073 vdd.n1072 9.3005
R19062 vdd.n1780 vdd.n1779 9.3005
R19063 vdd.n1781 vdd.n1071 9.3005
R19064 vdd.n1783 vdd.n1782 9.3005
R19065 vdd.n1062 vdd.n1061 9.3005
R19066 vdd.n1797 vdd.n1796 9.3005
R19067 vdd.n1798 vdd.n1060 9.3005
R19068 vdd.n1800 vdd.n1799 9.3005
R19069 vdd.n1050 vdd.n1049 9.3005
R19070 vdd.n1815 vdd.n1814 9.3005
R19071 vdd.n1816 vdd.n1048 9.3005
R19072 vdd.n2244 vdd.n2243 9.3005
R19073 vdd.n295 vdd.n294 9.3005
R19074 vdd.n290 vdd.n289 9.3005
R19075 vdd.n301 vdd.n300 9.3005
R19076 vdd.n303 vdd.n302 9.3005
R19077 vdd.n286 vdd.n285 9.3005
R19078 vdd.n309 vdd.n308 9.3005
R19079 vdd.n311 vdd.n310 9.3005
R19080 vdd.n283 vdd.n280 9.3005
R19081 vdd.n318 vdd.n317 9.3005
R19082 vdd.n240 vdd.n239 9.3005
R19083 vdd.n235 vdd.n234 9.3005
R19084 vdd.n246 vdd.n245 9.3005
R19085 vdd.n248 vdd.n247 9.3005
R19086 vdd.n231 vdd.n230 9.3005
R19087 vdd.n254 vdd.n253 9.3005
R19088 vdd.n256 vdd.n255 9.3005
R19089 vdd.n228 vdd.n225 9.3005
R19090 vdd.n263 vdd.n262 9.3005
R19091 vdd.n197 vdd.n196 9.3005
R19092 vdd.n192 vdd.n191 9.3005
R19093 vdd.n203 vdd.n202 9.3005
R19094 vdd.n205 vdd.n204 9.3005
R19095 vdd.n188 vdd.n187 9.3005
R19096 vdd.n211 vdd.n210 9.3005
R19097 vdd.n213 vdd.n212 9.3005
R19098 vdd.n185 vdd.n182 9.3005
R19099 vdd.n220 vdd.n219 9.3005
R19100 vdd.n142 vdd.n141 9.3005
R19101 vdd.n137 vdd.n136 9.3005
R19102 vdd.n148 vdd.n147 9.3005
R19103 vdd.n150 vdd.n149 9.3005
R19104 vdd.n133 vdd.n132 9.3005
R19105 vdd.n156 vdd.n155 9.3005
R19106 vdd.n158 vdd.n157 9.3005
R19107 vdd.n130 vdd.n127 9.3005
R19108 vdd.n165 vdd.n164 9.3005
R19109 vdd.n100 vdd.n99 9.3005
R19110 vdd.n95 vdd.n94 9.3005
R19111 vdd.n106 vdd.n105 9.3005
R19112 vdd.n108 vdd.n107 9.3005
R19113 vdd.n91 vdd.n90 9.3005
R19114 vdd.n114 vdd.n113 9.3005
R19115 vdd.n116 vdd.n115 9.3005
R19116 vdd.n88 vdd.n85 9.3005
R19117 vdd.n123 vdd.n122 9.3005
R19118 vdd.n45 vdd.n44 9.3005
R19119 vdd.n40 vdd.n39 9.3005
R19120 vdd.n51 vdd.n50 9.3005
R19121 vdd.n53 vdd.n52 9.3005
R19122 vdd.n36 vdd.n35 9.3005
R19123 vdd.n59 vdd.n58 9.3005
R19124 vdd.n61 vdd.n60 9.3005
R19125 vdd.n33 vdd.n30 9.3005
R19126 vdd.n68 vdd.n67 9.3005
R19127 vdd.n3059 vdd.n3058 9.3005
R19128 vdd.n3060 vdd.n721 9.3005
R19129 vdd.n720 vdd.n718 9.3005
R19130 vdd.n3066 vdd.n717 9.3005
R19131 vdd.n3067 vdd.n716 9.3005
R19132 vdd.n3068 vdd.n715 9.3005
R19133 vdd.n714 vdd.n712 9.3005
R19134 vdd.n3074 vdd.n711 9.3005
R19135 vdd.n3075 vdd.n710 9.3005
R19136 vdd.n3076 vdd.n709 9.3005
R19137 vdd.n708 vdd.n706 9.3005
R19138 vdd.n3082 vdd.n705 9.3005
R19139 vdd.n3083 vdd.n704 9.3005
R19140 vdd.n3084 vdd.n703 9.3005
R19141 vdd.n702 vdd.n700 9.3005
R19142 vdd.n3090 vdd.n699 9.3005
R19143 vdd.n3091 vdd.n698 9.3005
R19144 vdd.n3092 vdd.n697 9.3005
R19145 vdd.n696 vdd.n694 9.3005
R19146 vdd.n3098 vdd.n693 9.3005
R19147 vdd.n3099 vdd.n692 9.3005
R19148 vdd.n3100 vdd.n691 9.3005
R19149 vdd.n690 vdd.n688 9.3005
R19150 vdd.n3106 vdd.n685 9.3005
R19151 vdd.n3107 vdd.n684 9.3005
R19152 vdd.n3108 vdd.n683 9.3005
R19153 vdd.n682 vdd.n680 9.3005
R19154 vdd.n3114 vdd.n679 9.3005
R19155 vdd.n3115 vdd.n678 9.3005
R19156 vdd.n3116 vdd.n677 9.3005
R19157 vdd.n676 vdd.n674 9.3005
R19158 vdd.n3122 vdd.n673 9.3005
R19159 vdd.n3123 vdd.n672 9.3005
R19160 vdd.n3124 vdd.n671 9.3005
R19161 vdd.n670 vdd.n668 9.3005
R19162 vdd.n3129 vdd.n667 9.3005
R19163 vdd.n3139 vdd.n661 9.3005
R19164 vdd.n3141 vdd.n3140 9.3005
R19165 vdd.n652 vdd.n651 9.3005
R19166 vdd.n3156 vdd.n3155 9.3005
R19167 vdd.n3157 vdd.n650 9.3005
R19168 vdd.n3159 vdd.n3158 9.3005
R19169 vdd.n640 vdd.n639 9.3005
R19170 vdd.n3172 vdd.n3171 9.3005
R19171 vdd.n3173 vdd.n638 9.3005
R19172 vdd.n3175 vdd.n3174 9.3005
R19173 vdd.n628 vdd.n627 9.3005
R19174 vdd.n3189 vdd.n3188 9.3005
R19175 vdd.n3190 vdd.n626 9.3005
R19176 vdd.n3192 vdd.n3191 9.3005
R19177 vdd.n617 vdd.n616 9.3005
R19178 vdd.n3208 vdd.n3207 9.3005
R19179 vdd.n3209 vdd.n615 9.3005
R19180 vdd.n3211 vdd.n3210 9.3005
R19181 vdd.n324 vdd.n322 9.3005
R19182 vdd.n3143 vdd.n3142 9.3005
R19183 vdd.n3290 vdd.n3289 9.3005
R19184 vdd.n325 vdd.n323 9.3005
R19185 vdd.n3283 vdd.n334 9.3005
R19186 vdd.n3282 vdd.n335 9.3005
R19187 vdd.n3281 vdd.n336 9.3005
R19188 vdd.n343 vdd.n337 9.3005
R19189 vdd.n3275 vdd.n344 9.3005
R19190 vdd.n3274 vdd.n345 9.3005
R19191 vdd.n3273 vdd.n346 9.3005
R19192 vdd.n354 vdd.n347 9.3005
R19193 vdd.n3267 vdd.n355 9.3005
R19194 vdd.n3266 vdd.n356 9.3005
R19195 vdd.n3265 vdd.n357 9.3005
R19196 vdd.n365 vdd.n358 9.3005
R19197 vdd.n3259 vdd.n366 9.3005
R19198 vdd.n3258 vdd.n367 9.3005
R19199 vdd.n3257 vdd.n368 9.3005
R19200 vdd.n443 vdd.n369 9.3005
R19201 vdd.n447 vdd.n442 9.3005
R19202 vdd.n451 vdd.n450 9.3005
R19203 vdd.n452 vdd.n441 9.3005
R19204 vdd.n456 vdd.n453 9.3005
R19205 vdd.n457 vdd.n440 9.3005
R19206 vdd.n461 vdd.n460 9.3005
R19207 vdd.n462 vdd.n439 9.3005
R19208 vdd.n466 vdd.n463 9.3005
R19209 vdd.n467 vdd.n438 9.3005
R19210 vdd.n471 vdd.n470 9.3005
R19211 vdd.n472 vdd.n437 9.3005
R19212 vdd.n476 vdd.n473 9.3005
R19213 vdd.n477 vdd.n436 9.3005
R19214 vdd.n481 vdd.n480 9.3005
R19215 vdd.n482 vdd.n435 9.3005
R19216 vdd.n486 vdd.n483 9.3005
R19217 vdd.n487 vdd.n434 9.3005
R19218 vdd.n491 vdd.n490 9.3005
R19219 vdd.n492 vdd.n433 9.3005
R19220 vdd.n496 vdd.n493 9.3005
R19221 vdd.n497 vdd.n430 9.3005
R19222 vdd.n501 vdd.n500 9.3005
R19223 vdd.n502 vdd.n429 9.3005
R19224 vdd.n506 vdd.n503 9.3005
R19225 vdd.n507 vdd.n428 9.3005
R19226 vdd.n511 vdd.n510 9.3005
R19227 vdd.n512 vdd.n427 9.3005
R19228 vdd.n516 vdd.n513 9.3005
R19229 vdd.n517 vdd.n426 9.3005
R19230 vdd.n521 vdd.n520 9.3005
R19231 vdd.n522 vdd.n425 9.3005
R19232 vdd.n526 vdd.n523 9.3005
R19233 vdd.n527 vdd.n424 9.3005
R19234 vdd.n531 vdd.n530 9.3005
R19235 vdd.n532 vdd.n423 9.3005
R19236 vdd.n536 vdd.n533 9.3005
R19237 vdd.n537 vdd.n422 9.3005
R19238 vdd.n541 vdd.n540 9.3005
R19239 vdd.n542 vdd.n421 9.3005
R19240 vdd.n546 vdd.n543 9.3005
R19241 vdd.n547 vdd.n418 9.3005
R19242 vdd.n551 vdd.n550 9.3005
R19243 vdd.n552 vdd.n417 9.3005
R19244 vdd.n556 vdd.n553 9.3005
R19245 vdd.n557 vdd.n416 9.3005
R19246 vdd.n561 vdd.n560 9.3005
R19247 vdd.n562 vdd.n415 9.3005
R19248 vdd.n566 vdd.n563 9.3005
R19249 vdd.n567 vdd.n414 9.3005
R19250 vdd.n571 vdd.n570 9.3005
R19251 vdd.n572 vdd.n413 9.3005
R19252 vdd.n576 vdd.n573 9.3005
R19253 vdd.n577 vdd.n412 9.3005
R19254 vdd.n581 vdd.n580 9.3005
R19255 vdd.n582 vdd.n411 9.3005
R19256 vdd.n586 vdd.n583 9.3005
R19257 vdd.n587 vdd.n410 9.3005
R19258 vdd.n591 vdd.n590 9.3005
R19259 vdd.n592 vdd.n409 9.3005
R19260 vdd.n596 vdd.n593 9.3005
R19261 vdd.n598 vdd.n408 9.3005
R19262 vdd.n600 vdd.n599 9.3005
R19263 vdd.n3250 vdd.n3249 9.3005
R19264 vdd.n446 vdd.n444 9.3005
R19265 vdd.n3149 vdd.n655 9.3005
R19266 vdd.n3151 vdd.n3150 9.3005
R19267 vdd.n646 vdd.n645 9.3005
R19268 vdd.n3164 vdd.n3163 9.3005
R19269 vdd.n3165 vdd.n644 9.3005
R19270 vdd.n3167 vdd.n3166 9.3005
R19271 vdd.n633 vdd.n632 9.3005
R19272 vdd.n3180 vdd.n3179 9.3005
R19273 vdd.n3181 vdd.n631 9.3005
R19274 vdd.n3183 vdd.n3182 9.3005
R19275 vdd.n622 vdd.n621 9.3005
R19276 vdd.n3197 vdd.n3196 9.3005
R19277 vdd.n3198 vdd.n620 9.3005
R19278 vdd.n3203 vdd.n3199 9.3005
R19279 vdd.n3202 vdd.n3201 9.3005
R19280 vdd.n3200 vdd.n610 9.3005
R19281 vdd.n3216 vdd.n611 9.3005
R19282 vdd.n3217 vdd.n609 9.3005
R19283 vdd.n3219 vdd.n3218 9.3005
R19284 vdd.n3220 vdd.n608 9.3005
R19285 vdd.n3223 vdd.n3221 9.3005
R19286 vdd.n3224 vdd.n607 9.3005
R19287 vdd.n3226 vdd.n3225 9.3005
R19288 vdd.n3227 vdd.n606 9.3005
R19289 vdd.n3230 vdd.n3228 9.3005
R19290 vdd.n3231 vdd.n605 9.3005
R19291 vdd.n3233 vdd.n3232 9.3005
R19292 vdd.n3234 vdd.n604 9.3005
R19293 vdd.n3238 vdd.n3235 9.3005
R19294 vdd.n3239 vdd.n603 9.3005
R19295 vdd.n3241 vdd.n3240 9.3005
R19296 vdd.n3242 vdd.n602 9.3005
R19297 vdd.n3245 vdd.n3243 9.3005
R19298 vdd.n3246 vdd.n601 9.3005
R19299 vdd.n3248 vdd.n3247 9.3005
R19300 vdd.n3148 vdd.n3147 9.3005
R19301 vdd.n3012 vdd.n656 9.3005
R19302 vdd.n3017 vdd.n3011 9.3005
R19303 vdd.n3027 vdd.n748 9.3005
R19304 vdd.n3028 vdd.n747 9.3005
R19305 vdd.n746 vdd.n744 9.3005
R19306 vdd.n3034 vdd.n743 9.3005
R19307 vdd.n3035 vdd.n742 9.3005
R19308 vdd.n3036 vdd.n741 9.3005
R19309 vdd.n740 vdd.n738 9.3005
R19310 vdd.n3042 vdd.n737 9.3005
R19311 vdd.n3043 vdd.n736 9.3005
R19312 vdd.n3044 vdd.n735 9.3005
R19313 vdd.n734 vdd.n732 9.3005
R19314 vdd.n3049 vdd.n731 9.3005
R19315 vdd.n3050 vdd.n730 9.3005
R19316 vdd.n726 vdd.n725 9.3005
R19317 vdd.n3056 vdd.n3055 9.3005
R19318 vdd.n3057 vdd.n722 9.3005
R19319 vdd.n2254 vdd.n2253 9.3005
R19320 vdd.n2249 vdd.n1038 9.3005
R19321 vdd.n1380 vdd.n1379 9.3005
R19322 vdd.n1136 vdd.n1135 9.3005
R19323 vdd.n1393 vdd.n1392 9.3005
R19324 vdd.n1394 vdd.n1134 9.3005
R19325 vdd.n1396 vdd.n1395 9.3005
R19326 vdd.n1124 vdd.n1123 9.3005
R19327 vdd.n1410 vdd.n1409 9.3005
R19328 vdd.n1411 vdd.n1122 9.3005
R19329 vdd.n1413 vdd.n1412 9.3005
R19330 vdd.n1114 vdd.n1113 9.3005
R19331 vdd.n1427 vdd.n1426 9.3005
R19332 vdd.n1428 vdd.n1112 9.3005
R19333 vdd.n1430 vdd.n1429 9.3005
R19334 vdd.n1101 vdd.n1100 9.3005
R19335 vdd.n1443 vdd.n1442 9.3005
R19336 vdd.n1444 vdd.n1099 9.3005
R19337 vdd.n1446 vdd.n1445 9.3005
R19338 vdd.n1090 vdd.n1089 9.3005
R19339 vdd.n1755 vdd.n1754 9.3005
R19340 vdd.n1756 vdd.n1088 9.3005
R19341 vdd.n1758 vdd.n1757 9.3005
R19342 vdd.n1079 vdd.n1078 9.3005
R19343 vdd.n1771 vdd.n1770 9.3005
R19344 vdd.n1772 vdd.n1077 9.3005
R19345 vdd.n1774 vdd.n1773 9.3005
R19346 vdd.n1067 vdd.n1066 9.3005
R19347 vdd.n1788 vdd.n1787 9.3005
R19348 vdd.n1789 vdd.n1065 9.3005
R19349 vdd.n1791 vdd.n1790 9.3005
R19350 vdd.n1057 vdd.n1056 9.3005
R19351 vdd.n1805 vdd.n1804 9.3005
R19352 vdd.n1806 vdd.n1054 9.3005
R19353 vdd.n1810 vdd.n1809 9.3005
R19354 vdd.n1808 vdd.n1055 9.3005
R19355 vdd.n1807 vdd.n1043 9.3005
R19356 vdd.n1378 vdd.n1146 9.3005
R19357 vdd.n1271 vdd.n1147 9.3005
R19358 vdd.n1273 vdd.n1272 9.3005
R19359 vdd.n1274 vdd.n1266 9.3005
R19360 vdd.n1276 vdd.n1275 9.3005
R19361 vdd.n1277 vdd.n1265 9.3005
R19362 vdd.n1279 vdd.n1278 9.3005
R19363 vdd.n1280 vdd.n1260 9.3005
R19364 vdd.n1282 vdd.n1281 9.3005
R19365 vdd.n1283 vdd.n1259 9.3005
R19366 vdd.n1285 vdd.n1284 9.3005
R19367 vdd.n1286 vdd.n1254 9.3005
R19368 vdd.n1288 vdd.n1287 9.3005
R19369 vdd.n1289 vdd.n1253 9.3005
R19370 vdd.n1291 vdd.n1290 9.3005
R19371 vdd.n1292 vdd.n1248 9.3005
R19372 vdd.n1294 vdd.n1293 9.3005
R19373 vdd.n1295 vdd.n1247 9.3005
R19374 vdd.n1297 vdd.n1296 9.3005
R19375 vdd.n1298 vdd.n1242 9.3005
R19376 vdd.n1300 vdd.n1299 9.3005
R19377 vdd.n1301 vdd.n1241 9.3005
R19378 vdd.n1306 vdd.n1302 9.3005
R19379 vdd.n1307 vdd.n1237 9.3005
R19380 vdd.n1309 vdd.n1308 9.3005
R19381 vdd.n1310 vdd.n1236 9.3005
R19382 vdd.n1312 vdd.n1311 9.3005
R19383 vdd.n1313 vdd.n1231 9.3005
R19384 vdd.n1315 vdd.n1314 9.3005
R19385 vdd.n1316 vdd.n1230 9.3005
R19386 vdd.n1318 vdd.n1317 9.3005
R19387 vdd.n1319 vdd.n1225 9.3005
R19388 vdd.n1321 vdd.n1320 9.3005
R19389 vdd.n1322 vdd.n1224 9.3005
R19390 vdd.n1324 vdd.n1323 9.3005
R19391 vdd.n1325 vdd.n1219 9.3005
R19392 vdd.n1327 vdd.n1326 9.3005
R19393 vdd.n1328 vdd.n1218 9.3005
R19394 vdd.n1330 vdd.n1329 9.3005
R19395 vdd.n1331 vdd.n1213 9.3005
R19396 vdd.n1333 vdd.n1332 9.3005
R19397 vdd.n1334 vdd.n1212 9.3005
R19398 vdd.n1336 vdd.n1335 9.3005
R19399 vdd.n1337 vdd.n1209 9.3005
R19400 vdd.n1343 vdd.n1342 9.3005
R19401 vdd.n1344 vdd.n1208 9.3005
R19402 vdd.n1346 vdd.n1345 9.3005
R19403 vdd.n1347 vdd.n1203 9.3005
R19404 vdd.n1349 vdd.n1348 9.3005
R19405 vdd.n1350 vdd.n1202 9.3005
R19406 vdd.n1352 vdd.n1351 9.3005
R19407 vdd.n1353 vdd.n1197 9.3005
R19408 vdd.n1355 vdd.n1354 9.3005
R19409 vdd.n1356 vdd.n1196 9.3005
R19410 vdd.n1358 vdd.n1357 9.3005
R19411 vdd.n1359 vdd.n1191 9.3005
R19412 vdd.n1361 vdd.n1360 9.3005
R19413 vdd.n1362 vdd.n1190 9.3005
R19414 vdd.n1364 vdd.n1363 9.3005
R19415 vdd.n1365 vdd.n1186 9.3005
R19416 vdd.n1367 vdd.n1366 9.3005
R19417 vdd.n1368 vdd.n1185 9.3005
R19418 vdd.n1370 vdd.n1369 9.3005
R19419 vdd.n1371 vdd.n1184 9.3005
R19420 vdd.n1377 vdd.n1376 9.3005
R19421 vdd.n1385 vdd.n1384 9.3005
R19422 vdd.n1386 vdd.n1140 9.3005
R19423 vdd.n1388 vdd.n1387 9.3005
R19424 vdd.n1130 vdd.n1129 9.3005
R19425 vdd.n1402 vdd.n1401 9.3005
R19426 vdd.n1403 vdd.n1128 9.3005
R19427 vdd.n1405 vdd.n1404 9.3005
R19428 vdd.n1119 vdd.n1118 9.3005
R19429 vdd.n1419 vdd.n1418 9.3005
R19430 vdd.n1420 vdd.n1117 9.3005
R19431 vdd.n1422 vdd.n1421 9.3005
R19432 vdd.n1108 vdd.n1107 9.3005
R19433 vdd.n1435 vdd.n1434 9.3005
R19434 vdd.n1436 vdd.n1106 9.3005
R19435 vdd.n1438 vdd.n1437 9.3005
R19436 vdd.n1096 vdd.n1095 9.3005
R19437 vdd.n1452 vdd.n1451 9.3005
R19438 vdd.n1142 vdd.n1141 9.3005
R19439 vdd.n1664 vdd.n1663 9.3005
R19440 vdd.n1659 vdd.n1658 9.3005
R19441 vdd.n1670 vdd.n1669 9.3005
R19442 vdd.n1672 vdd.n1671 9.3005
R19443 vdd.n1655 vdd.n1654 9.3005
R19444 vdd.n1678 vdd.n1677 9.3005
R19445 vdd.n1680 vdd.n1679 9.3005
R19446 vdd.n1652 vdd.n1649 9.3005
R19447 vdd.n1687 vdd.n1686 9.3005
R19448 vdd.n1719 vdd.n1718 9.3005
R19449 vdd.n1714 vdd.n1713 9.3005
R19450 vdd.n1725 vdd.n1724 9.3005
R19451 vdd.n1727 vdd.n1726 9.3005
R19452 vdd.n1710 vdd.n1709 9.3005
R19453 vdd.n1733 vdd.n1732 9.3005
R19454 vdd.n1735 vdd.n1734 9.3005
R19455 vdd.n1707 vdd.n1704 9.3005
R19456 vdd.n1742 vdd.n1741 9.3005
R19457 vdd.n1566 vdd.n1565 9.3005
R19458 vdd.n1561 vdd.n1560 9.3005
R19459 vdd.n1572 vdd.n1571 9.3005
R19460 vdd.n1574 vdd.n1573 9.3005
R19461 vdd.n1557 vdd.n1556 9.3005
R19462 vdd.n1580 vdd.n1579 9.3005
R19463 vdd.n1582 vdd.n1581 9.3005
R19464 vdd.n1554 vdd.n1551 9.3005
R19465 vdd.n1589 vdd.n1588 9.3005
R19466 vdd.n1621 vdd.n1620 9.3005
R19467 vdd.n1616 vdd.n1615 9.3005
R19468 vdd.n1627 vdd.n1626 9.3005
R19469 vdd.n1629 vdd.n1628 9.3005
R19470 vdd.n1612 vdd.n1611 9.3005
R19471 vdd.n1635 vdd.n1634 9.3005
R19472 vdd.n1637 vdd.n1636 9.3005
R19473 vdd.n1609 vdd.n1606 9.3005
R19474 vdd.n1644 vdd.n1643 9.3005
R19475 vdd.n1469 vdd.n1468 9.3005
R19476 vdd.n1464 vdd.n1463 9.3005
R19477 vdd.n1475 vdd.n1474 9.3005
R19478 vdd.n1477 vdd.n1476 9.3005
R19479 vdd.n1460 vdd.n1459 9.3005
R19480 vdd.n1483 vdd.n1482 9.3005
R19481 vdd.n1485 vdd.n1484 9.3005
R19482 vdd.n1457 vdd.n1454 9.3005
R19483 vdd.n1492 vdd.n1491 9.3005
R19484 vdd.n1524 vdd.n1523 9.3005
R19485 vdd.n1519 vdd.n1518 9.3005
R19486 vdd.n1530 vdd.n1529 9.3005
R19487 vdd.n1532 vdd.n1531 9.3005
R19488 vdd.n1515 vdd.n1514 9.3005
R19489 vdd.n1538 vdd.n1537 9.3005
R19490 vdd.n1540 vdd.n1539 9.3005
R19491 vdd.n1512 vdd.n1509 9.3005
R19492 vdd.n1547 vdd.n1546 9.3005
R19493 vdd.n1398 vdd.t84 9.18308
R19494 vdd.n3236 vdd.t27 9.18308
R19495 vdd.n1424 vdd.t31 8.95635
R19496 vdd.t29 vdd.n3277 8.95635
R19497 vdd.n300 vdd.n299 8.92171
R19498 vdd.n245 vdd.n244 8.92171
R19499 vdd.n202 vdd.n201 8.92171
R19500 vdd.n147 vdd.n146 8.92171
R19501 vdd.n105 vdd.n104 8.92171
R19502 vdd.n50 vdd.n49 8.92171
R19503 vdd.n1669 vdd.n1668 8.92171
R19504 vdd.n1724 vdd.n1723 8.92171
R19505 vdd.n1571 vdd.n1570 8.92171
R19506 vdd.n1626 vdd.n1625 8.92171
R19507 vdd.n1474 vdd.n1473 8.92171
R19508 vdd.n1529 vdd.n1528 8.92171
R19509 vdd.n223 vdd.n125 8.81535
R19510 vdd.n1647 vdd.n1549 8.81535
R19511 vdd.n1104 vdd.t87 8.72962
R19512 vdd.t57 vdd.n3286 8.72962
R19513 vdd.n1760 vdd.t15 8.50289
R19514 vdd.n3205 vdd.t100 8.50289
R19515 vdd.n28 vdd.n14 8.42249
R19516 vdd.n1776 vdd.t25 8.27616
R19517 vdd.t74 vdd.n636 8.27616
R19518 vdd.n3292 vdd.n3291 8.16225
R19519 vdd.n1747 vdd.n1746 8.16225
R19520 vdd.n296 vdd.n290 8.14595
R19521 vdd.n241 vdd.n235 8.14595
R19522 vdd.n198 vdd.n192 8.14595
R19523 vdd.n143 vdd.n137 8.14595
R19524 vdd.n101 vdd.n95 8.14595
R19525 vdd.n46 vdd.n40 8.14595
R19526 vdd.n1665 vdd.n1659 8.14595
R19527 vdd.n1720 vdd.n1714 8.14595
R19528 vdd.n1567 vdd.n1561 8.14595
R19529 vdd.n1622 vdd.n1616 8.14595
R19530 vdd.n1470 vdd.n1464 8.14595
R19531 vdd.n1525 vdd.n1519 8.14595
R19532 vdd.n2840 vdd.n820 8.11757
R19533 vdd.n2314 vdd.n2313 8.11757
R19534 vdd.t185 vdd.n1138 7.8227
R19535 vdd.t189 vdd.n363 7.8227
R19536 vdd.n2292 vdd.n1014 7.70933
R19537 vdd.n2298 vdd.n1014 7.70933
R19538 vdd.n2304 vdd.n1008 7.70933
R19539 vdd.n2304 vdd.n1001 7.70933
R19540 vdd.n2310 vdd.n1001 7.70933
R19541 vdd.n2310 vdd.n1004 7.70933
R19542 vdd.n2317 vdd.n989 7.70933
R19543 vdd.n2323 vdd.n989 7.70933
R19544 vdd.n2329 vdd.n983 7.70933
R19545 vdd.n2335 vdd.n979 7.70933
R19546 vdd.n2341 vdd.n973 7.70933
R19547 vdd.n2353 vdd.n960 7.70933
R19548 vdd.n2359 vdd.n954 7.70933
R19549 vdd.n2359 vdd.n947 7.70933
R19550 vdd.n2367 vdd.n947 7.70933
R19551 vdd.n2374 vdd.t1 7.70933
R19552 vdd.n2449 vdd.t1 7.70933
R19553 vdd.n2781 vdd.t256 7.70933
R19554 vdd.n2787 vdd.t256 7.70933
R19555 vdd.n2793 vdd.n868 7.70933
R19556 vdd.n2799 vdd.n868 7.70933
R19557 vdd.n2799 vdd.n871 7.70933
R19558 vdd.n2805 vdd.n864 7.70933
R19559 vdd.n2817 vdd.n851 7.70933
R19560 vdd.n2823 vdd.n845 7.70933
R19561 vdd.n2829 vdd.n841 7.70933
R19562 vdd.n2835 vdd.n828 7.70933
R19563 vdd.n2843 vdd.n828 7.70933
R19564 vdd.n2849 vdd.n822 7.70933
R19565 vdd.n2849 vdd.n814 7.70933
R19566 vdd.n2900 vdd.n814 7.70933
R19567 vdd.n2900 vdd.n817 7.70933
R19568 vdd.n2906 vdd.n774 7.70933
R19569 vdd.n2976 vdd.n774 7.70933
R19570 vdd.n295 vdd.n292 7.3702
R19571 vdd.n240 vdd.n237 7.3702
R19572 vdd.n197 vdd.n194 7.3702
R19573 vdd.n142 vdd.n139 7.3702
R19574 vdd.n100 vdd.n97 7.3702
R19575 vdd.n45 vdd.n42 7.3702
R19576 vdd.n1664 vdd.n1661 7.3702
R19577 vdd.n1719 vdd.n1716 7.3702
R19578 vdd.n1566 vdd.n1563 7.3702
R19579 vdd.n1621 vdd.n1618 7.3702
R19580 vdd.n1469 vdd.n1466 7.3702
R19581 vdd.n1524 vdd.n1521 7.3702
R19582 vdd.n1307 vdd.n1306 6.98232
R19583 vdd.n1956 vdd.n1955 6.98232
R19584 vdd.n547 vdd.n546 6.98232
R19585 vdd.n3060 vdd.n3059 6.98232
R19586 vdd.n1794 vdd.t118 6.91577
R19587 vdd.n3169 vdd.t80 6.91577
R19588 vdd.t45 vdd.n1075 6.68904
R19589 vdd.n3185 vdd.t47 6.68904
R19590 vdd.n1752 vdd.t96 6.46231
R19591 vdd.n3213 vdd.t55 6.46231
R19592 vdd.n3292 vdd.n321 6.32949
R19593 vdd.n1746 vdd.n1745 6.32949
R19594 vdd.t59 vdd.n1103 6.23558
R19595 vdd.t50 vdd.n332 6.23558
R19596 vdd.n1416 vdd.t82 6.00885
R19597 vdd.n2329 vdd.t147 6.00885
R19598 vdd.n2829 vdd.t0 6.00885
R19599 vdd.n3271 vdd.t53 6.00885
R19600 vdd.n1004 vdd.t235 5.89549
R19601 vdd.t203 vdd.n822 5.89549
R19602 vdd.n296 vdd.n295 5.81868
R19603 vdd.n241 vdd.n240 5.81868
R19604 vdd.n198 vdd.n197 5.81868
R19605 vdd.n143 vdd.n142 5.81868
R19606 vdd.n101 vdd.n100 5.81868
R19607 vdd.n46 vdd.n45 5.81868
R19608 vdd.n1665 vdd.n1664 5.81868
R19609 vdd.n1720 vdd.n1719 5.81868
R19610 vdd.n1567 vdd.n1566 5.81868
R19611 vdd.n1622 vdd.n1621 5.81868
R19612 vdd.n1470 vdd.n1469 5.81868
R19613 vdd.n1525 vdd.n1524 5.81868
R19614 vdd.t231 vdd.n1008 5.78212
R19615 vdd.n2073 vdd.t216 5.78212
R19616 vdd.n2698 vdd.t224 5.78212
R19617 vdd.n817 vdd.t220 5.78212
R19618 vdd.n2457 vdd.n2456 5.77611
R19619 vdd.n2200 vdd.n2070 5.77611
R19620 vdd.n2711 vdd.n2710 5.77611
R19621 vdd.n2915 vdd.n806 5.77611
R19622 vdd.n2981 vdd.n770 5.77611
R19623 vdd.n2621 vdd.n2561 5.77611
R19624 vdd.n2382 vdd.n938 5.77611
R19625 vdd.n2130 vdd.n2129 5.77611
R19626 vdd.n1376 vdd.n1150 5.62474
R19627 vdd.n2252 vdd.n2249 5.62474
R19628 vdd.n3250 vdd.n407 5.62474
R19629 vdd.n3015 vdd.n3012 5.62474
R19630 vdd.t153 vdd.n960 5.44203
R19631 vdd.n864 vdd.t262 5.44203
R19632 vdd.n1126 vdd.t82 5.32866
R19633 vdd.t53 vdd.n3270 5.32866
R19634 vdd.n1432 vdd.t59 5.10193
R19635 vdd.t139 vdd.n983 5.10193
R19636 vdd.n973 vdd.t9 5.10193
R19637 vdd.t10 vdd.n851 5.10193
R19638 vdd.n841 vdd.t152 5.10193
R19639 vdd.n3279 vdd.t50 5.10193
R19640 vdd.n299 vdd.n290 5.04292
R19641 vdd.n244 vdd.n235 5.04292
R19642 vdd.n201 vdd.n192 5.04292
R19643 vdd.n146 vdd.n137 5.04292
R19644 vdd.n104 vdd.n95 5.04292
R19645 vdd.n49 vdd.n40 5.04292
R19646 vdd.n1668 vdd.n1659 5.04292
R19647 vdd.n1723 vdd.n1714 5.04292
R19648 vdd.n1570 vdd.n1561 5.04292
R19649 vdd.n1625 vdd.n1616 5.04292
R19650 vdd.n1473 vdd.n1464 5.04292
R19651 vdd.n1528 vdd.n1519 5.04292
R19652 vdd.n1448 vdd.t96 4.8752
R19653 vdd.t149 vdd.t150 4.8752
R19654 vdd.t148 vdd.t140 4.8752
R19655 vdd.t7 vdd.t6 4.8752
R19656 vdd.t155 vdd.t142 4.8752
R19657 vdd.t55 vdd.n328 4.8752
R19658 vdd.n2458 vdd.n2457 4.83952
R19659 vdd.n2070 vdd.n2066 4.83952
R19660 vdd.n2712 vdd.n2711 4.83952
R19661 vdd.n806 vdd.n801 4.83952
R19662 vdd.n770 vdd.n765 4.83952
R19663 vdd.n2618 vdd.n2561 4.83952
R19664 vdd.n2385 vdd.n938 4.83952
R19665 vdd.n2129 vdd.n2128 4.83952
R19666 vdd.n1924 vdd.n1036 4.74817
R19667 vdd.n1919 vdd.n1037 4.74817
R19668 vdd.n1821 vdd.n1818 4.74817
R19669 vdd.n2233 vdd.n1822 4.74817
R19670 vdd.n2235 vdd.n1821 4.74817
R19671 vdd.n2234 vdd.n2233 4.74817
R19672 vdd.n664 vdd.n662 4.74817
R19673 vdd.n3130 vdd.n665 4.74817
R19674 vdd.n3133 vdd.n665 4.74817
R19675 vdd.n3134 vdd.n664 4.74817
R19676 vdd.n3022 vdd.n749 4.74817
R19677 vdd.n3018 vdd.n751 4.74817
R19678 vdd.n3021 vdd.n751 4.74817
R19679 vdd.n3026 vdd.n749 4.74817
R19680 vdd.n1920 vdd.n1036 4.74817
R19681 vdd.n1039 vdd.n1037 4.74817
R19682 vdd.n321 vdd.n320 4.7074
R19683 vdd.n223 vdd.n222 4.7074
R19684 vdd.n1745 vdd.n1744 4.7074
R19685 vdd.n1647 vdd.n1646 4.7074
R19686 vdd.n1768 vdd.t45 4.64847
R19687 vdd.n3194 vdd.t47 4.64847
R19688 vdd.n2335 vdd.t162 4.53511
R19689 vdd.n2823 vdd.t145 4.53511
R19690 vdd.n1069 vdd.t118 4.42174
R19691 vdd.t80 vdd.n635 4.42174
R19692 vdd.n2367 vdd.t143 4.30838
R19693 vdd.n2793 vdd.t4 4.30838
R19694 vdd.n300 vdd.n288 4.26717
R19695 vdd.n245 vdd.n233 4.26717
R19696 vdd.n202 vdd.n190 4.26717
R19697 vdd.n147 vdd.n135 4.26717
R19698 vdd.n105 vdd.n93 4.26717
R19699 vdd.n50 vdd.n38 4.26717
R19700 vdd.n1669 vdd.n1657 4.26717
R19701 vdd.n1724 vdd.n1712 4.26717
R19702 vdd.n1571 vdd.n1559 4.26717
R19703 vdd.n1626 vdd.n1614 4.26717
R19704 vdd.n1474 vdd.n1462 4.26717
R19705 vdd.n1529 vdd.n1517 4.26717
R19706 vdd.n321 vdd.n223 4.10845
R19707 vdd.n1745 vdd.n1647 4.10845
R19708 vdd.n277 vdd.t133 4.06363
R19709 vdd.n277 vdd.t44 4.06363
R19710 vdd.n275 vdd.t65 4.06363
R19711 vdd.n275 vdd.t132 4.06363
R19712 vdd.n273 vdd.t134 4.06363
R19713 vdd.n273 vdd.t64 4.06363
R19714 vdd.n271 vdd.t69 4.06363
R19715 vdd.n271 vdd.t71 4.06363
R19716 vdd.n269 vdd.t110 4.06363
R19717 vdd.n269 vdd.t36 4.06363
R19718 vdd.n267 vdd.t39 4.06363
R19719 vdd.n267 vdd.t89 4.06363
R19720 vdd.n265 vdd.t91 4.06363
R19721 vdd.n265 vdd.t115 4.06363
R19722 vdd.n179 vdd.t122 4.06363
R19723 vdd.n179 vdd.t28 4.06363
R19724 vdd.n177 vdd.t52 4.06363
R19725 vdd.n177 vdd.t121 4.06363
R19726 vdd.n175 vdd.t125 4.06363
R19727 vdd.n175 vdd.t51 4.06363
R19728 vdd.n173 vdd.t56 4.06363
R19729 vdd.n173 vdd.t58 4.06363
R19730 vdd.n171 vdd.t101 4.06363
R19731 vdd.n171 vdd.t138 4.06363
R19732 vdd.n169 vdd.t18 4.06363
R19733 vdd.n169 vdd.t72 4.06363
R19734 vdd.n167 vdd.t81 4.06363
R19735 vdd.n167 vdd.t103 4.06363
R19736 vdd.n82 vdd.t54 4.06363
R19737 vdd.n82 vdd.t117 4.06363
R19738 vdd.n80 vdd.t30 4.06363
R19739 vdd.n80 vdd.t77 4.06363
R19740 vdd.n78 vdd.t22 4.06363
R19741 vdd.n78 vdd.t61 4.06363
R19742 vdd.n76 vdd.t131 4.06363
R19743 vdd.n76 vdd.t107 4.06363
R19744 vdd.n74 vdd.t111 4.06363
R19745 vdd.n74 vdd.t68 4.06363
R19746 vdd.n72 vdd.t136 4.06363
R19747 vdd.n72 vdd.t48 4.06363
R19748 vdd.n70 vdd.t123 4.06363
R19749 vdd.n70 vdd.t75 4.06363
R19750 vdd.n1689 vdd.t41 4.06363
R19751 vdd.n1689 vdd.t128 4.06363
R19752 vdd.n1691 vdd.t127 4.06363
R19753 vdd.n1691 vdd.t109 4.06363
R19754 vdd.n1693 vdd.t86 4.06363
R19755 vdd.n1693 vdd.t38 4.06363
R19756 vdd.n1695 vdd.t137 4.06363
R19757 vdd.n1695 vdd.t108 4.06363
R19758 vdd.n1697 vdd.t104 4.06363
R19759 vdd.n1697 vdd.t63 4.06363
R19760 vdd.n1699 vdd.t62 4.06363
R19761 vdd.n1699 vdd.t105 4.06363
R19762 vdd.n1701 vdd.t92 4.06363
R19763 vdd.n1701 vdd.t93 4.06363
R19764 vdd.n1591 vdd.t26 4.06363
R19765 vdd.n1591 vdd.t119 4.06363
R19766 vdd.n1593 vdd.t112 4.06363
R19767 vdd.n1593 vdd.t99 4.06363
R19768 vdd.n1595 vdd.t70 4.06363
R19769 vdd.n1595 vdd.t16 4.06363
R19770 vdd.n1597 vdd.t126 4.06363
R19771 vdd.n1597 vdd.t97 4.06363
R19772 vdd.n1599 vdd.t94 4.06363
R19773 vdd.n1599 vdd.t49 4.06363
R19774 vdd.n1601 vdd.t43 4.06363
R19775 vdd.n1601 vdd.t95 4.06363
R19776 vdd.n1603 vdd.t85 4.06363
R19777 vdd.n1603 vdd.t83 4.06363
R19778 vdd.n1494 vdd.t73 4.06363
R19779 vdd.n1494 vdd.t124 4.06363
R19780 vdd.n1496 vdd.t46 4.06363
R19781 vdd.n1496 vdd.t106 4.06363
R19782 vdd.n1498 vdd.t67 4.06363
R19783 vdd.n1498 vdd.t113 4.06363
R19784 vdd.n1500 vdd.t88 4.06363
R19785 vdd.n1500 vdd.t130 4.06363
R19786 vdd.n1502 vdd.t60 4.06363
R19787 vdd.n1502 vdd.t20 4.06363
R19788 vdd.n1504 vdd.t78 4.06363
R19789 vdd.n1504 vdd.t32 4.06363
R19790 vdd.n1506 vdd.t120 4.06363
R19791 vdd.n1506 vdd.t135 4.06363
R19792 vdd.n26 vdd.t171 3.9605
R19793 vdd.n26 vdd.t179 3.9605
R19794 vdd.n23 vdd.t172 3.9605
R19795 vdd.n23 vdd.t165 3.9605
R19796 vdd.n21 vdd.t168 3.9605
R19797 vdd.n21 vdd.t175 3.9605
R19798 vdd.n20 vdd.t174 3.9605
R19799 vdd.n20 vdd.t176 3.9605
R19800 vdd.n15 vdd.t167 3.9605
R19801 vdd.n15 vdd.t164 3.9605
R19802 vdd.n16 vdd.t169 3.9605
R19803 vdd.n16 vdd.t177 3.9605
R19804 vdd.n18 vdd.t166 3.9605
R19805 vdd.n18 vdd.t170 3.9605
R19806 vdd.n25 vdd.t173 3.9605
R19807 vdd.n25 vdd.t178 3.9605
R19808 vdd.n7 vdd.t156 3.61217
R19809 vdd.n7 vdd.t146 3.61217
R19810 vdd.n8 vdd.t8 3.61217
R19811 vdd.n8 vdd.t263 3.61217
R19812 vdd.n10 vdd.t257 3.61217
R19813 vdd.n10 vdd.t5 3.61217
R19814 vdd.n12 vdd.t161 3.61217
R19815 vdd.n12 vdd.t259 3.61217
R19816 vdd.n5 vdd.t261 3.61217
R19817 vdd.n5 vdd.t158 3.61217
R19818 vdd.n3 vdd.t144 3.61217
R19819 vdd.n3 vdd.t2 3.61217
R19820 vdd.n1 vdd.t154 3.61217
R19821 vdd.n1 vdd.t141 3.61217
R19822 vdd.n0 vdd.t163 3.61217
R19823 vdd.n0 vdd.t151 3.61217
R19824 vdd.n1382 vdd.t185 3.51482
R19825 vdd.n3255 vdd.t189 3.51482
R19826 vdd.n304 vdd.n303 3.49141
R19827 vdd.n249 vdd.n248 3.49141
R19828 vdd.n206 vdd.n205 3.49141
R19829 vdd.n151 vdd.n150 3.49141
R19830 vdd.n109 vdd.n108 3.49141
R19831 vdd.n54 vdd.n53 3.49141
R19832 vdd.n1673 vdd.n1672 3.49141
R19833 vdd.n1728 vdd.n1727 3.49141
R19834 vdd.n1575 vdd.n1574 3.49141
R19835 vdd.n1630 vdd.n1629 3.49141
R19836 vdd.n1478 vdd.n1477 3.49141
R19837 vdd.n1533 vdd.n1532 3.49141
R19838 vdd.n2073 vdd.t143 3.40145
R19839 vdd.n2521 vdd.t260 3.40145
R19840 vdd.n2774 vdd.t258 3.40145
R19841 vdd.n2698 vdd.t4 3.40145
R19842 vdd.n2174 vdd.t162 3.17472
R19843 vdd.n2677 vdd.t145 3.17472
R19844 vdd.n1785 vdd.t25 3.06136
R19845 vdd.n3177 vdd.t74 3.06136
R19846 vdd.t15 vdd.n1081 2.83463
R19847 vdd.n624 vdd.t100 2.83463
R19848 vdd.n307 vdd.n286 2.71565
R19849 vdd.n252 vdd.n231 2.71565
R19850 vdd.n209 vdd.n188 2.71565
R19851 vdd.n154 vdd.n133 2.71565
R19852 vdd.n112 vdd.n91 2.71565
R19853 vdd.n57 vdd.n36 2.71565
R19854 vdd.n1676 vdd.n1655 2.71565
R19855 vdd.n1731 vdd.n1710 2.71565
R19856 vdd.n1578 vdd.n1557 2.71565
R19857 vdd.n1633 vdd.n1612 2.71565
R19858 vdd.n1481 vdd.n1460 2.71565
R19859 vdd.n1536 vdd.n1515 2.71565
R19860 vdd.n1449 vdd.t87 2.6079
R19861 vdd.n2323 vdd.t139 2.6079
R19862 vdd.n2347 vdd.t9 2.6079
R19863 vdd.n2811 vdd.t10 2.6079
R19864 vdd.n2835 vdd.t152 2.6079
R19865 vdd.n3287 vdd.t57 2.6079
R19866 vdd.n2841 vdd.n2840 2.49806
R19867 vdd.n2315 vdd.n2314 2.49806
R19868 vdd.n294 vdd.n293 2.4129
R19869 vdd.n239 vdd.n238 2.4129
R19870 vdd.n196 vdd.n195 2.4129
R19871 vdd.n141 vdd.n140 2.4129
R19872 vdd.n99 vdd.n98 2.4129
R19873 vdd.n44 vdd.n43 2.4129
R19874 vdd.n1663 vdd.n1662 2.4129
R19875 vdd.n1718 vdd.n1717 2.4129
R19876 vdd.n1565 vdd.n1564 2.4129
R19877 vdd.n1620 vdd.n1619 2.4129
R19878 vdd.n1468 vdd.n1467 2.4129
R19879 vdd.n1523 vdd.n1522 2.4129
R19880 vdd.t31 vdd.n1110 2.38117
R19881 vdd.n3278 vdd.t29 2.38117
R19882 vdd.n2232 vdd.n1821 2.27742
R19883 vdd.n2233 vdd.n2232 2.27742
R19884 vdd.n2942 vdd.n665 2.27742
R19885 vdd.n2942 vdd.n664 2.27742
R19886 vdd.n3010 vdd.n751 2.27742
R19887 vdd.n3010 vdd.n749 2.27742
R19888 vdd.n2255 vdd.n1036 2.27742
R19889 vdd.n2255 vdd.n1037 2.27742
R19890 vdd.n2347 vdd.t153 2.2678
R19891 vdd.n2811 vdd.t262 2.2678
R19892 vdd.n1407 vdd.t84 2.15444
R19893 vdd.n3269 vdd.t27 2.15444
R19894 vdd.t140 vdd.n954 2.04107
R19895 vdd.n871 vdd.t7 2.04107
R19896 vdd.n308 vdd.n284 1.93989
R19897 vdd.n253 vdd.n229 1.93989
R19898 vdd.n210 vdd.n186 1.93989
R19899 vdd.n155 vdd.n131 1.93989
R19900 vdd.n113 vdd.n89 1.93989
R19901 vdd.n58 vdd.n34 1.93989
R19902 vdd.n1677 vdd.n1653 1.93989
R19903 vdd.n1732 vdd.n1708 1.93989
R19904 vdd.n1579 vdd.n1555 1.93989
R19905 vdd.n1634 vdd.n1610 1.93989
R19906 vdd.n1482 vdd.n1458 1.93989
R19907 vdd.n1537 vdd.n1513 1.93989
R19908 vdd.n2298 vdd.t231 1.92771
R19909 vdd.n2374 vdd.t216 1.92771
R19910 vdd.n2787 vdd.t224 1.92771
R19911 vdd.n2906 vdd.t220 1.92771
R19912 vdd.n1399 vdd.t23 1.70098
R19913 vdd.n2174 vdd.t147 1.70098
R19914 vdd.n979 vdd.t149 1.70098
R19915 vdd.t142 vdd.n845 1.70098
R19916 vdd.n2677 vdd.t0 1.70098
R19917 vdd.n3263 vdd.t33 1.70098
R19918 vdd.n1415 vdd.t42 1.47425
R19919 vdd.n349 vdd.t76 1.47425
R19920 vdd.n1440 vdd.t19 1.24752
R19921 vdd.t196 vdd.n1044 1.24752
R19922 vdd.n659 vdd.t181 1.24752
R19923 vdd.t21 vdd.n3285 1.24752
R19924 vdd.n319 vdd.n279 1.16414
R19925 vdd.n312 vdd.n311 1.16414
R19926 vdd.n264 vdd.n224 1.16414
R19927 vdd.n257 vdd.n256 1.16414
R19928 vdd.n221 vdd.n181 1.16414
R19929 vdd.n214 vdd.n213 1.16414
R19930 vdd.n166 vdd.n126 1.16414
R19931 vdd.n159 vdd.n158 1.16414
R19932 vdd.n124 vdd.n84 1.16414
R19933 vdd.n117 vdd.n116 1.16414
R19934 vdd.n69 vdd.n29 1.16414
R19935 vdd.n62 vdd.n61 1.16414
R19936 vdd.n1688 vdd.n1648 1.16414
R19937 vdd.n1681 vdd.n1680 1.16414
R19938 vdd.n1743 vdd.n1703 1.16414
R19939 vdd.n1736 vdd.n1735 1.16414
R19940 vdd.n1590 vdd.n1550 1.16414
R19941 vdd.n1583 vdd.n1582 1.16414
R19942 vdd.n1645 vdd.n1605 1.16414
R19943 vdd.n1638 vdd.n1637 1.16414
R19944 vdd.n1493 vdd.n1453 1.16414
R19945 vdd.n1486 vdd.n1485 1.16414
R19946 vdd.n1548 vdd.n1508 1.16414
R19947 vdd.n1541 vdd.n1540 1.16414
R19948 vdd.n2341 vdd.t150 1.13415
R19949 vdd.n2817 vdd.t155 1.13415
R19950 vdd.n1092 vdd.t66 1.02079
R19951 vdd.t235 vdd.t3 1.02079
R19952 vdd.t159 vdd.t203 1.02079
R19953 vdd.t35 vdd.n613 1.02079
R19954 vdd.n1271 vdd.n1150 0.970197
R19955 vdd.n2253 vdd.n2252 0.970197
R19956 vdd.n599 vdd.n407 0.970197
R19957 vdd.n3017 vdd.n3015 0.970197
R19958 vdd.n1746 vdd.n28 0.852297
R19959 vdd vdd.n3292 0.844463
R19960 vdd.n1777 vdd.t98 0.794056
R19961 vdd.n2317 vdd.t3 0.794056
R19962 vdd.n2353 vdd.t148 0.794056
R19963 vdd.n2805 vdd.t6 0.794056
R19964 vdd.n2843 vdd.t159 0.794056
R19965 vdd.n3186 vdd.t17 0.794056
R19966 vdd.n1793 vdd.t11 0.567326
R19967 vdd.t13 vdd.n642 0.567326
R19968 vdd.n2243 vdd.n2242 0.482207
R19969 vdd.n3142 vdd.n3141 0.482207
R19970 vdd.n444 vdd.n443 0.482207
R19971 vdd.n3249 vdd.n3248 0.482207
R19972 vdd.n3148 vdd.n656 0.482207
R19973 vdd.n1807 vdd.n1038 0.482207
R19974 vdd.n1378 vdd.n1377 0.482207
R19975 vdd.n1184 vdd.n1141 0.482207
R19976 vdd.n4 vdd.n2 0.459552
R19977 vdd.n11 vdd.n9 0.459552
R19978 vdd.n317 vdd.n316 0.388379
R19979 vdd.n283 vdd.n281 0.388379
R19980 vdd.n262 vdd.n261 0.388379
R19981 vdd.n228 vdd.n226 0.388379
R19982 vdd.n219 vdd.n218 0.388379
R19983 vdd.n185 vdd.n183 0.388379
R19984 vdd.n164 vdd.n163 0.388379
R19985 vdd.n130 vdd.n128 0.388379
R19986 vdd.n122 vdd.n121 0.388379
R19987 vdd.n88 vdd.n86 0.388379
R19988 vdd.n67 vdd.n66 0.388379
R19989 vdd.n33 vdd.n31 0.388379
R19990 vdd.n1686 vdd.n1685 0.388379
R19991 vdd.n1652 vdd.n1650 0.388379
R19992 vdd.n1741 vdd.n1740 0.388379
R19993 vdd.n1707 vdd.n1705 0.388379
R19994 vdd.n1588 vdd.n1587 0.388379
R19995 vdd.n1554 vdd.n1552 0.388379
R19996 vdd.n1643 vdd.n1642 0.388379
R19997 vdd.n1609 vdd.n1607 0.388379
R19998 vdd.n1491 vdd.n1490 0.388379
R19999 vdd.n1457 vdd.n1455 0.388379
R20000 vdd.n1546 vdd.n1545 0.388379
R20001 vdd.n1512 vdd.n1510 0.388379
R20002 vdd.n19 vdd.n17 0.387128
R20003 vdd.n24 vdd.n22 0.387128
R20004 vdd.n6 vdd.n4 0.358259
R20005 vdd.n13 vdd.n11 0.358259
R20006 vdd.n268 vdd.n266 0.358259
R20007 vdd.n270 vdd.n268 0.358259
R20008 vdd.n272 vdd.n270 0.358259
R20009 vdd.n274 vdd.n272 0.358259
R20010 vdd.n276 vdd.n274 0.358259
R20011 vdd.n278 vdd.n276 0.358259
R20012 vdd.n320 vdd.n278 0.358259
R20013 vdd.n170 vdd.n168 0.358259
R20014 vdd.n172 vdd.n170 0.358259
R20015 vdd.n174 vdd.n172 0.358259
R20016 vdd.n176 vdd.n174 0.358259
R20017 vdd.n178 vdd.n176 0.358259
R20018 vdd.n180 vdd.n178 0.358259
R20019 vdd.n222 vdd.n180 0.358259
R20020 vdd.n73 vdd.n71 0.358259
R20021 vdd.n75 vdd.n73 0.358259
R20022 vdd.n77 vdd.n75 0.358259
R20023 vdd.n79 vdd.n77 0.358259
R20024 vdd.n81 vdd.n79 0.358259
R20025 vdd.n83 vdd.n81 0.358259
R20026 vdd.n125 vdd.n83 0.358259
R20027 vdd.n1744 vdd.n1702 0.358259
R20028 vdd.n1702 vdd.n1700 0.358259
R20029 vdd.n1700 vdd.n1698 0.358259
R20030 vdd.n1698 vdd.n1696 0.358259
R20031 vdd.n1696 vdd.n1694 0.358259
R20032 vdd.n1694 vdd.n1692 0.358259
R20033 vdd.n1692 vdd.n1690 0.358259
R20034 vdd.n1646 vdd.n1604 0.358259
R20035 vdd.n1604 vdd.n1602 0.358259
R20036 vdd.n1602 vdd.n1600 0.358259
R20037 vdd.n1600 vdd.n1598 0.358259
R20038 vdd.n1598 vdd.n1596 0.358259
R20039 vdd.n1596 vdd.n1594 0.358259
R20040 vdd.n1594 vdd.n1592 0.358259
R20041 vdd.n1549 vdd.n1507 0.358259
R20042 vdd.n1507 vdd.n1505 0.358259
R20043 vdd.n1505 vdd.n1503 0.358259
R20044 vdd.n1503 vdd.n1501 0.358259
R20045 vdd.n1501 vdd.n1499 0.358259
R20046 vdd.n1499 vdd.n1497 0.358259
R20047 vdd.n1497 vdd.n1495 0.358259
R20048 vdd.n14 vdd.n6 0.334552
R20049 vdd.n14 vdd.n13 0.334552
R20050 vdd.n27 vdd.n19 0.21707
R20051 vdd.n27 vdd.n24 0.21707
R20052 vdd.n318 vdd.n280 0.155672
R20053 vdd.n310 vdd.n280 0.155672
R20054 vdd.n310 vdd.n309 0.155672
R20055 vdd.n309 vdd.n285 0.155672
R20056 vdd.n302 vdd.n285 0.155672
R20057 vdd.n302 vdd.n301 0.155672
R20058 vdd.n301 vdd.n289 0.155672
R20059 vdd.n294 vdd.n289 0.155672
R20060 vdd.n263 vdd.n225 0.155672
R20061 vdd.n255 vdd.n225 0.155672
R20062 vdd.n255 vdd.n254 0.155672
R20063 vdd.n254 vdd.n230 0.155672
R20064 vdd.n247 vdd.n230 0.155672
R20065 vdd.n247 vdd.n246 0.155672
R20066 vdd.n246 vdd.n234 0.155672
R20067 vdd.n239 vdd.n234 0.155672
R20068 vdd.n220 vdd.n182 0.155672
R20069 vdd.n212 vdd.n182 0.155672
R20070 vdd.n212 vdd.n211 0.155672
R20071 vdd.n211 vdd.n187 0.155672
R20072 vdd.n204 vdd.n187 0.155672
R20073 vdd.n204 vdd.n203 0.155672
R20074 vdd.n203 vdd.n191 0.155672
R20075 vdd.n196 vdd.n191 0.155672
R20076 vdd.n165 vdd.n127 0.155672
R20077 vdd.n157 vdd.n127 0.155672
R20078 vdd.n157 vdd.n156 0.155672
R20079 vdd.n156 vdd.n132 0.155672
R20080 vdd.n149 vdd.n132 0.155672
R20081 vdd.n149 vdd.n148 0.155672
R20082 vdd.n148 vdd.n136 0.155672
R20083 vdd.n141 vdd.n136 0.155672
R20084 vdd.n123 vdd.n85 0.155672
R20085 vdd.n115 vdd.n85 0.155672
R20086 vdd.n115 vdd.n114 0.155672
R20087 vdd.n114 vdd.n90 0.155672
R20088 vdd.n107 vdd.n90 0.155672
R20089 vdd.n107 vdd.n106 0.155672
R20090 vdd.n106 vdd.n94 0.155672
R20091 vdd.n99 vdd.n94 0.155672
R20092 vdd.n68 vdd.n30 0.155672
R20093 vdd.n60 vdd.n30 0.155672
R20094 vdd.n60 vdd.n59 0.155672
R20095 vdd.n59 vdd.n35 0.155672
R20096 vdd.n52 vdd.n35 0.155672
R20097 vdd.n52 vdd.n51 0.155672
R20098 vdd.n51 vdd.n39 0.155672
R20099 vdd.n44 vdd.n39 0.155672
R20100 vdd.n1687 vdd.n1649 0.155672
R20101 vdd.n1679 vdd.n1649 0.155672
R20102 vdd.n1679 vdd.n1678 0.155672
R20103 vdd.n1678 vdd.n1654 0.155672
R20104 vdd.n1671 vdd.n1654 0.155672
R20105 vdd.n1671 vdd.n1670 0.155672
R20106 vdd.n1670 vdd.n1658 0.155672
R20107 vdd.n1663 vdd.n1658 0.155672
R20108 vdd.n1742 vdd.n1704 0.155672
R20109 vdd.n1734 vdd.n1704 0.155672
R20110 vdd.n1734 vdd.n1733 0.155672
R20111 vdd.n1733 vdd.n1709 0.155672
R20112 vdd.n1726 vdd.n1709 0.155672
R20113 vdd.n1726 vdd.n1725 0.155672
R20114 vdd.n1725 vdd.n1713 0.155672
R20115 vdd.n1718 vdd.n1713 0.155672
R20116 vdd.n1589 vdd.n1551 0.155672
R20117 vdd.n1581 vdd.n1551 0.155672
R20118 vdd.n1581 vdd.n1580 0.155672
R20119 vdd.n1580 vdd.n1556 0.155672
R20120 vdd.n1573 vdd.n1556 0.155672
R20121 vdd.n1573 vdd.n1572 0.155672
R20122 vdd.n1572 vdd.n1560 0.155672
R20123 vdd.n1565 vdd.n1560 0.155672
R20124 vdd.n1644 vdd.n1606 0.155672
R20125 vdd.n1636 vdd.n1606 0.155672
R20126 vdd.n1636 vdd.n1635 0.155672
R20127 vdd.n1635 vdd.n1611 0.155672
R20128 vdd.n1628 vdd.n1611 0.155672
R20129 vdd.n1628 vdd.n1627 0.155672
R20130 vdd.n1627 vdd.n1615 0.155672
R20131 vdd.n1620 vdd.n1615 0.155672
R20132 vdd.n1492 vdd.n1454 0.155672
R20133 vdd.n1484 vdd.n1454 0.155672
R20134 vdd.n1484 vdd.n1483 0.155672
R20135 vdd.n1483 vdd.n1459 0.155672
R20136 vdd.n1476 vdd.n1459 0.155672
R20137 vdd.n1476 vdd.n1475 0.155672
R20138 vdd.n1475 vdd.n1463 0.155672
R20139 vdd.n1468 vdd.n1463 0.155672
R20140 vdd.n1547 vdd.n1509 0.155672
R20141 vdd.n1539 vdd.n1509 0.155672
R20142 vdd.n1539 vdd.n1538 0.155672
R20143 vdd.n1538 vdd.n1514 0.155672
R20144 vdd.n1531 vdd.n1514 0.155672
R20145 vdd.n1531 vdd.n1530 0.155672
R20146 vdd.n1530 vdd.n1518 0.155672
R20147 vdd.n1523 vdd.n1518 0.155672
R20148 vdd.n2018 vdd.n1823 0.152939
R20149 vdd.n1829 vdd.n1823 0.152939
R20150 vdd.n1830 vdd.n1829 0.152939
R20151 vdd.n1831 vdd.n1830 0.152939
R20152 vdd.n1832 vdd.n1831 0.152939
R20153 vdd.n1836 vdd.n1832 0.152939
R20154 vdd.n1837 vdd.n1836 0.152939
R20155 vdd.n1838 vdd.n1837 0.152939
R20156 vdd.n1839 vdd.n1838 0.152939
R20157 vdd.n1843 vdd.n1839 0.152939
R20158 vdd.n1844 vdd.n1843 0.152939
R20159 vdd.n1845 vdd.n1844 0.152939
R20160 vdd.n1993 vdd.n1845 0.152939
R20161 vdd.n1993 vdd.n1992 0.152939
R20162 vdd.n1992 vdd.n1991 0.152939
R20163 vdd.n1991 vdd.n1851 0.152939
R20164 vdd.n1856 vdd.n1851 0.152939
R20165 vdd.n1857 vdd.n1856 0.152939
R20166 vdd.n1858 vdd.n1857 0.152939
R20167 vdd.n1862 vdd.n1858 0.152939
R20168 vdd.n1863 vdd.n1862 0.152939
R20169 vdd.n1864 vdd.n1863 0.152939
R20170 vdd.n1865 vdd.n1864 0.152939
R20171 vdd.n1869 vdd.n1865 0.152939
R20172 vdd.n1870 vdd.n1869 0.152939
R20173 vdd.n1871 vdd.n1870 0.152939
R20174 vdd.n1872 vdd.n1871 0.152939
R20175 vdd.n1876 vdd.n1872 0.152939
R20176 vdd.n1877 vdd.n1876 0.152939
R20177 vdd.n1878 vdd.n1877 0.152939
R20178 vdd.n1879 vdd.n1878 0.152939
R20179 vdd.n1883 vdd.n1879 0.152939
R20180 vdd.n1884 vdd.n1883 0.152939
R20181 vdd.n1885 vdd.n1884 0.152939
R20182 vdd.n1954 vdd.n1885 0.152939
R20183 vdd.n1954 vdd.n1953 0.152939
R20184 vdd.n1953 vdd.n1952 0.152939
R20185 vdd.n1952 vdd.n1891 0.152939
R20186 vdd.n1896 vdd.n1891 0.152939
R20187 vdd.n1897 vdd.n1896 0.152939
R20188 vdd.n1898 vdd.n1897 0.152939
R20189 vdd.n1902 vdd.n1898 0.152939
R20190 vdd.n1903 vdd.n1902 0.152939
R20191 vdd.n1904 vdd.n1903 0.152939
R20192 vdd.n1905 vdd.n1904 0.152939
R20193 vdd.n1909 vdd.n1905 0.152939
R20194 vdd.n1910 vdd.n1909 0.152939
R20195 vdd.n1911 vdd.n1910 0.152939
R20196 vdd.n1912 vdd.n1911 0.152939
R20197 vdd.n1913 vdd.n1912 0.152939
R20198 vdd.n1913 vdd.n1035 0.152939
R20199 vdd.n2242 vdd.n1817 0.152939
R20200 vdd.n1749 vdd.n1748 0.152939
R20201 vdd.n1749 vdd.n1084 0.152939
R20202 vdd.n1763 vdd.n1084 0.152939
R20203 vdd.n1764 vdd.n1763 0.152939
R20204 vdd.n1765 vdd.n1764 0.152939
R20205 vdd.n1765 vdd.n1072 0.152939
R20206 vdd.n1780 vdd.n1072 0.152939
R20207 vdd.n1781 vdd.n1780 0.152939
R20208 vdd.n1782 vdd.n1781 0.152939
R20209 vdd.n1782 vdd.n1061 0.152939
R20210 vdd.n1797 vdd.n1061 0.152939
R20211 vdd.n1798 vdd.n1797 0.152939
R20212 vdd.n1799 vdd.n1798 0.152939
R20213 vdd.n1799 vdd.n1049 0.152939
R20214 vdd.n1815 vdd.n1049 0.152939
R20215 vdd.n1816 vdd.n1815 0.152939
R20216 vdd.n2243 vdd.n1816 0.152939
R20217 vdd.n670 vdd.n667 0.152939
R20218 vdd.n671 vdd.n670 0.152939
R20219 vdd.n672 vdd.n671 0.152939
R20220 vdd.n673 vdd.n672 0.152939
R20221 vdd.n676 vdd.n673 0.152939
R20222 vdd.n677 vdd.n676 0.152939
R20223 vdd.n678 vdd.n677 0.152939
R20224 vdd.n679 vdd.n678 0.152939
R20225 vdd.n682 vdd.n679 0.152939
R20226 vdd.n683 vdd.n682 0.152939
R20227 vdd.n684 vdd.n683 0.152939
R20228 vdd.n685 vdd.n684 0.152939
R20229 vdd.n690 vdd.n685 0.152939
R20230 vdd.n691 vdd.n690 0.152939
R20231 vdd.n692 vdd.n691 0.152939
R20232 vdd.n693 vdd.n692 0.152939
R20233 vdd.n696 vdd.n693 0.152939
R20234 vdd.n697 vdd.n696 0.152939
R20235 vdd.n698 vdd.n697 0.152939
R20236 vdd.n699 vdd.n698 0.152939
R20237 vdd.n702 vdd.n699 0.152939
R20238 vdd.n703 vdd.n702 0.152939
R20239 vdd.n704 vdd.n703 0.152939
R20240 vdd.n705 vdd.n704 0.152939
R20241 vdd.n708 vdd.n705 0.152939
R20242 vdd.n709 vdd.n708 0.152939
R20243 vdd.n710 vdd.n709 0.152939
R20244 vdd.n711 vdd.n710 0.152939
R20245 vdd.n714 vdd.n711 0.152939
R20246 vdd.n715 vdd.n714 0.152939
R20247 vdd.n716 vdd.n715 0.152939
R20248 vdd.n717 vdd.n716 0.152939
R20249 vdd.n720 vdd.n717 0.152939
R20250 vdd.n721 vdd.n720 0.152939
R20251 vdd.n3058 vdd.n721 0.152939
R20252 vdd.n3058 vdd.n3057 0.152939
R20253 vdd.n3057 vdd.n3056 0.152939
R20254 vdd.n3056 vdd.n725 0.152939
R20255 vdd.n730 vdd.n725 0.152939
R20256 vdd.n731 vdd.n730 0.152939
R20257 vdd.n734 vdd.n731 0.152939
R20258 vdd.n735 vdd.n734 0.152939
R20259 vdd.n736 vdd.n735 0.152939
R20260 vdd.n737 vdd.n736 0.152939
R20261 vdd.n740 vdd.n737 0.152939
R20262 vdd.n741 vdd.n740 0.152939
R20263 vdd.n742 vdd.n741 0.152939
R20264 vdd.n743 vdd.n742 0.152939
R20265 vdd.n746 vdd.n743 0.152939
R20266 vdd.n747 vdd.n746 0.152939
R20267 vdd.n748 vdd.n747 0.152939
R20268 vdd.n3141 vdd.n661 0.152939
R20269 vdd.n3142 vdd.n651 0.152939
R20270 vdd.n3156 vdd.n651 0.152939
R20271 vdd.n3157 vdd.n3156 0.152939
R20272 vdd.n3158 vdd.n3157 0.152939
R20273 vdd.n3158 vdd.n639 0.152939
R20274 vdd.n3172 vdd.n639 0.152939
R20275 vdd.n3173 vdd.n3172 0.152939
R20276 vdd.n3174 vdd.n3173 0.152939
R20277 vdd.n3174 vdd.n627 0.152939
R20278 vdd.n3189 vdd.n627 0.152939
R20279 vdd.n3190 vdd.n3189 0.152939
R20280 vdd.n3191 vdd.n3190 0.152939
R20281 vdd.n3191 vdd.n616 0.152939
R20282 vdd.n3208 vdd.n616 0.152939
R20283 vdd.n3209 vdd.n3208 0.152939
R20284 vdd.n3210 vdd.n3209 0.152939
R20285 vdd.n3210 vdd.n322 0.152939
R20286 vdd.n3290 vdd.n323 0.152939
R20287 vdd.n334 vdd.n323 0.152939
R20288 vdd.n335 vdd.n334 0.152939
R20289 vdd.n336 vdd.n335 0.152939
R20290 vdd.n343 vdd.n336 0.152939
R20291 vdd.n344 vdd.n343 0.152939
R20292 vdd.n345 vdd.n344 0.152939
R20293 vdd.n346 vdd.n345 0.152939
R20294 vdd.n354 vdd.n346 0.152939
R20295 vdd.n355 vdd.n354 0.152939
R20296 vdd.n356 vdd.n355 0.152939
R20297 vdd.n357 vdd.n356 0.152939
R20298 vdd.n365 vdd.n357 0.152939
R20299 vdd.n366 vdd.n365 0.152939
R20300 vdd.n367 vdd.n366 0.152939
R20301 vdd.n368 vdd.n367 0.152939
R20302 vdd.n443 vdd.n368 0.152939
R20303 vdd.n444 vdd.n442 0.152939
R20304 vdd.n451 vdd.n442 0.152939
R20305 vdd.n452 vdd.n451 0.152939
R20306 vdd.n453 vdd.n452 0.152939
R20307 vdd.n453 vdd.n440 0.152939
R20308 vdd.n461 vdd.n440 0.152939
R20309 vdd.n462 vdd.n461 0.152939
R20310 vdd.n463 vdd.n462 0.152939
R20311 vdd.n463 vdd.n438 0.152939
R20312 vdd.n471 vdd.n438 0.152939
R20313 vdd.n472 vdd.n471 0.152939
R20314 vdd.n473 vdd.n472 0.152939
R20315 vdd.n473 vdd.n436 0.152939
R20316 vdd.n481 vdd.n436 0.152939
R20317 vdd.n482 vdd.n481 0.152939
R20318 vdd.n483 vdd.n482 0.152939
R20319 vdd.n483 vdd.n434 0.152939
R20320 vdd.n491 vdd.n434 0.152939
R20321 vdd.n492 vdd.n491 0.152939
R20322 vdd.n493 vdd.n492 0.152939
R20323 vdd.n493 vdd.n430 0.152939
R20324 vdd.n501 vdd.n430 0.152939
R20325 vdd.n502 vdd.n501 0.152939
R20326 vdd.n503 vdd.n502 0.152939
R20327 vdd.n503 vdd.n428 0.152939
R20328 vdd.n511 vdd.n428 0.152939
R20329 vdd.n512 vdd.n511 0.152939
R20330 vdd.n513 vdd.n512 0.152939
R20331 vdd.n513 vdd.n426 0.152939
R20332 vdd.n521 vdd.n426 0.152939
R20333 vdd.n522 vdd.n521 0.152939
R20334 vdd.n523 vdd.n522 0.152939
R20335 vdd.n523 vdd.n424 0.152939
R20336 vdd.n531 vdd.n424 0.152939
R20337 vdd.n532 vdd.n531 0.152939
R20338 vdd.n533 vdd.n532 0.152939
R20339 vdd.n533 vdd.n422 0.152939
R20340 vdd.n541 vdd.n422 0.152939
R20341 vdd.n542 vdd.n541 0.152939
R20342 vdd.n543 vdd.n542 0.152939
R20343 vdd.n543 vdd.n418 0.152939
R20344 vdd.n551 vdd.n418 0.152939
R20345 vdd.n552 vdd.n551 0.152939
R20346 vdd.n553 vdd.n552 0.152939
R20347 vdd.n553 vdd.n416 0.152939
R20348 vdd.n561 vdd.n416 0.152939
R20349 vdd.n562 vdd.n561 0.152939
R20350 vdd.n563 vdd.n562 0.152939
R20351 vdd.n563 vdd.n414 0.152939
R20352 vdd.n571 vdd.n414 0.152939
R20353 vdd.n572 vdd.n571 0.152939
R20354 vdd.n573 vdd.n572 0.152939
R20355 vdd.n573 vdd.n412 0.152939
R20356 vdd.n581 vdd.n412 0.152939
R20357 vdd.n582 vdd.n581 0.152939
R20358 vdd.n583 vdd.n582 0.152939
R20359 vdd.n583 vdd.n410 0.152939
R20360 vdd.n591 vdd.n410 0.152939
R20361 vdd.n592 vdd.n591 0.152939
R20362 vdd.n593 vdd.n592 0.152939
R20363 vdd.n593 vdd.n408 0.152939
R20364 vdd.n600 vdd.n408 0.152939
R20365 vdd.n3249 vdd.n600 0.152939
R20366 vdd.n3149 vdd.n3148 0.152939
R20367 vdd.n3150 vdd.n3149 0.152939
R20368 vdd.n3150 vdd.n645 0.152939
R20369 vdd.n3164 vdd.n645 0.152939
R20370 vdd.n3165 vdd.n3164 0.152939
R20371 vdd.n3166 vdd.n3165 0.152939
R20372 vdd.n3166 vdd.n632 0.152939
R20373 vdd.n3180 vdd.n632 0.152939
R20374 vdd.n3181 vdd.n3180 0.152939
R20375 vdd.n3182 vdd.n3181 0.152939
R20376 vdd.n3182 vdd.n621 0.152939
R20377 vdd.n3197 vdd.n621 0.152939
R20378 vdd.n3198 vdd.n3197 0.152939
R20379 vdd.n3199 vdd.n3198 0.152939
R20380 vdd.n3201 vdd.n3199 0.152939
R20381 vdd.n3201 vdd.n3200 0.152939
R20382 vdd.n3200 vdd.n611 0.152939
R20383 vdd.n611 vdd.n609 0.152939
R20384 vdd.n3219 vdd.n609 0.152939
R20385 vdd.n3220 vdd.n3219 0.152939
R20386 vdd.n3221 vdd.n3220 0.152939
R20387 vdd.n3221 vdd.n607 0.152939
R20388 vdd.n3226 vdd.n607 0.152939
R20389 vdd.n3227 vdd.n3226 0.152939
R20390 vdd.n3228 vdd.n3227 0.152939
R20391 vdd.n3228 vdd.n605 0.152939
R20392 vdd.n3233 vdd.n605 0.152939
R20393 vdd.n3234 vdd.n3233 0.152939
R20394 vdd.n3235 vdd.n3234 0.152939
R20395 vdd.n3235 vdd.n603 0.152939
R20396 vdd.n3241 vdd.n603 0.152939
R20397 vdd.n3242 vdd.n3241 0.152939
R20398 vdd.n3243 vdd.n3242 0.152939
R20399 vdd.n3243 vdd.n601 0.152939
R20400 vdd.n3248 vdd.n601 0.152939
R20401 vdd.n3011 vdd.n656 0.152939
R20402 vdd.n2254 vdd.n1038 0.152939
R20403 vdd.n1379 vdd.n1378 0.152939
R20404 vdd.n1379 vdd.n1135 0.152939
R20405 vdd.n1393 vdd.n1135 0.152939
R20406 vdd.n1394 vdd.n1393 0.152939
R20407 vdd.n1395 vdd.n1394 0.152939
R20408 vdd.n1395 vdd.n1123 0.152939
R20409 vdd.n1410 vdd.n1123 0.152939
R20410 vdd.n1411 vdd.n1410 0.152939
R20411 vdd.n1412 vdd.n1411 0.152939
R20412 vdd.n1412 vdd.n1113 0.152939
R20413 vdd.n1427 vdd.n1113 0.152939
R20414 vdd.n1428 vdd.n1427 0.152939
R20415 vdd.n1429 vdd.n1428 0.152939
R20416 vdd.n1429 vdd.n1100 0.152939
R20417 vdd.n1443 vdd.n1100 0.152939
R20418 vdd.n1444 vdd.n1443 0.152939
R20419 vdd.n1445 vdd.n1444 0.152939
R20420 vdd.n1445 vdd.n1089 0.152939
R20421 vdd.n1755 vdd.n1089 0.152939
R20422 vdd.n1756 vdd.n1755 0.152939
R20423 vdd.n1757 vdd.n1756 0.152939
R20424 vdd.n1757 vdd.n1078 0.152939
R20425 vdd.n1771 vdd.n1078 0.152939
R20426 vdd.n1772 vdd.n1771 0.152939
R20427 vdd.n1773 vdd.n1772 0.152939
R20428 vdd.n1773 vdd.n1066 0.152939
R20429 vdd.n1788 vdd.n1066 0.152939
R20430 vdd.n1789 vdd.n1788 0.152939
R20431 vdd.n1790 vdd.n1789 0.152939
R20432 vdd.n1790 vdd.n1056 0.152939
R20433 vdd.n1805 vdd.n1056 0.152939
R20434 vdd.n1806 vdd.n1805 0.152939
R20435 vdd.n1809 vdd.n1806 0.152939
R20436 vdd.n1809 vdd.n1808 0.152939
R20437 vdd.n1808 vdd.n1807 0.152939
R20438 vdd.n1369 vdd.n1184 0.152939
R20439 vdd.n1369 vdd.n1368 0.152939
R20440 vdd.n1368 vdd.n1367 0.152939
R20441 vdd.n1367 vdd.n1186 0.152939
R20442 vdd.n1363 vdd.n1186 0.152939
R20443 vdd.n1363 vdd.n1362 0.152939
R20444 vdd.n1362 vdd.n1361 0.152939
R20445 vdd.n1361 vdd.n1191 0.152939
R20446 vdd.n1357 vdd.n1191 0.152939
R20447 vdd.n1357 vdd.n1356 0.152939
R20448 vdd.n1356 vdd.n1355 0.152939
R20449 vdd.n1355 vdd.n1197 0.152939
R20450 vdd.n1351 vdd.n1197 0.152939
R20451 vdd.n1351 vdd.n1350 0.152939
R20452 vdd.n1350 vdd.n1349 0.152939
R20453 vdd.n1349 vdd.n1203 0.152939
R20454 vdd.n1345 vdd.n1203 0.152939
R20455 vdd.n1345 vdd.n1344 0.152939
R20456 vdd.n1344 vdd.n1343 0.152939
R20457 vdd.n1343 vdd.n1209 0.152939
R20458 vdd.n1335 vdd.n1209 0.152939
R20459 vdd.n1335 vdd.n1334 0.152939
R20460 vdd.n1334 vdd.n1333 0.152939
R20461 vdd.n1333 vdd.n1213 0.152939
R20462 vdd.n1329 vdd.n1213 0.152939
R20463 vdd.n1329 vdd.n1328 0.152939
R20464 vdd.n1328 vdd.n1327 0.152939
R20465 vdd.n1327 vdd.n1219 0.152939
R20466 vdd.n1323 vdd.n1219 0.152939
R20467 vdd.n1323 vdd.n1322 0.152939
R20468 vdd.n1322 vdd.n1321 0.152939
R20469 vdd.n1321 vdd.n1225 0.152939
R20470 vdd.n1317 vdd.n1225 0.152939
R20471 vdd.n1317 vdd.n1316 0.152939
R20472 vdd.n1316 vdd.n1315 0.152939
R20473 vdd.n1315 vdd.n1231 0.152939
R20474 vdd.n1311 vdd.n1231 0.152939
R20475 vdd.n1311 vdd.n1310 0.152939
R20476 vdd.n1310 vdd.n1309 0.152939
R20477 vdd.n1309 vdd.n1237 0.152939
R20478 vdd.n1302 vdd.n1237 0.152939
R20479 vdd.n1302 vdd.n1301 0.152939
R20480 vdd.n1301 vdd.n1300 0.152939
R20481 vdd.n1300 vdd.n1242 0.152939
R20482 vdd.n1296 vdd.n1242 0.152939
R20483 vdd.n1296 vdd.n1295 0.152939
R20484 vdd.n1295 vdd.n1294 0.152939
R20485 vdd.n1294 vdd.n1248 0.152939
R20486 vdd.n1290 vdd.n1248 0.152939
R20487 vdd.n1290 vdd.n1289 0.152939
R20488 vdd.n1289 vdd.n1288 0.152939
R20489 vdd.n1288 vdd.n1254 0.152939
R20490 vdd.n1284 vdd.n1254 0.152939
R20491 vdd.n1284 vdd.n1283 0.152939
R20492 vdd.n1283 vdd.n1282 0.152939
R20493 vdd.n1282 vdd.n1260 0.152939
R20494 vdd.n1278 vdd.n1260 0.152939
R20495 vdd.n1278 vdd.n1277 0.152939
R20496 vdd.n1277 vdd.n1276 0.152939
R20497 vdd.n1276 vdd.n1266 0.152939
R20498 vdd.n1272 vdd.n1266 0.152939
R20499 vdd.n1272 vdd.n1147 0.152939
R20500 vdd.n1377 vdd.n1147 0.152939
R20501 vdd.n1385 vdd.n1141 0.152939
R20502 vdd.n1386 vdd.n1385 0.152939
R20503 vdd.n1387 vdd.n1386 0.152939
R20504 vdd.n1387 vdd.n1129 0.152939
R20505 vdd.n1402 vdd.n1129 0.152939
R20506 vdd.n1403 vdd.n1402 0.152939
R20507 vdd.n1404 vdd.n1403 0.152939
R20508 vdd.n1404 vdd.n1118 0.152939
R20509 vdd.n1419 vdd.n1118 0.152939
R20510 vdd.n1420 vdd.n1419 0.152939
R20511 vdd.n1421 vdd.n1420 0.152939
R20512 vdd.n1421 vdd.n1107 0.152939
R20513 vdd.n1435 vdd.n1107 0.152939
R20514 vdd.n1436 vdd.n1435 0.152939
R20515 vdd.n1437 vdd.n1436 0.152939
R20516 vdd.n1437 vdd.n1095 0.152939
R20517 vdd.n1452 vdd.n1095 0.152939
R20518 vdd.n2232 vdd.n1817 0.110256
R20519 vdd.n2942 vdd.n661 0.110256
R20520 vdd.n3011 vdd.n3010 0.110256
R20521 vdd.n2255 vdd.n2254 0.110256
R20522 vdd.n1748 vdd.n1747 0.0695946
R20523 vdd.n3291 vdd.n322 0.0695946
R20524 vdd.n3291 vdd.n3290 0.0695946
R20525 vdd.n1747 vdd.n1452 0.0695946
R20526 vdd.n2232 vdd.n2018 0.0431829
R20527 vdd.n2255 vdd.n1035 0.0431829
R20528 vdd.n2942 vdd.n667 0.0431829
R20529 vdd.n3010 vdd.n748 0.0431829
R20530 vdd vdd.n28 0.00833333
R20531 a_n2848_n452.n5 a_n2848_n452.t75 539.01
R20532 a_n2848_n452.n97 a_n2848_n452.t58 512.366
R20533 a_n2848_n452.n96 a_n2848_n452.t62 512.366
R20534 a_n2848_n452.n70 a_n2848_n452.t52 512.366
R20535 a_n2848_n452.n95 a_n2848_n452.t67 512.366
R20536 a_n2848_n452.n1 a_n2848_n452.t29 533.058
R20537 a_n2848_n452.n101 a_n2848_n452.t37 512.366
R20538 a_n2848_n452.n100 a_n2848_n452.t23 512.366
R20539 a_n2848_n452.n69 a_n2848_n452.t31 512.366
R20540 a_n2848_n452.n98 a_n2848_n452.t41 512.366
R20541 a_n2848_n452.n19 a_n2848_n452.t25 539.01
R20542 a_n2848_n452.n78 a_n2848_n452.t43 512.366
R20543 a_n2848_n452.n79 a_n2848_n452.t39 512.366
R20544 a_n2848_n452.n73 a_n2848_n452.t27 512.366
R20545 a_n2848_n452.n80 a_n2848_n452.t35 512.366
R20546 a_n2848_n452.n23 a_n2848_n452.t70 539.01
R20547 a_n2848_n452.n75 a_n2848_n452.t71 512.366
R20548 a_n2848_n452.n76 a_n2848_n452.t50 512.366
R20549 a_n2848_n452.n74 a_n2848_n452.t56 512.366
R20550 a_n2848_n452.n77 a_n2848_n452.t65 512.366
R20551 a_n2848_n452.n92 a_n2848_n452.t64 512.366
R20552 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R20553 a_n2848_n452.n93 a_n2848_n452.t49 512.366
R20554 a_n2848_n452.n90 a_n2848_n452.t72 512.366
R20555 a_n2848_n452.n83 a_n2848_n452.t61 512.366
R20556 a_n2848_n452.n91 a_n2848_n452.t60 512.366
R20557 a_n2848_n452.n88 a_n2848_n452.t68 512.366
R20558 a_n2848_n452.n84 a_n2848_n452.t53 512.366
R20559 a_n2848_n452.n89 a_n2848_n452.t54 512.366
R20560 a_n2848_n452.n86 a_n2848_n452.t57 512.366
R20561 a_n2848_n452.n85 a_n2848_n452.t66 512.366
R20562 a_n2848_n452.n87 a_n2848_n452.t48 512.366
R20563 a_n2848_n452.n50 a_n2848_n452.n3 70.3058
R20564 a_n2848_n452.n47 a_n2848_n452.n6 70.3058
R20565 a_n2848_n452.n16 a_n2848_n452.n37 70.3058
R20566 a_n2848_n452.n20 a_n2848_n452.n34 70.3058
R20567 a_n2848_n452.n33 a_n2848_n452.n21 70.1674
R20568 a_n2848_n452.n33 a_n2848_n452.n74 20.9683
R20569 a_n2848_n452.n21 a_n2848_n452.n32 75.0448
R20570 a_n2848_n452.n76 a_n2848_n452.n32 11.2134
R20571 a_n2848_n452.n22 a_n2848_n452.n23 44.8194
R20572 a_n2848_n452.n36 a_n2848_n452.n17 70.1674
R20573 a_n2848_n452.n36 a_n2848_n452.n73 20.9683
R20574 a_n2848_n452.n17 a_n2848_n452.n35 75.0448
R20575 a_n2848_n452.n79 a_n2848_n452.n35 11.2134
R20576 a_n2848_n452.n18 a_n2848_n452.n19 44.8194
R20577 a_n2848_n452.n7 a_n2848_n452.n45 70.1674
R20578 a_n2848_n452.n9 a_n2848_n452.n43 70.1674
R20579 a_n2848_n452.n11 a_n2848_n452.n41 70.1674
R20580 a_n2848_n452.n14 a_n2848_n452.n39 70.1674
R20581 a_n2848_n452.n87 a_n2848_n452.n39 20.9683
R20582 a_n2848_n452.n38 a_n2848_n452.n15 75.0448
R20583 a_n2848_n452.n38 a_n2848_n452.n85 11.2134
R20584 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R20585 a_n2848_n452.n89 a_n2848_n452.n41 20.9683
R20586 a_n2848_n452.n40 a_n2848_n452.n12 75.0448
R20587 a_n2848_n452.n40 a_n2848_n452.n84 11.2134
R20588 a_n2848_n452.n12 a_n2848_n452.n88 161.3
R20589 a_n2848_n452.n91 a_n2848_n452.n43 20.9683
R20590 a_n2848_n452.n42 a_n2848_n452.n10 75.0448
R20591 a_n2848_n452.n42 a_n2848_n452.n83 11.2134
R20592 a_n2848_n452.n10 a_n2848_n452.n90 161.3
R20593 a_n2848_n452.n93 a_n2848_n452.n45 20.9683
R20594 a_n2848_n452.n44 a_n2848_n452.n8 75.0448
R20595 a_n2848_n452.n44 a_n2848_n452.n82 11.2134
R20596 a_n2848_n452.n8 a_n2848_n452.n92 161.3
R20597 a_n2848_n452.n6 a_n2848_n452.n46 70.1674
R20598 a_n2848_n452.n46 a_n2848_n452.n69 20.9683
R20599 a_n2848_n452.n99 a_n2848_n452.n0 161.3
R20600 a_n2848_n452.n4 a_n2848_n452.n49 70.1674
R20601 a_n2848_n452.n49 a_n2848_n452.n70 20.9683
R20602 a_n2848_n452.n48 a_n2848_n452.n4 75.0448
R20603 a_n2848_n452.n96 a_n2848_n452.n48 11.2134
R20604 a_n2848_n452.n2 a_n2848_n452.n5 44.8194
R20605 a_n2848_n452.n100 a_n2848_n452.n51 20.9683
R20606 a_n2848_n452.n51 a_n2848_n452.n0 70.1674
R20607 a_n2848_n452.n0 a_n2848_n452.n1 70.3058
R20608 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R20609 a_n2848_n452.n58 a_n2848_n452.n56 81.4626
R20610 a_n2848_n452.n54 a_n2848_n452.n52 81.4626
R20611 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R20612 a_n2848_n452.n31 a_n2848_n452.n68 80.9324
R20613 a_n2848_n452.n30 a_n2848_n452.n64 80.9324
R20614 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R20615 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R20616 a_n2848_n452.n58 a_n2848_n452.n57 80.9324
R20617 a_n2848_n452.n29 a_n2848_n452.n59 80.9324
R20618 a_n2848_n452.n28 a_n2848_n452.n55 80.9324
R20619 a_n2848_n452.n54 a_n2848_n452.n53 80.9324
R20620 a_n2848_n452.n27 a_n2848_n452.t46 74.6477
R20621 a_n2848_n452.n24 a_n2848_n452.t26 74.6477
R20622 a_n2848_n452.n26 a_n2848_n452.t30 74.2899
R20623 a_n2848_n452.n25 a_n2848_n452.t34 74.2897
R20624 a_n2848_n452.n27 a_n2848_n452.n103 70.6783
R20625 a_n2848_n452.n25 a_n2848_n452.n72 70.6783
R20626 a_n2848_n452.n24 a_n2848_n452.n71 70.6783
R20627 a_n2848_n452.n104 a_n2848_n452.n27 70.6782
R20628 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R20629 a_n2848_n452.n95 a_n2848_n452.n49 20.9683
R20630 a_n2848_n452.n101 a_n2848_n452.n51 20.9683
R20631 a_n2848_n452.n98 a_n2848_n452.n46 20.9683
R20632 a_n2848_n452.n79 a_n2848_n452.n78 48.2005
R20633 a_n2848_n452.n80 a_n2848_n452.n36 20.9683
R20634 a_n2848_n452.n76 a_n2848_n452.n75 48.2005
R20635 a_n2848_n452.n77 a_n2848_n452.n33 20.9683
R20636 a_n2848_n452.n92 a_n2848_n452.n82 48.2005
R20637 a_n2848_n452.t69 a_n2848_n452.n45 533.335
R20638 a_n2848_n452.n90 a_n2848_n452.n83 48.2005
R20639 a_n2848_n452.t74 a_n2848_n452.n43 533.335
R20640 a_n2848_n452.n88 a_n2848_n452.n84 48.2005
R20641 a_n2848_n452.t63 a_n2848_n452.n41 533.335
R20642 a_n2848_n452.n86 a_n2848_n452.n85 48.2005
R20643 a_n2848_n452.t59 a_n2848_n452.n39 533.335
R20644 a_n2848_n452.n50 a_n2848_n452.t73 533.058
R20645 a_n2848_n452.n47 a_n2848_n452.t45 533.058
R20646 a_n2848_n452.t33 a_n2848_n452.n37 533.058
R20647 a_n2848_n452.t51 a_n2848_n452.n34 533.058
R20648 a_n2848_n452.n61 a_n2848_n452.n29 33.585
R20649 a_n2848_n452.n48 a_n2848_n452.n70 35.3134
R20650 a_n2848_n452.n100 a_n2848_n452.n99 24.1005
R20651 a_n2848_n452.n99 a_n2848_n452.n69 24.1005
R20652 a_n2848_n452.n73 a_n2848_n452.n35 35.3134
R20653 a_n2848_n452.n74 a_n2848_n452.n32 35.3134
R20654 a_n2848_n452.n93 a_n2848_n452.n44 35.3134
R20655 a_n2848_n452.n91 a_n2848_n452.n42 35.3134
R20656 a_n2848_n452.n89 a_n2848_n452.n40 35.3134
R20657 a_n2848_n452.n87 a_n2848_n452.n38 35.3134
R20658 a_n2848_n452.n0 a_n2848_n452.n31 23.891
R20659 a_n2848_n452.n22 a_n2848_n452.n13 12.046
R20660 a_n2848_n452.n3 a_n2848_n452.n94 11.8414
R20661 a_n2848_n452.n102 a_n2848_n452.n0 10.5365
R20662 a_n2848_n452.n81 a_n2848_n452.n25 9.50122
R20663 a_n2848_n452.n15 a_n2848_n452.n13 7.47588
R20664 a_n2848_n452.n94 a_n2848_n452.n7 7.47588
R20665 a_n2848_n452.n81 a_n2848_n452.n16 6.70126
R20666 a_n2848_n452.n26 a_n2848_n452.n102 5.65783
R20667 a_n2848_n452.n94 a_n2848_n452.n81 5.3452
R20668 a_n2848_n452.n18 a_n2848_n452.n20 3.95126
R20669 a_n2848_n452.n6 a_n2848_n452.n2 3.95126
R20670 a_n2848_n452.n103 a_n2848_n452.t32 3.61217
R20671 a_n2848_n452.n103 a_n2848_n452.t42 3.61217
R20672 a_n2848_n452.n72 a_n2848_n452.t28 3.61217
R20673 a_n2848_n452.n72 a_n2848_n452.t36 3.61217
R20674 a_n2848_n452.n71 a_n2848_n452.t44 3.61217
R20675 a_n2848_n452.n71 a_n2848_n452.t40 3.61217
R20676 a_n2848_n452.n104 a_n2848_n452.t38 3.61217
R20677 a_n2848_n452.t24 a_n2848_n452.n104 3.61217
R20678 a_n2848_n452.n65 a_n2848_n452.t6 2.82907
R20679 a_n2848_n452.n65 a_n2848_n452.t9 2.82907
R20680 a_n2848_n452.n66 a_n2848_n452.t1 2.82907
R20681 a_n2848_n452.n66 a_n2848_n452.t12 2.82907
R20682 a_n2848_n452.n68 a_n2848_n452.t15 2.82907
R20683 a_n2848_n452.n68 a_n2848_n452.t16 2.82907
R20684 a_n2848_n452.n64 a_n2848_n452.t10 2.82907
R20685 a_n2848_n452.n64 a_n2848_n452.t4 2.82907
R20686 a_n2848_n452.n62 a_n2848_n452.t0 2.82907
R20687 a_n2848_n452.n62 a_n2848_n452.t7 2.82907
R20688 a_n2848_n452.n60 a_n2848_n452.t14 2.82907
R20689 a_n2848_n452.n60 a_n2848_n452.t21 2.82907
R20690 a_n2848_n452.n56 a_n2848_n452.t20 2.82907
R20691 a_n2848_n452.n56 a_n2848_n452.t18 2.82907
R20692 a_n2848_n452.n57 a_n2848_n452.t11 2.82907
R20693 a_n2848_n452.n57 a_n2848_n452.t22 2.82907
R20694 a_n2848_n452.n59 a_n2848_n452.t8 2.82907
R20695 a_n2848_n452.n59 a_n2848_n452.t5 2.82907
R20696 a_n2848_n452.n55 a_n2848_n452.t47 2.82907
R20697 a_n2848_n452.n55 a_n2848_n452.t2 2.82907
R20698 a_n2848_n452.n53 a_n2848_n452.t13 2.82907
R20699 a_n2848_n452.n53 a_n2848_n452.t17 2.82907
R20700 a_n2848_n452.n52 a_n2848_n452.t3 2.82907
R20701 a_n2848_n452.n52 a_n2848_n452.t19 2.82907
R20702 a_n2848_n452.n102 a_n2848_n452.n13 1.30542
R20703 a_n2848_n452.n10 a_n2848_n452.n11 1.04595
R20704 a_n2848_n452.n5 a_n2848_n452.n97 13.657
R20705 a_n2848_n452.n95 a_n2848_n452.n50 21.4216
R20706 a_n2848_n452.n1 a_n2848_n452.n101 21.4216
R20707 a_n2848_n452.n98 a_n2848_n452.n47 21.4216
R20708 a_n2848_n452.n78 a_n2848_n452.n19 13.657
R20709 a_n2848_n452.n37 a_n2848_n452.n80 21.4216
R20710 a_n2848_n452.n75 a_n2848_n452.n23 13.657
R20711 a_n2848_n452.n34 a_n2848_n452.n77 21.4216
R20712 a_n2848_n452.n0 a_n2848_n452.n6 1.47777
R20713 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R20714 a_n2848_n452.n21 a_n2848_n452.n20 0.758076
R20715 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R20716 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R20717 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R20718 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R20719 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R20720 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R20721 a_n2848_n452.n4 a_n2848_n452.n2 0.758076
R20722 a_n2848_n452.n4 a_n2848_n452.n3 0.758076
R20723 a_n2848_n452.n27 a_n2848_n452.n26 0.716017
R20724 a_n2848_n452.n25 a_n2848_n452.n24 0.716017
R20725 a_n2848_n452.n12 a_n2848_n452.n14 0.67853
R20726 a_n2848_n452.n8 a_n2848_n452.n9 0.67853
R20727 a_n2848_n452.n28 a_n2848_n452.n54 0.530672
R20728 a_n2848_n452.n29 a_n2848_n452.n58 0.530672
R20729 a_n2848_n452.n63 a_n2848_n452.n61 0.530672
R20730 a_n2848_n452.n30 a_n2848_n452.n63 0.530672
R20731 a_n2848_n452.n31 a_n2848_n452.n67 0.530672
R20732 a_n2848_n452.n31 a_n2848_n452.n30 0.530672
R20733 a_n2848_n452.n29 a_n2848_n452.n28 0.530672
R20734 a_n1986_8322.n6 a_n1986_8322.t14 74.6477
R20735 a_n1986_8322.n1 a_n1986_8322.t1 74.6477
R20736 a_n1986_8322.n16 a_n1986_8322.t10 74.6474
R20737 a_n1986_8322.n14 a_n1986_8322.t3 74.2899
R20738 a_n1986_8322.n7 a_n1986_8322.t12 74.2899
R20739 a_n1986_8322.n8 a_n1986_8322.t15 74.2899
R20740 a_n1986_8322.n11 a_n1986_8322.t16 74.2899
R20741 a_n1986_8322.n4 a_n1986_8322.t0 74.2899
R20742 a_n1986_8322.n16 a_n1986_8322.n15 70.6783
R20743 a_n1986_8322.n6 a_n1986_8322.n5 70.6783
R20744 a_n1986_8322.n10 a_n1986_8322.n9 70.6783
R20745 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R20746 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R20747 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R20748 a_n1986_8322.n12 a_n1986_8322.n4 22.7556
R20749 a_n1986_8322.n13 a_n1986_8322.t22 9.7972
R20750 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R20751 a_n1986_8322.n14 a_n1986_8322.n13 5.83671
R20752 a_n1986_8322.n13 a_n1986_8322.n12 5.3452
R20753 a_n1986_8322.n15 a_n1986_8322.t8 3.61217
R20754 a_n1986_8322.n15 a_n1986_8322.t5 3.61217
R20755 a_n1986_8322.n5 a_n1986_8322.t18 3.61217
R20756 a_n1986_8322.n5 a_n1986_8322.t17 3.61217
R20757 a_n1986_8322.n9 a_n1986_8322.t13 3.61217
R20758 a_n1986_8322.n9 a_n1986_8322.t19 3.61217
R20759 a_n1986_8322.n0 a_n1986_8322.t9 3.61217
R20760 a_n1986_8322.n0 a_n1986_8322.t4 3.61217
R20761 a_n1986_8322.n2 a_n1986_8322.t7 3.61217
R20762 a_n1986_8322.n2 a_n1986_8322.t6 3.61217
R20763 a_n1986_8322.n18 a_n1986_8322.t2 3.61217
R20764 a_n1986_8322.t11 a_n1986_8322.n18 3.61217
R20765 a_n1986_8322.n11 a_n1986_8322.n10 0.358259
R20766 a_n1986_8322.n10 a_n1986_8322.n8 0.358259
R20767 a_n1986_8322.n7 a_n1986_8322.n6 0.358259
R20768 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R20769 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R20770 a_n1986_8322.n17 a_n1986_8322.n14 0.358259
R20771 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R20772 a_n1986_8322.n8 a_n1986_8322.n7 0.101793
R20773 a_n1986_8322.t23 a_n1986_8322.t20 0.0788333
R20774 a_n1986_8322.t21 a_n1986_8322.t23 0.0631667
R20775 a_n1986_8322.t22 a_n1986_8322.t21 0.0471944
R20776 a_n1986_8322.t22 a_n1986_8322.t20 0.0453889
R20777 a_n1808_13878.n5 a_n1808_13878.n3 98.9633
R20778 a_n1808_13878.n2 a_n1808_13878.n0 98.7517
R20779 a_n1808_13878.n2 a_n1808_13878.n1 98.6055
R20780 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20781 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20782 a_n1808_13878.n7 a_n1808_13878.n6 98.6054
R20783 a_n1808_13878.n9 a_n1808_13878.t13 74.6477
R20784 a_n1808_13878.n14 a_n1808_13878.t14 74.2899
R20785 a_n1808_13878.n11 a_n1808_13878.t15 74.2899
R20786 a_n1808_13878.n10 a_n1808_13878.t12 74.2899
R20787 a_n1808_13878.n13 a_n1808_13878.n12 70.6783
R20788 a_n1808_13878.n9 a_n1808_13878.n8 70.6783
R20789 a_n1808_13878.n16 a_n1808_13878.n15 13.5694
R20790 a_n1808_13878.n15 a_n1808_13878.n7 11.5762
R20791 a_n1808_13878.n15 a_n1808_13878.n14 6.2408
R20792 a_n1808_13878.n1 a_n1808_13878.t6 3.61217
R20793 a_n1808_13878.n1 a_n1808_13878.t1 3.61217
R20794 a_n1808_13878.n0 a_n1808_13878.t0 3.61217
R20795 a_n1808_13878.n0 a_n1808_13878.t2 3.61217
R20796 a_n1808_13878.n6 a_n1808_13878.t7 3.61217
R20797 a_n1808_13878.n6 a_n1808_13878.t8 3.61217
R20798 a_n1808_13878.n4 a_n1808_13878.t10 3.61217
R20799 a_n1808_13878.n4 a_n1808_13878.t3 3.61217
R20800 a_n1808_13878.n3 a_n1808_13878.t5 3.61217
R20801 a_n1808_13878.n3 a_n1808_13878.t9 3.61217
R20802 a_n1808_13878.n12 a_n1808_13878.t18 3.61217
R20803 a_n1808_13878.n12 a_n1808_13878.t19 3.61217
R20804 a_n1808_13878.n8 a_n1808_13878.t16 3.61217
R20805 a_n1808_13878.n8 a_n1808_13878.t17 3.61217
R20806 a_n1808_13878.n17 a_n1808_13878.t4 3.61217
R20807 a_n1808_13878.t11 a_n1808_13878.n17 3.61217
R20808 a_n1808_13878.n7 a_n1808_13878.n5 0.358259
R20809 a_n1808_13878.n10 a_n1808_13878.n9 0.358259
R20810 a_n1808_13878.n13 a_n1808_13878.n11 0.358259
R20811 a_n1808_13878.n14 a_n1808_13878.n13 0.358259
R20812 a_n1808_13878.n16 a_n1808_13878.n2 0.146627
R20813 a_n1808_13878.n11 a_n1808_13878.n10 0.101793
R20814 plus.n76 plus.t11 250.337
R20815 plus.n15 plus.t14 250.337
R20816 plus.n124 plus.t1 243.97
R20817 plus.n120 plus.t24 231.093
R20818 plus.n59 plus.t20 231.093
R20819 plus.n124 plus.n123 223.454
R20820 plus.n126 plus.n125 223.454
R20821 plus.n77 plus.t5 187.445
R20822 plus.n74 plus.t22 187.445
R20823 plus.n72 plus.t21 187.445
R20824 plus.n89 plus.t16 187.445
R20825 plus.n95 plus.t17 187.445
R20826 plus.n68 plus.t13 187.445
R20827 plus.n66 plus.t15 187.445
R20828 plus.n107 plus.t10 187.445
R20829 plus.n113 plus.t26 187.445
R20830 plus.n62 plus.t28 187.445
R20831 plus.n1 plus.t23 187.445
R20832 plus.n52 plus.t6 187.445
R20833 plus.n46 plus.t12 187.445
R20834 plus.n5 plus.t8 187.445
R20835 plus.n7 plus.t7 187.445
R20836 plus.n34 plus.t19 187.445
R20837 plus.n28 plus.t18 187.445
R20838 plus.n11 plus.t27 187.445
R20839 plus.n13 plus.t25 187.445
R20840 plus.n16 plus.t9 187.445
R20841 plus.n121 plus.n120 161.3
R20842 plus.n119 plus.n61 161.3
R20843 plus.n118 plus.n117 161.3
R20844 plus.n116 plus.n115 161.3
R20845 plus.n114 plus.n63 161.3
R20846 plus.n112 plus.n111 161.3
R20847 plus.n110 plus.n64 161.3
R20848 plus.n109 plus.n108 161.3
R20849 plus.n106 plus.n65 161.3
R20850 plus.n105 plus.n104 161.3
R20851 plus.n103 plus.n102 161.3
R20852 plus.n101 plus.n67 161.3
R20853 plus.n100 plus.n99 161.3
R20854 plus.n98 plus.n97 161.3
R20855 plus.n96 plus.n69 161.3
R20856 plus.n94 plus.n93 161.3
R20857 plus.n92 plus.n70 161.3
R20858 plus.n91 plus.n90 161.3
R20859 plus.n88 plus.n71 161.3
R20860 plus.n87 plus.n86 161.3
R20861 plus.n85 plus.n84 161.3
R20862 plus.n83 plus.n73 161.3
R20863 plus.n82 plus.n81 161.3
R20864 plus.n80 plus.n79 161.3
R20865 plus.n78 plus.n75 161.3
R20866 plus.n17 plus.n14 161.3
R20867 plus.n19 plus.n18 161.3
R20868 plus.n21 plus.n20 161.3
R20869 plus.n22 plus.n12 161.3
R20870 plus.n24 plus.n23 161.3
R20871 plus.n26 plus.n25 161.3
R20872 plus.n27 plus.n10 161.3
R20873 plus.n30 plus.n29 161.3
R20874 plus.n31 plus.n9 161.3
R20875 plus.n33 plus.n32 161.3
R20876 plus.n35 plus.n8 161.3
R20877 plus.n37 plus.n36 161.3
R20878 plus.n39 plus.n38 161.3
R20879 plus.n40 plus.n6 161.3
R20880 plus.n42 plus.n41 161.3
R20881 plus.n44 plus.n43 161.3
R20882 plus.n45 plus.n4 161.3
R20883 plus.n48 plus.n47 161.3
R20884 plus.n49 plus.n3 161.3
R20885 plus.n51 plus.n50 161.3
R20886 plus.n53 plus.n2 161.3
R20887 plus.n55 plus.n54 161.3
R20888 plus.n57 plus.n56 161.3
R20889 plus.n58 plus.n0 161.3
R20890 plus.n60 plus.n59 161.3
R20891 plus.n88 plus.n87 56.5617
R20892 plus.n97 plus.n96 56.5617
R20893 plus.n106 plus.n105 56.5617
R20894 plus.n45 plus.n44 56.5617
R20895 plus.n36 plus.n35 56.5617
R20896 plus.n27 plus.n26 56.5617
R20897 plus.n79 plus.n78 56.5617
R20898 plus.n115 plus.n114 56.5617
R20899 plus.n54 plus.n53 56.5617
R20900 plus.n18 plus.n17 56.5617
R20901 plus.n119 plus.n118 50.2647
R20902 plus.n58 plus.n57 50.2647
R20903 plus.n84 plus.n83 46.3896
R20904 plus.n108 plus.n64 46.3896
R20905 plus.n47 plus.n3 46.3896
R20906 plus.n23 plus.n22 46.3896
R20907 plus.n76 plus.n75 43.1929
R20908 plus.n15 plus.n14 43.1929
R20909 plus.n94 plus.n70 42.5146
R20910 plus.n101 plus.n100 42.5146
R20911 plus.n40 plus.n39 42.5146
R20912 plus.n33 plus.n9 42.5146
R20913 plus.n77 plus.n76 40.6041
R20914 plus.n16 plus.n15 40.6041
R20915 plus.n90 plus.n70 38.6395
R20916 plus.n102 plus.n101 38.6395
R20917 plus.n41 plus.n40 38.6395
R20918 plus.n29 plus.n9 38.6395
R20919 plus.n122 plus.n121 35.2031
R20920 plus.n83 plus.n82 34.7644
R20921 plus.n112 plus.n64 34.7644
R20922 plus.n51 plus.n3 34.7644
R20923 plus.n22 plus.n21 34.7644
R20924 plus.n79 plus.n74 21.8872
R20925 plus.n114 plus.n113 21.8872
R20926 plus.n53 plus.n52 21.8872
R20927 plus.n18 plus.n13 21.8872
R20928 plus.n89 plus.n88 19.9199
R20929 plus.n105 plus.n66 19.9199
R20930 plus.n44 plus.n5 19.9199
R20931 plus.n28 plus.n27 19.9199
R20932 plus.n123 plus.t2 19.8005
R20933 plus.n123 plus.t4 19.8005
R20934 plus.n125 plus.t3 19.8005
R20935 plus.n125 plus.t0 19.8005
R20936 plus.n96 plus.n95 17.9525
R20937 plus.n97 plus.n68 17.9525
R20938 plus.n36 plus.n7 17.9525
R20939 plus.n35 plus.n34 17.9525
R20940 plus.n87 plus.n72 15.9852
R20941 plus.n107 plus.n106 15.9852
R20942 plus.n46 plus.n45 15.9852
R20943 plus.n26 plus.n11 15.9852
R20944 plus plus.n127 14.4034
R20945 plus.n78 plus.n77 14.0178
R20946 plus.n115 plus.n62 14.0178
R20947 plus.n54 plus.n1 14.0178
R20948 plus.n17 plus.n16 14.0178
R20949 plus.n122 plus.n60 11.9342
R20950 plus.n118 plus.n62 10.575
R20951 plus.n57 plus.n1 10.575
R20952 plus.n120 plus.n119 9.49444
R20953 plus.n59 plus.n58 9.49444
R20954 plus.n84 plus.n72 8.60764
R20955 plus.n108 plus.n107 8.60764
R20956 plus.n47 plus.n46 8.60764
R20957 plus.n23 plus.n11 8.60764
R20958 plus.n95 plus.n94 6.6403
R20959 plus.n100 plus.n68 6.6403
R20960 plus.n39 plus.n7 6.6403
R20961 plus.n34 plus.n33 6.6403
R20962 plus.n127 plus.n126 5.40567
R20963 plus.n90 plus.n89 4.67295
R20964 plus.n102 plus.n66 4.67295
R20965 plus.n41 plus.n5 4.67295
R20966 plus.n29 plus.n28 4.67295
R20967 plus.n82 plus.n74 2.7056
R20968 plus.n113 plus.n112 2.7056
R20969 plus.n52 plus.n51 2.7056
R20970 plus.n21 plus.n13 2.7056
R20971 plus.n127 plus.n122 1.188
R20972 plus.n126 plus.n124 0.716017
R20973 plus.n80 plus.n75 0.189894
R20974 plus.n81 plus.n80 0.189894
R20975 plus.n81 plus.n73 0.189894
R20976 plus.n85 plus.n73 0.189894
R20977 plus.n86 plus.n85 0.189894
R20978 plus.n86 plus.n71 0.189894
R20979 plus.n91 plus.n71 0.189894
R20980 plus.n92 plus.n91 0.189894
R20981 plus.n93 plus.n92 0.189894
R20982 plus.n93 plus.n69 0.189894
R20983 plus.n98 plus.n69 0.189894
R20984 plus.n99 plus.n98 0.189894
R20985 plus.n99 plus.n67 0.189894
R20986 plus.n103 plus.n67 0.189894
R20987 plus.n104 plus.n103 0.189894
R20988 plus.n104 plus.n65 0.189894
R20989 plus.n109 plus.n65 0.189894
R20990 plus.n110 plus.n109 0.189894
R20991 plus.n111 plus.n110 0.189894
R20992 plus.n111 plus.n63 0.189894
R20993 plus.n116 plus.n63 0.189894
R20994 plus.n117 plus.n116 0.189894
R20995 plus.n117 plus.n61 0.189894
R20996 plus.n121 plus.n61 0.189894
R20997 plus.n60 plus.n0 0.189894
R20998 plus.n56 plus.n0 0.189894
R20999 plus.n56 plus.n55 0.189894
R21000 plus.n55 plus.n2 0.189894
R21001 plus.n50 plus.n2 0.189894
R21002 plus.n50 plus.n49 0.189894
R21003 plus.n49 plus.n48 0.189894
R21004 plus.n48 plus.n4 0.189894
R21005 plus.n43 plus.n4 0.189894
R21006 plus.n43 plus.n42 0.189894
R21007 plus.n42 plus.n6 0.189894
R21008 plus.n38 plus.n6 0.189894
R21009 plus.n38 plus.n37 0.189894
R21010 plus.n37 plus.n8 0.189894
R21011 plus.n32 plus.n8 0.189894
R21012 plus.n32 plus.n31 0.189894
R21013 plus.n31 plus.n30 0.189894
R21014 plus.n30 plus.n10 0.189894
R21015 plus.n25 plus.n10 0.189894
R21016 plus.n25 plus.n24 0.189894
R21017 plus.n24 plus.n12 0.189894
R21018 plus.n20 plus.n12 0.189894
R21019 plus.n20 plus.n19 0.189894
R21020 plus.n19 plus.n14 0.189894
R21021 a_n3106_n452.n1 a_n3106_n452.t31 214.321
R21022 a_n3106_n452.n14 a_n3106_n452.t40 214.321
R21023 a_n3106_n452.n15 a_n3106_n452.t32 214.321
R21024 a_n3106_n452.n16 a_n3106_n452.t39 214.321
R21025 a_n3106_n452.n17 a_n3106_n452.t28 214.321
R21026 a_n3106_n452.n18 a_n3106_n452.t0 214.321
R21027 a_n3106_n452.n19 a_n3106_n452.t43 214.321
R21028 a_n3106_n452.n20 a_n3106_n452.t41 214.321
R21029 a_n3106_n452.n0 a_n3106_n452.t21 55.8337
R21030 a_n3106_n452.n2 a_n3106_n452.t37 55.8337
R21031 a_n3106_n452.n13 a_n3106_n452.t46 55.8337
R21032 a_n3106_n452.n47 a_n3106_n452.t8 55.8335
R21033 a_n3106_n452.n45 a_n3106_n452.t50 55.8335
R21034 a_n3106_n452.n34 a_n3106_n452.t29 55.8335
R21035 a_n3106_n452.n33 a_n3106_n452.t18 55.8335
R21036 a_n3106_n452.n22 a_n3106_n452.t12 55.8335
R21037 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R21038 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R21039 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R21040 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R21041 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R21042 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R21043 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R21044 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R21045 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R21046 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R21047 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R21048 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R21049 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R21050 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R21051 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R21052 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R21053 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R21054 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R21055 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R21056 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R21057 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R21058 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R21059 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R21060 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R21061 a_n3106_n452.n48 a_n3106_n452.t6 2.82907
R21062 a_n3106_n452.n48 a_n3106_n452.t4 2.82907
R21063 a_n3106_n452.n50 a_n3106_n452.t17 2.82907
R21064 a_n3106_n452.n50 a_n3106_n452.t22 2.82907
R21065 a_n3106_n452.n52 a_n3106_n452.t15 2.82907
R21066 a_n3106_n452.n52 a_n3106_n452.t19 2.82907
R21067 a_n3106_n452.n54 a_n3106_n452.t11 2.82907
R21068 a_n3106_n452.n54 a_n3106_n452.t16 2.82907
R21069 a_n3106_n452.n3 a_n3106_n452.t44 2.82907
R21070 a_n3106_n452.n3 a_n3106_n452.t34 2.82907
R21071 a_n3106_n452.n5 a_n3106_n452.t48 2.82907
R21072 a_n3106_n452.n5 a_n3106_n452.t2 2.82907
R21073 a_n3106_n452.n7 a_n3106_n452.t30 2.82907
R21074 a_n3106_n452.n7 a_n3106_n452.t47 2.82907
R21075 a_n3106_n452.n9 a_n3106_n452.t35 2.82907
R21076 a_n3106_n452.n9 a_n3106_n452.t38 2.82907
R21077 a_n3106_n452.n11 a_n3106_n452.t53 2.82907
R21078 a_n3106_n452.n11 a_n3106_n452.t1 2.82907
R21079 a_n3106_n452.n43 a_n3106_n452.t54 2.82907
R21080 a_n3106_n452.n43 a_n3106_n452.t52 2.82907
R21081 a_n3106_n452.n41 a_n3106_n452.t33 2.82907
R21082 a_n3106_n452.n41 a_n3106_n452.t42 2.82907
R21083 a_n3106_n452.n39 a_n3106_n452.t3 2.82907
R21084 a_n3106_n452.n39 a_n3106_n452.t36 2.82907
R21085 a_n3106_n452.n37 a_n3106_n452.t49 2.82907
R21086 a_n3106_n452.n37 a_n3106_n452.t55 2.82907
R21087 a_n3106_n452.n35 a_n3106_n452.t51 2.82907
R21088 a_n3106_n452.n35 a_n3106_n452.t45 2.82907
R21089 a_n3106_n452.n31 a_n3106_n452.t7 2.82907
R21090 a_n3106_n452.n31 a_n3106_n452.t23 2.82907
R21091 a_n3106_n452.n29 a_n3106_n452.t14 2.82907
R21092 a_n3106_n452.n29 a_n3106_n452.t5 2.82907
R21093 a_n3106_n452.n27 a_n3106_n452.t25 2.82907
R21094 a_n3106_n452.n27 a_n3106_n452.t13 2.82907
R21095 a_n3106_n452.n25 a_n3106_n452.t20 2.82907
R21096 a_n3106_n452.n25 a_n3106_n452.t24 2.82907
R21097 a_n3106_n452.n23 a_n3106_n452.t9 2.82907
R21098 a_n3106_n452.n23 a_n3106_n452.t26 2.82907
R21099 a_n3106_n452.t27 a_n3106_n452.n57 2.82907
R21100 a_n3106_n452.n57 a_n3106_n452.t10 2.82907
R21101 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R21102 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R21103 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R21104 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R21105 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R21106 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R21107 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R21108 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R21109 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R21110 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R21111 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R21112 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R21113 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R21114 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R21115 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R21116 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R21117 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R21118 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R21119 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R21120 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R21121 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R21122 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R21123 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R21124 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R21125 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R21126 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R21127 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R21128 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R21129 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R21130 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R21131 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R21132 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R21133 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R21134 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R21135 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R21136 outputibias.n27 outputibias.n1 289.615
R21137 outputibias.n58 outputibias.n32 289.615
R21138 outputibias.n90 outputibias.n64 289.615
R21139 outputibias.n122 outputibias.n96 289.615
R21140 outputibias.n28 outputibias.n27 185
R21141 outputibias.n26 outputibias.n25 185
R21142 outputibias.n5 outputibias.n4 185
R21143 outputibias.n20 outputibias.n19 185
R21144 outputibias.n18 outputibias.n17 185
R21145 outputibias.n9 outputibias.n8 185
R21146 outputibias.n12 outputibias.n11 185
R21147 outputibias.n59 outputibias.n58 185
R21148 outputibias.n57 outputibias.n56 185
R21149 outputibias.n36 outputibias.n35 185
R21150 outputibias.n51 outputibias.n50 185
R21151 outputibias.n49 outputibias.n48 185
R21152 outputibias.n40 outputibias.n39 185
R21153 outputibias.n43 outputibias.n42 185
R21154 outputibias.n91 outputibias.n90 185
R21155 outputibias.n89 outputibias.n88 185
R21156 outputibias.n68 outputibias.n67 185
R21157 outputibias.n83 outputibias.n82 185
R21158 outputibias.n81 outputibias.n80 185
R21159 outputibias.n72 outputibias.n71 185
R21160 outputibias.n75 outputibias.n74 185
R21161 outputibias.n123 outputibias.n122 185
R21162 outputibias.n121 outputibias.n120 185
R21163 outputibias.n100 outputibias.n99 185
R21164 outputibias.n115 outputibias.n114 185
R21165 outputibias.n113 outputibias.n112 185
R21166 outputibias.n104 outputibias.n103 185
R21167 outputibias.n107 outputibias.n106 185
R21168 outputibias.n0 outputibias.t8 178.945
R21169 outputibias.n133 outputibias.t10 177.018
R21170 outputibias.n132 outputibias.t11 177.018
R21171 outputibias.n0 outputibias.t9 177.018
R21172 outputibias.t5 outputibias.n10 147.661
R21173 outputibias.t7 outputibias.n41 147.661
R21174 outputibias.t1 outputibias.n73 147.661
R21175 outputibias.t3 outputibias.n105 147.661
R21176 outputibias.n128 outputibias.t4 132.363
R21177 outputibias.n128 outputibias.t6 130.436
R21178 outputibias.n129 outputibias.t0 130.436
R21179 outputibias.n130 outputibias.t2 130.436
R21180 outputibias.n27 outputibias.n26 104.615
R21181 outputibias.n26 outputibias.n4 104.615
R21182 outputibias.n19 outputibias.n4 104.615
R21183 outputibias.n19 outputibias.n18 104.615
R21184 outputibias.n18 outputibias.n8 104.615
R21185 outputibias.n11 outputibias.n8 104.615
R21186 outputibias.n58 outputibias.n57 104.615
R21187 outputibias.n57 outputibias.n35 104.615
R21188 outputibias.n50 outputibias.n35 104.615
R21189 outputibias.n50 outputibias.n49 104.615
R21190 outputibias.n49 outputibias.n39 104.615
R21191 outputibias.n42 outputibias.n39 104.615
R21192 outputibias.n90 outputibias.n89 104.615
R21193 outputibias.n89 outputibias.n67 104.615
R21194 outputibias.n82 outputibias.n67 104.615
R21195 outputibias.n82 outputibias.n81 104.615
R21196 outputibias.n81 outputibias.n71 104.615
R21197 outputibias.n74 outputibias.n71 104.615
R21198 outputibias.n122 outputibias.n121 104.615
R21199 outputibias.n121 outputibias.n99 104.615
R21200 outputibias.n114 outputibias.n99 104.615
R21201 outputibias.n114 outputibias.n113 104.615
R21202 outputibias.n113 outputibias.n103 104.615
R21203 outputibias.n106 outputibias.n103 104.615
R21204 outputibias.n63 outputibias.n31 95.6354
R21205 outputibias.n63 outputibias.n62 94.6732
R21206 outputibias.n95 outputibias.n94 94.6732
R21207 outputibias.n127 outputibias.n126 94.6732
R21208 outputibias.n11 outputibias.t5 52.3082
R21209 outputibias.n42 outputibias.t7 52.3082
R21210 outputibias.n74 outputibias.t1 52.3082
R21211 outputibias.n106 outputibias.t3 52.3082
R21212 outputibias.n12 outputibias.n10 15.6674
R21213 outputibias.n43 outputibias.n41 15.6674
R21214 outputibias.n75 outputibias.n73 15.6674
R21215 outputibias.n107 outputibias.n105 15.6674
R21216 outputibias.n13 outputibias.n9 12.8005
R21217 outputibias.n44 outputibias.n40 12.8005
R21218 outputibias.n76 outputibias.n72 12.8005
R21219 outputibias.n108 outputibias.n104 12.8005
R21220 outputibias.n17 outputibias.n16 12.0247
R21221 outputibias.n48 outputibias.n47 12.0247
R21222 outputibias.n80 outputibias.n79 12.0247
R21223 outputibias.n112 outputibias.n111 12.0247
R21224 outputibias.n20 outputibias.n7 11.249
R21225 outputibias.n51 outputibias.n38 11.249
R21226 outputibias.n83 outputibias.n70 11.249
R21227 outputibias.n115 outputibias.n102 11.249
R21228 outputibias.n21 outputibias.n5 10.4732
R21229 outputibias.n52 outputibias.n36 10.4732
R21230 outputibias.n84 outputibias.n68 10.4732
R21231 outputibias.n116 outputibias.n100 10.4732
R21232 outputibias.n25 outputibias.n24 9.69747
R21233 outputibias.n56 outputibias.n55 9.69747
R21234 outputibias.n88 outputibias.n87 9.69747
R21235 outputibias.n120 outputibias.n119 9.69747
R21236 outputibias.n31 outputibias.n30 9.45567
R21237 outputibias.n62 outputibias.n61 9.45567
R21238 outputibias.n94 outputibias.n93 9.45567
R21239 outputibias.n126 outputibias.n125 9.45567
R21240 outputibias.n30 outputibias.n29 9.3005
R21241 outputibias.n3 outputibias.n2 9.3005
R21242 outputibias.n24 outputibias.n23 9.3005
R21243 outputibias.n22 outputibias.n21 9.3005
R21244 outputibias.n7 outputibias.n6 9.3005
R21245 outputibias.n16 outputibias.n15 9.3005
R21246 outputibias.n14 outputibias.n13 9.3005
R21247 outputibias.n61 outputibias.n60 9.3005
R21248 outputibias.n34 outputibias.n33 9.3005
R21249 outputibias.n55 outputibias.n54 9.3005
R21250 outputibias.n53 outputibias.n52 9.3005
R21251 outputibias.n38 outputibias.n37 9.3005
R21252 outputibias.n47 outputibias.n46 9.3005
R21253 outputibias.n45 outputibias.n44 9.3005
R21254 outputibias.n93 outputibias.n92 9.3005
R21255 outputibias.n66 outputibias.n65 9.3005
R21256 outputibias.n87 outputibias.n86 9.3005
R21257 outputibias.n85 outputibias.n84 9.3005
R21258 outputibias.n70 outputibias.n69 9.3005
R21259 outputibias.n79 outputibias.n78 9.3005
R21260 outputibias.n77 outputibias.n76 9.3005
R21261 outputibias.n125 outputibias.n124 9.3005
R21262 outputibias.n98 outputibias.n97 9.3005
R21263 outputibias.n119 outputibias.n118 9.3005
R21264 outputibias.n117 outputibias.n116 9.3005
R21265 outputibias.n102 outputibias.n101 9.3005
R21266 outputibias.n111 outputibias.n110 9.3005
R21267 outputibias.n109 outputibias.n108 9.3005
R21268 outputibias.n28 outputibias.n3 8.92171
R21269 outputibias.n59 outputibias.n34 8.92171
R21270 outputibias.n91 outputibias.n66 8.92171
R21271 outputibias.n123 outputibias.n98 8.92171
R21272 outputibias.n29 outputibias.n1 8.14595
R21273 outputibias.n60 outputibias.n32 8.14595
R21274 outputibias.n92 outputibias.n64 8.14595
R21275 outputibias.n124 outputibias.n96 8.14595
R21276 outputibias.n31 outputibias.n1 5.81868
R21277 outputibias.n62 outputibias.n32 5.81868
R21278 outputibias.n94 outputibias.n64 5.81868
R21279 outputibias.n126 outputibias.n96 5.81868
R21280 outputibias.n131 outputibias.n130 5.20947
R21281 outputibias.n29 outputibias.n28 5.04292
R21282 outputibias.n60 outputibias.n59 5.04292
R21283 outputibias.n92 outputibias.n91 5.04292
R21284 outputibias.n124 outputibias.n123 5.04292
R21285 outputibias.n131 outputibias.n127 4.42209
R21286 outputibias.n14 outputibias.n10 4.38594
R21287 outputibias.n45 outputibias.n41 4.38594
R21288 outputibias.n77 outputibias.n73 4.38594
R21289 outputibias.n109 outputibias.n105 4.38594
R21290 outputibias.n132 outputibias.n131 4.28454
R21291 outputibias.n25 outputibias.n3 4.26717
R21292 outputibias.n56 outputibias.n34 4.26717
R21293 outputibias.n88 outputibias.n66 4.26717
R21294 outputibias.n120 outputibias.n98 4.26717
R21295 outputibias.n24 outputibias.n5 3.49141
R21296 outputibias.n55 outputibias.n36 3.49141
R21297 outputibias.n87 outputibias.n68 3.49141
R21298 outputibias.n119 outputibias.n100 3.49141
R21299 outputibias.n21 outputibias.n20 2.71565
R21300 outputibias.n52 outputibias.n51 2.71565
R21301 outputibias.n84 outputibias.n83 2.71565
R21302 outputibias.n116 outputibias.n115 2.71565
R21303 outputibias.n17 outputibias.n7 1.93989
R21304 outputibias.n48 outputibias.n38 1.93989
R21305 outputibias.n80 outputibias.n70 1.93989
R21306 outputibias.n112 outputibias.n102 1.93989
R21307 outputibias.n130 outputibias.n129 1.9266
R21308 outputibias.n129 outputibias.n128 1.9266
R21309 outputibias.n133 outputibias.n132 1.92658
R21310 outputibias.n134 outputibias.n133 1.29913
R21311 outputibias.n16 outputibias.n9 1.16414
R21312 outputibias.n47 outputibias.n40 1.16414
R21313 outputibias.n79 outputibias.n72 1.16414
R21314 outputibias.n111 outputibias.n104 1.16414
R21315 outputibias.n127 outputibias.n95 0.962709
R21316 outputibias.n95 outputibias.n63 0.962709
R21317 outputibias.n13 outputibias.n12 0.388379
R21318 outputibias.n44 outputibias.n43 0.388379
R21319 outputibias.n76 outputibias.n75 0.388379
R21320 outputibias.n108 outputibias.n107 0.388379
R21321 outputibias.n134 outputibias.n0 0.337251
R21322 outputibias outputibias.n134 0.302375
R21323 outputibias.n30 outputibias.n2 0.155672
R21324 outputibias.n23 outputibias.n2 0.155672
R21325 outputibias.n23 outputibias.n22 0.155672
R21326 outputibias.n22 outputibias.n6 0.155672
R21327 outputibias.n15 outputibias.n6 0.155672
R21328 outputibias.n15 outputibias.n14 0.155672
R21329 outputibias.n61 outputibias.n33 0.155672
R21330 outputibias.n54 outputibias.n33 0.155672
R21331 outputibias.n54 outputibias.n53 0.155672
R21332 outputibias.n53 outputibias.n37 0.155672
R21333 outputibias.n46 outputibias.n37 0.155672
R21334 outputibias.n46 outputibias.n45 0.155672
R21335 outputibias.n93 outputibias.n65 0.155672
R21336 outputibias.n86 outputibias.n65 0.155672
R21337 outputibias.n86 outputibias.n85 0.155672
R21338 outputibias.n85 outputibias.n69 0.155672
R21339 outputibias.n78 outputibias.n69 0.155672
R21340 outputibias.n78 outputibias.n77 0.155672
R21341 outputibias.n125 outputibias.n97 0.155672
R21342 outputibias.n118 outputibias.n97 0.155672
R21343 outputibias.n118 outputibias.n117 0.155672
R21344 outputibias.n117 outputibias.n101 0.155672
R21345 outputibias.n110 outputibias.n101 0.155672
R21346 outputibias.n110 outputibias.n109 0.155672
R21347 output.n41 output.n15 289.615
R21348 output.n72 output.n46 289.615
R21349 output.n104 output.n78 289.615
R21350 output.n136 output.n110 289.615
R21351 output.n77 output.n45 197.26
R21352 output.n77 output.n76 196.298
R21353 output.n109 output.n108 196.298
R21354 output.n141 output.n140 196.298
R21355 output.n42 output.n41 185
R21356 output.n40 output.n39 185
R21357 output.n19 output.n18 185
R21358 output.n34 output.n33 185
R21359 output.n32 output.n31 185
R21360 output.n23 output.n22 185
R21361 output.n26 output.n25 185
R21362 output.n73 output.n72 185
R21363 output.n71 output.n70 185
R21364 output.n50 output.n49 185
R21365 output.n65 output.n64 185
R21366 output.n63 output.n62 185
R21367 output.n54 output.n53 185
R21368 output.n57 output.n56 185
R21369 output.n105 output.n104 185
R21370 output.n103 output.n102 185
R21371 output.n82 output.n81 185
R21372 output.n97 output.n96 185
R21373 output.n95 output.n94 185
R21374 output.n86 output.n85 185
R21375 output.n89 output.n88 185
R21376 output.n137 output.n136 185
R21377 output.n135 output.n134 185
R21378 output.n114 output.n113 185
R21379 output.n129 output.n128 185
R21380 output.n127 output.n126 185
R21381 output.n118 output.n117 185
R21382 output.n121 output.n120 185
R21383 output.t3 output.n24 147.661
R21384 output.t2 output.n55 147.661
R21385 output.t1 output.n87 147.661
R21386 output.t0 output.n119 147.661
R21387 output.n41 output.n40 104.615
R21388 output.n40 output.n18 104.615
R21389 output.n33 output.n18 104.615
R21390 output.n33 output.n32 104.615
R21391 output.n32 output.n22 104.615
R21392 output.n25 output.n22 104.615
R21393 output.n72 output.n71 104.615
R21394 output.n71 output.n49 104.615
R21395 output.n64 output.n49 104.615
R21396 output.n64 output.n63 104.615
R21397 output.n63 output.n53 104.615
R21398 output.n56 output.n53 104.615
R21399 output.n104 output.n103 104.615
R21400 output.n103 output.n81 104.615
R21401 output.n96 output.n81 104.615
R21402 output.n96 output.n95 104.615
R21403 output.n95 output.n85 104.615
R21404 output.n88 output.n85 104.615
R21405 output.n136 output.n135 104.615
R21406 output.n135 output.n113 104.615
R21407 output.n128 output.n113 104.615
R21408 output.n128 output.n127 104.615
R21409 output.n127 output.n117 104.615
R21410 output.n120 output.n117 104.615
R21411 output.n1 output.t19 77.056
R21412 output.n14 output.t4 76.6694
R21413 output.n1 output.n0 72.7095
R21414 output.n3 output.n2 72.7095
R21415 output.n5 output.n4 72.7095
R21416 output.n7 output.n6 72.7095
R21417 output.n9 output.n8 72.7095
R21418 output.n11 output.n10 72.7095
R21419 output.n13 output.n12 72.7095
R21420 output.n25 output.t3 52.3082
R21421 output.n56 output.t2 52.3082
R21422 output.n88 output.t1 52.3082
R21423 output.n120 output.t0 52.3082
R21424 output.n26 output.n24 15.6674
R21425 output.n57 output.n55 15.6674
R21426 output.n89 output.n87 15.6674
R21427 output.n121 output.n119 15.6674
R21428 output.n27 output.n23 12.8005
R21429 output.n58 output.n54 12.8005
R21430 output.n90 output.n86 12.8005
R21431 output.n122 output.n118 12.8005
R21432 output.n31 output.n30 12.0247
R21433 output.n62 output.n61 12.0247
R21434 output.n94 output.n93 12.0247
R21435 output.n126 output.n125 12.0247
R21436 output.n34 output.n21 11.249
R21437 output.n65 output.n52 11.249
R21438 output.n97 output.n84 11.249
R21439 output.n129 output.n116 11.249
R21440 output.n35 output.n19 10.4732
R21441 output.n66 output.n50 10.4732
R21442 output.n98 output.n82 10.4732
R21443 output.n130 output.n114 10.4732
R21444 output.n39 output.n38 9.69747
R21445 output.n70 output.n69 9.69747
R21446 output.n102 output.n101 9.69747
R21447 output.n134 output.n133 9.69747
R21448 output.n45 output.n44 9.45567
R21449 output.n76 output.n75 9.45567
R21450 output.n108 output.n107 9.45567
R21451 output.n140 output.n139 9.45567
R21452 output.n44 output.n43 9.3005
R21453 output.n17 output.n16 9.3005
R21454 output.n38 output.n37 9.3005
R21455 output.n36 output.n35 9.3005
R21456 output.n21 output.n20 9.3005
R21457 output.n30 output.n29 9.3005
R21458 output.n28 output.n27 9.3005
R21459 output.n75 output.n74 9.3005
R21460 output.n48 output.n47 9.3005
R21461 output.n69 output.n68 9.3005
R21462 output.n67 output.n66 9.3005
R21463 output.n52 output.n51 9.3005
R21464 output.n61 output.n60 9.3005
R21465 output.n59 output.n58 9.3005
R21466 output.n107 output.n106 9.3005
R21467 output.n80 output.n79 9.3005
R21468 output.n101 output.n100 9.3005
R21469 output.n99 output.n98 9.3005
R21470 output.n84 output.n83 9.3005
R21471 output.n93 output.n92 9.3005
R21472 output.n91 output.n90 9.3005
R21473 output.n139 output.n138 9.3005
R21474 output.n112 output.n111 9.3005
R21475 output.n133 output.n132 9.3005
R21476 output.n131 output.n130 9.3005
R21477 output.n116 output.n115 9.3005
R21478 output.n125 output.n124 9.3005
R21479 output.n123 output.n122 9.3005
R21480 output.n42 output.n17 8.92171
R21481 output.n73 output.n48 8.92171
R21482 output.n105 output.n80 8.92171
R21483 output.n137 output.n112 8.92171
R21484 output output.n141 8.15037
R21485 output.n43 output.n15 8.14595
R21486 output.n74 output.n46 8.14595
R21487 output.n106 output.n78 8.14595
R21488 output.n138 output.n110 8.14595
R21489 output.n45 output.n15 5.81868
R21490 output.n76 output.n46 5.81868
R21491 output.n108 output.n78 5.81868
R21492 output.n140 output.n110 5.81868
R21493 output.n43 output.n42 5.04292
R21494 output.n74 output.n73 5.04292
R21495 output.n106 output.n105 5.04292
R21496 output.n138 output.n137 5.04292
R21497 output.n28 output.n24 4.38594
R21498 output.n59 output.n55 4.38594
R21499 output.n91 output.n87 4.38594
R21500 output.n123 output.n119 4.38594
R21501 output.n39 output.n17 4.26717
R21502 output.n70 output.n48 4.26717
R21503 output.n102 output.n80 4.26717
R21504 output.n134 output.n112 4.26717
R21505 output.n0 output.t9 3.9605
R21506 output.n0 output.t13 3.9605
R21507 output.n2 output.t16 3.9605
R21508 output.n2 output.t5 3.9605
R21509 output.n4 output.t6 3.9605
R21510 output.n4 output.t11 3.9605
R21511 output.n6 output.t15 3.9605
R21512 output.n6 output.t7 3.9605
R21513 output.n8 output.t10 3.9605
R21514 output.n8 output.t8 3.9605
R21515 output.n10 output.t14 3.9605
R21516 output.n10 output.t17 3.9605
R21517 output.n12 output.t18 3.9605
R21518 output.n12 output.t12 3.9605
R21519 output.n38 output.n19 3.49141
R21520 output.n69 output.n50 3.49141
R21521 output.n101 output.n82 3.49141
R21522 output.n133 output.n114 3.49141
R21523 output.n35 output.n34 2.71565
R21524 output.n66 output.n65 2.71565
R21525 output.n98 output.n97 2.71565
R21526 output.n130 output.n129 2.71565
R21527 output.n31 output.n21 1.93989
R21528 output.n62 output.n52 1.93989
R21529 output.n94 output.n84 1.93989
R21530 output.n126 output.n116 1.93989
R21531 output.n30 output.n23 1.16414
R21532 output.n61 output.n54 1.16414
R21533 output.n93 output.n86 1.16414
R21534 output.n125 output.n118 1.16414
R21535 output.n141 output.n109 0.962709
R21536 output.n109 output.n77 0.962709
R21537 output.n27 output.n26 0.388379
R21538 output.n58 output.n57 0.388379
R21539 output.n90 output.n89 0.388379
R21540 output.n122 output.n121 0.388379
R21541 output.n14 output.n13 0.387128
R21542 output.n13 output.n11 0.387128
R21543 output.n11 output.n9 0.387128
R21544 output.n9 output.n7 0.387128
R21545 output.n7 output.n5 0.387128
R21546 output.n5 output.n3 0.387128
R21547 output.n3 output.n1 0.387128
R21548 output.n44 output.n16 0.155672
R21549 output.n37 output.n16 0.155672
R21550 output.n37 output.n36 0.155672
R21551 output.n36 output.n20 0.155672
R21552 output.n29 output.n20 0.155672
R21553 output.n29 output.n28 0.155672
R21554 output.n75 output.n47 0.155672
R21555 output.n68 output.n47 0.155672
R21556 output.n68 output.n67 0.155672
R21557 output.n67 output.n51 0.155672
R21558 output.n60 output.n51 0.155672
R21559 output.n60 output.n59 0.155672
R21560 output.n107 output.n79 0.155672
R21561 output.n100 output.n79 0.155672
R21562 output.n100 output.n99 0.155672
R21563 output.n99 output.n83 0.155672
R21564 output.n92 output.n83 0.155672
R21565 output.n92 output.n91 0.155672
R21566 output.n139 output.n111 0.155672
R21567 output.n132 output.n111 0.155672
R21568 output.n132 output.n131 0.155672
R21569 output.n131 output.n115 0.155672
R21570 output.n124 output.n115 0.155672
R21571 output.n124 output.n123 0.155672
R21572 output output.n14 0.126227
R21573 minus.n76 minus.t28 250.337
R21574 minus.n15 minus.t20 250.337
R21575 minus.n126 minus.t1 243.255
R21576 minus.n120 minus.t8 231.093
R21577 minus.n59 minus.t10 231.093
R21578 minus.n125 minus.n123 224.169
R21579 minus.n125 minus.n124 223.454
R21580 minus.n62 minus.t12 187.445
R21581 minus.n113 minus.t18 187.445
R21582 minus.n107 minus.t25 187.445
R21583 minus.n66 minus.t22 187.445
R21584 minus.n68 minus.t19 187.445
R21585 minus.n95 minus.t7 187.445
R21586 minus.n89 minus.t6 187.445
R21587 minus.n72 minus.t16 187.445
R21588 minus.n74 minus.t15 187.445
R21589 minus.n77 minus.t23 187.445
R21590 minus.n16 minus.t14 187.445
R21591 minus.n13 minus.t9 187.445
R21592 minus.n11 minus.t5 187.445
R21593 minus.n28 minus.t26 187.445
R21594 minus.n34 minus.t27 187.445
R21595 minus.n7 minus.t21 187.445
R21596 minus.n5 minus.t24 187.445
R21597 minus.n46 minus.t17 187.445
R21598 minus.n52 minus.t11 187.445
R21599 minus.n1 minus.t13 187.445
R21600 minus.n78 minus.n75 161.3
R21601 minus.n80 minus.n79 161.3
R21602 minus.n82 minus.n81 161.3
R21603 minus.n83 minus.n73 161.3
R21604 minus.n85 minus.n84 161.3
R21605 minus.n87 minus.n86 161.3
R21606 minus.n88 minus.n71 161.3
R21607 minus.n91 minus.n90 161.3
R21608 minus.n92 minus.n70 161.3
R21609 minus.n94 minus.n93 161.3
R21610 minus.n96 minus.n69 161.3
R21611 minus.n98 minus.n97 161.3
R21612 minus.n100 minus.n99 161.3
R21613 minus.n101 minus.n67 161.3
R21614 minus.n103 minus.n102 161.3
R21615 minus.n105 minus.n104 161.3
R21616 minus.n106 minus.n65 161.3
R21617 minus.n109 minus.n108 161.3
R21618 minus.n110 minus.n64 161.3
R21619 minus.n112 minus.n111 161.3
R21620 minus.n114 minus.n63 161.3
R21621 minus.n116 minus.n115 161.3
R21622 minus.n118 minus.n117 161.3
R21623 minus.n119 minus.n61 161.3
R21624 minus.n121 minus.n120 161.3
R21625 minus.n60 minus.n59 161.3
R21626 minus.n58 minus.n0 161.3
R21627 minus.n57 minus.n56 161.3
R21628 minus.n55 minus.n54 161.3
R21629 minus.n53 minus.n2 161.3
R21630 minus.n51 minus.n50 161.3
R21631 minus.n49 minus.n3 161.3
R21632 minus.n48 minus.n47 161.3
R21633 minus.n45 minus.n4 161.3
R21634 minus.n44 minus.n43 161.3
R21635 minus.n42 minus.n41 161.3
R21636 minus.n40 minus.n6 161.3
R21637 minus.n39 minus.n38 161.3
R21638 minus.n37 minus.n36 161.3
R21639 minus.n35 minus.n8 161.3
R21640 minus.n33 minus.n32 161.3
R21641 minus.n31 minus.n9 161.3
R21642 minus.n30 minus.n29 161.3
R21643 minus.n27 minus.n10 161.3
R21644 minus.n26 minus.n25 161.3
R21645 minus.n24 minus.n23 161.3
R21646 minus.n22 minus.n12 161.3
R21647 minus.n21 minus.n20 161.3
R21648 minus.n19 minus.n18 161.3
R21649 minus.n17 minus.n14 161.3
R21650 minus.n106 minus.n105 56.5617
R21651 minus.n97 minus.n96 56.5617
R21652 minus.n88 minus.n87 56.5617
R21653 minus.n27 minus.n26 56.5617
R21654 minus.n36 minus.n35 56.5617
R21655 minus.n45 minus.n44 56.5617
R21656 minus.n115 minus.n114 56.5617
R21657 minus.n79 minus.n78 56.5617
R21658 minus.n18 minus.n17 56.5617
R21659 minus.n54 minus.n53 56.5617
R21660 minus.n119 minus.n118 50.2647
R21661 minus.n58 minus.n57 50.2647
R21662 minus.n108 minus.n64 46.3896
R21663 minus.n84 minus.n83 46.3896
R21664 minus.n23 minus.n22 46.3896
R21665 minus.n47 minus.n3 46.3896
R21666 minus.n76 minus.n75 43.1929
R21667 minus.n15 minus.n14 43.1929
R21668 minus.n101 minus.n100 42.5146
R21669 minus.n94 minus.n70 42.5146
R21670 minus.n33 minus.n9 42.5146
R21671 minus.n40 minus.n39 42.5146
R21672 minus.n77 minus.n76 40.6041
R21673 minus.n16 minus.n15 40.6041
R21674 minus.n102 minus.n101 38.6395
R21675 minus.n90 minus.n70 38.6395
R21676 minus.n29 minus.n9 38.6395
R21677 minus.n41 minus.n40 38.6395
R21678 minus.n122 minus.n121 35.4191
R21679 minus.n112 minus.n64 34.7644
R21680 minus.n83 minus.n82 34.7644
R21681 minus.n22 minus.n21 34.7644
R21682 minus.n51 minus.n3 34.7644
R21683 minus.n114 minus.n113 21.8872
R21684 minus.n79 minus.n74 21.8872
R21685 minus.n18 minus.n13 21.8872
R21686 minus.n53 minus.n52 21.8872
R21687 minus.n105 minus.n66 19.9199
R21688 minus.n89 minus.n88 19.9199
R21689 minus.n28 minus.n27 19.9199
R21690 minus.n44 minus.n5 19.9199
R21691 minus.n124 minus.t0 19.8005
R21692 minus.n124 minus.t2 19.8005
R21693 minus.n123 minus.t4 19.8005
R21694 minus.n123 minus.t3 19.8005
R21695 minus.n97 minus.n68 17.9525
R21696 minus.n96 minus.n95 17.9525
R21697 minus.n35 minus.n34 17.9525
R21698 minus.n36 minus.n7 17.9525
R21699 minus.n107 minus.n106 15.9852
R21700 minus.n87 minus.n72 15.9852
R21701 minus.n26 minus.n11 15.9852
R21702 minus.n46 minus.n45 15.9852
R21703 minus.n115 minus.n62 14.0178
R21704 minus.n78 minus.n77 14.0178
R21705 minus.n17 minus.n16 14.0178
R21706 minus.n54 minus.n1 14.0178
R21707 minus.n122 minus.n60 12.1501
R21708 minus minus.n127 10.9162
R21709 minus.n118 minus.n62 10.575
R21710 minus.n57 minus.n1 10.575
R21711 minus.n120 minus.n119 9.49444
R21712 minus.n59 minus.n58 9.49444
R21713 minus.n108 minus.n107 8.60764
R21714 minus.n84 minus.n72 8.60764
R21715 minus.n23 minus.n11 8.60764
R21716 minus.n47 minus.n46 8.60764
R21717 minus.n100 minus.n68 6.6403
R21718 minus.n95 minus.n94 6.6403
R21719 minus.n34 minus.n33 6.6403
R21720 minus.n39 minus.n7 6.6403
R21721 minus.n127 minus.n126 4.80222
R21722 minus.n102 minus.n66 4.67295
R21723 minus.n90 minus.n89 4.67295
R21724 minus.n29 minus.n28 4.67295
R21725 minus.n41 minus.n5 4.67295
R21726 minus.n113 minus.n112 2.7056
R21727 minus.n82 minus.n74 2.7056
R21728 minus.n21 minus.n13 2.7056
R21729 minus.n52 minus.n51 2.7056
R21730 minus.n127 minus.n122 0.972091
R21731 minus.n126 minus.n125 0.716017
R21732 minus.n121 minus.n61 0.189894
R21733 minus.n117 minus.n61 0.189894
R21734 minus.n117 minus.n116 0.189894
R21735 minus.n116 minus.n63 0.189894
R21736 minus.n111 minus.n63 0.189894
R21737 minus.n111 minus.n110 0.189894
R21738 minus.n110 minus.n109 0.189894
R21739 minus.n109 minus.n65 0.189894
R21740 minus.n104 minus.n65 0.189894
R21741 minus.n104 minus.n103 0.189894
R21742 minus.n103 minus.n67 0.189894
R21743 minus.n99 minus.n67 0.189894
R21744 minus.n99 minus.n98 0.189894
R21745 minus.n98 minus.n69 0.189894
R21746 minus.n93 minus.n69 0.189894
R21747 minus.n93 minus.n92 0.189894
R21748 minus.n92 minus.n91 0.189894
R21749 minus.n91 minus.n71 0.189894
R21750 minus.n86 minus.n71 0.189894
R21751 minus.n86 minus.n85 0.189894
R21752 minus.n85 minus.n73 0.189894
R21753 minus.n81 minus.n73 0.189894
R21754 minus.n81 minus.n80 0.189894
R21755 minus.n80 minus.n75 0.189894
R21756 minus.n19 minus.n14 0.189894
R21757 minus.n20 minus.n19 0.189894
R21758 minus.n20 minus.n12 0.189894
R21759 minus.n24 minus.n12 0.189894
R21760 minus.n25 minus.n24 0.189894
R21761 minus.n25 minus.n10 0.189894
R21762 minus.n30 minus.n10 0.189894
R21763 minus.n31 minus.n30 0.189894
R21764 minus.n32 minus.n31 0.189894
R21765 minus.n32 minus.n8 0.189894
R21766 minus.n37 minus.n8 0.189894
R21767 minus.n38 minus.n37 0.189894
R21768 minus.n38 minus.n6 0.189894
R21769 minus.n42 minus.n6 0.189894
R21770 minus.n43 minus.n42 0.189894
R21771 minus.n43 minus.n4 0.189894
R21772 minus.n48 minus.n4 0.189894
R21773 minus.n49 minus.n48 0.189894
R21774 minus.n50 minus.n49 0.189894
R21775 minus.n50 minus.n2 0.189894
R21776 minus.n55 minus.n2 0.189894
R21777 minus.n56 minus.n55 0.189894
R21778 minus.n56 minus.n0 0.189894
R21779 minus.n60 minus.n0 0.189894
R21780 diffpairibias.n0 diffpairibias.t18 436.822
R21781 diffpairibias.n21 diffpairibias.t19 435.479
R21782 diffpairibias.n20 diffpairibias.t16 435.479
R21783 diffpairibias.n19 diffpairibias.t17 435.479
R21784 diffpairibias.n18 diffpairibias.t21 435.479
R21785 diffpairibias.n0 diffpairibias.t22 435.479
R21786 diffpairibias.n1 diffpairibias.t20 435.479
R21787 diffpairibias.n2 diffpairibias.t23 435.479
R21788 diffpairibias.n10 diffpairibias.t0 377.536
R21789 diffpairibias.n10 diffpairibias.t8 376.193
R21790 diffpairibias.n11 diffpairibias.t10 376.193
R21791 diffpairibias.n12 diffpairibias.t6 376.193
R21792 diffpairibias.n13 diffpairibias.t2 376.193
R21793 diffpairibias.n14 diffpairibias.t12 376.193
R21794 diffpairibias.n15 diffpairibias.t4 376.193
R21795 diffpairibias.n16 diffpairibias.t14 376.193
R21796 diffpairibias.n3 diffpairibias.t1 113.368
R21797 diffpairibias.n3 diffpairibias.t9 112.698
R21798 diffpairibias.n4 diffpairibias.t11 112.698
R21799 diffpairibias.n5 diffpairibias.t7 112.698
R21800 diffpairibias.n6 diffpairibias.t3 112.698
R21801 diffpairibias.n7 diffpairibias.t13 112.698
R21802 diffpairibias.n8 diffpairibias.t5 112.698
R21803 diffpairibias.n9 diffpairibias.t15 112.698
R21804 diffpairibias.n17 diffpairibias.n16 4.77242
R21805 diffpairibias.n17 diffpairibias.n9 4.30807
R21806 diffpairibias.n18 diffpairibias.n17 4.13945
R21807 diffpairibias.n16 diffpairibias.n15 1.34352
R21808 diffpairibias.n15 diffpairibias.n14 1.34352
R21809 diffpairibias.n14 diffpairibias.n13 1.34352
R21810 diffpairibias.n13 diffpairibias.n12 1.34352
R21811 diffpairibias.n12 diffpairibias.n11 1.34352
R21812 diffpairibias.n11 diffpairibias.n10 1.34352
R21813 diffpairibias.n2 diffpairibias.n1 1.34352
R21814 diffpairibias.n1 diffpairibias.n0 1.34352
R21815 diffpairibias.n19 diffpairibias.n18 1.34352
R21816 diffpairibias.n20 diffpairibias.n19 1.34352
R21817 diffpairibias.n21 diffpairibias.n20 1.34352
R21818 diffpairibias.n22 diffpairibias.n21 0.862419
R21819 diffpairibias diffpairibias.n22 0.684875
R21820 diffpairibias.n9 diffpairibias.n8 0.672012
R21821 diffpairibias.n8 diffpairibias.n7 0.672012
R21822 diffpairibias.n7 diffpairibias.n6 0.672012
R21823 diffpairibias.n6 diffpairibias.n5 0.672012
R21824 diffpairibias.n5 diffpairibias.n4 0.672012
R21825 diffpairibias.n4 diffpairibias.n3 0.672012
R21826 diffpairibias.n22 diffpairibias.n2 0.190907
C0 CSoutput outputibias 0.032386f
C1 vdd CSoutput 0.116309p
C2 commonsourceibias output 0.006808f
C3 minus diffpairibias 5.39e-19
C4 CSoutput minus 2.25384f
C5 vdd plus 0.088406f
C6 plus diffpairibias 4.4e-19
C7 commonsourceibias outputibias 0.003832f
C8 vdd commonsourceibias 0.004218f
C9 CSoutput plus 0.874948f
C10 commonsourceibias diffpairibias 0.052851f
C11 CSoutput commonsourceibias 29.0223f
C12 minus plus 9.674179f
C13 minus commonsourceibias 0.515369f
C14 plus commonsourceibias 0.498793f
C15 output outputibias 2.34152f
C16 vdd output 7.23429f
C17 CSoutput output 6.13571f
C18 diffpairibias gnd 48.95304f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.118072p
C22 plus gnd 37.5393f
C23 minus gnd 28.66661f
C24 CSoutput gnd 88.29008f
C25 vdd gnd 0.408085p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031832f
C74 minus.t13 gnd 0.535246f
C75 minus.n1 gnd 0.216477f
C76 minus.n2 gnd 0.031832f
C77 minus.t11 gnd 0.535246f
C78 minus.n3 gnd 0.027201f
C79 minus.n4 gnd 0.031832f
C80 minus.t17 gnd 0.535246f
C81 minus.t24 gnd 0.535246f
C82 minus.n5 gnd 0.216477f
C83 minus.n6 gnd 0.031832f
C84 minus.t21 gnd 0.535246f
C85 minus.n7 gnd 0.216477f
C86 minus.n8 gnd 0.031832f
C87 minus.t27 gnd 0.535246f
C88 minus.n9 gnd 0.025872f
C89 minus.n10 gnd 0.031832f
C90 minus.t26 gnd 0.535246f
C91 minus.t5 gnd 0.535246f
C92 minus.n11 gnd 0.216477f
C93 minus.n12 gnd 0.031832f
C94 minus.t9 gnd 0.535246f
C95 minus.n13 gnd 0.216477f
C96 minus.n14 gnd 0.135091f
C97 minus.t14 gnd 0.535246f
C98 minus.t20 gnd 0.59877f
C99 minus.n15 gnd 0.253084f
C100 minus.n16 gnd 0.247907f
C101 minus.n17 gnd 0.040787f
C102 minus.n18 gnd 0.036021f
C103 minus.n19 gnd 0.031832f
C104 minus.n20 gnd 0.031832f
C105 minus.n21 gnd 0.038039f
C106 minus.n22 gnd 0.027201f
C107 minus.n23 gnd 0.041457f
C108 minus.n24 gnd 0.031832f
C109 minus.n25 gnd 0.031832f
C110 minus.n26 gnd 0.039596f
C111 minus.n27 gnd 0.037213f
C112 minus.n28 gnd 0.216477f
C113 minus.n29 gnd 0.039874f
C114 minus.n30 gnd 0.031832f
C115 minus.n31 gnd 0.031832f
C116 minus.n32 gnd 0.031832f
C117 minus.n33 gnd 0.04095f
C118 minus.n34 gnd 0.216477f
C119 minus.n35 gnd 0.038404f
C120 minus.n36 gnd 0.038404f
C121 minus.n37 gnd 0.031832f
C122 minus.n38 gnd 0.031832f
C123 minus.n39 gnd 0.04095f
C124 minus.n40 gnd 0.025872f
C125 minus.n41 gnd 0.039874f
C126 minus.n42 gnd 0.031832f
C127 minus.n43 gnd 0.031832f
C128 minus.n44 gnd 0.037213f
C129 minus.n45 gnd 0.039596f
C130 minus.n46 gnd 0.216477f
C131 minus.n47 gnd 0.041457f
C132 minus.n48 gnd 0.031832f
C133 minus.n49 gnd 0.031832f
C134 minus.n50 gnd 0.031832f
C135 minus.n51 gnd 0.038039f
C136 minus.n52 gnd 0.216477f
C137 minus.n53 gnd 0.036021f
C138 minus.n54 gnd 0.040787f
C139 minus.n55 gnd 0.031832f
C140 minus.n56 gnd 0.031832f
C141 minus.n57 gnd 0.041526f
C142 minus.n58 gnd 0.011569f
C143 minus.t10 gnd 0.578869f
C144 minus.n59 gnd 0.250644f
C145 minus.n60 gnd 0.372897f
C146 minus.n61 gnd 0.031832f
C147 minus.t8 gnd 0.578869f
C148 minus.t12 gnd 0.535246f
C149 minus.n62 gnd 0.216477f
C150 minus.n63 gnd 0.031832f
C151 minus.t18 gnd 0.535246f
C152 minus.n64 gnd 0.027201f
C153 minus.n65 gnd 0.031832f
C154 minus.t25 gnd 0.535246f
C155 minus.t22 gnd 0.535246f
C156 minus.n66 gnd 0.216477f
C157 minus.n67 gnd 0.031832f
C158 minus.t19 gnd 0.535246f
C159 minus.n68 gnd 0.216477f
C160 minus.n69 gnd 0.031832f
C161 minus.t7 gnd 0.535246f
C162 minus.n70 gnd 0.025872f
C163 minus.n71 gnd 0.031832f
C164 minus.t6 gnd 0.535246f
C165 minus.t16 gnd 0.535246f
C166 minus.n72 gnd 0.216477f
C167 minus.n73 gnd 0.031832f
C168 minus.t15 gnd 0.535246f
C169 minus.n74 gnd 0.216477f
C170 minus.n75 gnd 0.135091f
C171 minus.t23 gnd 0.535246f
C172 minus.t28 gnd 0.59877f
C173 minus.n76 gnd 0.253084f
C174 minus.n77 gnd 0.247907f
C175 minus.n78 gnd 0.040787f
C176 minus.n79 gnd 0.036021f
C177 minus.n80 gnd 0.031832f
C178 minus.n81 gnd 0.031832f
C179 minus.n82 gnd 0.038039f
C180 minus.n83 gnd 0.027201f
C181 minus.n84 gnd 0.041457f
C182 minus.n85 gnd 0.031832f
C183 minus.n86 gnd 0.031832f
C184 minus.n87 gnd 0.039596f
C185 minus.n88 gnd 0.037213f
C186 minus.n89 gnd 0.216477f
C187 minus.n90 gnd 0.039874f
C188 minus.n91 gnd 0.031832f
C189 minus.n92 gnd 0.031832f
C190 minus.n93 gnd 0.031832f
C191 minus.n94 gnd 0.04095f
C192 minus.n95 gnd 0.216477f
C193 minus.n96 gnd 0.038404f
C194 minus.n97 gnd 0.038404f
C195 minus.n98 gnd 0.031832f
C196 minus.n99 gnd 0.031832f
C197 minus.n100 gnd 0.04095f
C198 minus.n101 gnd 0.025872f
C199 minus.n102 gnd 0.039874f
C200 minus.n103 gnd 0.031832f
C201 minus.n104 gnd 0.031832f
C202 minus.n105 gnd 0.037213f
C203 minus.n106 gnd 0.039596f
C204 minus.n107 gnd 0.216477f
C205 minus.n108 gnd 0.041457f
C206 minus.n109 gnd 0.031832f
C207 minus.n110 gnd 0.031832f
C208 minus.n111 gnd 0.031832f
C209 minus.n112 gnd 0.038039f
C210 minus.n113 gnd 0.216477f
C211 minus.n114 gnd 0.036021f
C212 minus.n115 gnd 0.040787f
C213 minus.n116 gnd 0.031832f
C214 minus.n117 gnd 0.031832f
C215 minus.n118 gnd 0.041526f
C216 minus.n119 gnd 0.011569f
C217 minus.n120 gnd 0.250644f
C218 minus.n121 gnd 1.16121f
C219 minus.n122 gnd 1.70573f
C220 minus.t4 gnd 0.009813f
C221 minus.t3 gnd 0.009813f
C222 minus.n123 gnd 0.032267f
C223 minus.t0 gnd 0.009813f
C224 minus.t2 gnd 0.009813f
C225 minus.n124 gnd 0.031825f
C226 minus.n125 gnd 0.271609f
C227 minus.t1 gnd 0.054617f
C228 minus.n126 gnd 0.148215f
C229 minus.n127 gnd 1.6183f
C230 output.t19 gnd 0.464308f
C231 output.t9 gnd 0.044422f
C232 output.t13 gnd 0.044422f
C233 output.n0 gnd 0.364624f
C234 output.n1 gnd 0.614102f
C235 output.t16 gnd 0.044422f
C236 output.t5 gnd 0.044422f
C237 output.n2 gnd 0.364624f
C238 output.n3 gnd 0.350265f
C239 output.t6 gnd 0.044422f
C240 output.t11 gnd 0.044422f
C241 output.n4 gnd 0.364624f
C242 output.n5 gnd 0.350265f
C243 output.t15 gnd 0.044422f
C244 output.t7 gnd 0.044422f
C245 output.n6 gnd 0.364624f
C246 output.n7 gnd 0.350265f
C247 output.t10 gnd 0.044422f
C248 output.t8 gnd 0.044422f
C249 output.n8 gnd 0.364624f
C250 output.n9 gnd 0.350265f
C251 output.t14 gnd 0.044422f
C252 output.t17 gnd 0.044422f
C253 output.n10 gnd 0.364624f
C254 output.n11 gnd 0.350265f
C255 output.t18 gnd 0.044422f
C256 output.t12 gnd 0.044422f
C257 output.n12 gnd 0.364624f
C258 output.n13 gnd 0.350265f
C259 output.t4 gnd 0.462979f
C260 output.n14 gnd 0.28994f
C261 output.n15 gnd 0.015803f
C262 output.n16 gnd 0.011243f
C263 output.n17 gnd 0.006041f
C264 output.n18 gnd 0.01428f
C265 output.n19 gnd 0.006397f
C266 output.n20 gnd 0.011243f
C267 output.n21 gnd 0.006041f
C268 output.n22 gnd 0.01428f
C269 output.n23 gnd 0.006397f
C270 output.n24 gnd 0.048111f
C271 output.t3 gnd 0.023274f
C272 output.n25 gnd 0.01071f
C273 output.n26 gnd 0.008435f
C274 output.n27 gnd 0.006041f
C275 output.n28 gnd 0.267512f
C276 output.n29 gnd 0.011243f
C277 output.n30 gnd 0.006041f
C278 output.n31 gnd 0.006397f
C279 output.n32 gnd 0.01428f
C280 output.n33 gnd 0.01428f
C281 output.n34 gnd 0.006397f
C282 output.n35 gnd 0.006041f
C283 output.n36 gnd 0.011243f
C284 output.n37 gnd 0.011243f
C285 output.n38 gnd 0.006041f
C286 output.n39 gnd 0.006397f
C287 output.n40 gnd 0.01428f
C288 output.n41 gnd 0.030913f
C289 output.n42 gnd 0.006397f
C290 output.n43 gnd 0.006041f
C291 output.n44 gnd 0.025987f
C292 output.n45 gnd 0.097665f
C293 output.n46 gnd 0.015803f
C294 output.n47 gnd 0.011243f
C295 output.n48 gnd 0.006041f
C296 output.n49 gnd 0.01428f
C297 output.n50 gnd 0.006397f
C298 output.n51 gnd 0.011243f
C299 output.n52 gnd 0.006041f
C300 output.n53 gnd 0.01428f
C301 output.n54 gnd 0.006397f
C302 output.n55 gnd 0.048111f
C303 output.t2 gnd 0.023274f
C304 output.n56 gnd 0.01071f
C305 output.n57 gnd 0.008435f
C306 output.n58 gnd 0.006041f
C307 output.n59 gnd 0.267512f
C308 output.n60 gnd 0.011243f
C309 output.n61 gnd 0.006041f
C310 output.n62 gnd 0.006397f
C311 output.n63 gnd 0.01428f
C312 output.n64 gnd 0.01428f
C313 output.n65 gnd 0.006397f
C314 output.n66 gnd 0.006041f
C315 output.n67 gnd 0.011243f
C316 output.n68 gnd 0.011243f
C317 output.n69 gnd 0.006041f
C318 output.n70 gnd 0.006397f
C319 output.n71 gnd 0.01428f
C320 output.n72 gnd 0.030913f
C321 output.n73 gnd 0.006397f
C322 output.n74 gnd 0.006041f
C323 output.n75 gnd 0.025987f
C324 output.n76 gnd 0.09306f
C325 output.n77 gnd 1.65264f
C326 output.n78 gnd 0.015803f
C327 output.n79 gnd 0.011243f
C328 output.n80 gnd 0.006041f
C329 output.n81 gnd 0.01428f
C330 output.n82 gnd 0.006397f
C331 output.n83 gnd 0.011243f
C332 output.n84 gnd 0.006041f
C333 output.n85 gnd 0.01428f
C334 output.n86 gnd 0.006397f
C335 output.n87 gnd 0.048111f
C336 output.t1 gnd 0.023274f
C337 output.n88 gnd 0.01071f
C338 output.n89 gnd 0.008435f
C339 output.n90 gnd 0.006041f
C340 output.n91 gnd 0.267512f
C341 output.n92 gnd 0.011243f
C342 output.n93 gnd 0.006041f
C343 output.n94 gnd 0.006397f
C344 output.n95 gnd 0.01428f
C345 output.n96 gnd 0.01428f
C346 output.n97 gnd 0.006397f
C347 output.n98 gnd 0.006041f
C348 output.n99 gnd 0.011243f
C349 output.n100 gnd 0.011243f
C350 output.n101 gnd 0.006041f
C351 output.n102 gnd 0.006397f
C352 output.n103 gnd 0.01428f
C353 output.n104 gnd 0.030913f
C354 output.n105 gnd 0.006397f
C355 output.n106 gnd 0.006041f
C356 output.n107 gnd 0.025987f
C357 output.n108 gnd 0.09306f
C358 output.n109 gnd 0.713089f
C359 output.n110 gnd 0.015803f
C360 output.n111 gnd 0.011243f
C361 output.n112 gnd 0.006041f
C362 output.n113 gnd 0.01428f
C363 output.n114 gnd 0.006397f
C364 output.n115 gnd 0.011243f
C365 output.n116 gnd 0.006041f
C366 output.n117 gnd 0.01428f
C367 output.n118 gnd 0.006397f
C368 output.n119 gnd 0.048111f
C369 output.t0 gnd 0.023274f
C370 output.n120 gnd 0.01071f
C371 output.n121 gnd 0.008435f
C372 output.n122 gnd 0.006041f
C373 output.n123 gnd 0.267512f
C374 output.n124 gnd 0.011243f
C375 output.n125 gnd 0.006041f
C376 output.n126 gnd 0.006397f
C377 output.n127 gnd 0.01428f
C378 output.n128 gnd 0.01428f
C379 output.n129 gnd 0.006397f
C380 output.n130 gnd 0.006041f
C381 output.n131 gnd 0.011243f
C382 output.n132 gnd 0.011243f
C383 output.n133 gnd 0.006041f
C384 output.n134 gnd 0.006397f
C385 output.n135 gnd 0.01428f
C386 output.n136 gnd 0.030913f
C387 output.n137 gnd 0.006397f
C388 output.n138 gnd 0.006041f
C389 output.n139 gnd 0.025987f
C390 output.n140 gnd 0.09306f
C391 output.n141 gnd 1.67353f
C392 outputibias.t9 gnd 0.11477f
C393 outputibias.t8 gnd 0.115567f
C394 outputibias.n0 gnd 0.130108f
C395 outputibias.n1 gnd 0.001372f
C396 outputibias.n2 gnd 9.76e-19
C397 outputibias.n3 gnd 5.24e-19
C398 outputibias.n4 gnd 0.001239f
C399 outputibias.n5 gnd 5.55e-19
C400 outputibias.n6 gnd 9.76e-19
C401 outputibias.n7 gnd 5.24e-19
C402 outputibias.n8 gnd 0.001239f
C403 outputibias.n9 gnd 5.55e-19
C404 outputibias.n10 gnd 0.004176f
C405 outputibias.t5 gnd 0.00202f
C406 outputibias.n11 gnd 9.3e-19
C407 outputibias.n12 gnd 7.32e-19
C408 outputibias.n13 gnd 5.24e-19
C409 outputibias.n14 gnd 0.02322f
C410 outputibias.n15 gnd 9.76e-19
C411 outputibias.n16 gnd 5.24e-19
C412 outputibias.n17 gnd 5.55e-19
C413 outputibias.n18 gnd 0.001239f
C414 outputibias.n19 gnd 0.001239f
C415 outputibias.n20 gnd 5.55e-19
C416 outputibias.n21 gnd 5.24e-19
C417 outputibias.n22 gnd 9.76e-19
C418 outputibias.n23 gnd 9.76e-19
C419 outputibias.n24 gnd 5.24e-19
C420 outputibias.n25 gnd 5.55e-19
C421 outputibias.n26 gnd 0.001239f
C422 outputibias.n27 gnd 0.002683f
C423 outputibias.n28 gnd 5.55e-19
C424 outputibias.n29 gnd 5.24e-19
C425 outputibias.n30 gnd 0.002256f
C426 outputibias.n31 gnd 0.005781f
C427 outputibias.n32 gnd 0.001372f
C428 outputibias.n33 gnd 9.76e-19
C429 outputibias.n34 gnd 5.24e-19
C430 outputibias.n35 gnd 0.001239f
C431 outputibias.n36 gnd 5.55e-19
C432 outputibias.n37 gnd 9.76e-19
C433 outputibias.n38 gnd 5.24e-19
C434 outputibias.n39 gnd 0.001239f
C435 outputibias.n40 gnd 5.55e-19
C436 outputibias.n41 gnd 0.004176f
C437 outputibias.t7 gnd 0.00202f
C438 outputibias.n42 gnd 9.3e-19
C439 outputibias.n43 gnd 7.32e-19
C440 outputibias.n44 gnd 5.24e-19
C441 outputibias.n45 gnd 0.02322f
C442 outputibias.n46 gnd 9.76e-19
C443 outputibias.n47 gnd 5.24e-19
C444 outputibias.n48 gnd 5.55e-19
C445 outputibias.n49 gnd 0.001239f
C446 outputibias.n50 gnd 0.001239f
C447 outputibias.n51 gnd 5.55e-19
C448 outputibias.n52 gnd 5.24e-19
C449 outputibias.n53 gnd 9.76e-19
C450 outputibias.n54 gnd 9.76e-19
C451 outputibias.n55 gnd 5.24e-19
C452 outputibias.n56 gnd 5.55e-19
C453 outputibias.n57 gnd 0.001239f
C454 outputibias.n58 gnd 0.002683f
C455 outputibias.n59 gnd 5.55e-19
C456 outputibias.n60 gnd 5.24e-19
C457 outputibias.n61 gnd 0.002256f
C458 outputibias.n62 gnd 0.005197f
C459 outputibias.n63 gnd 0.121892f
C460 outputibias.n64 gnd 0.001372f
C461 outputibias.n65 gnd 9.76e-19
C462 outputibias.n66 gnd 5.24e-19
C463 outputibias.n67 gnd 0.001239f
C464 outputibias.n68 gnd 5.55e-19
C465 outputibias.n69 gnd 9.76e-19
C466 outputibias.n70 gnd 5.24e-19
C467 outputibias.n71 gnd 0.001239f
C468 outputibias.n72 gnd 5.55e-19
C469 outputibias.n73 gnd 0.004176f
C470 outputibias.t1 gnd 0.00202f
C471 outputibias.n74 gnd 9.3e-19
C472 outputibias.n75 gnd 7.32e-19
C473 outputibias.n76 gnd 5.24e-19
C474 outputibias.n77 gnd 0.02322f
C475 outputibias.n78 gnd 9.76e-19
C476 outputibias.n79 gnd 5.24e-19
C477 outputibias.n80 gnd 5.55e-19
C478 outputibias.n81 gnd 0.001239f
C479 outputibias.n82 gnd 0.001239f
C480 outputibias.n83 gnd 5.55e-19
C481 outputibias.n84 gnd 5.24e-19
C482 outputibias.n85 gnd 9.76e-19
C483 outputibias.n86 gnd 9.76e-19
C484 outputibias.n87 gnd 5.24e-19
C485 outputibias.n88 gnd 5.55e-19
C486 outputibias.n89 gnd 0.001239f
C487 outputibias.n90 gnd 0.002683f
C488 outputibias.n91 gnd 5.55e-19
C489 outputibias.n92 gnd 5.24e-19
C490 outputibias.n93 gnd 0.002256f
C491 outputibias.n94 gnd 0.005197f
C492 outputibias.n95 gnd 0.064513f
C493 outputibias.n96 gnd 0.001372f
C494 outputibias.n97 gnd 9.76e-19
C495 outputibias.n98 gnd 5.24e-19
C496 outputibias.n99 gnd 0.001239f
C497 outputibias.n100 gnd 5.55e-19
C498 outputibias.n101 gnd 9.76e-19
C499 outputibias.n102 gnd 5.24e-19
C500 outputibias.n103 gnd 0.001239f
C501 outputibias.n104 gnd 5.55e-19
C502 outputibias.n105 gnd 0.004176f
C503 outputibias.t3 gnd 0.00202f
C504 outputibias.n106 gnd 9.3e-19
C505 outputibias.n107 gnd 7.32e-19
C506 outputibias.n108 gnd 5.24e-19
C507 outputibias.n109 gnd 0.02322f
C508 outputibias.n110 gnd 9.76e-19
C509 outputibias.n111 gnd 5.24e-19
C510 outputibias.n112 gnd 5.55e-19
C511 outputibias.n113 gnd 0.001239f
C512 outputibias.n114 gnd 0.001239f
C513 outputibias.n115 gnd 5.55e-19
C514 outputibias.n116 gnd 5.24e-19
C515 outputibias.n117 gnd 9.76e-19
C516 outputibias.n118 gnd 9.76e-19
C517 outputibias.n119 gnd 5.24e-19
C518 outputibias.n120 gnd 5.55e-19
C519 outputibias.n121 gnd 0.001239f
C520 outputibias.n122 gnd 0.002683f
C521 outputibias.n123 gnd 5.55e-19
C522 outputibias.n124 gnd 5.24e-19
C523 outputibias.n125 gnd 0.002256f
C524 outputibias.n126 gnd 0.005197f
C525 outputibias.n127 gnd 0.084814f
C526 outputibias.t2 gnd 0.108319f
C527 outputibias.t0 gnd 0.108319f
C528 outputibias.t6 gnd 0.108319f
C529 outputibias.t4 gnd 0.109238f
C530 outputibias.n128 gnd 0.134674f
C531 outputibias.n129 gnd 0.07244f
C532 outputibias.n130 gnd 0.079818f
C533 outputibias.n131 gnd 0.164901f
C534 outputibias.t11 gnd 0.11477f
C535 outputibias.n132 gnd 0.067481f
C536 outputibias.t10 gnd 0.11477f
C537 outputibias.n133 gnd 0.065115f
C538 outputibias.n134 gnd 0.029159f
C539 a_n3106_n452.t10 gnd 0.10001f
C540 a_n3106_n452.t21 gnd 1.03942f
C541 a_n3106_n452.n0 gnd 0.392946f
C542 a_n3106_n452.t31 gnd 1.29145f
C543 a_n3106_n452.n1 gnd 1.22854f
C544 a_n3106_n452.t37 gnd 1.03942f
C545 a_n3106_n452.n2 gnd 0.392946f
C546 a_n3106_n452.t44 gnd 0.10001f
C547 a_n3106_n452.t34 gnd 0.10001f
C548 a_n3106_n452.n3 gnd 0.816794f
C549 a_n3106_n452.n4 gnd 0.411618f
C550 a_n3106_n452.t48 gnd 0.10001f
C551 a_n3106_n452.t2 gnd 0.10001f
C552 a_n3106_n452.n5 gnd 0.816794f
C553 a_n3106_n452.n6 gnd 0.411618f
C554 a_n3106_n452.t30 gnd 0.10001f
C555 a_n3106_n452.t47 gnd 0.10001f
C556 a_n3106_n452.n7 gnd 0.816794f
C557 a_n3106_n452.n8 gnd 0.411618f
C558 a_n3106_n452.t35 gnd 0.10001f
C559 a_n3106_n452.t38 gnd 0.10001f
C560 a_n3106_n452.n9 gnd 0.816794f
C561 a_n3106_n452.n10 gnd 0.411618f
C562 a_n3106_n452.t53 gnd 0.10001f
C563 a_n3106_n452.t1 gnd 0.10001f
C564 a_n3106_n452.n11 gnd 0.816794f
C565 a_n3106_n452.n12 gnd 0.411618f
C566 a_n3106_n452.t46 gnd 1.03942f
C567 a_n3106_n452.n13 gnd 0.972974f
C568 a_n3106_n452.t40 gnd 1.29145f
C569 a_n3106_n452.n14 gnd 0.909591f
C570 a_n3106_n452.t32 gnd 1.29145f
C571 a_n3106_n452.n15 gnd 0.909591f
C572 a_n3106_n452.t39 gnd 1.29145f
C573 a_n3106_n452.n16 gnd 0.909591f
C574 a_n3106_n452.t28 gnd 1.29145f
C575 a_n3106_n452.n17 gnd 0.909591f
C576 a_n3106_n452.t0 gnd 1.29145f
C577 a_n3106_n452.n18 gnd 0.909591f
C578 a_n3106_n452.t43 gnd 1.29145f
C579 a_n3106_n452.n19 gnd 0.909591f
C580 a_n3106_n452.t41 gnd 1.29145f
C581 a_n3106_n452.n20 gnd 0.789472f
C582 a_n3106_n452.n21 gnd 0.948419f
C583 a_n3106_n452.t12 gnd 1.03941f
C584 a_n3106_n452.n22 gnd 0.645631f
C585 a_n3106_n452.t9 gnd 0.10001f
C586 a_n3106_n452.t26 gnd 0.10001f
C587 a_n3106_n452.n23 gnd 0.816793f
C588 a_n3106_n452.n24 gnd 0.41162f
C589 a_n3106_n452.t20 gnd 0.10001f
C590 a_n3106_n452.t24 gnd 0.10001f
C591 a_n3106_n452.n25 gnd 0.816793f
C592 a_n3106_n452.n26 gnd 0.41162f
C593 a_n3106_n452.t25 gnd 0.10001f
C594 a_n3106_n452.t13 gnd 0.10001f
C595 a_n3106_n452.n27 gnd 0.816793f
C596 a_n3106_n452.n28 gnd 0.41162f
C597 a_n3106_n452.t14 gnd 0.10001f
C598 a_n3106_n452.t5 gnd 0.10001f
C599 a_n3106_n452.n29 gnd 0.816793f
C600 a_n3106_n452.n30 gnd 0.41162f
C601 a_n3106_n452.t7 gnd 0.10001f
C602 a_n3106_n452.t23 gnd 0.10001f
C603 a_n3106_n452.n31 gnd 0.816793f
C604 a_n3106_n452.n32 gnd 0.41162f
C605 a_n3106_n452.t18 gnd 1.03941f
C606 a_n3106_n452.n33 gnd 0.39295f
C607 a_n3106_n452.t29 gnd 1.03941f
C608 a_n3106_n452.n34 gnd 0.39295f
C609 a_n3106_n452.t51 gnd 0.10001f
C610 a_n3106_n452.t45 gnd 0.10001f
C611 a_n3106_n452.n35 gnd 0.816793f
C612 a_n3106_n452.n36 gnd 0.41162f
C613 a_n3106_n452.t49 gnd 0.10001f
C614 a_n3106_n452.t55 gnd 0.10001f
C615 a_n3106_n452.n37 gnd 0.816793f
C616 a_n3106_n452.n38 gnd 0.41162f
C617 a_n3106_n452.t3 gnd 0.10001f
C618 a_n3106_n452.t36 gnd 0.10001f
C619 a_n3106_n452.n39 gnd 0.816793f
C620 a_n3106_n452.n40 gnd 0.41162f
C621 a_n3106_n452.t33 gnd 0.10001f
C622 a_n3106_n452.t42 gnd 0.10001f
C623 a_n3106_n452.n41 gnd 0.816793f
C624 a_n3106_n452.n42 gnd 0.41162f
C625 a_n3106_n452.t54 gnd 0.10001f
C626 a_n3106_n452.t52 gnd 0.10001f
C627 a_n3106_n452.n43 gnd 0.816793f
C628 a_n3106_n452.n44 gnd 0.41162f
C629 a_n3106_n452.t50 gnd 1.03941f
C630 a_n3106_n452.n45 gnd 0.645631f
C631 a_n3106_n452.n46 gnd 1.05146f
C632 a_n3106_n452.t8 gnd 1.03941f
C633 a_n3106_n452.n47 gnd 0.972978f
C634 a_n3106_n452.t6 gnd 0.10001f
C635 a_n3106_n452.t4 gnd 0.10001f
C636 a_n3106_n452.n48 gnd 0.816794f
C637 a_n3106_n452.n49 gnd 0.411618f
C638 a_n3106_n452.t17 gnd 0.10001f
C639 a_n3106_n452.t22 gnd 0.10001f
C640 a_n3106_n452.n50 gnd 0.816794f
C641 a_n3106_n452.n51 gnd 0.411618f
C642 a_n3106_n452.t15 gnd 0.10001f
C643 a_n3106_n452.t19 gnd 0.10001f
C644 a_n3106_n452.n52 gnd 0.816794f
C645 a_n3106_n452.n53 gnd 0.411618f
C646 a_n3106_n452.t11 gnd 0.10001f
C647 a_n3106_n452.t16 gnd 0.10001f
C648 a_n3106_n452.n54 gnd 0.816794f
C649 a_n3106_n452.n55 gnd 0.411618f
C650 a_n3106_n452.n56 gnd 0.411617f
C651 a_n3106_n452.n57 gnd 0.816796f
C652 a_n3106_n452.t27 gnd 0.10001f
C653 plus.n0 gnd 0.023652f
C654 plus.t20 gnd 0.430126f
C655 plus.t23 gnd 0.397712f
C656 plus.n1 gnd 0.160852f
C657 plus.n2 gnd 0.023652f
C658 plus.t6 gnd 0.397712f
C659 plus.n3 gnd 0.020211f
C660 plus.n4 gnd 0.023652f
C661 plus.t12 gnd 0.397712f
C662 plus.t8 gnd 0.397712f
C663 plus.n5 gnd 0.160852f
C664 plus.n6 gnd 0.023652f
C665 plus.t7 gnd 0.397712f
C666 plus.n7 gnd 0.160852f
C667 plus.n8 gnd 0.023652f
C668 plus.t19 gnd 0.397712f
C669 plus.n9 gnd 0.019224f
C670 plus.n10 gnd 0.023652f
C671 plus.t18 gnd 0.397712f
C672 plus.t27 gnd 0.397712f
C673 plus.n11 gnd 0.160852f
C674 plus.n12 gnd 0.023652f
C675 plus.t25 gnd 0.397712f
C676 plus.n13 gnd 0.160852f
C677 plus.n14 gnd 0.100378f
C678 plus.t9 gnd 0.397712f
C679 plus.t14 gnd 0.444913f
C680 plus.n15 gnd 0.188053f
C681 plus.n16 gnd 0.184206f
C682 plus.n17 gnd 0.030307f
C683 plus.n18 gnd 0.026765f
C684 plus.n19 gnd 0.023652f
C685 plus.n20 gnd 0.023652f
C686 plus.n21 gnd 0.028265f
C687 plus.n22 gnd 0.020211f
C688 plus.n23 gnd 0.030804f
C689 plus.n24 gnd 0.023652f
C690 plus.n25 gnd 0.023652f
C691 plus.n26 gnd 0.029422f
C692 plus.n27 gnd 0.027651f
C693 plus.n28 gnd 0.160852f
C694 plus.n29 gnd 0.029629f
C695 plus.n30 gnd 0.023652f
C696 plus.n31 gnd 0.023652f
C697 plus.n32 gnd 0.023652f
C698 plus.n33 gnd 0.030428f
C699 plus.n34 gnd 0.160852f
C700 plus.n35 gnd 0.028536f
C701 plus.n36 gnd 0.028536f
C702 plus.n37 gnd 0.023652f
C703 plus.n38 gnd 0.023652f
C704 plus.n39 gnd 0.030428f
C705 plus.n40 gnd 0.019224f
C706 plus.n41 gnd 0.029629f
C707 plus.n42 gnd 0.023652f
C708 plus.n43 gnd 0.023652f
C709 plus.n44 gnd 0.027651f
C710 plus.n45 gnd 0.029422f
C711 plus.n46 gnd 0.160852f
C712 plus.n47 gnd 0.030804f
C713 plus.n48 gnd 0.023652f
C714 plus.n49 gnd 0.023652f
C715 plus.n50 gnd 0.023652f
C716 plus.n51 gnd 0.028265f
C717 plus.n52 gnd 0.160852f
C718 plus.n53 gnd 0.026765f
C719 plus.n54 gnd 0.030307f
C720 plus.n55 gnd 0.023652f
C721 plus.n56 gnd 0.023652f
C722 plus.n57 gnd 0.030855f
C723 plus.n58 gnd 0.008596f
C724 plus.n59 gnd 0.18624f
C725 plus.n60 gnd 0.270994f
C726 plus.n61 gnd 0.023652f
C727 plus.t28 gnd 0.397712f
C728 plus.n62 gnd 0.160852f
C729 plus.n63 gnd 0.023652f
C730 plus.t26 gnd 0.397712f
C731 plus.n64 gnd 0.020211f
C732 plus.n65 gnd 0.023652f
C733 plus.t10 gnd 0.397712f
C734 plus.t15 gnd 0.397712f
C735 plus.n66 gnd 0.160852f
C736 plus.n67 gnd 0.023652f
C737 plus.t13 gnd 0.397712f
C738 plus.n68 gnd 0.160852f
C739 plus.n69 gnd 0.023652f
C740 plus.t17 gnd 0.397712f
C741 plus.n70 gnd 0.019224f
C742 plus.n71 gnd 0.023652f
C743 plus.t16 gnd 0.397712f
C744 plus.t21 gnd 0.397712f
C745 plus.n72 gnd 0.160852f
C746 plus.n73 gnd 0.023652f
C747 plus.t22 gnd 0.397712f
C748 plus.n74 gnd 0.160852f
C749 plus.n75 gnd 0.100378f
C750 plus.t5 gnd 0.397712f
C751 plus.t11 gnd 0.444913f
C752 plus.n76 gnd 0.188053f
C753 plus.n77 gnd 0.184206f
C754 plus.n78 gnd 0.030307f
C755 plus.n79 gnd 0.026765f
C756 plus.n80 gnd 0.023652f
C757 plus.n81 gnd 0.023652f
C758 plus.n82 gnd 0.028265f
C759 plus.n83 gnd 0.020211f
C760 plus.n84 gnd 0.030804f
C761 plus.n85 gnd 0.023652f
C762 plus.n86 gnd 0.023652f
C763 plus.n87 gnd 0.029422f
C764 plus.n88 gnd 0.027651f
C765 plus.n89 gnd 0.160852f
C766 plus.n90 gnd 0.029629f
C767 plus.n91 gnd 0.023652f
C768 plus.n92 gnd 0.023652f
C769 plus.n93 gnd 0.023652f
C770 plus.n94 gnd 0.030428f
C771 plus.n95 gnd 0.160852f
C772 plus.n96 gnd 0.028536f
C773 plus.n97 gnd 0.028536f
C774 plus.n98 gnd 0.023652f
C775 plus.n99 gnd 0.023652f
C776 plus.n100 gnd 0.030428f
C777 plus.n101 gnd 0.019224f
C778 plus.n102 gnd 0.029629f
C779 plus.n103 gnd 0.023652f
C780 plus.n104 gnd 0.023652f
C781 plus.n105 gnd 0.027651f
C782 plus.n106 gnd 0.029422f
C783 plus.n107 gnd 0.160852f
C784 plus.n108 gnd 0.030804f
C785 plus.n109 gnd 0.023652f
C786 plus.n110 gnd 0.023652f
C787 plus.n111 gnd 0.023652f
C788 plus.n112 gnd 0.028265f
C789 plus.n113 gnd 0.160852f
C790 plus.n114 gnd 0.026765f
C791 plus.n115 gnd 0.030307f
C792 plus.n116 gnd 0.023652f
C793 plus.n117 gnd 0.023652f
C794 plus.n118 gnd 0.030855f
C795 plus.n119 gnd 0.008596f
C796 plus.t24 gnd 0.430126f
C797 plus.n120 gnd 0.18624f
C798 plus.n121 gnd 0.853371f
C799 plus.n122 gnd 1.25804f
C800 plus.t1 gnd 0.040831f
C801 plus.t2 gnd 0.007291f
C802 plus.t4 gnd 0.007291f
C803 plus.n123 gnd 0.023647f
C804 plus.n124 gnd 0.183575f
C805 plus.t3 gnd 0.007291f
C806 plus.t0 gnd 0.007291f
C807 plus.n125 gnd 0.023647f
C808 plus.n126 gnd 0.137795f
C809 plus.n127 gnd 2.64316f
C810 a_n1808_13878.t4 gnd 0.185195f
C811 a_n1808_13878.t0 gnd 0.185195f
C812 a_n1808_13878.t2 gnd 0.185195f
C813 a_n1808_13878.n0 gnd 1.4598f
C814 a_n1808_13878.t6 gnd 0.185195f
C815 a_n1808_13878.t1 gnd 0.185195f
C816 a_n1808_13878.n1 gnd 1.45825f
C817 a_n1808_13878.n2 gnd 2.03762f
C818 a_n1808_13878.t5 gnd 0.185195f
C819 a_n1808_13878.t9 gnd 0.185195f
C820 a_n1808_13878.n3 gnd 1.46067f
C821 a_n1808_13878.t10 gnd 0.185195f
C822 a_n1808_13878.t3 gnd 0.185195f
C823 a_n1808_13878.n4 gnd 1.45825f
C824 a_n1808_13878.n5 gnd 1.31079f
C825 a_n1808_13878.t7 gnd 0.185195f
C826 a_n1808_13878.t8 gnd 0.185195f
C827 a_n1808_13878.n6 gnd 1.45825f
C828 a_n1808_13878.n7 gnd 1.80025f
C829 a_n1808_13878.t13 gnd 1.73408f
C830 a_n1808_13878.t16 gnd 0.185195f
C831 a_n1808_13878.t17 gnd 0.185195f
C832 a_n1808_13878.n8 gnd 1.30452f
C833 a_n1808_13878.n9 gnd 1.4576f
C834 a_n1808_13878.t12 gnd 1.73062f
C835 a_n1808_13878.n10 gnd 0.733487f
C836 a_n1808_13878.t15 gnd 1.73062f
C837 a_n1808_13878.n11 gnd 0.733487f
C838 a_n1808_13878.t18 gnd 0.185195f
C839 a_n1808_13878.t19 gnd 0.185195f
C840 a_n1808_13878.n12 gnd 1.30452f
C841 a_n1808_13878.n13 gnd 0.74059f
C842 a_n1808_13878.t14 gnd 1.73062f
C843 a_n1808_13878.n14 gnd 1.7272f
C844 a_n1808_13878.n15 gnd 2.51438f
C845 a_n1808_13878.n16 gnd 3.69301f
C846 a_n1808_13878.n17 gnd 1.45826f
C847 a_n1808_13878.t11 gnd 0.185195f
C848 a_n1986_8322.t20 gnd 38.672398f
C849 a_n1986_8322.t22 gnd 27.512402f
C850 a_n1986_8322.t23 gnd 19.268198f
C851 a_n1986_8322.t21 gnd 38.672398f
C852 a_n1986_8322.t2 gnd 0.093533f
C853 a_n1986_8322.t1 gnd 0.875792f
C854 a_n1986_8322.t9 gnd 0.093533f
C855 a_n1986_8322.t4 gnd 0.093533f
C856 a_n1986_8322.n0 gnd 0.658844f
C857 a_n1986_8322.n1 gnd 0.736161f
C858 a_n1986_8322.t7 gnd 0.093533f
C859 a_n1986_8322.t6 gnd 0.093533f
C860 a_n1986_8322.n2 gnd 0.658844f
C861 a_n1986_8322.n3 gnd 0.374034f
C862 a_n1986_8322.t0 gnd 0.874048f
C863 a_n1986_8322.n4 gnd 1.39896f
C864 a_n1986_8322.t14 gnd 0.875792f
C865 a_n1986_8322.t18 gnd 0.093533f
C866 a_n1986_8322.t17 gnd 0.093533f
C867 a_n1986_8322.n5 gnd 0.658844f
C868 a_n1986_8322.n6 gnd 0.736161f
C869 a_n1986_8322.t12 gnd 0.874048f
C870 a_n1986_8322.n7 gnd 0.370446f
C871 a_n1986_8322.t15 gnd 0.874048f
C872 a_n1986_8322.n8 gnd 0.370446f
C873 a_n1986_8322.t13 gnd 0.093533f
C874 a_n1986_8322.t19 gnd 0.093533f
C875 a_n1986_8322.n9 gnd 0.658844f
C876 a_n1986_8322.n10 gnd 0.374034f
C877 a_n1986_8322.t16 gnd 0.874048f
C878 a_n1986_8322.n11 gnd 0.872317f
C879 a_n1986_8322.n12 gnd 1.59071f
C880 a_n1986_8322.n13 gnd 3.20172f
C881 a_n1986_8322.t3 gnd 0.874048f
C882 a_n1986_8322.n14 gnd 0.76652f
C883 a_n1986_8322.t10 gnd 0.875789f
C884 a_n1986_8322.t8 gnd 0.093533f
C885 a_n1986_8322.t5 gnd 0.093533f
C886 a_n1986_8322.n15 gnd 0.658844f
C887 a_n1986_8322.n16 gnd 0.736163f
C888 a_n1986_8322.n17 gnd 0.374032f
C889 a_n1986_8322.n18 gnd 0.658845f
C890 a_n1986_8322.t11 gnd 0.093533f
C891 a_n2848_n452.n0 gnd 3.415f
C892 a_n2848_n452.n1 gnd 0.285666f
C893 a_n2848_n452.n2 gnd 0.492471f
C894 a_n2848_n452.n3 gnd 0.664435f
C895 a_n2848_n452.n4 gnd 0.215942f
C896 a_n2848_n452.n5 gnd 0.282512f
C897 a_n2848_n452.n6 gnd 0.546457f
C898 a_n2848_n452.n7 gnd 0.526038f
C899 a_n2848_n452.n8 gnd 0.204894f
C900 a_n2848_n452.n9 gnd 0.150908f
C901 a_n2848_n452.n10 gnd 0.23718f
C902 a_n2848_n452.n11 gnd 0.183194f
C903 a_n2848_n452.n12 gnd 0.204894f
C904 a_n2848_n452.n13 gnd 1.0063f
C905 a_n2848_n452.n14 gnd 0.150908f
C906 a_n2848_n452.n15 gnd 0.580023f
C907 a_n2848_n452.n16 gnd 0.432289f
C908 a_n2848_n452.n17 gnd 0.215942f
C909 a_n2848_n452.n18 gnd 0.492471f
C910 a_n2848_n452.n19 gnd 0.282512f
C911 a_n2848_n452.n20 gnd 0.438486f
C912 a_n2848_n452.n21 gnd 0.215942f
C913 a_n2848_n452.n22 gnd 0.731535f
C914 a_n2848_n452.n23 gnd 0.282512f
C915 a_n2848_n452.n24 gnd 1.17886f
C916 a_n2848_n452.n25 gnd 1.91568f
C917 a_n2848_n452.n26 gnd 1.14458f
C918 a_n2848_n452.n27 gnd 1.77783f
C919 a_n2848_n452.n28 gnd 0.377489f
C920 a_n2848_n452.n29 gnd 3.11576f
C921 a_n2848_n452.n30 gnd 0.377488f
C922 a_n2848_n452.n31 gnd 3.20158f
C923 a_n2848_n452.n32 gnd 0.008361f
C924 a_n2848_n452.n34 gnd 0.285666f
C925 a_n2848_n452.n35 gnd 0.008361f
C926 a_n2848_n452.n37 gnd 0.285666f
C927 a_n2848_n452.n38 gnd 0.008361f
C928 a_n2848_n452.n39 gnd 0.28526f
C929 a_n2848_n452.n40 gnd 0.008361f
C930 a_n2848_n452.n41 gnd 0.28526f
C931 a_n2848_n452.n42 gnd 0.008361f
C932 a_n2848_n452.n43 gnd 0.28526f
C933 a_n2848_n452.n44 gnd 0.008361f
C934 a_n2848_n452.n45 gnd 0.28526f
C935 a_n2848_n452.n47 gnd 0.285666f
C936 a_n2848_n452.n48 gnd 0.008361f
C937 a_n2848_n452.n50 gnd 0.285666f
C938 a_n2848_n452.t38 gnd 0.14978f
C939 a_n2848_n452.t29 gnd 0.708223f
C940 a_n2848_n452.t37 gnd 0.696704f
C941 a_n2848_n452.t23 gnd 0.696704f
C942 a_n2848_n452.t3 gnd 0.116496f
C943 a_n2848_n452.t19 gnd 0.116496f
C944 a_n2848_n452.n52 gnd 1.03243f
C945 a_n2848_n452.t13 gnd 0.116496f
C946 a_n2848_n452.t17 gnd 0.116496f
C947 a_n2848_n452.n53 gnd 1.0294f
C948 a_n2848_n452.n54 gnd 0.912817f
C949 a_n2848_n452.t47 gnd 0.116496f
C950 a_n2848_n452.t2 gnd 0.116496f
C951 a_n2848_n452.n55 gnd 1.0294f
C952 a_n2848_n452.t20 gnd 0.116496f
C953 a_n2848_n452.t18 gnd 0.116496f
C954 a_n2848_n452.n56 gnd 1.03243f
C955 a_n2848_n452.t11 gnd 0.116496f
C956 a_n2848_n452.t22 gnd 0.116496f
C957 a_n2848_n452.n57 gnd 1.0294f
C958 a_n2848_n452.n58 gnd 0.912817f
C959 a_n2848_n452.t8 gnd 0.116496f
C960 a_n2848_n452.t5 gnd 0.116496f
C961 a_n2848_n452.n59 gnd 1.0294f
C962 a_n2848_n452.t14 gnd 0.116496f
C963 a_n2848_n452.t21 gnd 0.116496f
C964 a_n2848_n452.n60 gnd 1.0294f
C965 a_n2848_n452.n61 gnd 3.15028f
C966 a_n2848_n452.t0 gnd 0.116496f
C967 a_n2848_n452.t7 gnd 0.116496f
C968 a_n2848_n452.n62 gnd 1.0294f
C969 a_n2848_n452.n63 gnd 0.449443f
C970 a_n2848_n452.t10 gnd 0.116496f
C971 a_n2848_n452.t4 gnd 0.116496f
C972 a_n2848_n452.n64 gnd 1.0294f
C973 a_n2848_n452.t6 gnd 0.116496f
C974 a_n2848_n452.t9 gnd 0.116496f
C975 a_n2848_n452.n65 gnd 1.03243f
C976 a_n2848_n452.t1 gnd 0.116496f
C977 a_n2848_n452.t12 gnd 0.116496f
C978 a_n2848_n452.n66 gnd 1.0294f
C979 a_n2848_n452.n67 gnd 0.912814f
C980 a_n2848_n452.t15 gnd 0.116496f
C981 a_n2848_n452.t16 gnd 0.116496f
C982 a_n2848_n452.n68 gnd 1.0294f
C983 a_n2848_n452.t31 gnd 0.696704f
C984 a_n2848_n452.n69 gnd 0.302425f
C985 a_n2848_n452.t41 gnd 0.696704f
C986 a_n2848_n452.t45 gnd 0.708223f
C987 a_n2848_n452.t75 gnd 0.711378f
C988 a_n2848_n452.t58 gnd 0.696704f
C989 a_n2848_n452.t62 gnd 0.696704f
C990 a_n2848_n452.t52 gnd 0.696704f
C991 a_n2848_n452.n70 gnd 0.306315f
C992 a_n2848_n452.t67 gnd 0.696704f
C993 a_n2848_n452.t73 gnd 0.708223f
C994 a_n2848_n452.t26 gnd 1.40246f
C995 a_n2848_n452.t44 gnd 0.14978f
C996 a_n2848_n452.t40 gnd 0.14978f
C997 a_n2848_n452.n71 gnd 1.05505f
C998 a_n2848_n452.t28 gnd 0.14978f
C999 a_n2848_n452.t36 gnd 0.14978f
C1000 a_n2848_n452.n72 gnd 1.05505f
C1001 a_n2848_n452.t34 gnd 1.39967f
C1002 a_n2848_n452.t27 gnd 0.696704f
C1003 a_n2848_n452.n73 gnd 0.306315f
C1004 a_n2848_n452.t35 gnd 0.696704f
C1005 a_n2848_n452.t43 gnd 0.696704f
C1006 a_n2848_n452.t56 gnd 0.696704f
C1007 a_n2848_n452.n74 gnd 0.306315f
C1008 a_n2848_n452.t65 gnd 0.696704f
C1009 a_n2848_n452.t71 gnd 0.696704f
C1010 a_n2848_n452.t70 gnd 0.711378f
C1011 a_n2848_n452.n75 gnd 0.308932f
C1012 a_n2848_n452.t50 gnd 0.696704f
C1013 a_n2848_n452.n76 gnd 0.302425f
C1014 a_n2848_n452.n77 gnd 0.308933f
C1015 a_n2848_n452.t51 gnd 0.708223f
C1016 a_n2848_n452.t25 gnd 0.711378f
C1017 a_n2848_n452.n78 gnd 0.308932f
C1018 a_n2848_n452.t39 gnd 0.696704f
C1019 a_n2848_n452.n79 gnd 0.302425f
C1020 a_n2848_n452.n80 gnd 0.308933f
C1021 a_n2848_n452.t33 gnd 0.708223f
C1022 a_n2848_n452.n81 gnd 1.13204f
C1023 a_n2848_n452.t55 gnd 0.696704f
C1024 a_n2848_n452.n82 gnd 0.302425f
C1025 a_n2848_n452.t61 gnd 0.696704f
C1026 a_n2848_n452.n83 gnd 0.302425f
C1027 a_n2848_n452.t53 gnd 0.696704f
C1028 a_n2848_n452.n84 gnd 0.302425f
C1029 a_n2848_n452.t66 gnd 0.696704f
C1030 a_n2848_n452.n85 gnd 0.302425f
C1031 a_n2848_n452.t57 gnd 0.696704f
C1032 a_n2848_n452.n86 gnd 0.296933f
C1033 a_n2848_n452.t48 gnd 0.696704f
C1034 a_n2848_n452.n87 gnd 0.306315f
C1035 a_n2848_n452.t59 gnd 0.708378f
C1036 a_n2848_n452.t68 gnd 0.696704f
C1037 a_n2848_n452.n88 gnd 0.296933f
C1038 a_n2848_n452.t54 gnd 0.696704f
C1039 a_n2848_n452.n89 gnd 0.306315f
C1040 a_n2848_n452.t63 gnd 0.708378f
C1041 a_n2848_n452.t72 gnd 0.696704f
C1042 a_n2848_n452.n90 gnd 0.296933f
C1043 a_n2848_n452.t60 gnd 0.696704f
C1044 a_n2848_n452.n91 gnd 0.306315f
C1045 a_n2848_n452.t74 gnd 0.708378f
C1046 a_n2848_n452.t64 gnd 0.696704f
C1047 a_n2848_n452.n92 gnd 0.296933f
C1048 a_n2848_n452.t49 gnd 0.696704f
C1049 a_n2848_n452.n93 gnd 0.306315f
C1050 a_n2848_n452.t69 gnd 0.708378f
C1051 a_n2848_n452.n94 gnd 1.33845f
C1052 a_n2848_n452.n95 gnd 0.308933f
C1053 a_n2848_n452.n96 gnd 0.302425f
C1054 a_n2848_n452.n97 gnd 0.308932f
C1055 a_n2848_n452.n98 gnd 0.308933f
C1056 a_n2848_n452.n99 gnd 0.01225f
C1057 a_n2848_n452.n100 gnd 0.302425f
C1058 a_n2848_n452.n101 gnd 0.308933f
C1059 a_n2848_n452.n102 gnd 0.786935f
C1060 a_n2848_n452.t30 gnd 1.39967f
C1061 a_n2848_n452.t46 gnd 1.40246f
C1062 a_n2848_n452.t32 gnd 0.14978f
C1063 a_n2848_n452.t42 gnd 0.14978f
C1064 a_n2848_n452.n103 gnd 1.05505f
C1065 a_n2848_n452.n104 gnd 1.05505f
C1066 a_n2848_n452.t24 gnd 0.14978f
C1067 vdd.t163 gnd 0.03834f
C1068 vdd.t151 gnd 0.03834f
C1069 vdd.n0 gnd 0.302391f
C1070 vdd.t154 gnd 0.03834f
C1071 vdd.t141 gnd 0.03834f
C1072 vdd.n1 gnd 0.301892f
C1073 vdd.n2 gnd 0.278402f
C1074 vdd.t144 gnd 0.03834f
C1075 vdd.t2 gnd 0.03834f
C1076 vdd.n3 gnd 0.301892f
C1077 vdd.n4 gnd 0.140798f
C1078 vdd.t261 gnd 0.03834f
C1079 vdd.t158 gnd 0.03834f
C1080 vdd.n5 gnd 0.301892f
C1081 vdd.n6 gnd 0.132113f
C1082 vdd.t156 gnd 0.03834f
C1083 vdd.t146 gnd 0.03834f
C1084 vdd.n7 gnd 0.302391f
C1085 vdd.t8 gnd 0.03834f
C1086 vdd.t263 gnd 0.03834f
C1087 vdd.n8 gnd 0.301892f
C1088 vdd.n9 gnd 0.278402f
C1089 vdd.t257 gnd 0.03834f
C1090 vdd.t5 gnd 0.03834f
C1091 vdd.n10 gnd 0.301892f
C1092 vdd.n11 gnd 0.140798f
C1093 vdd.t161 gnd 0.03834f
C1094 vdd.t259 gnd 0.03834f
C1095 vdd.n12 gnd 0.301892f
C1096 vdd.n13 gnd 0.132113f
C1097 vdd.n14 gnd 0.093402f
C1098 vdd.t167 gnd 0.0213f
C1099 vdd.t164 gnd 0.0213f
C1100 vdd.n15 gnd 0.196056f
C1101 vdd.t169 gnd 0.0213f
C1102 vdd.t177 gnd 0.0213f
C1103 vdd.n16 gnd 0.195482f
C1104 vdd.n17 gnd 0.3402f
C1105 vdd.t166 gnd 0.0213f
C1106 vdd.t170 gnd 0.0213f
C1107 vdd.n18 gnd 0.195482f
C1108 vdd.n19 gnd 0.140745f
C1109 vdd.t174 gnd 0.0213f
C1110 vdd.t176 gnd 0.0213f
C1111 vdd.n20 gnd 0.196056f
C1112 vdd.t168 gnd 0.0213f
C1113 vdd.t175 gnd 0.0213f
C1114 vdd.n21 gnd 0.195482f
C1115 vdd.n22 gnd 0.3402f
C1116 vdd.t172 gnd 0.0213f
C1117 vdd.t165 gnd 0.0213f
C1118 vdd.n23 gnd 0.195482f
C1119 vdd.n24 gnd 0.140745f
C1120 vdd.t173 gnd 0.0213f
C1121 vdd.t178 gnd 0.0213f
C1122 vdd.n25 gnd 0.195482f
C1123 vdd.t171 gnd 0.0213f
C1124 vdd.t179 gnd 0.0213f
C1125 vdd.n26 gnd 0.195482f
C1126 vdd.n27 gnd 22.286598f
C1127 vdd.n28 gnd 8.13899f
C1128 vdd.n29 gnd 0.005809f
C1129 vdd.n30 gnd 0.005391f
C1130 vdd.n31 gnd 0.002982f
C1131 vdd.n32 gnd 0.006847f
C1132 vdd.n33 gnd 0.002897f
C1133 vdd.n34 gnd 0.003067f
C1134 vdd.n35 gnd 0.005391f
C1135 vdd.n36 gnd 0.002897f
C1136 vdd.n37 gnd 0.006847f
C1137 vdd.n38 gnd 0.003067f
C1138 vdd.n39 gnd 0.005391f
C1139 vdd.n40 gnd 0.002897f
C1140 vdd.n41 gnd 0.005135f
C1141 vdd.n42 gnd 0.005151f
C1142 vdd.t14 gnd 0.01471f
C1143 vdd.n43 gnd 0.03273f
C1144 vdd.n44 gnd 0.170333f
C1145 vdd.n45 gnd 0.002897f
C1146 vdd.n46 gnd 0.003067f
C1147 vdd.n47 gnd 0.006847f
C1148 vdd.n48 gnd 0.006847f
C1149 vdd.n49 gnd 0.003067f
C1150 vdd.n50 gnd 0.002897f
C1151 vdd.n51 gnd 0.005391f
C1152 vdd.n52 gnd 0.005391f
C1153 vdd.n53 gnd 0.002897f
C1154 vdd.n54 gnd 0.003067f
C1155 vdd.n55 gnd 0.006847f
C1156 vdd.n56 gnd 0.006847f
C1157 vdd.n57 gnd 0.003067f
C1158 vdd.n58 gnd 0.002897f
C1159 vdd.n59 gnd 0.005391f
C1160 vdd.n60 gnd 0.005391f
C1161 vdd.n61 gnd 0.002897f
C1162 vdd.n62 gnd 0.003067f
C1163 vdd.n63 gnd 0.006847f
C1164 vdd.n64 gnd 0.006847f
C1165 vdd.n65 gnd 0.016188f
C1166 vdd.n66 gnd 0.002982f
C1167 vdd.n67 gnd 0.002897f
C1168 vdd.n68 gnd 0.013933f
C1169 vdd.n69 gnd 0.009728f
C1170 vdd.t123 gnd 0.03408f
C1171 vdd.t75 gnd 0.03408f
C1172 vdd.n70 gnd 0.234219f
C1173 vdd.n71 gnd 0.184178f
C1174 vdd.t136 gnd 0.03408f
C1175 vdd.t48 gnd 0.03408f
C1176 vdd.n72 gnd 0.234219f
C1177 vdd.n73 gnd 0.14863f
C1178 vdd.t111 gnd 0.03408f
C1179 vdd.t68 gnd 0.03408f
C1180 vdd.n74 gnd 0.234219f
C1181 vdd.n75 gnd 0.14863f
C1182 vdd.t131 gnd 0.03408f
C1183 vdd.t107 gnd 0.03408f
C1184 vdd.n76 gnd 0.234219f
C1185 vdd.n77 gnd 0.14863f
C1186 vdd.t22 gnd 0.03408f
C1187 vdd.t61 gnd 0.03408f
C1188 vdd.n78 gnd 0.234219f
C1189 vdd.n79 gnd 0.14863f
C1190 vdd.t30 gnd 0.03408f
C1191 vdd.t77 gnd 0.03408f
C1192 vdd.n80 gnd 0.234219f
C1193 vdd.n81 gnd 0.14863f
C1194 vdd.t54 gnd 0.03408f
C1195 vdd.t117 gnd 0.03408f
C1196 vdd.n82 gnd 0.234219f
C1197 vdd.n83 gnd 0.14863f
C1198 vdd.n84 gnd 0.005809f
C1199 vdd.n85 gnd 0.005391f
C1200 vdd.n86 gnd 0.002982f
C1201 vdd.n87 gnd 0.006847f
C1202 vdd.n88 gnd 0.002897f
C1203 vdd.n89 gnd 0.003067f
C1204 vdd.n90 gnd 0.005391f
C1205 vdd.n91 gnd 0.002897f
C1206 vdd.n92 gnd 0.006847f
C1207 vdd.n93 gnd 0.003067f
C1208 vdd.n94 gnd 0.005391f
C1209 vdd.n95 gnd 0.002897f
C1210 vdd.n96 gnd 0.005135f
C1211 vdd.n97 gnd 0.005151f
C1212 vdd.t34 gnd 0.01471f
C1213 vdd.n98 gnd 0.03273f
C1214 vdd.n99 gnd 0.170333f
C1215 vdd.n100 gnd 0.002897f
C1216 vdd.n101 gnd 0.003067f
C1217 vdd.n102 gnd 0.006847f
C1218 vdd.n103 gnd 0.006847f
C1219 vdd.n104 gnd 0.003067f
C1220 vdd.n105 gnd 0.002897f
C1221 vdd.n106 gnd 0.005391f
C1222 vdd.n107 gnd 0.005391f
C1223 vdd.n108 gnd 0.002897f
C1224 vdd.n109 gnd 0.003067f
C1225 vdd.n110 gnd 0.006847f
C1226 vdd.n111 gnd 0.006847f
C1227 vdd.n112 gnd 0.003067f
C1228 vdd.n113 gnd 0.002897f
C1229 vdd.n114 gnd 0.005391f
C1230 vdd.n115 gnd 0.005391f
C1231 vdd.n116 gnd 0.002897f
C1232 vdd.n117 gnd 0.003067f
C1233 vdd.n118 gnd 0.006847f
C1234 vdd.n119 gnd 0.006847f
C1235 vdd.n120 gnd 0.016188f
C1236 vdd.n121 gnd 0.002982f
C1237 vdd.n122 gnd 0.002897f
C1238 vdd.n123 gnd 0.013933f
C1239 vdd.n124 gnd 0.009422f
C1240 vdd.n125 gnd 0.110582f
C1241 vdd.n126 gnd 0.005809f
C1242 vdd.n127 gnd 0.005391f
C1243 vdd.n128 gnd 0.002982f
C1244 vdd.n129 gnd 0.006847f
C1245 vdd.n130 gnd 0.002897f
C1246 vdd.n131 gnd 0.003067f
C1247 vdd.n132 gnd 0.005391f
C1248 vdd.n133 gnd 0.002897f
C1249 vdd.n134 gnd 0.006847f
C1250 vdd.n135 gnd 0.003067f
C1251 vdd.n136 gnd 0.005391f
C1252 vdd.n137 gnd 0.002897f
C1253 vdd.n138 gnd 0.005135f
C1254 vdd.n139 gnd 0.005151f
C1255 vdd.t79 gnd 0.01471f
C1256 vdd.n140 gnd 0.03273f
C1257 vdd.n141 gnd 0.170333f
C1258 vdd.n142 gnd 0.002897f
C1259 vdd.n143 gnd 0.003067f
C1260 vdd.n144 gnd 0.006847f
C1261 vdd.n145 gnd 0.006847f
C1262 vdd.n146 gnd 0.003067f
C1263 vdd.n147 gnd 0.002897f
C1264 vdd.n148 gnd 0.005391f
C1265 vdd.n149 gnd 0.005391f
C1266 vdd.n150 gnd 0.002897f
C1267 vdd.n151 gnd 0.003067f
C1268 vdd.n152 gnd 0.006847f
C1269 vdd.n153 gnd 0.006847f
C1270 vdd.n154 gnd 0.003067f
C1271 vdd.n155 gnd 0.002897f
C1272 vdd.n156 gnd 0.005391f
C1273 vdd.n157 gnd 0.005391f
C1274 vdd.n158 gnd 0.002897f
C1275 vdd.n159 gnd 0.003067f
C1276 vdd.n160 gnd 0.006847f
C1277 vdd.n161 gnd 0.006847f
C1278 vdd.n162 gnd 0.016188f
C1279 vdd.n163 gnd 0.002982f
C1280 vdd.n164 gnd 0.002897f
C1281 vdd.n165 gnd 0.013933f
C1282 vdd.n166 gnd 0.009728f
C1283 vdd.t81 gnd 0.03408f
C1284 vdd.t103 gnd 0.03408f
C1285 vdd.n167 gnd 0.234219f
C1286 vdd.n168 gnd 0.184178f
C1287 vdd.t18 gnd 0.03408f
C1288 vdd.t72 gnd 0.03408f
C1289 vdd.n169 gnd 0.234219f
C1290 vdd.n170 gnd 0.14863f
C1291 vdd.t101 gnd 0.03408f
C1292 vdd.t138 gnd 0.03408f
C1293 vdd.n171 gnd 0.234219f
C1294 vdd.n172 gnd 0.14863f
C1295 vdd.t56 gnd 0.03408f
C1296 vdd.t58 gnd 0.03408f
C1297 vdd.n173 gnd 0.234219f
C1298 vdd.n174 gnd 0.14863f
C1299 vdd.t125 gnd 0.03408f
C1300 vdd.t51 gnd 0.03408f
C1301 vdd.n175 gnd 0.234219f
C1302 vdd.n176 gnd 0.14863f
C1303 vdd.t52 gnd 0.03408f
C1304 vdd.t121 gnd 0.03408f
C1305 vdd.n177 gnd 0.234219f
C1306 vdd.n178 gnd 0.14863f
C1307 vdd.t122 gnd 0.03408f
C1308 vdd.t28 gnd 0.03408f
C1309 vdd.n179 gnd 0.234219f
C1310 vdd.n180 gnd 0.14863f
C1311 vdd.n181 gnd 0.005809f
C1312 vdd.n182 gnd 0.005391f
C1313 vdd.n183 gnd 0.002982f
C1314 vdd.n184 gnd 0.006847f
C1315 vdd.n185 gnd 0.002897f
C1316 vdd.n186 gnd 0.003067f
C1317 vdd.n187 gnd 0.005391f
C1318 vdd.n188 gnd 0.002897f
C1319 vdd.n189 gnd 0.006847f
C1320 vdd.n190 gnd 0.003067f
C1321 vdd.n191 gnd 0.005391f
C1322 vdd.n192 gnd 0.002897f
C1323 vdd.n193 gnd 0.005135f
C1324 vdd.n194 gnd 0.005151f
C1325 vdd.t102 gnd 0.01471f
C1326 vdd.n195 gnd 0.03273f
C1327 vdd.n196 gnd 0.170333f
C1328 vdd.n197 gnd 0.002897f
C1329 vdd.n198 gnd 0.003067f
C1330 vdd.n199 gnd 0.006847f
C1331 vdd.n200 gnd 0.006847f
C1332 vdd.n201 gnd 0.003067f
C1333 vdd.n202 gnd 0.002897f
C1334 vdd.n203 gnd 0.005391f
C1335 vdd.n204 gnd 0.005391f
C1336 vdd.n205 gnd 0.002897f
C1337 vdd.n206 gnd 0.003067f
C1338 vdd.n207 gnd 0.006847f
C1339 vdd.n208 gnd 0.006847f
C1340 vdd.n209 gnd 0.003067f
C1341 vdd.n210 gnd 0.002897f
C1342 vdd.n211 gnd 0.005391f
C1343 vdd.n212 gnd 0.005391f
C1344 vdd.n213 gnd 0.002897f
C1345 vdd.n214 gnd 0.003067f
C1346 vdd.n215 gnd 0.006847f
C1347 vdd.n216 gnd 0.006847f
C1348 vdd.n217 gnd 0.016188f
C1349 vdd.n218 gnd 0.002982f
C1350 vdd.n219 gnd 0.002897f
C1351 vdd.n220 gnd 0.013933f
C1352 vdd.n221 gnd 0.009422f
C1353 vdd.n222 gnd 0.065785f
C1354 vdd.n223 gnd 0.237041f
C1355 vdd.n224 gnd 0.005809f
C1356 vdd.n225 gnd 0.005391f
C1357 vdd.n226 gnd 0.002982f
C1358 vdd.n227 gnd 0.006847f
C1359 vdd.n228 gnd 0.002897f
C1360 vdd.n229 gnd 0.003067f
C1361 vdd.n230 gnd 0.005391f
C1362 vdd.n231 gnd 0.002897f
C1363 vdd.n232 gnd 0.006847f
C1364 vdd.n233 gnd 0.003067f
C1365 vdd.n234 gnd 0.005391f
C1366 vdd.n235 gnd 0.002897f
C1367 vdd.n236 gnd 0.005135f
C1368 vdd.n237 gnd 0.005151f
C1369 vdd.t90 gnd 0.01471f
C1370 vdd.n238 gnd 0.03273f
C1371 vdd.n239 gnd 0.170333f
C1372 vdd.n240 gnd 0.002897f
C1373 vdd.n241 gnd 0.003067f
C1374 vdd.n242 gnd 0.006847f
C1375 vdd.n243 gnd 0.006847f
C1376 vdd.n244 gnd 0.003067f
C1377 vdd.n245 gnd 0.002897f
C1378 vdd.n246 gnd 0.005391f
C1379 vdd.n247 gnd 0.005391f
C1380 vdd.n248 gnd 0.002897f
C1381 vdd.n249 gnd 0.003067f
C1382 vdd.n250 gnd 0.006847f
C1383 vdd.n251 gnd 0.006847f
C1384 vdd.n252 gnd 0.003067f
C1385 vdd.n253 gnd 0.002897f
C1386 vdd.n254 gnd 0.005391f
C1387 vdd.n255 gnd 0.005391f
C1388 vdd.n256 gnd 0.002897f
C1389 vdd.n257 gnd 0.003067f
C1390 vdd.n258 gnd 0.006847f
C1391 vdd.n259 gnd 0.006847f
C1392 vdd.n260 gnd 0.016188f
C1393 vdd.n261 gnd 0.002982f
C1394 vdd.n262 gnd 0.002897f
C1395 vdd.n263 gnd 0.013933f
C1396 vdd.n264 gnd 0.009728f
C1397 vdd.t91 gnd 0.03408f
C1398 vdd.t115 gnd 0.03408f
C1399 vdd.n265 gnd 0.234219f
C1400 vdd.n266 gnd 0.184178f
C1401 vdd.t39 gnd 0.03408f
C1402 vdd.t89 gnd 0.03408f
C1403 vdd.n267 gnd 0.234219f
C1404 vdd.n268 gnd 0.14863f
C1405 vdd.t110 gnd 0.03408f
C1406 vdd.t36 gnd 0.03408f
C1407 vdd.n269 gnd 0.234219f
C1408 vdd.n270 gnd 0.14863f
C1409 vdd.t69 gnd 0.03408f
C1410 vdd.t71 gnd 0.03408f
C1411 vdd.n271 gnd 0.234219f
C1412 vdd.n272 gnd 0.14863f
C1413 vdd.t134 gnd 0.03408f
C1414 vdd.t64 gnd 0.03408f
C1415 vdd.n273 gnd 0.234219f
C1416 vdd.n274 gnd 0.14863f
C1417 vdd.t65 gnd 0.03408f
C1418 vdd.t132 gnd 0.03408f
C1419 vdd.n275 gnd 0.234219f
C1420 vdd.n276 gnd 0.14863f
C1421 vdd.t133 gnd 0.03408f
C1422 vdd.t44 gnd 0.03408f
C1423 vdd.n277 gnd 0.234219f
C1424 vdd.n278 gnd 0.14863f
C1425 vdd.n279 gnd 0.005809f
C1426 vdd.n280 gnd 0.005391f
C1427 vdd.n281 gnd 0.002982f
C1428 vdd.n282 gnd 0.006847f
C1429 vdd.n283 gnd 0.002897f
C1430 vdd.n284 gnd 0.003067f
C1431 vdd.n285 gnd 0.005391f
C1432 vdd.n286 gnd 0.002897f
C1433 vdd.n287 gnd 0.006847f
C1434 vdd.n288 gnd 0.003067f
C1435 vdd.n289 gnd 0.005391f
C1436 vdd.n290 gnd 0.002897f
C1437 vdd.n291 gnd 0.005135f
C1438 vdd.n292 gnd 0.005151f
C1439 vdd.t116 gnd 0.01471f
C1440 vdd.n293 gnd 0.03273f
C1441 vdd.n294 gnd 0.170333f
C1442 vdd.n295 gnd 0.002897f
C1443 vdd.n296 gnd 0.003067f
C1444 vdd.n297 gnd 0.006847f
C1445 vdd.n298 gnd 0.006847f
C1446 vdd.n299 gnd 0.003067f
C1447 vdd.n300 gnd 0.002897f
C1448 vdd.n301 gnd 0.005391f
C1449 vdd.n302 gnd 0.005391f
C1450 vdd.n303 gnd 0.002897f
C1451 vdd.n304 gnd 0.003067f
C1452 vdd.n305 gnd 0.006847f
C1453 vdd.n306 gnd 0.006847f
C1454 vdd.n307 gnd 0.003067f
C1455 vdd.n308 gnd 0.002897f
C1456 vdd.n309 gnd 0.005391f
C1457 vdd.n310 gnd 0.005391f
C1458 vdd.n311 gnd 0.002897f
C1459 vdd.n312 gnd 0.003067f
C1460 vdd.n313 gnd 0.006847f
C1461 vdd.n314 gnd 0.006847f
C1462 vdd.n315 gnd 0.016188f
C1463 vdd.n316 gnd 0.002982f
C1464 vdd.n317 gnd 0.002897f
C1465 vdd.n318 gnd 0.013933f
C1466 vdd.n319 gnd 0.009422f
C1467 vdd.n320 gnd 0.065785f
C1468 vdd.n321 gnd 0.265454f
C1469 vdd.n322 gnd 0.008136f
C1470 vdd.n323 gnd 0.010585f
C1471 vdd.n324 gnd 0.00852f
C1472 vdd.n325 gnd 0.00852f
C1473 vdd.n326 gnd 0.010585f
C1474 vdd.n327 gnd 0.010585f
C1475 vdd.n328 gnd 0.773468f
C1476 vdd.n329 gnd 0.010585f
C1477 vdd.n330 gnd 0.010585f
C1478 vdd.n331 gnd 0.010585f
C1479 vdd.n332 gnd 0.838374f
C1480 vdd.n333 gnd 0.010585f
C1481 vdd.n334 gnd 0.010585f
C1482 vdd.n335 gnd 0.010585f
C1483 vdd.n336 gnd 0.010585f
C1484 vdd.n337 gnd 0.00852f
C1485 vdd.n338 gnd 0.010585f
C1486 vdd.t50 gnd 0.540887f
C1487 vdd.n339 gnd 0.010585f
C1488 vdd.n340 gnd 0.010585f
C1489 vdd.n341 gnd 0.010585f
C1490 vdd.t76 gnd 0.540887f
C1491 vdd.n342 gnd 0.010585f
C1492 vdd.n343 gnd 0.010585f
C1493 vdd.n344 gnd 0.010585f
C1494 vdd.n345 gnd 0.010585f
C1495 vdd.n346 gnd 0.010585f
C1496 vdd.n347 gnd 0.00852f
C1497 vdd.n348 gnd 0.010585f
C1498 vdd.n349 gnd 0.611202f
C1499 vdd.n350 gnd 0.010585f
C1500 vdd.n351 gnd 0.010585f
C1501 vdd.n352 gnd 0.010585f
C1502 vdd.t27 gnd 0.540887f
C1503 vdd.n353 gnd 0.010585f
C1504 vdd.n354 gnd 0.010585f
C1505 vdd.n355 gnd 0.010585f
C1506 vdd.n356 gnd 0.010585f
C1507 vdd.n357 gnd 0.010585f
C1508 vdd.n358 gnd 0.00852f
C1509 vdd.n359 gnd 0.010585f
C1510 vdd.t33 gnd 0.540887f
C1511 vdd.n360 gnd 0.010585f
C1512 vdd.n361 gnd 0.010585f
C1513 vdd.n362 gnd 0.010585f
C1514 vdd.n363 gnd 0.914099f
C1515 vdd.n364 gnd 0.010585f
C1516 vdd.n365 gnd 0.010585f
C1517 vdd.n366 gnd 0.010585f
C1518 vdd.n367 gnd 0.010585f
C1519 vdd.n368 gnd 0.010585f
C1520 vdd.n369 gnd 0.007072f
C1521 vdd.n370 gnd 0.024105f
C1522 vdd.t189 gnd 0.540887f
C1523 vdd.n371 gnd 0.010585f
C1524 vdd.n372 gnd 0.024105f
C1525 vdd.n404 gnd 0.010585f
C1526 vdd.t191 gnd 0.130228f
C1527 vdd.t190 gnd 0.139178f
C1528 vdd.t188 gnd 0.170076f
C1529 vdd.n405 gnd 0.218013f
C1530 vdd.n406 gnd 0.184022f
C1531 vdd.n407 gnd 0.013973f
C1532 vdd.n408 gnd 0.010585f
C1533 vdd.n409 gnd 0.00852f
C1534 vdd.n410 gnd 0.010585f
C1535 vdd.n411 gnd 0.00852f
C1536 vdd.n412 gnd 0.010585f
C1537 vdd.n413 gnd 0.00852f
C1538 vdd.n414 gnd 0.010585f
C1539 vdd.n415 gnd 0.00852f
C1540 vdd.n416 gnd 0.010585f
C1541 vdd.n417 gnd 0.00852f
C1542 vdd.n418 gnd 0.010585f
C1543 vdd.t246 gnd 0.130228f
C1544 vdd.t245 gnd 0.139178f
C1545 vdd.t244 gnd 0.170076f
C1546 vdd.n419 gnd 0.218013f
C1547 vdd.n420 gnd 0.184022f
C1548 vdd.n421 gnd 0.00852f
C1549 vdd.n422 gnd 0.010585f
C1550 vdd.n423 gnd 0.00852f
C1551 vdd.n424 gnd 0.010585f
C1552 vdd.n425 gnd 0.00852f
C1553 vdd.n426 gnd 0.010585f
C1554 vdd.n427 gnd 0.00852f
C1555 vdd.n428 gnd 0.010585f
C1556 vdd.n429 gnd 0.00852f
C1557 vdd.n430 gnd 0.010585f
C1558 vdd.t252 gnd 0.130228f
C1559 vdd.t251 gnd 0.139178f
C1560 vdd.t250 gnd 0.170076f
C1561 vdd.n431 gnd 0.218013f
C1562 vdd.n432 gnd 0.184022f
C1563 vdd.n433 gnd 0.018233f
C1564 vdd.n434 gnd 0.010585f
C1565 vdd.n435 gnd 0.00852f
C1566 vdd.n436 gnd 0.010585f
C1567 vdd.n437 gnd 0.00852f
C1568 vdd.n438 gnd 0.010585f
C1569 vdd.n439 gnd 0.00852f
C1570 vdd.n440 gnd 0.010585f
C1571 vdd.n441 gnd 0.00852f
C1572 vdd.n442 gnd 0.010585f
C1573 vdd.n443 gnd 0.024105f
C1574 vdd.n444 gnd 0.02427f
C1575 vdd.n445 gnd 0.02427f
C1576 vdd.n446 gnd 0.007072f
C1577 vdd.n447 gnd 0.00852f
C1578 vdd.n448 gnd 0.010585f
C1579 vdd.n449 gnd 0.010585f
C1580 vdd.n450 gnd 0.00852f
C1581 vdd.n451 gnd 0.010585f
C1582 vdd.n452 gnd 0.010585f
C1583 vdd.n453 gnd 0.010585f
C1584 vdd.n454 gnd 0.010585f
C1585 vdd.n455 gnd 0.010585f
C1586 vdd.n456 gnd 0.00852f
C1587 vdd.n457 gnd 0.00852f
C1588 vdd.n458 gnd 0.010585f
C1589 vdd.n459 gnd 0.010585f
C1590 vdd.n460 gnd 0.00852f
C1591 vdd.n461 gnd 0.010585f
C1592 vdd.n462 gnd 0.010585f
C1593 vdd.n463 gnd 0.010585f
C1594 vdd.n464 gnd 0.010585f
C1595 vdd.n465 gnd 0.010585f
C1596 vdd.n466 gnd 0.00852f
C1597 vdd.n467 gnd 0.00852f
C1598 vdd.n468 gnd 0.010585f
C1599 vdd.n469 gnd 0.010585f
C1600 vdd.n470 gnd 0.00852f
C1601 vdd.n471 gnd 0.010585f
C1602 vdd.n472 gnd 0.010585f
C1603 vdd.n473 gnd 0.010585f
C1604 vdd.n474 gnd 0.010585f
C1605 vdd.n475 gnd 0.010585f
C1606 vdd.n476 gnd 0.00852f
C1607 vdd.n477 gnd 0.00852f
C1608 vdd.n478 gnd 0.010585f
C1609 vdd.n479 gnd 0.010585f
C1610 vdd.n480 gnd 0.00852f
C1611 vdd.n481 gnd 0.010585f
C1612 vdd.n482 gnd 0.010585f
C1613 vdd.n483 gnd 0.010585f
C1614 vdd.n484 gnd 0.010585f
C1615 vdd.n485 gnd 0.010585f
C1616 vdd.n486 gnd 0.00852f
C1617 vdd.n487 gnd 0.00852f
C1618 vdd.n488 gnd 0.010585f
C1619 vdd.n489 gnd 0.010585f
C1620 vdd.n490 gnd 0.007114f
C1621 vdd.n491 gnd 0.010585f
C1622 vdd.n492 gnd 0.010585f
C1623 vdd.n493 gnd 0.010585f
C1624 vdd.n494 gnd 0.010585f
C1625 vdd.n495 gnd 0.010585f
C1626 vdd.n496 gnd 0.007114f
C1627 vdd.n497 gnd 0.00852f
C1628 vdd.n498 gnd 0.010585f
C1629 vdd.n499 gnd 0.010585f
C1630 vdd.n500 gnd 0.00852f
C1631 vdd.n501 gnd 0.010585f
C1632 vdd.n502 gnd 0.010585f
C1633 vdd.n503 gnd 0.010585f
C1634 vdd.n504 gnd 0.010585f
C1635 vdd.n505 gnd 0.010585f
C1636 vdd.n506 gnd 0.00852f
C1637 vdd.n507 gnd 0.00852f
C1638 vdd.n508 gnd 0.010585f
C1639 vdd.n509 gnd 0.010585f
C1640 vdd.n510 gnd 0.00852f
C1641 vdd.n511 gnd 0.010585f
C1642 vdd.n512 gnd 0.010585f
C1643 vdd.n513 gnd 0.010585f
C1644 vdd.n514 gnd 0.010585f
C1645 vdd.n515 gnd 0.010585f
C1646 vdd.n516 gnd 0.00852f
C1647 vdd.n517 gnd 0.00852f
C1648 vdd.n518 gnd 0.010585f
C1649 vdd.n519 gnd 0.010585f
C1650 vdd.n520 gnd 0.00852f
C1651 vdd.n521 gnd 0.010585f
C1652 vdd.n522 gnd 0.010585f
C1653 vdd.n523 gnd 0.010585f
C1654 vdd.n524 gnd 0.010585f
C1655 vdd.n525 gnd 0.010585f
C1656 vdd.n526 gnd 0.00852f
C1657 vdd.n527 gnd 0.00852f
C1658 vdd.n528 gnd 0.010585f
C1659 vdd.n529 gnd 0.010585f
C1660 vdd.n530 gnd 0.00852f
C1661 vdd.n531 gnd 0.010585f
C1662 vdd.n532 gnd 0.010585f
C1663 vdd.n533 gnd 0.010585f
C1664 vdd.n534 gnd 0.010585f
C1665 vdd.n535 gnd 0.010585f
C1666 vdd.n536 gnd 0.00852f
C1667 vdd.n537 gnd 0.00852f
C1668 vdd.n538 gnd 0.010585f
C1669 vdd.n539 gnd 0.010585f
C1670 vdd.n540 gnd 0.00852f
C1671 vdd.n541 gnd 0.010585f
C1672 vdd.n542 gnd 0.010585f
C1673 vdd.n543 gnd 0.010585f
C1674 vdd.n544 gnd 0.010585f
C1675 vdd.n545 gnd 0.010585f
C1676 vdd.n546 gnd 0.005794f
C1677 vdd.n547 gnd 0.018233f
C1678 vdd.n548 gnd 0.010585f
C1679 vdd.n549 gnd 0.010585f
C1680 vdd.n550 gnd 0.008435f
C1681 vdd.n551 gnd 0.010585f
C1682 vdd.n552 gnd 0.010585f
C1683 vdd.n553 gnd 0.010585f
C1684 vdd.n554 gnd 0.010585f
C1685 vdd.n555 gnd 0.010585f
C1686 vdd.n556 gnd 0.00852f
C1687 vdd.n557 gnd 0.00852f
C1688 vdd.n558 gnd 0.010585f
C1689 vdd.n559 gnd 0.010585f
C1690 vdd.n560 gnd 0.00852f
C1691 vdd.n561 gnd 0.010585f
C1692 vdd.n562 gnd 0.010585f
C1693 vdd.n563 gnd 0.010585f
C1694 vdd.n564 gnd 0.010585f
C1695 vdd.n565 gnd 0.010585f
C1696 vdd.n566 gnd 0.00852f
C1697 vdd.n567 gnd 0.00852f
C1698 vdd.n568 gnd 0.010585f
C1699 vdd.n569 gnd 0.010585f
C1700 vdd.n570 gnd 0.00852f
C1701 vdd.n571 gnd 0.010585f
C1702 vdd.n572 gnd 0.010585f
C1703 vdd.n573 gnd 0.010585f
C1704 vdd.n574 gnd 0.010585f
C1705 vdd.n575 gnd 0.010585f
C1706 vdd.n576 gnd 0.00852f
C1707 vdd.n577 gnd 0.00852f
C1708 vdd.n578 gnd 0.010585f
C1709 vdd.n579 gnd 0.010585f
C1710 vdd.n580 gnd 0.00852f
C1711 vdd.n581 gnd 0.010585f
C1712 vdd.n582 gnd 0.010585f
C1713 vdd.n583 gnd 0.010585f
C1714 vdd.n584 gnd 0.010585f
C1715 vdd.n585 gnd 0.010585f
C1716 vdd.n586 gnd 0.00852f
C1717 vdd.n587 gnd 0.00852f
C1718 vdd.n588 gnd 0.010585f
C1719 vdd.n589 gnd 0.010585f
C1720 vdd.n590 gnd 0.00852f
C1721 vdd.n591 gnd 0.010585f
C1722 vdd.n592 gnd 0.010585f
C1723 vdd.n593 gnd 0.010585f
C1724 vdd.n594 gnd 0.010585f
C1725 vdd.n595 gnd 0.010585f
C1726 vdd.n596 gnd 0.00852f
C1727 vdd.n597 gnd 0.010585f
C1728 vdd.n598 gnd 0.00852f
C1729 vdd.n599 gnd 0.004473f
C1730 vdd.n600 gnd 0.010585f
C1731 vdd.n601 gnd 0.010585f
C1732 vdd.n602 gnd 0.00852f
C1733 vdd.n603 gnd 0.010585f
C1734 vdd.n604 gnd 0.00852f
C1735 vdd.n605 gnd 0.010585f
C1736 vdd.n606 gnd 0.00852f
C1737 vdd.n607 gnd 0.010585f
C1738 vdd.n608 gnd 0.00852f
C1739 vdd.n609 gnd 0.010585f
C1740 vdd.n610 gnd 0.00852f
C1741 vdd.n611 gnd 0.010585f
C1742 vdd.n612 gnd 0.010585f
C1743 vdd.n613 gnd 0.589566f
C1744 vdd.t55 gnd 0.540887f
C1745 vdd.n614 gnd 0.010585f
C1746 vdd.n615 gnd 0.00852f
C1747 vdd.n616 gnd 0.010585f
C1748 vdd.n617 gnd 0.00852f
C1749 vdd.n618 gnd 0.010585f
C1750 vdd.t100 gnd 0.540887f
C1751 vdd.n619 gnd 0.010585f
C1752 vdd.n620 gnd 0.00852f
C1753 vdd.n621 gnd 0.010585f
C1754 vdd.n622 gnd 0.00852f
C1755 vdd.n623 gnd 0.010585f
C1756 vdd.t47 gnd 0.540887f
C1757 vdd.n624 gnd 0.676108f
C1758 vdd.n625 gnd 0.010585f
C1759 vdd.n626 gnd 0.00852f
C1760 vdd.n627 gnd 0.010585f
C1761 vdd.n628 gnd 0.00852f
C1762 vdd.n629 gnd 0.010585f
C1763 vdd.t17 gnd 0.540887f
C1764 vdd.n630 gnd 0.010585f
C1765 vdd.n631 gnd 0.00852f
C1766 vdd.n632 gnd 0.010585f
C1767 vdd.n633 gnd 0.00852f
C1768 vdd.n634 gnd 0.010585f
C1769 vdd.n635 gnd 0.751832f
C1770 vdd.n636 gnd 0.897872f
C1771 vdd.t74 gnd 0.540887f
C1772 vdd.n637 gnd 0.010585f
C1773 vdd.n638 gnd 0.00852f
C1774 vdd.n639 gnd 0.010585f
C1775 vdd.n640 gnd 0.00852f
C1776 vdd.n641 gnd 0.010585f
C1777 vdd.n642 gnd 0.567931f
C1778 vdd.n643 gnd 0.010585f
C1779 vdd.n644 gnd 0.00852f
C1780 vdd.n645 gnd 0.010585f
C1781 vdd.n646 gnd 0.00852f
C1782 vdd.n647 gnd 0.010585f
C1783 vdd.n648 gnd 1.08177f
C1784 vdd.t13 gnd 0.540887f
C1785 vdd.n649 gnd 0.010585f
C1786 vdd.n650 gnd 0.00852f
C1787 vdd.n651 gnd 0.010585f
C1788 vdd.n652 gnd 0.00852f
C1789 vdd.n653 gnd 0.010585f
C1790 vdd.t181 gnd 0.540887f
C1791 vdd.n654 gnd 0.010585f
C1792 vdd.n655 gnd 0.00852f
C1793 vdd.n656 gnd 0.02427f
C1794 vdd.n657 gnd 0.02427f
C1795 vdd.n658 gnd 7.64814f
C1796 vdd.n659 gnd 0.600384f
C1797 vdd.n660 gnd 0.02427f
C1798 vdd.n661 gnd 0.009103f
C1799 vdd.n662 gnd 0.00852f
C1800 vdd.n667 gnd 0.006775f
C1801 vdd.n668 gnd 0.00852f
C1802 vdd.n669 gnd 0.010585f
C1803 vdd.n670 gnd 0.010585f
C1804 vdd.n671 gnd 0.010585f
C1805 vdd.n672 gnd 0.010585f
C1806 vdd.n673 gnd 0.010585f
C1807 vdd.n674 gnd 0.00852f
C1808 vdd.n675 gnd 0.010585f
C1809 vdd.n676 gnd 0.010585f
C1810 vdd.n677 gnd 0.010585f
C1811 vdd.n678 gnd 0.010585f
C1812 vdd.n679 gnd 0.010585f
C1813 vdd.n680 gnd 0.00852f
C1814 vdd.n681 gnd 0.010585f
C1815 vdd.n682 gnd 0.010585f
C1816 vdd.n683 gnd 0.010585f
C1817 vdd.n684 gnd 0.010585f
C1818 vdd.n685 gnd 0.010585f
C1819 vdd.t193 gnd 0.130228f
C1820 vdd.t194 gnd 0.139178f
C1821 vdd.t192 gnd 0.170076f
C1822 vdd.n686 gnd 0.218013f
C1823 vdd.n687 gnd 0.18317f
C1824 vdd.n688 gnd 0.017381f
C1825 vdd.n689 gnd 0.010585f
C1826 vdd.n690 gnd 0.010585f
C1827 vdd.n691 gnd 0.010585f
C1828 vdd.n692 gnd 0.010585f
C1829 vdd.n693 gnd 0.010585f
C1830 vdd.n694 gnd 0.00852f
C1831 vdd.n695 gnd 0.010585f
C1832 vdd.n696 gnd 0.010585f
C1833 vdd.n697 gnd 0.010585f
C1834 vdd.n698 gnd 0.010585f
C1835 vdd.n699 gnd 0.010585f
C1836 vdd.n700 gnd 0.00852f
C1837 vdd.n701 gnd 0.010585f
C1838 vdd.n702 gnd 0.010585f
C1839 vdd.n703 gnd 0.010585f
C1840 vdd.n704 gnd 0.010585f
C1841 vdd.n705 gnd 0.010585f
C1842 vdd.n706 gnd 0.00852f
C1843 vdd.n707 gnd 0.010585f
C1844 vdd.n708 gnd 0.010585f
C1845 vdd.n709 gnd 0.010585f
C1846 vdd.n710 gnd 0.010585f
C1847 vdd.n711 gnd 0.010585f
C1848 vdd.n712 gnd 0.00852f
C1849 vdd.n713 gnd 0.010585f
C1850 vdd.n714 gnd 0.010585f
C1851 vdd.n715 gnd 0.010585f
C1852 vdd.n716 gnd 0.010585f
C1853 vdd.n717 gnd 0.010585f
C1854 vdd.n718 gnd 0.00852f
C1855 vdd.n719 gnd 0.010585f
C1856 vdd.n720 gnd 0.010585f
C1857 vdd.n721 gnd 0.010585f
C1858 vdd.n722 gnd 0.008435f
C1859 vdd.t182 gnd 0.130228f
C1860 vdd.t183 gnd 0.139178f
C1861 vdd.t180 gnd 0.170076f
C1862 vdd.n723 gnd 0.218013f
C1863 vdd.n724 gnd 0.18317f
C1864 vdd.n725 gnd 0.010585f
C1865 vdd.n726 gnd 0.00852f
C1866 vdd.n728 gnd 0.010585f
C1867 vdd.n730 gnd 0.010585f
C1868 vdd.n731 gnd 0.010585f
C1869 vdd.n732 gnd 0.00852f
C1870 vdd.n733 gnd 0.010585f
C1871 vdd.n734 gnd 0.010585f
C1872 vdd.n735 gnd 0.010585f
C1873 vdd.n736 gnd 0.010585f
C1874 vdd.n737 gnd 0.010585f
C1875 vdd.n738 gnd 0.00852f
C1876 vdd.n739 gnd 0.010585f
C1877 vdd.n740 gnd 0.010585f
C1878 vdd.n741 gnd 0.010585f
C1879 vdd.n742 gnd 0.010585f
C1880 vdd.n743 gnd 0.010585f
C1881 vdd.n744 gnd 0.00852f
C1882 vdd.n745 gnd 0.010585f
C1883 vdd.n746 gnd 0.010585f
C1884 vdd.n747 gnd 0.010585f
C1885 vdd.n748 gnd 0.006775f
C1886 vdd.n753 gnd 0.007198f
C1887 vdd.n754 gnd 0.007198f
C1888 vdd.n755 gnd 0.007198f
C1889 vdd.n756 gnd 7.45342f
C1890 vdd.n757 gnd 0.007198f
C1891 vdd.n758 gnd 0.007198f
C1892 vdd.n759 gnd 0.007198f
C1893 vdd.n761 gnd 0.007198f
C1894 vdd.n762 gnd 0.007198f
C1895 vdd.n764 gnd 0.007198f
C1896 vdd.n765 gnd 0.00524f
C1897 vdd.n767 gnd 0.007198f
C1898 vdd.t229 gnd 0.290872f
C1899 vdd.t228 gnd 0.297744f
C1900 vdd.t227 gnd 0.189892f
C1901 vdd.n768 gnd 0.102626f
C1902 vdd.n769 gnd 0.058213f
C1903 vdd.n770 gnd 0.010287f
C1904 vdd.n771 gnd 0.016823f
C1905 vdd.n773 gnd 0.007198f
C1906 vdd.n774 gnd 0.735606f
C1907 vdd.n775 gnd 0.015947f
C1908 vdd.n776 gnd 0.015947f
C1909 vdd.n777 gnd 0.007198f
C1910 vdd.n778 gnd 0.01708f
C1911 vdd.n779 gnd 0.007198f
C1912 vdd.n780 gnd 0.007198f
C1913 vdd.n781 gnd 0.007198f
C1914 vdd.n782 gnd 0.007198f
C1915 vdd.n783 gnd 0.007198f
C1916 vdd.n785 gnd 0.007198f
C1917 vdd.n786 gnd 0.007198f
C1918 vdd.n788 gnd 0.007198f
C1919 vdd.n789 gnd 0.007198f
C1920 vdd.n791 gnd 0.007198f
C1921 vdd.n792 gnd 0.007198f
C1922 vdd.n794 gnd 0.007198f
C1923 vdd.n795 gnd 0.007198f
C1924 vdd.n797 gnd 0.007198f
C1925 vdd.n798 gnd 0.007198f
C1926 vdd.n800 gnd 0.007198f
C1927 vdd.n801 gnd 0.00524f
C1928 vdd.n803 gnd 0.007198f
C1929 vdd.t222 gnd 0.290872f
C1930 vdd.t221 gnd 0.297744f
C1931 vdd.t219 gnd 0.189892f
C1932 vdd.n804 gnd 0.102626f
C1933 vdd.n805 gnd 0.058213f
C1934 vdd.n806 gnd 0.010287f
C1935 vdd.n807 gnd 0.007198f
C1936 vdd.n808 gnd 0.007198f
C1937 vdd.t220 gnd 0.367803f
C1938 vdd.n809 gnd 0.007198f
C1939 vdd.n810 gnd 0.007198f
C1940 vdd.n811 gnd 0.007198f
C1941 vdd.n812 gnd 0.007198f
C1942 vdd.n813 gnd 0.007198f
C1943 vdd.n814 gnd 0.735606f
C1944 vdd.n815 gnd 0.007198f
C1945 vdd.n816 gnd 0.007198f
C1946 vdd.n817 gnd 0.643655f
C1947 vdd.n818 gnd 0.007198f
C1948 vdd.n819 gnd 0.007198f
C1949 vdd.n820 gnd 0.006351f
C1950 vdd.n821 gnd 0.007198f
C1951 vdd.n822 gnd 0.649064f
C1952 vdd.n823 gnd 0.007198f
C1953 vdd.n824 gnd 0.007198f
C1954 vdd.n825 gnd 0.007198f
C1955 vdd.n826 gnd 0.007198f
C1956 vdd.n827 gnd 0.007198f
C1957 vdd.n828 gnd 0.735606f
C1958 vdd.n829 gnd 0.007198f
C1959 vdd.n830 gnd 0.007198f
C1960 vdd.t203 gnd 0.329941f
C1961 vdd.t159 gnd 0.086542f
C1962 vdd.n831 gnd 0.007198f
C1963 vdd.n832 gnd 0.007198f
C1964 vdd.n833 gnd 0.007198f
C1965 vdd.t152 gnd 0.367803f
C1966 vdd.n834 gnd 0.007198f
C1967 vdd.n835 gnd 0.007198f
C1968 vdd.n836 gnd 0.007198f
C1969 vdd.n837 gnd 0.007198f
C1970 vdd.n838 gnd 0.007198f
C1971 vdd.t0 gnd 0.367803f
C1972 vdd.n839 gnd 0.007198f
C1973 vdd.n840 gnd 0.007198f
C1974 vdd.n841 gnd 0.611202f
C1975 vdd.n842 gnd 0.007198f
C1976 vdd.n843 gnd 0.007198f
C1977 vdd.n844 gnd 0.007198f
C1978 vdd.n845 gnd 0.448936f
C1979 vdd.n846 gnd 0.007198f
C1980 vdd.n847 gnd 0.007198f
C1981 vdd.t145 gnd 0.367803f
C1982 vdd.n848 gnd 0.007198f
C1983 vdd.n849 gnd 0.007198f
C1984 vdd.n850 gnd 0.007198f
C1985 vdd.n851 gnd 0.611202f
C1986 vdd.n852 gnd 0.007198f
C1987 vdd.n853 gnd 0.007198f
C1988 vdd.t142 gnd 0.313714f
C1989 vdd.t155 gnd 0.28667f
C1990 vdd.n854 gnd 0.007198f
C1991 vdd.n855 gnd 0.007198f
C1992 vdd.n856 gnd 0.007198f
C1993 vdd.t262 gnd 0.367803f
C1994 vdd.n857 gnd 0.007198f
C1995 vdd.n858 gnd 0.007198f
C1996 vdd.t10 gnd 0.367803f
C1997 vdd.n859 gnd 0.007198f
C1998 vdd.n860 gnd 0.007198f
C1999 vdd.n861 gnd 0.007198f
C2000 vdd.t6 gnd 0.270443f
C2001 vdd.n862 gnd 0.007198f
C2002 vdd.n863 gnd 0.007198f
C2003 vdd.n864 gnd 0.627429f
C2004 vdd.n865 gnd 0.007198f
C2005 vdd.n866 gnd 0.007198f
C2006 vdd.n867 gnd 0.007198f
C2007 vdd.n868 gnd 0.735606f
C2008 vdd.n869 gnd 0.007198f
C2009 vdd.n870 gnd 0.007198f
C2010 vdd.t7 gnd 0.329941f
C2011 vdd.n871 gnd 0.465163f
C2012 vdd.n872 gnd 0.007198f
C2013 vdd.n873 gnd 0.007198f
C2014 vdd.n874 gnd 0.007198f
C2015 vdd.t4 gnd 0.367803f
C2016 vdd.n875 gnd 0.007198f
C2017 vdd.n876 gnd 0.007198f
C2018 vdd.n877 gnd 0.007198f
C2019 vdd.n878 gnd 0.007198f
C2020 vdd.n879 gnd 0.007198f
C2021 vdd.t256 gnd 0.735606f
C2022 vdd.n880 gnd 0.007198f
C2023 vdd.n881 gnd 0.007198f
C2024 vdd.t224 gnd 0.367803f
C2025 vdd.n882 gnd 0.007198f
C2026 vdd.n883 gnd 0.01708f
C2027 vdd.n884 gnd 0.01708f
C2028 vdd.t258 gnd 0.692335f
C2029 vdd.n885 gnd 0.015947f
C2030 vdd.n886 gnd 0.015947f
C2031 vdd.n887 gnd 0.01708f
C2032 vdd.n888 gnd 0.007198f
C2033 vdd.n889 gnd 0.007198f
C2034 vdd.t260 gnd 0.692335f
C2035 vdd.n907 gnd 0.01708f
C2036 vdd.n925 gnd 0.015947f
C2037 vdd.n926 gnd 0.007198f
C2038 vdd.n927 gnd 0.015947f
C2039 vdd.t243 gnd 0.290872f
C2040 vdd.t242 gnd 0.297744f
C2041 vdd.t241 gnd 0.189892f
C2042 vdd.n928 gnd 0.102626f
C2043 vdd.n929 gnd 0.058213f
C2044 vdd.n930 gnd 0.016823f
C2045 vdd.n931 gnd 0.007198f
C2046 vdd.t1 gnd 0.735606f
C2047 vdd.n932 gnd 0.015947f
C2048 vdd.n933 gnd 0.007198f
C2049 vdd.n934 gnd 0.01708f
C2050 vdd.n935 gnd 0.007198f
C2051 vdd.t218 gnd 0.290872f
C2052 vdd.t217 gnd 0.297744f
C2053 vdd.t215 gnd 0.189892f
C2054 vdd.n936 gnd 0.102626f
C2055 vdd.n937 gnd 0.058213f
C2056 vdd.n938 gnd 0.010287f
C2057 vdd.n939 gnd 0.007198f
C2058 vdd.n940 gnd 0.007198f
C2059 vdd.t216 gnd 0.367803f
C2060 vdd.n941 gnd 0.007198f
C2061 vdd.n942 gnd 0.007198f
C2062 vdd.n943 gnd 0.007198f
C2063 vdd.n944 gnd 0.007198f
C2064 vdd.n945 gnd 0.007198f
C2065 vdd.n946 gnd 0.007198f
C2066 vdd.n947 gnd 0.735606f
C2067 vdd.n948 gnd 0.007198f
C2068 vdd.n949 gnd 0.007198f
C2069 vdd.t143 gnd 0.367803f
C2070 vdd.n950 gnd 0.007198f
C2071 vdd.n951 gnd 0.007198f
C2072 vdd.n952 gnd 0.007198f
C2073 vdd.n953 gnd 0.007198f
C2074 vdd.n954 gnd 0.465163f
C2075 vdd.n955 gnd 0.007198f
C2076 vdd.n956 gnd 0.007198f
C2077 vdd.n957 gnd 0.007198f
C2078 vdd.n958 gnd 0.007198f
C2079 vdd.n959 gnd 0.007198f
C2080 vdd.n960 gnd 0.627429f
C2081 vdd.n961 gnd 0.007198f
C2082 vdd.n962 gnd 0.007198f
C2083 vdd.t140 gnd 0.329941f
C2084 vdd.t148 gnd 0.270443f
C2085 vdd.n963 gnd 0.007198f
C2086 vdd.n964 gnd 0.007198f
C2087 vdd.n965 gnd 0.007198f
C2088 vdd.t9 gnd 0.367803f
C2089 vdd.n966 gnd 0.007198f
C2090 vdd.n967 gnd 0.007198f
C2091 vdd.t153 gnd 0.367803f
C2092 vdd.n968 gnd 0.007198f
C2093 vdd.n969 gnd 0.007198f
C2094 vdd.n970 gnd 0.007198f
C2095 vdd.t150 gnd 0.28667f
C2096 vdd.n971 gnd 0.007198f
C2097 vdd.n972 gnd 0.007198f
C2098 vdd.n973 gnd 0.611202f
C2099 vdd.n974 gnd 0.007198f
C2100 vdd.n975 gnd 0.007198f
C2101 vdd.n976 gnd 0.007198f
C2102 vdd.t162 gnd 0.367803f
C2103 vdd.n977 gnd 0.007198f
C2104 vdd.n978 gnd 0.007198f
C2105 vdd.t149 gnd 0.313714f
C2106 vdd.n979 gnd 0.448936f
C2107 vdd.n980 gnd 0.007198f
C2108 vdd.n981 gnd 0.007198f
C2109 vdd.n982 gnd 0.007198f
C2110 vdd.n983 gnd 0.611202f
C2111 vdd.n984 gnd 0.007198f
C2112 vdd.n985 gnd 0.007198f
C2113 vdd.t147 gnd 0.367803f
C2114 vdd.n986 gnd 0.007198f
C2115 vdd.n987 gnd 0.007198f
C2116 vdd.n988 gnd 0.007198f
C2117 vdd.n989 gnd 0.735606f
C2118 vdd.n990 gnd 0.007198f
C2119 vdd.n991 gnd 0.007198f
C2120 vdd.t139 gnd 0.367803f
C2121 vdd.n992 gnd 0.007198f
C2122 vdd.n993 gnd 0.007198f
C2123 vdd.n994 gnd 0.007198f
C2124 vdd.t3 gnd 0.086542f
C2125 vdd.n995 gnd 0.007198f
C2126 vdd.n996 gnd 0.007198f
C2127 vdd.n997 gnd 0.007198f
C2128 vdd.t236 gnd 0.297744f
C2129 vdd.t234 gnd 0.189892f
C2130 vdd.t237 gnd 0.297744f
C2131 vdd.n998 gnd 0.167344f
C2132 vdd.n999 gnd 0.007198f
C2133 vdd.n1000 gnd 0.007198f
C2134 vdd.n1001 gnd 0.735606f
C2135 vdd.n1002 gnd 0.007198f
C2136 vdd.n1003 gnd 0.007198f
C2137 vdd.t235 gnd 0.329941f
C2138 vdd.n1004 gnd 0.649064f
C2139 vdd.n1005 gnd 0.007198f
C2140 vdd.n1006 gnd 0.007198f
C2141 vdd.n1007 gnd 0.007198f
C2142 vdd.n1008 gnd 0.643655f
C2143 vdd.n1009 gnd 0.007198f
C2144 vdd.n1010 gnd 0.007198f
C2145 vdd.n1011 gnd 0.007198f
C2146 vdd.n1012 gnd 0.007198f
C2147 vdd.n1013 gnd 0.007198f
C2148 vdd.n1014 gnd 0.735606f
C2149 vdd.n1015 gnd 0.007198f
C2150 vdd.n1016 gnd 0.007198f
C2151 vdd.t231 gnd 0.367803f
C2152 vdd.n1017 gnd 0.007198f
C2153 vdd.n1018 gnd 0.01708f
C2154 vdd.n1019 gnd 0.01708f
C2155 vdd.n1020 gnd 7.45342f
C2156 vdd.n1021 gnd 0.015947f
C2157 vdd.n1022 gnd 0.015947f
C2158 vdd.n1023 gnd 0.01708f
C2159 vdd.n1024 gnd 0.007198f
C2160 vdd.n1025 gnd 0.007198f
C2161 vdd.n1026 gnd 0.007198f
C2162 vdd.n1027 gnd 0.007198f
C2163 vdd.n1028 gnd 0.007198f
C2164 vdd.n1029 gnd 0.007198f
C2165 vdd.n1030 gnd 0.007198f
C2166 vdd.n1031 gnd 0.007198f
C2167 vdd.n1033 gnd 0.007198f
C2168 vdd.n1034 gnd 0.007198f
C2169 vdd.n1035 gnd 0.006775f
C2170 vdd.n1038 gnd 0.02427f
C2171 vdd.n1039 gnd 0.00852f
C2172 vdd.n1040 gnd 0.010585f
C2173 vdd.n1042 gnd 0.010585f
C2174 vdd.n1043 gnd 0.007072f
C2175 vdd.n1044 gnd 0.600384f
C2176 vdd.n1045 gnd 7.64814f
C2177 vdd.n1046 gnd 0.010585f
C2178 vdd.n1047 gnd 0.02427f
C2179 vdd.n1048 gnd 0.00852f
C2180 vdd.n1049 gnd 0.010585f
C2181 vdd.n1050 gnd 0.00852f
C2182 vdd.n1051 gnd 0.010585f
C2183 vdd.n1052 gnd 1.08177f
C2184 vdd.n1053 gnd 0.010585f
C2185 vdd.n1054 gnd 0.00852f
C2186 vdd.n1055 gnd 0.00852f
C2187 vdd.n1056 gnd 0.010585f
C2188 vdd.n1057 gnd 0.00852f
C2189 vdd.n1058 gnd 0.010585f
C2190 vdd.t11 gnd 0.540887f
C2191 vdd.n1059 gnd 0.010585f
C2192 vdd.n1060 gnd 0.00852f
C2193 vdd.n1061 gnd 0.010585f
C2194 vdd.n1062 gnd 0.00852f
C2195 vdd.n1063 gnd 0.010585f
C2196 vdd.t118 gnd 0.540887f
C2197 vdd.n1064 gnd 0.010585f
C2198 vdd.n1065 gnd 0.00852f
C2199 vdd.n1066 gnd 0.010585f
C2200 vdd.n1067 gnd 0.00852f
C2201 vdd.n1068 gnd 0.010585f
C2202 vdd.t25 gnd 0.540887f
C2203 vdd.n1069 gnd 0.751832f
C2204 vdd.n1070 gnd 0.010585f
C2205 vdd.n1071 gnd 0.00852f
C2206 vdd.n1072 gnd 0.010585f
C2207 vdd.n1073 gnd 0.00852f
C2208 vdd.n1074 gnd 0.010585f
C2209 vdd.n1075 gnd 0.86001f
C2210 vdd.n1076 gnd 0.010585f
C2211 vdd.n1077 gnd 0.00852f
C2212 vdd.n1078 gnd 0.010585f
C2213 vdd.n1079 gnd 0.00852f
C2214 vdd.n1080 gnd 0.010585f
C2215 vdd.n1081 gnd 0.676108f
C2216 vdd.t45 gnd 0.540887f
C2217 vdd.n1082 gnd 0.010585f
C2218 vdd.n1083 gnd 0.00852f
C2219 vdd.n1084 gnd 0.010585f
C2220 vdd.n1085 gnd 0.00852f
C2221 vdd.n1086 gnd 0.010585f
C2222 vdd.t66 gnd 0.540887f
C2223 vdd.n1087 gnd 0.010585f
C2224 vdd.n1088 gnd 0.00852f
C2225 vdd.n1089 gnd 0.010585f
C2226 vdd.n1090 gnd 0.00852f
C2227 vdd.n1091 gnd 0.010585f
C2228 vdd.t96 gnd 0.540887f
C2229 vdd.n1092 gnd 0.589566f
C2230 vdd.n1093 gnd 0.010585f
C2231 vdd.n1094 gnd 0.00852f
C2232 vdd.n1095 gnd 0.010585f
C2233 vdd.n1096 gnd 0.00852f
C2234 vdd.n1097 gnd 0.010585f
C2235 vdd.t87 gnd 0.540887f
C2236 vdd.n1098 gnd 0.010585f
C2237 vdd.n1099 gnd 0.00852f
C2238 vdd.n1100 gnd 0.010585f
C2239 vdd.n1101 gnd 0.00852f
C2240 vdd.n1102 gnd 0.010585f
C2241 vdd.n1103 gnd 0.838374f
C2242 vdd.n1104 gnd 0.897872f
C2243 vdd.t19 gnd 0.540887f
C2244 vdd.n1105 gnd 0.010585f
C2245 vdd.n1106 gnd 0.00852f
C2246 vdd.n1107 gnd 0.010585f
C2247 vdd.n1108 gnd 0.00852f
C2248 vdd.n1109 gnd 0.010585f
C2249 vdd.n1110 gnd 0.654473f
C2250 vdd.n1111 gnd 0.010585f
C2251 vdd.n1112 gnd 0.00852f
C2252 vdd.n1113 gnd 0.010585f
C2253 vdd.n1114 gnd 0.00852f
C2254 vdd.n1115 gnd 0.010585f
C2255 vdd.t42 gnd 0.540887f
C2256 vdd.t31 gnd 0.540887f
C2257 vdd.n1116 gnd 0.010585f
C2258 vdd.n1117 gnd 0.00852f
C2259 vdd.n1118 gnd 0.010585f
C2260 vdd.n1119 gnd 0.00852f
C2261 vdd.n1120 gnd 0.010585f
C2262 vdd.t82 gnd 0.540887f
C2263 vdd.n1121 gnd 0.010585f
C2264 vdd.n1122 gnd 0.00852f
C2265 vdd.n1123 gnd 0.010585f
C2266 vdd.n1124 gnd 0.00852f
C2267 vdd.n1125 gnd 0.010585f
C2268 vdd.t84 gnd 0.540887f
C2269 vdd.n1126 gnd 0.795103f
C2270 vdd.n1127 gnd 0.010585f
C2271 vdd.n1128 gnd 0.00852f
C2272 vdd.n1129 gnd 0.010585f
C2273 vdd.n1130 gnd 0.00852f
C2274 vdd.n1131 gnd 0.010585f
C2275 vdd.n1132 gnd 1.08177f
C2276 vdd.n1133 gnd 0.010585f
C2277 vdd.n1134 gnd 0.00852f
C2278 vdd.n1135 gnd 0.010585f
C2279 vdd.n1136 gnd 0.00852f
C2280 vdd.n1137 gnd 0.010585f
C2281 vdd.n1138 gnd 0.914099f
C2282 vdd.n1139 gnd 0.010585f
C2283 vdd.n1140 gnd 0.00852f
C2284 vdd.n1141 gnd 0.024105f
C2285 vdd.n1142 gnd 0.007072f
C2286 vdd.n1143 gnd 0.024105f
C2287 vdd.n1144 gnd 1.42794f
C2288 vdd.n1145 gnd 0.024105f
C2289 vdd.n1146 gnd 0.007072f
C2290 vdd.n1147 gnd 0.010585f
C2291 vdd.t186 gnd 0.130228f
C2292 vdd.t187 gnd 0.139178f
C2293 vdd.t184 gnd 0.170076f
C2294 vdd.n1148 gnd 0.218013f
C2295 vdd.n1149 gnd 0.184022f
C2296 vdd.n1150 gnd 0.013973f
C2297 vdd.n1151 gnd 0.010585f
C2298 vdd.n1182 gnd 0.010585f
C2299 vdd.n1183 gnd 0.010585f
C2300 vdd.n1184 gnd 0.02427f
C2301 vdd.n1185 gnd 0.00852f
C2302 vdd.n1186 gnd 0.010585f
C2303 vdd.n1187 gnd 0.010585f
C2304 vdd.n1188 gnd 0.010585f
C2305 vdd.n1189 gnd 0.010585f
C2306 vdd.n1190 gnd 0.00852f
C2307 vdd.n1191 gnd 0.010585f
C2308 vdd.n1192 gnd 0.010585f
C2309 vdd.n1193 gnd 0.010585f
C2310 vdd.n1194 gnd 0.010585f
C2311 vdd.n1195 gnd 0.010585f
C2312 vdd.n1196 gnd 0.00852f
C2313 vdd.n1197 gnd 0.010585f
C2314 vdd.n1198 gnd 0.010585f
C2315 vdd.n1199 gnd 0.010585f
C2316 vdd.n1200 gnd 0.010585f
C2317 vdd.n1201 gnd 0.010585f
C2318 vdd.n1202 gnd 0.00852f
C2319 vdd.n1203 gnd 0.010585f
C2320 vdd.n1204 gnd 0.010585f
C2321 vdd.n1205 gnd 0.010585f
C2322 vdd.n1206 gnd 0.010585f
C2323 vdd.n1207 gnd 0.010585f
C2324 vdd.n1208 gnd 0.007114f
C2325 vdd.n1209 gnd 0.010585f
C2326 vdd.n1210 gnd 0.010585f
C2327 vdd.n1211 gnd 0.010585f
C2328 vdd.n1212 gnd 0.00852f
C2329 vdd.n1213 gnd 0.010585f
C2330 vdd.n1214 gnd 0.010585f
C2331 vdd.n1215 gnd 0.010585f
C2332 vdd.n1216 gnd 0.010585f
C2333 vdd.n1217 gnd 0.010585f
C2334 vdd.n1218 gnd 0.00852f
C2335 vdd.n1219 gnd 0.010585f
C2336 vdd.n1220 gnd 0.010585f
C2337 vdd.n1221 gnd 0.010585f
C2338 vdd.n1222 gnd 0.010585f
C2339 vdd.n1223 gnd 0.010585f
C2340 vdd.n1224 gnd 0.00852f
C2341 vdd.n1225 gnd 0.010585f
C2342 vdd.n1226 gnd 0.010585f
C2343 vdd.n1227 gnd 0.010585f
C2344 vdd.n1228 gnd 0.010585f
C2345 vdd.n1229 gnd 0.010585f
C2346 vdd.n1230 gnd 0.00852f
C2347 vdd.n1231 gnd 0.010585f
C2348 vdd.n1232 gnd 0.010585f
C2349 vdd.n1233 gnd 0.010585f
C2350 vdd.n1234 gnd 0.010585f
C2351 vdd.n1235 gnd 0.010585f
C2352 vdd.n1236 gnd 0.00852f
C2353 vdd.n1237 gnd 0.010585f
C2354 vdd.n1238 gnd 0.010585f
C2355 vdd.n1239 gnd 0.010585f
C2356 vdd.n1240 gnd 0.010585f
C2357 vdd.n1241 gnd 0.008435f
C2358 vdd.n1242 gnd 0.010585f
C2359 vdd.n1243 gnd 0.010585f
C2360 vdd.n1244 gnd 0.010585f
C2361 vdd.n1245 gnd 0.010585f
C2362 vdd.n1246 gnd 0.010585f
C2363 vdd.n1247 gnd 0.00852f
C2364 vdd.n1248 gnd 0.010585f
C2365 vdd.n1249 gnd 0.010585f
C2366 vdd.n1250 gnd 0.010585f
C2367 vdd.n1251 gnd 0.010585f
C2368 vdd.n1252 gnd 0.010585f
C2369 vdd.n1253 gnd 0.00852f
C2370 vdd.n1254 gnd 0.010585f
C2371 vdd.n1255 gnd 0.010585f
C2372 vdd.n1256 gnd 0.010585f
C2373 vdd.n1257 gnd 0.010585f
C2374 vdd.n1258 gnd 0.010585f
C2375 vdd.n1259 gnd 0.00852f
C2376 vdd.n1260 gnd 0.010585f
C2377 vdd.n1261 gnd 0.010585f
C2378 vdd.n1262 gnd 0.010585f
C2379 vdd.n1263 gnd 0.010585f
C2380 vdd.n1264 gnd 0.010585f
C2381 vdd.n1265 gnd 0.00852f
C2382 vdd.n1266 gnd 0.010585f
C2383 vdd.n1267 gnd 0.010585f
C2384 vdd.n1268 gnd 0.010585f
C2385 vdd.n1269 gnd 0.010585f
C2386 vdd.n1270 gnd 0.010585f
C2387 vdd.n1271 gnd 0.004473f
C2388 vdd.n1272 gnd 0.010585f
C2389 vdd.n1273 gnd 0.00852f
C2390 vdd.n1274 gnd 0.00852f
C2391 vdd.n1275 gnd 0.00852f
C2392 vdd.n1276 gnd 0.010585f
C2393 vdd.n1277 gnd 0.010585f
C2394 vdd.n1278 gnd 0.010585f
C2395 vdd.n1279 gnd 0.00852f
C2396 vdd.n1280 gnd 0.00852f
C2397 vdd.n1281 gnd 0.00852f
C2398 vdd.n1282 gnd 0.010585f
C2399 vdd.n1283 gnd 0.010585f
C2400 vdd.n1284 gnd 0.010585f
C2401 vdd.n1285 gnd 0.00852f
C2402 vdd.n1286 gnd 0.00852f
C2403 vdd.n1287 gnd 0.00852f
C2404 vdd.n1288 gnd 0.010585f
C2405 vdd.n1289 gnd 0.010585f
C2406 vdd.n1290 gnd 0.010585f
C2407 vdd.n1291 gnd 0.00852f
C2408 vdd.n1292 gnd 0.00852f
C2409 vdd.n1293 gnd 0.00852f
C2410 vdd.n1294 gnd 0.010585f
C2411 vdd.n1295 gnd 0.010585f
C2412 vdd.n1296 gnd 0.010585f
C2413 vdd.n1297 gnd 0.00852f
C2414 vdd.n1298 gnd 0.00852f
C2415 vdd.n1299 gnd 0.00852f
C2416 vdd.n1300 gnd 0.010585f
C2417 vdd.n1301 gnd 0.010585f
C2418 vdd.n1302 gnd 0.010585f
C2419 vdd.n1303 gnd 0.010585f
C2420 vdd.t200 gnd 0.130228f
C2421 vdd.t201 gnd 0.139178f
C2422 vdd.t199 gnd 0.170076f
C2423 vdd.n1304 gnd 0.218013f
C2424 vdd.n1305 gnd 0.184022f
C2425 vdd.n1306 gnd 0.018233f
C2426 vdd.n1307 gnd 0.005794f
C2427 vdd.n1308 gnd 0.00852f
C2428 vdd.n1309 gnd 0.010585f
C2429 vdd.n1310 gnd 0.010585f
C2430 vdd.n1311 gnd 0.010585f
C2431 vdd.n1312 gnd 0.00852f
C2432 vdd.n1313 gnd 0.00852f
C2433 vdd.n1314 gnd 0.00852f
C2434 vdd.n1315 gnd 0.010585f
C2435 vdd.n1316 gnd 0.010585f
C2436 vdd.n1317 gnd 0.010585f
C2437 vdd.n1318 gnd 0.00852f
C2438 vdd.n1319 gnd 0.00852f
C2439 vdd.n1320 gnd 0.00852f
C2440 vdd.n1321 gnd 0.010585f
C2441 vdd.n1322 gnd 0.010585f
C2442 vdd.n1323 gnd 0.010585f
C2443 vdd.n1324 gnd 0.00852f
C2444 vdd.n1325 gnd 0.00852f
C2445 vdd.n1326 gnd 0.00852f
C2446 vdd.n1327 gnd 0.010585f
C2447 vdd.n1328 gnd 0.010585f
C2448 vdd.n1329 gnd 0.010585f
C2449 vdd.n1330 gnd 0.00852f
C2450 vdd.n1331 gnd 0.00852f
C2451 vdd.n1332 gnd 0.00852f
C2452 vdd.n1333 gnd 0.010585f
C2453 vdd.n1334 gnd 0.010585f
C2454 vdd.n1335 gnd 0.010585f
C2455 vdd.n1336 gnd 0.00852f
C2456 vdd.n1337 gnd 0.007114f
C2457 vdd.n1338 gnd 0.010585f
C2458 vdd.n1339 gnd 0.010585f
C2459 vdd.t207 gnd 0.130228f
C2460 vdd.t208 gnd 0.139178f
C2461 vdd.t206 gnd 0.170076f
C2462 vdd.n1340 gnd 0.218013f
C2463 vdd.n1341 gnd 0.184022f
C2464 vdd.n1342 gnd 0.018233f
C2465 vdd.n1343 gnd 0.010585f
C2466 vdd.n1344 gnd 0.010585f
C2467 vdd.n1345 gnd 0.010585f
C2468 vdd.n1346 gnd 0.00852f
C2469 vdd.n1347 gnd 0.00852f
C2470 vdd.n1348 gnd 0.00852f
C2471 vdd.n1349 gnd 0.010585f
C2472 vdd.n1350 gnd 0.010585f
C2473 vdd.n1351 gnd 0.010585f
C2474 vdd.n1352 gnd 0.00852f
C2475 vdd.n1353 gnd 0.00852f
C2476 vdd.n1354 gnd 0.00852f
C2477 vdd.n1355 gnd 0.010585f
C2478 vdd.n1356 gnd 0.010585f
C2479 vdd.n1357 gnd 0.010585f
C2480 vdd.n1358 gnd 0.00852f
C2481 vdd.n1359 gnd 0.00852f
C2482 vdd.n1360 gnd 0.00852f
C2483 vdd.n1361 gnd 0.010585f
C2484 vdd.n1362 gnd 0.010585f
C2485 vdd.n1363 gnd 0.010585f
C2486 vdd.n1364 gnd 0.00852f
C2487 vdd.n1365 gnd 0.00852f
C2488 vdd.n1366 gnd 0.00852f
C2489 vdd.n1367 gnd 0.010585f
C2490 vdd.n1368 gnd 0.010585f
C2491 vdd.n1369 gnd 0.010585f
C2492 vdd.n1370 gnd 0.00852f
C2493 vdd.n1371 gnd 0.007072f
C2494 vdd.n1372 gnd 0.02427f
C2495 vdd.n1374 gnd 2.39072f
C2496 vdd.n1375 gnd 0.02427f
C2497 vdd.n1376 gnd 0.004047f
C2498 vdd.n1377 gnd 0.02427f
C2499 vdd.n1378 gnd 0.024105f
C2500 vdd.n1379 gnd 0.010585f
C2501 vdd.n1380 gnd 0.00852f
C2502 vdd.n1381 gnd 0.010585f
C2503 vdd.t185 gnd 0.540887f
C2504 vdd.n1382 gnd 0.708562f
C2505 vdd.n1383 gnd 0.010585f
C2506 vdd.n1384 gnd 0.00852f
C2507 vdd.n1385 gnd 0.010585f
C2508 vdd.n1386 gnd 0.010585f
C2509 vdd.n1387 gnd 0.010585f
C2510 vdd.n1388 gnd 0.00852f
C2511 vdd.n1389 gnd 0.010585f
C2512 vdd.n1390 gnd 1.08177f
C2513 vdd.n1391 gnd 0.010585f
C2514 vdd.n1392 gnd 0.00852f
C2515 vdd.n1393 gnd 0.010585f
C2516 vdd.n1394 gnd 0.010585f
C2517 vdd.n1395 gnd 0.010585f
C2518 vdd.n1396 gnd 0.00852f
C2519 vdd.n1397 gnd 0.010585f
C2520 vdd.n1398 gnd 0.897872f
C2521 vdd.t23 gnd 0.540887f
C2522 vdd.n1399 gnd 0.62202f
C2523 vdd.n1400 gnd 0.010585f
C2524 vdd.n1401 gnd 0.00852f
C2525 vdd.n1402 gnd 0.010585f
C2526 vdd.n1403 gnd 0.010585f
C2527 vdd.n1404 gnd 0.010585f
C2528 vdd.n1405 gnd 0.00852f
C2529 vdd.n1406 gnd 0.010585f
C2530 vdd.n1407 gnd 0.643655f
C2531 vdd.n1408 gnd 0.010585f
C2532 vdd.n1409 gnd 0.00852f
C2533 vdd.n1410 gnd 0.010585f
C2534 vdd.n1411 gnd 0.010585f
C2535 vdd.n1412 gnd 0.010585f
C2536 vdd.n1413 gnd 0.00852f
C2537 vdd.n1414 gnd 0.010585f
C2538 vdd.n1415 gnd 0.611202f
C2539 vdd.n1416 gnd 0.827557f
C2540 vdd.n1417 gnd 0.010585f
C2541 vdd.n1418 gnd 0.00852f
C2542 vdd.n1419 gnd 0.010585f
C2543 vdd.n1420 gnd 0.010585f
C2544 vdd.n1421 gnd 0.010585f
C2545 vdd.n1422 gnd 0.00852f
C2546 vdd.n1423 gnd 0.010585f
C2547 vdd.n1424 gnd 0.897872f
C2548 vdd.n1425 gnd 0.010585f
C2549 vdd.n1426 gnd 0.00852f
C2550 vdd.n1427 gnd 0.010585f
C2551 vdd.n1428 gnd 0.010585f
C2552 vdd.n1429 gnd 0.010585f
C2553 vdd.n1430 gnd 0.00852f
C2554 vdd.n1431 gnd 0.010585f
C2555 vdd.t59 gnd 0.540887f
C2556 vdd.n1432 gnd 0.784286f
C2557 vdd.n1433 gnd 0.010585f
C2558 vdd.n1434 gnd 0.00852f
C2559 vdd.n1435 gnd 0.010585f
C2560 vdd.n1436 gnd 0.010585f
C2561 vdd.n1437 gnd 0.010585f
C2562 vdd.n1438 gnd 0.00852f
C2563 vdd.n1439 gnd 0.010585f
C2564 vdd.n1440 gnd 0.600384f
C2565 vdd.n1441 gnd 0.010585f
C2566 vdd.n1442 gnd 0.00852f
C2567 vdd.n1443 gnd 0.010585f
C2568 vdd.n1444 gnd 0.010585f
C2569 vdd.n1445 gnd 0.010585f
C2570 vdd.n1446 gnd 0.00852f
C2571 vdd.n1447 gnd 0.010585f
C2572 vdd.n1448 gnd 0.773468f
C2573 vdd.n1449 gnd 0.665291f
C2574 vdd.n1450 gnd 0.010585f
C2575 vdd.n1451 gnd 0.00852f
C2576 vdd.n1452 gnd 0.008136f
C2577 vdd.n1453 gnd 0.005809f
C2578 vdd.n1454 gnd 0.005391f
C2579 vdd.n1455 gnd 0.002982f
C2580 vdd.n1456 gnd 0.006847f
C2581 vdd.n1457 gnd 0.002897f
C2582 vdd.n1458 gnd 0.003067f
C2583 vdd.n1459 gnd 0.005391f
C2584 vdd.n1460 gnd 0.002897f
C2585 vdd.n1461 gnd 0.006847f
C2586 vdd.n1462 gnd 0.003067f
C2587 vdd.n1463 gnd 0.005391f
C2588 vdd.n1464 gnd 0.002897f
C2589 vdd.n1465 gnd 0.005135f
C2590 vdd.n1466 gnd 0.005151f
C2591 vdd.t12 gnd 0.01471f
C2592 vdd.n1467 gnd 0.03273f
C2593 vdd.n1468 gnd 0.170333f
C2594 vdd.n1469 gnd 0.002897f
C2595 vdd.n1470 gnd 0.003067f
C2596 vdd.n1471 gnd 0.006847f
C2597 vdd.n1472 gnd 0.006847f
C2598 vdd.n1473 gnd 0.003067f
C2599 vdd.n1474 gnd 0.002897f
C2600 vdd.n1475 gnd 0.005391f
C2601 vdd.n1476 gnd 0.005391f
C2602 vdd.n1477 gnd 0.002897f
C2603 vdd.n1478 gnd 0.003067f
C2604 vdd.n1479 gnd 0.006847f
C2605 vdd.n1480 gnd 0.006847f
C2606 vdd.n1481 gnd 0.003067f
C2607 vdd.n1482 gnd 0.002897f
C2608 vdd.n1483 gnd 0.005391f
C2609 vdd.n1484 gnd 0.005391f
C2610 vdd.n1485 gnd 0.002897f
C2611 vdd.n1486 gnd 0.003067f
C2612 vdd.n1487 gnd 0.006847f
C2613 vdd.n1488 gnd 0.006847f
C2614 vdd.n1489 gnd 0.016188f
C2615 vdd.n1490 gnd 0.002982f
C2616 vdd.n1491 gnd 0.002897f
C2617 vdd.n1492 gnd 0.013933f
C2618 vdd.n1493 gnd 0.009728f
C2619 vdd.t73 gnd 0.03408f
C2620 vdd.t124 gnd 0.03408f
C2621 vdd.n1494 gnd 0.234219f
C2622 vdd.n1495 gnd 0.184178f
C2623 vdd.t46 gnd 0.03408f
C2624 vdd.t106 gnd 0.03408f
C2625 vdd.n1496 gnd 0.234219f
C2626 vdd.n1497 gnd 0.14863f
C2627 vdd.t67 gnd 0.03408f
C2628 vdd.t113 gnd 0.03408f
C2629 vdd.n1498 gnd 0.234219f
C2630 vdd.n1499 gnd 0.14863f
C2631 vdd.t88 gnd 0.03408f
C2632 vdd.t130 gnd 0.03408f
C2633 vdd.n1500 gnd 0.234219f
C2634 vdd.n1501 gnd 0.14863f
C2635 vdd.t60 gnd 0.03408f
C2636 vdd.t20 gnd 0.03408f
C2637 vdd.n1502 gnd 0.234219f
C2638 vdd.n1503 gnd 0.14863f
C2639 vdd.t78 gnd 0.03408f
C2640 vdd.t32 gnd 0.03408f
C2641 vdd.n1504 gnd 0.234219f
C2642 vdd.n1505 gnd 0.14863f
C2643 vdd.t120 gnd 0.03408f
C2644 vdd.t135 gnd 0.03408f
C2645 vdd.n1506 gnd 0.234219f
C2646 vdd.n1507 gnd 0.14863f
C2647 vdd.n1508 gnd 0.005809f
C2648 vdd.n1509 gnd 0.005391f
C2649 vdd.n1510 gnd 0.002982f
C2650 vdd.n1511 gnd 0.006847f
C2651 vdd.n1512 gnd 0.002897f
C2652 vdd.n1513 gnd 0.003067f
C2653 vdd.n1514 gnd 0.005391f
C2654 vdd.n1515 gnd 0.002897f
C2655 vdd.n1516 gnd 0.006847f
C2656 vdd.n1517 gnd 0.003067f
C2657 vdd.n1518 gnd 0.005391f
C2658 vdd.n1519 gnd 0.002897f
C2659 vdd.n1520 gnd 0.005135f
C2660 vdd.n1521 gnd 0.005151f
C2661 vdd.t37 gnd 0.01471f
C2662 vdd.n1522 gnd 0.03273f
C2663 vdd.n1523 gnd 0.170333f
C2664 vdd.n1524 gnd 0.002897f
C2665 vdd.n1525 gnd 0.003067f
C2666 vdd.n1526 gnd 0.006847f
C2667 vdd.n1527 gnd 0.006847f
C2668 vdd.n1528 gnd 0.003067f
C2669 vdd.n1529 gnd 0.002897f
C2670 vdd.n1530 gnd 0.005391f
C2671 vdd.n1531 gnd 0.005391f
C2672 vdd.n1532 gnd 0.002897f
C2673 vdd.n1533 gnd 0.003067f
C2674 vdd.n1534 gnd 0.006847f
C2675 vdd.n1535 gnd 0.006847f
C2676 vdd.n1536 gnd 0.003067f
C2677 vdd.n1537 gnd 0.002897f
C2678 vdd.n1538 gnd 0.005391f
C2679 vdd.n1539 gnd 0.005391f
C2680 vdd.n1540 gnd 0.002897f
C2681 vdd.n1541 gnd 0.003067f
C2682 vdd.n1542 gnd 0.006847f
C2683 vdd.n1543 gnd 0.006847f
C2684 vdd.n1544 gnd 0.016188f
C2685 vdd.n1545 gnd 0.002982f
C2686 vdd.n1546 gnd 0.002897f
C2687 vdd.n1547 gnd 0.013933f
C2688 vdd.n1548 gnd 0.009422f
C2689 vdd.n1549 gnd 0.110582f
C2690 vdd.n1550 gnd 0.005809f
C2691 vdd.n1551 gnd 0.005391f
C2692 vdd.n1552 gnd 0.002982f
C2693 vdd.n1553 gnd 0.006847f
C2694 vdd.n1554 gnd 0.002897f
C2695 vdd.n1555 gnd 0.003067f
C2696 vdd.n1556 gnd 0.005391f
C2697 vdd.n1557 gnd 0.002897f
C2698 vdd.n1558 gnd 0.006847f
C2699 vdd.n1559 gnd 0.003067f
C2700 vdd.n1560 gnd 0.005391f
C2701 vdd.n1561 gnd 0.002897f
C2702 vdd.n1562 gnd 0.005135f
C2703 vdd.n1563 gnd 0.005151f
C2704 vdd.t114 gnd 0.01471f
C2705 vdd.n1564 gnd 0.03273f
C2706 vdd.n1565 gnd 0.170333f
C2707 vdd.n1566 gnd 0.002897f
C2708 vdd.n1567 gnd 0.003067f
C2709 vdd.n1568 gnd 0.006847f
C2710 vdd.n1569 gnd 0.006847f
C2711 vdd.n1570 gnd 0.003067f
C2712 vdd.n1571 gnd 0.002897f
C2713 vdd.n1572 gnd 0.005391f
C2714 vdd.n1573 gnd 0.005391f
C2715 vdd.n1574 gnd 0.002897f
C2716 vdd.n1575 gnd 0.003067f
C2717 vdd.n1576 gnd 0.006847f
C2718 vdd.n1577 gnd 0.006847f
C2719 vdd.n1578 gnd 0.003067f
C2720 vdd.n1579 gnd 0.002897f
C2721 vdd.n1580 gnd 0.005391f
C2722 vdd.n1581 gnd 0.005391f
C2723 vdd.n1582 gnd 0.002897f
C2724 vdd.n1583 gnd 0.003067f
C2725 vdd.n1584 gnd 0.006847f
C2726 vdd.n1585 gnd 0.006847f
C2727 vdd.n1586 gnd 0.016188f
C2728 vdd.n1587 gnd 0.002982f
C2729 vdd.n1588 gnd 0.002897f
C2730 vdd.n1589 gnd 0.013933f
C2731 vdd.n1590 gnd 0.009728f
C2732 vdd.t26 gnd 0.03408f
C2733 vdd.t119 gnd 0.03408f
C2734 vdd.n1591 gnd 0.234219f
C2735 vdd.n1592 gnd 0.184178f
C2736 vdd.t112 gnd 0.03408f
C2737 vdd.t99 gnd 0.03408f
C2738 vdd.n1593 gnd 0.234219f
C2739 vdd.n1594 gnd 0.14863f
C2740 vdd.t70 gnd 0.03408f
C2741 vdd.t16 gnd 0.03408f
C2742 vdd.n1595 gnd 0.234219f
C2743 vdd.n1596 gnd 0.14863f
C2744 vdd.t126 gnd 0.03408f
C2745 vdd.t97 gnd 0.03408f
C2746 vdd.n1597 gnd 0.234219f
C2747 vdd.n1598 gnd 0.14863f
C2748 vdd.t94 gnd 0.03408f
C2749 vdd.t49 gnd 0.03408f
C2750 vdd.n1599 gnd 0.234219f
C2751 vdd.n1600 gnd 0.14863f
C2752 vdd.t43 gnd 0.03408f
C2753 vdd.t95 gnd 0.03408f
C2754 vdd.n1601 gnd 0.234219f
C2755 vdd.n1602 gnd 0.14863f
C2756 vdd.t85 gnd 0.03408f
C2757 vdd.t83 gnd 0.03408f
C2758 vdd.n1603 gnd 0.234219f
C2759 vdd.n1604 gnd 0.14863f
C2760 vdd.n1605 gnd 0.005809f
C2761 vdd.n1606 gnd 0.005391f
C2762 vdd.n1607 gnd 0.002982f
C2763 vdd.n1608 gnd 0.006847f
C2764 vdd.n1609 gnd 0.002897f
C2765 vdd.n1610 gnd 0.003067f
C2766 vdd.n1611 gnd 0.005391f
C2767 vdd.n1612 gnd 0.002897f
C2768 vdd.n1613 gnd 0.006847f
C2769 vdd.n1614 gnd 0.003067f
C2770 vdd.n1615 gnd 0.005391f
C2771 vdd.n1616 gnd 0.002897f
C2772 vdd.n1617 gnd 0.005135f
C2773 vdd.n1618 gnd 0.005151f
C2774 vdd.t24 gnd 0.01471f
C2775 vdd.n1619 gnd 0.03273f
C2776 vdd.n1620 gnd 0.170333f
C2777 vdd.n1621 gnd 0.002897f
C2778 vdd.n1622 gnd 0.003067f
C2779 vdd.n1623 gnd 0.006847f
C2780 vdd.n1624 gnd 0.006847f
C2781 vdd.n1625 gnd 0.003067f
C2782 vdd.n1626 gnd 0.002897f
C2783 vdd.n1627 gnd 0.005391f
C2784 vdd.n1628 gnd 0.005391f
C2785 vdd.n1629 gnd 0.002897f
C2786 vdd.n1630 gnd 0.003067f
C2787 vdd.n1631 gnd 0.006847f
C2788 vdd.n1632 gnd 0.006847f
C2789 vdd.n1633 gnd 0.003067f
C2790 vdd.n1634 gnd 0.002897f
C2791 vdd.n1635 gnd 0.005391f
C2792 vdd.n1636 gnd 0.005391f
C2793 vdd.n1637 gnd 0.002897f
C2794 vdd.n1638 gnd 0.003067f
C2795 vdd.n1639 gnd 0.006847f
C2796 vdd.n1640 gnd 0.006847f
C2797 vdd.n1641 gnd 0.016188f
C2798 vdd.n1642 gnd 0.002982f
C2799 vdd.n1643 gnd 0.002897f
C2800 vdd.n1644 gnd 0.013933f
C2801 vdd.n1645 gnd 0.009422f
C2802 vdd.n1646 gnd 0.065785f
C2803 vdd.n1647 gnd 0.237041f
C2804 vdd.n1648 gnd 0.005809f
C2805 vdd.n1649 gnd 0.005391f
C2806 vdd.n1650 gnd 0.002982f
C2807 vdd.n1651 gnd 0.006847f
C2808 vdd.n1652 gnd 0.002897f
C2809 vdd.n1653 gnd 0.003067f
C2810 vdd.n1654 gnd 0.005391f
C2811 vdd.n1655 gnd 0.002897f
C2812 vdd.n1656 gnd 0.006847f
C2813 vdd.n1657 gnd 0.003067f
C2814 vdd.n1658 gnd 0.005391f
C2815 vdd.n1659 gnd 0.002897f
C2816 vdd.n1660 gnd 0.005135f
C2817 vdd.n1661 gnd 0.005151f
C2818 vdd.t129 gnd 0.01471f
C2819 vdd.n1662 gnd 0.03273f
C2820 vdd.n1663 gnd 0.170333f
C2821 vdd.n1664 gnd 0.002897f
C2822 vdd.n1665 gnd 0.003067f
C2823 vdd.n1666 gnd 0.006847f
C2824 vdd.n1667 gnd 0.006847f
C2825 vdd.n1668 gnd 0.003067f
C2826 vdd.n1669 gnd 0.002897f
C2827 vdd.n1670 gnd 0.005391f
C2828 vdd.n1671 gnd 0.005391f
C2829 vdd.n1672 gnd 0.002897f
C2830 vdd.n1673 gnd 0.003067f
C2831 vdd.n1674 gnd 0.006847f
C2832 vdd.n1675 gnd 0.006847f
C2833 vdd.n1676 gnd 0.003067f
C2834 vdd.n1677 gnd 0.002897f
C2835 vdd.n1678 gnd 0.005391f
C2836 vdd.n1679 gnd 0.005391f
C2837 vdd.n1680 gnd 0.002897f
C2838 vdd.n1681 gnd 0.003067f
C2839 vdd.n1682 gnd 0.006847f
C2840 vdd.n1683 gnd 0.006847f
C2841 vdd.n1684 gnd 0.016188f
C2842 vdd.n1685 gnd 0.002982f
C2843 vdd.n1686 gnd 0.002897f
C2844 vdd.n1687 gnd 0.013933f
C2845 vdd.n1688 gnd 0.009728f
C2846 vdd.t41 gnd 0.03408f
C2847 vdd.t128 gnd 0.03408f
C2848 vdd.n1689 gnd 0.234219f
C2849 vdd.n1690 gnd 0.184178f
C2850 vdd.t127 gnd 0.03408f
C2851 vdd.t109 gnd 0.03408f
C2852 vdd.n1691 gnd 0.234219f
C2853 vdd.n1692 gnd 0.14863f
C2854 vdd.t86 gnd 0.03408f
C2855 vdd.t38 gnd 0.03408f
C2856 vdd.n1693 gnd 0.234219f
C2857 vdd.n1694 gnd 0.14863f
C2858 vdd.t137 gnd 0.03408f
C2859 vdd.t108 gnd 0.03408f
C2860 vdd.n1695 gnd 0.234219f
C2861 vdd.n1696 gnd 0.14863f
C2862 vdd.t104 gnd 0.03408f
C2863 vdd.t63 gnd 0.03408f
C2864 vdd.n1697 gnd 0.234219f
C2865 vdd.n1698 gnd 0.14863f
C2866 vdd.t62 gnd 0.03408f
C2867 vdd.t105 gnd 0.03408f
C2868 vdd.n1699 gnd 0.234219f
C2869 vdd.n1700 gnd 0.14863f
C2870 vdd.t92 gnd 0.03408f
C2871 vdd.t93 gnd 0.03408f
C2872 vdd.n1701 gnd 0.234219f
C2873 vdd.n1702 gnd 0.14863f
C2874 vdd.n1703 gnd 0.005809f
C2875 vdd.n1704 gnd 0.005391f
C2876 vdd.n1705 gnd 0.002982f
C2877 vdd.n1706 gnd 0.006847f
C2878 vdd.n1707 gnd 0.002897f
C2879 vdd.n1708 gnd 0.003067f
C2880 vdd.n1709 gnd 0.005391f
C2881 vdd.n1710 gnd 0.002897f
C2882 vdd.n1711 gnd 0.006847f
C2883 vdd.n1712 gnd 0.003067f
C2884 vdd.n1713 gnd 0.005391f
C2885 vdd.n1714 gnd 0.002897f
C2886 vdd.n1715 gnd 0.005135f
C2887 vdd.n1716 gnd 0.005151f
C2888 vdd.t40 gnd 0.01471f
C2889 vdd.n1717 gnd 0.03273f
C2890 vdd.n1718 gnd 0.170333f
C2891 vdd.n1719 gnd 0.002897f
C2892 vdd.n1720 gnd 0.003067f
C2893 vdd.n1721 gnd 0.006847f
C2894 vdd.n1722 gnd 0.006847f
C2895 vdd.n1723 gnd 0.003067f
C2896 vdd.n1724 gnd 0.002897f
C2897 vdd.n1725 gnd 0.005391f
C2898 vdd.n1726 gnd 0.005391f
C2899 vdd.n1727 gnd 0.002897f
C2900 vdd.n1728 gnd 0.003067f
C2901 vdd.n1729 gnd 0.006847f
C2902 vdd.n1730 gnd 0.006847f
C2903 vdd.n1731 gnd 0.003067f
C2904 vdd.n1732 gnd 0.002897f
C2905 vdd.n1733 gnd 0.005391f
C2906 vdd.n1734 gnd 0.005391f
C2907 vdd.n1735 gnd 0.002897f
C2908 vdd.n1736 gnd 0.003067f
C2909 vdd.n1737 gnd 0.006847f
C2910 vdd.n1738 gnd 0.006847f
C2911 vdd.n1739 gnd 0.016188f
C2912 vdd.n1740 gnd 0.002982f
C2913 vdd.n1741 gnd 0.002897f
C2914 vdd.n1742 gnd 0.013933f
C2915 vdd.n1743 gnd 0.009422f
C2916 vdd.n1744 gnd 0.065785f
C2917 vdd.n1745 gnd 0.265454f
C2918 vdd.n1746 gnd 2.53217f
C2919 vdd.n1747 gnd 0.624365f
C2920 vdd.n1748 gnd 0.008136f
C2921 vdd.n1749 gnd 0.010585f
C2922 vdd.n1750 gnd 0.00852f
C2923 vdd.n1751 gnd 0.010585f
C2924 vdd.n1752 gnd 0.849192f
C2925 vdd.n1753 gnd 0.010585f
C2926 vdd.n1754 gnd 0.00852f
C2927 vdd.n1755 gnd 0.010585f
C2928 vdd.n1756 gnd 0.010585f
C2929 vdd.n1757 gnd 0.010585f
C2930 vdd.n1758 gnd 0.00852f
C2931 vdd.n1759 gnd 0.010585f
C2932 vdd.t15 gnd 0.540887f
C2933 vdd.n1760 gnd 0.897872f
C2934 vdd.n1761 gnd 0.010585f
C2935 vdd.n1762 gnd 0.00852f
C2936 vdd.n1763 gnd 0.010585f
C2937 vdd.n1764 gnd 0.010585f
C2938 vdd.n1765 gnd 0.010585f
C2939 vdd.n1766 gnd 0.00852f
C2940 vdd.n1767 gnd 0.010585f
C2941 vdd.n1768 gnd 0.76265f
C2942 vdd.n1769 gnd 0.010585f
C2943 vdd.n1770 gnd 0.00852f
C2944 vdd.n1771 gnd 0.010585f
C2945 vdd.n1772 gnd 0.010585f
C2946 vdd.n1773 gnd 0.010585f
C2947 vdd.n1774 gnd 0.00852f
C2948 vdd.n1775 gnd 0.010585f
C2949 vdd.n1776 gnd 0.897872f
C2950 vdd.t98 gnd 0.540887f
C2951 vdd.n1777 gnd 0.578749f
C2952 vdd.n1778 gnd 0.010585f
C2953 vdd.n1779 gnd 0.00852f
C2954 vdd.n1780 gnd 0.010585f
C2955 vdd.n1781 gnd 0.010585f
C2956 vdd.n1782 gnd 0.010585f
C2957 vdd.n1783 gnd 0.00852f
C2958 vdd.n1784 gnd 0.010585f
C2959 vdd.n1785 gnd 0.686926f
C2960 vdd.n1786 gnd 0.010585f
C2961 vdd.n1787 gnd 0.00852f
C2962 vdd.n1788 gnd 0.010585f
C2963 vdd.n1789 gnd 0.010585f
C2964 vdd.n1790 gnd 0.010585f
C2965 vdd.n1791 gnd 0.00852f
C2966 vdd.n1792 gnd 0.010585f
C2967 vdd.n1793 gnd 0.567931f
C2968 vdd.n1794 gnd 0.870828f
C2969 vdd.n1795 gnd 0.010585f
C2970 vdd.n1796 gnd 0.00852f
C2971 vdd.n1797 gnd 0.010585f
C2972 vdd.n1798 gnd 0.010585f
C2973 vdd.n1799 gnd 0.010585f
C2974 vdd.n1800 gnd 0.00852f
C2975 vdd.n1801 gnd 0.010585f
C2976 vdd.n1802 gnd 1.05473f
C2977 vdd.n1803 gnd 0.010585f
C2978 vdd.n1804 gnd 0.00852f
C2979 vdd.n1805 gnd 0.010585f
C2980 vdd.n1806 gnd 0.010585f
C2981 vdd.n1807 gnd 0.024105f
C2982 vdd.n1808 gnd 0.010585f
C2983 vdd.n1809 gnd 0.010585f
C2984 vdd.n1810 gnd 0.00852f
C2985 vdd.n1811 gnd 0.010585f
C2986 vdd.t196 gnd 0.540887f
C2987 vdd.n1812 gnd 1.02228f
C2988 vdd.n1813 gnd 0.010585f
C2989 vdd.n1814 gnd 0.00852f
C2990 vdd.n1815 gnd 0.010585f
C2991 vdd.n1816 gnd 0.010585f
C2992 vdd.n1817 gnd 0.009103f
C2993 vdd.n1818 gnd 0.00852f
C2994 vdd.n1820 gnd 0.010585f
C2995 vdd.n1822 gnd 0.00852f
C2996 vdd.n1823 gnd 0.010585f
C2997 vdd.n1824 gnd 0.00852f
C2998 vdd.n1826 gnd 0.010585f
C2999 vdd.n1827 gnd 0.00852f
C3000 vdd.n1828 gnd 0.010585f
C3001 vdd.n1829 gnd 0.010585f
C3002 vdd.n1830 gnd 0.010585f
C3003 vdd.n1831 gnd 0.010585f
C3004 vdd.n1832 gnd 0.010585f
C3005 vdd.n1833 gnd 0.00852f
C3006 vdd.n1835 gnd 0.010585f
C3007 vdd.n1836 gnd 0.010585f
C3008 vdd.n1837 gnd 0.010585f
C3009 vdd.n1838 gnd 0.010585f
C3010 vdd.n1839 gnd 0.010585f
C3011 vdd.n1840 gnd 0.00852f
C3012 vdd.n1842 gnd 0.010585f
C3013 vdd.n1843 gnd 0.010585f
C3014 vdd.n1844 gnd 0.010585f
C3015 vdd.n1845 gnd 0.010585f
C3016 vdd.n1846 gnd 0.007114f
C3017 vdd.t214 gnd 0.130228f
C3018 vdd.t213 gnd 0.139178f
C3019 vdd.t212 gnd 0.170076f
C3020 vdd.n1847 gnd 0.218013f
C3021 vdd.n1848 gnd 0.18317f
C3022 vdd.n1850 gnd 0.010585f
C3023 vdd.n1851 gnd 0.010585f
C3024 vdd.n1852 gnd 0.00852f
C3025 vdd.n1853 gnd 0.010585f
C3026 vdd.n1855 gnd 0.010585f
C3027 vdd.n1856 gnd 0.010585f
C3028 vdd.n1857 gnd 0.010585f
C3029 vdd.n1858 gnd 0.010585f
C3030 vdd.n1859 gnd 0.00852f
C3031 vdd.n1861 gnd 0.010585f
C3032 vdd.n1862 gnd 0.010585f
C3033 vdd.n1863 gnd 0.010585f
C3034 vdd.n1864 gnd 0.010585f
C3035 vdd.n1865 gnd 0.010585f
C3036 vdd.n1866 gnd 0.00852f
C3037 vdd.n1868 gnd 0.010585f
C3038 vdd.n1869 gnd 0.010585f
C3039 vdd.n1870 gnd 0.010585f
C3040 vdd.n1871 gnd 0.010585f
C3041 vdd.n1872 gnd 0.010585f
C3042 vdd.n1873 gnd 0.00852f
C3043 vdd.n1875 gnd 0.010585f
C3044 vdd.n1876 gnd 0.010585f
C3045 vdd.n1877 gnd 0.010585f
C3046 vdd.n1878 gnd 0.010585f
C3047 vdd.n1879 gnd 0.010585f
C3048 vdd.n1880 gnd 0.00852f
C3049 vdd.n1882 gnd 0.010585f
C3050 vdd.n1883 gnd 0.010585f
C3051 vdd.n1884 gnd 0.010585f
C3052 vdd.n1885 gnd 0.010585f
C3053 vdd.n1886 gnd 0.008435f
C3054 vdd.t211 gnd 0.130228f
C3055 vdd.t210 gnd 0.139178f
C3056 vdd.t209 gnd 0.170076f
C3057 vdd.n1887 gnd 0.218013f
C3058 vdd.n1888 gnd 0.18317f
C3059 vdd.n1890 gnd 0.010585f
C3060 vdd.n1891 gnd 0.010585f
C3061 vdd.n1892 gnd 0.00852f
C3062 vdd.n1893 gnd 0.010585f
C3063 vdd.n1895 gnd 0.010585f
C3064 vdd.n1896 gnd 0.010585f
C3065 vdd.n1897 gnd 0.010585f
C3066 vdd.n1898 gnd 0.010585f
C3067 vdd.n1899 gnd 0.00852f
C3068 vdd.n1901 gnd 0.010585f
C3069 vdd.n1902 gnd 0.010585f
C3070 vdd.n1903 gnd 0.010585f
C3071 vdd.n1904 gnd 0.010585f
C3072 vdd.n1905 gnd 0.010585f
C3073 vdd.n1906 gnd 0.00852f
C3074 vdd.n1908 gnd 0.010585f
C3075 vdd.n1909 gnd 0.010585f
C3076 vdd.n1910 gnd 0.010585f
C3077 vdd.n1911 gnd 0.010585f
C3078 vdd.n1912 gnd 0.010585f
C3079 vdd.n1913 gnd 0.010585f
C3080 vdd.n1914 gnd 0.00852f
C3081 vdd.n1916 gnd 0.010585f
C3082 vdd.n1918 gnd 0.010585f
C3083 vdd.n1919 gnd 0.00852f
C3084 vdd.n1920 gnd 0.00852f
C3085 vdd.n1921 gnd 0.010585f
C3086 vdd.n1923 gnd 0.010585f
C3087 vdd.n1924 gnd 0.00852f
C3088 vdd.n1925 gnd 0.00852f
C3089 vdd.n1926 gnd 0.010585f
C3090 vdd.n1928 gnd 0.010585f
C3091 vdd.n1929 gnd 0.010585f
C3092 vdd.n1930 gnd 0.00852f
C3093 vdd.n1931 gnd 0.00852f
C3094 vdd.n1932 gnd 0.00852f
C3095 vdd.n1933 gnd 0.010585f
C3096 vdd.n1935 gnd 0.010585f
C3097 vdd.n1936 gnd 0.010585f
C3098 vdd.n1937 gnd 0.00852f
C3099 vdd.n1938 gnd 0.00852f
C3100 vdd.n1939 gnd 0.00852f
C3101 vdd.n1940 gnd 0.010585f
C3102 vdd.n1942 gnd 0.010585f
C3103 vdd.n1943 gnd 0.010585f
C3104 vdd.n1944 gnd 0.00852f
C3105 vdd.n1945 gnd 0.00852f
C3106 vdd.n1946 gnd 0.00852f
C3107 vdd.n1947 gnd 0.010585f
C3108 vdd.n1949 gnd 0.010585f
C3109 vdd.n1950 gnd 0.010585f
C3110 vdd.n1951 gnd 0.00852f
C3111 vdd.n1952 gnd 0.010585f
C3112 vdd.n1953 gnd 0.010585f
C3113 vdd.n1954 gnd 0.010585f
C3114 vdd.n1955 gnd 0.017381f
C3115 vdd.n1956 gnd 0.005794f
C3116 vdd.n1957 gnd 0.00852f
C3117 vdd.n1958 gnd 0.010585f
C3118 vdd.n1960 gnd 0.010585f
C3119 vdd.n1961 gnd 0.010585f
C3120 vdd.n1962 gnd 0.00852f
C3121 vdd.n1963 gnd 0.00852f
C3122 vdd.n1964 gnd 0.00852f
C3123 vdd.n1965 gnd 0.010585f
C3124 vdd.n1967 gnd 0.010585f
C3125 vdd.n1968 gnd 0.010585f
C3126 vdd.n1969 gnd 0.00852f
C3127 vdd.n1970 gnd 0.00852f
C3128 vdd.n1971 gnd 0.00852f
C3129 vdd.n1972 gnd 0.010585f
C3130 vdd.n1974 gnd 0.010585f
C3131 vdd.n1975 gnd 0.010585f
C3132 vdd.n1976 gnd 0.00852f
C3133 vdd.n1977 gnd 0.00852f
C3134 vdd.n1978 gnd 0.00852f
C3135 vdd.n1979 gnd 0.010585f
C3136 vdd.n1981 gnd 0.010585f
C3137 vdd.n1982 gnd 0.010585f
C3138 vdd.n1983 gnd 0.00852f
C3139 vdd.n1984 gnd 0.00852f
C3140 vdd.n1985 gnd 0.00852f
C3141 vdd.n1986 gnd 0.010585f
C3142 vdd.n1988 gnd 0.010585f
C3143 vdd.n1989 gnd 0.010585f
C3144 vdd.n1990 gnd 0.00852f
C3145 vdd.n1991 gnd 0.010585f
C3146 vdd.n1992 gnd 0.010585f
C3147 vdd.n1993 gnd 0.010585f
C3148 vdd.n1994 gnd 0.017381f
C3149 vdd.n1995 gnd 0.007114f
C3150 vdd.n1996 gnd 0.00852f
C3151 vdd.n1997 gnd 0.010585f
C3152 vdd.n1999 gnd 0.010585f
C3153 vdd.n2000 gnd 0.010585f
C3154 vdd.n2001 gnd 0.00852f
C3155 vdd.n2002 gnd 0.00852f
C3156 vdd.n2003 gnd 0.00852f
C3157 vdd.n2004 gnd 0.010585f
C3158 vdd.n2006 gnd 0.010585f
C3159 vdd.n2007 gnd 0.010585f
C3160 vdd.n2008 gnd 0.00852f
C3161 vdd.n2009 gnd 0.00852f
C3162 vdd.n2010 gnd 0.00852f
C3163 vdd.n2011 gnd 0.010585f
C3164 vdd.n2013 gnd 0.010585f
C3165 vdd.n2014 gnd 0.010585f
C3166 vdd.n2016 gnd 0.010585f
C3167 vdd.n2017 gnd 0.00852f
C3168 vdd.n2018 gnd 0.006775f
C3169 vdd.n2019 gnd 0.007198f
C3170 vdd.n2020 gnd 0.007198f
C3171 vdd.n2021 gnd 0.007198f
C3172 vdd.n2022 gnd 0.007198f
C3173 vdd.n2023 gnd 0.007198f
C3174 vdd.n2024 gnd 0.007198f
C3175 vdd.n2025 gnd 0.007198f
C3176 vdd.n2026 gnd 0.007198f
C3177 vdd.n2028 gnd 0.007198f
C3178 vdd.n2029 gnd 0.007198f
C3179 vdd.n2030 gnd 0.007198f
C3180 vdd.n2031 gnd 0.007198f
C3181 vdd.n2032 gnd 0.007198f
C3182 vdd.n2034 gnd 0.007198f
C3183 vdd.n2036 gnd 0.007198f
C3184 vdd.n2037 gnd 0.007198f
C3185 vdd.n2038 gnd 0.007198f
C3186 vdd.n2039 gnd 0.007198f
C3187 vdd.n2040 gnd 0.007198f
C3188 vdd.n2042 gnd 0.007198f
C3189 vdd.n2044 gnd 0.007198f
C3190 vdd.n2045 gnd 0.007198f
C3191 vdd.n2046 gnd 0.007198f
C3192 vdd.n2047 gnd 0.007198f
C3193 vdd.n2048 gnd 0.007198f
C3194 vdd.n2050 gnd 0.007198f
C3195 vdd.n2052 gnd 0.007198f
C3196 vdd.n2053 gnd 0.007198f
C3197 vdd.n2054 gnd 0.007198f
C3198 vdd.n2055 gnd 0.007198f
C3199 vdd.n2056 gnd 0.007198f
C3200 vdd.n2058 gnd 0.007198f
C3201 vdd.n2059 gnd 0.007198f
C3202 vdd.n2060 gnd 0.007198f
C3203 vdd.n2061 gnd 0.007198f
C3204 vdd.n2062 gnd 0.007198f
C3205 vdd.n2063 gnd 0.007198f
C3206 vdd.n2064 gnd 0.007198f
C3207 vdd.n2065 gnd 0.007198f
C3208 vdd.n2066 gnd 0.00524f
C3209 vdd.n2067 gnd 0.007198f
C3210 vdd.t254 gnd 0.290872f
C3211 vdd.t255 gnd 0.297744f
C3212 vdd.t253 gnd 0.189892f
C3213 vdd.n2068 gnd 0.102626f
C3214 vdd.n2069 gnd 0.058213f
C3215 vdd.n2070 gnd 0.010287f
C3216 vdd.n2071 gnd 0.007198f
C3217 vdd.n2072 gnd 0.007198f
C3218 vdd.n2073 gnd 0.438118f
C3219 vdd.n2074 gnd 0.007198f
C3220 vdd.n2075 gnd 0.007198f
C3221 vdd.n2076 gnd 0.007198f
C3222 vdd.n2077 gnd 0.007198f
C3223 vdd.n2078 gnd 0.007198f
C3224 vdd.n2079 gnd 0.007198f
C3225 vdd.n2080 gnd 0.007198f
C3226 vdd.n2081 gnd 0.007198f
C3227 vdd.n2082 gnd 0.007198f
C3228 vdd.n2083 gnd 0.007198f
C3229 vdd.n2084 gnd 0.007198f
C3230 vdd.n2085 gnd 0.007198f
C3231 vdd.n2086 gnd 0.007198f
C3232 vdd.n2087 gnd 0.007198f
C3233 vdd.n2088 gnd 0.007198f
C3234 vdd.n2089 gnd 0.007198f
C3235 vdd.n2090 gnd 0.007198f
C3236 vdd.n2091 gnd 0.007198f
C3237 vdd.n2092 gnd 0.007198f
C3238 vdd.n2093 gnd 0.007198f
C3239 vdd.t232 gnd 0.290872f
C3240 vdd.t233 gnd 0.297744f
C3241 vdd.t230 gnd 0.189892f
C3242 vdd.n2094 gnd 0.102626f
C3243 vdd.n2095 gnd 0.058213f
C3244 vdd.n2096 gnd 0.007198f
C3245 vdd.n2097 gnd 0.007198f
C3246 vdd.n2098 gnd 0.007198f
C3247 vdd.n2099 gnd 0.007198f
C3248 vdd.n2100 gnd 0.007198f
C3249 vdd.n2101 gnd 0.007198f
C3250 vdd.n2103 gnd 0.007198f
C3251 vdd.n2104 gnd 0.007198f
C3252 vdd.n2105 gnd 0.007198f
C3253 vdd.n2106 gnd 0.007198f
C3254 vdd.n2108 gnd 0.007198f
C3255 vdd.n2110 gnd 0.007198f
C3256 vdd.n2111 gnd 0.007198f
C3257 vdd.n2112 gnd 0.007198f
C3258 vdd.n2113 gnd 0.007198f
C3259 vdd.n2114 gnd 0.007198f
C3260 vdd.n2116 gnd 0.007198f
C3261 vdd.n2118 gnd 0.007198f
C3262 vdd.n2119 gnd 0.007198f
C3263 vdd.n2120 gnd 0.007198f
C3264 vdd.n2121 gnd 0.007198f
C3265 vdd.n2122 gnd 0.007198f
C3266 vdd.n2124 gnd 0.007198f
C3267 vdd.n2126 gnd 0.007198f
C3268 vdd.n2127 gnd 0.007198f
C3269 vdd.n2128 gnd 0.00524f
C3270 vdd.n2129 gnd 0.010287f
C3271 vdd.n2130 gnd 0.005557f
C3272 vdd.n2131 gnd 0.007198f
C3273 vdd.n2133 gnd 0.007198f
C3274 vdd.n2134 gnd 0.01708f
C3275 vdd.n2135 gnd 0.01708f
C3276 vdd.n2136 gnd 0.015947f
C3277 vdd.n2137 gnd 0.007198f
C3278 vdd.n2138 gnd 0.007198f
C3279 vdd.n2139 gnd 0.007198f
C3280 vdd.n2140 gnd 0.007198f
C3281 vdd.n2141 gnd 0.007198f
C3282 vdd.n2142 gnd 0.007198f
C3283 vdd.n2143 gnd 0.007198f
C3284 vdd.n2144 gnd 0.007198f
C3285 vdd.n2145 gnd 0.007198f
C3286 vdd.n2146 gnd 0.007198f
C3287 vdd.n2147 gnd 0.007198f
C3288 vdd.n2148 gnd 0.007198f
C3289 vdd.n2149 gnd 0.007198f
C3290 vdd.n2150 gnd 0.007198f
C3291 vdd.n2151 gnd 0.007198f
C3292 vdd.n2152 gnd 0.007198f
C3293 vdd.n2153 gnd 0.007198f
C3294 vdd.n2154 gnd 0.007198f
C3295 vdd.n2155 gnd 0.007198f
C3296 vdd.n2156 gnd 0.007198f
C3297 vdd.n2157 gnd 0.007198f
C3298 vdd.n2158 gnd 0.007198f
C3299 vdd.n2159 gnd 0.007198f
C3300 vdd.n2160 gnd 0.007198f
C3301 vdd.n2161 gnd 0.007198f
C3302 vdd.n2162 gnd 0.007198f
C3303 vdd.n2163 gnd 0.007198f
C3304 vdd.n2164 gnd 0.007198f
C3305 vdd.n2165 gnd 0.007198f
C3306 vdd.n2166 gnd 0.007198f
C3307 vdd.n2167 gnd 0.007198f
C3308 vdd.n2168 gnd 0.007198f
C3309 vdd.n2169 gnd 0.007198f
C3310 vdd.n2170 gnd 0.007198f
C3311 vdd.n2171 gnd 0.007198f
C3312 vdd.n2172 gnd 0.007198f
C3313 vdd.n2173 gnd 0.007198f
C3314 vdd.n2174 gnd 0.232581f
C3315 vdd.n2175 gnd 0.007198f
C3316 vdd.n2176 gnd 0.007198f
C3317 vdd.n2177 gnd 0.007198f
C3318 vdd.n2178 gnd 0.007198f
C3319 vdd.n2179 gnd 0.007198f
C3320 vdd.n2180 gnd 0.007198f
C3321 vdd.n2181 gnd 0.007198f
C3322 vdd.n2182 gnd 0.007198f
C3323 vdd.n2183 gnd 0.007198f
C3324 vdd.n2184 gnd 0.007198f
C3325 vdd.n2185 gnd 0.007198f
C3326 vdd.n2186 gnd 0.007198f
C3327 vdd.n2187 gnd 0.007198f
C3328 vdd.n2188 gnd 0.007198f
C3329 vdd.n2189 gnd 0.007198f
C3330 vdd.n2190 gnd 0.007198f
C3331 vdd.n2191 gnd 0.007198f
C3332 vdd.n2192 gnd 0.007198f
C3333 vdd.n2193 gnd 0.007198f
C3334 vdd.n2194 gnd 0.007198f
C3335 vdd.n2195 gnd 0.015947f
C3336 vdd.n2197 gnd 0.01708f
C3337 vdd.n2198 gnd 0.01708f
C3338 vdd.n2199 gnd 0.007198f
C3339 vdd.n2200 gnd 0.005557f
C3340 vdd.n2201 gnd 0.007198f
C3341 vdd.n2203 gnd 0.007198f
C3342 vdd.n2205 gnd 0.007198f
C3343 vdd.n2206 gnd 0.007198f
C3344 vdd.n2207 gnd 0.007198f
C3345 vdd.n2208 gnd 0.007198f
C3346 vdd.n2209 gnd 0.007198f
C3347 vdd.n2211 gnd 0.007198f
C3348 vdd.n2213 gnd 0.007198f
C3349 vdd.n2214 gnd 0.007198f
C3350 vdd.n2215 gnd 0.007198f
C3351 vdd.n2216 gnd 0.007198f
C3352 vdd.n2217 gnd 0.007198f
C3353 vdd.n2219 gnd 0.007198f
C3354 vdd.n2221 gnd 0.007198f
C3355 vdd.n2222 gnd 0.007198f
C3356 vdd.n2223 gnd 0.007198f
C3357 vdd.n2224 gnd 0.007198f
C3358 vdd.n2225 gnd 0.007198f
C3359 vdd.n2227 gnd 0.007198f
C3360 vdd.n2229 gnd 0.007198f
C3361 vdd.n2230 gnd 0.007198f
C3362 vdd.n2231 gnd 0.02147f
C3363 vdd.n2232 gnd 0.63647f
C3364 vdd.n2234 gnd 0.00852f
C3365 vdd.n2235 gnd 0.00852f
C3366 vdd.n2236 gnd 0.010585f
C3367 vdd.n2238 gnd 0.010585f
C3368 vdd.n2239 gnd 0.010585f
C3369 vdd.n2240 gnd 0.00852f
C3370 vdd.n2241 gnd 0.007072f
C3371 vdd.n2242 gnd 0.02427f
C3372 vdd.n2243 gnd 0.024105f
C3373 vdd.n2244 gnd 0.007072f
C3374 vdd.n2245 gnd 0.024105f
C3375 vdd.n2246 gnd 1.42794f
C3376 vdd.n2247 gnd 0.024105f
C3377 vdd.n2248 gnd 0.02427f
C3378 vdd.n2249 gnd 0.004047f
C3379 vdd.t198 gnd 0.130228f
C3380 vdd.t197 gnd 0.139178f
C3381 vdd.t195 gnd 0.170076f
C3382 vdd.n2250 gnd 0.218013f
C3383 vdd.n2251 gnd 0.18317f
C3384 vdd.n2252 gnd 0.013121f
C3385 vdd.n2253 gnd 0.004473f
C3386 vdd.n2254 gnd 0.009103f
C3387 vdd.n2255 gnd 0.63647f
C3388 vdd.n2256 gnd 0.02147f
C3389 vdd.n2257 gnd 0.007198f
C3390 vdd.n2258 gnd 0.007198f
C3391 vdd.n2259 gnd 0.007198f
C3392 vdd.n2261 gnd 0.007198f
C3393 vdd.n2263 gnd 0.007198f
C3394 vdd.n2264 gnd 0.007198f
C3395 vdd.n2265 gnd 0.007198f
C3396 vdd.n2266 gnd 0.007198f
C3397 vdd.n2267 gnd 0.007198f
C3398 vdd.n2269 gnd 0.007198f
C3399 vdd.n2271 gnd 0.007198f
C3400 vdd.n2272 gnd 0.007198f
C3401 vdd.n2273 gnd 0.007198f
C3402 vdd.n2274 gnd 0.007198f
C3403 vdd.n2275 gnd 0.007198f
C3404 vdd.n2277 gnd 0.007198f
C3405 vdd.n2279 gnd 0.007198f
C3406 vdd.n2280 gnd 0.007198f
C3407 vdd.n2281 gnd 0.007198f
C3408 vdd.n2282 gnd 0.007198f
C3409 vdd.n2283 gnd 0.007198f
C3410 vdd.n2285 gnd 0.007198f
C3411 vdd.n2287 gnd 0.007198f
C3412 vdd.n2288 gnd 0.007198f
C3413 vdd.n2289 gnd 0.01708f
C3414 vdd.n2290 gnd 0.015947f
C3415 vdd.n2291 gnd 0.015947f
C3416 vdd.n2292 gnd 1.06014f
C3417 vdd.n2293 gnd 0.015947f
C3418 vdd.n2294 gnd 0.015947f
C3419 vdd.n2295 gnd 0.007198f
C3420 vdd.n2296 gnd 0.007198f
C3421 vdd.n2297 gnd 0.007198f
C3422 vdd.n2298 gnd 0.459754f
C3423 vdd.n2299 gnd 0.007198f
C3424 vdd.n2300 gnd 0.007198f
C3425 vdd.n2301 gnd 0.007198f
C3426 vdd.n2302 gnd 0.007198f
C3427 vdd.n2303 gnd 0.007198f
C3428 vdd.n2304 gnd 0.735606f
C3429 vdd.n2305 gnd 0.007198f
C3430 vdd.n2306 gnd 0.007198f
C3431 vdd.n2307 gnd 0.007198f
C3432 vdd.n2308 gnd 0.007198f
C3433 vdd.n2309 gnd 0.007198f
C3434 vdd.n2310 gnd 0.735606f
C3435 vdd.n2311 gnd 0.007198f
C3436 vdd.n2312 gnd 0.007198f
C3437 vdd.n2313 gnd 0.006351f
C3438 vdd.n2314 gnd 0.020852f
C3439 vdd.n2315 gnd 0.004446f
C3440 vdd.n2316 gnd 0.007198f
C3441 vdd.n2317 gnd 0.405665f
C3442 vdd.n2318 gnd 0.007198f
C3443 vdd.n2319 gnd 0.007198f
C3444 vdd.n2320 gnd 0.007198f
C3445 vdd.n2321 gnd 0.007198f
C3446 vdd.n2322 gnd 0.007198f
C3447 vdd.n2323 gnd 0.492207f
C3448 vdd.n2324 gnd 0.007198f
C3449 vdd.n2325 gnd 0.007198f
C3450 vdd.n2326 gnd 0.007198f
C3451 vdd.n2327 gnd 0.007198f
C3452 vdd.n2328 gnd 0.007198f
C3453 vdd.n2329 gnd 0.654473f
C3454 vdd.n2330 gnd 0.007198f
C3455 vdd.n2331 gnd 0.007198f
C3456 vdd.n2332 gnd 0.007198f
C3457 vdd.n2333 gnd 0.007198f
C3458 vdd.n2334 gnd 0.007198f
C3459 vdd.n2335 gnd 0.584158f
C3460 vdd.n2336 gnd 0.007198f
C3461 vdd.n2337 gnd 0.007198f
C3462 vdd.n2338 gnd 0.007198f
C3463 vdd.n2339 gnd 0.007198f
C3464 vdd.n2340 gnd 0.007198f
C3465 vdd.n2341 gnd 0.421892f
C3466 vdd.n2342 gnd 0.007198f
C3467 vdd.n2343 gnd 0.007198f
C3468 vdd.n2344 gnd 0.007198f
C3469 vdd.n2345 gnd 0.007198f
C3470 vdd.n2346 gnd 0.007198f
C3471 vdd.n2347 gnd 0.232581f
C3472 vdd.n2348 gnd 0.007198f
C3473 vdd.n2349 gnd 0.007198f
C3474 vdd.n2350 gnd 0.007198f
C3475 vdd.n2351 gnd 0.007198f
C3476 vdd.n2352 gnd 0.007198f
C3477 vdd.n2353 gnd 0.405665f
C3478 vdd.n2354 gnd 0.007198f
C3479 vdd.n2355 gnd 0.007198f
C3480 vdd.n2356 gnd 0.007198f
C3481 vdd.n2357 gnd 0.007198f
C3482 vdd.n2358 gnd 0.007198f
C3483 vdd.n2359 gnd 0.735606f
C3484 vdd.n2360 gnd 0.007198f
C3485 vdd.n2361 gnd 0.007198f
C3486 vdd.n2362 gnd 0.007198f
C3487 vdd.n2363 gnd 0.007198f
C3488 vdd.n2364 gnd 0.007198f
C3489 vdd.n2365 gnd 0.007198f
C3490 vdd.n2366 gnd 0.007198f
C3491 vdd.n2367 gnd 0.57334f
C3492 vdd.n2368 gnd 0.007198f
C3493 vdd.n2369 gnd 0.007198f
C3494 vdd.n2370 gnd 0.007198f
C3495 vdd.n2371 gnd 0.007198f
C3496 vdd.n2372 gnd 0.007198f
C3497 vdd.n2373 gnd 0.007198f
C3498 vdd.n2374 gnd 0.459754f
C3499 vdd.n2375 gnd 0.007198f
C3500 vdd.n2376 gnd 0.007198f
C3501 vdd.n2377 gnd 0.007198f
C3502 vdd.n2378 gnd 0.016823f
C3503 vdd.n2379 gnd 0.016203f
C3504 vdd.n2380 gnd 0.007198f
C3505 vdd.n2381 gnd 0.007198f
C3506 vdd.n2382 gnd 0.005557f
C3507 vdd.n2383 gnd 0.007198f
C3508 vdd.n2384 gnd 0.007198f
C3509 vdd.n2385 gnd 0.00524f
C3510 vdd.n2386 gnd 0.007198f
C3511 vdd.n2387 gnd 0.007198f
C3512 vdd.n2388 gnd 0.007198f
C3513 vdd.n2389 gnd 0.007198f
C3514 vdd.n2390 gnd 0.007198f
C3515 vdd.n2391 gnd 0.007198f
C3516 vdd.n2392 gnd 0.007198f
C3517 vdd.n2393 gnd 0.007198f
C3518 vdd.n2394 gnd 0.007198f
C3519 vdd.n2395 gnd 0.007198f
C3520 vdd.n2396 gnd 0.007198f
C3521 vdd.n2397 gnd 0.007198f
C3522 vdd.n2398 gnd 0.007198f
C3523 vdd.n2399 gnd 0.007198f
C3524 vdd.n2400 gnd 0.007198f
C3525 vdd.n2401 gnd 0.007198f
C3526 vdd.n2402 gnd 0.007198f
C3527 vdd.n2403 gnd 0.007198f
C3528 vdd.n2404 gnd 0.007198f
C3529 vdd.n2405 gnd 0.007198f
C3530 vdd.n2406 gnd 0.007198f
C3531 vdd.n2407 gnd 0.007198f
C3532 vdd.n2408 gnd 0.007198f
C3533 vdd.n2409 gnd 0.007198f
C3534 vdd.n2410 gnd 0.007198f
C3535 vdd.n2411 gnd 0.007198f
C3536 vdd.n2412 gnd 0.007198f
C3537 vdd.n2413 gnd 0.007198f
C3538 vdd.n2414 gnd 0.007198f
C3539 vdd.n2415 gnd 0.007198f
C3540 vdd.n2416 gnd 0.007198f
C3541 vdd.n2417 gnd 0.007198f
C3542 vdd.n2418 gnd 0.007198f
C3543 vdd.n2419 gnd 0.007198f
C3544 vdd.n2420 gnd 0.007198f
C3545 vdd.n2421 gnd 0.007198f
C3546 vdd.n2422 gnd 0.007198f
C3547 vdd.n2423 gnd 0.007198f
C3548 vdd.n2424 gnd 0.007198f
C3549 vdd.n2425 gnd 0.007198f
C3550 vdd.n2426 gnd 0.007198f
C3551 vdd.n2427 gnd 0.007198f
C3552 vdd.n2428 gnd 0.007198f
C3553 vdd.n2429 gnd 0.007198f
C3554 vdd.n2430 gnd 0.007198f
C3555 vdd.n2431 gnd 0.007198f
C3556 vdd.n2432 gnd 0.007198f
C3557 vdd.n2433 gnd 0.007198f
C3558 vdd.n2434 gnd 0.007198f
C3559 vdd.n2435 gnd 0.007198f
C3560 vdd.n2436 gnd 0.007198f
C3561 vdd.n2437 gnd 0.007198f
C3562 vdd.n2438 gnd 0.007198f
C3563 vdd.n2439 gnd 0.007198f
C3564 vdd.n2440 gnd 0.007198f
C3565 vdd.n2441 gnd 0.007198f
C3566 vdd.n2442 gnd 0.007198f
C3567 vdd.n2443 gnd 0.007198f
C3568 vdd.n2444 gnd 0.007198f
C3569 vdd.n2445 gnd 0.007198f
C3570 vdd.n2446 gnd 0.01708f
C3571 vdd.n2447 gnd 0.015947f
C3572 vdd.n2448 gnd 0.015947f
C3573 vdd.n2449 gnd 0.897872f
C3574 vdd.n2450 gnd 0.015947f
C3575 vdd.n2451 gnd 0.01708f
C3576 vdd.n2452 gnd 0.016203f
C3577 vdd.n2453 gnd 0.007198f
C3578 vdd.n2454 gnd 0.007198f
C3579 vdd.n2455 gnd 0.007198f
C3580 vdd.n2456 gnd 0.005557f
C3581 vdd.n2457 gnd 0.010287f
C3582 vdd.n2458 gnd 0.00524f
C3583 vdd.n2459 gnd 0.007198f
C3584 vdd.n2460 gnd 0.007198f
C3585 vdd.n2461 gnd 0.007198f
C3586 vdd.n2462 gnd 0.007198f
C3587 vdd.n2463 gnd 0.007198f
C3588 vdd.n2464 gnd 0.007198f
C3589 vdd.n2465 gnd 0.007198f
C3590 vdd.n2466 gnd 0.007198f
C3591 vdd.n2467 gnd 0.007198f
C3592 vdd.n2468 gnd 0.007198f
C3593 vdd.n2469 gnd 0.007198f
C3594 vdd.n2470 gnd 0.007198f
C3595 vdd.n2471 gnd 0.007198f
C3596 vdd.n2472 gnd 0.007198f
C3597 vdd.n2473 gnd 0.007198f
C3598 vdd.n2474 gnd 0.007198f
C3599 vdd.n2475 gnd 0.007198f
C3600 vdd.n2476 gnd 0.007198f
C3601 vdd.n2477 gnd 0.007198f
C3602 vdd.n2478 gnd 0.007198f
C3603 vdd.n2479 gnd 0.007198f
C3604 vdd.n2480 gnd 0.007198f
C3605 vdd.n2481 gnd 0.007198f
C3606 vdd.n2482 gnd 0.007198f
C3607 vdd.n2483 gnd 0.007198f
C3608 vdd.n2484 gnd 0.007198f
C3609 vdd.n2485 gnd 0.007198f
C3610 vdd.n2486 gnd 0.007198f
C3611 vdd.n2487 gnd 0.007198f
C3612 vdd.n2488 gnd 0.007198f
C3613 vdd.n2489 gnd 0.007198f
C3614 vdd.n2490 gnd 0.007198f
C3615 vdd.n2491 gnd 0.007198f
C3616 vdd.n2492 gnd 0.007198f
C3617 vdd.n2493 gnd 0.007198f
C3618 vdd.n2494 gnd 0.007198f
C3619 vdd.n2495 gnd 0.007198f
C3620 vdd.n2496 gnd 0.007198f
C3621 vdd.n2497 gnd 0.007198f
C3622 vdd.n2498 gnd 0.007198f
C3623 vdd.n2499 gnd 0.007198f
C3624 vdd.n2500 gnd 0.007198f
C3625 vdd.n2501 gnd 0.007198f
C3626 vdd.n2502 gnd 0.007198f
C3627 vdd.n2503 gnd 0.007198f
C3628 vdd.n2504 gnd 0.007198f
C3629 vdd.n2505 gnd 0.007198f
C3630 vdd.n2506 gnd 0.007198f
C3631 vdd.n2507 gnd 0.007198f
C3632 vdd.n2508 gnd 0.007198f
C3633 vdd.n2509 gnd 0.007198f
C3634 vdd.n2510 gnd 0.007198f
C3635 vdd.n2511 gnd 0.007198f
C3636 vdd.n2512 gnd 0.007198f
C3637 vdd.n2513 gnd 0.007198f
C3638 vdd.n2514 gnd 0.007198f
C3639 vdd.n2515 gnd 0.007198f
C3640 vdd.n2516 gnd 0.007198f
C3641 vdd.n2517 gnd 0.007198f
C3642 vdd.n2518 gnd 0.007198f
C3643 vdd.n2519 gnd 0.01708f
C3644 vdd.n2520 gnd 0.01708f
C3645 vdd.n2521 gnd 0.897872f
C3646 vdd.t157 gnd 3.19123f
C3647 vdd.t160 gnd 3.19123f
C3648 vdd.n2554 gnd 0.01708f
C3649 vdd.n2555 gnd 0.007198f
C3650 vdd.t225 gnd 0.290872f
C3651 vdd.t226 gnd 0.297744f
C3652 vdd.t223 gnd 0.189892f
C3653 vdd.n2556 gnd 0.102626f
C3654 vdd.n2557 gnd 0.058213f
C3655 vdd.n2558 gnd 0.007198f
C3656 vdd.t239 gnd 0.290872f
C3657 vdd.t240 gnd 0.297744f
C3658 vdd.t238 gnd 0.189892f
C3659 vdd.n2559 gnd 0.102626f
C3660 vdd.n2560 gnd 0.058213f
C3661 vdd.n2561 gnd 0.010287f
C3662 vdd.n2562 gnd 0.007198f
C3663 vdd.n2563 gnd 0.007198f
C3664 vdd.n2564 gnd 0.007198f
C3665 vdd.n2565 gnd 0.007198f
C3666 vdd.n2566 gnd 0.007198f
C3667 vdd.n2567 gnd 0.007198f
C3668 vdd.n2568 gnd 0.007198f
C3669 vdd.n2569 gnd 0.007198f
C3670 vdd.n2570 gnd 0.007198f
C3671 vdd.n2571 gnd 0.007198f
C3672 vdd.n2572 gnd 0.007198f
C3673 vdd.n2573 gnd 0.007198f
C3674 vdd.n2574 gnd 0.007198f
C3675 vdd.n2575 gnd 0.007198f
C3676 vdd.n2576 gnd 0.007198f
C3677 vdd.n2577 gnd 0.007198f
C3678 vdd.n2578 gnd 0.007198f
C3679 vdd.n2579 gnd 0.007198f
C3680 vdd.n2580 gnd 0.007198f
C3681 vdd.n2581 gnd 0.007198f
C3682 vdd.n2582 gnd 0.007198f
C3683 vdd.n2583 gnd 0.007198f
C3684 vdd.n2584 gnd 0.007198f
C3685 vdd.n2585 gnd 0.007198f
C3686 vdd.n2586 gnd 0.007198f
C3687 vdd.n2587 gnd 0.007198f
C3688 vdd.n2588 gnd 0.007198f
C3689 vdd.n2589 gnd 0.007198f
C3690 vdd.n2590 gnd 0.007198f
C3691 vdd.n2591 gnd 0.007198f
C3692 vdd.n2592 gnd 0.007198f
C3693 vdd.n2593 gnd 0.007198f
C3694 vdd.n2594 gnd 0.007198f
C3695 vdd.n2595 gnd 0.007198f
C3696 vdd.n2596 gnd 0.007198f
C3697 vdd.n2597 gnd 0.007198f
C3698 vdd.n2598 gnd 0.007198f
C3699 vdd.n2599 gnd 0.007198f
C3700 vdd.n2600 gnd 0.007198f
C3701 vdd.n2601 gnd 0.007198f
C3702 vdd.n2602 gnd 0.007198f
C3703 vdd.n2603 gnd 0.007198f
C3704 vdd.n2604 gnd 0.007198f
C3705 vdd.n2605 gnd 0.007198f
C3706 vdd.n2606 gnd 0.007198f
C3707 vdd.n2607 gnd 0.007198f
C3708 vdd.n2608 gnd 0.007198f
C3709 vdd.n2609 gnd 0.007198f
C3710 vdd.n2610 gnd 0.007198f
C3711 vdd.n2611 gnd 0.007198f
C3712 vdd.n2612 gnd 0.007198f
C3713 vdd.n2613 gnd 0.007198f
C3714 vdd.n2614 gnd 0.007198f
C3715 vdd.n2615 gnd 0.007198f
C3716 vdd.n2616 gnd 0.007198f
C3717 vdd.n2617 gnd 0.007198f
C3718 vdd.n2618 gnd 0.00524f
C3719 vdd.n2619 gnd 0.007198f
C3720 vdd.n2620 gnd 0.007198f
C3721 vdd.n2621 gnd 0.005557f
C3722 vdd.n2622 gnd 0.007198f
C3723 vdd.n2623 gnd 0.007198f
C3724 vdd.n2624 gnd 0.01708f
C3725 vdd.n2625 gnd 0.015947f
C3726 vdd.n2626 gnd 0.007198f
C3727 vdd.n2627 gnd 0.007198f
C3728 vdd.n2628 gnd 0.007198f
C3729 vdd.n2629 gnd 0.007198f
C3730 vdd.n2630 gnd 0.007198f
C3731 vdd.n2631 gnd 0.007198f
C3732 vdd.n2632 gnd 0.007198f
C3733 vdd.n2633 gnd 0.007198f
C3734 vdd.n2634 gnd 0.007198f
C3735 vdd.n2635 gnd 0.007198f
C3736 vdd.n2636 gnd 0.007198f
C3737 vdd.n2637 gnd 0.007198f
C3738 vdd.n2638 gnd 0.007198f
C3739 vdd.n2639 gnd 0.007198f
C3740 vdd.n2640 gnd 0.007198f
C3741 vdd.n2641 gnd 0.007198f
C3742 vdd.n2642 gnd 0.007198f
C3743 vdd.n2643 gnd 0.007198f
C3744 vdd.n2644 gnd 0.007198f
C3745 vdd.n2645 gnd 0.007198f
C3746 vdd.n2646 gnd 0.007198f
C3747 vdd.n2647 gnd 0.007198f
C3748 vdd.n2648 gnd 0.007198f
C3749 vdd.n2649 gnd 0.007198f
C3750 vdd.n2650 gnd 0.007198f
C3751 vdd.n2651 gnd 0.007198f
C3752 vdd.n2652 gnd 0.007198f
C3753 vdd.n2653 gnd 0.007198f
C3754 vdd.n2654 gnd 0.007198f
C3755 vdd.n2655 gnd 0.007198f
C3756 vdd.n2656 gnd 0.007198f
C3757 vdd.n2657 gnd 0.007198f
C3758 vdd.n2658 gnd 0.007198f
C3759 vdd.n2659 gnd 0.007198f
C3760 vdd.n2660 gnd 0.007198f
C3761 vdd.n2661 gnd 0.007198f
C3762 vdd.n2662 gnd 0.007198f
C3763 vdd.n2663 gnd 0.007198f
C3764 vdd.n2664 gnd 0.007198f
C3765 vdd.n2665 gnd 0.007198f
C3766 vdd.n2666 gnd 0.007198f
C3767 vdd.n2667 gnd 0.007198f
C3768 vdd.n2668 gnd 0.007198f
C3769 vdd.n2669 gnd 0.007198f
C3770 vdd.n2670 gnd 0.007198f
C3771 vdd.n2671 gnd 0.007198f
C3772 vdd.n2672 gnd 0.007198f
C3773 vdd.n2673 gnd 0.007198f
C3774 vdd.n2674 gnd 0.007198f
C3775 vdd.n2675 gnd 0.007198f
C3776 vdd.n2676 gnd 0.007198f
C3777 vdd.n2677 gnd 0.232581f
C3778 vdd.n2678 gnd 0.007198f
C3779 vdd.n2679 gnd 0.007198f
C3780 vdd.n2680 gnd 0.007198f
C3781 vdd.n2681 gnd 0.007198f
C3782 vdd.n2682 gnd 0.007198f
C3783 vdd.n2683 gnd 0.007198f
C3784 vdd.n2684 gnd 0.007198f
C3785 vdd.n2685 gnd 0.007198f
C3786 vdd.n2686 gnd 0.007198f
C3787 vdd.n2687 gnd 0.007198f
C3788 vdd.n2688 gnd 0.007198f
C3789 vdd.n2689 gnd 0.007198f
C3790 vdd.n2690 gnd 0.007198f
C3791 vdd.n2691 gnd 0.007198f
C3792 vdd.n2692 gnd 0.007198f
C3793 vdd.n2693 gnd 0.007198f
C3794 vdd.n2694 gnd 0.007198f
C3795 vdd.n2695 gnd 0.007198f
C3796 vdd.n2696 gnd 0.007198f
C3797 vdd.n2697 gnd 0.007198f
C3798 vdd.n2698 gnd 0.438118f
C3799 vdd.n2699 gnd 0.007198f
C3800 vdd.n2700 gnd 0.007198f
C3801 vdd.n2701 gnd 0.007198f
C3802 vdd.n2702 gnd 0.007198f
C3803 vdd.n2703 gnd 0.007198f
C3804 vdd.n2704 gnd 0.015947f
C3805 vdd.n2705 gnd 0.01708f
C3806 vdd.n2706 gnd 0.01708f
C3807 vdd.n2707 gnd 0.007198f
C3808 vdd.n2708 gnd 0.007198f
C3809 vdd.n2709 gnd 0.007198f
C3810 vdd.n2710 gnd 0.005557f
C3811 vdd.n2711 gnd 0.010287f
C3812 vdd.n2712 gnd 0.00524f
C3813 vdd.n2713 gnd 0.007198f
C3814 vdd.n2714 gnd 0.007198f
C3815 vdd.n2715 gnd 0.007198f
C3816 vdd.n2716 gnd 0.007198f
C3817 vdd.n2717 gnd 0.007198f
C3818 vdd.n2718 gnd 0.007198f
C3819 vdd.n2719 gnd 0.007198f
C3820 vdd.n2720 gnd 0.007198f
C3821 vdd.n2721 gnd 0.007198f
C3822 vdd.n2722 gnd 0.007198f
C3823 vdd.n2723 gnd 0.007198f
C3824 vdd.n2724 gnd 0.007198f
C3825 vdd.n2725 gnd 0.007198f
C3826 vdd.n2726 gnd 0.007198f
C3827 vdd.n2727 gnd 0.007198f
C3828 vdd.n2728 gnd 0.007198f
C3829 vdd.n2729 gnd 0.007198f
C3830 vdd.n2730 gnd 0.007198f
C3831 vdd.n2731 gnd 0.007198f
C3832 vdd.n2732 gnd 0.007198f
C3833 vdd.n2733 gnd 0.007198f
C3834 vdd.n2734 gnd 0.007198f
C3835 vdd.n2735 gnd 0.007198f
C3836 vdd.n2736 gnd 0.007198f
C3837 vdd.n2737 gnd 0.007198f
C3838 vdd.n2738 gnd 0.007198f
C3839 vdd.n2739 gnd 0.007198f
C3840 vdd.n2740 gnd 0.007198f
C3841 vdd.n2741 gnd 0.007198f
C3842 vdd.n2742 gnd 0.007198f
C3843 vdd.n2743 gnd 0.007198f
C3844 vdd.n2744 gnd 0.007198f
C3845 vdd.n2745 gnd 0.007198f
C3846 vdd.n2746 gnd 0.007198f
C3847 vdd.n2747 gnd 0.007198f
C3848 vdd.n2748 gnd 0.007198f
C3849 vdd.n2749 gnd 0.007198f
C3850 vdd.n2750 gnd 0.007198f
C3851 vdd.n2751 gnd 0.007198f
C3852 vdd.n2752 gnd 0.007198f
C3853 vdd.n2753 gnd 0.007198f
C3854 vdd.n2754 gnd 0.007198f
C3855 vdd.n2755 gnd 0.007198f
C3856 vdd.n2756 gnd 0.007198f
C3857 vdd.n2757 gnd 0.007198f
C3858 vdd.n2758 gnd 0.007198f
C3859 vdd.n2759 gnd 0.007198f
C3860 vdd.n2760 gnd 0.007198f
C3861 vdd.n2761 gnd 0.007198f
C3862 vdd.n2762 gnd 0.007198f
C3863 vdd.n2763 gnd 0.007198f
C3864 vdd.n2764 gnd 0.007198f
C3865 vdd.n2765 gnd 0.007198f
C3866 vdd.n2766 gnd 0.007198f
C3867 vdd.n2767 gnd 0.007198f
C3868 vdd.n2768 gnd 0.007198f
C3869 vdd.n2769 gnd 0.007198f
C3870 vdd.n2770 gnd 0.007198f
C3871 vdd.n2771 gnd 0.007198f
C3872 vdd.n2772 gnd 0.007198f
C3873 vdd.n2774 gnd 0.897872f
C3874 vdd.n2776 gnd 0.007198f
C3875 vdd.n2777 gnd 0.007198f
C3876 vdd.n2778 gnd 0.01708f
C3877 vdd.n2779 gnd 0.015947f
C3878 vdd.n2780 gnd 0.015947f
C3879 vdd.n2781 gnd 0.897872f
C3880 vdd.n2782 gnd 0.015947f
C3881 vdd.n2783 gnd 0.015947f
C3882 vdd.n2784 gnd 0.007198f
C3883 vdd.n2785 gnd 0.007198f
C3884 vdd.n2786 gnd 0.007198f
C3885 vdd.n2787 gnd 0.459754f
C3886 vdd.n2788 gnd 0.007198f
C3887 vdd.n2789 gnd 0.007198f
C3888 vdd.n2790 gnd 0.007198f
C3889 vdd.n2791 gnd 0.007198f
C3890 vdd.n2792 gnd 0.007198f
C3891 vdd.n2793 gnd 0.57334f
C3892 vdd.n2794 gnd 0.007198f
C3893 vdd.n2795 gnd 0.007198f
C3894 vdd.n2796 gnd 0.007198f
C3895 vdd.n2797 gnd 0.007198f
C3896 vdd.n2798 gnd 0.007198f
C3897 vdd.n2799 gnd 0.735606f
C3898 vdd.n2800 gnd 0.007198f
C3899 vdd.n2801 gnd 0.007198f
C3900 vdd.n2802 gnd 0.007198f
C3901 vdd.n2803 gnd 0.007198f
C3902 vdd.n2804 gnd 0.007198f
C3903 vdd.n2805 gnd 0.405665f
C3904 vdd.n2806 gnd 0.007198f
C3905 vdd.n2807 gnd 0.007198f
C3906 vdd.n2808 gnd 0.007198f
C3907 vdd.n2809 gnd 0.007198f
C3908 vdd.n2810 gnd 0.007198f
C3909 vdd.n2811 gnd 0.232581f
C3910 vdd.n2812 gnd 0.007198f
C3911 vdd.n2813 gnd 0.007198f
C3912 vdd.n2814 gnd 0.007198f
C3913 vdd.n2815 gnd 0.007198f
C3914 vdd.n2816 gnd 0.007198f
C3915 vdd.n2817 gnd 0.421892f
C3916 vdd.n2818 gnd 0.007198f
C3917 vdd.n2819 gnd 0.007198f
C3918 vdd.n2820 gnd 0.007198f
C3919 vdd.n2821 gnd 0.007198f
C3920 vdd.n2822 gnd 0.007198f
C3921 vdd.n2823 gnd 0.584158f
C3922 vdd.n2824 gnd 0.007198f
C3923 vdd.n2825 gnd 0.007198f
C3924 vdd.n2826 gnd 0.007198f
C3925 vdd.n2827 gnd 0.007198f
C3926 vdd.n2828 gnd 0.007198f
C3927 vdd.n2829 gnd 0.654473f
C3928 vdd.n2830 gnd 0.007198f
C3929 vdd.n2831 gnd 0.007198f
C3930 vdd.n2832 gnd 0.007198f
C3931 vdd.n2833 gnd 0.007198f
C3932 vdd.n2834 gnd 0.007198f
C3933 vdd.n2835 gnd 0.492207f
C3934 vdd.n2836 gnd 0.007198f
C3935 vdd.n2837 gnd 0.007198f
C3936 vdd.n2838 gnd 0.007198f
C3937 vdd.t204 gnd 0.297744f
C3938 vdd.t202 gnd 0.189892f
C3939 vdd.t205 gnd 0.297744f
C3940 vdd.n2839 gnd 0.167344f
C3941 vdd.n2840 gnd 0.020852f
C3942 vdd.n2841 gnd 0.004446f
C3943 vdd.n2842 gnd 0.007198f
C3944 vdd.n2843 gnd 0.405665f
C3945 vdd.n2844 gnd 0.007198f
C3946 vdd.n2845 gnd 0.007198f
C3947 vdd.n2846 gnd 0.007198f
C3948 vdd.n2847 gnd 0.007198f
C3949 vdd.n2848 gnd 0.007198f
C3950 vdd.n2849 gnd 0.735606f
C3951 vdd.n2850 gnd 0.007198f
C3952 vdd.n2851 gnd 0.007198f
C3953 vdd.n2852 gnd 0.007198f
C3954 vdd.n2853 gnd 0.007198f
C3955 vdd.n2854 gnd 0.007198f
C3956 vdd.n2855 gnd 0.007198f
C3957 vdd.n2857 gnd 0.007198f
C3958 vdd.n2858 gnd 0.007198f
C3959 vdd.n2860 gnd 0.007198f
C3960 vdd.n2861 gnd 0.007198f
C3961 vdd.n2864 gnd 0.007198f
C3962 vdd.n2865 gnd 0.007198f
C3963 vdd.n2866 gnd 0.007198f
C3964 vdd.n2867 gnd 0.007198f
C3965 vdd.n2869 gnd 0.007198f
C3966 vdd.n2870 gnd 0.007198f
C3967 vdd.n2871 gnd 0.007198f
C3968 vdd.n2872 gnd 0.007198f
C3969 vdd.n2873 gnd 0.007198f
C3970 vdd.n2874 gnd 0.007198f
C3971 vdd.n2876 gnd 0.007198f
C3972 vdd.n2877 gnd 0.007198f
C3973 vdd.n2878 gnd 0.007198f
C3974 vdd.n2879 gnd 0.007198f
C3975 vdd.n2880 gnd 0.007198f
C3976 vdd.n2881 gnd 0.007198f
C3977 vdd.n2883 gnd 0.007198f
C3978 vdd.n2884 gnd 0.007198f
C3979 vdd.n2885 gnd 0.007198f
C3980 vdd.n2886 gnd 0.007198f
C3981 vdd.n2887 gnd 0.007198f
C3982 vdd.n2888 gnd 0.007198f
C3983 vdd.n2890 gnd 0.007198f
C3984 vdd.n2891 gnd 0.01708f
C3985 vdd.n2892 gnd 0.01708f
C3986 vdd.n2893 gnd 0.015947f
C3987 vdd.n2894 gnd 0.007198f
C3988 vdd.n2895 gnd 0.007198f
C3989 vdd.n2896 gnd 0.007198f
C3990 vdd.n2897 gnd 0.007198f
C3991 vdd.n2898 gnd 0.007198f
C3992 vdd.n2899 gnd 0.007198f
C3993 vdd.n2900 gnd 0.735606f
C3994 vdd.n2901 gnd 0.007198f
C3995 vdd.n2902 gnd 0.007198f
C3996 vdd.n2903 gnd 0.007198f
C3997 vdd.n2904 gnd 0.007198f
C3998 vdd.n2905 gnd 0.007198f
C3999 vdd.n2906 gnd 0.459754f
C4000 vdd.n2907 gnd 0.007198f
C4001 vdd.n2908 gnd 0.007198f
C4002 vdd.n2909 gnd 0.007198f
C4003 vdd.n2910 gnd 0.016823f
C4004 vdd.n2912 gnd 0.01708f
C4005 vdd.n2913 gnd 0.016203f
C4006 vdd.n2914 gnd 0.007198f
C4007 vdd.n2915 gnd 0.005557f
C4008 vdd.n2916 gnd 0.007198f
C4009 vdd.n2918 gnd 0.007198f
C4010 vdd.n2919 gnd 0.007198f
C4011 vdd.n2920 gnd 0.007198f
C4012 vdd.n2921 gnd 0.007198f
C4013 vdd.n2922 gnd 0.007198f
C4014 vdd.n2923 gnd 0.007198f
C4015 vdd.n2925 gnd 0.007198f
C4016 vdd.n2926 gnd 0.007198f
C4017 vdd.n2927 gnd 0.007198f
C4018 vdd.n2928 gnd 0.007198f
C4019 vdd.n2929 gnd 0.007198f
C4020 vdd.n2930 gnd 0.007198f
C4021 vdd.n2932 gnd 0.007198f
C4022 vdd.n2933 gnd 0.007198f
C4023 vdd.n2934 gnd 0.007198f
C4024 vdd.n2935 gnd 0.007198f
C4025 vdd.n2936 gnd 0.007198f
C4026 vdd.n2937 gnd 0.007198f
C4027 vdd.n2939 gnd 0.007198f
C4028 vdd.n2940 gnd 0.007198f
C4029 vdd.n2941 gnd 0.007198f
C4030 vdd.n2942 gnd 0.640643f
C4031 vdd.n2943 gnd 0.017297f
C4032 vdd.n2944 gnd 0.007198f
C4033 vdd.n2945 gnd 0.007198f
C4034 vdd.n2947 gnd 0.007198f
C4035 vdd.n2948 gnd 0.007198f
C4036 vdd.n2949 gnd 0.007198f
C4037 vdd.n2950 gnd 0.007198f
C4038 vdd.n2951 gnd 0.007198f
C4039 vdd.n2952 gnd 0.007198f
C4040 vdd.n2954 gnd 0.007198f
C4041 vdd.n2955 gnd 0.007198f
C4042 vdd.n2956 gnd 0.007198f
C4043 vdd.n2957 gnd 0.007198f
C4044 vdd.n2958 gnd 0.007198f
C4045 vdd.n2959 gnd 0.007198f
C4046 vdd.n2961 gnd 0.007198f
C4047 vdd.n2962 gnd 0.007198f
C4048 vdd.n2963 gnd 0.007198f
C4049 vdd.n2964 gnd 0.007198f
C4050 vdd.n2965 gnd 0.007198f
C4051 vdd.n2966 gnd 0.007198f
C4052 vdd.n2968 gnd 0.007198f
C4053 vdd.n2969 gnd 0.007198f
C4054 vdd.n2971 gnd 0.007198f
C4055 vdd.n2972 gnd 0.007198f
C4056 vdd.n2973 gnd 0.01708f
C4057 vdd.n2974 gnd 0.015947f
C4058 vdd.n2975 gnd 0.015947f
C4059 vdd.n2976 gnd 1.06014f
C4060 vdd.n2977 gnd 0.015947f
C4061 vdd.n2978 gnd 0.01708f
C4062 vdd.n2979 gnd 0.016203f
C4063 vdd.n2980 gnd 0.007198f
C4064 vdd.n2981 gnd 0.005557f
C4065 vdd.n2982 gnd 0.007198f
C4066 vdd.n2984 gnd 0.007198f
C4067 vdd.n2985 gnd 0.007198f
C4068 vdd.n2986 gnd 0.007198f
C4069 vdd.n2987 gnd 0.007198f
C4070 vdd.n2988 gnd 0.007198f
C4071 vdd.n2989 gnd 0.007198f
C4072 vdd.n2991 gnd 0.007198f
C4073 vdd.n2992 gnd 0.007198f
C4074 vdd.n2993 gnd 0.007198f
C4075 vdd.n2994 gnd 0.007198f
C4076 vdd.n2995 gnd 0.007198f
C4077 vdd.n2996 gnd 0.007198f
C4078 vdd.n2998 gnd 0.007198f
C4079 vdd.n2999 gnd 0.007198f
C4080 vdd.n3000 gnd 0.007198f
C4081 vdd.n3001 gnd 0.007198f
C4082 vdd.n3002 gnd 0.007198f
C4083 vdd.n3003 gnd 0.007198f
C4084 vdd.n3005 gnd 0.007198f
C4085 vdd.n3006 gnd 0.007198f
C4086 vdd.n3008 gnd 0.007198f
C4087 vdd.n3009 gnd 0.017297f
C4088 vdd.n3010 gnd 0.640643f
C4089 vdd.n3011 gnd 0.009103f
C4090 vdd.n3012 gnd 0.004047f
C4091 vdd.t248 gnd 0.130228f
C4092 vdd.t249 gnd 0.139178f
C4093 vdd.t247 gnd 0.170076f
C4094 vdd.n3013 gnd 0.218013f
C4095 vdd.n3014 gnd 0.18317f
C4096 vdd.n3015 gnd 0.013121f
C4097 vdd.n3016 gnd 0.010585f
C4098 vdd.n3017 gnd 0.004473f
C4099 vdd.n3018 gnd 0.00852f
C4100 vdd.n3019 gnd 0.010585f
C4101 vdd.n3020 gnd 0.010585f
C4102 vdd.n3021 gnd 0.00852f
C4103 vdd.n3022 gnd 0.00852f
C4104 vdd.n3023 gnd 0.010585f
C4105 vdd.n3025 gnd 0.010585f
C4106 vdd.n3026 gnd 0.00852f
C4107 vdd.n3027 gnd 0.00852f
C4108 vdd.n3028 gnd 0.00852f
C4109 vdd.n3029 gnd 0.010585f
C4110 vdd.n3031 gnd 0.010585f
C4111 vdd.n3033 gnd 0.010585f
C4112 vdd.n3034 gnd 0.00852f
C4113 vdd.n3035 gnd 0.00852f
C4114 vdd.n3036 gnd 0.00852f
C4115 vdd.n3037 gnd 0.010585f
C4116 vdd.n3039 gnd 0.010585f
C4117 vdd.n3041 gnd 0.010585f
C4118 vdd.n3042 gnd 0.00852f
C4119 vdd.n3043 gnd 0.00852f
C4120 vdd.n3044 gnd 0.00852f
C4121 vdd.n3045 gnd 0.010585f
C4122 vdd.n3047 gnd 0.010585f
C4123 vdd.n3048 gnd 0.010585f
C4124 vdd.n3049 gnd 0.00852f
C4125 vdd.n3050 gnd 0.00852f
C4126 vdd.n3051 gnd 0.010585f
C4127 vdd.n3052 gnd 0.010585f
C4128 vdd.n3054 gnd 0.010585f
C4129 vdd.n3055 gnd 0.00852f
C4130 vdd.n3056 gnd 0.010585f
C4131 vdd.n3057 gnd 0.010585f
C4132 vdd.n3058 gnd 0.010585f
C4133 vdd.n3059 gnd 0.017381f
C4134 vdd.n3060 gnd 0.005794f
C4135 vdd.n3061 gnd 0.010585f
C4136 vdd.n3063 gnd 0.010585f
C4137 vdd.n3065 gnd 0.010585f
C4138 vdd.n3066 gnd 0.00852f
C4139 vdd.n3067 gnd 0.00852f
C4140 vdd.n3068 gnd 0.00852f
C4141 vdd.n3069 gnd 0.010585f
C4142 vdd.n3071 gnd 0.010585f
C4143 vdd.n3073 gnd 0.010585f
C4144 vdd.n3074 gnd 0.00852f
C4145 vdd.n3075 gnd 0.00852f
C4146 vdd.n3076 gnd 0.00852f
C4147 vdd.n3077 gnd 0.010585f
C4148 vdd.n3079 gnd 0.010585f
C4149 vdd.n3081 gnd 0.010585f
C4150 vdd.n3082 gnd 0.00852f
C4151 vdd.n3083 gnd 0.00852f
C4152 vdd.n3084 gnd 0.00852f
C4153 vdd.n3085 gnd 0.010585f
C4154 vdd.n3087 gnd 0.010585f
C4155 vdd.n3089 gnd 0.010585f
C4156 vdd.n3090 gnd 0.00852f
C4157 vdd.n3091 gnd 0.00852f
C4158 vdd.n3092 gnd 0.00852f
C4159 vdd.n3093 gnd 0.010585f
C4160 vdd.n3095 gnd 0.010585f
C4161 vdd.n3097 gnd 0.010585f
C4162 vdd.n3098 gnd 0.00852f
C4163 vdd.n3099 gnd 0.00852f
C4164 vdd.n3100 gnd 0.007114f
C4165 vdd.n3101 gnd 0.010585f
C4166 vdd.n3103 gnd 0.010585f
C4167 vdd.n3105 gnd 0.010585f
C4168 vdd.n3106 gnd 0.007114f
C4169 vdd.n3107 gnd 0.00852f
C4170 vdd.n3108 gnd 0.00852f
C4171 vdd.n3109 gnd 0.010585f
C4172 vdd.n3111 gnd 0.010585f
C4173 vdd.n3113 gnd 0.010585f
C4174 vdd.n3114 gnd 0.00852f
C4175 vdd.n3115 gnd 0.00852f
C4176 vdd.n3116 gnd 0.00852f
C4177 vdd.n3117 gnd 0.010585f
C4178 vdd.n3119 gnd 0.010585f
C4179 vdd.n3121 gnd 0.010585f
C4180 vdd.n3122 gnd 0.00852f
C4181 vdd.n3123 gnd 0.00852f
C4182 vdd.n3124 gnd 0.00852f
C4183 vdd.n3125 gnd 0.010585f
C4184 vdd.n3127 gnd 0.010585f
C4185 vdd.n3128 gnd 0.010585f
C4186 vdd.n3129 gnd 0.00852f
C4187 vdd.n3130 gnd 0.00852f
C4188 vdd.n3131 gnd 0.010585f
C4189 vdd.n3132 gnd 0.010585f
C4190 vdd.n3133 gnd 0.00852f
C4191 vdd.n3134 gnd 0.00852f
C4192 vdd.n3135 gnd 0.010585f
C4193 vdd.n3136 gnd 0.010585f
C4194 vdd.n3138 gnd 0.010585f
C4195 vdd.n3139 gnd 0.00852f
C4196 vdd.n3140 gnd 0.007072f
C4197 vdd.n3141 gnd 0.02427f
C4198 vdd.n3142 gnd 0.024105f
C4199 vdd.n3143 gnd 0.007072f
C4200 vdd.n3144 gnd 0.024105f
C4201 vdd.n3145 gnd 1.42794f
C4202 vdd.n3146 gnd 0.024105f
C4203 vdd.n3147 gnd 0.007072f
C4204 vdd.n3148 gnd 0.024105f
C4205 vdd.n3149 gnd 0.010585f
C4206 vdd.n3150 gnd 0.010585f
C4207 vdd.n3151 gnd 0.00852f
C4208 vdd.n3152 gnd 0.010585f
C4209 vdd.n3153 gnd 1.02228f
C4210 vdd.n3154 gnd 0.010585f
C4211 vdd.n3155 gnd 0.00852f
C4212 vdd.n3156 gnd 0.010585f
C4213 vdd.n3157 gnd 0.010585f
C4214 vdd.n3158 gnd 0.010585f
C4215 vdd.n3159 gnd 0.00852f
C4216 vdd.n3160 gnd 0.010585f
C4217 vdd.n3161 gnd 1.05473f
C4218 vdd.n3162 gnd 0.010585f
C4219 vdd.n3163 gnd 0.00852f
C4220 vdd.n3164 gnd 0.010585f
C4221 vdd.n3165 gnd 0.010585f
C4222 vdd.n3166 gnd 0.010585f
C4223 vdd.n3167 gnd 0.00852f
C4224 vdd.n3168 gnd 0.010585f
C4225 vdd.t80 gnd 0.540887f
C4226 vdd.n3169 gnd 0.870828f
C4227 vdd.n3170 gnd 0.010585f
C4228 vdd.n3171 gnd 0.00852f
C4229 vdd.n3172 gnd 0.010585f
C4230 vdd.n3173 gnd 0.010585f
C4231 vdd.n3174 gnd 0.010585f
C4232 vdd.n3175 gnd 0.00852f
C4233 vdd.n3176 gnd 0.010585f
C4234 vdd.n3177 gnd 0.686926f
C4235 vdd.n3178 gnd 0.010585f
C4236 vdd.n3179 gnd 0.00852f
C4237 vdd.n3180 gnd 0.010585f
C4238 vdd.n3181 gnd 0.010585f
C4239 vdd.n3182 gnd 0.010585f
C4240 vdd.n3183 gnd 0.00852f
C4241 vdd.n3184 gnd 0.010585f
C4242 vdd.n3185 gnd 0.86001f
C4243 vdd.n3186 gnd 0.578749f
C4244 vdd.n3187 gnd 0.010585f
C4245 vdd.n3188 gnd 0.00852f
C4246 vdd.n3189 gnd 0.010585f
C4247 vdd.n3190 gnd 0.010585f
C4248 vdd.n3191 gnd 0.010585f
C4249 vdd.n3192 gnd 0.00852f
C4250 vdd.n3193 gnd 0.010585f
C4251 vdd.n3194 gnd 0.76265f
C4252 vdd.n3195 gnd 0.010585f
C4253 vdd.n3196 gnd 0.00852f
C4254 vdd.n3197 gnd 0.010585f
C4255 vdd.n3198 gnd 0.010585f
C4256 vdd.n3199 gnd 0.010585f
C4257 vdd.n3200 gnd 0.010585f
C4258 vdd.n3201 gnd 0.010585f
C4259 vdd.n3202 gnd 0.00852f
C4260 vdd.n3203 gnd 0.00852f
C4261 vdd.n3204 gnd 0.010585f
C4262 vdd.t35 gnd 0.540887f
C4263 vdd.n3205 gnd 0.897872f
C4264 vdd.n3206 gnd 0.010585f
C4265 vdd.n3207 gnd 0.00852f
C4266 vdd.n3208 gnd 0.010585f
C4267 vdd.n3209 gnd 0.010585f
C4268 vdd.n3210 gnd 0.010585f
C4269 vdd.n3211 gnd 0.00852f
C4270 vdd.n3212 gnd 0.010585f
C4271 vdd.n3213 gnd 0.849192f
C4272 vdd.n3214 gnd 0.010585f
C4273 vdd.n3215 gnd 0.010585f
C4274 vdd.n3216 gnd 0.00852f
C4275 vdd.n3217 gnd 0.00852f
C4276 vdd.n3218 gnd 0.00852f
C4277 vdd.n3219 gnd 0.010585f
C4278 vdd.n3220 gnd 0.010585f
C4279 vdd.n3221 gnd 0.010585f
C4280 vdd.n3222 gnd 0.010585f
C4281 vdd.n3223 gnd 0.00852f
C4282 vdd.n3224 gnd 0.00852f
C4283 vdd.n3225 gnd 0.00852f
C4284 vdd.n3226 gnd 0.010585f
C4285 vdd.n3227 gnd 0.010585f
C4286 vdd.n3228 gnd 0.010585f
C4287 vdd.n3229 gnd 0.010585f
C4288 vdd.n3230 gnd 0.00852f
C4289 vdd.n3231 gnd 0.00852f
C4290 vdd.n3232 gnd 0.00852f
C4291 vdd.n3233 gnd 0.010585f
C4292 vdd.n3234 gnd 0.010585f
C4293 vdd.n3235 gnd 0.010585f
C4294 vdd.n3236 gnd 0.897872f
C4295 vdd.n3237 gnd 0.010585f
C4296 vdd.n3238 gnd 0.00852f
C4297 vdd.n3239 gnd 0.00852f
C4298 vdd.n3240 gnd 0.00852f
C4299 vdd.n3241 gnd 0.010585f
C4300 vdd.n3242 gnd 0.010585f
C4301 vdd.n3243 gnd 0.010585f
C4302 vdd.n3244 gnd 0.010585f
C4303 vdd.n3245 gnd 0.00852f
C4304 vdd.n3246 gnd 0.00852f
C4305 vdd.n3247 gnd 0.007072f
C4306 vdd.n3248 gnd 0.024105f
C4307 vdd.n3249 gnd 0.02427f
C4308 vdd.n3250 gnd 0.004047f
C4309 vdd.n3251 gnd 0.02427f
C4310 vdd.n3253 gnd 2.39072f
C4311 vdd.n3254 gnd 1.42794f
C4312 vdd.n3255 gnd 0.708562f
C4313 vdd.n3256 gnd 0.010585f
C4314 vdd.n3257 gnd 0.00852f
C4315 vdd.n3258 gnd 0.00852f
C4316 vdd.n3259 gnd 0.00852f
C4317 vdd.n3260 gnd 0.010585f
C4318 vdd.n3261 gnd 1.08177f
C4319 vdd.n3262 gnd 1.08177f
C4320 vdd.n3263 gnd 0.62202f
C4321 vdd.n3264 gnd 0.010585f
C4322 vdd.n3265 gnd 0.00852f
C4323 vdd.n3266 gnd 0.00852f
C4324 vdd.n3267 gnd 0.00852f
C4325 vdd.n3268 gnd 0.010585f
C4326 vdd.n3269 gnd 0.643655f
C4327 vdd.n3270 gnd 0.795103f
C4328 vdd.t53 gnd 0.540887f
C4329 vdd.n3271 gnd 0.827557f
C4330 vdd.n3272 gnd 0.010585f
C4331 vdd.n3273 gnd 0.00852f
C4332 vdd.n3274 gnd 0.00852f
C4333 vdd.n3275 gnd 0.00852f
C4334 vdd.n3276 gnd 0.010585f
C4335 vdd.n3277 gnd 0.897872f
C4336 vdd.t29 gnd 0.540887f
C4337 vdd.n3278 gnd 0.654473f
C4338 vdd.n3279 gnd 0.784286f
C4339 vdd.n3280 gnd 0.010585f
C4340 vdd.n3281 gnd 0.00852f
C4341 vdd.n3282 gnd 0.00852f
C4342 vdd.n3283 gnd 0.00852f
C4343 vdd.n3284 gnd 0.010585f
C4344 vdd.n3285 gnd 0.600384f
C4345 vdd.t21 gnd 0.540887f
C4346 vdd.n3286 gnd 0.897872f
C4347 vdd.t57 gnd 0.540887f
C4348 vdd.n3287 gnd 0.665291f
C4349 vdd.n3288 gnd 0.010585f
C4350 vdd.n3289 gnd 0.00852f
C4351 vdd.n3290 gnd 0.008136f
C4352 vdd.n3291 gnd 0.624364f
C4353 vdd.n3292 gnd 2.52013f
C4354 a_n6972_8799.n0 gnd 0.207737f
C4355 a_n6972_8799.n1 gnd 0.290352f
C4356 a_n6972_8799.n2 gnd 0.207737f
C4357 a_n6972_8799.n3 gnd 0.207737f
C4358 a_n6972_8799.n4 gnd 0.207737f
C4359 a_n6972_8799.n5 gnd 0.273684f
C4360 a_n6972_8799.n6 gnd 0.207737f
C4361 a_n6972_8799.n7 gnd 0.290352f
C4362 a_n6972_8799.n8 gnd 0.207737f
C4363 a_n6972_8799.n9 gnd 0.207737f
C4364 a_n6972_8799.n10 gnd 0.207737f
C4365 a_n6972_8799.n11 gnd 0.273684f
C4366 a_n6972_8799.n12 gnd 0.207737f
C4367 a_n6972_8799.n13 gnd 0.455038f
C4368 a_n6972_8799.n14 gnd 0.207737f
C4369 a_n6972_8799.n15 gnd 0.207737f
C4370 a_n6972_8799.n16 gnd 0.207737f
C4371 a_n6972_8799.n17 gnd 0.273684f
C4372 a_n6972_8799.n18 gnd 0.325619f
C4373 a_n6972_8799.n19 gnd 0.207737f
C4374 a_n6972_8799.n20 gnd 0.207737f
C4375 a_n6972_8799.n21 gnd 0.207737f
C4376 a_n6972_8799.n22 gnd 0.207737f
C4377 a_n6972_8799.n23 gnd 0.238418f
C4378 a_n6972_8799.n24 gnd 0.325619f
C4379 a_n6972_8799.n25 gnd 0.207737f
C4380 a_n6972_8799.n26 gnd 0.207737f
C4381 a_n6972_8799.n27 gnd 0.207737f
C4382 a_n6972_8799.n28 gnd 0.207737f
C4383 a_n6972_8799.n29 gnd 0.238418f
C4384 a_n6972_8799.n30 gnd 0.325619f
C4385 a_n6972_8799.n31 gnd 0.207737f
C4386 a_n6972_8799.n32 gnd 0.207737f
C4387 a_n6972_8799.n33 gnd 0.207737f
C4388 a_n6972_8799.n34 gnd 0.207737f
C4389 a_n6972_8799.n35 gnd 0.403104f
C4390 a_n6972_8799.n36 gnd 4.02811f
C4391 a_n6972_8799.n37 gnd 2.79029f
C4392 a_n6972_8799.n38 gnd 0.363145f
C4393 a_n6972_8799.n39 gnd 3.04349f
C4394 a_n6972_8799.n40 gnd 0.363144f
C4395 a_n6972_8799.n41 gnd 0.8559f
C4396 a_n6972_8799.n42 gnd 0.008616f
C4397 a_n6972_8799.n43 gnd 0.001157f
C4398 a_n6972_8799.n45 gnd 0.007738f
C4399 a_n6972_8799.n46 gnd 0.011695f
C4400 a_n6972_8799.n47 gnd 0.008043f
C4401 a_n6972_8799.n49 gnd 4.02e-19
C4402 a_n6972_8799.n50 gnd 0.008335f
C4403 a_n6972_8799.n51 gnd 0.011513f
C4404 a_n6972_8799.n52 gnd 0.007418f
C4405 a_n6972_8799.n53 gnd 0.008616f
C4406 a_n6972_8799.n54 gnd 0.001157f
C4407 a_n6972_8799.n56 gnd 0.007738f
C4408 a_n6972_8799.n57 gnd 0.011695f
C4409 a_n6972_8799.n58 gnd 0.008043f
C4410 a_n6972_8799.n60 gnd 4.02e-19
C4411 a_n6972_8799.n61 gnd 0.008335f
C4412 a_n6972_8799.n62 gnd 0.011513f
C4413 a_n6972_8799.n63 gnd 0.007418f
C4414 a_n6972_8799.n64 gnd 0.008616f
C4415 a_n6972_8799.n65 gnd 0.001157f
C4416 a_n6972_8799.n67 gnd 0.007738f
C4417 a_n6972_8799.n68 gnd 0.011695f
C4418 a_n6972_8799.n69 gnd 0.008043f
C4419 a_n6972_8799.n71 gnd 4.02e-19
C4420 a_n6972_8799.n72 gnd 0.008335f
C4421 a_n6972_8799.n73 gnd 0.011513f
C4422 a_n6972_8799.n74 gnd 0.007418f
C4423 a_n6972_8799.n75 gnd 0.001157f
C4424 a_n6972_8799.n77 gnd 0.007738f
C4425 a_n6972_8799.n78 gnd 0.011695f
C4426 a_n6972_8799.n79 gnd 0.008043f
C4427 a_n6972_8799.n81 gnd 4.02e-19
C4428 a_n6972_8799.n82 gnd 0.008335f
C4429 a_n6972_8799.n83 gnd 0.011513f
C4430 a_n6972_8799.n84 gnd 0.007418f
C4431 a_n6972_8799.n85 gnd 0.250096f
C4432 a_n6972_8799.n86 gnd 0.001157f
C4433 a_n6972_8799.n88 gnd 0.007738f
C4434 a_n6972_8799.n89 gnd 0.011695f
C4435 a_n6972_8799.n90 gnd 0.008043f
C4436 a_n6972_8799.n92 gnd 4.02e-19
C4437 a_n6972_8799.n93 gnd 0.008335f
C4438 a_n6972_8799.n94 gnd 0.011513f
C4439 a_n6972_8799.n95 gnd 0.007418f
C4440 a_n6972_8799.n96 gnd 0.250096f
C4441 a_n6972_8799.n97 gnd 0.001157f
C4442 a_n6972_8799.n99 gnd 0.007738f
C4443 a_n6972_8799.n100 gnd 0.011695f
C4444 a_n6972_8799.n101 gnd 0.008043f
C4445 a_n6972_8799.n103 gnd 4.02e-19
C4446 a_n6972_8799.n104 gnd 0.008335f
C4447 a_n6972_8799.n105 gnd 0.011513f
C4448 a_n6972_8799.n106 gnd 0.007418f
C4449 a_n6972_8799.n107 gnd 0.250096f
C4450 a_n6972_8799.t18 gnd 0.144089f
C4451 a_n6972_8799.t3 gnd 0.144089f
C4452 a_n6972_8799.t9 gnd 0.144089f
C4453 a_n6972_8799.n108 gnd 1.13645f
C4454 a_n6972_8799.t4 gnd 0.144089f
C4455 a_n6972_8799.t13 gnd 0.144089f
C4456 a_n6972_8799.n109 gnd 1.13645f
C4457 a_n6972_8799.t12 gnd 0.144089f
C4458 a_n6972_8799.t22 gnd 0.144089f
C4459 a_n6972_8799.n110 gnd 1.13457f
C4460 a_n6972_8799.t7 gnd 0.144089f
C4461 a_n6972_8799.t8 gnd 0.144089f
C4462 a_n6972_8799.n111 gnd 1.13457f
C4463 a_n6972_8799.t15 gnd 0.112069f
C4464 a_n6972_8799.t20 gnd 0.112069f
C4465 a_n6972_8799.n112 gnd 0.993201f
C4466 a_n6972_8799.t28 gnd 0.112069f
C4467 a_n6972_8799.t30 gnd 0.112069f
C4468 a_n6972_8799.n113 gnd 0.990281f
C4469 a_n6972_8799.n114 gnd 0.878129f
C4470 a_n6972_8799.t35 gnd 0.112069f
C4471 a_n6972_8799.t0 gnd 0.112069f
C4472 a_n6972_8799.n115 gnd 0.990281f
C4473 a_n6972_8799.t1 gnd 0.112069f
C4474 a_n6972_8799.t29 gnd 0.112069f
C4475 a_n6972_8799.n116 gnd 0.9932f
C4476 a_n6972_8799.t11 gnd 0.112069f
C4477 a_n6972_8799.t16 gnd 0.112069f
C4478 a_n6972_8799.n117 gnd 0.99028f
C4479 a_n6972_8799.n118 gnd 0.878131f
C4480 a_n6972_8799.t32 gnd 0.112069f
C4481 a_n6972_8799.t5 gnd 0.112069f
C4482 a_n6972_8799.n119 gnd 0.99028f
C4483 a_n6972_8799.t17 gnd 0.112069f
C4484 a_n6972_8799.t33 gnd 0.112069f
C4485 a_n6972_8799.n120 gnd 0.9932f
C4486 a_n6972_8799.t34 gnd 0.112069f
C4487 a_n6972_8799.t6 gnd 0.112069f
C4488 a_n6972_8799.n121 gnd 0.99028f
C4489 a_n6972_8799.n122 gnd 0.878131f
C4490 a_n6972_8799.t24 gnd 0.112069f
C4491 a_n6972_8799.t27 gnd 0.112069f
C4492 a_n6972_8799.n123 gnd 0.99028f
C4493 a_n6972_8799.t19 gnd 0.112069f
C4494 a_n6972_8799.t10 gnd 0.112069f
C4495 a_n6972_8799.n124 gnd 0.990281f
C4496 a_n6972_8799.n125 gnd 3.08917f
C4497 a_n6972_8799.t26 gnd 0.112069f
C4498 a_n6972_8799.t25 gnd 0.112069f
C4499 a_n6972_8799.n126 gnd 0.990281f
C4500 a_n6972_8799.n127 gnd 0.432365f
C4501 a_n6972_8799.t31 gnd 0.112069f
C4502 a_n6972_8799.t23 gnd 0.112069f
C4503 a_n6972_8799.n128 gnd 0.990281f
C4504 a_n6972_8799.t114 gnd 0.597459f
C4505 a_n6972_8799.n129 gnd 0.267109f
C4506 a_n6972_8799.t47 gnd 0.597459f
C4507 a_n6972_8799.t65 gnd 0.597459f
C4508 a_n6972_8799.n130 gnd 0.270418f
C4509 a_n6972_8799.t83 gnd 0.597459f
C4510 a_n6972_8799.t100 gnd 0.597459f
C4511 a_n6972_8799.t101 gnd 0.597459f
C4512 a_n6972_8799.n131 gnd 0.272502f
C4513 a_n6972_8799.t68 gnd 0.597459f
C4514 a_n6972_8799.t78 gnd 0.597459f
C4515 a_n6972_8799.n132 gnd 0.266036f
C4516 a_n6972_8799.t115 gnd 0.608767f
C4517 a_n6972_8799.n133 gnd 0.250481f
C4518 a_n6972_8799.n134 gnd 0.011785f
C4519 a_n6972_8799.t77 gnd 0.597459f
C4520 a_n6972_8799.n135 gnd 0.266836f
C4521 a_n6972_8799.n136 gnd 0.270404f
C4522 a_n6972_8799.t69 gnd 0.597459f
C4523 a_n6972_8799.n137 gnd 0.266926f
C4524 a_n6972_8799.n138 gnd 0.261553f
C4525 a_n6972_8799.t37 gnd 0.597459f
C4526 a_n6972_8799.n139 gnd 0.266676f
C4527 a_n6972_8799.n140 gnd 0.272936f
C4528 a_n6972_8799.t117 gnd 0.597459f
C4529 a_n6972_8799.n141 gnd 0.270286f
C4530 a_n6972_8799.n142 gnd 0.266356f
C4531 a_n6972_8799.t64 gnd 0.597459f
C4532 a_n6972_8799.n143 gnd 0.261873f
C4533 a_n6972_8799.t46 gnd 0.597459f
C4534 a_n6972_8799.n144 gnd 0.270403f
C4535 a_n6972_8799.t45 gnd 0.608756f
C4536 a_n6972_8799.t124 gnd 0.597459f
C4537 a_n6972_8799.n145 gnd 0.267109f
C4538 a_n6972_8799.t61 gnd 0.597459f
C4539 a_n6972_8799.t74 gnd 0.597459f
C4540 a_n6972_8799.n146 gnd 0.270418f
C4541 a_n6972_8799.t94 gnd 0.597459f
C4542 a_n6972_8799.t109 gnd 0.597459f
C4543 a_n6972_8799.t113 gnd 0.597459f
C4544 a_n6972_8799.n147 gnd 0.272502f
C4545 a_n6972_8799.t75 gnd 0.597459f
C4546 a_n6972_8799.t84 gnd 0.597459f
C4547 a_n6972_8799.n148 gnd 0.266036f
C4548 a_n6972_8799.t125 gnd 0.608767f
C4549 a_n6972_8799.n149 gnd 0.250481f
C4550 a_n6972_8799.n150 gnd 0.011785f
C4551 a_n6972_8799.t85 gnd 0.597459f
C4552 a_n6972_8799.n151 gnd 0.266836f
C4553 a_n6972_8799.n152 gnd 0.270404f
C4554 a_n6972_8799.t76 gnd 0.597459f
C4555 a_n6972_8799.n153 gnd 0.266926f
C4556 a_n6972_8799.n154 gnd 0.261553f
C4557 a_n6972_8799.t48 gnd 0.597459f
C4558 a_n6972_8799.n155 gnd 0.266676f
C4559 a_n6972_8799.n156 gnd 0.272936f
C4560 a_n6972_8799.t129 gnd 0.597459f
C4561 a_n6972_8799.n157 gnd 0.270286f
C4562 a_n6972_8799.n158 gnd 0.266356f
C4563 a_n6972_8799.t73 gnd 0.597459f
C4564 a_n6972_8799.n159 gnd 0.261873f
C4565 a_n6972_8799.t55 gnd 0.597459f
C4566 a_n6972_8799.n160 gnd 0.270403f
C4567 a_n6972_8799.t59 gnd 0.608756f
C4568 a_n6972_8799.n161 gnd 0.899839f
C4569 a_n6972_8799.t91 gnd 0.597459f
C4570 a_n6972_8799.n162 gnd 0.267109f
C4571 a_n6972_8799.t111 gnd 0.597459f
C4572 a_n6972_8799.t44 gnd 0.597459f
C4573 a_n6972_8799.n163 gnd 0.270418f
C4574 a_n6972_8799.t97 gnd 0.597459f
C4575 a_n6972_8799.t127 gnd 0.597459f
C4576 a_n6972_8799.t88 gnd 0.597459f
C4577 a_n6972_8799.n164 gnd 0.272502f
C4578 a_n6972_8799.t121 gnd 0.597459f
C4579 a_n6972_8799.t54 gnd 0.597459f
C4580 a_n6972_8799.n165 gnd 0.266036f
C4581 a_n6972_8799.t118 gnd 0.608767f
C4582 a_n6972_8799.n166 gnd 0.250481f
C4583 a_n6972_8799.n167 gnd 0.011785f
C4584 a_n6972_8799.t39 gnd 0.597459f
C4585 a_n6972_8799.n168 gnd 0.266836f
C4586 a_n6972_8799.n169 gnd 0.270404f
C4587 a_n6972_8799.t103 gnd 0.597459f
C4588 a_n6972_8799.n170 gnd 0.266926f
C4589 a_n6972_8799.n171 gnd 0.261553f
C4590 a_n6972_8799.t82 gnd 0.597459f
C4591 a_n6972_8799.n172 gnd 0.266676f
C4592 a_n6972_8799.n173 gnd 0.272936f
C4593 a_n6972_8799.t60 gnd 0.597459f
C4594 a_n6972_8799.n174 gnd 0.270286f
C4595 a_n6972_8799.n175 gnd 0.266356f
C4596 a_n6972_8799.t67 gnd 0.597459f
C4597 a_n6972_8799.n176 gnd 0.261873f
C4598 a_n6972_8799.t50 gnd 0.597459f
C4599 a_n6972_8799.n177 gnd 0.270403f
C4600 a_n6972_8799.t131 gnd 0.608756f
C4601 a_n6972_8799.n178 gnd 1.53901f
C4602 a_n6972_8799.t80 gnd 0.597459f
C4603 a_n6972_8799.t79 gnd 0.597459f
C4604 a_n6972_8799.t58 gnd 0.597459f
C4605 a_n6972_8799.n179 gnd 0.270005f
C4606 a_n6972_8799.t116 gnd 0.597459f
C4607 a_n6972_8799.t81 gnd 0.597459f
C4608 a_n6972_8799.t63 gnd 0.597459f
C4609 a_n6972_8799.n180 gnd 0.266926f
C4610 a_n6972_8799.t119 gnd 0.597459f
C4611 a_n6972_8799.t95 gnd 0.597459f
C4612 a_n6972_8799.t93 gnd 0.597459f
C4613 a_n6972_8799.n181 gnd 0.270418f
C4614 a_n6972_8799.t40 gnd 0.597459f
C4615 a_n6972_8799.t99 gnd 0.597459f
C4616 a_n6972_8799.t98 gnd 0.597459f
C4617 a_n6972_8799.n182 gnd 0.266356f
C4618 a_n6972_8799.t42 gnd 0.597459f
C4619 a_n6972_8799.t41 gnd 0.597459f
C4620 a_n6972_8799.t112 gnd 0.597459f
C4621 a_n6972_8799.n183 gnd 0.270403f
C4622 a_n6972_8799.t57 gnd 0.608767f
C4623 a_n6972_8799.n184 gnd 0.250481f
C4624 a_n6972_8799.n185 gnd 0.267109f
C4625 a_n6972_8799.n186 gnd 0.261873f
C4626 a_n6972_8799.n187 gnd 0.270286f
C4627 a_n6972_8799.n188 gnd 0.272936f
C4628 a_n6972_8799.n189 gnd 0.266676f
C4629 a_n6972_8799.n190 gnd 0.261553f
C4630 a_n6972_8799.n191 gnd 0.270404f
C4631 a_n6972_8799.n192 gnd 0.272502f
C4632 a_n6972_8799.n193 gnd 0.266036f
C4633 a_n6972_8799.n194 gnd 0.261393f
C4634 a_n6972_8799.t87 gnd 0.597459f
C4635 a_n6972_8799.t86 gnd 0.597459f
C4636 a_n6972_8799.t70 gnd 0.597459f
C4637 a_n6972_8799.n195 gnd 0.270005f
C4638 a_n6972_8799.t128 gnd 0.597459f
C4639 a_n6972_8799.t92 gnd 0.597459f
C4640 a_n6972_8799.t72 gnd 0.597459f
C4641 a_n6972_8799.n196 gnd 0.266926f
C4642 a_n6972_8799.t36 gnd 0.597459f
C4643 a_n6972_8799.t105 gnd 0.597459f
C4644 a_n6972_8799.t104 gnd 0.597459f
C4645 a_n6972_8799.n197 gnd 0.270418f
C4646 a_n6972_8799.t49 gnd 0.597459f
C4647 a_n6972_8799.t108 gnd 0.597459f
C4648 a_n6972_8799.t107 gnd 0.597459f
C4649 a_n6972_8799.n198 gnd 0.266356f
C4650 a_n6972_8799.t53 gnd 0.597459f
C4651 a_n6972_8799.t52 gnd 0.597459f
C4652 a_n6972_8799.t123 gnd 0.597459f
C4653 a_n6972_8799.n199 gnd 0.270403f
C4654 a_n6972_8799.t71 gnd 0.608767f
C4655 a_n6972_8799.n200 gnd 0.250481f
C4656 a_n6972_8799.n201 gnd 0.267109f
C4657 a_n6972_8799.n202 gnd 0.261873f
C4658 a_n6972_8799.n203 gnd 0.270286f
C4659 a_n6972_8799.n204 gnd 0.272936f
C4660 a_n6972_8799.n205 gnd 0.266676f
C4661 a_n6972_8799.n206 gnd 0.261553f
C4662 a_n6972_8799.n207 gnd 0.270404f
C4663 a_n6972_8799.n208 gnd 0.272502f
C4664 a_n6972_8799.n209 gnd 0.266036f
C4665 a_n6972_8799.n210 gnd 0.261393f
C4666 a_n6972_8799.n211 gnd 0.899839f
C4667 a_n6972_8799.t130 gnd 0.597459f
C4668 a_n6972_8799.t51 gnd 0.597459f
C4669 a_n6972_8799.t90 gnd 0.597459f
C4670 a_n6972_8799.n212 gnd 0.270005f
C4671 a_n6972_8799.t38 gnd 0.597459f
C4672 a_n6972_8799.t110 gnd 0.597459f
C4673 a_n6972_8799.t62 gnd 0.597459f
C4674 a_n6972_8799.n213 gnd 0.266926f
C4675 a_n6972_8799.t96 gnd 0.597459f
C4676 a_n6972_8799.t43 gnd 0.597459f
C4677 a_n6972_8799.t66 gnd 0.597459f
C4678 a_n6972_8799.n214 gnd 0.270418f
C4679 a_n6972_8799.t126 gnd 0.597459f
C4680 a_n6972_8799.t102 gnd 0.597459f
C4681 a_n6972_8799.t122 gnd 0.597459f
C4682 a_n6972_8799.n215 gnd 0.266356f
C4683 a_n6972_8799.t89 gnd 0.597459f
C4684 a_n6972_8799.t106 gnd 0.597459f
C4685 a_n6972_8799.t56 gnd 0.597459f
C4686 a_n6972_8799.n216 gnd 0.270403f
C4687 a_n6972_8799.t120 gnd 0.608767f
C4688 a_n6972_8799.n217 gnd 0.250481f
C4689 a_n6972_8799.n218 gnd 0.267109f
C4690 a_n6972_8799.n219 gnd 0.261873f
C4691 a_n6972_8799.n220 gnd 0.270286f
C4692 a_n6972_8799.n221 gnd 0.272936f
C4693 a_n6972_8799.n222 gnd 0.266676f
C4694 a_n6972_8799.n223 gnd 0.261553f
C4695 a_n6972_8799.n224 gnd 0.270404f
C4696 a_n6972_8799.n225 gnd 0.272502f
C4697 a_n6972_8799.n226 gnd 0.266036f
C4698 a_n6972_8799.n227 gnd 0.261393f
C4699 a_n6972_8799.n228 gnd 1.08613f
C4700 a_n6972_8799.n229 gnd 12.2028f
C4701 a_n6972_8799.n230 gnd 4.37253f
C4702 a_n6972_8799.n231 gnd 5.6731f
C4703 a_n6972_8799.t14 gnd 0.144089f
C4704 a_n6972_8799.t21 gnd 0.144089f
C4705 a_n6972_8799.n232 gnd 1.13457f
C4706 a_n6972_8799.n233 gnd 1.13458f
C4707 a_n6972_8799.t2 gnd 0.144089f
C4708 CSoutput.n0 gnd 0.044705f
C4709 CSoutput.t154 gnd 0.295714f
C4710 CSoutput.n1 gnd 0.133529f
C4711 CSoutput.n2 gnd 0.044705f
C4712 CSoutput.t159 gnd 0.295714f
C4713 CSoutput.n3 gnd 0.035432f
C4714 CSoutput.n4 gnd 0.044705f
C4715 CSoutput.t148 gnd 0.295714f
C4716 CSoutput.n5 gnd 0.030554f
C4717 CSoutput.n6 gnd 0.044705f
C4718 CSoutput.t156 gnd 0.295714f
C4719 CSoutput.t162 gnd 0.295714f
C4720 CSoutput.n7 gnd 0.132074f
C4721 CSoutput.n8 gnd 0.044705f
C4722 CSoutput.t161 gnd 0.295714f
C4723 CSoutput.n9 gnd 0.029131f
C4724 CSoutput.n10 gnd 0.044705f
C4725 CSoutput.t149 gnd 0.295714f
C4726 CSoutput.t160 gnd 0.295714f
C4727 CSoutput.n11 gnd 0.132074f
C4728 CSoutput.n12 gnd 0.044705f
C4729 CSoutput.t158 gnd 0.295714f
C4730 CSoutput.n13 gnd 0.030554f
C4731 CSoutput.n14 gnd 0.044705f
C4732 CSoutput.t147 gnd 0.295714f
C4733 CSoutput.t151 gnd 0.295714f
C4734 CSoutput.n15 gnd 0.132074f
C4735 CSoutput.n16 gnd 0.044705f
C4736 CSoutput.t155 gnd 0.295714f
C4737 CSoutput.n17 gnd 0.032633f
C4738 CSoutput.t165 gnd 0.353386f
C4739 CSoutput.t145 gnd 0.295714f
C4740 CSoutput.n18 gnd 0.168607f
C4741 CSoutput.n19 gnd 0.163607f
C4742 CSoutput.n20 gnd 0.189804f
C4743 CSoutput.n21 gnd 0.044705f
C4744 CSoutput.n22 gnd 0.037311f
C4745 CSoutput.n23 gnd 0.132074f
C4746 CSoutput.n24 gnd 0.035967f
C4747 CSoutput.n25 gnd 0.035432f
C4748 CSoutput.n26 gnd 0.044705f
C4749 CSoutput.n27 gnd 0.044705f
C4750 CSoutput.n28 gnd 0.037024f
C4751 CSoutput.n29 gnd 0.031435f
C4752 CSoutput.n30 gnd 0.135014f
C4753 CSoutput.n31 gnd 0.031868f
C4754 CSoutput.n32 gnd 0.044705f
C4755 CSoutput.n33 gnd 0.044705f
C4756 CSoutput.n34 gnd 0.044705f
C4757 CSoutput.n35 gnd 0.03663f
C4758 CSoutput.n36 gnd 0.132074f
C4759 CSoutput.n37 gnd 0.035031f
C4760 CSoutput.n38 gnd 0.036368f
C4761 CSoutput.n39 gnd 0.044705f
C4762 CSoutput.n40 gnd 0.044705f
C4763 CSoutput.n41 gnd 0.037304f
C4764 CSoutput.n42 gnd 0.034096f
C4765 CSoutput.n43 gnd 0.132074f
C4766 CSoutput.n44 gnd 0.03496f
C4767 CSoutput.n45 gnd 0.044705f
C4768 CSoutput.n46 gnd 0.044705f
C4769 CSoutput.n47 gnd 0.044705f
C4770 CSoutput.n48 gnd 0.03496f
C4771 CSoutput.n49 gnd 0.132074f
C4772 CSoutput.n50 gnd 0.034096f
C4773 CSoutput.n51 gnd 0.037304f
C4774 CSoutput.n52 gnd 0.044705f
C4775 CSoutput.n53 gnd 0.044705f
C4776 CSoutput.n54 gnd 0.036368f
C4777 CSoutput.n55 gnd 0.035031f
C4778 CSoutput.n56 gnd 0.132074f
C4779 CSoutput.n57 gnd 0.03663f
C4780 CSoutput.n58 gnd 0.044705f
C4781 CSoutput.n59 gnd 0.044705f
C4782 CSoutput.n60 gnd 0.044705f
C4783 CSoutput.n61 gnd 0.031868f
C4784 CSoutput.n62 gnd 0.135014f
C4785 CSoutput.n63 gnd 0.031435f
C4786 CSoutput.t164 gnd 0.295714f
C4787 CSoutput.n64 gnd 0.132074f
C4788 CSoutput.n65 gnd 0.037024f
C4789 CSoutput.n66 gnd 0.044705f
C4790 CSoutput.n67 gnd 0.044705f
C4791 CSoutput.n68 gnd 0.044705f
C4792 CSoutput.n69 gnd 0.035967f
C4793 CSoutput.n70 gnd 0.132074f
C4794 CSoutput.n71 gnd 0.037311f
C4795 CSoutput.n72 gnd 0.032633f
C4796 CSoutput.n73 gnd 0.044705f
C4797 CSoutput.n74 gnd 0.044705f
C4798 CSoutput.n75 gnd 0.033843f
C4799 CSoutput.n76 gnd 0.020099f
C4800 CSoutput.t144 gnd 0.332255f
C4801 CSoutput.n77 gnd 0.165051f
C4802 CSoutput.n78 gnd 0.706239f
C4803 CSoutput.t2 gnd 0.055763f
C4804 CSoutput.t13 gnd 0.055763f
C4805 CSoutput.n79 gnd 0.431737f
C4806 CSoutput.t40 gnd 0.055763f
C4807 CSoutput.t55 gnd 0.055763f
C4808 CSoutput.n80 gnd 0.430967f
C4809 CSoutput.n81 gnd 0.437431f
C4810 CSoutput.t34 gnd 0.055763f
C4811 CSoutput.t33 gnd 0.055763f
C4812 CSoutput.n82 gnd 0.430967f
C4813 CSoutput.n83 gnd 0.215548f
C4814 CSoutput.t0 gnd 0.055763f
C4815 CSoutput.t57 gnd 0.055763f
C4816 CSoutput.n84 gnd 0.430967f
C4817 CSoutput.n85 gnd 0.215548f
C4818 CSoutput.t62 gnd 0.055763f
C4819 CSoutput.t35 gnd 0.055763f
C4820 CSoutput.n86 gnd 0.430967f
C4821 CSoutput.n87 gnd 0.215548f
C4822 CSoutput.t12 gnd 0.055763f
C4823 CSoutput.t3 gnd 0.055763f
C4824 CSoutput.n88 gnd 0.430967f
C4825 CSoutput.n89 gnd 0.215548f
C4826 CSoutput.t44 gnd 0.055763f
C4827 CSoutput.t17 gnd 0.055763f
C4828 CSoutput.n90 gnd 0.430967f
C4829 CSoutput.n91 gnd 0.215548f
C4830 CSoutput.t64 gnd 0.055763f
C4831 CSoutput.t130 gnd 0.055763f
C4832 CSoutput.n92 gnd 0.430967f
C4833 CSoutput.n93 gnd 0.395264f
C4834 CSoutput.t22 gnd 0.055763f
C4835 CSoutput.t23 gnd 0.055763f
C4836 CSoutput.n94 gnd 0.431737f
C4837 CSoutput.t28 gnd 0.055763f
C4838 CSoutput.t136 gnd 0.055763f
C4839 CSoutput.n95 gnd 0.430967f
C4840 CSoutput.n96 gnd 0.437431f
C4841 CSoutput.t18 gnd 0.055763f
C4842 CSoutput.t133 gnd 0.055763f
C4843 CSoutput.n97 gnd 0.430967f
C4844 CSoutput.n98 gnd 0.215548f
C4845 CSoutput.t143 gnd 0.055763f
C4846 CSoutput.t73 gnd 0.055763f
C4847 CSoutput.n99 gnd 0.430967f
C4848 CSoutput.n100 gnd 0.215548f
C4849 CSoutput.t7 gnd 0.055763f
C4850 CSoutput.t128 gnd 0.055763f
C4851 CSoutput.n101 gnd 0.430967f
C4852 CSoutput.n102 gnd 0.215548f
C4853 CSoutput.t49 gnd 0.055763f
C4854 CSoutput.t30 gnd 0.055763f
C4855 CSoutput.n103 gnd 0.430967f
C4856 CSoutput.n104 gnd 0.215548f
C4857 CSoutput.t36 gnd 0.055763f
C4858 CSoutput.t15 gnd 0.055763f
C4859 CSoutput.n105 gnd 0.430967f
C4860 CSoutput.n106 gnd 0.215548f
C4861 CSoutput.t60 gnd 0.055763f
C4862 CSoutput.t59 gnd 0.055763f
C4863 CSoutput.n107 gnd 0.430967f
C4864 CSoutput.n108 gnd 0.321436f
C4865 CSoutput.n109 gnd 0.405328f
C4866 CSoutput.t42 gnd 0.055763f
C4867 CSoutput.t67 gnd 0.055763f
C4868 CSoutput.n110 gnd 0.431737f
C4869 CSoutput.t29 gnd 0.055763f
C4870 CSoutput.t139 gnd 0.055763f
C4871 CSoutput.n111 gnd 0.430967f
C4872 CSoutput.n112 gnd 0.437431f
C4873 CSoutput.t5 gnd 0.055763f
C4874 CSoutput.t24 gnd 0.055763f
C4875 CSoutput.n113 gnd 0.430967f
C4876 CSoutput.n114 gnd 0.215548f
C4877 CSoutput.t141 gnd 0.055763f
C4878 CSoutput.t142 gnd 0.055763f
C4879 CSoutput.n115 gnd 0.430967f
C4880 CSoutput.n116 gnd 0.215548f
C4881 CSoutput.t72 gnd 0.055763f
C4882 CSoutput.t76 gnd 0.055763f
C4883 CSoutput.n117 gnd 0.430967f
C4884 CSoutput.n118 gnd 0.215548f
C4885 CSoutput.t54 gnd 0.055763f
C4886 CSoutput.t58 gnd 0.055763f
C4887 CSoutput.n119 gnd 0.430967f
C4888 CSoutput.n120 gnd 0.215548f
C4889 CSoutput.t138 gnd 0.055763f
C4890 CSoutput.t9 gnd 0.055763f
C4891 CSoutput.n121 gnd 0.430967f
C4892 CSoutput.n122 gnd 0.215548f
C4893 CSoutput.t61 gnd 0.055763f
C4894 CSoutput.t32 gnd 0.055763f
C4895 CSoutput.n123 gnd 0.430967f
C4896 CSoutput.n124 gnd 0.321436f
C4897 CSoutput.n125 gnd 0.453053f
C4898 CSoutput.n126 gnd 7.74234f
C4899 CSoutput.n128 gnd 0.790823f
C4900 CSoutput.n129 gnd 0.593117f
C4901 CSoutput.n130 gnd 0.790823f
C4902 CSoutput.n131 gnd 0.790823f
C4903 CSoutput.n132 gnd 2.12914f
C4904 CSoutput.n133 gnd 0.790823f
C4905 CSoutput.n134 gnd 0.790823f
C4906 CSoutput.t163 gnd 0.988529f
C4907 CSoutput.n135 gnd 0.790823f
C4908 CSoutput.n136 gnd 0.790823f
C4909 CSoutput.n140 gnd 0.790823f
C4910 CSoutput.n144 gnd 0.790823f
C4911 CSoutput.n145 gnd 0.790823f
C4912 CSoutput.n147 gnd 0.790823f
C4913 CSoutput.n152 gnd 0.790823f
C4914 CSoutput.n154 gnd 0.790823f
C4915 CSoutput.n155 gnd 0.790823f
C4916 CSoutput.n157 gnd 0.790823f
C4917 CSoutput.n158 gnd 0.790823f
C4918 CSoutput.n160 gnd 0.790823f
C4919 CSoutput.t152 gnd 13.2146f
C4920 CSoutput.n162 gnd 0.790823f
C4921 CSoutput.n163 gnd 0.593117f
C4922 CSoutput.n164 gnd 0.790823f
C4923 CSoutput.n165 gnd 0.790823f
C4924 CSoutput.n166 gnd 2.12914f
C4925 CSoutput.n167 gnd 0.790823f
C4926 CSoutput.n168 gnd 0.790823f
C4927 CSoutput.t150 gnd 0.988529f
C4928 CSoutput.n169 gnd 0.790823f
C4929 CSoutput.n170 gnd 0.790823f
C4930 CSoutput.n174 gnd 0.790823f
C4931 CSoutput.n178 gnd 0.790823f
C4932 CSoutput.n179 gnd 0.790823f
C4933 CSoutput.n181 gnd 0.790823f
C4934 CSoutput.n186 gnd 0.790823f
C4935 CSoutput.n188 gnd 0.790823f
C4936 CSoutput.n189 gnd 0.790823f
C4937 CSoutput.n191 gnd 0.790823f
C4938 CSoutput.n192 gnd 0.790823f
C4939 CSoutput.n194 gnd 0.790823f
C4940 CSoutput.n195 gnd 0.593117f
C4941 CSoutput.n197 gnd 0.790823f
C4942 CSoutput.n198 gnd 0.593117f
C4943 CSoutput.n199 gnd 0.790823f
C4944 CSoutput.n200 gnd 0.790823f
C4945 CSoutput.n201 gnd 2.12914f
C4946 CSoutput.n202 gnd 0.790823f
C4947 CSoutput.n203 gnd 0.790823f
C4948 CSoutput.t146 gnd 0.988529f
C4949 CSoutput.n204 gnd 0.790823f
C4950 CSoutput.n205 gnd 2.12914f
C4951 CSoutput.n207 gnd 0.790823f
C4952 CSoutput.n208 gnd 0.790823f
C4953 CSoutput.n210 gnd 0.790823f
C4954 CSoutput.n211 gnd 0.790823f
C4955 CSoutput.t153 gnd 12.9992f
C4956 CSoutput.t157 gnd 13.2146f
C4957 CSoutput.n217 gnd 2.48093f
C4958 CSoutput.n218 gnd 10.1064f
C4959 CSoutput.n219 gnd 10.5293f
C4960 CSoutput.n224 gnd 2.68751f
C4961 CSoutput.n230 gnd 0.790823f
C4962 CSoutput.n232 gnd 0.790823f
C4963 CSoutput.n234 gnd 0.790823f
C4964 CSoutput.n236 gnd 0.790823f
C4965 CSoutput.n238 gnd 0.790823f
C4966 CSoutput.n244 gnd 0.790823f
C4967 CSoutput.n251 gnd 1.45086f
C4968 CSoutput.n252 gnd 1.45086f
C4969 CSoutput.n253 gnd 0.790823f
C4970 CSoutput.n254 gnd 0.790823f
C4971 CSoutput.n256 gnd 0.593117f
C4972 CSoutput.n257 gnd 0.507952f
C4973 CSoutput.n259 gnd 0.593117f
C4974 CSoutput.n260 gnd 0.507952f
C4975 CSoutput.n261 gnd 0.593117f
C4976 CSoutput.n263 gnd 0.790823f
C4977 CSoutput.n265 gnd 2.12914f
C4978 CSoutput.n266 gnd 2.48093f
C4979 CSoutput.n267 gnd 9.29529f
C4980 CSoutput.n269 gnd 0.593117f
C4981 CSoutput.n270 gnd 1.52613f
C4982 CSoutput.n271 gnd 0.593117f
C4983 CSoutput.n273 gnd 0.790823f
C4984 CSoutput.n275 gnd 2.12914f
C4985 CSoutput.n276 gnd 4.63761f
C4986 CSoutput.t26 gnd 0.055763f
C4987 CSoutput.t78 gnd 0.055763f
C4988 CSoutput.n277 gnd 0.431737f
C4989 CSoutput.t8 gnd 0.055763f
C4990 CSoutput.t56 gnd 0.055763f
C4991 CSoutput.n278 gnd 0.430967f
C4992 CSoutput.n279 gnd 0.437431f
C4993 CSoutput.t14 gnd 0.055763f
C4994 CSoutput.t50 gnd 0.055763f
C4995 CSoutput.n280 gnd 0.430967f
C4996 CSoutput.n281 gnd 0.215548f
C4997 CSoutput.t38 gnd 0.055763f
C4998 CSoutput.t74 gnd 0.055763f
C4999 CSoutput.n282 gnd 0.430967f
C5000 CSoutput.n283 gnd 0.215548f
C5001 CSoutput.t51 gnd 0.055763f
C5002 CSoutput.t16 gnd 0.055763f
C5003 CSoutput.n284 gnd 0.430967f
C5004 CSoutput.n285 gnd 0.215548f
C5005 CSoutput.t1 gnd 0.055763f
C5006 CSoutput.t66 gnd 0.055763f
C5007 CSoutput.n286 gnd 0.430967f
C5008 CSoutput.n287 gnd 0.215548f
C5009 CSoutput.t43 gnd 0.055763f
C5010 CSoutput.t31 gnd 0.055763f
C5011 CSoutput.n288 gnd 0.430967f
C5012 CSoutput.n289 gnd 0.215548f
C5013 CSoutput.t131 gnd 0.055763f
C5014 CSoutput.t65 gnd 0.055763f
C5015 CSoutput.n290 gnd 0.430967f
C5016 CSoutput.n291 gnd 0.395264f
C5017 CSoutput.t41 gnd 0.055763f
C5018 CSoutput.t37 gnd 0.055763f
C5019 CSoutput.n292 gnd 0.431737f
C5020 CSoutput.t45 gnd 0.055763f
C5021 CSoutput.t48 gnd 0.055763f
C5022 CSoutput.n293 gnd 0.430967f
C5023 CSoutput.n294 gnd 0.437431f
C5024 CSoutput.t11 gnd 0.055763f
C5025 CSoutput.t79 gnd 0.055763f
C5026 CSoutput.n295 gnd 0.430967f
C5027 CSoutput.n296 gnd 0.215548f
C5028 CSoutput.t63 gnd 0.055763f
C5029 CSoutput.t75 gnd 0.055763f
C5030 CSoutput.n297 gnd 0.430967f
C5031 CSoutput.n298 gnd 0.215548f
C5032 CSoutput.t132 gnd 0.055763f
C5033 CSoutput.t4 gnd 0.055763f
C5034 CSoutput.n299 gnd 0.430967f
C5035 CSoutput.n300 gnd 0.215548f
C5036 CSoutput.t6 gnd 0.055763f
C5037 CSoutput.t21 gnd 0.055763f
C5038 CSoutput.n301 gnd 0.430967f
C5039 CSoutput.n302 gnd 0.215548f
C5040 CSoutput.t129 gnd 0.055763f
C5041 CSoutput.t71 gnd 0.055763f
C5042 CSoutput.n303 gnd 0.430967f
C5043 CSoutput.n304 gnd 0.215548f
C5044 CSoutput.t25 gnd 0.055763f
C5045 CSoutput.t77 gnd 0.055763f
C5046 CSoutput.n305 gnd 0.430967f
C5047 CSoutput.n306 gnd 0.321436f
C5048 CSoutput.n307 gnd 0.405328f
C5049 CSoutput.t137 gnd 0.055763f
C5050 CSoutput.t46 gnd 0.055763f
C5051 CSoutput.n308 gnd 0.431737f
C5052 CSoutput.t10 gnd 0.055763f
C5053 CSoutput.t52 gnd 0.055763f
C5054 CSoutput.n309 gnd 0.430967f
C5055 CSoutput.n310 gnd 0.437431f
C5056 CSoutput.t27 gnd 0.055763f
C5057 CSoutput.t39 gnd 0.055763f
C5058 CSoutput.n311 gnd 0.430967f
C5059 CSoutput.n312 gnd 0.215548f
C5060 CSoutput.t68 gnd 0.055763f
C5061 CSoutput.t19 gnd 0.055763f
C5062 CSoutput.n313 gnd 0.430967f
C5063 CSoutput.n314 gnd 0.215548f
C5064 CSoutput.t70 gnd 0.055763f
C5065 CSoutput.t20 gnd 0.055763f
C5066 CSoutput.n315 gnd 0.430967f
C5067 CSoutput.n316 gnd 0.215548f
C5068 CSoutput.t53 gnd 0.055763f
C5069 CSoutput.t140 gnd 0.055763f
C5070 CSoutput.n317 gnd 0.430967f
C5071 CSoutput.n318 gnd 0.215548f
C5072 CSoutput.t134 gnd 0.055763f
C5073 CSoutput.t69 gnd 0.055763f
C5074 CSoutput.n319 gnd 0.430967f
C5075 CSoutput.n320 gnd 0.215548f
C5076 CSoutput.t47 gnd 0.055763f
C5077 CSoutput.t135 gnd 0.055763f
C5078 CSoutput.n321 gnd 0.430965f
C5079 CSoutput.n322 gnd 0.321437f
C5080 CSoutput.n323 gnd 0.453053f
C5081 CSoutput.n324 gnd 11.346299f
C5082 CSoutput.t104 gnd 0.048793f
C5083 CSoutput.t94 gnd 0.048793f
C5084 CSoutput.n325 gnd 0.432593f
C5085 CSoutput.t120 gnd 0.048793f
C5086 CSoutput.t122 gnd 0.048793f
C5087 CSoutput.n326 gnd 0.43115f
C5088 CSoutput.n327 gnd 0.401751f
C5089 CSoutput.t99 gnd 0.048793f
C5090 CSoutput.t89 gnd 0.048793f
C5091 CSoutput.n328 gnd 0.43115f
C5092 CSoutput.n329 gnd 0.198044f
C5093 CSoutput.t125 gnd 0.048793f
C5094 CSoutput.t106 gnd 0.048793f
C5095 CSoutput.n330 gnd 0.43115f
C5096 CSoutput.n331 gnd 0.198044f
C5097 CSoutput.t108 gnd 0.048793f
C5098 CSoutput.t97 gnd 0.048793f
C5099 CSoutput.n332 gnd 0.43115f
C5100 CSoutput.n333 gnd 0.198044f
C5101 CSoutput.t111 gnd 0.048793f
C5102 CSoutput.t113 gnd 0.048793f
C5103 CSoutput.n334 gnd 0.43115f
C5104 CSoutput.n335 gnd 0.365234f
C5105 CSoutput.t114 gnd 0.048793f
C5106 CSoutput.t103 gnd 0.048793f
C5107 CSoutput.n336 gnd 0.432593f
C5108 CSoutput.t126 gnd 0.048793f
C5109 CSoutput.t80 gnd 0.048793f
C5110 CSoutput.n337 gnd 0.43115f
C5111 CSoutput.n338 gnd 0.401751f
C5112 CSoutput.t109 gnd 0.048793f
C5113 CSoutput.t98 gnd 0.048793f
C5114 CSoutput.n339 gnd 0.43115f
C5115 CSoutput.n340 gnd 0.198044f
C5116 CSoutput.t84 gnd 0.048793f
C5117 CSoutput.t115 gnd 0.048793f
C5118 CSoutput.n341 gnd 0.43115f
C5119 CSoutput.n342 gnd 0.198044f
C5120 CSoutput.t117 gnd 0.048793f
C5121 CSoutput.t107 gnd 0.048793f
C5122 CSoutput.n343 gnd 0.43115f
C5123 CSoutput.n344 gnd 0.198044f
C5124 CSoutput.t118 gnd 0.048793f
C5125 CSoutput.t121 gnd 0.048793f
C5126 CSoutput.n345 gnd 0.43115f
C5127 CSoutput.n346 gnd 0.300674f
C5128 CSoutput.n347 gnd 0.558675f
C5129 CSoutput.n348 gnd 11.651f
C5130 CSoutput.t83 gnd 0.048793f
C5131 CSoutput.t91 gnd 0.048793f
C5132 CSoutput.n349 gnd 0.432593f
C5133 CSoutput.t112 gnd 0.048793f
C5134 CSoutput.t124 gnd 0.048793f
C5135 CSoutput.n350 gnd 0.43115f
C5136 CSoutput.n351 gnd 0.401751f
C5137 CSoutput.t127 gnd 0.048793f
C5138 CSoutput.t87 gnd 0.048793f
C5139 CSoutput.n352 gnd 0.43115f
C5140 CSoutput.n353 gnd 0.198044f
C5141 CSoutput.t92 gnd 0.048793f
C5142 CSoutput.t81 gnd 0.048793f
C5143 CSoutput.n354 gnd 0.43115f
C5144 CSoutput.n355 gnd 0.198044f
C5145 CSoutput.t85 gnd 0.048793f
C5146 CSoutput.t95 gnd 0.048793f
C5147 CSoutput.n356 gnd 0.43115f
C5148 CSoutput.n357 gnd 0.198044f
C5149 CSoutput.t100 gnd 0.048793f
C5150 CSoutput.t116 gnd 0.048793f
C5151 CSoutput.n358 gnd 0.43115f
C5152 CSoutput.n359 gnd 0.365234f
C5153 CSoutput.t90 gnd 0.048793f
C5154 CSoutput.t102 gnd 0.048793f
C5155 CSoutput.n360 gnd 0.432593f
C5156 CSoutput.t119 gnd 0.048793f
C5157 CSoutput.t82 gnd 0.048793f
C5158 CSoutput.n361 gnd 0.43115f
C5159 CSoutput.n362 gnd 0.401751f
C5160 CSoutput.t86 gnd 0.048793f
C5161 CSoutput.t96 gnd 0.048793f
C5162 CSoutput.n363 gnd 0.43115f
C5163 CSoutput.n364 gnd 0.198044f
C5164 CSoutput.t101 gnd 0.048793f
C5165 CSoutput.t88 gnd 0.048793f
C5166 CSoutput.n365 gnd 0.43115f
C5167 CSoutput.n366 gnd 0.198044f
C5168 CSoutput.t93 gnd 0.048793f
C5169 CSoutput.t105 gnd 0.048793f
C5170 CSoutput.n367 gnd 0.43115f
C5171 CSoutput.n368 gnd 0.198044f
C5172 CSoutput.t110 gnd 0.048793f
C5173 CSoutput.t123 gnd 0.048793f
C5174 CSoutput.n369 gnd 0.43115f
C5175 CSoutput.n370 gnd 0.300674f
C5176 CSoutput.n371 gnd 0.558675f
C5177 CSoutput.n372 gnd 6.50657f
C5178 CSoutput.n373 gnd 14.331701f
C5179 commonsourceibias.n0 gnd 0.010301f
C5180 commonsourceibias.t71 gnd 0.155981f
C5181 commonsourceibias.t81 gnd 0.144227f
C5182 commonsourceibias.n1 gnd 0.057546f
C5183 commonsourceibias.n2 gnd 0.00772f
C5184 commonsourceibias.t55 gnd 0.144227f
C5185 commonsourceibias.n3 gnd 0.006245f
C5186 commonsourceibias.n4 gnd 0.00772f
C5187 commonsourceibias.t53 gnd 0.144227f
C5188 commonsourceibias.n5 gnd 0.007453f
C5189 commonsourceibias.n6 gnd 0.00772f
C5190 commonsourceibias.t76 gnd 0.144227f
C5191 commonsourceibias.n7 gnd 0.057546f
C5192 commonsourceibias.t86 gnd 0.144227f
C5193 commonsourceibias.n8 gnd 0.006235f
C5194 commonsourceibias.n9 gnd 0.010301f
C5195 commonsourceibias.t32 gnd 0.155981f
C5196 commonsourceibias.t14 gnd 0.144227f
C5197 commonsourceibias.n10 gnd 0.057546f
C5198 commonsourceibias.n11 gnd 0.00772f
C5199 commonsourceibias.t24 gnd 0.144227f
C5200 commonsourceibias.n12 gnd 0.006245f
C5201 commonsourceibias.n13 gnd 0.00772f
C5202 commonsourceibias.t30 gnd 0.144227f
C5203 commonsourceibias.n14 gnd 0.007453f
C5204 commonsourceibias.n15 gnd 0.00772f
C5205 commonsourceibias.t20 gnd 0.144227f
C5206 commonsourceibias.n16 gnd 0.057546f
C5207 commonsourceibias.t36 gnd 0.144227f
C5208 commonsourceibias.n17 gnd 0.006235f
C5209 commonsourceibias.n18 gnd 0.00772f
C5210 commonsourceibias.t44 gnd 0.144227f
C5211 commonsourceibias.t26 gnd 0.144227f
C5212 commonsourceibias.n19 gnd 0.057546f
C5213 commonsourceibias.n20 gnd 0.00772f
C5214 commonsourceibias.t34 gnd 0.144227f
C5215 commonsourceibias.n21 gnd 0.057546f
C5216 commonsourceibias.n22 gnd 0.00772f
C5217 commonsourceibias.t10 gnd 0.144227f
C5218 commonsourceibias.n23 gnd 0.057546f
C5219 commonsourceibias.n24 gnd 0.038863f
C5220 commonsourceibias.t40 gnd 0.144227f
C5221 commonsourceibias.t46 gnd 0.162743f
C5222 commonsourceibias.n25 gnd 0.066782f
C5223 commonsourceibias.n26 gnd 0.069137f
C5224 commonsourceibias.n27 gnd 0.009515f
C5225 commonsourceibias.n28 gnd 0.010526f
C5226 commonsourceibias.n29 gnd 0.00772f
C5227 commonsourceibias.n30 gnd 0.00772f
C5228 commonsourceibias.n31 gnd 0.010457f
C5229 commonsourceibias.n32 gnd 0.006245f
C5230 commonsourceibias.n33 gnd 0.010587f
C5231 commonsourceibias.n34 gnd 0.00772f
C5232 commonsourceibias.n35 gnd 0.00772f
C5233 commonsourceibias.n36 gnd 0.010651f
C5234 commonsourceibias.n37 gnd 0.009185f
C5235 commonsourceibias.n38 gnd 0.007453f
C5236 commonsourceibias.n39 gnd 0.00772f
C5237 commonsourceibias.n40 gnd 0.00772f
C5238 commonsourceibias.n41 gnd 0.009442f
C5239 commonsourceibias.n42 gnd 0.010598f
C5240 commonsourceibias.n43 gnd 0.057546f
C5241 commonsourceibias.n44 gnd 0.010527f
C5242 commonsourceibias.n45 gnd 0.00772f
C5243 commonsourceibias.n46 gnd 0.00772f
C5244 commonsourceibias.n47 gnd 0.00772f
C5245 commonsourceibias.n48 gnd 0.010527f
C5246 commonsourceibias.n49 gnd 0.057546f
C5247 commonsourceibias.n50 gnd 0.010598f
C5248 commonsourceibias.n51 gnd 0.009442f
C5249 commonsourceibias.n52 gnd 0.00772f
C5250 commonsourceibias.n53 gnd 0.00772f
C5251 commonsourceibias.n54 gnd 0.00772f
C5252 commonsourceibias.n55 gnd 0.009185f
C5253 commonsourceibias.n56 gnd 0.010651f
C5254 commonsourceibias.n57 gnd 0.057546f
C5255 commonsourceibias.n58 gnd 0.010587f
C5256 commonsourceibias.n59 gnd 0.00772f
C5257 commonsourceibias.n60 gnd 0.00772f
C5258 commonsourceibias.n61 gnd 0.00772f
C5259 commonsourceibias.n62 gnd 0.010457f
C5260 commonsourceibias.n63 gnd 0.057546f
C5261 commonsourceibias.n64 gnd 0.010526f
C5262 commonsourceibias.n65 gnd 0.009515f
C5263 commonsourceibias.n66 gnd 0.00772f
C5264 commonsourceibias.n67 gnd 0.00772f
C5265 commonsourceibias.n68 gnd 0.007831f
C5266 commonsourceibias.n69 gnd 0.008096f
C5267 commonsourceibias.n70 gnd 0.068855f
C5268 commonsourceibias.n71 gnd 0.076384f
C5269 commonsourceibias.t33 gnd 0.016658f
C5270 commonsourceibias.t15 gnd 0.016658f
C5271 commonsourceibias.n72 gnd 0.147197f
C5272 commonsourceibias.n73 gnd 0.12719f
C5273 commonsourceibias.t25 gnd 0.016658f
C5274 commonsourceibias.t31 gnd 0.016658f
C5275 commonsourceibias.n74 gnd 0.147197f
C5276 commonsourceibias.n75 gnd 0.067614f
C5277 commonsourceibias.t21 gnd 0.016658f
C5278 commonsourceibias.t37 gnd 0.016658f
C5279 commonsourceibias.n76 gnd 0.147197f
C5280 commonsourceibias.n77 gnd 0.056488f
C5281 commonsourceibias.t41 gnd 0.016658f
C5282 commonsourceibias.t47 gnd 0.016658f
C5283 commonsourceibias.n78 gnd 0.14769f
C5284 commonsourceibias.t35 gnd 0.016658f
C5285 commonsourceibias.t11 gnd 0.016658f
C5286 commonsourceibias.n79 gnd 0.147197f
C5287 commonsourceibias.n80 gnd 0.13716f
C5288 commonsourceibias.t45 gnd 0.016658f
C5289 commonsourceibias.t27 gnd 0.016658f
C5290 commonsourceibias.n81 gnd 0.147197f
C5291 commonsourceibias.n82 gnd 0.056488f
C5292 commonsourceibias.n83 gnd 0.068401f
C5293 commonsourceibias.n84 gnd 0.00772f
C5294 commonsourceibias.t50 gnd 0.144227f
C5295 commonsourceibias.t69 gnd 0.144227f
C5296 commonsourceibias.n85 gnd 0.057546f
C5297 commonsourceibias.n86 gnd 0.00772f
C5298 commonsourceibias.t67 gnd 0.144227f
C5299 commonsourceibias.n87 gnd 0.057546f
C5300 commonsourceibias.n88 gnd 0.00772f
C5301 commonsourceibias.t78 gnd 0.144227f
C5302 commonsourceibias.n89 gnd 0.057546f
C5303 commonsourceibias.n90 gnd 0.038863f
C5304 commonsourceibias.t64 gnd 0.144227f
C5305 commonsourceibias.t62 gnd 0.162743f
C5306 commonsourceibias.n91 gnd 0.066782f
C5307 commonsourceibias.n92 gnd 0.069137f
C5308 commonsourceibias.n93 gnd 0.009515f
C5309 commonsourceibias.n94 gnd 0.010526f
C5310 commonsourceibias.n95 gnd 0.00772f
C5311 commonsourceibias.n96 gnd 0.00772f
C5312 commonsourceibias.n97 gnd 0.010457f
C5313 commonsourceibias.n98 gnd 0.006245f
C5314 commonsourceibias.n99 gnd 0.010587f
C5315 commonsourceibias.n100 gnd 0.00772f
C5316 commonsourceibias.n101 gnd 0.00772f
C5317 commonsourceibias.n102 gnd 0.010651f
C5318 commonsourceibias.n103 gnd 0.009185f
C5319 commonsourceibias.n104 gnd 0.007453f
C5320 commonsourceibias.n105 gnd 0.00772f
C5321 commonsourceibias.n106 gnd 0.00772f
C5322 commonsourceibias.n107 gnd 0.009442f
C5323 commonsourceibias.n108 gnd 0.010598f
C5324 commonsourceibias.n109 gnd 0.057546f
C5325 commonsourceibias.n110 gnd 0.010527f
C5326 commonsourceibias.n111 gnd 0.007683f
C5327 commonsourceibias.n112 gnd 0.055804f
C5328 commonsourceibias.n113 gnd 0.007683f
C5329 commonsourceibias.n114 gnd 0.010527f
C5330 commonsourceibias.n115 gnd 0.057546f
C5331 commonsourceibias.n116 gnd 0.010598f
C5332 commonsourceibias.n117 gnd 0.009442f
C5333 commonsourceibias.n118 gnd 0.00772f
C5334 commonsourceibias.n119 gnd 0.00772f
C5335 commonsourceibias.n120 gnd 0.00772f
C5336 commonsourceibias.n121 gnd 0.009185f
C5337 commonsourceibias.n122 gnd 0.010651f
C5338 commonsourceibias.n123 gnd 0.057546f
C5339 commonsourceibias.n124 gnd 0.010587f
C5340 commonsourceibias.n125 gnd 0.00772f
C5341 commonsourceibias.n126 gnd 0.00772f
C5342 commonsourceibias.n127 gnd 0.00772f
C5343 commonsourceibias.n128 gnd 0.010457f
C5344 commonsourceibias.n129 gnd 0.057546f
C5345 commonsourceibias.n130 gnd 0.010526f
C5346 commonsourceibias.n131 gnd 0.009515f
C5347 commonsourceibias.n132 gnd 0.00772f
C5348 commonsourceibias.n133 gnd 0.00772f
C5349 commonsourceibias.n134 gnd 0.007831f
C5350 commonsourceibias.n135 gnd 0.008096f
C5351 commonsourceibias.n136 gnd 0.068855f
C5352 commonsourceibias.n137 gnd 0.04456f
C5353 commonsourceibias.n138 gnd 0.010301f
C5354 commonsourceibias.t72 gnd 0.144227f
C5355 commonsourceibias.n139 gnd 0.057546f
C5356 commonsourceibias.n140 gnd 0.00772f
C5357 commonsourceibias.t49 gnd 0.144227f
C5358 commonsourceibias.n141 gnd 0.006245f
C5359 commonsourceibias.n142 gnd 0.00772f
C5360 commonsourceibias.t95 gnd 0.144227f
C5361 commonsourceibias.n143 gnd 0.007453f
C5362 commonsourceibias.n144 gnd 0.00772f
C5363 commonsourceibias.t66 gnd 0.144227f
C5364 commonsourceibias.n145 gnd 0.057546f
C5365 commonsourceibias.t77 gnd 0.144227f
C5366 commonsourceibias.n146 gnd 0.006235f
C5367 commonsourceibias.n147 gnd 0.00772f
C5368 commonsourceibias.t91 gnd 0.144227f
C5369 commonsourceibias.t60 gnd 0.144227f
C5370 commonsourceibias.n148 gnd 0.057546f
C5371 commonsourceibias.n149 gnd 0.00772f
C5372 commonsourceibias.t58 gnd 0.144227f
C5373 commonsourceibias.n150 gnd 0.057546f
C5374 commonsourceibias.n151 gnd 0.00772f
C5375 commonsourceibias.t68 gnd 0.144227f
C5376 commonsourceibias.n152 gnd 0.057546f
C5377 commonsourceibias.n153 gnd 0.038863f
C5378 commonsourceibias.t57 gnd 0.144227f
C5379 commonsourceibias.t54 gnd 0.162743f
C5380 commonsourceibias.n154 gnd 0.066782f
C5381 commonsourceibias.n155 gnd 0.069137f
C5382 commonsourceibias.n156 gnd 0.009515f
C5383 commonsourceibias.n157 gnd 0.010526f
C5384 commonsourceibias.n158 gnd 0.00772f
C5385 commonsourceibias.n159 gnd 0.00772f
C5386 commonsourceibias.n160 gnd 0.010457f
C5387 commonsourceibias.n161 gnd 0.006245f
C5388 commonsourceibias.n162 gnd 0.010587f
C5389 commonsourceibias.n163 gnd 0.00772f
C5390 commonsourceibias.n164 gnd 0.00772f
C5391 commonsourceibias.n165 gnd 0.010651f
C5392 commonsourceibias.n166 gnd 0.009185f
C5393 commonsourceibias.n167 gnd 0.007453f
C5394 commonsourceibias.n168 gnd 0.00772f
C5395 commonsourceibias.n169 gnd 0.00772f
C5396 commonsourceibias.n170 gnd 0.009442f
C5397 commonsourceibias.n171 gnd 0.010598f
C5398 commonsourceibias.n172 gnd 0.057546f
C5399 commonsourceibias.n173 gnd 0.010527f
C5400 commonsourceibias.n174 gnd 0.00772f
C5401 commonsourceibias.n175 gnd 0.00772f
C5402 commonsourceibias.n176 gnd 0.00772f
C5403 commonsourceibias.n177 gnd 0.010527f
C5404 commonsourceibias.n178 gnd 0.057546f
C5405 commonsourceibias.n179 gnd 0.010598f
C5406 commonsourceibias.n180 gnd 0.009442f
C5407 commonsourceibias.n181 gnd 0.00772f
C5408 commonsourceibias.n182 gnd 0.00772f
C5409 commonsourceibias.n183 gnd 0.00772f
C5410 commonsourceibias.n184 gnd 0.009185f
C5411 commonsourceibias.n185 gnd 0.010651f
C5412 commonsourceibias.n186 gnd 0.057546f
C5413 commonsourceibias.n187 gnd 0.010587f
C5414 commonsourceibias.n188 gnd 0.00772f
C5415 commonsourceibias.n189 gnd 0.00772f
C5416 commonsourceibias.n190 gnd 0.00772f
C5417 commonsourceibias.n191 gnd 0.010457f
C5418 commonsourceibias.n192 gnd 0.057546f
C5419 commonsourceibias.n193 gnd 0.010526f
C5420 commonsourceibias.n194 gnd 0.009515f
C5421 commonsourceibias.n195 gnd 0.00772f
C5422 commonsourceibias.n196 gnd 0.00772f
C5423 commonsourceibias.n197 gnd 0.007831f
C5424 commonsourceibias.n198 gnd 0.008096f
C5425 commonsourceibias.t61 gnd 0.155981f
C5426 commonsourceibias.n199 gnd 0.068855f
C5427 commonsourceibias.n200 gnd 0.023432f
C5428 commonsourceibias.n201 gnd 0.388694f
C5429 commonsourceibias.n202 gnd 0.010301f
C5430 commonsourceibias.t84 gnd 0.155981f
C5431 commonsourceibias.t92 gnd 0.144227f
C5432 commonsourceibias.n203 gnd 0.057546f
C5433 commonsourceibias.n204 gnd 0.00772f
C5434 commonsourceibias.t51 gnd 0.144227f
C5435 commonsourceibias.n205 gnd 0.006245f
C5436 commonsourceibias.n206 gnd 0.00772f
C5437 commonsourceibias.t63 gnd 0.144227f
C5438 commonsourceibias.n207 gnd 0.007453f
C5439 commonsourceibias.n208 gnd 0.00772f
C5440 commonsourceibias.t48 gnd 0.144227f
C5441 commonsourceibias.n209 gnd 0.006235f
C5442 commonsourceibias.n210 gnd 0.00772f
C5443 commonsourceibias.t94 gnd 0.144227f
C5444 commonsourceibias.t83 gnd 0.144227f
C5445 commonsourceibias.n211 gnd 0.057546f
C5446 commonsourceibias.n212 gnd 0.00772f
C5447 commonsourceibias.t80 gnd 0.144227f
C5448 commonsourceibias.n213 gnd 0.057546f
C5449 commonsourceibias.n214 gnd 0.00772f
C5450 commonsourceibias.t90 gnd 0.144227f
C5451 commonsourceibias.n215 gnd 0.057546f
C5452 commonsourceibias.n216 gnd 0.038863f
C5453 commonsourceibias.t59 gnd 0.144227f
C5454 commonsourceibias.t75 gnd 0.162743f
C5455 commonsourceibias.n217 gnd 0.066782f
C5456 commonsourceibias.n218 gnd 0.069137f
C5457 commonsourceibias.n219 gnd 0.009515f
C5458 commonsourceibias.n220 gnd 0.010526f
C5459 commonsourceibias.n221 gnd 0.00772f
C5460 commonsourceibias.n222 gnd 0.00772f
C5461 commonsourceibias.n223 gnd 0.010457f
C5462 commonsourceibias.n224 gnd 0.006245f
C5463 commonsourceibias.n225 gnd 0.010587f
C5464 commonsourceibias.n226 gnd 0.00772f
C5465 commonsourceibias.n227 gnd 0.00772f
C5466 commonsourceibias.n228 gnd 0.010651f
C5467 commonsourceibias.n229 gnd 0.009185f
C5468 commonsourceibias.n230 gnd 0.007453f
C5469 commonsourceibias.n231 gnd 0.00772f
C5470 commonsourceibias.n232 gnd 0.00772f
C5471 commonsourceibias.n233 gnd 0.009442f
C5472 commonsourceibias.n234 gnd 0.010598f
C5473 commonsourceibias.n235 gnd 0.057546f
C5474 commonsourceibias.n236 gnd 0.010527f
C5475 commonsourceibias.n237 gnd 0.007683f
C5476 commonsourceibias.t17 gnd 0.016658f
C5477 commonsourceibias.t9 gnd 0.016658f
C5478 commonsourceibias.n238 gnd 0.14769f
C5479 commonsourceibias.t19 gnd 0.016658f
C5480 commonsourceibias.t5 gnd 0.016658f
C5481 commonsourceibias.n239 gnd 0.147197f
C5482 commonsourceibias.n240 gnd 0.13716f
C5483 commonsourceibias.t43 gnd 0.016658f
C5484 commonsourceibias.t13 gnd 0.016658f
C5485 commonsourceibias.n241 gnd 0.147197f
C5486 commonsourceibias.n242 gnd 0.056488f
C5487 commonsourceibias.n243 gnd 0.010301f
C5488 commonsourceibias.t22 gnd 0.144227f
C5489 commonsourceibias.n244 gnd 0.057546f
C5490 commonsourceibias.n245 gnd 0.00772f
C5491 commonsourceibias.t38 gnd 0.144227f
C5492 commonsourceibias.n246 gnd 0.006245f
C5493 commonsourceibias.n247 gnd 0.00772f
C5494 commonsourceibias.t0 gnd 0.144227f
C5495 commonsourceibias.n248 gnd 0.007453f
C5496 commonsourceibias.n249 gnd 0.00772f
C5497 commonsourceibias.t6 gnd 0.144227f
C5498 commonsourceibias.n250 gnd 0.006235f
C5499 commonsourceibias.n251 gnd 0.00772f
C5500 commonsourceibias.t12 gnd 0.144227f
C5501 commonsourceibias.t42 gnd 0.144227f
C5502 commonsourceibias.n252 gnd 0.057546f
C5503 commonsourceibias.n253 gnd 0.00772f
C5504 commonsourceibias.t4 gnd 0.144227f
C5505 commonsourceibias.n254 gnd 0.057546f
C5506 commonsourceibias.n255 gnd 0.00772f
C5507 commonsourceibias.t18 gnd 0.144227f
C5508 commonsourceibias.n256 gnd 0.057546f
C5509 commonsourceibias.n257 gnd 0.038863f
C5510 commonsourceibias.t8 gnd 0.144227f
C5511 commonsourceibias.t16 gnd 0.162743f
C5512 commonsourceibias.n258 gnd 0.066782f
C5513 commonsourceibias.n259 gnd 0.069137f
C5514 commonsourceibias.n260 gnd 0.009515f
C5515 commonsourceibias.n261 gnd 0.010526f
C5516 commonsourceibias.n262 gnd 0.00772f
C5517 commonsourceibias.n263 gnd 0.00772f
C5518 commonsourceibias.n264 gnd 0.010457f
C5519 commonsourceibias.n265 gnd 0.006245f
C5520 commonsourceibias.n266 gnd 0.010587f
C5521 commonsourceibias.n267 gnd 0.00772f
C5522 commonsourceibias.n268 gnd 0.00772f
C5523 commonsourceibias.n269 gnd 0.010651f
C5524 commonsourceibias.n270 gnd 0.009185f
C5525 commonsourceibias.n271 gnd 0.007453f
C5526 commonsourceibias.n272 gnd 0.00772f
C5527 commonsourceibias.n273 gnd 0.00772f
C5528 commonsourceibias.n274 gnd 0.009442f
C5529 commonsourceibias.n275 gnd 0.010598f
C5530 commonsourceibias.n276 gnd 0.057546f
C5531 commonsourceibias.n277 gnd 0.010527f
C5532 commonsourceibias.n278 gnd 0.00772f
C5533 commonsourceibias.n279 gnd 0.00772f
C5534 commonsourceibias.n280 gnd 0.00772f
C5535 commonsourceibias.n281 gnd 0.010527f
C5536 commonsourceibias.n282 gnd 0.057546f
C5537 commonsourceibias.n283 gnd 0.010598f
C5538 commonsourceibias.t28 gnd 0.144227f
C5539 commonsourceibias.n284 gnd 0.057546f
C5540 commonsourceibias.n285 gnd 0.009442f
C5541 commonsourceibias.n286 gnd 0.00772f
C5542 commonsourceibias.n287 gnd 0.00772f
C5543 commonsourceibias.n288 gnd 0.00772f
C5544 commonsourceibias.n289 gnd 0.009185f
C5545 commonsourceibias.n290 gnd 0.010651f
C5546 commonsourceibias.n291 gnd 0.057546f
C5547 commonsourceibias.n292 gnd 0.010587f
C5548 commonsourceibias.n293 gnd 0.00772f
C5549 commonsourceibias.n294 gnd 0.00772f
C5550 commonsourceibias.n295 gnd 0.00772f
C5551 commonsourceibias.n296 gnd 0.010457f
C5552 commonsourceibias.n297 gnd 0.057546f
C5553 commonsourceibias.n298 gnd 0.010526f
C5554 commonsourceibias.n299 gnd 0.009515f
C5555 commonsourceibias.n300 gnd 0.00772f
C5556 commonsourceibias.n301 gnd 0.00772f
C5557 commonsourceibias.n302 gnd 0.007831f
C5558 commonsourceibias.n303 gnd 0.008096f
C5559 commonsourceibias.t2 gnd 0.155981f
C5560 commonsourceibias.n304 gnd 0.068855f
C5561 commonsourceibias.n305 gnd 0.076384f
C5562 commonsourceibias.t23 gnd 0.016658f
C5563 commonsourceibias.t3 gnd 0.016658f
C5564 commonsourceibias.n306 gnd 0.147197f
C5565 commonsourceibias.n307 gnd 0.12719f
C5566 commonsourceibias.t1 gnd 0.016658f
C5567 commonsourceibias.t39 gnd 0.016658f
C5568 commonsourceibias.n308 gnd 0.147197f
C5569 commonsourceibias.n309 gnd 0.067614f
C5570 commonsourceibias.t7 gnd 0.016658f
C5571 commonsourceibias.t29 gnd 0.016658f
C5572 commonsourceibias.n310 gnd 0.147197f
C5573 commonsourceibias.n311 gnd 0.056488f
C5574 commonsourceibias.n312 gnd 0.068401f
C5575 commonsourceibias.n313 gnd 0.055804f
C5576 commonsourceibias.n314 gnd 0.007683f
C5577 commonsourceibias.n315 gnd 0.010527f
C5578 commonsourceibias.n316 gnd 0.057546f
C5579 commonsourceibias.n317 gnd 0.010598f
C5580 commonsourceibias.t88 gnd 0.144227f
C5581 commonsourceibias.n318 gnd 0.057546f
C5582 commonsourceibias.n319 gnd 0.009442f
C5583 commonsourceibias.n320 gnd 0.00772f
C5584 commonsourceibias.n321 gnd 0.00772f
C5585 commonsourceibias.n322 gnd 0.00772f
C5586 commonsourceibias.n323 gnd 0.009185f
C5587 commonsourceibias.n324 gnd 0.010651f
C5588 commonsourceibias.n325 gnd 0.057546f
C5589 commonsourceibias.n326 gnd 0.010587f
C5590 commonsourceibias.n327 gnd 0.00772f
C5591 commonsourceibias.n328 gnd 0.00772f
C5592 commonsourceibias.n329 gnd 0.00772f
C5593 commonsourceibias.n330 gnd 0.010457f
C5594 commonsourceibias.n331 gnd 0.057546f
C5595 commonsourceibias.n332 gnd 0.010526f
C5596 commonsourceibias.n333 gnd 0.009515f
C5597 commonsourceibias.n334 gnd 0.00772f
C5598 commonsourceibias.n335 gnd 0.00772f
C5599 commonsourceibias.n336 gnd 0.007831f
C5600 commonsourceibias.n337 gnd 0.008096f
C5601 commonsourceibias.n338 gnd 0.068855f
C5602 commonsourceibias.n339 gnd 0.04456f
C5603 commonsourceibias.n340 gnd 0.010301f
C5604 commonsourceibias.t85 gnd 0.144227f
C5605 commonsourceibias.n341 gnd 0.057546f
C5606 commonsourceibias.n342 gnd 0.00772f
C5607 commonsourceibias.t93 gnd 0.144227f
C5608 commonsourceibias.n343 gnd 0.006245f
C5609 commonsourceibias.n344 gnd 0.00772f
C5610 commonsourceibias.t56 gnd 0.144227f
C5611 commonsourceibias.n345 gnd 0.007453f
C5612 commonsourceibias.n346 gnd 0.00772f
C5613 commonsourceibias.t89 gnd 0.144227f
C5614 commonsourceibias.n347 gnd 0.006235f
C5615 commonsourceibias.n348 gnd 0.00772f
C5616 commonsourceibias.t87 gnd 0.144227f
C5617 commonsourceibias.t74 gnd 0.144227f
C5618 commonsourceibias.n349 gnd 0.057546f
C5619 commonsourceibias.n350 gnd 0.00772f
C5620 commonsourceibias.t70 gnd 0.144227f
C5621 commonsourceibias.n351 gnd 0.057546f
C5622 commonsourceibias.n352 gnd 0.00772f
C5623 commonsourceibias.t82 gnd 0.144227f
C5624 commonsourceibias.n353 gnd 0.057546f
C5625 commonsourceibias.n354 gnd 0.038863f
C5626 commonsourceibias.t52 gnd 0.144227f
C5627 commonsourceibias.t65 gnd 0.162743f
C5628 commonsourceibias.n355 gnd 0.066782f
C5629 commonsourceibias.n356 gnd 0.069137f
C5630 commonsourceibias.n357 gnd 0.009515f
C5631 commonsourceibias.n358 gnd 0.010526f
C5632 commonsourceibias.n359 gnd 0.00772f
C5633 commonsourceibias.n360 gnd 0.00772f
C5634 commonsourceibias.n361 gnd 0.010457f
C5635 commonsourceibias.n362 gnd 0.006245f
C5636 commonsourceibias.n363 gnd 0.010587f
C5637 commonsourceibias.n364 gnd 0.00772f
C5638 commonsourceibias.n365 gnd 0.00772f
C5639 commonsourceibias.n366 gnd 0.010651f
C5640 commonsourceibias.n367 gnd 0.009185f
C5641 commonsourceibias.n368 gnd 0.007453f
C5642 commonsourceibias.n369 gnd 0.00772f
C5643 commonsourceibias.n370 gnd 0.00772f
C5644 commonsourceibias.n371 gnd 0.009442f
C5645 commonsourceibias.n372 gnd 0.010598f
C5646 commonsourceibias.n373 gnd 0.057546f
C5647 commonsourceibias.n374 gnd 0.010527f
C5648 commonsourceibias.n375 gnd 0.00772f
C5649 commonsourceibias.n376 gnd 0.00772f
C5650 commonsourceibias.n377 gnd 0.00772f
C5651 commonsourceibias.n378 gnd 0.010527f
C5652 commonsourceibias.n379 gnd 0.057546f
C5653 commonsourceibias.n380 gnd 0.010598f
C5654 commonsourceibias.t79 gnd 0.144227f
C5655 commonsourceibias.n381 gnd 0.057546f
C5656 commonsourceibias.n382 gnd 0.009442f
C5657 commonsourceibias.n383 gnd 0.00772f
C5658 commonsourceibias.n384 gnd 0.00772f
C5659 commonsourceibias.n385 gnd 0.00772f
C5660 commonsourceibias.n386 gnd 0.009185f
C5661 commonsourceibias.n387 gnd 0.010651f
C5662 commonsourceibias.n388 gnd 0.057546f
C5663 commonsourceibias.n389 gnd 0.010587f
C5664 commonsourceibias.n390 gnd 0.00772f
C5665 commonsourceibias.n391 gnd 0.00772f
C5666 commonsourceibias.n392 gnd 0.00772f
C5667 commonsourceibias.n393 gnd 0.010457f
C5668 commonsourceibias.n394 gnd 0.057546f
C5669 commonsourceibias.n395 gnd 0.010526f
C5670 commonsourceibias.n396 gnd 0.009515f
C5671 commonsourceibias.n397 gnd 0.00772f
C5672 commonsourceibias.n398 gnd 0.00772f
C5673 commonsourceibias.n399 gnd 0.007831f
C5674 commonsourceibias.n400 gnd 0.008096f
C5675 commonsourceibias.t73 gnd 0.155981f
C5676 commonsourceibias.n401 gnd 0.068855f
C5677 commonsourceibias.n402 gnd 0.023432f
C5678 commonsourceibias.n403 gnd 0.212991f
C5679 commonsourceibias.n404 gnd 4.01312f
.ends

