* NGSPICE file created from diffpair.ext - technology: sky130A

.subckt diffpair minus drain_right drain_left source plus
X0 source.t15 plus.t0 drain_left.t7 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X1 a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=18.72 ps=102.24 w=6 l=1
X2 drain_left.t2 plus.t1 source.t14 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X3 drain_left.t0 plus.t2 source.t13 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X4 a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X5 source.t12 plus.t3 drain_left.t6 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X6 source.t11 plus.t4 drain_left.t1 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X7 drain_right.t7 minus.t0 source.t3 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X8 drain_left.t4 plus.t5 source.t10 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X9 drain_right.t6 minus.t1 source.t0 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X10 source.t4 minus.t2 drain_right.t5 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X11 a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X12 drain_right.t4 minus.t3 source.t6 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X13 drain_right.t3 minus.t4 source.t1 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=2.34 ps=12.78 w=6 l=1
X14 drain_left.t3 plus.t6 source.t9 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X15 a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=1
X16 source.t2 minus.t5 drain_right.t2 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X17 source.t7 minus.t6 drain_right.t1 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=0.99 pd=6.33 as=0.99 ps=6.33 w=6 l=1
X18 source.t5 minus.t7 drain_right.t0 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
X19 source.t8 plus.t7 drain_left.t5 a_n2046_n2088# sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0.99 ps=6.33 w=6 l=1
R0 plus.n2 plus.t7 199.144
R1 plus.n15 plus.t5 199.144
R2 plus.n11 plus.t2 183.883
R3 plus.n24 plus.t3 183.883
R4 plus.n5 plus.n4 161.3
R5 plus.n6 plus.n1 161.3
R6 plus.n8 plus.n7 161.3
R7 plus.n10 plus.n0 161.3
R8 plus.n18 plus.n17 161.3
R9 plus.n19 plus.n14 161.3
R10 plus.n21 plus.n20 161.3
R11 plus.n23 plus.n13 161.3
R12 plus.n9 plus.t0 144.601
R13 plus.n3 plus.t1 144.601
R14 plus.n22 plus.t6 144.601
R15 plus.n16 plus.t4 144.601
R16 plus.n12 plus.n11 80.6037
R17 plus.n25 plus.n24 80.6037
R18 plus.n11 plus.n10 56.3158
R19 plus.n24 plus.n23 56.3158
R20 plus.n3 plus.n2 46.9082
R21 plus.n16 plus.n15 46.9082
R22 plus.n5 plus.n2 43.8991
R23 plus.n18 plus.n15 43.8991
R24 plus.n8 plus.n1 40.577
R25 plus.n4 plus.n1 40.577
R26 plus.n21 plus.n14 40.577
R27 plus.n17 plus.n14 40.577
R28 plus plus.n25 28.8593
R29 plus.n10 plus.n9 16.477
R30 plus.n23 plus.n22 16.477
R31 plus plus.n12 10.2509
R32 plus.n9 plus.n8 8.11581
R33 plus.n4 plus.n3 8.11581
R34 plus.n22 plus.n21 8.11581
R35 plus.n17 plus.n16 8.11581
R36 plus.n12 plus.n0 0.285035
R37 plus.n25 plus.n13 0.285035
R38 plus.n6 plus.n5 0.189894
R39 plus.n7 plus.n6 0.189894
R40 plus.n7 plus.n0 0.189894
R41 plus.n20 plus.n13 0.189894
R42 plus.n20 plus.n19 0.189894
R43 plus.n19 plus.n18 0.189894
R44 drain_left.n5 drain_left.n3 68.3374
R45 drain_left.n2 drain_left.n1 67.7086
R46 drain_left.n2 drain_left.n0 67.7086
R47 drain_left.n5 drain_left.n4 67.1907
R48 drain_left drain_left.n2 26.8346
R49 drain_left drain_left.n5 6.79977
R50 drain_left.n1 drain_left.t1 3.3005
R51 drain_left.n1 drain_left.t4 3.3005
R52 drain_left.n0 drain_left.t6 3.3005
R53 drain_left.n0 drain_left.t3 3.3005
R54 drain_left.n4 drain_left.t7 3.3005
R55 drain_left.n4 drain_left.t0 3.3005
R56 drain_left.n3 drain_left.t5 3.3005
R57 drain_left.n3 drain_left.t2 3.3005
R58 source.n258 source.n232 289.615
R59 source.n224 source.n198 289.615
R60 source.n192 source.n166 289.615
R61 source.n158 source.n132 289.615
R62 source.n26 source.n0 289.615
R63 source.n60 source.n34 289.615
R64 source.n92 source.n66 289.615
R65 source.n126 source.n100 289.615
R66 source.n243 source.n242 185
R67 source.n240 source.n239 185
R68 source.n249 source.n248 185
R69 source.n251 source.n250 185
R70 source.n236 source.n235 185
R71 source.n257 source.n256 185
R72 source.n259 source.n258 185
R73 source.n209 source.n208 185
R74 source.n206 source.n205 185
R75 source.n215 source.n214 185
R76 source.n217 source.n216 185
R77 source.n202 source.n201 185
R78 source.n223 source.n222 185
R79 source.n225 source.n224 185
R80 source.n177 source.n176 185
R81 source.n174 source.n173 185
R82 source.n183 source.n182 185
R83 source.n185 source.n184 185
R84 source.n170 source.n169 185
R85 source.n191 source.n190 185
R86 source.n193 source.n192 185
R87 source.n143 source.n142 185
R88 source.n140 source.n139 185
R89 source.n149 source.n148 185
R90 source.n151 source.n150 185
R91 source.n136 source.n135 185
R92 source.n157 source.n156 185
R93 source.n159 source.n158 185
R94 source.n27 source.n26 185
R95 source.n25 source.n24 185
R96 source.n4 source.n3 185
R97 source.n19 source.n18 185
R98 source.n17 source.n16 185
R99 source.n8 source.n7 185
R100 source.n11 source.n10 185
R101 source.n61 source.n60 185
R102 source.n59 source.n58 185
R103 source.n38 source.n37 185
R104 source.n53 source.n52 185
R105 source.n51 source.n50 185
R106 source.n42 source.n41 185
R107 source.n45 source.n44 185
R108 source.n93 source.n92 185
R109 source.n91 source.n90 185
R110 source.n70 source.n69 185
R111 source.n85 source.n84 185
R112 source.n83 source.n82 185
R113 source.n74 source.n73 185
R114 source.n77 source.n76 185
R115 source.n127 source.n126 185
R116 source.n125 source.n124 185
R117 source.n104 source.n103 185
R118 source.n119 source.n118 185
R119 source.n117 source.n116 185
R120 source.n108 source.n107 185
R121 source.n111 source.n110 185
R122 source.t1 source.n241 147.661
R123 source.t4 source.n207 147.661
R124 source.t10 source.n175 147.661
R125 source.t12 source.n141 147.661
R126 source.t13 source.n9 147.661
R127 source.t8 source.n43 147.661
R128 source.t0 source.n75 147.661
R129 source.t5 source.n109 147.661
R130 source.n242 source.n239 104.615
R131 source.n249 source.n239 104.615
R132 source.n250 source.n249 104.615
R133 source.n250 source.n235 104.615
R134 source.n257 source.n235 104.615
R135 source.n258 source.n257 104.615
R136 source.n208 source.n205 104.615
R137 source.n215 source.n205 104.615
R138 source.n216 source.n215 104.615
R139 source.n216 source.n201 104.615
R140 source.n223 source.n201 104.615
R141 source.n224 source.n223 104.615
R142 source.n176 source.n173 104.615
R143 source.n183 source.n173 104.615
R144 source.n184 source.n183 104.615
R145 source.n184 source.n169 104.615
R146 source.n191 source.n169 104.615
R147 source.n192 source.n191 104.615
R148 source.n142 source.n139 104.615
R149 source.n149 source.n139 104.615
R150 source.n150 source.n149 104.615
R151 source.n150 source.n135 104.615
R152 source.n157 source.n135 104.615
R153 source.n158 source.n157 104.615
R154 source.n26 source.n25 104.615
R155 source.n25 source.n3 104.615
R156 source.n18 source.n3 104.615
R157 source.n18 source.n17 104.615
R158 source.n17 source.n7 104.615
R159 source.n10 source.n7 104.615
R160 source.n60 source.n59 104.615
R161 source.n59 source.n37 104.615
R162 source.n52 source.n37 104.615
R163 source.n52 source.n51 104.615
R164 source.n51 source.n41 104.615
R165 source.n44 source.n41 104.615
R166 source.n92 source.n91 104.615
R167 source.n91 source.n69 104.615
R168 source.n84 source.n69 104.615
R169 source.n84 source.n83 104.615
R170 source.n83 source.n73 104.615
R171 source.n76 source.n73 104.615
R172 source.n126 source.n125 104.615
R173 source.n125 source.n103 104.615
R174 source.n118 source.n103 104.615
R175 source.n118 source.n117 104.615
R176 source.n117 source.n107 104.615
R177 source.n110 source.n107 104.615
R178 source.n242 source.t1 52.3082
R179 source.n208 source.t4 52.3082
R180 source.n176 source.t10 52.3082
R181 source.n142 source.t12 52.3082
R182 source.n10 source.t13 52.3082
R183 source.n44 source.t8 52.3082
R184 source.n76 source.t0 52.3082
R185 source.n110 source.t5 52.3082
R186 source.n33 source.n32 50.512
R187 source.n99 source.n98 50.512
R188 source.n231 source.n230 50.5119
R189 source.n165 source.n164 50.5119
R190 source.n263 source.n262 32.1853
R191 source.n229 source.n228 32.1853
R192 source.n197 source.n196 32.1853
R193 source.n163 source.n162 32.1853
R194 source.n31 source.n30 32.1853
R195 source.n65 source.n64 32.1853
R196 source.n97 source.n96 32.1853
R197 source.n131 source.n130 32.1853
R198 source.n163 source.n131 17.8888
R199 source.n243 source.n241 15.6674
R200 source.n209 source.n207 15.6674
R201 source.n177 source.n175 15.6674
R202 source.n143 source.n141 15.6674
R203 source.n11 source.n9 15.6674
R204 source.n45 source.n43 15.6674
R205 source.n77 source.n75 15.6674
R206 source.n111 source.n109 15.6674
R207 source.n244 source.n240 12.8005
R208 source.n210 source.n206 12.8005
R209 source.n178 source.n174 12.8005
R210 source.n144 source.n140 12.8005
R211 source.n12 source.n8 12.8005
R212 source.n46 source.n42 12.8005
R213 source.n78 source.n74 12.8005
R214 source.n112 source.n108 12.8005
R215 source.n264 source.n31 12.0526
R216 source.n248 source.n247 12.0247
R217 source.n214 source.n213 12.0247
R218 source.n182 source.n181 12.0247
R219 source.n148 source.n147 12.0247
R220 source.n16 source.n15 12.0247
R221 source.n50 source.n49 12.0247
R222 source.n82 source.n81 12.0247
R223 source.n116 source.n115 12.0247
R224 source.n251 source.n238 11.249
R225 source.n217 source.n204 11.249
R226 source.n185 source.n172 11.249
R227 source.n151 source.n138 11.249
R228 source.n19 source.n6 11.249
R229 source.n53 source.n40 11.249
R230 source.n85 source.n72 11.249
R231 source.n119 source.n106 11.249
R232 source.n252 source.n236 10.4732
R233 source.n218 source.n202 10.4732
R234 source.n186 source.n170 10.4732
R235 source.n152 source.n136 10.4732
R236 source.n20 source.n4 10.4732
R237 source.n54 source.n38 10.4732
R238 source.n86 source.n70 10.4732
R239 source.n120 source.n104 10.4732
R240 source.n256 source.n255 9.69747
R241 source.n222 source.n221 9.69747
R242 source.n190 source.n189 9.69747
R243 source.n156 source.n155 9.69747
R244 source.n24 source.n23 9.69747
R245 source.n58 source.n57 9.69747
R246 source.n90 source.n89 9.69747
R247 source.n124 source.n123 9.69747
R248 source.n262 source.n261 9.45567
R249 source.n228 source.n227 9.45567
R250 source.n196 source.n195 9.45567
R251 source.n162 source.n161 9.45567
R252 source.n30 source.n29 9.45567
R253 source.n64 source.n63 9.45567
R254 source.n96 source.n95 9.45567
R255 source.n130 source.n129 9.45567
R256 source.n261 source.n260 9.3005
R257 source.n234 source.n233 9.3005
R258 source.n255 source.n254 9.3005
R259 source.n253 source.n252 9.3005
R260 source.n238 source.n237 9.3005
R261 source.n247 source.n246 9.3005
R262 source.n245 source.n244 9.3005
R263 source.n227 source.n226 9.3005
R264 source.n200 source.n199 9.3005
R265 source.n221 source.n220 9.3005
R266 source.n219 source.n218 9.3005
R267 source.n204 source.n203 9.3005
R268 source.n213 source.n212 9.3005
R269 source.n211 source.n210 9.3005
R270 source.n195 source.n194 9.3005
R271 source.n168 source.n167 9.3005
R272 source.n189 source.n188 9.3005
R273 source.n187 source.n186 9.3005
R274 source.n172 source.n171 9.3005
R275 source.n181 source.n180 9.3005
R276 source.n179 source.n178 9.3005
R277 source.n161 source.n160 9.3005
R278 source.n134 source.n133 9.3005
R279 source.n155 source.n154 9.3005
R280 source.n153 source.n152 9.3005
R281 source.n138 source.n137 9.3005
R282 source.n147 source.n146 9.3005
R283 source.n145 source.n144 9.3005
R284 source.n29 source.n28 9.3005
R285 source.n2 source.n1 9.3005
R286 source.n23 source.n22 9.3005
R287 source.n21 source.n20 9.3005
R288 source.n6 source.n5 9.3005
R289 source.n15 source.n14 9.3005
R290 source.n13 source.n12 9.3005
R291 source.n63 source.n62 9.3005
R292 source.n36 source.n35 9.3005
R293 source.n57 source.n56 9.3005
R294 source.n55 source.n54 9.3005
R295 source.n40 source.n39 9.3005
R296 source.n49 source.n48 9.3005
R297 source.n47 source.n46 9.3005
R298 source.n95 source.n94 9.3005
R299 source.n68 source.n67 9.3005
R300 source.n89 source.n88 9.3005
R301 source.n87 source.n86 9.3005
R302 source.n72 source.n71 9.3005
R303 source.n81 source.n80 9.3005
R304 source.n79 source.n78 9.3005
R305 source.n129 source.n128 9.3005
R306 source.n102 source.n101 9.3005
R307 source.n123 source.n122 9.3005
R308 source.n121 source.n120 9.3005
R309 source.n106 source.n105 9.3005
R310 source.n115 source.n114 9.3005
R311 source.n113 source.n112 9.3005
R312 source.n259 source.n234 8.92171
R313 source.n225 source.n200 8.92171
R314 source.n193 source.n168 8.92171
R315 source.n159 source.n134 8.92171
R316 source.n27 source.n2 8.92171
R317 source.n61 source.n36 8.92171
R318 source.n93 source.n68 8.92171
R319 source.n127 source.n102 8.92171
R320 source.n260 source.n232 8.14595
R321 source.n226 source.n198 8.14595
R322 source.n194 source.n166 8.14595
R323 source.n160 source.n132 8.14595
R324 source.n28 source.n0 8.14595
R325 source.n62 source.n34 8.14595
R326 source.n94 source.n66 8.14595
R327 source.n128 source.n100 8.14595
R328 source.n264 source.n263 5.83671
R329 source.n262 source.n232 5.81868
R330 source.n228 source.n198 5.81868
R331 source.n196 source.n166 5.81868
R332 source.n162 source.n132 5.81868
R333 source.n30 source.n0 5.81868
R334 source.n64 source.n34 5.81868
R335 source.n96 source.n66 5.81868
R336 source.n130 source.n100 5.81868
R337 source.n260 source.n259 5.04292
R338 source.n226 source.n225 5.04292
R339 source.n194 source.n193 5.04292
R340 source.n160 source.n159 5.04292
R341 source.n28 source.n27 5.04292
R342 source.n62 source.n61 5.04292
R343 source.n94 source.n93 5.04292
R344 source.n128 source.n127 5.04292
R345 source.n245 source.n241 4.38594
R346 source.n211 source.n207 4.38594
R347 source.n179 source.n175 4.38594
R348 source.n145 source.n141 4.38594
R349 source.n13 source.n9 4.38594
R350 source.n47 source.n43 4.38594
R351 source.n79 source.n75 4.38594
R352 source.n113 source.n109 4.38594
R353 source.n256 source.n234 4.26717
R354 source.n222 source.n200 4.26717
R355 source.n190 source.n168 4.26717
R356 source.n156 source.n134 4.26717
R357 source.n24 source.n2 4.26717
R358 source.n58 source.n36 4.26717
R359 source.n90 source.n68 4.26717
R360 source.n124 source.n102 4.26717
R361 source.n255 source.n236 3.49141
R362 source.n221 source.n202 3.49141
R363 source.n189 source.n170 3.49141
R364 source.n155 source.n136 3.49141
R365 source.n23 source.n4 3.49141
R366 source.n57 source.n38 3.49141
R367 source.n89 source.n70 3.49141
R368 source.n123 source.n104 3.49141
R369 source.n230 source.t3 3.3005
R370 source.n230 source.t7 3.3005
R371 source.n164 source.t9 3.3005
R372 source.n164 source.t11 3.3005
R373 source.n32 source.t14 3.3005
R374 source.n32 source.t15 3.3005
R375 source.n98 source.t6 3.3005
R376 source.n98 source.t2 3.3005
R377 source.n252 source.n251 2.71565
R378 source.n218 source.n217 2.71565
R379 source.n186 source.n185 2.71565
R380 source.n152 source.n151 2.71565
R381 source.n20 source.n19 2.71565
R382 source.n54 source.n53 2.71565
R383 source.n86 source.n85 2.71565
R384 source.n120 source.n119 2.71565
R385 source.n248 source.n238 1.93989
R386 source.n214 source.n204 1.93989
R387 source.n182 source.n172 1.93989
R388 source.n148 source.n138 1.93989
R389 source.n16 source.n6 1.93989
R390 source.n50 source.n40 1.93989
R391 source.n82 source.n72 1.93989
R392 source.n116 source.n106 1.93989
R393 source.n247 source.n240 1.16414
R394 source.n213 source.n206 1.16414
R395 source.n181 source.n174 1.16414
R396 source.n147 source.n140 1.16414
R397 source.n15 source.n8 1.16414
R398 source.n49 source.n42 1.16414
R399 source.n81 source.n74 1.16414
R400 source.n115 source.n108 1.16414
R401 source.n131 source.n99 1.14705
R402 source.n99 source.n97 1.14705
R403 source.n65 source.n33 1.14705
R404 source.n33 source.n31 1.14705
R405 source.n165 source.n163 1.14705
R406 source.n197 source.n165 1.14705
R407 source.n231 source.n229 1.14705
R408 source.n263 source.n231 1.14705
R409 source.n97 source.n65 0.470328
R410 source.n229 source.n197 0.470328
R411 source.n244 source.n243 0.388379
R412 source.n210 source.n209 0.388379
R413 source.n178 source.n177 0.388379
R414 source.n144 source.n143 0.388379
R415 source.n12 source.n11 0.388379
R416 source.n46 source.n45 0.388379
R417 source.n78 source.n77 0.388379
R418 source.n112 source.n111 0.388379
R419 source source.n264 0.188
R420 source.n246 source.n245 0.155672
R421 source.n246 source.n237 0.155672
R422 source.n253 source.n237 0.155672
R423 source.n254 source.n253 0.155672
R424 source.n254 source.n233 0.155672
R425 source.n261 source.n233 0.155672
R426 source.n212 source.n211 0.155672
R427 source.n212 source.n203 0.155672
R428 source.n219 source.n203 0.155672
R429 source.n220 source.n219 0.155672
R430 source.n220 source.n199 0.155672
R431 source.n227 source.n199 0.155672
R432 source.n180 source.n179 0.155672
R433 source.n180 source.n171 0.155672
R434 source.n187 source.n171 0.155672
R435 source.n188 source.n187 0.155672
R436 source.n188 source.n167 0.155672
R437 source.n195 source.n167 0.155672
R438 source.n146 source.n145 0.155672
R439 source.n146 source.n137 0.155672
R440 source.n153 source.n137 0.155672
R441 source.n154 source.n153 0.155672
R442 source.n154 source.n133 0.155672
R443 source.n161 source.n133 0.155672
R444 source.n29 source.n1 0.155672
R445 source.n22 source.n1 0.155672
R446 source.n22 source.n21 0.155672
R447 source.n21 source.n5 0.155672
R448 source.n14 source.n5 0.155672
R449 source.n14 source.n13 0.155672
R450 source.n63 source.n35 0.155672
R451 source.n56 source.n35 0.155672
R452 source.n56 source.n55 0.155672
R453 source.n55 source.n39 0.155672
R454 source.n48 source.n39 0.155672
R455 source.n48 source.n47 0.155672
R456 source.n95 source.n67 0.155672
R457 source.n88 source.n67 0.155672
R458 source.n88 source.n87 0.155672
R459 source.n87 source.n71 0.155672
R460 source.n80 source.n71 0.155672
R461 source.n80 source.n79 0.155672
R462 source.n129 source.n101 0.155672
R463 source.n122 source.n101 0.155672
R464 source.n122 source.n121 0.155672
R465 source.n121 source.n105 0.155672
R466 source.n114 source.n105 0.155672
R467 source.n114 source.n113 0.155672
R468 minus.n2 minus.t1 199.144
R469 minus.n15 minus.t2 199.144
R470 minus.n11 minus.t7 183.883
R471 minus.n24 minus.t4 183.883
R472 minus.n10 minus.n0 161.3
R473 minus.n8 minus.n7 161.3
R474 minus.n6 minus.n1 161.3
R475 minus.n5 minus.n4 161.3
R476 minus.n23 minus.n13 161.3
R477 minus.n21 minus.n20 161.3
R478 minus.n19 minus.n14 161.3
R479 minus.n18 minus.n17 161.3
R480 minus.n3 minus.t5 144.601
R481 minus.n9 minus.t3 144.601
R482 minus.n16 minus.t0 144.601
R483 minus.n22 minus.t6 144.601
R484 minus.n12 minus.n11 80.6037
R485 minus.n25 minus.n24 80.6037
R486 minus.n11 minus.n10 56.3158
R487 minus.n24 minus.n23 56.3158
R488 minus.n3 minus.n2 46.9082
R489 minus.n16 minus.n15 46.9082
R490 minus.n5 minus.n2 43.8991
R491 minus.n18 minus.n15 43.8991
R492 minus.n4 minus.n1 40.577
R493 minus.n8 minus.n1 40.577
R494 minus.n17 minus.n14 40.577
R495 minus.n21 minus.n14 40.577
R496 minus.n26 minus.n12 32.7055
R497 minus.n10 minus.n9 16.477
R498 minus.n23 minus.n22 16.477
R499 minus.n4 minus.n3 8.11581
R500 minus.n9 minus.n8 8.11581
R501 minus.n17 minus.n16 8.11581
R502 minus.n22 minus.n21 8.11581
R503 minus.n26 minus.n25 6.87973
R504 minus.n12 minus.n0 0.285035
R505 minus.n25 minus.n13 0.285035
R506 minus.n7 minus.n0 0.189894
R507 minus.n7 minus.n6 0.189894
R508 minus.n6 minus.n5 0.189894
R509 minus.n19 minus.n18 0.189894
R510 minus.n20 minus.n19 0.189894
R511 minus.n20 minus.n13 0.189894
R512 minus minus.n26 0.188
R513 drain_right.n5 drain_right.n3 68.3372
R514 drain_right.n2 drain_right.n1 67.7086
R515 drain_right.n2 drain_right.n0 67.7086
R516 drain_right.n5 drain_right.n4 67.1908
R517 drain_right drain_right.n2 26.2813
R518 drain_right drain_right.n5 6.79977
R519 drain_right.n1 drain_right.t1 3.3005
R520 drain_right.n1 drain_right.t3 3.3005
R521 drain_right.n0 drain_right.t5 3.3005
R522 drain_right.n0 drain_right.t7 3.3005
R523 drain_right.n3 drain_right.t2 3.3005
R524 drain_right.n3 drain_right.t6 3.3005
R525 drain_right.n4 drain_right.t0 3.3005
R526 drain_right.n4 drain_right.t4 3.3005
C0 drain_right minus 3.46293f
C1 plus minus 4.57166f
C2 drain_left minus 0.172134f
C3 drain_right source 6.0968f
C4 source plus 3.67766f
C5 drain_right plus 0.355422f
C6 drain_left source 6.09324f
C7 drain_right drain_left 0.975109f
C8 source minus 3.66364f
C9 drain_left plus 3.663f
C10 drain_right a_n2046_n2088# 4.76271f
C11 drain_left a_n2046_n2088# 5.05962f
C12 source a_n2046_n2088# 5.589285f
C13 minus a_n2046_n2088# 7.431395f
C14 plus a_n2046_n2088# 8.733979f
C15 drain_right.t5 a_n2046_n2088# 0.120858f
C16 drain_right.t7 a_n2046_n2088# 0.120858f
C17 drain_right.n0 a_n2046_n2088# 1.01067f
C18 drain_right.t1 a_n2046_n2088# 0.120858f
C19 drain_right.t3 a_n2046_n2088# 0.120858f
C20 drain_right.n1 a_n2046_n2088# 1.01067f
C21 drain_right.n2 a_n2046_n2088# 1.66162f
C22 drain_right.t2 a_n2046_n2088# 0.120858f
C23 drain_right.t6 a_n2046_n2088# 0.120858f
C24 drain_right.n3 a_n2046_n2088# 1.01476f
C25 drain_right.t0 a_n2046_n2088# 0.120858f
C26 drain_right.t4 a_n2046_n2088# 0.120858f
C27 drain_right.n4 a_n2046_n2088# 1.00796f
C28 drain_right.n5 a_n2046_n2088# 1.02846f
C29 minus.n0 a_n2046_n2088# 0.053307f
C30 minus.t3 a_n2046_n2088# 0.634422f
C31 minus.n1 a_n2046_n2088# 0.032266f
C32 minus.t1 a_n2046_n2088# 0.719971f
C33 minus.n2 a_n2046_n2088# 0.317661f
C34 minus.t5 a_n2046_n2088# 0.634422f
C35 minus.n3 a_n2046_n2088# 0.296035f
C36 minus.n4 a_n2046_n2088# 0.054477f
C37 minus.n5 a_n2046_n2088# 0.171022f
C38 minus.n6 a_n2046_n2088# 0.039949f
C39 minus.n7 a_n2046_n2088# 0.039949f
C40 minus.n8 a_n2046_n2088# 0.054477f
C41 minus.n9 a_n2046_n2088# 0.260486f
C42 minus.n10 a_n2046_n2088# 0.054796f
C43 minus.t7 a_n2046_n2088# 0.695252f
C44 minus.n11 a_n2046_n2088# 0.322287f
C45 minus.n12 a_n2046_n2088# 1.22771f
C46 minus.n13 a_n2046_n2088# 0.053307f
C47 minus.t6 a_n2046_n2088# 0.634422f
C48 minus.n14 a_n2046_n2088# 0.032266f
C49 minus.t2 a_n2046_n2088# 0.719971f
C50 minus.n15 a_n2046_n2088# 0.317661f
C51 minus.t0 a_n2046_n2088# 0.634422f
C52 minus.n16 a_n2046_n2088# 0.296035f
C53 minus.n17 a_n2046_n2088# 0.054477f
C54 minus.n18 a_n2046_n2088# 0.171022f
C55 minus.n19 a_n2046_n2088# 0.039949f
C56 minus.n20 a_n2046_n2088# 0.039949f
C57 minus.n21 a_n2046_n2088# 0.054477f
C58 minus.n22 a_n2046_n2088# 0.260486f
C59 minus.n23 a_n2046_n2088# 0.054796f
C60 minus.t4 a_n2046_n2088# 0.695252f
C61 minus.n24 a_n2046_n2088# 0.322287f
C62 minus.n25 a_n2046_n2088# 0.31023f
C63 minus.n26 a_n2046_n2088# 1.47427f
C64 source.n0 a_n2046_n2088# 0.030265f
C65 source.n1 a_n2046_n2088# 0.021532f
C66 source.n2 a_n2046_n2088# 0.01157f
C67 source.n3 a_n2046_n2088# 0.027348f
C68 source.n4 a_n2046_n2088# 0.012251f
C69 source.n5 a_n2046_n2088# 0.021532f
C70 source.n6 a_n2046_n2088# 0.01157f
C71 source.n7 a_n2046_n2088# 0.027348f
C72 source.n8 a_n2046_n2088# 0.012251f
C73 source.n9 a_n2046_n2088# 0.09214f
C74 source.t13 a_n2046_n2088# 0.044573f
C75 source.n10 a_n2046_n2088# 0.020511f
C76 source.n11 a_n2046_n2088# 0.016154f
C77 source.n12 a_n2046_n2088# 0.01157f
C78 source.n13 a_n2046_n2088# 0.512324f
C79 source.n14 a_n2046_n2088# 0.021532f
C80 source.n15 a_n2046_n2088# 0.01157f
C81 source.n16 a_n2046_n2088# 0.012251f
C82 source.n17 a_n2046_n2088# 0.027348f
C83 source.n18 a_n2046_n2088# 0.027348f
C84 source.n19 a_n2046_n2088# 0.012251f
C85 source.n20 a_n2046_n2088# 0.01157f
C86 source.n21 a_n2046_n2088# 0.021532f
C87 source.n22 a_n2046_n2088# 0.021532f
C88 source.n23 a_n2046_n2088# 0.01157f
C89 source.n24 a_n2046_n2088# 0.012251f
C90 source.n25 a_n2046_n2088# 0.027348f
C91 source.n26 a_n2046_n2088# 0.059203f
C92 source.n27 a_n2046_n2088# 0.012251f
C93 source.n28 a_n2046_n2088# 0.01157f
C94 source.n29 a_n2046_n2088# 0.049769f
C95 source.n30 a_n2046_n2088# 0.033126f
C96 source.n31 a_n2046_n2088# 0.593096f
C97 source.t14 a_n2046_n2088# 0.10209f
C98 source.t15 a_n2046_n2088# 0.10209f
C99 source.n32 a_n2046_n2088# 0.795082f
C100 source.n33 a_n2046_n2088# 0.360933f
C101 source.n34 a_n2046_n2088# 0.030265f
C102 source.n35 a_n2046_n2088# 0.021532f
C103 source.n36 a_n2046_n2088# 0.01157f
C104 source.n37 a_n2046_n2088# 0.027348f
C105 source.n38 a_n2046_n2088# 0.012251f
C106 source.n39 a_n2046_n2088# 0.021532f
C107 source.n40 a_n2046_n2088# 0.01157f
C108 source.n41 a_n2046_n2088# 0.027348f
C109 source.n42 a_n2046_n2088# 0.012251f
C110 source.n43 a_n2046_n2088# 0.09214f
C111 source.t8 a_n2046_n2088# 0.044573f
C112 source.n44 a_n2046_n2088# 0.020511f
C113 source.n45 a_n2046_n2088# 0.016154f
C114 source.n46 a_n2046_n2088# 0.01157f
C115 source.n47 a_n2046_n2088# 0.512324f
C116 source.n48 a_n2046_n2088# 0.021532f
C117 source.n49 a_n2046_n2088# 0.01157f
C118 source.n50 a_n2046_n2088# 0.012251f
C119 source.n51 a_n2046_n2088# 0.027348f
C120 source.n52 a_n2046_n2088# 0.027348f
C121 source.n53 a_n2046_n2088# 0.012251f
C122 source.n54 a_n2046_n2088# 0.01157f
C123 source.n55 a_n2046_n2088# 0.021532f
C124 source.n56 a_n2046_n2088# 0.021532f
C125 source.n57 a_n2046_n2088# 0.01157f
C126 source.n58 a_n2046_n2088# 0.012251f
C127 source.n59 a_n2046_n2088# 0.027348f
C128 source.n60 a_n2046_n2088# 0.059203f
C129 source.n61 a_n2046_n2088# 0.012251f
C130 source.n62 a_n2046_n2088# 0.01157f
C131 source.n63 a_n2046_n2088# 0.049769f
C132 source.n64 a_n2046_n2088# 0.033126f
C133 source.n65 a_n2046_n2088# 0.130533f
C134 source.n66 a_n2046_n2088# 0.030265f
C135 source.n67 a_n2046_n2088# 0.021532f
C136 source.n68 a_n2046_n2088# 0.01157f
C137 source.n69 a_n2046_n2088# 0.027348f
C138 source.n70 a_n2046_n2088# 0.012251f
C139 source.n71 a_n2046_n2088# 0.021532f
C140 source.n72 a_n2046_n2088# 0.01157f
C141 source.n73 a_n2046_n2088# 0.027348f
C142 source.n74 a_n2046_n2088# 0.012251f
C143 source.n75 a_n2046_n2088# 0.09214f
C144 source.t0 a_n2046_n2088# 0.044573f
C145 source.n76 a_n2046_n2088# 0.020511f
C146 source.n77 a_n2046_n2088# 0.016154f
C147 source.n78 a_n2046_n2088# 0.01157f
C148 source.n79 a_n2046_n2088# 0.512324f
C149 source.n80 a_n2046_n2088# 0.021532f
C150 source.n81 a_n2046_n2088# 0.01157f
C151 source.n82 a_n2046_n2088# 0.012251f
C152 source.n83 a_n2046_n2088# 0.027348f
C153 source.n84 a_n2046_n2088# 0.027348f
C154 source.n85 a_n2046_n2088# 0.012251f
C155 source.n86 a_n2046_n2088# 0.01157f
C156 source.n87 a_n2046_n2088# 0.021532f
C157 source.n88 a_n2046_n2088# 0.021532f
C158 source.n89 a_n2046_n2088# 0.01157f
C159 source.n90 a_n2046_n2088# 0.012251f
C160 source.n91 a_n2046_n2088# 0.027348f
C161 source.n92 a_n2046_n2088# 0.059203f
C162 source.n93 a_n2046_n2088# 0.012251f
C163 source.n94 a_n2046_n2088# 0.01157f
C164 source.n95 a_n2046_n2088# 0.049769f
C165 source.n96 a_n2046_n2088# 0.033126f
C166 source.n97 a_n2046_n2088# 0.130533f
C167 source.t6 a_n2046_n2088# 0.10209f
C168 source.t2 a_n2046_n2088# 0.10209f
C169 source.n98 a_n2046_n2088# 0.795082f
C170 source.n99 a_n2046_n2088# 0.360933f
C171 source.n100 a_n2046_n2088# 0.030265f
C172 source.n101 a_n2046_n2088# 0.021532f
C173 source.n102 a_n2046_n2088# 0.01157f
C174 source.n103 a_n2046_n2088# 0.027348f
C175 source.n104 a_n2046_n2088# 0.012251f
C176 source.n105 a_n2046_n2088# 0.021532f
C177 source.n106 a_n2046_n2088# 0.01157f
C178 source.n107 a_n2046_n2088# 0.027348f
C179 source.n108 a_n2046_n2088# 0.012251f
C180 source.n109 a_n2046_n2088# 0.09214f
C181 source.t5 a_n2046_n2088# 0.044573f
C182 source.n110 a_n2046_n2088# 0.020511f
C183 source.n111 a_n2046_n2088# 0.016154f
C184 source.n112 a_n2046_n2088# 0.01157f
C185 source.n113 a_n2046_n2088# 0.512324f
C186 source.n114 a_n2046_n2088# 0.021532f
C187 source.n115 a_n2046_n2088# 0.01157f
C188 source.n116 a_n2046_n2088# 0.012251f
C189 source.n117 a_n2046_n2088# 0.027348f
C190 source.n118 a_n2046_n2088# 0.027348f
C191 source.n119 a_n2046_n2088# 0.012251f
C192 source.n120 a_n2046_n2088# 0.01157f
C193 source.n121 a_n2046_n2088# 0.021532f
C194 source.n122 a_n2046_n2088# 0.021532f
C195 source.n123 a_n2046_n2088# 0.01157f
C196 source.n124 a_n2046_n2088# 0.012251f
C197 source.n125 a_n2046_n2088# 0.027348f
C198 source.n126 a_n2046_n2088# 0.059203f
C199 source.n127 a_n2046_n2088# 0.012251f
C200 source.n128 a_n2046_n2088# 0.01157f
C201 source.n129 a_n2046_n2088# 0.049769f
C202 source.n130 a_n2046_n2088# 0.033126f
C203 source.n131 a_n2046_n2088# 0.88247f
C204 source.n132 a_n2046_n2088# 0.030265f
C205 source.n133 a_n2046_n2088# 0.021532f
C206 source.n134 a_n2046_n2088# 0.01157f
C207 source.n135 a_n2046_n2088# 0.027348f
C208 source.n136 a_n2046_n2088# 0.012251f
C209 source.n137 a_n2046_n2088# 0.021532f
C210 source.n138 a_n2046_n2088# 0.01157f
C211 source.n139 a_n2046_n2088# 0.027348f
C212 source.n140 a_n2046_n2088# 0.012251f
C213 source.n141 a_n2046_n2088# 0.09214f
C214 source.t12 a_n2046_n2088# 0.044573f
C215 source.n142 a_n2046_n2088# 0.020511f
C216 source.n143 a_n2046_n2088# 0.016154f
C217 source.n144 a_n2046_n2088# 0.01157f
C218 source.n145 a_n2046_n2088# 0.512324f
C219 source.n146 a_n2046_n2088# 0.021532f
C220 source.n147 a_n2046_n2088# 0.01157f
C221 source.n148 a_n2046_n2088# 0.012251f
C222 source.n149 a_n2046_n2088# 0.027348f
C223 source.n150 a_n2046_n2088# 0.027348f
C224 source.n151 a_n2046_n2088# 0.012251f
C225 source.n152 a_n2046_n2088# 0.01157f
C226 source.n153 a_n2046_n2088# 0.021532f
C227 source.n154 a_n2046_n2088# 0.021532f
C228 source.n155 a_n2046_n2088# 0.01157f
C229 source.n156 a_n2046_n2088# 0.012251f
C230 source.n157 a_n2046_n2088# 0.027348f
C231 source.n158 a_n2046_n2088# 0.059203f
C232 source.n159 a_n2046_n2088# 0.012251f
C233 source.n160 a_n2046_n2088# 0.01157f
C234 source.n161 a_n2046_n2088# 0.049769f
C235 source.n162 a_n2046_n2088# 0.033126f
C236 source.n163 a_n2046_n2088# 0.88247f
C237 source.t9 a_n2046_n2088# 0.10209f
C238 source.t11 a_n2046_n2088# 0.10209f
C239 source.n164 a_n2046_n2088# 0.795077f
C240 source.n165 a_n2046_n2088# 0.360938f
C241 source.n166 a_n2046_n2088# 0.030265f
C242 source.n167 a_n2046_n2088# 0.021532f
C243 source.n168 a_n2046_n2088# 0.01157f
C244 source.n169 a_n2046_n2088# 0.027348f
C245 source.n170 a_n2046_n2088# 0.012251f
C246 source.n171 a_n2046_n2088# 0.021532f
C247 source.n172 a_n2046_n2088# 0.01157f
C248 source.n173 a_n2046_n2088# 0.027348f
C249 source.n174 a_n2046_n2088# 0.012251f
C250 source.n175 a_n2046_n2088# 0.09214f
C251 source.t10 a_n2046_n2088# 0.044573f
C252 source.n176 a_n2046_n2088# 0.020511f
C253 source.n177 a_n2046_n2088# 0.016154f
C254 source.n178 a_n2046_n2088# 0.01157f
C255 source.n179 a_n2046_n2088# 0.512324f
C256 source.n180 a_n2046_n2088# 0.021532f
C257 source.n181 a_n2046_n2088# 0.01157f
C258 source.n182 a_n2046_n2088# 0.012251f
C259 source.n183 a_n2046_n2088# 0.027348f
C260 source.n184 a_n2046_n2088# 0.027348f
C261 source.n185 a_n2046_n2088# 0.012251f
C262 source.n186 a_n2046_n2088# 0.01157f
C263 source.n187 a_n2046_n2088# 0.021532f
C264 source.n188 a_n2046_n2088# 0.021532f
C265 source.n189 a_n2046_n2088# 0.01157f
C266 source.n190 a_n2046_n2088# 0.012251f
C267 source.n191 a_n2046_n2088# 0.027348f
C268 source.n192 a_n2046_n2088# 0.059203f
C269 source.n193 a_n2046_n2088# 0.012251f
C270 source.n194 a_n2046_n2088# 0.01157f
C271 source.n195 a_n2046_n2088# 0.049769f
C272 source.n196 a_n2046_n2088# 0.033126f
C273 source.n197 a_n2046_n2088# 0.130533f
C274 source.n198 a_n2046_n2088# 0.030265f
C275 source.n199 a_n2046_n2088# 0.021532f
C276 source.n200 a_n2046_n2088# 0.01157f
C277 source.n201 a_n2046_n2088# 0.027348f
C278 source.n202 a_n2046_n2088# 0.012251f
C279 source.n203 a_n2046_n2088# 0.021532f
C280 source.n204 a_n2046_n2088# 0.01157f
C281 source.n205 a_n2046_n2088# 0.027348f
C282 source.n206 a_n2046_n2088# 0.012251f
C283 source.n207 a_n2046_n2088# 0.09214f
C284 source.t4 a_n2046_n2088# 0.044573f
C285 source.n208 a_n2046_n2088# 0.020511f
C286 source.n209 a_n2046_n2088# 0.016154f
C287 source.n210 a_n2046_n2088# 0.01157f
C288 source.n211 a_n2046_n2088# 0.512324f
C289 source.n212 a_n2046_n2088# 0.021532f
C290 source.n213 a_n2046_n2088# 0.01157f
C291 source.n214 a_n2046_n2088# 0.012251f
C292 source.n215 a_n2046_n2088# 0.027348f
C293 source.n216 a_n2046_n2088# 0.027348f
C294 source.n217 a_n2046_n2088# 0.012251f
C295 source.n218 a_n2046_n2088# 0.01157f
C296 source.n219 a_n2046_n2088# 0.021532f
C297 source.n220 a_n2046_n2088# 0.021532f
C298 source.n221 a_n2046_n2088# 0.01157f
C299 source.n222 a_n2046_n2088# 0.012251f
C300 source.n223 a_n2046_n2088# 0.027348f
C301 source.n224 a_n2046_n2088# 0.059203f
C302 source.n225 a_n2046_n2088# 0.012251f
C303 source.n226 a_n2046_n2088# 0.01157f
C304 source.n227 a_n2046_n2088# 0.049769f
C305 source.n228 a_n2046_n2088# 0.033126f
C306 source.n229 a_n2046_n2088# 0.130533f
C307 source.t3 a_n2046_n2088# 0.10209f
C308 source.t7 a_n2046_n2088# 0.10209f
C309 source.n230 a_n2046_n2088# 0.795077f
C310 source.n231 a_n2046_n2088# 0.360938f
C311 source.n232 a_n2046_n2088# 0.030265f
C312 source.n233 a_n2046_n2088# 0.021532f
C313 source.n234 a_n2046_n2088# 0.01157f
C314 source.n235 a_n2046_n2088# 0.027348f
C315 source.n236 a_n2046_n2088# 0.012251f
C316 source.n237 a_n2046_n2088# 0.021532f
C317 source.n238 a_n2046_n2088# 0.01157f
C318 source.n239 a_n2046_n2088# 0.027348f
C319 source.n240 a_n2046_n2088# 0.012251f
C320 source.n241 a_n2046_n2088# 0.09214f
C321 source.t1 a_n2046_n2088# 0.044573f
C322 source.n242 a_n2046_n2088# 0.020511f
C323 source.n243 a_n2046_n2088# 0.016154f
C324 source.n244 a_n2046_n2088# 0.01157f
C325 source.n245 a_n2046_n2088# 0.512324f
C326 source.n246 a_n2046_n2088# 0.021532f
C327 source.n247 a_n2046_n2088# 0.01157f
C328 source.n248 a_n2046_n2088# 0.012251f
C329 source.n249 a_n2046_n2088# 0.027348f
C330 source.n250 a_n2046_n2088# 0.027348f
C331 source.n251 a_n2046_n2088# 0.012251f
C332 source.n252 a_n2046_n2088# 0.01157f
C333 source.n253 a_n2046_n2088# 0.021532f
C334 source.n254 a_n2046_n2088# 0.021532f
C335 source.n255 a_n2046_n2088# 0.01157f
C336 source.n256 a_n2046_n2088# 0.012251f
C337 source.n257 a_n2046_n2088# 0.027348f
C338 source.n258 a_n2046_n2088# 0.059203f
C339 source.n259 a_n2046_n2088# 0.012251f
C340 source.n260 a_n2046_n2088# 0.01157f
C341 source.n261 a_n2046_n2088# 0.049769f
C342 source.n262 a_n2046_n2088# 0.033126f
C343 source.n263 a_n2046_n2088# 0.284895f
C344 source.n264 a_n2046_n2088# 0.902264f
C345 drain_left.t6 a_n2046_n2088# 0.122108f
C346 drain_left.t3 a_n2046_n2088# 0.122108f
C347 drain_left.n0 a_n2046_n2088# 1.02112f
C348 drain_left.t1 a_n2046_n2088# 0.122108f
C349 drain_left.t4 a_n2046_n2088# 0.122108f
C350 drain_left.n1 a_n2046_n2088# 1.02112f
C351 drain_left.n2 a_n2046_n2088# 1.73093f
C352 drain_left.t5 a_n2046_n2088# 0.122108f
C353 drain_left.t2 a_n2046_n2088# 0.122108f
C354 drain_left.n3 a_n2046_n2088# 1.02526f
C355 drain_left.t7 a_n2046_n2088# 0.122108f
C356 drain_left.t0 a_n2046_n2088# 0.122108f
C357 drain_left.n4 a_n2046_n2088# 1.01838f
C358 drain_left.n5 a_n2046_n2088# 1.0391f
C359 plus.n0 a_n2046_n2088# 0.054585f
C360 plus.t2 a_n2046_n2088# 0.71191f
C361 plus.t0 a_n2046_n2088# 0.649623f
C362 plus.n1 a_n2046_n2088# 0.033039f
C363 plus.t7 a_n2046_n2088# 0.737221f
C364 plus.n2 a_n2046_n2088# 0.325271f
C365 plus.t1 a_n2046_n2088# 0.649623f
C366 plus.n3 a_n2046_n2088# 0.303128f
C367 plus.n4 a_n2046_n2088# 0.055783f
C368 plus.n5 a_n2046_n2088# 0.17512f
C369 plus.n6 a_n2046_n2088# 0.040907f
C370 plus.n7 a_n2046_n2088# 0.040907f
C371 plus.n8 a_n2046_n2088# 0.055783f
C372 plus.n9 a_n2046_n2088# 0.266727f
C373 plus.n10 a_n2046_n2088# 0.056109f
C374 plus.n11 a_n2046_n2088# 0.330009f
C375 plus.n12 a_n2046_n2088# 0.402574f
C376 plus.n13 a_n2046_n2088# 0.054585f
C377 plus.t3 a_n2046_n2088# 0.71191f
C378 plus.t6 a_n2046_n2088# 0.649623f
C379 plus.n14 a_n2046_n2088# 0.033039f
C380 plus.t5 a_n2046_n2088# 0.737221f
C381 plus.n15 a_n2046_n2088# 0.325271f
C382 plus.t4 a_n2046_n2088# 0.649623f
C383 plus.n16 a_n2046_n2088# 0.303128f
C384 plus.n17 a_n2046_n2088# 0.055783f
C385 plus.n18 a_n2046_n2088# 0.17512f
C386 plus.n19 a_n2046_n2088# 0.040907f
C387 plus.n20 a_n2046_n2088# 0.040907f
C388 plus.n21 a_n2046_n2088# 0.055783f
C389 plus.n22 a_n2046_n2088# 0.266727f
C390 plus.n23 a_n2046_n2088# 0.056109f
C391 plus.n24 a_n2046_n2088# 0.330009f
C392 plus.n25 a_n2046_n2088# 1.14032f
.ends

