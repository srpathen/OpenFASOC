* NGSPICE file created from opamp426.ext - technology: sky130A

.subckt opamp426 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 gnd.t349 commonsourceibias.t80 CSoutput.t114 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X1 CSoutput.t48 a_n8300_8799.t36 vdd.t299 vdd.t243 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X2 a_n2140_13878.t23 a_n2318_13878.t31 a_n2318_13878.t32 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 commonsourceibias.t13 commonsourceibias.t12 gnd.t348 gnd.t313 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X4 a_n2140_13878.t7 a_n2318_13878.t52 vdd.t24 vdd.t23 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X5 vdd.t298 a_n8300_8799.t37 CSoutput.t0 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 outputibias.t7 outputibias.t6 gnd.t58 gnd.t57 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X7 gnd.t189 gnd.t187 gnd.t188 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 CSoutput.t53 a_n8300_8799.t38 vdd.t297 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X9 CSoutput.t188 a_n8300_8799.t39 vdd.t296 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X10 gnd.t347 commonsourceibias.t81 CSoutput.t113 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X11 CSoutput.t200 a_n2318_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X12 gnd.t346 commonsourceibias.t82 CSoutput.t112 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X13 gnd.t345 commonsourceibias.t10 commonsourceibias.t11 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X14 gnd.t344 commonsourceibias.t83 CSoutput.t111 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 a_n2318_8322.t27 a_n2318_13878.t53 a_n8300_8799.t5 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X16 gnd.t343 commonsourceibias.t84 CSoutput.t110 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X17 output.t15 CSoutput.t201 vdd.t13 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X18 CSoutput.t82 a_n8300_8799.t40 vdd.t295 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 outputibias.t5 outputibias.t4 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X20 gnd.t186 gnd.t184 plus.t4 gnd.t185 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X21 a_n8300_8799.t31 plus.t5 a_n2903_n3924.t25 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X22 gnd.t342 commonsourceibias.t85 CSoutput.t109 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 vdd.t294 a_n8300_8799.t41 CSoutput.t76 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 minus.t4 gnd.t181 gnd.t183 gnd.t182 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X25 gnd.t341 commonsourceibias.t8 commonsourceibias.t9 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X26 a_n8300_8799.t14 a_n2318_13878.t54 a_n2318_8322.t26 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X27 vdd.t293 a_n8300_8799.t42 CSoutput.t194 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X28 vdd.t292 a_n8300_8799.t43 CSoutput.t29 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X29 CSoutput.t2 a_n8300_8799.t44 vdd.t291 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X30 vdd.t290 a_n8300_8799.t45 CSoutput.t75 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X31 a_n8300_8799.t15 a_n2318_13878.t55 a_n2318_8322.t25 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X32 a_n8300_8799.t3 plus.t6 a_n2903_n3924.t24 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X33 CSoutput.t108 commonsourceibias.t86 gnd.t340 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X34 gnd.t339 commonsourceibias.t50 commonsourceibias.t51 gnd.t302 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 vdd.t101 vdd.t99 vdd.t100 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X36 CSoutput.t149 commonsourceibias.t87 gnd.t338 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X37 CSoutput.t61 a_n8300_8799.t46 vdd.t289 vdd.t243 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X38 vdd.t11 CSoutput.t202 output.t14 gnd.t17 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X39 CSoutput.t148 commonsourceibias.t88 gnd.t337 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 CSoutput.t80 a_n8300_8799.t47 vdd.t288 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X41 CSoutput.t147 commonsourceibias.t89 gnd.t336 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 a_n2903_n3924.t41 diffpairibias.t16 gnd.t65 gnd.t64 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X43 a_n2903_n3924.t3 minus.t5 a_n2318_13878.t3 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X44 CSoutput.t43 a_n8300_8799.t48 vdd.t287 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X45 a_n2903_n3924.t23 plus.t7 a_n8300_8799.t32 gnd.t350 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X46 vdd.t286 a_n8300_8799.t49 CSoutput.t27 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X47 a_n2318_13878.t49 minus.t6 a_n2903_n3924.t45 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X48 CSoutput.t146 commonsourceibias.t90 gnd.t335 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 a_n2903_n3924.t22 plus.t8 a_n8300_8799.t34 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X50 a_n2903_n3924.t4 minus.t7 a_n2318_13878.t4 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X51 CSoutput.t42 a_n8300_8799.t50 vdd.t285 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X52 gnd.t334 commonsourceibias.t48 commonsourceibias.t49 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X53 outputibias.t3 outputibias.t2 gnd.t36 gnd.t35 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X54 output.t13 CSoutput.t203 vdd.t6 gnd.t16 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X55 a_n2140_13878.t22 a_n2318_13878.t37 a_n2318_13878.t38 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X56 CSoutput.t145 commonsourceibias.t91 gnd.t333 gnd.t313 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X57 a_n2318_13878.t18 a_n2318_13878.t17 a_n2140_13878.t21 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X58 commonsourceibias.t47 commonsourceibias.t46 gnd.t332 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X59 CSoutput.t204 a_n2318_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X60 CSoutput.t26 a_n8300_8799.t51 vdd.t284 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 vdd.t98 vdd.t96 vdd.t97 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X62 a_n2903_n3924.t33 minus.t8 a_n2318_13878.t9 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X63 vdd.t283 a_n8300_8799.t52 CSoutput.t66 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 diffpairibias.t15 diffpairibias.t14 gnd.t78 gnd.t77 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X65 a_n8300_8799.t20 a_n2318_13878.t56 a_n2318_8322.t24 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X66 gnd.t180 gnd.t178 gnd.t179 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X67 gnd.t177 gnd.t175 gnd.t176 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X68 CSoutput.t180 a_n8300_8799.t53 vdd.t282 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X69 gnd.t174 gnd.t173 plus.t3 gnd.t111 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X70 vdd.t281 a_n8300_8799.t54 CSoutput.t47 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X71 vdd.t280 a_n8300_8799.t55 CSoutput.t25 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 minus.t3 gnd.t170 gnd.t172 gnd.t171 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X73 gnd.t331 commonsourceibias.t92 CSoutput.t144 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 diffpairibias.t13 diffpairibias.t12 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X75 gnd.t330 commonsourceibias.t93 CSoutput.t143 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 CSoutput.t88 a_n8300_8799.t56 vdd.t279 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 output.t12 CSoutput.t205 vdd.t16 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X78 commonsourceibias.t45 commonsourceibias.t44 gnd.t329 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 gnd.t328 commonsourceibias.t94 CSoutput.t142 gnd.t302 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 vdd.t278 a_n8300_8799.t57 CSoutput.t62 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X81 CSoutput.t81 a_n8300_8799.t58 vdd.t277 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 vdd.t95 vdd.t93 vdd.t94 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X83 CSoutput.t10 a_n8300_8799.t59 vdd.t276 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X84 CSoutput.t74 a_n8300_8799.t60 vdd.t275 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X85 CSoutput.t46 a_n8300_8799.t61 vdd.t274 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 commonsourceibias.t43 commonsourceibias.t42 gnd.t327 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X87 gnd.t326 commonsourceibias.t95 CSoutput.t141 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 output.t11 CSoutput.t206 vdd.t7 gnd.t14 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X89 commonsourceibias.t41 commonsourceibias.t40 gnd.t325 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X90 a_n8300_8799.t17 plus.t9 a_n2903_n3924.t21 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X91 gnd.t324 commonsourceibias.t96 CSoutput.t122 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 CSoutput.t121 commonsourceibias.t97 gnd.t323 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X93 gnd.t322 commonsourceibias.t24 commonsourceibias.t25 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 a_n2903_n3924.t27 diffpairibias.t17 gnd.t28 gnd.t27 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X95 CSoutput.t207 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X96 vdd.t273 a_n8300_8799.t62 CSoutput.t86 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 a_n2903_n3924.t31 minus.t9 a_n2318_13878.t7 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X98 vdd.t272 a_n8300_8799.t63 CSoutput.t185 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 a_n2318_13878.t26 a_n2318_13878.t25 a_n2140_13878.t20 vdd.t19 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X100 vdd.t271 a_n8300_8799.t64 CSoutput.t11 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 vdd.t270 a_n8300_8799.t65 CSoutput.t8 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X102 a_n8300_8799.t21 a_n2318_13878.t57 a_n2318_8322.t23 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X103 vdd.t269 a_n8300_8799.t66 CSoutput.t19 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X104 a_n2318_13878.t24 a_n2318_13878.t23 a_n2140_13878.t19 vdd.t127 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X105 gnd.t321 commonsourceibias.t22 commonsourceibias.t23 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X106 a_n2318_13878.t50 minus.t10 a_n2903_n3924.t46 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X107 a_n2903_n3924.t20 plus.t10 a_n8300_8799.t29 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X108 commonsourceibias.t21 commonsourceibias.t20 gnd.t320 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 CSoutput.t157 commonsourceibias.t98 gnd.t285 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t268 a_n8300_8799.t67 CSoutput.t183 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 CSoutput.t184 a_n8300_8799.t68 vdd.t267 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X112 CSoutput.t120 commonsourceibias.t99 gnd.t319 gnd.t281 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X113 vdd.t4 CSoutput.t208 output.t10 gnd.t13 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X114 a_n2903_n3924.t38 minus.t11 a_n2318_13878.t12 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X115 vdd.t92 vdd.t90 vdd.t91 vdd.t39 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X116 vdd.t89 vdd.t87 vdd.t88 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X117 CSoutput.t119 commonsourceibias.t100 gnd.t318 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 CSoutput.t96 a_n8300_8799.t69 vdd.t266 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X119 vdd.t86 vdd.t83 vdd.t85 vdd.t84 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X120 gnd.t317 commonsourceibias.t101 CSoutput.t118 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X121 commonsourceibias.t19 commonsourceibias.t18 gnd.t316 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 CSoutput.t117 commonsourceibias.t102 gnd.t315 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X123 CSoutput.t116 commonsourceibias.t103 gnd.t314 gnd.t313 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 CSoutput.t4 a_n8300_8799.t70 vdd.t265 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 vdd.t264 a_n8300_8799.t71 CSoutput.t54 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X126 vdd.t119 a_n2318_13878.t58 a_n2318_8322.t11 vdd.t118 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X127 a_n2318_13878.t36 a_n2318_13878.t35 a_n2140_13878.t18 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X128 vdd.t82 vdd.t80 vdd.t81 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X129 a_n2318_8322.t10 a_n2318_13878.t59 vdd.t121 vdd.t120 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X130 a_n2903_n3924.t35 diffpairibias.t18 gnd.t47 gnd.t46 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X131 CSoutput.t85 a_n8300_8799.t72 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X132 CSoutput.t20 a_n8300_8799.t73 vdd.t261 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X133 a_n2318_13878.t8 minus.t12 a_n2903_n3924.t32 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X134 gnd.t312 commonsourceibias.t104 CSoutput.t115 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X135 commonsourceibias.t17 commonsourceibias.t16 gnd.t311 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X136 commonsourceibias.t15 commonsourceibias.t14 gnd.t310 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X137 a_n2903_n3924.t19 plus.t11 a_n8300_8799.t2 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X138 vdd.t111 a_n2318_13878.t60 a_n2140_13878.t6 vdd.t110 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X139 vdd.t79 vdd.t76 vdd.t78 vdd.t77 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X140 gnd.t309 commonsourceibias.t6 commonsourceibias.t7 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X141 vdd.t260 a_n8300_8799.t74 CSoutput.t57 vdd.t259 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X142 vdd.t258 a_n8300_8799.t75 CSoutput.t52 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X143 gnd.t308 commonsourceibias.t105 CSoutput.t107 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X144 vdd.t257 a_n8300_8799.t76 CSoutput.t24 vdd.t256 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X145 gnd.t307 commonsourceibias.t4 commonsourceibias.t5 gnd.t306 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 outputibias.t1 outputibias.t0 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X147 a_n8300_8799.t0 plus.t12 a_n2903_n3924.t18 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X148 vdd.t75 vdd.t72 vdd.t74 vdd.t73 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X149 a_n2318_8322.t9 a_n2318_13878.t61 vdd.t113 vdd.t112 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X150 a_n8300_8799.t12 a_n2318_13878.t62 a_n2318_8322.t22 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X151 commonsourceibias.t3 commonsourceibias.t2 gnd.t305 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X152 gnd.t304 commonsourceibias.t106 CSoutput.t106 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 a_n2318_13878.t6 minus.t13 a_n2903_n3924.t30 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X154 gnd.t303 commonsourceibias.t107 CSoutput.t105 gnd.t302 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X155 gnd.t301 commonsourceibias.t108 CSoutput.t104 gnd.t258 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X156 CSoutput.t72 a_n8300_8799.t77 vdd.t255 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X157 diffpairibias.t11 diffpairibias.t10 gnd.t69 gnd.t68 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 vdd.t254 a_n8300_8799.t78 CSoutput.t97 vdd.t253 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X159 a_n2318_13878.t28 a_n2318_13878.t27 a_n2140_13878.t17 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X160 vdd.t252 a_n8300_8799.t79 CSoutput.t69 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X161 a_n8300_8799.t13 a_n2318_13878.t63 a_n2318_8322.t21 vdd.t109 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X162 CSoutput.t91 a_n8300_8799.t80 vdd.t251 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 gnd.t300 commonsourceibias.t109 CSoutput.t103 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 a_n2140_13878.t16 a_n2318_13878.t29 a_n2318_13878.t30 vdd.t25 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X165 output.t19 outputibias.t8 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X166 vdd.t71 vdd.t69 vdd.t70 vdd.t39 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X167 gnd.t299 commonsourceibias.t110 CSoutput.t102 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X168 CSoutput.t101 commonsourceibias.t111 gnd.t297 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X169 plus.t2 gnd.t167 gnd.t169 gnd.t168 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X170 commonsourceibias.t1 commonsourceibias.t0 gnd.t296 gnd.t295 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 gnd.t166 gnd.t164 minus.t2 gnd.t165 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X172 CSoutput.t92 a_n8300_8799.t81 vdd.t250 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 a_n2318_13878.t1 minus.t14 a_n2903_n3924.t1 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X174 gnd.t294 commonsourceibias.t112 CSoutput.t100 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X175 vdd.t105 a_n2318_13878.t64 a_n2318_8322.t8 vdd.t104 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X176 a_n2140_13878.t15 a_n2318_13878.t47 a_n2318_13878.t48 vdd.t114 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X177 CSoutput.t163 commonsourceibias.t113 gnd.t293 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 vdd.t249 a_n8300_8799.t82 CSoutput.t93 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 a_n2318_13878.t42 a_n2318_13878.t41 a_n2140_13878.t14 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X180 vdd.t248 a_n8300_8799.t83 CSoutput.t94 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X181 CSoutput.t162 commonsourceibias.t114 gnd.t292 gnd.t281 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X182 a_n2903_n3924.t29 diffpairibias.t19 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X183 gnd.t163 gnd.t160 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 a_n2903_n3924.t40 diffpairibias.t20 gnd.t63 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X185 a_n2318_13878.t11 minus.t15 a_n2903_n3924.t37 gnd.t51 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X186 vdd.t9 CSoutput.t209 output.t9 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X187 CSoutput.t161 commonsourceibias.t115 gnd.t291 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X188 CSoutput.t160 commonsourceibias.t116 gnd.t290 gnd.t289 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X189 vdd.t247 a_n8300_8799.t84 CSoutput.t95 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 vdd.t246 a_n8300_8799.t85 CSoutput.t98 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X191 gnd.t288 commonsourceibias.t117 CSoutput.t159 gnd.t287 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X192 gnd.t286 commonsourceibias.t118 CSoutput.t158 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 CSoutput.t156 commonsourceibias.t119 gnd.t284 gnd.t283 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X194 gnd.t159 gnd.t157 minus.t1 gnd.t158 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X195 commonsourceibias.t65 commonsourceibias.t64 gnd.t282 gnd.t281 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 CSoutput.t155 commonsourceibias.t120 gnd.t280 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X197 gnd.t156 gnd.t154 gnd.t155 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X198 gnd.t153 gnd.t150 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X199 gnd.t149 gnd.t147 gnd.t148 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X200 CSoutput.t71 a_n8300_8799.t86 vdd.t245 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 gnd.t279 commonsourceibias.t121 CSoutput.t154 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X202 CSoutput.t186 a_n8300_8799.t87 vdd.t244 vdd.t243 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X203 a_n2318_13878.t0 minus.t16 a_n2903_n3924.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X204 CSoutput.t37 a_n8300_8799.t88 vdd.t242 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X205 gnd.t146 gnd.t144 gnd.t145 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X206 CSoutput.t150 commonsourceibias.t122 gnd.t197 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 diffpairibias.t9 diffpairibias.t8 gnd.t32 gnd.t31 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X208 a_n2140_13878.t5 a_n2318_13878.t65 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X209 vdd.t103 a_n2318_13878.t66 a_n2140_13878.t4 vdd.t102 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X210 CSoutput.t193 a_n8300_8799.t89 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X211 a_n2903_n3924.t17 plus.t13 a_n8300_8799.t1 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X212 vdd.t239 a_n8300_8799.t90 CSoutput.t41 vdd.t238 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X213 vdd.t237 a_n8300_8799.t91 CSoutput.t99 vdd.t236 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X214 gnd.t278 commonsourceibias.t123 CSoutput.t153 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 CSoutput.t133 commonsourceibias.t124 gnd.t277 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X216 CSoutput.t15 a_n8300_8799.t92 vdd.t235 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X217 a_n2903_n3924.t36 minus.t17 a_n2318_13878.t10 gnd.t50 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X218 a_n2140_13878.t13 a_n2318_13878.t43 a_n2318_13878.t44 vdd.t122 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X219 gnd.t276 commonsourceibias.t30 commonsourceibias.t31 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X220 a_n2903_n3924.t16 plus.t14 a_n8300_8799.t30 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X221 gnd.t275 commonsourceibias.t125 CSoutput.t132 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 gnd.t273 commonsourceibias.t126 CSoutput.t130 gnd.t258 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X223 a_n2903_n3924.t43 minus.t18 a_n2318_13878.t15 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X224 a_n8300_8799.t7 plus.t15 a_n2903_n3924.t15 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X225 vdd.t234 a_n8300_8799.t93 CSoutput.t16 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 gnd.t274 commonsourceibias.t127 CSoutput.t131 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 a_n2318_8322.t20 a_n2318_13878.t67 a_n8300_8799.t11 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X228 vdd.t17 CSoutput.t210 output.t8 gnd.t11 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X229 CSoutput.t65 a_n8300_8799.t94 vdd.t233 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X230 diffpairibias.t7 diffpairibias.t6 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X231 CSoutput.t129 commonsourceibias.t128 gnd.t272 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X232 vdd.t232 a_n8300_8799.t95 CSoutput.t36 vdd.t231 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X233 vdd.t68 vdd.t66 vdd.t67 vdd.t49 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X234 vdd.t137 a_n2318_13878.t68 a_n2318_8322.t7 vdd.t136 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X235 gnd.t271 commonsourceibias.t28 commonsourceibias.t29 gnd.t270 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 vdd.t230 a_n8300_8799.t96 CSoutput.t17 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X237 vdd.t229 a_n8300_8799.t97 CSoutput.t90 vdd.t228 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X238 gnd.t143 gnd.t141 gnd.t142 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X239 CSoutput.t128 commonsourceibias.t129 gnd.t269 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 gnd.t268 commonsourceibias.t130 CSoutput.t127 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 CSoutput.t126 commonsourceibias.t131 gnd.t267 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X242 CSoutput.t5 a_n8300_8799.t98 vdd.t227 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X243 a_n2140_13878.t3 a_n2318_13878.t69 vdd.t139 vdd.t138 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X244 vdd.t65 vdd.t62 vdd.t64 vdd.t63 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X245 vdd.t61 vdd.t59 vdd.t60 vdd.t49 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X246 plus.t1 gnd.t138 gnd.t140 gnd.t139 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X247 vdd.t226 a_n8300_8799.t99 CSoutput.t12 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X248 CSoutput.t18 a_n8300_8799.t100 vdd.t225 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X249 CSoutput.t13 a_n8300_8799.t101 vdd.t224 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X250 CSoutput.t6 a_n8300_8799.t102 vdd.t223 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X251 gnd.t266 commonsourceibias.t26 commonsourceibias.t27 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X252 gnd.t137 gnd.t135 minus.t0 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X253 gnd.t134 gnd.t131 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X254 vdd.t222 a_n8300_8799.t103 CSoutput.t28 vdd.t196 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X255 a_n2903_n3924.t26 diffpairibias.t21 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X256 CSoutput.t125 commonsourceibias.t132 gnd.t265 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 a_n2318_8322.t19 a_n2318_13878.t70 a_n8300_8799.t28 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X258 vdd.t135 a_n2318_13878.t71 a_n2318_8322.t6 vdd.t134 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X259 CSoutput.t211 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X260 CSoutput.t60 a_n8300_8799.t104 vdd.t221 vdd.t220 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X261 vdd.t219 a_n8300_8799.t105 CSoutput.t70 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X262 CSoutput.t22 a_n8300_8799.t106 vdd.t218 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 CSoutput.t124 commonsourceibias.t133 gnd.t264 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 vdd.t217 a_n8300_8799.t107 CSoutput.t7 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 gnd.t263 commonsourceibias.t134 CSoutput.t123 gnd.t262 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X266 vdd.t216 a_n8300_8799.t108 CSoutput.t181 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X267 gnd.t261 commonsourceibias.t38 commonsourceibias.t39 gnd.t260 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X268 gnd.t259 commonsourceibias.t36 commonsourceibias.t37 gnd.t258 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X269 vdd.t12 CSoutput.t212 output.t7 gnd.t10 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X270 CSoutput.t140 commonsourceibias.t135 gnd.t257 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X271 vdd.t58 vdd.t56 vdd.t57 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X272 output.t6 CSoutput.t213 vdd.t15 gnd.t9 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X273 CSoutput.t139 commonsourceibias.t136 gnd.t256 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X274 gnd.t255 commonsourceibias.t137 CSoutput.t138 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X275 a_n2903_n3924.t14 plus.t16 a_n8300_8799.t4 gnd.t39 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X276 vdd.t55 vdd.t52 vdd.t54 vdd.t53 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X277 gnd.t130 gnd.t128 gnd.t129 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X278 vdd.t215 a_n8300_8799.t109 CSoutput.t73 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X279 gnd.t127 gnd.t124 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X280 a_n8300_8799.t8 plus.t17 a_n2903_n3924.t13 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X281 CSoutput.t34 a_n8300_8799.t110 vdd.t214 vdd.t213 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X282 a_n2903_n3924.t42 minus.t19 a_n2318_13878.t14 gnd.t76 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X283 a_n2140_13878.t12 a_n2318_13878.t33 a_n2318_13878.t34 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X284 CSoutput.t182 a_n8300_8799.t111 vdd.t212 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 gnd.t123 gnd.t121 gnd.t122 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X286 CSoutput.t137 commonsourceibias.t138 gnd.t254 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X287 a_n2318_8322.t18 a_n2318_13878.t72 a_n8300_8799.t27 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X288 vdd.t51 vdd.t48 vdd.t50 vdd.t49 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X289 diffpairibias.t5 diffpairibias.t4 gnd.t67 gnd.t66 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X290 CSoutput.t214 a_n2318_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X291 a_n2903_n3924.t47 minus.t20 a_n2318_13878.t51 gnd.t350 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X292 a_n8300_8799.t6 plus.t18 a_n2903_n3924.t12 gnd.t41 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X293 commonsourceibias.t35 commonsourceibias.t34 gnd.t253 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 CSoutput.t21 a_n8300_8799.t112 vdd.t211 vdd.t210 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X295 CSoutput.t89 a_n8300_8799.t113 vdd.t209 vdd.t208 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X296 CSoutput.t32 a_n8300_8799.t114 vdd.t207 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X297 vdd.t206 a_n8300_8799.t115 CSoutput.t51 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X298 gnd.t252 commonsourceibias.t139 CSoutput.t136 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 CSoutput.t135 commonsourceibias.t140 gnd.t250 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X300 vdd.t205 a_n8300_8799.t116 CSoutput.t1 vdd.t204 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X301 a_n2318_8322.t5 a_n2318_13878.t73 vdd.t133 vdd.t132 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X302 gnd.t249 commonsourceibias.t32 commonsourceibias.t33 gnd.t248 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X303 gnd.t247 commonsourceibias.t141 CSoutput.t134 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 CSoutput.t23 a_n8300_8799.t117 vdd.t203 vdd.t202 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X305 CSoutput.t35 a_n8300_8799.t118 vdd.t201 vdd.t200 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 a_n2903_n3924.t11 plus.t19 a_n8300_8799.t35 gnd.t43 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X307 vdd.t47 vdd.t45 vdd.t46 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X308 vdd.t199 a_n8300_8799.t119 CSoutput.t14 vdd.t196 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X309 gnd.t120 gnd.t118 gnd.t119 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X310 output.t18 outputibias.t9 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X311 CSoutput.t58 a_n8300_8799.t120 vdd.t198 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X312 CSoutput.t177 commonsourceibias.t142 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 vdd.t126 a_n2318_13878.t74 a_n2140_13878.t2 vdd.t125 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X314 vdd.t197 a_n8300_8799.t121 CSoutput.t187 vdd.t196 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X315 CSoutput.t33 a_n8300_8799.t122 vdd.t195 vdd.t194 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 output.t5 CSoutput.t215 vdd.t14 gnd.t8 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X317 CSoutput.t198 a_n8300_8799.t123 vdd.t193 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X318 gnd.t117 gnd.t114 gnd.t116 gnd.t115 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X319 vdd.t5 CSoutput.t216 output.t4 gnd.t7 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X320 gnd.t195 commonsourceibias.t143 CSoutput.t179 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X321 gnd.t113 gnd.t110 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X322 CSoutput.t176 commonsourceibias.t144 gnd.t244 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 CSoutput.t175 commonsourceibias.t145 gnd.t243 gnd.t242 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X324 vdd.t192 a_n8300_8799.t124 CSoutput.t38 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X325 gnd.t241 commonsourceibias.t76 commonsourceibias.t77 gnd.t240 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 vdd.t190 a_n8300_8799.t125 CSoutput.t192 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X327 output.t17 outputibias.t10 gnd.t75 gnd.t74 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X328 a_n2903_n3924.t39 minus.t21 a_n2318_13878.t13 gnd.t24 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X329 vdd.t44 vdd.t42 vdd.t43 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X330 a_n2318_8322.t17 a_n2318_13878.t75 a_n8300_8799.t22 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X331 CSoutput.t9 a_n8300_8799.t126 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X332 a_n8300_8799.t26 a_n2318_13878.t76 a_n2318_8322.t16 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X333 vdd.t187 a_n8300_8799.t127 CSoutput.t39 vdd.t186 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X334 a_n2140_13878.t1 a_n2318_13878.t77 vdd.t131 vdd.t130 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X335 output.t16 outputibias.t11 gnd.t56 gnd.t55 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X336 vdd.t10 CSoutput.t217 output.t3 gnd.t6 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X337 vdd.t185 a_n8300_8799.t128 CSoutput.t30 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X338 CSoutput.t83 a_n8300_8799.t129 vdd.t184 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 a_n8300_8799.t16 plus.t20 a_n2903_n3924.t10 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X340 CSoutput.t174 commonsourceibias.t146 gnd.t239 gnd.t238 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X341 gnd.t109 gnd.t106 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X342 a_n2318_8322.t15 a_n2318_13878.t78 a_n8300_8799.t24 vdd.t18 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X343 a_n2318_13878.t16 minus.t22 a_n2903_n3924.t44 gnd.t59 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X344 vdd.t182 a_n8300_8799.t130 CSoutput.t50 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 CSoutput.t64 a_n8300_8799.t131 vdd.t180 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X346 CSoutput.t189 a_n8300_8799.t132 vdd.t178 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X347 CSoutput.t195 a_n8300_8799.t133 vdd.t177 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 output.t2 CSoutput.t218 vdd.t3 gnd.t5 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X349 a_n2140_13878.t11 a_n2318_13878.t45 a_n2318_13878.t46 vdd.t108 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X350 commonsourceibias.t75 commonsourceibias.t74 gnd.t237 gnd.t236 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X351 gnd.t226 commonsourceibias.t147 CSoutput.t169 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 vdd.t176 a_n8300_8799.t134 CSoutput.t63 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X353 gnd.t235 commonsourceibias.t72 commonsourceibias.t73 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X354 vdd.t41 vdd.t38 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X355 CSoutput.t173 commonsourceibias.t148 gnd.t234 gnd.t233 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 gnd.t232 commonsourceibias.t149 CSoutput.t172 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 vdd.t37 vdd.t34 vdd.t36 vdd.t35 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X358 a_n8300_8799.t10 plus.t21 a_n2903_n3924.t9 gnd.t2 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X359 a_n2903_n3924.t34 diffpairibias.t22 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X360 output.t1 CSoutput.t219 vdd.t8 gnd.t4 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X361 gnd.t230 commonsourceibias.t150 CSoutput.t171 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 vdd.t175 a_n8300_8799.t135 CSoutput.t40 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 vdd.t174 a_n8300_8799.t136 CSoutput.t3 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 gnd.t105 gnd.t102 gnd.t104 gnd.t103 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X365 gnd.t228 commonsourceibias.t151 CSoutput.t170 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 CSoutput.t45 a_n8300_8799.t137 vdd.t173 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 a_n2318_13878.t22 a_n2318_13878.t21 a_n2140_13878.t10 vdd.t22 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X368 commonsourceibias.t71 commonsourceibias.t70 gnd.t225 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X369 a_n8300_8799.t25 a_n2318_13878.t79 a_n2318_8322.t14 vdd.t123 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X370 gnd.t101 gnd.t98 gnd.t100 gnd.t99 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X371 gnd.t224 commonsourceibias.t152 CSoutput.t168 gnd.t223 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X372 vdd.t172 a_n8300_8799.t138 CSoutput.t68 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X373 CSoutput.t44 a_n8300_8799.t139 vdd.t171 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X374 a_n2903_n3924.t8 plus.t22 a_n8300_8799.t18 gnd.t54 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X375 vdd.t169 a_n8300_8799.t140 CSoutput.t191 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X376 diffpairibias.t3 diffpairibias.t2 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X377 vdd.t168 a_n8300_8799.t141 CSoutput.t56 vdd.t167 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X378 CSoutput.t78 a_n8300_8799.t142 vdd.t166 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X379 CSoutput.t55 a_n8300_8799.t143 vdd.t165 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X380 a_n2318_8322.t13 a_n2318_13878.t80 a_n8300_8799.t19 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X381 commonsourceibias.t69 commonsourceibias.t68 gnd.t222 gnd.t221 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X382 vdd.t163 a_n8300_8799.t144 CSoutput.t67 vdd.t162 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X383 gnd.t220 commonsourceibias.t153 CSoutput.t167 gnd.t219 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X384 CSoutput.t87 a_n8300_8799.t145 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X385 diffpairibias.t1 diffpairibias.t0 gnd.t20 gnd.t19 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X386 a_n8300_8799.t33 plus.t23 a_n2903_n3924.t7 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.5
X387 CSoutput.t220 a_n2318_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X388 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X389 CSoutput.t166 commonsourceibias.t154 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X390 gnd.t93 gnd.t90 gnd.t92 gnd.t91 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.5
X391 vdd.t33 vdd.t30 vdd.t32 vdd.t31 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X392 vdd.t116 a_n2318_13878.t81 a_n2140_13878.t0 vdd.t115 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X393 commonsourceibias.t67 commonsourceibias.t66 gnd.t216 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X394 gnd.t89 gnd.t86 gnd.t88 gnd.t87 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X395 CSoutput.t77 a_n8300_8799.t146 vdd.t159 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X396 gnd.t215 commonsourceibias.t155 CSoutput.t165 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X397 vdd.t29 vdd.t26 vdd.t28 vdd.t27 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X398 CSoutput.t164 commonsourceibias.t156 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X399 CSoutput.t178 commonsourceibias.t157 gnd.t193 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 vdd.t157 a_n8300_8799.t147 CSoutput.t196 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X401 commonsourceibias.t63 commonsourceibias.t62 gnd.t212 gnd.t211 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X402 vdd.t155 a_n8300_8799.t148 CSoutput.t31 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X403 CSoutput.t152 commonsourceibias.t158 gnd.t210 gnd.t209 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X404 CSoutput.t197 a_n8300_8799.t149 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X405 gnd.t208 commonsourceibias.t60 commonsourceibias.t61 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 vdd.t2 CSoutput.t221 output.t0 gnd.t3 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X407 a_n2318_13878.t2 minus.t23 a_n2903_n3924.t2 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X408 CSoutput.t151 commonsourceibias.t159 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X409 a_n2318_8322.t12 a_n2318_13878.t82 a_n8300_8799.t23 vdd.t127 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X410 gnd.t205 commonsourceibias.t58 commonsourceibias.t59 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X411 vdd.t151 a_n8300_8799.t150 CSoutput.t79 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X412 vdd.t149 a_n8300_8799.t151 CSoutput.t190 vdd.t148 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X413 vdd.t147 a_n8300_8799.t152 CSoutput.t84 vdd.t146 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X414 CSoutput.t199 a_n8300_8799.t153 vdd.t145 vdd.t144 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 commonsourceibias.t57 commonsourceibias.t56 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X416 gnd.t85 gnd.t83 plus.t0 gnd.t84 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X417 gnd.t201 commonsourceibias.t54 commonsourceibias.t55 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X418 a_n2903_n3924.t6 plus.t24 a_n8300_8799.t9 gnd.t53 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.5
X419 a_n2318_8322.t4 a_n2318_13878.t83 vdd.t129 vdd.t128 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X420 a_n2318_13878.t5 minus.t24 a_n2903_n3924.t5 gnd.t23 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.5
X421 a_n2140_13878.t9 a_n2318_13878.t39 a_n2318_13878.t40 vdd.t20 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X422 vdd.t143 a_n8300_8799.t154 CSoutput.t59 vdd.t142 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X423 commonsourceibias.t53 commonsourceibias.t52 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X424 a_n2903_n3924.t28 diffpairibias.t23 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X425 CSoutput.t49 a_n8300_8799.t155 vdd.t141 vdd.t140 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X426 gnd.t191 commonsourceibias.t78 commonsourceibias.t79 gnd.t190 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X427 a_n2318_13878.t20 a_n2318_13878.t19 a_n2140_13878.t8 vdd.t1 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
R0 commonsourceibias.n281 commonsourceibias.t102 222.032
R1 commonsourceibias.n44 commonsourceibias.t46 222.032
R2 commonsourceibias.n166 commonsourceibias.t119 222.032
R3 commonsourceibias.n643 commonsourceibias.t108 222.032
R4 commonsourceibias.n413 commonsourceibias.t36 222.032
R5 commonsourceibias.n529 commonsourceibias.t126 222.032
R6 commonsourceibias.n364 commonsourceibias.t101 207.983
R7 commonsourceibias.n127 commonsourceibias.t22 207.983
R8 commonsourceibias.n249 commonsourceibias.t117 207.983
R9 commonsourceibias.n731 commonsourceibias.t124 207.983
R10 commonsourceibias.n501 commonsourceibias.t52 207.983
R11 commonsourceibias.n616 commonsourceibias.t140 207.983
R12 commonsourceibias.n280 commonsourceibias.t152 168.701
R13 commonsourceibias.n286 commonsourceibias.t157 168.701
R14 commonsourceibias.n292 commonsourceibias.t112 168.701
R15 commonsourceibias.n276 commonsourceibias.t97 168.701
R16 commonsourceibias.n300 commonsourceibias.t85 168.701
R17 commonsourceibias.n306 commonsourceibias.t122 168.701
R18 commonsourceibias.n271 commonsourceibias.t104 168.701
R19 commonsourceibias.n314 commonsourceibias.t91 168.701
R20 commonsourceibias.n320 commonsourceibias.t94 168.701
R21 commonsourceibias.n266 commonsourceibias.t113 168.701
R22 commonsourceibias.n328 commonsourceibias.t96 168.701
R23 commonsourceibias.n334 commonsourceibias.t100 168.701
R24 commonsourceibias.n261 commonsourceibias.t151 168.701
R25 commonsourceibias.n342 commonsourceibias.t129 168.701
R26 commonsourceibias.n348 commonsourceibias.t109 168.701
R27 commonsourceibias.n256 commonsourceibias.t159 168.701
R28 commonsourceibias.n356 commonsourceibias.t81 168.701
R29 commonsourceibias.n362 commonsourceibias.t120 168.701
R30 commonsourceibias.n125 commonsourceibias.t74 168.701
R31 commonsourceibias.n119 commonsourceibias.t4 168.701
R32 commonsourceibias.n19 commonsourceibias.t20 168.701
R33 commonsourceibias.n111 commonsourceibias.t28 168.701
R34 commonsourceibias.n105 commonsourceibias.t40 168.701
R35 commonsourceibias.n24 commonsourceibias.t10 168.701
R36 commonsourceibias.n97 commonsourceibias.t16 168.701
R37 commonsourceibias.n91 commonsourceibias.t24 168.701
R38 commonsourceibias.n29 commonsourceibias.t68 168.701
R39 commonsourceibias.n83 commonsourceibias.t50 168.701
R40 commonsourceibias.n77 commonsourceibias.t12 168.701
R41 commonsourceibias.n34 commonsourceibias.t38 168.701
R42 commonsourceibias.n69 commonsourceibias.t42 168.701
R43 commonsourceibias.n63 commonsourceibias.t76 168.701
R44 commonsourceibias.n39 commonsourceibias.t0 168.701
R45 commonsourceibias.n55 commonsourceibias.t54 168.701
R46 commonsourceibias.n49 commonsourceibias.t66 168.701
R47 commonsourceibias.n43 commonsourceibias.t72 168.701
R48 commonsourceibias.n247 commonsourceibias.t135 168.701
R49 commonsourceibias.n241 commonsourceibias.t92 168.701
R50 commonsourceibias.n5 commonsourceibias.t90 168.701
R51 commonsourceibias.n233 commonsourceibias.t127 168.701
R52 commonsourceibias.n227 commonsourceibias.t145 168.701
R53 commonsourceibias.n10 commonsourceibias.t83 168.701
R54 commonsourceibias.n219 commonsourceibias.t116 168.701
R55 commonsourceibias.n213 commonsourceibias.t110 168.701
R56 commonsourceibias.n150 commonsourceibias.t131 168.701
R57 commonsourceibias.n151 commonsourceibias.t107 168.701
R58 commonsourceibias.n153 commonsourceibias.t103 168.701
R59 commonsourceibias.n155 commonsourceibias.t121 168.701
R60 commonsourceibias.n191 commonsourceibias.t138 168.701
R61 commonsourceibias.n185 commonsourceibias.t95 168.701
R62 commonsourceibias.n161 commonsourceibias.t111 168.701
R63 commonsourceibias.n177 commonsourceibias.t130 168.701
R64 commonsourceibias.n171 commonsourceibias.t87 168.701
R65 commonsourceibias.n165 commonsourceibias.t84 168.701
R66 commonsourceibias.n642 commonsourceibias.t158 168.701
R67 commonsourceibias.n648 commonsourceibias.t150 168.701
R68 commonsourceibias.n654 commonsourceibias.t136 168.701
R69 commonsourceibias.n656 commonsourceibias.t118 168.701
R70 commonsourceibias.n663 commonsourceibias.t99 168.701
R71 commonsourceibias.n669 commonsourceibias.t143 168.701
R72 commonsourceibias.n671 commonsourceibias.t128 168.701
R73 commonsourceibias.n678 commonsourceibias.t106 168.701
R74 commonsourceibias.n684 commonsourceibias.t88 168.701
R75 commonsourceibias.n686 commonsourceibias.t137 168.701
R76 commonsourceibias.n693 commonsourceibias.t115 168.701
R77 commonsourceibias.n699 commonsourceibias.t123 168.701
R78 commonsourceibias.n701 commonsourceibias.t144 168.701
R79 commonsourceibias.n708 commonsourceibias.t147 168.701
R80 commonsourceibias.n714 commonsourceibias.t132 168.701
R81 commonsourceibias.n716 commonsourceibias.t93 168.701
R82 commonsourceibias.n723 commonsourceibias.t154 168.701
R83 commonsourceibias.n729 commonsourceibias.t141 168.701
R84 commonsourceibias.n412 commonsourceibias.t14 168.701
R85 commonsourceibias.n418 commonsourceibias.t6 168.701
R86 commonsourceibias.n424 commonsourceibias.t34 168.701
R87 commonsourceibias.n426 commonsourceibias.t48 168.701
R88 commonsourceibias.n433 commonsourceibias.t64 168.701
R89 commonsourceibias.n439 commonsourceibias.t60 168.701
R90 commonsourceibias.n441 commonsourceibias.t2 168.701
R91 commonsourceibias.n448 commonsourceibias.t32 168.701
R92 commonsourceibias.n454 commonsourceibias.t62 168.701
R93 commonsourceibias.n456 commonsourceibias.t26 168.701
R94 commonsourceibias.n463 commonsourceibias.t56 168.701
R95 commonsourceibias.n469 commonsourceibias.t8 168.701
R96 commonsourceibias.n471 commonsourceibias.t70 168.701
R97 commonsourceibias.n478 commonsourceibias.t58 168.701
R98 commonsourceibias.n484 commonsourceibias.t18 168.701
R99 commonsourceibias.n486 commonsourceibias.t78 168.701
R100 commonsourceibias.n493 commonsourceibias.t44 168.701
R101 commonsourceibias.n499 commonsourceibias.t30 168.701
R102 commonsourceibias.n614 commonsourceibias.t153 168.701
R103 commonsourceibias.n608 commonsourceibias.t86 168.701
R104 commonsourceibias.n601 commonsourceibias.t105 168.701
R105 commonsourceibias.n599 commonsourceibias.t146 168.701
R106 commonsourceibias.n593 commonsourceibias.t80 168.701
R107 commonsourceibias.n586 commonsourceibias.t156 168.701
R108 commonsourceibias.n584 commonsourceibias.t139 168.701
R109 commonsourceibias.n578 commonsourceibias.t133 168.701
R110 commonsourceibias.n571 commonsourceibias.t149 168.701
R111 commonsourceibias.n528 commonsourceibias.t89 168.701
R112 commonsourceibias.n534 commonsourceibias.t82 168.701
R113 commonsourceibias.n540 commonsourceibias.t148 168.701
R114 commonsourceibias.n542 commonsourceibias.t134 168.701
R115 commonsourceibias.n549 commonsourceibias.t114 168.701
R116 commonsourceibias.n555 commonsourceibias.t155 168.701
R117 commonsourceibias.n519 commonsourceibias.t142 168.701
R118 commonsourceibias.n517 commonsourceibias.t125 168.701
R119 commonsourceibias.n515 commonsourceibias.t98 168.701
R120 commonsourceibias.n363 commonsourceibias.n251 161.3
R121 commonsourceibias.n361 commonsourceibias.n360 161.3
R122 commonsourceibias.n359 commonsourceibias.n252 161.3
R123 commonsourceibias.n358 commonsourceibias.n357 161.3
R124 commonsourceibias.n355 commonsourceibias.n253 161.3
R125 commonsourceibias.n354 commonsourceibias.n353 161.3
R126 commonsourceibias.n352 commonsourceibias.n254 161.3
R127 commonsourceibias.n351 commonsourceibias.n350 161.3
R128 commonsourceibias.n349 commonsourceibias.n255 161.3
R129 commonsourceibias.n347 commonsourceibias.n346 161.3
R130 commonsourceibias.n345 commonsourceibias.n257 161.3
R131 commonsourceibias.n344 commonsourceibias.n343 161.3
R132 commonsourceibias.n341 commonsourceibias.n258 161.3
R133 commonsourceibias.n340 commonsourceibias.n339 161.3
R134 commonsourceibias.n338 commonsourceibias.n259 161.3
R135 commonsourceibias.n337 commonsourceibias.n336 161.3
R136 commonsourceibias.n335 commonsourceibias.n260 161.3
R137 commonsourceibias.n333 commonsourceibias.n332 161.3
R138 commonsourceibias.n331 commonsourceibias.n262 161.3
R139 commonsourceibias.n330 commonsourceibias.n329 161.3
R140 commonsourceibias.n327 commonsourceibias.n263 161.3
R141 commonsourceibias.n326 commonsourceibias.n325 161.3
R142 commonsourceibias.n324 commonsourceibias.n264 161.3
R143 commonsourceibias.n323 commonsourceibias.n322 161.3
R144 commonsourceibias.n321 commonsourceibias.n265 161.3
R145 commonsourceibias.n319 commonsourceibias.n318 161.3
R146 commonsourceibias.n317 commonsourceibias.n267 161.3
R147 commonsourceibias.n316 commonsourceibias.n315 161.3
R148 commonsourceibias.n313 commonsourceibias.n268 161.3
R149 commonsourceibias.n312 commonsourceibias.n311 161.3
R150 commonsourceibias.n310 commonsourceibias.n269 161.3
R151 commonsourceibias.n309 commonsourceibias.n308 161.3
R152 commonsourceibias.n307 commonsourceibias.n270 161.3
R153 commonsourceibias.n305 commonsourceibias.n304 161.3
R154 commonsourceibias.n303 commonsourceibias.n272 161.3
R155 commonsourceibias.n302 commonsourceibias.n301 161.3
R156 commonsourceibias.n299 commonsourceibias.n273 161.3
R157 commonsourceibias.n298 commonsourceibias.n297 161.3
R158 commonsourceibias.n296 commonsourceibias.n274 161.3
R159 commonsourceibias.n295 commonsourceibias.n294 161.3
R160 commonsourceibias.n293 commonsourceibias.n275 161.3
R161 commonsourceibias.n291 commonsourceibias.n290 161.3
R162 commonsourceibias.n289 commonsourceibias.n277 161.3
R163 commonsourceibias.n288 commonsourceibias.n287 161.3
R164 commonsourceibias.n285 commonsourceibias.n278 161.3
R165 commonsourceibias.n284 commonsourceibias.n283 161.3
R166 commonsourceibias.n282 commonsourceibias.n279 161.3
R167 commonsourceibias.n45 commonsourceibias.n42 161.3
R168 commonsourceibias.n47 commonsourceibias.n46 161.3
R169 commonsourceibias.n48 commonsourceibias.n41 161.3
R170 commonsourceibias.n51 commonsourceibias.n50 161.3
R171 commonsourceibias.n52 commonsourceibias.n40 161.3
R172 commonsourceibias.n54 commonsourceibias.n53 161.3
R173 commonsourceibias.n56 commonsourceibias.n38 161.3
R174 commonsourceibias.n58 commonsourceibias.n57 161.3
R175 commonsourceibias.n59 commonsourceibias.n37 161.3
R176 commonsourceibias.n61 commonsourceibias.n60 161.3
R177 commonsourceibias.n62 commonsourceibias.n36 161.3
R178 commonsourceibias.n65 commonsourceibias.n64 161.3
R179 commonsourceibias.n66 commonsourceibias.n35 161.3
R180 commonsourceibias.n68 commonsourceibias.n67 161.3
R181 commonsourceibias.n70 commonsourceibias.n33 161.3
R182 commonsourceibias.n72 commonsourceibias.n71 161.3
R183 commonsourceibias.n73 commonsourceibias.n32 161.3
R184 commonsourceibias.n75 commonsourceibias.n74 161.3
R185 commonsourceibias.n76 commonsourceibias.n31 161.3
R186 commonsourceibias.n79 commonsourceibias.n78 161.3
R187 commonsourceibias.n80 commonsourceibias.n30 161.3
R188 commonsourceibias.n82 commonsourceibias.n81 161.3
R189 commonsourceibias.n84 commonsourceibias.n28 161.3
R190 commonsourceibias.n86 commonsourceibias.n85 161.3
R191 commonsourceibias.n87 commonsourceibias.n27 161.3
R192 commonsourceibias.n89 commonsourceibias.n88 161.3
R193 commonsourceibias.n90 commonsourceibias.n26 161.3
R194 commonsourceibias.n93 commonsourceibias.n92 161.3
R195 commonsourceibias.n94 commonsourceibias.n25 161.3
R196 commonsourceibias.n96 commonsourceibias.n95 161.3
R197 commonsourceibias.n98 commonsourceibias.n23 161.3
R198 commonsourceibias.n100 commonsourceibias.n99 161.3
R199 commonsourceibias.n101 commonsourceibias.n22 161.3
R200 commonsourceibias.n103 commonsourceibias.n102 161.3
R201 commonsourceibias.n104 commonsourceibias.n21 161.3
R202 commonsourceibias.n107 commonsourceibias.n106 161.3
R203 commonsourceibias.n108 commonsourceibias.n20 161.3
R204 commonsourceibias.n110 commonsourceibias.n109 161.3
R205 commonsourceibias.n112 commonsourceibias.n18 161.3
R206 commonsourceibias.n114 commonsourceibias.n113 161.3
R207 commonsourceibias.n115 commonsourceibias.n17 161.3
R208 commonsourceibias.n117 commonsourceibias.n116 161.3
R209 commonsourceibias.n118 commonsourceibias.n16 161.3
R210 commonsourceibias.n121 commonsourceibias.n120 161.3
R211 commonsourceibias.n122 commonsourceibias.n15 161.3
R212 commonsourceibias.n124 commonsourceibias.n123 161.3
R213 commonsourceibias.n126 commonsourceibias.n14 161.3
R214 commonsourceibias.n167 commonsourceibias.n164 161.3
R215 commonsourceibias.n169 commonsourceibias.n168 161.3
R216 commonsourceibias.n170 commonsourceibias.n163 161.3
R217 commonsourceibias.n173 commonsourceibias.n172 161.3
R218 commonsourceibias.n174 commonsourceibias.n162 161.3
R219 commonsourceibias.n176 commonsourceibias.n175 161.3
R220 commonsourceibias.n178 commonsourceibias.n160 161.3
R221 commonsourceibias.n180 commonsourceibias.n179 161.3
R222 commonsourceibias.n181 commonsourceibias.n159 161.3
R223 commonsourceibias.n183 commonsourceibias.n182 161.3
R224 commonsourceibias.n184 commonsourceibias.n158 161.3
R225 commonsourceibias.n187 commonsourceibias.n186 161.3
R226 commonsourceibias.n188 commonsourceibias.n157 161.3
R227 commonsourceibias.n190 commonsourceibias.n189 161.3
R228 commonsourceibias.n192 commonsourceibias.n156 161.3
R229 commonsourceibias.n194 commonsourceibias.n193 161.3
R230 commonsourceibias.n196 commonsourceibias.n195 161.3
R231 commonsourceibias.n197 commonsourceibias.n154 161.3
R232 commonsourceibias.n199 commonsourceibias.n198 161.3
R233 commonsourceibias.n201 commonsourceibias.n200 161.3
R234 commonsourceibias.n202 commonsourceibias.n152 161.3
R235 commonsourceibias.n204 commonsourceibias.n203 161.3
R236 commonsourceibias.n206 commonsourceibias.n205 161.3
R237 commonsourceibias.n208 commonsourceibias.n207 161.3
R238 commonsourceibias.n209 commonsourceibias.n13 161.3
R239 commonsourceibias.n211 commonsourceibias.n210 161.3
R240 commonsourceibias.n212 commonsourceibias.n12 161.3
R241 commonsourceibias.n215 commonsourceibias.n214 161.3
R242 commonsourceibias.n216 commonsourceibias.n11 161.3
R243 commonsourceibias.n218 commonsourceibias.n217 161.3
R244 commonsourceibias.n220 commonsourceibias.n9 161.3
R245 commonsourceibias.n222 commonsourceibias.n221 161.3
R246 commonsourceibias.n223 commonsourceibias.n8 161.3
R247 commonsourceibias.n225 commonsourceibias.n224 161.3
R248 commonsourceibias.n226 commonsourceibias.n7 161.3
R249 commonsourceibias.n229 commonsourceibias.n228 161.3
R250 commonsourceibias.n230 commonsourceibias.n6 161.3
R251 commonsourceibias.n232 commonsourceibias.n231 161.3
R252 commonsourceibias.n234 commonsourceibias.n4 161.3
R253 commonsourceibias.n236 commonsourceibias.n235 161.3
R254 commonsourceibias.n237 commonsourceibias.n3 161.3
R255 commonsourceibias.n239 commonsourceibias.n238 161.3
R256 commonsourceibias.n240 commonsourceibias.n2 161.3
R257 commonsourceibias.n243 commonsourceibias.n242 161.3
R258 commonsourceibias.n244 commonsourceibias.n1 161.3
R259 commonsourceibias.n246 commonsourceibias.n245 161.3
R260 commonsourceibias.n248 commonsourceibias.n0 161.3
R261 commonsourceibias.n730 commonsourceibias.n618 161.3
R262 commonsourceibias.n728 commonsourceibias.n727 161.3
R263 commonsourceibias.n726 commonsourceibias.n619 161.3
R264 commonsourceibias.n725 commonsourceibias.n724 161.3
R265 commonsourceibias.n722 commonsourceibias.n620 161.3
R266 commonsourceibias.n721 commonsourceibias.n720 161.3
R267 commonsourceibias.n719 commonsourceibias.n621 161.3
R268 commonsourceibias.n718 commonsourceibias.n717 161.3
R269 commonsourceibias.n715 commonsourceibias.n622 161.3
R270 commonsourceibias.n713 commonsourceibias.n712 161.3
R271 commonsourceibias.n711 commonsourceibias.n623 161.3
R272 commonsourceibias.n710 commonsourceibias.n709 161.3
R273 commonsourceibias.n707 commonsourceibias.n624 161.3
R274 commonsourceibias.n706 commonsourceibias.n705 161.3
R275 commonsourceibias.n704 commonsourceibias.n625 161.3
R276 commonsourceibias.n703 commonsourceibias.n702 161.3
R277 commonsourceibias.n700 commonsourceibias.n626 161.3
R278 commonsourceibias.n698 commonsourceibias.n697 161.3
R279 commonsourceibias.n696 commonsourceibias.n627 161.3
R280 commonsourceibias.n695 commonsourceibias.n694 161.3
R281 commonsourceibias.n692 commonsourceibias.n628 161.3
R282 commonsourceibias.n691 commonsourceibias.n690 161.3
R283 commonsourceibias.n689 commonsourceibias.n629 161.3
R284 commonsourceibias.n688 commonsourceibias.n687 161.3
R285 commonsourceibias.n685 commonsourceibias.n630 161.3
R286 commonsourceibias.n683 commonsourceibias.n682 161.3
R287 commonsourceibias.n681 commonsourceibias.n631 161.3
R288 commonsourceibias.n680 commonsourceibias.n679 161.3
R289 commonsourceibias.n677 commonsourceibias.n632 161.3
R290 commonsourceibias.n676 commonsourceibias.n675 161.3
R291 commonsourceibias.n674 commonsourceibias.n633 161.3
R292 commonsourceibias.n673 commonsourceibias.n672 161.3
R293 commonsourceibias.n670 commonsourceibias.n634 161.3
R294 commonsourceibias.n668 commonsourceibias.n667 161.3
R295 commonsourceibias.n666 commonsourceibias.n635 161.3
R296 commonsourceibias.n665 commonsourceibias.n664 161.3
R297 commonsourceibias.n662 commonsourceibias.n636 161.3
R298 commonsourceibias.n661 commonsourceibias.n660 161.3
R299 commonsourceibias.n659 commonsourceibias.n637 161.3
R300 commonsourceibias.n658 commonsourceibias.n657 161.3
R301 commonsourceibias.n655 commonsourceibias.n638 161.3
R302 commonsourceibias.n653 commonsourceibias.n652 161.3
R303 commonsourceibias.n651 commonsourceibias.n639 161.3
R304 commonsourceibias.n650 commonsourceibias.n649 161.3
R305 commonsourceibias.n647 commonsourceibias.n640 161.3
R306 commonsourceibias.n646 commonsourceibias.n645 161.3
R307 commonsourceibias.n644 commonsourceibias.n641 161.3
R308 commonsourceibias.n500 commonsourceibias.n388 161.3
R309 commonsourceibias.n498 commonsourceibias.n497 161.3
R310 commonsourceibias.n496 commonsourceibias.n389 161.3
R311 commonsourceibias.n495 commonsourceibias.n494 161.3
R312 commonsourceibias.n492 commonsourceibias.n390 161.3
R313 commonsourceibias.n491 commonsourceibias.n490 161.3
R314 commonsourceibias.n489 commonsourceibias.n391 161.3
R315 commonsourceibias.n488 commonsourceibias.n487 161.3
R316 commonsourceibias.n485 commonsourceibias.n392 161.3
R317 commonsourceibias.n483 commonsourceibias.n482 161.3
R318 commonsourceibias.n481 commonsourceibias.n393 161.3
R319 commonsourceibias.n480 commonsourceibias.n479 161.3
R320 commonsourceibias.n477 commonsourceibias.n394 161.3
R321 commonsourceibias.n476 commonsourceibias.n475 161.3
R322 commonsourceibias.n474 commonsourceibias.n395 161.3
R323 commonsourceibias.n473 commonsourceibias.n472 161.3
R324 commonsourceibias.n470 commonsourceibias.n396 161.3
R325 commonsourceibias.n468 commonsourceibias.n467 161.3
R326 commonsourceibias.n466 commonsourceibias.n397 161.3
R327 commonsourceibias.n465 commonsourceibias.n464 161.3
R328 commonsourceibias.n462 commonsourceibias.n398 161.3
R329 commonsourceibias.n461 commonsourceibias.n460 161.3
R330 commonsourceibias.n459 commonsourceibias.n399 161.3
R331 commonsourceibias.n458 commonsourceibias.n457 161.3
R332 commonsourceibias.n455 commonsourceibias.n400 161.3
R333 commonsourceibias.n453 commonsourceibias.n452 161.3
R334 commonsourceibias.n451 commonsourceibias.n401 161.3
R335 commonsourceibias.n450 commonsourceibias.n449 161.3
R336 commonsourceibias.n447 commonsourceibias.n402 161.3
R337 commonsourceibias.n446 commonsourceibias.n445 161.3
R338 commonsourceibias.n444 commonsourceibias.n403 161.3
R339 commonsourceibias.n443 commonsourceibias.n442 161.3
R340 commonsourceibias.n440 commonsourceibias.n404 161.3
R341 commonsourceibias.n438 commonsourceibias.n437 161.3
R342 commonsourceibias.n436 commonsourceibias.n405 161.3
R343 commonsourceibias.n435 commonsourceibias.n434 161.3
R344 commonsourceibias.n432 commonsourceibias.n406 161.3
R345 commonsourceibias.n431 commonsourceibias.n430 161.3
R346 commonsourceibias.n429 commonsourceibias.n407 161.3
R347 commonsourceibias.n428 commonsourceibias.n427 161.3
R348 commonsourceibias.n425 commonsourceibias.n408 161.3
R349 commonsourceibias.n423 commonsourceibias.n422 161.3
R350 commonsourceibias.n421 commonsourceibias.n409 161.3
R351 commonsourceibias.n420 commonsourceibias.n419 161.3
R352 commonsourceibias.n417 commonsourceibias.n410 161.3
R353 commonsourceibias.n416 commonsourceibias.n415 161.3
R354 commonsourceibias.n414 commonsourceibias.n411 161.3
R355 commonsourceibias.n570 commonsourceibias.n569 161.3
R356 commonsourceibias.n568 commonsourceibias.n567 161.3
R357 commonsourceibias.n566 commonsourceibias.n516 161.3
R358 commonsourceibias.n565 commonsourceibias.n564 161.3
R359 commonsourceibias.n563 commonsourceibias.n562 161.3
R360 commonsourceibias.n561 commonsourceibias.n518 161.3
R361 commonsourceibias.n560 commonsourceibias.n559 161.3
R362 commonsourceibias.n558 commonsourceibias.n557 161.3
R363 commonsourceibias.n556 commonsourceibias.n520 161.3
R364 commonsourceibias.n554 commonsourceibias.n553 161.3
R365 commonsourceibias.n552 commonsourceibias.n521 161.3
R366 commonsourceibias.n551 commonsourceibias.n550 161.3
R367 commonsourceibias.n548 commonsourceibias.n522 161.3
R368 commonsourceibias.n547 commonsourceibias.n546 161.3
R369 commonsourceibias.n545 commonsourceibias.n523 161.3
R370 commonsourceibias.n544 commonsourceibias.n543 161.3
R371 commonsourceibias.n541 commonsourceibias.n524 161.3
R372 commonsourceibias.n539 commonsourceibias.n538 161.3
R373 commonsourceibias.n537 commonsourceibias.n525 161.3
R374 commonsourceibias.n536 commonsourceibias.n535 161.3
R375 commonsourceibias.n533 commonsourceibias.n526 161.3
R376 commonsourceibias.n532 commonsourceibias.n531 161.3
R377 commonsourceibias.n530 commonsourceibias.n527 161.3
R378 commonsourceibias.n615 commonsourceibias.n367 161.3
R379 commonsourceibias.n613 commonsourceibias.n612 161.3
R380 commonsourceibias.n611 commonsourceibias.n368 161.3
R381 commonsourceibias.n610 commonsourceibias.n609 161.3
R382 commonsourceibias.n607 commonsourceibias.n369 161.3
R383 commonsourceibias.n606 commonsourceibias.n605 161.3
R384 commonsourceibias.n604 commonsourceibias.n370 161.3
R385 commonsourceibias.n603 commonsourceibias.n602 161.3
R386 commonsourceibias.n600 commonsourceibias.n371 161.3
R387 commonsourceibias.n598 commonsourceibias.n597 161.3
R388 commonsourceibias.n596 commonsourceibias.n372 161.3
R389 commonsourceibias.n595 commonsourceibias.n594 161.3
R390 commonsourceibias.n592 commonsourceibias.n373 161.3
R391 commonsourceibias.n591 commonsourceibias.n590 161.3
R392 commonsourceibias.n589 commonsourceibias.n374 161.3
R393 commonsourceibias.n588 commonsourceibias.n587 161.3
R394 commonsourceibias.n585 commonsourceibias.n375 161.3
R395 commonsourceibias.n583 commonsourceibias.n582 161.3
R396 commonsourceibias.n581 commonsourceibias.n376 161.3
R397 commonsourceibias.n580 commonsourceibias.n579 161.3
R398 commonsourceibias.n577 commonsourceibias.n377 161.3
R399 commonsourceibias.n576 commonsourceibias.n575 161.3
R400 commonsourceibias.n574 commonsourceibias.n378 161.3
R401 commonsourceibias.n573 commonsourceibias.n572 161.3
R402 commonsourceibias.n141 commonsourceibias.n139 81.5057
R403 commonsourceibias.n381 commonsourceibias.n379 81.5057
R404 commonsourceibias.n141 commonsourceibias.n140 80.9324
R405 commonsourceibias.n143 commonsourceibias.n142 80.9324
R406 commonsourceibias.n145 commonsourceibias.n144 80.9324
R407 commonsourceibias.n147 commonsourceibias.n146 80.9324
R408 commonsourceibias.n138 commonsourceibias.n137 80.9324
R409 commonsourceibias.n136 commonsourceibias.n135 80.9324
R410 commonsourceibias.n134 commonsourceibias.n133 80.9324
R411 commonsourceibias.n132 commonsourceibias.n131 80.9324
R412 commonsourceibias.n130 commonsourceibias.n129 80.9324
R413 commonsourceibias.n504 commonsourceibias.n503 80.9324
R414 commonsourceibias.n506 commonsourceibias.n505 80.9324
R415 commonsourceibias.n508 commonsourceibias.n507 80.9324
R416 commonsourceibias.n510 commonsourceibias.n509 80.9324
R417 commonsourceibias.n512 commonsourceibias.n511 80.9324
R418 commonsourceibias.n387 commonsourceibias.n386 80.9324
R419 commonsourceibias.n385 commonsourceibias.n384 80.9324
R420 commonsourceibias.n383 commonsourceibias.n382 80.9324
R421 commonsourceibias.n381 commonsourceibias.n380 80.9324
R422 commonsourceibias.n365 commonsourceibias.n364 80.6037
R423 commonsourceibias.n128 commonsourceibias.n127 80.6037
R424 commonsourceibias.n250 commonsourceibias.n249 80.6037
R425 commonsourceibias.n732 commonsourceibias.n731 80.6037
R426 commonsourceibias.n502 commonsourceibias.n501 80.6037
R427 commonsourceibias.n617 commonsourceibias.n616 80.6037
R428 commonsourceibias.n322 commonsourceibias.n321 56.5617
R429 commonsourceibias.n336 commonsourceibias.n335 56.5617
R430 commonsourceibias.n85 commonsourceibias.n84 56.5617
R431 commonsourceibias.n71 commonsourceibias.n70 56.5617
R432 commonsourceibias.n207 commonsourceibias.n206 56.5617
R433 commonsourceibias.n193 commonsourceibias.n192 56.5617
R434 commonsourceibias.n687 commonsourceibias.n685 56.5617
R435 commonsourceibias.n702 commonsourceibias.n700 56.5617
R436 commonsourceibias.n457 commonsourceibias.n455 56.5617
R437 commonsourceibias.n472 commonsourceibias.n470 56.5617
R438 commonsourceibias.n572 commonsourceibias.n570 56.5617
R439 commonsourceibias.n294 commonsourceibias.n293 56.5617
R440 commonsourceibias.n308 commonsourceibias.n307 56.5617
R441 commonsourceibias.n350 commonsourceibias.n349 56.5617
R442 commonsourceibias.n113 commonsourceibias.n112 56.5617
R443 commonsourceibias.n99 commonsourceibias.n98 56.5617
R444 commonsourceibias.n57 commonsourceibias.n56 56.5617
R445 commonsourceibias.n235 commonsourceibias.n234 56.5617
R446 commonsourceibias.n221 commonsourceibias.n220 56.5617
R447 commonsourceibias.n179 commonsourceibias.n178 56.5617
R448 commonsourceibias.n657 commonsourceibias.n655 56.5617
R449 commonsourceibias.n672 commonsourceibias.n670 56.5617
R450 commonsourceibias.n717 commonsourceibias.n715 56.5617
R451 commonsourceibias.n427 commonsourceibias.n425 56.5617
R452 commonsourceibias.n442 commonsourceibias.n440 56.5617
R453 commonsourceibias.n487 commonsourceibias.n485 56.5617
R454 commonsourceibias.n602 commonsourceibias.n600 56.5617
R455 commonsourceibias.n587 commonsourceibias.n585 56.5617
R456 commonsourceibias.n543 commonsourceibias.n541 56.5617
R457 commonsourceibias.n557 commonsourceibias.n556 56.5617
R458 commonsourceibias.n285 commonsourceibias.n284 51.2335
R459 commonsourceibias.n357 commonsourceibias.n252 51.2335
R460 commonsourceibias.n120 commonsourceibias.n15 51.2335
R461 commonsourceibias.n48 commonsourceibias.n47 51.2335
R462 commonsourceibias.n242 commonsourceibias.n1 51.2335
R463 commonsourceibias.n170 commonsourceibias.n169 51.2335
R464 commonsourceibias.n647 commonsourceibias.n646 51.2335
R465 commonsourceibias.n724 commonsourceibias.n619 51.2335
R466 commonsourceibias.n417 commonsourceibias.n416 51.2335
R467 commonsourceibias.n494 commonsourceibias.n389 51.2335
R468 commonsourceibias.n609 commonsourceibias.n368 51.2335
R469 commonsourceibias.n533 commonsourceibias.n532 51.2335
R470 commonsourceibias.n364 commonsourceibias.n363 50.9056
R471 commonsourceibias.n127 commonsourceibias.n126 50.9056
R472 commonsourceibias.n249 commonsourceibias.n248 50.9056
R473 commonsourceibias.n731 commonsourceibias.n730 50.9056
R474 commonsourceibias.n501 commonsourceibias.n500 50.9056
R475 commonsourceibias.n616 commonsourceibias.n615 50.9056
R476 commonsourceibias.n299 commonsourceibias.n298 50.2647
R477 commonsourceibias.n343 commonsourceibias.n257 50.2647
R478 commonsourceibias.n106 commonsourceibias.n20 50.2647
R479 commonsourceibias.n62 commonsourceibias.n61 50.2647
R480 commonsourceibias.n228 commonsourceibias.n6 50.2647
R481 commonsourceibias.n184 commonsourceibias.n183 50.2647
R482 commonsourceibias.n662 commonsourceibias.n661 50.2647
R483 commonsourceibias.n709 commonsourceibias.n623 50.2647
R484 commonsourceibias.n432 commonsourceibias.n431 50.2647
R485 commonsourceibias.n479 commonsourceibias.n393 50.2647
R486 commonsourceibias.n594 commonsourceibias.n372 50.2647
R487 commonsourceibias.n548 commonsourceibias.n547 50.2647
R488 commonsourceibias.n281 commonsourceibias.n280 49.9027
R489 commonsourceibias.n44 commonsourceibias.n43 49.9027
R490 commonsourceibias.n166 commonsourceibias.n165 49.9027
R491 commonsourceibias.n643 commonsourceibias.n642 49.9027
R492 commonsourceibias.n413 commonsourceibias.n412 49.9027
R493 commonsourceibias.n529 commonsourceibias.n528 49.9027
R494 commonsourceibias.n313 commonsourceibias.n312 49.296
R495 commonsourceibias.n329 commonsourceibias.n262 49.296
R496 commonsourceibias.n92 commonsourceibias.n25 49.296
R497 commonsourceibias.n76 commonsourceibias.n75 49.296
R498 commonsourceibias.n214 commonsourceibias.n11 49.296
R499 commonsourceibias.n198 commonsourceibias.n197 49.296
R500 commonsourceibias.n677 commonsourceibias.n676 49.296
R501 commonsourceibias.n694 commonsourceibias.n627 49.296
R502 commonsourceibias.n447 commonsourceibias.n446 49.296
R503 commonsourceibias.n464 commonsourceibias.n397 49.296
R504 commonsourceibias.n579 commonsourceibias.n376 49.296
R505 commonsourceibias.n562 commonsourceibias.n561 49.296
R506 commonsourceibias.n315 commonsourceibias.n267 48.3272
R507 commonsourceibias.n327 commonsourceibias.n326 48.3272
R508 commonsourceibias.n90 commonsourceibias.n89 48.3272
R509 commonsourceibias.n78 commonsourceibias.n30 48.3272
R510 commonsourceibias.n212 commonsourceibias.n211 48.3272
R511 commonsourceibias.n202 commonsourceibias.n201 48.3272
R512 commonsourceibias.n679 commonsourceibias.n631 48.3272
R513 commonsourceibias.n692 commonsourceibias.n691 48.3272
R514 commonsourceibias.n449 commonsourceibias.n401 48.3272
R515 commonsourceibias.n462 commonsourceibias.n461 48.3272
R516 commonsourceibias.n577 commonsourceibias.n576 48.3272
R517 commonsourceibias.n566 commonsourceibias.n565 48.3272
R518 commonsourceibias.n301 commonsourceibias.n272 47.3584
R519 commonsourceibias.n341 commonsourceibias.n340 47.3584
R520 commonsourceibias.n104 commonsourceibias.n103 47.3584
R521 commonsourceibias.n64 commonsourceibias.n35 47.3584
R522 commonsourceibias.n226 commonsourceibias.n225 47.3584
R523 commonsourceibias.n186 commonsourceibias.n157 47.3584
R524 commonsourceibias.n664 commonsourceibias.n635 47.3584
R525 commonsourceibias.n707 commonsourceibias.n706 47.3584
R526 commonsourceibias.n434 commonsourceibias.n405 47.3584
R527 commonsourceibias.n477 commonsourceibias.n476 47.3584
R528 commonsourceibias.n592 commonsourceibias.n591 47.3584
R529 commonsourceibias.n550 commonsourceibias.n521 47.3584
R530 commonsourceibias.n287 commonsourceibias.n277 46.3896
R531 commonsourceibias.n355 commonsourceibias.n354 46.3896
R532 commonsourceibias.n118 commonsourceibias.n117 46.3896
R533 commonsourceibias.n50 commonsourceibias.n40 46.3896
R534 commonsourceibias.n240 commonsourceibias.n239 46.3896
R535 commonsourceibias.n172 commonsourceibias.n162 46.3896
R536 commonsourceibias.n649 commonsourceibias.n639 46.3896
R537 commonsourceibias.n722 commonsourceibias.n721 46.3896
R538 commonsourceibias.n419 commonsourceibias.n409 46.3896
R539 commonsourceibias.n492 commonsourceibias.n491 46.3896
R540 commonsourceibias.n607 commonsourceibias.n606 46.3896
R541 commonsourceibias.n535 commonsourceibias.n525 46.3896
R542 commonsourceibias.n282 commonsourceibias.n281 44.7059
R543 commonsourceibias.n644 commonsourceibias.n643 44.7059
R544 commonsourceibias.n414 commonsourceibias.n413 44.7059
R545 commonsourceibias.n530 commonsourceibias.n529 44.7059
R546 commonsourceibias.n45 commonsourceibias.n44 44.7059
R547 commonsourceibias.n167 commonsourceibias.n166 44.7059
R548 commonsourceibias.n291 commonsourceibias.n277 34.7644
R549 commonsourceibias.n354 commonsourceibias.n254 34.7644
R550 commonsourceibias.n117 commonsourceibias.n17 34.7644
R551 commonsourceibias.n54 commonsourceibias.n40 34.7644
R552 commonsourceibias.n239 commonsourceibias.n3 34.7644
R553 commonsourceibias.n176 commonsourceibias.n162 34.7644
R554 commonsourceibias.n653 commonsourceibias.n639 34.7644
R555 commonsourceibias.n721 commonsourceibias.n621 34.7644
R556 commonsourceibias.n423 commonsourceibias.n409 34.7644
R557 commonsourceibias.n491 commonsourceibias.n391 34.7644
R558 commonsourceibias.n606 commonsourceibias.n370 34.7644
R559 commonsourceibias.n539 commonsourceibias.n525 34.7644
R560 commonsourceibias.n305 commonsourceibias.n272 33.7956
R561 commonsourceibias.n340 commonsourceibias.n259 33.7956
R562 commonsourceibias.n103 commonsourceibias.n22 33.7956
R563 commonsourceibias.n68 commonsourceibias.n35 33.7956
R564 commonsourceibias.n225 commonsourceibias.n8 33.7956
R565 commonsourceibias.n190 commonsourceibias.n157 33.7956
R566 commonsourceibias.n668 commonsourceibias.n635 33.7956
R567 commonsourceibias.n706 commonsourceibias.n625 33.7956
R568 commonsourceibias.n438 commonsourceibias.n405 33.7956
R569 commonsourceibias.n476 commonsourceibias.n395 33.7956
R570 commonsourceibias.n591 commonsourceibias.n374 33.7956
R571 commonsourceibias.n554 commonsourceibias.n521 33.7956
R572 commonsourceibias.n319 commonsourceibias.n267 32.8269
R573 commonsourceibias.n326 commonsourceibias.n264 32.8269
R574 commonsourceibias.n89 commonsourceibias.n27 32.8269
R575 commonsourceibias.n82 commonsourceibias.n30 32.8269
R576 commonsourceibias.n211 commonsourceibias.n13 32.8269
R577 commonsourceibias.n203 commonsourceibias.n202 32.8269
R578 commonsourceibias.n683 commonsourceibias.n631 32.8269
R579 commonsourceibias.n691 commonsourceibias.n629 32.8269
R580 commonsourceibias.n453 commonsourceibias.n401 32.8269
R581 commonsourceibias.n461 commonsourceibias.n399 32.8269
R582 commonsourceibias.n576 commonsourceibias.n378 32.8269
R583 commonsourceibias.n567 commonsourceibias.n566 32.8269
R584 commonsourceibias.n312 commonsourceibias.n269 31.8581
R585 commonsourceibias.n333 commonsourceibias.n262 31.8581
R586 commonsourceibias.n96 commonsourceibias.n25 31.8581
R587 commonsourceibias.n75 commonsourceibias.n32 31.8581
R588 commonsourceibias.n218 commonsourceibias.n11 31.8581
R589 commonsourceibias.n197 commonsourceibias.n196 31.8581
R590 commonsourceibias.n676 commonsourceibias.n633 31.8581
R591 commonsourceibias.n698 commonsourceibias.n627 31.8581
R592 commonsourceibias.n446 commonsourceibias.n403 31.8581
R593 commonsourceibias.n468 commonsourceibias.n397 31.8581
R594 commonsourceibias.n583 commonsourceibias.n376 31.8581
R595 commonsourceibias.n561 commonsourceibias.n560 31.8581
R596 commonsourceibias.n298 commonsourceibias.n274 30.8893
R597 commonsourceibias.n347 commonsourceibias.n257 30.8893
R598 commonsourceibias.n110 commonsourceibias.n20 30.8893
R599 commonsourceibias.n61 commonsourceibias.n37 30.8893
R600 commonsourceibias.n232 commonsourceibias.n6 30.8893
R601 commonsourceibias.n183 commonsourceibias.n159 30.8893
R602 commonsourceibias.n661 commonsourceibias.n637 30.8893
R603 commonsourceibias.n713 commonsourceibias.n623 30.8893
R604 commonsourceibias.n431 commonsourceibias.n407 30.8893
R605 commonsourceibias.n483 commonsourceibias.n393 30.8893
R606 commonsourceibias.n598 commonsourceibias.n372 30.8893
R607 commonsourceibias.n547 commonsourceibias.n523 30.8893
R608 commonsourceibias.n284 commonsourceibias.n279 29.9206
R609 commonsourceibias.n361 commonsourceibias.n252 29.9206
R610 commonsourceibias.n124 commonsourceibias.n15 29.9206
R611 commonsourceibias.n47 commonsourceibias.n42 29.9206
R612 commonsourceibias.n246 commonsourceibias.n1 29.9206
R613 commonsourceibias.n169 commonsourceibias.n164 29.9206
R614 commonsourceibias.n646 commonsourceibias.n641 29.9206
R615 commonsourceibias.n728 commonsourceibias.n619 29.9206
R616 commonsourceibias.n416 commonsourceibias.n411 29.9206
R617 commonsourceibias.n498 commonsourceibias.n389 29.9206
R618 commonsourceibias.n613 commonsourceibias.n368 29.9206
R619 commonsourceibias.n532 commonsourceibias.n527 29.9206
R620 commonsourceibias.n363 commonsourceibias.n362 21.8872
R621 commonsourceibias.n126 commonsourceibias.n125 21.8872
R622 commonsourceibias.n248 commonsourceibias.n247 21.8872
R623 commonsourceibias.n730 commonsourceibias.n729 21.8872
R624 commonsourceibias.n500 commonsourceibias.n499 21.8872
R625 commonsourceibias.n615 commonsourceibias.n614 21.8872
R626 commonsourceibias.n294 commonsourceibias.n276 21.3954
R627 commonsourceibias.n349 commonsourceibias.n348 21.3954
R628 commonsourceibias.n112 commonsourceibias.n111 21.3954
R629 commonsourceibias.n57 commonsourceibias.n39 21.3954
R630 commonsourceibias.n234 commonsourceibias.n233 21.3954
R631 commonsourceibias.n179 commonsourceibias.n161 21.3954
R632 commonsourceibias.n657 commonsourceibias.n656 21.3954
R633 commonsourceibias.n715 commonsourceibias.n714 21.3954
R634 commonsourceibias.n427 commonsourceibias.n426 21.3954
R635 commonsourceibias.n485 commonsourceibias.n484 21.3954
R636 commonsourceibias.n600 commonsourceibias.n599 21.3954
R637 commonsourceibias.n543 commonsourceibias.n542 21.3954
R638 commonsourceibias.n308 commonsourceibias.n271 20.9036
R639 commonsourceibias.n335 commonsourceibias.n334 20.9036
R640 commonsourceibias.n98 commonsourceibias.n97 20.9036
R641 commonsourceibias.n71 commonsourceibias.n34 20.9036
R642 commonsourceibias.n220 commonsourceibias.n219 20.9036
R643 commonsourceibias.n193 commonsourceibias.n155 20.9036
R644 commonsourceibias.n672 commonsourceibias.n671 20.9036
R645 commonsourceibias.n700 commonsourceibias.n699 20.9036
R646 commonsourceibias.n442 commonsourceibias.n441 20.9036
R647 commonsourceibias.n470 commonsourceibias.n469 20.9036
R648 commonsourceibias.n585 commonsourceibias.n584 20.9036
R649 commonsourceibias.n557 commonsourceibias.n519 20.9036
R650 commonsourceibias.n321 commonsourceibias.n320 20.4117
R651 commonsourceibias.n322 commonsourceibias.n266 20.4117
R652 commonsourceibias.n85 commonsourceibias.n29 20.4117
R653 commonsourceibias.n84 commonsourceibias.n83 20.4117
R654 commonsourceibias.n207 commonsourceibias.n150 20.4117
R655 commonsourceibias.n206 commonsourceibias.n151 20.4117
R656 commonsourceibias.n685 commonsourceibias.n684 20.4117
R657 commonsourceibias.n687 commonsourceibias.n686 20.4117
R658 commonsourceibias.n455 commonsourceibias.n454 20.4117
R659 commonsourceibias.n457 commonsourceibias.n456 20.4117
R660 commonsourceibias.n572 commonsourceibias.n571 20.4117
R661 commonsourceibias.n570 commonsourceibias.n515 20.4117
R662 commonsourceibias.n307 commonsourceibias.n306 19.9199
R663 commonsourceibias.n336 commonsourceibias.n261 19.9199
R664 commonsourceibias.n99 commonsourceibias.n24 19.9199
R665 commonsourceibias.n70 commonsourceibias.n69 19.9199
R666 commonsourceibias.n221 commonsourceibias.n10 19.9199
R667 commonsourceibias.n192 commonsourceibias.n191 19.9199
R668 commonsourceibias.n670 commonsourceibias.n669 19.9199
R669 commonsourceibias.n702 commonsourceibias.n701 19.9199
R670 commonsourceibias.n440 commonsourceibias.n439 19.9199
R671 commonsourceibias.n472 commonsourceibias.n471 19.9199
R672 commonsourceibias.n587 commonsourceibias.n586 19.9199
R673 commonsourceibias.n556 commonsourceibias.n555 19.9199
R674 commonsourceibias.n293 commonsourceibias.n292 19.4281
R675 commonsourceibias.n350 commonsourceibias.n256 19.4281
R676 commonsourceibias.n113 commonsourceibias.n19 19.4281
R677 commonsourceibias.n56 commonsourceibias.n55 19.4281
R678 commonsourceibias.n235 commonsourceibias.n5 19.4281
R679 commonsourceibias.n178 commonsourceibias.n177 19.4281
R680 commonsourceibias.n655 commonsourceibias.n654 19.4281
R681 commonsourceibias.n717 commonsourceibias.n716 19.4281
R682 commonsourceibias.n425 commonsourceibias.n424 19.4281
R683 commonsourceibias.n487 commonsourceibias.n486 19.4281
R684 commonsourceibias.n602 commonsourceibias.n601 19.4281
R685 commonsourceibias.n541 commonsourceibias.n540 19.4281
R686 commonsourceibias.n286 commonsourceibias.n285 13.526
R687 commonsourceibias.n357 commonsourceibias.n356 13.526
R688 commonsourceibias.n120 commonsourceibias.n119 13.526
R689 commonsourceibias.n49 commonsourceibias.n48 13.526
R690 commonsourceibias.n242 commonsourceibias.n241 13.526
R691 commonsourceibias.n171 commonsourceibias.n170 13.526
R692 commonsourceibias.n648 commonsourceibias.n647 13.526
R693 commonsourceibias.n724 commonsourceibias.n723 13.526
R694 commonsourceibias.n418 commonsourceibias.n417 13.526
R695 commonsourceibias.n494 commonsourceibias.n493 13.526
R696 commonsourceibias.n609 commonsourceibias.n608 13.526
R697 commonsourceibias.n534 commonsourceibias.n533 13.526
R698 commonsourceibias.n130 commonsourceibias.n128 13.2322
R699 commonsourceibias.n504 commonsourceibias.n502 13.2322
R700 commonsourceibias.n300 commonsourceibias.n299 13.0342
R701 commonsourceibias.n343 commonsourceibias.n342 13.0342
R702 commonsourceibias.n106 commonsourceibias.n105 13.0342
R703 commonsourceibias.n63 commonsourceibias.n62 13.0342
R704 commonsourceibias.n228 commonsourceibias.n227 13.0342
R705 commonsourceibias.n185 commonsourceibias.n184 13.0342
R706 commonsourceibias.n663 commonsourceibias.n662 13.0342
R707 commonsourceibias.n709 commonsourceibias.n708 13.0342
R708 commonsourceibias.n433 commonsourceibias.n432 13.0342
R709 commonsourceibias.n479 commonsourceibias.n478 13.0342
R710 commonsourceibias.n594 commonsourceibias.n593 13.0342
R711 commonsourceibias.n549 commonsourceibias.n548 13.0342
R712 commonsourceibias.n314 commonsourceibias.n313 12.5423
R713 commonsourceibias.n329 commonsourceibias.n328 12.5423
R714 commonsourceibias.n92 commonsourceibias.n91 12.5423
R715 commonsourceibias.n77 commonsourceibias.n76 12.5423
R716 commonsourceibias.n214 commonsourceibias.n213 12.5423
R717 commonsourceibias.n198 commonsourceibias.n153 12.5423
R718 commonsourceibias.n678 commonsourceibias.n677 12.5423
R719 commonsourceibias.n694 commonsourceibias.n693 12.5423
R720 commonsourceibias.n448 commonsourceibias.n447 12.5423
R721 commonsourceibias.n464 commonsourceibias.n463 12.5423
R722 commonsourceibias.n579 commonsourceibias.n578 12.5423
R723 commonsourceibias.n562 commonsourceibias.n517 12.5423
R724 commonsourceibias.n315 commonsourceibias.n314 12.0505
R725 commonsourceibias.n328 commonsourceibias.n327 12.0505
R726 commonsourceibias.n91 commonsourceibias.n90 12.0505
R727 commonsourceibias.n78 commonsourceibias.n77 12.0505
R728 commonsourceibias.n213 commonsourceibias.n212 12.0505
R729 commonsourceibias.n201 commonsourceibias.n153 12.0505
R730 commonsourceibias.n679 commonsourceibias.n678 12.0505
R731 commonsourceibias.n693 commonsourceibias.n692 12.0505
R732 commonsourceibias.n449 commonsourceibias.n448 12.0505
R733 commonsourceibias.n463 commonsourceibias.n462 12.0505
R734 commonsourceibias.n578 commonsourceibias.n577 12.0505
R735 commonsourceibias.n565 commonsourceibias.n517 12.0505
R736 commonsourceibias.n734 commonsourceibias.n366 11.9876
R737 commonsourceibias.n301 commonsourceibias.n300 11.5587
R738 commonsourceibias.n342 commonsourceibias.n341 11.5587
R739 commonsourceibias.n105 commonsourceibias.n104 11.5587
R740 commonsourceibias.n64 commonsourceibias.n63 11.5587
R741 commonsourceibias.n227 commonsourceibias.n226 11.5587
R742 commonsourceibias.n186 commonsourceibias.n185 11.5587
R743 commonsourceibias.n664 commonsourceibias.n663 11.5587
R744 commonsourceibias.n708 commonsourceibias.n707 11.5587
R745 commonsourceibias.n434 commonsourceibias.n433 11.5587
R746 commonsourceibias.n478 commonsourceibias.n477 11.5587
R747 commonsourceibias.n593 commonsourceibias.n592 11.5587
R748 commonsourceibias.n550 commonsourceibias.n549 11.5587
R749 commonsourceibias.n287 commonsourceibias.n286 11.0668
R750 commonsourceibias.n356 commonsourceibias.n355 11.0668
R751 commonsourceibias.n119 commonsourceibias.n118 11.0668
R752 commonsourceibias.n50 commonsourceibias.n49 11.0668
R753 commonsourceibias.n241 commonsourceibias.n240 11.0668
R754 commonsourceibias.n172 commonsourceibias.n171 11.0668
R755 commonsourceibias.n649 commonsourceibias.n648 11.0668
R756 commonsourceibias.n723 commonsourceibias.n722 11.0668
R757 commonsourceibias.n419 commonsourceibias.n418 11.0668
R758 commonsourceibias.n493 commonsourceibias.n492 11.0668
R759 commonsourceibias.n608 commonsourceibias.n607 11.0668
R760 commonsourceibias.n535 commonsourceibias.n534 11.0668
R761 commonsourceibias.n734 commonsourceibias.n733 10.3347
R762 commonsourceibias.n149 commonsourceibias.n148 9.50363
R763 commonsourceibias.n514 commonsourceibias.n513 9.50363
R764 commonsourceibias.n366 commonsourceibias.n250 8.75852
R765 commonsourceibias.n733 commonsourceibias.n617 8.75852
R766 commonsourceibias.n292 commonsourceibias.n291 5.16479
R767 commonsourceibias.n256 commonsourceibias.n254 5.16479
R768 commonsourceibias.n19 commonsourceibias.n17 5.16479
R769 commonsourceibias.n55 commonsourceibias.n54 5.16479
R770 commonsourceibias.n5 commonsourceibias.n3 5.16479
R771 commonsourceibias.n177 commonsourceibias.n176 5.16479
R772 commonsourceibias.n654 commonsourceibias.n653 5.16479
R773 commonsourceibias.n716 commonsourceibias.n621 5.16479
R774 commonsourceibias.n424 commonsourceibias.n423 5.16479
R775 commonsourceibias.n486 commonsourceibias.n391 5.16479
R776 commonsourceibias.n601 commonsourceibias.n370 5.16479
R777 commonsourceibias.n540 commonsourceibias.n539 5.16479
R778 commonsourceibias.n366 commonsourceibias.n365 5.03125
R779 commonsourceibias.n733 commonsourceibias.n732 5.03125
R780 commonsourceibias.n306 commonsourceibias.n305 4.67295
R781 commonsourceibias.n261 commonsourceibias.n259 4.67295
R782 commonsourceibias.n24 commonsourceibias.n22 4.67295
R783 commonsourceibias.n69 commonsourceibias.n68 4.67295
R784 commonsourceibias.n10 commonsourceibias.n8 4.67295
R785 commonsourceibias.n191 commonsourceibias.n190 4.67295
R786 commonsourceibias.n669 commonsourceibias.n668 4.67295
R787 commonsourceibias.n701 commonsourceibias.n625 4.67295
R788 commonsourceibias.n439 commonsourceibias.n438 4.67295
R789 commonsourceibias.n471 commonsourceibias.n395 4.67295
R790 commonsourceibias.n586 commonsourceibias.n374 4.67295
R791 commonsourceibias.n555 commonsourceibias.n554 4.67295
R792 commonsourceibias commonsourceibias.n734 4.20978
R793 commonsourceibias.n320 commonsourceibias.n319 4.18111
R794 commonsourceibias.n266 commonsourceibias.n264 4.18111
R795 commonsourceibias.n29 commonsourceibias.n27 4.18111
R796 commonsourceibias.n83 commonsourceibias.n82 4.18111
R797 commonsourceibias.n150 commonsourceibias.n13 4.18111
R798 commonsourceibias.n203 commonsourceibias.n151 4.18111
R799 commonsourceibias.n684 commonsourceibias.n683 4.18111
R800 commonsourceibias.n686 commonsourceibias.n629 4.18111
R801 commonsourceibias.n454 commonsourceibias.n453 4.18111
R802 commonsourceibias.n456 commonsourceibias.n399 4.18111
R803 commonsourceibias.n571 commonsourceibias.n378 4.18111
R804 commonsourceibias.n567 commonsourceibias.n515 4.18111
R805 commonsourceibias.n271 commonsourceibias.n269 3.68928
R806 commonsourceibias.n334 commonsourceibias.n333 3.68928
R807 commonsourceibias.n97 commonsourceibias.n96 3.68928
R808 commonsourceibias.n34 commonsourceibias.n32 3.68928
R809 commonsourceibias.n219 commonsourceibias.n218 3.68928
R810 commonsourceibias.n196 commonsourceibias.n155 3.68928
R811 commonsourceibias.n671 commonsourceibias.n633 3.68928
R812 commonsourceibias.n699 commonsourceibias.n698 3.68928
R813 commonsourceibias.n441 commonsourceibias.n403 3.68928
R814 commonsourceibias.n469 commonsourceibias.n468 3.68928
R815 commonsourceibias.n584 commonsourceibias.n583 3.68928
R816 commonsourceibias.n560 commonsourceibias.n519 3.68928
R817 commonsourceibias.n276 commonsourceibias.n274 3.19744
R818 commonsourceibias.n348 commonsourceibias.n347 3.19744
R819 commonsourceibias.n111 commonsourceibias.n110 3.19744
R820 commonsourceibias.n39 commonsourceibias.n37 3.19744
R821 commonsourceibias.n233 commonsourceibias.n232 3.19744
R822 commonsourceibias.n161 commonsourceibias.n159 3.19744
R823 commonsourceibias.n656 commonsourceibias.n637 3.19744
R824 commonsourceibias.n714 commonsourceibias.n713 3.19744
R825 commonsourceibias.n426 commonsourceibias.n407 3.19744
R826 commonsourceibias.n484 commonsourceibias.n483 3.19744
R827 commonsourceibias.n599 commonsourceibias.n598 3.19744
R828 commonsourceibias.n542 commonsourceibias.n523 3.19744
R829 commonsourceibias.n139 commonsourceibias.t73 2.82907
R830 commonsourceibias.n139 commonsourceibias.t47 2.82907
R831 commonsourceibias.n140 commonsourceibias.t55 2.82907
R832 commonsourceibias.n140 commonsourceibias.t67 2.82907
R833 commonsourceibias.n142 commonsourceibias.t77 2.82907
R834 commonsourceibias.n142 commonsourceibias.t1 2.82907
R835 commonsourceibias.n144 commonsourceibias.t39 2.82907
R836 commonsourceibias.n144 commonsourceibias.t43 2.82907
R837 commonsourceibias.n146 commonsourceibias.t51 2.82907
R838 commonsourceibias.n146 commonsourceibias.t13 2.82907
R839 commonsourceibias.n137 commonsourceibias.t25 2.82907
R840 commonsourceibias.n137 commonsourceibias.t69 2.82907
R841 commonsourceibias.n135 commonsourceibias.t11 2.82907
R842 commonsourceibias.n135 commonsourceibias.t17 2.82907
R843 commonsourceibias.n133 commonsourceibias.t29 2.82907
R844 commonsourceibias.n133 commonsourceibias.t41 2.82907
R845 commonsourceibias.n131 commonsourceibias.t5 2.82907
R846 commonsourceibias.n131 commonsourceibias.t21 2.82907
R847 commonsourceibias.n129 commonsourceibias.t23 2.82907
R848 commonsourceibias.n129 commonsourceibias.t75 2.82907
R849 commonsourceibias.n503 commonsourceibias.t31 2.82907
R850 commonsourceibias.n503 commonsourceibias.t53 2.82907
R851 commonsourceibias.n505 commonsourceibias.t79 2.82907
R852 commonsourceibias.n505 commonsourceibias.t45 2.82907
R853 commonsourceibias.n507 commonsourceibias.t59 2.82907
R854 commonsourceibias.n507 commonsourceibias.t19 2.82907
R855 commonsourceibias.n509 commonsourceibias.t9 2.82907
R856 commonsourceibias.n509 commonsourceibias.t71 2.82907
R857 commonsourceibias.n511 commonsourceibias.t27 2.82907
R858 commonsourceibias.n511 commonsourceibias.t57 2.82907
R859 commonsourceibias.n386 commonsourceibias.t33 2.82907
R860 commonsourceibias.n386 commonsourceibias.t63 2.82907
R861 commonsourceibias.n384 commonsourceibias.t61 2.82907
R862 commonsourceibias.n384 commonsourceibias.t3 2.82907
R863 commonsourceibias.n382 commonsourceibias.t49 2.82907
R864 commonsourceibias.n382 commonsourceibias.t65 2.82907
R865 commonsourceibias.n380 commonsourceibias.t7 2.82907
R866 commonsourceibias.n380 commonsourceibias.t35 2.82907
R867 commonsourceibias.n379 commonsourceibias.t37 2.82907
R868 commonsourceibias.n379 commonsourceibias.t15 2.82907
R869 commonsourceibias.n280 commonsourceibias.n279 2.7056
R870 commonsourceibias.n362 commonsourceibias.n361 2.7056
R871 commonsourceibias.n125 commonsourceibias.n124 2.7056
R872 commonsourceibias.n43 commonsourceibias.n42 2.7056
R873 commonsourceibias.n247 commonsourceibias.n246 2.7056
R874 commonsourceibias.n165 commonsourceibias.n164 2.7056
R875 commonsourceibias.n642 commonsourceibias.n641 2.7056
R876 commonsourceibias.n729 commonsourceibias.n728 2.7056
R877 commonsourceibias.n412 commonsourceibias.n411 2.7056
R878 commonsourceibias.n499 commonsourceibias.n498 2.7056
R879 commonsourceibias.n614 commonsourceibias.n613 2.7056
R880 commonsourceibias.n528 commonsourceibias.n527 2.7056
R881 commonsourceibias.n132 commonsourceibias.n130 0.573776
R882 commonsourceibias.n134 commonsourceibias.n132 0.573776
R883 commonsourceibias.n136 commonsourceibias.n134 0.573776
R884 commonsourceibias.n138 commonsourceibias.n136 0.573776
R885 commonsourceibias.n147 commonsourceibias.n145 0.573776
R886 commonsourceibias.n145 commonsourceibias.n143 0.573776
R887 commonsourceibias.n143 commonsourceibias.n141 0.573776
R888 commonsourceibias.n383 commonsourceibias.n381 0.573776
R889 commonsourceibias.n385 commonsourceibias.n383 0.573776
R890 commonsourceibias.n387 commonsourceibias.n385 0.573776
R891 commonsourceibias.n512 commonsourceibias.n510 0.573776
R892 commonsourceibias.n510 commonsourceibias.n508 0.573776
R893 commonsourceibias.n508 commonsourceibias.n506 0.573776
R894 commonsourceibias.n506 commonsourceibias.n504 0.573776
R895 commonsourceibias.n148 commonsourceibias.n138 0.287138
R896 commonsourceibias.n148 commonsourceibias.n147 0.287138
R897 commonsourceibias.n513 commonsourceibias.n387 0.287138
R898 commonsourceibias.n513 commonsourceibias.n512 0.287138
R899 commonsourceibias.n365 commonsourceibias.n251 0.285035
R900 commonsourceibias.n128 commonsourceibias.n14 0.285035
R901 commonsourceibias.n250 commonsourceibias.n0 0.285035
R902 commonsourceibias.n732 commonsourceibias.n618 0.285035
R903 commonsourceibias.n502 commonsourceibias.n388 0.285035
R904 commonsourceibias.n617 commonsourceibias.n367 0.285035
R905 commonsourceibias.n360 commonsourceibias.n251 0.189894
R906 commonsourceibias.n360 commonsourceibias.n359 0.189894
R907 commonsourceibias.n359 commonsourceibias.n358 0.189894
R908 commonsourceibias.n358 commonsourceibias.n253 0.189894
R909 commonsourceibias.n353 commonsourceibias.n253 0.189894
R910 commonsourceibias.n353 commonsourceibias.n352 0.189894
R911 commonsourceibias.n352 commonsourceibias.n351 0.189894
R912 commonsourceibias.n351 commonsourceibias.n255 0.189894
R913 commonsourceibias.n346 commonsourceibias.n255 0.189894
R914 commonsourceibias.n346 commonsourceibias.n345 0.189894
R915 commonsourceibias.n345 commonsourceibias.n344 0.189894
R916 commonsourceibias.n344 commonsourceibias.n258 0.189894
R917 commonsourceibias.n339 commonsourceibias.n258 0.189894
R918 commonsourceibias.n339 commonsourceibias.n338 0.189894
R919 commonsourceibias.n338 commonsourceibias.n337 0.189894
R920 commonsourceibias.n337 commonsourceibias.n260 0.189894
R921 commonsourceibias.n332 commonsourceibias.n260 0.189894
R922 commonsourceibias.n332 commonsourceibias.n331 0.189894
R923 commonsourceibias.n331 commonsourceibias.n330 0.189894
R924 commonsourceibias.n330 commonsourceibias.n263 0.189894
R925 commonsourceibias.n325 commonsourceibias.n263 0.189894
R926 commonsourceibias.n325 commonsourceibias.n324 0.189894
R927 commonsourceibias.n324 commonsourceibias.n323 0.189894
R928 commonsourceibias.n323 commonsourceibias.n265 0.189894
R929 commonsourceibias.n318 commonsourceibias.n265 0.189894
R930 commonsourceibias.n318 commonsourceibias.n317 0.189894
R931 commonsourceibias.n317 commonsourceibias.n316 0.189894
R932 commonsourceibias.n316 commonsourceibias.n268 0.189894
R933 commonsourceibias.n311 commonsourceibias.n268 0.189894
R934 commonsourceibias.n311 commonsourceibias.n310 0.189894
R935 commonsourceibias.n310 commonsourceibias.n309 0.189894
R936 commonsourceibias.n309 commonsourceibias.n270 0.189894
R937 commonsourceibias.n304 commonsourceibias.n270 0.189894
R938 commonsourceibias.n304 commonsourceibias.n303 0.189894
R939 commonsourceibias.n303 commonsourceibias.n302 0.189894
R940 commonsourceibias.n302 commonsourceibias.n273 0.189894
R941 commonsourceibias.n297 commonsourceibias.n273 0.189894
R942 commonsourceibias.n297 commonsourceibias.n296 0.189894
R943 commonsourceibias.n296 commonsourceibias.n295 0.189894
R944 commonsourceibias.n295 commonsourceibias.n275 0.189894
R945 commonsourceibias.n290 commonsourceibias.n275 0.189894
R946 commonsourceibias.n290 commonsourceibias.n289 0.189894
R947 commonsourceibias.n289 commonsourceibias.n288 0.189894
R948 commonsourceibias.n288 commonsourceibias.n278 0.189894
R949 commonsourceibias.n283 commonsourceibias.n278 0.189894
R950 commonsourceibias.n283 commonsourceibias.n282 0.189894
R951 commonsourceibias.n123 commonsourceibias.n14 0.189894
R952 commonsourceibias.n123 commonsourceibias.n122 0.189894
R953 commonsourceibias.n122 commonsourceibias.n121 0.189894
R954 commonsourceibias.n121 commonsourceibias.n16 0.189894
R955 commonsourceibias.n116 commonsourceibias.n16 0.189894
R956 commonsourceibias.n116 commonsourceibias.n115 0.189894
R957 commonsourceibias.n115 commonsourceibias.n114 0.189894
R958 commonsourceibias.n114 commonsourceibias.n18 0.189894
R959 commonsourceibias.n109 commonsourceibias.n18 0.189894
R960 commonsourceibias.n109 commonsourceibias.n108 0.189894
R961 commonsourceibias.n108 commonsourceibias.n107 0.189894
R962 commonsourceibias.n107 commonsourceibias.n21 0.189894
R963 commonsourceibias.n102 commonsourceibias.n21 0.189894
R964 commonsourceibias.n102 commonsourceibias.n101 0.189894
R965 commonsourceibias.n101 commonsourceibias.n100 0.189894
R966 commonsourceibias.n100 commonsourceibias.n23 0.189894
R967 commonsourceibias.n95 commonsourceibias.n23 0.189894
R968 commonsourceibias.n95 commonsourceibias.n94 0.189894
R969 commonsourceibias.n94 commonsourceibias.n93 0.189894
R970 commonsourceibias.n93 commonsourceibias.n26 0.189894
R971 commonsourceibias.n88 commonsourceibias.n26 0.189894
R972 commonsourceibias.n88 commonsourceibias.n87 0.189894
R973 commonsourceibias.n87 commonsourceibias.n86 0.189894
R974 commonsourceibias.n86 commonsourceibias.n28 0.189894
R975 commonsourceibias.n81 commonsourceibias.n28 0.189894
R976 commonsourceibias.n81 commonsourceibias.n80 0.189894
R977 commonsourceibias.n80 commonsourceibias.n79 0.189894
R978 commonsourceibias.n79 commonsourceibias.n31 0.189894
R979 commonsourceibias.n74 commonsourceibias.n31 0.189894
R980 commonsourceibias.n74 commonsourceibias.n73 0.189894
R981 commonsourceibias.n73 commonsourceibias.n72 0.189894
R982 commonsourceibias.n72 commonsourceibias.n33 0.189894
R983 commonsourceibias.n67 commonsourceibias.n33 0.189894
R984 commonsourceibias.n67 commonsourceibias.n66 0.189894
R985 commonsourceibias.n66 commonsourceibias.n65 0.189894
R986 commonsourceibias.n65 commonsourceibias.n36 0.189894
R987 commonsourceibias.n60 commonsourceibias.n36 0.189894
R988 commonsourceibias.n60 commonsourceibias.n59 0.189894
R989 commonsourceibias.n59 commonsourceibias.n58 0.189894
R990 commonsourceibias.n58 commonsourceibias.n38 0.189894
R991 commonsourceibias.n53 commonsourceibias.n38 0.189894
R992 commonsourceibias.n53 commonsourceibias.n52 0.189894
R993 commonsourceibias.n52 commonsourceibias.n51 0.189894
R994 commonsourceibias.n51 commonsourceibias.n41 0.189894
R995 commonsourceibias.n46 commonsourceibias.n41 0.189894
R996 commonsourceibias.n46 commonsourceibias.n45 0.189894
R997 commonsourceibias.n205 commonsourceibias.n204 0.189894
R998 commonsourceibias.n204 commonsourceibias.n152 0.189894
R999 commonsourceibias.n200 commonsourceibias.n152 0.189894
R1000 commonsourceibias.n200 commonsourceibias.n199 0.189894
R1001 commonsourceibias.n199 commonsourceibias.n154 0.189894
R1002 commonsourceibias.n195 commonsourceibias.n154 0.189894
R1003 commonsourceibias.n195 commonsourceibias.n194 0.189894
R1004 commonsourceibias.n194 commonsourceibias.n156 0.189894
R1005 commonsourceibias.n189 commonsourceibias.n156 0.189894
R1006 commonsourceibias.n189 commonsourceibias.n188 0.189894
R1007 commonsourceibias.n188 commonsourceibias.n187 0.189894
R1008 commonsourceibias.n187 commonsourceibias.n158 0.189894
R1009 commonsourceibias.n182 commonsourceibias.n158 0.189894
R1010 commonsourceibias.n182 commonsourceibias.n181 0.189894
R1011 commonsourceibias.n181 commonsourceibias.n180 0.189894
R1012 commonsourceibias.n180 commonsourceibias.n160 0.189894
R1013 commonsourceibias.n175 commonsourceibias.n160 0.189894
R1014 commonsourceibias.n175 commonsourceibias.n174 0.189894
R1015 commonsourceibias.n174 commonsourceibias.n173 0.189894
R1016 commonsourceibias.n173 commonsourceibias.n163 0.189894
R1017 commonsourceibias.n168 commonsourceibias.n163 0.189894
R1018 commonsourceibias.n168 commonsourceibias.n167 0.189894
R1019 commonsourceibias.n245 commonsourceibias.n0 0.189894
R1020 commonsourceibias.n245 commonsourceibias.n244 0.189894
R1021 commonsourceibias.n244 commonsourceibias.n243 0.189894
R1022 commonsourceibias.n243 commonsourceibias.n2 0.189894
R1023 commonsourceibias.n238 commonsourceibias.n2 0.189894
R1024 commonsourceibias.n238 commonsourceibias.n237 0.189894
R1025 commonsourceibias.n237 commonsourceibias.n236 0.189894
R1026 commonsourceibias.n236 commonsourceibias.n4 0.189894
R1027 commonsourceibias.n231 commonsourceibias.n4 0.189894
R1028 commonsourceibias.n231 commonsourceibias.n230 0.189894
R1029 commonsourceibias.n230 commonsourceibias.n229 0.189894
R1030 commonsourceibias.n229 commonsourceibias.n7 0.189894
R1031 commonsourceibias.n224 commonsourceibias.n7 0.189894
R1032 commonsourceibias.n224 commonsourceibias.n223 0.189894
R1033 commonsourceibias.n223 commonsourceibias.n222 0.189894
R1034 commonsourceibias.n222 commonsourceibias.n9 0.189894
R1035 commonsourceibias.n217 commonsourceibias.n9 0.189894
R1036 commonsourceibias.n217 commonsourceibias.n216 0.189894
R1037 commonsourceibias.n216 commonsourceibias.n215 0.189894
R1038 commonsourceibias.n215 commonsourceibias.n12 0.189894
R1039 commonsourceibias.n210 commonsourceibias.n12 0.189894
R1040 commonsourceibias.n210 commonsourceibias.n209 0.189894
R1041 commonsourceibias.n209 commonsourceibias.n208 0.189894
R1042 commonsourceibias.n645 commonsourceibias.n644 0.189894
R1043 commonsourceibias.n645 commonsourceibias.n640 0.189894
R1044 commonsourceibias.n650 commonsourceibias.n640 0.189894
R1045 commonsourceibias.n651 commonsourceibias.n650 0.189894
R1046 commonsourceibias.n652 commonsourceibias.n651 0.189894
R1047 commonsourceibias.n652 commonsourceibias.n638 0.189894
R1048 commonsourceibias.n658 commonsourceibias.n638 0.189894
R1049 commonsourceibias.n659 commonsourceibias.n658 0.189894
R1050 commonsourceibias.n660 commonsourceibias.n659 0.189894
R1051 commonsourceibias.n660 commonsourceibias.n636 0.189894
R1052 commonsourceibias.n665 commonsourceibias.n636 0.189894
R1053 commonsourceibias.n666 commonsourceibias.n665 0.189894
R1054 commonsourceibias.n667 commonsourceibias.n666 0.189894
R1055 commonsourceibias.n667 commonsourceibias.n634 0.189894
R1056 commonsourceibias.n673 commonsourceibias.n634 0.189894
R1057 commonsourceibias.n674 commonsourceibias.n673 0.189894
R1058 commonsourceibias.n675 commonsourceibias.n674 0.189894
R1059 commonsourceibias.n675 commonsourceibias.n632 0.189894
R1060 commonsourceibias.n680 commonsourceibias.n632 0.189894
R1061 commonsourceibias.n681 commonsourceibias.n680 0.189894
R1062 commonsourceibias.n682 commonsourceibias.n681 0.189894
R1063 commonsourceibias.n682 commonsourceibias.n630 0.189894
R1064 commonsourceibias.n688 commonsourceibias.n630 0.189894
R1065 commonsourceibias.n689 commonsourceibias.n688 0.189894
R1066 commonsourceibias.n690 commonsourceibias.n689 0.189894
R1067 commonsourceibias.n690 commonsourceibias.n628 0.189894
R1068 commonsourceibias.n695 commonsourceibias.n628 0.189894
R1069 commonsourceibias.n696 commonsourceibias.n695 0.189894
R1070 commonsourceibias.n697 commonsourceibias.n696 0.189894
R1071 commonsourceibias.n697 commonsourceibias.n626 0.189894
R1072 commonsourceibias.n703 commonsourceibias.n626 0.189894
R1073 commonsourceibias.n704 commonsourceibias.n703 0.189894
R1074 commonsourceibias.n705 commonsourceibias.n704 0.189894
R1075 commonsourceibias.n705 commonsourceibias.n624 0.189894
R1076 commonsourceibias.n710 commonsourceibias.n624 0.189894
R1077 commonsourceibias.n711 commonsourceibias.n710 0.189894
R1078 commonsourceibias.n712 commonsourceibias.n711 0.189894
R1079 commonsourceibias.n712 commonsourceibias.n622 0.189894
R1080 commonsourceibias.n718 commonsourceibias.n622 0.189894
R1081 commonsourceibias.n719 commonsourceibias.n718 0.189894
R1082 commonsourceibias.n720 commonsourceibias.n719 0.189894
R1083 commonsourceibias.n720 commonsourceibias.n620 0.189894
R1084 commonsourceibias.n725 commonsourceibias.n620 0.189894
R1085 commonsourceibias.n726 commonsourceibias.n725 0.189894
R1086 commonsourceibias.n727 commonsourceibias.n726 0.189894
R1087 commonsourceibias.n727 commonsourceibias.n618 0.189894
R1088 commonsourceibias.n415 commonsourceibias.n414 0.189894
R1089 commonsourceibias.n415 commonsourceibias.n410 0.189894
R1090 commonsourceibias.n420 commonsourceibias.n410 0.189894
R1091 commonsourceibias.n421 commonsourceibias.n420 0.189894
R1092 commonsourceibias.n422 commonsourceibias.n421 0.189894
R1093 commonsourceibias.n422 commonsourceibias.n408 0.189894
R1094 commonsourceibias.n428 commonsourceibias.n408 0.189894
R1095 commonsourceibias.n429 commonsourceibias.n428 0.189894
R1096 commonsourceibias.n430 commonsourceibias.n429 0.189894
R1097 commonsourceibias.n430 commonsourceibias.n406 0.189894
R1098 commonsourceibias.n435 commonsourceibias.n406 0.189894
R1099 commonsourceibias.n436 commonsourceibias.n435 0.189894
R1100 commonsourceibias.n437 commonsourceibias.n436 0.189894
R1101 commonsourceibias.n437 commonsourceibias.n404 0.189894
R1102 commonsourceibias.n443 commonsourceibias.n404 0.189894
R1103 commonsourceibias.n444 commonsourceibias.n443 0.189894
R1104 commonsourceibias.n445 commonsourceibias.n444 0.189894
R1105 commonsourceibias.n445 commonsourceibias.n402 0.189894
R1106 commonsourceibias.n450 commonsourceibias.n402 0.189894
R1107 commonsourceibias.n451 commonsourceibias.n450 0.189894
R1108 commonsourceibias.n452 commonsourceibias.n451 0.189894
R1109 commonsourceibias.n452 commonsourceibias.n400 0.189894
R1110 commonsourceibias.n458 commonsourceibias.n400 0.189894
R1111 commonsourceibias.n459 commonsourceibias.n458 0.189894
R1112 commonsourceibias.n460 commonsourceibias.n459 0.189894
R1113 commonsourceibias.n460 commonsourceibias.n398 0.189894
R1114 commonsourceibias.n465 commonsourceibias.n398 0.189894
R1115 commonsourceibias.n466 commonsourceibias.n465 0.189894
R1116 commonsourceibias.n467 commonsourceibias.n466 0.189894
R1117 commonsourceibias.n467 commonsourceibias.n396 0.189894
R1118 commonsourceibias.n473 commonsourceibias.n396 0.189894
R1119 commonsourceibias.n474 commonsourceibias.n473 0.189894
R1120 commonsourceibias.n475 commonsourceibias.n474 0.189894
R1121 commonsourceibias.n475 commonsourceibias.n394 0.189894
R1122 commonsourceibias.n480 commonsourceibias.n394 0.189894
R1123 commonsourceibias.n481 commonsourceibias.n480 0.189894
R1124 commonsourceibias.n482 commonsourceibias.n481 0.189894
R1125 commonsourceibias.n482 commonsourceibias.n392 0.189894
R1126 commonsourceibias.n488 commonsourceibias.n392 0.189894
R1127 commonsourceibias.n489 commonsourceibias.n488 0.189894
R1128 commonsourceibias.n490 commonsourceibias.n489 0.189894
R1129 commonsourceibias.n490 commonsourceibias.n390 0.189894
R1130 commonsourceibias.n495 commonsourceibias.n390 0.189894
R1131 commonsourceibias.n496 commonsourceibias.n495 0.189894
R1132 commonsourceibias.n497 commonsourceibias.n496 0.189894
R1133 commonsourceibias.n497 commonsourceibias.n388 0.189894
R1134 commonsourceibias.n531 commonsourceibias.n530 0.189894
R1135 commonsourceibias.n531 commonsourceibias.n526 0.189894
R1136 commonsourceibias.n536 commonsourceibias.n526 0.189894
R1137 commonsourceibias.n537 commonsourceibias.n536 0.189894
R1138 commonsourceibias.n538 commonsourceibias.n537 0.189894
R1139 commonsourceibias.n538 commonsourceibias.n524 0.189894
R1140 commonsourceibias.n544 commonsourceibias.n524 0.189894
R1141 commonsourceibias.n545 commonsourceibias.n544 0.189894
R1142 commonsourceibias.n546 commonsourceibias.n545 0.189894
R1143 commonsourceibias.n546 commonsourceibias.n522 0.189894
R1144 commonsourceibias.n551 commonsourceibias.n522 0.189894
R1145 commonsourceibias.n552 commonsourceibias.n551 0.189894
R1146 commonsourceibias.n553 commonsourceibias.n552 0.189894
R1147 commonsourceibias.n553 commonsourceibias.n520 0.189894
R1148 commonsourceibias.n558 commonsourceibias.n520 0.189894
R1149 commonsourceibias.n559 commonsourceibias.n558 0.189894
R1150 commonsourceibias.n559 commonsourceibias.n518 0.189894
R1151 commonsourceibias.n563 commonsourceibias.n518 0.189894
R1152 commonsourceibias.n564 commonsourceibias.n563 0.189894
R1153 commonsourceibias.n564 commonsourceibias.n516 0.189894
R1154 commonsourceibias.n568 commonsourceibias.n516 0.189894
R1155 commonsourceibias.n569 commonsourceibias.n568 0.189894
R1156 commonsourceibias.n574 commonsourceibias.n573 0.189894
R1157 commonsourceibias.n575 commonsourceibias.n574 0.189894
R1158 commonsourceibias.n575 commonsourceibias.n377 0.189894
R1159 commonsourceibias.n580 commonsourceibias.n377 0.189894
R1160 commonsourceibias.n581 commonsourceibias.n580 0.189894
R1161 commonsourceibias.n582 commonsourceibias.n581 0.189894
R1162 commonsourceibias.n582 commonsourceibias.n375 0.189894
R1163 commonsourceibias.n588 commonsourceibias.n375 0.189894
R1164 commonsourceibias.n589 commonsourceibias.n588 0.189894
R1165 commonsourceibias.n590 commonsourceibias.n589 0.189894
R1166 commonsourceibias.n590 commonsourceibias.n373 0.189894
R1167 commonsourceibias.n595 commonsourceibias.n373 0.189894
R1168 commonsourceibias.n596 commonsourceibias.n595 0.189894
R1169 commonsourceibias.n597 commonsourceibias.n596 0.189894
R1170 commonsourceibias.n597 commonsourceibias.n371 0.189894
R1171 commonsourceibias.n603 commonsourceibias.n371 0.189894
R1172 commonsourceibias.n604 commonsourceibias.n603 0.189894
R1173 commonsourceibias.n605 commonsourceibias.n604 0.189894
R1174 commonsourceibias.n605 commonsourceibias.n369 0.189894
R1175 commonsourceibias.n610 commonsourceibias.n369 0.189894
R1176 commonsourceibias.n611 commonsourceibias.n610 0.189894
R1177 commonsourceibias.n612 commonsourceibias.n611 0.189894
R1178 commonsourceibias.n612 commonsourceibias.n367 0.189894
R1179 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R1180 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R1181 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R1182 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R1183 CSoutput.n19 CSoutput.t206 184.661
R1184 CSoutput.n78 CSoutput.n77 165.8
R1185 CSoutput.n76 CSoutput.n0 165.8
R1186 CSoutput.n75 CSoutput.n74 165.8
R1187 CSoutput.n73 CSoutput.n72 165.8
R1188 CSoutput.n71 CSoutput.n2 165.8
R1189 CSoutput.n69 CSoutput.n68 165.8
R1190 CSoutput.n67 CSoutput.n3 165.8
R1191 CSoutput.n66 CSoutput.n65 165.8
R1192 CSoutput.n63 CSoutput.n4 165.8
R1193 CSoutput.n61 CSoutput.n60 165.8
R1194 CSoutput.n59 CSoutput.n5 165.8
R1195 CSoutput.n58 CSoutput.n57 165.8
R1196 CSoutput.n55 CSoutput.n6 165.8
R1197 CSoutput.n54 CSoutput.n53 165.8
R1198 CSoutput.n52 CSoutput.n51 165.8
R1199 CSoutput.n50 CSoutput.n8 165.8
R1200 CSoutput.n48 CSoutput.n47 165.8
R1201 CSoutput.n46 CSoutput.n9 165.8
R1202 CSoutput.n45 CSoutput.n44 165.8
R1203 CSoutput.n42 CSoutput.n10 165.8
R1204 CSoutput.n41 CSoutput.n40 165.8
R1205 CSoutput.n39 CSoutput.n38 165.8
R1206 CSoutput.n37 CSoutput.n12 165.8
R1207 CSoutput.n35 CSoutput.n34 165.8
R1208 CSoutput.n33 CSoutput.n13 165.8
R1209 CSoutput.n32 CSoutput.n31 165.8
R1210 CSoutput.n29 CSoutput.n14 165.8
R1211 CSoutput.n28 CSoutput.n27 165.8
R1212 CSoutput.n26 CSoutput.n25 165.8
R1213 CSoutput.n24 CSoutput.n16 165.8
R1214 CSoutput.n22 CSoutput.n21 165.8
R1215 CSoutput.n20 CSoutput.n17 165.8
R1216 CSoutput.n77 CSoutput.t208 162.194
R1217 CSoutput.n18 CSoutput.t217 120.501
R1218 CSoutput.n23 CSoutput.t219 120.501
R1219 CSoutput.n15 CSoutput.t212 120.501
R1220 CSoutput.n30 CSoutput.t203 120.501
R1221 CSoutput.n36 CSoutput.t221 120.501
R1222 CSoutput.n11 CSoutput.t215 120.501
R1223 CSoutput.n43 CSoutput.t210 120.501
R1224 CSoutput.n49 CSoutput.t201 120.501
R1225 CSoutput.n7 CSoutput.t202 120.501
R1226 CSoutput.n56 CSoutput.t213 120.501
R1227 CSoutput.n62 CSoutput.t209 120.501
R1228 CSoutput.n64 CSoutput.t205 120.501
R1229 CSoutput.n70 CSoutput.t216 120.501
R1230 CSoutput.n1 CSoutput.t218 120.501
R1231 CSoutput.n330 CSoutput.n328 103.469
R1232 CSoutput.n310 CSoutput.n308 103.469
R1233 CSoutput.n291 CSoutput.n289 103.469
R1234 CSoutput.n120 CSoutput.n118 103.469
R1235 CSoutput.n100 CSoutput.n98 103.469
R1236 CSoutput.n81 CSoutput.n79 103.469
R1237 CSoutput.n344 CSoutput.n343 103.111
R1238 CSoutput.n342 CSoutput.n341 103.111
R1239 CSoutput.n340 CSoutput.n339 103.111
R1240 CSoutput.n338 CSoutput.n337 103.111
R1241 CSoutput.n336 CSoutput.n335 103.111
R1242 CSoutput.n334 CSoutput.n333 103.111
R1243 CSoutput.n332 CSoutput.n331 103.111
R1244 CSoutput.n330 CSoutput.n329 103.111
R1245 CSoutput.n326 CSoutput.n325 103.111
R1246 CSoutput.n324 CSoutput.n323 103.111
R1247 CSoutput.n322 CSoutput.n321 103.111
R1248 CSoutput.n320 CSoutput.n319 103.111
R1249 CSoutput.n318 CSoutput.n317 103.111
R1250 CSoutput.n316 CSoutput.n315 103.111
R1251 CSoutput.n314 CSoutput.n313 103.111
R1252 CSoutput.n312 CSoutput.n311 103.111
R1253 CSoutput.n310 CSoutput.n309 103.111
R1254 CSoutput.n307 CSoutput.n306 103.111
R1255 CSoutput.n305 CSoutput.n304 103.111
R1256 CSoutput.n303 CSoutput.n302 103.111
R1257 CSoutput.n301 CSoutput.n300 103.111
R1258 CSoutput.n299 CSoutput.n298 103.111
R1259 CSoutput.n297 CSoutput.n296 103.111
R1260 CSoutput.n295 CSoutput.n294 103.111
R1261 CSoutput.n293 CSoutput.n292 103.111
R1262 CSoutput.n291 CSoutput.n290 103.111
R1263 CSoutput.n120 CSoutput.n119 103.111
R1264 CSoutput.n122 CSoutput.n121 103.111
R1265 CSoutput.n124 CSoutput.n123 103.111
R1266 CSoutput.n126 CSoutput.n125 103.111
R1267 CSoutput.n128 CSoutput.n127 103.111
R1268 CSoutput.n130 CSoutput.n129 103.111
R1269 CSoutput.n132 CSoutput.n131 103.111
R1270 CSoutput.n134 CSoutput.n133 103.111
R1271 CSoutput.n136 CSoutput.n135 103.111
R1272 CSoutput.n100 CSoutput.n99 103.111
R1273 CSoutput.n102 CSoutput.n101 103.111
R1274 CSoutput.n104 CSoutput.n103 103.111
R1275 CSoutput.n106 CSoutput.n105 103.111
R1276 CSoutput.n108 CSoutput.n107 103.111
R1277 CSoutput.n110 CSoutput.n109 103.111
R1278 CSoutput.n112 CSoutput.n111 103.111
R1279 CSoutput.n114 CSoutput.n113 103.111
R1280 CSoutput.n116 CSoutput.n115 103.111
R1281 CSoutput.n81 CSoutput.n80 103.111
R1282 CSoutput.n83 CSoutput.n82 103.111
R1283 CSoutput.n85 CSoutput.n84 103.111
R1284 CSoutput.n87 CSoutput.n86 103.111
R1285 CSoutput.n89 CSoutput.n88 103.111
R1286 CSoutput.n91 CSoutput.n90 103.111
R1287 CSoutput.n93 CSoutput.n92 103.111
R1288 CSoutput.n95 CSoutput.n94 103.111
R1289 CSoutput.n97 CSoutput.n96 103.111
R1290 CSoutput.n346 CSoutput.n345 103.111
R1291 CSoutput.n370 CSoutput.n368 81.5057
R1292 CSoutput.n351 CSoutput.n349 81.5057
R1293 CSoutput.n410 CSoutput.n408 81.5057
R1294 CSoutput.n391 CSoutput.n389 81.5057
R1295 CSoutput.n386 CSoutput.n385 80.9324
R1296 CSoutput.n384 CSoutput.n383 80.9324
R1297 CSoutput.n382 CSoutput.n381 80.9324
R1298 CSoutput.n380 CSoutput.n379 80.9324
R1299 CSoutput.n378 CSoutput.n377 80.9324
R1300 CSoutput.n376 CSoutput.n375 80.9324
R1301 CSoutput.n374 CSoutput.n373 80.9324
R1302 CSoutput.n372 CSoutput.n371 80.9324
R1303 CSoutput.n370 CSoutput.n369 80.9324
R1304 CSoutput.n367 CSoutput.n366 80.9324
R1305 CSoutput.n365 CSoutput.n364 80.9324
R1306 CSoutput.n363 CSoutput.n362 80.9324
R1307 CSoutput.n361 CSoutput.n360 80.9324
R1308 CSoutput.n359 CSoutput.n358 80.9324
R1309 CSoutput.n357 CSoutput.n356 80.9324
R1310 CSoutput.n355 CSoutput.n354 80.9324
R1311 CSoutput.n353 CSoutput.n352 80.9324
R1312 CSoutput.n351 CSoutput.n350 80.9324
R1313 CSoutput.n410 CSoutput.n409 80.9324
R1314 CSoutput.n412 CSoutput.n411 80.9324
R1315 CSoutput.n414 CSoutput.n413 80.9324
R1316 CSoutput.n416 CSoutput.n415 80.9324
R1317 CSoutput.n418 CSoutput.n417 80.9324
R1318 CSoutput.n420 CSoutput.n419 80.9324
R1319 CSoutput.n422 CSoutput.n421 80.9324
R1320 CSoutput.n424 CSoutput.n423 80.9324
R1321 CSoutput.n426 CSoutput.n425 80.9324
R1322 CSoutput.n391 CSoutput.n390 80.9324
R1323 CSoutput.n393 CSoutput.n392 80.9324
R1324 CSoutput.n395 CSoutput.n394 80.9324
R1325 CSoutput.n397 CSoutput.n396 80.9324
R1326 CSoutput.n399 CSoutput.n398 80.9324
R1327 CSoutput.n401 CSoutput.n400 80.9324
R1328 CSoutput.n403 CSoutput.n402 80.9324
R1329 CSoutput.n405 CSoutput.n404 80.9324
R1330 CSoutput.n407 CSoutput.n406 80.9324
R1331 CSoutput.n25 CSoutput.n24 48.1486
R1332 CSoutput.n69 CSoutput.n3 48.1486
R1333 CSoutput.n38 CSoutput.n37 48.1486
R1334 CSoutput.n42 CSoutput.n41 48.1486
R1335 CSoutput.n51 CSoutput.n50 48.1486
R1336 CSoutput.n55 CSoutput.n54 48.1486
R1337 CSoutput.n22 CSoutput.n17 46.462
R1338 CSoutput.n72 CSoutput.n71 46.462
R1339 CSoutput.n20 CSoutput.n19 44.9055
R1340 CSoutput.n29 CSoutput.n28 43.7635
R1341 CSoutput.n65 CSoutput.n63 43.7635
R1342 CSoutput.n35 CSoutput.n13 41.7396
R1343 CSoutput.n57 CSoutput.n5 41.7396
R1344 CSoutput.n44 CSoutput.n9 37.0171
R1345 CSoutput.n48 CSoutput.n9 37.0171
R1346 CSoutput.n76 CSoutput.n75 34.9932
R1347 CSoutput.n31 CSoutput.n13 32.2947
R1348 CSoutput.n61 CSoutput.n5 32.2947
R1349 CSoutput.n30 CSoutput.n29 29.6014
R1350 CSoutput.n63 CSoutput.n62 29.6014
R1351 CSoutput.n19 CSoutput.n18 28.4085
R1352 CSoutput.n18 CSoutput.n17 25.1176
R1353 CSoutput.n72 CSoutput.n1 25.1176
R1354 CSoutput.n43 CSoutput.n42 22.0922
R1355 CSoutput.n50 CSoutput.n49 22.0922
R1356 CSoutput.n77 CSoutput.n76 21.8586
R1357 CSoutput.n37 CSoutput.n36 18.9681
R1358 CSoutput.n56 CSoutput.n55 18.9681
R1359 CSoutput.n25 CSoutput.n15 17.6292
R1360 CSoutput.n64 CSoutput.n3 17.6292
R1361 CSoutput.n24 CSoutput.n23 15.844
R1362 CSoutput.n70 CSoutput.n69 15.844
R1363 CSoutput.n38 CSoutput.n11 14.5051
R1364 CSoutput.n54 CSoutput.n7 14.5051
R1365 CSoutput.n429 CSoutput.n78 11.6139
R1366 CSoutput.n41 CSoutput.n11 11.3811
R1367 CSoutput.n51 CSoutput.n7 11.3811
R1368 CSoutput.n23 CSoutput.n22 10.0422
R1369 CSoutput.n71 CSoutput.n70 10.0422
R1370 CSoutput.n327 CSoutput.n307 9.25285
R1371 CSoutput.n117 CSoutput.n97 9.25285
R1372 CSoutput.n387 CSoutput.n367 8.97993
R1373 CSoutput.n427 CSoutput.n407 8.97993
R1374 CSoutput.n388 CSoutput.n348 8.84557
R1375 CSoutput.n28 CSoutput.n15 8.25698
R1376 CSoutput.n65 CSoutput.n64 8.25698
R1377 CSoutput.n388 CSoutput.n387 7.89345
R1378 CSoutput.n428 CSoutput.n427 7.89345
R1379 CSoutput.n348 CSoutput.n347 7.12641
R1380 CSoutput.n138 CSoutput.n137 7.12641
R1381 CSoutput.n36 CSoutput.n35 6.91809
R1382 CSoutput.n57 CSoutput.n56 6.91809
R1383 CSoutput.n429 CSoutput.n138 5.25314
R1384 CSoutput.n387 CSoutput.n386 5.25266
R1385 CSoutput.n427 CSoutput.n426 5.25266
R1386 CSoutput.n347 CSoutput.n346 5.1449
R1387 CSoutput.n327 CSoutput.n326 5.1449
R1388 CSoutput.n137 CSoutput.n136 5.1449
R1389 CSoutput.n117 CSoutput.n116 5.1449
R1390 CSoutput.n229 CSoutput.n182 4.5005
R1391 CSoutput.n198 CSoutput.n182 4.5005
R1392 CSoutput.n193 CSoutput.n177 4.5005
R1393 CSoutput.n193 CSoutput.n179 4.5005
R1394 CSoutput.n193 CSoutput.n176 4.5005
R1395 CSoutput.n193 CSoutput.n180 4.5005
R1396 CSoutput.n193 CSoutput.n175 4.5005
R1397 CSoutput.n193 CSoutput.t220 4.5005
R1398 CSoutput.n193 CSoutput.n174 4.5005
R1399 CSoutput.n193 CSoutput.n181 4.5005
R1400 CSoutput.n193 CSoutput.n182 4.5005
R1401 CSoutput.n191 CSoutput.n177 4.5005
R1402 CSoutput.n191 CSoutput.n179 4.5005
R1403 CSoutput.n191 CSoutput.n176 4.5005
R1404 CSoutput.n191 CSoutput.n180 4.5005
R1405 CSoutput.n191 CSoutput.n175 4.5005
R1406 CSoutput.n191 CSoutput.t220 4.5005
R1407 CSoutput.n191 CSoutput.n174 4.5005
R1408 CSoutput.n191 CSoutput.n181 4.5005
R1409 CSoutput.n191 CSoutput.n182 4.5005
R1410 CSoutput.n190 CSoutput.n177 4.5005
R1411 CSoutput.n190 CSoutput.n179 4.5005
R1412 CSoutput.n190 CSoutput.n176 4.5005
R1413 CSoutput.n190 CSoutput.n180 4.5005
R1414 CSoutput.n190 CSoutput.n175 4.5005
R1415 CSoutput.n190 CSoutput.t220 4.5005
R1416 CSoutput.n190 CSoutput.n174 4.5005
R1417 CSoutput.n190 CSoutput.n181 4.5005
R1418 CSoutput.n190 CSoutput.n182 4.5005
R1419 CSoutput.n275 CSoutput.n177 4.5005
R1420 CSoutput.n275 CSoutput.n179 4.5005
R1421 CSoutput.n275 CSoutput.n176 4.5005
R1422 CSoutput.n275 CSoutput.n180 4.5005
R1423 CSoutput.n275 CSoutput.n175 4.5005
R1424 CSoutput.n275 CSoutput.t220 4.5005
R1425 CSoutput.n275 CSoutput.n174 4.5005
R1426 CSoutput.n275 CSoutput.n181 4.5005
R1427 CSoutput.n275 CSoutput.n182 4.5005
R1428 CSoutput.n273 CSoutput.n177 4.5005
R1429 CSoutput.n273 CSoutput.n179 4.5005
R1430 CSoutput.n273 CSoutput.n176 4.5005
R1431 CSoutput.n273 CSoutput.n180 4.5005
R1432 CSoutput.n273 CSoutput.n175 4.5005
R1433 CSoutput.n273 CSoutput.t220 4.5005
R1434 CSoutput.n273 CSoutput.n174 4.5005
R1435 CSoutput.n273 CSoutput.n181 4.5005
R1436 CSoutput.n271 CSoutput.n177 4.5005
R1437 CSoutput.n271 CSoutput.n179 4.5005
R1438 CSoutput.n271 CSoutput.n176 4.5005
R1439 CSoutput.n271 CSoutput.n180 4.5005
R1440 CSoutput.n271 CSoutput.n175 4.5005
R1441 CSoutput.n271 CSoutput.t220 4.5005
R1442 CSoutput.n271 CSoutput.n174 4.5005
R1443 CSoutput.n271 CSoutput.n181 4.5005
R1444 CSoutput.n201 CSoutput.n177 4.5005
R1445 CSoutput.n201 CSoutput.n179 4.5005
R1446 CSoutput.n201 CSoutput.n176 4.5005
R1447 CSoutput.n201 CSoutput.n180 4.5005
R1448 CSoutput.n201 CSoutput.n175 4.5005
R1449 CSoutput.n201 CSoutput.t220 4.5005
R1450 CSoutput.n201 CSoutput.n174 4.5005
R1451 CSoutput.n201 CSoutput.n181 4.5005
R1452 CSoutput.n201 CSoutput.n182 4.5005
R1453 CSoutput.n200 CSoutput.n177 4.5005
R1454 CSoutput.n200 CSoutput.n179 4.5005
R1455 CSoutput.n200 CSoutput.n176 4.5005
R1456 CSoutput.n200 CSoutput.n180 4.5005
R1457 CSoutput.n200 CSoutput.n175 4.5005
R1458 CSoutput.n200 CSoutput.t220 4.5005
R1459 CSoutput.n200 CSoutput.n174 4.5005
R1460 CSoutput.n200 CSoutput.n181 4.5005
R1461 CSoutput.n200 CSoutput.n182 4.5005
R1462 CSoutput.n204 CSoutput.n177 4.5005
R1463 CSoutput.n204 CSoutput.n179 4.5005
R1464 CSoutput.n204 CSoutput.n176 4.5005
R1465 CSoutput.n204 CSoutput.n180 4.5005
R1466 CSoutput.n204 CSoutput.n175 4.5005
R1467 CSoutput.n204 CSoutput.t220 4.5005
R1468 CSoutput.n204 CSoutput.n174 4.5005
R1469 CSoutput.n204 CSoutput.n181 4.5005
R1470 CSoutput.n204 CSoutput.n182 4.5005
R1471 CSoutput.n203 CSoutput.n177 4.5005
R1472 CSoutput.n203 CSoutput.n179 4.5005
R1473 CSoutput.n203 CSoutput.n176 4.5005
R1474 CSoutput.n203 CSoutput.n180 4.5005
R1475 CSoutput.n203 CSoutput.n175 4.5005
R1476 CSoutput.n203 CSoutput.t220 4.5005
R1477 CSoutput.n203 CSoutput.n174 4.5005
R1478 CSoutput.n203 CSoutput.n181 4.5005
R1479 CSoutput.n203 CSoutput.n182 4.5005
R1480 CSoutput.n186 CSoutput.n177 4.5005
R1481 CSoutput.n186 CSoutput.n179 4.5005
R1482 CSoutput.n186 CSoutput.n176 4.5005
R1483 CSoutput.n186 CSoutput.n180 4.5005
R1484 CSoutput.n186 CSoutput.n175 4.5005
R1485 CSoutput.n186 CSoutput.t220 4.5005
R1486 CSoutput.n186 CSoutput.n174 4.5005
R1487 CSoutput.n186 CSoutput.n181 4.5005
R1488 CSoutput.n186 CSoutput.n182 4.5005
R1489 CSoutput.n278 CSoutput.n177 4.5005
R1490 CSoutput.n278 CSoutput.n179 4.5005
R1491 CSoutput.n278 CSoutput.n176 4.5005
R1492 CSoutput.n278 CSoutput.n180 4.5005
R1493 CSoutput.n278 CSoutput.n175 4.5005
R1494 CSoutput.n278 CSoutput.t220 4.5005
R1495 CSoutput.n278 CSoutput.n174 4.5005
R1496 CSoutput.n278 CSoutput.n181 4.5005
R1497 CSoutput.n278 CSoutput.n182 4.5005
R1498 CSoutput.n265 CSoutput.n236 4.5005
R1499 CSoutput.n265 CSoutput.n242 4.5005
R1500 CSoutput.n223 CSoutput.n212 4.5005
R1501 CSoutput.n223 CSoutput.n214 4.5005
R1502 CSoutput.n223 CSoutput.n211 4.5005
R1503 CSoutput.n223 CSoutput.n215 4.5005
R1504 CSoutput.n223 CSoutput.n210 4.5005
R1505 CSoutput.n223 CSoutput.t214 4.5005
R1506 CSoutput.n223 CSoutput.n209 4.5005
R1507 CSoutput.n223 CSoutput.n216 4.5005
R1508 CSoutput.n265 CSoutput.n223 4.5005
R1509 CSoutput.n244 CSoutput.n212 4.5005
R1510 CSoutput.n244 CSoutput.n214 4.5005
R1511 CSoutput.n244 CSoutput.n211 4.5005
R1512 CSoutput.n244 CSoutput.n215 4.5005
R1513 CSoutput.n244 CSoutput.n210 4.5005
R1514 CSoutput.n244 CSoutput.t214 4.5005
R1515 CSoutput.n244 CSoutput.n209 4.5005
R1516 CSoutput.n244 CSoutput.n216 4.5005
R1517 CSoutput.n265 CSoutput.n244 4.5005
R1518 CSoutput.n222 CSoutput.n212 4.5005
R1519 CSoutput.n222 CSoutput.n214 4.5005
R1520 CSoutput.n222 CSoutput.n211 4.5005
R1521 CSoutput.n222 CSoutput.n215 4.5005
R1522 CSoutput.n222 CSoutput.n210 4.5005
R1523 CSoutput.n222 CSoutput.t214 4.5005
R1524 CSoutput.n222 CSoutput.n209 4.5005
R1525 CSoutput.n222 CSoutput.n216 4.5005
R1526 CSoutput.n265 CSoutput.n222 4.5005
R1527 CSoutput.n246 CSoutput.n212 4.5005
R1528 CSoutput.n246 CSoutput.n214 4.5005
R1529 CSoutput.n246 CSoutput.n211 4.5005
R1530 CSoutput.n246 CSoutput.n215 4.5005
R1531 CSoutput.n246 CSoutput.n210 4.5005
R1532 CSoutput.n246 CSoutput.t214 4.5005
R1533 CSoutput.n246 CSoutput.n209 4.5005
R1534 CSoutput.n246 CSoutput.n216 4.5005
R1535 CSoutput.n265 CSoutput.n246 4.5005
R1536 CSoutput.n212 CSoutput.n207 4.5005
R1537 CSoutput.n214 CSoutput.n207 4.5005
R1538 CSoutput.n211 CSoutput.n207 4.5005
R1539 CSoutput.n215 CSoutput.n207 4.5005
R1540 CSoutput.n210 CSoutput.n207 4.5005
R1541 CSoutput.t214 CSoutput.n207 4.5005
R1542 CSoutput.n209 CSoutput.n207 4.5005
R1543 CSoutput.n216 CSoutput.n207 4.5005
R1544 CSoutput.n268 CSoutput.n212 4.5005
R1545 CSoutput.n268 CSoutput.n214 4.5005
R1546 CSoutput.n268 CSoutput.n211 4.5005
R1547 CSoutput.n268 CSoutput.n215 4.5005
R1548 CSoutput.n268 CSoutput.n210 4.5005
R1549 CSoutput.n268 CSoutput.t214 4.5005
R1550 CSoutput.n268 CSoutput.n209 4.5005
R1551 CSoutput.n268 CSoutput.n216 4.5005
R1552 CSoutput.n266 CSoutput.n212 4.5005
R1553 CSoutput.n266 CSoutput.n214 4.5005
R1554 CSoutput.n266 CSoutput.n211 4.5005
R1555 CSoutput.n266 CSoutput.n215 4.5005
R1556 CSoutput.n266 CSoutput.n210 4.5005
R1557 CSoutput.n266 CSoutput.t214 4.5005
R1558 CSoutput.n266 CSoutput.n209 4.5005
R1559 CSoutput.n266 CSoutput.n216 4.5005
R1560 CSoutput.n266 CSoutput.n265 4.5005
R1561 CSoutput.n248 CSoutput.n212 4.5005
R1562 CSoutput.n248 CSoutput.n214 4.5005
R1563 CSoutput.n248 CSoutput.n211 4.5005
R1564 CSoutput.n248 CSoutput.n215 4.5005
R1565 CSoutput.n248 CSoutput.n210 4.5005
R1566 CSoutput.n248 CSoutput.t214 4.5005
R1567 CSoutput.n248 CSoutput.n209 4.5005
R1568 CSoutput.n248 CSoutput.n216 4.5005
R1569 CSoutput.n265 CSoutput.n248 4.5005
R1570 CSoutput.n220 CSoutput.n212 4.5005
R1571 CSoutput.n220 CSoutput.n214 4.5005
R1572 CSoutput.n220 CSoutput.n211 4.5005
R1573 CSoutput.n220 CSoutput.n215 4.5005
R1574 CSoutput.n220 CSoutput.n210 4.5005
R1575 CSoutput.n220 CSoutput.t214 4.5005
R1576 CSoutput.n220 CSoutput.n209 4.5005
R1577 CSoutput.n220 CSoutput.n216 4.5005
R1578 CSoutput.n265 CSoutput.n220 4.5005
R1579 CSoutput.n250 CSoutput.n212 4.5005
R1580 CSoutput.n250 CSoutput.n214 4.5005
R1581 CSoutput.n250 CSoutput.n211 4.5005
R1582 CSoutput.n250 CSoutput.n215 4.5005
R1583 CSoutput.n250 CSoutput.n210 4.5005
R1584 CSoutput.n250 CSoutput.t214 4.5005
R1585 CSoutput.n250 CSoutput.n209 4.5005
R1586 CSoutput.n250 CSoutput.n216 4.5005
R1587 CSoutput.n265 CSoutput.n250 4.5005
R1588 CSoutput.n219 CSoutput.n212 4.5005
R1589 CSoutput.n219 CSoutput.n214 4.5005
R1590 CSoutput.n219 CSoutput.n211 4.5005
R1591 CSoutput.n219 CSoutput.n215 4.5005
R1592 CSoutput.n219 CSoutput.n210 4.5005
R1593 CSoutput.n219 CSoutput.t214 4.5005
R1594 CSoutput.n219 CSoutput.n209 4.5005
R1595 CSoutput.n219 CSoutput.n216 4.5005
R1596 CSoutput.n265 CSoutput.n219 4.5005
R1597 CSoutput.n264 CSoutput.n212 4.5005
R1598 CSoutput.n264 CSoutput.n214 4.5005
R1599 CSoutput.n264 CSoutput.n211 4.5005
R1600 CSoutput.n264 CSoutput.n215 4.5005
R1601 CSoutput.n264 CSoutput.n210 4.5005
R1602 CSoutput.n264 CSoutput.t214 4.5005
R1603 CSoutput.n264 CSoutput.n209 4.5005
R1604 CSoutput.n264 CSoutput.n216 4.5005
R1605 CSoutput.n265 CSoutput.n264 4.5005
R1606 CSoutput.n263 CSoutput.n148 4.5005
R1607 CSoutput.n164 CSoutput.n148 4.5005
R1608 CSoutput.n159 CSoutput.n143 4.5005
R1609 CSoutput.n159 CSoutput.n145 4.5005
R1610 CSoutput.n159 CSoutput.n142 4.5005
R1611 CSoutput.n159 CSoutput.n146 4.5005
R1612 CSoutput.n159 CSoutput.n141 4.5005
R1613 CSoutput.n159 CSoutput.t211 4.5005
R1614 CSoutput.n159 CSoutput.n140 4.5005
R1615 CSoutput.n159 CSoutput.n147 4.5005
R1616 CSoutput.n159 CSoutput.n148 4.5005
R1617 CSoutput.n157 CSoutput.n143 4.5005
R1618 CSoutput.n157 CSoutput.n145 4.5005
R1619 CSoutput.n157 CSoutput.n142 4.5005
R1620 CSoutput.n157 CSoutput.n146 4.5005
R1621 CSoutput.n157 CSoutput.n141 4.5005
R1622 CSoutput.n157 CSoutput.t211 4.5005
R1623 CSoutput.n157 CSoutput.n140 4.5005
R1624 CSoutput.n157 CSoutput.n147 4.5005
R1625 CSoutput.n157 CSoutput.n148 4.5005
R1626 CSoutput.n156 CSoutput.n143 4.5005
R1627 CSoutput.n156 CSoutput.n145 4.5005
R1628 CSoutput.n156 CSoutput.n142 4.5005
R1629 CSoutput.n156 CSoutput.n146 4.5005
R1630 CSoutput.n156 CSoutput.n141 4.5005
R1631 CSoutput.n156 CSoutput.t211 4.5005
R1632 CSoutput.n156 CSoutput.n140 4.5005
R1633 CSoutput.n156 CSoutput.n147 4.5005
R1634 CSoutput.n156 CSoutput.n148 4.5005
R1635 CSoutput.n285 CSoutput.n143 4.5005
R1636 CSoutput.n285 CSoutput.n145 4.5005
R1637 CSoutput.n285 CSoutput.n142 4.5005
R1638 CSoutput.n285 CSoutput.n146 4.5005
R1639 CSoutput.n285 CSoutput.n141 4.5005
R1640 CSoutput.n285 CSoutput.t211 4.5005
R1641 CSoutput.n285 CSoutput.n140 4.5005
R1642 CSoutput.n285 CSoutput.n147 4.5005
R1643 CSoutput.n285 CSoutput.n148 4.5005
R1644 CSoutput.n283 CSoutput.n143 4.5005
R1645 CSoutput.n283 CSoutput.n145 4.5005
R1646 CSoutput.n283 CSoutput.n142 4.5005
R1647 CSoutput.n283 CSoutput.n146 4.5005
R1648 CSoutput.n283 CSoutput.n141 4.5005
R1649 CSoutput.n283 CSoutput.t211 4.5005
R1650 CSoutput.n283 CSoutput.n140 4.5005
R1651 CSoutput.n283 CSoutput.n147 4.5005
R1652 CSoutput.n281 CSoutput.n143 4.5005
R1653 CSoutput.n281 CSoutput.n145 4.5005
R1654 CSoutput.n281 CSoutput.n142 4.5005
R1655 CSoutput.n281 CSoutput.n146 4.5005
R1656 CSoutput.n281 CSoutput.n141 4.5005
R1657 CSoutput.n281 CSoutput.t211 4.5005
R1658 CSoutput.n281 CSoutput.n140 4.5005
R1659 CSoutput.n281 CSoutput.n147 4.5005
R1660 CSoutput.n167 CSoutput.n143 4.5005
R1661 CSoutput.n167 CSoutput.n145 4.5005
R1662 CSoutput.n167 CSoutput.n142 4.5005
R1663 CSoutput.n167 CSoutput.n146 4.5005
R1664 CSoutput.n167 CSoutput.n141 4.5005
R1665 CSoutput.n167 CSoutput.t211 4.5005
R1666 CSoutput.n167 CSoutput.n140 4.5005
R1667 CSoutput.n167 CSoutput.n147 4.5005
R1668 CSoutput.n167 CSoutput.n148 4.5005
R1669 CSoutput.n166 CSoutput.n143 4.5005
R1670 CSoutput.n166 CSoutput.n145 4.5005
R1671 CSoutput.n166 CSoutput.n142 4.5005
R1672 CSoutput.n166 CSoutput.n146 4.5005
R1673 CSoutput.n166 CSoutput.n141 4.5005
R1674 CSoutput.n166 CSoutput.t211 4.5005
R1675 CSoutput.n166 CSoutput.n140 4.5005
R1676 CSoutput.n166 CSoutput.n147 4.5005
R1677 CSoutput.n166 CSoutput.n148 4.5005
R1678 CSoutput.n170 CSoutput.n143 4.5005
R1679 CSoutput.n170 CSoutput.n145 4.5005
R1680 CSoutput.n170 CSoutput.n142 4.5005
R1681 CSoutput.n170 CSoutput.n146 4.5005
R1682 CSoutput.n170 CSoutput.n141 4.5005
R1683 CSoutput.n170 CSoutput.t211 4.5005
R1684 CSoutput.n170 CSoutput.n140 4.5005
R1685 CSoutput.n170 CSoutput.n147 4.5005
R1686 CSoutput.n170 CSoutput.n148 4.5005
R1687 CSoutput.n169 CSoutput.n143 4.5005
R1688 CSoutput.n169 CSoutput.n145 4.5005
R1689 CSoutput.n169 CSoutput.n142 4.5005
R1690 CSoutput.n169 CSoutput.n146 4.5005
R1691 CSoutput.n169 CSoutput.n141 4.5005
R1692 CSoutput.n169 CSoutput.t211 4.5005
R1693 CSoutput.n169 CSoutput.n140 4.5005
R1694 CSoutput.n169 CSoutput.n147 4.5005
R1695 CSoutput.n169 CSoutput.n148 4.5005
R1696 CSoutput.n152 CSoutput.n143 4.5005
R1697 CSoutput.n152 CSoutput.n145 4.5005
R1698 CSoutput.n152 CSoutput.n142 4.5005
R1699 CSoutput.n152 CSoutput.n146 4.5005
R1700 CSoutput.n152 CSoutput.n141 4.5005
R1701 CSoutput.n152 CSoutput.t211 4.5005
R1702 CSoutput.n152 CSoutput.n140 4.5005
R1703 CSoutput.n152 CSoutput.n147 4.5005
R1704 CSoutput.n152 CSoutput.n148 4.5005
R1705 CSoutput.n288 CSoutput.n143 4.5005
R1706 CSoutput.n288 CSoutput.n145 4.5005
R1707 CSoutput.n288 CSoutput.n142 4.5005
R1708 CSoutput.n288 CSoutput.n146 4.5005
R1709 CSoutput.n288 CSoutput.n141 4.5005
R1710 CSoutput.n288 CSoutput.t211 4.5005
R1711 CSoutput.n288 CSoutput.n140 4.5005
R1712 CSoutput.n288 CSoutput.n147 4.5005
R1713 CSoutput.n288 CSoutput.n148 4.5005
R1714 CSoutput.n347 CSoutput.n327 4.10845
R1715 CSoutput.n137 CSoutput.n117 4.10845
R1716 CSoutput.n345 CSoutput.t185 4.06363
R1717 CSoutput.n345 CSoutput.t87 4.06363
R1718 CSoutput.n343 CSoutput.t84 4.06363
R1719 CSoutput.n343 CSoutput.t13 4.06363
R1720 CSoutput.n341 CSoutput.t95 4.06363
R1721 CSoutput.n341 CSoutput.t74 4.06363
R1722 CSoutput.n339 CSoutput.t75 4.06363
R1723 CSoutput.n339 CSoutput.t189 4.06363
R1724 CSoutput.n337 CSoutput.t30 4.06363
R1725 CSoutput.n337 CSoutput.t88 4.06363
R1726 CSoutput.n335 CSoutput.t76 4.06363
R1727 CSoutput.n335 CSoutput.t82 4.06363
R1728 CSoutput.n333 CSoutput.t7 4.06363
R1729 CSoutput.n333 CSoutput.t22 4.06363
R1730 CSoutput.n331 CSoutput.t12 4.06363
R1731 CSoutput.n331 CSoutput.t188 4.06363
R1732 CSoutput.n329 CSoutput.t191 4.06363
R1733 CSoutput.n329 CSoutput.t6 4.06363
R1734 CSoutput.n328 CSoutput.t98 4.06363
R1735 CSoutput.n328 CSoutput.t46 4.06363
R1736 CSoutput.n325 CSoutput.t57 4.06363
R1737 CSoutput.n325 CSoutput.t53 4.06363
R1738 CSoutput.n323 CSoutput.t29 4.06363
R1739 CSoutput.n323 CSoutput.t35 4.06363
R1740 CSoutput.n321 CSoutput.t90 4.06363
R1741 CSoutput.n321 CSoutput.t20 4.06363
R1742 CSoutput.n319 CSoutput.t25 4.06363
R1743 CSoutput.n319 CSoutput.t77 4.06363
R1744 CSoutput.n317 CSoutput.t67 4.06363
R1745 CSoutput.n317 CSoutput.t96 4.06363
R1746 CSoutput.n315 CSoutput.t66 4.06363
R1747 CSoutput.n315 CSoutput.t26 4.06363
R1748 CSoutput.n313 CSoutput.t38 4.06363
R1749 CSoutput.n313 CSoutput.t198 4.06363
R1750 CSoutput.n311 CSoutput.t1 4.06363
R1751 CSoutput.n311 CSoutput.t42 4.06363
R1752 CSoutput.n309 CSoutput.t59 4.06363
R1753 CSoutput.n309 CSoutput.t23 4.06363
R1754 CSoutput.n308 CSoutput.t17 4.06363
R1755 CSoutput.n308 CSoutput.t85 4.06363
R1756 CSoutput.n306 CSoutput.t54 4.06363
R1757 CSoutput.n306 CSoutput.t58 4.06363
R1758 CSoutput.n304 CSoutput.t27 4.06363
R1759 CSoutput.n304 CSoutput.t15 4.06363
R1760 CSoutput.n302 CSoutput.t86 4.06363
R1761 CSoutput.n302 CSoutput.t34 4.06363
R1762 CSoutput.n300 CSoutput.t97 4.06363
R1763 CSoutput.n300 CSoutput.t195 4.06363
R1764 CSoutput.n298 CSoutput.t47 4.06363
R1765 CSoutput.n298 CSoutput.t44 4.06363
R1766 CSoutput.n296 CSoutput.t36 4.06363
R1767 CSoutput.n296 CSoutput.t33 4.06363
R1768 CSoutput.n294 CSoutput.t51 4.06363
R1769 CSoutput.n294 CSoutput.t55 4.06363
R1770 CSoutput.n292 CSoutput.t11 4.06363
R1771 CSoutput.n292 CSoutput.t197 4.06363
R1772 CSoutput.n290 CSoutput.t70 4.06363
R1773 CSoutput.n290 CSoutput.t2 4.06363
R1774 CSoutput.n289 CSoutput.t39 4.06363
R1775 CSoutput.n289 CSoutput.t81 4.06363
R1776 CSoutput.n118 CSoutput.t3 4.06363
R1777 CSoutput.n118 CSoutput.t80 4.06363
R1778 CSoutput.n119 CSoutput.t19 4.06363
R1779 CSoutput.n119 CSoutput.t37 4.06363
R1780 CSoutput.n121 CSoutput.t181 4.06363
R1781 CSoutput.n121 CSoutput.t48 4.06363
R1782 CSoutput.n123 CSoutput.t183 4.06363
R1783 CSoutput.n123 CSoutput.t184 4.06363
R1784 CSoutput.n125 CSoutput.t93 4.06363
R1785 CSoutput.n125 CSoutput.t182 4.06363
R1786 CSoutput.n127 CSoutput.t63 4.06363
R1787 CSoutput.n127 CSoutput.t92 4.06363
R1788 CSoutput.n129 CSoutput.t94 4.06363
R1789 CSoutput.n129 CSoutput.t32 4.06363
R1790 CSoutput.n131 CSoutput.t40 4.06363
R1791 CSoutput.n131 CSoutput.t45 4.06363
R1792 CSoutput.n133 CSoutput.t8 4.06363
R1793 CSoutput.n133 CSoutput.t5 4.06363
R1794 CSoutput.n135 CSoutput.t28 4.06363
R1795 CSoutput.n135 CSoutput.t78 4.06363
R1796 CSoutput.n98 CSoutput.t190 4.06363
R1797 CSoutput.n98 CSoutput.t10 4.06363
R1798 CSoutput.n99 CSoutput.t24 4.06363
R1799 CSoutput.n99 CSoutput.t18 4.06363
R1800 CSoutput.n101 CSoutput.t192 4.06363
R1801 CSoutput.n101 CSoutput.t61 4.06363
R1802 CSoutput.n103 CSoutput.t69 4.06363
R1803 CSoutput.n103 CSoutput.t91 4.06363
R1804 CSoutput.n105 CSoutput.t41 4.06363
R1805 CSoutput.n105 CSoutput.t83 4.06363
R1806 CSoutput.n107 CSoutput.t31 4.06363
R1807 CSoutput.n107 CSoutput.t193 4.06363
R1808 CSoutput.n109 CSoutput.t16 4.06363
R1809 CSoutput.n109 CSoutput.t64 4.06363
R1810 CSoutput.n111 CSoutput.t79 4.06363
R1811 CSoutput.n111 CSoutput.t199 4.06363
R1812 CSoutput.n113 CSoutput.t52 4.06363
R1813 CSoutput.n113 CSoutput.t21 4.06363
R1814 CSoutput.n115 CSoutput.t14 4.06363
R1815 CSoutput.n115 CSoutput.t49 4.06363
R1816 CSoutput.n79 CSoutput.t62 4.06363
R1817 CSoutput.n79 CSoutput.t9 4.06363
R1818 CSoutput.n80 CSoutput.t194 4.06363
R1819 CSoutput.n80 CSoutput.t60 4.06363
R1820 CSoutput.n82 CSoutput.t196 4.06363
R1821 CSoutput.n82 CSoutput.t186 4.06363
R1822 CSoutput.n84 CSoutput.t56 4.06363
R1823 CSoutput.n84 CSoutput.t89 4.06363
R1824 CSoutput.n86 CSoutput.t0 4.06363
R1825 CSoutput.n86 CSoutput.t65 4.06363
R1826 CSoutput.n88 CSoutput.t68 4.06363
R1827 CSoutput.n88 CSoutput.t180 4.06363
R1828 CSoutput.n90 CSoutput.t50 4.06363
R1829 CSoutput.n90 CSoutput.t72 4.06363
R1830 CSoutput.n92 CSoutput.t73 4.06363
R1831 CSoutput.n92 CSoutput.t71 4.06363
R1832 CSoutput.n94 CSoutput.t99 4.06363
R1833 CSoutput.n94 CSoutput.t43 4.06363
R1834 CSoutput.n96 CSoutput.t187 4.06363
R1835 CSoutput.n96 CSoutput.t4 4.06363
R1836 CSoutput.n44 CSoutput.n43 3.79402
R1837 CSoutput.n49 CSoutput.n48 3.79402
R1838 CSoutput.n429 CSoutput.n428 3.57343
R1839 CSoutput.n428 CSoutput.n388 3.42304
R1840 CSoutput.n385 CSoutput.t168 2.82907
R1841 CSoutput.n385 CSoutput.t117 2.82907
R1842 CSoutput.n383 CSoutput.t100 2.82907
R1843 CSoutput.n383 CSoutput.t178 2.82907
R1844 CSoutput.n381 CSoutput.t109 2.82907
R1845 CSoutput.n381 CSoutput.t121 2.82907
R1846 CSoutput.n379 CSoutput.t115 2.82907
R1847 CSoutput.n379 CSoutput.t150 2.82907
R1848 CSoutput.n377 CSoutput.t142 2.82907
R1849 CSoutput.n377 CSoutput.t145 2.82907
R1850 CSoutput.n375 CSoutput.t122 2.82907
R1851 CSoutput.n375 CSoutput.t163 2.82907
R1852 CSoutput.n373 CSoutput.t170 2.82907
R1853 CSoutput.n373 CSoutput.t119 2.82907
R1854 CSoutput.n371 CSoutput.t103 2.82907
R1855 CSoutput.n371 CSoutput.t128 2.82907
R1856 CSoutput.n369 CSoutput.t113 2.82907
R1857 CSoutput.n369 CSoutput.t151 2.82907
R1858 CSoutput.n368 CSoutput.t118 2.82907
R1859 CSoutput.n368 CSoutput.t155 2.82907
R1860 CSoutput.n366 CSoutput.t110 2.82907
R1861 CSoutput.n366 CSoutput.t156 2.82907
R1862 CSoutput.n364 CSoutput.t127 2.82907
R1863 CSoutput.n364 CSoutput.t149 2.82907
R1864 CSoutput.n362 CSoutput.t141 2.82907
R1865 CSoutput.n362 CSoutput.t101 2.82907
R1866 CSoutput.n360 CSoutput.t154 2.82907
R1867 CSoutput.n360 CSoutput.t137 2.82907
R1868 CSoutput.n358 CSoutput.t105 2.82907
R1869 CSoutput.n358 CSoutput.t116 2.82907
R1870 CSoutput.n356 CSoutput.t102 2.82907
R1871 CSoutput.n356 CSoutput.t126 2.82907
R1872 CSoutput.n354 CSoutput.t111 2.82907
R1873 CSoutput.n354 CSoutput.t160 2.82907
R1874 CSoutput.n352 CSoutput.t131 2.82907
R1875 CSoutput.n352 CSoutput.t175 2.82907
R1876 CSoutput.n350 CSoutput.t144 2.82907
R1877 CSoutput.n350 CSoutput.t146 2.82907
R1878 CSoutput.n349 CSoutput.t159 2.82907
R1879 CSoutput.n349 CSoutput.t140 2.82907
R1880 CSoutput.n408 CSoutput.t134 2.82907
R1881 CSoutput.n408 CSoutput.t133 2.82907
R1882 CSoutput.n409 CSoutput.t143 2.82907
R1883 CSoutput.n409 CSoutput.t166 2.82907
R1884 CSoutput.n411 CSoutput.t169 2.82907
R1885 CSoutput.n411 CSoutput.t125 2.82907
R1886 CSoutput.n413 CSoutput.t153 2.82907
R1887 CSoutput.n413 CSoutput.t176 2.82907
R1888 CSoutput.n415 CSoutput.t138 2.82907
R1889 CSoutput.n415 CSoutput.t161 2.82907
R1890 CSoutput.n417 CSoutput.t106 2.82907
R1891 CSoutput.n417 CSoutput.t148 2.82907
R1892 CSoutput.n419 CSoutput.t179 2.82907
R1893 CSoutput.n419 CSoutput.t129 2.82907
R1894 CSoutput.n421 CSoutput.t158 2.82907
R1895 CSoutput.n421 CSoutput.t120 2.82907
R1896 CSoutput.n423 CSoutput.t171 2.82907
R1897 CSoutput.n423 CSoutput.t139 2.82907
R1898 CSoutput.n425 CSoutput.t104 2.82907
R1899 CSoutput.n425 CSoutput.t152 2.82907
R1900 CSoutput.n389 CSoutput.t167 2.82907
R1901 CSoutput.n389 CSoutput.t135 2.82907
R1902 CSoutput.n390 CSoutput.t107 2.82907
R1903 CSoutput.n390 CSoutput.t108 2.82907
R1904 CSoutput.n392 CSoutput.t114 2.82907
R1905 CSoutput.n392 CSoutput.t174 2.82907
R1906 CSoutput.n394 CSoutput.t136 2.82907
R1907 CSoutput.n394 CSoutput.t164 2.82907
R1908 CSoutput.n396 CSoutput.t172 2.82907
R1909 CSoutput.n396 CSoutput.t124 2.82907
R1910 CSoutput.n398 CSoutput.t132 2.82907
R1911 CSoutput.n398 CSoutput.t157 2.82907
R1912 CSoutput.n400 CSoutput.t165 2.82907
R1913 CSoutput.n400 CSoutput.t177 2.82907
R1914 CSoutput.n402 CSoutput.t123 2.82907
R1915 CSoutput.n402 CSoutput.t162 2.82907
R1916 CSoutput.n404 CSoutput.t112 2.82907
R1917 CSoutput.n404 CSoutput.t173 2.82907
R1918 CSoutput.n406 CSoutput.t130 2.82907
R1919 CSoutput.n406 CSoutput.t147 2.82907
R1920 CSoutput.n348 CSoutput.n138 2.78353
R1921 CSoutput.n75 CSoutput.n1 2.45513
R1922 CSoutput.n229 CSoutput.n227 2.251
R1923 CSoutput.n229 CSoutput.n226 2.251
R1924 CSoutput.n229 CSoutput.n225 2.251
R1925 CSoutput.n229 CSoutput.n224 2.251
R1926 CSoutput.n198 CSoutput.n197 2.251
R1927 CSoutput.n198 CSoutput.n196 2.251
R1928 CSoutput.n198 CSoutput.n195 2.251
R1929 CSoutput.n198 CSoutput.n194 2.251
R1930 CSoutput.n271 CSoutput.n270 2.251
R1931 CSoutput.n236 CSoutput.n234 2.251
R1932 CSoutput.n236 CSoutput.n233 2.251
R1933 CSoutput.n236 CSoutput.n232 2.251
R1934 CSoutput.n254 CSoutput.n236 2.251
R1935 CSoutput.n242 CSoutput.n241 2.251
R1936 CSoutput.n242 CSoutput.n240 2.251
R1937 CSoutput.n242 CSoutput.n239 2.251
R1938 CSoutput.n242 CSoutput.n238 2.251
R1939 CSoutput.n268 CSoutput.n208 2.251
R1940 CSoutput.n263 CSoutput.n261 2.251
R1941 CSoutput.n263 CSoutput.n260 2.251
R1942 CSoutput.n263 CSoutput.n259 2.251
R1943 CSoutput.n263 CSoutput.n258 2.251
R1944 CSoutput.n164 CSoutput.n163 2.251
R1945 CSoutput.n164 CSoutput.n162 2.251
R1946 CSoutput.n164 CSoutput.n161 2.251
R1947 CSoutput.n164 CSoutput.n160 2.251
R1948 CSoutput.n281 CSoutput.n280 2.251
R1949 CSoutput.n198 CSoutput.n178 2.2505
R1950 CSoutput.n193 CSoutput.n178 2.2505
R1951 CSoutput.n191 CSoutput.n178 2.2505
R1952 CSoutput.n190 CSoutput.n178 2.2505
R1953 CSoutput.n275 CSoutput.n178 2.2505
R1954 CSoutput.n273 CSoutput.n178 2.2505
R1955 CSoutput.n271 CSoutput.n178 2.2505
R1956 CSoutput.n201 CSoutput.n178 2.2505
R1957 CSoutput.n200 CSoutput.n178 2.2505
R1958 CSoutput.n204 CSoutput.n178 2.2505
R1959 CSoutput.n203 CSoutput.n178 2.2505
R1960 CSoutput.n186 CSoutput.n178 2.2505
R1961 CSoutput.n278 CSoutput.n178 2.2505
R1962 CSoutput.n278 CSoutput.n277 2.2505
R1963 CSoutput.n242 CSoutput.n213 2.2505
R1964 CSoutput.n223 CSoutput.n213 2.2505
R1965 CSoutput.n244 CSoutput.n213 2.2505
R1966 CSoutput.n222 CSoutput.n213 2.2505
R1967 CSoutput.n246 CSoutput.n213 2.2505
R1968 CSoutput.n213 CSoutput.n207 2.2505
R1969 CSoutput.n268 CSoutput.n213 2.2505
R1970 CSoutput.n266 CSoutput.n213 2.2505
R1971 CSoutput.n248 CSoutput.n213 2.2505
R1972 CSoutput.n220 CSoutput.n213 2.2505
R1973 CSoutput.n250 CSoutput.n213 2.2505
R1974 CSoutput.n219 CSoutput.n213 2.2505
R1975 CSoutput.n264 CSoutput.n213 2.2505
R1976 CSoutput.n264 CSoutput.n217 2.2505
R1977 CSoutput.n164 CSoutput.n144 2.2505
R1978 CSoutput.n159 CSoutput.n144 2.2505
R1979 CSoutput.n157 CSoutput.n144 2.2505
R1980 CSoutput.n156 CSoutput.n144 2.2505
R1981 CSoutput.n285 CSoutput.n144 2.2505
R1982 CSoutput.n283 CSoutput.n144 2.2505
R1983 CSoutput.n281 CSoutput.n144 2.2505
R1984 CSoutput.n167 CSoutput.n144 2.2505
R1985 CSoutput.n166 CSoutput.n144 2.2505
R1986 CSoutput.n170 CSoutput.n144 2.2505
R1987 CSoutput.n169 CSoutput.n144 2.2505
R1988 CSoutput.n152 CSoutput.n144 2.2505
R1989 CSoutput.n288 CSoutput.n144 2.2505
R1990 CSoutput.n288 CSoutput.n287 2.2505
R1991 CSoutput.n206 CSoutput.n199 2.25024
R1992 CSoutput.n206 CSoutput.n192 2.25024
R1993 CSoutput.n274 CSoutput.n206 2.25024
R1994 CSoutput.n206 CSoutput.n202 2.25024
R1995 CSoutput.n206 CSoutput.n205 2.25024
R1996 CSoutput.n206 CSoutput.n173 2.25024
R1997 CSoutput.n256 CSoutput.n253 2.25024
R1998 CSoutput.n256 CSoutput.n252 2.25024
R1999 CSoutput.n256 CSoutput.n251 2.25024
R2000 CSoutput.n256 CSoutput.n218 2.25024
R2001 CSoutput.n256 CSoutput.n255 2.25024
R2002 CSoutput.n257 CSoutput.n256 2.25024
R2003 CSoutput.n172 CSoutput.n165 2.25024
R2004 CSoutput.n172 CSoutput.n158 2.25024
R2005 CSoutput.n284 CSoutput.n172 2.25024
R2006 CSoutput.n172 CSoutput.n168 2.25024
R2007 CSoutput.n172 CSoutput.n171 2.25024
R2008 CSoutput.n172 CSoutput.n139 2.25024
R2009 CSoutput.n273 CSoutput.n183 1.50111
R2010 CSoutput.n221 CSoutput.n207 1.50111
R2011 CSoutput.n283 CSoutput.n149 1.50111
R2012 CSoutput.n229 CSoutput.n228 1.501
R2013 CSoutput.n236 CSoutput.n235 1.501
R2014 CSoutput.n263 CSoutput.n262 1.501
R2015 CSoutput.n277 CSoutput.n188 1.12536
R2016 CSoutput.n277 CSoutput.n189 1.12536
R2017 CSoutput.n277 CSoutput.n276 1.12536
R2018 CSoutput.n237 CSoutput.n217 1.12536
R2019 CSoutput.n243 CSoutput.n217 1.12536
R2020 CSoutput.n245 CSoutput.n217 1.12536
R2021 CSoutput.n287 CSoutput.n154 1.12536
R2022 CSoutput.n287 CSoutput.n155 1.12536
R2023 CSoutput.n287 CSoutput.n286 1.12536
R2024 CSoutput.n277 CSoutput.n184 1.12536
R2025 CSoutput.n277 CSoutput.n185 1.12536
R2026 CSoutput.n277 CSoutput.n187 1.12536
R2027 CSoutput.n267 CSoutput.n217 1.12536
R2028 CSoutput.n247 CSoutput.n217 1.12536
R2029 CSoutput.n249 CSoutput.n217 1.12536
R2030 CSoutput.n287 CSoutput.n150 1.12536
R2031 CSoutput.n287 CSoutput.n151 1.12536
R2032 CSoutput.n287 CSoutput.n153 1.12536
R2033 CSoutput.n31 CSoutput.n30 0.669944
R2034 CSoutput.n62 CSoutput.n61 0.669944
R2035 CSoutput.n372 CSoutput.n370 0.573776
R2036 CSoutput.n374 CSoutput.n372 0.573776
R2037 CSoutput.n376 CSoutput.n374 0.573776
R2038 CSoutput.n378 CSoutput.n376 0.573776
R2039 CSoutput.n380 CSoutput.n378 0.573776
R2040 CSoutput.n382 CSoutput.n380 0.573776
R2041 CSoutput.n384 CSoutput.n382 0.573776
R2042 CSoutput.n386 CSoutput.n384 0.573776
R2043 CSoutput.n353 CSoutput.n351 0.573776
R2044 CSoutput.n355 CSoutput.n353 0.573776
R2045 CSoutput.n357 CSoutput.n355 0.573776
R2046 CSoutput.n359 CSoutput.n357 0.573776
R2047 CSoutput.n361 CSoutput.n359 0.573776
R2048 CSoutput.n363 CSoutput.n361 0.573776
R2049 CSoutput.n365 CSoutput.n363 0.573776
R2050 CSoutput.n367 CSoutput.n365 0.573776
R2051 CSoutput.n426 CSoutput.n424 0.573776
R2052 CSoutput.n424 CSoutput.n422 0.573776
R2053 CSoutput.n422 CSoutput.n420 0.573776
R2054 CSoutput.n420 CSoutput.n418 0.573776
R2055 CSoutput.n418 CSoutput.n416 0.573776
R2056 CSoutput.n416 CSoutput.n414 0.573776
R2057 CSoutput.n414 CSoutput.n412 0.573776
R2058 CSoutput.n412 CSoutput.n410 0.573776
R2059 CSoutput.n407 CSoutput.n405 0.573776
R2060 CSoutput.n405 CSoutput.n403 0.573776
R2061 CSoutput.n403 CSoutput.n401 0.573776
R2062 CSoutput.n401 CSoutput.n399 0.573776
R2063 CSoutput.n399 CSoutput.n397 0.573776
R2064 CSoutput.n397 CSoutput.n395 0.573776
R2065 CSoutput.n395 CSoutput.n393 0.573776
R2066 CSoutput.n393 CSoutput.n391 0.573776
R2067 CSoutput.n429 CSoutput.n288 0.53442
R2068 CSoutput.n332 CSoutput.n330 0.358259
R2069 CSoutput.n334 CSoutput.n332 0.358259
R2070 CSoutput.n336 CSoutput.n334 0.358259
R2071 CSoutput.n338 CSoutput.n336 0.358259
R2072 CSoutput.n340 CSoutput.n338 0.358259
R2073 CSoutput.n342 CSoutput.n340 0.358259
R2074 CSoutput.n344 CSoutput.n342 0.358259
R2075 CSoutput.n346 CSoutput.n344 0.358259
R2076 CSoutput.n312 CSoutput.n310 0.358259
R2077 CSoutput.n314 CSoutput.n312 0.358259
R2078 CSoutput.n316 CSoutput.n314 0.358259
R2079 CSoutput.n318 CSoutput.n316 0.358259
R2080 CSoutput.n320 CSoutput.n318 0.358259
R2081 CSoutput.n322 CSoutput.n320 0.358259
R2082 CSoutput.n324 CSoutput.n322 0.358259
R2083 CSoutput.n326 CSoutput.n324 0.358259
R2084 CSoutput.n293 CSoutput.n291 0.358259
R2085 CSoutput.n295 CSoutput.n293 0.358259
R2086 CSoutput.n297 CSoutput.n295 0.358259
R2087 CSoutput.n299 CSoutput.n297 0.358259
R2088 CSoutput.n301 CSoutput.n299 0.358259
R2089 CSoutput.n303 CSoutput.n301 0.358259
R2090 CSoutput.n305 CSoutput.n303 0.358259
R2091 CSoutput.n307 CSoutput.n305 0.358259
R2092 CSoutput.n136 CSoutput.n134 0.358259
R2093 CSoutput.n134 CSoutput.n132 0.358259
R2094 CSoutput.n132 CSoutput.n130 0.358259
R2095 CSoutput.n130 CSoutput.n128 0.358259
R2096 CSoutput.n128 CSoutput.n126 0.358259
R2097 CSoutput.n126 CSoutput.n124 0.358259
R2098 CSoutput.n124 CSoutput.n122 0.358259
R2099 CSoutput.n122 CSoutput.n120 0.358259
R2100 CSoutput.n116 CSoutput.n114 0.358259
R2101 CSoutput.n114 CSoutput.n112 0.358259
R2102 CSoutput.n112 CSoutput.n110 0.358259
R2103 CSoutput.n110 CSoutput.n108 0.358259
R2104 CSoutput.n108 CSoutput.n106 0.358259
R2105 CSoutput.n106 CSoutput.n104 0.358259
R2106 CSoutput.n104 CSoutput.n102 0.358259
R2107 CSoutput.n102 CSoutput.n100 0.358259
R2108 CSoutput.n97 CSoutput.n95 0.358259
R2109 CSoutput.n95 CSoutput.n93 0.358259
R2110 CSoutput.n93 CSoutput.n91 0.358259
R2111 CSoutput.n91 CSoutput.n89 0.358259
R2112 CSoutput.n89 CSoutput.n87 0.358259
R2113 CSoutput.n87 CSoutput.n85 0.358259
R2114 CSoutput.n85 CSoutput.n83 0.358259
R2115 CSoutput.n83 CSoutput.n81 0.358259
R2116 CSoutput.n21 CSoutput.n20 0.169105
R2117 CSoutput.n21 CSoutput.n16 0.169105
R2118 CSoutput.n26 CSoutput.n16 0.169105
R2119 CSoutput.n27 CSoutput.n26 0.169105
R2120 CSoutput.n27 CSoutput.n14 0.169105
R2121 CSoutput.n32 CSoutput.n14 0.169105
R2122 CSoutput.n33 CSoutput.n32 0.169105
R2123 CSoutput.n34 CSoutput.n33 0.169105
R2124 CSoutput.n34 CSoutput.n12 0.169105
R2125 CSoutput.n39 CSoutput.n12 0.169105
R2126 CSoutput.n40 CSoutput.n39 0.169105
R2127 CSoutput.n40 CSoutput.n10 0.169105
R2128 CSoutput.n45 CSoutput.n10 0.169105
R2129 CSoutput.n46 CSoutput.n45 0.169105
R2130 CSoutput.n47 CSoutput.n46 0.169105
R2131 CSoutput.n47 CSoutput.n8 0.169105
R2132 CSoutput.n52 CSoutput.n8 0.169105
R2133 CSoutput.n53 CSoutput.n52 0.169105
R2134 CSoutput.n53 CSoutput.n6 0.169105
R2135 CSoutput.n58 CSoutput.n6 0.169105
R2136 CSoutput.n59 CSoutput.n58 0.169105
R2137 CSoutput.n60 CSoutput.n59 0.169105
R2138 CSoutput.n60 CSoutput.n4 0.169105
R2139 CSoutput.n66 CSoutput.n4 0.169105
R2140 CSoutput.n67 CSoutput.n66 0.169105
R2141 CSoutput.n68 CSoutput.n67 0.169105
R2142 CSoutput.n68 CSoutput.n2 0.169105
R2143 CSoutput.n73 CSoutput.n2 0.169105
R2144 CSoutput.n74 CSoutput.n73 0.169105
R2145 CSoutput.n74 CSoutput.n0 0.169105
R2146 CSoutput.n78 CSoutput.n0 0.169105
R2147 CSoutput.n231 CSoutput.n230 0.0910737
R2148 CSoutput.n282 CSoutput.n279 0.0723685
R2149 CSoutput.n236 CSoutput.n231 0.0522944
R2150 CSoutput.n279 CSoutput.n278 0.0499135
R2151 CSoutput.n230 CSoutput.n229 0.0499135
R2152 CSoutput.n264 CSoutput.n263 0.0464294
R2153 CSoutput.n272 CSoutput.n269 0.0391444
R2154 CSoutput.n231 CSoutput.t200 0.023435
R2155 CSoutput.n279 CSoutput.t204 0.02262
R2156 CSoutput.n230 CSoutput.t207 0.02262
R2157 CSoutput CSoutput.n429 0.0052
R2158 CSoutput.n201 CSoutput.n184 0.00365111
R2159 CSoutput.n204 CSoutput.n185 0.00365111
R2160 CSoutput.n187 CSoutput.n186 0.00365111
R2161 CSoutput.n229 CSoutput.n188 0.00365111
R2162 CSoutput.n193 CSoutput.n189 0.00365111
R2163 CSoutput.n276 CSoutput.n190 0.00365111
R2164 CSoutput.n267 CSoutput.n266 0.00365111
R2165 CSoutput.n247 CSoutput.n220 0.00365111
R2166 CSoutput.n249 CSoutput.n219 0.00365111
R2167 CSoutput.n237 CSoutput.n236 0.00365111
R2168 CSoutput.n243 CSoutput.n223 0.00365111
R2169 CSoutput.n245 CSoutput.n222 0.00365111
R2170 CSoutput.n167 CSoutput.n150 0.00365111
R2171 CSoutput.n170 CSoutput.n151 0.00365111
R2172 CSoutput.n153 CSoutput.n152 0.00365111
R2173 CSoutput.n263 CSoutput.n154 0.00365111
R2174 CSoutput.n159 CSoutput.n155 0.00365111
R2175 CSoutput.n286 CSoutput.n156 0.00365111
R2176 CSoutput.n198 CSoutput.n188 0.00340054
R2177 CSoutput.n191 CSoutput.n189 0.00340054
R2178 CSoutput.n276 CSoutput.n275 0.00340054
R2179 CSoutput.n271 CSoutput.n184 0.00340054
R2180 CSoutput.n200 CSoutput.n185 0.00340054
R2181 CSoutput.n203 CSoutput.n187 0.00340054
R2182 CSoutput.n242 CSoutput.n237 0.00340054
R2183 CSoutput.n244 CSoutput.n243 0.00340054
R2184 CSoutput.n246 CSoutput.n245 0.00340054
R2185 CSoutput.n268 CSoutput.n267 0.00340054
R2186 CSoutput.n248 CSoutput.n247 0.00340054
R2187 CSoutput.n250 CSoutput.n249 0.00340054
R2188 CSoutput.n164 CSoutput.n154 0.00340054
R2189 CSoutput.n157 CSoutput.n155 0.00340054
R2190 CSoutput.n286 CSoutput.n285 0.00340054
R2191 CSoutput.n281 CSoutput.n150 0.00340054
R2192 CSoutput.n166 CSoutput.n151 0.00340054
R2193 CSoutput.n169 CSoutput.n153 0.00340054
R2194 CSoutput.n199 CSoutput.n193 0.00252698
R2195 CSoutput.n192 CSoutput.n190 0.00252698
R2196 CSoutput.n274 CSoutput.n273 0.00252698
R2197 CSoutput.n202 CSoutput.n200 0.00252698
R2198 CSoutput.n205 CSoutput.n203 0.00252698
R2199 CSoutput.n278 CSoutput.n173 0.00252698
R2200 CSoutput.n199 CSoutput.n198 0.00252698
R2201 CSoutput.n192 CSoutput.n191 0.00252698
R2202 CSoutput.n275 CSoutput.n274 0.00252698
R2203 CSoutput.n202 CSoutput.n201 0.00252698
R2204 CSoutput.n205 CSoutput.n204 0.00252698
R2205 CSoutput.n186 CSoutput.n173 0.00252698
R2206 CSoutput.n253 CSoutput.n223 0.00252698
R2207 CSoutput.n252 CSoutput.n222 0.00252698
R2208 CSoutput.n251 CSoutput.n207 0.00252698
R2209 CSoutput.n248 CSoutput.n218 0.00252698
R2210 CSoutput.n255 CSoutput.n250 0.00252698
R2211 CSoutput.n264 CSoutput.n257 0.00252698
R2212 CSoutput.n253 CSoutput.n242 0.00252698
R2213 CSoutput.n252 CSoutput.n244 0.00252698
R2214 CSoutput.n251 CSoutput.n246 0.00252698
R2215 CSoutput.n266 CSoutput.n218 0.00252698
R2216 CSoutput.n255 CSoutput.n220 0.00252698
R2217 CSoutput.n257 CSoutput.n219 0.00252698
R2218 CSoutput.n165 CSoutput.n159 0.00252698
R2219 CSoutput.n158 CSoutput.n156 0.00252698
R2220 CSoutput.n284 CSoutput.n283 0.00252698
R2221 CSoutput.n168 CSoutput.n166 0.00252698
R2222 CSoutput.n171 CSoutput.n169 0.00252698
R2223 CSoutput.n288 CSoutput.n139 0.00252698
R2224 CSoutput.n165 CSoutput.n164 0.00252698
R2225 CSoutput.n158 CSoutput.n157 0.00252698
R2226 CSoutput.n285 CSoutput.n284 0.00252698
R2227 CSoutput.n168 CSoutput.n167 0.00252698
R2228 CSoutput.n171 CSoutput.n170 0.00252698
R2229 CSoutput.n152 CSoutput.n139 0.00252698
R2230 CSoutput.n273 CSoutput.n272 0.0020275
R2231 CSoutput.n272 CSoutput.n271 0.0020275
R2232 CSoutput.n269 CSoutput.n207 0.0020275
R2233 CSoutput.n269 CSoutput.n268 0.0020275
R2234 CSoutput.n283 CSoutput.n282 0.0020275
R2235 CSoutput.n282 CSoutput.n281 0.0020275
R2236 CSoutput.n183 CSoutput.n182 0.00166668
R2237 CSoutput.n265 CSoutput.n221 0.00166668
R2238 CSoutput.n149 CSoutput.n148 0.00166668
R2239 CSoutput.n287 CSoutput.n149 0.00133328
R2240 CSoutput.n221 CSoutput.n217 0.00133328
R2241 CSoutput.n277 CSoutput.n183 0.00133328
R2242 CSoutput.n280 CSoutput.n172 0.001
R2243 CSoutput.n258 CSoutput.n172 0.001
R2244 CSoutput.n160 CSoutput.n140 0.001
R2245 CSoutput.n259 CSoutput.n140 0.001
R2246 CSoutput.n161 CSoutput.n141 0.001
R2247 CSoutput.n260 CSoutput.n141 0.001
R2248 CSoutput.n162 CSoutput.n142 0.001
R2249 CSoutput.n261 CSoutput.n142 0.001
R2250 CSoutput.n163 CSoutput.n143 0.001
R2251 CSoutput.n262 CSoutput.n143 0.001
R2252 CSoutput.n256 CSoutput.n208 0.001
R2253 CSoutput.n256 CSoutput.n254 0.001
R2254 CSoutput.n238 CSoutput.n209 0.001
R2255 CSoutput.n232 CSoutput.n209 0.001
R2256 CSoutput.n239 CSoutput.n210 0.001
R2257 CSoutput.n233 CSoutput.n210 0.001
R2258 CSoutput.n240 CSoutput.n211 0.001
R2259 CSoutput.n234 CSoutput.n211 0.001
R2260 CSoutput.n241 CSoutput.n212 0.001
R2261 CSoutput.n235 CSoutput.n212 0.001
R2262 CSoutput.n270 CSoutput.n206 0.001
R2263 CSoutput.n224 CSoutput.n206 0.001
R2264 CSoutput.n194 CSoutput.n174 0.001
R2265 CSoutput.n225 CSoutput.n174 0.001
R2266 CSoutput.n195 CSoutput.n175 0.001
R2267 CSoutput.n226 CSoutput.n175 0.001
R2268 CSoutput.n196 CSoutput.n176 0.001
R2269 CSoutput.n227 CSoutput.n176 0.001
R2270 CSoutput.n197 CSoutput.n177 0.001
R2271 CSoutput.n228 CSoutput.n177 0.001
R2272 CSoutput.n228 CSoutput.n178 0.001
R2273 CSoutput.n227 CSoutput.n179 0.001
R2274 CSoutput.n226 CSoutput.n180 0.001
R2275 CSoutput.n225 CSoutput.t220 0.001
R2276 CSoutput.n224 CSoutput.n181 0.001
R2277 CSoutput.n197 CSoutput.n179 0.001
R2278 CSoutput.n196 CSoutput.n180 0.001
R2279 CSoutput.n195 CSoutput.t220 0.001
R2280 CSoutput.n194 CSoutput.n181 0.001
R2281 CSoutput.n270 CSoutput.n182 0.001
R2282 CSoutput.n235 CSoutput.n213 0.001
R2283 CSoutput.n234 CSoutput.n214 0.001
R2284 CSoutput.n233 CSoutput.n215 0.001
R2285 CSoutput.n232 CSoutput.t214 0.001
R2286 CSoutput.n254 CSoutput.n216 0.001
R2287 CSoutput.n241 CSoutput.n214 0.001
R2288 CSoutput.n240 CSoutput.n215 0.001
R2289 CSoutput.n239 CSoutput.t214 0.001
R2290 CSoutput.n238 CSoutput.n216 0.001
R2291 CSoutput.n265 CSoutput.n208 0.001
R2292 CSoutput.n262 CSoutput.n144 0.001
R2293 CSoutput.n261 CSoutput.n145 0.001
R2294 CSoutput.n260 CSoutput.n146 0.001
R2295 CSoutput.n259 CSoutput.t211 0.001
R2296 CSoutput.n258 CSoutput.n147 0.001
R2297 CSoutput.n163 CSoutput.n145 0.001
R2298 CSoutput.n162 CSoutput.n146 0.001
R2299 CSoutput.n161 CSoutput.t211 0.001
R2300 CSoutput.n160 CSoutput.n147 0.001
R2301 CSoutput.n280 CSoutput.n148 0.001
R2302 gnd.n7153 gnd.n520 1257.24
R2303 gnd.n6511 gnd.n5107 939.716
R2304 gnd.n3229 gnd.n2564 771.183
R2305 gnd.n4626 gnd.n1611 771.183
R2306 gnd.n3233 gnd.n2561 771.183
R2307 gnd.n1992 gnd.n1613 771.183
R2308 gnd.n6405 gnd.n998 766.379
R2309 gnd.n6427 gnd.n6426 766.379
R2310 gnd.n5627 gnd.n5526 766.379
R2311 gnd.n5625 gnd.n5528 766.379
R2312 gnd.n6513 gnd.n995 756.769
R2313 gnd.n5134 gnd.n997 756.769
R2314 gnd.n5759 gnd.n5488 756.769
R2315 gnd.n5745 gnd.n5477 756.769
R2316 gnd.n7510 gnd.n125 751.963
R2317 gnd.n7668 gnd.n7667 751.963
R2318 gnd.n4277 gnd.n4276 751.963
R2319 gnd.n1882 gnd.n1881 751.963
R2320 gnd.n1413 gnd.n1401 751.963
R2321 gnd.n3331 gnd.n3330 751.963
R2322 gnd.n2913 gnd.n1039 751.963
R2323 gnd.n2975 gnd.n2914 751.963
R2324 gnd.n7665 gnd.n127 732.745
R2325 gnd.n195 gnd.n123 732.745
R2326 gnd.n2174 gnd.n2172 732.745
R2327 gnd.n2098 gnd.n1638 732.745
R2328 gnd.n4830 gnd.n1406 732.745
R2329 gnd.n3328 gnd.n2624 732.745
R2330 gnd.n5029 gnd.n5028 732.745
R2331 gnd.n5105 gnd.n1043 732.745
R2332 gnd.n6700 gnd.n795 670.282
R2333 gnd.n7154 gnd.n521 670.282
R2334 gnd.n7371 gnd.n395 670.282
R2335 gnd.n2755 gnd.n2752 670.282
R2336 gnd.n6700 gnd.n6699 585
R2337 gnd.n6701 gnd.n6700 585
R2338 gnd.n6698 gnd.n797 585
R2339 gnd.n797 gnd.n796 585
R2340 gnd.n6697 gnd.n6696 585
R2341 gnd.n6696 gnd.n6695 585
R2342 gnd.n802 gnd.n801 585
R2343 gnd.n6694 gnd.n802 585
R2344 gnd.n6692 gnd.n6691 585
R2345 gnd.n6693 gnd.n6692 585
R2346 gnd.n6690 gnd.n804 585
R2347 gnd.n804 gnd.n803 585
R2348 gnd.n6689 gnd.n6688 585
R2349 gnd.n6688 gnd.n6687 585
R2350 gnd.n810 gnd.n809 585
R2351 gnd.n6686 gnd.n810 585
R2352 gnd.n6684 gnd.n6683 585
R2353 gnd.n6685 gnd.n6684 585
R2354 gnd.n6682 gnd.n812 585
R2355 gnd.n812 gnd.n811 585
R2356 gnd.n6681 gnd.n6680 585
R2357 gnd.n6680 gnd.n6679 585
R2358 gnd.n818 gnd.n817 585
R2359 gnd.n6678 gnd.n818 585
R2360 gnd.n6676 gnd.n6675 585
R2361 gnd.n6677 gnd.n6676 585
R2362 gnd.n6674 gnd.n820 585
R2363 gnd.n820 gnd.n819 585
R2364 gnd.n6673 gnd.n6672 585
R2365 gnd.n6672 gnd.n6671 585
R2366 gnd.n826 gnd.n825 585
R2367 gnd.n6670 gnd.n826 585
R2368 gnd.n6668 gnd.n6667 585
R2369 gnd.n6669 gnd.n6668 585
R2370 gnd.n6666 gnd.n828 585
R2371 gnd.n828 gnd.n827 585
R2372 gnd.n6665 gnd.n6664 585
R2373 gnd.n6664 gnd.n6663 585
R2374 gnd.n834 gnd.n833 585
R2375 gnd.n6662 gnd.n834 585
R2376 gnd.n6660 gnd.n6659 585
R2377 gnd.n6661 gnd.n6660 585
R2378 gnd.n6658 gnd.n836 585
R2379 gnd.n836 gnd.n835 585
R2380 gnd.n6657 gnd.n6656 585
R2381 gnd.n6656 gnd.n6655 585
R2382 gnd.n842 gnd.n841 585
R2383 gnd.n6654 gnd.n842 585
R2384 gnd.n6652 gnd.n6651 585
R2385 gnd.n6653 gnd.n6652 585
R2386 gnd.n6650 gnd.n844 585
R2387 gnd.n844 gnd.n843 585
R2388 gnd.n6649 gnd.n6648 585
R2389 gnd.n6648 gnd.n6647 585
R2390 gnd.n850 gnd.n849 585
R2391 gnd.n6646 gnd.n850 585
R2392 gnd.n6644 gnd.n6643 585
R2393 gnd.n6645 gnd.n6644 585
R2394 gnd.n6642 gnd.n852 585
R2395 gnd.n852 gnd.n851 585
R2396 gnd.n6641 gnd.n6640 585
R2397 gnd.n6640 gnd.n6639 585
R2398 gnd.n858 gnd.n857 585
R2399 gnd.n6638 gnd.n858 585
R2400 gnd.n6636 gnd.n6635 585
R2401 gnd.n6637 gnd.n6636 585
R2402 gnd.n6634 gnd.n860 585
R2403 gnd.n860 gnd.n859 585
R2404 gnd.n6633 gnd.n6632 585
R2405 gnd.n6632 gnd.n6631 585
R2406 gnd.n866 gnd.n865 585
R2407 gnd.n6630 gnd.n866 585
R2408 gnd.n6628 gnd.n6627 585
R2409 gnd.n6629 gnd.n6628 585
R2410 gnd.n6626 gnd.n868 585
R2411 gnd.n868 gnd.n867 585
R2412 gnd.n6625 gnd.n6624 585
R2413 gnd.n6624 gnd.n6623 585
R2414 gnd.n874 gnd.n873 585
R2415 gnd.n6622 gnd.n874 585
R2416 gnd.n6620 gnd.n6619 585
R2417 gnd.n6621 gnd.n6620 585
R2418 gnd.n6618 gnd.n876 585
R2419 gnd.n876 gnd.n875 585
R2420 gnd.n6617 gnd.n6616 585
R2421 gnd.n6616 gnd.n6615 585
R2422 gnd.n882 gnd.n881 585
R2423 gnd.n6614 gnd.n882 585
R2424 gnd.n6612 gnd.n6611 585
R2425 gnd.n6613 gnd.n6612 585
R2426 gnd.n6610 gnd.n884 585
R2427 gnd.n884 gnd.n883 585
R2428 gnd.n6609 gnd.n6608 585
R2429 gnd.n6608 gnd.n6607 585
R2430 gnd.n890 gnd.n889 585
R2431 gnd.n6606 gnd.n890 585
R2432 gnd.n6604 gnd.n6603 585
R2433 gnd.n6605 gnd.n6604 585
R2434 gnd.n6602 gnd.n892 585
R2435 gnd.n892 gnd.n891 585
R2436 gnd.n6601 gnd.n6600 585
R2437 gnd.n6600 gnd.n6599 585
R2438 gnd.n898 gnd.n897 585
R2439 gnd.n6598 gnd.n898 585
R2440 gnd.n6596 gnd.n6595 585
R2441 gnd.n6597 gnd.n6596 585
R2442 gnd.n6594 gnd.n900 585
R2443 gnd.n900 gnd.n899 585
R2444 gnd.n6593 gnd.n6592 585
R2445 gnd.n6592 gnd.n6591 585
R2446 gnd.n906 gnd.n905 585
R2447 gnd.n6590 gnd.n906 585
R2448 gnd.n6588 gnd.n6587 585
R2449 gnd.n6589 gnd.n6588 585
R2450 gnd.n6586 gnd.n908 585
R2451 gnd.n908 gnd.n907 585
R2452 gnd.n6585 gnd.n6584 585
R2453 gnd.n6584 gnd.n6583 585
R2454 gnd.n914 gnd.n913 585
R2455 gnd.n6582 gnd.n914 585
R2456 gnd.n6580 gnd.n6579 585
R2457 gnd.n6581 gnd.n6580 585
R2458 gnd.n6578 gnd.n916 585
R2459 gnd.n916 gnd.n915 585
R2460 gnd.n6577 gnd.n6576 585
R2461 gnd.n6576 gnd.n6575 585
R2462 gnd.n922 gnd.n921 585
R2463 gnd.n6574 gnd.n922 585
R2464 gnd.n6572 gnd.n6571 585
R2465 gnd.n6573 gnd.n6572 585
R2466 gnd.n6570 gnd.n924 585
R2467 gnd.n924 gnd.n923 585
R2468 gnd.n6569 gnd.n6568 585
R2469 gnd.n6568 gnd.n6567 585
R2470 gnd.n930 gnd.n929 585
R2471 gnd.n6566 gnd.n930 585
R2472 gnd.n6564 gnd.n6563 585
R2473 gnd.n6565 gnd.n6564 585
R2474 gnd.n6562 gnd.n932 585
R2475 gnd.n932 gnd.n931 585
R2476 gnd.n6561 gnd.n6560 585
R2477 gnd.n6560 gnd.n6559 585
R2478 gnd.n938 gnd.n937 585
R2479 gnd.n6558 gnd.n938 585
R2480 gnd.n6556 gnd.n6555 585
R2481 gnd.n6557 gnd.n6556 585
R2482 gnd.n6554 gnd.n940 585
R2483 gnd.n940 gnd.n939 585
R2484 gnd.n6553 gnd.n6552 585
R2485 gnd.n6552 gnd.n6551 585
R2486 gnd.n946 gnd.n945 585
R2487 gnd.n6550 gnd.n946 585
R2488 gnd.n6548 gnd.n6547 585
R2489 gnd.n6549 gnd.n6548 585
R2490 gnd.n6546 gnd.n948 585
R2491 gnd.n948 gnd.n947 585
R2492 gnd.n6545 gnd.n6544 585
R2493 gnd.n6544 gnd.n6543 585
R2494 gnd.n954 gnd.n953 585
R2495 gnd.n6542 gnd.n954 585
R2496 gnd.n6540 gnd.n6539 585
R2497 gnd.n6541 gnd.n6540 585
R2498 gnd.n6538 gnd.n956 585
R2499 gnd.n956 gnd.n955 585
R2500 gnd.n6537 gnd.n6536 585
R2501 gnd.n6536 gnd.n6535 585
R2502 gnd.n962 gnd.n961 585
R2503 gnd.n6534 gnd.n962 585
R2504 gnd.n795 gnd.n794 585
R2505 gnd.n6702 gnd.n795 585
R2506 gnd.n6705 gnd.n6704 585
R2507 gnd.n6704 gnd.n6703 585
R2508 gnd.n792 gnd.n791 585
R2509 gnd.n791 gnd.n790 585
R2510 gnd.n6710 gnd.n6709 585
R2511 gnd.n6711 gnd.n6710 585
R2512 gnd.n789 gnd.n788 585
R2513 gnd.n6712 gnd.n789 585
R2514 gnd.n6715 gnd.n6714 585
R2515 gnd.n6714 gnd.n6713 585
R2516 gnd.n786 gnd.n785 585
R2517 gnd.n785 gnd.n784 585
R2518 gnd.n6720 gnd.n6719 585
R2519 gnd.n6721 gnd.n6720 585
R2520 gnd.n783 gnd.n782 585
R2521 gnd.n6722 gnd.n783 585
R2522 gnd.n6725 gnd.n6724 585
R2523 gnd.n6724 gnd.n6723 585
R2524 gnd.n780 gnd.n779 585
R2525 gnd.n779 gnd.n778 585
R2526 gnd.n6730 gnd.n6729 585
R2527 gnd.n6731 gnd.n6730 585
R2528 gnd.n777 gnd.n776 585
R2529 gnd.n6732 gnd.n777 585
R2530 gnd.n6735 gnd.n6734 585
R2531 gnd.n6734 gnd.n6733 585
R2532 gnd.n774 gnd.n773 585
R2533 gnd.n773 gnd.n772 585
R2534 gnd.n6740 gnd.n6739 585
R2535 gnd.n6741 gnd.n6740 585
R2536 gnd.n771 gnd.n770 585
R2537 gnd.n6742 gnd.n771 585
R2538 gnd.n6745 gnd.n6744 585
R2539 gnd.n6744 gnd.n6743 585
R2540 gnd.n768 gnd.n767 585
R2541 gnd.n767 gnd.n766 585
R2542 gnd.n6750 gnd.n6749 585
R2543 gnd.n6751 gnd.n6750 585
R2544 gnd.n765 gnd.n764 585
R2545 gnd.n6752 gnd.n765 585
R2546 gnd.n6755 gnd.n6754 585
R2547 gnd.n6754 gnd.n6753 585
R2548 gnd.n762 gnd.n761 585
R2549 gnd.n761 gnd.n760 585
R2550 gnd.n6760 gnd.n6759 585
R2551 gnd.n6761 gnd.n6760 585
R2552 gnd.n759 gnd.n758 585
R2553 gnd.n6762 gnd.n759 585
R2554 gnd.n6765 gnd.n6764 585
R2555 gnd.n6764 gnd.n6763 585
R2556 gnd.n756 gnd.n755 585
R2557 gnd.n755 gnd.n754 585
R2558 gnd.n6770 gnd.n6769 585
R2559 gnd.n6771 gnd.n6770 585
R2560 gnd.n753 gnd.n752 585
R2561 gnd.n6772 gnd.n753 585
R2562 gnd.n6775 gnd.n6774 585
R2563 gnd.n6774 gnd.n6773 585
R2564 gnd.n750 gnd.n749 585
R2565 gnd.n749 gnd.n748 585
R2566 gnd.n6780 gnd.n6779 585
R2567 gnd.n6781 gnd.n6780 585
R2568 gnd.n747 gnd.n746 585
R2569 gnd.n6782 gnd.n747 585
R2570 gnd.n6785 gnd.n6784 585
R2571 gnd.n6784 gnd.n6783 585
R2572 gnd.n744 gnd.n743 585
R2573 gnd.n743 gnd.n742 585
R2574 gnd.n6790 gnd.n6789 585
R2575 gnd.n6791 gnd.n6790 585
R2576 gnd.n741 gnd.n740 585
R2577 gnd.n6792 gnd.n741 585
R2578 gnd.n6795 gnd.n6794 585
R2579 gnd.n6794 gnd.n6793 585
R2580 gnd.n738 gnd.n737 585
R2581 gnd.n737 gnd.n736 585
R2582 gnd.n6800 gnd.n6799 585
R2583 gnd.n6801 gnd.n6800 585
R2584 gnd.n735 gnd.n734 585
R2585 gnd.n6802 gnd.n735 585
R2586 gnd.n6805 gnd.n6804 585
R2587 gnd.n6804 gnd.n6803 585
R2588 gnd.n732 gnd.n731 585
R2589 gnd.n731 gnd.n730 585
R2590 gnd.n6810 gnd.n6809 585
R2591 gnd.n6811 gnd.n6810 585
R2592 gnd.n729 gnd.n728 585
R2593 gnd.n6812 gnd.n729 585
R2594 gnd.n6815 gnd.n6814 585
R2595 gnd.n6814 gnd.n6813 585
R2596 gnd.n726 gnd.n725 585
R2597 gnd.n725 gnd.n724 585
R2598 gnd.n6820 gnd.n6819 585
R2599 gnd.n6821 gnd.n6820 585
R2600 gnd.n723 gnd.n722 585
R2601 gnd.n6822 gnd.n723 585
R2602 gnd.n6825 gnd.n6824 585
R2603 gnd.n6824 gnd.n6823 585
R2604 gnd.n720 gnd.n719 585
R2605 gnd.n719 gnd.n718 585
R2606 gnd.n6830 gnd.n6829 585
R2607 gnd.n6831 gnd.n6830 585
R2608 gnd.n717 gnd.n716 585
R2609 gnd.n6832 gnd.n717 585
R2610 gnd.n6835 gnd.n6834 585
R2611 gnd.n6834 gnd.n6833 585
R2612 gnd.n714 gnd.n713 585
R2613 gnd.n713 gnd.n712 585
R2614 gnd.n6840 gnd.n6839 585
R2615 gnd.n6841 gnd.n6840 585
R2616 gnd.n711 gnd.n710 585
R2617 gnd.n6842 gnd.n711 585
R2618 gnd.n6845 gnd.n6844 585
R2619 gnd.n6844 gnd.n6843 585
R2620 gnd.n708 gnd.n707 585
R2621 gnd.n707 gnd.n706 585
R2622 gnd.n6850 gnd.n6849 585
R2623 gnd.n6851 gnd.n6850 585
R2624 gnd.n705 gnd.n704 585
R2625 gnd.n6852 gnd.n705 585
R2626 gnd.n6855 gnd.n6854 585
R2627 gnd.n6854 gnd.n6853 585
R2628 gnd.n702 gnd.n701 585
R2629 gnd.n701 gnd.n700 585
R2630 gnd.n6860 gnd.n6859 585
R2631 gnd.n6861 gnd.n6860 585
R2632 gnd.n699 gnd.n698 585
R2633 gnd.n6862 gnd.n699 585
R2634 gnd.n6865 gnd.n6864 585
R2635 gnd.n6864 gnd.n6863 585
R2636 gnd.n696 gnd.n695 585
R2637 gnd.n695 gnd.n694 585
R2638 gnd.n6870 gnd.n6869 585
R2639 gnd.n6871 gnd.n6870 585
R2640 gnd.n693 gnd.n692 585
R2641 gnd.n6872 gnd.n693 585
R2642 gnd.n6875 gnd.n6874 585
R2643 gnd.n6874 gnd.n6873 585
R2644 gnd.n690 gnd.n689 585
R2645 gnd.n689 gnd.n688 585
R2646 gnd.n6880 gnd.n6879 585
R2647 gnd.n6881 gnd.n6880 585
R2648 gnd.n687 gnd.n686 585
R2649 gnd.n6882 gnd.n687 585
R2650 gnd.n6885 gnd.n6884 585
R2651 gnd.n6884 gnd.n6883 585
R2652 gnd.n684 gnd.n683 585
R2653 gnd.n683 gnd.n682 585
R2654 gnd.n6890 gnd.n6889 585
R2655 gnd.n6891 gnd.n6890 585
R2656 gnd.n681 gnd.n680 585
R2657 gnd.n6892 gnd.n681 585
R2658 gnd.n6895 gnd.n6894 585
R2659 gnd.n6894 gnd.n6893 585
R2660 gnd.n678 gnd.n677 585
R2661 gnd.n677 gnd.n676 585
R2662 gnd.n6900 gnd.n6899 585
R2663 gnd.n6901 gnd.n6900 585
R2664 gnd.n675 gnd.n674 585
R2665 gnd.n6902 gnd.n675 585
R2666 gnd.n6905 gnd.n6904 585
R2667 gnd.n6904 gnd.n6903 585
R2668 gnd.n672 gnd.n671 585
R2669 gnd.n671 gnd.n670 585
R2670 gnd.n6910 gnd.n6909 585
R2671 gnd.n6911 gnd.n6910 585
R2672 gnd.n669 gnd.n668 585
R2673 gnd.n6912 gnd.n669 585
R2674 gnd.n6915 gnd.n6914 585
R2675 gnd.n6914 gnd.n6913 585
R2676 gnd.n666 gnd.n665 585
R2677 gnd.n665 gnd.n664 585
R2678 gnd.n6920 gnd.n6919 585
R2679 gnd.n6921 gnd.n6920 585
R2680 gnd.n663 gnd.n662 585
R2681 gnd.n6922 gnd.n663 585
R2682 gnd.n6925 gnd.n6924 585
R2683 gnd.n6924 gnd.n6923 585
R2684 gnd.n660 gnd.n659 585
R2685 gnd.n659 gnd.n658 585
R2686 gnd.n6930 gnd.n6929 585
R2687 gnd.n6931 gnd.n6930 585
R2688 gnd.n657 gnd.n656 585
R2689 gnd.n6932 gnd.n657 585
R2690 gnd.n6935 gnd.n6934 585
R2691 gnd.n6934 gnd.n6933 585
R2692 gnd.n654 gnd.n653 585
R2693 gnd.n653 gnd.n652 585
R2694 gnd.n6940 gnd.n6939 585
R2695 gnd.n6941 gnd.n6940 585
R2696 gnd.n651 gnd.n650 585
R2697 gnd.n6942 gnd.n651 585
R2698 gnd.n6945 gnd.n6944 585
R2699 gnd.n6944 gnd.n6943 585
R2700 gnd.n648 gnd.n647 585
R2701 gnd.n647 gnd.n646 585
R2702 gnd.n6950 gnd.n6949 585
R2703 gnd.n6951 gnd.n6950 585
R2704 gnd.n645 gnd.n644 585
R2705 gnd.n6952 gnd.n645 585
R2706 gnd.n6955 gnd.n6954 585
R2707 gnd.n6954 gnd.n6953 585
R2708 gnd.n642 gnd.n641 585
R2709 gnd.n641 gnd.n640 585
R2710 gnd.n6960 gnd.n6959 585
R2711 gnd.n6961 gnd.n6960 585
R2712 gnd.n639 gnd.n638 585
R2713 gnd.n6962 gnd.n639 585
R2714 gnd.n6965 gnd.n6964 585
R2715 gnd.n6964 gnd.n6963 585
R2716 gnd.n636 gnd.n635 585
R2717 gnd.n635 gnd.n634 585
R2718 gnd.n6970 gnd.n6969 585
R2719 gnd.n6971 gnd.n6970 585
R2720 gnd.n633 gnd.n632 585
R2721 gnd.n6972 gnd.n633 585
R2722 gnd.n6975 gnd.n6974 585
R2723 gnd.n6974 gnd.n6973 585
R2724 gnd.n630 gnd.n629 585
R2725 gnd.n629 gnd.n628 585
R2726 gnd.n6980 gnd.n6979 585
R2727 gnd.n6981 gnd.n6980 585
R2728 gnd.n627 gnd.n626 585
R2729 gnd.n6982 gnd.n627 585
R2730 gnd.n6985 gnd.n6984 585
R2731 gnd.n6984 gnd.n6983 585
R2732 gnd.n624 gnd.n623 585
R2733 gnd.n623 gnd.n622 585
R2734 gnd.n6990 gnd.n6989 585
R2735 gnd.n6991 gnd.n6990 585
R2736 gnd.n621 gnd.n620 585
R2737 gnd.n6992 gnd.n621 585
R2738 gnd.n6995 gnd.n6994 585
R2739 gnd.n6994 gnd.n6993 585
R2740 gnd.n618 gnd.n617 585
R2741 gnd.n617 gnd.n616 585
R2742 gnd.n7000 gnd.n6999 585
R2743 gnd.n7001 gnd.n7000 585
R2744 gnd.n615 gnd.n614 585
R2745 gnd.n7002 gnd.n615 585
R2746 gnd.n7005 gnd.n7004 585
R2747 gnd.n7004 gnd.n7003 585
R2748 gnd.n612 gnd.n611 585
R2749 gnd.n611 gnd.n610 585
R2750 gnd.n7010 gnd.n7009 585
R2751 gnd.n7011 gnd.n7010 585
R2752 gnd.n609 gnd.n608 585
R2753 gnd.n7012 gnd.n609 585
R2754 gnd.n7015 gnd.n7014 585
R2755 gnd.n7014 gnd.n7013 585
R2756 gnd.n606 gnd.n605 585
R2757 gnd.n605 gnd.n604 585
R2758 gnd.n7020 gnd.n7019 585
R2759 gnd.n7021 gnd.n7020 585
R2760 gnd.n603 gnd.n602 585
R2761 gnd.n7022 gnd.n603 585
R2762 gnd.n7025 gnd.n7024 585
R2763 gnd.n7024 gnd.n7023 585
R2764 gnd.n600 gnd.n599 585
R2765 gnd.n599 gnd.n598 585
R2766 gnd.n7030 gnd.n7029 585
R2767 gnd.n7031 gnd.n7030 585
R2768 gnd.n597 gnd.n596 585
R2769 gnd.n7032 gnd.n597 585
R2770 gnd.n7035 gnd.n7034 585
R2771 gnd.n7034 gnd.n7033 585
R2772 gnd.n594 gnd.n593 585
R2773 gnd.n593 gnd.n592 585
R2774 gnd.n7040 gnd.n7039 585
R2775 gnd.n7041 gnd.n7040 585
R2776 gnd.n591 gnd.n590 585
R2777 gnd.n7042 gnd.n591 585
R2778 gnd.n7045 gnd.n7044 585
R2779 gnd.n7044 gnd.n7043 585
R2780 gnd.n588 gnd.n587 585
R2781 gnd.n587 gnd.n586 585
R2782 gnd.n7050 gnd.n7049 585
R2783 gnd.n7051 gnd.n7050 585
R2784 gnd.n585 gnd.n584 585
R2785 gnd.n7052 gnd.n585 585
R2786 gnd.n7055 gnd.n7054 585
R2787 gnd.n7054 gnd.n7053 585
R2788 gnd.n582 gnd.n581 585
R2789 gnd.n581 gnd.n580 585
R2790 gnd.n7060 gnd.n7059 585
R2791 gnd.n7061 gnd.n7060 585
R2792 gnd.n579 gnd.n578 585
R2793 gnd.n7062 gnd.n579 585
R2794 gnd.n7065 gnd.n7064 585
R2795 gnd.n7064 gnd.n7063 585
R2796 gnd.n576 gnd.n575 585
R2797 gnd.n575 gnd.n574 585
R2798 gnd.n7070 gnd.n7069 585
R2799 gnd.n7071 gnd.n7070 585
R2800 gnd.n573 gnd.n572 585
R2801 gnd.n7072 gnd.n573 585
R2802 gnd.n7075 gnd.n7074 585
R2803 gnd.n7074 gnd.n7073 585
R2804 gnd.n570 gnd.n569 585
R2805 gnd.n569 gnd.n568 585
R2806 gnd.n7080 gnd.n7079 585
R2807 gnd.n7081 gnd.n7080 585
R2808 gnd.n567 gnd.n566 585
R2809 gnd.n7082 gnd.n567 585
R2810 gnd.n7085 gnd.n7084 585
R2811 gnd.n7084 gnd.n7083 585
R2812 gnd.n564 gnd.n563 585
R2813 gnd.n563 gnd.n562 585
R2814 gnd.n7090 gnd.n7089 585
R2815 gnd.n7091 gnd.n7090 585
R2816 gnd.n561 gnd.n560 585
R2817 gnd.n7092 gnd.n561 585
R2818 gnd.n7095 gnd.n7094 585
R2819 gnd.n7094 gnd.n7093 585
R2820 gnd.n558 gnd.n557 585
R2821 gnd.n557 gnd.n556 585
R2822 gnd.n7100 gnd.n7099 585
R2823 gnd.n7101 gnd.n7100 585
R2824 gnd.n555 gnd.n554 585
R2825 gnd.n7102 gnd.n555 585
R2826 gnd.n7105 gnd.n7104 585
R2827 gnd.n7104 gnd.n7103 585
R2828 gnd.n552 gnd.n551 585
R2829 gnd.n551 gnd.n550 585
R2830 gnd.n7110 gnd.n7109 585
R2831 gnd.n7111 gnd.n7110 585
R2832 gnd.n549 gnd.n548 585
R2833 gnd.n7112 gnd.n549 585
R2834 gnd.n7115 gnd.n7114 585
R2835 gnd.n7114 gnd.n7113 585
R2836 gnd.n546 gnd.n545 585
R2837 gnd.n545 gnd.n544 585
R2838 gnd.n7120 gnd.n7119 585
R2839 gnd.n7121 gnd.n7120 585
R2840 gnd.n543 gnd.n542 585
R2841 gnd.n7122 gnd.n543 585
R2842 gnd.n7125 gnd.n7124 585
R2843 gnd.n7124 gnd.n7123 585
R2844 gnd.n540 gnd.n539 585
R2845 gnd.n539 gnd.n538 585
R2846 gnd.n7130 gnd.n7129 585
R2847 gnd.n7131 gnd.n7130 585
R2848 gnd.n537 gnd.n536 585
R2849 gnd.n7132 gnd.n537 585
R2850 gnd.n7135 gnd.n7134 585
R2851 gnd.n7134 gnd.n7133 585
R2852 gnd.n534 gnd.n533 585
R2853 gnd.n533 gnd.n532 585
R2854 gnd.n7140 gnd.n7139 585
R2855 gnd.n7141 gnd.n7140 585
R2856 gnd.n531 gnd.n530 585
R2857 gnd.n7142 gnd.n531 585
R2858 gnd.n7145 gnd.n7144 585
R2859 gnd.n7144 gnd.n7143 585
R2860 gnd.n528 gnd.n527 585
R2861 gnd.n527 gnd.n526 585
R2862 gnd.n7150 gnd.n7149 585
R2863 gnd.n7151 gnd.n7150 585
R2864 gnd.n525 gnd.n524 585
R2865 gnd.n7152 gnd.n525 585
R2866 gnd.n7155 gnd.n7154 585
R2867 gnd.n7154 gnd.n7153 585
R2868 gnd.n7366 gnd.n7365 585
R2869 gnd.n7365 gnd.n7364 585
R2870 gnd.n399 gnd.n398 585
R2871 gnd.n7363 gnd.n399 585
R2872 gnd.n7361 gnd.n7360 585
R2873 gnd.n7362 gnd.n7361 585
R2874 gnd.n402 gnd.n401 585
R2875 gnd.n401 gnd.n400 585
R2876 gnd.n7355 gnd.n7354 585
R2877 gnd.n7354 gnd.n7353 585
R2878 gnd.n405 gnd.n404 585
R2879 gnd.n7352 gnd.n405 585
R2880 gnd.n7350 gnd.n7349 585
R2881 gnd.n7351 gnd.n7350 585
R2882 gnd.n408 gnd.n407 585
R2883 gnd.n407 gnd.n406 585
R2884 gnd.n7345 gnd.n7344 585
R2885 gnd.n7344 gnd.n7343 585
R2886 gnd.n411 gnd.n410 585
R2887 gnd.n7342 gnd.n411 585
R2888 gnd.n7340 gnd.n7339 585
R2889 gnd.n7341 gnd.n7340 585
R2890 gnd.n414 gnd.n413 585
R2891 gnd.n413 gnd.n412 585
R2892 gnd.n7335 gnd.n7334 585
R2893 gnd.n7334 gnd.n7333 585
R2894 gnd.n417 gnd.n416 585
R2895 gnd.n7332 gnd.n417 585
R2896 gnd.n7330 gnd.n7329 585
R2897 gnd.n7331 gnd.n7330 585
R2898 gnd.n420 gnd.n419 585
R2899 gnd.n419 gnd.n418 585
R2900 gnd.n7325 gnd.n7324 585
R2901 gnd.n7324 gnd.n7323 585
R2902 gnd.n423 gnd.n422 585
R2903 gnd.n7322 gnd.n423 585
R2904 gnd.n7320 gnd.n7319 585
R2905 gnd.n7321 gnd.n7320 585
R2906 gnd.n426 gnd.n425 585
R2907 gnd.n425 gnd.n424 585
R2908 gnd.n7315 gnd.n7314 585
R2909 gnd.n7314 gnd.n7313 585
R2910 gnd.n429 gnd.n428 585
R2911 gnd.n7312 gnd.n429 585
R2912 gnd.n7310 gnd.n7309 585
R2913 gnd.n7311 gnd.n7310 585
R2914 gnd.n432 gnd.n431 585
R2915 gnd.n431 gnd.n430 585
R2916 gnd.n7305 gnd.n7304 585
R2917 gnd.n7304 gnd.n7303 585
R2918 gnd.n435 gnd.n434 585
R2919 gnd.n7302 gnd.n435 585
R2920 gnd.n7300 gnd.n7299 585
R2921 gnd.n7301 gnd.n7300 585
R2922 gnd.n438 gnd.n437 585
R2923 gnd.n437 gnd.n436 585
R2924 gnd.n7295 gnd.n7294 585
R2925 gnd.n7294 gnd.n7293 585
R2926 gnd.n441 gnd.n440 585
R2927 gnd.n7292 gnd.n441 585
R2928 gnd.n7290 gnd.n7289 585
R2929 gnd.n7291 gnd.n7290 585
R2930 gnd.n444 gnd.n443 585
R2931 gnd.n443 gnd.n442 585
R2932 gnd.n7285 gnd.n7284 585
R2933 gnd.n7284 gnd.n7283 585
R2934 gnd.n447 gnd.n446 585
R2935 gnd.n7282 gnd.n447 585
R2936 gnd.n7280 gnd.n7279 585
R2937 gnd.n7281 gnd.n7280 585
R2938 gnd.n450 gnd.n449 585
R2939 gnd.n449 gnd.n448 585
R2940 gnd.n7275 gnd.n7274 585
R2941 gnd.n7274 gnd.n7273 585
R2942 gnd.n453 gnd.n452 585
R2943 gnd.n7272 gnd.n453 585
R2944 gnd.n7270 gnd.n7269 585
R2945 gnd.n7271 gnd.n7270 585
R2946 gnd.n456 gnd.n455 585
R2947 gnd.n455 gnd.n454 585
R2948 gnd.n7265 gnd.n7264 585
R2949 gnd.n7264 gnd.n7263 585
R2950 gnd.n459 gnd.n458 585
R2951 gnd.n7262 gnd.n459 585
R2952 gnd.n7260 gnd.n7259 585
R2953 gnd.n7261 gnd.n7260 585
R2954 gnd.n462 gnd.n461 585
R2955 gnd.n461 gnd.n460 585
R2956 gnd.n7255 gnd.n7254 585
R2957 gnd.n7254 gnd.n7253 585
R2958 gnd.n465 gnd.n464 585
R2959 gnd.n7252 gnd.n465 585
R2960 gnd.n7250 gnd.n7249 585
R2961 gnd.n7251 gnd.n7250 585
R2962 gnd.n468 gnd.n467 585
R2963 gnd.n467 gnd.n466 585
R2964 gnd.n7245 gnd.n7244 585
R2965 gnd.n7244 gnd.n7243 585
R2966 gnd.n471 gnd.n470 585
R2967 gnd.n7242 gnd.n471 585
R2968 gnd.n7240 gnd.n7239 585
R2969 gnd.n7241 gnd.n7240 585
R2970 gnd.n474 gnd.n473 585
R2971 gnd.n473 gnd.n472 585
R2972 gnd.n7235 gnd.n7234 585
R2973 gnd.n7234 gnd.n7233 585
R2974 gnd.n477 gnd.n476 585
R2975 gnd.n7232 gnd.n477 585
R2976 gnd.n7230 gnd.n7229 585
R2977 gnd.n7231 gnd.n7230 585
R2978 gnd.n480 gnd.n479 585
R2979 gnd.n479 gnd.n478 585
R2980 gnd.n7225 gnd.n7224 585
R2981 gnd.n7224 gnd.n7223 585
R2982 gnd.n483 gnd.n482 585
R2983 gnd.n7222 gnd.n483 585
R2984 gnd.n7220 gnd.n7219 585
R2985 gnd.n7221 gnd.n7220 585
R2986 gnd.n486 gnd.n485 585
R2987 gnd.n485 gnd.n484 585
R2988 gnd.n7215 gnd.n7214 585
R2989 gnd.n7214 gnd.n7213 585
R2990 gnd.n489 gnd.n488 585
R2991 gnd.n7212 gnd.n489 585
R2992 gnd.n7210 gnd.n7209 585
R2993 gnd.n7211 gnd.n7210 585
R2994 gnd.n492 gnd.n491 585
R2995 gnd.n491 gnd.n490 585
R2996 gnd.n7205 gnd.n7204 585
R2997 gnd.n7204 gnd.n7203 585
R2998 gnd.n495 gnd.n494 585
R2999 gnd.n7202 gnd.n495 585
R3000 gnd.n7200 gnd.n7199 585
R3001 gnd.n7201 gnd.n7200 585
R3002 gnd.n498 gnd.n497 585
R3003 gnd.n497 gnd.n496 585
R3004 gnd.n7195 gnd.n7194 585
R3005 gnd.n7194 gnd.n7193 585
R3006 gnd.n501 gnd.n500 585
R3007 gnd.n7192 gnd.n501 585
R3008 gnd.n7190 gnd.n7189 585
R3009 gnd.n7191 gnd.n7190 585
R3010 gnd.n504 gnd.n503 585
R3011 gnd.n503 gnd.n502 585
R3012 gnd.n7185 gnd.n7184 585
R3013 gnd.n7184 gnd.n7183 585
R3014 gnd.n507 gnd.n506 585
R3015 gnd.n7182 gnd.n507 585
R3016 gnd.n7180 gnd.n7179 585
R3017 gnd.n7181 gnd.n7180 585
R3018 gnd.n510 gnd.n509 585
R3019 gnd.n509 gnd.n508 585
R3020 gnd.n7175 gnd.n7174 585
R3021 gnd.n7174 gnd.n7173 585
R3022 gnd.n513 gnd.n512 585
R3023 gnd.n7172 gnd.n513 585
R3024 gnd.n7170 gnd.n7169 585
R3025 gnd.n7171 gnd.n7170 585
R3026 gnd.n516 gnd.n515 585
R3027 gnd.n515 gnd.n514 585
R3028 gnd.n7165 gnd.n7164 585
R3029 gnd.n7164 gnd.n7163 585
R3030 gnd.n519 gnd.n518 585
R3031 gnd.n7162 gnd.n519 585
R3032 gnd.n7160 gnd.n7159 585
R3033 gnd.n7161 gnd.n7160 585
R3034 gnd.n522 gnd.n521 585
R3035 gnd.n521 gnd.n520 585
R3036 gnd.n1401 gnd.n1400 585
R3037 gnd.n3329 gnd.n1401 585
R3038 gnd.n4839 gnd.n4838 585
R3039 gnd.n4838 gnd.n4837 585
R3040 gnd.n4840 gnd.n1395 585
R3041 gnd.n3258 gnd.n1395 585
R3042 gnd.n4842 gnd.n4841 585
R3043 gnd.n4843 gnd.n4842 585
R3044 gnd.n1379 gnd.n1378 585
R3045 gnd.n3188 gnd.n1379 585
R3046 gnd.n4851 gnd.n4850 585
R3047 gnd.n4850 gnd.n4849 585
R3048 gnd.n4852 gnd.n1373 585
R3049 gnd.n3196 gnd.n1373 585
R3050 gnd.n4854 gnd.n4853 585
R3051 gnd.n4855 gnd.n4854 585
R3052 gnd.n1358 gnd.n1357 585
R3053 gnd.n3178 gnd.n1358 585
R3054 gnd.n4863 gnd.n4862 585
R3055 gnd.n4862 gnd.n4861 585
R3056 gnd.n4864 gnd.n1352 585
R3057 gnd.n3170 gnd.n1352 585
R3058 gnd.n4866 gnd.n4865 585
R3059 gnd.n4867 gnd.n4866 585
R3060 gnd.n1337 gnd.n1336 585
R3061 gnd.n3161 gnd.n1337 585
R3062 gnd.n4875 gnd.n4874 585
R3063 gnd.n4874 gnd.n4873 585
R3064 gnd.n4876 gnd.n1331 585
R3065 gnd.n3153 gnd.n1331 585
R3066 gnd.n4878 gnd.n4877 585
R3067 gnd.n4879 gnd.n4878 585
R3068 gnd.n1316 gnd.n1315 585
R3069 gnd.n3145 gnd.n1316 585
R3070 gnd.n4887 gnd.n4886 585
R3071 gnd.n4886 gnd.n4885 585
R3072 gnd.n4888 gnd.n1310 585
R3073 gnd.n3137 gnd.n1310 585
R3074 gnd.n4890 gnd.n4889 585
R3075 gnd.n4891 gnd.n4890 585
R3076 gnd.n1295 gnd.n1294 585
R3077 gnd.n3129 gnd.n1295 585
R3078 gnd.n4899 gnd.n4898 585
R3079 gnd.n4898 gnd.n4897 585
R3080 gnd.n4900 gnd.n1289 585
R3081 gnd.n3121 gnd.n1289 585
R3082 gnd.n4902 gnd.n4901 585
R3083 gnd.n4903 gnd.n4902 585
R3084 gnd.n1274 gnd.n1273 585
R3085 gnd.n3113 gnd.n1274 585
R3086 gnd.n4911 gnd.n4910 585
R3087 gnd.n4910 gnd.n4909 585
R3088 gnd.n4912 gnd.n1268 585
R3089 gnd.n3105 gnd.n1268 585
R3090 gnd.n4914 gnd.n4913 585
R3091 gnd.n4915 gnd.n4914 585
R3092 gnd.n1255 gnd.n1254 585
R3093 gnd.n3097 gnd.n1255 585
R3094 gnd.n4924 gnd.n4923 585
R3095 gnd.n4923 gnd.n4922 585
R3096 gnd.n4925 gnd.n1250 585
R3097 gnd.n3089 gnd.n1250 585
R3098 gnd.n4927 gnd.n4926 585
R3099 gnd.n4928 gnd.n4927 585
R3100 gnd.n1238 gnd.n1237 585
R3101 gnd.n3081 gnd.n1238 585
R3102 gnd.n4937 gnd.n4936 585
R3103 gnd.n4936 gnd.n4935 585
R3104 gnd.n4938 gnd.n1232 585
R3105 gnd.n3073 gnd.n1232 585
R3106 gnd.n4940 gnd.n4939 585
R3107 gnd.n4941 gnd.n4940 585
R3108 gnd.n1218 gnd.n1217 585
R3109 gnd.n3065 gnd.n1218 585
R3110 gnd.n4950 gnd.n4949 585
R3111 gnd.n4949 gnd.n4948 585
R3112 gnd.n4951 gnd.n1212 585
R3113 gnd.n3057 gnd.n1212 585
R3114 gnd.n4953 gnd.n4952 585
R3115 gnd.n4954 gnd.n4953 585
R3116 gnd.n1197 gnd.n1196 585
R3117 gnd.n3049 gnd.n1197 585
R3118 gnd.n4962 gnd.n4961 585
R3119 gnd.n4961 gnd.n4960 585
R3120 gnd.n4963 gnd.n1191 585
R3121 gnd.n3041 gnd.n1191 585
R3122 gnd.n4965 gnd.n4964 585
R3123 gnd.n4966 gnd.n4965 585
R3124 gnd.n1175 gnd.n1174 585
R3125 gnd.n3033 gnd.n1175 585
R3126 gnd.n4974 gnd.n4973 585
R3127 gnd.n4973 gnd.n4972 585
R3128 gnd.n4975 gnd.n1169 585
R3129 gnd.n1176 gnd.n1169 585
R3130 gnd.n4977 gnd.n4976 585
R3131 gnd.n4978 gnd.n4977 585
R3132 gnd.n1156 gnd.n1155 585
R3133 gnd.n1159 gnd.n1156 585
R3134 gnd.n4986 gnd.n4985 585
R3135 gnd.n4985 gnd.n4984 585
R3136 gnd.n4987 gnd.n1150 585
R3137 gnd.n1150 gnd.n1149 585
R3138 gnd.n4989 gnd.n4988 585
R3139 gnd.n4990 gnd.n4989 585
R3140 gnd.n1135 gnd.n1134 585
R3141 gnd.n1139 gnd.n1135 585
R3142 gnd.n4998 gnd.n4997 585
R3143 gnd.n4997 gnd.n4996 585
R3144 gnd.n4999 gnd.n1129 585
R3145 gnd.n1136 gnd.n1129 585
R3146 gnd.n5001 gnd.n5000 585
R3147 gnd.n5002 gnd.n5001 585
R3148 gnd.n1116 gnd.n1115 585
R3149 gnd.n1119 gnd.n1116 585
R3150 gnd.n5010 gnd.n5009 585
R3151 gnd.n5009 gnd.n5008 585
R3152 gnd.n5011 gnd.n1110 585
R3153 gnd.n1110 gnd.n1108 585
R3154 gnd.n5013 gnd.n5012 585
R3155 gnd.n5014 gnd.n5013 585
R3156 gnd.n1111 gnd.n1109 585
R3157 gnd.n1109 gnd.n1096 585
R3158 gnd.n2980 gnd.n1097 585
R3159 gnd.n5020 gnd.n1097 585
R3160 gnd.n2917 gnd.n2915 585
R3161 gnd.n2915 gnd.n1094 585
R3162 gnd.n2985 gnd.n2984 585
R3163 gnd.n2992 gnd.n2985 585
R3164 gnd.n2916 gnd.n2914 585
R3165 gnd.n2914 gnd.n1040 585
R3166 gnd.n2976 gnd.n2975 585
R3167 gnd.n2974 gnd.n2973 585
R3168 gnd.n2972 gnd.n2971 585
R3169 gnd.n2970 gnd.n2969 585
R3170 gnd.n2968 gnd.n2967 585
R3171 gnd.n2966 gnd.n2965 585
R3172 gnd.n2964 gnd.n2963 585
R3173 gnd.n2962 gnd.n2961 585
R3174 gnd.n2960 gnd.n2959 585
R3175 gnd.n2958 gnd.n2957 585
R3176 gnd.n2956 gnd.n2955 585
R3177 gnd.n2954 gnd.n2953 585
R3178 gnd.n2952 gnd.n2951 585
R3179 gnd.n2950 gnd.n2949 585
R3180 gnd.n2948 gnd.n2947 585
R3181 gnd.n2946 gnd.n2945 585
R3182 gnd.n2944 gnd.n2943 585
R3183 gnd.n2936 gnd.n2933 585
R3184 gnd.n2939 gnd.n1039 585
R3185 gnd.n5107 gnd.n1039 585
R3186 gnd.n3332 gnd.n3331 585
R3187 gnd.n3333 gnd.n2621 585
R3188 gnd.n3334 gnd.n2617 585
R3189 gnd.n2611 gnd.n2610 585
R3190 gnd.n3341 gnd.n2609 585
R3191 gnd.n3342 gnd.n2608 585
R3192 gnd.n2607 gnd.n2601 585
R3193 gnd.n3349 gnd.n2600 585
R3194 gnd.n3350 gnd.n2599 585
R3195 gnd.n2593 gnd.n2592 585
R3196 gnd.n3357 gnd.n2591 585
R3197 gnd.n3358 gnd.n2590 585
R3198 gnd.n2589 gnd.n2583 585
R3199 gnd.n3365 gnd.n2582 585
R3200 gnd.n3366 gnd.n2581 585
R3201 gnd.n2573 gnd.n2572 585
R3202 gnd.n3373 gnd.n2571 585
R3203 gnd.n3374 gnd.n2570 585
R3204 gnd.n3375 gnd.n1413 585
R3205 gnd.n4829 gnd.n1413 585
R3206 gnd.n3330 gnd.n2623 585
R3207 gnd.n3330 gnd.n3329 585
R3208 gnd.n2629 gnd.n1404 585
R3209 gnd.n4837 gnd.n1404 585
R3210 gnd.n3257 gnd.n3256 585
R3211 gnd.n3258 gnd.n3257 585
R3212 gnd.n2628 gnd.n1393 585
R3213 gnd.n4843 gnd.n1393 585
R3214 gnd.n3190 gnd.n3189 585
R3215 gnd.n3189 gnd.n3188 585
R3216 gnd.n2690 gnd.n1382 585
R3217 gnd.n4849 gnd.n1382 585
R3218 gnd.n3195 gnd.n3194 585
R3219 gnd.n3196 gnd.n3195 585
R3220 gnd.n2689 gnd.n1372 585
R3221 gnd.n4855 gnd.n1372 585
R3222 gnd.n3177 gnd.n3176 585
R3223 gnd.n3178 gnd.n3177 585
R3224 gnd.n2696 gnd.n1361 585
R3225 gnd.n4861 gnd.n1361 585
R3226 gnd.n3172 gnd.n3171 585
R3227 gnd.n3171 gnd.n3170 585
R3228 gnd.n2698 gnd.n1350 585
R3229 gnd.n4867 gnd.n1350 585
R3230 gnd.n3160 gnd.n3159 585
R3231 gnd.n3161 gnd.n3160 585
R3232 gnd.n2703 gnd.n1340 585
R3233 gnd.n4873 gnd.n1340 585
R3234 gnd.n3155 gnd.n3154 585
R3235 gnd.n3154 gnd.n3153 585
R3236 gnd.n2705 gnd.n1330 585
R3237 gnd.n4879 gnd.n1330 585
R3238 gnd.n3144 gnd.n3143 585
R3239 gnd.n3145 gnd.n3144 585
R3240 gnd.n2710 gnd.n1319 585
R3241 gnd.n4885 gnd.n1319 585
R3242 gnd.n3139 gnd.n3138 585
R3243 gnd.n3138 gnd.n3137 585
R3244 gnd.n2712 gnd.n1308 585
R3245 gnd.n4891 gnd.n1308 585
R3246 gnd.n3128 gnd.n3127 585
R3247 gnd.n3129 gnd.n3128 585
R3248 gnd.n2717 gnd.n1298 585
R3249 gnd.n4897 gnd.n1298 585
R3250 gnd.n3123 gnd.n3122 585
R3251 gnd.n3122 gnd.n3121 585
R3252 gnd.n2719 gnd.n1288 585
R3253 gnd.n4903 gnd.n1288 585
R3254 gnd.n3112 gnd.n3111 585
R3255 gnd.n3113 gnd.n3112 585
R3256 gnd.n2724 gnd.n1277 585
R3257 gnd.n4909 gnd.n1277 585
R3258 gnd.n3107 gnd.n3106 585
R3259 gnd.n3106 gnd.n3105 585
R3260 gnd.n2726 gnd.n1266 585
R3261 gnd.n4915 gnd.n1266 585
R3262 gnd.n3096 gnd.n3095 585
R3263 gnd.n3097 gnd.n3096 585
R3264 gnd.n2730 gnd.n1258 585
R3265 gnd.n4922 gnd.n1258 585
R3266 gnd.n3091 gnd.n3090 585
R3267 gnd.n3090 gnd.n3089 585
R3268 gnd.n2732 gnd.n1249 585
R3269 gnd.n4928 gnd.n1249 585
R3270 gnd.n3080 gnd.n3079 585
R3271 gnd.n3081 gnd.n3080 585
R3272 gnd.n2738 gnd.n1241 585
R3273 gnd.n4935 gnd.n1241 585
R3274 gnd.n3075 gnd.n3074 585
R3275 gnd.n3074 gnd.n3073 585
R3276 gnd.n2740 gnd.n1230 585
R3277 gnd.n4941 gnd.n1230 585
R3278 gnd.n3064 gnd.n3063 585
R3279 gnd.n3065 gnd.n3064 585
R3280 gnd.n2744 gnd.n1221 585
R3281 gnd.n4948 gnd.n1221 585
R3282 gnd.n3059 gnd.n3058 585
R3283 gnd.n3058 gnd.n3057 585
R3284 gnd.n2746 gnd.n1211 585
R3285 gnd.n4954 gnd.n1211 585
R3286 gnd.n3048 gnd.n3047 585
R3287 gnd.n3049 gnd.n3048 585
R3288 gnd.n2861 gnd.n1200 585
R3289 gnd.n4960 gnd.n1200 585
R3290 gnd.n3043 gnd.n3042 585
R3291 gnd.n3042 gnd.n3041 585
R3292 gnd.n2863 gnd.n1189 585
R3293 gnd.n4966 gnd.n1189 585
R3294 gnd.n3032 gnd.n3031 585
R3295 gnd.n3033 gnd.n3032 585
R3296 gnd.n2902 gnd.n1178 585
R3297 gnd.n4972 gnd.n1178 585
R3298 gnd.n3027 gnd.n3026 585
R3299 gnd.n3026 gnd.n1176 585
R3300 gnd.n3025 gnd.n1168 585
R3301 gnd.n4978 gnd.n1168 585
R3302 gnd.n3024 gnd.n3023 585
R3303 gnd.n3023 gnd.n1159 585
R3304 gnd.n2904 gnd.n1158 585
R3305 gnd.n4984 gnd.n1158 585
R3306 gnd.n3019 gnd.n3018 585
R3307 gnd.n3018 gnd.n1149 585
R3308 gnd.n3017 gnd.n1148 585
R3309 gnd.n4990 gnd.n1148 585
R3310 gnd.n3016 gnd.n3015 585
R3311 gnd.n3015 gnd.n1139 585
R3312 gnd.n2906 gnd.n1138 585
R3313 gnd.n4996 gnd.n1138 585
R3314 gnd.n3011 gnd.n3010 585
R3315 gnd.n3010 gnd.n1136 585
R3316 gnd.n3009 gnd.n1128 585
R3317 gnd.n5002 gnd.n1128 585
R3318 gnd.n3008 gnd.n3007 585
R3319 gnd.n3007 gnd.n1119 585
R3320 gnd.n2908 gnd.n1118 585
R3321 gnd.n5008 gnd.n1118 585
R3322 gnd.n3003 gnd.n3002 585
R3323 gnd.n3002 gnd.n1108 585
R3324 gnd.n3001 gnd.n1107 585
R3325 gnd.n5014 gnd.n1107 585
R3326 gnd.n3000 gnd.n2999 585
R3327 gnd.n2999 gnd.n1096 585
R3328 gnd.n2910 gnd.n1095 585
R3329 gnd.n5020 gnd.n1095 585
R3330 gnd.n2995 gnd.n2994 585
R3331 gnd.n2994 gnd.n1094 585
R3332 gnd.n2993 gnd.n2912 585
R3333 gnd.n2993 gnd.n2992 585
R3334 gnd.n2937 gnd.n2913 585
R3335 gnd.n2913 gnd.n1040 585
R3336 gnd.n7570 gnd.n125 585
R3337 gnd.n7666 gnd.n125 585
R3338 gnd.n7571 gnd.n7508 585
R3339 gnd.n7508 gnd.n122 585
R3340 gnd.n7572 gnd.n203 585
R3341 gnd.n7586 gnd.n203 585
R3342 gnd.n216 gnd.n214 585
R3343 gnd.n214 gnd.n212 585
R3344 gnd.n7577 gnd.n7576 585
R3345 gnd.n7578 gnd.n7577 585
R3346 gnd.n215 gnd.n213 585
R3347 gnd.n213 gnd.n209 585
R3348 gnd.n7504 gnd.n7503 585
R3349 gnd.n7503 gnd.n7502 585
R3350 gnd.n219 gnd.n218 585
R3351 gnd.n229 gnd.n219 585
R3352 gnd.n7493 gnd.n7492 585
R3353 gnd.n7494 gnd.n7493 585
R3354 gnd.n231 gnd.n230 585
R3355 gnd.n230 gnd.n226 585
R3356 gnd.n7488 gnd.n7487 585
R3357 gnd.n7487 gnd.n7486 585
R3358 gnd.n234 gnd.n233 585
R3359 gnd.n235 gnd.n234 585
R3360 gnd.n7477 gnd.n7476 585
R3361 gnd.n7478 gnd.n7477 585
R3362 gnd.n245 gnd.n244 585
R3363 gnd.n250 gnd.n244 585
R3364 gnd.n7472 gnd.n7471 585
R3365 gnd.n7471 gnd.n7470 585
R3366 gnd.n248 gnd.n247 585
R3367 gnd.n259 gnd.n248 585
R3368 gnd.n7461 gnd.n7460 585
R3369 gnd.n7462 gnd.n7461 585
R3370 gnd.n261 gnd.n260 585
R3371 gnd.n260 gnd.n256 585
R3372 gnd.n7456 gnd.n7455 585
R3373 gnd.n7455 gnd.n7454 585
R3374 gnd.n264 gnd.n263 585
R3375 gnd.n265 gnd.n264 585
R3376 gnd.n7445 gnd.n7444 585
R3377 gnd.n7446 gnd.n7445 585
R3378 gnd.n276 gnd.n275 585
R3379 gnd.n7373 gnd.n275 585
R3380 gnd.n7440 gnd.n7439 585
R3381 gnd.n7439 gnd.n7438 585
R3382 gnd.n279 gnd.n278 585
R3383 gnd.n7379 gnd.n279 585
R3384 gnd.n7429 gnd.n7428 585
R3385 gnd.n7430 gnd.n7429 585
R3386 gnd.n292 gnd.n291 585
R3387 gnd.n4511 gnd.n291 585
R3388 gnd.n7424 gnd.n7423 585
R3389 gnd.n7423 gnd.n7422 585
R3390 gnd.n295 gnd.n294 585
R3391 gnd.n4515 gnd.n295 585
R3392 gnd.n7400 gnd.n7399 585
R3393 gnd.n7399 gnd.n7398 585
R3394 gnd.n7401 gnd.n325 585
R3395 gnd.n7394 gnd.n325 585
R3396 gnd.n4522 gnd.n323 585
R3397 gnd.n4523 gnd.n4522 585
R3398 gnd.n7405 gnd.n322 585
R3399 gnd.n1704 gnd.n322 585
R3400 gnd.n7406 gnd.n321 585
R3401 gnd.n4542 gnd.n321 585
R3402 gnd.n7407 gnd.n320 585
R3403 gnd.n4547 gnd.n320 585
R3404 gnd.n317 gnd.n315 585
R3405 gnd.n4531 gnd.n315 585
R3406 gnd.n7412 gnd.n7411 585
R3407 gnd.n7413 gnd.n7412 585
R3408 gnd.n316 gnd.n314 585
R3409 gnd.n4495 gnd.n314 585
R3410 gnd.n4565 gnd.n4563 585
R3411 gnd.n4563 gnd.n4562 585
R3412 gnd.n4566 gnd.n1682 585
R3413 gnd.n4559 gnd.n1682 585
R3414 gnd.n4567 gnd.n1681 585
R3415 gnd.n4468 gnd.n1681 585
R3416 gnd.n1719 gnd.n1679 585
R3417 gnd.n4487 gnd.n1719 585
R3418 gnd.n4571 gnd.n1678 585
R3419 gnd.n4439 gnd.n1678 585
R3420 gnd.n4572 gnd.n1677 585
R3421 gnd.n4477 gnd.n1677 585
R3422 gnd.n4573 gnd.n1676 585
R3423 gnd.n4448 gnd.n1676 585
R3424 gnd.n1734 gnd.n1674 585
R3425 gnd.n1735 gnd.n1734 585
R3426 gnd.n4577 gnd.n1673 585
R3427 gnd.n4433 gnd.n1673 585
R3428 gnd.n4578 gnd.n1672 585
R3429 gnd.n4313 gnd.n1672 585
R3430 gnd.n4579 gnd.n1671 585
R3431 gnd.n4423 gnd.n1671 585
R3432 gnd.n4410 gnd.n1669 585
R3433 gnd.n4411 gnd.n4410 585
R3434 gnd.n4583 gnd.n1668 585
R3435 gnd.n1761 gnd.n1668 585
R3436 gnd.n4584 gnd.n1667 585
R3437 gnd.n4401 gnd.n1667 585
R3438 gnd.n4585 gnd.n1666 585
R3439 gnd.n4321 gnd.n1666 585
R3440 gnd.n4390 gnd.n1664 585
R3441 gnd.n4391 gnd.n4390 585
R3442 gnd.n4589 gnd.n1663 585
R3443 gnd.n4378 gnd.n1663 585
R3444 gnd.n4590 gnd.n1662 585
R3445 gnd.n1787 gnd.n1662 585
R3446 gnd.n4591 gnd.n1661 585
R3447 gnd.n4369 gnd.n1661 585
R3448 gnd.n1806 gnd.n1659 585
R3449 gnd.n1807 gnd.n1806 585
R3450 gnd.n4595 gnd.n1658 585
R3451 gnd.n4359 gnd.n1658 585
R3452 gnd.n4596 gnd.n1657 585
R3453 gnd.n4347 gnd.n1657 585
R3454 gnd.n4597 gnd.n1656 585
R3455 gnd.n1825 gnd.n1656 585
R3456 gnd.n1653 gnd.n1651 585
R3457 gnd.n4337 gnd.n1651 585
R3458 gnd.n4602 gnd.n4601 585
R3459 gnd.n4603 gnd.n4602 585
R3460 gnd.n1652 gnd.n1650 585
R3461 gnd.n4284 gnd.n1650 585
R3462 gnd.n1883 gnd.n1637 585
R3463 gnd.n4609 gnd.n1637 585
R3464 gnd.n1884 gnd.n1882 585
R3465 gnd.n1882 gnd.n1633 585
R3466 gnd.n1881 gnd.n1878 585
R3467 gnd.n1877 gnd.n1876 585
R3468 gnd.n1899 gnd.n1898 585
R3469 gnd.n1901 gnd.n1875 585
R3470 gnd.n1904 gnd.n1903 585
R3471 gnd.n1868 gnd.n1867 585
R3472 gnd.n1918 gnd.n1917 585
R3473 gnd.n1920 gnd.n1866 585
R3474 gnd.n1923 gnd.n1922 585
R3475 gnd.n1859 gnd.n1858 585
R3476 gnd.n1937 gnd.n1936 585
R3477 gnd.n1939 gnd.n1857 585
R3478 gnd.n1942 gnd.n1941 585
R3479 gnd.n1850 gnd.n1849 585
R3480 gnd.n1956 gnd.n1955 585
R3481 gnd.n1958 gnd.n1848 585
R3482 gnd.n1961 gnd.n1960 585
R3483 gnd.n1841 gnd.n1838 585
R3484 gnd.n4276 gnd.n4275 585
R3485 gnd.n4276 gnd.n1624 585
R3486 gnd.n7669 gnd.n7668 585
R3487 gnd.n7541 gnd.n120 585
R3488 gnd.n7543 gnd.n7542 585
R3489 gnd.n7539 gnd.n7538 585
R3490 gnd.n7547 gnd.n7537 585
R3491 gnd.n7548 gnd.n7535 585
R3492 gnd.n7549 gnd.n7534 585
R3493 gnd.n7532 gnd.n7530 585
R3494 gnd.n7553 gnd.n7529 585
R3495 gnd.n7554 gnd.n7527 585
R3496 gnd.n7555 gnd.n7526 585
R3497 gnd.n7524 gnd.n7522 585
R3498 gnd.n7559 gnd.n7521 585
R3499 gnd.n7560 gnd.n7519 585
R3500 gnd.n7561 gnd.n7518 585
R3501 gnd.n7516 gnd.n7514 585
R3502 gnd.n7565 gnd.n7513 585
R3503 gnd.n7566 gnd.n7511 585
R3504 gnd.n7567 gnd.n7510 585
R3505 gnd.n7510 gnd.n124 585
R3506 gnd.n7667 gnd.n116 585
R3507 gnd.n7667 gnd.n7666 585
R3508 gnd.n7673 gnd.n115 585
R3509 gnd.n122 gnd.n115 585
R3510 gnd.n7674 gnd.n114 585
R3511 gnd.n7586 gnd.n114 585
R3512 gnd.n7675 gnd.n113 585
R3513 gnd.n212 gnd.n113 585
R3514 gnd.n211 gnd.n111 585
R3515 gnd.n7578 gnd.n211 585
R3516 gnd.n7679 gnd.n110 585
R3517 gnd.n209 gnd.n110 585
R3518 gnd.n7680 gnd.n109 585
R3519 gnd.n7502 gnd.n109 585
R3520 gnd.n7681 gnd.n108 585
R3521 gnd.n229 gnd.n108 585
R3522 gnd.n228 gnd.n106 585
R3523 gnd.n7494 gnd.n228 585
R3524 gnd.n7685 gnd.n105 585
R3525 gnd.n226 gnd.n105 585
R3526 gnd.n7686 gnd.n104 585
R3527 gnd.n7486 gnd.n104 585
R3528 gnd.n7687 gnd.n103 585
R3529 gnd.n235 gnd.n103 585
R3530 gnd.n243 gnd.n101 585
R3531 gnd.n7478 gnd.n243 585
R3532 gnd.n7691 gnd.n100 585
R3533 gnd.n250 gnd.n100 585
R3534 gnd.n7692 gnd.n99 585
R3535 gnd.n7470 gnd.n99 585
R3536 gnd.n7693 gnd.n98 585
R3537 gnd.n259 gnd.n98 585
R3538 gnd.n258 gnd.n96 585
R3539 gnd.n7462 gnd.n258 585
R3540 gnd.n7697 gnd.n95 585
R3541 gnd.n256 gnd.n95 585
R3542 gnd.n7698 gnd.n94 585
R3543 gnd.n7454 gnd.n94 585
R3544 gnd.n7699 gnd.n93 585
R3545 gnd.n265 gnd.n93 585
R3546 gnd.n273 gnd.n91 585
R3547 gnd.n7446 gnd.n273 585
R3548 gnd.n7703 gnd.n90 585
R3549 gnd.n7373 gnd.n90 585
R3550 gnd.n7704 gnd.n89 585
R3551 gnd.n7438 gnd.n89 585
R3552 gnd.n7705 gnd.n88 585
R3553 gnd.n7379 gnd.n88 585
R3554 gnd.n289 gnd.n86 585
R3555 gnd.n7430 gnd.n289 585
R3556 gnd.n7709 gnd.n85 585
R3557 gnd.n4511 gnd.n85 585
R3558 gnd.n7710 gnd.n84 585
R3559 gnd.n7422 gnd.n84 585
R3560 gnd.n7711 gnd.n83 585
R3561 gnd.n4515 gnd.n83 585
R3562 gnd.n327 gnd.n81 585
R3563 gnd.n7398 gnd.n327 585
R3564 gnd.n7715 gnd.n80 585
R3565 gnd.n7394 gnd.n80 585
R3566 gnd.n7716 gnd.n79 585
R3567 gnd.n4523 gnd.n79 585
R3568 gnd.n7717 gnd.n78 585
R3569 gnd.n1704 gnd.n78 585
R3570 gnd.n1697 gnd.n76 585
R3571 gnd.n4542 gnd.n1697 585
R3572 gnd.n4549 gnd.n4548 585
R3573 gnd.n4548 gnd.n4547 585
R3574 gnd.n4551 gnd.n1696 585
R3575 gnd.n4531 gnd.n1696 585
R3576 gnd.n4552 gnd.n312 585
R3577 gnd.n7413 gnd.n312 585
R3578 gnd.n4553 gnd.n1695 585
R3579 gnd.n4495 gnd.n1695 585
R3580 gnd.n1692 gnd.n1685 585
R3581 gnd.n4562 gnd.n1685 585
R3582 gnd.n4558 gnd.n4557 585
R3583 gnd.n4559 gnd.n4558 585
R3584 gnd.n1691 gnd.n1690 585
R3585 gnd.n4468 gnd.n1690 585
R3586 gnd.n4441 gnd.n1717 585
R3587 gnd.n4487 gnd.n1717 585
R3588 gnd.n4442 gnd.n4440 585
R3589 gnd.n4440 gnd.n4439 585
R3590 gnd.n1739 gnd.n1727 585
R3591 gnd.n4477 gnd.n1727 585
R3592 gnd.n4447 gnd.n4446 585
R3593 gnd.n4448 gnd.n4447 585
R3594 gnd.n1738 gnd.n1737 585
R3595 gnd.n1737 gnd.n1735 585
R3596 gnd.n4435 gnd.n4434 585
R3597 gnd.n4434 gnd.n4433 585
R3598 gnd.n1742 gnd.n1741 585
R3599 gnd.n4313 gnd.n1742 585
R3600 gnd.n1765 gnd.n1754 585
R3601 gnd.n4423 gnd.n1754 585
R3602 gnd.n4409 gnd.n4408 585
R3603 gnd.n4411 gnd.n4409 585
R3604 gnd.n1764 gnd.n1763 585
R3605 gnd.n1763 gnd.n1761 585
R3606 gnd.n4403 gnd.n4402 585
R3607 gnd.n4402 gnd.n4401 585
R3608 gnd.n1768 gnd.n1767 585
R3609 gnd.n4321 gnd.n1768 585
R3610 gnd.n1791 gnd.n1780 585
R3611 gnd.n4391 gnd.n1780 585
R3612 gnd.n4377 gnd.n4376 585
R3613 gnd.n4378 gnd.n4377 585
R3614 gnd.n1790 gnd.n1789 585
R3615 gnd.n1789 gnd.n1787 585
R3616 gnd.n4371 gnd.n4370 585
R3617 gnd.n4370 gnd.n4369 585
R3618 gnd.n1794 gnd.n1793 585
R3619 gnd.n1807 gnd.n1794 585
R3620 gnd.n1829 gnd.n1805 585
R3621 gnd.n4359 gnd.n1805 585
R3622 gnd.n4345 gnd.n4344 585
R3623 gnd.n4347 gnd.n4345 585
R3624 gnd.n1828 gnd.n1827 585
R3625 gnd.n1827 gnd.n1825 585
R3626 gnd.n4339 gnd.n4338 585
R3627 gnd.n4338 gnd.n4337 585
R3628 gnd.n1831 gnd.n1648 585
R3629 gnd.n4603 gnd.n1648 585
R3630 gnd.n4283 gnd.n4282 585
R3631 gnd.n4284 gnd.n4283 585
R3632 gnd.n1836 gnd.n1635 585
R3633 gnd.n4609 gnd.n1635 585
R3634 gnd.n4278 gnd.n4277 585
R3635 gnd.n4277 gnd.n1633 585
R3636 gnd.n6406 gnd.n6405 585
R3637 gnd.n6405 gnd.n996 585
R3638 gnd.n984 gnd.n983 585
R3639 gnd.n6410 gnd.n984 585
R3640 gnd.n6521 gnd.n6520 585
R3641 gnd.n6520 gnd.n6519 585
R3642 gnd.n6522 gnd.n978 585
R3643 gnd.n6418 gnd.n978 585
R3644 gnd.n6524 gnd.n6523 585
R3645 gnd.n6525 gnd.n6524 585
R3646 gnd.n979 gnd.n977 585
R3647 gnd.n977 gnd.n973 585
R3648 gnd.n6138 gnd.n6137 585
R3649 gnd.n6137 gnd.n6136 585
R3650 gnd.n5177 gnd.n5176 585
R3651 gnd.n5177 gnd.n963 585
R3652 gnd.n6122 gnd.n6121 585
R3653 gnd.n6123 gnd.n6122 585
R3654 gnd.n5187 gnd.n5186 585
R3655 gnd.n5195 gnd.n5186 585
R3656 gnd.n6099 gnd.n5207 585
R3657 gnd.n5207 gnd.n5194 585
R3658 gnd.n6101 gnd.n6100 585
R3659 gnd.n6102 gnd.n6101 585
R3660 gnd.n5208 gnd.n5206 585
R3661 gnd.n5206 gnd.n5202 585
R3662 gnd.n6088 gnd.n6087 585
R3663 gnd.n6087 gnd.n6086 585
R3664 gnd.n5213 gnd.n5212 585
R3665 gnd.n6057 gnd.n5213 585
R3666 gnd.n6077 gnd.n6076 585
R3667 gnd.n6076 gnd.n6075 585
R3668 gnd.n5220 gnd.n5219 585
R3669 gnd.n6063 gnd.n5220 585
R3670 gnd.n6036 gnd.n5240 585
R3671 gnd.n5240 gnd.n5239 585
R3672 gnd.n6038 gnd.n6037 585
R3673 gnd.n6039 gnd.n6038 585
R3674 gnd.n5241 gnd.n5238 585
R3675 gnd.n5249 gnd.n5238 585
R3676 gnd.n6014 gnd.n5261 585
R3677 gnd.n5261 gnd.n5248 585
R3678 gnd.n6016 gnd.n6015 585
R3679 gnd.n6017 gnd.n6016 585
R3680 gnd.n5262 gnd.n5260 585
R3681 gnd.n5260 gnd.n5256 585
R3682 gnd.n6002 gnd.n6001 585
R3683 gnd.n6001 gnd.n6000 585
R3684 gnd.n5267 gnd.n5266 585
R3685 gnd.n5277 gnd.n5267 585
R3686 gnd.n5991 gnd.n5990 585
R3687 gnd.n5990 gnd.n5989 585
R3688 gnd.n5274 gnd.n5273 585
R3689 gnd.n5977 gnd.n5274 585
R3690 gnd.n5951 gnd.n5355 585
R3691 gnd.n5355 gnd.n5284 585
R3692 gnd.n5953 gnd.n5952 585
R3693 gnd.n5954 gnd.n5953 585
R3694 gnd.n5356 gnd.n5354 585
R3695 gnd.n5364 gnd.n5354 585
R3696 gnd.n5929 gnd.n5376 585
R3697 gnd.n5376 gnd.n5363 585
R3698 gnd.n5931 gnd.n5930 585
R3699 gnd.n5932 gnd.n5931 585
R3700 gnd.n5377 gnd.n5375 585
R3701 gnd.n5375 gnd.n5371 585
R3702 gnd.n5917 gnd.n5916 585
R3703 gnd.n5916 gnd.n5915 585
R3704 gnd.n5382 gnd.n5381 585
R3705 gnd.n5391 gnd.n5382 585
R3706 gnd.n5906 gnd.n5905 585
R3707 gnd.n5905 gnd.n5904 585
R3708 gnd.n5389 gnd.n5388 585
R3709 gnd.n5892 gnd.n5389 585
R3710 gnd.n5864 gnd.n5863 585
R3711 gnd.n5863 gnd.n5398 585
R3712 gnd.n5865 gnd.n5409 585
R3713 gnd.n5856 gnd.n5409 585
R3714 gnd.n5867 gnd.n5866 585
R3715 gnd.n5868 gnd.n5867 585
R3716 gnd.n5410 gnd.n5408 585
R3717 gnd.n5424 gnd.n5408 585
R3718 gnd.n5848 gnd.n5847 585
R3719 gnd.n5847 gnd.n5846 585
R3720 gnd.n5421 gnd.n5420 585
R3721 gnd.n5831 gnd.n5421 585
R3722 gnd.n5818 gnd.n5441 585
R3723 gnd.n5441 gnd.n5431 585
R3724 gnd.n5820 gnd.n5819 585
R3725 gnd.n5821 gnd.n5820 585
R3726 gnd.n5442 gnd.n5440 585
R3727 gnd.n5450 gnd.n5440 585
R3728 gnd.n5794 gnd.n5462 585
R3729 gnd.n5462 gnd.n5449 585
R3730 gnd.n5796 gnd.n5795 585
R3731 gnd.n5797 gnd.n5796 585
R3732 gnd.n5463 gnd.n5461 585
R3733 gnd.n5461 gnd.n5457 585
R3734 gnd.n5782 gnd.n5781 585
R3735 gnd.n5781 gnd.n5780 585
R3736 gnd.n5468 gnd.n5467 585
R3737 gnd.n5472 gnd.n5468 585
R3738 gnd.n5766 gnd.n5765 585
R3739 gnd.n5767 gnd.n5766 585
R3740 gnd.n5483 gnd.n5482 585
R3741 gnd.n5482 gnd.n5478 585
R3742 gnd.n5756 gnd.n5755 585
R3743 gnd.n5757 gnd.n5756 585
R3744 gnd.n5492 gnd.n5491 585
R3745 gnd.n5491 gnd.n5489 585
R3746 gnd.n5750 gnd.n5749 585
R3747 gnd.n5749 gnd.n5748 585
R3748 gnd.n5496 gnd.n5495 585
R3749 gnd.n5504 gnd.n5496 585
R3750 gnd.n5657 gnd.n5656 585
R3751 gnd.n5658 gnd.n5657 585
R3752 gnd.n5506 gnd.n5505 585
R3753 gnd.n5505 gnd.n5503 585
R3754 gnd.n5652 gnd.n5651 585
R3755 gnd.n5651 gnd.n5650 585
R3756 gnd.n5509 gnd.n5508 585
R3757 gnd.n5510 gnd.n5509 585
R3758 gnd.n5641 gnd.n5640 585
R3759 gnd.n5642 gnd.n5641 585
R3760 gnd.n5518 gnd.n5517 585
R3761 gnd.n5517 gnd.n5516 585
R3762 gnd.n5636 gnd.n5635 585
R3763 gnd.n5635 gnd.n5634 585
R3764 gnd.n5521 gnd.n5520 585
R3765 gnd.n5522 gnd.n5521 585
R3766 gnd.n5625 gnd.n5624 585
R3767 gnd.n5626 gnd.n5625 585
R3768 gnd.n5621 gnd.n5528 585
R3769 gnd.n5620 gnd.n5619 585
R3770 gnd.n5617 gnd.n5530 585
R3771 gnd.n5617 gnd.n5527 585
R3772 gnd.n5616 gnd.n5615 585
R3773 gnd.n5614 gnd.n5613 585
R3774 gnd.n5612 gnd.n5535 585
R3775 gnd.n5610 gnd.n5609 585
R3776 gnd.n5608 gnd.n5536 585
R3777 gnd.n5607 gnd.n5606 585
R3778 gnd.n5604 gnd.n5541 585
R3779 gnd.n5602 gnd.n5601 585
R3780 gnd.n5600 gnd.n5542 585
R3781 gnd.n5599 gnd.n5598 585
R3782 gnd.n5596 gnd.n5547 585
R3783 gnd.n5594 gnd.n5593 585
R3784 gnd.n5592 gnd.n5548 585
R3785 gnd.n5591 gnd.n5590 585
R3786 gnd.n5588 gnd.n5553 585
R3787 gnd.n5586 gnd.n5585 585
R3788 gnd.n5584 gnd.n5554 585
R3789 gnd.n5583 gnd.n5582 585
R3790 gnd.n5580 gnd.n5559 585
R3791 gnd.n5578 gnd.n5577 585
R3792 gnd.n5575 gnd.n5560 585
R3793 gnd.n5574 gnd.n5573 585
R3794 gnd.n5571 gnd.n5569 585
R3795 gnd.n5567 gnd.n5526 585
R3796 gnd.n6428 gnd.n6427 585
R3797 gnd.n6430 gnd.n6429 585
R3798 gnd.n6432 gnd.n6431 585
R3799 gnd.n6434 gnd.n6433 585
R3800 gnd.n6436 gnd.n6435 585
R3801 gnd.n6438 gnd.n6437 585
R3802 gnd.n6440 gnd.n6439 585
R3803 gnd.n6442 gnd.n6441 585
R3804 gnd.n6444 gnd.n6443 585
R3805 gnd.n6446 gnd.n6445 585
R3806 gnd.n6448 gnd.n6447 585
R3807 gnd.n6450 gnd.n6449 585
R3808 gnd.n6452 gnd.n6451 585
R3809 gnd.n6454 gnd.n6453 585
R3810 gnd.n6456 gnd.n6455 585
R3811 gnd.n6458 gnd.n6457 585
R3812 gnd.n6460 gnd.n6459 585
R3813 gnd.n6462 gnd.n6461 585
R3814 gnd.n6464 gnd.n6463 585
R3815 gnd.n6466 gnd.n6465 585
R3816 gnd.n6468 gnd.n6467 585
R3817 gnd.n6470 gnd.n6469 585
R3818 gnd.n6472 gnd.n6471 585
R3819 gnd.n6474 gnd.n6473 585
R3820 gnd.n6476 gnd.n6475 585
R3821 gnd.n6477 gnd.n5140 585
R3822 gnd.n6478 gnd.n998 585
R3823 gnd.n6511 gnd.n998 585
R3824 gnd.n6426 gnd.n6425 585
R3825 gnd.n6426 gnd.n996 585
R3826 gnd.n5170 gnd.n5169 585
R3827 gnd.n6410 gnd.n5169 585
R3828 gnd.n6421 gnd.n985 585
R3829 gnd.n6519 gnd.n985 585
R3830 gnd.n6420 gnd.n6419 585
R3831 gnd.n6419 gnd.n6418 585
R3832 gnd.n5172 gnd.n975 585
R3833 gnd.n6525 gnd.n975 585
R3834 gnd.n6131 gnd.n5179 585
R3835 gnd.n5179 gnd.n973 585
R3836 gnd.n6133 gnd.n6132 585
R3837 gnd.n6136 gnd.n6133 585
R3838 gnd.n5180 gnd.n5178 585
R3839 gnd.n5178 gnd.n963 585
R3840 gnd.n6125 gnd.n6124 585
R3841 gnd.n6124 gnd.n6123 585
R3842 gnd.n5183 gnd.n5182 585
R3843 gnd.n5195 gnd.n5183 585
R3844 gnd.n6052 gnd.n6051 585
R3845 gnd.n6051 gnd.n5194 585
R3846 gnd.n6053 gnd.n5204 585
R3847 gnd.n6102 gnd.n5204 585
R3848 gnd.n6055 gnd.n6054 585
R3849 gnd.n6054 gnd.n5202 585
R3850 gnd.n6056 gnd.n5215 585
R3851 gnd.n6086 gnd.n5215 585
R3852 gnd.n6059 gnd.n6058 585
R3853 gnd.n6058 gnd.n6057 585
R3854 gnd.n6060 gnd.n5222 585
R3855 gnd.n6075 gnd.n5222 585
R3856 gnd.n6062 gnd.n6061 585
R3857 gnd.n6063 gnd.n6062 585
R3858 gnd.n5232 gnd.n5231 585
R3859 gnd.n5239 gnd.n5231 585
R3860 gnd.n6041 gnd.n6040 585
R3861 gnd.n6040 gnd.n6039 585
R3862 gnd.n5235 gnd.n5234 585
R3863 gnd.n5249 gnd.n5235 585
R3864 gnd.n5967 gnd.n5966 585
R3865 gnd.n5966 gnd.n5248 585
R3866 gnd.n5968 gnd.n5258 585
R3867 gnd.n6017 gnd.n5258 585
R3868 gnd.n5970 gnd.n5969 585
R3869 gnd.n5969 gnd.n5256 585
R3870 gnd.n5971 gnd.n5269 585
R3871 gnd.n6000 gnd.n5269 585
R3872 gnd.n5973 gnd.n5972 585
R3873 gnd.n5972 gnd.n5277 585
R3874 gnd.n5974 gnd.n5276 585
R3875 gnd.n5989 gnd.n5276 585
R3876 gnd.n5976 gnd.n5975 585
R3877 gnd.n5977 gnd.n5976 585
R3878 gnd.n5288 gnd.n5287 585
R3879 gnd.n5287 gnd.n5284 585
R3880 gnd.n5956 gnd.n5955 585
R3881 gnd.n5955 gnd.n5954 585
R3882 gnd.n5351 gnd.n5350 585
R3883 gnd.n5364 gnd.n5351 585
R3884 gnd.n5877 gnd.n5876 585
R3885 gnd.n5876 gnd.n5363 585
R3886 gnd.n5878 gnd.n5373 585
R3887 gnd.n5932 gnd.n5373 585
R3888 gnd.n5881 gnd.n5880 585
R3889 gnd.n5880 gnd.n5371 585
R3890 gnd.n5882 gnd.n5384 585
R3891 gnd.n5915 gnd.n5384 585
R3892 gnd.n5885 gnd.n5884 585
R3893 gnd.n5884 gnd.n5391 585
R3894 gnd.n5886 gnd.n5390 585
R3895 gnd.n5904 gnd.n5390 585
R3896 gnd.n5889 gnd.n5888 585
R3897 gnd.n5892 gnd.n5889 585
R3898 gnd.n5874 gnd.n5400 585
R3899 gnd.n5400 gnd.n5398 585
R3900 gnd.n5405 gnd.n5401 585
R3901 gnd.n5856 gnd.n5405 585
R3902 gnd.n5870 gnd.n5869 585
R3903 gnd.n5869 gnd.n5868 585
R3904 gnd.n5404 gnd.n5403 585
R3905 gnd.n5424 gnd.n5404 585
R3906 gnd.n5828 gnd.n5423 585
R3907 gnd.n5846 gnd.n5423 585
R3908 gnd.n5830 gnd.n5829 585
R3909 gnd.n5831 gnd.n5830 585
R3910 gnd.n5434 gnd.n5433 585
R3911 gnd.n5433 gnd.n5431 585
R3912 gnd.n5823 gnd.n5822 585
R3913 gnd.n5822 gnd.n5821 585
R3914 gnd.n5437 gnd.n5436 585
R3915 gnd.n5450 gnd.n5437 585
R3916 gnd.n5674 gnd.n5673 585
R3917 gnd.n5673 gnd.n5449 585
R3918 gnd.n5675 gnd.n5459 585
R3919 gnd.n5797 gnd.n5459 585
R3920 gnd.n5677 gnd.n5676 585
R3921 gnd.n5676 gnd.n5457 585
R3922 gnd.n5678 gnd.n5469 585
R3923 gnd.n5780 gnd.n5469 585
R3924 gnd.n5680 gnd.n5679 585
R3925 gnd.n5679 gnd.n5472 585
R3926 gnd.n5681 gnd.n5480 585
R3927 gnd.n5767 gnd.n5480 585
R3928 gnd.n5683 gnd.n5682 585
R3929 gnd.n5682 gnd.n5478 585
R3930 gnd.n5684 gnd.n5490 585
R3931 gnd.n5757 gnd.n5490 585
R3932 gnd.n5685 gnd.n5498 585
R3933 gnd.n5498 gnd.n5489 585
R3934 gnd.n5687 gnd.n5686 585
R3935 gnd.n5748 gnd.n5687 585
R3936 gnd.n5499 gnd.n5497 585
R3937 gnd.n5504 gnd.n5497 585
R3938 gnd.n5660 gnd.n5659 585
R3939 gnd.n5659 gnd.n5658 585
R3940 gnd.n5502 gnd.n5501 585
R3941 gnd.n5503 gnd.n5502 585
R3942 gnd.n5649 gnd.n5648 585
R3943 gnd.n5650 gnd.n5649 585
R3944 gnd.n5512 gnd.n5511 585
R3945 gnd.n5511 gnd.n5510 585
R3946 gnd.n5644 gnd.n5643 585
R3947 gnd.n5643 gnd.n5642 585
R3948 gnd.n5515 gnd.n5514 585
R3949 gnd.n5516 gnd.n5515 585
R3950 gnd.n5633 gnd.n5632 585
R3951 gnd.n5634 gnd.n5633 585
R3952 gnd.n5524 gnd.n5523 585
R3953 gnd.n5523 gnd.n5522 585
R3954 gnd.n5628 gnd.n5627 585
R3955 gnd.n5627 gnd.n5626 585
R3956 gnd.n6514 gnd.n6513 585
R3957 gnd.n6513 gnd.n6512 585
R3958 gnd.n6515 gnd.n988 585
R3959 gnd.n6411 gnd.n988 585
R3960 gnd.n6517 gnd.n6516 585
R3961 gnd.n6518 gnd.n6517 585
R3962 gnd.n989 gnd.n987 585
R3963 gnd.n6417 gnd.n987 585
R3964 gnd.n972 gnd.n971 585
R3965 gnd.n976 gnd.n972 585
R3966 gnd.n6528 gnd.n6527 585
R3967 gnd.n6527 gnd.n6526 585
R3968 gnd.n6529 gnd.n966 585
R3969 gnd.n6135 gnd.n966 585
R3970 gnd.n6531 gnd.n6530 585
R3971 gnd.n6532 gnd.n6531 585
R3972 gnd.n967 gnd.n965 585
R3973 gnd.n5185 gnd.n965 585
R3974 gnd.n6111 gnd.n5197 585
R3975 gnd.n5197 gnd.n5184 585
R3976 gnd.n6113 gnd.n6112 585
R3977 gnd.n6114 gnd.n6113 585
R3978 gnd.n5198 gnd.n5196 585
R3979 gnd.n5205 gnd.n5196 585
R3980 gnd.n6105 gnd.n6104 585
R3981 gnd.n6104 gnd.n6103 585
R3982 gnd.n5201 gnd.n5200 585
R3983 gnd.n6085 gnd.n5201 585
R3984 gnd.n6071 gnd.n5224 585
R3985 gnd.n5224 gnd.n5214 585
R3986 gnd.n6073 gnd.n6072 585
R3987 gnd.n6074 gnd.n6073 585
R3988 gnd.n5225 gnd.n5223 585
R3989 gnd.n5223 gnd.n5221 585
R3990 gnd.n6066 gnd.n6065 585
R3991 gnd.n6065 gnd.n6064 585
R3992 gnd.n5228 gnd.n5227 585
R3993 gnd.n5237 gnd.n5228 585
R3994 gnd.n6025 gnd.n5251 585
R3995 gnd.n5251 gnd.n5236 585
R3996 gnd.n6027 gnd.n6026 585
R3997 gnd.n6028 gnd.n6027 585
R3998 gnd.n5252 gnd.n5250 585
R3999 gnd.n5259 gnd.n5250 585
R4000 gnd.n6020 gnd.n6019 585
R4001 gnd.n6019 gnd.n6018 585
R4002 gnd.n5255 gnd.n5254 585
R4003 gnd.n5999 gnd.n5255 585
R4004 gnd.n5985 gnd.n5279 585
R4005 gnd.n5279 gnd.n5268 585
R4006 gnd.n5987 gnd.n5986 585
R4007 gnd.n5988 gnd.n5987 585
R4008 gnd.n5280 gnd.n5278 585
R4009 gnd.n5278 gnd.n5275 585
R4010 gnd.n5980 gnd.n5979 585
R4011 gnd.n5979 gnd.n5978 585
R4012 gnd.n5283 gnd.n5282 585
R4013 gnd.n5353 gnd.n5283 585
R4014 gnd.n5940 gnd.n5366 585
R4015 gnd.n5366 gnd.n5352 585
R4016 gnd.n5942 gnd.n5941 585
R4017 gnd.n5943 gnd.n5942 585
R4018 gnd.n5367 gnd.n5365 585
R4019 gnd.n5374 gnd.n5365 585
R4020 gnd.n5935 gnd.n5934 585
R4021 gnd.n5934 gnd.n5933 585
R4022 gnd.n5370 gnd.n5369 585
R4023 gnd.n5914 gnd.n5370 585
R4024 gnd.n5900 gnd.n5393 585
R4025 gnd.n5393 gnd.n5383 585
R4026 gnd.n5902 gnd.n5901 585
R4027 gnd.n5903 gnd.n5902 585
R4028 gnd.n5394 gnd.n5392 585
R4029 gnd.n5891 gnd.n5392 585
R4030 gnd.n5895 gnd.n5894 585
R4031 gnd.n5894 gnd.n5893 585
R4032 gnd.n5397 gnd.n5396 585
R4033 gnd.n5857 gnd.n5397 585
R4034 gnd.n5841 gnd.n5840 585
R4035 gnd.n5840 gnd.n5407 585
R4036 gnd.n5842 gnd.n5426 585
R4037 gnd.n5426 gnd.n5406 585
R4038 gnd.n5844 gnd.n5843 585
R4039 gnd.n5845 gnd.n5844 585
R4040 gnd.n5427 gnd.n5425 585
R4041 gnd.n5425 gnd.n5422 585
R4042 gnd.n5834 gnd.n5833 585
R4043 gnd.n5833 gnd.n5832 585
R4044 gnd.n5430 gnd.n5429 585
R4045 gnd.n5439 gnd.n5430 585
R4046 gnd.n5805 gnd.n5452 585
R4047 gnd.n5452 gnd.n5438 585
R4048 gnd.n5807 gnd.n5806 585
R4049 gnd.n5808 gnd.n5807 585
R4050 gnd.n5453 gnd.n5451 585
R4051 gnd.n5460 gnd.n5451 585
R4052 gnd.n5800 gnd.n5799 585
R4053 gnd.n5799 gnd.n5798 585
R4054 gnd.n5456 gnd.n5455 585
R4055 gnd.n5779 gnd.n5456 585
R4056 gnd.n5775 gnd.n5774 585
R4057 gnd.n5776 gnd.n5775 585
R4058 gnd.n5474 gnd.n5473 585
R4059 gnd.n5481 gnd.n5473 585
R4060 gnd.n5770 gnd.n5769 585
R4061 gnd.n5769 gnd.n5768 585
R4062 gnd.n5477 gnd.n5476 585
R4063 gnd.n5758 gnd.n5477 585
R4064 gnd.n5745 gnd.n5744 585
R4065 gnd.n5743 gnd.n5696 585
R4066 gnd.n5742 gnd.n5695 585
R4067 gnd.n5747 gnd.n5695 585
R4068 gnd.n5741 gnd.n5740 585
R4069 gnd.n5739 gnd.n5738 585
R4070 gnd.n5737 gnd.n5736 585
R4071 gnd.n5735 gnd.n5734 585
R4072 gnd.n5733 gnd.n5732 585
R4073 gnd.n5731 gnd.n5730 585
R4074 gnd.n5729 gnd.n5728 585
R4075 gnd.n5727 gnd.n5726 585
R4076 gnd.n5725 gnd.n5724 585
R4077 gnd.n5723 gnd.n5722 585
R4078 gnd.n5721 gnd.n5720 585
R4079 gnd.n5719 gnd.n5718 585
R4080 gnd.n5717 gnd.n5716 585
R4081 gnd.n5712 gnd.n5488 585
R4082 gnd.n5135 gnd.n5134 585
R4083 gnd.n6484 gnd.n6483 585
R4084 gnd.n6486 gnd.n6485 585
R4085 gnd.n6488 gnd.n6487 585
R4086 gnd.n6490 gnd.n6489 585
R4087 gnd.n6492 gnd.n6491 585
R4088 gnd.n6494 gnd.n6493 585
R4089 gnd.n6496 gnd.n6495 585
R4090 gnd.n6498 gnd.n6497 585
R4091 gnd.n6500 gnd.n6499 585
R4092 gnd.n6502 gnd.n6501 585
R4093 gnd.n6504 gnd.n6503 585
R4094 gnd.n6506 gnd.n6505 585
R4095 gnd.n6507 gnd.n5116 585
R4096 gnd.n6509 gnd.n6508 585
R4097 gnd.n5117 gnd.n5115 585
R4098 gnd.n5118 gnd.n995 585
R4099 gnd.n6511 gnd.n995 585
R4100 gnd.n6409 gnd.n997 585
R4101 gnd.n6512 gnd.n997 585
R4102 gnd.n6413 gnd.n6412 585
R4103 gnd.n6412 gnd.n6411 585
R4104 gnd.n6414 gnd.n986 585
R4105 gnd.n6518 gnd.n986 585
R4106 gnd.n6416 gnd.n6415 585
R4107 gnd.n6417 gnd.n6416 585
R4108 gnd.n6401 gnd.n5173 585
R4109 gnd.n5173 gnd.n976 585
R4110 gnd.n6399 gnd.n974 585
R4111 gnd.n6526 gnd.n974 585
R4112 gnd.n6134 gnd.n5174 585
R4113 gnd.n6135 gnd.n6134 585
R4114 gnd.n5191 gnd.n964 585
R4115 gnd.n6532 gnd.n964 585
R4116 gnd.n6118 gnd.n6117 585
R4117 gnd.n6117 gnd.n5185 585
R4118 gnd.n6116 gnd.n5190 585
R4119 gnd.n6116 gnd.n5184 585
R4120 gnd.n6115 gnd.n5193 585
R4121 gnd.n6115 gnd.n6114 585
R4122 gnd.n6094 gnd.n5192 585
R4123 gnd.n5205 gnd.n5192 585
R4124 gnd.n6093 gnd.n5203 585
R4125 gnd.n6103 gnd.n5203 585
R4126 gnd.n6084 gnd.n5210 585
R4127 gnd.n6085 gnd.n6084 585
R4128 gnd.n6083 gnd.n6082 585
R4129 gnd.n6083 gnd.n5214 585
R4130 gnd.n6081 gnd.n5216 585
R4131 gnd.n6074 gnd.n5216 585
R4132 gnd.n5229 gnd.n5217 585
R4133 gnd.n5229 gnd.n5221 585
R4134 gnd.n6033 gnd.n5230 585
R4135 gnd.n6064 gnd.n5230 585
R4136 gnd.n6032 gnd.n6031 585
R4137 gnd.n6031 gnd.n5237 585
R4138 gnd.n6030 gnd.n5245 585
R4139 gnd.n6030 gnd.n5236 585
R4140 gnd.n6029 gnd.n5247 585
R4141 gnd.n6029 gnd.n6028 585
R4142 gnd.n6008 gnd.n5246 585
R4143 gnd.n5259 gnd.n5246 585
R4144 gnd.n6007 gnd.n5257 585
R4145 gnd.n6018 gnd.n5257 585
R4146 gnd.n5998 gnd.n5264 585
R4147 gnd.n5999 gnd.n5998 585
R4148 gnd.n5997 gnd.n5996 585
R4149 gnd.n5997 gnd.n5268 585
R4150 gnd.n5995 gnd.n5270 585
R4151 gnd.n5988 gnd.n5270 585
R4152 gnd.n5285 gnd.n5271 585
R4153 gnd.n5285 gnd.n5275 585
R4154 gnd.n5948 gnd.n5286 585
R4155 gnd.n5978 gnd.n5286 585
R4156 gnd.n5947 gnd.n5946 585
R4157 gnd.n5946 gnd.n5353 585
R4158 gnd.n5945 gnd.n5360 585
R4159 gnd.n5945 gnd.n5352 585
R4160 gnd.n5944 gnd.n5362 585
R4161 gnd.n5944 gnd.n5943 585
R4162 gnd.n5923 gnd.n5361 585
R4163 gnd.n5374 gnd.n5361 585
R4164 gnd.n5922 gnd.n5372 585
R4165 gnd.n5933 gnd.n5372 585
R4166 gnd.n5913 gnd.n5379 585
R4167 gnd.n5914 gnd.n5913 585
R4168 gnd.n5912 gnd.n5911 585
R4169 gnd.n5912 gnd.n5383 585
R4170 gnd.n5910 gnd.n5385 585
R4171 gnd.n5903 gnd.n5385 585
R4172 gnd.n5890 gnd.n5386 585
R4173 gnd.n5891 gnd.n5890 585
R4174 gnd.n5860 gnd.n5399 585
R4175 gnd.n5893 gnd.n5399 585
R4176 gnd.n5859 gnd.n5858 585
R4177 gnd.n5858 gnd.n5857 585
R4178 gnd.n5855 gnd.n5416 585
R4179 gnd.n5855 gnd.n5407 585
R4180 gnd.n5854 gnd.n5853 585
R4181 gnd.n5854 gnd.n5406 585
R4182 gnd.n5418 gnd.n5417 585
R4183 gnd.n5845 gnd.n5417 585
R4184 gnd.n5814 gnd.n5813 585
R4185 gnd.n5813 gnd.n5422 585
R4186 gnd.n5815 gnd.n5432 585
R4187 gnd.n5832 gnd.n5432 585
R4188 gnd.n5812 gnd.n5811 585
R4189 gnd.n5811 gnd.n5439 585
R4190 gnd.n5810 gnd.n5446 585
R4191 gnd.n5810 gnd.n5438 585
R4192 gnd.n5809 gnd.n5448 585
R4193 gnd.n5809 gnd.n5808 585
R4194 gnd.n5788 gnd.n5447 585
R4195 gnd.n5460 gnd.n5447 585
R4196 gnd.n5787 gnd.n5458 585
R4197 gnd.n5798 gnd.n5458 585
R4198 gnd.n5778 gnd.n5465 585
R4199 gnd.n5779 gnd.n5778 585
R4200 gnd.n5777 gnd.n5471 585
R4201 gnd.n5777 gnd.n5776 585
R4202 gnd.n5762 gnd.n5470 585
R4203 gnd.n5481 gnd.n5470 585
R4204 gnd.n5761 gnd.n5479 585
R4205 gnd.n5768 gnd.n5479 585
R4206 gnd.n5760 gnd.n5759 585
R4207 gnd.n5759 gnd.n5758 585
R4208 gnd.n4834 gnd.n1406 585
R4209 gnd.n3329 gnd.n1406 585
R4210 gnd.n4836 gnd.n4835 585
R4211 gnd.n4837 gnd.n4836 585
R4212 gnd.n1390 gnd.n1389 585
R4213 gnd.n3258 gnd.n1390 585
R4214 gnd.n4845 gnd.n4844 585
R4215 gnd.n4844 gnd.n4843 585
R4216 gnd.n4846 gnd.n1384 585
R4217 gnd.n3188 gnd.n1384 585
R4218 gnd.n4848 gnd.n4847 585
R4219 gnd.n4849 gnd.n4848 585
R4220 gnd.n1369 gnd.n1368 585
R4221 gnd.n3196 gnd.n1369 585
R4222 gnd.n4857 gnd.n4856 585
R4223 gnd.n4856 gnd.n4855 585
R4224 gnd.n4858 gnd.n1363 585
R4225 gnd.n3178 gnd.n1363 585
R4226 gnd.n4860 gnd.n4859 585
R4227 gnd.n4861 gnd.n4860 585
R4228 gnd.n1347 gnd.n1346 585
R4229 gnd.n3170 gnd.n1347 585
R4230 gnd.n4869 gnd.n4868 585
R4231 gnd.n4868 gnd.n4867 585
R4232 gnd.n4870 gnd.n1341 585
R4233 gnd.n3161 gnd.n1341 585
R4234 gnd.n4872 gnd.n4871 585
R4235 gnd.n4873 gnd.n4872 585
R4236 gnd.n1327 gnd.n1326 585
R4237 gnd.n3153 gnd.n1327 585
R4238 gnd.n4881 gnd.n4880 585
R4239 gnd.n4880 gnd.n4879 585
R4240 gnd.n4882 gnd.n1321 585
R4241 gnd.n3145 gnd.n1321 585
R4242 gnd.n4884 gnd.n4883 585
R4243 gnd.n4885 gnd.n4884 585
R4244 gnd.n1305 gnd.n1304 585
R4245 gnd.n3137 gnd.n1305 585
R4246 gnd.n4893 gnd.n4892 585
R4247 gnd.n4892 gnd.n4891 585
R4248 gnd.n4894 gnd.n1299 585
R4249 gnd.n3129 gnd.n1299 585
R4250 gnd.n4896 gnd.n4895 585
R4251 gnd.n4897 gnd.n4896 585
R4252 gnd.n1285 gnd.n1284 585
R4253 gnd.n3121 gnd.n1285 585
R4254 gnd.n4905 gnd.n4904 585
R4255 gnd.n4904 gnd.n4903 585
R4256 gnd.n4906 gnd.n1279 585
R4257 gnd.n3113 gnd.n1279 585
R4258 gnd.n4908 gnd.n4907 585
R4259 gnd.n4909 gnd.n4908 585
R4260 gnd.n1263 gnd.n1262 585
R4261 gnd.n3105 gnd.n1263 585
R4262 gnd.n4917 gnd.n4916 585
R4263 gnd.n4916 gnd.n4915 585
R4264 gnd.n4918 gnd.n1260 585
R4265 gnd.n3097 gnd.n1260 585
R4266 gnd.n4921 gnd.n4920 585
R4267 gnd.n4922 gnd.n4921 585
R4268 gnd.n1261 gnd.n1246 585
R4269 gnd.n3089 gnd.n1246 585
R4270 gnd.n4930 gnd.n4929 585
R4271 gnd.n4929 gnd.n4928 585
R4272 gnd.n4931 gnd.n1243 585
R4273 gnd.n3081 gnd.n1243 585
R4274 gnd.n4934 gnd.n4933 585
R4275 gnd.n4935 gnd.n4934 585
R4276 gnd.n1244 gnd.n1227 585
R4277 gnd.n3073 gnd.n1227 585
R4278 gnd.n4943 gnd.n4942 585
R4279 gnd.n4942 gnd.n4941 585
R4280 gnd.n4944 gnd.n1223 585
R4281 gnd.n3065 gnd.n1223 585
R4282 gnd.n4947 gnd.n4946 585
R4283 gnd.n4948 gnd.n4947 585
R4284 gnd.n1208 gnd.n1207 585
R4285 gnd.n3057 gnd.n1208 585
R4286 gnd.n4956 gnd.n4955 585
R4287 gnd.n4955 gnd.n4954 585
R4288 gnd.n4957 gnd.n1202 585
R4289 gnd.n3049 gnd.n1202 585
R4290 gnd.n4959 gnd.n4958 585
R4291 gnd.n4960 gnd.n4959 585
R4292 gnd.n1186 gnd.n1185 585
R4293 gnd.n3041 gnd.n1186 585
R4294 gnd.n4968 gnd.n4967 585
R4295 gnd.n4967 gnd.n4966 585
R4296 gnd.n4969 gnd.n1180 585
R4297 gnd.n3033 gnd.n1180 585
R4298 gnd.n4971 gnd.n4970 585
R4299 gnd.n4972 gnd.n4971 585
R4300 gnd.n1166 gnd.n1165 585
R4301 gnd.n1176 gnd.n1166 585
R4302 gnd.n4980 gnd.n4979 585
R4303 gnd.n4979 gnd.n4978 585
R4304 gnd.n4981 gnd.n1160 585
R4305 gnd.n1160 gnd.n1159 585
R4306 gnd.n4983 gnd.n4982 585
R4307 gnd.n4984 gnd.n4983 585
R4308 gnd.n1146 gnd.n1145 585
R4309 gnd.n1149 gnd.n1146 585
R4310 gnd.n4992 gnd.n4991 585
R4311 gnd.n4991 gnd.n4990 585
R4312 gnd.n4993 gnd.n1140 585
R4313 gnd.n1140 gnd.n1139 585
R4314 gnd.n4995 gnd.n4994 585
R4315 gnd.n4996 gnd.n4995 585
R4316 gnd.n1126 gnd.n1125 585
R4317 gnd.n1136 gnd.n1126 585
R4318 gnd.n5004 gnd.n5003 585
R4319 gnd.n5003 gnd.n5002 585
R4320 gnd.n5005 gnd.n1120 585
R4321 gnd.n1120 gnd.n1119 585
R4322 gnd.n5007 gnd.n5006 585
R4323 gnd.n5008 gnd.n5007 585
R4324 gnd.n1105 gnd.n1104 585
R4325 gnd.n1108 gnd.n1105 585
R4326 gnd.n5016 gnd.n5015 585
R4327 gnd.n5015 gnd.n5014 585
R4328 gnd.n5017 gnd.n1099 585
R4329 gnd.n1099 gnd.n1096 585
R4330 gnd.n5019 gnd.n5018 585
R4331 gnd.n5020 gnd.n5019 585
R4332 gnd.n1100 gnd.n1098 585
R4333 gnd.n1098 gnd.n1094 585
R4334 gnd.n2991 gnd.n2990 585
R4335 gnd.n2992 gnd.n2991 585
R4336 gnd.n2986 gnd.n1043 585
R4337 gnd.n1043 gnd.n1040 585
R4338 gnd.n5105 gnd.n5104 585
R4339 gnd.n5103 gnd.n1042 585
R4340 gnd.n5102 gnd.n1041 585
R4341 gnd.n5107 gnd.n1041 585
R4342 gnd.n5101 gnd.n5100 585
R4343 gnd.n5099 gnd.n5098 585
R4344 gnd.n5097 gnd.n5096 585
R4345 gnd.n5095 gnd.n5094 585
R4346 gnd.n5093 gnd.n5092 585
R4347 gnd.n5091 gnd.n5090 585
R4348 gnd.n5089 gnd.n5088 585
R4349 gnd.n5087 gnd.n5086 585
R4350 gnd.n5085 gnd.n5084 585
R4351 gnd.n5083 gnd.n5082 585
R4352 gnd.n5081 gnd.n5080 585
R4353 gnd.n5079 gnd.n5078 585
R4354 gnd.n5077 gnd.n5076 585
R4355 gnd.n5075 gnd.n5074 585
R4356 gnd.n5073 gnd.n5072 585
R4357 gnd.n5070 gnd.n5069 585
R4358 gnd.n5068 gnd.n5067 585
R4359 gnd.n5066 gnd.n5065 585
R4360 gnd.n5064 gnd.n5063 585
R4361 gnd.n5062 gnd.n5061 585
R4362 gnd.n5060 gnd.n5059 585
R4363 gnd.n5058 gnd.n5057 585
R4364 gnd.n5056 gnd.n5055 585
R4365 gnd.n5054 gnd.n5053 585
R4366 gnd.n5052 gnd.n5051 585
R4367 gnd.n5050 gnd.n5049 585
R4368 gnd.n5048 gnd.n5047 585
R4369 gnd.n5046 gnd.n5045 585
R4370 gnd.n5044 gnd.n5043 585
R4371 gnd.n5042 gnd.n5041 585
R4372 gnd.n5040 gnd.n5039 585
R4373 gnd.n5038 gnd.n5037 585
R4374 gnd.n5036 gnd.n5035 585
R4375 gnd.n5034 gnd.n1082 585
R4376 gnd.n1086 gnd.n1083 585
R4377 gnd.n5030 gnd.n5029 585
R4378 gnd.n3324 gnd.n2624 585
R4379 gnd.n3323 gnd.n3266 585
R4380 gnd.n3322 gnd.n3321 585
R4381 gnd.n3315 gnd.n3267 585
R4382 gnd.n3317 gnd.n3316 585
R4383 gnd.n3314 gnd.n3313 585
R4384 gnd.n3312 gnd.n3311 585
R4385 gnd.n3305 gnd.n3269 585
R4386 gnd.n3307 gnd.n3306 585
R4387 gnd.n3304 gnd.n3303 585
R4388 gnd.n3302 gnd.n3301 585
R4389 gnd.n3295 gnd.n3271 585
R4390 gnd.n3297 gnd.n3296 585
R4391 gnd.n3294 gnd.n3293 585
R4392 gnd.n3292 gnd.n3291 585
R4393 gnd.n3285 gnd.n3273 585
R4394 gnd.n3287 gnd.n3286 585
R4395 gnd.n3284 gnd.n3283 585
R4396 gnd.n3282 gnd.n3281 585
R4397 gnd.n3277 gnd.n3276 585
R4398 gnd.n3275 gnd.n1457 585
R4399 gnd.n4802 gnd.n4801 585
R4400 gnd.n4804 gnd.n4803 585
R4401 gnd.n4806 gnd.n4805 585
R4402 gnd.n4808 gnd.n4807 585
R4403 gnd.n4810 gnd.n4809 585
R4404 gnd.n4812 gnd.n4811 585
R4405 gnd.n4814 gnd.n4813 585
R4406 gnd.n4816 gnd.n4815 585
R4407 gnd.n4818 gnd.n4817 585
R4408 gnd.n4820 gnd.n4819 585
R4409 gnd.n4822 gnd.n4821 585
R4410 gnd.n4824 gnd.n4823 585
R4411 gnd.n4825 gnd.n1442 585
R4412 gnd.n4827 gnd.n4826 585
R4413 gnd.n1411 gnd.n1410 585
R4414 gnd.n4831 gnd.n4830 585
R4415 gnd.n4830 gnd.n4829 585
R4416 gnd.n3328 gnd.n3327 585
R4417 gnd.n3329 gnd.n3328 585
R4418 gnd.n2625 gnd.n1403 585
R4419 gnd.n4837 gnd.n1403 585
R4420 gnd.n3260 gnd.n3259 585
R4421 gnd.n3259 gnd.n3258 585
R4422 gnd.n2627 gnd.n1392 585
R4423 gnd.n4843 gnd.n1392 585
R4424 gnd.n3187 gnd.n3186 585
R4425 gnd.n3188 gnd.n3187 585
R4426 gnd.n2692 gnd.n1381 585
R4427 gnd.n4849 gnd.n1381 585
R4428 gnd.n3182 gnd.n2688 585
R4429 gnd.n3196 gnd.n2688 585
R4430 gnd.n3181 gnd.n1371 585
R4431 gnd.n4855 gnd.n1371 585
R4432 gnd.n3180 gnd.n3179 585
R4433 gnd.n3179 gnd.n3178 585
R4434 gnd.n2694 gnd.n1360 585
R4435 gnd.n4861 gnd.n1360 585
R4436 gnd.n3169 gnd.n3168 585
R4437 gnd.n3170 gnd.n3169 585
R4438 gnd.n2699 gnd.n1349 585
R4439 gnd.n4867 gnd.n1349 585
R4440 gnd.n3163 gnd.n3162 585
R4441 gnd.n3162 gnd.n3161 585
R4442 gnd.n2701 gnd.n1339 585
R4443 gnd.n4873 gnd.n1339 585
R4444 gnd.n3152 gnd.n3151 585
R4445 gnd.n3153 gnd.n3152 585
R4446 gnd.n2707 gnd.n1329 585
R4447 gnd.n4879 gnd.n1329 585
R4448 gnd.n3147 gnd.n3146 585
R4449 gnd.n3146 gnd.n3145 585
R4450 gnd.n2709 gnd.n1318 585
R4451 gnd.n4885 gnd.n1318 585
R4452 gnd.n3136 gnd.n3135 585
R4453 gnd.n3137 gnd.n3136 585
R4454 gnd.n2713 gnd.n1307 585
R4455 gnd.n4891 gnd.n1307 585
R4456 gnd.n3131 gnd.n3130 585
R4457 gnd.n3130 gnd.n3129 585
R4458 gnd.n2715 gnd.n1297 585
R4459 gnd.n4897 gnd.n1297 585
R4460 gnd.n3120 gnd.n3119 585
R4461 gnd.n3121 gnd.n3120 585
R4462 gnd.n2721 gnd.n1287 585
R4463 gnd.n4903 gnd.n1287 585
R4464 gnd.n3115 gnd.n3114 585
R4465 gnd.n3114 gnd.n3113 585
R4466 gnd.n2723 gnd.n1276 585
R4467 gnd.n4909 gnd.n1276 585
R4468 gnd.n3104 gnd.n3103 585
R4469 gnd.n3105 gnd.n3104 585
R4470 gnd.n2727 gnd.n1265 585
R4471 gnd.n4915 gnd.n1265 585
R4472 gnd.n3099 gnd.n3098 585
R4473 gnd.n3098 gnd.n3097 585
R4474 gnd.n2729 gnd.n1257 585
R4475 gnd.n4922 gnd.n1257 585
R4476 gnd.n3088 gnd.n3087 585
R4477 gnd.n3089 gnd.n3088 585
R4478 gnd.n2734 gnd.n1248 585
R4479 gnd.n4928 gnd.n1248 585
R4480 gnd.n3083 gnd.n3082 585
R4481 gnd.n3082 gnd.n3081 585
R4482 gnd.n2737 gnd.n1240 585
R4483 gnd.n4935 gnd.n1240 585
R4484 gnd.n3072 gnd.n3071 585
R4485 gnd.n3073 gnd.n3072 585
R4486 gnd.n2741 gnd.n1229 585
R4487 gnd.n4941 gnd.n1229 585
R4488 gnd.n3067 gnd.n3066 585
R4489 gnd.n3066 gnd.n3065 585
R4490 gnd.n2743 gnd.n1220 585
R4491 gnd.n4948 gnd.n1220 585
R4492 gnd.n3056 gnd.n3055 585
R4493 gnd.n3057 gnd.n3056 585
R4494 gnd.n2858 gnd.n1210 585
R4495 gnd.n4954 gnd.n1210 585
R4496 gnd.n3051 gnd.n3050 585
R4497 gnd.n3050 gnd.n3049 585
R4498 gnd.n2860 gnd.n1199 585
R4499 gnd.n4960 gnd.n1199 585
R4500 gnd.n3040 gnd.n3039 585
R4501 gnd.n3041 gnd.n3040 585
R4502 gnd.n2864 gnd.n1188 585
R4503 gnd.n4966 gnd.n1188 585
R4504 gnd.n3035 gnd.n3034 585
R4505 gnd.n3034 gnd.n3033 585
R4506 gnd.n2901 gnd.n1177 585
R4507 gnd.n4972 gnd.n1177 585
R4508 gnd.n2900 gnd.n2899 585
R4509 gnd.n2899 gnd.n1176 585
R4510 gnd.n2866 gnd.n1167 585
R4511 gnd.n4978 gnd.n1167 585
R4512 gnd.n2895 gnd.n2894 585
R4513 gnd.n2894 gnd.n1159 585
R4514 gnd.n2893 gnd.n1157 585
R4515 gnd.n4984 gnd.n1157 585
R4516 gnd.n2892 gnd.n2891 585
R4517 gnd.n2891 gnd.n1149 585
R4518 gnd.n2868 gnd.n1147 585
R4519 gnd.n4990 gnd.n1147 585
R4520 gnd.n2887 gnd.n2886 585
R4521 gnd.n2886 gnd.n1139 585
R4522 gnd.n2885 gnd.n1137 585
R4523 gnd.n4996 gnd.n1137 585
R4524 gnd.n2884 gnd.n2883 585
R4525 gnd.n2883 gnd.n1136 585
R4526 gnd.n2870 gnd.n1127 585
R4527 gnd.n5002 gnd.n1127 585
R4528 gnd.n2879 gnd.n2878 585
R4529 gnd.n2878 gnd.n1119 585
R4530 gnd.n2877 gnd.n1117 585
R4531 gnd.n5008 gnd.n1117 585
R4532 gnd.n2876 gnd.n2875 585
R4533 gnd.n2875 gnd.n1108 585
R4534 gnd.n2872 gnd.n1106 585
R4535 gnd.n5014 gnd.n1106 585
R4536 gnd.n1093 gnd.n1091 585
R4537 gnd.n1096 gnd.n1093 585
R4538 gnd.n5022 gnd.n5021 585
R4539 gnd.n5021 gnd.n5020 585
R4540 gnd.n1092 gnd.n1089 585
R4541 gnd.n1094 gnd.n1092 585
R4542 gnd.n5026 gnd.n1088 585
R4543 gnd.n2992 gnd.n1088 585
R4544 gnd.n5028 gnd.n5027 585
R4545 gnd.n5028 gnd.n1040 585
R4546 gnd.n7665 gnd.n7664 585
R4547 gnd.n7666 gnd.n7665 585
R4548 gnd.n128 gnd.n126 585
R4549 gnd.n126 gnd.n122 585
R4550 gnd.n7585 gnd.n7584 585
R4551 gnd.n7586 gnd.n7585 585
R4552 gnd.n205 gnd.n204 585
R4553 gnd.n212 gnd.n204 585
R4554 gnd.n7580 gnd.n7579 585
R4555 gnd.n7579 gnd.n7578 585
R4556 gnd.n208 gnd.n207 585
R4557 gnd.n209 gnd.n208 585
R4558 gnd.n7501 gnd.n7500 585
R4559 gnd.n7502 gnd.n7501 585
R4560 gnd.n222 gnd.n221 585
R4561 gnd.n229 gnd.n221 585
R4562 gnd.n7496 gnd.n7495 585
R4563 gnd.n7495 gnd.n7494 585
R4564 gnd.n225 gnd.n224 585
R4565 gnd.n226 gnd.n225 585
R4566 gnd.n7485 gnd.n7484 585
R4567 gnd.n7486 gnd.n7485 585
R4568 gnd.n238 gnd.n237 585
R4569 gnd.n237 gnd.n235 585
R4570 gnd.n7480 gnd.n7479 585
R4571 gnd.n7479 gnd.n7478 585
R4572 gnd.n241 gnd.n240 585
R4573 gnd.n250 gnd.n241 585
R4574 gnd.n7469 gnd.n7468 585
R4575 gnd.n7470 gnd.n7469 585
R4576 gnd.n252 gnd.n251 585
R4577 gnd.n259 gnd.n251 585
R4578 gnd.n7464 gnd.n7463 585
R4579 gnd.n7463 gnd.n7462 585
R4580 gnd.n255 gnd.n254 585
R4581 gnd.n256 gnd.n255 585
R4582 gnd.n7453 gnd.n7452 585
R4583 gnd.n7454 gnd.n7453 585
R4584 gnd.n268 gnd.n267 585
R4585 gnd.n267 gnd.n265 585
R4586 gnd.n7448 gnd.n7447 585
R4587 gnd.n7447 gnd.n7446 585
R4588 gnd.n271 gnd.n270 585
R4589 gnd.n7373 gnd.n271 585
R4590 gnd.n7437 gnd.n7436 585
R4591 gnd.n7438 gnd.n7437 585
R4592 gnd.n283 gnd.n282 585
R4593 gnd.n7379 gnd.n282 585
R4594 gnd.n7432 gnd.n7431 585
R4595 gnd.n7431 gnd.n7430 585
R4596 gnd.n286 gnd.n285 585
R4597 gnd.n4511 gnd.n286 585
R4598 gnd.n7421 gnd.n7420 585
R4599 gnd.n7422 gnd.n7421 585
R4600 gnd.n300 gnd.n299 585
R4601 gnd.n4515 gnd.n299 585
R4602 gnd.n7397 gnd.n7396 585
R4603 gnd.n7398 gnd.n7397 585
R4604 gnd.n7395 gnd.n331 585
R4605 gnd.n7395 gnd.n7394 585
R4606 gnd.n330 gnd.n329 585
R4607 gnd.n4523 gnd.n329 585
R4608 gnd.n1701 gnd.n1700 585
R4609 gnd.n1704 gnd.n1700 585
R4610 gnd.n4543 gnd.n1702 585
R4611 gnd.n4543 gnd.n4542 585
R4612 gnd.n4546 gnd.n4545 585
R4613 gnd.n4547 gnd.n4546 585
R4614 gnd.n4544 gnd.n309 585
R4615 gnd.n4531 gnd.n309 585
R4616 gnd.n7415 gnd.n7414 585
R4617 gnd.n7414 gnd.n7413 585
R4618 gnd.n7416 gnd.n308 585
R4619 gnd.n4495 gnd.n308 585
R4620 gnd.n4561 gnd.n307 585
R4621 gnd.n4562 gnd.n4561 585
R4622 gnd.n4560 gnd.n1688 585
R4623 gnd.n4560 gnd.n4559 585
R4624 gnd.n4484 gnd.n1687 585
R4625 gnd.n4468 gnd.n1687 585
R4626 gnd.n4486 gnd.n4485 585
R4627 gnd.n4487 gnd.n4486 585
R4628 gnd.n1721 gnd.n1720 585
R4629 gnd.n4439 gnd.n1720 585
R4630 gnd.n4479 gnd.n4478 585
R4631 gnd.n4478 gnd.n4477 585
R4632 gnd.n1724 gnd.n1723 585
R4633 gnd.n4448 gnd.n1724 585
R4634 gnd.n4430 gnd.n1747 585
R4635 gnd.n1747 gnd.n1735 585
R4636 gnd.n4432 gnd.n4431 585
R4637 gnd.n4433 gnd.n4432 585
R4638 gnd.n1748 gnd.n1746 585
R4639 gnd.n4313 gnd.n1746 585
R4640 gnd.n4425 gnd.n4424 585
R4641 gnd.n4424 gnd.n4423 585
R4642 gnd.n1751 gnd.n1750 585
R4643 gnd.n4411 gnd.n1751 585
R4644 gnd.n4398 gnd.n1773 585
R4645 gnd.n1773 gnd.n1761 585
R4646 gnd.n4400 gnd.n4399 585
R4647 gnd.n4401 gnd.n4400 585
R4648 gnd.n1774 gnd.n1772 585
R4649 gnd.n4321 gnd.n1772 585
R4650 gnd.n4393 gnd.n4392 585
R4651 gnd.n4392 gnd.n4391 585
R4652 gnd.n1777 gnd.n1776 585
R4653 gnd.n4378 gnd.n1777 585
R4654 gnd.n4366 gnd.n1799 585
R4655 gnd.n1799 gnd.n1787 585
R4656 gnd.n4368 gnd.n4367 585
R4657 gnd.n4369 gnd.n4368 585
R4658 gnd.n1800 gnd.n1798 585
R4659 gnd.n1807 gnd.n1798 585
R4660 gnd.n4361 gnd.n4360 585
R4661 gnd.n4360 gnd.n4359 585
R4662 gnd.n1803 gnd.n1802 585
R4663 gnd.n4347 gnd.n1803 585
R4664 gnd.n1824 gnd.n1823 585
R4665 gnd.n1825 gnd.n1824 585
R4666 gnd.n1645 gnd.n1644 585
R4667 gnd.n4337 gnd.n1645 585
R4668 gnd.n4605 gnd.n4604 585
R4669 gnd.n4604 gnd.n4603 585
R4670 gnd.n4606 gnd.n1639 585
R4671 gnd.n4284 gnd.n1639 585
R4672 gnd.n4608 gnd.n4607 585
R4673 gnd.n4609 gnd.n4608 585
R4674 gnd.n1640 gnd.n1638 585
R4675 gnd.n1638 gnd.n1633 585
R4676 gnd.n2098 gnd.n2097 585
R4677 gnd.n2101 gnd.n2100 585
R4678 gnd.n2094 gnd.n2093 585
R4679 gnd.n2093 gnd.n1624 585
R4680 gnd.n2106 gnd.n2105 585
R4681 gnd.n2108 gnd.n2092 585
R4682 gnd.n2111 gnd.n2110 585
R4683 gnd.n2090 gnd.n2089 585
R4684 gnd.n2116 gnd.n2115 585
R4685 gnd.n2118 gnd.n2088 585
R4686 gnd.n2121 gnd.n2120 585
R4687 gnd.n2086 gnd.n2085 585
R4688 gnd.n2127 gnd.n2126 585
R4689 gnd.n2129 gnd.n2084 585
R4690 gnd.n2130 gnd.n2081 585
R4691 gnd.n2133 gnd.n2132 585
R4692 gnd.n2083 gnd.n2078 585
R4693 gnd.n2217 gnd.n2216 585
R4694 gnd.n2214 gnd.n2140 585
R4695 gnd.n2212 gnd.n2211 585
R4696 gnd.n2210 gnd.n2141 585
R4697 gnd.n2209 gnd.n2208 585
R4698 gnd.n2206 gnd.n2146 585
R4699 gnd.n2204 gnd.n2203 585
R4700 gnd.n2202 gnd.n2147 585
R4701 gnd.n2201 gnd.n2200 585
R4702 gnd.n2198 gnd.n2152 585
R4703 gnd.n2196 gnd.n2195 585
R4704 gnd.n2194 gnd.n2153 585
R4705 gnd.n2193 gnd.n2192 585
R4706 gnd.n2190 gnd.n2158 585
R4707 gnd.n2188 gnd.n2187 585
R4708 gnd.n2186 gnd.n2159 585
R4709 gnd.n2185 gnd.n2184 585
R4710 gnd.n2182 gnd.n2164 585
R4711 gnd.n2180 gnd.n2179 585
R4712 gnd.n2168 gnd.n2165 585
R4713 gnd.n2175 gnd.n2174 585
R4714 gnd.n196 gnd.n195 585
R4715 gnd.n7594 gnd.n191 585
R4716 gnd.n7596 gnd.n7595 585
R4717 gnd.n7598 gnd.n189 585
R4718 gnd.n7600 gnd.n7599 585
R4719 gnd.n7601 gnd.n184 585
R4720 gnd.n7603 gnd.n7602 585
R4721 gnd.n7605 gnd.n182 585
R4722 gnd.n7607 gnd.n7606 585
R4723 gnd.n7608 gnd.n177 585
R4724 gnd.n7610 gnd.n7609 585
R4725 gnd.n7612 gnd.n175 585
R4726 gnd.n7614 gnd.n7613 585
R4727 gnd.n7615 gnd.n170 585
R4728 gnd.n7617 gnd.n7616 585
R4729 gnd.n7619 gnd.n168 585
R4730 gnd.n7621 gnd.n7620 585
R4731 gnd.n7622 gnd.n163 585
R4732 gnd.n7624 gnd.n7623 585
R4733 gnd.n7626 gnd.n161 585
R4734 gnd.n7628 gnd.n7627 585
R4735 gnd.n7632 gnd.n156 585
R4736 gnd.n7634 gnd.n7633 585
R4737 gnd.n7636 gnd.n154 585
R4738 gnd.n7638 gnd.n7637 585
R4739 gnd.n7639 gnd.n149 585
R4740 gnd.n7641 gnd.n7640 585
R4741 gnd.n7643 gnd.n147 585
R4742 gnd.n7645 gnd.n7644 585
R4743 gnd.n7646 gnd.n142 585
R4744 gnd.n7648 gnd.n7647 585
R4745 gnd.n7650 gnd.n140 585
R4746 gnd.n7652 gnd.n7651 585
R4747 gnd.n7653 gnd.n135 585
R4748 gnd.n7655 gnd.n7654 585
R4749 gnd.n7657 gnd.n133 585
R4750 gnd.n7659 gnd.n7658 585
R4751 gnd.n7660 gnd.n131 585
R4752 gnd.n7661 gnd.n127 585
R4753 gnd.n127 gnd.n124 585
R4754 gnd.n7590 gnd.n123 585
R4755 gnd.n7666 gnd.n123 585
R4756 gnd.n7589 gnd.n7588 585
R4757 gnd.n7588 gnd.n122 585
R4758 gnd.n7587 gnd.n200 585
R4759 gnd.n7587 gnd.n7586 585
R4760 gnd.n369 gnd.n201 585
R4761 gnd.n212 gnd.n201 585
R4762 gnd.n370 gnd.n210 585
R4763 gnd.n7578 gnd.n210 585
R4764 gnd.n372 gnd.n371 585
R4765 gnd.n371 gnd.n209 585
R4766 gnd.n373 gnd.n220 585
R4767 gnd.n7502 gnd.n220 585
R4768 gnd.n375 gnd.n374 585
R4769 gnd.n374 gnd.n229 585
R4770 gnd.n376 gnd.n227 585
R4771 gnd.n7494 gnd.n227 585
R4772 gnd.n378 gnd.n377 585
R4773 gnd.n377 gnd.n226 585
R4774 gnd.n379 gnd.n236 585
R4775 gnd.n7486 gnd.n236 585
R4776 gnd.n381 gnd.n380 585
R4777 gnd.n380 gnd.n235 585
R4778 gnd.n382 gnd.n242 585
R4779 gnd.n7478 gnd.n242 585
R4780 gnd.n384 gnd.n383 585
R4781 gnd.n383 gnd.n250 585
R4782 gnd.n385 gnd.n249 585
R4783 gnd.n7470 gnd.n249 585
R4784 gnd.n387 gnd.n386 585
R4785 gnd.n386 gnd.n259 585
R4786 gnd.n388 gnd.n257 585
R4787 gnd.n7462 gnd.n257 585
R4788 gnd.n390 gnd.n389 585
R4789 gnd.n389 gnd.n256 585
R4790 gnd.n391 gnd.n266 585
R4791 gnd.n7454 gnd.n266 585
R4792 gnd.n393 gnd.n392 585
R4793 gnd.n392 gnd.n265 585
R4794 gnd.n394 gnd.n272 585
R4795 gnd.n7446 gnd.n272 585
R4796 gnd.n7375 gnd.n7374 585
R4797 gnd.n7374 gnd.n7373 585
R4798 gnd.n7376 gnd.n280 585
R4799 gnd.n7438 gnd.n280 585
R4800 gnd.n7378 gnd.n7377 585
R4801 gnd.n7379 gnd.n7378 585
R4802 gnd.n346 gnd.n288 585
R4803 gnd.n7430 gnd.n288 585
R4804 gnd.n4513 gnd.n4512 585
R4805 gnd.n4512 gnd.n4511 585
R4806 gnd.n4514 gnd.n297 585
R4807 gnd.n7422 gnd.n297 585
R4808 gnd.n4517 gnd.n4516 585
R4809 gnd.n4516 gnd.n4515 585
R4810 gnd.n4518 gnd.n326 585
R4811 gnd.n7398 gnd.n326 585
R4812 gnd.n4519 gnd.n333 585
R4813 gnd.n7394 gnd.n333 585
R4814 gnd.n4524 gnd.n4520 585
R4815 gnd.n4524 gnd.n4523 585
R4816 gnd.n4526 gnd.n4525 585
R4817 gnd.n4525 gnd.n1704 585
R4818 gnd.n4527 gnd.n1703 585
R4819 gnd.n4542 gnd.n1703 585
R4820 gnd.n4528 gnd.n1698 585
R4821 gnd.n4547 gnd.n1698 585
R4822 gnd.n4530 gnd.n4529 585
R4823 gnd.n4531 gnd.n4530 585
R4824 gnd.n1709 gnd.n311 585
R4825 gnd.n7413 gnd.n311 585
R4826 gnd.n4497 gnd.n4496 585
R4827 gnd.n4496 gnd.n4495 585
R4828 gnd.n4494 gnd.n1684 585
R4829 gnd.n4562 gnd.n1684 585
R4830 gnd.n4493 gnd.n1689 585
R4831 gnd.n4559 gnd.n1689 585
R4832 gnd.n1715 gnd.n1711 585
R4833 gnd.n4468 gnd.n1715 585
R4834 gnd.n4489 gnd.n4488 585
R4835 gnd.n4488 gnd.n4487 585
R4836 gnd.n1714 gnd.n1713 585
R4837 gnd.n4439 gnd.n1714 585
R4838 gnd.n4308 gnd.n1726 585
R4839 gnd.n4477 gnd.n1726 585
R4840 gnd.n4309 gnd.n1736 585
R4841 gnd.n4448 gnd.n1736 585
R4842 gnd.n4311 gnd.n4310 585
R4843 gnd.n4310 gnd.n1735 585
R4844 gnd.n4312 gnd.n1744 585
R4845 gnd.n4433 gnd.n1744 585
R4846 gnd.n4315 gnd.n4314 585
R4847 gnd.n4314 gnd.n4313 585
R4848 gnd.n4316 gnd.n1753 585
R4849 gnd.n4423 gnd.n1753 585
R4850 gnd.n4317 gnd.n1762 585
R4851 gnd.n4411 gnd.n1762 585
R4852 gnd.n4319 gnd.n4318 585
R4853 gnd.n4318 gnd.n1761 585
R4854 gnd.n4320 gnd.n1770 585
R4855 gnd.n4401 gnd.n1770 585
R4856 gnd.n4323 gnd.n4322 585
R4857 gnd.n4322 gnd.n4321 585
R4858 gnd.n4324 gnd.n1779 585
R4859 gnd.n4391 gnd.n1779 585
R4860 gnd.n4325 gnd.n1788 585
R4861 gnd.n4378 gnd.n1788 585
R4862 gnd.n4327 gnd.n4326 585
R4863 gnd.n4326 gnd.n1787 585
R4864 gnd.n4328 gnd.n1796 585
R4865 gnd.n4369 gnd.n1796 585
R4866 gnd.n4330 gnd.n4329 585
R4867 gnd.n4329 gnd.n1807 585
R4868 gnd.n4331 gnd.n1804 585
R4869 gnd.n4359 gnd.n1804 585
R4870 gnd.n4332 gnd.n1826 585
R4871 gnd.n4347 gnd.n1826 585
R4872 gnd.n4333 gnd.n1832 585
R4873 gnd.n1832 gnd.n1825 585
R4874 gnd.n4335 gnd.n4334 585
R4875 gnd.n4337 gnd.n4335 585
R4876 gnd.n1833 gnd.n1647 585
R4877 gnd.n4603 gnd.n1647 585
R4878 gnd.n4286 gnd.n4285 585
R4879 gnd.n4285 gnd.n4284 585
R4880 gnd.n1835 gnd.n1634 585
R4881 gnd.n4609 gnd.n1634 585
R4882 gnd.n2172 gnd.n2171 585
R4883 gnd.n2172 gnd.n1633 585
R4884 gnd.n4090 gnd.n2227 585
R4885 gnd.n2227 gnd.n2043 585
R4886 gnd.n4092 gnd.n4091 585
R4887 gnd.n4093 gnd.n4092 585
R4888 gnd.n4001 gnd.n2226 585
R4889 gnd.n3995 gnd.n2226 585
R4890 gnd.n4000 gnd.n3999 585
R4891 gnd.n3999 gnd.n3998 585
R4892 gnd.n2229 gnd.n2228 585
R4893 gnd.n3982 gnd.n2229 585
R4894 gnd.n3971 gnd.n2247 585
R4895 gnd.n2247 gnd.n2239 585
R4896 gnd.n3973 gnd.n3972 585
R4897 gnd.n3974 gnd.n3973 585
R4898 gnd.n3970 gnd.n2246 585
R4899 gnd.n3933 gnd.n2246 585
R4900 gnd.n3969 gnd.n3968 585
R4901 gnd.n3968 gnd.n3967 585
R4902 gnd.n2249 gnd.n2248 585
R4903 gnd.n2297 gnd.n2249 585
R4904 gnd.n3956 gnd.n3955 585
R4905 gnd.n3957 gnd.n3956 585
R4906 gnd.n3954 gnd.n2262 585
R4907 gnd.n2262 gnd.n2258 585
R4908 gnd.n3953 gnd.n3952 585
R4909 gnd.n3952 gnd.n3951 585
R4910 gnd.n2264 gnd.n2263 585
R4911 gnd.n2305 gnd.n2264 585
R4912 gnd.n3923 gnd.n3922 585
R4913 gnd.n3924 gnd.n3923 585
R4914 gnd.n3921 gnd.n2276 585
R4915 gnd.n2276 gnd.n2273 585
R4916 gnd.n3920 gnd.n3919 585
R4917 gnd.n3919 gnd.n3918 585
R4918 gnd.n2278 gnd.n2277 585
R4919 gnd.n3891 gnd.n2278 585
R4920 gnd.n3904 gnd.n3903 585
R4921 gnd.n3905 gnd.n3904 585
R4922 gnd.n3902 gnd.n2289 585
R4923 gnd.n3897 gnd.n2289 585
R4924 gnd.n3901 gnd.n3900 585
R4925 gnd.n3900 gnd.n3899 585
R4926 gnd.n2291 gnd.n2290 585
R4927 gnd.n2318 gnd.n2291 585
R4928 gnd.n3867 gnd.n2328 585
R4929 gnd.n2328 gnd.n2317 585
R4930 gnd.n3869 gnd.n3868 585
R4931 gnd.n3870 gnd.n3869 585
R4932 gnd.n3866 gnd.n2327 585
R4933 gnd.n2327 gnd.n2324 585
R4934 gnd.n3865 gnd.n3864 585
R4935 gnd.n3864 gnd.n3863 585
R4936 gnd.n2330 gnd.n2329 585
R4937 gnd.n3810 gnd.n2330 585
R4938 gnd.n3851 gnd.n3850 585
R4939 gnd.n3852 gnd.n3851 585
R4940 gnd.n3849 gnd.n2342 585
R4941 gnd.n2342 gnd.n2339 585
R4942 gnd.n3848 gnd.n3847 585
R4943 gnd.n3847 gnd.n3846 585
R4944 gnd.n2344 gnd.n2343 585
R4945 gnd.n3818 gnd.n2344 585
R4946 gnd.n3833 gnd.n3832 585
R4947 gnd.n3834 gnd.n3833 585
R4948 gnd.n3831 gnd.n2355 585
R4949 gnd.n3824 gnd.n2355 585
R4950 gnd.n3830 gnd.n3829 585
R4951 gnd.n3829 gnd.n3828 585
R4952 gnd.n2357 gnd.n2356 585
R4953 gnd.n3796 gnd.n2357 585
R4954 gnd.n3782 gnd.n3781 585
R4955 gnd.n3781 gnd.n2363 585
R4956 gnd.n3783 gnd.n2372 585
R4957 gnd.n3715 gnd.n2372 585
R4958 gnd.n3785 gnd.n3784 585
R4959 gnd.n3786 gnd.n3785 585
R4960 gnd.n3780 gnd.n2371 585
R4961 gnd.n3775 gnd.n2371 585
R4962 gnd.n3779 gnd.n3778 585
R4963 gnd.n3778 gnd.n3777 585
R4964 gnd.n2374 gnd.n2373 585
R4965 gnd.n2386 gnd.n2374 585
R4966 gnd.n3739 gnd.n3738 585
R4967 gnd.n3738 gnd.n2385 585
R4968 gnd.n3740 gnd.n2396 585
R4969 gnd.n3726 gnd.n2396 585
R4970 gnd.n3742 gnd.n3741 585
R4971 gnd.n3743 gnd.n3742 585
R4972 gnd.n3737 gnd.n2395 585
R4973 gnd.n3732 gnd.n2395 585
R4974 gnd.n3736 gnd.n3735 585
R4975 gnd.n3735 gnd.n3734 585
R4976 gnd.n2398 gnd.n2397 585
R4977 gnd.n3709 gnd.n2398 585
R4978 gnd.n3695 gnd.n2413 585
R4979 gnd.n3673 gnd.n2413 585
R4980 gnd.n3697 gnd.n3696 585
R4981 gnd.n3698 gnd.n3697 585
R4982 gnd.n3694 gnd.n2412 585
R4983 gnd.n3688 gnd.n2412 585
R4984 gnd.n3693 gnd.n3692 585
R4985 gnd.n3692 gnd.n3691 585
R4986 gnd.n2415 gnd.n2414 585
R4987 gnd.n3681 gnd.n2415 585
R4988 gnd.n3657 gnd.n2432 585
R4989 gnd.n2432 gnd.n2431 585
R4990 gnd.n3659 gnd.n3658 585
R4991 gnd.n3660 gnd.n3659 585
R4992 gnd.n3656 gnd.n2429 585
R4993 gnd.n2429 gnd.n2426 585
R4994 gnd.n3655 gnd.n3654 585
R4995 gnd.n3654 gnd.n3653 585
R4996 gnd.n2434 gnd.n2433 585
R4997 gnd.n3569 gnd.n2434 585
R4998 gnd.n3637 gnd.n3636 585
R4999 gnd.n3638 gnd.n3637 585
R5000 gnd.n3635 gnd.n2447 585
R5001 gnd.n3630 gnd.n2447 585
R5002 gnd.n3634 gnd.n3633 585
R5003 gnd.n3633 gnd.n3632 585
R5004 gnd.n2449 gnd.n2448 585
R5005 gnd.n3618 gnd.n2449 585
R5006 gnd.n3605 gnd.n2470 585
R5007 gnd.n2470 gnd.n2459 585
R5008 gnd.n3607 gnd.n3606 585
R5009 gnd.n3608 gnd.n3607 585
R5010 gnd.n3604 gnd.n2469 585
R5011 gnd.n2469 gnd.t168 585
R5012 gnd.n3603 gnd.n3602 585
R5013 gnd.n3602 gnd.n3601 585
R5014 gnd.n2472 gnd.n2471 585
R5015 gnd.n3584 gnd.n2472 585
R5016 gnd.n3590 gnd.n3589 585
R5017 gnd.n3591 gnd.n3590 585
R5018 gnd.n3588 gnd.n3587 585
R5019 gnd.n3587 gnd.n2480 585
R5020 gnd.n1522 gnd.n1521 585
R5021 gnd.n3560 gnd.n1522 585
R5022 gnd.n4728 gnd.n4727 585
R5023 gnd.n4727 gnd.n4726 585
R5024 gnd.n4729 gnd.n1500 585
R5025 gnd.n3549 gnd.n1500 585
R5026 gnd.n4794 gnd.n4793 585
R5027 gnd.n4792 gnd.n1499 585
R5028 gnd.n4791 gnd.n1498 585
R5029 gnd.n4796 gnd.n1498 585
R5030 gnd.n4790 gnd.n4789 585
R5031 gnd.n4788 gnd.n4787 585
R5032 gnd.n4786 gnd.n4785 585
R5033 gnd.n4784 gnd.n4783 585
R5034 gnd.n4782 gnd.n4781 585
R5035 gnd.n4780 gnd.n4779 585
R5036 gnd.n4778 gnd.n4777 585
R5037 gnd.n4776 gnd.n4775 585
R5038 gnd.n4774 gnd.n4773 585
R5039 gnd.n4772 gnd.n4771 585
R5040 gnd.n4770 gnd.n4769 585
R5041 gnd.n4768 gnd.n4767 585
R5042 gnd.n4766 gnd.n4765 585
R5043 gnd.n4764 gnd.n4763 585
R5044 gnd.n4762 gnd.n4761 585
R5045 gnd.n4760 gnd.n4759 585
R5046 gnd.n4758 gnd.n4757 585
R5047 gnd.n4756 gnd.n4755 585
R5048 gnd.n4754 gnd.n4753 585
R5049 gnd.n4752 gnd.n4751 585
R5050 gnd.n4750 gnd.n4749 585
R5051 gnd.n4748 gnd.n4747 585
R5052 gnd.n4746 gnd.n4745 585
R5053 gnd.n4744 gnd.n4743 585
R5054 gnd.n4742 gnd.n4741 585
R5055 gnd.n4740 gnd.n4739 585
R5056 gnd.n4738 gnd.n4737 585
R5057 gnd.n4736 gnd.n4735 585
R5058 gnd.n4734 gnd.n1463 585
R5059 gnd.n4799 gnd.n4798 585
R5060 gnd.n1465 gnd.n1462 585
R5061 gnd.n3485 gnd.n3484 585
R5062 gnd.n3487 gnd.n3486 585
R5063 gnd.n3490 gnd.n3489 585
R5064 gnd.n3492 gnd.n3491 585
R5065 gnd.n3494 gnd.n3493 585
R5066 gnd.n3496 gnd.n3495 585
R5067 gnd.n3498 gnd.n3497 585
R5068 gnd.n3500 gnd.n3499 585
R5069 gnd.n3502 gnd.n3501 585
R5070 gnd.n3504 gnd.n3503 585
R5071 gnd.n3506 gnd.n3505 585
R5072 gnd.n3508 gnd.n3507 585
R5073 gnd.n3510 gnd.n3509 585
R5074 gnd.n3512 gnd.n3511 585
R5075 gnd.n3514 gnd.n3513 585
R5076 gnd.n3516 gnd.n3515 585
R5077 gnd.n3518 gnd.n3517 585
R5078 gnd.n3520 gnd.n3519 585
R5079 gnd.n3522 gnd.n3521 585
R5080 gnd.n3524 gnd.n3523 585
R5081 gnd.n3526 gnd.n3525 585
R5082 gnd.n3528 gnd.n3527 585
R5083 gnd.n3530 gnd.n3529 585
R5084 gnd.n3532 gnd.n3531 585
R5085 gnd.n3534 gnd.n3533 585
R5086 gnd.n3536 gnd.n3535 585
R5087 gnd.n3538 gnd.n3537 585
R5088 gnd.n3540 gnd.n3539 585
R5089 gnd.n3542 gnd.n3541 585
R5090 gnd.n3544 gnd.n3543 585
R5091 gnd.n3545 gnd.n3481 585
R5092 gnd.n4097 gnd.n4096 585
R5093 gnd.n4099 gnd.n4098 585
R5094 gnd.n4101 gnd.n4100 585
R5095 gnd.n4103 gnd.n4102 585
R5096 gnd.n4105 gnd.n4104 585
R5097 gnd.n4107 gnd.n4106 585
R5098 gnd.n4109 gnd.n4108 585
R5099 gnd.n4111 gnd.n4110 585
R5100 gnd.n4113 gnd.n4112 585
R5101 gnd.n4115 gnd.n4114 585
R5102 gnd.n4117 gnd.n4116 585
R5103 gnd.n4119 gnd.n4118 585
R5104 gnd.n4121 gnd.n4120 585
R5105 gnd.n4123 gnd.n4122 585
R5106 gnd.n4125 gnd.n4124 585
R5107 gnd.n4127 gnd.n4126 585
R5108 gnd.n4129 gnd.n4128 585
R5109 gnd.n4131 gnd.n4130 585
R5110 gnd.n4133 gnd.n4132 585
R5111 gnd.n4135 gnd.n4134 585
R5112 gnd.n4137 gnd.n4136 585
R5113 gnd.n4139 gnd.n4138 585
R5114 gnd.n4141 gnd.n4140 585
R5115 gnd.n4143 gnd.n4142 585
R5116 gnd.n4145 gnd.n4144 585
R5117 gnd.n4147 gnd.n4146 585
R5118 gnd.n4149 gnd.n4148 585
R5119 gnd.n4151 gnd.n4150 585
R5120 gnd.n4153 gnd.n4152 585
R5121 gnd.n4156 gnd.n4155 585
R5122 gnd.n4158 gnd.n4157 585
R5123 gnd.n4160 gnd.n4159 585
R5124 gnd.n4162 gnd.n4161 585
R5125 gnd.n4023 gnd.n2219 585
R5126 gnd.n4025 gnd.n4024 585
R5127 gnd.n4027 gnd.n4026 585
R5128 gnd.n4029 gnd.n4028 585
R5129 gnd.n4032 gnd.n4031 585
R5130 gnd.n4034 gnd.n4033 585
R5131 gnd.n4036 gnd.n4035 585
R5132 gnd.n4038 gnd.n4037 585
R5133 gnd.n4040 gnd.n4039 585
R5134 gnd.n4042 gnd.n4041 585
R5135 gnd.n4044 gnd.n4043 585
R5136 gnd.n4046 gnd.n4045 585
R5137 gnd.n4048 gnd.n4047 585
R5138 gnd.n4050 gnd.n4049 585
R5139 gnd.n4052 gnd.n4051 585
R5140 gnd.n4054 gnd.n4053 585
R5141 gnd.n4056 gnd.n4055 585
R5142 gnd.n4058 gnd.n4057 585
R5143 gnd.n4060 gnd.n4059 585
R5144 gnd.n4062 gnd.n4061 585
R5145 gnd.n4064 gnd.n4063 585
R5146 gnd.n4066 gnd.n4065 585
R5147 gnd.n4068 gnd.n4067 585
R5148 gnd.n4070 gnd.n4069 585
R5149 gnd.n4072 gnd.n4071 585
R5150 gnd.n4074 gnd.n4073 585
R5151 gnd.n4076 gnd.n4075 585
R5152 gnd.n4078 gnd.n4077 585
R5153 gnd.n4080 gnd.n4079 585
R5154 gnd.n4082 gnd.n4081 585
R5155 gnd.n4084 gnd.n4083 585
R5156 gnd.n4086 gnd.n4085 585
R5157 gnd.n4088 gnd.n4087 585
R5158 gnd.n4095 gnd.n2222 585
R5159 gnd.n4095 gnd.n2043 585
R5160 gnd.n4094 gnd.n2224 585
R5161 gnd.n4094 gnd.n4093 585
R5162 gnd.n3978 gnd.n2223 585
R5163 gnd.n3995 gnd.n2223 585
R5164 gnd.n3979 gnd.n2231 585
R5165 gnd.n3998 gnd.n2231 585
R5166 gnd.n3981 gnd.n3980 585
R5167 gnd.n3982 gnd.n3981 585
R5168 gnd.n3977 gnd.n2241 585
R5169 gnd.n2241 gnd.n2239 585
R5170 gnd.n3976 gnd.n3975 585
R5171 gnd.n3975 gnd.n3974 585
R5172 gnd.n2243 gnd.n2242 585
R5173 gnd.n3933 gnd.n2243 585
R5174 gnd.n2296 gnd.n2252 585
R5175 gnd.n3967 gnd.n2252 585
R5176 gnd.n2299 gnd.n2298 585
R5177 gnd.n2298 gnd.n2297 585
R5178 gnd.n2300 gnd.n2259 585
R5179 gnd.n3957 gnd.n2259 585
R5180 gnd.n2302 gnd.n2301 585
R5181 gnd.n2301 gnd.n2258 585
R5182 gnd.n2303 gnd.n2266 585
R5183 gnd.n3951 gnd.n2266 585
R5184 gnd.n2307 gnd.n2306 585
R5185 gnd.n2306 gnd.n2305 585
R5186 gnd.n2308 gnd.n2274 585
R5187 gnd.n3924 gnd.n2274 585
R5188 gnd.n2310 gnd.n2309 585
R5189 gnd.n2309 gnd.n2273 585
R5190 gnd.n2311 gnd.n2280 585
R5191 gnd.n3918 gnd.n2280 585
R5192 gnd.n3893 gnd.n3892 585
R5193 gnd.n3892 gnd.n3891 585
R5194 gnd.n3894 gnd.n2288 585
R5195 gnd.n3905 gnd.n2288 585
R5196 gnd.n3896 gnd.n3895 585
R5197 gnd.n3897 gnd.n3896 585
R5198 gnd.n2295 gnd.n2294 585
R5199 gnd.n3899 gnd.n2294 585
R5200 gnd.n3801 gnd.n3800 585
R5201 gnd.n3801 gnd.n2318 585
R5202 gnd.n3803 gnd.n3802 585
R5203 gnd.n3802 gnd.n2317 585
R5204 gnd.n3804 gnd.n2325 585
R5205 gnd.n3870 gnd.n2325 585
R5206 gnd.n3806 gnd.n3805 585
R5207 gnd.n3805 gnd.n2324 585
R5208 gnd.n3807 gnd.n2332 585
R5209 gnd.n3863 gnd.n2332 585
R5210 gnd.n3812 gnd.n3811 585
R5211 gnd.n3811 gnd.n3810 585
R5212 gnd.n3813 gnd.n2340 585
R5213 gnd.n3852 gnd.n2340 585
R5214 gnd.n3815 gnd.n3814 585
R5215 gnd.n3814 gnd.n2339 585
R5216 gnd.n3816 gnd.n2346 585
R5217 gnd.n3846 gnd.n2346 585
R5218 gnd.n3820 gnd.n3819 585
R5219 gnd.n3819 gnd.n3818 585
R5220 gnd.n3821 gnd.n2353 585
R5221 gnd.n3834 gnd.n2353 585
R5222 gnd.n3823 gnd.n3822 585
R5223 gnd.n3824 gnd.n3823 585
R5224 gnd.n3799 gnd.n2359 585
R5225 gnd.n3828 gnd.n2359 585
R5226 gnd.n3798 gnd.n3797 585
R5227 gnd.n3797 gnd.n3796 585
R5228 gnd.n2362 gnd.n2361 585
R5229 gnd.n2363 gnd.n2362 585
R5230 gnd.n3717 gnd.n3716 585
R5231 gnd.n3716 gnd.n3715 585
R5232 gnd.n3718 gnd.n2369 585
R5233 gnd.n3786 gnd.n2369 585
R5234 gnd.n3719 gnd.n2377 585
R5235 gnd.n3775 gnd.n2377 585
R5236 gnd.n3720 gnd.n2376 585
R5237 gnd.n3777 gnd.n2376 585
R5238 gnd.n3722 gnd.n3721 585
R5239 gnd.n3722 gnd.n2386 585
R5240 gnd.n3723 gnd.n3713 585
R5241 gnd.n3723 gnd.n2385 585
R5242 gnd.n3728 gnd.n3727 585
R5243 gnd.n3727 gnd.n3726 585
R5244 gnd.n3729 gnd.n2394 585
R5245 gnd.n3743 gnd.n2394 585
R5246 gnd.n3731 gnd.n3730 585
R5247 gnd.n3732 gnd.n3731 585
R5248 gnd.n3712 gnd.n2399 585
R5249 gnd.n3734 gnd.n2399 585
R5250 gnd.n3711 gnd.n3710 585
R5251 gnd.n3710 gnd.n3709 585
R5252 gnd.n2401 gnd.n2400 585
R5253 gnd.n3673 gnd.n2401 585
R5254 gnd.n3685 gnd.n2411 585
R5255 gnd.n3698 gnd.n2411 585
R5256 gnd.n3687 gnd.n3686 585
R5257 gnd.n3688 gnd.n3687 585
R5258 gnd.n3684 gnd.n2416 585
R5259 gnd.n3691 gnd.n2416 585
R5260 gnd.n3683 gnd.n3682 585
R5261 gnd.n3682 gnd.n3681 585
R5262 gnd.n2418 gnd.n2417 585
R5263 gnd.n2431 gnd.n2418 585
R5264 gnd.n3565 gnd.n2427 585
R5265 gnd.n3660 gnd.n2427 585
R5266 gnd.n3567 gnd.n3566 585
R5267 gnd.n3566 gnd.n2426 585
R5268 gnd.n3568 gnd.n2437 585
R5269 gnd.n3653 gnd.n2437 585
R5270 gnd.n3571 gnd.n3570 585
R5271 gnd.n3570 gnd.n3569 585
R5272 gnd.n3572 gnd.n2445 585
R5273 gnd.n3638 gnd.n2445 585
R5274 gnd.n3573 gnd.n2452 585
R5275 gnd.n3630 gnd.n2452 585
R5276 gnd.n3574 gnd.n2451 585
R5277 gnd.n3632 gnd.n2451 585
R5278 gnd.n3575 gnd.n2460 585
R5279 gnd.n3618 gnd.n2460 585
R5280 gnd.n3577 gnd.n3576 585
R5281 gnd.n3576 gnd.n2459 585
R5282 gnd.n3578 gnd.n2466 585
R5283 gnd.n3608 gnd.n2466 585
R5284 gnd.n3580 gnd.n3579 585
R5285 gnd.n3579 gnd.t168 585
R5286 gnd.n3581 gnd.n2474 585
R5287 gnd.n3601 gnd.n2474 585
R5288 gnd.n3583 gnd.n3582 585
R5289 gnd.n3584 gnd.n3583 585
R5290 gnd.n3564 gnd.n2481 585
R5291 gnd.n3591 gnd.n2481 585
R5292 gnd.n3563 gnd.n3562 585
R5293 gnd.n3562 gnd.n2480 585
R5294 gnd.n3561 gnd.n2483 585
R5295 gnd.n3561 gnd.n3560 585
R5296 gnd.n3546 gnd.n1524 585
R5297 gnd.n4726 gnd.n1524 585
R5298 gnd.n3548 gnd.n3547 585
R5299 gnd.n3549 gnd.n3548 585
R5300 gnd.n2756 gnd.n2755 585
R5301 gnd.n2755 gnd.n1179 585
R5302 gnd.n7367 gnd.n395 585
R5303 gnd.n395 gnd.n274 585
R5304 gnd.n7371 gnd.n7370 585
R5305 gnd.n7372 gnd.n7371 585
R5306 gnd.n345 gnd.n344 585
R5307 gnd.n345 gnd.n281 585
R5308 gnd.n7382 gnd.n7381 585
R5309 gnd.n7381 gnd.n7380 585
R5310 gnd.n7383 gnd.n339 585
R5311 gnd.n339 gnd.n290 585
R5312 gnd.n7385 gnd.n7384 585
R5313 gnd.n7385 gnd.n287 585
R5314 gnd.n7386 gnd.n338 585
R5315 gnd.n7386 gnd.n298 585
R5316 gnd.n7388 gnd.n7387 585
R5317 gnd.n7387 gnd.n296 585
R5318 gnd.n7389 gnd.n335 585
R5319 gnd.n335 gnd.n328 585
R5320 gnd.n7392 gnd.n7391 585
R5321 gnd.n7393 gnd.n7392 585
R5322 gnd.n336 gnd.n334 585
R5323 gnd.n334 gnd.n332 585
R5324 gnd.n4538 gnd.n1706 585
R5325 gnd.n4521 gnd.n1706 585
R5326 gnd.n4540 gnd.n4539 585
R5327 gnd.n4541 gnd.n4540 585
R5328 gnd.n4535 gnd.n1705 585
R5329 gnd.n1705 gnd.n1699 585
R5330 gnd.n4534 gnd.n4533 585
R5331 gnd.n4533 gnd.n4532 585
R5332 gnd.n4461 gnd.n1708 585
R5333 gnd.n1708 gnd.n313 585
R5334 gnd.n4463 gnd.n4462 585
R5335 gnd.n4462 gnd.n310 585
R5336 gnd.n4465 gnd.n4458 585
R5337 gnd.n4458 gnd.n1686 585
R5338 gnd.n4467 gnd.n4466 585
R5339 gnd.n4467 gnd.n1683 585
R5340 gnd.n4470 gnd.n4457 585
R5341 gnd.n4470 gnd.n4469 585
R5342 gnd.n4472 gnd.n4471 585
R5343 gnd.n4471 gnd.n1718 585
R5344 gnd.n4473 gnd.n1729 585
R5345 gnd.n1729 gnd.n1716 585
R5346 gnd.n4475 gnd.n4474 585
R5347 gnd.n4476 gnd.n4475 585
R5348 gnd.n1730 gnd.n1728 585
R5349 gnd.n1728 gnd.n1725 585
R5350 gnd.n4451 gnd.n4450 585
R5351 gnd.n4450 gnd.n4449 585
R5352 gnd.n1733 gnd.n1732 585
R5353 gnd.n1745 gnd.n1733 585
R5354 gnd.n4419 gnd.n1756 585
R5355 gnd.n1756 gnd.n1743 585
R5356 gnd.n4421 gnd.n4420 585
R5357 gnd.n4422 gnd.n4421 585
R5358 gnd.n1757 gnd.n1755 585
R5359 gnd.n1755 gnd.n1752 585
R5360 gnd.n4414 gnd.n4413 585
R5361 gnd.n4413 gnd.n4412 585
R5362 gnd.n1760 gnd.n1759 585
R5363 gnd.n1771 gnd.n1760 585
R5364 gnd.n4386 gnd.n1782 585
R5365 gnd.n1782 gnd.n1769 585
R5366 gnd.n4388 gnd.n4387 585
R5367 gnd.n4389 gnd.n4388 585
R5368 gnd.n1783 gnd.n1781 585
R5369 gnd.n1781 gnd.n1778 585
R5370 gnd.n4381 gnd.n4380 585
R5371 gnd.n4380 gnd.n4379 585
R5372 gnd.n1786 gnd.n1785 585
R5373 gnd.n1797 gnd.n1786 585
R5374 gnd.n4355 gnd.n1809 585
R5375 gnd.n1809 gnd.n1795 585
R5376 gnd.n4357 gnd.n4356 585
R5377 gnd.n4358 gnd.n4357 585
R5378 gnd.n1810 gnd.n1808 585
R5379 gnd.n4346 gnd.n1808 585
R5380 gnd.n4350 gnd.n4349 585
R5381 gnd.n4349 gnd.n4348 585
R5382 gnd.n1820 gnd.n1812 585
R5383 gnd.n4336 gnd.n1820 585
R5384 gnd.n1819 gnd.n1818 585
R5385 gnd.n1819 gnd.n1649 585
R5386 gnd.n1814 gnd.n1813 585
R5387 gnd.n1813 gnd.n1646 585
R5388 gnd.n1631 gnd.n1630 585
R5389 gnd.n1636 gnd.n1631 585
R5390 gnd.n4612 gnd.n4611 585
R5391 gnd.n4611 gnd.n4610 585
R5392 gnd.n4613 gnd.n1625 585
R5393 gnd.n1632 gnd.n1625 585
R5394 gnd.n4615 gnd.n4614 585
R5395 gnd.n4616 gnd.n4615 585
R5396 gnd.n1622 gnd.n1621 585
R5397 gnd.n4617 gnd.n1622 585
R5398 gnd.n4620 gnd.n4619 585
R5399 gnd.n4619 gnd.n4618 585
R5400 gnd.n4621 gnd.n1616 585
R5401 gnd.n1616 gnd.n1614 585
R5402 gnd.n4623 gnd.n4622 585
R5403 gnd.n4624 gnd.n4623 585
R5404 gnd.n1617 gnd.n1615 585
R5405 gnd.n1615 gnd.n1612 585
R5406 gnd.n4249 gnd.n4248 585
R5407 gnd.n4250 gnd.n4249 585
R5408 gnd.n1998 gnd.n1997 585
R5409 gnd.n4238 gnd.n1997 585
R5410 gnd.n4243 gnd.n4242 585
R5411 gnd.n4242 gnd.n4241 585
R5412 gnd.n2001 gnd.n2000 585
R5413 gnd.n4227 gnd.n2001 585
R5414 gnd.n4225 gnd.n4224 585
R5415 gnd.n4226 gnd.n4225 585
R5416 gnd.n2010 gnd.n2009 585
R5417 gnd.n4215 gnd.n2009 585
R5418 gnd.n4220 gnd.n4219 585
R5419 gnd.n4219 gnd.n4218 585
R5420 gnd.n2013 gnd.n2012 585
R5421 gnd.n4206 gnd.n2013 585
R5422 gnd.n4204 gnd.n4203 585
R5423 gnd.n4205 gnd.n4204 585
R5424 gnd.n2022 gnd.n2021 585
R5425 gnd.n4194 gnd.n2021 585
R5426 gnd.n4199 gnd.n4198 585
R5427 gnd.n4198 gnd.n4197 585
R5428 gnd.n2025 gnd.n2024 585
R5429 gnd.n4185 gnd.n2025 585
R5430 gnd.n4183 gnd.n4182 585
R5431 gnd.n4184 gnd.n4183 585
R5432 gnd.n2034 gnd.n2033 585
R5433 gnd.n4173 gnd.n2033 585
R5434 gnd.n4178 gnd.n4177 585
R5435 gnd.n4177 gnd.n4176 585
R5436 gnd.n2037 gnd.n2036 585
R5437 gnd.n4164 gnd.n2037 585
R5438 gnd.n3991 gnd.n2234 585
R5439 gnd.n2234 gnd.t182 585
R5440 gnd.n3993 gnd.n3992 585
R5441 gnd.n3994 gnd.n3993 585
R5442 gnd.n2235 gnd.n2233 585
R5443 gnd.n2233 gnd.n2230 585
R5444 gnd.n3986 gnd.n3985 585
R5445 gnd.n3985 gnd.n3984 585
R5446 gnd.n2238 gnd.n2237 585
R5447 gnd.n2244 gnd.n2238 585
R5448 gnd.n3965 gnd.n3964 585
R5449 gnd.n3966 gnd.n3965 585
R5450 gnd.n2254 gnd.n2253 585
R5451 gnd.n2261 gnd.n2253 585
R5452 gnd.n3960 gnd.n3959 585
R5453 gnd.n3959 gnd.n3958 585
R5454 gnd.n2257 gnd.n2256 585
R5455 gnd.n2265 gnd.n2257 585
R5456 gnd.n3913 gnd.n2282 585
R5457 gnd.n2282 gnd.n2275 585
R5458 gnd.n3915 gnd.n3914 585
R5459 gnd.n3916 gnd.n3915 585
R5460 gnd.n2283 gnd.n2281 585
R5461 gnd.n2281 gnd.n2279 585
R5462 gnd.n3908 gnd.n3907 585
R5463 gnd.n3907 gnd.n3906 585
R5464 gnd.n2286 gnd.n2285 585
R5465 gnd.n3898 gnd.n2286 585
R5466 gnd.n3879 gnd.n3878 585
R5467 gnd.n3880 gnd.n3879 585
R5468 gnd.n2320 gnd.n2319 585
R5469 gnd.n2326 gnd.n2319 585
R5470 gnd.n3874 gnd.n3873 585
R5471 gnd.n3873 gnd.n3872 585
R5472 gnd.n2323 gnd.n2322 585
R5473 gnd.n2331 gnd.n2323 585
R5474 gnd.n3842 gnd.n2348 585
R5475 gnd.n2348 gnd.n2341 585
R5476 gnd.n3844 gnd.n3843 585
R5477 gnd.n3845 gnd.n3844 585
R5478 gnd.n2349 gnd.n2347 585
R5479 gnd.n3817 gnd.n2347 585
R5480 gnd.n3837 gnd.n3836 585
R5481 gnd.n3836 gnd.n3835 585
R5482 gnd.n2352 gnd.n2351 585
R5483 gnd.n3827 gnd.n2352 585
R5484 gnd.n3794 gnd.n3793 585
R5485 gnd.n3795 gnd.n3794 585
R5486 gnd.n2365 gnd.n2364 585
R5487 gnd.n3714 gnd.n2364 585
R5488 gnd.n3789 gnd.n3788 585
R5489 gnd.n3788 gnd.n3787 585
R5490 gnd.n2368 gnd.n2367 585
R5491 gnd.n3776 gnd.n2368 585
R5492 gnd.n3751 gnd.n3750 585
R5493 gnd.n3752 gnd.n3751 585
R5494 gnd.n2388 gnd.n2387 585
R5495 gnd.n3725 gnd.n2387 585
R5496 gnd.n3746 gnd.n3745 585
R5497 gnd.n3745 gnd.n3744 585
R5498 gnd.n2391 gnd.n2390 585
R5499 gnd.n3733 gnd.n2391 585
R5500 gnd.n3671 gnd.n3670 585
R5501 gnd.n3671 gnd.n2402 585
R5502 gnd.n3676 gnd.n3675 585
R5503 gnd.n3675 gnd.n3674 585
R5504 gnd.n3677 gnd.n2421 585
R5505 gnd.n2421 gnd.n2410 585
R5506 gnd.n3679 gnd.n3678 585
R5507 gnd.n3680 gnd.n3679 585
R5508 gnd.n2422 gnd.n2420 585
R5509 gnd.n2430 gnd.n2420 585
R5510 gnd.n3663 gnd.n3662 585
R5511 gnd.n3662 gnd.n3661 585
R5512 gnd.n2425 gnd.n2424 585
R5513 gnd.n3652 gnd.n2425 585
R5514 gnd.n3626 gnd.n2454 585
R5515 gnd.n2454 gnd.n2446 585
R5516 gnd.n3628 gnd.n3627 585
R5517 gnd.n3629 gnd.n3628 585
R5518 gnd.n2455 gnd.n2453 585
R5519 gnd.n2453 gnd.n2450 585
R5520 gnd.n3621 gnd.n3620 585
R5521 gnd.n3620 gnd.n3619 585
R5522 gnd.n2458 gnd.n2457 585
R5523 gnd.n3609 gnd.n2458 585
R5524 gnd.n3599 gnd.n3598 585
R5525 gnd.n3600 gnd.n3599 585
R5526 gnd.n2476 gnd.n2475 585
R5527 gnd.n3585 gnd.n2475 585
R5528 gnd.n3594 gnd.n3593 585
R5529 gnd.n3593 gnd.n3592 585
R5530 gnd.n2479 gnd.n2478 585
R5531 gnd.n2479 gnd.n1526 585
R5532 gnd.n3477 gnd.n2490 585
R5533 gnd.n2490 gnd.n1523 585
R5534 gnd.n3479 gnd.n3478 585
R5535 gnd.n3480 gnd.n3479 585
R5536 gnd.n2491 gnd.n2489 585
R5537 gnd.n2497 gnd.n2489 585
R5538 gnd.n3472 gnd.n3471 585
R5539 gnd.n3471 gnd.n3470 585
R5540 gnd.n2494 gnd.n2493 585
R5541 gnd.n3459 gnd.n2494 585
R5542 gnd.n3433 gnd.n3432 585
R5543 gnd.n3433 gnd.n2505 585
R5544 gnd.n3435 gnd.n3434 585
R5545 gnd.n3434 gnd.n2514 585
R5546 gnd.n3436 gnd.n2525 585
R5547 gnd.n2525 gnd.n2524 585
R5548 gnd.n3438 gnd.n3437 585
R5549 gnd.n3439 gnd.n3438 585
R5550 gnd.n2526 gnd.n2523 585
R5551 gnd.n2523 gnd.n2520 585
R5552 gnd.n3425 gnd.n3424 585
R5553 gnd.n3424 gnd.n3423 585
R5554 gnd.n2529 gnd.n2528 585
R5555 gnd.n2538 gnd.n2529 585
R5556 gnd.n3400 gnd.n2550 585
R5557 gnd.n2550 gnd.n2537 585
R5558 gnd.n3402 gnd.n3401 585
R5559 gnd.n3403 gnd.n3402 585
R5560 gnd.n2551 gnd.n2549 585
R5561 gnd.n2549 gnd.n2546 585
R5562 gnd.n3395 gnd.n3394 585
R5563 gnd.n3394 gnd.n3393 585
R5564 gnd.n2554 gnd.n2553 585
R5565 gnd.n2563 gnd.n2554 585
R5566 gnd.n3224 gnd.n3223 585
R5567 gnd.n3223 gnd.n2562 585
R5568 gnd.n3225 gnd.n2675 585
R5569 gnd.n2675 gnd.n2673 585
R5570 gnd.n3227 gnd.n3226 585
R5571 gnd.n3228 gnd.n3227 585
R5572 gnd.n2676 gnd.n2674 585
R5573 gnd.n2674 gnd.n2649 585
R5574 gnd.n3217 gnd.n3216 585
R5575 gnd.n3216 gnd.n3215 585
R5576 gnd.n3214 gnd.n2678 585
R5577 gnd.n3214 gnd.n1423 585
R5578 gnd.n3213 gnd.n3212 585
R5579 gnd.n3213 gnd.n1412 585
R5580 gnd.n2680 gnd.n2679 585
R5581 gnd.n2679 gnd.n1405 585
R5582 gnd.n3208 gnd.n3207 585
R5583 gnd.n3207 gnd.n1402 585
R5584 gnd.n3206 gnd.n2682 585
R5585 gnd.n3206 gnd.n1394 585
R5586 gnd.n3205 gnd.n3204 585
R5587 gnd.n3205 gnd.n1391 585
R5588 gnd.n2684 gnd.n2683 585
R5589 gnd.n2683 gnd.n1383 585
R5590 gnd.n3200 gnd.n3199 585
R5591 gnd.n3199 gnd.n1380 585
R5592 gnd.n3198 gnd.n2686 585
R5593 gnd.n3198 gnd.n3197 585
R5594 gnd.n2805 gnd.n2687 585
R5595 gnd.n2687 gnd.n1370 585
R5596 gnd.n2807 gnd.n2806 585
R5597 gnd.n2807 gnd.n1362 585
R5598 gnd.n2809 gnd.n2808 585
R5599 gnd.n2808 gnd.n1359 585
R5600 gnd.n2810 gnd.n2798 585
R5601 gnd.n2798 gnd.n1351 585
R5602 gnd.n2812 gnd.n2811 585
R5603 gnd.n2812 gnd.n1348 585
R5604 gnd.n2813 gnd.n2797 585
R5605 gnd.n2813 gnd.n2702 585
R5606 gnd.n2815 gnd.n2814 585
R5607 gnd.n2814 gnd.n1338 585
R5608 gnd.n2816 gnd.n2792 585
R5609 gnd.n2792 gnd.n2706 585
R5610 gnd.n2818 gnd.n2817 585
R5611 gnd.n2818 gnd.n1328 585
R5612 gnd.n2819 gnd.n2791 585
R5613 gnd.n2819 gnd.n1320 585
R5614 gnd.n2821 gnd.n2820 585
R5615 gnd.n2820 gnd.n1317 585
R5616 gnd.n2822 gnd.n2786 585
R5617 gnd.n2786 gnd.n1309 585
R5618 gnd.n2824 gnd.n2823 585
R5619 gnd.n2824 gnd.n1306 585
R5620 gnd.n2825 gnd.n2785 585
R5621 gnd.n2825 gnd.n2716 585
R5622 gnd.n2827 gnd.n2826 585
R5623 gnd.n2826 gnd.n1296 585
R5624 gnd.n2828 gnd.n2780 585
R5625 gnd.n2780 gnd.n2720 585
R5626 gnd.n2830 gnd.n2829 585
R5627 gnd.n2830 gnd.n1286 585
R5628 gnd.n2831 gnd.n2779 585
R5629 gnd.n2831 gnd.n1278 585
R5630 gnd.n2833 gnd.n2832 585
R5631 gnd.n2832 gnd.n1275 585
R5632 gnd.n2834 gnd.n2777 585
R5633 gnd.n2777 gnd.n1267 585
R5634 gnd.n2836 gnd.n2835 585
R5635 gnd.n2836 gnd.n1264 585
R5636 gnd.n2838 gnd.n2837 585
R5637 gnd.n2837 gnd.n1259 585
R5638 gnd.n2840 gnd.n2839 585
R5639 gnd.n2840 gnd.n1256 585
R5640 gnd.n2842 gnd.n2841 585
R5641 gnd.n2841 gnd.n2733 585
R5642 gnd.n2844 gnd.n2843 585
R5643 gnd.n2844 gnd.n1247 585
R5644 gnd.n2846 gnd.n2845 585
R5645 gnd.n2846 gnd.n1242 585
R5646 gnd.n2847 gnd.n2775 585
R5647 gnd.n2847 gnd.n1239 585
R5648 gnd.n2849 gnd.n2848 585
R5649 gnd.n2848 gnd.n1231 585
R5650 gnd.n2776 gnd.n2770 585
R5651 gnd.n2776 gnd.n1228 585
R5652 gnd.n2853 gnd.n2769 585
R5653 gnd.n2769 gnd.n1222 585
R5654 gnd.n2854 gnd.n2748 585
R5655 gnd.n2748 gnd.n1219 585
R5656 gnd.n2856 gnd.n2855 585
R5657 gnd.n2857 gnd.n2856 585
R5658 gnd.n2749 gnd.n2747 585
R5659 gnd.n2747 gnd.n1209 585
R5660 gnd.n2764 gnd.n2763 585
R5661 gnd.n2763 gnd.n1201 585
R5662 gnd.n2762 gnd.n2751 585
R5663 gnd.n2762 gnd.n1198 585
R5664 gnd.n2761 gnd.n2760 585
R5665 gnd.n2761 gnd.n1190 585
R5666 gnd.n2753 gnd.n2752 585
R5667 gnd.n2752 gnd.n1187 585
R5668 gnd.n4627 gnd.n4626 585
R5669 gnd.n4626 gnd.n4625 585
R5670 gnd.n4628 gnd.n1609 585
R5671 gnd.n4251 gnd.n1609 585
R5672 gnd.n4629 gnd.n1608 585
R5673 gnd.n4237 gnd.n1608 585
R5674 gnd.n4239 gnd.n1606 585
R5675 gnd.n4240 gnd.n4239 585
R5676 gnd.n4633 gnd.n1605 585
R5677 gnd.n2002 gnd.n1605 585
R5678 gnd.n4634 gnd.n1604 585
R5679 gnd.n4228 gnd.n1604 585
R5680 gnd.n4635 gnd.n1603 585
R5681 gnd.n2008 gnd.n1603 585
R5682 gnd.n4216 gnd.n1601 585
R5683 gnd.n4217 gnd.n4216 585
R5684 gnd.n4639 gnd.n1600 585
R5685 gnd.n2014 gnd.n1600 585
R5686 gnd.n4640 gnd.n1599 585
R5687 gnd.n4207 gnd.n1599 585
R5688 gnd.n4641 gnd.n1598 585
R5689 gnd.n2020 gnd.n1598 585
R5690 gnd.n4195 gnd.n1596 585
R5691 gnd.n4196 gnd.n4195 585
R5692 gnd.n4645 gnd.n1595 585
R5693 gnd.n2026 gnd.n1595 585
R5694 gnd.n4646 gnd.n1594 585
R5695 gnd.n4186 gnd.n1594 585
R5696 gnd.n4647 gnd.n1593 585
R5697 gnd.n2032 gnd.n1593 585
R5698 gnd.n4174 gnd.n1591 585
R5699 gnd.n4175 gnd.n4174 585
R5700 gnd.n4651 gnd.n1590 585
R5701 gnd.n4163 gnd.n1590 585
R5702 gnd.n4652 gnd.n1589 585
R5703 gnd.n4165 gnd.n1589 585
R5704 gnd.n4653 gnd.n1588 585
R5705 gnd.n2225 gnd.n1588 585
R5706 gnd.n3996 gnd.n1586 585
R5707 gnd.n3997 gnd.n3996 585
R5708 gnd.n4657 gnd.n1585 585
R5709 gnd.n3983 gnd.n1585 585
R5710 gnd.n4658 gnd.n1584 585
R5711 gnd.n2245 gnd.n1584 585
R5712 gnd.n4659 gnd.n1583 585
R5713 gnd.n3934 gnd.n1583 585
R5714 gnd.n2250 gnd.n1581 585
R5715 gnd.n2251 gnd.n2250 585
R5716 gnd.n4663 gnd.n1580 585
R5717 gnd.n3957 gnd.n1580 585
R5718 gnd.n4664 gnd.n1579 585
R5719 gnd.n3950 gnd.n1579 585
R5720 gnd.n4665 gnd.n1578 585
R5721 gnd.n2304 gnd.n1578 585
R5722 gnd.n3925 gnd.n1576 585
R5723 gnd.n3926 gnd.n3925 585
R5724 gnd.n4669 gnd.n1575 585
R5725 gnd.n3917 gnd.n1575 585
R5726 gnd.n4670 gnd.n1574 585
R5727 gnd.n3890 gnd.n1574 585
R5728 gnd.n4671 gnd.n1573 585
R5729 gnd.n2287 gnd.n1573 585
R5730 gnd.n2292 gnd.n1571 585
R5731 gnd.n2293 gnd.n2292 585
R5732 gnd.n4675 gnd.n1570 585
R5733 gnd.n3881 gnd.n1570 585
R5734 gnd.n4676 gnd.n1569 585
R5735 gnd.n3871 gnd.n1569 585
R5736 gnd.n4677 gnd.n1568 585
R5737 gnd.n3862 gnd.n1568 585
R5738 gnd.n3808 gnd.n1566 585
R5739 gnd.n3809 gnd.n3808 585
R5740 gnd.n4681 gnd.n1565 585
R5741 gnd.n3853 gnd.n1565 585
R5742 gnd.n4682 gnd.n1564 585
R5743 gnd.n2345 gnd.n1564 585
R5744 gnd.n4683 gnd.n1563 585
R5745 gnd.n2354 gnd.n1563 585
R5746 gnd.n3825 gnd.n1561 585
R5747 gnd.n3826 gnd.n3825 585
R5748 gnd.n4687 gnd.n1560 585
R5749 gnd.n2358 gnd.n1560 585
R5750 gnd.n4688 gnd.n1559 585
R5751 gnd.n2363 gnd.n1559 585
R5752 gnd.n4689 gnd.n1558 585
R5753 gnd.n2370 gnd.n1558 585
R5754 gnd.n3773 gnd.n1556 585
R5755 gnd.n3774 gnd.n3773 585
R5756 gnd.n4693 gnd.n1555 585
R5757 gnd.n2375 gnd.n1555 585
R5758 gnd.n4694 gnd.n1554 585
R5759 gnd.n3753 gnd.n1554 585
R5760 gnd.n4695 gnd.n1553 585
R5761 gnd.n3724 gnd.n1553 585
R5762 gnd.n2392 gnd.n1551 585
R5763 gnd.n2393 gnd.n2392 585
R5764 gnd.n4699 gnd.n1550 585
R5765 gnd.n3708 gnd.n1550 585
R5766 gnd.n4700 gnd.n1549 585
R5767 gnd.n3672 gnd.n1549 585
R5768 gnd.n4701 gnd.n1548 585
R5769 gnd.n3699 gnd.n1548 585
R5770 gnd.n3689 gnd.n1546 585
R5771 gnd.n3690 gnd.n3689 585
R5772 gnd.n4705 gnd.n1545 585
R5773 gnd.n2419 gnd.n1545 585
R5774 gnd.n4706 gnd.n1544 585
R5775 gnd.n2428 gnd.n1544 585
R5776 gnd.n4707 gnd.n1543 585
R5777 gnd.n3651 gnd.n1543 585
R5778 gnd.n2435 gnd.n1541 585
R5779 gnd.n2436 gnd.n2435 585
R5780 gnd.n4711 gnd.n1540 585
R5781 gnd.n3639 gnd.n1540 585
R5782 gnd.n4712 gnd.n1539 585
R5783 gnd.n3631 gnd.n1539 585
R5784 gnd.n4713 gnd.n1538 585
R5785 gnd.n3618 gnd.n1538 585
R5786 gnd.n2467 gnd.n1536 585
R5787 gnd.n2468 gnd.n2467 585
R5788 gnd.n4717 gnd.n1535 585
R5789 gnd.n3610 gnd.n1535 585
R5790 gnd.n4718 gnd.n1534 585
R5791 gnd.n2473 gnd.n1534 585
R5792 gnd.n4719 gnd.n1533 585
R5793 gnd.n3586 gnd.n1533 585
R5794 gnd.n1530 gnd.n1528 585
R5795 gnd.n3559 gnd.n1528 585
R5796 gnd.n4724 gnd.n4723 585
R5797 gnd.n4725 gnd.n4724 585
R5798 gnd.n1529 gnd.n1527 585
R5799 gnd.n3550 gnd.n1527 585
R5800 gnd.n2501 gnd.n2499 585
R5801 gnd.n2499 gnd.n1497 585
R5802 gnd.n3468 gnd.n3467 585
R5803 gnd.n3469 gnd.n3468 585
R5804 gnd.n2500 gnd.n2498 585
R5805 gnd.n2498 gnd.n2495 585
R5806 gnd.n3462 gnd.n3461 585
R5807 gnd.n3461 gnd.n3460 585
R5808 gnd.n2504 gnd.n2503 585
R5809 gnd.n2513 gnd.n2504 585
R5810 gnd.n3447 gnd.n3446 585
R5811 gnd.n3448 gnd.n3447 585
R5812 gnd.n2516 gnd.n2515 585
R5813 gnd.n2522 gnd.n2515 585
R5814 gnd.n3442 gnd.n3441 585
R5815 gnd.n3441 gnd.n3440 585
R5816 gnd.n2519 gnd.n2518 585
R5817 gnd.n3422 gnd.n2519 585
R5818 gnd.n2542 gnd.n2540 585
R5819 gnd.n2540 gnd.n2530 585
R5820 gnd.n3412 gnd.n3411 585
R5821 gnd.n3413 gnd.n3412 585
R5822 gnd.n2541 gnd.n2539 585
R5823 gnd.n2548 gnd.n2539 585
R5824 gnd.n3406 gnd.n3405 585
R5825 gnd.n3405 gnd.n3404 585
R5826 gnd.n2545 gnd.n2544 585
R5827 gnd.n3392 gnd.n2545 585
R5828 gnd.n2567 gnd.n2565 585
R5829 gnd.n2565 gnd.n2555 585
R5830 gnd.n3382 gnd.n3381 585
R5831 gnd.n3383 gnd.n3382 585
R5832 gnd.n2566 gnd.n2564 585
R5833 gnd.n2672 gnd.n2564 585
R5834 gnd.n3229 gnd.n2576 585
R5835 gnd.n3370 gnd.n2577 585
R5836 gnd.n3369 gnd.n2578 585
R5837 gnd.n3231 gnd.n2578 585
R5838 gnd.n2650 gnd.n2579 585
R5839 gnd.n3362 gnd.n2585 585
R5840 gnd.n3361 gnd.n2586 585
R5841 gnd.n2652 gnd.n2587 585
R5842 gnd.n3354 gnd.n2595 585
R5843 gnd.n3353 gnd.n2596 585
R5844 gnd.n2655 gnd.n2597 585
R5845 gnd.n3346 gnd.n2603 585
R5846 gnd.n3345 gnd.n2604 585
R5847 gnd.n2657 gnd.n2605 585
R5848 gnd.n3338 gnd.n2613 585
R5849 gnd.n3337 gnd.n2614 585
R5850 gnd.n2660 gnd.n2615 585
R5851 gnd.n2664 gnd.n2663 585
R5852 gnd.n2665 gnd.n2633 585
R5853 gnd.n3250 gnd.n2634 585
R5854 gnd.n3249 gnd.n2635 585
R5855 gnd.n3248 gnd.n2636 585
R5856 gnd.n2668 gnd.n2637 585
R5857 gnd.n3244 gnd.n2639 585
R5858 gnd.n3243 gnd.n2640 585
R5859 gnd.n3242 gnd.n2641 585
R5860 gnd.n3239 gnd.n2646 585
R5861 gnd.n3238 gnd.n2647 585
R5862 gnd.n3237 gnd.n2648 585
R5863 gnd.n3234 gnd.n3233 585
R5864 gnd.n4254 gnd.n1613 585
R5865 gnd.n4625 gnd.n1613 585
R5866 gnd.n4253 gnd.n4252 585
R5867 gnd.n4252 gnd.n4251 585
R5868 gnd.n1996 gnd.n1995 585
R5869 gnd.n4237 gnd.n1996 585
R5870 gnd.n4236 gnd.n4235 585
R5871 gnd.n4240 gnd.n4236 585
R5872 gnd.n2004 gnd.n2003 585
R5873 gnd.n2003 gnd.n2002 585
R5874 gnd.n4230 gnd.n4229 585
R5875 gnd.n4229 gnd.n4228 585
R5876 gnd.n2007 gnd.n2006 585
R5877 gnd.n2008 gnd.n2007 585
R5878 gnd.n4214 gnd.n4213 585
R5879 gnd.n4217 gnd.n4214 585
R5880 gnd.n2016 gnd.n2015 585
R5881 gnd.n2015 gnd.n2014 585
R5882 gnd.n4209 gnd.n4208 585
R5883 gnd.n4208 gnd.n4207 585
R5884 gnd.n2019 gnd.n2018 585
R5885 gnd.n2020 gnd.n2019 585
R5886 gnd.n4193 gnd.n4192 585
R5887 gnd.n4196 gnd.n4193 585
R5888 gnd.n2028 gnd.n2027 585
R5889 gnd.n2027 gnd.n2026 585
R5890 gnd.n4188 gnd.n4187 585
R5891 gnd.n4187 gnd.n4186 585
R5892 gnd.n2031 gnd.n2030 585
R5893 gnd.n2032 gnd.n2031 585
R5894 gnd.n4172 gnd.n4171 585
R5895 gnd.n4175 gnd.n4172 585
R5896 gnd.n2039 gnd.n2038 585
R5897 gnd.n4163 gnd.n2038 585
R5898 gnd.n4167 gnd.n4166 585
R5899 gnd.n4166 gnd.n4165 585
R5900 gnd.n2042 gnd.n2041 585
R5901 gnd.n2225 gnd.n2042 585
R5902 gnd.n3938 gnd.n2232 585
R5903 gnd.n3997 gnd.n2232 585
R5904 gnd.n3937 gnd.n2240 585
R5905 gnd.n3983 gnd.n2240 585
R5906 gnd.n3942 gnd.n3936 585
R5907 gnd.n3936 gnd.n2245 585
R5908 gnd.n3943 gnd.n3935 585
R5909 gnd.n3935 gnd.n3934 585
R5910 gnd.n3944 gnd.n3932 585
R5911 gnd.n3932 gnd.n2251 585
R5912 gnd.n2269 gnd.n2260 585
R5913 gnd.n3957 gnd.n2260 585
R5914 gnd.n3949 gnd.n3948 585
R5915 gnd.n3950 gnd.n3949 585
R5916 gnd.n2268 gnd.n2267 585
R5917 gnd.n2304 gnd.n2267 585
R5918 gnd.n3928 gnd.n3927 585
R5919 gnd.n3927 gnd.n3926 585
R5920 gnd.n2272 gnd.n2271 585
R5921 gnd.n3917 gnd.n2272 585
R5922 gnd.n3889 gnd.n3888 585
R5923 gnd.n3890 gnd.n3889 585
R5924 gnd.n2313 gnd.n2312 585
R5925 gnd.n2312 gnd.n2287 585
R5926 gnd.n3884 gnd.n3883 585
R5927 gnd.n3883 gnd.n2293 585
R5928 gnd.n3882 gnd.n2315 585
R5929 gnd.n3882 gnd.n3881 585
R5930 gnd.n2335 gnd.n2316 585
R5931 gnd.n3871 gnd.n2316 585
R5932 gnd.n3861 gnd.n3860 585
R5933 gnd.n3862 gnd.n3861 585
R5934 gnd.n2334 gnd.n2333 585
R5935 gnd.n3809 gnd.n2333 585
R5936 gnd.n3855 gnd.n3854 585
R5937 gnd.n3854 gnd.n3853 585
R5938 gnd.n2338 gnd.n2337 585
R5939 gnd.n2345 gnd.n2338 585
R5940 gnd.n3762 gnd.n3761 585
R5941 gnd.n3761 gnd.n2354 585
R5942 gnd.n3765 gnd.n2360 585
R5943 gnd.n3826 gnd.n2360 585
R5944 gnd.n3766 gnd.n3760 585
R5945 gnd.n3760 gnd.n2358 585
R5946 gnd.n3767 gnd.n3759 585
R5947 gnd.n3759 gnd.n2363 585
R5948 gnd.n2381 gnd.n2379 585
R5949 gnd.n2379 gnd.n2370 585
R5950 gnd.n3772 gnd.n3771 585
R5951 gnd.n3774 gnd.n3772 585
R5952 gnd.n2380 gnd.n2378 585
R5953 gnd.n2378 gnd.n2375 585
R5954 gnd.n3755 gnd.n3754 585
R5955 gnd.n3754 gnd.n3753 585
R5956 gnd.n2384 gnd.n2383 585
R5957 gnd.n3724 gnd.n2384 585
R5958 gnd.n2406 gnd.n2404 585
R5959 gnd.n2404 gnd.n2393 585
R5960 gnd.n3707 gnd.n3706 585
R5961 gnd.n3708 gnd.n3707 585
R5962 gnd.n2405 gnd.n2403 585
R5963 gnd.n3672 gnd.n2403 585
R5964 gnd.n3701 gnd.n3700 585
R5965 gnd.n3700 gnd.n3699 585
R5966 gnd.n2409 gnd.n2408 585
R5967 gnd.n3690 gnd.n2409 585
R5968 gnd.n3645 gnd.n3644 585
R5969 gnd.n3644 gnd.n2419 585
R5970 gnd.n2441 gnd.n2439 585
R5971 gnd.n2439 gnd.n2428 585
R5972 gnd.n3650 gnd.n3649 585
R5973 gnd.n3651 gnd.n3650 585
R5974 gnd.n2440 gnd.n2438 585
R5975 gnd.n2438 gnd.n2436 585
R5976 gnd.n3641 gnd.n3640 585
R5977 gnd.n3640 gnd.n3639 585
R5978 gnd.n2444 gnd.n2443 585
R5979 gnd.n3631 gnd.n2444 585
R5980 gnd.n3617 gnd.n3616 585
R5981 gnd.n3618 gnd.n3617 585
R5982 gnd.n2462 gnd.n2461 585
R5983 gnd.n2468 gnd.n2461 585
R5984 gnd.n3612 gnd.n3611 585
R5985 gnd.n3611 gnd.n3610 585
R5986 gnd.n2465 gnd.n2464 585
R5987 gnd.n2473 gnd.n2465 585
R5988 gnd.n2485 gnd.n2482 585
R5989 gnd.n3586 gnd.n2482 585
R5990 gnd.n3558 gnd.n3557 585
R5991 gnd.n3559 gnd.n3558 585
R5992 gnd.n2484 gnd.n1525 585
R5993 gnd.n4725 gnd.n1525 585
R5994 gnd.n3552 gnd.n3551 585
R5995 gnd.n3551 gnd.n3550 585
R5996 gnd.n2488 gnd.n2487 585
R5997 gnd.n2488 gnd.n1497 585
R5998 gnd.n3453 gnd.n2496 585
R5999 gnd.n3469 gnd.n2496 585
R6000 gnd.n2509 gnd.n2507 585
R6001 gnd.n2507 gnd.n2495 585
R6002 gnd.n3458 gnd.n3457 585
R6003 gnd.n3460 gnd.n3458 585
R6004 gnd.n2508 gnd.n2506 585
R6005 gnd.n2513 gnd.n2506 585
R6006 gnd.n3450 gnd.n3449 585
R6007 gnd.n3449 gnd.n3448 585
R6008 gnd.n2512 gnd.n2511 585
R6009 gnd.n2522 gnd.n2512 585
R6010 gnd.n2533 gnd.n2521 585
R6011 gnd.n3440 gnd.n2521 585
R6012 gnd.n3421 gnd.n3420 585
R6013 gnd.n3422 gnd.n3421 585
R6014 gnd.n2532 gnd.n2531 585
R6015 gnd.n2531 gnd.n2530 585
R6016 gnd.n3415 gnd.n3414 585
R6017 gnd.n3414 gnd.n3413 585
R6018 gnd.n2536 gnd.n2535 585
R6019 gnd.n2548 gnd.n2536 585
R6020 gnd.n2558 gnd.n2547 585
R6021 gnd.n3404 gnd.n2547 585
R6022 gnd.n3391 gnd.n3390 585
R6023 gnd.n3392 gnd.n3391 585
R6024 gnd.n2557 gnd.n2556 585
R6025 gnd.n2556 gnd.n2555 585
R6026 gnd.n3385 gnd.n3384 585
R6027 gnd.n3384 gnd.n3383 585
R6028 gnd.n2561 gnd.n2560 585
R6029 gnd.n2672 gnd.n2561 585
R6030 gnd.n1993 gnd.n1992 585
R6031 gnd.n1992 gnd.n1623 585
R6032 gnd.n4258 gnd.n1991 585
R6033 gnd.n4259 gnd.n1989 585
R6034 gnd.n4260 gnd.n1988 585
R6035 gnd.n1986 gnd.n1981 585
R6036 gnd.n4264 gnd.n1980 585
R6037 gnd.n4265 gnd.n1978 585
R6038 gnd.n4266 gnd.n1977 585
R6039 gnd.n1975 gnd.n1973 585
R6040 gnd.n4270 gnd.n1972 585
R6041 gnd.n4271 gnd.n1970 585
R6042 gnd.n4272 gnd.n1969 585
R6043 gnd.n1967 gnd.n1844 585
R6044 gnd.n1966 gnd.n1965 585
R6045 gnd.n1950 gnd.n1846 585
R6046 gnd.n1952 gnd.n1951 585
R6047 gnd.n1948 gnd.n1853 585
R6048 gnd.n1947 gnd.n1946 585
R6049 gnd.n1931 gnd.n1855 585
R6050 gnd.n1933 gnd.n1932 585
R6051 gnd.n1929 gnd.n1862 585
R6052 gnd.n1928 gnd.n1927 585
R6053 gnd.n1912 gnd.n1864 585
R6054 gnd.n1914 gnd.n1913 585
R6055 gnd.n1910 gnd.n1871 585
R6056 gnd.n1909 gnd.n1908 585
R6057 gnd.n1893 gnd.n1873 585
R6058 gnd.n1895 gnd.n1894 585
R6059 gnd.n1891 gnd.n1611 585
R6060 gnd.n3482 gnd.t178 543.808
R6061 gnd.n2220 gnd.t90 543.808
R6062 gnd.n4731 gnd.t110 543.808
R6063 gnd.n4021 gnd.t147 543.808
R6064 gnd.n4087 gnd.n2227 478.086
R6065 gnd.n4096 gnd.n4095 478.086
R6066 gnd.n3548 gnd.n3481 478.086
R6067 gnd.n4794 gnd.n1500 478.086
R6068 gnd.n6702 gnd.n6701 400.269
R6069 gnd.n2642 gnd.t160 371.625
R6070 gnd.n118 gnd.t98 371.625
R6071 gnd.n1839 gnd.t128 371.625
R6072 gnd.n2618 gnd.t144 371.625
R6073 gnd.n2137 gnd.t121 371.625
R6074 gnd.n2166 gnd.t102 371.625
R6075 gnd.n197 gnd.t175 371.625
R6076 gnd.n7629 gnd.t187 371.625
R6077 gnd.n1062 gnd.t118 371.625
R6078 gnd.n1084 gnd.t94 371.625
R6079 gnd.n2934 gnd.t154 371.625
R6080 gnd.n3264 gnd.t114 371.625
R6081 gnd.n1458 gnd.t141 371.625
R6082 gnd.n1983 gnd.t131 371.625
R6083 gnd.n5713 gnd.t86 323.425
R6084 gnd.n5136 gnd.t124 323.425
R6085 gnd.n6390 gnd.n6364 289.615
R6086 gnd.n6358 gnd.n6332 289.615
R6087 gnd.n6326 gnd.n6300 289.615
R6088 gnd.n6295 gnd.n6269 289.615
R6089 gnd.n6263 gnd.n6237 289.615
R6090 gnd.n6231 gnd.n6205 289.615
R6091 gnd.n6199 gnd.n6173 289.615
R6092 gnd.n6168 gnd.n6142 289.615
R6093 gnd.n5563 gnd.t150 279.217
R6094 gnd.n5162 gnd.t106 279.217
R6095 gnd.n1507 gnd.t186 260.649
R6096 gnd.n4013 gnd.t166 260.649
R6097 gnd.n4796 gnd.n4795 256.663
R6098 gnd.n4796 gnd.n1466 256.663
R6099 gnd.n4796 gnd.n1467 256.663
R6100 gnd.n4796 gnd.n1468 256.663
R6101 gnd.n4796 gnd.n1469 256.663
R6102 gnd.n4796 gnd.n1470 256.663
R6103 gnd.n4796 gnd.n1471 256.663
R6104 gnd.n4796 gnd.n1472 256.663
R6105 gnd.n4796 gnd.n1473 256.663
R6106 gnd.n4796 gnd.n1474 256.663
R6107 gnd.n4796 gnd.n1475 256.663
R6108 gnd.n4796 gnd.n1476 256.663
R6109 gnd.n4796 gnd.n1477 256.663
R6110 gnd.n4796 gnd.n1478 256.663
R6111 gnd.n4796 gnd.n1479 256.663
R6112 gnd.n4796 gnd.n1480 256.663
R6113 gnd.n4799 gnd.n1464 256.663
R6114 gnd.n4797 gnd.n4796 256.663
R6115 gnd.n4796 gnd.n1481 256.663
R6116 gnd.n4796 gnd.n1482 256.663
R6117 gnd.n4796 gnd.n1483 256.663
R6118 gnd.n4796 gnd.n1484 256.663
R6119 gnd.n4796 gnd.n1485 256.663
R6120 gnd.n4796 gnd.n1486 256.663
R6121 gnd.n4796 gnd.n1487 256.663
R6122 gnd.n4796 gnd.n1488 256.663
R6123 gnd.n4796 gnd.n1489 256.663
R6124 gnd.n4796 gnd.n1490 256.663
R6125 gnd.n4796 gnd.n1491 256.663
R6126 gnd.n4796 gnd.n1492 256.663
R6127 gnd.n4796 gnd.n1493 256.663
R6128 gnd.n4796 gnd.n1494 256.663
R6129 gnd.n4796 gnd.n1495 256.663
R6130 gnd.n4796 gnd.n1496 256.663
R6131 gnd.n4162 gnd.n2061 256.663
R6132 gnd.n4162 gnd.n2062 256.663
R6133 gnd.n4162 gnd.n2063 256.663
R6134 gnd.n4162 gnd.n2064 256.663
R6135 gnd.n4162 gnd.n2065 256.663
R6136 gnd.n4162 gnd.n2066 256.663
R6137 gnd.n4162 gnd.n2067 256.663
R6138 gnd.n4162 gnd.n2068 256.663
R6139 gnd.n4162 gnd.n2069 256.663
R6140 gnd.n4162 gnd.n2070 256.663
R6141 gnd.n4162 gnd.n2071 256.663
R6142 gnd.n4162 gnd.n2072 256.663
R6143 gnd.n4162 gnd.n2073 256.663
R6144 gnd.n4162 gnd.n2074 256.663
R6145 gnd.n4162 gnd.n2075 256.663
R6146 gnd.n4162 gnd.n2076 256.663
R6147 gnd.n2219 gnd.n2077 256.663
R6148 gnd.n4162 gnd.n2060 256.663
R6149 gnd.n4162 gnd.n2059 256.663
R6150 gnd.n4162 gnd.n2058 256.663
R6151 gnd.n4162 gnd.n2057 256.663
R6152 gnd.n4162 gnd.n2056 256.663
R6153 gnd.n4162 gnd.n2055 256.663
R6154 gnd.n4162 gnd.n2054 256.663
R6155 gnd.n4162 gnd.n2053 256.663
R6156 gnd.n4162 gnd.n2052 256.663
R6157 gnd.n4162 gnd.n2051 256.663
R6158 gnd.n4162 gnd.n2050 256.663
R6159 gnd.n4162 gnd.n2049 256.663
R6160 gnd.n4162 gnd.n2048 256.663
R6161 gnd.n4162 gnd.n2047 256.663
R6162 gnd.n4162 gnd.n2046 256.663
R6163 gnd.n4162 gnd.n2045 256.663
R6164 gnd.n4162 gnd.n2044 256.663
R6165 gnd.n5107 gnd.n1030 242.672
R6166 gnd.n5107 gnd.n1031 242.672
R6167 gnd.n5107 gnd.n1032 242.672
R6168 gnd.n5107 gnd.n1033 242.672
R6169 gnd.n5107 gnd.n1034 242.672
R6170 gnd.n5107 gnd.n1035 242.672
R6171 gnd.n5107 gnd.n1036 242.672
R6172 gnd.n5107 gnd.n1037 242.672
R6173 gnd.n5107 gnd.n1038 242.672
R6174 gnd.n4829 gnd.n1422 242.672
R6175 gnd.n4829 gnd.n1421 242.672
R6176 gnd.n4829 gnd.n1420 242.672
R6177 gnd.n4829 gnd.n1419 242.672
R6178 gnd.n4829 gnd.n1418 242.672
R6179 gnd.n4829 gnd.n1417 242.672
R6180 gnd.n4829 gnd.n1416 242.672
R6181 gnd.n4829 gnd.n1415 242.672
R6182 gnd.n4829 gnd.n1414 242.672
R6183 gnd.n1880 gnd.n1624 242.672
R6184 gnd.n1900 gnd.n1624 242.672
R6185 gnd.n1902 gnd.n1624 242.672
R6186 gnd.n1919 gnd.n1624 242.672
R6187 gnd.n1921 gnd.n1624 242.672
R6188 gnd.n1938 gnd.n1624 242.672
R6189 gnd.n1940 gnd.n1624 242.672
R6190 gnd.n1957 gnd.n1624 242.672
R6191 gnd.n1959 gnd.n1624 242.672
R6192 gnd.n124 gnd.n121 242.672
R6193 gnd.n7540 gnd.n124 242.672
R6194 gnd.n7536 gnd.n124 242.672
R6195 gnd.n7533 gnd.n124 242.672
R6196 gnd.n7528 gnd.n124 242.672
R6197 gnd.n7525 gnd.n124 242.672
R6198 gnd.n7520 gnd.n124 242.672
R6199 gnd.n7517 gnd.n124 242.672
R6200 gnd.n7512 gnd.n124 242.672
R6201 gnd.n5618 gnd.n5527 242.672
R6202 gnd.n5531 gnd.n5527 242.672
R6203 gnd.n5611 gnd.n5527 242.672
R6204 gnd.n5605 gnd.n5527 242.672
R6205 gnd.n5603 gnd.n5527 242.672
R6206 gnd.n5597 gnd.n5527 242.672
R6207 gnd.n5595 gnd.n5527 242.672
R6208 gnd.n5589 gnd.n5527 242.672
R6209 gnd.n5587 gnd.n5527 242.672
R6210 gnd.n5581 gnd.n5527 242.672
R6211 gnd.n5579 gnd.n5527 242.672
R6212 gnd.n5572 gnd.n5527 242.672
R6213 gnd.n5570 gnd.n5527 242.672
R6214 gnd.n6511 gnd.n1011 242.672
R6215 gnd.n6511 gnd.n1010 242.672
R6216 gnd.n6511 gnd.n1009 242.672
R6217 gnd.n6511 gnd.n1008 242.672
R6218 gnd.n6511 gnd.n1007 242.672
R6219 gnd.n6511 gnd.n1006 242.672
R6220 gnd.n6511 gnd.n1005 242.672
R6221 gnd.n6511 gnd.n1004 242.672
R6222 gnd.n6511 gnd.n1003 242.672
R6223 gnd.n6511 gnd.n1002 242.672
R6224 gnd.n6511 gnd.n1001 242.672
R6225 gnd.n6511 gnd.n1000 242.672
R6226 gnd.n6511 gnd.n999 242.672
R6227 gnd.n5747 gnd.n5746 242.672
R6228 gnd.n5747 gnd.n5688 242.672
R6229 gnd.n5747 gnd.n5689 242.672
R6230 gnd.n5747 gnd.n5690 242.672
R6231 gnd.n5747 gnd.n5691 242.672
R6232 gnd.n5747 gnd.n5692 242.672
R6233 gnd.n5747 gnd.n5693 242.672
R6234 gnd.n5747 gnd.n5694 242.672
R6235 gnd.n6511 gnd.n5108 242.672
R6236 gnd.n6511 gnd.n5109 242.672
R6237 gnd.n6511 gnd.n5110 242.672
R6238 gnd.n6511 gnd.n5111 242.672
R6239 gnd.n6511 gnd.n5112 242.672
R6240 gnd.n6511 gnd.n5113 242.672
R6241 gnd.n6511 gnd.n5114 242.672
R6242 gnd.n6511 gnd.n6510 242.672
R6243 gnd.n5107 gnd.n5106 242.672
R6244 gnd.n5107 gnd.n1012 242.672
R6245 gnd.n5107 gnd.n1013 242.672
R6246 gnd.n5107 gnd.n1014 242.672
R6247 gnd.n5107 gnd.n1015 242.672
R6248 gnd.n5107 gnd.n1016 242.672
R6249 gnd.n5107 gnd.n1017 242.672
R6250 gnd.n5107 gnd.n1018 242.672
R6251 gnd.n5107 gnd.n1019 242.672
R6252 gnd.n5107 gnd.n1020 242.672
R6253 gnd.n5107 gnd.n1021 242.672
R6254 gnd.n5107 gnd.n1022 242.672
R6255 gnd.n5107 gnd.n1023 242.672
R6256 gnd.n5107 gnd.n1024 242.672
R6257 gnd.n5107 gnd.n1025 242.672
R6258 gnd.n5107 gnd.n1026 242.672
R6259 gnd.n5107 gnd.n1027 242.672
R6260 gnd.n5107 gnd.n1028 242.672
R6261 gnd.n5107 gnd.n1029 242.672
R6262 gnd.n4829 gnd.n1424 242.672
R6263 gnd.n4829 gnd.n1425 242.672
R6264 gnd.n4829 gnd.n1426 242.672
R6265 gnd.n4829 gnd.n1427 242.672
R6266 gnd.n4829 gnd.n1428 242.672
R6267 gnd.n4829 gnd.n1429 242.672
R6268 gnd.n4829 gnd.n1430 242.672
R6269 gnd.n4829 gnd.n1431 242.672
R6270 gnd.n4829 gnd.n1432 242.672
R6271 gnd.n4829 gnd.n1433 242.672
R6272 gnd.n4829 gnd.n1434 242.672
R6273 gnd.n4800 gnd.n1460 242.672
R6274 gnd.n4829 gnd.n1435 242.672
R6275 gnd.n4829 gnd.n1436 242.672
R6276 gnd.n4829 gnd.n1437 242.672
R6277 gnd.n4829 gnd.n1438 242.672
R6278 gnd.n4829 gnd.n1439 242.672
R6279 gnd.n4829 gnd.n1440 242.672
R6280 gnd.n4829 gnd.n1441 242.672
R6281 gnd.n4829 gnd.n4828 242.672
R6282 gnd.n2099 gnd.n1624 242.672
R6283 gnd.n2107 gnd.n1624 242.672
R6284 gnd.n2109 gnd.n1624 242.672
R6285 gnd.n2117 gnd.n1624 242.672
R6286 gnd.n2119 gnd.n1624 242.672
R6287 gnd.n2128 gnd.n1624 242.672
R6288 gnd.n2131 gnd.n1624 242.672
R6289 gnd.n2082 gnd.n1624 242.672
R6290 gnd.n2218 gnd.n2079 242.672
R6291 gnd.n2215 gnd.n1624 242.672
R6292 gnd.n2213 gnd.n1624 242.672
R6293 gnd.n2207 gnd.n1624 242.672
R6294 gnd.n2205 gnd.n1624 242.672
R6295 gnd.n2199 gnd.n1624 242.672
R6296 gnd.n2197 gnd.n1624 242.672
R6297 gnd.n2191 gnd.n1624 242.672
R6298 gnd.n2189 gnd.n1624 242.672
R6299 gnd.n2183 gnd.n1624 242.672
R6300 gnd.n2181 gnd.n1624 242.672
R6301 gnd.n2173 gnd.n1624 242.672
R6302 gnd.n194 gnd.n124 242.672
R6303 gnd.n7597 gnd.n124 242.672
R6304 gnd.n190 gnd.n124 242.672
R6305 gnd.n7604 gnd.n124 242.672
R6306 gnd.n183 gnd.n124 242.672
R6307 gnd.n7611 gnd.n124 242.672
R6308 gnd.n176 gnd.n124 242.672
R6309 gnd.n7618 gnd.n124 242.672
R6310 gnd.n169 gnd.n124 242.672
R6311 gnd.n7625 gnd.n124 242.672
R6312 gnd.n162 gnd.n124 242.672
R6313 gnd.n7635 gnd.n124 242.672
R6314 gnd.n155 gnd.n124 242.672
R6315 gnd.n7642 gnd.n124 242.672
R6316 gnd.n148 gnd.n124 242.672
R6317 gnd.n7649 gnd.n124 242.672
R6318 gnd.n141 gnd.n124 242.672
R6319 gnd.n7656 gnd.n124 242.672
R6320 gnd.n134 gnd.n124 242.672
R6321 gnd.n3231 gnd.n3230 242.672
R6322 gnd.n3231 gnd.n2651 242.672
R6323 gnd.n3231 gnd.n2653 242.672
R6324 gnd.n3231 gnd.n2654 242.672
R6325 gnd.n3231 gnd.n2656 242.672
R6326 gnd.n3231 gnd.n2658 242.672
R6327 gnd.n3231 gnd.n2659 242.672
R6328 gnd.n3231 gnd.n2661 242.672
R6329 gnd.n3231 gnd.n2666 242.672
R6330 gnd.n3231 gnd.n2667 242.672
R6331 gnd.n3231 gnd.n2669 242.672
R6332 gnd.n3231 gnd.n2670 242.672
R6333 gnd.n3231 gnd.n2671 242.672
R6334 gnd.n3232 gnd.n3231 242.672
R6335 gnd.n1990 gnd.n1623 242.672
R6336 gnd.n1987 gnd.n1623 242.672
R6337 gnd.n1979 gnd.n1623 242.672
R6338 gnd.n1976 gnd.n1623 242.672
R6339 gnd.n1971 gnd.n1623 242.672
R6340 gnd.n1968 gnd.n1623 242.672
R6341 gnd.n1845 gnd.n1623 242.672
R6342 gnd.n1949 gnd.n1623 242.672
R6343 gnd.n1854 gnd.n1623 242.672
R6344 gnd.n1930 gnd.n1623 242.672
R6345 gnd.n1863 gnd.n1623 242.672
R6346 gnd.n1911 gnd.n1623 242.672
R6347 gnd.n1872 gnd.n1623 242.672
R6348 gnd.n1892 gnd.n1623 242.672
R6349 gnd.n131 gnd.n127 240.244
R6350 gnd.n7658 gnd.n7657 240.244
R6351 gnd.n7655 gnd.n135 240.244
R6352 gnd.n7651 gnd.n7650 240.244
R6353 gnd.n7648 gnd.n142 240.244
R6354 gnd.n7644 gnd.n7643 240.244
R6355 gnd.n7641 gnd.n149 240.244
R6356 gnd.n7637 gnd.n7636 240.244
R6357 gnd.n7634 gnd.n156 240.244
R6358 gnd.n7627 gnd.n7626 240.244
R6359 gnd.n7624 gnd.n163 240.244
R6360 gnd.n7620 gnd.n7619 240.244
R6361 gnd.n7617 gnd.n170 240.244
R6362 gnd.n7613 gnd.n7612 240.244
R6363 gnd.n7610 gnd.n177 240.244
R6364 gnd.n7606 gnd.n7605 240.244
R6365 gnd.n7603 gnd.n184 240.244
R6366 gnd.n7599 gnd.n7598 240.244
R6367 gnd.n7596 gnd.n191 240.244
R6368 gnd.n2172 gnd.n1634 240.244
R6369 gnd.n4285 gnd.n1634 240.244
R6370 gnd.n4285 gnd.n1647 240.244
R6371 gnd.n4335 gnd.n1647 240.244
R6372 gnd.n4335 gnd.n1832 240.244
R6373 gnd.n1832 gnd.n1826 240.244
R6374 gnd.n1826 gnd.n1804 240.244
R6375 gnd.n4329 gnd.n1804 240.244
R6376 gnd.n4329 gnd.n1796 240.244
R6377 gnd.n4326 gnd.n1796 240.244
R6378 gnd.n4326 gnd.n1788 240.244
R6379 gnd.n1788 gnd.n1779 240.244
R6380 gnd.n4322 gnd.n1779 240.244
R6381 gnd.n4322 gnd.n1770 240.244
R6382 gnd.n4318 gnd.n1770 240.244
R6383 gnd.n4318 gnd.n1762 240.244
R6384 gnd.n1762 gnd.n1753 240.244
R6385 gnd.n4314 gnd.n1753 240.244
R6386 gnd.n4314 gnd.n1744 240.244
R6387 gnd.n4310 gnd.n1744 240.244
R6388 gnd.n4310 gnd.n1736 240.244
R6389 gnd.n1736 gnd.n1726 240.244
R6390 gnd.n1726 gnd.n1714 240.244
R6391 gnd.n4488 gnd.n1714 240.244
R6392 gnd.n4488 gnd.n1715 240.244
R6393 gnd.n1715 gnd.n1689 240.244
R6394 gnd.n1689 gnd.n1684 240.244
R6395 gnd.n4496 gnd.n1684 240.244
R6396 gnd.n4496 gnd.n311 240.244
R6397 gnd.n4530 gnd.n311 240.244
R6398 gnd.n4530 gnd.n1698 240.244
R6399 gnd.n1703 gnd.n1698 240.244
R6400 gnd.n4525 gnd.n1703 240.244
R6401 gnd.n4525 gnd.n4524 240.244
R6402 gnd.n4524 gnd.n333 240.244
R6403 gnd.n333 gnd.n326 240.244
R6404 gnd.n4516 gnd.n326 240.244
R6405 gnd.n4516 gnd.n297 240.244
R6406 gnd.n4512 gnd.n297 240.244
R6407 gnd.n4512 gnd.n288 240.244
R6408 gnd.n7378 gnd.n288 240.244
R6409 gnd.n7378 gnd.n280 240.244
R6410 gnd.n7374 gnd.n280 240.244
R6411 gnd.n7374 gnd.n272 240.244
R6412 gnd.n392 gnd.n272 240.244
R6413 gnd.n392 gnd.n266 240.244
R6414 gnd.n389 gnd.n266 240.244
R6415 gnd.n389 gnd.n257 240.244
R6416 gnd.n386 gnd.n257 240.244
R6417 gnd.n386 gnd.n249 240.244
R6418 gnd.n383 gnd.n249 240.244
R6419 gnd.n383 gnd.n242 240.244
R6420 gnd.n380 gnd.n242 240.244
R6421 gnd.n380 gnd.n236 240.244
R6422 gnd.n377 gnd.n236 240.244
R6423 gnd.n377 gnd.n227 240.244
R6424 gnd.n374 gnd.n227 240.244
R6425 gnd.n374 gnd.n220 240.244
R6426 gnd.n371 gnd.n220 240.244
R6427 gnd.n371 gnd.n210 240.244
R6428 gnd.n210 gnd.n201 240.244
R6429 gnd.n7587 gnd.n201 240.244
R6430 gnd.n7588 gnd.n7587 240.244
R6431 gnd.n7588 gnd.n123 240.244
R6432 gnd.n2100 gnd.n2093 240.244
R6433 gnd.n2106 gnd.n2093 240.244
R6434 gnd.n2110 gnd.n2108 240.244
R6435 gnd.n2116 gnd.n2089 240.244
R6436 gnd.n2120 gnd.n2118 240.244
R6437 gnd.n2127 gnd.n2085 240.244
R6438 gnd.n2130 gnd.n2129 240.244
R6439 gnd.n2132 gnd.n2083 240.244
R6440 gnd.n2216 gnd.n2214 240.244
R6441 gnd.n2212 gnd.n2141 240.244
R6442 gnd.n2208 gnd.n2206 240.244
R6443 gnd.n2204 gnd.n2147 240.244
R6444 gnd.n2200 gnd.n2198 240.244
R6445 gnd.n2196 gnd.n2153 240.244
R6446 gnd.n2192 gnd.n2190 240.244
R6447 gnd.n2188 gnd.n2159 240.244
R6448 gnd.n2184 gnd.n2182 240.244
R6449 gnd.n2180 gnd.n2165 240.244
R6450 gnd.n4608 gnd.n1638 240.244
R6451 gnd.n4608 gnd.n1639 240.244
R6452 gnd.n4604 gnd.n1639 240.244
R6453 gnd.n4604 gnd.n1645 240.244
R6454 gnd.n1824 gnd.n1645 240.244
R6455 gnd.n1824 gnd.n1803 240.244
R6456 gnd.n4360 gnd.n1803 240.244
R6457 gnd.n4360 gnd.n1798 240.244
R6458 gnd.n4368 gnd.n1798 240.244
R6459 gnd.n4368 gnd.n1799 240.244
R6460 gnd.n1799 gnd.n1777 240.244
R6461 gnd.n4392 gnd.n1777 240.244
R6462 gnd.n4392 gnd.n1772 240.244
R6463 gnd.n4400 gnd.n1772 240.244
R6464 gnd.n4400 gnd.n1773 240.244
R6465 gnd.n1773 gnd.n1751 240.244
R6466 gnd.n4424 gnd.n1751 240.244
R6467 gnd.n4424 gnd.n1746 240.244
R6468 gnd.n4432 gnd.n1746 240.244
R6469 gnd.n4432 gnd.n1747 240.244
R6470 gnd.n1747 gnd.n1724 240.244
R6471 gnd.n4478 gnd.n1724 240.244
R6472 gnd.n4478 gnd.n1720 240.244
R6473 gnd.n4486 gnd.n1720 240.244
R6474 gnd.n4486 gnd.n1687 240.244
R6475 gnd.n4560 gnd.n1687 240.244
R6476 gnd.n4561 gnd.n4560 240.244
R6477 gnd.n4561 gnd.n308 240.244
R6478 gnd.n7414 gnd.n308 240.244
R6479 gnd.n7414 gnd.n309 240.244
R6480 gnd.n4546 gnd.n309 240.244
R6481 gnd.n4546 gnd.n4543 240.244
R6482 gnd.n4543 gnd.n1700 240.244
R6483 gnd.n1700 gnd.n329 240.244
R6484 gnd.n7395 gnd.n329 240.244
R6485 gnd.n7397 gnd.n7395 240.244
R6486 gnd.n7397 gnd.n299 240.244
R6487 gnd.n7421 gnd.n299 240.244
R6488 gnd.n7421 gnd.n286 240.244
R6489 gnd.n7431 gnd.n286 240.244
R6490 gnd.n7431 gnd.n282 240.244
R6491 gnd.n7437 gnd.n282 240.244
R6492 gnd.n7437 gnd.n271 240.244
R6493 gnd.n7447 gnd.n271 240.244
R6494 gnd.n7447 gnd.n267 240.244
R6495 gnd.n7453 gnd.n267 240.244
R6496 gnd.n7453 gnd.n255 240.244
R6497 gnd.n7463 gnd.n255 240.244
R6498 gnd.n7463 gnd.n251 240.244
R6499 gnd.n7469 gnd.n251 240.244
R6500 gnd.n7469 gnd.n241 240.244
R6501 gnd.n7479 gnd.n241 240.244
R6502 gnd.n7479 gnd.n237 240.244
R6503 gnd.n7485 gnd.n237 240.244
R6504 gnd.n7485 gnd.n225 240.244
R6505 gnd.n7495 gnd.n225 240.244
R6506 gnd.n7495 gnd.n221 240.244
R6507 gnd.n7501 gnd.n221 240.244
R6508 gnd.n7501 gnd.n208 240.244
R6509 gnd.n7579 gnd.n208 240.244
R6510 gnd.n7579 gnd.n204 240.244
R6511 gnd.n7585 gnd.n204 240.244
R6512 gnd.n7585 gnd.n126 240.244
R6513 gnd.n7665 gnd.n126 240.244
R6514 gnd.n4830 gnd.n1411 240.244
R6515 gnd.n4827 gnd.n1442 240.244
R6516 gnd.n4823 gnd.n4822 240.244
R6517 gnd.n4819 gnd.n4818 240.244
R6518 gnd.n4815 gnd.n4814 240.244
R6519 gnd.n4811 gnd.n4810 240.244
R6520 gnd.n4807 gnd.n4806 240.244
R6521 gnd.n4803 gnd.n4802 240.244
R6522 gnd.n3276 gnd.n3275 240.244
R6523 gnd.n3283 gnd.n3282 240.244
R6524 gnd.n3286 gnd.n3285 240.244
R6525 gnd.n3293 gnd.n3292 240.244
R6526 gnd.n3296 gnd.n3295 240.244
R6527 gnd.n3303 gnd.n3302 240.244
R6528 gnd.n3306 gnd.n3305 240.244
R6529 gnd.n3313 gnd.n3312 240.244
R6530 gnd.n3316 gnd.n3315 240.244
R6531 gnd.n3321 gnd.n3266 240.244
R6532 gnd.n5028 gnd.n1088 240.244
R6533 gnd.n1092 gnd.n1088 240.244
R6534 gnd.n5021 gnd.n1092 240.244
R6535 gnd.n5021 gnd.n1093 240.244
R6536 gnd.n1106 gnd.n1093 240.244
R6537 gnd.n2875 gnd.n1106 240.244
R6538 gnd.n2875 gnd.n1117 240.244
R6539 gnd.n2878 gnd.n1117 240.244
R6540 gnd.n2878 gnd.n1127 240.244
R6541 gnd.n2883 gnd.n1127 240.244
R6542 gnd.n2883 gnd.n1137 240.244
R6543 gnd.n2886 gnd.n1137 240.244
R6544 gnd.n2886 gnd.n1147 240.244
R6545 gnd.n2891 gnd.n1147 240.244
R6546 gnd.n2891 gnd.n1157 240.244
R6547 gnd.n2894 gnd.n1157 240.244
R6548 gnd.n2894 gnd.n1167 240.244
R6549 gnd.n2899 gnd.n1167 240.244
R6550 gnd.n2899 gnd.n1177 240.244
R6551 gnd.n3034 gnd.n1177 240.244
R6552 gnd.n3034 gnd.n1188 240.244
R6553 gnd.n3040 gnd.n1188 240.244
R6554 gnd.n3040 gnd.n1199 240.244
R6555 gnd.n3050 gnd.n1199 240.244
R6556 gnd.n3050 gnd.n1210 240.244
R6557 gnd.n3056 gnd.n1210 240.244
R6558 gnd.n3056 gnd.n1220 240.244
R6559 gnd.n3066 gnd.n1220 240.244
R6560 gnd.n3066 gnd.n1229 240.244
R6561 gnd.n3072 gnd.n1229 240.244
R6562 gnd.n3072 gnd.n1240 240.244
R6563 gnd.n3082 gnd.n1240 240.244
R6564 gnd.n3082 gnd.n1248 240.244
R6565 gnd.n3088 gnd.n1248 240.244
R6566 gnd.n3088 gnd.n1257 240.244
R6567 gnd.n3098 gnd.n1257 240.244
R6568 gnd.n3098 gnd.n1265 240.244
R6569 gnd.n3104 gnd.n1265 240.244
R6570 gnd.n3104 gnd.n1276 240.244
R6571 gnd.n3114 gnd.n1276 240.244
R6572 gnd.n3114 gnd.n1287 240.244
R6573 gnd.n3120 gnd.n1287 240.244
R6574 gnd.n3120 gnd.n1297 240.244
R6575 gnd.n3130 gnd.n1297 240.244
R6576 gnd.n3130 gnd.n1307 240.244
R6577 gnd.n3136 gnd.n1307 240.244
R6578 gnd.n3136 gnd.n1318 240.244
R6579 gnd.n3146 gnd.n1318 240.244
R6580 gnd.n3146 gnd.n1329 240.244
R6581 gnd.n3152 gnd.n1329 240.244
R6582 gnd.n3152 gnd.n1339 240.244
R6583 gnd.n3162 gnd.n1339 240.244
R6584 gnd.n3162 gnd.n1349 240.244
R6585 gnd.n3169 gnd.n1349 240.244
R6586 gnd.n3169 gnd.n1360 240.244
R6587 gnd.n3179 gnd.n1360 240.244
R6588 gnd.n3179 gnd.n1371 240.244
R6589 gnd.n2688 gnd.n1371 240.244
R6590 gnd.n2688 gnd.n1381 240.244
R6591 gnd.n3187 gnd.n1381 240.244
R6592 gnd.n3187 gnd.n1392 240.244
R6593 gnd.n3259 gnd.n1392 240.244
R6594 gnd.n3259 gnd.n1403 240.244
R6595 gnd.n3328 gnd.n1403 240.244
R6596 gnd.n1042 gnd.n1041 240.244
R6597 gnd.n5100 gnd.n1041 240.244
R6598 gnd.n5098 gnd.n5097 240.244
R6599 gnd.n5094 gnd.n5093 240.244
R6600 gnd.n5090 gnd.n5089 240.244
R6601 gnd.n5086 gnd.n5085 240.244
R6602 gnd.n5082 gnd.n5081 240.244
R6603 gnd.n5078 gnd.n5077 240.244
R6604 gnd.n5074 gnd.n5073 240.244
R6605 gnd.n5069 gnd.n5068 240.244
R6606 gnd.n5065 gnd.n5064 240.244
R6607 gnd.n5061 gnd.n5060 240.244
R6608 gnd.n5057 gnd.n5056 240.244
R6609 gnd.n5053 gnd.n5052 240.244
R6610 gnd.n5049 gnd.n5048 240.244
R6611 gnd.n5045 gnd.n5044 240.244
R6612 gnd.n5041 gnd.n5040 240.244
R6613 gnd.n5037 gnd.n5036 240.244
R6614 gnd.n1083 gnd.n1082 240.244
R6615 gnd.n2991 gnd.n1043 240.244
R6616 gnd.n2991 gnd.n1098 240.244
R6617 gnd.n5019 gnd.n1098 240.244
R6618 gnd.n5019 gnd.n1099 240.244
R6619 gnd.n5015 gnd.n1099 240.244
R6620 gnd.n5015 gnd.n1105 240.244
R6621 gnd.n5007 gnd.n1105 240.244
R6622 gnd.n5007 gnd.n1120 240.244
R6623 gnd.n5003 gnd.n1120 240.244
R6624 gnd.n5003 gnd.n1126 240.244
R6625 gnd.n4995 gnd.n1126 240.244
R6626 gnd.n4995 gnd.n1140 240.244
R6627 gnd.n4991 gnd.n1140 240.244
R6628 gnd.n4991 gnd.n1146 240.244
R6629 gnd.n4983 gnd.n1146 240.244
R6630 gnd.n4983 gnd.n1160 240.244
R6631 gnd.n4979 gnd.n1160 240.244
R6632 gnd.n4979 gnd.n1166 240.244
R6633 gnd.n4971 gnd.n1166 240.244
R6634 gnd.n4971 gnd.n1180 240.244
R6635 gnd.n4967 gnd.n1180 240.244
R6636 gnd.n4967 gnd.n1186 240.244
R6637 gnd.n4959 gnd.n1186 240.244
R6638 gnd.n4959 gnd.n1202 240.244
R6639 gnd.n4955 gnd.n1202 240.244
R6640 gnd.n4955 gnd.n1208 240.244
R6641 gnd.n4947 gnd.n1208 240.244
R6642 gnd.n4947 gnd.n1223 240.244
R6643 gnd.n4942 gnd.n1223 240.244
R6644 gnd.n4942 gnd.n1227 240.244
R6645 gnd.n4934 gnd.n1227 240.244
R6646 gnd.n4934 gnd.n1243 240.244
R6647 gnd.n4929 gnd.n1243 240.244
R6648 gnd.n4929 gnd.n1246 240.244
R6649 gnd.n4921 gnd.n1246 240.244
R6650 gnd.n4921 gnd.n1260 240.244
R6651 gnd.n4916 gnd.n1260 240.244
R6652 gnd.n4916 gnd.n1263 240.244
R6653 gnd.n4908 gnd.n1263 240.244
R6654 gnd.n4908 gnd.n1279 240.244
R6655 gnd.n4904 gnd.n1279 240.244
R6656 gnd.n4904 gnd.n1285 240.244
R6657 gnd.n4896 gnd.n1285 240.244
R6658 gnd.n4896 gnd.n1299 240.244
R6659 gnd.n4892 gnd.n1299 240.244
R6660 gnd.n4892 gnd.n1305 240.244
R6661 gnd.n4884 gnd.n1305 240.244
R6662 gnd.n4884 gnd.n1321 240.244
R6663 gnd.n4880 gnd.n1321 240.244
R6664 gnd.n4880 gnd.n1327 240.244
R6665 gnd.n4872 gnd.n1327 240.244
R6666 gnd.n4872 gnd.n1341 240.244
R6667 gnd.n4868 gnd.n1341 240.244
R6668 gnd.n4868 gnd.n1347 240.244
R6669 gnd.n4860 gnd.n1347 240.244
R6670 gnd.n4860 gnd.n1363 240.244
R6671 gnd.n4856 gnd.n1363 240.244
R6672 gnd.n4856 gnd.n1369 240.244
R6673 gnd.n4848 gnd.n1369 240.244
R6674 gnd.n4848 gnd.n1384 240.244
R6675 gnd.n4844 gnd.n1384 240.244
R6676 gnd.n4844 gnd.n1390 240.244
R6677 gnd.n4836 gnd.n1390 240.244
R6678 gnd.n4836 gnd.n1406 240.244
R6679 gnd.n5115 gnd.n995 240.244
R6680 gnd.n6509 gnd.n5116 240.244
R6681 gnd.n6505 gnd.n6504 240.244
R6682 gnd.n6501 gnd.n6500 240.244
R6683 gnd.n6497 gnd.n6496 240.244
R6684 gnd.n6493 gnd.n6492 240.244
R6685 gnd.n6489 gnd.n6488 240.244
R6686 gnd.n6485 gnd.n6484 240.244
R6687 gnd.n5759 gnd.n5479 240.244
R6688 gnd.n5479 gnd.n5470 240.244
R6689 gnd.n5777 gnd.n5470 240.244
R6690 gnd.n5778 gnd.n5777 240.244
R6691 gnd.n5778 gnd.n5458 240.244
R6692 gnd.n5458 gnd.n5447 240.244
R6693 gnd.n5809 gnd.n5447 240.244
R6694 gnd.n5810 gnd.n5809 240.244
R6695 gnd.n5811 gnd.n5810 240.244
R6696 gnd.n5811 gnd.n5432 240.244
R6697 gnd.n5813 gnd.n5432 240.244
R6698 gnd.n5813 gnd.n5417 240.244
R6699 gnd.n5854 gnd.n5417 240.244
R6700 gnd.n5855 gnd.n5854 240.244
R6701 gnd.n5858 gnd.n5855 240.244
R6702 gnd.n5858 gnd.n5399 240.244
R6703 gnd.n5890 gnd.n5399 240.244
R6704 gnd.n5890 gnd.n5385 240.244
R6705 gnd.n5912 gnd.n5385 240.244
R6706 gnd.n5913 gnd.n5912 240.244
R6707 gnd.n5913 gnd.n5372 240.244
R6708 gnd.n5372 gnd.n5361 240.244
R6709 gnd.n5944 gnd.n5361 240.244
R6710 gnd.n5945 gnd.n5944 240.244
R6711 gnd.n5946 gnd.n5945 240.244
R6712 gnd.n5946 gnd.n5286 240.244
R6713 gnd.n5286 gnd.n5285 240.244
R6714 gnd.n5285 gnd.n5270 240.244
R6715 gnd.n5997 gnd.n5270 240.244
R6716 gnd.n5998 gnd.n5997 240.244
R6717 gnd.n5998 gnd.n5257 240.244
R6718 gnd.n5257 gnd.n5246 240.244
R6719 gnd.n6029 gnd.n5246 240.244
R6720 gnd.n6030 gnd.n6029 240.244
R6721 gnd.n6031 gnd.n6030 240.244
R6722 gnd.n6031 gnd.n5230 240.244
R6723 gnd.n5230 gnd.n5229 240.244
R6724 gnd.n5229 gnd.n5216 240.244
R6725 gnd.n6083 gnd.n5216 240.244
R6726 gnd.n6084 gnd.n6083 240.244
R6727 gnd.n6084 gnd.n5203 240.244
R6728 gnd.n5203 gnd.n5192 240.244
R6729 gnd.n6115 gnd.n5192 240.244
R6730 gnd.n6116 gnd.n6115 240.244
R6731 gnd.n6117 gnd.n6116 240.244
R6732 gnd.n6117 gnd.n964 240.244
R6733 gnd.n6134 gnd.n964 240.244
R6734 gnd.n6134 gnd.n974 240.244
R6735 gnd.n5173 gnd.n974 240.244
R6736 gnd.n6416 gnd.n5173 240.244
R6737 gnd.n6416 gnd.n986 240.244
R6738 gnd.n6412 gnd.n986 240.244
R6739 gnd.n6412 gnd.n997 240.244
R6740 gnd.n5696 gnd.n5695 240.244
R6741 gnd.n5740 gnd.n5695 240.244
R6742 gnd.n5738 gnd.n5737 240.244
R6743 gnd.n5734 gnd.n5733 240.244
R6744 gnd.n5730 gnd.n5729 240.244
R6745 gnd.n5726 gnd.n5725 240.244
R6746 gnd.n5722 gnd.n5721 240.244
R6747 gnd.n5718 gnd.n5717 240.244
R6748 gnd.n5769 gnd.n5477 240.244
R6749 gnd.n5769 gnd.n5473 240.244
R6750 gnd.n5775 gnd.n5473 240.244
R6751 gnd.n5775 gnd.n5456 240.244
R6752 gnd.n5799 gnd.n5456 240.244
R6753 gnd.n5799 gnd.n5451 240.244
R6754 gnd.n5807 gnd.n5451 240.244
R6755 gnd.n5807 gnd.n5452 240.244
R6756 gnd.n5452 gnd.n5430 240.244
R6757 gnd.n5833 gnd.n5430 240.244
R6758 gnd.n5833 gnd.n5425 240.244
R6759 gnd.n5844 gnd.n5425 240.244
R6760 gnd.n5844 gnd.n5426 240.244
R6761 gnd.n5840 gnd.n5426 240.244
R6762 gnd.n5840 gnd.n5397 240.244
R6763 gnd.n5894 gnd.n5397 240.244
R6764 gnd.n5894 gnd.n5392 240.244
R6765 gnd.n5902 gnd.n5392 240.244
R6766 gnd.n5902 gnd.n5393 240.244
R6767 gnd.n5393 gnd.n5370 240.244
R6768 gnd.n5934 gnd.n5370 240.244
R6769 gnd.n5934 gnd.n5365 240.244
R6770 gnd.n5942 gnd.n5365 240.244
R6771 gnd.n5942 gnd.n5366 240.244
R6772 gnd.n5366 gnd.n5283 240.244
R6773 gnd.n5979 gnd.n5283 240.244
R6774 gnd.n5979 gnd.n5278 240.244
R6775 gnd.n5987 gnd.n5278 240.244
R6776 gnd.n5987 gnd.n5279 240.244
R6777 gnd.n5279 gnd.n5255 240.244
R6778 gnd.n6019 gnd.n5255 240.244
R6779 gnd.n6019 gnd.n5250 240.244
R6780 gnd.n6027 gnd.n5250 240.244
R6781 gnd.n6027 gnd.n5251 240.244
R6782 gnd.n5251 gnd.n5228 240.244
R6783 gnd.n6065 gnd.n5228 240.244
R6784 gnd.n6065 gnd.n5223 240.244
R6785 gnd.n6073 gnd.n5223 240.244
R6786 gnd.n6073 gnd.n5224 240.244
R6787 gnd.n5224 gnd.n5201 240.244
R6788 gnd.n6104 gnd.n5201 240.244
R6789 gnd.n6104 gnd.n5196 240.244
R6790 gnd.n6113 gnd.n5196 240.244
R6791 gnd.n6113 gnd.n5197 240.244
R6792 gnd.n5197 gnd.n965 240.244
R6793 gnd.n6531 gnd.n965 240.244
R6794 gnd.n6531 gnd.n966 240.244
R6795 gnd.n6527 gnd.n966 240.244
R6796 gnd.n6527 gnd.n972 240.244
R6797 gnd.n987 gnd.n972 240.244
R6798 gnd.n6517 gnd.n987 240.244
R6799 gnd.n6517 gnd.n988 240.244
R6800 gnd.n6513 gnd.n988 240.244
R6801 gnd.n5140 gnd.n998 240.244
R6802 gnd.n6475 gnd.n6474 240.244
R6803 gnd.n6471 gnd.n6470 240.244
R6804 gnd.n6467 gnd.n6466 240.244
R6805 gnd.n6463 gnd.n6462 240.244
R6806 gnd.n6459 gnd.n6458 240.244
R6807 gnd.n6455 gnd.n6454 240.244
R6808 gnd.n6451 gnd.n6450 240.244
R6809 gnd.n6447 gnd.n6446 240.244
R6810 gnd.n6443 gnd.n6442 240.244
R6811 gnd.n6439 gnd.n6438 240.244
R6812 gnd.n6435 gnd.n6434 240.244
R6813 gnd.n6431 gnd.n6430 240.244
R6814 gnd.n5627 gnd.n5523 240.244
R6815 gnd.n5633 gnd.n5523 240.244
R6816 gnd.n5633 gnd.n5515 240.244
R6817 gnd.n5643 gnd.n5515 240.244
R6818 gnd.n5643 gnd.n5511 240.244
R6819 gnd.n5649 gnd.n5511 240.244
R6820 gnd.n5649 gnd.n5502 240.244
R6821 gnd.n5659 gnd.n5502 240.244
R6822 gnd.n5659 gnd.n5497 240.244
R6823 gnd.n5687 gnd.n5497 240.244
R6824 gnd.n5687 gnd.n5498 240.244
R6825 gnd.n5498 gnd.n5490 240.244
R6826 gnd.n5682 gnd.n5490 240.244
R6827 gnd.n5682 gnd.n5480 240.244
R6828 gnd.n5679 gnd.n5480 240.244
R6829 gnd.n5679 gnd.n5469 240.244
R6830 gnd.n5676 gnd.n5469 240.244
R6831 gnd.n5676 gnd.n5459 240.244
R6832 gnd.n5673 gnd.n5459 240.244
R6833 gnd.n5673 gnd.n5437 240.244
R6834 gnd.n5822 gnd.n5437 240.244
R6835 gnd.n5822 gnd.n5433 240.244
R6836 gnd.n5830 gnd.n5433 240.244
R6837 gnd.n5830 gnd.n5423 240.244
R6838 gnd.n5423 gnd.n5404 240.244
R6839 gnd.n5869 gnd.n5404 240.244
R6840 gnd.n5869 gnd.n5405 240.244
R6841 gnd.n5405 gnd.n5400 240.244
R6842 gnd.n5889 gnd.n5400 240.244
R6843 gnd.n5889 gnd.n5390 240.244
R6844 gnd.n5884 gnd.n5390 240.244
R6845 gnd.n5884 gnd.n5384 240.244
R6846 gnd.n5880 gnd.n5384 240.244
R6847 gnd.n5880 gnd.n5373 240.244
R6848 gnd.n5876 gnd.n5373 240.244
R6849 gnd.n5876 gnd.n5351 240.244
R6850 gnd.n5955 gnd.n5351 240.244
R6851 gnd.n5955 gnd.n5287 240.244
R6852 gnd.n5976 gnd.n5287 240.244
R6853 gnd.n5976 gnd.n5276 240.244
R6854 gnd.n5972 gnd.n5276 240.244
R6855 gnd.n5972 gnd.n5269 240.244
R6856 gnd.n5969 gnd.n5269 240.244
R6857 gnd.n5969 gnd.n5258 240.244
R6858 gnd.n5966 gnd.n5258 240.244
R6859 gnd.n5966 gnd.n5235 240.244
R6860 gnd.n6040 gnd.n5235 240.244
R6861 gnd.n6040 gnd.n5231 240.244
R6862 gnd.n6062 gnd.n5231 240.244
R6863 gnd.n6062 gnd.n5222 240.244
R6864 gnd.n6058 gnd.n5222 240.244
R6865 gnd.n6058 gnd.n5215 240.244
R6866 gnd.n6054 gnd.n5215 240.244
R6867 gnd.n6054 gnd.n5204 240.244
R6868 gnd.n6051 gnd.n5204 240.244
R6869 gnd.n6051 gnd.n5183 240.244
R6870 gnd.n6124 gnd.n5183 240.244
R6871 gnd.n6124 gnd.n5178 240.244
R6872 gnd.n6133 gnd.n5178 240.244
R6873 gnd.n6133 gnd.n5179 240.244
R6874 gnd.n5179 gnd.n975 240.244
R6875 gnd.n6419 gnd.n975 240.244
R6876 gnd.n6419 gnd.n985 240.244
R6877 gnd.n5169 gnd.n985 240.244
R6878 gnd.n6426 gnd.n5169 240.244
R6879 gnd.n5619 gnd.n5617 240.244
R6880 gnd.n5617 gnd.n5616 240.244
R6881 gnd.n5613 gnd.n5612 240.244
R6882 gnd.n5610 gnd.n5536 240.244
R6883 gnd.n5606 gnd.n5604 240.244
R6884 gnd.n5602 gnd.n5542 240.244
R6885 gnd.n5598 gnd.n5596 240.244
R6886 gnd.n5594 gnd.n5548 240.244
R6887 gnd.n5590 gnd.n5588 240.244
R6888 gnd.n5586 gnd.n5554 240.244
R6889 gnd.n5582 gnd.n5580 240.244
R6890 gnd.n5578 gnd.n5560 240.244
R6891 gnd.n5573 gnd.n5571 240.244
R6892 gnd.n5625 gnd.n5521 240.244
R6893 gnd.n5635 gnd.n5521 240.244
R6894 gnd.n5635 gnd.n5517 240.244
R6895 gnd.n5641 gnd.n5517 240.244
R6896 gnd.n5641 gnd.n5509 240.244
R6897 gnd.n5651 gnd.n5509 240.244
R6898 gnd.n5651 gnd.n5505 240.244
R6899 gnd.n5657 gnd.n5505 240.244
R6900 gnd.n5657 gnd.n5496 240.244
R6901 gnd.n5749 gnd.n5496 240.244
R6902 gnd.n5749 gnd.n5491 240.244
R6903 gnd.n5756 gnd.n5491 240.244
R6904 gnd.n5756 gnd.n5482 240.244
R6905 gnd.n5766 gnd.n5482 240.244
R6906 gnd.n5766 gnd.n5468 240.244
R6907 gnd.n5781 gnd.n5468 240.244
R6908 gnd.n5781 gnd.n5461 240.244
R6909 gnd.n5796 gnd.n5461 240.244
R6910 gnd.n5796 gnd.n5462 240.244
R6911 gnd.n5462 gnd.n5440 240.244
R6912 gnd.n5820 gnd.n5440 240.244
R6913 gnd.n5820 gnd.n5441 240.244
R6914 gnd.n5441 gnd.n5421 240.244
R6915 gnd.n5847 gnd.n5421 240.244
R6916 gnd.n5847 gnd.n5408 240.244
R6917 gnd.n5867 gnd.n5408 240.244
R6918 gnd.n5867 gnd.n5409 240.244
R6919 gnd.n5863 gnd.n5409 240.244
R6920 gnd.n5863 gnd.n5389 240.244
R6921 gnd.n5905 gnd.n5389 240.244
R6922 gnd.n5905 gnd.n5382 240.244
R6923 gnd.n5916 gnd.n5382 240.244
R6924 gnd.n5916 gnd.n5375 240.244
R6925 gnd.n5931 gnd.n5375 240.244
R6926 gnd.n5931 gnd.n5376 240.244
R6927 gnd.n5376 gnd.n5354 240.244
R6928 gnd.n5953 gnd.n5354 240.244
R6929 gnd.n5953 gnd.n5355 240.244
R6930 gnd.n5355 gnd.n5274 240.244
R6931 gnd.n5990 gnd.n5274 240.244
R6932 gnd.n5990 gnd.n5267 240.244
R6933 gnd.n6001 gnd.n5267 240.244
R6934 gnd.n6001 gnd.n5260 240.244
R6935 gnd.n6016 gnd.n5260 240.244
R6936 gnd.n6016 gnd.n5261 240.244
R6937 gnd.n5261 gnd.n5238 240.244
R6938 gnd.n6038 gnd.n5238 240.244
R6939 gnd.n6038 gnd.n5240 240.244
R6940 gnd.n5240 gnd.n5220 240.244
R6941 gnd.n6076 gnd.n5220 240.244
R6942 gnd.n6076 gnd.n5213 240.244
R6943 gnd.n6087 gnd.n5213 240.244
R6944 gnd.n6087 gnd.n5206 240.244
R6945 gnd.n6101 gnd.n5206 240.244
R6946 gnd.n6101 gnd.n5207 240.244
R6947 gnd.n5207 gnd.n5186 240.244
R6948 gnd.n6122 gnd.n5186 240.244
R6949 gnd.n6122 gnd.n5177 240.244
R6950 gnd.n6137 gnd.n5177 240.244
R6951 gnd.n6137 gnd.n977 240.244
R6952 gnd.n6524 gnd.n977 240.244
R6953 gnd.n6524 gnd.n978 240.244
R6954 gnd.n6520 gnd.n978 240.244
R6955 gnd.n6520 gnd.n984 240.244
R6956 gnd.n6405 gnd.n984 240.244
R6957 gnd.n7511 gnd.n7510 240.244
R6958 gnd.n7516 gnd.n7513 240.244
R6959 gnd.n7519 gnd.n7518 240.244
R6960 gnd.n7524 gnd.n7521 240.244
R6961 gnd.n7527 gnd.n7526 240.244
R6962 gnd.n7532 gnd.n7529 240.244
R6963 gnd.n7535 gnd.n7534 240.244
R6964 gnd.n7539 gnd.n7537 240.244
R6965 gnd.n7542 gnd.n7541 240.244
R6966 gnd.n4277 gnd.n1635 240.244
R6967 gnd.n4283 gnd.n1635 240.244
R6968 gnd.n4283 gnd.n1648 240.244
R6969 gnd.n4338 gnd.n1648 240.244
R6970 gnd.n4338 gnd.n1827 240.244
R6971 gnd.n4345 gnd.n1827 240.244
R6972 gnd.n4345 gnd.n1805 240.244
R6973 gnd.n1805 gnd.n1794 240.244
R6974 gnd.n4370 gnd.n1794 240.244
R6975 gnd.n4370 gnd.n1789 240.244
R6976 gnd.n4377 gnd.n1789 240.244
R6977 gnd.n4377 gnd.n1780 240.244
R6978 gnd.n1780 gnd.n1768 240.244
R6979 gnd.n4402 gnd.n1768 240.244
R6980 gnd.n4402 gnd.n1763 240.244
R6981 gnd.n4409 gnd.n1763 240.244
R6982 gnd.n4409 gnd.n1754 240.244
R6983 gnd.n1754 gnd.n1742 240.244
R6984 gnd.n4434 gnd.n1742 240.244
R6985 gnd.n4434 gnd.n1737 240.244
R6986 gnd.n4447 gnd.n1737 240.244
R6987 gnd.n4447 gnd.n1727 240.244
R6988 gnd.n4440 gnd.n1727 240.244
R6989 gnd.n4440 gnd.n1717 240.244
R6990 gnd.n1717 gnd.n1690 240.244
R6991 gnd.n4558 gnd.n1690 240.244
R6992 gnd.n4558 gnd.n1685 240.244
R6993 gnd.n1695 gnd.n1685 240.244
R6994 gnd.n1695 gnd.n312 240.244
R6995 gnd.n1696 gnd.n312 240.244
R6996 gnd.n4548 gnd.n1696 240.244
R6997 gnd.n4548 gnd.n1697 240.244
R6998 gnd.n1697 gnd.n78 240.244
R6999 gnd.n79 gnd.n78 240.244
R7000 gnd.n80 gnd.n79 240.244
R7001 gnd.n327 gnd.n80 240.244
R7002 gnd.n327 gnd.n83 240.244
R7003 gnd.n84 gnd.n83 240.244
R7004 gnd.n85 gnd.n84 240.244
R7005 gnd.n289 gnd.n85 240.244
R7006 gnd.n289 gnd.n88 240.244
R7007 gnd.n89 gnd.n88 240.244
R7008 gnd.n90 gnd.n89 240.244
R7009 gnd.n273 gnd.n90 240.244
R7010 gnd.n273 gnd.n93 240.244
R7011 gnd.n94 gnd.n93 240.244
R7012 gnd.n95 gnd.n94 240.244
R7013 gnd.n258 gnd.n95 240.244
R7014 gnd.n258 gnd.n98 240.244
R7015 gnd.n99 gnd.n98 240.244
R7016 gnd.n100 gnd.n99 240.244
R7017 gnd.n243 gnd.n100 240.244
R7018 gnd.n243 gnd.n103 240.244
R7019 gnd.n104 gnd.n103 240.244
R7020 gnd.n105 gnd.n104 240.244
R7021 gnd.n228 gnd.n105 240.244
R7022 gnd.n228 gnd.n108 240.244
R7023 gnd.n109 gnd.n108 240.244
R7024 gnd.n110 gnd.n109 240.244
R7025 gnd.n211 gnd.n110 240.244
R7026 gnd.n211 gnd.n113 240.244
R7027 gnd.n114 gnd.n113 240.244
R7028 gnd.n115 gnd.n114 240.244
R7029 gnd.n7667 gnd.n115 240.244
R7030 gnd.n1899 gnd.n1876 240.244
R7031 gnd.n1903 gnd.n1901 240.244
R7032 gnd.n1918 gnd.n1867 240.244
R7033 gnd.n1922 gnd.n1920 240.244
R7034 gnd.n1937 gnd.n1858 240.244
R7035 gnd.n1941 gnd.n1939 240.244
R7036 gnd.n1956 gnd.n1849 240.244
R7037 gnd.n1960 gnd.n1958 240.244
R7038 gnd.n4276 gnd.n1838 240.244
R7039 gnd.n1882 gnd.n1637 240.244
R7040 gnd.n1650 gnd.n1637 240.244
R7041 gnd.n4602 gnd.n1650 240.244
R7042 gnd.n4602 gnd.n1651 240.244
R7043 gnd.n1656 gnd.n1651 240.244
R7044 gnd.n1657 gnd.n1656 240.244
R7045 gnd.n1658 gnd.n1657 240.244
R7046 gnd.n1806 gnd.n1658 240.244
R7047 gnd.n1806 gnd.n1661 240.244
R7048 gnd.n1662 gnd.n1661 240.244
R7049 gnd.n1663 gnd.n1662 240.244
R7050 gnd.n4390 gnd.n1663 240.244
R7051 gnd.n4390 gnd.n1666 240.244
R7052 gnd.n1667 gnd.n1666 240.244
R7053 gnd.n1668 gnd.n1667 240.244
R7054 gnd.n4410 gnd.n1668 240.244
R7055 gnd.n4410 gnd.n1671 240.244
R7056 gnd.n1672 gnd.n1671 240.244
R7057 gnd.n1673 gnd.n1672 240.244
R7058 gnd.n1734 gnd.n1673 240.244
R7059 gnd.n1734 gnd.n1676 240.244
R7060 gnd.n1677 gnd.n1676 240.244
R7061 gnd.n1678 gnd.n1677 240.244
R7062 gnd.n1719 gnd.n1678 240.244
R7063 gnd.n1719 gnd.n1681 240.244
R7064 gnd.n1682 gnd.n1681 240.244
R7065 gnd.n4563 gnd.n1682 240.244
R7066 gnd.n4563 gnd.n314 240.244
R7067 gnd.n7412 gnd.n314 240.244
R7068 gnd.n7412 gnd.n315 240.244
R7069 gnd.n320 gnd.n315 240.244
R7070 gnd.n321 gnd.n320 240.244
R7071 gnd.n322 gnd.n321 240.244
R7072 gnd.n4522 gnd.n322 240.244
R7073 gnd.n4522 gnd.n325 240.244
R7074 gnd.n7399 gnd.n325 240.244
R7075 gnd.n7399 gnd.n295 240.244
R7076 gnd.n7423 gnd.n295 240.244
R7077 gnd.n7423 gnd.n291 240.244
R7078 gnd.n7429 gnd.n291 240.244
R7079 gnd.n7429 gnd.n279 240.244
R7080 gnd.n7439 gnd.n279 240.244
R7081 gnd.n7439 gnd.n275 240.244
R7082 gnd.n7445 gnd.n275 240.244
R7083 gnd.n7445 gnd.n264 240.244
R7084 gnd.n7455 gnd.n264 240.244
R7085 gnd.n7455 gnd.n260 240.244
R7086 gnd.n7461 gnd.n260 240.244
R7087 gnd.n7461 gnd.n248 240.244
R7088 gnd.n7471 gnd.n248 240.244
R7089 gnd.n7471 gnd.n244 240.244
R7090 gnd.n7477 gnd.n244 240.244
R7091 gnd.n7477 gnd.n234 240.244
R7092 gnd.n7487 gnd.n234 240.244
R7093 gnd.n7487 gnd.n230 240.244
R7094 gnd.n7493 gnd.n230 240.244
R7095 gnd.n7493 gnd.n219 240.244
R7096 gnd.n7503 gnd.n219 240.244
R7097 gnd.n7503 gnd.n213 240.244
R7098 gnd.n7577 gnd.n213 240.244
R7099 gnd.n7577 gnd.n214 240.244
R7100 gnd.n214 gnd.n203 240.244
R7101 gnd.n7508 gnd.n203 240.244
R7102 gnd.n7508 gnd.n125 240.244
R7103 gnd.n2570 gnd.n1413 240.244
R7104 gnd.n2572 gnd.n2571 240.244
R7105 gnd.n2582 gnd.n2581 240.244
R7106 gnd.n2590 gnd.n2589 240.244
R7107 gnd.n2592 gnd.n2591 240.244
R7108 gnd.n2600 gnd.n2599 240.244
R7109 gnd.n2608 gnd.n2607 240.244
R7110 gnd.n2610 gnd.n2609 240.244
R7111 gnd.n2621 gnd.n2617 240.244
R7112 gnd.n2993 gnd.n2913 240.244
R7113 gnd.n2994 gnd.n2993 240.244
R7114 gnd.n2994 gnd.n1095 240.244
R7115 gnd.n2999 gnd.n1095 240.244
R7116 gnd.n2999 gnd.n1107 240.244
R7117 gnd.n3002 gnd.n1107 240.244
R7118 gnd.n3002 gnd.n1118 240.244
R7119 gnd.n3007 gnd.n1118 240.244
R7120 gnd.n3007 gnd.n1128 240.244
R7121 gnd.n3010 gnd.n1128 240.244
R7122 gnd.n3010 gnd.n1138 240.244
R7123 gnd.n3015 gnd.n1138 240.244
R7124 gnd.n3015 gnd.n1148 240.244
R7125 gnd.n3018 gnd.n1148 240.244
R7126 gnd.n3018 gnd.n1158 240.244
R7127 gnd.n3023 gnd.n1158 240.244
R7128 gnd.n3023 gnd.n1168 240.244
R7129 gnd.n3026 gnd.n1168 240.244
R7130 gnd.n3026 gnd.n1178 240.244
R7131 gnd.n3032 gnd.n1178 240.244
R7132 gnd.n3032 gnd.n1189 240.244
R7133 gnd.n3042 gnd.n1189 240.244
R7134 gnd.n3042 gnd.n1200 240.244
R7135 gnd.n3048 gnd.n1200 240.244
R7136 gnd.n3048 gnd.n1211 240.244
R7137 gnd.n3058 gnd.n1211 240.244
R7138 gnd.n3058 gnd.n1221 240.244
R7139 gnd.n3064 gnd.n1221 240.244
R7140 gnd.n3064 gnd.n1230 240.244
R7141 gnd.n3074 gnd.n1230 240.244
R7142 gnd.n3074 gnd.n1241 240.244
R7143 gnd.n3080 gnd.n1241 240.244
R7144 gnd.n3080 gnd.n1249 240.244
R7145 gnd.n3090 gnd.n1249 240.244
R7146 gnd.n3090 gnd.n1258 240.244
R7147 gnd.n3096 gnd.n1258 240.244
R7148 gnd.n3096 gnd.n1266 240.244
R7149 gnd.n3106 gnd.n1266 240.244
R7150 gnd.n3106 gnd.n1277 240.244
R7151 gnd.n3112 gnd.n1277 240.244
R7152 gnd.n3112 gnd.n1288 240.244
R7153 gnd.n3122 gnd.n1288 240.244
R7154 gnd.n3122 gnd.n1298 240.244
R7155 gnd.n3128 gnd.n1298 240.244
R7156 gnd.n3128 gnd.n1308 240.244
R7157 gnd.n3138 gnd.n1308 240.244
R7158 gnd.n3138 gnd.n1319 240.244
R7159 gnd.n3144 gnd.n1319 240.244
R7160 gnd.n3144 gnd.n1330 240.244
R7161 gnd.n3154 gnd.n1330 240.244
R7162 gnd.n3154 gnd.n1340 240.244
R7163 gnd.n3160 gnd.n1340 240.244
R7164 gnd.n3160 gnd.n1350 240.244
R7165 gnd.n3171 gnd.n1350 240.244
R7166 gnd.n3171 gnd.n1361 240.244
R7167 gnd.n3177 gnd.n1361 240.244
R7168 gnd.n3177 gnd.n1372 240.244
R7169 gnd.n3195 gnd.n1372 240.244
R7170 gnd.n3195 gnd.n1382 240.244
R7171 gnd.n3189 gnd.n1382 240.244
R7172 gnd.n3189 gnd.n1393 240.244
R7173 gnd.n3257 gnd.n1393 240.244
R7174 gnd.n3257 gnd.n1404 240.244
R7175 gnd.n3330 gnd.n1404 240.244
R7176 gnd.n2973 gnd.n2972 240.244
R7177 gnd.n2969 gnd.n2968 240.244
R7178 gnd.n2965 gnd.n2964 240.244
R7179 gnd.n2961 gnd.n2960 240.244
R7180 gnd.n2957 gnd.n2956 240.244
R7181 gnd.n2953 gnd.n2952 240.244
R7182 gnd.n2949 gnd.n2948 240.244
R7183 gnd.n2945 gnd.n2944 240.244
R7184 gnd.n2933 gnd.n1039 240.244
R7185 gnd.n2985 gnd.n2914 240.244
R7186 gnd.n2985 gnd.n2915 240.244
R7187 gnd.n2915 gnd.n1097 240.244
R7188 gnd.n1109 gnd.n1097 240.244
R7189 gnd.n5013 gnd.n1109 240.244
R7190 gnd.n5013 gnd.n1110 240.244
R7191 gnd.n5009 gnd.n1110 240.244
R7192 gnd.n5009 gnd.n1116 240.244
R7193 gnd.n5001 gnd.n1116 240.244
R7194 gnd.n5001 gnd.n1129 240.244
R7195 gnd.n4997 gnd.n1129 240.244
R7196 gnd.n4997 gnd.n1135 240.244
R7197 gnd.n4989 gnd.n1135 240.244
R7198 gnd.n4989 gnd.n1150 240.244
R7199 gnd.n4985 gnd.n1150 240.244
R7200 gnd.n4985 gnd.n1156 240.244
R7201 gnd.n4977 gnd.n1156 240.244
R7202 gnd.n4977 gnd.n1169 240.244
R7203 gnd.n4973 gnd.n1169 240.244
R7204 gnd.n4973 gnd.n1175 240.244
R7205 gnd.n4965 gnd.n1175 240.244
R7206 gnd.n4965 gnd.n1191 240.244
R7207 gnd.n4961 gnd.n1191 240.244
R7208 gnd.n4961 gnd.n1197 240.244
R7209 gnd.n4953 gnd.n1197 240.244
R7210 gnd.n4953 gnd.n1212 240.244
R7211 gnd.n4949 gnd.n1212 240.244
R7212 gnd.n4949 gnd.n1218 240.244
R7213 gnd.n4940 gnd.n1218 240.244
R7214 gnd.n4940 gnd.n1232 240.244
R7215 gnd.n4936 gnd.n1232 240.244
R7216 gnd.n4936 gnd.n1238 240.244
R7217 gnd.n4927 gnd.n1238 240.244
R7218 gnd.n4927 gnd.n1250 240.244
R7219 gnd.n4923 gnd.n1250 240.244
R7220 gnd.n4923 gnd.n1255 240.244
R7221 gnd.n4914 gnd.n1255 240.244
R7222 gnd.n4914 gnd.n1268 240.244
R7223 gnd.n4910 gnd.n1268 240.244
R7224 gnd.n4910 gnd.n1274 240.244
R7225 gnd.n4902 gnd.n1274 240.244
R7226 gnd.n4902 gnd.n1289 240.244
R7227 gnd.n4898 gnd.n1289 240.244
R7228 gnd.n4898 gnd.n1295 240.244
R7229 gnd.n4890 gnd.n1295 240.244
R7230 gnd.n4890 gnd.n1310 240.244
R7231 gnd.n4886 gnd.n1310 240.244
R7232 gnd.n4886 gnd.n1316 240.244
R7233 gnd.n4878 gnd.n1316 240.244
R7234 gnd.n4878 gnd.n1331 240.244
R7235 gnd.n4874 gnd.n1331 240.244
R7236 gnd.n4874 gnd.n1337 240.244
R7237 gnd.n4866 gnd.n1337 240.244
R7238 gnd.n4866 gnd.n1352 240.244
R7239 gnd.n4862 gnd.n1352 240.244
R7240 gnd.n4862 gnd.n1358 240.244
R7241 gnd.n4854 gnd.n1358 240.244
R7242 gnd.n4854 gnd.n1373 240.244
R7243 gnd.n4850 gnd.n1373 240.244
R7244 gnd.n4850 gnd.n1379 240.244
R7245 gnd.n4842 gnd.n1379 240.244
R7246 gnd.n4842 gnd.n1395 240.244
R7247 gnd.n4838 gnd.n1395 240.244
R7248 gnd.n4838 gnd.n1401 240.244
R7249 gnd.n6704 gnd.n795 240.244
R7250 gnd.n6704 gnd.n791 240.244
R7251 gnd.n6710 gnd.n791 240.244
R7252 gnd.n6710 gnd.n789 240.244
R7253 gnd.n6714 gnd.n789 240.244
R7254 gnd.n6714 gnd.n785 240.244
R7255 gnd.n6720 gnd.n785 240.244
R7256 gnd.n6720 gnd.n783 240.244
R7257 gnd.n6724 gnd.n783 240.244
R7258 gnd.n6724 gnd.n779 240.244
R7259 gnd.n6730 gnd.n779 240.244
R7260 gnd.n6730 gnd.n777 240.244
R7261 gnd.n6734 gnd.n777 240.244
R7262 gnd.n6734 gnd.n773 240.244
R7263 gnd.n6740 gnd.n773 240.244
R7264 gnd.n6740 gnd.n771 240.244
R7265 gnd.n6744 gnd.n771 240.244
R7266 gnd.n6744 gnd.n767 240.244
R7267 gnd.n6750 gnd.n767 240.244
R7268 gnd.n6750 gnd.n765 240.244
R7269 gnd.n6754 gnd.n765 240.244
R7270 gnd.n6754 gnd.n761 240.244
R7271 gnd.n6760 gnd.n761 240.244
R7272 gnd.n6760 gnd.n759 240.244
R7273 gnd.n6764 gnd.n759 240.244
R7274 gnd.n6764 gnd.n755 240.244
R7275 gnd.n6770 gnd.n755 240.244
R7276 gnd.n6770 gnd.n753 240.244
R7277 gnd.n6774 gnd.n753 240.244
R7278 gnd.n6774 gnd.n749 240.244
R7279 gnd.n6780 gnd.n749 240.244
R7280 gnd.n6780 gnd.n747 240.244
R7281 gnd.n6784 gnd.n747 240.244
R7282 gnd.n6784 gnd.n743 240.244
R7283 gnd.n6790 gnd.n743 240.244
R7284 gnd.n6790 gnd.n741 240.244
R7285 gnd.n6794 gnd.n741 240.244
R7286 gnd.n6794 gnd.n737 240.244
R7287 gnd.n6800 gnd.n737 240.244
R7288 gnd.n6800 gnd.n735 240.244
R7289 gnd.n6804 gnd.n735 240.244
R7290 gnd.n6804 gnd.n731 240.244
R7291 gnd.n6810 gnd.n731 240.244
R7292 gnd.n6810 gnd.n729 240.244
R7293 gnd.n6814 gnd.n729 240.244
R7294 gnd.n6814 gnd.n725 240.244
R7295 gnd.n6820 gnd.n725 240.244
R7296 gnd.n6820 gnd.n723 240.244
R7297 gnd.n6824 gnd.n723 240.244
R7298 gnd.n6824 gnd.n719 240.244
R7299 gnd.n6830 gnd.n719 240.244
R7300 gnd.n6830 gnd.n717 240.244
R7301 gnd.n6834 gnd.n717 240.244
R7302 gnd.n6834 gnd.n713 240.244
R7303 gnd.n6840 gnd.n713 240.244
R7304 gnd.n6840 gnd.n711 240.244
R7305 gnd.n6844 gnd.n711 240.244
R7306 gnd.n6844 gnd.n707 240.244
R7307 gnd.n6850 gnd.n707 240.244
R7308 gnd.n6850 gnd.n705 240.244
R7309 gnd.n6854 gnd.n705 240.244
R7310 gnd.n6854 gnd.n701 240.244
R7311 gnd.n6860 gnd.n701 240.244
R7312 gnd.n6860 gnd.n699 240.244
R7313 gnd.n6864 gnd.n699 240.244
R7314 gnd.n6864 gnd.n695 240.244
R7315 gnd.n6870 gnd.n695 240.244
R7316 gnd.n6870 gnd.n693 240.244
R7317 gnd.n6874 gnd.n693 240.244
R7318 gnd.n6874 gnd.n689 240.244
R7319 gnd.n6880 gnd.n689 240.244
R7320 gnd.n6880 gnd.n687 240.244
R7321 gnd.n6884 gnd.n687 240.244
R7322 gnd.n6884 gnd.n683 240.244
R7323 gnd.n6890 gnd.n683 240.244
R7324 gnd.n6890 gnd.n681 240.244
R7325 gnd.n6894 gnd.n681 240.244
R7326 gnd.n6894 gnd.n677 240.244
R7327 gnd.n6900 gnd.n677 240.244
R7328 gnd.n6900 gnd.n675 240.244
R7329 gnd.n6904 gnd.n675 240.244
R7330 gnd.n6904 gnd.n671 240.244
R7331 gnd.n6910 gnd.n671 240.244
R7332 gnd.n6910 gnd.n669 240.244
R7333 gnd.n6914 gnd.n669 240.244
R7334 gnd.n6914 gnd.n665 240.244
R7335 gnd.n6920 gnd.n665 240.244
R7336 gnd.n6920 gnd.n663 240.244
R7337 gnd.n6924 gnd.n663 240.244
R7338 gnd.n6924 gnd.n659 240.244
R7339 gnd.n6930 gnd.n659 240.244
R7340 gnd.n6930 gnd.n657 240.244
R7341 gnd.n6934 gnd.n657 240.244
R7342 gnd.n6934 gnd.n653 240.244
R7343 gnd.n6940 gnd.n653 240.244
R7344 gnd.n6940 gnd.n651 240.244
R7345 gnd.n6944 gnd.n651 240.244
R7346 gnd.n6944 gnd.n647 240.244
R7347 gnd.n6950 gnd.n647 240.244
R7348 gnd.n6950 gnd.n645 240.244
R7349 gnd.n6954 gnd.n645 240.244
R7350 gnd.n6954 gnd.n641 240.244
R7351 gnd.n6960 gnd.n641 240.244
R7352 gnd.n6960 gnd.n639 240.244
R7353 gnd.n6964 gnd.n639 240.244
R7354 gnd.n6964 gnd.n635 240.244
R7355 gnd.n6970 gnd.n635 240.244
R7356 gnd.n6970 gnd.n633 240.244
R7357 gnd.n6974 gnd.n633 240.244
R7358 gnd.n6974 gnd.n629 240.244
R7359 gnd.n6980 gnd.n629 240.244
R7360 gnd.n6980 gnd.n627 240.244
R7361 gnd.n6984 gnd.n627 240.244
R7362 gnd.n6984 gnd.n623 240.244
R7363 gnd.n6990 gnd.n623 240.244
R7364 gnd.n6990 gnd.n621 240.244
R7365 gnd.n6994 gnd.n621 240.244
R7366 gnd.n6994 gnd.n617 240.244
R7367 gnd.n7000 gnd.n617 240.244
R7368 gnd.n7000 gnd.n615 240.244
R7369 gnd.n7004 gnd.n615 240.244
R7370 gnd.n7004 gnd.n611 240.244
R7371 gnd.n7010 gnd.n611 240.244
R7372 gnd.n7010 gnd.n609 240.244
R7373 gnd.n7014 gnd.n609 240.244
R7374 gnd.n7014 gnd.n605 240.244
R7375 gnd.n7020 gnd.n605 240.244
R7376 gnd.n7020 gnd.n603 240.244
R7377 gnd.n7024 gnd.n603 240.244
R7378 gnd.n7024 gnd.n599 240.244
R7379 gnd.n7030 gnd.n599 240.244
R7380 gnd.n7030 gnd.n597 240.244
R7381 gnd.n7034 gnd.n597 240.244
R7382 gnd.n7034 gnd.n593 240.244
R7383 gnd.n7040 gnd.n593 240.244
R7384 gnd.n7040 gnd.n591 240.244
R7385 gnd.n7044 gnd.n591 240.244
R7386 gnd.n7044 gnd.n587 240.244
R7387 gnd.n7050 gnd.n587 240.244
R7388 gnd.n7050 gnd.n585 240.244
R7389 gnd.n7054 gnd.n585 240.244
R7390 gnd.n7054 gnd.n581 240.244
R7391 gnd.n7060 gnd.n581 240.244
R7392 gnd.n7060 gnd.n579 240.244
R7393 gnd.n7064 gnd.n579 240.244
R7394 gnd.n7064 gnd.n575 240.244
R7395 gnd.n7070 gnd.n575 240.244
R7396 gnd.n7070 gnd.n573 240.244
R7397 gnd.n7074 gnd.n573 240.244
R7398 gnd.n7074 gnd.n569 240.244
R7399 gnd.n7080 gnd.n569 240.244
R7400 gnd.n7080 gnd.n567 240.244
R7401 gnd.n7084 gnd.n567 240.244
R7402 gnd.n7084 gnd.n563 240.244
R7403 gnd.n7090 gnd.n563 240.244
R7404 gnd.n7090 gnd.n561 240.244
R7405 gnd.n7094 gnd.n561 240.244
R7406 gnd.n7094 gnd.n557 240.244
R7407 gnd.n7100 gnd.n557 240.244
R7408 gnd.n7100 gnd.n555 240.244
R7409 gnd.n7104 gnd.n555 240.244
R7410 gnd.n7104 gnd.n551 240.244
R7411 gnd.n7110 gnd.n551 240.244
R7412 gnd.n7110 gnd.n549 240.244
R7413 gnd.n7114 gnd.n549 240.244
R7414 gnd.n7114 gnd.n545 240.244
R7415 gnd.n7120 gnd.n545 240.244
R7416 gnd.n7120 gnd.n543 240.244
R7417 gnd.n7124 gnd.n543 240.244
R7418 gnd.n7124 gnd.n539 240.244
R7419 gnd.n7130 gnd.n539 240.244
R7420 gnd.n7130 gnd.n537 240.244
R7421 gnd.n7134 gnd.n537 240.244
R7422 gnd.n7134 gnd.n533 240.244
R7423 gnd.n7140 gnd.n533 240.244
R7424 gnd.n7140 gnd.n531 240.244
R7425 gnd.n7144 gnd.n531 240.244
R7426 gnd.n7144 gnd.n527 240.244
R7427 gnd.n7150 gnd.n527 240.244
R7428 gnd.n7150 gnd.n525 240.244
R7429 gnd.n7154 gnd.n525 240.244
R7430 gnd.n7160 gnd.n521 240.244
R7431 gnd.n7160 gnd.n519 240.244
R7432 gnd.n7164 gnd.n519 240.244
R7433 gnd.n7164 gnd.n515 240.244
R7434 gnd.n7170 gnd.n515 240.244
R7435 gnd.n7170 gnd.n513 240.244
R7436 gnd.n7174 gnd.n513 240.244
R7437 gnd.n7174 gnd.n509 240.244
R7438 gnd.n7180 gnd.n509 240.244
R7439 gnd.n7180 gnd.n507 240.244
R7440 gnd.n7184 gnd.n507 240.244
R7441 gnd.n7184 gnd.n503 240.244
R7442 gnd.n7190 gnd.n503 240.244
R7443 gnd.n7190 gnd.n501 240.244
R7444 gnd.n7194 gnd.n501 240.244
R7445 gnd.n7194 gnd.n497 240.244
R7446 gnd.n7200 gnd.n497 240.244
R7447 gnd.n7200 gnd.n495 240.244
R7448 gnd.n7204 gnd.n495 240.244
R7449 gnd.n7204 gnd.n491 240.244
R7450 gnd.n7210 gnd.n491 240.244
R7451 gnd.n7210 gnd.n489 240.244
R7452 gnd.n7214 gnd.n489 240.244
R7453 gnd.n7214 gnd.n485 240.244
R7454 gnd.n7220 gnd.n485 240.244
R7455 gnd.n7220 gnd.n483 240.244
R7456 gnd.n7224 gnd.n483 240.244
R7457 gnd.n7224 gnd.n479 240.244
R7458 gnd.n7230 gnd.n479 240.244
R7459 gnd.n7230 gnd.n477 240.244
R7460 gnd.n7234 gnd.n477 240.244
R7461 gnd.n7234 gnd.n473 240.244
R7462 gnd.n7240 gnd.n473 240.244
R7463 gnd.n7240 gnd.n471 240.244
R7464 gnd.n7244 gnd.n471 240.244
R7465 gnd.n7244 gnd.n467 240.244
R7466 gnd.n7250 gnd.n467 240.244
R7467 gnd.n7250 gnd.n465 240.244
R7468 gnd.n7254 gnd.n465 240.244
R7469 gnd.n7254 gnd.n461 240.244
R7470 gnd.n7260 gnd.n461 240.244
R7471 gnd.n7260 gnd.n459 240.244
R7472 gnd.n7264 gnd.n459 240.244
R7473 gnd.n7264 gnd.n455 240.244
R7474 gnd.n7270 gnd.n455 240.244
R7475 gnd.n7270 gnd.n453 240.244
R7476 gnd.n7274 gnd.n453 240.244
R7477 gnd.n7274 gnd.n449 240.244
R7478 gnd.n7280 gnd.n449 240.244
R7479 gnd.n7280 gnd.n447 240.244
R7480 gnd.n7284 gnd.n447 240.244
R7481 gnd.n7284 gnd.n443 240.244
R7482 gnd.n7290 gnd.n443 240.244
R7483 gnd.n7290 gnd.n441 240.244
R7484 gnd.n7294 gnd.n441 240.244
R7485 gnd.n7294 gnd.n437 240.244
R7486 gnd.n7300 gnd.n437 240.244
R7487 gnd.n7300 gnd.n435 240.244
R7488 gnd.n7304 gnd.n435 240.244
R7489 gnd.n7304 gnd.n431 240.244
R7490 gnd.n7310 gnd.n431 240.244
R7491 gnd.n7310 gnd.n429 240.244
R7492 gnd.n7314 gnd.n429 240.244
R7493 gnd.n7314 gnd.n425 240.244
R7494 gnd.n7320 gnd.n425 240.244
R7495 gnd.n7320 gnd.n423 240.244
R7496 gnd.n7324 gnd.n423 240.244
R7497 gnd.n7324 gnd.n419 240.244
R7498 gnd.n7330 gnd.n419 240.244
R7499 gnd.n7330 gnd.n417 240.244
R7500 gnd.n7334 gnd.n417 240.244
R7501 gnd.n7334 gnd.n413 240.244
R7502 gnd.n7340 gnd.n413 240.244
R7503 gnd.n7340 gnd.n411 240.244
R7504 gnd.n7344 gnd.n411 240.244
R7505 gnd.n7344 gnd.n407 240.244
R7506 gnd.n7350 gnd.n407 240.244
R7507 gnd.n7350 gnd.n405 240.244
R7508 gnd.n7354 gnd.n405 240.244
R7509 gnd.n7354 gnd.n401 240.244
R7510 gnd.n7361 gnd.n401 240.244
R7511 gnd.n7361 gnd.n399 240.244
R7512 gnd.n7365 gnd.n399 240.244
R7513 gnd.n7365 gnd.n395 240.244
R7514 gnd.n2761 gnd.n2752 240.244
R7515 gnd.n2762 gnd.n2761 240.244
R7516 gnd.n2763 gnd.n2762 240.244
R7517 gnd.n2763 gnd.n2747 240.244
R7518 gnd.n2856 gnd.n2747 240.244
R7519 gnd.n2856 gnd.n2748 240.244
R7520 gnd.n2769 gnd.n2748 240.244
R7521 gnd.n2776 gnd.n2769 240.244
R7522 gnd.n2848 gnd.n2776 240.244
R7523 gnd.n2848 gnd.n2847 240.244
R7524 gnd.n2847 gnd.n2846 240.244
R7525 gnd.n2846 gnd.n2844 240.244
R7526 gnd.n2844 gnd.n2841 240.244
R7527 gnd.n2841 gnd.n2840 240.244
R7528 gnd.n2840 gnd.n2837 240.244
R7529 gnd.n2837 gnd.n2836 240.244
R7530 gnd.n2836 gnd.n2777 240.244
R7531 gnd.n2832 gnd.n2777 240.244
R7532 gnd.n2832 gnd.n2831 240.244
R7533 gnd.n2831 gnd.n2830 240.244
R7534 gnd.n2830 gnd.n2780 240.244
R7535 gnd.n2826 gnd.n2780 240.244
R7536 gnd.n2826 gnd.n2825 240.244
R7537 gnd.n2825 gnd.n2824 240.244
R7538 gnd.n2824 gnd.n2786 240.244
R7539 gnd.n2820 gnd.n2786 240.244
R7540 gnd.n2820 gnd.n2819 240.244
R7541 gnd.n2819 gnd.n2818 240.244
R7542 gnd.n2818 gnd.n2792 240.244
R7543 gnd.n2814 gnd.n2792 240.244
R7544 gnd.n2814 gnd.n2813 240.244
R7545 gnd.n2813 gnd.n2812 240.244
R7546 gnd.n2812 gnd.n2798 240.244
R7547 gnd.n2808 gnd.n2798 240.244
R7548 gnd.n2808 gnd.n2807 240.244
R7549 gnd.n2807 gnd.n2687 240.244
R7550 gnd.n3198 gnd.n2687 240.244
R7551 gnd.n3199 gnd.n3198 240.244
R7552 gnd.n3199 gnd.n2683 240.244
R7553 gnd.n3205 gnd.n2683 240.244
R7554 gnd.n3206 gnd.n3205 240.244
R7555 gnd.n3207 gnd.n3206 240.244
R7556 gnd.n3207 gnd.n2679 240.244
R7557 gnd.n3213 gnd.n2679 240.244
R7558 gnd.n3214 gnd.n3213 240.244
R7559 gnd.n3216 gnd.n3214 240.244
R7560 gnd.n3216 gnd.n2674 240.244
R7561 gnd.n3227 gnd.n2674 240.244
R7562 gnd.n3227 gnd.n2675 240.244
R7563 gnd.n3223 gnd.n2675 240.244
R7564 gnd.n3223 gnd.n2554 240.244
R7565 gnd.n3394 gnd.n2554 240.244
R7566 gnd.n3394 gnd.n2549 240.244
R7567 gnd.n3402 gnd.n2549 240.244
R7568 gnd.n3402 gnd.n2550 240.244
R7569 gnd.n2550 gnd.n2529 240.244
R7570 gnd.n3424 gnd.n2529 240.244
R7571 gnd.n3424 gnd.n2523 240.244
R7572 gnd.n3438 gnd.n2523 240.244
R7573 gnd.n3438 gnd.n2525 240.244
R7574 gnd.n3434 gnd.n2525 240.244
R7575 gnd.n3434 gnd.n3433 240.244
R7576 gnd.n3433 gnd.n2494 240.244
R7577 gnd.n3471 gnd.n2494 240.244
R7578 gnd.n3471 gnd.n2489 240.244
R7579 gnd.n3479 gnd.n2489 240.244
R7580 gnd.n3479 gnd.n2490 240.244
R7581 gnd.n2490 gnd.n2479 240.244
R7582 gnd.n3593 gnd.n2479 240.244
R7583 gnd.n3593 gnd.n2475 240.244
R7584 gnd.n3599 gnd.n2475 240.244
R7585 gnd.n3599 gnd.n2458 240.244
R7586 gnd.n3620 gnd.n2458 240.244
R7587 gnd.n3620 gnd.n2453 240.244
R7588 gnd.n3628 gnd.n2453 240.244
R7589 gnd.n3628 gnd.n2454 240.244
R7590 gnd.n2454 gnd.n2425 240.244
R7591 gnd.n3662 gnd.n2425 240.244
R7592 gnd.n3662 gnd.n2420 240.244
R7593 gnd.n3679 gnd.n2420 240.244
R7594 gnd.n3679 gnd.n2421 240.244
R7595 gnd.n3675 gnd.n2421 240.244
R7596 gnd.n3675 gnd.n3671 240.244
R7597 gnd.n3671 gnd.n2391 240.244
R7598 gnd.n3745 gnd.n2391 240.244
R7599 gnd.n3745 gnd.n2387 240.244
R7600 gnd.n3751 gnd.n2387 240.244
R7601 gnd.n3751 gnd.n2368 240.244
R7602 gnd.n3788 gnd.n2368 240.244
R7603 gnd.n3788 gnd.n2364 240.244
R7604 gnd.n3794 gnd.n2364 240.244
R7605 gnd.n3794 gnd.n2352 240.244
R7606 gnd.n3836 gnd.n2352 240.244
R7607 gnd.n3836 gnd.n2347 240.244
R7608 gnd.n3844 gnd.n2347 240.244
R7609 gnd.n3844 gnd.n2348 240.244
R7610 gnd.n2348 gnd.n2323 240.244
R7611 gnd.n3873 gnd.n2323 240.244
R7612 gnd.n3873 gnd.n2319 240.244
R7613 gnd.n3879 gnd.n2319 240.244
R7614 gnd.n3879 gnd.n2286 240.244
R7615 gnd.n3907 gnd.n2286 240.244
R7616 gnd.n3907 gnd.n2281 240.244
R7617 gnd.n3915 gnd.n2281 240.244
R7618 gnd.n3915 gnd.n2282 240.244
R7619 gnd.n2282 gnd.n2257 240.244
R7620 gnd.n3959 gnd.n2257 240.244
R7621 gnd.n3959 gnd.n2253 240.244
R7622 gnd.n3965 gnd.n2253 240.244
R7623 gnd.n3965 gnd.n2238 240.244
R7624 gnd.n3985 gnd.n2238 240.244
R7625 gnd.n3985 gnd.n2233 240.244
R7626 gnd.n3993 gnd.n2233 240.244
R7627 gnd.n3993 gnd.n2234 240.244
R7628 gnd.n2234 gnd.n2037 240.244
R7629 gnd.n4177 gnd.n2037 240.244
R7630 gnd.n4177 gnd.n2033 240.244
R7631 gnd.n4183 gnd.n2033 240.244
R7632 gnd.n4183 gnd.n2025 240.244
R7633 gnd.n4198 gnd.n2025 240.244
R7634 gnd.n4198 gnd.n2021 240.244
R7635 gnd.n4204 gnd.n2021 240.244
R7636 gnd.n4204 gnd.n2013 240.244
R7637 gnd.n4219 gnd.n2013 240.244
R7638 gnd.n4219 gnd.n2009 240.244
R7639 gnd.n4225 gnd.n2009 240.244
R7640 gnd.n4225 gnd.n2001 240.244
R7641 gnd.n4242 gnd.n2001 240.244
R7642 gnd.n4242 gnd.n1997 240.244
R7643 gnd.n4249 gnd.n1997 240.244
R7644 gnd.n4249 gnd.n1615 240.244
R7645 gnd.n4623 gnd.n1615 240.244
R7646 gnd.n4623 gnd.n1616 240.244
R7647 gnd.n4619 gnd.n1616 240.244
R7648 gnd.n4619 gnd.n1622 240.244
R7649 gnd.n4615 gnd.n1622 240.244
R7650 gnd.n4615 gnd.n1625 240.244
R7651 gnd.n4611 gnd.n1625 240.244
R7652 gnd.n4611 gnd.n1631 240.244
R7653 gnd.n1813 gnd.n1631 240.244
R7654 gnd.n1819 gnd.n1813 240.244
R7655 gnd.n1820 gnd.n1819 240.244
R7656 gnd.n4349 gnd.n1820 240.244
R7657 gnd.n4349 gnd.n1808 240.244
R7658 gnd.n4357 gnd.n1808 240.244
R7659 gnd.n4357 gnd.n1809 240.244
R7660 gnd.n1809 gnd.n1786 240.244
R7661 gnd.n4380 gnd.n1786 240.244
R7662 gnd.n4380 gnd.n1781 240.244
R7663 gnd.n4388 gnd.n1781 240.244
R7664 gnd.n4388 gnd.n1782 240.244
R7665 gnd.n1782 gnd.n1760 240.244
R7666 gnd.n4413 gnd.n1760 240.244
R7667 gnd.n4413 gnd.n1755 240.244
R7668 gnd.n4421 gnd.n1755 240.244
R7669 gnd.n4421 gnd.n1756 240.244
R7670 gnd.n1756 gnd.n1733 240.244
R7671 gnd.n4450 gnd.n1733 240.244
R7672 gnd.n4450 gnd.n1728 240.244
R7673 gnd.n4475 gnd.n1728 240.244
R7674 gnd.n4475 gnd.n1729 240.244
R7675 gnd.n4471 gnd.n1729 240.244
R7676 gnd.n4471 gnd.n4470 240.244
R7677 gnd.n4470 gnd.n4467 240.244
R7678 gnd.n4467 gnd.n4458 240.244
R7679 gnd.n4462 gnd.n4458 240.244
R7680 gnd.n4462 gnd.n1708 240.244
R7681 gnd.n4533 gnd.n1708 240.244
R7682 gnd.n4533 gnd.n1705 240.244
R7683 gnd.n4540 gnd.n1705 240.244
R7684 gnd.n4540 gnd.n1706 240.244
R7685 gnd.n1706 gnd.n334 240.244
R7686 gnd.n7392 gnd.n334 240.244
R7687 gnd.n7392 gnd.n335 240.244
R7688 gnd.n7387 gnd.n335 240.244
R7689 gnd.n7387 gnd.n7386 240.244
R7690 gnd.n7386 gnd.n7385 240.244
R7691 gnd.n7385 gnd.n339 240.244
R7692 gnd.n7381 gnd.n339 240.244
R7693 gnd.n7381 gnd.n345 240.244
R7694 gnd.n7371 gnd.n345 240.244
R7695 gnd.n6700 gnd.n797 240.244
R7696 gnd.n6696 gnd.n797 240.244
R7697 gnd.n6696 gnd.n802 240.244
R7698 gnd.n6692 gnd.n802 240.244
R7699 gnd.n6692 gnd.n804 240.244
R7700 gnd.n6688 gnd.n804 240.244
R7701 gnd.n6688 gnd.n810 240.244
R7702 gnd.n6684 gnd.n810 240.244
R7703 gnd.n6684 gnd.n812 240.244
R7704 gnd.n6680 gnd.n812 240.244
R7705 gnd.n6680 gnd.n818 240.244
R7706 gnd.n6676 gnd.n818 240.244
R7707 gnd.n6676 gnd.n820 240.244
R7708 gnd.n6672 gnd.n820 240.244
R7709 gnd.n6672 gnd.n826 240.244
R7710 gnd.n6668 gnd.n826 240.244
R7711 gnd.n6668 gnd.n828 240.244
R7712 gnd.n6664 gnd.n828 240.244
R7713 gnd.n6664 gnd.n834 240.244
R7714 gnd.n6660 gnd.n834 240.244
R7715 gnd.n6660 gnd.n836 240.244
R7716 gnd.n6656 gnd.n836 240.244
R7717 gnd.n6656 gnd.n842 240.244
R7718 gnd.n6652 gnd.n842 240.244
R7719 gnd.n6652 gnd.n844 240.244
R7720 gnd.n6648 gnd.n844 240.244
R7721 gnd.n6648 gnd.n850 240.244
R7722 gnd.n6644 gnd.n850 240.244
R7723 gnd.n6644 gnd.n852 240.244
R7724 gnd.n6640 gnd.n852 240.244
R7725 gnd.n6640 gnd.n858 240.244
R7726 gnd.n6636 gnd.n858 240.244
R7727 gnd.n6636 gnd.n860 240.244
R7728 gnd.n6632 gnd.n860 240.244
R7729 gnd.n6632 gnd.n866 240.244
R7730 gnd.n6628 gnd.n866 240.244
R7731 gnd.n6628 gnd.n868 240.244
R7732 gnd.n6624 gnd.n868 240.244
R7733 gnd.n6624 gnd.n874 240.244
R7734 gnd.n6620 gnd.n874 240.244
R7735 gnd.n6620 gnd.n876 240.244
R7736 gnd.n6616 gnd.n876 240.244
R7737 gnd.n6616 gnd.n882 240.244
R7738 gnd.n6612 gnd.n882 240.244
R7739 gnd.n6612 gnd.n884 240.244
R7740 gnd.n6608 gnd.n884 240.244
R7741 gnd.n6608 gnd.n890 240.244
R7742 gnd.n6604 gnd.n890 240.244
R7743 gnd.n6604 gnd.n892 240.244
R7744 gnd.n6600 gnd.n892 240.244
R7745 gnd.n6600 gnd.n898 240.244
R7746 gnd.n6596 gnd.n898 240.244
R7747 gnd.n6596 gnd.n900 240.244
R7748 gnd.n6592 gnd.n900 240.244
R7749 gnd.n6592 gnd.n906 240.244
R7750 gnd.n6588 gnd.n906 240.244
R7751 gnd.n6588 gnd.n908 240.244
R7752 gnd.n6584 gnd.n908 240.244
R7753 gnd.n6584 gnd.n914 240.244
R7754 gnd.n6580 gnd.n914 240.244
R7755 gnd.n6580 gnd.n916 240.244
R7756 gnd.n6576 gnd.n916 240.244
R7757 gnd.n6576 gnd.n922 240.244
R7758 gnd.n6572 gnd.n922 240.244
R7759 gnd.n6572 gnd.n924 240.244
R7760 gnd.n6568 gnd.n924 240.244
R7761 gnd.n6568 gnd.n930 240.244
R7762 gnd.n6564 gnd.n930 240.244
R7763 gnd.n6564 gnd.n932 240.244
R7764 gnd.n6560 gnd.n932 240.244
R7765 gnd.n6560 gnd.n938 240.244
R7766 gnd.n6556 gnd.n938 240.244
R7767 gnd.n6556 gnd.n940 240.244
R7768 gnd.n6552 gnd.n940 240.244
R7769 gnd.n6552 gnd.n946 240.244
R7770 gnd.n6548 gnd.n946 240.244
R7771 gnd.n6548 gnd.n948 240.244
R7772 gnd.n6544 gnd.n948 240.244
R7773 gnd.n6544 gnd.n954 240.244
R7774 gnd.n6540 gnd.n954 240.244
R7775 gnd.n6540 gnd.n956 240.244
R7776 gnd.n6536 gnd.n956 240.244
R7777 gnd.n6536 gnd.n962 240.244
R7778 gnd.n2755 gnd.n962 240.244
R7779 gnd.n3382 gnd.n2564 240.244
R7780 gnd.n3382 gnd.n2565 240.244
R7781 gnd.n2565 gnd.n2545 240.244
R7782 gnd.n3405 gnd.n2545 240.244
R7783 gnd.n3405 gnd.n2539 240.244
R7784 gnd.n3412 gnd.n2539 240.244
R7785 gnd.n3412 gnd.n2540 240.244
R7786 gnd.n2540 gnd.n2519 240.244
R7787 gnd.n3441 gnd.n2519 240.244
R7788 gnd.n3441 gnd.n2515 240.244
R7789 gnd.n3447 gnd.n2515 240.244
R7790 gnd.n3447 gnd.n2504 240.244
R7791 gnd.n3461 gnd.n2504 240.244
R7792 gnd.n3461 gnd.n2498 240.244
R7793 gnd.n3468 gnd.n2498 240.244
R7794 gnd.n3468 gnd.n2499 240.244
R7795 gnd.n2499 gnd.n1527 240.244
R7796 gnd.n4724 gnd.n1527 240.244
R7797 gnd.n4724 gnd.n1528 240.244
R7798 gnd.n1533 gnd.n1528 240.244
R7799 gnd.n1534 gnd.n1533 240.244
R7800 gnd.n1535 gnd.n1534 240.244
R7801 gnd.n2467 gnd.n1535 240.244
R7802 gnd.n2467 gnd.n1538 240.244
R7803 gnd.n1539 gnd.n1538 240.244
R7804 gnd.n1540 gnd.n1539 240.244
R7805 gnd.n2435 gnd.n1540 240.244
R7806 gnd.n2435 gnd.n1543 240.244
R7807 gnd.n1544 gnd.n1543 240.244
R7808 gnd.n1545 gnd.n1544 240.244
R7809 gnd.n3689 gnd.n1545 240.244
R7810 gnd.n3689 gnd.n1548 240.244
R7811 gnd.n1549 gnd.n1548 240.244
R7812 gnd.n1550 gnd.n1549 240.244
R7813 gnd.n2392 gnd.n1550 240.244
R7814 gnd.n2392 gnd.n1553 240.244
R7815 gnd.n1554 gnd.n1553 240.244
R7816 gnd.n1555 gnd.n1554 240.244
R7817 gnd.n3773 gnd.n1555 240.244
R7818 gnd.n3773 gnd.n1558 240.244
R7819 gnd.n1559 gnd.n1558 240.244
R7820 gnd.n1560 gnd.n1559 240.244
R7821 gnd.n3825 gnd.n1560 240.244
R7822 gnd.n3825 gnd.n1563 240.244
R7823 gnd.n1564 gnd.n1563 240.244
R7824 gnd.n1565 gnd.n1564 240.244
R7825 gnd.n3808 gnd.n1565 240.244
R7826 gnd.n3808 gnd.n1568 240.244
R7827 gnd.n1569 gnd.n1568 240.244
R7828 gnd.n1570 gnd.n1569 240.244
R7829 gnd.n2292 gnd.n1570 240.244
R7830 gnd.n2292 gnd.n1573 240.244
R7831 gnd.n1574 gnd.n1573 240.244
R7832 gnd.n1575 gnd.n1574 240.244
R7833 gnd.n3925 gnd.n1575 240.244
R7834 gnd.n3925 gnd.n1578 240.244
R7835 gnd.n1579 gnd.n1578 240.244
R7836 gnd.n1580 gnd.n1579 240.244
R7837 gnd.n2250 gnd.n1580 240.244
R7838 gnd.n2250 gnd.n1583 240.244
R7839 gnd.n1584 gnd.n1583 240.244
R7840 gnd.n1585 gnd.n1584 240.244
R7841 gnd.n3996 gnd.n1585 240.244
R7842 gnd.n3996 gnd.n1588 240.244
R7843 gnd.n1589 gnd.n1588 240.244
R7844 gnd.n1590 gnd.n1589 240.244
R7845 gnd.n4174 gnd.n1590 240.244
R7846 gnd.n4174 gnd.n1593 240.244
R7847 gnd.n1594 gnd.n1593 240.244
R7848 gnd.n1595 gnd.n1594 240.244
R7849 gnd.n4195 gnd.n1595 240.244
R7850 gnd.n4195 gnd.n1598 240.244
R7851 gnd.n1599 gnd.n1598 240.244
R7852 gnd.n1600 gnd.n1599 240.244
R7853 gnd.n4216 gnd.n1600 240.244
R7854 gnd.n4216 gnd.n1603 240.244
R7855 gnd.n1604 gnd.n1603 240.244
R7856 gnd.n1605 gnd.n1604 240.244
R7857 gnd.n4239 gnd.n1605 240.244
R7858 gnd.n4239 gnd.n1608 240.244
R7859 gnd.n1609 gnd.n1608 240.244
R7860 gnd.n4626 gnd.n1609 240.244
R7861 gnd.n2578 gnd.n2577 240.244
R7862 gnd.n2650 gnd.n2578 240.244
R7863 gnd.n2586 gnd.n2585 240.244
R7864 gnd.n2652 gnd.n2595 240.244
R7865 gnd.n2655 gnd.n2596 240.244
R7866 gnd.n2604 gnd.n2603 240.244
R7867 gnd.n2657 gnd.n2613 240.244
R7868 gnd.n2660 gnd.n2614 240.244
R7869 gnd.n2665 gnd.n2664 240.244
R7870 gnd.n2635 gnd.n2634 240.244
R7871 gnd.n2668 gnd.n2636 240.244
R7872 gnd.n2640 gnd.n2639 240.244
R7873 gnd.n2646 gnd.n2641 240.244
R7874 gnd.n2648 gnd.n2647 240.244
R7875 gnd.n3384 gnd.n2561 240.244
R7876 gnd.n3384 gnd.n2556 240.244
R7877 gnd.n3391 gnd.n2556 240.244
R7878 gnd.n3391 gnd.n2547 240.244
R7879 gnd.n2547 gnd.n2536 240.244
R7880 gnd.n3414 gnd.n2536 240.244
R7881 gnd.n3414 gnd.n2531 240.244
R7882 gnd.n3421 gnd.n2531 240.244
R7883 gnd.n3421 gnd.n2521 240.244
R7884 gnd.n2521 gnd.n2512 240.244
R7885 gnd.n3449 gnd.n2512 240.244
R7886 gnd.n3449 gnd.n2506 240.244
R7887 gnd.n3458 gnd.n2506 240.244
R7888 gnd.n3458 gnd.n2507 240.244
R7889 gnd.n2507 gnd.n2496 240.244
R7890 gnd.n2496 gnd.n2488 240.244
R7891 gnd.n3551 gnd.n2488 240.244
R7892 gnd.n3551 gnd.n1525 240.244
R7893 gnd.n3558 gnd.n1525 240.244
R7894 gnd.n3558 gnd.n2482 240.244
R7895 gnd.n2482 gnd.n2465 240.244
R7896 gnd.n3611 gnd.n2465 240.244
R7897 gnd.n3611 gnd.n2461 240.244
R7898 gnd.n3617 gnd.n2461 240.244
R7899 gnd.n3617 gnd.n2444 240.244
R7900 gnd.n3640 gnd.n2444 240.244
R7901 gnd.n3640 gnd.n2438 240.244
R7902 gnd.n3650 gnd.n2438 240.244
R7903 gnd.n3650 gnd.n2439 240.244
R7904 gnd.n3644 gnd.n2439 240.244
R7905 gnd.n3644 gnd.n2409 240.244
R7906 gnd.n3700 gnd.n2409 240.244
R7907 gnd.n3700 gnd.n2403 240.244
R7908 gnd.n3707 gnd.n2403 240.244
R7909 gnd.n3707 gnd.n2404 240.244
R7910 gnd.n2404 gnd.n2384 240.244
R7911 gnd.n3754 gnd.n2384 240.244
R7912 gnd.n3754 gnd.n2378 240.244
R7913 gnd.n3772 gnd.n2378 240.244
R7914 gnd.n3772 gnd.n2379 240.244
R7915 gnd.n3759 gnd.n2379 240.244
R7916 gnd.n3760 gnd.n3759 240.244
R7917 gnd.n3760 gnd.n2360 240.244
R7918 gnd.n3761 gnd.n2360 240.244
R7919 gnd.n3761 gnd.n2338 240.244
R7920 gnd.n3854 gnd.n2338 240.244
R7921 gnd.n3854 gnd.n2333 240.244
R7922 gnd.n3861 gnd.n2333 240.244
R7923 gnd.n3861 gnd.n2316 240.244
R7924 gnd.n3882 gnd.n2316 240.244
R7925 gnd.n3883 gnd.n3882 240.244
R7926 gnd.n3883 gnd.n2312 240.244
R7927 gnd.n3889 gnd.n2312 240.244
R7928 gnd.n3889 gnd.n2272 240.244
R7929 gnd.n3927 gnd.n2272 240.244
R7930 gnd.n3927 gnd.n2267 240.244
R7931 gnd.n3949 gnd.n2267 240.244
R7932 gnd.n3949 gnd.n2260 240.244
R7933 gnd.n3932 gnd.n2260 240.244
R7934 gnd.n3935 gnd.n3932 240.244
R7935 gnd.n3936 gnd.n3935 240.244
R7936 gnd.n3936 gnd.n2240 240.244
R7937 gnd.n2240 gnd.n2232 240.244
R7938 gnd.n2232 gnd.n2042 240.244
R7939 gnd.n4166 gnd.n2042 240.244
R7940 gnd.n4166 gnd.n2038 240.244
R7941 gnd.n4172 gnd.n2038 240.244
R7942 gnd.n4172 gnd.n2031 240.244
R7943 gnd.n4187 gnd.n2031 240.244
R7944 gnd.n4187 gnd.n2027 240.244
R7945 gnd.n4193 gnd.n2027 240.244
R7946 gnd.n4193 gnd.n2019 240.244
R7947 gnd.n4208 gnd.n2019 240.244
R7948 gnd.n4208 gnd.n2015 240.244
R7949 gnd.n4214 gnd.n2015 240.244
R7950 gnd.n4214 gnd.n2007 240.244
R7951 gnd.n4229 gnd.n2007 240.244
R7952 gnd.n4229 gnd.n2003 240.244
R7953 gnd.n4236 gnd.n2003 240.244
R7954 gnd.n4236 gnd.n1996 240.244
R7955 gnd.n4252 gnd.n1996 240.244
R7956 gnd.n4252 gnd.n1613 240.244
R7957 gnd.n1894 gnd.n1893 240.244
R7958 gnd.n1910 gnd.n1909 240.244
R7959 gnd.n1913 gnd.n1912 240.244
R7960 gnd.n1929 gnd.n1928 240.244
R7961 gnd.n1932 gnd.n1931 240.244
R7962 gnd.n1948 gnd.n1947 240.244
R7963 gnd.n1951 gnd.n1950 240.244
R7964 gnd.n1967 gnd.n1966 240.244
R7965 gnd.n1970 gnd.n1969 240.244
R7966 gnd.n1975 gnd.n1972 240.244
R7967 gnd.n1978 gnd.n1977 240.244
R7968 gnd.n1986 gnd.n1980 240.244
R7969 gnd.n1989 gnd.n1988 240.244
R7970 gnd.n1992 gnd.n1991 240.244
R7971 gnd.n1507 gnd.n1506 240.132
R7972 gnd.n4013 gnd.n4012 240.132
R7973 gnd.n6703 gnd.n6702 225.874
R7974 gnd.n6703 gnd.n790 225.874
R7975 gnd.n6711 gnd.n790 225.874
R7976 gnd.n6712 gnd.n6711 225.874
R7977 gnd.n6713 gnd.n6712 225.874
R7978 gnd.n6713 gnd.n784 225.874
R7979 gnd.n6721 gnd.n784 225.874
R7980 gnd.n6722 gnd.n6721 225.874
R7981 gnd.n6723 gnd.n6722 225.874
R7982 gnd.n6723 gnd.n778 225.874
R7983 gnd.n6731 gnd.n778 225.874
R7984 gnd.n6732 gnd.n6731 225.874
R7985 gnd.n6733 gnd.n6732 225.874
R7986 gnd.n6733 gnd.n772 225.874
R7987 gnd.n6741 gnd.n772 225.874
R7988 gnd.n6742 gnd.n6741 225.874
R7989 gnd.n6743 gnd.n6742 225.874
R7990 gnd.n6743 gnd.n766 225.874
R7991 gnd.n6751 gnd.n766 225.874
R7992 gnd.n6752 gnd.n6751 225.874
R7993 gnd.n6753 gnd.n6752 225.874
R7994 gnd.n6753 gnd.n760 225.874
R7995 gnd.n6761 gnd.n760 225.874
R7996 gnd.n6762 gnd.n6761 225.874
R7997 gnd.n6763 gnd.n6762 225.874
R7998 gnd.n6763 gnd.n754 225.874
R7999 gnd.n6771 gnd.n754 225.874
R8000 gnd.n6772 gnd.n6771 225.874
R8001 gnd.n6773 gnd.n6772 225.874
R8002 gnd.n6773 gnd.n748 225.874
R8003 gnd.n6781 gnd.n748 225.874
R8004 gnd.n6782 gnd.n6781 225.874
R8005 gnd.n6783 gnd.n6782 225.874
R8006 gnd.n6783 gnd.n742 225.874
R8007 gnd.n6791 gnd.n742 225.874
R8008 gnd.n6792 gnd.n6791 225.874
R8009 gnd.n6793 gnd.n6792 225.874
R8010 gnd.n6793 gnd.n736 225.874
R8011 gnd.n6801 gnd.n736 225.874
R8012 gnd.n6802 gnd.n6801 225.874
R8013 gnd.n6803 gnd.n6802 225.874
R8014 gnd.n6803 gnd.n730 225.874
R8015 gnd.n6811 gnd.n730 225.874
R8016 gnd.n6812 gnd.n6811 225.874
R8017 gnd.n6813 gnd.n6812 225.874
R8018 gnd.n6813 gnd.n724 225.874
R8019 gnd.n6821 gnd.n724 225.874
R8020 gnd.n6822 gnd.n6821 225.874
R8021 gnd.n6823 gnd.n6822 225.874
R8022 gnd.n6823 gnd.n718 225.874
R8023 gnd.n6831 gnd.n718 225.874
R8024 gnd.n6832 gnd.n6831 225.874
R8025 gnd.n6833 gnd.n6832 225.874
R8026 gnd.n6833 gnd.n712 225.874
R8027 gnd.n6841 gnd.n712 225.874
R8028 gnd.n6842 gnd.n6841 225.874
R8029 gnd.n6843 gnd.n6842 225.874
R8030 gnd.n6843 gnd.n706 225.874
R8031 gnd.n6851 gnd.n706 225.874
R8032 gnd.n6852 gnd.n6851 225.874
R8033 gnd.n6853 gnd.n6852 225.874
R8034 gnd.n6853 gnd.n700 225.874
R8035 gnd.n6861 gnd.n700 225.874
R8036 gnd.n6862 gnd.n6861 225.874
R8037 gnd.n6863 gnd.n6862 225.874
R8038 gnd.n6863 gnd.n694 225.874
R8039 gnd.n6871 gnd.n694 225.874
R8040 gnd.n6872 gnd.n6871 225.874
R8041 gnd.n6873 gnd.n6872 225.874
R8042 gnd.n6873 gnd.n688 225.874
R8043 gnd.n6881 gnd.n688 225.874
R8044 gnd.n6882 gnd.n6881 225.874
R8045 gnd.n6883 gnd.n6882 225.874
R8046 gnd.n6883 gnd.n682 225.874
R8047 gnd.n6891 gnd.n682 225.874
R8048 gnd.n6892 gnd.n6891 225.874
R8049 gnd.n6893 gnd.n6892 225.874
R8050 gnd.n6893 gnd.n676 225.874
R8051 gnd.n6901 gnd.n676 225.874
R8052 gnd.n6902 gnd.n6901 225.874
R8053 gnd.n6903 gnd.n6902 225.874
R8054 gnd.n6903 gnd.n670 225.874
R8055 gnd.n6911 gnd.n670 225.874
R8056 gnd.n6912 gnd.n6911 225.874
R8057 gnd.n6913 gnd.n6912 225.874
R8058 gnd.n6913 gnd.n664 225.874
R8059 gnd.n6921 gnd.n664 225.874
R8060 gnd.n6922 gnd.n6921 225.874
R8061 gnd.n6923 gnd.n6922 225.874
R8062 gnd.n6923 gnd.n658 225.874
R8063 gnd.n6931 gnd.n658 225.874
R8064 gnd.n6932 gnd.n6931 225.874
R8065 gnd.n6933 gnd.n6932 225.874
R8066 gnd.n6933 gnd.n652 225.874
R8067 gnd.n6941 gnd.n652 225.874
R8068 gnd.n6942 gnd.n6941 225.874
R8069 gnd.n6943 gnd.n6942 225.874
R8070 gnd.n6943 gnd.n646 225.874
R8071 gnd.n6951 gnd.n646 225.874
R8072 gnd.n6952 gnd.n6951 225.874
R8073 gnd.n6953 gnd.n6952 225.874
R8074 gnd.n6953 gnd.n640 225.874
R8075 gnd.n6961 gnd.n640 225.874
R8076 gnd.n6962 gnd.n6961 225.874
R8077 gnd.n6963 gnd.n6962 225.874
R8078 gnd.n6963 gnd.n634 225.874
R8079 gnd.n6971 gnd.n634 225.874
R8080 gnd.n6972 gnd.n6971 225.874
R8081 gnd.n6973 gnd.n6972 225.874
R8082 gnd.n6973 gnd.n628 225.874
R8083 gnd.n6981 gnd.n628 225.874
R8084 gnd.n6982 gnd.n6981 225.874
R8085 gnd.n6983 gnd.n6982 225.874
R8086 gnd.n6983 gnd.n622 225.874
R8087 gnd.n6991 gnd.n622 225.874
R8088 gnd.n6992 gnd.n6991 225.874
R8089 gnd.n6993 gnd.n6992 225.874
R8090 gnd.n6993 gnd.n616 225.874
R8091 gnd.n7001 gnd.n616 225.874
R8092 gnd.n7002 gnd.n7001 225.874
R8093 gnd.n7003 gnd.n7002 225.874
R8094 gnd.n7003 gnd.n610 225.874
R8095 gnd.n7011 gnd.n610 225.874
R8096 gnd.n7012 gnd.n7011 225.874
R8097 gnd.n7013 gnd.n7012 225.874
R8098 gnd.n7013 gnd.n604 225.874
R8099 gnd.n7021 gnd.n604 225.874
R8100 gnd.n7022 gnd.n7021 225.874
R8101 gnd.n7023 gnd.n7022 225.874
R8102 gnd.n7023 gnd.n598 225.874
R8103 gnd.n7031 gnd.n598 225.874
R8104 gnd.n7032 gnd.n7031 225.874
R8105 gnd.n7033 gnd.n7032 225.874
R8106 gnd.n7033 gnd.n592 225.874
R8107 gnd.n7041 gnd.n592 225.874
R8108 gnd.n7042 gnd.n7041 225.874
R8109 gnd.n7043 gnd.n7042 225.874
R8110 gnd.n7043 gnd.n586 225.874
R8111 gnd.n7051 gnd.n586 225.874
R8112 gnd.n7052 gnd.n7051 225.874
R8113 gnd.n7053 gnd.n7052 225.874
R8114 gnd.n7053 gnd.n580 225.874
R8115 gnd.n7061 gnd.n580 225.874
R8116 gnd.n7062 gnd.n7061 225.874
R8117 gnd.n7063 gnd.n7062 225.874
R8118 gnd.n7063 gnd.n574 225.874
R8119 gnd.n7071 gnd.n574 225.874
R8120 gnd.n7072 gnd.n7071 225.874
R8121 gnd.n7073 gnd.n7072 225.874
R8122 gnd.n7073 gnd.n568 225.874
R8123 gnd.n7081 gnd.n568 225.874
R8124 gnd.n7082 gnd.n7081 225.874
R8125 gnd.n7083 gnd.n7082 225.874
R8126 gnd.n7083 gnd.n562 225.874
R8127 gnd.n7091 gnd.n562 225.874
R8128 gnd.n7092 gnd.n7091 225.874
R8129 gnd.n7093 gnd.n7092 225.874
R8130 gnd.n7093 gnd.n556 225.874
R8131 gnd.n7101 gnd.n556 225.874
R8132 gnd.n7102 gnd.n7101 225.874
R8133 gnd.n7103 gnd.n7102 225.874
R8134 gnd.n7103 gnd.n550 225.874
R8135 gnd.n7111 gnd.n550 225.874
R8136 gnd.n7112 gnd.n7111 225.874
R8137 gnd.n7113 gnd.n7112 225.874
R8138 gnd.n7113 gnd.n544 225.874
R8139 gnd.n7121 gnd.n544 225.874
R8140 gnd.n7122 gnd.n7121 225.874
R8141 gnd.n7123 gnd.n7122 225.874
R8142 gnd.n7123 gnd.n538 225.874
R8143 gnd.n7131 gnd.n538 225.874
R8144 gnd.n7132 gnd.n7131 225.874
R8145 gnd.n7133 gnd.n7132 225.874
R8146 gnd.n7133 gnd.n532 225.874
R8147 gnd.n7141 gnd.n532 225.874
R8148 gnd.n7142 gnd.n7141 225.874
R8149 gnd.n7143 gnd.n7142 225.874
R8150 gnd.n7143 gnd.n526 225.874
R8151 gnd.n7151 gnd.n526 225.874
R8152 gnd.n7152 gnd.n7151 225.874
R8153 gnd.n7153 gnd.n7152 225.874
R8154 gnd.n5563 gnd.t153 224.174
R8155 gnd.n5162 gnd.t108 224.174
R8156 gnd.n2082 gnd.n2079 199.319
R8157 gnd.n2215 gnd.n2079 199.319
R8158 gnd.n1460 gnd.n1435 199.319
R8159 gnd.n1460 gnd.n1434 199.319
R8160 gnd.n1508 gnd.n1505 186.49
R8161 gnd.n4014 gnd.n4011 186.49
R8162 gnd.n6391 gnd.n6390 185
R8163 gnd.n6389 gnd.n6388 185
R8164 gnd.n6368 gnd.n6367 185
R8165 gnd.n6383 gnd.n6382 185
R8166 gnd.n6381 gnd.n6380 185
R8167 gnd.n6372 gnd.n6371 185
R8168 gnd.n6375 gnd.n6374 185
R8169 gnd.n6359 gnd.n6358 185
R8170 gnd.n6357 gnd.n6356 185
R8171 gnd.n6336 gnd.n6335 185
R8172 gnd.n6351 gnd.n6350 185
R8173 gnd.n6349 gnd.n6348 185
R8174 gnd.n6340 gnd.n6339 185
R8175 gnd.n6343 gnd.n6342 185
R8176 gnd.n6327 gnd.n6326 185
R8177 gnd.n6325 gnd.n6324 185
R8178 gnd.n6304 gnd.n6303 185
R8179 gnd.n6319 gnd.n6318 185
R8180 gnd.n6317 gnd.n6316 185
R8181 gnd.n6308 gnd.n6307 185
R8182 gnd.n6311 gnd.n6310 185
R8183 gnd.n6296 gnd.n6295 185
R8184 gnd.n6294 gnd.n6293 185
R8185 gnd.n6273 gnd.n6272 185
R8186 gnd.n6288 gnd.n6287 185
R8187 gnd.n6286 gnd.n6285 185
R8188 gnd.n6277 gnd.n6276 185
R8189 gnd.n6280 gnd.n6279 185
R8190 gnd.n6264 gnd.n6263 185
R8191 gnd.n6262 gnd.n6261 185
R8192 gnd.n6241 gnd.n6240 185
R8193 gnd.n6256 gnd.n6255 185
R8194 gnd.n6254 gnd.n6253 185
R8195 gnd.n6245 gnd.n6244 185
R8196 gnd.n6248 gnd.n6247 185
R8197 gnd.n6232 gnd.n6231 185
R8198 gnd.n6230 gnd.n6229 185
R8199 gnd.n6209 gnd.n6208 185
R8200 gnd.n6224 gnd.n6223 185
R8201 gnd.n6222 gnd.n6221 185
R8202 gnd.n6213 gnd.n6212 185
R8203 gnd.n6216 gnd.n6215 185
R8204 gnd.n6200 gnd.n6199 185
R8205 gnd.n6198 gnd.n6197 185
R8206 gnd.n6177 gnd.n6176 185
R8207 gnd.n6192 gnd.n6191 185
R8208 gnd.n6190 gnd.n6189 185
R8209 gnd.n6181 gnd.n6180 185
R8210 gnd.n6184 gnd.n6183 185
R8211 gnd.n6169 gnd.n6168 185
R8212 gnd.n6167 gnd.n6166 185
R8213 gnd.n6146 gnd.n6145 185
R8214 gnd.n6161 gnd.n6160 185
R8215 gnd.n6159 gnd.n6158 185
R8216 gnd.n6150 gnd.n6149 185
R8217 gnd.n6153 gnd.n6152 185
R8218 gnd.n5564 gnd.t152 178.987
R8219 gnd.n5163 gnd.t109 178.987
R8220 gnd.n1 gnd.t26 170.774
R8221 gnd.n7 gnd.t47 170.103
R8222 gnd.n6 gnd.t45 170.103
R8223 gnd.n5 gnd.t63 170.103
R8224 gnd.n4 gnd.t30 170.103
R8225 gnd.n3 gnd.t34 170.103
R8226 gnd.n2 gnd.t65 170.103
R8227 gnd.n1 gnd.t28 170.103
R8228 gnd.n4085 gnd.n4084 163.367
R8229 gnd.n4081 gnd.n4080 163.367
R8230 gnd.n4077 gnd.n4076 163.367
R8231 gnd.n4073 gnd.n4072 163.367
R8232 gnd.n4069 gnd.n4068 163.367
R8233 gnd.n4065 gnd.n4064 163.367
R8234 gnd.n4061 gnd.n4060 163.367
R8235 gnd.n4057 gnd.n4056 163.367
R8236 gnd.n4053 gnd.n4052 163.367
R8237 gnd.n4049 gnd.n4048 163.367
R8238 gnd.n4045 gnd.n4044 163.367
R8239 gnd.n4041 gnd.n4040 163.367
R8240 gnd.n4037 gnd.n4036 163.367
R8241 gnd.n4033 gnd.n4032 163.367
R8242 gnd.n4028 gnd.n4027 163.367
R8243 gnd.n4024 gnd.n4023 163.367
R8244 gnd.n4161 gnd.n4160 163.367
R8245 gnd.n4157 gnd.n4156 163.367
R8246 gnd.n4152 gnd.n4151 163.367
R8247 gnd.n4148 gnd.n4147 163.367
R8248 gnd.n4144 gnd.n4143 163.367
R8249 gnd.n4140 gnd.n4139 163.367
R8250 gnd.n4136 gnd.n4135 163.367
R8251 gnd.n4132 gnd.n4131 163.367
R8252 gnd.n4128 gnd.n4127 163.367
R8253 gnd.n4124 gnd.n4123 163.367
R8254 gnd.n4120 gnd.n4119 163.367
R8255 gnd.n4116 gnd.n4115 163.367
R8256 gnd.n4112 gnd.n4111 163.367
R8257 gnd.n4108 gnd.n4107 163.367
R8258 gnd.n4104 gnd.n4103 163.367
R8259 gnd.n4100 gnd.n4099 163.367
R8260 gnd.n3548 gnd.n1524 163.367
R8261 gnd.n3561 gnd.n1524 163.367
R8262 gnd.n3562 gnd.n3561 163.367
R8263 gnd.n3562 gnd.n2481 163.367
R8264 gnd.n3583 gnd.n2481 163.367
R8265 gnd.n3583 gnd.n2474 163.367
R8266 gnd.n3579 gnd.n2474 163.367
R8267 gnd.n3579 gnd.n2466 163.367
R8268 gnd.n3576 gnd.n2466 163.367
R8269 gnd.n3576 gnd.n2460 163.367
R8270 gnd.n2460 gnd.n2451 163.367
R8271 gnd.n2452 gnd.n2451 163.367
R8272 gnd.n2452 gnd.n2445 163.367
R8273 gnd.n3570 gnd.n2445 163.367
R8274 gnd.n3570 gnd.n2437 163.367
R8275 gnd.n3566 gnd.n2437 163.367
R8276 gnd.n3566 gnd.n2427 163.367
R8277 gnd.n2427 gnd.n2418 163.367
R8278 gnd.n3682 gnd.n2418 163.367
R8279 gnd.n3682 gnd.n2416 163.367
R8280 gnd.n3687 gnd.n2416 163.367
R8281 gnd.n3687 gnd.n2411 163.367
R8282 gnd.n2411 gnd.n2401 163.367
R8283 gnd.n3710 gnd.n2401 163.367
R8284 gnd.n3710 gnd.n2399 163.367
R8285 gnd.n3731 gnd.n2399 163.367
R8286 gnd.n3731 gnd.n2394 163.367
R8287 gnd.n3727 gnd.n2394 163.367
R8288 gnd.n3727 gnd.n3723 163.367
R8289 gnd.n3723 gnd.n3722 163.367
R8290 gnd.n3722 gnd.n2376 163.367
R8291 gnd.n2377 gnd.n2376 163.367
R8292 gnd.n2377 gnd.n2369 163.367
R8293 gnd.n3716 gnd.n2369 163.367
R8294 gnd.n3716 gnd.n2362 163.367
R8295 gnd.n3797 gnd.n2362 163.367
R8296 gnd.n3797 gnd.n2359 163.367
R8297 gnd.n3823 gnd.n2359 163.367
R8298 gnd.n3823 gnd.n2353 163.367
R8299 gnd.n3819 gnd.n2353 163.367
R8300 gnd.n3819 gnd.n2346 163.367
R8301 gnd.n3814 gnd.n2346 163.367
R8302 gnd.n3814 gnd.n2340 163.367
R8303 gnd.n3811 gnd.n2340 163.367
R8304 gnd.n3811 gnd.n2332 163.367
R8305 gnd.n3805 gnd.n2332 163.367
R8306 gnd.n3805 gnd.n2325 163.367
R8307 gnd.n3802 gnd.n2325 163.367
R8308 gnd.n3802 gnd.n3801 163.367
R8309 gnd.n3801 gnd.n2294 163.367
R8310 gnd.n3896 gnd.n2294 163.367
R8311 gnd.n3896 gnd.n2288 163.367
R8312 gnd.n3892 gnd.n2288 163.367
R8313 gnd.n3892 gnd.n2280 163.367
R8314 gnd.n2309 gnd.n2280 163.367
R8315 gnd.n2309 gnd.n2274 163.367
R8316 gnd.n2306 gnd.n2274 163.367
R8317 gnd.n2306 gnd.n2266 163.367
R8318 gnd.n2301 gnd.n2266 163.367
R8319 gnd.n2301 gnd.n2259 163.367
R8320 gnd.n2298 gnd.n2259 163.367
R8321 gnd.n2298 gnd.n2252 163.367
R8322 gnd.n2252 gnd.n2243 163.367
R8323 gnd.n3975 gnd.n2243 163.367
R8324 gnd.n3975 gnd.n2241 163.367
R8325 gnd.n3981 gnd.n2241 163.367
R8326 gnd.n3981 gnd.n2231 163.367
R8327 gnd.n2231 gnd.n2223 163.367
R8328 gnd.n4094 gnd.n2223 163.367
R8329 gnd.n4095 gnd.n4094 163.367
R8330 gnd.n1499 gnd.n1498 163.367
R8331 gnd.n4789 gnd.n1498 163.367
R8332 gnd.n4787 gnd.n4786 163.367
R8333 gnd.n4783 gnd.n4782 163.367
R8334 gnd.n4779 gnd.n4778 163.367
R8335 gnd.n4775 gnd.n4774 163.367
R8336 gnd.n4771 gnd.n4770 163.367
R8337 gnd.n4767 gnd.n4766 163.367
R8338 gnd.n4763 gnd.n4762 163.367
R8339 gnd.n4759 gnd.n4758 163.367
R8340 gnd.n4755 gnd.n4754 163.367
R8341 gnd.n4751 gnd.n4750 163.367
R8342 gnd.n4747 gnd.n4746 163.367
R8343 gnd.n4743 gnd.n4742 163.367
R8344 gnd.n4739 gnd.n4738 163.367
R8345 gnd.n4735 gnd.n4734 163.367
R8346 gnd.n4798 gnd.n1465 163.367
R8347 gnd.n3486 gnd.n3485 163.367
R8348 gnd.n3491 gnd.n3490 163.367
R8349 gnd.n3495 gnd.n3494 163.367
R8350 gnd.n3499 gnd.n3498 163.367
R8351 gnd.n3503 gnd.n3502 163.367
R8352 gnd.n3507 gnd.n3506 163.367
R8353 gnd.n3511 gnd.n3510 163.367
R8354 gnd.n3515 gnd.n3514 163.367
R8355 gnd.n3519 gnd.n3518 163.367
R8356 gnd.n3523 gnd.n3522 163.367
R8357 gnd.n3527 gnd.n3526 163.367
R8358 gnd.n3531 gnd.n3530 163.367
R8359 gnd.n3535 gnd.n3534 163.367
R8360 gnd.n3539 gnd.n3538 163.367
R8361 gnd.n3543 gnd.n3542 163.367
R8362 gnd.n4727 gnd.n1500 163.367
R8363 gnd.n4727 gnd.n1522 163.367
R8364 gnd.n3587 gnd.n1522 163.367
R8365 gnd.n3590 gnd.n3587 163.367
R8366 gnd.n3590 gnd.n2472 163.367
R8367 gnd.n3602 gnd.n2472 163.367
R8368 gnd.n3602 gnd.n2469 163.367
R8369 gnd.n3607 gnd.n2469 163.367
R8370 gnd.n3607 gnd.n2470 163.367
R8371 gnd.n2470 gnd.n2449 163.367
R8372 gnd.n3633 gnd.n2449 163.367
R8373 gnd.n3633 gnd.n2447 163.367
R8374 gnd.n3637 gnd.n2447 163.367
R8375 gnd.n3637 gnd.n2434 163.367
R8376 gnd.n3654 gnd.n2434 163.367
R8377 gnd.n3654 gnd.n2429 163.367
R8378 gnd.n3659 gnd.n2429 163.367
R8379 gnd.n3659 gnd.n2432 163.367
R8380 gnd.n2432 gnd.n2415 163.367
R8381 gnd.n3692 gnd.n2415 163.367
R8382 gnd.n3692 gnd.n2412 163.367
R8383 gnd.n3697 gnd.n2412 163.367
R8384 gnd.n3697 gnd.n2413 163.367
R8385 gnd.n2413 gnd.n2398 163.367
R8386 gnd.n3735 gnd.n2398 163.367
R8387 gnd.n3735 gnd.n2395 163.367
R8388 gnd.n3742 gnd.n2395 163.367
R8389 gnd.n3742 gnd.n2396 163.367
R8390 gnd.n3738 gnd.n2396 163.367
R8391 gnd.n3738 gnd.n2374 163.367
R8392 gnd.n3778 gnd.n2374 163.367
R8393 gnd.n3778 gnd.n2371 163.367
R8394 gnd.n3785 gnd.n2371 163.367
R8395 gnd.n3785 gnd.n2372 163.367
R8396 gnd.n3781 gnd.n2372 163.367
R8397 gnd.n3781 gnd.n2357 163.367
R8398 gnd.n3829 gnd.n2357 163.367
R8399 gnd.n3829 gnd.n2355 163.367
R8400 gnd.n3833 gnd.n2355 163.367
R8401 gnd.n3833 gnd.n2344 163.367
R8402 gnd.n3847 gnd.n2344 163.367
R8403 gnd.n3847 gnd.n2342 163.367
R8404 gnd.n3851 gnd.n2342 163.367
R8405 gnd.n3851 gnd.n2330 163.367
R8406 gnd.n3864 gnd.n2330 163.367
R8407 gnd.n3864 gnd.n2327 163.367
R8408 gnd.n3869 gnd.n2327 163.367
R8409 gnd.n3869 gnd.n2328 163.367
R8410 gnd.n2328 gnd.n2291 163.367
R8411 gnd.n3900 gnd.n2291 163.367
R8412 gnd.n3900 gnd.n2289 163.367
R8413 gnd.n3904 gnd.n2289 163.367
R8414 gnd.n3904 gnd.n2278 163.367
R8415 gnd.n3919 gnd.n2278 163.367
R8416 gnd.n3919 gnd.n2276 163.367
R8417 gnd.n3923 gnd.n2276 163.367
R8418 gnd.n3923 gnd.n2264 163.367
R8419 gnd.n3952 gnd.n2264 163.367
R8420 gnd.n3952 gnd.n2262 163.367
R8421 gnd.n3956 gnd.n2262 163.367
R8422 gnd.n3956 gnd.n2249 163.367
R8423 gnd.n3968 gnd.n2249 163.367
R8424 gnd.n3968 gnd.n2246 163.367
R8425 gnd.n3973 gnd.n2246 163.367
R8426 gnd.n3973 gnd.n2247 163.367
R8427 gnd.n2247 gnd.n2229 163.367
R8428 gnd.n3999 gnd.n2229 163.367
R8429 gnd.n3999 gnd.n2226 163.367
R8430 gnd.n4092 gnd.n2226 163.367
R8431 gnd.n4092 gnd.n2227 163.367
R8432 gnd.n4020 gnd.n4019 156.462
R8433 gnd.n6331 gnd.n6299 153.042
R8434 gnd.n6395 gnd.n6394 152.079
R8435 gnd.n6363 gnd.n6362 152.079
R8436 gnd.n6331 gnd.n6330 152.079
R8437 gnd.n1513 gnd.n1512 152
R8438 gnd.n1514 gnd.n1503 152
R8439 gnd.n1516 gnd.n1515 152
R8440 gnd.n1518 gnd.n1501 152
R8441 gnd.n1520 gnd.n1519 152
R8442 gnd.n4018 gnd.n4002 152
R8443 gnd.n4010 gnd.n4003 152
R8444 gnd.n4009 gnd.n4008 152
R8445 gnd.n4007 gnd.n4004 152
R8446 gnd.n4005 gnd.t164 150.546
R8447 gnd.t80 gnd.n6373 147.661
R8448 gnd.t61 gnd.n6341 147.661
R8449 gnd.t75 gnd.n6309 147.661
R8450 gnd.t56 gnd.n6278 147.661
R8451 gnd.t58 gnd.n6246 147.661
R8452 gnd.t73 gnd.n6214 147.661
R8453 gnd.t36 gnd.n6182 147.661
R8454 gnd.t82 gnd.n6151 147.661
R8455 gnd.n2077 gnd.n2060 143.351
R8456 gnd.n1480 gnd.n1464 143.351
R8457 gnd.n4797 gnd.n1464 143.351
R8458 gnd.n2219 gnd.n2218 133.44
R8459 gnd.n4800 gnd.n4799 133.44
R8460 gnd.n1510 gnd.t83 130.484
R8461 gnd.n1519 gnd.t184 126.766
R8462 gnd.n1517 gnd.t138 126.766
R8463 gnd.n1503 gnd.t173 126.766
R8464 gnd.n1511 gnd.t167 126.766
R8465 gnd.n4006 gnd.t170 126.766
R8466 gnd.n4008 gnd.t135 126.766
R8467 gnd.n4017 gnd.t181 126.766
R8468 gnd.n4019 gnd.t157 126.766
R8469 gnd.n7161 gnd.n520 122.392
R8470 gnd.n7162 gnd.n7161 122.392
R8471 gnd.n7163 gnd.n7162 122.392
R8472 gnd.n7163 gnd.n514 122.392
R8473 gnd.n7171 gnd.n514 122.392
R8474 gnd.n7172 gnd.n7171 122.392
R8475 gnd.n7173 gnd.n7172 122.392
R8476 gnd.n7173 gnd.n508 122.392
R8477 gnd.n7181 gnd.n508 122.392
R8478 gnd.n7182 gnd.n7181 122.392
R8479 gnd.n7183 gnd.n7182 122.392
R8480 gnd.n7183 gnd.n502 122.392
R8481 gnd.n7191 gnd.n502 122.392
R8482 gnd.n7192 gnd.n7191 122.392
R8483 gnd.n7193 gnd.n7192 122.392
R8484 gnd.n7193 gnd.n496 122.392
R8485 gnd.n7201 gnd.n496 122.392
R8486 gnd.n7202 gnd.n7201 122.392
R8487 gnd.n7203 gnd.n7202 122.392
R8488 gnd.n7203 gnd.n490 122.392
R8489 gnd.n7211 gnd.n490 122.392
R8490 gnd.n7212 gnd.n7211 122.392
R8491 gnd.n7213 gnd.n7212 122.392
R8492 gnd.n7213 gnd.n484 122.392
R8493 gnd.n7221 gnd.n484 122.392
R8494 gnd.n7222 gnd.n7221 122.392
R8495 gnd.n7223 gnd.n7222 122.392
R8496 gnd.n7223 gnd.n478 122.392
R8497 gnd.n7231 gnd.n478 122.392
R8498 gnd.n7232 gnd.n7231 122.392
R8499 gnd.n7233 gnd.n7232 122.392
R8500 gnd.n7233 gnd.n472 122.392
R8501 gnd.n7241 gnd.n472 122.392
R8502 gnd.n7242 gnd.n7241 122.392
R8503 gnd.n7243 gnd.n7242 122.392
R8504 gnd.n7243 gnd.n466 122.392
R8505 gnd.n7251 gnd.n466 122.392
R8506 gnd.n7252 gnd.n7251 122.392
R8507 gnd.n7253 gnd.n7252 122.392
R8508 gnd.n7253 gnd.n460 122.392
R8509 gnd.n7261 gnd.n460 122.392
R8510 gnd.n7262 gnd.n7261 122.392
R8511 gnd.n7263 gnd.n7262 122.392
R8512 gnd.n7263 gnd.n454 122.392
R8513 gnd.n7271 gnd.n454 122.392
R8514 gnd.n7272 gnd.n7271 122.392
R8515 gnd.n7273 gnd.n7272 122.392
R8516 gnd.n7273 gnd.n448 122.392
R8517 gnd.n7281 gnd.n448 122.392
R8518 gnd.n7282 gnd.n7281 122.392
R8519 gnd.n7283 gnd.n7282 122.392
R8520 gnd.n7283 gnd.n442 122.392
R8521 gnd.n7291 gnd.n442 122.392
R8522 gnd.n7292 gnd.n7291 122.392
R8523 gnd.n7293 gnd.n7292 122.392
R8524 gnd.n7293 gnd.n436 122.392
R8525 gnd.n7301 gnd.n436 122.392
R8526 gnd.n7302 gnd.n7301 122.392
R8527 gnd.n7303 gnd.n7302 122.392
R8528 gnd.n7303 gnd.n430 122.392
R8529 gnd.n7311 gnd.n430 122.392
R8530 gnd.n7312 gnd.n7311 122.392
R8531 gnd.n7313 gnd.n7312 122.392
R8532 gnd.n7313 gnd.n424 122.392
R8533 gnd.n7321 gnd.n424 122.392
R8534 gnd.n7322 gnd.n7321 122.392
R8535 gnd.n7323 gnd.n7322 122.392
R8536 gnd.n7323 gnd.n418 122.392
R8537 gnd.n7331 gnd.n418 122.392
R8538 gnd.n7332 gnd.n7331 122.392
R8539 gnd.n7333 gnd.n7332 122.392
R8540 gnd.n7333 gnd.n412 122.392
R8541 gnd.n7341 gnd.n412 122.392
R8542 gnd.n7342 gnd.n7341 122.392
R8543 gnd.n7343 gnd.n7342 122.392
R8544 gnd.n7343 gnd.n406 122.392
R8545 gnd.n7351 gnd.n406 122.392
R8546 gnd.n7352 gnd.n7351 122.392
R8547 gnd.n7353 gnd.n7352 122.392
R8548 gnd.n7353 gnd.n400 122.392
R8549 gnd.n7362 gnd.n400 122.392
R8550 gnd.n7363 gnd.n7362 122.392
R8551 gnd.n7364 gnd.n7363 122.392
R8552 gnd.n6390 gnd.n6389 104.615
R8553 gnd.n6389 gnd.n6367 104.615
R8554 gnd.n6382 gnd.n6367 104.615
R8555 gnd.n6382 gnd.n6381 104.615
R8556 gnd.n6381 gnd.n6371 104.615
R8557 gnd.n6374 gnd.n6371 104.615
R8558 gnd.n6358 gnd.n6357 104.615
R8559 gnd.n6357 gnd.n6335 104.615
R8560 gnd.n6350 gnd.n6335 104.615
R8561 gnd.n6350 gnd.n6349 104.615
R8562 gnd.n6349 gnd.n6339 104.615
R8563 gnd.n6342 gnd.n6339 104.615
R8564 gnd.n6326 gnd.n6325 104.615
R8565 gnd.n6325 gnd.n6303 104.615
R8566 gnd.n6318 gnd.n6303 104.615
R8567 gnd.n6318 gnd.n6317 104.615
R8568 gnd.n6317 gnd.n6307 104.615
R8569 gnd.n6310 gnd.n6307 104.615
R8570 gnd.n6295 gnd.n6294 104.615
R8571 gnd.n6294 gnd.n6272 104.615
R8572 gnd.n6287 gnd.n6272 104.615
R8573 gnd.n6287 gnd.n6286 104.615
R8574 gnd.n6286 gnd.n6276 104.615
R8575 gnd.n6279 gnd.n6276 104.615
R8576 gnd.n6263 gnd.n6262 104.615
R8577 gnd.n6262 gnd.n6240 104.615
R8578 gnd.n6255 gnd.n6240 104.615
R8579 gnd.n6255 gnd.n6254 104.615
R8580 gnd.n6254 gnd.n6244 104.615
R8581 gnd.n6247 gnd.n6244 104.615
R8582 gnd.n6231 gnd.n6230 104.615
R8583 gnd.n6230 gnd.n6208 104.615
R8584 gnd.n6223 gnd.n6208 104.615
R8585 gnd.n6223 gnd.n6222 104.615
R8586 gnd.n6222 gnd.n6212 104.615
R8587 gnd.n6215 gnd.n6212 104.615
R8588 gnd.n6199 gnd.n6198 104.615
R8589 gnd.n6198 gnd.n6176 104.615
R8590 gnd.n6191 gnd.n6176 104.615
R8591 gnd.n6191 gnd.n6190 104.615
R8592 gnd.n6190 gnd.n6180 104.615
R8593 gnd.n6183 gnd.n6180 104.615
R8594 gnd.n6168 gnd.n6167 104.615
R8595 gnd.n6167 gnd.n6145 104.615
R8596 gnd.n6160 gnd.n6145 104.615
R8597 gnd.n6160 gnd.n6159 104.615
R8598 gnd.n6159 gnd.n6149 104.615
R8599 gnd.n6152 gnd.n6149 104.615
R8600 gnd.n5713 gnd.t89 100.632
R8601 gnd.n5136 gnd.t126 100.632
R8602 gnd.n7658 gnd.n134 99.6594
R8603 gnd.n7656 gnd.n7655 99.6594
R8604 gnd.n7651 gnd.n141 99.6594
R8605 gnd.n7649 gnd.n7648 99.6594
R8606 gnd.n7644 gnd.n148 99.6594
R8607 gnd.n7642 gnd.n7641 99.6594
R8608 gnd.n7637 gnd.n155 99.6594
R8609 gnd.n7635 gnd.n7634 99.6594
R8610 gnd.n7627 gnd.n162 99.6594
R8611 gnd.n7625 gnd.n7624 99.6594
R8612 gnd.n7620 gnd.n169 99.6594
R8613 gnd.n7618 gnd.n7617 99.6594
R8614 gnd.n7613 gnd.n176 99.6594
R8615 gnd.n7611 gnd.n7610 99.6594
R8616 gnd.n7606 gnd.n183 99.6594
R8617 gnd.n7604 gnd.n7603 99.6594
R8618 gnd.n7599 gnd.n190 99.6594
R8619 gnd.n7597 gnd.n7596 99.6594
R8620 gnd.n195 gnd.n194 99.6594
R8621 gnd.n2099 gnd.n2098 99.6594
R8622 gnd.n2107 gnd.n2106 99.6594
R8623 gnd.n2110 gnd.n2109 99.6594
R8624 gnd.n2117 gnd.n2116 99.6594
R8625 gnd.n2120 gnd.n2119 99.6594
R8626 gnd.n2128 gnd.n2127 99.6594
R8627 gnd.n2131 gnd.n2130 99.6594
R8628 gnd.n2083 gnd.n2082 99.6594
R8629 gnd.n2214 gnd.n2213 99.6594
R8630 gnd.n2207 gnd.n2141 99.6594
R8631 gnd.n2206 gnd.n2205 99.6594
R8632 gnd.n2199 gnd.n2147 99.6594
R8633 gnd.n2198 gnd.n2197 99.6594
R8634 gnd.n2191 gnd.n2153 99.6594
R8635 gnd.n2190 gnd.n2189 99.6594
R8636 gnd.n2183 gnd.n2159 99.6594
R8637 gnd.n2182 gnd.n2181 99.6594
R8638 gnd.n2173 gnd.n2165 99.6594
R8639 gnd.n4828 gnd.n4827 99.6594
R8640 gnd.n4823 gnd.n1441 99.6594
R8641 gnd.n4819 gnd.n1440 99.6594
R8642 gnd.n4815 gnd.n1439 99.6594
R8643 gnd.n4811 gnd.n1438 99.6594
R8644 gnd.n4807 gnd.n1437 99.6594
R8645 gnd.n4803 gnd.n1436 99.6594
R8646 gnd.n3275 gnd.n1434 99.6594
R8647 gnd.n3282 gnd.n1433 99.6594
R8648 gnd.n3286 gnd.n1432 99.6594
R8649 gnd.n3292 gnd.n1431 99.6594
R8650 gnd.n3296 gnd.n1430 99.6594
R8651 gnd.n3302 gnd.n1429 99.6594
R8652 gnd.n3306 gnd.n1428 99.6594
R8653 gnd.n3312 gnd.n1427 99.6594
R8654 gnd.n3316 gnd.n1426 99.6594
R8655 gnd.n3321 gnd.n1425 99.6594
R8656 gnd.n2624 gnd.n1424 99.6594
R8657 gnd.n5106 gnd.n5105 99.6594
R8658 gnd.n5100 gnd.n1012 99.6594
R8659 gnd.n5097 gnd.n1013 99.6594
R8660 gnd.n5093 gnd.n1014 99.6594
R8661 gnd.n5089 gnd.n1015 99.6594
R8662 gnd.n5085 gnd.n1016 99.6594
R8663 gnd.n5081 gnd.n1017 99.6594
R8664 gnd.n5077 gnd.n1018 99.6594
R8665 gnd.n5073 gnd.n1019 99.6594
R8666 gnd.n5068 gnd.n1020 99.6594
R8667 gnd.n5064 gnd.n1021 99.6594
R8668 gnd.n5060 gnd.n1022 99.6594
R8669 gnd.n5056 gnd.n1023 99.6594
R8670 gnd.n5052 gnd.n1024 99.6594
R8671 gnd.n5048 gnd.n1025 99.6594
R8672 gnd.n5044 gnd.n1026 99.6594
R8673 gnd.n5040 gnd.n1027 99.6594
R8674 gnd.n5036 gnd.n1028 99.6594
R8675 gnd.n1083 gnd.n1029 99.6594
R8676 gnd.n6510 gnd.n6509 99.6594
R8677 gnd.n6505 gnd.n5114 99.6594
R8678 gnd.n6501 gnd.n5113 99.6594
R8679 gnd.n6497 gnd.n5112 99.6594
R8680 gnd.n6493 gnd.n5111 99.6594
R8681 gnd.n6489 gnd.n5110 99.6594
R8682 gnd.n6485 gnd.n5109 99.6594
R8683 gnd.n5134 gnd.n5108 99.6594
R8684 gnd.n5746 gnd.n5745 99.6594
R8685 gnd.n5740 gnd.n5688 99.6594
R8686 gnd.n5737 gnd.n5689 99.6594
R8687 gnd.n5733 gnd.n5690 99.6594
R8688 gnd.n5729 gnd.n5691 99.6594
R8689 gnd.n5725 gnd.n5692 99.6594
R8690 gnd.n5721 gnd.n5693 99.6594
R8691 gnd.n5717 gnd.n5694 99.6594
R8692 gnd.n6475 gnd.n999 99.6594
R8693 gnd.n6471 gnd.n1000 99.6594
R8694 gnd.n6467 gnd.n1001 99.6594
R8695 gnd.n6463 gnd.n1002 99.6594
R8696 gnd.n6459 gnd.n1003 99.6594
R8697 gnd.n6455 gnd.n1004 99.6594
R8698 gnd.n6451 gnd.n1005 99.6594
R8699 gnd.n6447 gnd.n1006 99.6594
R8700 gnd.n6443 gnd.n1007 99.6594
R8701 gnd.n6439 gnd.n1008 99.6594
R8702 gnd.n6435 gnd.n1009 99.6594
R8703 gnd.n6431 gnd.n1010 99.6594
R8704 gnd.n6427 gnd.n1011 99.6594
R8705 gnd.n5618 gnd.n5528 99.6594
R8706 gnd.n5616 gnd.n5531 99.6594
R8707 gnd.n5612 gnd.n5611 99.6594
R8708 gnd.n5605 gnd.n5536 99.6594
R8709 gnd.n5604 gnd.n5603 99.6594
R8710 gnd.n5597 gnd.n5542 99.6594
R8711 gnd.n5596 gnd.n5595 99.6594
R8712 gnd.n5589 gnd.n5548 99.6594
R8713 gnd.n5588 gnd.n5587 99.6594
R8714 gnd.n5581 gnd.n5554 99.6594
R8715 gnd.n5580 gnd.n5579 99.6594
R8716 gnd.n5572 gnd.n5560 99.6594
R8717 gnd.n5571 gnd.n5570 99.6594
R8718 gnd.n7513 gnd.n7512 99.6594
R8719 gnd.n7518 gnd.n7517 99.6594
R8720 gnd.n7521 gnd.n7520 99.6594
R8721 gnd.n7526 gnd.n7525 99.6594
R8722 gnd.n7529 gnd.n7528 99.6594
R8723 gnd.n7534 gnd.n7533 99.6594
R8724 gnd.n7537 gnd.n7536 99.6594
R8725 gnd.n7542 gnd.n7540 99.6594
R8726 gnd.n7668 gnd.n121 99.6594
R8727 gnd.n1881 gnd.n1880 99.6594
R8728 gnd.n1900 gnd.n1899 99.6594
R8729 gnd.n1903 gnd.n1902 99.6594
R8730 gnd.n1919 gnd.n1918 99.6594
R8731 gnd.n1922 gnd.n1921 99.6594
R8732 gnd.n1938 gnd.n1937 99.6594
R8733 gnd.n1941 gnd.n1940 99.6594
R8734 gnd.n1957 gnd.n1956 99.6594
R8735 gnd.n1960 gnd.n1959 99.6594
R8736 gnd.n2571 gnd.n1414 99.6594
R8737 gnd.n2581 gnd.n1415 99.6594
R8738 gnd.n2589 gnd.n1416 99.6594
R8739 gnd.n2591 gnd.n1417 99.6594
R8740 gnd.n2599 gnd.n1418 99.6594
R8741 gnd.n2607 gnd.n1419 99.6594
R8742 gnd.n2609 gnd.n1420 99.6594
R8743 gnd.n2617 gnd.n1421 99.6594
R8744 gnd.n3331 gnd.n1422 99.6594
R8745 gnd.n2975 gnd.n1030 99.6594
R8746 gnd.n2972 gnd.n1031 99.6594
R8747 gnd.n2968 gnd.n1032 99.6594
R8748 gnd.n2964 gnd.n1033 99.6594
R8749 gnd.n2960 gnd.n1034 99.6594
R8750 gnd.n2956 gnd.n1035 99.6594
R8751 gnd.n2952 gnd.n1036 99.6594
R8752 gnd.n2948 gnd.n1037 99.6594
R8753 gnd.n2944 gnd.n1038 99.6594
R8754 gnd.n2973 gnd.n1030 99.6594
R8755 gnd.n2969 gnd.n1031 99.6594
R8756 gnd.n2965 gnd.n1032 99.6594
R8757 gnd.n2961 gnd.n1033 99.6594
R8758 gnd.n2957 gnd.n1034 99.6594
R8759 gnd.n2953 gnd.n1035 99.6594
R8760 gnd.n2949 gnd.n1036 99.6594
R8761 gnd.n2945 gnd.n1037 99.6594
R8762 gnd.n2933 gnd.n1038 99.6594
R8763 gnd.n2621 gnd.n1422 99.6594
R8764 gnd.n2610 gnd.n1421 99.6594
R8765 gnd.n2608 gnd.n1420 99.6594
R8766 gnd.n2600 gnd.n1419 99.6594
R8767 gnd.n2592 gnd.n1418 99.6594
R8768 gnd.n2590 gnd.n1417 99.6594
R8769 gnd.n2582 gnd.n1416 99.6594
R8770 gnd.n2572 gnd.n1415 99.6594
R8771 gnd.n2570 gnd.n1414 99.6594
R8772 gnd.n1880 gnd.n1876 99.6594
R8773 gnd.n1901 gnd.n1900 99.6594
R8774 gnd.n1902 gnd.n1867 99.6594
R8775 gnd.n1920 gnd.n1919 99.6594
R8776 gnd.n1921 gnd.n1858 99.6594
R8777 gnd.n1939 gnd.n1938 99.6594
R8778 gnd.n1940 gnd.n1849 99.6594
R8779 gnd.n1958 gnd.n1957 99.6594
R8780 gnd.n1959 gnd.n1838 99.6594
R8781 gnd.n7541 gnd.n121 99.6594
R8782 gnd.n7540 gnd.n7539 99.6594
R8783 gnd.n7536 gnd.n7535 99.6594
R8784 gnd.n7533 gnd.n7532 99.6594
R8785 gnd.n7528 gnd.n7527 99.6594
R8786 gnd.n7525 gnd.n7524 99.6594
R8787 gnd.n7520 gnd.n7519 99.6594
R8788 gnd.n7517 gnd.n7516 99.6594
R8789 gnd.n7512 gnd.n7511 99.6594
R8790 gnd.n5619 gnd.n5618 99.6594
R8791 gnd.n5613 gnd.n5531 99.6594
R8792 gnd.n5611 gnd.n5610 99.6594
R8793 gnd.n5606 gnd.n5605 99.6594
R8794 gnd.n5603 gnd.n5602 99.6594
R8795 gnd.n5598 gnd.n5597 99.6594
R8796 gnd.n5595 gnd.n5594 99.6594
R8797 gnd.n5590 gnd.n5589 99.6594
R8798 gnd.n5587 gnd.n5586 99.6594
R8799 gnd.n5582 gnd.n5581 99.6594
R8800 gnd.n5579 gnd.n5578 99.6594
R8801 gnd.n5573 gnd.n5572 99.6594
R8802 gnd.n5570 gnd.n5526 99.6594
R8803 gnd.n6430 gnd.n1011 99.6594
R8804 gnd.n6434 gnd.n1010 99.6594
R8805 gnd.n6438 gnd.n1009 99.6594
R8806 gnd.n6442 gnd.n1008 99.6594
R8807 gnd.n6446 gnd.n1007 99.6594
R8808 gnd.n6450 gnd.n1006 99.6594
R8809 gnd.n6454 gnd.n1005 99.6594
R8810 gnd.n6458 gnd.n1004 99.6594
R8811 gnd.n6462 gnd.n1003 99.6594
R8812 gnd.n6466 gnd.n1002 99.6594
R8813 gnd.n6470 gnd.n1001 99.6594
R8814 gnd.n6474 gnd.n1000 99.6594
R8815 gnd.n5140 gnd.n999 99.6594
R8816 gnd.n5746 gnd.n5696 99.6594
R8817 gnd.n5738 gnd.n5688 99.6594
R8818 gnd.n5734 gnd.n5689 99.6594
R8819 gnd.n5730 gnd.n5690 99.6594
R8820 gnd.n5726 gnd.n5691 99.6594
R8821 gnd.n5722 gnd.n5692 99.6594
R8822 gnd.n5718 gnd.n5693 99.6594
R8823 gnd.n5694 gnd.n5488 99.6594
R8824 gnd.n6484 gnd.n5108 99.6594
R8825 gnd.n6488 gnd.n5109 99.6594
R8826 gnd.n6492 gnd.n5110 99.6594
R8827 gnd.n6496 gnd.n5111 99.6594
R8828 gnd.n6500 gnd.n5112 99.6594
R8829 gnd.n6504 gnd.n5113 99.6594
R8830 gnd.n5116 gnd.n5114 99.6594
R8831 gnd.n6510 gnd.n5115 99.6594
R8832 gnd.n5106 gnd.n1042 99.6594
R8833 gnd.n5098 gnd.n1012 99.6594
R8834 gnd.n5094 gnd.n1013 99.6594
R8835 gnd.n5090 gnd.n1014 99.6594
R8836 gnd.n5086 gnd.n1015 99.6594
R8837 gnd.n5082 gnd.n1016 99.6594
R8838 gnd.n5078 gnd.n1017 99.6594
R8839 gnd.n5074 gnd.n1018 99.6594
R8840 gnd.n5069 gnd.n1019 99.6594
R8841 gnd.n5065 gnd.n1020 99.6594
R8842 gnd.n5061 gnd.n1021 99.6594
R8843 gnd.n5057 gnd.n1022 99.6594
R8844 gnd.n5053 gnd.n1023 99.6594
R8845 gnd.n5049 gnd.n1024 99.6594
R8846 gnd.n5045 gnd.n1025 99.6594
R8847 gnd.n5041 gnd.n1026 99.6594
R8848 gnd.n5037 gnd.n1027 99.6594
R8849 gnd.n1082 gnd.n1028 99.6594
R8850 gnd.n5029 gnd.n1029 99.6594
R8851 gnd.n3266 gnd.n1424 99.6594
R8852 gnd.n3315 gnd.n1425 99.6594
R8853 gnd.n3313 gnd.n1426 99.6594
R8854 gnd.n3305 gnd.n1427 99.6594
R8855 gnd.n3303 gnd.n1428 99.6594
R8856 gnd.n3295 gnd.n1429 99.6594
R8857 gnd.n3293 gnd.n1430 99.6594
R8858 gnd.n3285 gnd.n1431 99.6594
R8859 gnd.n3283 gnd.n1432 99.6594
R8860 gnd.n3276 gnd.n1433 99.6594
R8861 gnd.n4802 gnd.n1435 99.6594
R8862 gnd.n4806 gnd.n1436 99.6594
R8863 gnd.n4810 gnd.n1437 99.6594
R8864 gnd.n4814 gnd.n1438 99.6594
R8865 gnd.n4818 gnd.n1439 99.6594
R8866 gnd.n4822 gnd.n1440 99.6594
R8867 gnd.n1442 gnd.n1441 99.6594
R8868 gnd.n4828 gnd.n1411 99.6594
R8869 gnd.n2100 gnd.n2099 99.6594
R8870 gnd.n2108 gnd.n2107 99.6594
R8871 gnd.n2109 gnd.n2089 99.6594
R8872 gnd.n2118 gnd.n2117 99.6594
R8873 gnd.n2119 gnd.n2085 99.6594
R8874 gnd.n2129 gnd.n2128 99.6594
R8875 gnd.n2132 gnd.n2131 99.6594
R8876 gnd.n2216 gnd.n2215 99.6594
R8877 gnd.n2213 gnd.n2212 99.6594
R8878 gnd.n2208 gnd.n2207 99.6594
R8879 gnd.n2205 gnd.n2204 99.6594
R8880 gnd.n2200 gnd.n2199 99.6594
R8881 gnd.n2197 gnd.n2196 99.6594
R8882 gnd.n2192 gnd.n2191 99.6594
R8883 gnd.n2189 gnd.n2188 99.6594
R8884 gnd.n2184 gnd.n2183 99.6594
R8885 gnd.n2181 gnd.n2180 99.6594
R8886 gnd.n2174 gnd.n2173 99.6594
R8887 gnd.n194 gnd.n191 99.6594
R8888 gnd.n7598 gnd.n7597 99.6594
R8889 gnd.n190 gnd.n184 99.6594
R8890 gnd.n7605 gnd.n7604 99.6594
R8891 gnd.n183 gnd.n177 99.6594
R8892 gnd.n7612 gnd.n7611 99.6594
R8893 gnd.n176 gnd.n170 99.6594
R8894 gnd.n7619 gnd.n7618 99.6594
R8895 gnd.n169 gnd.n163 99.6594
R8896 gnd.n7626 gnd.n7625 99.6594
R8897 gnd.n162 gnd.n156 99.6594
R8898 gnd.n7636 gnd.n7635 99.6594
R8899 gnd.n155 gnd.n149 99.6594
R8900 gnd.n7643 gnd.n7642 99.6594
R8901 gnd.n148 gnd.n142 99.6594
R8902 gnd.n7650 gnd.n7649 99.6594
R8903 gnd.n141 gnd.n135 99.6594
R8904 gnd.n7657 gnd.n7656 99.6594
R8905 gnd.n134 gnd.n131 99.6594
R8906 gnd.n3230 gnd.n3229 99.6594
R8907 gnd.n2651 gnd.n2650 99.6594
R8908 gnd.n2653 gnd.n2586 99.6594
R8909 gnd.n2654 gnd.n2595 99.6594
R8910 gnd.n2656 gnd.n2655 99.6594
R8911 gnd.n2658 gnd.n2604 99.6594
R8912 gnd.n2659 gnd.n2613 99.6594
R8913 gnd.n2661 gnd.n2660 99.6594
R8914 gnd.n2666 gnd.n2665 99.6594
R8915 gnd.n2667 gnd.n2635 99.6594
R8916 gnd.n2669 gnd.n2668 99.6594
R8917 gnd.n2670 gnd.n2640 99.6594
R8918 gnd.n2671 gnd.n2646 99.6594
R8919 gnd.n3232 gnd.n2648 99.6594
R8920 gnd.n3230 gnd.n2577 99.6594
R8921 gnd.n2651 gnd.n2585 99.6594
R8922 gnd.n2653 gnd.n2652 99.6594
R8923 gnd.n2654 gnd.n2596 99.6594
R8924 gnd.n2656 gnd.n2603 99.6594
R8925 gnd.n2658 gnd.n2657 99.6594
R8926 gnd.n2659 gnd.n2614 99.6594
R8927 gnd.n2664 gnd.n2661 99.6594
R8928 gnd.n2666 gnd.n2634 99.6594
R8929 gnd.n2667 gnd.n2636 99.6594
R8930 gnd.n2669 gnd.n2639 99.6594
R8931 gnd.n2670 gnd.n2641 99.6594
R8932 gnd.n2671 gnd.n2647 99.6594
R8933 gnd.n3233 gnd.n3232 99.6594
R8934 gnd.n1894 gnd.n1892 99.6594
R8935 gnd.n1909 gnd.n1872 99.6594
R8936 gnd.n1913 gnd.n1911 99.6594
R8937 gnd.n1928 gnd.n1863 99.6594
R8938 gnd.n1932 gnd.n1930 99.6594
R8939 gnd.n1947 gnd.n1854 99.6594
R8940 gnd.n1951 gnd.n1949 99.6594
R8941 gnd.n1966 gnd.n1845 99.6594
R8942 gnd.n1969 gnd.n1968 99.6594
R8943 gnd.n1972 gnd.n1971 99.6594
R8944 gnd.n1977 gnd.n1976 99.6594
R8945 gnd.n1980 gnd.n1979 99.6594
R8946 gnd.n1988 gnd.n1987 99.6594
R8947 gnd.n1991 gnd.n1990 99.6594
R8948 gnd.n1990 gnd.n1989 99.6594
R8949 gnd.n1987 gnd.n1986 99.6594
R8950 gnd.n1979 gnd.n1978 99.6594
R8951 gnd.n1976 gnd.n1975 99.6594
R8952 gnd.n1971 gnd.n1970 99.6594
R8953 gnd.n1968 gnd.n1967 99.6594
R8954 gnd.n1950 gnd.n1845 99.6594
R8955 gnd.n1949 gnd.n1948 99.6594
R8956 gnd.n1931 gnd.n1854 99.6594
R8957 gnd.n1930 gnd.n1929 99.6594
R8958 gnd.n1912 gnd.n1863 99.6594
R8959 gnd.n1911 gnd.n1910 99.6594
R8960 gnd.n1893 gnd.n1872 99.6594
R8961 gnd.n1892 gnd.n1611 99.6594
R8962 gnd.n2642 gnd.t163 98.63
R8963 gnd.n118 gnd.t100 98.63
R8964 gnd.n1839 gnd.t130 98.63
R8965 gnd.n2618 gnd.t145 98.63
R8966 gnd.n2137 gnd.t123 98.63
R8967 gnd.n2166 gnd.t105 98.63
R8968 gnd.n197 gnd.t176 98.63
R8969 gnd.n7629 gnd.t188 98.63
R8970 gnd.n1062 gnd.t120 98.63
R8971 gnd.n1084 gnd.t97 98.63
R8972 gnd.n2934 gnd.t156 98.63
R8973 gnd.n3264 gnd.t116 98.63
R8974 gnd.n1458 gnd.t142 98.63
R8975 gnd.n1983 gnd.t133 98.63
R8976 gnd.n3482 gnd.t180 88.9408
R8977 gnd.n2220 gnd.t92 88.9408
R8978 gnd.n4731 gnd.t113 88.933
R8979 gnd.n4021 gnd.t148 88.933
R8980 gnd.n1510 gnd.n1509 81.8399
R8981 gnd.n5714 gnd.t88 74.8376
R8982 gnd.n5137 gnd.t127 74.8376
R8983 gnd.n7364 gnd.n202 73.4358
R8984 gnd.n3483 gnd.t179 72.8438
R8985 gnd.n2221 gnd.t93 72.8438
R8986 gnd.n1511 gnd.n1504 72.8411
R8987 gnd.n1517 gnd.n1502 72.8411
R8988 gnd.n4017 gnd.n4016 72.8411
R8989 gnd.n2643 gnd.t162 72.836
R8990 gnd.n4732 gnd.t112 72.836
R8991 gnd.n4022 gnd.t149 72.836
R8992 gnd.n119 gnd.t101 72.836
R8993 gnd.n1840 gnd.t129 72.836
R8994 gnd.n2619 gnd.t146 72.836
R8995 gnd.n2138 gnd.t122 72.836
R8996 gnd.n2167 gnd.t104 72.836
R8997 gnd.n198 gnd.t177 72.836
R8998 gnd.n7630 gnd.t189 72.836
R8999 gnd.n1063 gnd.t119 72.836
R9000 gnd.n1085 gnd.t96 72.836
R9001 gnd.n2935 gnd.t155 72.836
R9002 gnd.n3265 gnd.t117 72.836
R9003 gnd.n1459 gnd.t143 72.836
R9004 gnd.n1984 gnd.t134 72.836
R9005 gnd.n4085 gnd.n2044 71.676
R9006 gnd.n4081 gnd.n2045 71.676
R9007 gnd.n4077 gnd.n2046 71.676
R9008 gnd.n4073 gnd.n2047 71.676
R9009 gnd.n4069 gnd.n2048 71.676
R9010 gnd.n4065 gnd.n2049 71.676
R9011 gnd.n4061 gnd.n2050 71.676
R9012 gnd.n4057 gnd.n2051 71.676
R9013 gnd.n4053 gnd.n2052 71.676
R9014 gnd.n4049 gnd.n2053 71.676
R9015 gnd.n4045 gnd.n2054 71.676
R9016 gnd.n4041 gnd.n2055 71.676
R9017 gnd.n4037 gnd.n2056 71.676
R9018 gnd.n4033 gnd.n2057 71.676
R9019 gnd.n4028 gnd.n2058 71.676
R9020 gnd.n4024 gnd.n2059 71.676
R9021 gnd.n4161 gnd.n2077 71.676
R9022 gnd.n4157 gnd.n2076 71.676
R9023 gnd.n4152 gnd.n2075 71.676
R9024 gnd.n4148 gnd.n2074 71.676
R9025 gnd.n4144 gnd.n2073 71.676
R9026 gnd.n4140 gnd.n2072 71.676
R9027 gnd.n4136 gnd.n2071 71.676
R9028 gnd.n4132 gnd.n2070 71.676
R9029 gnd.n4128 gnd.n2069 71.676
R9030 gnd.n4124 gnd.n2068 71.676
R9031 gnd.n4120 gnd.n2067 71.676
R9032 gnd.n4116 gnd.n2066 71.676
R9033 gnd.n4112 gnd.n2065 71.676
R9034 gnd.n4108 gnd.n2064 71.676
R9035 gnd.n4104 gnd.n2063 71.676
R9036 gnd.n4100 gnd.n2062 71.676
R9037 gnd.n4096 gnd.n2061 71.676
R9038 gnd.n4795 gnd.n4794 71.676
R9039 gnd.n4789 gnd.n1466 71.676
R9040 gnd.n4786 gnd.n1467 71.676
R9041 gnd.n4782 gnd.n1468 71.676
R9042 gnd.n4778 gnd.n1469 71.676
R9043 gnd.n4774 gnd.n1470 71.676
R9044 gnd.n4770 gnd.n1471 71.676
R9045 gnd.n4766 gnd.n1472 71.676
R9046 gnd.n4762 gnd.n1473 71.676
R9047 gnd.n4758 gnd.n1474 71.676
R9048 gnd.n4754 gnd.n1475 71.676
R9049 gnd.n4750 gnd.n1476 71.676
R9050 gnd.n4746 gnd.n1477 71.676
R9051 gnd.n4742 gnd.n1478 71.676
R9052 gnd.n4738 gnd.n1479 71.676
R9053 gnd.n4734 gnd.n1480 71.676
R9054 gnd.n1481 gnd.n1465 71.676
R9055 gnd.n3486 gnd.n1482 71.676
R9056 gnd.n3491 gnd.n1483 71.676
R9057 gnd.n3495 gnd.n1484 71.676
R9058 gnd.n3499 gnd.n1485 71.676
R9059 gnd.n3503 gnd.n1486 71.676
R9060 gnd.n3507 gnd.n1487 71.676
R9061 gnd.n3511 gnd.n1488 71.676
R9062 gnd.n3515 gnd.n1489 71.676
R9063 gnd.n3519 gnd.n1490 71.676
R9064 gnd.n3523 gnd.n1491 71.676
R9065 gnd.n3527 gnd.n1492 71.676
R9066 gnd.n3531 gnd.n1493 71.676
R9067 gnd.n3535 gnd.n1494 71.676
R9068 gnd.n3539 gnd.n1495 71.676
R9069 gnd.n3543 gnd.n1496 71.676
R9070 gnd.n4795 gnd.n1499 71.676
R9071 gnd.n4787 gnd.n1466 71.676
R9072 gnd.n4783 gnd.n1467 71.676
R9073 gnd.n4779 gnd.n1468 71.676
R9074 gnd.n4775 gnd.n1469 71.676
R9075 gnd.n4771 gnd.n1470 71.676
R9076 gnd.n4767 gnd.n1471 71.676
R9077 gnd.n4763 gnd.n1472 71.676
R9078 gnd.n4759 gnd.n1473 71.676
R9079 gnd.n4755 gnd.n1474 71.676
R9080 gnd.n4751 gnd.n1475 71.676
R9081 gnd.n4747 gnd.n1476 71.676
R9082 gnd.n4743 gnd.n1477 71.676
R9083 gnd.n4739 gnd.n1478 71.676
R9084 gnd.n4735 gnd.n1479 71.676
R9085 gnd.n4798 gnd.n4797 71.676
R9086 gnd.n3485 gnd.n1481 71.676
R9087 gnd.n3490 gnd.n1482 71.676
R9088 gnd.n3494 gnd.n1483 71.676
R9089 gnd.n3498 gnd.n1484 71.676
R9090 gnd.n3502 gnd.n1485 71.676
R9091 gnd.n3506 gnd.n1486 71.676
R9092 gnd.n3510 gnd.n1487 71.676
R9093 gnd.n3514 gnd.n1488 71.676
R9094 gnd.n3518 gnd.n1489 71.676
R9095 gnd.n3522 gnd.n1490 71.676
R9096 gnd.n3526 gnd.n1491 71.676
R9097 gnd.n3530 gnd.n1492 71.676
R9098 gnd.n3534 gnd.n1493 71.676
R9099 gnd.n3538 gnd.n1494 71.676
R9100 gnd.n3542 gnd.n1495 71.676
R9101 gnd.n3481 gnd.n1496 71.676
R9102 gnd.n4099 gnd.n2061 71.676
R9103 gnd.n4103 gnd.n2062 71.676
R9104 gnd.n4107 gnd.n2063 71.676
R9105 gnd.n4111 gnd.n2064 71.676
R9106 gnd.n4115 gnd.n2065 71.676
R9107 gnd.n4119 gnd.n2066 71.676
R9108 gnd.n4123 gnd.n2067 71.676
R9109 gnd.n4127 gnd.n2068 71.676
R9110 gnd.n4131 gnd.n2069 71.676
R9111 gnd.n4135 gnd.n2070 71.676
R9112 gnd.n4139 gnd.n2071 71.676
R9113 gnd.n4143 gnd.n2072 71.676
R9114 gnd.n4147 gnd.n2073 71.676
R9115 gnd.n4151 gnd.n2074 71.676
R9116 gnd.n4156 gnd.n2075 71.676
R9117 gnd.n4160 gnd.n2076 71.676
R9118 gnd.n4023 gnd.n2060 71.676
R9119 gnd.n4027 gnd.n2059 71.676
R9120 gnd.n4032 gnd.n2058 71.676
R9121 gnd.n4036 gnd.n2057 71.676
R9122 gnd.n4040 gnd.n2056 71.676
R9123 gnd.n4044 gnd.n2055 71.676
R9124 gnd.n4048 gnd.n2054 71.676
R9125 gnd.n4052 gnd.n2053 71.676
R9126 gnd.n4056 gnd.n2052 71.676
R9127 gnd.n4060 gnd.n2051 71.676
R9128 gnd.n4064 gnd.n2050 71.676
R9129 gnd.n4068 gnd.n2049 71.676
R9130 gnd.n4072 gnd.n2048 71.676
R9131 gnd.n4076 gnd.n2047 71.676
R9132 gnd.n4080 gnd.n2046 71.676
R9133 gnd.n4084 gnd.n2045 71.676
R9134 gnd.n4087 gnd.n2044 71.676
R9135 gnd.n8 gnd.t78 69.1507
R9136 gnd.n14 gnd.t20 68.4792
R9137 gnd.n13 gnd.t32 68.4792
R9138 gnd.n12 gnd.t69 68.4792
R9139 gnd.n11 gnd.t71 68.4792
R9140 gnd.n10 gnd.t38 68.4792
R9141 gnd.n9 gnd.t49 68.4792
R9142 gnd.n8 gnd.t67 68.4792
R9143 gnd.n5626 gnd.n5527 64.369
R9144 gnd.n3488 gnd.n3483 59.5399
R9145 gnd.n4154 gnd.n2221 59.5399
R9146 gnd.n4733 gnd.n4732 59.5399
R9147 gnd.n4030 gnd.n4022 59.5399
R9148 gnd.n4730 gnd.n1520 59.1804
R9149 gnd.n6512 gnd.n6511 57.3586
R9150 gnd.n5329 gnd.t199 56.607
R9151 gnd.n56 gnd.t321 56.607
R9152 gnd.n5290 gnd.t277 56.407
R9153 gnd.n5309 gnd.t250 56.407
R9154 gnd.n17 gnd.t317 56.407
R9155 gnd.n36 gnd.t288 56.407
R9156 gnd.n5346 gnd.t259 55.8337
R9157 gnd.n5307 gnd.t301 55.8337
R9158 gnd.n5326 gnd.t273 55.8337
R9159 gnd.n73 gnd.t332 55.8337
R9160 gnd.n34 gnd.t315 55.8337
R9161 gnd.n53 gnd.t284 55.8337
R9162 gnd.n1508 gnd.n1507 54.358
R9163 gnd.n4014 gnd.n4013 54.358
R9164 gnd.n5329 gnd.n5328 53.0052
R9165 gnd.n5331 gnd.n5330 53.0052
R9166 gnd.n5333 gnd.n5332 53.0052
R9167 gnd.n5335 gnd.n5334 53.0052
R9168 gnd.n5337 gnd.n5336 53.0052
R9169 gnd.n5339 gnd.n5338 53.0052
R9170 gnd.n5341 gnd.n5340 53.0052
R9171 gnd.n5343 gnd.n5342 53.0052
R9172 gnd.n5345 gnd.n5344 53.0052
R9173 gnd.n5290 gnd.n5289 53.0052
R9174 gnd.n5292 gnd.n5291 53.0052
R9175 gnd.n5294 gnd.n5293 53.0052
R9176 gnd.n5296 gnd.n5295 53.0052
R9177 gnd.n5298 gnd.n5297 53.0052
R9178 gnd.n5300 gnd.n5299 53.0052
R9179 gnd.n5302 gnd.n5301 53.0052
R9180 gnd.n5304 gnd.n5303 53.0052
R9181 gnd.n5306 gnd.n5305 53.0052
R9182 gnd.n5309 gnd.n5308 53.0052
R9183 gnd.n5311 gnd.n5310 53.0052
R9184 gnd.n5313 gnd.n5312 53.0052
R9185 gnd.n5315 gnd.n5314 53.0052
R9186 gnd.n5317 gnd.n5316 53.0052
R9187 gnd.n5319 gnd.n5318 53.0052
R9188 gnd.n5321 gnd.n5320 53.0052
R9189 gnd.n5323 gnd.n5322 53.0052
R9190 gnd.n5325 gnd.n5324 53.0052
R9191 gnd.n72 gnd.n71 53.0052
R9192 gnd.n70 gnd.n69 53.0052
R9193 gnd.n68 gnd.n67 53.0052
R9194 gnd.n66 gnd.n65 53.0052
R9195 gnd.n64 gnd.n63 53.0052
R9196 gnd.n62 gnd.n61 53.0052
R9197 gnd.n60 gnd.n59 53.0052
R9198 gnd.n58 gnd.n57 53.0052
R9199 gnd.n56 gnd.n55 53.0052
R9200 gnd.n33 gnd.n32 53.0052
R9201 gnd.n31 gnd.n30 53.0052
R9202 gnd.n29 gnd.n28 53.0052
R9203 gnd.n27 gnd.n26 53.0052
R9204 gnd.n25 gnd.n24 53.0052
R9205 gnd.n23 gnd.n22 53.0052
R9206 gnd.n21 gnd.n20 53.0052
R9207 gnd.n19 gnd.n18 53.0052
R9208 gnd.n17 gnd.n16 53.0052
R9209 gnd.n52 gnd.n51 53.0052
R9210 gnd.n50 gnd.n49 53.0052
R9211 gnd.n48 gnd.n47 53.0052
R9212 gnd.n46 gnd.n45 53.0052
R9213 gnd.n44 gnd.n43 53.0052
R9214 gnd.n42 gnd.n41 53.0052
R9215 gnd.n40 gnd.n39 53.0052
R9216 gnd.n38 gnd.n37 53.0052
R9217 gnd.n36 gnd.n35 53.0052
R9218 gnd.n4005 gnd.n4004 52.4801
R9219 gnd.n6374 gnd.t80 52.3082
R9220 gnd.n6342 gnd.t61 52.3082
R9221 gnd.n6310 gnd.t75 52.3082
R9222 gnd.n6279 gnd.t56 52.3082
R9223 gnd.n6247 gnd.t58 52.3082
R9224 gnd.n6215 gnd.t73 52.3082
R9225 gnd.n6183 gnd.t36 52.3082
R9226 gnd.n6152 gnd.t82 52.3082
R9227 gnd.n5107 gnd.n1040 51.6227
R9228 gnd.n7666 gnd.n124 51.6227
R9229 gnd.n6204 gnd.n6172 51.4173
R9230 gnd.n6268 gnd.n6267 50.455
R9231 gnd.n6236 gnd.n6235 50.455
R9232 gnd.n6204 gnd.n6203 50.455
R9233 gnd.n5564 gnd.n5563 45.1884
R9234 gnd.n5163 gnd.n5162 45.1884
R9235 gnd.n4089 gnd.n4020 44.3322
R9236 gnd.n1511 gnd.n1510 44.3189
R9237 gnd.n2644 gnd.n2643 42.2793
R9238 gnd.n5576 gnd.n5564 42.2793
R9239 gnd.n5164 gnd.n5163 42.2793
R9240 gnd.n5716 gnd.n5714 42.2793
R9241 gnd.n6483 gnd.n5137 42.2793
R9242 gnd.n120 gnd.n119 42.2793
R9243 gnd.n1841 gnd.n1840 42.2793
R9244 gnd.n3333 gnd.n2619 42.2793
R9245 gnd.n2168 gnd.n2167 42.2793
R9246 gnd.n7594 gnd.n198 42.2793
R9247 gnd.n7631 gnd.n7630 42.2793
R9248 gnd.n5071 gnd.n1063 42.2793
R9249 gnd.n1086 gnd.n1085 42.2793
R9250 gnd.n2936 gnd.n2935 42.2793
R9251 gnd.n3323 gnd.n3265 42.2793
R9252 gnd.n1985 gnd.n1984 42.2793
R9253 gnd.n1509 gnd.n1508 41.6274
R9254 gnd.n4015 gnd.n4014 41.6274
R9255 gnd.n1518 gnd.n1517 40.8975
R9256 gnd.n4018 gnd.n4017 40.8975
R9257 gnd.n2218 gnd.n2138 36.9518
R9258 gnd.n4800 gnd.n1459 36.9518
R9259 gnd.n6701 gnd.n796 36.1788
R9260 gnd.n6695 gnd.n796 36.1788
R9261 gnd.n6695 gnd.n6694 36.1788
R9262 gnd.n6694 gnd.n6693 36.1788
R9263 gnd.n6693 gnd.n803 36.1788
R9264 gnd.n6687 gnd.n803 36.1788
R9265 gnd.n6687 gnd.n6686 36.1788
R9266 gnd.n6686 gnd.n6685 36.1788
R9267 gnd.n6685 gnd.n811 36.1788
R9268 gnd.n6679 gnd.n811 36.1788
R9269 gnd.n6679 gnd.n6678 36.1788
R9270 gnd.n6678 gnd.n6677 36.1788
R9271 gnd.n6677 gnd.n819 36.1788
R9272 gnd.n6671 gnd.n819 36.1788
R9273 gnd.n6671 gnd.n6670 36.1788
R9274 gnd.n6670 gnd.n6669 36.1788
R9275 gnd.n6669 gnd.n827 36.1788
R9276 gnd.n6663 gnd.n827 36.1788
R9277 gnd.n6663 gnd.n6662 36.1788
R9278 gnd.n6662 gnd.n6661 36.1788
R9279 gnd.n6661 gnd.n835 36.1788
R9280 gnd.n6655 gnd.n835 36.1788
R9281 gnd.n6655 gnd.n6654 36.1788
R9282 gnd.n6654 gnd.n6653 36.1788
R9283 gnd.n6653 gnd.n843 36.1788
R9284 gnd.n6647 gnd.n843 36.1788
R9285 gnd.n6647 gnd.n6646 36.1788
R9286 gnd.n6646 gnd.n6645 36.1788
R9287 gnd.n6645 gnd.n851 36.1788
R9288 gnd.n6639 gnd.n851 36.1788
R9289 gnd.n6639 gnd.n6638 36.1788
R9290 gnd.n6638 gnd.n6637 36.1788
R9291 gnd.n6637 gnd.n859 36.1788
R9292 gnd.n6631 gnd.n859 36.1788
R9293 gnd.n6631 gnd.n6630 36.1788
R9294 gnd.n6630 gnd.n6629 36.1788
R9295 gnd.n6629 gnd.n867 36.1788
R9296 gnd.n6623 gnd.n867 36.1788
R9297 gnd.n6623 gnd.n6622 36.1788
R9298 gnd.n6622 gnd.n6621 36.1788
R9299 gnd.n6621 gnd.n875 36.1788
R9300 gnd.n6615 gnd.n875 36.1788
R9301 gnd.n6615 gnd.n6614 36.1788
R9302 gnd.n6614 gnd.n6613 36.1788
R9303 gnd.n6613 gnd.n883 36.1788
R9304 gnd.n6607 gnd.n883 36.1788
R9305 gnd.n6607 gnd.n6606 36.1788
R9306 gnd.n6606 gnd.n6605 36.1788
R9307 gnd.n6605 gnd.n891 36.1788
R9308 gnd.n6599 gnd.n891 36.1788
R9309 gnd.n6599 gnd.n6598 36.1788
R9310 gnd.n6598 gnd.n6597 36.1788
R9311 gnd.n6597 gnd.n899 36.1788
R9312 gnd.n6591 gnd.n899 36.1788
R9313 gnd.n6591 gnd.n6590 36.1788
R9314 gnd.n6590 gnd.n6589 36.1788
R9315 gnd.n6589 gnd.n907 36.1788
R9316 gnd.n6583 gnd.n907 36.1788
R9317 gnd.n6583 gnd.n6582 36.1788
R9318 gnd.n6582 gnd.n6581 36.1788
R9319 gnd.n6581 gnd.n915 36.1788
R9320 gnd.n6575 gnd.n915 36.1788
R9321 gnd.n6575 gnd.n6574 36.1788
R9322 gnd.n6574 gnd.n6573 36.1788
R9323 gnd.n6573 gnd.n923 36.1788
R9324 gnd.n6567 gnd.n923 36.1788
R9325 gnd.n6567 gnd.n6566 36.1788
R9326 gnd.n6566 gnd.n6565 36.1788
R9327 gnd.n6565 gnd.n931 36.1788
R9328 gnd.n6559 gnd.n931 36.1788
R9329 gnd.n6559 gnd.n6558 36.1788
R9330 gnd.n6558 gnd.n6557 36.1788
R9331 gnd.n6557 gnd.n939 36.1788
R9332 gnd.n6551 gnd.n939 36.1788
R9333 gnd.n6551 gnd.n6550 36.1788
R9334 gnd.n6550 gnd.n6549 36.1788
R9335 gnd.n6549 gnd.n947 36.1788
R9336 gnd.n6543 gnd.n947 36.1788
R9337 gnd.n6543 gnd.n6542 36.1788
R9338 gnd.n6542 gnd.n6541 36.1788
R9339 gnd.n6541 gnd.n955 36.1788
R9340 gnd.n6535 gnd.n955 36.1788
R9341 gnd.n6535 gnd.n6534 36.1788
R9342 gnd.n1517 gnd.n1516 35.055
R9343 gnd.n1512 gnd.n1511 35.055
R9344 gnd.n4007 gnd.n4006 35.055
R9345 gnd.n4017 gnd.n4003 35.055
R9346 gnd.n5626 gnd.n5522 31.8661
R9347 gnd.n5634 gnd.n5522 31.8661
R9348 gnd.n5642 gnd.n5516 31.8661
R9349 gnd.n5642 gnd.n5510 31.8661
R9350 gnd.n5650 gnd.n5510 31.8661
R9351 gnd.n5650 gnd.n5503 31.8661
R9352 gnd.n5658 gnd.n5503 31.8661
R9353 gnd.n5658 gnd.n5504 31.8661
R9354 gnd.n5757 gnd.n5489 31.8661
R9355 gnd.n2992 gnd.n1040 31.8661
R9356 gnd.n5020 gnd.n1094 31.8661
R9357 gnd.n5020 gnd.n1096 31.8661
R9358 gnd.n5014 gnd.n1096 31.8661
R9359 gnd.n5014 gnd.n1108 31.8661
R9360 gnd.n5008 gnd.n1119 31.8661
R9361 gnd.n5002 gnd.n1119 31.8661
R9362 gnd.n4996 gnd.n1136 31.8661
R9363 gnd.n4996 gnd.n1139 31.8661
R9364 gnd.n4990 gnd.n1149 31.8661
R9365 gnd.n4984 gnd.n1159 31.8661
R9366 gnd.n4978 gnd.n1159 31.8661
R9367 gnd.n4972 gnd.n1176 31.8661
R9368 gnd.n3215 gnd.n1423 31.8661
R9369 gnd.n3215 gnd.n2649 31.8661
R9370 gnd.n3228 gnd.n2673 31.8661
R9371 gnd.n4624 gnd.n1614 31.8661
R9372 gnd.n4618 gnd.n4617 31.8661
R9373 gnd.n4617 gnd.n4616 31.8661
R9374 gnd.n7454 gnd.n265 31.8661
R9375 gnd.n7462 gnd.n256 31.8661
R9376 gnd.n7462 gnd.n259 31.8661
R9377 gnd.n7470 gnd.n250 31.8661
R9378 gnd.n7478 gnd.n235 31.8661
R9379 gnd.n7486 gnd.n235 31.8661
R9380 gnd.n7494 gnd.n226 31.8661
R9381 gnd.n7494 gnd.n229 31.8661
R9382 gnd.n7502 gnd.n209 31.8661
R9383 gnd.n7578 gnd.n209 31.8661
R9384 gnd.n7578 gnd.n212 31.8661
R9385 gnd.n7666 gnd.n122 31.8661
R9386 gnd.n4966 gnd.n1190 31.2288
R9387 gnd.n4960 gnd.n1201 31.2288
R9388 gnd.n3049 gnd.n1209 31.2288
R9389 gnd.n3057 gnd.n1219 31.2288
R9390 gnd.n4948 gnd.n1222 31.2288
R9391 gnd.n4941 gnd.n1231 31.2288
R9392 gnd.n4935 gnd.n1242 31.2288
R9393 gnd.n3081 gnd.n1247 31.2288
R9394 gnd.n3089 gnd.n1256 31.2288
R9395 gnd.n4922 gnd.n1259 31.2288
R9396 gnd.n3097 gnd.n1264 31.2288
R9397 gnd.n4915 gnd.n1267 31.2288
R9398 gnd.n4909 gnd.n1278 31.2288
R9399 gnd.n3113 gnd.n1286 31.2288
R9400 gnd.n3121 gnd.n1296 31.2288
R9401 gnd.n3129 gnd.n1306 31.2288
R9402 gnd.n4891 gnd.n1309 31.2288
R9403 gnd.n4885 gnd.n1320 31.2288
R9404 gnd.n3145 gnd.n1328 31.2288
R9405 gnd.n3153 gnd.n1338 31.2288
R9406 gnd.n3161 gnd.n1348 31.2288
R9407 gnd.n4867 gnd.n1351 31.2288
R9408 gnd.n4861 gnd.n1362 31.2288
R9409 gnd.n3178 gnd.n1370 31.2288
R9410 gnd.n3196 gnd.n1380 31.2288
R9411 gnd.n4849 gnd.n1383 31.2288
R9412 gnd.n3188 gnd.n1391 31.2288
R9413 gnd.n4843 gnd.n1394 31.2288
R9414 gnd.n4837 gnd.n1405 31.2288
R9415 gnd.n3329 gnd.n1412 31.2288
R9416 gnd.n1633 gnd.n1632 31.2288
R9417 gnd.n4610 gnd.n4609 31.2288
R9418 gnd.n4603 gnd.n1646 31.2288
R9419 gnd.n4337 gnd.n1649 31.2288
R9420 gnd.n4336 gnd.n1825 31.2288
R9421 gnd.n4348 gnd.n4347 31.2288
R9422 gnd.n4358 gnd.n1807 31.2288
R9423 gnd.n4369 gnd.n1795 31.2288
R9424 gnd.n4379 gnd.n4378 31.2288
R9425 gnd.n4391 gnd.n1778 31.2288
R9426 gnd.n4401 gnd.n1769 31.2288
R9427 gnd.n4412 gnd.n4411 31.2288
R9428 gnd.n4423 gnd.n1752 31.2288
R9429 gnd.n4433 gnd.n1743 31.2288
R9430 gnd.n1745 gnd.n1735 31.2288
R9431 gnd.n4477 gnd.n1725 31.2288
R9432 gnd.n4487 gnd.n1716 31.2288
R9433 gnd.n4468 gnd.n1718 31.2288
R9434 gnd.n4562 gnd.n1683 31.2288
R9435 gnd.n4495 gnd.n1686 31.2288
R9436 gnd.n7413 gnd.n310 31.2288
R9437 gnd.n4531 gnd.n313 31.2288
R9438 gnd.n4542 gnd.n1699 31.2288
R9439 gnd.n4541 gnd.n1704 31.2288
R9440 gnd.n7394 gnd.n332 31.2288
R9441 gnd.n4515 gnd.n328 31.2288
R9442 gnd.n7422 gnd.n296 31.2288
R9443 gnd.n7430 gnd.n287 31.2288
R9444 gnd.n7379 gnd.n290 31.2288
R9445 gnd.n7373 gnd.n281 31.2288
R9446 gnd.n4097 gnd.n2222 31.0639
R9447 gnd.n3547 gnd.n3545 31.0639
R9448 gnd.t248 gnd.n1228 30.9101
R9449 gnd.n4897 gnd.t204 30.9101
R9450 gnd.t242 gnd.n4448 30.9101
R9451 gnd.n7393 gnd.t313 30.9101
R9452 gnd.n4990 gnd.t229 30.2728
R9453 gnd.t281 gnd.n1187 30.2728
R9454 gnd.n4873 gnd.t217 30.2728
R9455 gnd.n4321 gnd.t306 30.2728
R9456 gnd.n7372 gnd.t240 30.2728
R9457 gnd.n250 gnd.t192 30.2728
R9458 gnd.n2992 gnd.t95 28.3609
R9459 gnd.t99 gnd.n122 28.3609
R9460 gnd.t115 gnd.n1402 27.7236
R9461 gnd.t103 gnd.n1636 27.7236
R9462 gnd.n7586 gnd.n202 26.1303
R9463 gnd.n2643 gnd.n2642 25.7944
R9464 gnd.n5714 gnd.n5713 25.7944
R9465 gnd.n5137 gnd.n5136 25.7944
R9466 gnd.n119 gnd.n118 25.7944
R9467 gnd.n1840 gnd.n1839 25.7944
R9468 gnd.n2619 gnd.n2618 25.7944
R9469 gnd.n2138 gnd.n2137 25.7944
R9470 gnd.n2167 gnd.n2166 25.7944
R9471 gnd.n198 gnd.n197 25.7944
R9472 gnd.n7630 gnd.n7629 25.7944
R9473 gnd.n1063 gnd.n1062 25.7944
R9474 gnd.n1085 gnd.n1084 25.7944
R9475 gnd.n2935 gnd.n2934 25.7944
R9476 gnd.n3265 gnd.n3264 25.7944
R9477 gnd.n1459 gnd.n1458 25.7944
R9478 gnd.n1984 gnd.n1983 25.7944
R9479 gnd.n5758 gnd.n5478 24.8557
R9480 gnd.n5481 gnd.n5472 24.8557
R9481 gnd.n5779 gnd.n5457 24.8557
R9482 gnd.n5798 gnd.n5797 24.8557
R9483 gnd.n5808 gnd.n5450 24.8557
R9484 gnd.n5821 gnd.n5438 24.8557
R9485 gnd.n5846 gnd.n5422 24.8557
R9486 gnd.n5845 gnd.n5424 24.8557
R9487 gnd.n5868 gnd.n5406 24.8557
R9488 gnd.n5857 gnd.n5398 24.8557
R9489 gnd.n5893 gnd.n5892 24.8557
R9490 gnd.n5903 gnd.n5391 24.8557
R9491 gnd.n5915 gnd.n5383 24.8557
R9492 gnd.n5914 gnd.n5371 24.8557
R9493 gnd.n5933 gnd.n5932 24.8557
R9494 gnd.n5954 gnd.n5352 24.8557
R9495 gnd.n5978 gnd.n5977 24.8557
R9496 gnd.n5989 gnd.n5275 24.8557
R9497 gnd.n5988 gnd.n5277 24.8557
R9498 gnd.n6000 gnd.n5268 24.8557
R9499 gnd.n6018 gnd.n6017 24.8557
R9500 gnd.n5259 gnd.n5248 24.8557
R9501 gnd.n6039 gnd.n5236 24.8557
R9502 gnd.n5239 gnd.n5237 24.8557
R9503 gnd.n6064 gnd.n6063 24.8557
R9504 gnd.n6075 gnd.n5221 24.8557
R9505 gnd.n6086 gnd.n5214 24.8557
R9506 gnd.n6085 gnd.n5202 24.8557
R9507 gnd.n5205 gnd.n5194 24.8557
R9508 gnd.n6123 gnd.n5184 24.8557
R9509 gnd.n5185 gnd.n963 24.8557
R9510 gnd.n6135 gnd.n973 24.8557
R9511 gnd.n6526 gnd.n6525 24.8557
R9512 gnd.n6418 gnd.n976 24.8557
R9513 gnd.n6411 gnd.n996 24.8557
R9514 gnd.n5776 gnd.t81 23.2624
R9515 gnd.t258 gnd.n1108 23.2624
R9516 gnd.n7502 gnd.t283 23.2624
R9517 gnd.n5768 gnd.t87 22.6251
R9518 gnd.t233 gnd.n1149 22.6251
R9519 gnd.n3197 gnd.t198 22.6251
R9520 gnd.n4346 gnd.t287 22.6251
R9521 gnd.n7470 gnd.t200 22.6251
R9522 gnd.n3041 gnd.t194 21.9878
R9523 gnd.n2706 gnd.t190 21.9878
R9524 gnd.n1771 gnd.t206 21.9878
R9525 gnd.n7438 gnd.t196 21.9878
R9526 gnd.n6534 gnd.n6533 21.7075
R9527 gnd.n5748 gnd.t55 21.3504
R9528 gnd.n3073 gnd.t211 21.3504
R9529 gnd.n2720 gnd.t213 21.3504
R9530 gnd.n4476 gnd.t227 21.3504
R9531 gnd.n4523 gnd.t302 21.3504
R9532 gnd.t7 gnd.n6102 20.7131
R9533 gnd.n2733 gnd.t231 20.7131
R9534 gnd.n3105 gnd.t251 20.7131
R9535 gnd.n4559 gnd.t289 20.7131
R9536 gnd.n4532 gnd.t221 20.7131
R9537 gnd.n4829 gnd.n1412 20.3945
R9538 gnd.n1632 gnd.n1624 20.3945
R9539 gnd.t9 gnd.n5249 20.0758
R9540 gnd.n1176 gnd.t262 20.0758
R9541 gnd.n2857 gnd.t245 20.0758
R9542 gnd.n3137 gnd.t238 20.0758
R9543 gnd.n4313 gnd.t270 20.0758
R9544 gnd.t260 gnd.n298 20.0758
R9545 gnd.n7454 gnd.t295 20.0758
R9546 gnd.n1505 gnd.t169 19.8005
R9547 gnd.n1505 gnd.t85 19.8005
R9548 gnd.n1506 gnd.t140 19.8005
R9549 gnd.n1506 gnd.t174 19.8005
R9550 gnd.n4011 gnd.t183 19.8005
R9551 gnd.n4011 gnd.t159 19.8005
R9552 gnd.n4012 gnd.t172 19.8005
R9553 gnd.n4012 gnd.t137 19.8005
R9554 gnd.n1502 gnd.n1501 19.5087
R9555 gnd.n1515 gnd.n1502 19.5087
R9556 gnd.n1513 gnd.n1504 19.5087
R9557 gnd.n4016 gnd.n4010 19.5087
R9558 gnd.t11 gnd.n5284 19.4385
R9559 gnd.n1136 gnd.t209 19.4385
R9560 gnd.n3033 gnd.n1179 19.4385
R9561 gnd.n3170 gnd.t219 19.4385
R9562 gnd.t236 gnd.n1787 19.4385
R9563 gnd.n7446 gnd.n274 19.4385
R9564 gnd.n7486 gnd.t223 19.4385
R9565 gnd.n3385 gnd.n2560 19.3944
R9566 gnd.n3385 gnd.n2557 19.3944
R9567 gnd.n3390 gnd.n2557 19.3944
R9568 gnd.n3390 gnd.n2558 19.3944
R9569 gnd.n2558 gnd.n2535 19.3944
R9570 gnd.n3415 gnd.n2535 19.3944
R9571 gnd.n3415 gnd.n2532 19.3944
R9572 gnd.n3420 gnd.n2532 19.3944
R9573 gnd.n3420 gnd.n2533 19.3944
R9574 gnd.n2533 gnd.n2511 19.3944
R9575 gnd.n3450 gnd.n2511 19.3944
R9576 gnd.n3450 gnd.n2508 19.3944
R9577 gnd.n3457 gnd.n2508 19.3944
R9578 gnd.n3457 gnd.n2509 19.3944
R9579 gnd.n3453 gnd.n2509 19.3944
R9580 gnd.n3453 gnd.n2487 19.3944
R9581 gnd.n3552 gnd.n2487 19.3944
R9582 gnd.n3552 gnd.n2484 19.3944
R9583 gnd.n3557 gnd.n2484 19.3944
R9584 gnd.n3557 gnd.n2485 19.3944
R9585 gnd.n2485 gnd.n2464 19.3944
R9586 gnd.n3612 gnd.n2464 19.3944
R9587 gnd.n3612 gnd.n2462 19.3944
R9588 gnd.n3616 gnd.n2462 19.3944
R9589 gnd.n3616 gnd.n2443 19.3944
R9590 gnd.n3641 gnd.n2443 19.3944
R9591 gnd.n3641 gnd.n2440 19.3944
R9592 gnd.n3649 gnd.n2440 19.3944
R9593 gnd.n3649 gnd.n2441 19.3944
R9594 gnd.n3645 gnd.n2441 19.3944
R9595 gnd.n3645 gnd.n2408 19.3944
R9596 gnd.n3701 gnd.n2408 19.3944
R9597 gnd.n3701 gnd.n2405 19.3944
R9598 gnd.n3706 gnd.n2405 19.3944
R9599 gnd.n3706 gnd.n2406 19.3944
R9600 gnd.n2406 gnd.n2383 19.3944
R9601 gnd.n3755 gnd.n2383 19.3944
R9602 gnd.n3755 gnd.n2380 19.3944
R9603 gnd.n3771 gnd.n2380 19.3944
R9604 gnd.n3771 gnd.n2381 19.3944
R9605 gnd.n3767 gnd.n2381 19.3944
R9606 gnd.n3767 gnd.n3766 19.3944
R9607 gnd.n3766 gnd.n3765 19.3944
R9608 gnd.n3765 gnd.n3762 19.3944
R9609 gnd.n3762 gnd.n2337 19.3944
R9610 gnd.n3855 gnd.n2337 19.3944
R9611 gnd.n3855 gnd.n2334 19.3944
R9612 gnd.n3860 gnd.n2334 19.3944
R9613 gnd.n3860 gnd.n2335 19.3944
R9614 gnd.n2335 gnd.n2315 19.3944
R9615 gnd.n3884 gnd.n2315 19.3944
R9616 gnd.n3884 gnd.n2313 19.3944
R9617 gnd.n3888 gnd.n2313 19.3944
R9618 gnd.n3888 gnd.n2271 19.3944
R9619 gnd.n3928 gnd.n2271 19.3944
R9620 gnd.n3928 gnd.n2268 19.3944
R9621 gnd.n3948 gnd.n2268 19.3944
R9622 gnd.n3948 gnd.n2269 19.3944
R9623 gnd.n3944 gnd.n2269 19.3944
R9624 gnd.n3944 gnd.n3943 19.3944
R9625 gnd.n3943 gnd.n3942 19.3944
R9626 gnd.n3942 gnd.n3937 19.3944
R9627 gnd.n3938 gnd.n3937 19.3944
R9628 gnd.n3938 gnd.n2041 19.3944
R9629 gnd.n4167 gnd.n2041 19.3944
R9630 gnd.n4167 gnd.n2039 19.3944
R9631 gnd.n4171 gnd.n2039 19.3944
R9632 gnd.n4171 gnd.n2030 19.3944
R9633 gnd.n4188 gnd.n2030 19.3944
R9634 gnd.n4188 gnd.n2028 19.3944
R9635 gnd.n4192 gnd.n2028 19.3944
R9636 gnd.n4192 gnd.n2018 19.3944
R9637 gnd.n4209 gnd.n2018 19.3944
R9638 gnd.n4209 gnd.n2016 19.3944
R9639 gnd.n4213 gnd.n2016 19.3944
R9640 gnd.n4213 gnd.n2006 19.3944
R9641 gnd.n4230 gnd.n2006 19.3944
R9642 gnd.n4230 gnd.n2004 19.3944
R9643 gnd.n4235 gnd.n2004 19.3944
R9644 gnd.n4235 gnd.n1995 19.3944
R9645 gnd.n4253 gnd.n1995 19.3944
R9646 gnd.n4254 gnd.n4253 19.3944
R9647 gnd.n3239 gnd.n3238 19.3944
R9648 gnd.n3238 gnd.n3237 19.3944
R9649 gnd.n3237 gnd.n3234 19.3944
R9650 gnd.n3370 gnd.n2576 19.3944
R9651 gnd.n3370 gnd.n3369 19.3944
R9652 gnd.n3369 gnd.n2579 19.3944
R9653 gnd.n3362 gnd.n2579 19.3944
R9654 gnd.n3362 gnd.n3361 19.3944
R9655 gnd.n3361 gnd.n2587 19.3944
R9656 gnd.n3354 gnd.n2587 19.3944
R9657 gnd.n3354 gnd.n3353 19.3944
R9658 gnd.n3353 gnd.n2597 19.3944
R9659 gnd.n3346 gnd.n2597 19.3944
R9660 gnd.n3346 gnd.n3345 19.3944
R9661 gnd.n3345 gnd.n2605 19.3944
R9662 gnd.n3338 gnd.n2605 19.3944
R9663 gnd.n3338 gnd.n3337 19.3944
R9664 gnd.n3337 gnd.n2615 19.3944
R9665 gnd.n2663 gnd.n2615 19.3944
R9666 gnd.n2663 gnd.n2633 19.3944
R9667 gnd.n3250 gnd.n2633 19.3944
R9668 gnd.n3250 gnd.n3249 19.3944
R9669 gnd.n3249 gnd.n3248 19.3944
R9670 gnd.n3248 gnd.n2637 19.3944
R9671 gnd.n3244 gnd.n2637 19.3944
R9672 gnd.n3244 gnd.n3243 19.3944
R9673 gnd.n3243 gnd.n3242 19.3944
R9674 gnd.n5621 gnd.n5620 19.3944
R9675 gnd.n5620 gnd.n5530 19.3944
R9676 gnd.n5615 gnd.n5530 19.3944
R9677 gnd.n5615 gnd.n5614 19.3944
R9678 gnd.n5614 gnd.n5535 19.3944
R9679 gnd.n5609 gnd.n5535 19.3944
R9680 gnd.n5609 gnd.n5608 19.3944
R9681 gnd.n5608 gnd.n5607 19.3944
R9682 gnd.n5607 gnd.n5541 19.3944
R9683 gnd.n5601 gnd.n5541 19.3944
R9684 gnd.n5601 gnd.n5600 19.3944
R9685 gnd.n5600 gnd.n5599 19.3944
R9686 gnd.n5599 gnd.n5547 19.3944
R9687 gnd.n5593 gnd.n5547 19.3944
R9688 gnd.n5593 gnd.n5592 19.3944
R9689 gnd.n5592 gnd.n5591 19.3944
R9690 gnd.n5591 gnd.n5553 19.3944
R9691 gnd.n5585 gnd.n5553 19.3944
R9692 gnd.n5585 gnd.n5584 19.3944
R9693 gnd.n5584 gnd.n5583 19.3944
R9694 gnd.n5583 gnd.n5559 19.3944
R9695 gnd.n5577 gnd.n5559 19.3944
R9696 gnd.n5575 gnd.n5574 19.3944
R9697 gnd.n5574 gnd.n5569 19.3944
R9698 gnd.n5569 gnd.n5567 19.3944
R9699 gnd.n6433 gnd.n6432 19.3944
R9700 gnd.n6432 gnd.n6429 19.3944
R9701 gnd.n6429 gnd.n6428 19.3944
R9702 gnd.n6478 gnd.n6477 19.3944
R9703 gnd.n6477 gnd.n6476 19.3944
R9704 gnd.n6476 gnd.n6473 19.3944
R9705 gnd.n6473 gnd.n6472 19.3944
R9706 gnd.n6472 gnd.n6469 19.3944
R9707 gnd.n6469 gnd.n6468 19.3944
R9708 gnd.n6468 gnd.n6465 19.3944
R9709 gnd.n6465 gnd.n6464 19.3944
R9710 gnd.n6464 gnd.n6461 19.3944
R9711 gnd.n6461 gnd.n6460 19.3944
R9712 gnd.n6460 gnd.n6457 19.3944
R9713 gnd.n6457 gnd.n6456 19.3944
R9714 gnd.n6456 gnd.n6453 19.3944
R9715 gnd.n6453 gnd.n6452 19.3944
R9716 gnd.n6452 gnd.n6449 19.3944
R9717 gnd.n6449 gnd.n6448 19.3944
R9718 gnd.n6448 gnd.n6445 19.3944
R9719 gnd.n6445 gnd.n6444 19.3944
R9720 gnd.n6444 gnd.n6441 19.3944
R9721 gnd.n6441 gnd.n6440 19.3944
R9722 gnd.n6440 gnd.n6437 19.3944
R9723 gnd.n6437 gnd.n6436 19.3944
R9724 gnd.n5761 gnd.n5760 19.3944
R9725 gnd.n5762 gnd.n5761 19.3944
R9726 gnd.n5762 gnd.n5471 19.3944
R9727 gnd.n5471 gnd.n5465 19.3944
R9728 gnd.n5787 gnd.n5465 19.3944
R9729 gnd.n5788 gnd.n5787 19.3944
R9730 gnd.n5788 gnd.n5448 19.3944
R9731 gnd.n5448 gnd.n5446 19.3944
R9732 gnd.n5812 gnd.n5446 19.3944
R9733 gnd.n5815 gnd.n5812 19.3944
R9734 gnd.n5815 gnd.n5814 19.3944
R9735 gnd.n5814 gnd.n5418 19.3944
R9736 gnd.n5853 gnd.n5418 19.3944
R9737 gnd.n5853 gnd.n5416 19.3944
R9738 gnd.n5859 gnd.n5416 19.3944
R9739 gnd.n5860 gnd.n5859 19.3944
R9740 gnd.n5860 gnd.n5386 19.3944
R9741 gnd.n5910 gnd.n5386 19.3944
R9742 gnd.n5911 gnd.n5910 19.3944
R9743 gnd.n5911 gnd.n5379 19.3944
R9744 gnd.n5922 gnd.n5379 19.3944
R9745 gnd.n5923 gnd.n5922 19.3944
R9746 gnd.n5923 gnd.n5362 19.3944
R9747 gnd.n5362 gnd.n5360 19.3944
R9748 gnd.n5947 gnd.n5360 19.3944
R9749 gnd.n5948 gnd.n5947 19.3944
R9750 gnd.n5948 gnd.n5271 19.3944
R9751 gnd.n5995 gnd.n5271 19.3944
R9752 gnd.n5996 gnd.n5995 19.3944
R9753 gnd.n5996 gnd.n5264 19.3944
R9754 gnd.n6007 gnd.n5264 19.3944
R9755 gnd.n6008 gnd.n6007 19.3944
R9756 gnd.n6008 gnd.n5247 19.3944
R9757 gnd.n5247 gnd.n5245 19.3944
R9758 gnd.n6032 gnd.n5245 19.3944
R9759 gnd.n6033 gnd.n6032 19.3944
R9760 gnd.n6033 gnd.n5217 19.3944
R9761 gnd.n6081 gnd.n5217 19.3944
R9762 gnd.n6082 gnd.n6081 19.3944
R9763 gnd.n6082 gnd.n5210 19.3944
R9764 gnd.n6093 gnd.n5210 19.3944
R9765 gnd.n6094 gnd.n6093 19.3944
R9766 gnd.n6094 gnd.n5193 19.3944
R9767 gnd.n5193 gnd.n5190 19.3944
R9768 gnd.n6118 gnd.n5190 19.3944
R9769 gnd.n6118 gnd.n5191 19.3944
R9770 gnd.n5191 gnd.n5174 19.3944
R9771 gnd.n6399 gnd.n5174 19.3944
R9772 gnd.n6401 gnd.n6399 19.3944
R9773 gnd.n6415 gnd.n6401 19.3944
R9774 gnd.n6415 gnd.n6414 19.3944
R9775 gnd.n6414 gnd.n6413 19.3944
R9776 gnd.n6413 gnd.n6409 19.3944
R9777 gnd.n5744 gnd.n5743 19.3944
R9778 gnd.n5743 gnd.n5742 19.3944
R9779 gnd.n5742 gnd.n5741 19.3944
R9780 gnd.n5741 gnd.n5739 19.3944
R9781 gnd.n5739 gnd.n5736 19.3944
R9782 gnd.n5736 gnd.n5735 19.3944
R9783 gnd.n5735 gnd.n5732 19.3944
R9784 gnd.n5732 gnd.n5731 19.3944
R9785 gnd.n5731 gnd.n5728 19.3944
R9786 gnd.n5728 gnd.n5727 19.3944
R9787 gnd.n5727 gnd.n5724 19.3944
R9788 gnd.n5724 gnd.n5723 19.3944
R9789 gnd.n5723 gnd.n5720 19.3944
R9790 gnd.n5720 gnd.n5719 19.3944
R9791 gnd.n5770 gnd.n5476 19.3944
R9792 gnd.n5770 gnd.n5474 19.3944
R9793 gnd.n5774 gnd.n5474 19.3944
R9794 gnd.n5774 gnd.n5455 19.3944
R9795 gnd.n5800 gnd.n5455 19.3944
R9796 gnd.n5800 gnd.n5453 19.3944
R9797 gnd.n5806 gnd.n5453 19.3944
R9798 gnd.n5806 gnd.n5805 19.3944
R9799 gnd.n5805 gnd.n5429 19.3944
R9800 gnd.n5834 gnd.n5429 19.3944
R9801 gnd.n5834 gnd.n5427 19.3944
R9802 gnd.n5843 gnd.n5427 19.3944
R9803 gnd.n5843 gnd.n5842 19.3944
R9804 gnd.n5842 gnd.n5841 19.3944
R9805 gnd.n5841 gnd.n5396 19.3944
R9806 gnd.n5895 gnd.n5396 19.3944
R9807 gnd.n5895 gnd.n5394 19.3944
R9808 gnd.n5901 gnd.n5394 19.3944
R9809 gnd.n5901 gnd.n5900 19.3944
R9810 gnd.n5900 gnd.n5369 19.3944
R9811 gnd.n5935 gnd.n5369 19.3944
R9812 gnd.n5935 gnd.n5367 19.3944
R9813 gnd.n5941 gnd.n5367 19.3944
R9814 gnd.n5941 gnd.n5940 19.3944
R9815 gnd.n5940 gnd.n5282 19.3944
R9816 gnd.n5980 gnd.n5282 19.3944
R9817 gnd.n5980 gnd.n5280 19.3944
R9818 gnd.n5986 gnd.n5280 19.3944
R9819 gnd.n5986 gnd.n5985 19.3944
R9820 gnd.n5985 gnd.n5254 19.3944
R9821 gnd.n6020 gnd.n5254 19.3944
R9822 gnd.n6020 gnd.n5252 19.3944
R9823 gnd.n6026 gnd.n5252 19.3944
R9824 gnd.n6026 gnd.n6025 19.3944
R9825 gnd.n6025 gnd.n5227 19.3944
R9826 gnd.n6066 gnd.n5227 19.3944
R9827 gnd.n6066 gnd.n5225 19.3944
R9828 gnd.n6072 gnd.n5225 19.3944
R9829 gnd.n6072 gnd.n6071 19.3944
R9830 gnd.n6071 gnd.n5200 19.3944
R9831 gnd.n6105 gnd.n5200 19.3944
R9832 gnd.n6105 gnd.n5198 19.3944
R9833 gnd.n6112 gnd.n5198 19.3944
R9834 gnd.n6112 gnd.n6111 19.3944
R9835 gnd.n6111 gnd.n967 19.3944
R9836 gnd.n6530 gnd.n967 19.3944
R9837 gnd.n6530 gnd.n6529 19.3944
R9838 gnd.n6529 gnd.n6528 19.3944
R9839 gnd.n6528 gnd.n971 19.3944
R9840 gnd.n989 gnd.n971 19.3944
R9841 gnd.n6516 gnd.n989 19.3944
R9842 gnd.n6516 gnd.n6515 19.3944
R9843 gnd.n6515 gnd.n6514 19.3944
R9844 gnd.n5118 gnd.n5117 19.3944
R9845 gnd.n6508 gnd.n5117 19.3944
R9846 gnd.n6508 gnd.n6507 19.3944
R9847 gnd.n6507 gnd.n6506 19.3944
R9848 gnd.n6506 gnd.n6503 19.3944
R9849 gnd.n6503 gnd.n6502 19.3944
R9850 gnd.n6502 gnd.n6499 19.3944
R9851 gnd.n6499 gnd.n6498 19.3944
R9852 gnd.n6498 gnd.n6495 19.3944
R9853 gnd.n6495 gnd.n6494 19.3944
R9854 gnd.n6494 gnd.n6491 19.3944
R9855 gnd.n6491 gnd.n6490 19.3944
R9856 gnd.n6490 gnd.n6487 19.3944
R9857 gnd.n6487 gnd.n6486 19.3944
R9858 gnd.n5628 gnd.n5524 19.3944
R9859 gnd.n5632 gnd.n5524 19.3944
R9860 gnd.n5632 gnd.n5514 19.3944
R9861 gnd.n5644 gnd.n5514 19.3944
R9862 gnd.n5644 gnd.n5512 19.3944
R9863 gnd.n5648 gnd.n5512 19.3944
R9864 gnd.n5648 gnd.n5501 19.3944
R9865 gnd.n5660 gnd.n5501 19.3944
R9866 gnd.n5660 gnd.n5499 19.3944
R9867 gnd.n5686 gnd.n5499 19.3944
R9868 gnd.n5686 gnd.n5685 19.3944
R9869 gnd.n5685 gnd.n5684 19.3944
R9870 gnd.n5684 gnd.n5683 19.3944
R9871 gnd.n5683 gnd.n5681 19.3944
R9872 gnd.n5681 gnd.n5680 19.3944
R9873 gnd.n5680 gnd.n5678 19.3944
R9874 gnd.n5678 gnd.n5677 19.3944
R9875 gnd.n5677 gnd.n5675 19.3944
R9876 gnd.n5675 gnd.n5674 19.3944
R9877 gnd.n5674 gnd.n5436 19.3944
R9878 gnd.n5823 gnd.n5436 19.3944
R9879 gnd.n5823 gnd.n5434 19.3944
R9880 gnd.n5829 gnd.n5434 19.3944
R9881 gnd.n5829 gnd.n5828 19.3944
R9882 gnd.n5828 gnd.n5403 19.3944
R9883 gnd.n5870 gnd.n5403 19.3944
R9884 gnd.n5870 gnd.n5401 19.3944
R9885 gnd.n5874 gnd.n5401 19.3944
R9886 gnd.n5888 gnd.n5874 19.3944
R9887 gnd.n5886 gnd.n5885 19.3944
R9888 gnd.n5882 gnd.n5881 19.3944
R9889 gnd.n5878 gnd.n5877 19.3944
R9890 gnd.n5956 gnd.n5350 19.3944
R9891 gnd.n5956 gnd.n5288 19.3944
R9892 gnd.n5975 gnd.n5288 19.3944
R9893 gnd.n5975 gnd.n5974 19.3944
R9894 gnd.n5974 gnd.n5973 19.3944
R9895 gnd.n5973 gnd.n5971 19.3944
R9896 gnd.n5971 gnd.n5970 19.3944
R9897 gnd.n5970 gnd.n5968 19.3944
R9898 gnd.n5968 gnd.n5967 19.3944
R9899 gnd.n5967 gnd.n5234 19.3944
R9900 gnd.n6041 gnd.n5234 19.3944
R9901 gnd.n6041 gnd.n5232 19.3944
R9902 gnd.n6061 gnd.n5232 19.3944
R9903 gnd.n6061 gnd.n6060 19.3944
R9904 gnd.n6060 gnd.n6059 19.3944
R9905 gnd.n6059 gnd.n6056 19.3944
R9906 gnd.n6056 gnd.n6055 19.3944
R9907 gnd.n6055 gnd.n6053 19.3944
R9908 gnd.n6053 gnd.n6052 19.3944
R9909 gnd.n6052 gnd.n5182 19.3944
R9910 gnd.n6125 gnd.n5182 19.3944
R9911 gnd.n6125 gnd.n5180 19.3944
R9912 gnd.n6132 gnd.n5180 19.3944
R9913 gnd.n6132 gnd.n6131 19.3944
R9914 gnd.n6131 gnd.n5172 19.3944
R9915 gnd.n6420 gnd.n5172 19.3944
R9916 gnd.n6421 gnd.n6420 19.3944
R9917 gnd.n6421 gnd.n5170 19.3944
R9918 gnd.n6425 gnd.n5170 19.3944
R9919 gnd.n5624 gnd.n5520 19.3944
R9920 gnd.n5636 gnd.n5520 19.3944
R9921 gnd.n5636 gnd.n5518 19.3944
R9922 gnd.n5640 gnd.n5518 19.3944
R9923 gnd.n5640 gnd.n5508 19.3944
R9924 gnd.n5652 gnd.n5508 19.3944
R9925 gnd.n5652 gnd.n5506 19.3944
R9926 gnd.n5656 gnd.n5506 19.3944
R9927 gnd.n5656 gnd.n5495 19.3944
R9928 gnd.n5750 gnd.n5495 19.3944
R9929 gnd.n5750 gnd.n5492 19.3944
R9930 gnd.n5755 gnd.n5492 19.3944
R9931 gnd.n5755 gnd.n5483 19.3944
R9932 gnd.n5765 gnd.n5483 19.3944
R9933 gnd.n5765 gnd.n5467 19.3944
R9934 gnd.n5782 gnd.n5467 19.3944
R9935 gnd.n5782 gnd.n5463 19.3944
R9936 gnd.n5795 gnd.n5463 19.3944
R9937 gnd.n5795 gnd.n5794 19.3944
R9938 gnd.n5794 gnd.n5442 19.3944
R9939 gnd.n5819 gnd.n5442 19.3944
R9940 gnd.n5819 gnd.n5818 19.3944
R9941 gnd.n5818 gnd.n5420 19.3944
R9942 gnd.n5848 gnd.n5420 19.3944
R9943 gnd.n5848 gnd.n5410 19.3944
R9944 gnd.n5866 gnd.n5410 19.3944
R9945 gnd.n5866 gnd.n5865 19.3944
R9946 gnd.n5865 gnd.n5864 19.3944
R9947 gnd.n5864 gnd.n5388 19.3944
R9948 gnd.n5906 gnd.n5388 19.3944
R9949 gnd.n5906 gnd.n5381 19.3944
R9950 gnd.n5917 gnd.n5381 19.3944
R9951 gnd.n5917 gnd.n5377 19.3944
R9952 gnd.n5930 gnd.n5377 19.3944
R9953 gnd.n5930 gnd.n5929 19.3944
R9954 gnd.n5929 gnd.n5356 19.3944
R9955 gnd.n5952 gnd.n5356 19.3944
R9956 gnd.n5952 gnd.n5951 19.3944
R9957 gnd.n5951 gnd.n5273 19.3944
R9958 gnd.n5991 gnd.n5273 19.3944
R9959 gnd.n5991 gnd.n5266 19.3944
R9960 gnd.n6002 gnd.n5266 19.3944
R9961 gnd.n6002 gnd.n5262 19.3944
R9962 gnd.n6015 gnd.n5262 19.3944
R9963 gnd.n6015 gnd.n6014 19.3944
R9964 gnd.n6014 gnd.n5241 19.3944
R9965 gnd.n6037 gnd.n5241 19.3944
R9966 gnd.n6037 gnd.n6036 19.3944
R9967 gnd.n6036 gnd.n5219 19.3944
R9968 gnd.n6077 gnd.n5219 19.3944
R9969 gnd.n6077 gnd.n5212 19.3944
R9970 gnd.n6088 gnd.n5212 19.3944
R9971 gnd.n6088 gnd.n5208 19.3944
R9972 gnd.n6100 gnd.n5208 19.3944
R9973 gnd.n6100 gnd.n6099 19.3944
R9974 gnd.n6099 gnd.n5187 19.3944
R9975 gnd.n6121 gnd.n5187 19.3944
R9976 gnd.n6121 gnd.n5176 19.3944
R9977 gnd.n6138 gnd.n5176 19.3944
R9978 gnd.n6138 gnd.n979 19.3944
R9979 gnd.n6523 gnd.n979 19.3944
R9980 gnd.n6523 gnd.n6522 19.3944
R9981 gnd.n6522 gnd.n6521 19.3944
R9982 gnd.n6521 gnd.n983 19.3944
R9983 gnd.n6406 gnd.n983 19.3944
R9984 gnd.n4278 gnd.n1836 19.3944
R9985 gnd.n4282 gnd.n1836 19.3944
R9986 gnd.n4282 gnd.n1831 19.3944
R9987 gnd.n4339 gnd.n1831 19.3944
R9988 gnd.n4339 gnd.n1828 19.3944
R9989 gnd.n4344 gnd.n1828 19.3944
R9990 gnd.n4344 gnd.n1829 19.3944
R9991 gnd.n1829 gnd.n1793 19.3944
R9992 gnd.n4371 gnd.n1793 19.3944
R9993 gnd.n4371 gnd.n1790 19.3944
R9994 gnd.n4376 gnd.n1790 19.3944
R9995 gnd.n4376 gnd.n1791 19.3944
R9996 gnd.n1791 gnd.n1767 19.3944
R9997 gnd.n4403 gnd.n1767 19.3944
R9998 gnd.n4403 gnd.n1764 19.3944
R9999 gnd.n4408 gnd.n1764 19.3944
R10000 gnd.n4408 gnd.n1765 19.3944
R10001 gnd.n1765 gnd.n1741 19.3944
R10002 gnd.n4435 gnd.n1741 19.3944
R10003 gnd.n4435 gnd.n1738 19.3944
R10004 gnd.n4446 gnd.n1738 19.3944
R10005 gnd.n4446 gnd.n1739 19.3944
R10006 gnd.n4442 gnd.n1739 19.3944
R10007 gnd.n4442 gnd.n4441 19.3944
R10008 gnd.n4441 gnd.n1691 19.3944
R10009 gnd.n4557 gnd.n1691 19.3944
R10010 gnd.n4557 gnd.n1692 19.3944
R10011 gnd.n4553 gnd.n1692 19.3944
R10012 gnd.n4553 gnd.n4552 19.3944
R10013 gnd.n4552 gnd.n4551 19.3944
R10014 gnd.n4551 gnd.n4549 19.3944
R10015 gnd.n4549 gnd.n76 19.3944
R10016 gnd.n7717 gnd.n76 19.3944
R10017 gnd.n7717 gnd.n7716 19.3944
R10018 gnd.n7716 gnd.n7715 19.3944
R10019 gnd.n7715 gnd.n81 19.3944
R10020 gnd.n7711 gnd.n81 19.3944
R10021 gnd.n7711 gnd.n7710 19.3944
R10022 gnd.n7710 gnd.n7709 19.3944
R10023 gnd.n7709 gnd.n86 19.3944
R10024 gnd.n7705 gnd.n86 19.3944
R10025 gnd.n7705 gnd.n7704 19.3944
R10026 gnd.n7704 gnd.n7703 19.3944
R10027 gnd.n7703 gnd.n91 19.3944
R10028 gnd.n7699 gnd.n91 19.3944
R10029 gnd.n7699 gnd.n7698 19.3944
R10030 gnd.n7698 gnd.n7697 19.3944
R10031 gnd.n7697 gnd.n96 19.3944
R10032 gnd.n7693 gnd.n96 19.3944
R10033 gnd.n7693 gnd.n7692 19.3944
R10034 gnd.n7692 gnd.n7691 19.3944
R10035 gnd.n7691 gnd.n101 19.3944
R10036 gnd.n7687 gnd.n101 19.3944
R10037 gnd.n7687 gnd.n7686 19.3944
R10038 gnd.n7686 gnd.n7685 19.3944
R10039 gnd.n7685 gnd.n106 19.3944
R10040 gnd.n7681 gnd.n106 19.3944
R10041 gnd.n7681 gnd.n7680 19.3944
R10042 gnd.n7680 gnd.n7679 19.3944
R10043 gnd.n7679 gnd.n111 19.3944
R10044 gnd.n7675 gnd.n111 19.3944
R10045 gnd.n7675 gnd.n7674 19.3944
R10046 gnd.n7674 gnd.n7673 19.3944
R10047 gnd.n7673 gnd.n116 19.3944
R10048 gnd.n7567 gnd.n7566 19.3944
R10049 gnd.n7566 gnd.n7565 19.3944
R10050 gnd.n7565 gnd.n7514 19.3944
R10051 gnd.n7561 gnd.n7514 19.3944
R10052 gnd.n7561 gnd.n7560 19.3944
R10053 gnd.n7560 gnd.n7559 19.3944
R10054 gnd.n7559 gnd.n7522 19.3944
R10055 gnd.n7555 gnd.n7522 19.3944
R10056 gnd.n7555 gnd.n7554 19.3944
R10057 gnd.n7554 gnd.n7553 19.3944
R10058 gnd.n7553 gnd.n7530 19.3944
R10059 gnd.n7549 gnd.n7530 19.3944
R10060 gnd.n7549 gnd.n7548 19.3944
R10061 gnd.n7548 gnd.n7547 19.3944
R10062 gnd.n7547 gnd.n7538 19.3944
R10063 gnd.n7543 gnd.n7538 19.3944
R10064 gnd.n1878 gnd.n1877 19.3944
R10065 gnd.n1898 gnd.n1877 19.3944
R10066 gnd.n1898 gnd.n1875 19.3944
R10067 gnd.n1904 gnd.n1875 19.3944
R10068 gnd.n1904 gnd.n1868 19.3944
R10069 gnd.n1917 gnd.n1868 19.3944
R10070 gnd.n1917 gnd.n1866 19.3944
R10071 gnd.n1923 gnd.n1866 19.3944
R10072 gnd.n1923 gnd.n1859 19.3944
R10073 gnd.n1936 gnd.n1859 19.3944
R10074 gnd.n1936 gnd.n1857 19.3944
R10075 gnd.n1942 gnd.n1857 19.3944
R10076 gnd.n1942 gnd.n1850 19.3944
R10077 gnd.n1955 gnd.n1850 19.3944
R10078 gnd.n1955 gnd.n1848 19.3944
R10079 gnd.n1961 gnd.n1848 19.3944
R10080 gnd.n1884 gnd.n1883 19.3944
R10081 gnd.n1883 gnd.n1652 19.3944
R10082 gnd.n4601 gnd.n1652 19.3944
R10083 gnd.n4601 gnd.n1653 19.3944
R10084 gnd.n4597 gnd.n1653 19.3944
R10085 gnd.n4597 gnd.n4596 19.3944
R10086 gnd.n4596 gnd.n4595 19.3944
R10087 gnd.n4595 gnd.n1659 19.3944
R10088 gnd.n4591 gnd.n1659 19.3944
R10089 gnd.n4591 gnd.n4590 19.3944
R10090 gnd.n4590 gnd.n4589 19.3944
R10091 gnd.n4589 gnd.n1664 19.3944
R10092 gnd.n4585 gnd.n1664 19.3944
R10093 gnd.n4585 gnd.n4584 19.3944
R10094 gnd.n4584 gnd.n4583 19.3944
R10095 gnd.n4583 gnd.n1669 19.3944
R10096 gnd.n4579 gnd.n1669 19.3944
R10097 gnd.n4579 gnd.n4578 19.3944
R10098 gnd.n4578 gnd.n4577 19.3944
R10099 gnd.n4577 gnd.n1674 19.3944
R10100 gnd.n4573 gnd.n1674 19.3944
R10101 gnd.n4573 gnd.n4572 19.3944
R10102 gnd.n4572 gnd.n4571 19.3944
R10103 gnd.n4571 gnd.n1679 19.3944
R10104 gnd.n4567 gnd.n1679 19.3944
R10105 gnd.n4567 gnd.n4566 19.3944
R10106 gnd.n4566 gnd.n4565 19.3944
R10107 gnd.n4565 gnd.n316 19.3944
R10108 gnd.n7411 gnd.n316 19.3944
R10109 gnd.n7411 gnd.n317 19.3944
R10110 gnd.n7407 gnd.n317 19.3944
R10111 gnd.n7407 gnd.n7406 19.3944
R10112 gnd.n7406 gnd.n7405 19.3944
R10113 gnd.n7405 gnd.n323 19.3944
R10114 gnd.n7401 gnd.n323 19.3944
R10115 gnd.n7401 gnd.n7400 19.3944
R10116 gnd.n7400 gnd.n294 19.3944
R10117 gnd.n7424 gnd.n294 19.3944
R10118 gnd.n7424 gnd.n292 19.3944
R10119 gnd.n7428 gnd.n292 19.3944
R10120 gnd.n7428 gnd.n278 19.3944
R10121 gnd.n7440 gnd.n278 19.3944
R10122 gnd.n7440 gnd.n276 19.3944
R10123 gnd.n7444 gnd.n276 19.3944
R10124 gnd.n7444 gnd.n263 19.3944
R10125 gnd.n7456 gnd.n263 19.3944
R10126 gnd.n7456 gnd.n261 19.3944
R10127 gnd.n7460 gnd.n261 19.3944
R10128 gnd.n7460 gnd.n247 19.3944
R10129 gnd.n7472 gnd.n247 19.3944
R10130 gnd.n7472 gnd.n245 19.3944
R10131 gnd.n7476 gnd.n245 19.3944
R10132 gnd.n7476 gnd.n233 19.3944
R10133 gnd.n7488 gnd.n233 19.3944
R10134 gnd.n7488 gnd.n231 19.3944
R10135 gnd.n7492 gnd.n231 19.3944
R10136 gnd.n7492 gnd.n218 19.3944
R10137 gnd.n7504 gnd.n218 19.3944
R10138 gnd.n7504 gnd.n215 19.3944
R10139 gnd.n7576 gnd.n215 19.3944
R10140 gnd.n7576 gnd.n216 19.3944
R10141 gnd.n7572 gnd.n216 19.3944
R10142 gnd.n7572 gnd.n7571 19.3944
R10143 gnd.n7571 gnd.n7570 19.3944
R10144 gnd.n3375 gnd.n3374 19.3944
R10145 gnd.n3374 gnd.n3373 19.3944
R10146 gnd.n3373 gnd.n2573 19.3944
R10147 gnd.n3366 gnd.n2573 19.3944
R10148 gnd.n3366 gnd.n3365 19.3944
R10149 gnd.n3365 gnd.n2583 19.3944
R10150 gnd.n3358 gnd.n2583 19.3944
R10151 gnd.n3358 gnd.n3357 19.3944
R10152 gnd.n3357 gnd.n2593 19.3944
R10153 gnd.n3350 gnd.n2593 19.3944
R10154 gnd.n3350 gnd.n3349 19.3944
R10155 gnd.n3349 gnd.n2601 19.3944
R10156 gnd.n3342 gnd.n2601 19.3944
R10157 gnd.n3342 gnd.n3341 19.3944
R10158 gnd.n3341 gnd.n2611 19.3944
R10159 gnd.n3334 gnd.n2611 19.3944
R10160 gnd.n7159 gnd.n522 19.3944
R10161 gnd.n7159 gnd.n518 19.3944
R10162 gnd.n7165 gnd.n518 19.3944
R10163 gnd.n7165 gnd.n516 19.3944
R10164 gnd.n7169 gnd.n516 19.3944
R10165 gnd.n7169 gnd.n512 19.3944
R10166 gnd.n7175 gnd.n512 19.3944
R10167 gnd.n7175 gnd.n510 19.3944
R10168 gnd.n7179 gnd.n510 19.3944
R10169 gnd.n7179 gnd.n506 19.3944
R10170 gnd.n7185 gnd.n506 19.3944
R10171 gnd.n7185 gnd.n504 19.3944
R10172 gnd.n7189 gnd.n504 19.3944
R10173 gnd.n7189 gnd.n500 19.3944
R10174 gnd.n7195 gnd.n500 19.3944
R10175 gnd.n7195 gnd.n498 19.3944
R10176 gnd.n7199 gnd.n498 19.3944
R10177 gnd.n7199 gnd.n494 19.3944
R10178 gnd.n7205 gnd.n494 19.3944
R10179 gnd.n7205 gnd.n492 19.3944
R10180 gnd.n7209 gnd.n492 19.3944
R10181 gnd.n7209 gnd.n488 19.3944
R10182 gnd.n7215 gnd.n488 19.3944
R10183 gnd.n7215 gnd.n486 19.3944
R10184 gnd.n7219 gnd.n486 19.3944
R10185 gnd.n7219 gnd.n482 19.3944
R10186 gnd.n7225 gnd.n482 19.3944
R10187 gnd.n7225 gnd.n480 19.3944
R10188 gnd.n7229 gnd.n480 19.3944
R10189 gnd.n7229 gnd.n476 19.3944
R10190 gnd.n7235 gnd.n476 19.3944
R10191 gnd.n7235 gnd.n474 19.3944
R10192 gnd.n7239 gnd.n474 19.3944
R10193 gnd.n7239 gnd.n470 19.3944
R10194 gnd.n7245 gnd.n470 19.3944
R10195 gnd.n7245 gnd.n468 19.3944
R10196 gnd.n7249 gnd.n468 19.3944
R10197 gnd.n7249 gnd.n464 19.3944
R10198 gnd.n7255 gnd.n464 19.3944
R10199 gnd.n7255 gnd.n462 19.3944
R10200 gnd.n7259 gnd.n462 19.3944
R10201 gnd.n7259 gnd.n458 19.3944
R10202 gnd.n7265 gnd.n458 19.3944
R10203 gnd.n7265 gnd.n456 19.3944
R10204 gnd.n7269 gnd.n456 19.3944
R10205 gnd.n7269 gnd.n452 19.3944
R10206 gnd.n7275 gnd.n452 19.3944
R10207 gnd.n7275 gnd.n450 19.3944
R10208 gnd.n7279 gnd.n450 19.3944
R10209 gnd.n7279 gnd.n446 19.3944
R10210 gnd.n7285 gnd.n446 19.3944
R10211 gnd.n7285 gnd.n444 19.3944
R10212 gnd.n7289 gnd.n444 19.3944
R10213 gnd.n7289 gnd.n440 19.3944
R10214 gnd.n7295 gnd.n440 19.3944
R10215 gnd.n7295 gnd.n438 19.3944
R10216 gnd.n7299 gnd.n438 19.3944
R10217 gnd.n7299 gnd.n434 19.3944
R10218 gnd.n7305 gnd.n434 19.3944
R10219 gnd.n7305 gnd.n432 19.3944
R10220 gnd.n7309 gnd.n432 19.3944
R10221 gnd.n7309 gnd.n428 19.3944
R10222 gnd.n7315 gnd.n428 19.3944
R10223 gnd.n7315 gnd.n426 19.3944
R10224 gnd.n7319 gnd.n426 19.3944
R10225 gnd.n7319 gnd.n422 19.3944
R10226 gnd.n7325 gnd.n422 19.3944
R10227 gnd.n7325 gnd.n420 19.3944
R10228 gnd.n7329 gnd.n420 19.3944
R10229 gnd.n7329 gnd.n416 19.3944
R10230 gnd.n7335 gnd.n416 19.3944
R10231 gnd.n7335 gnd.n414 19.3944
R10232 gnd.n7339 gnd.n414 19.3944
R10233 gnd.n7339 gnd.n410 19.3944
R10234 gnd.n7345 gnd.n410 19.3944
R10235 gnd.n7345 gnd.n408 19.3944
R10236 gnd.n7349 gnd.n408 19.3944
R10237 gnd.n7349 gnd.n404 19.3944
R10238 gnd.n7355 gnd.n404 19.3944
R10239 gnd.n7355 gnd.n402 19.3944
R10240 gnd.n7360 gnd.n402 19.3944
R10241 gnd.n7360 gnd.n398 19.3944
R10242 gnd.n7366 gnd.n398 19.3944
R10243 gnd.n7367 gnd.n7366 19.3944
R10244 gnd.n6705 gnd.n794 19.3944
R10245 gnd.n6705 gnd.n792 19.3944
R10246 gnd.n6709 gnd.n792 19.3944
R10247 gnd.n6709 gnd.n788 19.3944
R10248 gnd.n6715 gnd.n788 19.3944
R10249 gnd.n6715 gnd.n786 19.3944
R10250 gnd.n6719 gnd.n786 19.3944
R10251 gnd.n6719 gnd.n782 19.3944
R10252 gnd.n6725 gnd.n782 19.3944
R10253 gnd.n6725 gnd.n780 19.3944
R10254 gnd.n6729 gnd.n780 19.3944
R10255 gnd.n6729 gnd.n776 19.3944
R10256 gnd.n6735 gnd.n776 19.3944
R10257 gnd.n6735 gnd.n774 19.3944
R10258 gnd.n6739 gnd.n774 19.3944
R10259 gnd.n6739 gnd.n770 19.3944
R10260 gnd.n6745 gnd.n770 19.3944
R10261 gnd.n6745 gnd.n768 19.3944
R10262 gnd.n6749 gnd.n768 19.3944
R10263 gnd.n6749 gnd.n764 19.3944
R10264 gnd.n6755 gnd.n764 19.3944
R10265 gnd.n6755 gnd.n762 19.3944
R10266 gnd.n6759 gnd.n762 19.3944
R10267 gnd.n6759 gnd.n758 19.3944
R10268 gnd.n6765 gnd.n758 19.3944
R10269 gnd.n6765 gnd.n756 19.3944
R10270 gnd.n6769 gnd.n756 19.3944
R10271 gnd.n6769 gnd.n752 19.3944
R10272 gnd.n6775 gnd.n752 19.3944
R10273 gnd.n6775 gnd.n750 19.3944
R10274 gnd.n6779 gnd.n750 19.3944
R10275 gnd.n6779 gnd.n746 19.3944
R10276 gnd.n6785 gnd.n746 19.3944
R10277 gnd.n6785 gnd.n744 19.3944
R10278 gnd.n6789 gnd.n744 19.3944
R10279 gnd.n6789 gnd.n740 19.3944
R10280 gnd.n6795 gnd.n740 19.3944
R10281 gnd.n6795 gnd.n738 19.3944
R10282 gnd.n6799 gnd.n738 19.3944
R10283 gnd.n6799 gnd.n734 19.3944
R10284 gnd.n6805 gnd.n734 19.3944
R10285 gnd.n6805 gnd.n732 19.3944
R10286 gnd.n6809 gnd.n732 19.3944
R10287 gnd.n6809 gnd.n728 19.3944
R10288 gnd.n6815 gnd.n728 19.3944
R10289 gnd.n6815 gnd.n726 19.3944
R10290 gnd.n6819 gnd.n726 19.3944
R10291 gnd.n6819 gnd.n722 19.3944
R10292 gnd.n6825 gnd.n722 19.3944
R10293 gnd.n6825 gnd.n720 19.3944
R10294 gnd.n6829 gnd.n720 19.3944
R10295 gnd.n6829 gnd.n716 19.3944
R10296 gnd.n6835 gnd.n716 19.3944
R10297 gnd.n6835 gnd.n714 19.3944
R10298 gnd.n6839 gnd.n714 19.3944
R10299 gnd.n6839 gnd.n710 19.3944
R10300 gnd.n6845 gnd.n710 19.3944
R10301 gnd.n6845 gnd.n708 19.3944
R10302 gnd.n6849 gnd.n708 19.3944
R10303 gnd.n6849 gnd.n704 19.3944
R10304 gnd.n6855 gnd.n704 19.3944
R10305 gnd.n6855 gnd.n702 19.3944
R10306 gnd.n6859 gnd.n702 19.3944
R10307 gnd.n6859 gnd.n698 19.3944
R10308 gnd.n6865 gnd.n698 19.3944
R10309 gnd.n6865 gnd.n696 19.3944
R10310 gnd.n6869 gnd.n696 19.3944
R10311 gnd.n6869 gnd.n692 19.3944
R10312 gnd.n6875 gnd.n692 19.3944
R10313 gnd.n6875 gnd.n690 19.3944
R10314 gnd.n6879 gnd.n690 19.3944
R10315 gnd.n6879 gnd.n686 19.3944
R10316 gnd.n6885 gnd.n686 19.3944
R10317 gnd.n6885 gnd.n684 19.3944
R10318 gnd.n6889 gnd.n684 19.3944
R10319 gnd.n6889 gnd.n680 19.3944
R10320 gnd.n6895 gnd.n680 19.3944
R10321 gnd.n6895 gnd.n678 19.3944
R10322 gnd.n6899 gnd.n678 19.3944
R10323 gnd.n6899 gnd.n674 19.3944
R10324 gnd.n6905 gnd.n674 19.3944
R10325 gnd.n6905 gnd.n672 19.3944
R10326 gnd.n6909 gnd.n672 19.3944
R10327 gnd.n6909 gnd.n668 19.3944
R10328 gnd.n6915 gnd.n668 19.3944
R10329 gnd.n6915 gnd.n666 19.3944
R10330 gnd.n6919 gnd.n666 19.3944
R10331 gnd.n6919 gnd.n662 19.3944
R10332 gnd.n6925 gnd.n662 19.3944
R10333 gnd.n6925 gnd.n660 19.3944
R10334 gnd.n6929 gnd.n660 19.3944
R10335 gnd.n6929 gnd.n656 19.3944
R10336 gnd.n6935 gnd.n656 19.3944
R10337 gnd.n6935 gnd.n654 19.3944
R10338 gnd.n6939 gnd.n654 19.3944
R10339 gnd.n6939 gnd.n650 19.3944
R10340 gnd.n6945 gnd.n650 19.3944
R10341 gnd.n6945 gnd.n648 19.3944
R10342 gnd.n6949 gnd.n648 19.3944
R10343 gnd.n6949 gnd.n644 19.3944
R10344 gnd.n6955 gnd.n644 19.3944
R10345 gnd.n6955 gnd.n642 19.3944
R10346 gnd.n6959 gnd.n642 19.3944
R10347 gnd.n6959 gnd.n638 19.3944
R10348 gnd.n6965 gnd.n638 19.3944
R10349 gnd.n6965 gnd.n636 19.3944
R10350 gnd.n6969 gnd.n636 19.3944
R10351 gnd.n6969 gnd.n632 19.3944
R10352 gnd.n6975 gnd.n632 19.3944
R10353 gnd.n6975 gnd.n630 19.3944
R10354 gnd.n6979 gnd.n630 19.3944
R10355 gnd.n6979 gnd.n626 19.3944
R10356 gnd.n6985 gnd.n626 19.3944
R10357 gnd.n6985 gnd.n624 19.3944
R10358 gnd.n6989 gnd.n624 19.3944
R10359 gnd.n6989 gnd.n620 19.3944
R10360 gnd.n6995 gnd.n620 19.3944
R10361 gnd.n6995 gnd.n618 19.3944
R10362 gnd.n6999 gnd.n618 19.3944
R10363 gnd.n6999 gnd.n614 19.3944
R10364 gnd.n7005 gnd.n614 19.3944
R10365 gnd.n7005 gnd.n612 19.3944
R10366 gnd.n7009 gnd.n612 19.3944
R10367 gnd.n7009 gnd.n608 19.3944
R10368 gnd.n7015 gnd.n608 19.3944
R10369 gnd.n7015 gnd.n606 19.3944
R10370 gnd.n7019 gnd.n606 19.3944
R10371 gnd.n7019 gnd.n602 19.3944
R10372 gnd.n7025 gnd.n602 19.3944
R10373 gnd.n7025 gnd.n600 19.3944
R10374 gnd.n7029 gnd.n600 19.3944
R10375 gnd.n7029 gnd.n596 19.3944
R10376 gnd.n7035 gnd.n596 19.3944
R10377 gnd.n7035 gnd.n594 19.3944
R10378 gnd.n7039 gnd.n594 19.3944
R10379 gnd.n7039 gnd.n590 19.3944
R10380 gnd.n7045 gnd.n590 19.3944
R10381 gnd.n7045 gnd.n588 19.3944
R10382 gnd.n7049 gnd.n588 19.3944
R10383 gnd.n7049 gnd.n584 19.3944
R10384 gnd.n7055 gnd.n584 19.3944
R10385 gnd.n7055 gnd.n582 19.3944
R10386 gnd.n7059 gnd.n582 19.3944
R10387 gnd.n7059 gnd.n578 19.3944
R10388 gnd.n7065 gnd.n578 19.3944
R10389 gnd.n7065 gnd.n576 19.3944
R10390 gnd.n7069 gnd.n576 19.3944
R10391 gnd.n7069 gnd.n572 19.3944
R10392 gnd.n7075 gnd.n572 19.3944
R10393 gnd.n7075 gnd.n570 19.3944
R10394 gnd.n7079 gnd.n570 19.3944
R10395 gnd.n7079 gnd.n566 19.3944
R10396 gnd.n7085 gnd.n566 19.3944
R10397 gnd.n7085 gnd.n564 19.3944
R10398 gnd.n7089 gnd.n564 19.3944
R10399 gnd.n7089 gnd.n560 19.3944
R10400 gnd.n7095 gnd.n560 19.3944
R10401 gnd.n7095 gnd.n558 19.3944
R10402 gnd.n7099 gnd.n558 19.3944
R10403 gnd.n7099 gnd.n554 19.3944
R10404 gnd.n7105 gnd.n554 19.3944
R10405 gnd.n7105 gnd.n552 19.3944
R10406 gnd.n7109 gnd.n552 19.3944
R10407 gnd.n7109 gnd.n548 19.3944
R10408 gnd.n7115 gnd.n548 19.3944
R10409 gnd.n7115 gnd.n546 19.3944
R10410 gnd.n7119 gnd.n546 19.3944
R10411 gnd.n7119 gnd.n542 19.3944
R10412 gnd.n7125 gnd.n542 19.3944
R10413 gnd.n7125 gnd.n540 19.3944
R10414 gnd.n7129 gnd.n540 19.3944
R10415 gnd.n7129 gnd.n536 19.3944
R10416 gnd.n7135 gnd.n536 19.3944
R10417 gnd.n7135 gnd.n534 19.3944
R10418 gnd.n7139 gnd.n534 19.3944
R10419 gnd.n7139 gnd.n530 19.3944
R10420 gnd.n7145 gnd.n530 19.3944
R10421 gnd.n7145 gnd.n528 19.3944
R10422 gnd.n7149 gnd.n528 19.3944
R10423 gnd.n7149 gnd.n524 19.3944
R10424 gnd.n7155 gnd.n524 19.3944
R10425 gnd.n2101 gnd.n2097 19.3944
R10426 gnd.n2101 gnd.n2094 19.3944
R10427 gnd.n2105 gnd.n2094 19.3944
R10428 gnd.n2105 gnd.n2092 19.3944
R10429 gnd.n2111 gnd.n2092 19.3944
R10430 gnd.n2111 gnd.n2090 19.3944
R10431 gnd.n2115 gnd.n2090 19.3944
R10432 gnd.n2115 gnd.n2088 19.3944
R10433 gnd.n2121 gnd.n2088 19.3944
R10434 gnd.n2121 gnd.n2086 19.3944
R10435 gnd.n2126 gnd.n2086 19.3944
R10436 gnd.n2126 gnd.n2084 19.3944
R10437 gnd.n2084 gnd.n2081 19.3944
R10438 gnd.n2133 gnd.n2081 19.3944
R10439 gnd.n2133 gnd.n2078 19.3944
R10440 gnd.n2217 gnd.n2140 19.3944
R10441 gnd.n2211 gnd.n2140 19.3944
R10442 gnd.n2211 gnd.n2210 19.3944
R10443 gnd.n2210 gnd.n2209 19.3944
R10444 gnd.n2209 gnd.n2146 19.3944
R10445 gnd.n2203 gnd.n2146 19.3944
R10446 gnd.n2203 gnd.n2202 19.3944
R10447 gnd.n2202 gnd.n2201 19.3944
R10448 gnd.n2201 gnd.n2152 19.3944
R10449 gnd.n2195 gnd.n2152 19.3944
R10450 gnd.n2195 gnd.n2194 19.3944
R10451 gnd.n2194 gnd.n2193 19.3944
R10452 gnd.n2193 gnd.n2158 19.3944
R10453 gnd.n2187 gnd.n2158 19.3944
R10454 gnd.n2187 gnd.n2186 19.3944
R10455 gnd.n2186 gnd.n2185 19.3944
R10456 gnd.n2185 gnd.n2164 19.3944
R10457 gnd.n2179 gnd.n2164 19.3944
R10458 gnd.n2171 gnd.n1835 19.3944
R10459 gnd.n4286 gnd.n1835 19.3944
R10460 gnd.n4286 gnd.n1833 19.3944
R10461 gnd.n4334 gnd.n1833 19.3944
R10462 gnd.n4334 gnd.n4333 19.3944
R10463 gnd.n4333 gnd.n4332 19.3944
R10464 gnd.n4332 gnd.n4331 19.3944
R10465 gnd.n4331 gnd.n4330 19.3944
R10466 gnd.n4330 gnd.n4328 19.3944
R10467 gnd.n4328 gnd.n4327 19.3944
R10468 gnd.n4327 gnd.n4325 19.3944
R10469 gnd.n4325 gnd.n4324 19.3944
R10470 gnd.n4324 gnd.n4323 19.3944
R10471 gnd.n4323 gnd.n4320 19.3944
R10472 gnd.n4320 gnd.n4319 19.3944
R10473 gnd.n4319 gnd.n4317 19.3944
R10474 gnd.n4317 gnd.n4316 19.3944
R10475 gnd.n4316 gnd.n4315 19.3944
R10476 gnd.n4315 gnd.n4312 19.3944
R10477 gnd.n4312 gnd.n4311 19.3944
R10478 gnd.n4311 gnd.n4309 19.3944
R10479 gnd.n4309 gnd.n4308 19.3944
R10480 gnd.n4308 gnd.n1713 19.3944
R10481 gnd.n4489 gnd.n1713 19.3944
R10482 gnd.n4489 gnd.n1711 19.3944
R10483 gnd.n4493 gnd.n1711 19.3944
R10484 gnd.n4494 gnd.n4493 19.3944
R10485 gnd.n4497 gnd.n4494 19.3944
R10486 gnd.n4497 gnd.n1709 19.3944
R10487 gnd.n4529 gnd.n1709 19.3944
R10488 gnd.n4529 gnd.n4528 19.3944
R10489 gnd.n4528 gnd.n4527 19.3944
R10490 gnd.n4527 gnd.n4526 19.3944
R10491 gnd.n4526 gnd.n4520 19.3944
R10492 gnd.n4520 gnd.n4519 19.3944
R10493 gnd.n4519 gnd.n4518 19.3944
R10494 gnd.n4518 gnd.n4517 19.3944
R10495 gnd.n4517 gnd.n4514 19.3944
R10496 gnd.n4514 gnd.n4513 19.3944
R10497 gnd.n4513 gnd.n346 19.3944
R10498 gnd.n7377 gnd.n346 19.3944
R10499 gnd.n7377 gnd.n7376 19.3944
R10500 gnd.n7376 gnd.n7375 19.3944
R10501 gnd.n7375 gnd.n394 19.3944
R10502 gnd.n394 gnd.n393 19.3944
R10503 gnd.n393 gnd.n391 19.3944
R10504 gnd.n391 gnd.n390 19.3944
R10505 gnd.n390 gnd.n388 19.3944
R10506 gnd.n388 gnd.n387 19.3944
R10507 gnd.n387 gnd.n385 19.3944
R10508 gnd.n385 gnd.n384 19.3944
R10509 gnd.n384 gnd.n382 19.3944
R10510 gnd.n382 gnd.n381 19.3944
R10511 gnd.n381 gnd.n379 19.3944
R10512 gnd.n379 gnd.n378 19.3944
R10513 gnd.n378 gnd.n376 19.3944
R10514 gnd.n376 gnd.n375 19.3944
R10515 gnd.n375 gnd.n373 19.3944
R10516 gnd.n373 gnd.n372 19.3944
R10517 gnd.n372 gnd.n370 19.3944
R10518 gnd.n370 gnd.n369 19.3944
R10519 gnd.n369 gnd.n200 19.3944
R10520 gnd.n7589 gnd.n200 19.3944
R10521 gnd.n7590 gnd.n7589 19.3944
R10522 gnd.n7628 gnd.n161 19.3944
R10523 gnd.n7623 gnd.n161 19.3944
R10524 gnd.n7623 gnd.n7622 19.3944
R10525 gnd.n7622 gnd.n7621 19.3944
R10526 gnd.n7621 gnd.n168 19.3944
R10527 gnd.n7616 gnd.n168 19.3944
R10528 gnd.n7616 gnd.n7615 19.3944
R10529 gnd.n7615 gnd.n7614 19.3944
R10530 gnd.n7614 gnd.n175 19.3944
R10531 gnd.n7609 gnd.n175 19.3944
R10532 gnd.n7609 gnd.n7608 19.3944
R10533 gnd.n7608 gnd.n7607 19.3944
R10534 gnd.n7607 gnd.n182 19.3944
R10535 gnd.n7602 gnd.n182 19.3944
R10536 gnd.n7602 gnd.n7601 19.3944
R10537 gnd.n7601 gnd.n7600 19.3944
R10538 gnd.n7600 gnd.n189 19.3944
R10539 gnd.n7595 gnd.n189 19.3944
R10540 gnd.n7661 gnd.n7660 19.3944
R10541 gnd.n7660 gnd.n7659 19.3944
R10542 gnd.n7659 gnd.n133 19.3944
R10543 gnd.n7654 gnd.n133 19.3944
R10544 gnd.n7654 gnd.n7653 19.3944
R10545 gnd.n7653 gnd.n7652 19.3944
R10546 gnd.n7652 gnd.n140 19.3944
R10547 gnd.n7647 gnd.n140 19.3944
R10548 gnd.n7647 gnd.n7646 19.3944
R10549 gnd.n7646 gnd.n7645 19.3944
R10550 gnd.n7645 gnd.n147 19.3944
R10551 gnd.n7640 gnd.n147 19.3944
R10552 gnd.n7640 gnd.n7639 19.3944
R10553 gnd.n7639 gnd.n7638 19.3944
R10554 gnd.n7638 gnd.n154 19.3944
R10555 gnd.n7633 gnd.n154 19.3944
R10556 gnd.n7633 gnd.n7632 19.3944
R10557 gnd.n4607 gnd.n1640 19.3944
R10558 gnd.n4607 gnd.n4606 19.3944
R10559 gnd.n4606 gnd.n4605 19.3944
R10560 gnd.n4605 gnd.n1644 19.3944
R10561 gnd.n1823 gnd.n1644 19.3944
R10562 gnd.n1823 gnd.n1802 19.3944
R10563 gnd.n4361 gnd.n1802 19.3944
R10564 gnd.n4361 gnd.n1800 19.3944
R10565 gnd.n4367 gnd.n1800 19.3944
R10566 gnd.n4367 gnd.n4366 19.3944
R10567 gnd.n4366 gnd.n1776 19.3944
R10568 gnd.n4393 gnd.n1776 19.3944
R10569 gnd.n4393 gnd.n1774 19.3944
R10570 gnd.n4399 gnd.n1774 19.3944
R10571 gnd.n4399 gnd.n4398 19.3944
R10572 gnd.n4398 gnd.n1750 19.3944
R10573 gnd.n4425 gnd.n1750 19.3944
R10574 gnd.n4425 gnd.n1748 19.3944
R10575 gnd.n4431 gnd.n1748 19.3944
R10576 gnd.n4431 gnd.n4430 19.3944
R10577 gnd.n4430 gnd.n1723 19.3944
R10578 gnd.n4479 gnd.n1723 19.3944
R10579 gnd.n4479 gnd.n1721 19.3944
R10580 gnd.n4485 gnd.n1721 19.3944
R10581 gnd.n4485 gnd.n4484 19.3944
R10582 gnd.n4484 gnd.n1688 19.3944
R10583 gnd.n1688 gnd.n307 19.3944
R10584 gnd.n7416 gnd.n7415 19.3944
R10585 gnd.n4545 gnd.n4544 19.3944
R10586 gnd.n1702 gnd.n1701 19.3944
R10587 gnd.n331 gnd.n330 19.3944
R10588 gnd.n7396 gnd.n300 19.3944
R10589 gnd.n7420 gnd.n300 19.3944
R10590 gnd.n7420 gnd.n285 19.3944
R10591 gnd.n7432 gnd.n285 19.3944
R10592 gnd.n7432 gnd.n283 19.3944
R10593 gnd.n7436 gnd.n283 19.3944
R10594 gnd.n7436 gnd.n270 19.3944
R10595 gnd.n7448 gnd.n270 19.3944
R10596 gnd.n7448 gnd.n268 19.3944
R10597 gnd.n7452 gnd.n268 19.3944
R10598 gnd.n7452 gnd.n254 19.3944
R10599 gnd.n7464 gnd.n254 19.3944
R10600 gnd.n7464 gnd.n252 19.3944
R10601 gnd.n7468 gnd.n252 19.3944
R10602 gnd.n7468 gnd.n240 19.3944
R10603 gnd.n7480 gnd.n240 19.3944
R10604 gnd.n7480 gnd.n238 19.3944
R10605 gnd.n7484 gnd.n238 19.3944
R10606 gnd.n7484 gnd.n224 19.3944
R10607 gnd.n7496 gnd.n224 19.3944
R10608 gnd.n7496 gnd.n222 19.3944
R10609 gnd.n7500 gnd.n222 19.3944
R10610 gnd.n7500 gnd.n207 19.3944
R10611 gnd.n7580 gnd.n207 19.3944
R10612 gnd.n7580 gnd.n205 19.3944
R10613 gnd.n7584 gnd.n205 19.3944
R10614 gnd.n7584 gnd.n128 19.3944
R10615 gnd.n7664 gnd.n128 19.3944
R10616 gnd.n2760 gnd.n2753 19.3944
R10617 gnd.n2760 gnd.n2751 19.3944
R10618 gnd.n2764 gnd.n2751 19.3944
R10619 gnd.n2764 gnd.n2749 19.3944
R10620 gnd.n2855 gnd.n2749 19.3944
R10621 gnd.n2855 gnd.n2854 19.3944
R10622 gnd.n2854 gnd.n2853 19.3944
R10623 gnd.n2849 gnd.n2770 19.3944
R10624 gnd.n2845 gnd.n2775 19.3944
R10625 gnd.n2843 gnd.n2842 19.3944
R10626 gnd.n2839 gnd.n2838 19.3944
R10627 gnd.n2835 gnd.n2834 19.3944
R10628 gnd.n2834 gnd.n2833 19.3944
R10629 gnd.n2833 gnd.n2779 19.3944
R10630 gnd.n2829 gnd.n2779 19.3944
R10631 gnd.n2829 gnd.n2828 19.3944
R10632 gnd.n2828 gnd.n2827 19.3944
R10633 gnd.n2827 gnd.n2785 19.3944
R10634 gnd.n2823 gnd.n2785 19.3944
R10635 gnd.n2823 gnd.n2822 19.3944
R10636 gnd.n2822 gnd.n2821 19.3944
R10637 gnd.n2821 gnd.n2791 19.3944
R10638 gnd.n2817 gnd.n2791 19.3944
R10639 gnd.n2817 gnd.n2816 19.3944
R10640 gnd.n2816 gnd.n2815 19.3944
R10641 gnd.n2815 gnd.n2797 19.3944
R10642 gnd.n2811 gnd.n2797 19.3944
R10643 gnd.n2811 gnd.n2810 19.3944
R10644 gnd.n2810 gnd.n2809 19.3944
R10645 gnd.n2809 gnd.n2806 19.3944
R10646 gnd.n2806 gnd.n2805 19.3944
R10647 gnd.n2805 gnd.n2686 19.3944
R10648 gnd.n3200 gnd.n2686 19.3944
R10649 gnd.n3200 gnd.n2684 19.3944
R10650 gnd.n3204 gnd.n2684 19.3944
R10651 gnd.n3204 gnd.n2682 19.3944
R10652 gnd.n3208 gnd.n2682 19.3944
R10653 gnd.n3208 gnd.n2680 19.3944
R10654 gnd.n3212 gnd.n2680 19.3944
R10655 gnd.n3212 gnd.n2678 19.3944
R10656 gnd.n3217 gnd.n2678 19.3944
R10657 gnd.n3217 gnd.n2676 19.3944
R10658 gnd.n3226 gnd.n2676 19.3944
R10659 gnd.n3226 gnd.n3225 19.3944
R10660 gnd.n3225 gnd.n3224 19.3944
R10661 gnd.n3224 gnd.n2553 19.3944
R10662 gnd.n3395 gnd.n2553 19.3944
R10663 gnd.n3395 gnd.n2551 19.3944
R10664 gnd.n3401 gnd.n2551 19.3944
R10665 gnd.n3401 gnd.n3400 19.3944
R10666 gnd.n3400 gnd.n2528 19.3944
R10667 gnd.n3425 gnd.n2528 19.3944
R10668 gnd.n3425 gnd.n2526 19.3944
R10669 gnd.n3437 gnd.n2526 19.3944
R10670 gnd.n3437 gnd.n3436 19.3944
R10671 gnd.n3436 gnd.n3435 19.3944
R10672 gnd.n3435 gnd.n3432 19.3944
R10673 gnd.n3432 gnd.n2493 19.3944
R10674 gnd.n3472 gnd.n2493 19.3944
R10675 gnd.n3472 gnd.n2491 19.3944
R10676 gnd.n3478 gnd.n2491 19.3944
R10677 gnd.n3478 gnd.n3477 19.3944
R10678 gnd.n3477 gnd.n2478 19.3944
R10679 gnd.n3594 gnd.n2478 19.3944
R10680 gnd.n3594 gnd.n2476 19.3944
R10681 gnd.n3598 gnd.n2476 19.3944
R10682 gnd.n3598 gnd.n2457 19.3944
R10683 gnd.n3621 gnd.n2457 19.3944
R10684 gnd.n3621 gnd.n2455 19.3944
R10685 gnd.n3627 gnd.n2455 19.3944
R10686 gnd.n3627 gnd.n3626 19.3944
R10687 gnd.n3626 gnd.n2424 19.3944
R10688 gnd.n3663 gnd.n2424 19.3944
R10689 gnd.n3663 gnd.n2422 19.3944
R10690 gnd.n3678 gnd.n2422 19.3944
R10691 gnd.n3678 gnd.n3677 19.3944
R10692 gnd.n3677 gnd.n3676 19.3944
R10693 gnd.n3676 gnd.n3670 19.3944
R10694 gnd.n3670 gnd.n2390 19.3944
R10695 gnd.n3746 gnd.n2390 19.3944
R10696 gnd.n3746 gnd.n2388 19.3944
R10697 gnd.n3750 gnd.n2388 19.3944
R10698 gnd.n3750 gnd.n2367 19.3944
R10699 gnd.n3789 gnd.n2367 19.3944
R10700 gnd.n3789 gnd.n2365 19.3944
R10701 gnd.n3793 gnd.n2365 19.3944
R10702 gnd.n3793 gnd.n2351 19.3944
R10703 gnd.n3837 gnd.n2351 19.3944
R10704 gnd.n3837 gnd.n2349 19.3944
R10705 gnd.n3843 gnd.n2349 19.3944
R10706 gnd.n3843 gnd.n3842 19.3944
R10707 gnd.n3842 gnd.n2322 19.3944
R10708 gnd.n3874 gnd.n2322 19.3944
R10709 gnd.n3874 gnd.n2320 19.3944
R10710 gnd.n3878 gnd.n2320 19.3944
R10711 gnd.n3878 gnd.n2285 19.3944
R10712 gnd.n3908 gnd.n2285 19.3944
R10713 gnd.n3908 gnd.n2283 19.3944
R10714 gnd.n3914 gnd.n2283 19.3944
R10715 gnd.n3914 gnd.n3913 19.3944
R10716 gnd.n3913 gnd.n2256 19.3944
R10717 gnd.n3960 gnd.n2256 19.3944
R10718 gnd.n3960 gnd.n2254 19.3944
R10719 gnd.n3964 gnd.n2254 19.3944
R10720 gnd.n3964 gnd.n2237 19.3944
R10721 gnd.n3986 gnd.n2237 19.3944
R10722 gnd.n3986 gnd.n2235 19.3944
R10723 gnd.n3992 gnd.n2235 19.3944
R10724 gnd.n3992 gnd.n3991 19.3944
R10725 gnd.n3991 gnd.n2036 19.3944
R10726 gnd.n4178 gnd.n2036 19.3944
R10727 gnd.n4178 gnd.n2034 19.3944
R10728 gnd.n4182 gnd.n2034 19.3944
R10729 gnd.n4182 gnd.n2024 19.3944
R10730 gnd.n4199 gnd.n2024 19.3944
R10731 gnd.n4199 gnd.n2022 19.3944
R10732 gnd.n4203 gnd.n2022 19.3944
R10733 gnd.n4203 gnd.n2012 19.3944
R10734 gnd.n4220 gnd.n2012 19.3944
R10735 gnd.n4220 gnd.n2010 19.3944
R10736 gnd.n4224 gnd.n2010 19.3944
R10737 gnd.n4224 gnd.n2000 19.3944
R10738 gnd.n4243 gnd.n2000 19.3944
R10739 gnd.n4243 gnd.n1998 19.3944
R10740 gnd.n4248 gnd.n1998 19.3944
R10741 gnd.n4248 gnd.n1617 19.3944
R10742 gnd.n4622 gnd.n1617 19.3944
R10743 gnd.n4622 gnd.n4621 19.3944
R10744 gnd.n4621 gnd.n4620 19.3944
R10745 gnd.n4620 gnd.n1621 19.3944
R10746 gnd.n4614 gnd.n1621 19.3944
R10747 gnd.n4614 gnd.n4613 19.3944
R10748 gnd.n4613 gnd.n4612 19.3944
R10749 gnd.n4612 gnd.n1630 19.3944
R10750 gnd.n1814 gnd.n1630 19.3944
R10751 gnd.n1818 gnd.n1814 19.3944
R10752 gnd.n1818 gnd.n1812 19.3944
R10753 gnd.n4350 gnd.n1812 19.3944
R10754 gnd.n4350 gnd.n1810 19.3944
R10755 gnd.n4356 gnd.n1810 19.3944
R10756 gnd.n4356 gnd.n4355 19.3944
R10757 gnd.n4355 gnd.n1785 19.3944
R10758 gnd.n4381 gnd.n1785 19.3944
R10759 gnd.n4381 gnd.n1783 19.3944
R10760 gnd.n4387 gnd.n1783 19.3944
R10761 gnd.n4387 gnd.n4386 19.3944
R10762 gnd.n4386 gnd.n1759 19.3944
R10763 gnd.n4414 gnd.n1759 19.3944
R10764 gnd.n4414 gnd.n1757 19.3944
R10765 gnd.n4420 gnd.n1757 19.3944
R10766 gnd.n4420 gnd.n4419 19.3944
R10767 gnd.n4419 gnd.n1732 19.3944
R10768 gnd.n4451 gnd.n1732 19.3944
R10769 gnd.n4451 gnd.n1730 19.3944
R10770 gnd.n4474 gnd.n1730 19.3944
R10771 gnd.n4474 gnd.n4473 19.3944
R10772 gnd.n4473 gnd.n4472 19.3944
R10773 gnd.n4472 gnd.n4457 19.3944
R10774 gnd.n4466 gnd.n4457 19.3944
R10775 gnd.n4466 gnd.n4465 19.3944
R10776 gnd.n4463 gnd.n4461 19.3944
R10777 gnd.n4535 gnd.n4534 19.3944
R10778 gnd.n4539 gnd.n4538 19.3944
R10779 gnd.n7391 gnd.n336 19.3944
R10780 gnd.n7389 gnd.n7388 19.3944
R10781 gnd.n7388 gnd.n338 19.3944
R10782 gnd.n7384 gnd.n338 19.3944
R10783 gnd.n7384 gnd.n7383 19.3944
R10784 gnd.n7383 gnd.n7382 19.3944
R10785 gnd.n7382 gnd.n344 19.3944
R10786 gnd.n7370 gnd.n344 19.3944
R10787 gnd.n5104 gnd.n5103 19.3944
R10788 gnd.n5103 gnd.n5102 19.3944
R10789 gnd.n5102 gnd.n5101 19.3944
R10790 gnd.n5101 gnd.n5099 19.3944
R10791 gnd.n5099 gnd.n5096 19.3944
R10792 gnd.n5096 gnd.n5095 19.3944
R10793 gnd.n5095 gnd.n5092 19.3944
R10794 gnd.n5092 gnd.n5091 19.3944
R10795 gnd.n5091 gnd.n5088 19.3944
R10796 gnd.n5088 gnd.n5087 19.3944
R10797 gnd.n5087 gnd.n5084 19.3944
R10798 gnd.n5084 gnd.n5083 19.3944
R10799 gnd.n5083 gnd.n5080 19.3944
R10800 gnd.n5080 gnd.n5079 19.3944
R10801 gnd.n5079 gnd.n5076 19.3944
R10802 gnd.n5076 gnd.n5075 19.3944
R10803 gnd.n5075 gnd.n5072 19.3944
R10804 gnd.n5070 gnd.n5067 19.3944
R10805 gnd.n5067 gnd.n5066 19.3944
R10806 gnd.n5066 gnd.n5063 19.3944
R10807 gnd.n5063 gnd.n5062 19.3944
R10808 gnd.n5062 gnd.n5059 19.3944
R10809 gnd.n5059 gnd.n5058 19.3944
R10810 gnd.n5058 gnd.n5055 19.3944
R10811 gnd.n5055 gnd.n5054 19.3944
R10812 gnd.n5054 gnd.n5051 19.3944
R10813 gnd.n5051 gnd.n5050 19.3944
R10814 gnd.n5050 gnd.n5047 19.3944
R10815 gnd.n5047 gnd.n5046 19.3944
R10816 gnd.n5046 gnd.n5043 19.3944
R10817 gnd.n5043 gnd.n5042 19.3944
R10818 gnd.n5042 gnd.n5039 19.3944
R10819 gnd.n5039 gnd.n5038 19.3944
R10820 gnd.n5038 gnd.n5035 19.3944
R10821 gnd.n5035 gnd.n5034 19.3944
R10822 gnd.n2984 gnd.n2916 19.3944
R10823 gnd.n2984 gnd.n2917 19.3944
R10824 gnd.n2980 gnd.n2917 19.3944
R10825 gnd.n2980 gnd.n1111 19.3944
R10826 gnd.n5012 gnd.n1111 19.3944
R10827 gnd.n5012 gnd.n5011 19.3944
R10828 gnd.n5011 gnd.n5010 19.3944
R10829 gnd.n5010 gnd.n1115 19.3944
R10830 gnd.n5000 gnd.n1115 19.3944
R10831 gnd.n5000 gnd.n4999 19.3944
R10832 gnd.n4999 gnd.n4998 19.3944
R10833 gnd.n4998 gnd.n1134 19.3944
R10834 gnd.n4988 gnd.n1134 19.3944
R10835 gnd.n4988 gnd.n4987 19.3944
R10836 gnd.n4987 gnd.n4986 19.3944
R10837 gnd.n4986 gnd.n1155 19.3944
R10838 gnd.n4976 gnd.n1155 19.3944
R10839 gnd.n4976 gnd.n4975 19.3944
R10840 gnd.n4975 gnd.n4974 19.3944
R10841 gnd.n4974 gnd.n1174 19.3944
R10842 gnd.n4964 gnd.n1174 19.3944
R10843 gnd.n4964 gnd.n4963 19.3944
R10844 gnd.n4963 gnd.n4962 19.3944
R10845 gnd.n4962 gnd.n1196 19.3944
R10846 gnd.n4952 gnd.n1196 19.3944
R10847 gnd.n4952 gnd.n4951 19.3944
R10848 gnd.n4951 gnd.n4950 19.3944
R10849 gnd.n4950 gnd.n1217 19.3944
R10850 gnd.n4939 gnd.n1217 19.3944
R10851 gnd.n4939 gnd.n4938 19.3944
R10852 gnd.n4938 gnd.n4937 19.3944
R10853 gnd.n4937 gnd.n1237 19.3944
R10854 gnd.n4926 gnd.n1237 19.3944
R10855 gnd.n4926 gnd.n4925 19.3944
R10856 gnd.n4925 gnd.n4924 19.3944
R10857 gnd.n4924 gnd.n1254 19.3944
R10858 gnd.n4913 gnd.n1254 19.3944
R10859 gnd.n4913 gnd.n4912 19.3944
R10860 gnd.n4912 gnd.n4911 19.3944
R10861 gnd.n4911 gnd.n1273 19.3944
R10862 gnd.n4901 gnd.n1273 19.3944
R10863 gnd.n4901 gnd.n4900 19.3944
R10864 gnd.n4900 gnd.n4899 19.3944
R10865 gnd.n4899 gnd.n1294 19.3944
R10866 gnd.n4889 gnd.n1294 19.3944
R10867 gnd.n4889 gnd.n4888 19.3944
R10868 gnd.n4888 gnd.n4887 19.3944
R10869 gnd.n4887 gnd.n1315 19.3944
R10870 gnd.n4877 gnd.n1315 19.3944
R10871 gnd.n4877 gnd.n4876 19.3944
R10872 gnd.n4876 gnd.n4875 19.3944
R10873 gnd.n4875 gnd.n1336 19.3944
R10874 gnd.n4865 gnd.n1336 19.3944
R10875 gnd.n4865 gnd.n4864 19.3944
R10876 gnd.n4864 gnd.n4863 19.3944
R10877 gnd.n4863 gnd.n1357 19.3944
R10878 gnd.n4853 gnd.n1357 19.3944
R10879 gnd.n4853 gnd.n4852 19.3944
R10880 gnd.n4852 gnd.n4851 19.3944
R10881 gnd.n4851 gnd.n1378 19.3944
R10882 gnd.n4841 gnd.n1378 19.3944
R10883 gnd.n4841 gnd.n4840 19.3944
R10884 gnd.n4840 gnd.n4839 19.3944
R10885 gnd.n4839 gnd.n1400 19.3944
R10886 gnd.n2976 gnd.n2974 19.3944
R10887 gnd.n2974 gnd.n2971 19.3944
R10888 gnd.n2971 gnd.n2970 19.3944
R10889 gnd.n2970 gnd.n2967 19.3944
R10890 gnd.n2967 gnd.n2966 19.3944
R10891 gnd.n2966 gnd.n2963 19.3944
R10892 gnd.n2963 gnd.n2962 19.3944
R10893 gnd.n2962 gnd.n2959 19.3944
R10894 gnd.n2959 gnd.n2958 19.3944
R10895 gnd.n2958 gnd.n2955 19.3944
R10896 gnd.n2955 gnd.n2954 19.3944
R10897 gnd.n2954 gnd.n2951 19.3944
R10898 gnd.n2951 gnd.n2950 19.3944
R10899 gnd.n2950 gnd.n2947 19.3944
R10900 gnd.n2947 gnd.n2946 19.3944
R10901 gnd.n2946 gnd.n2943 19.3944
R10902 gnd.n2937 gnd.n2912 19.3944
R10903 gnd.n2995 gnd.n2912 19.3944
R10904 gnd.n2995 gnd.n2910 19.3944
R10905 gnd.n3000 gnd.n2910 19.3944
R10906 gnd.n3001 gnd.n3000 19.3944
R10907 gnd.n3003 gnd.n3001 19.3944
R10908 gnd.n3003 gnd.n2908 19.3944
R10909 gnd.n3008 gnd.n2908 19.3944
R10910 gnd.n3009 gnd.n3008 19.3944
R10911 gnd.n3011 gnd.n3009 19.3944
R10912 gnd.n3011 gnd.n2906 19.3944
R10913 gnd.n3016 gnd.n2906 19.3944
R10914 gnd.n3017 gnd.n3016 19.3944
R10915 gnd.n3019 gnd.n3017 19.3944
R10916 gnd.n3019 gnd.n2904 19.3944
R10917 gnd.n3024 gnd.n2904 19.3944
R10918 gnd.n3025 gnd.n3024 19.3944
R10919 gnd.n3027 gnd.n3025 19.3944
R10920 gnd.n3027 gnd.n2902 19.3944
R10921 gnd.n3031 gnd.n2902 19.3944
R10922 gnd.n3031 gnd.n2863 19.3944
R10923 gnd.n3043 gnd.n2863 19.3944
R10924 gnd.n3043 gnd.n2861 19.3944
R10925 gnd.n3047 gnd.n2861 19.3944
R10926 gnd.n3047 gnd.n2746 19.3944
R10927 gnd.n3059 gnd.n2746 19.3944
R10928 gnd.n3059 gnd.n2744 19.3944
R10929 gnd.n3063 gnd.n2744 19.3944
R10930 gnd.n3063 gnd.n2740 19.3944
R10931 gnd.n3075 gnd.n2740 19.3944
R10932 gnd.n3075 gnd.n2738 19.3944
R10933 gnd.n3079 gnd.n2738 19.3944
R10934 gnd.n3079 gnd.n2732 19.3944
R10935 gnd.n3091 gnd.n2732 19.3944
R10936 gnd.n3091 gnd.n2730 19.3944
R10937 gnd.n3095 gnd.n2730 19.3944
R10938 gnd.n3095 gnd.n2726 19.3944
R10939 gnd.n3107 gnd.n2726 19.3944
R10940 gnd.n3107 gnd.n2724 19.3944
R10941 gnd.n3111 gnd.n2724 19.3944
R10942 gnd.n3111 gnd.n2719 19.3944
R10943 gnd.n3123 gnd.n2719 19.3944
R10944 gnd.n3123 gnd.n2717 19.3944
R10945 gnd.n3127 gnd.n2717 19.3944
R10946 gnd.n3127 gnd.n2712 19.3944
R10947 gnd.n3139 gnd.n2712 19.3944
R10948 gnd.n3139 gnd.n2710 19.3944
R10949 gnd.n3143 gnd.n2710 19.3944
R10950 gnd.n3143 gnd.n2705 19.3944
R10951 gnd.n3155 gnd.n2705 19.3944
R10952 gnd.n3155 gnd.n2703 19.3944
R10953 gnd.n3159 gnd.n2703 19.3944
R10954 gnd.n3159 gnd.n2698 19.3944
R10955 gnd.n3172 gnd.n2698 19.3944
R10956 gnd.n3172 gnd.n2696 19.3944
R10957 gnd.n3176 gnd.n2696 19.3944
R10958 gnd.n3176 gnd.n2689 19.3944
R10959 gnd.n3194 gnd.n2689 19.3944
R10960 gnd.n3194 gnd.n2690 19.3944
R10961 gnd.n3190 gnd.n2690 19.3944
R10962 gnd.n3190 gnd.n2628 19.3944
R10963 gnd.n3256 gnd.n2628 19.3944
R10964 gnd.n3256 gnd.n2629 19.3944
R10965 gnd.n2629 gnd.n2623 19.3944
R10966 gnd.n5027 gnd.n5026 19.3944
R10967 gnd.n5026 gnd.n1089 19.3944
R10968 gnd.n5022 gnd.n1089 19.3944
R10969 gnd.n5022 gnd.n1091 19.3944
R10970 gnd.n2872 gnd.n1091 19.3944
R10971 gnd.n2876 gnd.n2872 19.3944
R10972 gnd.n2877 gnd.n2876 19.3944
R10973 gnd.n2879 gnd.n2877 19.3944
R10974 gnd.n2879 gnd.n2870 19.3944
R10975 gnd.n2884 gnd.n2870 19.3944
R10976 gnd.n2885 gnd.n2884 19.3944
R10977 gnd.n2887 gnd.n2885 19.3944
R10978 gnd.n2887 gnd.n2868 19.3944
R10979 gnd.n2892 gnd.n2868 19.3944
R10980 gnd.n2893 gnd.n2892 19.3944
R10981 gnd.n2895 gnd.n2893 19.3944
R10982 gnd.n2895 gnd.n2866 19.3944
R10983 gnd.n2900 gnd.n2866 19.3944
R10984 gnd.n2901 gnd.n2900 19.3944
R10985 gnd.n3035 gnd.n2901 19.3944
R10986 gnd.n3035 gnd.n2864 19.3944
R10987 gnd.n3039 gnd.n2864 19.3944
R10988 gnd.n3039 gnd.n2860 19.3944
R10989 gnd.n3051 gnd.n2860 19.3944
R10990 gnd.n3051 gnd.n2858 19.3944
R10991 gnd.n3055 gnd.n2858 19.3944
R10992 gnd.n3055 gnd.n2743 19.3944
R10993 gnd.n3067 gnd.n2743 19.3944
R10994 gnd.n3067 gnd.n2741 19.3944
R10995 gnd.n3071 gnd.n2741 19.3944
R10996 gnd.n3071 gnd.n2737 19.3944
R10997 gnd.n3083 gnd.n2737 19.3944
R10998 gnd.n3083 gnd.n2734 19.3944
R10999 gnd.n3087 gnd.n2734 19.3944
R11000 gnd.n3087 gnd.n2729 19.3944
R11001 gnd.n3099 gnd.n2729 19.3944
R11002 gnd.n3099 gnd.n2727 19.3944
R11003 gnd.n3103 gnd.n2727 19.3944
R11004 gnd.n3103 gnd.n2723 19.3944
R11005 gnd.n3115 gnd.n2723 19.3944
R11006 gnd.n3115 gnd.n2721 19.3944
R11007 gnd.n3119 gnd.n2721 19.3944
R11008 gnd.n3119 gnd.n2715 19.3944
R11009 gnd.n3131 gnd.n2715 19.3944
R11010 gnd.n3131 gnd.n2713 19.3944
R11011 gnd.n3135 gnd.n2713 19.3944
R11012 gnd.n3135 gnd.n2709 19.3944
R11013 gnd.n3147 gnd.n2709 19.3944
R11014 gnd.n3147 gnd.n2707 19.3944
R11015 gnd.n3151 gnd.n2707 19.3944
R11016 gnd.n3151 gnd.n2701 19.3944
R11017 gnd.n3163 gnd.n2701 19.3944
R11018 gnd.n3163 gnd.n2699 19.3944
R11019 gnd.n3168 gnd.n2699 19.3944
R11020 gnd.n3168 gnd.n2694 19.3944
R11021 gnd.n3180 gnd.n2694 19.3944
R11022 gnd.n3181 gnd.n3180 19.3944
R11023 gnd.n3182 gnd.n3181 19.3944
R11024 gnd.n3182 gnd.n2692 19.3944
R11025 gnd.n3186 gnd.n2692 19.3944
R11026 gnd.n3186 gnd.n2627 19.3944
R11027 gnd.n3260 gnd.n2627 19.3944
R11028 gnd.n3260 gnd.n2625 19.3944
R11029 gnd.n3327 gnd.n2625 19.3944
R11030 gnd.n3277 gnd.n1457 19.3944
R11031 gnd.n3281 gnd.n3277 19.3944
R11032 gnd.n3284 gnd.n3281 19.3944
R11033 gnd.n3287 gnd.n3284 19.3944
R11034 gnd.n3287 gnd.n3273 19.3944
R11035 gnd.n3291 gnd.n3273 19.3944
R11036 gnd.n3294 gnd.n3291 19.3944
R11037 gnd.n3297 gnd.n3294 19.3944
R11038 gnd.n3297 gnd.n3271 19.3944
R11039 gnd.n3301 gnd.n3271 19.3944
R11040 gnd.n3304 gnd.n3301 19.3944
R11041 gnd.n3307 gnd.n3304 19.3944
R11042 gnd.n3307 gnd.n3269 19.3944
R11043 gnd.n3311 gnd.n3269 19.3944
R11044 gnd.n3314 gnd.n3311 19.3944
R11045 gnd.n3317 gnd.n3314 19.3944
R11046 gnd.n3317 gnd.n3267 19.3944
R11047 gnd.n3322 gnd.n3267 19.3944
R11048 gnd.n4831 gnd.n1410 19.3944
R11049 gnd.n4826 gnd.n1410 19.3944
R11050 gnd.n4826 gnd.n4825 19.3944
R11051 gnd.n4825 gnd.n4824 19.3944
R11052 gnd.n4824 gnd.n4821 19.3944
R11053 gnd.n4821 gnd.n4820 19.3944
R11054 gnd.n4820 gnd.n4817 19.3944
R11055 gnd.n4817 gnd.n4816 19.3944
R11056 gnd.n4816 gnd.n4813 19.3944
R11057 gnd.n4813 gnd.n4812 19.3944
R11058 gnd.n4812 gnd.n4809 19.3944
R11059 gnd.n4809 gnd.n4808 19.3944
R11060 gnd.n4808 gnd.n4805 19.3944
R11061 gnd.n4805 gnd.n4804 19.3944
R11062 gnd.n4804 gnd.n4801 19.3944
R11063 gnd.n2990 gnd.n2986 19.3944
R11064 gnd.n2990 gnd.n1100 19.3944
R11065 gnd.n5018 gnd.n1100 19.3944
R11066 gnd.n5018 gnd.n5017 19.3944
R11067 gnd.n5017 gnd.n5016 19.3944
R11068 gnd.n5016 gnd.n1104 19.3944
R11069 gnd.n5006 gnd.n1104 19.3944
R11070 gnd.n5006 gnd.n5005 19.3944
R11071 gnd.n5005 gnd.n5004 19.3944
R11072 gnd.n5004 gnd.n1125 19.3944
R11073 gnd.n4994 gnd.n1125 19.3944
R11074 gnd.n4994 gnd.n4993 19.3944
R11075 gnd.n4993 gnd.n4992 19.3944
R11076 gnd.n4992 gnd.n1145 19.3944
R11077 gnd.n4982 gnd.n1145 19.3944
R11078 gnd.n4982 gnd.n4981 19.3944
R11079 gnd.n4981 gnd.n4980 19.3944
R11080 gnd.n4980 gnd.n1165 19.3944
R11081 gnd.n4970 gnd.n1165 19.3944
R11082 gnd.n4970 gnd.n4969 19.3944
R11083 gnd.n4969 gnd.n4968 19.3944
R11084 gnd.n4968 gnd.n1185 19.3944
R11085 gnd.n4958 gnd.n1185 19.3944
R11086 gnd.n4958 gnd.n4957 19.3944
R11087 gnd.n4957 gnd.n4956 19.3944
R11088 gnd.n4956 gnd.n1207 19.3944
R11089 gnd.n4946 gnd.n1207 19.3944
R11090 gnd.n4944 gnd.n4943 19.3944
R11091 gnd.n4933 gnd.n1244 19.3944
R11092 gnd.n4931 gnd.n4930 19.3944
R11093 gnd.n4920 gnd.n1261 19.3944
R11094 gnd.n4918 gnd.n4917 19.3944
R11095 gnd.n4917 gnd.n1262 19.3944
R11096 gnd.n4907 gnd.n1262 19.3944
R11097 gnd.n4907 gnd.n4906 19.3944
R11098 gnd.n4906 gnd.n4905 19.3944
R11099 gnd.n4905 gnd.n1284 19.3944
R11100 gnd.n4895 gnd.n1284 19.3944
R11101 gnd.n4895 gnd.n4894 19.3944
R11102 gnd.n4894 gnd.n4893 19.3944
R11103 gnd.n4893 gnd.n1304 19.3944
R11104 gnd.n4883 gnd.n1304 19.3944
R11105 gnd.n4883 gnd.n4882 19.3944
R11106 gnd.n4882 gnd.n4881 19.3944
R11107 gnd.n4881 gnd.n1326 19.3944
R11108 gnd.n4871 gnd.n1326 19.3944
R11109 gnd.n4871 gnd.n4870 19.3944
R11110 gnd.n4870 gnd.n4869 19.3944
R11111 gnd.n4869 gnd.n1346 19.3944
R11112 gnd.n4859 gnd.n1346 19.3944
R11113 gnd.n4859 gnd.n4858 19.3944
R11114 gnd.n4858 gnd.n4857 19.3944
R11115 gnd.n4857 gnd.n1368 19.3944
R11116 gnd.n4847 gnd.n1368 19.3944
R11117 gnd.n4847 gnd.n4846 19.3944
R11118 gnd.n4846 gnd.n4845 19.3944
R11119 gnd.n4845 gnd.n1389 19.3944
R11120 gnd.n4835 gnd.n1389 19.3944
R11121 gnd.n4835 gnd.n4834 19.3944
R11122 gnd.n6699 gnd.n6698 19.3944
R11123 gnd.n6698 gnd.n6697 19.3944
R11124 gnd.n6697 gnd.n801 19.3944
R11125 gnd.n6691 gnd.n801 19.3944
R11126 gnd.n6691 gnd.n6690 19.3944
R11127 gnd.n6690 gnd.n6689 19.3944
R11128 gnd.n6689 gnd.n809 19.3944
R11129 gnd.n6683 gnd.n809 19.3944
R11130 gnd.n6683 gnd.n6682 19.3944
R11131 gnd.n6682 gnd.n6681 19.3944
R11132 gnd.n6681 gnd.n817 19.3944
R11133 gnd.n6675 gnd.n817 19.3944
R11134 gnd.n6675 gnd.n6674 19.3944
R11135 gnd.n6674 gnd.n6673 19.3944
R11136 gnd.n6673 gnd.n825 19.3944
R11137 gnd.n6667 gnd.n825 19.3944
R11138 gnd.n6667 gnd.n6666 19.3944
R11139 gnd.n6666 gnd.n6665 19.3944
R11140 gnd.n6665 gnd.n833 19.3944
R11141 gnd.n6659 gnd.n833 19.3944
R11142 gnd.n6659 gnd.n6658 19.3944
R11143 gnd.n6658 gnd.n6657 19.3944
R11144 gnd.n6657 gnd.n841 19.3944
R11145 gnd.n6651 gnd.n841 19.3944
R11146 gnd.n6651 gnd.n6650 19.3944
R11147 gnd.n6650 gnd.n6649 19.3944
R11148 gnd.n6649 gnd.n849 19.3944
R11149 gnd.n6643 gnd.n849 19.3944
R11150 gnd.n6643 gnd.n6642 19.3944
R11151 gnd.n6642 gnd.n6641 19.3944
R11152 gnd.n6641 gnd.n857 19.3944
R11153 gnd.n6635 gnd.n857 19.3944
R11154 gnd.n6635 gnd.n6634 19.3944
R11155 gnd.n6634 gnd.n6633 19.3944
R11156 gnd.n6633 gnd.n865 19.3944
R11157 gnd.n6627 gnd.n865 19.3944
R11158 gnd.n6627 gnd.n6626 19.3944
R11159 gnd.n6626 gnd.n6625 19.3944
R11160 gnd.n6625 gnd.n873 19.3944
R11161 gnd.n6619 gnd.n873 19.3944
R11162 gnd.n6619 gnd.n6618 19.3944
R11163 gnd.n6618 gnd.n6617 19.3944
R11164 gnd.n6617 gnd.n881 19.3944
R11165 gnd.n6611 gnd.n881 19.3944
R11166 gnd.n6611 gnd.n6610 19.3944
R11167 gnd.n6610 gnd.n6609 19.3944
R11168 gnd.n6609 gnd.n889 19.3944
R11169 gnd.n6603 gnd.n889 19.3944
R11170 gnd.n6603 gnd.n6602 19.3944
R11171 gnd.n6602 gnd.n6601 19.3944
R11172 gnd.n6601 gnd.n897 19.3944
R11173 gnd.n6595 gnd.n897 19.3944
R11174 gnd.n6595 gnd.n6594 19.3944
R11175 gnd.n6594 gnd.n6593 19.3944
R11176 gnd.n6593 gnd.n905 19.3944
R11177 gnd.n6587 gnd.n905 19.3944
R11178 gnd.n6587 gnd.n6586 19.3944
R11179 gnd.n6586 gnd.n6585 19.3944
R11180 gnd.n6585 gnd.n913 19.3944
R11181 gnd.n6579 gnd.n913 19.3944
R11182 gnd.n6579 gnd.n6578 19.3944
R11183 gnd.n6578 gnd.n6577 19.3944
R11184 gnd.n6577 gnd.n921 19.3944
R11185 gnd.n6571 gnd.n921 19.3944
R11186 gnd.n6571 gnd.n6570 19.3944
R11187 gnd.n6570 gnd.n6569 19.3944
R11188 gnd.n6569 gnd.n929 19.3944
R11189 gnd.n6563 gnd.n929 19.3944
R11190 gnd.n6563 gnd.n6562 19.3944
R11191 gnd.n6562 gnd.n6561 19.3944
R11192 gnd.n6561 gnd.n937 19.3944
R11193 gnd.n6555 gnd.n937 19.3944
R11194 gnd.n6555 gnd.n6554 19.3944
R11195 gnd.n6554 gnd.n6553 19.3944
R11196 gnd.n6553 gnd.n945 19.3944
R11197 gnd.n6547 gnd.n945 19.3944
R11198 gnd.n6547 gnd.n6546 19.3944
R11199 gnd.n6546 gnd.n6545 19.3944
R11200 gnd.n6545 gnd.n953 19.3944
R11201 gnd.n6539 gnd.n953 19.3944
R11202 gnd.n6539 gnd.n6538 19.3944
R11203 gnd.n6538 gnd.n6537 19.3944
R11204 gnd.n6537 gnd.n961 19.3944
R11205 gnd.n2756 gnd.n961 19.3944
R11206 gnd.n3381 gnd.n2566 19.3944
R11207 gnd.n3381 gnd.n2567 19.3944
R11208 gnd.n2567 gnd.n2544 19.3944
R11209 gnd.n3406 gnd.n2544 19.3944
R11210 gnd.n3406 gnd.n2541 19.3944
R11211 gnd.n3411 gnd.n2541 19.3944
R11212 gnd.n3411 gnd.n2542 19.3944
R11213 gnd.n2542 gnd.n2518 19.3944
R11214 gnd.n3442 gnd.n2518 19.3944
R11215 gnd.n3442 gnd.n2516 19.3944
R11216 gnd.n3446 gnd.n2516 19.3944
R11217 gnd.n3446 gnd.n2503 19.3944
R11218 gnd.n3462 gnd.n2503 19.3944
R11219 gnd.n3462 gnd.n2500 19.3944
R11220 gnd.n3467 gnd.n2500 19.3944
R11221 gnd.n3467 gnd.n2501 19.3944
R11222 gnd.n2501 gnd.n1529 19.3944
R11223 gnd.n4723 gnd.n1529 19.3944
R11224 gnd.n4723 gnd.n1530 19.3944
R11225 gnd.n4719 gnd.n1530 19.3944
R11226 gnd.n4719 gnd.n4718 19.3944
R11227 gnd.n4718 gnd.n4717 19.3944
R11228 gnd.n4717 gnd.n1536 19.3944
R11229 gnd.n4713 gnd.n1536 19.3944
R11230 gnd.n4713 gnd.n4712 19.3944
R11231 gnd.n4712 gnd.n4711 19.3944
R11232 gnd.n4711 gnd.n1541 19.3944
R11233 gnd.n4707 gnd.n1541 19.3944
R11234 gnd.n4707 gnd.n4706 19.3944
R11235 gnd.n4706 gnd.n4705 19.3944
R11236 gnd.n4705 gnd.n1546 19.3944
R11237 gnd.n4701 gnd.n1546 19.3944
R11238 gnd.n4701 gnd.n4700 19.3944
R11239 gnd.n4700 gnd.n4699 19.3944
R11240 gnd.n4699 gnd.n1551 19.3944
R11241 gnd.n4695 gnd.n1551 19.3944
R11242 gnd.n4695 gnd.n4694 19.3944
R11243 gnd.n4694 gnd.n4693 19.3944
R11244 gnd.n4693 gnd.n1556 19.3944
R11245 gnd.n4689 gnd.n1556 19.3944
R11246 gnd.n4689 gnd.n4688 19.3944
R11247 gnd.n4688 gnd.n4687 19.3944
R11248 gnd.n4687 gnd.n1561 19.3944
R11249 gnd.n4683 gnd.n1561 19.3944
R11250 gnd.n4683 gnd.n4682 19.3944
R11251 gnd.n4682 gnd.n4681 19.3944
R11252 gnd.n4681 gnd.n1566 19.3944
R11253 gnd.n4677 gnd.n1566 19.3944
R11254 gnd.n4677 gnd.n4676 19.3944
R11255 gnd.n4676 gnd.n4675 19.3944
R11256 gnd.n4675 gnd.n1571 19.3944
R11257 gnd.n4671 gnd.n1571 19.3944
R11258 gnd.n4671 gnd.n4670 19.3944
R11259 gnd.n4670 gnd.n4669 19.3944
R11260 gnd.n4669 gnd.n1576 19.3944
R11261 gnd.n4665 gnd.n1576 19.3944
R11262 gnd.n4665 gnd.n4664 19.3944
R11263 gnd.n4664 gnd.n4663 19.3944
R11264 gnd.n4663 gnd.n1581 19.3944
R11265 gnd.n4659 gnd.n1581 19.3944
R11266 gnd.n4659 gnd.n4658 19.3944
R11267 gnd.n4658 gnd.n4657 19.3944
R11268 gnd.n4657 gnd.n1586 19.3944
R11269 gnd.n4653 gnd.n1586 19.3944
R11270 gnd.n4653 gnd.n4652 19.3944
R11271 gnd.n4652 gnd.n4651 19.3944
R11272 gnd.n4651 gnd.n1591 19.3944
R11273 gnd.n4647 gnd.n1591 19.3944
R11274 gnd.n4647 gnd.n4646 19.3944
R11275 gnd.n4646 gnd.n4645 19.3944
R11276 gnd.n4645 gnd.n1596 19.3944
R11277 gnd.n4641 gnd.n1596 19.3944
R11278 gnd.n4641 gnd.n4640 19.3944
R11279 gnd.n4640 gnd.n4639 19.3944
R11280 gnd.n4639 gnd.n1601 19.3944
R11281 gnd.n4635 gnd.n1601 19.3944
R11282 gnd.n4635 gnd.n4634 19.3944
R11283 gnd.n4634 gnd.n4633 19.3944
R11284 gnd.n4633 gnd.n1606 19.3944
R11285 gnd.n4629 gnd.n1606 19.3944
R11286 gnd.n4629 gnd.n4628 19.3944
R11287 gnd.n4628 gnd.n4627 19.3944
R11288 gnd.n4260 gnd.n4259 19.3944
R11289 gnd.n4259 gnd.n4258 19.3944
R11290 gnd.n4258 gnd.n1993 19.3944
R11291 gnd.n1895 gnd.n1891 19.3944
R11292 gnd.n1895 gnd.n1873 19.3944
R11293 gnd.n1908 gnd.n1873 19.3944
R11294 gnd.n1908 gnd.n1871 19.3944
R11295 gnd.n1914 gnd.n1871 19.3944
R11296 gnd.n1914 gnd.n1864 19.3944
R11297 gnd.n1927 gnd.n1864 19.3944
R11298 gnd.n1927 gnd.n1862 19.3944
R11299 gnd.n1933 gnd.n1862 19.3944
R11300 gnd.n1933 gnd.n1855 19.3944
R11301 gnd.n1946 gnd.n1855 19.3944
R11302 gnd.n1946 gnd.n1853 19.3944
R11303 gnd.n1952 gnd.n1853 19.3944
R11304 gnd.n1952 gnd.n1846 19.3944
R11305 gnd.n1965 gnd.n1846 19.3944
R11306 gnd.n1965 gnd.n1844 19.3944
R11307 gnd.n4272 gnd.n1844 19.3944
R11308 gnd.n4272 gnd.n4271 19.3944
R11309 gnd.n4271 gnd.n4270 19.3944
R11310 gnd.n4270 gnd.n1973 19.3944
R11311 gnd.n4266 gnd.n1973 19.3944
R11312 gnd.n4266 gnd.n4265 19.3944
R11313 gnd.n4265 gnd.n4264 19.3944
R11314 gnd.n4264 gnd.n1981 19.3944
R11315 gnd.n4730 gnd.n4729 18.8883
R11316 gnd.n4090 gnd.n4089 18.8883
R11317 gnd.n5904 gnd.t16 18.8012
R11318 gnd.n5943 gnd.t60 18.8012
R11319 gnd.n5747 gnd.n5489 18.4825
R11320 gnd.n2218 gnd.n2078 18.4247
R11321 gnd.n4801 gnd.n4800 18.4247
R11322 gnd.n7543 gnd.n120 18.2308
R11323 gnd.n1961 gnd.n1841 18.2308
R11324 gnd.n3334 gnd.n3333 18.2308
R11325 gnd.n2943 gnd.n2936 18.2308
R11326 gnd.t6 gnd.n5431 18.1639
R11327 gnd.n5460 gnd.t14 17.5266
R11328 gnd.t10 gnd.n5407 16.8893
R11329 gnd.t151 gnd.n5516 16.2519
R11330 gnd.n5374 gnd.t8 16.2519
R11331 gnd.n3483 gnd.n3482 16.0975
R11332 gnd.n2221 gnd.n2220 16.0975
R11333 gnd.n4732 gnd.n4731 16.0975
R11334 gnd.n4022 gnd.n4021 16.0975
R11335 gnd.n3231 gnd.n2649 15.9333
R11336 gnd.n3231 gnd.n3228 15.9333
R11337 gnd.n2673 gnd.n2672 15.9333
R11338 gnd.n2672 gnd.n2562 15.9333
R11339 gnd.n3383 gnd.n2562 15.9333
R11340 gnd.n3383 gnd.n2563 15.9333
R11341 gnd.n3393 gnd.n2555 15.9333
R11342 gnd.n3393 gnd.n3392 15.9333
R11343 gnd.n3392 gnd.n2546 15.9333
R11344 gnd.n3404 gnd.n2546 15.9333
R11345 gnd.n3404 gnd.n3403 15.9333
R11346 gnd.n3403 gnd.n2548 15.9333
R11347 gnd.n2548 gnd.n2537 15.9333
R11348 gnd.n3413 gnd.n2537 15.9333
R11349 gnd.n2538 gnd.n2530 15.9333
R11350 gnd.n3423 gnd.n2530 15.9333
R11351 gnd.n3423 gnd.n3422 15.9333
R11352 gnd.n3422 gnd.n2520 15.9333
R11353 gnd.n3440 gnd.n2520 15.9333
R11354 gnd.n3440 gnd.n3439 15.9333
R11355 gnd.n3439 gnd.n2522 15.9333
R11356 gnd.n2524 gnd.n2522 15.9333
R11357 gnd.n3448 gnd.n2514 15.9333
R11358 gnd.n2514 gnd.n2513 15.9333
R11359 gnd.n2513 gnd.n2505 15.9333
R11360 gnd.n3460 gnd.n2505 15.9333
R11361 gnd.n3460 gnd.n3459 15.9333
R11362 gnd.n3459 gnd.n2495 15.9333
R11363 gnd.n3470 gnd.n2495 15.9333
R11364 gnd.n3470 gnd.n3469 15.9333
R11365 gnd.n3469 gnd.n2497 15.9333
R11366 gnd.n3480 gnd.n1497 15.9333
R11367 gnd.n4725 gnd.n1526 15.9333
R11368 gnd.n3610 gnd.n3609 15.9333
R11369 gnd.n3652 gnd.n3651 15.9333
R11370 gnd.n2430 gnd.n2419 15.9333
R11371 gnd.n3699 gnd.n2410 15.9333
R11372 gnd.n3672 gnd.n2402 15.9333
R11373 gnd.n3744 gnd.n2393 15.9333
R11374 gnd.n3714 gnd.n2363 15.9333
R11375 gnd.n3795 gnd.n2363 15.9333
R11376 gnd.n3809 gnd.n2341 15.9333
R11377 gnd.n3872 gnd.n3871 15.9333
R11378 gnd.n3881 gnd.n3880 15.9333
R11379 gnd.n3906 gnd.n2287 15.9333
R11380 gnd.n3917 gnd.n3916 15.9333
R11381 gnd.n3957 gnd.n2261 15.9333
R11382 gnd.n3994 gnd.n2225 15.9333
R11383 gnd.n4165 gnd.n4164 15.9333
R11384 gnd.n4164 gnd.n4163 15.9333
R11385 gnd.n4176 gnd.n4175 15.9333
R11386 gnd.n4175 gnd.n4173 15.9333
R11387 gnd.n4173 gnd.n2032 15.9333
R11388 gnd.n4184 gnd.n2032 15.9333
R11389 gnd.n4186 gnd.n4184 15.9333
R11390 gnd.n4186 gnd.n4185 15.9333
R11391 gnd.n4185 gnd.n2026 15.9333
R11392 gnd.n4197 gnd.n2026 15.9333
R11393 gnd.n4197 gnd.n4196 15.9333
R11394 gnd.n4194 gnd.n2020 15.9333
R11395 gnd.n4205 gnd.n2020 15.9333
R11396 gnd.n4207 gnd.n4205 15.9333
R11397 gnd.n4207 gnd.n4206 15.9333
R11398 gnd.n4206 gnd.n2014 15.9333
R11399 gnd.n4218 gnd.n2014 15.9333
R11400 gnd.n4218 gnd.n4217 15.9333
R11401 gnd.n4217 gnd.n4215 15.9333
R11402 gnd.n4226 gnd.n2008 15.9333
R11403 gnd.n4228 gnd.n4226 15.9333
R11404 gnd.n4228 gnd.n4227 15.9333
R11405 gnd.n4227 gnd.n2002 15.9333
R11406 gnd.n4241 gnd.n2002 15.9333
R11407 gnd.n4241 gnd.n4240 15.9333
R11408 gnd.n4240 gnd.n4238 15.9333
R11409 gnd.n4238 gnd.n4237 15.9333
R11410 gnd.n4251 gnd.n4250 15.9333
R11411 gnd.n4251 gnd.n1612 15.9333
R11412 gnd.n4625 gnd.n1612 15.9333
R11413 gnd.n4625 gnd.n4624 15.9333
R11414 gnd.n1623 gnd.n1614 15.9333
R11415 gnd.n4618 gnd.n1623 15.9333
R11416 gnd.n6375 gnd.n6373 15.6674
R11417 gnd.n6343 gnd.n6341 15.6674
R11418 gnd.n6311 gnd.n6309 15.6674
R11419 gnd.n6280 gnd.n6278 15.6674
R11420 gnd.n6248 gnd.n6246 15.6674
R11421 gnd.n6216 gnd.n6214 15.6674
R11422 gnd.n6184 gnd.n6182 15.6674
R11423 gnd.n6153 gnd.n6151 15.6674
R11424 gnd.n5634 gnd.t151 15.6146
R11425 gnd.n6519 gnd.t107 15.6146
R11426 gnd.n6410 gnd.t125 15.6146
R11427 gnd.t161 gnd.n2555 15.6146
R11428 gnd.n4237 gnd.t132 15.6146
R11429 gnd.t185 gnd.n3480 15.296
R11430 gnd.n3690 gnd.n3688 15.296
R11431 gnd.n3709 gnd.n3708 15.296
R11432 gnd.n3862 gnd.n2324 15.296
R11433 gnd.n2318 gnd.n2293 15.296
R11434 gnd.n3934 gnd.t165 15.296
R11435 gnd.n4006 gnd.n4005 15.0827
R11436 gnd.n1509 gnd.n1504 15.0481
R11437 gnd.n4016 gnd.n4015 15.0481
R11438 gnd.n6074 gnd.t15 14.9773
R11439 gnd.n2524 gnd.t77 14.9773
R11440 gnd.t46 gnd.n4194 14.9773
R11441 gnd.n3600 gnd.t168 14.6587
R11442 gnd.n3638 gnd.n2446 14.6587
R11443 gnd.n2305 gnd.n2275 14.6587
R11444 gnd.n3933 gnd.n2244 14.6587
R11445 gnd.n6114 gnd.t57 14.34
R11446 gnd.n6532 gnd.t13 14.34
R11447 gnd.n3997 gnd.n3995 14.0214
R11448 gnd.t74 gnd.n5831 13.7027
R11449 gnd.n5716 gnd.n5712 13.5763
R11450 gnd.n6483 gnd.n5135 13.5763
R11451 gnd.n2179 gnd.n2168 13.5763
R11452 gnd.n7595 gnd.n7594 13.5763
R11453 gnd.n5034 gnd.n1086 13.5763
R11454 gnd.n3323 gnd.n3322 13.5763
R11455 gnd.n5748 gnd.n5747 13.384
R11456 gnd.n3592 gnd.n3591 13.384
R11457 gnd.n3661 gnd.n2426 13.384
R11458 gnd.n3725 gnd.n2385 13.384
R11459 gnd.n3753 gnd.t22 13.384
R11460 gnd.n3787 gnd.t1 13.384
R11461 gnd.n3827 gnd.t54 13.384
R11462 gnd.t51 gnd.n2345 13.384
R11463 gnd.n3846 gnd.n3845 13.384
R11464 gnd.n3918 gnd.n2279 13.384
R11465 gnd.n3982 gnd.n2230 13.384
R11466 gnd.n1520 gnd.n1501 13.1884
R11467 gnd.n1515 gnd.n1514 13.1884
R11468 gnd.n1514 gnd.n1513 13.1884
R11469 gnd.n4009 gnd.n4004 13.1884
R11470 gnd.n4010 gnd.n4009 13.1884
R11471 gnd.n1516 gnd.n1503 13.146
R11472 gnd.n1512 gnd.n1503 13.146
R11473 gnd.n4008 gnd.n4007 13.146
R11474 gnd.n4008 gnd.n4003 13.146
R11475 gnd.n6376 gnd.n6372 12.8005
R11476 gnd.n6344 gnd.n6340 12.8005
R11477 gnd.n6312 gnd.n6308 12.8005
R11478 gnd.n6281 gnd.n6277 12.8005
R11479 gnd.n6249 gnd.n6245 12.8005
R11480 gnd.n6217 gnd.n6213 12.8005
R11481 gnd.n6185 gnd.n6181 12.8005
R11482 gnd.n6154 gnd.n6150 12.8005
R11483 gnd.n4796 gnd.t27 12.7467
R11484 gnd.n3584 gnd.n2473 12.7467
R11485 gnd.n3653 gnd.n2436 12.7467
R11486 gnd.n2386 gnd.n2375 12.7467
R11487 gnd.n3818 gnd.n2354 12.7467
R11488 gnd.n3926 gnd.n2273 12.7467
R11489 gnd.n5002 gnd.t209 12.4281
R11490 gnd.n4972 gnd.n1179 12.4281
R11491 gnd.n274 gnd.n265 12.4281
R11492 gnd.t223 gnd.n226 12.4281
R11493 gnd.n5719 gnd.n5716 12.4126
R11494 gnd.n6486 gnd.n6483 12.4126
R11495 gnd.n2175 gnd.n2168 12.4126
R11496 gnd.n7594 gnd.n196 12.4126
R11497 gnd.n5030 gnd.n1086 12.4126
R11498 gnd.n3324 gnd.n3323 12.4126
R11499 gnd.n4793 gnd.n4730 12.1761
R11500 gnd.n4089 gnd.n4088 12.1761
R11501 gnd.n4726 gnd.n1523 12.1094
R11502 gnd.t84 gnd.n3618 12.1094
R11503 gnd.n3681 gnd.n3680 12.1094
R11504 gnd.n3733 gnd.n3732 12.1094
R11505 gnd.n3810 gnd.n2331 12.1094
R11506 gnd.n3898 gnd.n3897 12.1094
R11507 gnd.n4093 gnd.t182 12.1094
R11508 gnd.n6380 gnd.n6379 12.0247
R11509 gnd.n6348 gnd.n6347 12.0247
R11510 gnd.n6316 gnd.n6315 12.0247
R11511 gnd.n6285 gnd.n6284 12.0247
R11512 gnd.n6253 gnd.n6252 12.0247
R11513 gnd.n6221 gnd.n6220 12.0247
R11514 gnd.n6189 gnd.n6188 12.0247
R11515 gnd.n6158 gnd.n6157 12.0247
R11516 gnd.n4978 gnd.t262 11.7908
R11517 gnd.t219 gnd.n1359 11.7908
R11518 gnd.n1797 gnd.t236 11.7908
R11519 gnd.t295 gnd.n256 11.7908
R11520 gnd.n4829 gnd.n1423 11.4721
R11521 gnd.t139 gnd.n3559 11.4721
R11522 gnd.n3608 gnd.n2468 11.4721
R11523 gnd.t53 gnd.n2450 11.4721
R11524 gnd.n3631 gnd.n3630 11.4721
R11525 gnd.n3786 gnd.n2370 11.4721
R11526 gnd.n3828 gnd.n2358 11.4721
R11527 gnd.n3951 gnd.n3950 11.4721
R11528 gnd.n3958 gnd.t23 11.4721
R11529 gnd.n3967 gnd.n2251 11.4721
R11530 gnd.n4616 gnd.n1624 11.4721
R11531 gnd.n6383 gnd.n6370 11.249
R11532 gnd.n6351 gnd.n6338 11.249
R11533 gnd.n6319 gnd.n6306 11.249
R11534 gnd.n6288 gnd.n6275 11.249
R11535 gnd.n6256 gnd.n6243 11.249
R11536 gnd.n6224 gnd.n6211 11.249
R11537 gnd.n6192 gnd.n6179 11.249
R11538 gnd.n6161 gnd.n6148 11.249
R11539 gnd.n5832 gnd.t74 11.1535
R11540 gnd.n4954 gnd.t245 11.1535
R11541 gnd.t238 gnd.n1317 11.1535
R11542 gnd.n3413 gnd.t25 11.1535
R11543 gnd.t19 gnd.n2008 11.1535
R11544 gnd.n4422 gnd.t270 11.1535
R11545 gnd.n4511 gnd.t260 11.1535
R11546 gnd.n3674 gnd.n3673 10.8348
R11547 gnd.n3870 gnd.n2326 10.8348
R11548 gnd.n4159 gnd.n4158 10.6151
R11549 gnd.n4158 gnd.n4155 10.6151
R11550 gnd.n4153 gnd.n4150 10.6151
R11551 gnd.n4150 gnd.n4149 10.6151
R11552 gnd.n4149 gnd.n4146 10.6151
R11553 gnd.n4146 gnd.n4145 10.6151
R11554 gnd.n4145 gnd.n4142 10.6151
R11555 gnd.n4142 gnd.n4141 10.6151
R11556 gnd.n4141 gnd.n4138 10.6151
R11557 gnd.n4138 gnd.n4137 10.6151
R11558 gnd.n4137 gnd.n4134 10.6151
R11559 gnd.n4134 gnd.n4133 10.6151
R11560 gnd.n4133 gnd.n4130 10.6151
R11561 gnd.n4130 gnd.n4129 10.6151
R11562 gnd.n4129 gnd.n4126 10.6151
R11563 gnd.n4126 gnd.n4125 10.6151
R11564 gnd.n4125 gnd.n4122 10.6151
R11565 gnd.n4122 gnd.n4121 10.6151
R11566 gnd.n4121 gnd.n4118 10.6151
R11567 gnd.n4118 gnd.n4117 10.6151
R11568 gnd.n4117 gnd.n4114 10.6151
R11569 gnd.n4114 gnd.n4113 10.6151
R11570 gnd.n4113 gnd.n4110 10.6151
R11571 gnd.n4110 gnd.n4109 10.6151
R11572 gnd.n4109 gnd.n4106 10.6151
R11573 gnd.n4106 gnd.n4105 10.6151
R11574 gnd.n4105 gnd.n4102 10.6151
R11575 gnd.n4102 gnd.n4101 10.6151
R11576 gnd.n4101 gnd.n4098 10.6151
R11577 gnd.n4098 gnd.n4097 10.6151
R11578 gnd.n3547 gnd.n3546 10.6151
R11579 gnd.n3546 gnd.n2483 10.6151
R11580 gnd.n3563 gnd.n2483 10.6151
R11581 gnd.n3564 gnd.n3563 10.6151
R11582 gnd.n3582 gnd.n3564 10.6151
R11583 gnd.n3582 gnd.n3581 10.6151
R11584 gnd.n3581 gnd.n3580 10.6151
R11585 gnd.n3580 gnd.n3578 10.6151
R11586 gnd.n3578 gnd.n3577 10.6151
R11587 gnd.n3577 gnd.n3575 10.6151
R11588 gnd.n3575 gnd.n3574 10.6151
R11589 gnd.n3574 gnd.n3573 10.6151
R11590 gnd.n3573 gnd.n3572 10.6151
R11591 gnd.n3572 gnd.n3571 10.6151
R11592 gnd.n3571 gnd.n3568 10.6151
R11593 gnd.n3568 gnd.n3567 10.6151
R11594 gnd.n3567 gnd.n3565 10.6151
R11595 gnd.n3565 gnd.n2417 10.6151
R11596 gnd.n3683 gnd.n2417 10.6151
R11597 gnd.n3684 gnd.n3683 10.6151
R11598 gnd.n3686 gnd.n3684 10.6151
R11599 gnd.n3686 gnd.n3685 10.6151
R11600 gnd.n3685 gnd.n2400 10.6151
R11601 gnd.n3711 gnd.n2400 10.6151
R11602 gnd.n3712 gnd.n3711 10.6151
R11603 gnd.n3730 gnd.n3712 10.6151
R11604 gnd.n3730 gnd.n3729 10.6151
R11605 gnd.n3729 gnd.n3728 10.6151
R11606 gnd.n3728 gnd.n3713 10.6151
R11607 gnd.n3721 gnd.n3713 10.6151
R11608 gnd.n3721 gnd.n3720 10.6151
R11609 gnd.n3720 gnd.n3719 10.6151
R11610 gnd.n3719 gnd.n3718 10.6151
R11611 gnd.n3718 gnd.n3717 10.6151
R11612 gnd.n3717 gnd.n2361 10.6151
R11613 gnd.n3798 gnd.n2361 10.6151
R11614 gnd.n3799 gnd.n3798 10.6151
R11615 gnd.n3822 gnd.n3799 10.6151
R11616 gnd.n3822 gnd.n3821 10.6151
R11617 gnd.n3821 gnd.n3820 10.6151
R11618 gnd.n3820 gnd.n3816 10.6151
R11619 gnd.n3816 gnd.n3815 10.6151
R11620 gnd.n3815 gnd.n3813 10.6151
R11621 gnd.n3813 gnd.n3812 10.6151
R11622 gnd.n3812 gnd.n3807 10.6151
R11623 gnd.n3807 gnd.n3806 10.6151
R11624 gnd.n3806 gnd.n3804 10.6151
R11625 gnd.n3804 gnd.n3803 10.6151
R11626 gnd.n3803 gnd.n3800 10.6151
R11627 gnd.n3800 gnd.n2295 10.6151
R11628 gnd.n3895 gnd.n2295 10.6151
R11629 gnd.n3895 gnd.n3894 10.6151
R11630 gnd.n3894 gnd.n3893 10.6151
R11631 gnd.n3893 gnd.n2311 10.6151
R11632 gnd.n2311 gnd.n2310 10.6151
R11633 gnd.n2310 gnd.n2308 10.6151
R11634 gnd.n2308 gnd.n2307 10.6151
R11635 gnd.n2307 gnd.n2303 10.6151
R11636 gnd.n2303 gnd.n2302 10.6151
R11637 gnd.n2302 gnd.n2300 10.6151
R11638 gnd.n2300 gnd.n2299 10.6151
R11639 gnd.n2299 gnd.n2296 10.6151
R11640 gnd.n2296 gnd.n2242 10.6151
R11641 gnd.n3976 gnd.n2242 10.6151
R11642 gnd.n3977 gnd.n3976 10.6151
R11643 gnd.n3980 gnd.n3977 10.6151
R11644 gnd.n3980 gnd.n3979 10.6151
R11645 gnd.n3979 gnd.n3978 10.6151
R11646 gnd.n3978 gnd.n2224 10.6151
R11647 gnd.n2224 gnd.n2222 10.6151
R11648 gnd.n3484 gnd.n1462 10.6151
R11649 gnd.n3487 gnd.n3484 10.6151
R11650 gnd.n3492 gnd.n3489 10.6151
R11651 gnd.n3493 gnd.n3492 10.6151
R11652 gnd.n3496 gnd.n3493 10.6151
R11653 gnd.n3497 gnd.n3496 10.6151
R11654 gnd.n3500 gnd.n3497 10.6151
R11655 gnd.n3501 gnd.n3500 10.6151
R11656 gnd.n3504 gnd.n3501 10.6151
R11657 gnd.n3505 gnd.n3504 10.6151
R11658 gnd.n3508 gnd.n3505 10.6151
R11659 gnd.n3509 gnd.n3508 10.6151
R11660 gnd.n3512 gnd.n3509 10.6151
R11661 gnd.n3513 gnd.n3512 10.6151
R11662 gnd.n3516 gnd.n3513 10.6151
R11663 gnd.n3517 gnd.n3516 10.6151
R11664 gnd.n3520 gnd.n3517 10.6151
R11665 gnd.n3521 gnd.n3520 10.6151
R11666 gnd.n3524 gnd.n3521 10.6151
R11667 gnd.n3525 gnd.n3524 10.6151
R11668 gnd.n3528 gnd.n3525 10.6151
R11669 gnd.n3529 gnd.n3528 10.6151
R11670 gnd.n3532 gnd.n3529 10.6151
R11671 gnd.n3533 gnd.n3532 10.6151
R11672 gnd.n3536 gnd.n3533 10.6151
R11673 gnd.n3537 gnd.n3536 10.6151
R11674 gnd.n3540 gnd.n3537 10.6151
R11675 gnd.n3541 gnd.n3540 10.6151
R11676 gnd.n3544 gnd.n3541 10.6151
R11677 gnd.n3545 gnd.n3544 10.6151
R11678 gnd.n4793 gnd.n4792 10.6151
R11679 gnd.n4792 gnd.n4791 10.6151
R11680 gnd.n4791 gnd.n4790 10.6151
R11681 gnd.n4790 gnd.n4788 10.6151
R11682 gnd.n4788 gnd.n4785 10.6151
R11683 gnd.n4785 gnd.n4784 10.6151
R11684 gnd.n4784 gnd.n4781 10.6151
R11685 gnd.n4781 gnd.n4780 10.6151
R11686 gnd.n4780 gnd.n4777 10.6151
R11687 gnd.n4777 gnd.n4776 10.6151
R11688 gnd.n4776 gnd.n4773 10.6151
R11689 gnd.n4773 gnd.n4772 10.6151
R11690 gnd.n4772 gnd.n4769 10.6151
R11691 gnd.n4769 gnd.n4768 10.6151
R11692 gnd.n4768 gnd.n4765 10.6151
R11693 gnd.n4765 gnd.n4764 10.6151
R11694 gnd.n4764 gnd.n4761 10.6151
R11695 gnd.n4761 gnd.n4760 10.6151
R11696 gnd.n4760 gnd.n4757 10.6151
R11697 gnd.n4757 gnd.n4756 10.6151
R11698 gnd.n4756 gnd.n4753 10.6151
R11699 gnd.n4753 gnd.n4752 10.6151
R11700 gnd.n4752 gnd.n4749 10.6151
R11701 gnd.n4749 gnd.n4748 10.6151
R11702 gnd.n4748 gnd.n4745 10.6151
R11703 gnd.n4745 gnd.n4744 10.6151
R11704 gnd.n4744 gnd.n4741 10.6151
R11705 gnd.n4741 gnd.n4740 10.6151
R11706 gnd.n4737 gnd.n4736 10.6151
R11707 gnd.n4736 gnd.n1463 10.6151
R11708 gnd.n4088 gnd.n4086 10.6151
R11709 gnd.n4086 gnd.n4083 10.6151
R11710 gnd.n4083 gnd.n4082 10.6151
R11711 gnd.n4082 gnd.n4079 10.6151
R11712 gnd.n4079 gnd.n4078 10.6151
R11713 gnd.n4078 gnd.n4075 10.6151
R11714 gnd.n4075 gnd.n4074 10.6151
R11715 gnd.n4074 gnd.n4071 10.6151
R11716 gnd.n4071 gnd.n4070 10.6151
R11717 gnd.n4070 gnd.n4067 10.6151
R11718 gnd.n4067 gnd.n4066 10.6151
R11719 gnd.n4066 gnd.n4063 10.6151
R11720 gnd.n4063 gnd.n4062 10.6151
R11721 gnd.n4062 gnd.n4059 10.6151
R11722 gnd.n4059 gnd.n4058 10.6151
R11723 gnd.n4058 gnd.n4055 10.6151
R11724 gnd.n4055 gnd.n4054 10.6151
R11725 gnd.n4054 gnd.n4051 10.6151
R11726 gnd.n4051 gnd.n4050 10.6151
R11727 gnd.n4050 gnd.n4047 10.6151
R11728 gnd.n4047 gnd.n4046 10.6151
R11729 gnd.n4046 gnd.n4043 10.6151
R11730 gnd.n4043 gnd.n4042 10.6151
R11731 gnd.n4042 gnd.n4039 10.6151
R11732 gnd.n4039 gnd.n4038 10.6151
R11733 gnd.n4038 gnd.n4035 10.6151
R11734 gnd.n4035 gnd.n4034 10.6151
R11735 gnd.n4034 gnd.n4031 10.6151
R11736 gnd.n4029 gnd.n4026 10.6151
R11737 gnd.n4026 gnd.n4025 10.6151
R11738 gnd.n4729 gnd.n4728 10.6151
R11739 gnd.n4728 gnd.n1521 10.6151
R11740 gnd.n3588 gnd.n1521 10.6151
R11741 gnd.n3589 gnd.n3588 10.6151
R11742 gnd.n3589 gnd.n2471 10.6151
R11743 gnd.n3603 gnd.n2471 10.6151
R11744 gnd.n3604 gnd.n3603 10.6151
R11745 gnd.n3606 gnd.n3604 10.6151
R11746 gnd.n3606 gnd.n3605 10.6151
R11747 gnd.n3605 gnd.n2448 10.6151
R11748 gnd.n3634 gnd.n2448 10.6151
R11749 gnd.n3635 gnd.n3634 10.6151
R11750 gnd.n3636 gnd.n3635 10.6151
R11751 gnd.n3636 gnd.n2433 10.6151
R11752 gnd.n3655 gnd.n2433 10.6151
R11753 gnd.n3656 gnd.n3655 10.6151
R11754 gnd.n3658 gnd.n3656 10.6151
R11755 gnd.n3658 gnd.n3657 10.6151
R11756 gnd.n3657 gnd.n2414 10.6151
R11757 gnd.n3693 gnd.n2414 10.6151
R11758 gnd.n3694 gnd.n3693 10.6151
R11759 gnd.n3696 gnd.n3694 10.6151
R11760 gnd.n3696 gnd.n3695 10.6151
R11761 gnd.n3695 gnd.n2397 10.6151
R11762 gnd.n3736 gnd.n2397 10.6151
R11763 gnd.n3737 gnd.n3736 10.6151
R11764 gnd.n3741 gnd.n3737 10.6151
R11765 gnd.n3741 gnd.n3740 10.6151
R11766 gnd.n3740 gnd.n3739 10.6151
R11767 gnd.n3739 gnd.n2373 10.6151
R11768 gnd.n3779 gnd.n2373 10.6151
R11769 gnd.n3780 gnd.n3779 10.6151
R11770 gnd.n3784 gnd.n3780 10.6151
R11771 gnd.n3784 gnd.n3783 10.6151
R11772 gnd.n3783 gnd.n3782 10.6151
R11773 gnd.n3782 gnd.n2356 10.6151
R11774 gnd.n3830 gnd.n2356 10.6151
R11775 gnd.n3831 gnd.n3830 10.6151
R11776 gnd.n3832 gnd.n3831 10.6151
R11777 gnd.n3832 gnd.n2343 10.6151
R11778 gnd.n3848 gnd.n2343 10.6151
R11779 gnd.n3849 gnd.n3848 10.6151
R11780 gnd.n3850 gnd.n3849 10.6151
R11781 gnd.n3850 gnd.n2329 10.6151
R11782 gnd.n3865 gnd.n2329 10.6151
R11783 gnd.n3866 gnd.n3865 10.6151
R11784 gnd.n3868 gnd.n3866 10.6151
R11785 gnd.n3868 gnd.n3867 10.6151
R11786 gnd.n3867 gnd.n2290 10.6151
R11787 gnd.n3901 gnd.n2290 10.6151
R11788 gnd.n3902 gnd.n3901 10.6151
R11789 gnd.n3903 gnd.n3902 10.6151
R11790 gnd.n3903 gnd.n2277 10.6151
R11791 gnd.n3920 gnd.n2277 10.6151
R11792 gnd.n3921 gnd.n3920 10.6151
R11793 gnd.n3922 gnd.n3921 10.6151
R11794 gnd.n3922 gnd.n2263 10.6151
R11795 gnd.n3953 gnd.n2263 10.6151
R11796 gnd.n3954 gnd.n3953 10.6151
R11797 gnd.n3955 gnd.n3954 10.6151
R11798 gnd.n3955 gnd.n2248 10.6151
R11799 gnd.n3969 gnd.n2248 10.6151
R11800 gnd.n3970 gnd.n3969 10.6151
R11801 gnd.n3972 gnd.n3970 10.6151
R11802 gnd.n3972 gnd.n3971 10.6151
R11803 gnd.n3971 gnd.n2228 10.6151
R11804 gnd.n4000 gnd.n2228 10.6151
R11805 gnd.n4001 gnd.n4000 10.6151
R11806 gnd.n4091 gnd.n4001 10.6151
R11807 gnd.n4091 gnd.n4090 10.6151
R11808 gnd.n5504 gnd.t55 10.5161
R11809 gnd.t57 gnd.n5195 10.5161
R11810 gnd.n6136 gnd.t13 10.5161
R11811 gnd.n4928 gnd.t231 10.5161
R11812 gnd.t251 gnd.n1275 10.5161
R11813 gnd.n4469 gnd.t289 10.5161
R11814 gnd.n4547 gnd.t221 10.5161
R11815 gnd.n6384 gnd.n6368 10.4732
R11816 gnd.n6352 gnd.n6336 10.4732
R11817 gnd.n6320 gnd.n6304 10.4732
R11818 gnd.n6289 gnd.n6273 10.4732
R11819 gnd.n6257 gnd.n6241 10.4732
R11820 gnd.n6225 gnd.n6209 10.4732
R11821 gnd.n6193 gnd.n6177 10.4732
R11822 gnd.n6162 gnd.n6146 10.4732
R11823 gnd.n2468 gnd.n2459 10.1975
R11824 gnd.n2431 gnd.t52 10.1975
R11825 gnd.n3715 gnd.n2370 10.1975
R11826 gnd.n3796 gnd.n2358 10.1975
R11827 gnd.n3905 gnd.t76 10.1975
R11828 gnd.n2297 gnd.n2251 10.1975
R11829 gnd.n6057 gnd.t15 9.87883
R11830 gnd.t211 gnd.n1239 9.87883
R11831 gnd.n4903 gnd.t213 9.87883
R11832 gnd.n4439 gnd.t227 9.87883
R11833 gnd.t302 gnd.n4521 9.87883
R11834 gnd.n7720 gnd.n74 9.81789
R11835 gnd.n6388 gnd.n6387 9.69747
R11836 gnd.n6356 gnd.n6355 9.69747
R11837 gnd.n6324 gnd.n6323 9.69747
R11838 gnd.n6293 gnd.n6292 9.69747
R11839 gnd.n6261 gnd.n6260 9.69747
R11840 gnd.n6229 gnd.n6228 9.69747
R11841 gnd.n6197 gnd.n6196 9.69747
R11842 gnd.n6166 gnd.n6165 9.69747
R11843 gnd.n3549 gnd.n1523 9.56018
R11844 gnd.n3629 gnd.t40 9.56018
R11845 gnd.n3734 gnd.n3733 9.56018
R11846 gnd.n3863 gnd.n2331 9.56018
R11847 gnd.t50 gnd.n2265 9.56018
R11848 gnd.t182 gnd.n2043 9.56018
R11849 gnd.n3376 gnd.n3375 9.45599
R11850 gnd.n1886 gnd.n1878 9.45599
R11851 gnd.n6394 gnd.n6393 9.45567
R11852 gnd.n6362 gnd.n6361 9.45567
R11853 gnd.n6330 gnd.n6329 9.45567
R11854 gnd.n6299 gnd.n6298 9.45567
R11855 gnd.n6267 gnd.n6266 9.45567
R11856 gnd.n6235 gnd.n6234 9.45567
R11857 gnd.n6203 gnd.n6202 9.45567
R11858 gnd.n6172 gnd.n6171 9.45567
R11859 gnd.n5348 gnd.n5347 9.39724
R11860 gnd.n6393 gnd.n6392 9.3005
R11861 gnd.n6366 gnd.n6365 9.3005
R11862 gnd.n6387 gnd.n6386 9.3005
R11863 gnd.n6385 gnd.n6384 9.3005
R11864 gnd.n6370 gnd.n6369 9.3005
R11865 gnd.n6379 gnd.n6378 9.3005
R11866 gnd.n6377 gnd.n6376 9.3005
R11867 gnd.n6361 gnd.n6360 9.3005
R11868 gnd.n6334 gnd.n6333 9.3005
R11869 gnd.n6355 gnd.n6354 9.3005
R11870 gnd.n6353 gnd.n6352 9.3005
R11871 gnd.n6338 gnd.n6337 9.3005
R11872 gnd.n6347 gnd.n6346 9.3005
R11873 gnd.n6345 gnd.n6344 9.3005
R11874 gnd.n6329 gnd.n6328 9.3005
R11875 gnd.n6302 gnd.n6301 9.3005
R11876 gnd.n6323 gnd.n6322 9.3005
R11877 gnd.n6321 gnd.n6320 9.3005
R11878 gnd.n6306 gnd.n6305 9.3005
R11879 gnd.n6315 gnd.n6314 9.3005
R11880 gnd.n6313 gnd.n6312 9.3005
R11881 gnd.n6298 gnd.n6297 9.3005
R11882 gnd.n6271 gnd.n6270 9.3005
R11883 gnd.n6292 gnd.n6291 9.3005
R11884 gnd.n6290 gnd.n6289 9.3005
R11885 gnd.n6275 gnd.n6274 9.3005
R11886 gnd.n6284 gnd.n6283 9.3005
R11887 gnd.n6282 gnd.n6281 9.3005
R11888 gnd.n6266 gnd.n6265 9.3005
R11889 gnd.n6239 gnd.n6238 9.3005
R11890 gnd.n6260 gnd.n6259 9.3005
R11891 gnd.n6258 gnd.n6257 9.3005
R11892 gnd.n6243 gnd.n6242 9.3005
R11893 gnd.n6252 gnd.n6251 9.3005
R11894 gnd.n6250 gnd.n6249 9.3005
R11895 gnd.n6234 gnd.n6233 9.3005
R11896 gnd.n6207 gnd.n6206 9.3005
R11897 gnd.n6228 gnd.n6227 9.3005
R11898 gnd.n6226 gnd.n6225 9.3005
R11899 gnd.n6211 gnd.n6210 9.3005
R11900 gnd.n6220 gnd.n6219 9.3005
R11901 gnd.n6218 gnd.n6217 9.3005
R11902 gnd.n6202 gnd.n6201 9.3005
R11903 gnd.n6175 gnd.n6174 9.3005
R11904 gnd.n6196 gnd.n6195 9.3005
R11905 gnd.n6194 gnd.n6193 9.3005
R11906 gnd.n6179 gnd.n6178 9.3005
R11907 gnd.n6188 gnd.n6187 9.3005
R11908 gnd.n6186 gnd.n6185 9.3005
R11909 gnd.n6171 gnd.n6170 9.3005
R11910 gnd.n6144 gnd.n6143 9.3005
R11911 gnd.n6165 gnd.n6164 9.3005
R11912 gnd.n6163 gnd.n6162 9.3005
R11913 gnd.n6148 gnd.n6147 9.3005
R11914 gnd.n6157 gnd.n6156 9.3005
R11915 gnd.n6155 gnd.n6154 9.3005
R11916 gnd.n5120 gnd.n5117 9.3005
R11917 gnd.n6508 gnd.n5121 9.3005
R11918 gnd.n6507 gnd.n5122 9.3005
R11919 gnd.n6506 gnd.n5123 9.3005
R11920 gnd.n6503 gnd.n5124 9.3005
R11921 gnd.n6502 gnd.n5125 9.3005
R11922 gnd.n6499 gnd.n5126 9.3005
R11923 gnd.n6498 gnd.n5127 9.3005
R11924 gnd.n6495 gnd.n5128 9.3005
R11925 gnd.n6494 gnd.n5129 9.3005
R11926 gnd.n6491 gnd.n5130 9.3005
R11927 gnd.n6490 gnd.n5131 9.3005
R11928 gnd.n6487 gnd.n5132 9.3005
R11929 gnd.n6486 gnd.n5133 9.3005
R11930 gnd.n6483 gnd.n6482 9.3005
R11931 gnd.n6481 gnd.n5135 9.3005
R11932 gnd.n5119 gnd.n5118 9.3005
R11933 gnd.n5771 gnd.n5770 9.3005
R11934 gnd.n5772 gnd.n5474 9.3005
R11935 gnd.n5774 gnd.n5773 9.3005
R11936 gnd.n5455 gnd.n5454 9.3005
R11937 gnd.n5801 gnd.n5800 9.3005
R11938 gnd.n5802 gnd.n5453 9.3005
R11939 gnd.n5806 gnd.n5803 9.3005
R11940 gnd.n5805 gnd.n5804 9.3005
R11941 gnd.n5429 gnd.n5428 9.3005
R11942 gnd.n5835 gnd.n5834 9.3005
R11943 gnd.n5836 gnd.n5427 9.3005
R11944 gnd.n5843 gnd.n5837 9.3005
R11945 gnd.n5842 gnd.n5838 9.3005
R11946 gnd.n5841 gnd.n5839 9.3005
R11947 gnd.n5396 gnd.n5395 9.3005
R11948 gnd.n5896 gnd.n5895 9.3005
R11949 gnd.n5897 gnd.n5394 9.3005
R11950 gnd.n5901 gnd.n5898 9.3005
R11951 gnd.n5900 gnd.n5899 9.3005
R11952 gnd.n5369 gnd.n5368 9.3005
R11953 gnd.n5936 gnd.n5935 9.3005
R11954 gnd.n5937 gnd.n5367 9.3005
R11955 gnd.n5941 gnd.n5938 9.3005
R11956 gnd.n5940 gnd.n5939 9.3005
R11957 gnd.n5282 gnd.n5281 9.3005
R11958 gnd.n5981 gnd.n5980 9.3005
R11959 gnd.n5982 gnd.n5280 9.3005
R11960 gnd.n5986 gnd.n5983 9.3005
R11961 gnd.n5985 gnd.n5984 9.3005
R11962 gnd.n5254 gnd.n5253 9.3005
R11963 gnd.n6021 gnd.n6020 9.3005
R11964 gnd.n6022 gnd.n5252 9.3005
R11965 gnd.n6026 gnd.n6023 9.3005
R11966 gnd.n6025 gnd.n6024 9.3005
R11967 gnd.n5227 gnd.n5226 9.3005
R11968 gnd.n6067 gnd.n6066 9.3005
R11969 gnd.n6068 gnd.n5225 9.3005
R11970 gnd.n6072 gnd.n6069 9.3005
R11971 gnd.n6071 gnd.n6070 9.3005
R11972 gnd.n5200 gnd.n5199 9.3005
R11973 gnd.n6106 gnd.n6105 9.3005
R11974 gnd.n6107 gnd.n5198 9.3005
R11975 gnd.n6112 gnd.n6108 9.3005
R11976 gnd.n6111 gnd.n6110 9.3005
R11977 gnd.n6109 gnd.n967 9.3005
R11978 gnd.n6530 gnd.n968 9.3005
R11979 gnd.n6529 gnd.n969 9.3005
R11980 gnd.n6528 gnd.n970 9.3005
R11981 gnd.n990 gnd.n971 9.3005
R11982 gnd.n991 gnd.n989 9.3005
R11983 gnd.n6516 gnd.n992 9.3005
R11984 gnd.n6515 gnd.n993 9.3005
R11985 gnd.n6514 gnd.n994 9.3005
R11986 gnd.n5476 gnd.n5475 9.3005
R11987 gnd.n5716 gnd.n5715 9.3005
R11988 gnd.n5719 gnd.n5711 9.3005
R11989 gnd.n5720 gnd.n5710 9.3005
R11990 gnd.n5723 gnd.n5709 9.3005
R11991 gnd.n5724 gnd.n5708 9.3005
R11992 gnd.n5727 gnd.n5707 9.3005
R11993 gnd.n5728 gnd.n5706 9.3005
R11994 gnd.n5731 gnd.n5705 9.3005
R11995 gnd.n5732 gnd.n5704 9.3005
R11996 gnd.n5735 gnd.n5703 9.3005
R11997 gnd.n5736 gnd.n5702 9.3005
R11998 gnd.n5739 gnd.n5701 9.3005
R11999 gnd.n5741 gnd.n5700 9.3005
R12000 gnd.n5742 gnd.n5699 9.3005
R12001 gnd.n5743 gnd.n5698 9.3005
R12002 gnd.n5744 gnd.n5697 9.3005
R12003 gnd.n5712 gnd.n5493 9.3005
R12004 gnd.n5761 gnd.n5484 9.3005
R12005 gnd.n5763 gnd.n5762 9.3005
R12006 gnd.n5471 gnd.n5466 9.3005
R12007 gnd.n5784 gnd.n5465 9.3005
R12008 gnd.n5787 gnd.n5786 9.3005
R12009 gnd.n5789 gnd.n5788 9.3005
R12010 gnd.n5792 gnd.n5448 9.3005
R12011 gnd.n5790 gnd.n5446 9.3005
R12012 gnd.n5812 gnd.n5444 9.3005
R12013 gnd.n5816 gnd.n5815 9.3005
R12014 gnd.n5814 gnd.n5419 9.3005
R12015 gnd.n5850 gnd.n5418 9.3005
R12016 gnd.n5853 gnd.n5852 9.3005
R12017 gnd.n5416 gnd.n5415 9.3005
R12018 gnd.n5859 gnd.n5413 9.3005
R12019 gnd.n5861 gnd.n5860 9.3005
R12020 gnd.n5387 gnd.n5386 9.3005
R12021 gnd.n5910 gnd.n5909 9.3005
R12022 gnd.n5911 gnd.n5380 9.3005
R12023 gnd.n5919 gnd.n5379 9.3005
R12024 gnd.n5922 gnd.n5921 9.3005
R12025 gnd.n5924 gnd.n5923 9.3005
R12026 gnd.n5927 gnd.n5362 9.3005
R12027 gnd.n5925 gnd.n5360 9.3005
R12028 gnd.n5947 gnd.n5358 9.3005
R12029 gnd.n5949 gnd.n5948 9.3005
R12030 gnd.n5272 gnd.n5271 9.3005
R12031 gnd.n5995 gnd.n5994 9.3005
R12032 gnd.n5996 gnd.n5265 9.3005
R12033 gnd.n6004 gnd.n5264 9.3005
R12034 gnd.n6007 gnd.n6006 9.3005
R12035 gnd.n6009 gnd.n6008 9.3005
R12036 gnd.n6012 gnd.n5247 9.3005
R12037 gnd.n6010 gnd.n5245 9.3005
R12038 gnd.n6032 gnd.n5243 9.3005
R12039 gnd.n6034 gnd.n6033 9.3005
R12040 gnd.n5218 gnd.n5217 9.3005
R12041 gnd.n6081 gnd.n6080 9.3005
R12042 gnd.n6082 gnd.n5211 9.3005
R12043 gnd.n6090 gnd.n5210 9.3005
R12044 gnd.n6093 gnd.n6092 9.3005
R12045 gnd.n6095 gnd.n6094 9.3005
R12046 gnd.n6097 gnd.n5193 9.3005
R12047 gnd.n5190 gnd.n5188 9.3005
R12048 gnd.n6119 gnd.n6118 9.3005
R12049 gnd.n5191 gnd.n5175 9.3005
R12050 gnd.n6140 gnd.n5174 9.3005
R12051 gnd.n6399 gnd.n6398 9.3005
R12052 gnd.n6401 gnd.n6400 9.3005
R12053 gnd.n6415 gnd.n6402 9.3005
R12054 gnd.n6414 gnd.n6403 9.3005
R12055 gnd.n6413 gnd.n6408 9.3005
R12056 gnd.n6409 gnd.n5138 9.3005
R12057 gnd.n5760 gnd.n5487 9.3005
R12058 gnd.n6477 gnd.n5139 9.3005
R12059 gnd.n6476 gnd.n5141 9.3005
R12060 gnd.n6473 gnd.n5142 9.3005
R12061 gnd.n6472 gnd.n5143 9.3005
R12062 gnd.n6469 gnd.n5144 9.3005
R12063 gnd.n6468 gnd.n5145 9.3005
R12064 gnd.n6465 gnd.n5146 9.3005
R12065 gnd.n6464 gnd.n5147 9.3005
R12066 gnd.n6461 gnd.n5148 9.3005
R12067 gnd.n6460 gnd.n5149 9.3005
R12068 gnd.n6457 gnd.n5150 9.3005
R12069 gnd.n6456 gnd.n5151 9.3005
R12070 gnd.n6453 gnd.n5152 9.3005
R12071 gnd.n6452 gnd.n5153 9.3005
R12072 gnd.n6449 gnd.n5154 9.3005
R12073 gnd.n6448 gnd.n5155 9.3005
R12074 gnd.n6445 gnd.n5156 9.3005
R12075 gnd.n6444 gnd.n5157 9.3005
R12076 gnd.n6441 gnd.n5158 9.3005
R12077 gnd.n6440 gnd.n5159 9.3005
R12078 gnd.n6437 gnd.n5160 9.3005
R12079 gnd.n6436 gnd.n5161 9.3005
R12080 gnd.n6433 gnd.n5165 9.3005
R12081 gnd.n6432 gnd.n5166 9.3005
R12082 gnd.n6429 gnd.n5167 9.3005
R12083 gnd.n6428 gnd.n5168 9.3005
R12084 gnd.n6479 gnd.n6478 9.3005
R12085 gnd.n5957 gnd.n5956 9.3005
R12086 gnd.n5958 gnd.n5288 9.3005
R12087 gnd.n5975 gnd.n5959 9.3005
R12088 gnd.n5974 gnd.n5960 9.3005
R12089 gnd.n5973 gnd.n5961 9.3005
R12090 gnd.n5971 gnd.n5962 9.3005
R12091 gnd.n5970 gnd.n5963 9.3005
R12092 gnd.n5968 gnd.n5964 9.3005
R12093 gnd.n5967 gnd.n5965 9.3005
R12094 gnd.n5234 gnd.n5233 9.3005
R12095 gnd.n6042 gnd.n6041 9.3005
R12096 gnd.n6043 gnd.n5232 9.3005
R12097 gnd.n6061 gnd.n6044 9.3005
R12098 gnd.n6060 gnd.n6045 9.3005
R12099 gnd.n6059 gnd.n6046 9.3005
R12100 gnd.n6056 gnd.n6047 9.3005
R12101 gnd.n6055 gnd.n6048 9.3005
R12102 gnd.n6053 gnd.n6049 9.3005
R12103 gnd.n6052 gnd.n6050 9.3005
R12104 gnd.n5182 gnd.n5181 9.3005
R12105 gnd.n6126 gnd.n6125 9.3005
R12106 gnd.n6127 gnd.n5180 9.3005
R12107 gnd.n6132 gnd.n6128 9.3005
R12108 gnd.n6131 gnd.n6130 9.3005
R12109 gnd.n6129 gnd.n5172 9.3005
R12110 gnd.n6420 gnd.n5171 9.3005
R12111 gnd.n6422 gnd.n6421 9.3005
R12112 gnd.n6423 gnd.n5170 9.3005
R12113 gnd.n6425 gnd.n6424 9.3005
R12114 gnd.n5630 gnd.n5524 9.3005
R12115 gnd.n5632 gnd.n5631 9.3005
R12116 gnd.n5514 gnd.n5513 9.3005
R12117 gnd.n5645 gnd.n5644 9.3005
R12118 gnd.n5646 gnd.n5512 9.3005
R12119 gnd.n5648 gnd.n5647 9.3005
R12120 gnd.n5501 gnd.n5500 9.3005
R12121 gnd.n5661 gnd.n5660 9.3005
R12122 gnd.n5662 gnd.n5499 9.3005
R12123 gnd.n5686 gnd.n5663 9.3005
R12124 gnd.n5685 gnd.n5664 9.3005
R12125 gnd.n5684 gnd.n5665 9.3005
R12126 gnd.n5683 gnd.n5666 9.3005
R12127 gnd.n5681 gnd.n5667 9.3005
R12128 gnd.n5680 gnd.n5668 9.3005
R12129 gnd.n5678 gnd.n5669 9.3005
R12130 gnd.n5677 gnd.n5670 9.3005
R12131 gnd.n5675 gnd.n5671 9.3005
R12132 gnd.n5674 gnd.n5672 9.3005
R12133 gnd.n5436 gnd.n5435 9.3005
R12134 gnd.n5824 gnd.n5823 9.3005
R12135 gnd.n5825 gnd.n5434 9.3005
R12136 gnd.n5829 gnd.n5826 9.3005
R12137 gnd.n5828 gnd.n5827 9.3005
R12138 gnd.n5403 gnd.n5402 9.3005
R12139 gnd.n5871 gnd.n5870 9.3005
R12140 gnd.n5872 gnd.n5401 9.3005
R12141 gnd.n5874 gnd.n5873 9.3005
R12142 gnd.n5629 gnd.n5628 9.3005
R12143 gnd.n5569 gnd.n5568 9.3005
R12144 gnd.n5574 gnd.n5566 9.3005
R12145 gnd.n5575 gnd.n5565 9.3005
R12146 gnd.n5577 gnd.n5562 9.3005
R12147 gnd.n5561 gnd.n5559 9.3005
R12148 gnd.n5583 gnd.n5558 9.3005
R12149 gnd.n5584 gnd.n5557 9.3005
R12150 gnd.n5585 gnd.n5556 9.3005
R12151 gnd.n5555 gnd.n5553 9.3005
R12152 gnd.n5591 gnd.n5552 9.3005
R12153 gnd.n5592 gnd.n5551 9.3005
R12154 gnd.n5593 gnd.n5550 9.3005
R12155 gnd.n5549 gnd.n5547 9.3005
R12156 gnd.n5599 gnd.n5546 9.3005
R12157 gnd.n5600 gnd.n5545 9.3005
R12158 gnd.n5601 gnd.n5544 9.3005
R12159 gnd.n5543 gnd.n5541 9.3005
R12160 gnd.n5607 gnd.n5540 9.3005
R12161 gnd.n5608 gnd.n5539 9.3005
R12162 gnd.n5609 gnd.n5538 9.3005
R12163 gnd.n5537 gnd.n5535 9.3005
R12164 gnd.n5614 gnd.n5534 9.3005
R12165 gnd.n5615 gnd.n5533 9.3005
R12166 gnd.n5532 gnd.n5530 9.3005
R12167 gnd.n5620 gnd.n5529 9.3005
R12168 gnd.n5622 gnd.n5621 9.3005
R12169 gnd.n5567 gnd.n5525 9.3005
R12170 gnd.n5520 gnd.n5519 9.3005
R12171 gnd.n5637 gnd.n5636 9.3005
R12172 gnd.n5638 gnd.n5518 9.3005
R12173 gnd.n5640 gnd.n5639 9.3005
R12174 gnd.n5508 gnd.n5507 9.3005
R12175 gnd.n5653 gnd.n5652 9.3005
R12176 gnd.n5654 gnd.n5506 9.3005
R12177 gnd.n5656 gnd.n5655 9.3005
R12178 gnd.n5495 gnd.n5494 9.3005
R12179 gnd.n5751 gnd.n5750 9.3005
R12180 gnd.n5753 gnd.n5492 9.3005
R12181 gnd.n5755 gnd.n5754 9.3005
R12182 gnd.n5486 gnd.n5483 9.3005
R12183 gnd.n5765 gnd.n5764 9.3005
R12184 gnd.n5485 gnd.n5467 9.3005
R12185 gnd.n5783 gnd.n5782 9.3005
R12186 gnd.n5785 gnd.n5463 9.3005
R12187 gnd.n5795 gnd.n5464 9.3005
R12188 gnd.n5794 gnd.n5793 9.3005
R12189 gnd.n5791 gnd.n5442 9.3005
R12190 gnd.n5819 gnd.n5443 9.3005
R12191 gnd.n5818 gnd.n5817 9.3005
R12192 gnd.n5445 gnd.n5420 9.3005
R12193 gnd.n5849 gnd.n5848 9.3005
R12194 gnd.n5851 gnd.n5410 9.3005
R12195 gnd.n5866 gnd.n5411 9.3005
R12196 gnd.n5865 gnd.n5412 9.3005
R12197 gnd.n5864 gnd.n5862 9.3005
R12198 gnd.n5414 gnd.n5388 9.3005
R12199 gnd.n5907 gnd.n5906 9.3005
R12200 gnd.n5908 gnd.n5381 9.3005
R12201 gnd.n5918 gnd.n5917 9.3005
R12202 gnd.n5920 gnd.n5377 9.3005
R12203 gnd.n5930 gnd.n5378 9.3005
R12204 gnd.n5929 gnd.n5928 9.3005
R12205 gnd.n5926 gnd.n5356 9.3005
R12206 gnd.n5952 gnd.n5357 9.3005
R12207 gnd.n5951 gnd.n5950 9.3005
R12208 gnd.n5359 gnd.n5273 9.3005
R12209 gnd.n5992 gnd.n5991 9.3005
R12210 gnd.n5993 gnd.n5266 9.3005
R12211 gnd.n6003 gnd.n6002 9.3005
R12212 gnd.n6005 gnd.n5262 9.3005
R12213 gnd.n6015 gnd.n5263 9.3005
R12214 gnd.n6014 gnd.n6013 9.3005
R12215 gnd.n6011 gnd.n5241 9.3005
R12216 gnd.n6037 gnd.n5242 9.3005
R12217 gnd.n6036 gnd.n6035 9.3005
R12218 gnd.n5244 gnd.n5219 9.3005
R12219 gnd.n6078 gnd.n6077 9.3005
R12220 gnd.n6079 gnd.n5212 9.3005
R12221 gnd.n6089 gnd.n6088 9.3005
R12222 gnd.n6091 gnd.n5208 9.3005
R12223 gnd.n6100 gnd.n5209 9.3005
R12224 gnd.n6099 gnd.n6098 9.3005
R12225 gnd.n6096 gnd.n5187 9.3005
R12226 gnd.n6121 gnd.n6120 9.3005
R12227 gnd.n5189 gnd.n5176 9.3005
R12228 gnd.n6139 gnd.n6138 9.3005
R12229 gnd.n6141 gnd.n979 9.3005
R12230 gnd.n6523 gnd.n980 9.3005
R12231 gnd.n6522 gnd.n981 9.3005
R12232 gnd.n6521 gnd.n982 9.3005
R12233 gnd.n6404 gnd.n983 9.3005
R12234 gnd.n6407 gnd.n6406 9.3005
R12235 gnd.n5624 gnd.n5623 9.3005
R12236 gnd.n794 gnd.n793 9.3005
R12237 gnd.n6706 gnd.n6705 9.3005
R12238 gnd.n6707 gnd.n792 9.3005
R12239 gnd.n6709 gnd.n6708 9.3005
R12240 gnd.n788 gnd.n787 9.3005
R12241 gnd.n6716 gnd.n6715 9.3005
R12242 gnd.n6717 gnd.n786 9.3005
R12243 gnd.n6719 gnd.n6718 9.3005
R12244 gnd.n782 gnd.n781 9.3005
R12245 gnd.n6726 gnd.n6725 9.3005
R12246 gnd.n6727 gnd.n780 9.3005
R12247 gnd.n6729 gnd.n6728 9.3005
R12248 gnd.n776 gnd.n775 9.3005
R12249 gnd.n6736 gnd.n6735 9.3005
R12250 gnd.n6737 gnd.n774 9.3005
R12251 gnd.n6739 gnd.n6738 9.3005
R12252 gnd.n770 gnd.n769 9.3005
R12253 gnd.n6746 gnd.n6745 9.3005
R12254 gnd.n6747 gnd.n768 9.3005
R12255 gnd.n6749 gnd.n6748 9.3005
R12256 gnd.n764 gnd.n763 9.3005
R12257 gnd.n6756 gnd.n6755 9.3005
R12258 gnd.n6757 gnd.n762 9.3005
R12259 gnd.n6759 gnd.n6758 9.3005
R12260 gnd.n758 gnd.n757 9.3005
R12261 gnd.n6766 gnd.n6765 9.3005
R12262 gnd.n6767 gnd.n756 9.3005
R12263 gnd.n6769 gnd.n6768 9.3005
R12264 gnd.n752 gnd.n751 9.3005
R12265 gnd.n6776 gnd.n6775 9.3005
R12266 gnd.n6777 gnd.n750 9.3005
R12267 gnd.n6779 gnd.n6778 9.3005
R12268 gnd.n746 gnd.n745 9.3005
R12269 gnd.n6786 gnd.n6785 9.3005
R12270 gnd.n6787 gnd.n744 9.3005
R12271 gnd.n6789 gnd.n6788 9.3005
R12272 gnd.n740 gnd.n739 9.3005
R12273 gnd.n6796 gnd.n6795 9.3005
R12274 gnd.n6797 gnd.n738 9.3005
R12275 gnd.n6799 gnd.n6798 9.3005
R12276 gnd.n734 gnd.n733 9.3005
R12277 gnd.n6806 gnd.n6805 9.3005
R12278 gnd.n6807 gnd.n732 9.3005
R12279 gnd.n6809 gnd.n6808 9.3005
R12280 gnd.n728 gnd.n727 9.3005
R12281 gnd.n6816 gnd.n6815 9.3005
R12282 gnd.n6817 gnd.n726 9.3005
R12283 gnd.n6819 gnd.n6818 9.3005
R12284 gnd.n722 gnd.n721 9.3005
R12285 gnd.n6826 gnd.n6825 9.3005
R12286 gnd.n6827 gnd.n720 9.3005
R12287 gnd.n6829 gnd.n6828 9.3005
R12288 gnd.n716 gnd.n715 9.3005
R12289 gnd.n6836 gnd.n6835 9.3005
R12290 gnd.n6837 gnd.n714 9.3005
R12291 gnd.n6839 gnd.n6838 9.3005
R12292 gnd.n710 gnd.n709 9.3005
R12293 gnd.n6846 gnd.n6845 9.3005
R12294 gnd.n6847 gnd.n708 9.3005
R12295 gnd.n6849 gnd.n6848 9.3005
R12296 gnd.n704 gnd.n703 9.3005
R12297 gnd.n6856 gnd.n6855 9.3005
R12298 gnd.n6857 gnd.n702 9.3005
R12299 gnd.n6859 gnd.n6858 9.3005
R12300 gnd.n698 gnd.n697 9.3005
R12301 gnd.n6866 gnd.n6865 9.3005
R12302 gnd.n6867 gnd.n696 9.3005
R12303 gnd.n6869 gnd.n6868 9.3005
R12304 gnd.n692 gnd.n691 9.3005
R12305 gnd.n6876 gnd.n6875 9.3005
R12306 gnd.n6877 gnd.n690 9.3005
R12307 gnd.n6879 gnd.n6878 9.3005
R12308 gnd.n686 gnd.n685 9.3005
R12309 gnd.n6886 gnd.n6885 9.3005
R12310 gnd.n6887 gnd.n684 9.3005
R12311 gnd.n6889 gnd.n6888 9.3005
R12312 gnd.n680 gnd.n679 9.3005
R12313 gnd.n6896 gnd.n6895 9.3005
R12314 gnd.n6897 gnd.n678 9.3005
R12315 gnd.n6899 gnd.n6898 9.3005
R12316 gnd.n674 gnd.n673 9.3005
R12317 gnd.n6906 gnd.n6905 9.3005
R12318 gnd.n6907 gnd.n672 9.3005
R12319 gnd.n6909 gnd.n6908 9.3005
R12320 gnd.n668 gnd.n667 9.3005
R12321 gnd.n6916 gnd.n6915 9.3005
R12322 gnd.n6917 gnd.n666 9.3005
R12323 gnd.n6919 gnd.n6918 9.3005
R12324 gnd.n662 gnd.n661 9.3005
R12325 gnd.n6926 gnd.n6925 9.3005
R12326 gnd.n6927 gnd.n660 9.3005
R12327 gnd.n6929 gnd.n6928 9.3005
R12328 gnd.n656 gnd.n655 9.3005
R12329 gnd.n6936 gnd.n6935 9.3005
R12330 gnd.n6937 gnd.n654 9.3005
R12331 gnd.n6939 gnd.n6938 9.3005
R12332 gnd.n650 gnd.n649 9.3005
R12333 gnd.n6946 gnd.n6945 9.3005
R12334 gnd.n6947 gnd.n648 9.3005
R12335 gnd.n6949 gnd.n6948 9.3005
R12336 gnd.n644 gnd.n643 9.3005
R12337 gnd.n6956 gnd.n6955 9.3005
R12338 gnd.n6957 gnd.n642 9.3005
R12339 gnd.n6959 gnd.n6958 9.3005
R12340 gnd.n638 gnd.n637 9.3005
R12341 gnd.n6966 gnd.n6965 9.3005
R12342 gnd.n6967 gnd.n636 9.3005
R12343 gnd.n6969 gnd.n6968 9.3005
R12344 gnd.n632 gnd.n631 9.3005
R12345 gnd.n6976 gnd.n6975 9.3005
R12346 gnd.n6977 gnd.n630 9.3005
R12347 gnd.n6979 gnd.n6978 9.3005
R12348 gnd.n626 gnd.n625 9.3005
R12349 gnd.n6986 gnd.n6985 9.3005
R12350 gnd.n6987 gnd.n624 9.3005
R12351 gnd.n6989 gnd.n6988 9.3005
R12352 gnd.n620 gnd.n619 9.3005
R12353 gnd.n6996 gnd.n6995 9.3005
R12354 gnd.n6997 gnd.n618 9.3005
R12355 gnd.n6999 gnd.n6998 9.3005
R12356 gnd.n614 gnd.n613 9.3005
R12357 gnd.n7006 gnd.n7005 9.3005
R12358 gnd.n7007 gnd.n612 9.3005
R12359 gnd.n7009 gnd.n7008 9.3005
R12360 gnd.n608 gnd.n607 9.3005
R12361 gnd.n7016 gnd.n7015 9.3005
R12362 gnd.n7017 gnd.n606 9.3005
R12363 gnd.n7019 gnd.n7018 9.3005
R12364 gnd.n602 gnd.n601 9.3005
R12365 gnd.n7026 gnd.n7025 9.3005
R12366 gnd.n7027 gnd.n600 9.3005
R12367 gnd.n7029 gnd.n7028 9.3005
R12368 gnd.n596 gnd.n595 9.3005
R12369 gnd.n7036 gnd.n7035 9.3005
R12370 gnd.n7037 gnd.n594 9.3005
R12371 gnd.n7039 gnd.n7038 9.3005
R12372 gnd.n590 gnd.n589 9.3005
R12373 gnd.n7046 gnd.n7045 9.3005
R12374 gnd.n7047 gnd.n588 9.3005
R12375 gnd.n7049 gnd.n7048 9.3005
R12376 gnd.n584 gnd.n583 9.3005
R12377 gnd.n7056 gnd.n7055 9.3005
R12378 gnd.n7057 gnd.n582 9.3005
R12379 gnd.n7059 gnd.n7058 9.3005
R12380 gnd.n578 gnd.n577 9.3005
R12381 gnd.n7066 gnd.n7065 9.3005
R12382 gnd.n7067 gnd.n576 9.3005
R12383 gnd.n7069 gnd.n7068 9.3005
R12384 gnd.n572 gnd.n571 9.3005
R12385 gnd.n7076 gnd.n7075 9.3005
R12386 gnd.n7077 gnd.n570 9.3005
R12387 gnd.n7079 gnd.n7078 9.3005
R12388 gnd.n566 gnd.n565 9.3005
R12389 gnd.n7086 gnd.n7085 9.3005
R12390 gnd.n7087 gnd.n564 9.3005
R12391 gnd.n7089 gnd.n7088 9.3005
R12392 gnd.n560 gnd.n559 9.3005
R12393 gnd.n7096 gnd.n7095 9.3005
R12394 gnd.n7097 gnd.n558 9.3005
R12395 gnd.n7099 gnd.n7098 9.3005
R12396 gnd.n554 gnd.n553 9.3005
R12397 gnd.n7106 gnd.n7105 9.3005
R12398 gnd.n7107 gnd.n552 9.3005
R12399 gnd.n7109 gnd.n7108 9.3005
R12400 gnd.n548 gnd.n547 9.3005
R12401 gnd.n7116 gnd.n7115 9.3005
R12402 gnd.n7117 gnd.n546 9.3005
R12403 gnd.n7119 gnd.n7118 9.3005
R12404 gnd.n542 gnd.n541 9.3005
R12405 gnd.n7126 gnd.n7125 9.3005
R12406 gnd.n7127 gnd.n540 9.3005
R12407 gnd.n7129 gnd.n7128 9.3005
R12408 gnd.n536 gnd.n535 9.3005
R12409 gnd.n7136 gnd.n7135 9.3005
R12410 gnd.n7137 gnd.n534 9.3005
R12411 gnd.n7139 gnd.n7138 9.3005
R12412 gnd.n530 gnd.n529 9.3005
R12413 gnd.n7146 gnd.n7145 9.3005
R12414 gnd.n7147 gnd.n528 9.3005
R12415 gnd.n7149 gnd.n7148 9.3005
R12416 gnd.n524 gnd.n523 9.3005
R12417 gnd.n7156 gnd.n7155 9.3005
R12418 gnd.n7159 gnd.n7158 9.3005
R12419 gnd.n518 gnd.n517 9.3005
R12420 gnd.n7166 gnd.n7165 9.3005
R12421 gnd.n7167 gnd.n516 9.3005
R12422 gnd.n7169 gnd.n7168 9.3005
R12423 gnd.n512 gnd.n511 9.3005
R12424 gnd.n7176 gnd.n7175 9.3005
R12425 gnd.n7177 gnd.n510 9.3005
R12426 gnd.n7179 gnd.n7178 9.3005
R12427 gnd.n506 gnd.n505 9.3005
R12428 gnd.n7186 gnd.n7185 9.3005
R12429 gnd.n7187 gnd.n504 9.3005
R12430 gnd.n7189 gnd.n7188 9.3005
R12431 gnd.n500 gnd.n499 9.3005
R12432 gnd.n7196 gnd.n7195 9.3005
R12433 gnd.n7197 gnd.n498 9.3005
R12434 gnd.n7199 gnd.n7198 9.3005
R12435 gnd.n494 gnd.n493 9.3005
R12436 gnd.n7206 gnd.n7205 9.3005
R12437 gnd.n7207 gnd.n492 9.3005
R12438 gnd.n7209 gnd.n7208 9.3005
R12439 gnd.n488 gnd.n487 9.3005
R12440 gnd.n7216 gnd.n7215 9.3005
R12441 gnd.n7217 gnd.n486 9.3005
R12442 gnd.n7219 gnd.n7218 9.3005
R12443 gnd.n482 gnd.n481 9.3005
R12444 gnd.n7226 gnd.n7225 9.3005
R12445 gnd.n7227 gnd.n480 9.3005
R12446 gnd.n7229 gnd.n7228 9.3005
R12447 gnd.n476 gnd.n475 9.3005
R12448 gnd.n7236 gnd.n7235 9.3005
R12449 gnd.n7237 gnd.n474 9.3005
R12450 gnd.n7239 gnd.n7238 9.3005
R12451 gnd.n470 gnd.n469 9.3005
R12452 gnd.n7246 gnd.n7245 9.3005
R12453 gnd.n7247 gnd.n468 9.3005
R12454 gnd.n7249 gnd.n7248 9.3005
R12455 gnd.n464 gnd.n463 9.3005
R12456 gnd.n7256 gnd.n7255 9.3005
R12457 gnd.n7257 gnd.n462 9.3005
R12458 gnd.n7259 gnd.n7258 9.3005
R12459 gnd.n458 gnd.n457 9.3005
R12460 gnd.n7266 gnd.n7265 9.3005
R12461 gnd.n7267 gnd.n456 9.3005
R12462 gnd.n7269 gnd.n7268 9.3005
R12463 gnd.n452 gnd.n451 9.3005
R12464 gnd.n7276 gnd.n7275 9.3005
R12465 gnd.n7277 gnd.n450 9.3005
R12466 gnd.n7279 gnd.n7278 9.3005
R12467 gnd.n446 gnd.n445 9.3005
R12468 gnd.n7286 gnd.n7285 9.3005
R12469 gnd.n7287 gnd.n444 9.3005
R12470 gnd.n7289 gnd.n7288 9.3005
R12471 gnd.n440 gnd.n439 9.3005
R12472 gnd.n7296 gnd.n7295 9.3005
R12473 gnd.n7297 gnd.n438 9.3005
R12474 gnd.n7299 gnd.n7298 9.3005
R12475 gnd.n434 gnd.n433 9.3005
R12476 gnd.n7306 gnd.n7305 9.3005
R12477 gnd.n7307 gnd.n432 9.3005
R12478 gnd.n7309 gnd.n7308 9.3005
R12479 gnd.n428 gnd.n427 9.3005
R12480 gnd.n7316 gnd.n7315 9.3005
R12481 gnd.n7317 gnd.n426 9.3005
R12482 gnd.n7319 gnd.n7318 9.3005
R12483 gnd.n422 gnd.n421 9.3005
R12484 gnd.n7326 gnd.n7325 9.3005
R12485 gnd.n7327 gnd.n420 9.3005
R12486 gnd.n7329 gnd.n7328 9.3005
R12487 gnd.n416 gnd.n415 9.3005
R12488 gnd.n7336 gnd.n7335 9.3005
R12489 gnd.n7337 gnd.n414 9.3005
R12490 gnd.n7339 gnd.n7338 9.3005
R12491 gnd.n410 gnd.n409 9.3005
R12492 gnd.n7346 gnd.n7345 9.3005
R12493 gnd.n7347 gnd.n408 9.3005
R12494 gnd.n7349 gnd.n7348 9.3005
R12495 gnd.n404 gnd.n403 9.3005
R12496 gnd.n7356 gnd.n7355 9.3005
R12497 gnd.n7357 gnd.n402 9.3005
R12498 gnd.n7360 gnd.n7359 9.3005
R12499 gnd.n7358 gnd.n398 9.3005
R12500 gnd.n7366 gnd.n397 9.3005
R12501 gnd.n7368 gnd.n7367 9.3005
R12502 gnd.n7157 gnd.n522 9.3005
R12503 gnd.n7660 gnd.n130 9.3005
R12504 gnd.n7659 gnd.n132 9.3005
R12505 gnd.n136 gnd.n133 9.3005
R12506 gnd.n7654 gnd.n137 9.3005
R12507 gnd.n7653 gnd.n138 9.3005
R12508 gnd.n7652 gnd.n139 9.3005
R12509 gnd.n143 gnd.n140 9.3005
R12510 gnd.n7647 gnd.n144 9.3005
R12511 gnd.n7646 gnd.n145 9.3005
R12512 gnd.n7645 gnd.n146 9.3005
R12513 gnd.n150 gnd.n147 9.3005
R12514 gnd.n7640 gnd.n151 9.3005
R12515 gnd.n7639 gnd.n152 9.3005
R12516 gnd.n7638 gnd.n153 9.3005
R12517 gnd.n157 gnd.n154 9.3005
R12518 gnd.n7633 gnd.n158 9.3005
R12519 gnd.n7632 gnd.n159 9.3005
R12520 gnd.n7628 gnd.n160 9.3005
R12521 gnd.n164 gnd.n161 9.3005
R12522 gnd.n7623 gnd.n165 9.3005
R12523 gnd.n7622 gnd.n166 9.3005
R12524 gnd.n7621 gnd.n167 9.3005
R12525 gnd.n171 gnd.n168 9.3005
R12526 gnd.n7616 gnd.n172 9.3005
R12527 gnd.n7615 gnd.n173 9.3005
R12528 gnd.n7614 gnd.n174 9.3005
R12529 gnd.n178 gnd.n175 9.3005
R12530 gnd.n7609 gnd.n179 9.3005
R12531 gnd.n7608 gnd.n180 9.3005
R12532 gnd.n7607 gnd.n181 9.3005
R12533 gnd.n185 gnd.n182 9.3005
R12534 gnd.n7602 gnd.n186 9.3005
R12535 gnd.n7601 gnd.n187 9.3005
R12536 gnd.n7600 gnd.n188 9.3005
R12537 gnd.n192 gnd.n189 9.3005
R12538 gnd.n7595 gnd.n193 9.3005
R12539 gnd.n7594 gnd.n7593 9.3005
R12540 gnd.n7592 gnd.n196 9.3005
R12541 gnd.n7662 gnd.n7661 9.3005
R12542 gnd.n1835 gnd.n1834 9.3005
R12543 gnd.n4287 gnd.n4286 9.3005
R12544 gnd.n4288 gnd.n1833 9.3005
R12545 gnd.n4334 gnd.n4289 9.3005
R12546 gnd.n4333 gnd.n4290 9.3005
R12547 gnd.n4332 gnd.n4291 9.3005
R12548 gnd.n4331 gnd.n4292 9.3005
R12549 gnd.n4330 gnd.n4293 9.3005
R12550 gnd.n4328 gnd.n4294 9.3005
R12551 gnd.n4327 gnd.n4295 9.3005
R12552 gnd.n4325 gnd.n4296 9.3005
R12553 gnd.n4324 gnd.n4297 9.3005
R12554 gnd.n4323 gnd.n4298 9.3005
R12555 gnd.n4320 gnd.n4299 9.3005
R12556 gnd.n4319 gnd.n4300 9.3005
R12557 gnd.n4317 gnd.n4301 9.3005
R12558 gnd.n4316 gnd.n4302 9.3005
R12559 gnd.n4315 gnd.n4303 9.3005
R12560 gnd.n4312 gnd.n4304 9.3005
R12561 gnd.n4311 gnd.n4305 9.3005
R12562 gnd.n4309 gnd.n4306 9.3005
R12563 gnd.n4308 gnd.n4307 9.3005
R12564 gnd.n1713 gnd.n1712 9.3005
R12565 gnd.n4490 gnd.n4489 9.3005
R12566 gnd.n4491 gnd.n1711 9.3005
R12567 gnd.n4493 gnd.n4492 9.3005
R12568 gnd.n4494 gnd.n1710 9.3005
R12569 gnd.n4498 gnd.n4497 9.3005
R12570 gnd.n4499 gnd.n1709 9.3005
R12571 gnd.n4529 gnd.n4500 9.3005
R12572 gnd.n4528 gnd.n4501 9.3005
R12573 gnd.n4527 gnd.n4502 9.3005
R12574 gnd.n4526 gnd.n4503 9.3005
R12575 gnd.n4520 gnd.n4504 9.3005
R12576 gnd.n4519 gnd.n4505 9.3005
R12577 gnd.n4518 gnd.n4506 9.3005
R12578 gnd.n4517 gnd.n4507 9.3005
R12579 gnd.n4514 gnd.n4508 9.3005
R12580 gnd.n4513 gnd.n4510 9.3005
R12581 gnd.n4509 gnd.n346 9.3005
R12582 gnd.n7377 gnd.n347 9.3005
R12583 gnd.n7376 gnd.n348 9.3005
R12584 gnd.n7375 gnd.n349 9.3005
R12585 gnd.n394 gnd.n350 9.3005
R12586 gnd.n393 gnd.n351 9.3005
R12587 gnd.n391 gnd.n352 9.3005
R12588 gnd.n390 gnd.n353 9.3005
R12589 gnd.n388 gnd.n354 9.3005
R12590 gnd.n387 gnd.n355 9.3005
R12591 gnd.n385 gnd.n356 9.3005
R12592 gnd.n384 gnd.n357 9.3005
R12593 gnd.n382 gnd.n358 9.3005
R12594 gnd.n381 gnd.n359 9.3005
R12595 gnd.n379 gnd.n360 9.3005
R12596 gnd.n378 gnd.n361 9.3005
R12597 gnd.n376 gnd.n362 9.3005
R12598 gnd.n375 gnd.n363 9.3005
R12599 gnd.n373 gnd.n364 9.3005
R12600 gnd.n372 gnd.n365 9.3005
R12601 gnd.n370 gnd.n366 9.3005
R12602 gnd.n369 gnd.n368 9.3005
R12603 gnd.n367 gnd.n200 9.3005
R12604 gnd.n7589 gnd.n199 9.3005
R12605 gnd.n7591 gnd.n7590 9.3005
R12606 gnd.n2171 gnd.n2170 9.3005
R12607 gnd.n2179 gnd.n2178 9.3005
R12608 gnd.n2169 gnd.n2164 9.3005
R12609 gnd.n2185 gnd.n2163 9.3005
R12610 gnd.n2186 gnd.n2162 9.3005
R12611 gnd.n2187 gnd.n2161 9.3005
R12612 gnd.n2160 gnd.n2158 9.3005
R12613 gnd.n2193 gnd.n2157 9.3005
R12614 gnd.n2194 gnd.n2156 9.3005
R12615 gnd.n2195 gnd.n2155 9.3005
R12616 gnd.n2154 gnd.n2152 9.3005
R12617 gnd.n2201 gnd.n2151 9.3005
R12618 gnd.n2202 gnd.n2150 9.3005
R12619 gnd.n2203 gnd.n2149 9.3005
R12620 gnd.n2148 gnd.n2146 9.3005
R12621 gnd.n2209 gnd.n2145 9.3005
R12622 gnd.n2210 gnd.n2144 9.3005
R12623 gnd.n2211 gnd.n2143 9.3005
R12624 gnd.n2142 gnd.n2140 9.3005
R12625 gnd.n2217 gnd.n2139 9.3005
R12626 gnd.n2135 gnd.n2078 9.3005
R12627 gnd.n2134 gnd.n2133 9.3005
R12628 gnd.n2081 gnd.n2080 9.3005
R12629 gnd.n2124 gnd.n2084 9.3005
R12630 gnd.n2126 gnd.n2125 9.3005
R12631 gnd.n2123 gnd.n2086 9.3005
R12632 gnd.n2122 gnd.n2121 9.3005
R12633 gnd.n2088 gnd.n2087 9.3005
R12634 gnd.n2115 gnd.n2114 9.3005
R12635 gnd.n2113 gnd.n2090 9.3005
R12636 gnd.n2112 gnd.n2111 9.3005
R12637 gnd.n2092 gnd.n2091 9.3005
R12638 gnd.n2105 gnd.n2104 9.3005
R12639 gnd.n2103 gnd.n2094 9.3005
R12640 gnd.n2102 gnd.n2101 9.3005
R12641 gnd.n2097 gnd.n2096 9.3005
R12642 gnd.n2177 gnd.n2168 9.3005
R12643 gnd.n2176 gnd.n2175 9.3005
R12644 gnd.n4607 gnd.n1641 9.3005
R12645 gnd.n4606 gnd.n1642 9.3005
R12646 gnd.n4605 gnd.n1643 9.3005
R12647 gnd.n1821 gnd.n1644 9.3005
R12648 gnd.n1823 gnd.n1822 9.3005
R12649 gnd.n1802 gnd.n1801 9.3005
R12650 gnd.n4362 gnd.n4361 9.3005
R12651 gnd.n4363 gnd.n1800 9.3005
R12652 gnd.n4367 gnd.n4364 9.3005
R12653 gnd.n4366 gnd.n4365 9.3005
R12654 gnd.n1776 gnd.n1775 9.3005
R12655 gnd.n4394 gnd.n4393 9.3005
R12656 gnd.n4395 gnd.n1774 9.3005
R12657 gnd.n4399 gnd.n4396 9.3005
R12658 gnd.n4398 gnd.n4397 9.3005
R12659 gnd.n1750 gnd.n1749 9.3005
R12660 gnd.n4426 gnd.n4425 9.3005
R12661 gnd.n4427 gnd.n1748 9.3005
R12662 gnd.n4431 gnd.n4428 9.3005
R12663 gnd.n4430 gnd.n4429 9.3005
R12664 gnd.n1723 gnd.n1722 9.3005
R12665 gnd.n4480 gnd.n4479 9.3005
R12666 gnd.n4481 gnd.n1721 9.3005
R12667 gnd.n4485 gnd.n4482 9.3005
R12668 gnd.n4484 gnd.n4483 9.3005
R12669 gnd.n1688 gnd.n301 9.3005
R12670 gnd.n7420 gnd.n7419 9.3005
R12671 gnd.n285 gnd.n284 9.3005
R12672 gnd.n7433 gnd.n7432 9.3005
R12673 gnd.n7434 gnd.n283 9.3005
R12674 gnd.n7436 gnd.n7435 9.3005
R12675 gnd.n270 gnd.n269 9.3005
R12676 gnd.n7449 gnd.n7448 9.3005
R12677 gnd.n7450 gnd.n268 9.3005
R12678 gnd.n7452 gnd.n7451 9.3005
R12679 gnd.n254 gnd.n253 9.3005
R12680 gnd.n7465 gnd.n7464 9.3005
R12681 gnd.n7466 gnd.n252 9.3005
R12682 gnd.n7468 gnd.n7467 9.3005
R12683 gnd.n240 gnd.n239 9.3005
R12684 gnd.n7481 gnd.n7480 9.3005
R12685 gnd.n7482 gnd.n238 9.3005
R12686 gnd.n7484 gnd.n7483 9.3005
R12687 gnd.n224 gnd.n223 9.3005
R12688 gnd.n7497 gnd.n7496 9.3005
R12689 gnd.n7498 gnd.n222 9.3005
R12690 gnd.n7500 gnd.n7499 9.3005
R12691 gnd.n207 gnd.n206 9.3005
R12692 gnd.n7581 gnd.n7580 9.3005
R12693 gnd.n7582 gnd.n205 9.3005
R12694 gnd.n7584 gnd.n7583 9.3005
R12695 gnd.n129 gnd.n128 9.3005
R12696 gnd.n7664 gnd.n7663 9.3005
R12697 gnd.n2095 gnd.n1640 9.3005
R12698 gnd.n7418 gnd.n300 9.3005
R12699 gnd.n2834 gnd.n2771 9.3005
R12700 gnd.n2833 gnd.n2778 9.3005
R12701 gnd.n2781 gnd.n2779 9.3005
R12702 gnd.n2829 gnd.n2782 9.3005
R12703 gnd.n2828 gnd.n2783 9.3005
R12704 gnd.n2827 gnd.n2784 9.3005
R12705 gnd.n2787 gnd.n2785 9.3005
R12706 gnd.n2823 gnd.n2788 9.3005
R12707 gnd.n2822 gnd.n2789 9.3005
R12708 gnd.n2821 gnd.n2790 9.3005
R12709 gnd.n2793 gnd.n2791 9.3005
R12710 gnd.n2817 gnd.n2794 9.3005
R12711 gnd.n2816 gnd.n2795 9.3005
R12712 gnd.n2815 gnd.n2796 9.3005
R12713 gnd.n2799 gnd.n2797 9.3005
R12714 gnd.n2811 gnd.n2800 9.3005
R12715 gnd.n2810 gnd.n2801 9.3005
R12716 gnd.n2809 gnd.n2802 9.3005
R12717 gnd.n2806 gnd.n2803 9.3005
R12718 gnd.n2805 gnd.n2804 9.3005
R12719 gnd.n2686 gnd.n2685 9.3005
R12720 gnd.n3201 gnd.n3200 9.3005
R12721 gnd.n3202 gnd.n2684 9.3005
R12722 gnd.n3204 gnd.n3203 9.3005
R12723 gnd.n2682 gnd.n2681 9.3005
R12724 gnd.n3209 gnd.n3208 9.3005
R12725 gnd.n3210 gnd.n2680 9.3005
R12726 gnd.n3212 gnd.n3211 9.3005
R12727 gnd.n2678 gnd.n2677 9.3005
R12728 gnd.n3218 gnd.n3217 9.3005
R12729 gnd.n3219 gnd.n2676 9.3005
R12730 gnd.n3226 gnd.n3220 9.3005
R12731 gnd.n3225 gnd.n3221 9.3005
R12732 gnd.n3224 gnd.n3222 9.3005
R12733 gnd.n2553 gnd.n2552 9.3005
R12734 gnd.n3396 gnd.n3395 9.3005
R12735 gnd.n3397 gnd.n2551 9.3005
R12736 gnd.n3401 gnd.n3398 9.3005
R12737 gnd.n3400 gnd.n3399 9.3005
R12738 gnd.n2528 gnd.n2527 9.3005
R12739 gnd.n3426 gnd.n3425 9.3005
R12740 gnd.n3427 gnd.n2526 9.3005
R12741 gnd.n3437 gnd.n3428 9.3005
R12742 gnd.n3436 gnd.n3429 9.3005
R12743 gnd.n3435 gnd.n3430 9.3005
R12744 gnd.n3432 gnd.n3431 9.3005
R12745 gnd.n2493 gnd.n2492 9.3005
R12746 gnd.n3473 gnd.n3472 9.3005
R12747 gnd.n3474 gnd.n2491 9.3005
R12748 gnd.n3478 gnd.n3475 9.3005
R12749 gnd.n3477 gnd.n3476 9.3005
R12750 gnd.n2478 gnd.n2477 9.3005
R12751 gnd.n3595 gnd.n3594 9.3005
R12752 gnd.n3596 gnd.n2476 9.3005
R12753 gnd.n3598 gnd.n3597 9.3005
R12754 gnd.n2457 gnd.n2456 9.3005
R12755 gnd.n3622 gnd.n3621 9.3005
R12756 gnd.n3623 gnd.n2455 9.3005
R12757 gnd.n3627 gnd.n3624 9.3005
R12758 gnd.n3626 gnd.n3625 9.3005
R12759 gnd.n2424 gnd.n2423 9.3005
R12760 gnd.n3664 gnd.n3663 9.3005
R12761 gnd.n3665 gnd.n2422 9.3005
R12762 gnd.n3678 gnd.n3666 9.3005
R12763 gnd.n3677 gnd.n3667 9.3005
R12764 gnd.n3676 gnd.n3668 9.3005
R12765 gnd.n3670 gnd.n3669 9.3005
R12766 gnd.n2390 gnd.n2389 9.3005
R12767 gnd.n3747 gnd.n3746 9.3005
R12768 gnd.n3748 gnd.n2388 9.3005
R12769 gnd.n3750 gnd.n3749 9.3005
R12770 gnd.n2367 gnd.n2366 9.3005
R12771 gnd.n3790 gnd.n3789 9.3005
R12772 gnd.n3791 gnd.n2365 9.3005
R12773 gnd.n3793 gnd.n3792 9.3005
R12774 gnd.n2351 gnd.n2350 9.3005
R12775 gnd.n3838 gnd.n3837 9.3005
R12776 gnd.n3839 gnd.n2349 9.3005
R12777 gnd.n3843 gnd.n3840 9.3005
R12778 gnd.n3842 gnd.n3841 9.3005
R12779 gnd.n2322 gnd.n2321 9.3005
R12780 gnd.n3875 gnd.n3874 9.3005
R12781 gnd.n3876 gnd.n2320 9.3005
R12782 gnd.n3878 gnd.n3877 9.3005
R12783 gnd.n2285 gnd.n2284 9.3005
R12784 gnd.n3909 gnd.n3908 9.3005
R12785 gnd.n3910 gnd.n2283 9.3005
R12786 gnd.n3914 gnd.n3911 9.3005
R12787 gnd.n3913 gnd.n3912 9.3005
R12788 gnd.n2256 gnd.n2255 9.3005
R12789 gnd.n3961 gnd.n3960 9.3005
R12790 gnd.n3962 gnd.n2254 9.3005
R12791 gnd.n3964 gnd.n3963 9.3005
R12792 gnd.n2237 gnd.n2236 9.3005
R12793 gnd.n3987 gnd.n3986 9.3005
R12794 gnd.n3988 gnd.n2235 9.3005
R12795 gnd.n3992 gnd.n3989 9.3005
R12796 gnd.n3991 gnd.n3990 9.3005
R12797 gnd.n2036 gnd.n2035 9.3005
R12798 gnd.n4179 gnd.n4178 9.3005
R12799 gnd.n4180 gnd.n2034 9.3005
R12800 gnd.n4182 gnd.n4181 9.3005
R12801 gnd.n2024 gnd.n2023 9.3005
R12802 gnd.n4200 gnd.n4199 9.3005
R12803 gnd.n4201 gnd.n2022 9.3005
R12804 gnd.n4203 gnd.n4202 9.3005
R12805 gnd.n2012 gnd.n2011 9.3005
R12806 gnd.n4221 gnd.n4220 9.3005
R12807 gnd.n4222 gnd.n2010 9.3005
R12808 gnd.n4224 gnd.n4223 9.3005
R12809 gnd.n2000 gnd.n1999 9.3005
R12810 gnd.n4244 gnd.n4243 9.3005
R12811 gnd.n4245 gnd.n1998 9.3005
R12812 gnd.n4248 gnd.n4247 9.3005
R12813 gnd.n4246 gnd.n1617 9.3005
R12814 gnd.n4622 gnd.n1618 9.3005
R12815 gnd.n4621 gnd.n1619 9.3005
R12816 gnd.n4620 gnd.n1620 9.3005
R12817 gnd.n1626 gnd.n1621 9.3005
R12818 gnd.n4614 gnd.n1627 9.3005
R12819 gnd.n4613 gnd.n1628 9.3005
R12820 gnd.n4612 gnd.n1629 9.3005
R12821 gnd.n1815 gnd.n1630 9.3005
R12822 gnd.n1816 gnd.n1814 9.3005
R12823 gnd.n1818 gnd.n1817 9.3005
R12824 gnd.n1812 gnd.n1811 9.3005
R12825 gnd.n4351 gnd.n4350 9.3005
R12826 gnd.n4352 gnd.n1810 9.3005
R12827 gnd.n4356 gnd.n4353 9.3005
R12828 gnd.n4355 gnd.n4354 9.3005
R12829 gnd.n1785 gnd.n1784 9.3005
R12830 gnd.n4382 gnd.n4381 9.3005
R12831 gnd.n4383 gnd.n1783 9.3005
R12832 gnd.n4387 gnd.n4384 9.3005
R12833 gnd.n4386 gnd.n4385 9.3005
R12834 gnd.n1759 gnd.n1758 9.3005
R12835 gnd.n4415 gnd.n4414 9.3005
R12836 gnd.n4416 gnd.n1757 9.3005
R12837 gnd.n4420 gnd.n4417 9.3005
R12838 gnd.n4419 gnd.n4418 9.3005
R12839 gnd.n1732 gnd.n1731 9.3005
R12840 gnd.n4452 gnd.n4451 9.3005
R12841 gnd.n4453 gnd.n1730 9.3005
R12842 gnd.n4474 gnd.n4454 9.3005
R12843 gnd.n4473 gnd.n4455 9.3005
R12844 gnd.n4472 gnd.n4456 9.3005
R12845 gnd.n4459 gnd.n4457 9.3005
R12846 gnd.n4466 gnd.n4460 9.3005
R12847 gnd.n7388 gnd.n337 9.3005
R12848 gnd.n340 gnd.n338 9.3005
R12849 gnd.n7384 gnd.n341 9.3005
R12850 gnd.n7383 gnd.n342 9.3005
R12851 gnd.n7382 gnd.n343 9.3005
R12852 gnd.n396 gnd.n344 9.3005
R12853 gnd.n7370 gnd.n7369 9.3005
R12854 gnd.n3079 gnd.n3078 9.3005
R12855 gnd.n2912 gnd.n2911 9.3005
R12856 gnd.n2996 gnd.n2995 9.3005
R12857 gnd.n2997 gnd.n2910 9.3005
R12858 gnd.n3000 gnd.n2998 9.3005
R12859 gnd.n3001 gnd.n2909 9.3005
R12860 gnd.n3004 gnd.n3003 9.3005
R12861 gnd.n3005 gnd.n2908 9.3005
R12862 gnd.n3008 gnd.n3006 9.3005
R12863 gnd.n3009 gnd.n2907 9.3005
R12864 gnd.n3012 gnd.n3011 9.3005
R12865 gnd.n3013 gnd.n2906 9.3005
R12866 gnd.n3016 gnd.n3014 9.3005
R12867 gnd.n3017 gnd.n2905 9.3005
R12868 gnd.n3020 gnd.n3019 9.3005
R12869 gnd.n3021 gnd.n2904 9.3005
R12870 gnd.n3024 gnd.n3022 9.3005
R12871 gnd.n3025 gnd.n2903 9.3005
R12872 gnd.n3028 gnd.n3027 9.3005
R12873 gnd.n3029 gnd.n2902 9.3005
R12874 gnd.n3031 gnd.n3030 9.3005
R12875 gnd.n2863 gnd.n2862 9.3005
R12876 gnd.n3044 gnd.n3043 9.3005
R12877 gnd.n3045 gnd.n2861 9.3005
R12878 gnd.n3047 gnd.n3046 9.3005
R12879 gnd.n2746 gnd.n2745 9.3005
R12880 gnd.n3060 gnd.n3059 9.3005
R12881 gnd.n3061 gnd.n2744 9.3005
R12882 gnd.n3063 gnd.n3062 9.3005
R12883 gnd.n2740 gnd.n2739 9.3005
R12884 gnd.n3076 gnd.n3075 9.3005
R12885 gnd.n3077 gnd.n2738 9.3005
R12886 gnd.n2938 gnd.n2937 9.3005
R12887 gnd.n2943 gnd.n2942 9.3005
R12888 gnd.n2946 gnd.n2932 9.3005
R12889 gnd.n2947 gnd.n2931 9.3005
R12890 gnd.n2950 gnd.n2930 9.3005
R12891 gnd.n2951 gnd.n2929 9.3005
R12892 gnd.n2954 gnd.n2928 9.3005
R12893 gnd.n2955 gnd.n2927 9.3005
R12894 gnd.n2958 gnd.n2926 9.3005
R12895 gnd.n2959 gnd.n2925 9.3005
R12896 gnd.n2962 gnd.n2924 9.3005
R12897 gnd.n2963 gnd.n2923 9.3005
R12898 gnd.n2966 gnd.n2922 9.3005
R12899 gnd.n2967 gnd.n2921 9.3005
R12900 gnd.n2970 gnd.n2920 9.3005
R12901 gnd.n2971 gnd.n2919 9.3005
R12902 gnd.n2974 gnd.n2918 9.3005
R12903 gnd.n2977 gnd.n2976 9.3005
R12904 gnd.n2941 gnd.n2936 9.3005
R12905 gnd.n2940 gnd.n2939 9.3005
R12906 gnd.n2984 gnd.n2983 9.3005
R12907 gnd.n2982 gnd.n2917 9.3005
R12908 gnd.n2981 gnd.n2980 9.3005
R12909 gnd.n2979 gnd.n1111 9.3005
R12910 gnd.n5012 gnd.n1112 9.3005
R12911 gnd.n5011 gnd.n1113 9.3005
R12912 gnd.n5010 gnd.n1114 9.3005
R12913 gnd.n1130 gnd.n1115 9.3005
R12914 gnd.n5000 gnd.n1131 9.3005
R12915 gnd.n4999 gnd.n1132 9.3005
R12916 gnd.n4998 gnd.n1133 9.3005
R12917 gnd.n1151 gnd.n1134 9.3005
R12918 gnd.n4988 gnd.n1152 9.3005
R12919 gnd.n4987 gnd.n1153 9.3005
R12920 gnd.n4986 gnd.n1154 9.3005
R12921 gnd.n1170 gnd.n1155 9.3005
R12922 gnd.n4976 gnd.n1171 9.3005
R12923 gnd.n4975 gnd.n1172 9.3005
R12924 gnd.n4974 gnd.n1173 9.3005
R12925 gnd.n1192 gnd.n1174 9.3005
R12926 gnd.n4964 gnd.n1193 9.3005
R12927 gnd.n4963 gnd.n1194 9.3005
R12928 gnd.n4962 gnd.n1195 9.3005
R12929 gnd.n1213 gnd.n1196 9.3005
R12930 gnd.n4952 gnd.n1214 9.3005
R12931 gnd.n4951 gnd.n1215 9.3005
R12932 gnd.n4950 gnd.n1216 9.3005
R12933 gnd.n1233 gnd.n1217 9.3005
R12934 gnd.n4939 gnd.n1234 9.3005
R12935 gnd.n4938 gnd.n1235 9.3005
R12936 gnd.n4937 gnd.n1236 9.3005
R12937 gnd.n2735 gnd.n1237 9.3005
R12938 gnd.n4926 gnd.n1251 9.3005
R12939 gnd.n4925 gnd.n1252 9.3005
R12940 gnd.n4924 gnd.n1253 9.3005
R12941 gnd.n1269 gnd.n1254 9.3005
R12942 gnd.n4913 gnd.n1270 9.3005
R12943 gnd.n4912 gnd.n1271 9.3005
R12944 gnd.n4911 gnd.n1272 9.3005
R12945 gnd.n1290 gnd.n1273 9.3005
R12946 gnd.n4901 gnd.n1291 9.3005
R12947 gnd.n4900 gnd.n1292 9.3005
R12948 gnd.n4899 gnd.n1293 9.3005
R12949 gnd.n1311 gnd.n1294 9.3005
R12950 gnd.n4889 gnd.n1312 9.3005
R12951 gnd.n4888 gnd.n1313 9.3005
R12952 gnd.n4887 gnd.n1314 9.3005
R12953 gnd.n1332 gnd.n1315 9.3005
R12954 gnd.n4877 gnd.n1333 9.3005
R12955 gnd.n4876 gnd.n1334 9.3005
R12956 gnd.n4875 gnd.n1335 9.3005
R12957 gnd.n1353 gnd.n1336 9.3005
R12958 gnd.n4865 gnd.n1354 9.3005
R12959 gnd.n4864 gnd.n1355 9.3005
R12960 gnd.n4863 gnd.n1356 9.3005
R12961 gnd.n1374 gnd.n1357 9.3005
R12962 gnd.n4853 gnd.n1375 9.3005
R12963 gnd.n4852 gnd.n1376 9.3005
R12964 gnd.n4851 gnd.n1377 9.3005
R12965 gnd.n1396 gnd.n1378 9.3005
R12966 gnd.n4841 gnd.n1397 9.3005
R12967 gnd.n4840 gnd.n1398 9.3005
R12968 gnd.n4839 gnd.n1399 9.3005
R12969 gnd.n2569 gnd.n1400 9.3005
R12970 gnd.n2978 gnd.n2916 9.3005
R12971 gnd.n4801 gnd.n1456 9.3005
R12972 gnd.n4804 gnd.n1455 9.3005
R12973 gnd.n4805 gnd.n1454 9.3005
R12974 gnd.n4808 gnd.n1453 9.3005
R12975 gnd.n4809 gnd.n1452 9.3005
R12976 gnd.n4812 gnd.n1451 9.3005
R12977 gnd.n4813 gnd.n1450 9.3005
R12978 gnd.n4816 gnd.n1449 9.3005
R12979 gnd.n4817 gnd.n1448 9.3005
R12980 gnd.n4820 gnd.n1447 9.3005
R12981 gnd.n4821 gnd.n1446 9.3005
R12982 gnd.n4824 gnd.n1445 9.3005
R12983 gnd.n4825 gnd.n1444 9.3005
R12984 gnd.n4826 gnd.n1443 9.3005
R12985 gnd.n1410 gnd.n1409 9.3005
R12986 gnd.n4832 gnd.n4831 9.3005
R12987 gnd.n3279 gnd.n3277 9.3005
R12988 gnd.n3281 gnd.n3280 9.3005
R12989 gnd.n3284 gnd.n3274 9.3005
R12990 gnd.n3288 gnd.n3287 9.3005
R12991 gnd.n3289 gnd.n3273 9.3005
R12992 gnd.n3291 gnd.n3290 9.3005
R12993 gnd.n3294 gnd.n3272 9.3005
R12994 gnd.n3298 gnd.n3297 9.3005
R12995 gnd.n3299 gnd.n3271 9.3005
R12996 gnd.n3301 gnd.n3300 9.3005
R12997 gnd.n3304 gnd.n3270 9.3005
R12998 gnd.n3308 gnd.n3307 9.3005
R12999 gnd.n3309 gnd.n3269 9.3005
R13000 gnd.n3311 gnd.n3310 9.3005
R13001 gnd.n3314 gnd.n3268 9.3005
R13002 gnd.n3318 gnd.n3317 9.3005
R13003 gnd.n3319 gnd.n3267 9.3005
R13004 gnd.n3322 gnd.n3320 9.3005
R13005 gnd.n3323 gnd.n3263 9.3005
R13006 gnd.n3325 gnd.n3324 9.3005
R13007 gnd.n3278 gnd.n1457 9.3005
R13008 gnd.n5026 gnd.n5025 9.3005
R13009 gnd.n5024 gnd.n1089 9.3005
R13010 gnd.n5023 gnd.n5022 9.3005
R13011 gnd.n1091 gnd.n1090 9.3005
R13012 gnd.n2873 gnd.n2872 9.3005
R13013 gnd.n2876 gnd.n2874 9.3005
R13014 gnd.n2877 gnd.n2871 9.3005
R13015 gnd.n2880 gnd.n2879 9.3005
R13016 gnd.n2881 gnd.n2870 9.3005
R13017 gnd.n2884 gnd.n2882 9.3005
R13018 gnd.n2885 gnd.n2869 9.3005
R13019 gnd.n2888 gnd.n2887 9.3005
R13020 gnd.n2889 gnd.n2868 9.3005
R13021 gnd.n2892 gnd.n2890 9.3005
R13022 gnd.n2893 gnd.n2867 9.3005
R13023 gnd.n2896 gnd.n2895 9.3005
R13024 gnd.n2897 gnd.n2866 9.3005
R13025 gnd.n2900 gnd.n2898 9.3005
R13026 gnd.n2901 gnd.n2865 9.3005
R13027 gnd.n3036 gnd.n3035 9.3005
R13028 gnd.n3037 gnd.n2864 9.3005
R13029 gnd.n3039 gnd.n3038 9.3005
R13030 gnd.n2860 gnd.n2859 9.3005
R13031 gnd.n3052 gnd.n3051 9.3005
R13032 gnd.n3053 gnd.n2858 9.3005
R13033 gnd.n3055 gnd.n3054 9.3005
R13034 gnd.n2743 gnd.n2742 9.3005
R13035 gnd.n3068 gnd.n3067 9.3005
R13036 gnd.n3069 gnd.n2741 9.3005
R13037 gnd.n3071 gnd.n3070 9.3005
R13038 gnd.n2737 gnd.n2736 9.3005
R13039 gnd.n3084 gnd.n3083 9.3005
R13040 gnd.n3085 gnd.n2734 9.3005
R13041 gnd.n3087 gnd.n3086 9.3005
R13042 gnd.n2729 gnd.n2728 9.3005
R13043 gnd.n3100 gnd.n3099 9.3005
R13044 gnd.n3101 gnd.n2727 9.3005
R13045 gnd.n3103 gnd.n3102 9.3005
R13046 gnd.n2723 gnd.n2722 9.3005
R13047 gnd.n3116 gnd.n3115 9.3005
R13048 gnd.n3117 gnd.n2721 9.3005
R13049 gnd.n3119 gnd.n3118 9.3005
R13050 gnd.n2715 gnd.n2714 9.3005
R13051 gnd.n3132 gnd.n3131 9.3005
R13052 gnd.n3133 gnd.n2713 9.3005
R13053 gnd.n3135 gnd.n3134 9.3005
R13054 gnd.n2709 gnd.n2708 9.3005
R13055 gnd.n3148 gnd.n3147 9.3005
R13056 gnd.n3149 gnd.n2707 9.3005
R13057 gnd.n3151 gnd.n3150 9.3005
R13058 gnd.n2701 gnd.n2700 9.3005
R13059 gnd.n3164 gnd.n3163 9.3005
R13060 gnd.n3165 gnd.n2699 9.3005
R13061 gnd.n3168 gnd.n3167 9.3005
R13062 gnd.n3166 gnd.n2694 9.3005
R13063 gnd.n3180 gnd.n2695 9.3005
R13064 gnd.n3181 gnd.n2693 9.3005
R13065 gnd.n3183 gnd.n3182 9.3005
R13066 gnd.n3184 gnd.n2692 9.3005
R13067 gnd.n3186 gnd.n3185 9.3005
R13068 gnd.n2627 gnd.n2626 9.3005
R13069 gnd.n3261 gnd.n3260 9.3005
R13070 gnd.n3262 gnd.n2625 9.3005
R13071 gnd.n3327 gnd.n3326 9.3005
R13072 gnd.n5027 gnd.n1087 9.3005
R13073 gnd.n5034 gnd.n5033 9.3005
R13074 gnd.n5035 gnd.n1081 9.3005
R13075 gnd.n5038 gnd.n1080 9.3005
R13076 gnd.n5039 gnd.n1079 9.3005
R13077 gnd.n5042 gnd.n1078 9.3005
R13078 gnd.n5043 gnd.n1077 9.3005
R13079 gnd.n5046 gnd.n1076 9.3005
R13080 gnd.n5047 gnd.n1075 9.3005
R13081 gnd.n5050 gnd.n1074 9.3005
R13082 gnd.n5051 gnd.n1073 9.3005
R13083 gnd.n5054 gnd.n1072 9.3005
R13084 gnd.n5055 gnd.n1071 9.3005
R13085 gnd.n5058 gnd.n1070 9.3005
R13086 gnd.n5059 gnd.n1069 9.3005
R13087 gnd.n5062 gnd.n1068 9.3005
R13088 gnd.n5063 gnd.n1067 9.3005
R13089 gnd.n5066 gnd.n1066 9.3005
R13090 gnd.n5067 gnd.n1065 9.3005
R13091 gnd.n5070 gnd.n1064 9.3005
R13092 gnd.n5072 gnd.n1061 9.3005
R13093 gnd.n5075 gnd.n1060 9.3005
R13094 gnd.n5076 gnd.n1059 9.3005
R13095 gnd.n5079 gnd.n1058 9.3005
R13096 gnd.n5080 gnd.n1057 9.3005
R13097 gnd.n5083 gnd.n1056 9.3005
R13098 gnd.n5084 gnd.n1055 9.3005
R13099 gnd.n5087 gnd.n1054 9.3005
R13100 gnd.n5088 gnd.n1053 9.3005
R13101 gnd.n5091 gnd.n1052 9.3005
R13102 gnd.n5092 gnd.n1051 9.3005
R13103 gnd.n5095 gnd.n1050 9.3005
R13104 gnd.n5096 gnd.n1049 9.3005
R13105 gnd.n5099 gnd.n1048 9.3005
R13106 gnd.n5101 gnd.n1047 9.3005
R13107 gnd.n5102 gnd.n1046 9.3005
R13108 gnd.n5103 gnd.n1045 9.3005
R13109 gnd.n5104 gnd.n1044 9.3005
R13110 gnd.n5032 gnd.n1086 9.3005
R13111 gnd.n5031 gnd.n5030 9.3005
R13112 gnd.n2990 gnd.n2989 9.3005
R13113 gnd.n2988 gnd.n1100 9.3005
R13114 gnd.n5018 gnd.n1101 9.3005
R13115 gnd.n5017 gnd.n1102 9.3005
R13116 gnd.n5016 gnd.n1103 9.3005
R13117 gnd.n1121 gnd.n1104 9.3005
R13118 gnd.n5006 gnd.n1122 9.3005
R13119 gnd.n5005 gnd.n1123 9.3005
R13120 gnd.n5004 gnd.n1124 9.3005
R13121 gnd.n1141 gnd.n1125 9.3005
R13122 gnd.n4994 gnd.n1142 9.3005
R13123 gnd.n4993 gnd.n1143 9.3005
R13124 gnd.n4992 gnd.n1144 9.3005
R13125 gnd.n1161 gnd.n1145 9.3005
R13126 gnd.n4982 gnd.n1162 9.3005
R13127 gnd.n4981 gnd.n1163 9.3005
R13128 gnd.n4980 gnd.n1164 9.3005
R13129 gnd.n1181 gnd.n1165 9.3005
R13130 gnd.n4970 gnd.n1182 9.3005
R13131 gnd.n4969 gnd.n1183 9.3005
R13132 gnd.n4968 gnd.n1184 9.3005
R13133 gnd.n1203 gnd.n1185 9.3005
R13134 gnd.n4958 gnd.n1204 9.3005
R13135 gnd.n4957 gnd.n1205 9.3005
R13136 gnd.n4956 gnd.n1206 9.3005
R13137 gnd.n1224 gnd.n1207 9.3005
R13138 gnd.n1280 gnd.n1262 9.3005
R13139 gnd.n4907 gnd.n1281 9.3005
R13140 gnd.n4906 gnd.n1282 9.3005
R13141 gnd.n4905 gnd.n1283 9.3005
R13142 gnd.n1300 gnd.n1284 9.3005
R13143 gnd.n4895 gnd.n1301 9.3005
R13144 gnd.n4894 gnd.n1302 9.3005
R13145 gnd.n4893 gnd.n1303 9.3005
R13146 gnd.n1322 gnd.n1304 9.3005
R13147 gnd.n4883 gnd.n1323 9.3005
R13148 gnd.n4882 gnd.n1324 9.3005
R13149 gnd.n4881 gnd.n1325 9.3005
R13150 gnd.n1342 gnd.n1326 9.3005
R13151 gnd.n4871 gnd.n1343 9.3005
R13152 gnd.n4870 gnd.n1344 9.3005
R13153 gnd.n4869 gnd.n1345 9.3005
R13154 gnd.n1364 gnd.n1346 9.3005
R13155 gnd.n4859 gnd.n1365 9.3005
R13156 gnd.n4858 gnd.n1366 9.3005
R13157 gnd.n4857 gnd.n1367 9.3005
R13158 gnd.n1385 gnd.n1368 9.3005
R13159 gnd.n4847 gnd.n1386 9.3005
R13160 gnd.n4846 gnd.n1387 9.3005
R13161 gnd.n4845 gnd.n1388 9.3005
R13162 gnd.n1407 gnd.n1389 9.3005
R13163 gnd.n4835 gnd.n1408 9.3005
R13164 gnd.n4834 gnd.n4833 9.3005
R13165 gnd.n2987 gnd.n2986 9.3005
R13166 gnd.n4917 gnd.n1225 9.3005
R13167 gnd.n2760 gnd.n2759 9.3005
R13168 gnd.n2751 gnd.n2750 9.3005
R13169 gnd.n2765 gnd.n2764 9.3005
R13170 gnd.n2766 gnd.n2749 9.3005
R13171 gnd.n2855 gnd.n2767 9.3005
R13172 gnd.n2854 gnd.n2768 9.3005
R13173 gnd.n2758 gnd.n2753 9.3005
R13174 gnd.n2754 gnd.n961 9.3005
R13175 gnd.n6537 gnd.n960 9.3005
R13176 gnd.n6538 gnd.n959 9.3005
R13177 gnd.n6539 gnd.n958 9.3005
R13178 gnd.n957 gnd.n953 9.3005
R13179 gnd.n6545 gnd.n952 9.3005
R13180 gnd.n6546 gnd.n951 9.3005
R13181 gnd.n6547 gnd.n950 9.3005
R13182 gnd.n949 gnd.n945 9.3005
R13183 gnd.n6553 gnd.n944 9.3005
R13184 gnd.n6554 gnd.n943 9.3005
R13185 gnd.n6555 gnd.n942 9.3005
R13186 gnd.n941 gnd.n937 9.3005
R13187 gnd.n6561 gnd.n936 9.3005
R13188 gnd.n6562 gnd.n935 9.3005
R13189 gnd.n6563 gnd.n934 9.3005
R13190 gnd.n933 gnd.n929 9.3005
R13191 gnd.n6569 gnd.n928 9.3005
R13192 gnd.n6570 gnd.n927 9.3005
R13193 gnd.n6571 gnd.n926 9.3005
R13194 gnd.n925 gnd.n921 9.3005
R13195 gnd.n6577 gnd.n920 9.3005
R13196 gnd.n6578 gnd.n919 9.3005
R13197 gnd.n6579 gnd.n918 9.3005
R13198 gnd.n917 gnd.n913 9.3005
R13199 gnd.n6585 gnd.n912 9.3005
R13200 gnd.n6586 gnd.n911 9.3005
R13201 gnd.n6587 gnd.n910 9.3005
R13202 gnd.n909 gnd.n905 9.3005
R13203 gnd.n6593 gnd.n904 9.3005
R13204 gnd.n6594 gnd.n903 9.3005
R13205 gnd.n6595 gnd.n902 9.3005
R13206 gnd.n901 gnd.n897 9.3005
R13207 gnd.n6601 gnd.n896 9.3005
R13208 gnd.n6602 gnd.n895 9.3005
R13209 gnd.n6603 gnd.n894 9.3005
R13210 gnd.n893 gnd.n889 9.3005
R13211 gnd.n6609 gnd.n888 9.3005
R13212 gnd.n6610 gnd.n887 9.3005
R13213 gnd.n6611 gnd.n886 9.3005
R13214 gnd.n885 gnd.n881 9.3005
R13215 gnd.n6617 gnd.n880 9.3005
R13216 gnd.n6618 gnd.n879 9.3005
R13217 gnd.n6619 gnd.n878 9.3005
R13218 gnd.n877 gnd.n873 9.3005
R13219 gnd.n6625 gnd.n872 9.3005
R13220 gnd.n6626 gnd.n871 9.3005
R13221 gnd.n6627 gnd.n870 9.3005
R13222 gnd.n869 gnd.n865 9.3005
R13223 gnd.n6633 gnd.n864 9.3005
R13224 gnd.n6634 gnd.n863 9.3005
R13225 gnd.n6635 gnd.n862 9.3005
R13226 gnd.n861 gnd.n857 9.3005
R13227 gnd.n6641 gnd.n856 9.3005
R13228 gnd.n6642 gnd.n855 9.3005
R13229 gnd.n6643 gnd.n854 9.3005
R13230 gnd.n853 gnd.n849 9.3005
R13231 gnd.n6649 gnd.n848 9.3005
R13232 gnd.n6650 gnd.n847 9.3005
R13233 gnd.n6651 gnd.n846 9.3005
R13234 gnd.n845 gnd.n841 9.3005
R13235 gnd.n6657 gnd.n840 9.3005
R13236 gnd.n6658 gnd.n839 9.3005
R13237 gnd.n6659 gnd.n838 9.3005
R13238 gnd.n837 gnd.n833 9.3005
R13239 gnd.n6665 gnd.n832 9.3005
R13240 gnd.n6666 gnd.n831 9.3005
R13241 gnd.n6667 gnd.n830 9.3005
R13242 gnd.n829 gnd.n825 9.3005
R13243 gnd.n6673 gnd.n824 9.3005
R13244 gnd.n6674 gnd.n823 9.3005
R13245 gnd.n6675 gnd.n822 9.3005
R13246 gnd.n821 gnd.n817 9.3005
R13247 gnd.n6681 gnd.n816 9.3005
R13248 gnd.n6682 gnd.n815 9.3005
R13249 gnd.n6683 gnd.n814 9.3005
R13250 gnd.n813 gnd.n809 9.3005
R13251 gnd.n6689 gnd.n808 9.3005
R13252 gnd.n6690 gnd.n807 9.3005
R13253 gnd.n6691 gnd.n806 9.3005
R13254 gnd.n805 gnd.n801 9.3005
R13255 gnd.n6697 gnd.n800 9.3005
R13256 gnd.n6698 gnd.n799 9.3005
R13257 gnd.n6699 gnd.n798 9.3005
R13258 gnd.n2757 gnd.n2756 9.3005
R13259 gnd.n1896 gnd.n1895 9.3005
R13260 gnd.n1874 gnd.n1873 9.3005
R13261 gnd.n1908 gnd.n1907 9.3005
R13262 gnd.n1871 gnd.n1869 9.3005
R13263 gnd.n1915 gnd.n1914 9.3005
R13264 gnd.n1865 gnd.n1864 9.3005
R13265 gnd.n1927 gnd.n1926 9.3005
R13266 gnd.n1862 gnd.n1860 9.3005
R13267 gnd.n1934 gnd.n1933 9.3005
R13268 gnd.n1856 gnd.n1855 9.3005
R13269 gnd.n1946 gnd.n1945 9.3005
R13270 gnd.n1853 gnd.n1851 9.3005
R13271 gnd.n1953 gnd.n1952 9.3005
R13272 gnd.n1847 gnd.n1846 9.3005
R13273 gnd.n1965 gnd.n1964 9.3005
R13274 gnd.n1844 gnd.n1842 9.3005
R13275 gnd.n4273 gnd.n4272 9.3005
R13276 gnd.n4271 gnd.n1843 9.3005
R13277 gnd.n1891 gnd.n1889 9.3005
R13278 gnd.n1962 gnd.n1961 9.3005
R13279 gnd.n1852 gnd.n1848 9.3005
R13280 gnd.n1955 gnd.n1954 9.3005
R13281 gnd.n1944 gnd.n1850 9.3005
R13282 gnd.n1943 gnd.n1942 9.3005
R13283 gnd.n1861 gnd.n1857 9.3005
R13284 gnd.n1936 gnd.n1935 9.3005
R13285 gnd.n1925 gnd.n1859 9.3005
R13286 gnd.n1924 gnd.n1923 9.3005
R13287 gnd.n1870 gnd.n1866 9.3005
R13288 gnd.n1917 gnd.n1916 9.3005
R13289 gnd.n1906 gnd.n1868 9.3005
R13290 gnd.n1905 gnd.n1904 9.3005
R13291 gnd.n1890 gnd.n1875 9.3005
R13292 gnd.n1898 gnd.n1897 9.3005
R13293 gnd.n1888 gnd.n1877 9.3005
R13294 gnd.n1963 gnd.n1841 9.3005
R13295 gnd.n4275 gnd.n4274 9.3005
R13296 gnd.n4270 gnd.n4269 9.3005
R13297 gnd.n4268 gnd.n1973 9.3005
R13298 gnd.n4267 gnd.n4266 9.3005
R13299 gnd.n4265 gnd.n1974 9.3005
R13300 gnd.n4264 gnd.n4263 9.3005
R13301 gnd.n4262 gnd.n1981 9.3005
R13302 gnd.n4261 gnd.n4260 9.3005
R13303 gnd.n4259 gnd.n1982 9.3005
R13304 gnd.n4258 gnd.n4257 9.3005
R13305 gnd.n4256 gnd.n1993 9.3005
R13306 gnd.n3386 gnd.n3385 9.3005
R13307 gnd.n3387 gnd.n2557 9.3005
R13308 gnd.n3390 gnd.n3389 9.3005
R13309 gnd.n3388 gnd.n2558 9.3005
R13310 gnd.n2535 gnd.n2534 9.3005
R13311 gnd.n3416 gnd.n3415 9.3005
R13312 gnd.n3417 gnd.n2532 9.3005
R13313 gnd.n3420 gnd.n3419 9.3005
R13314 gnd.n3418 gnd.n2533 9.3005
R13315 gnd.n2511 gnd.n2510 9.3005
R13316 gnd.n3451 gnd.n3450 9.3005
R13317 gnd.n3452 gnd.n2508 9.3005
R13318 gnd.n3457 gnd.n3456 9.3005
R13319 gnd.n3455 gnd.n2509 9.3005
R13320 gnd.n3454 gnd.n3453 9.3005
R13321 gnd.n2487 gnd.n2486 9.3005
R13322 gnd.n3553 gnd.n3552 9.3005
R13323 gnd.n3554 gnd.n2484 9.3005
R13324 gnd.n3557 gnd.n3556 9.3005
R13325 gnd.n3555 gnd.n2485 9.3005
R13326 gnd.n2464 gnd.n2463 9.3005
R13327 gnd.n3613 gnd.n3612 9.3005
R13328 gnd.n3614 gnd.n2462 9.3005
R13329 gnd.n3616 gnd.n3615 9.3005
R13330 gnd.n2443 gnd.n2442 9.3005
R13331 gnd.n3642 gnd.n3641 9.3005
R13332 gnd.n3643 gnd.n2440 9.3005
R13333 gnd.n3649 gnd.n3648 9.3005
R13334 gnd.n3647 gnd.n2441 9.3005
R13335 gnd.n3646 gnd.n3645 9.3005
R13336 gnd.n2408 gnd.n2407 9.3005
R13337 gnd.n3702 gnd.n3701 9.3005
R13338 gnd.n3703 gnd.n2405 9.3005
R13339 gnd.n3706 gnd.n3705 9.3005
R13340 gnd.n3704 gnd.n2406 9.3005
R13341 gnd.n2383 gnd.n2382 9.3005
R13342 gnd.n3756 gnd.n3755 9.3005
R13343 gnd.n3757 gnd.n2380 9.3005
R13344 gnd.n3771 gnd.n3770 9.3005
R13345 gnd.n3769 gnd.n2381 9.3005
R13346 gnd.n3768 gnd.n3767 9.3005
R13347 gnd.n3766 gnd.n3758 9.3005
R13348 gnd.n3765 gnd.n3764 9.3005
R13349 gnd.n3763 gnd.n3762 9.3005
R13350 gnd.n2337 gnd.n2336 9.3005
R13351 gnd.n3856 gnd.n3855 9.3005
R13352 gnd.n3857 gnd.n2334 9.3005
R13353 gnd.n3860 gnd.n3859 9.3005
R13354 gnd.n3858 gnd.n2335 9.3005
R13355 gnd.n2315 gnd.n2314 9.3005
R13356 gnd.n3885 gnd.n3884 9.3005
R13357 gnd.n3886 gnd.n2313 9.3005
R13358 gnd.n3888 gnd.n3887 9.3005
R13359 gnd.n2271 gnd.n2270 9.3005
R13360 gnd.n3929 gnd.n3928 9.3005
R13361 gnd.n3930 gnd.n2268 9.3005
R13362 gnd.n3948 gnd.n3947 9.3005
R13363 gnd.n3946 gnd.n2269 9.3005
R13364 gnd.n3945 gnd.n3944 9.3005
R13365 gnd.n3943 gnd.n3931 9.3005
R13366 gnd.n3942 gnd.n3941 9.3005
R13367 gnd.n3940 gnd.n3937 9.3005
R13368 gnd.n3939 gnd.n3938 9.3005
R13369 gnd.n2041 gnd.n2040 9.3005
R13370 gnd.n4168 gnd.n4167 9.3005
R13371 gnd.n4169 gnd.n2039 9.3005
R13372 gnd.n4171 gnd.n4170 9.3005
R13373 gnd.n2030 gnd.n2029 9.3005
R13374 gnd.n4189 gnd.n4188 9.3005
R13375 gnd.n4190 gnd.n2028 9.3005
R13376 gnd.n4192 gnd.n4191 9.3005
R13377 gnd.n2018 gnd.n2017 9.3005
R13378 gnd.n4210 gnd.n4209 9.3005
R13379 gnd.n4211 gnd.n2016 9.3005
R13380 gnd.n4213 gnd.n4212 9.3005
R13381 gnd.n2006 gnd.n2005 9.3005
R13382 gnd.n4231 gnd.n4230 9.3005
R13383 gnd.n4232 gnd.n2004 9.3005
R13384 gnd.n4235 gnd.n4234 9.3005
R13385 gnd.n4233 gnd.n1995 9.3005
R13386 gnd.n4253 gnd.n1994 9.3005
R13387 gnd.n4255 gnd.n4254 9.3005
R13388 gnd.n2560 gnd.n2559 9.3005
R13389 gnd.n3237 gnd.n3236 9.3005
R13390 gnd.n3238 gnd.n2645 9.3005
R13391 gnd.n3240 gnd.n3239 9.3005
R13392 gnd.n3242 gnd.n3241 9.3005
R13393 gnd.n3243 gnd.n2638 9.3005
R13394 gnd.n3245 gnd.n3244 9.3005
R13395 gnd.n3246 gnd.n2637 9.3005
R13396 gnd.n3248 gnd.n3247 9.3005
R13397 gnd.n3249 gnd.n2631 9.3005
R13398 gnd.n3235 gnd.n3234 9.3005
R13399 gnd.n2732 gnd.n2731 9.3005
R13400 gnd.n3092 gnd.n3091 9.3005
R13401 gnd.n3093 gnd.n2730 9.3005
R13402 gnd.n3095 gnd.n3094 9.3005
R13403 gnd.n2726 gnd.n2725 9.3005
R13404 gnd.n3108 gnd.n3107 9.3005
R13405 gnd.n3109 gnd.n2724 9.3005
R13406 gnd.n3111 gnd.n3110 9.3005
R13407 gnd.n2719 gnd.n2718 9.3005
R13408 gnd.n3124 gnd.n3123 9.3005
R13409 gnd.n3125 gnd.n2717 9.3005
R13410 gnd.n3127 gnd.n3126 9.3005
R13411 gnd.n2712 gnd.n2711 9.3005
R13412 gnd.n3140 gnd.n3139 9.3005
R13413 gnd.n3141 gnd.n2710 9.3005
R13414 gnd.n3143 gnd.n3142 9.3005
R13415 gnd.n2705 gnd.n2704 9.3005
R13416 gnd.n3156 gnd.n3155 9.3005
R13417 gnd.n3157 gnd.n2703 9.3005
R13418 gnd.n3159 gnd.n3158 9.3005
R13419 gnd.n2698 gnd.n2697 9.3005
R13420 gnd.n3173 gnd.n3172 9.3005
R13421 gnd.n3174 gnd.n2696 9.3005
R13422 gnd.n3176 gnd.n3175 9.3005
R13423 gnd.n2691 gnd.n2689 9.3005
R13424 gnd.n3194 gnd.n3193 9.3005
R13425 gnd.n3192 gnd.n2690 9.3005
R13426 gnd.n3191 gnd.n3190 9.3005
R13427 gnd.n2630 gnd.n2628 9.3005
R13428 gnd.n3256 gnd.n3255 9.3005
R13429 gnd.n3254 gnd.n2629 9.3005
R13430 gnd.n3253 gnd.n2623 9.3005
R13431 gnd.n3251 gnd.n3250 9.3005
R13432 gnd.n2633 gnd.n2632 9.3005
R13433 gnd.n2663 gnd.n2662 9.3005
R13434 gnd.n2616 gnd.n2615 9.3005
R13435 gnd.n3337 gnd.n3336 9.3005
R13436 gnd.n3339 gnd.n3338 9.3005
R13437 gnd.n2606 gnd.n2605 9.3005
R13438 gnd.n3345 gnd.n3344 9.3005
R13439 gnd.n3347 gnd.n3346 9.3005
R13440 gnd.n2598 gnd.n2597 9.3005
R13441 gnd.n3353 gnd.n3352 9.3005
R13442 gnd.n3355 gnd.n3354 9.3005
R13443 gnd.n2588 gnd.n2587 9.3005
R13444 gnd.n3361 gnd.n3360 9.3005
R13445 gnd.n3363 gnd.n3362 9.3005
R13446 gnd.n2580 gnd.n2579 9.3005
R13447 gnd.n3369 gnd.n3368 9.3005
R13448 gnd.n3371 gnd.n3370 9.3005
R13449 gnd.n2576 gnd.n2574 9.3005
R13450 gnd.n3374 gnd.n2568 9.3005
R13451 gnd.n3373 gnd.n3372 9.3005
R13452 gnd.n2575 gnd.n2573 9.3005
R13453 gnd.n3367 gnd.n3366 9.3005
R13454 gnd.n3365 gnd.n3364 9.3005
R13455 gnd.n2584 gnd.n2583 9.3005
R13456 gnd.n3359 gnd.n3358 9.3005
R13457 gnd.n3357 gnd.n3356 9.3005
R13458 gnd.n2594 gnd.n2593 9.3005
R13459 gnd.n3351 gnd.n3350 9.3005
R13460 gnd.n3349 gnd.n3348 9.3005
R13461 gnd.n2602 gnd.n2601 9.3005
R13462 gnd.n3343 gnd.n3342 9.3005
R13463 gnd.n3341 gnd.n3340 9.3005
R13464 gnd.n2612 gnd.n2611 9.3005
R13465 gnd.n3335 gnd.n3334 9.3005
R13466 gnd.n3333 gnd.n2620 9.3005
R13467 gnd.n3332 gnd.n2622 9.3005
R13468 gnd.n3381 gnd.n3380 9.3005
R13469 gnd.n3379 gnd.n2567 9.3005
R13470 gnd.n2544 gnd.n2543 9.3005
R13471 gnd.n3407 gnd.n3406 9.3005
R13472 gnd.n3408 gnd.n2541 9.3005
R13473 gnd.n3411 gnd.n3410 9.3005
R13474 gnd.n3409 gnd.n2542 9.3005
R13475 gnd.n2518 gnd.n2517 9.3005
R13476 gnd.n3443 gnd.n3442 9.3005
R13477 gnd.n3444 gnd.n2516 9.3005
R13478 gnd.n3446 gnd.n3445 9.3005
R13479 gnd.n2503 gnd.n2502 9.3005
R13480 gnd.n3463 gnd.n3462 9.3005
R13481 gnd.n3464 gnd.n2500 9.3005
R13482 gnd.n3467 gnd.n3466 9.3005
R13483 gnd.n3465 gnd.n2501 9.3005
R13484 gnd.n1531 gnd.n1529 9.3005
R13485 gnd.n4723 gnd.n4722 9.3005
R13486 gnd.n4721 gnd.n1530 9.3005
R13487 gnd.n4720 gnd.n4719 9.3005
R13488 gnd.n4718 gnd.n1532 9.3005
R13489 gnd.n4717 gnd.n4716 9.3005
R13490 gnd.n4715 gnd.n1536 9.3005
R13491 gnd.n4714 gnd.n4713 9.3005
R13492 gnd.n4712 gnd.n1537 9.3005
R13493 gnd.n4711 gnd.n4710 9.3005
R13494 gnd.n4709 gnd.n1541 9.3005
R13495 gnd.n4708 gnd.n4707 9.3005
R13496 gnd.n4706 gnd.n1542 9.3005
R13497 gnd.n4705 gnd.n4704 9.3005
R13498 gnd.n4703 gnd.n1546 9.3005
R13499 gnd.n4702 gnd.n4701 9.3005
R13500 gnd.n4700 gnd.n1547 9.3005
R13501 gnd.n4699 gnd.n4698 9.3005
R13502 gnd.n4697 gnd.n1551 9.3005
R13503 gnd.n4696 gnd.n4695 9.3005
R13504 gnd.n4694 gnd.n1552 9.3005
R13505 gnd.n4693 gnd.n4692 9.3005
R13506 gnd.n4691 gnd.n1556 9.3005
R13507 gnd.n4690 gnd.n4689 9.3005
R13508 gnd.n4688 gnd.n1557 9.3005
R13509 gnd.n4687 gnd.n4686 9.3005
R13510 gnd.n4685 gnd.n1561 9.3005
R13511 gnd.n4684 gnd.n4683 9.3005
R13512 gnd.n4682 gnd.n1562 9.3005
R13513 gnd.n4681 gnd.n4680 9.3005
R13514 gnd.n4679 gnd.n1566 9.3005
R13515 gnd.n4678 gnd.n4677 9.3005
R13516 gnd.n4676 gnd.n1567 9.3005
R13517 gnd.n4675 gnd.n4674 9.3005
R13518 gnd.n4673 gnd.n1571 9.3005
R13519 gnd.n4672 gnd.n4671 9.3005
R13520 gnd.n4670 gnd.n1572 9.3005
R13521 gnd.n4669 gnd.n4668 9.3005
R13522 gnd.n4667 gnd.n1576 9.3005
R13523 gnd.n4666 gnd.n4665 9.3005
R13524 gnd.n4664 gnd.n1577 9.3005
R13525 gnd.n4663 gnd.n4662 9.3005
R13526 gnd.n4661 gnd.n1581 9.3005
R13527 gnd.n4660 gnd.n4659 9.3005
R13528 gnd.n4658 gnd.n1582 9.3005
R13529 gnd.n4657 gnd.n4656 9.3005
R13530 gnd.n4655 gnd.n1586 9.3005
R13531 gnd.n4654 gnd.n4653 9.3005
R13532 gnd.n4652 gnd.n1587 9.3005
R13533 gnd.n4651 gnd.n4650 9.3005
R13534 gnd.n4649 gnd.n1591 9.3005
R13535 gnd.n4648 gnd.n4647 9.3005
R13536 gnd.n4646 gnd.n1592 9.3005
R13537 gnd.n4645 gnd.n4644 9.3005
R13538 gnd.n4643 gnd.n1596 9.3005
R13539 gnd.n4642 gnd.n4641 9.3005
R13540 gnd.n4640 gnd.n1597 9.3005
R13541 gnd.n4639 gnd.n4638 9.3005
R13542 gnd.n4637 gnd.n1601 9.3005
R13543 gnd.n4636 gnd.n4635 9.3005
R13544 gnd.n4634 gnd.n1602 9.3005
R13545 gnd.n4633 gnd.n4632 9.3005
R13546 gnd.n4631 gnd.n1606 9.3005
R13547 gnd.n4630 gnd.n4629 9.3005
R13548 gnd.n4628 gnd.n1607 9.3005
R13549 gnd.n4627 gnd.n1610 9.3005
R13550 gnd.n3378 gnd.n2566 9.3005
R13551 gnd.n1883 gnd.n1879 9.3005
R13552 gnd.n1654 gnd.n1652 9.3005
R13553 gnd.n4601 gnd.n4600 9.3005
R13554 gnd.n4599 gnd.n1653 9.3005
R13555 gnd.n4598 gnd.n4597 9.3005
R13556 gnd.n4596 gnd.n1655 9.3005
R13557 gnd.n4595 gnd.n4594 9.3005
R13558 gnd.n4593 gnd.n1659 9.3005
R13559 gnd.n4592 gnd.n4591 9.3005
R13560 gnd.n4590 gnd.n1660 9.3005
R13561 gnd.n4589 gnd.n4588 9.3005
R13562 gnd.n4587 gnd.n1664 9.3005
R13563 gnd.n4586 gnd.n4585 9.3005
R13564 gnd.n4584 gnd.n1665 9.3005
R13565 gnd.n4583 gnd.n4582 9.3005
R13566 gnd.n4581 gnd.n1669 9.3005
R13567 gnd.n4580 gnd.n4579 9.3005
R13568 gnd.n4578 gnd.n1670 9.3005
R13569 gnd.n4577 gnd.n4576 9.3005
R13570 gnd.n4575 gnd.n1674 9.3005
R13571 gnd.n4574 gnd.n4573 9.3005
R13572 gnd.n4572 gnd.n1675 9.3005
R13573 gnd.n4571 gnd.n4570 9.3005
R13574 gnd.n4569 gnd.n1679 9.3005
R13575 gnd.n4568 gnd.n4567 9.3005
R13576 gnd.n4566 gnd.n1680 9.3005
R13577 gnd.n4565 gnd.n4564 9.3005
R13578 gnd.n318 gnd.n316 9.3005
R13579 gnd.n7411 gnd.n7410 9.3005
R13580 gnd.n7409 gnd.n317 9.3005
R13581 gnd.n7408 gnd.n7407 9.3005
R13582 gnd.n7406 gnd.n319 9.3005
R13583 gnd.n7405 gnd.n7404 9.3005
R13584 gnd.n7403 gnd.n323 9.3005
R13585 gnd.n7402 gnd.n7401 9.3005
R13586 gnd.n7400 gnd.n324 9.3005
R13587 gnd.n294 gnd.n293 9.3005
R13588 gnd.n7425 gnd.n7424 9.3005
R13589 gnd.n7426 gnd.n292 9.3005
R13590 gnd.n7428 gnd.n7427 9.3005
R13591 gnd.n278 gnd.n277 9.3005
R13592 gnd.n7441 gnd.n7440 9.3005
R13593 gnd.n7442 gnd.n276 9.3005
R13594 gnd.n7444 gnd.n7443 9.3005
R13595 gnd.n263 gnd.n262 9.3005
R13596 gnd.n7457 gnd.n7456 9.3005
R13597 gnd.n7458 gnd.n261 9.3005
R13598 gnd.n7460 gnd.n7459 9.3005
R13599 gnd.n247 gnd.n246 9.3005
R13600 gnd.n7473 gnd.n7472 9.3005
R13601 gnd.n7474 gnd.n245 9.3005
R13602 gnd.n7476 gnd.n7475 9.3005
R13603 gnd.n233 gnd.n232 9.3005
R13604 gnd.n7489 gnd.n7488 9.3005
R13605 gnd.n7490 gnd.n231 9.3005
R13606 gnd.n7492 gnd.n7491 9.3005
R13607 gnd.n218 gnd.n217 9.3005
R13608 gnd.n7505 gnd.n7504 9.3005
R13609 gnd.n7506 gnd.n215 9.3005
R13610 gnd.n7576 gnd.n7575 9.3005
R13611 gnd.n7574 gnd.n216 9.3005
R13612 gnd.n7573 gnd.n7572 9.3005
R13613 gnd.n7571 gnd.n7507 9.3005
R13614 gnd.n7570 gnd.n7569 9.3005
R13615 gnd.n1885 gnd.n1884 9.3005
R13616 gnd.n7566 gnd.n7509 9.3005
R13617 gnd.n7565 gnd.n7564 9.3005
R13618 gnd.n7563 gnd.n7514 9.3005
R13619 gnd.n7562 gnd.n7561 9.3005
R13620 gnd.n7560 gnd.n7515 9.3005
R13621 gnd.n7559 gnd.n7558 9.3005
R13622 gnd.n7557 gnd.n7522 9.3005
R13623 gnd.n7556 gnd.n7555 9.3005
R13624 gnd.n7554 gnd.n7523 9.3005
R13625 gnd.n7553 gnd.n7552 9.3005
R13626 gnd.n7551 gnd.n7530 9.3005
R13627 gnd.n7550 gnd.n7549 9.3005
R13628 gnd.n7548 gnd.n7531 9.3005
R13629 gnd.n7547 gnd.n7546 9.3005
R13630 gnd.n7545 gnd.n7538 9.3005
R13631 gnd.n7544 gnd.n7543 9.3005
R13632 gnd.n120 gnd.n117 9.3005
R13633 gnd.n7670 gnd.n7669 9.3005
R13634 gnd.n7568 gnd.n7567 9.3005
R13635 gnd.n4280 gnd.n1836 9.3005
R13636 gnd.n4282 gnd.n4281 9.3005
R13637 gnd.n1831 gnd.n1830 9.3005
R13638 gnd.n4340 gnd.n4339 9.3005
R13639 gnd.n4341 gnd.n1828 9.3005
R13640 gnd.n4344 gnd.n4343 9.3005
R13641 gnd.n4342 gnd.n1829 9.3005
R13642 gnd.n1793 gnd.n1792 9.3005
R13643 gnd.n4372 gnd.n4371 9.3005
R13644 gnd.n4373 gnd.n1790 9.3005
R13645 gnd.n4376 gnd.n4375 9.3005
R13646 gnd.n4374 gnd.n1791 9.3005
R13647 gnd.n1767 gnd.n1766 9.3005
R13648 gnd.n4404 gnd.n4403 9.3005
R13649 gnd.n4405 gnd.n1764 9.3005
R13650 gnd.n4408 gnd.n4407 9.3005
R13651 gnd.n4406 gnd.n1765 9.3005
R13652 gnd.n1741 gnd.n1740 9.3005
R13653 gnd.n4436 gnd.n4435 9.3005
R13654 gnd.n4437 gnd.n1738 9.3005
R13655 gnd.n4446 gnd.n4445 9.3005
R13656 gnd.n4444 gnd.n1739 9.3005
R13657 gnd.n4443 gnd.n4442 9.3005
R13658 gnd.n4441 gnd.n4438 9.3005
R13659 gnd.n1693 gnd.n1691 9.3005
R13660 gnd.n4557 gnd.n4556 9.3005
R13661 gnd.n4555 gnd.n1692 9.3005
R13662 gnd.n4554 gnd.n4553 9.3005
R13663 gnd.n4552 gnd.n1694 9.3005
R13664 gnd.n4551 gnd.n4550 9.3005
R13665 gnd.n4549 gnd.n75 9.3005
R13666 gnd.n7719 gnd.n76 9.3005
R13667 gnd.n7718 gnd.n7717 9.3005
R13668 gnd.n7716 gnd.n77 9.3005
R13669 gnd.n7715 gnd.n7714 9.3005
R13670 gnd.n7713 gnd.n81 9.3005
R13671 gnd.n7712 gnd.n7711 9.3005
R13672 gnd.n7710 gnd.n82 9.3005
R13673 gnd.n7709 gnd.n7708 9.3005
R13674 gnd.n7707 gnd.n86 9.3005
R13675 gnd.n7706 gnd.n7705 9.3005
R13676 gnd.n7704 gnd.n87 9.3005
R13677 gnd.n7703 gnd.n7702 9.3005
R13678 gnd.n7701 gnd.n91 9.3005
R13679 gnd.n7700 gnd.n7699 9.3005
R13680 gnd.n7698 gnd.n92 9.3005
R13681 gnd.n7697 gnd.n7696 9.3005
R13682 gnd.n7695 gnd.n96 9.3005
R13683 gnd.n7694 gnd.n7693 9.3005
R13684 gnd.n7692 gnd.n97 9.3005
R13685 gnd.n7691 gnd.n7690 9.3005
R13686 gnd.n7689 gnd.n101 9.3005
R13687 gnd.n7688 gnd.n7687 9.3005
R13688 gnd.n7686 gnd.n102 9.3005
R13689 gnd.n7685 gnd.n7684 9.3005
R13690 gnd.n7683 gnd.n106 9.3005
R13691 gnd.n7682 gnd.n7681 9.3005
R13692 gnd.n7680 gnd.n107 9.3005
R13693 gnd.n7679 gnd.n7678 9.3005
R13694 gnd.n7677 gnd.n111 9.3005
R13695 gnd.n7676 gnd.n7675 9.3005
R13696 gnd.n7674 gnd.n112 9.3005
R13697 gnd.n7673 gnd.n7672 9.3005
R13698 gnd.n7671 gnd.n116 9.3005
R13699 gnd.n4279 gnd.n4278 9.3005
R13700 gnd.t17 gnd.n5256 9.24152
R13701 gnd.n6417 gnd.t107 9.24152
R13702 gnd.n6518 gnd.t125 9.24152
R13703 gnd.n4984 gnd.t233 9.24152
R13704 gnd.t194 gnd.n1198 9.24152
R13705 gnd.n4879 gnd.t190 9.24152
R13706 gnd.t206 gnd.n1761 9.24152
R13707 gnd.n7380 gnd.t196 9.24152
R13708 gnd.n259 gnd.t200 9.24152
R13709 gnd.t72 gnd.t17 8.92286
R13710 gnd.n3601 gnd.n2473 8.92286
R13711 gnd.n3569 gnd.n2436 8.92286
R13712 gnd.n3680 gnd.t21 8.92286
R13713 gnd.n3698 gnd.t2 8.92286
R13714 gnd.n3777 gnd.n2375 8.92286
R13715 gnd.n3834 gnd.n2354 8.92286
R13716 gnd.t24 gnd.n2317 8.92286
R13717 gnd.t0 gnd.n3898 8.92286
R13718 gnd.n3926 gnd.n3924 8.92286
R13719 gnd.n3974 gnd.n2245 8.92286
R13720 gnd.n6391 gnd.n6366 8.92171
R13721 gnd.n6359 gnd.n6334 8.92171
R13722 gnd.n6327 gnd.n6302 8.92171
R13723 gnd.n6296 gnd.n6271 8.92171
R13724 gnd.n6264 gnd.n6239 8.92171
R13725 gnd.n6232 gnd.n6207 8.92171
R13726 gnd.n6200 gnd.n6175 8.92171
R13727 gnd.n6169 gnd.n6144 8.92171
R13728 gnd.n4020 gnd.n4002 8.72777
R13729 gnd.t8 gnd.n5363 8.60421
R13730 gnd.n5008 gnd.t258 8.60421
R13731 gnd.n4855 gnd.t198 8.60421
R13732 gnd.t37 gnd.n3775 8.60421
R13733 gnd.n3824 gnd.t29 8.60421
R13734 gnd.n4359 gnd.t287 8.60421
R13735 gnd.n229 gnd.t283 8.60421
R13736 gnd.n5327 gnd.n5307 8.43467
R13737 gnd.n54 gnd.n34 8.43467
R13738 gnd.n3078 gnd.n0 8.41456
R13739 gnd.n7720 gnd.n7719 8.41456
R13740 gnd.n3592 gnd.n2480 8.28555
R13741 gnd.n3661 gnd.n3660 8.28555
R13742 gnd.n3726 gnd.n3725 8.28555
R13743 gnd.n3845 gnd.n2339 8.28555
R13744 gnd.n3891 gnd.n2279 8.28555
R13745 gnd.n3998 gnd.n2230 8.28555
R13746 gnd.n6392 gnd.n6364 8.14595
R13747 gnd.n6360 gnd.n6332 8.14595
R13748 gnd.n6328 gnd.n6300 8.14595
R13749 gnd.n6297 gnd.n6269 8.14595
R13750 gnd.n6265 gnd.n6237 8.14595
R13751 gnd.n6233 gnd.n6205 8.14595
R13752 gnd.n6201 gnd.n6173 8.14595
R13753 gnd.n6170 gnd.n6142 8.14595
R13754 gnd.n6397 gnd.n6396 7.97301
R13755 gnd.n5856 gnd.t10 7.9669
R13756 gnd.t158 gnd.t31 7.9669
R13757 gnd.n7669 gnd.n120 7.75808
R13758 gnd.n4275 gnd.n1841 7.75808
R13759 gnd.n3333 gnd.n3332 7.75808
R13760 gnd.n2939 gnd.n2936 7.75808
R13761 gnd.n3559 gnd.n2480 7.64824
R13762 gnd.n3660 gnd.n2428 7.64824
R13763 gnd.n3724 gnd.t59 7.64824
R13764 gnd.n3726 gnd.n3724 7.64824
R13765 gnd.n3853 gnd.n2339 7.64824
R13766 gnd.n3853 gnd.t43 7.64824
R13767 gnd.n3891 gnd.n3890 7.64824
R13768 gnd.t14 gnd.n5449 7.32958
R13769 gnd.n1519 gnd.n1518 7.30353
R13770 gnd.n4019 gnd.n4018 7.30353
R13771 gnd.n5758 gnd.n5757 7.01093
R13772 gnd.n5768 gnd.n5478 7.01093
R13773 gnd.n5767 gnd.n5481 7.01093
R13774 gnd.n5776 gnd.n5472 7.01093
R13775 gnd.n5780 gnd.n5779 7.01093
R13776 gnd.n5798 gnd.n5457 7.01093
R13777 gnd.n5797 gnd.n5460 7.01093
R13778 gnd.n5808 gnd.n5449 7.01093
R13779 gnd.n5450 gnd.n5438 7.01093
R13780 gnd.n5821 gnd.n5439 7.01093
R13781 gnd.n5832 gnd.n5431 7.01093
R13782 gnd.n5831 gnd.n5422 7.01093
R13783 gnd.n5424 gnd.n5406 7.01093
R13784 gnd.n5868 gnd.n5407 7.01093
R13785 gnd.n5857 gnd.n5856 7.01093
R13786 gnd.n5893 gnd.n5398 7.01093
R13787 gnd.n5904 gnd.n5903 7.01093
R13788 gnd.n5391 gnd.n5383 7.01093
R13789 gnd.n5933 gnd.n5371 7.01093
R13790 gnd.n5932 gnd.n5374 7.01093
R13791 gnd.n5943 gnd.n5363 7.01093
R13792 gnd.n5364 gnd.n5352 7.01093
R13793 gnd.n5954 gnd.n5353 7.01093
R13794 gnd.n5978 gnd.n5284 7.01093
R13795 gnd.n5977 gnd.n5275 7.01093
R13796 gnd.n5277 gnd.n5268 7.01093
R13797 gnd.n6000 gnd.n5999 7.01093
R13798 gnd.n6018 gnd.n5256 7.01093
R13799 gnd.n6017 gnd.n5259 7.01093
R13800 gnd.n6028 gnd.n5248 7.01093
R13801 gnd.n5249 gnd.n5236 7.01093
R13802 gnd.n6039 gnd.n5237 7.01093
R13803 gnd.n6075 gnd.n6074 7.01093
R13804 gnd.n6057 gnd.n5214 7.01093
R13805 gnd.n6086 gnd.n6085 7.01093
R13806 gnd.n6103 gnd.n5202 7.01093
R13807 gnd.n6102 gnd.n5205 7.01093
R13808 gnd.n6114 gnd.n5194 7.01093
R13809 gnd.n6123 gnd.n5185 7.01093
R13810 gnd.n6136 gnd.n6135 7.01093
R13811 gnd.n6526 gnd.n973 7.01093
R13812 gnd.n6525 gnd.n976 7.01093
R13813 gnd.n6418 gnd.n6417 7.01093
R13814 gnd.n6519 gnd.n6518 7.01093
R13815 gnd.n6411 gnd.n6410 7.01093
R13816 gnd.n6512 gnd.n996 7.01093
R13817 gnd.n3601 gnd.n3600 7.01093
R13818 gnd.n3569 gnd.n2446 7.01093
R13819 gnd.n3777 gnd.n3776 7.01093
R13820 gnd.n3835 gnd.n3834 7.01093
R13821 gnd.n3924 gnd.n2275 7.01093
R13822 gnd.n3974 gnd.n2244 7.01093
R13823 gnd.t171 gnd.n2239 7.01093
R13824 gnd.n5439 gnd.t6 6.69227
R13825 gnd.n5999 gnd.t72 6.69227
R13826 gnd.t5 gnd.n5184 6.69227
R13827 gnd.n3586 gnd.t66 6.69227
R13828 gnd.t44 gnd.n3983 6.69227
R13829 gnd.n4155 gnd.n4154 6.5566
R13830 gnd.n3488 gnd.n3487 6.5566
R13831 gnd.n4737 gnd.n4733 6.5566
R13832 gnd.n4030 gnd.n4029 6.5566
R13833 gnd.n3550 gnd.n3549 6.37362
R13834 gnd.t111 gnd.n3585 6.37362
R13835 gnd.n3639 gnd.t40 6.37362
R13836 gnd.n3691 gnd.n3690 6.37362
R13837 gnd.n3743 gnd.t59 6.37362
R13838 gnd.t43 gnd.n3852 6.37362
R13839 gnd.n3899 gnd.n2293 6.37362
R13840 gnd.n2304 gnd.t50 6.37362
R13841 gnd.n3984 gnd.t91 6.37362
R13842 gnd.n4165 gnd.n2043 6.37362
R13843 gnd.n3239 gnd.n2644 6.20656
R13844 gnd.n7631 gnd.n7628 6.20656
R13845 gnd.n5071 gnd.n5070 6.20656
R13846 gnd.n4260 gnd.n1985 6.20656
R13847 gnd.n5892 gnd.t35 6.05496
R13848 gnd.n5891 gnd.t16 6.05496
R13849 gnd.t60 gnd.n5364 6.05496
R13850 gnd.n6064 gnd.t12 6.05496
R13851 gnd.n3776 gnd.t37 6.05496
R13852 gnd.n3835 gnd.t29 6.05496
R13853 gnd.n6394 gnd.n6364 5.81868
R13854 gnd.n6362 gnd.n6332 5.81868
R13855 gnd.n6330 gnd.n6300 5.81868
R13856 gnd.n6299 gnd.n6269 5.81868
R13857 gnd.n6267 gnd.n6237 5.81868
R13858 gnd.n6235 gnd.n6205 5.81868
R13859 gnd.n6203 gnd.n6173 5.81868
R13860 gnd.n6172 gnd.n6142 5.81868
R13861 gnd.n3619 gnd.n2459 5.73631
R13862 gnd.n3632 gnd.n2450 5.73631
R13863 gnd.n3715 gnd.n3714 5.73631
R13864 gnd.n3796 gnd.n3795 5.73631
R13865 gnd.n3958 gnd.n2258 5.73631
R13866 gnd.n2297 gnd.n2261 5.73631
R13867 gnd.n2245 gnd.t171 5.73631
R13868 gnd.n212 gnd.n202 5.73631
R13869 gnd.n4159 gnd.n2219 5.62001
R13870 gnd.n4799 gnd.n1462 5.62001
R13871 gnd.n4799 gnd.n1463 5.62001
R13872 gnd.n4025 gnd.n2219 5.62001
R13873 gnd.n5576 gnd.n5575 5.4308
R13874 gnd.n6433 gnd.n5164 5.4308
R13875 gnd.n5353 gnd.t11 5.41765
R13876 gnd.t18 gnd.n5988 5.41765
R13877 gnd.t79 gnd.n5221 5.41765
R13878 gnd.t64 gnd.n3631 5.41765
R13879 gnd.n3950 gnd.t68 5.41765
R13880 gnd.n3699 gnd.n3698 5.09899
R13881 gnd.n3673 gnd.n3672 5.09899
R13882 gnd.n3871 gnd.n3870 5.09899
R13883 gnd.n3881 gnd.n2317 5.09899
R13884 gnd.t136 gnd.n3997 5.09899
R13885 gnd.n6392 gnd.n6391 5.04292
R13886 gnd.n6360 gnd.n6359 5.04292
R13887 gnd.n6328 gnd.n6327 5.04292
R13888 gnd.n6297 gnd.n6296 5.04292
R13889 gnd.n6265 gnd.n6264 5.04292
R13890 gnd.n6233 gnd.n6232 5.04292
R13891 gnd.n6201 gnd.n6200 5.04292
R13892 gnd.n6170 gnd.n6169 5.04292
R13893 gnd.n5347 gnd.n5346 4.82753
R13894 gnd.n74 gnd.n73 4.82753
R13895 gnd.t3 gnd.n5914 4.78034
R13896 gnd.n6028 gnd.t9 4.78034
R13897 gnd.t25 gnd.n2538 4.78034
R13898 gnd.n3632 gnd.t64 4.78034
R13899 gnd.t68 gnd.n2258 4.78034
R13900 gnd.n4162 gnd.t158 4.78034
R13901 gnd.n4215 gnd.t19 4.78034
R13902 gnd.n5888 gnd.n5887 4.74817
R13903 gnd.n5883 gnd.n5882 4.74817
R13904 gnd.n5879 gnd.n5878 4.74817
R13905 gnd.n5875 gnd.n5350 4.74817
R13906 gnd.n5887 gnd.n5886 4.74817
R13907 gnd.n5885 gnd.n5883 4.74817
R13908 gnd.n5881 gnd.n5879 4.74817
R13909 gnd.n5877 gnd.n5875 4.74817
R13910 gnd.n7417 gnd.n7416 4.74817
R13911 gnd.n4544 gnd.n306 4.74817
R13912 gnd.n1702 gnd.n305 4.74817
R13913 gnd.n330 gnd.n304 4.74817
R13914 gnd.n7396 gnd.n303 4.74817
R13915 gnd.n7417 gnd.n307 4.74817
R13916 gnd.n7415 gnd.n306 4.74817
R13917 gnd.n4545 gnd.n305 4.74817
R13918 gnd.n1701 gnd.n304 4.74817
R13919 gnd.n331 gnd.n303 4.74817
R13920 gnd.n2853 gnd.n2852 4.74817
R13921 gnd.n2850 gnd.n2775 4.74817
R13922 gnd.n2843 gnd.n2774 4.74817
R13923 gnd.n2839 gnd.n2773 4.74817
R13924 gnd.n2835 gnd.n2772 4.74817
R13925 gnd.n4464 gnd.n4463 4.74817
R13926 gnd.n4534 gnd.n1707 4.74817
R13927 gnd.n4539 gnd.n4536 4.74817
R13928 gnd.n4537 gnd.n336 4.74817
R13929 gnd.n7390 gnd.n7389 4.74817
R13930 gnd.n4465 gnd.n4464 4.74817
R13931 gnd.n4461 gnd.n1707 4.74817
R13932 gnd.n4536 gnd.n4535 4.74817
R13933 gnd.n4538 gnd.n4537 4.74817
R13934 gnd.n7391 gnd.n7390 4.74817
R13935 gnd.n4945 gnd.n4944 4.74817
R13936 gnd.n1244 gnd.n1226 4.74817
R13937 gnd.n4932 gnd.n4931 4.74817
R13938 gnd.n1261 gnd.n1245 4.74817
R13939 gnd.n4919 gnd.n4918 4.74817
R13940 gnd.n4946 gnd.n4945 4.74817
R13941 gnd.n4943 gnd.n1226 4.74817
R13942 gnd.n4933 gnd.n4932 4.74817
R13943 gnd.n4930 gnd.n1245 4.74817
R13944 gnd.n4920 gnd.n4919 4.74817
R13945 gnd.n2852 gnd.n2770 4.74817
R13946 gnd.n2850 gnd.n2849 4.74817
R13947 gnd.n2845 gnd.n2774 4.74817
R13948 gnd.n2842 gnd.n2773 4.74817
R13949 gnd.n2838 gnd.n2772 4.74817
R13950 gnd.n5327 gnd.n5326 4.7074
R13951 gnd.n54 gnd.n53 4.7074
R13952 gnd.n5347 gnd.n5327 4.65959
R13953 gnd.n74 gnd.n54 4.65959
R13954 gnd.n2218 gnd.n2136 4.6132
R13955 gnd.n4800 gnd.n1461 4.6132
R13956 gnd.n3609 gnd.n3608 4.46168
R13957 gnd.n3618 gnd.t53 4.46168
R13958 gnd.n3630 gnd.n3629 4.46168
R13959 gnd.n3787 gnd.n3786 4.46168
R13960 gnd.n3828 gnd.n3827 4.46168
R13961 gnd.n3951 gnd.n2265 4.46168
R13962 gnd.t23 gnd.n3957 4.46168
R13963 gnd.n3967 gnd.n3966 4.46168
R13964 gnd.n4015 gnd.n4002 4.46111
R13965 gnd.n6377 gnd.n6373 4.38594
R13966 gnd.n6345 gnd.n6341 4.38594
R13967 gnd.n6313 gnd.n6309 4.38594
R13968 gnd.n6282 gnd.n6278 4.38594
R13969 gnd.n6250 gnd.n6246 4.38594
R13970 gnd.n6218 gnd.n6214 4.38594
R13971 gnd.n6186 gnd.n6182 4.38594
R13972 gnd.n6155 gnd.n6151 4.38594
R13973 gnd.n6388 gnd.n6366 4.26717
R13974 gnd.n6356 gnd.n6334 4.26717
R13975 gnd.n6324 gnd.n6302 4.26717
R13976 gnd.n6293 gnd.n6271 4.26717
R13977 gnd.n6261 gnd.n6239 4.26717
R13978 gnd.n6229 gnd.n6207 4.26717
R13979 gnd.n6197 gnd.n6175 4.26717
R13980 gnd.n6166 gnd.n6144 4.26717
R13981 gnd.t4 gnd.n5845 4.14303
R13982 gnd.n6103 gnd.t7 4.14303
R13983 gnd.n6396 gnd.n6395 4.08274
R13984 gnd.n4154 gnd.n4153 4.05904
R13985 gnd.n3489 gnd.n3488 4.05904
R13986 gnd.n4740 gnd.n4733 4.05904
R13987 gnd.n4031 gnd.n4030 4.05904
R13988 gnd.n15 gnd.n7 3.99943
R13989 gnd.n6533 gnd.n963 3.82437
R13990 gnd.n4726 gnd.n4725 3.82437
R13991 gnd.n3619 gnd.t84 3.82437
R13992 gnd.t52 gnd.n2428 3.82437
R13993 gnd.n3681 gnd.n2419 3.82437
R13994 gnd.n3732 gnd.n2393 3.82437
R13995 gnd.n3810 gnd.n3809 3.82437
R13996 gnd.n3897 gnd.n2287 3.82437
R13997 gnd.n3890 gnd.t76 3.82437
R13998 gnd.n4093 gnd.n2225 3.82437
R13999 gnd.n6396 gnd.n6268 3.70378
R14000 gnd.n5349 gnd.n5348 3.65935
R14001 gnd.n15 gnd.n14 3.60163
R14002 gnd.t95 gnd.n1094 3.50571
R14003 gnd.n3258 gnd.t115 3.50571
R14004 gnd.n4284 gnd.t103 3.50571
R14005 gnd.n7586 gnd.t99 3.50571
R14006 gnd.n6387 gnd.n6368 3.49141
R14007 gnd.n6355 gnd.n6336 3.49141
R14008 gnd.n6323 gnd.n6304 3.49141
R14009 gnd.n6292 gnd.n6273 3.49141
R14010 gnd.n6260 gnd.n6241 3.49141
R14011 gnd.n6228 gnd.n6209 3.49141
R14012 gnd.n6196 gnd.n6177 3.49141
R14013 gnd.n6165 gnd.n6146 3.49141
R14014 gnd.n6533 gnd.n6532 3.18706
R14015 gnd.n3585 gnd.n3584 3.18706
R14016 gnd.n3734 gnd.t39 3.18706
R14017 gnd.n3752 gnd.n2386 3.18706
R14018 gnd.n3818 gnd.n3817 3.18706
R14019 gnd.n3863 gnd.t42 3.18706
R14020 gnd.n3984 gnd.n2239 3.18706
R14021 gnd.n5846 gnd.t4 2.8684
R14022 gnd.n2497 gnd.t27 2.8684
R14023 gnd.t66 gnd.t111 2.8684
R14024 gnd.t91 gnd.t44 2.8684
R14025 gnd.n4176 gnd.t31 2.8684
R14026 gnd.n5328 gnd.t329 2.82907
R14027 gnd.n5328 gnd.t276 2.82907
R14028 gnd.n5330 gnd.t316 2.82907
R14029 gnd.n5330 gnd.t191 2.82907
R14030 gnd.n5332 gnd.t225 2.82907
R14031 gnd.n5332 gnd.t205 2.82907
R14032 gnd.n5334 gnd.t203 2.82907
R14033 gnd.n5334 gnd.t341 2.82907
R14034 gnd.n5336 gnd.t212 2.82907
R14035 gnd.n5336 gnd.t266 2.82907
R14036 gnd.n5338 gnd.t305 2.82907
R14037 gnd.n5338 gnd.t249 2.82907
R14038 gnd.n5340 gnd.t282 2.82907
R14039 gnd.n5340 gnd.t208 2.82907
R14040 gnd.n5342 gnd.t253 2.82907
R14041 gnd.n5342 gnd.t334 2.82907
R14042 gnd.n5344 gnd.t310 2.82907
R14043 gnd.n5344 gnd.t309 2.82907
R14044 gnd.n5289 gnd.t218 2.82907
R14045 gnd.n5289 gnd.t247 2.82907
R14046 gnd.n5291 gnd.t265 2.82907
R14047 gnd.n5291 gnd.t330 2.82907
R14048 gnd.n5293 gnd.t244 2.82907
R14049 gnd.n5293 gnd.t226 2.82907
R14050 gnd.n5295 gnd.t291 2.82907
R14051 gnd.n5295 gnd.t278 2.82907
R14052 gnd.n5297 gnd.t337 2.82907
R14053 gnd.n5297 gnd.t255 2.82907
R14054 gnd.n5299 gnd.t272 2.82907
R14055 gnd.n5299 gnd.t304 2.82907
R14056 gnd.n5301 gnd.t319 2.82907
R14057 gnd.n5301 gnd.t195 2.82907
R14058 gnd.n5303 gnd.t256 2.82907
R14059 gnd.n5303 gnd.t286 2.82907
R14060 gnd.n5305 gnd.t210 2.82907
R14061 gnd.n5305 gnd.t230 2.82907
R14062 gnd.n5308 gnd.t340 2.82907
R14063 gnd.n5308 gnd.t220 2.82907
R14064 gnd.n5310 gnd.t239 2.82907
R14065 gnd.n5310 gnd.t308 2.82907
R14066 gnd.n5312 gnd.t214 2.82907
R14067 gnd.n5312 gnd.t349 2.82907
R14068 gnd.n5314 gnd.t264 2.82907
R14069 gnd.n5314 gnd.t252 2.82907
R14070 gnd.n5316 gnd.t285 2.82907
R14071 gnd.n5316 gnd.t232 2.82907
R14072 gnd.n5318 gnd.t246 2.82907
R14073 gnd.n5318 gnd.t275 2.82907
R14074 gnd.n5320 gnd.t292 2.82907
R14075 gnd.n5320 gnd.t215 2.82907
R14076 gnd.n5322 gnd.t234 2.82907
R14077 gnd.n5322 gnd.t263 2.82907
R14078 gnd.n5324 gnd.t336 2.82907
R14079 gnd.n5324 gnd.t346 2.82907
R14080 gnd.n71 gnd.t216 2.82907
R14081 gnd.n71 gnd.t235 2.82907
R14082 gnd.n69 gnd.t296 2.82907
R14083 gnd.n69 gnd.t201 2.82907
R14084 gnd.n67 gnd.t327 2.82907
R14085 gnd.n67 gnd.t241 2.82907
R14086 gnd.n65 gnd.t348 2.82907
R14087 gnd.n65 gnd.t261 2.82907
R14088 gnd.n63 gnd.t222 2.82907
R14089 gnd.n63 gnd.t339 2.82907
R14090 gnd.n61 gnd.t311 2.82907
R14091 gnd.n61 gnd.t322 2.82907
R14092 gnd.n59 gnd.t325 2.82907
R14093 gnd.n59 gnd.t345 2.82907
R14094 gnd.n57 gnd.t320 2.82907
R14095 gnd.n57 gnd.t271 2.82907
R14096 gnd.n55 gnd.t237 2.82907
R14097 gnd.n55 gnd.t307 2.82907
R14098 gnd.n32 gnd.t193 2.82907
R14099 gnd.n32 gnd.t224 2.82907
R14100 gnd.n30 gnd.t323 2.82907
R14101 gnd.n30 gnd.t294 2.82907
R14102 gnd.n28 gnd.t197 2.82907
R14103 gnd.n28 gnd.t342 2.82907
R14104 gnd.n26 gnd.t333 2.82907
R14105 gnd.n26 gnd.t312 2.82907
R14106 gnd.n24 gnd.t293 2.82907
R14107 gnd.n24 gnd.t328 2.82907
R14108 gnd.n22 gnd.t318 2.82907
R14109 gnd.n22 gnd.t324 2.82907
R14110 gnd.n20 gnd.t269 2.82907
R14111 gnd.n20 gnd.t228 2.82907
R14112 gnd.n18 gnd.t207 2.82907
R14113 gnd.n18 gnd.t300 2.82907
R14114 gnd.n16 gnd.t280 2.82907
R14115 gnd.n16 gnd.t347 2.82907
R14116 gnd.n51 gnd.t338 2.82907
R14117 gnd.n51 gnd.t343 2.82907
R14118 gnd.n49 gnd.t297 2.82907
R14119 gnd.n49 gnd.t268 2.82907
R14120 gnd.n47 gnd.t254 2.82907
R14121 gnd.n47 gnd.t326 2.82907
R14122 gnd.n45 gnd.t314 2.82907
R14123 gnd.n45 gnd.t279 2.82907
R14124 gnd.n43 gnd.t267 2.82907
R14125 gnd.n43 gnd.t303 2.82907
R14126 gnd.n41 gnd.t290 2.82907
R14127 gnd.n41 gnd.t299 2.82907
R14128 gnd.n39 gnd.t243 2.82907
R14129 gnd.n39 gnd.t344 2.82907
R14130 gnd.n37 gnd.t335 2.82907
R14131 gnd.n37 gnd.t274 2.82907
R14132 gnd.n35 gnd.t257 2.82907
R14133 gnd.n35 gnd.t331 2.82907
R14134 gnd.n6384 gnd.n6383 2.71565
R14135 gnd.n6352 gnd.n6351 2.71565
R14136 gnd.n6320 gnd.n6319 2.71565
R14137 gnd.n6289 gnd.n6288 2.71565
R14138 gnd.n6257 gnd.n6256 2.71565
R14139 gnd.n6225 gnd.n6224 2.71565
R14140 gnd.n6193 gnd.n6192 2.71565
R14141 gnd.n6162 gnd.n6161 2.71565
R14142 gnd.n3560 gnd.t139 2.54975
R14143 gnd.n3591 gnd.n3586 2.54975
R14144 gnd.n3651 gnd.n2426 2.54975
R14145 gnd.n3753 gnd.n2385 2.54975
R14146 gnd.t22 gnd.n3752 2.54975
R14147 gnd.n3774 gnd.t1 2.54975
R14148 gnd.t54 gnd.n3826 2.54975
R14149 gnd.n3817 gnd.t51 2.54975
R14150 gnd.n3846 gnd.n2345 2.54975
R14151 gnd.n3918 gnd.n3917 2.54975
R14152 gnd.n3983 gnd.n3982 2.54975
R14153 gnd.n3998 gnd.t136 2.54975
R14154 gnd.n5887 gnd.n5349 2.27742
R14155 gnd.n5883 gnd.n5349 2.27742
R14156 gnd.n5879 gnd.n5349 2.27742
R14157 gnd.n5875 gnd.n5349 2.27742
R14158 gnd.n7418 gnd.n7417 2.27742
R14159 gnd.n7418 gnd.n306 2.27742
R14160 gnd.n7418 gnd.n305 2.27742
R14161 gnd.n7418 gnd.n304 2.27742
R14162 gnd.n7418 gnd.n303 2.27742
R14163 gnd.n4464 gnd.n302 2.27742
R14164 gnd.n1707 gnd.n302 2.27742
R14165 gnd.n4536 gnd.n302 2.27742
R14166 gnd.n4537 gnd.n302 2.27742
R14167 gnd.n7390 gnd.n302 2.27742
R14168 gnd.n4945 gnd.n1225 2.27742
R14169 gnd.n1226 gnd.n1225 2.27742
R14170 gnd.n4932 gnd.n1225 2.27742
R14171 gnd.n1245 gnd.n1225 2.27742
R14172 gnd.n4919 gnd.n1225 2.27742
R14173 gnd.n2852 gnd.n2851 2.27742
R14174 gnd.n2851 gnd.n2850 2.27742
R14175 gnd.n2851 gnd.n2774 2.27742
R14176 gnd.n2851 gnd.n2773 2.27742
R14177 gnd.n2851 gnd.n2772 2.27742
R14178 gnd.t87 gnd.n5767 2.23109
R14179 gnd.n5915 gnd.t3 2.23109
R14180 gnd.n3708 gnd.t33 2.23109
R14181 gnd.t70 gnd.n3862 2.23109
R14182 gnd.n6380 gnd.n6370 1.93989
R14183 gnd.n6348 gnd.n6338 1.93989
R14184 gnd.n6316 gnd.n6306 1.93989
R14185 gnd.n6285 gnd.n6275 1.93989
R14186 gnd.n6253 gnd.n6243 1.93989
R14187 gnd.n6221 gnd.n6211 1.93989
R14188 gnd.n6189 gnd.n6179 1.93989
R14189 gnd.n6158 gnd.n6148 1.93989
R14190 gnd.n3560 gnd.n1526 1.91244
R14191 gnd.n3653 gnd.t350 1.91244
R14192 gnd.n3674 gnd.t2 1.91244
R14193 gnd.n3744 gnd.n3743 1.91244
R14194 gnd.n3852 gnd.n2341 1.91244
R14195 gnd.n2326 gnd.t24 1.91244
R14196 gnd.t41 gnd.n2273 1.91244
R14197 gnd.n3995 gnd.n3994 1.91244
R14198 gnd.n5780 gnd.t81 1.59378
R14199 gnd.n5989 gnd.t18 1.59378
R14200 gnd.n6063 gnd.t79 1.59378
R14201 gnd.t229 gnd.n1139 1.59378
R14202 gnd.t48 gnd.n2430 1.59378
R14203 gnd.n3906 gnd.t62 1.59378
R14204 gnd.n7478 gnd.t192 1.59378
R14205 gnd.n3610 gnd.t168 1.27512
R14206 gnd.n3639 gnd.n3638 1.27512
R14207 gnd.t350 gnd.n3652 1.27512
R14208 gnd.n3775 gnd.n3774 1.27512
R14209 gnd.n3826 gnd.n3824 1.27512
R14210 gnd.n3916 gnd.t41 1.27512
R14211 gnd.n2305 gnd.n2304 1.27512
R14212 gnd.n3934 gnd.n3933 1.27512
R14213 gnd.n5577 gnd.n5576 1.16414
R14214 gnd.n6436 gnd.n5164 1.16414
R14215 gnd.n6379 gnd.n6372 1.16414
R14216 gnd.n6347 gnd.n6340 1.16414
R14217 gnd.n6315 gnd.n6308 1.16414
R14218 gnd.n6284 gnd.n6277 1.16414
R14219 gnd.n6252 gnd.n6245 1.16414
R14220 gnd.n6220 gnd.n6213 1.16414
R14221 gnd.n6188 gnd.n6181 1.16414
R14222 gnd.n6157 gnd.n6150 1.16414
R14223 gnd.n2218 gnd.n2217 0.970197
R14224 gnd.n4800 gnd.n1457 0.970197
R14225 gnd.n6363 gnd.n6331 0.962709
R14226 gnd.n6395 gnd.n6363 0.962709
R14227 gnd.n6236 gnd.n6204 0.962709
R14228 gnd.n6268 gnd.n6236 0.962709
R14229 gnd.t35 gnd.n5891 0.956468
R14230 gnd.n5239 gnd.t12 0.956468
R14231 gnd.n3033 gnd.t281 0.956468
R14232 gnd.n2702 gnd.t217 0.956468
R14233 gnd.n3448 gnd.t77 0.956468
R14234 gnd.t33 gnd.t39 0.956468
R14235 gnd.t42 gnd.t70 0.956468
R14236 gnd.n4196 gnd.t46 0.956468
R14237 gnd.n4389 gnd.t306 0.956468
R14238 gnd.n7446 gnd.t240 0.956468
R14239 gnd.n5339 gnd.n5337 0.773756
R14240 gnd.n66 gnd.n64 0.773756
R14241 gnd.n5346 gnd.n5345 0.773756
R14242 gnd.n5345 gnd.n5343 0.773756
R14243 gnd.n5343 gnd.n5341 0.773756
R14244 gnd.n5341 gnd.n5339 0.773756
R14245 gnd.n5337 gnd.n5335 0.773756
R14246 gnd.n5335 gnd.n5333 0.773756
R14247 gnd.n5333 gnd.n5331 0.773756
R14248 gnd.n5331 gnd.n5329 0.773756
R14249 gnd.n58 gnd.n56 0.773756
R14250 gnd.n60 gnd.n58 0.773756
R14251 gnd.n62 gnd.n60 0.773756
R14252 gnd.n64 gnd.n62 0.773756
R14253 gnd.n68 gnd.n66 0.773756
R14254 gnd.n70 gnd.n68 0.773756
R14255 gnd.n72 gnd.n70 0.773756
R14256 gnd.n73 gnd.n72 0.773756
R14257 gnd.n2 gnd.n1 0.672012
R14258 gnd.n3 gnd.n2 0.672012
R14259 gnd.n4 gnd.n3 0.672012
R14260 gnd.n5 gnd.n4 0.672012
R14261 gnd.n6 gnd.n5 0.672012
R14262 gnd.n7 gnd.n6 0.672012
R14263 gnd.n9 gnd.n8 0.672012
R14264 gnd.n10 gnd.n9 0.672012
R14265 gnd.n11 gnd.n10 0.672012
R14266 gnd.n12 gnd.n11 0.672012
R14267 gnd.n13 gnd.n12 0.672012
R14268 gnd.n14 gnd.n13 0.672012
R14269 gnd.n4966 gnd.n1187 0.637812
R14270 gnd.n3041 gnd.n1190 0.637812
R14271 gnd.n4960 gnd.n1198 0.637812
R14272 gnd.n3049 gnd.n1201 0.637812
R14273 gnd.n4954 gnd.n1209 0.637812
R14274 gnd.n3057 gnd.n2857 0.637812
R14275 gnd.n4948 gnd.n1219 0.637812
R14276 gnd.n3065 gnd.n1222 0.637812
R14277 gnd.n4941 gnd.n1228 0.637812
R14278 gnd.n3073 gnd.n1231 0.637812
R14279 gnd.n4935 gnd.n1239 0.637812
R14280 gnd.n3081 gnd.n1242 0.637812
R14281 gnd.n4928 gnd.n1247 0.637812
R14282 gnd.n3089 gnd.n2733 0.637812
R14283 gnd.n4922 gnd.n1256 0.637812
R14284 gnd.n4915 gnd.n1264 0.637812
R14285 gnd.n3105 gnd.n1267 0.637812
R14286 gnd.n4909 gnd.n1275 0.637812
R14287 gnd.n3113 gnd.n1278 0.637812
R14288 gnd.n4903 gnd.n1286 0.637812
R14289 gnd.n3121 gnd.n2720 0.637812
R14290 gnd.n4897 gnd.n1296 0.637812
R14291 gnd.n3129 gnd.n2716 0.637812
R14292 gnd.n4891 gnd.n1306 0.637812
R14293 gnd.n3137 gnd.n1309 0.637812
R14294 gnd.n4885 gnd.n1317 0.637812
R14295 gnd.n3145 gnd.n1320 0.637812
R14296 gnd.n4879 gnd.n1328 0.637812
R14297 gnd.n3153 gnd.n2706 0.637812
R14298 gnd.n4873 gnd.n1338 0.637812
R14299 gnd.n3161 gnd.n2702 0.637812
R14300 gnd.n4867 gnd.n1348 0.637812
R14301 gnd.n3170 gnd.n1351 0.637812
R14302 gnd.n4861 gnd.n1359 0.637812
R14303 gnd.n3178 gnd.n1362 0.637812
R14304 gnd.n4855 gnd.n1370 0.637812
R14305 gnd.n3197 gnd.n3196 0.637812
R14306 gnd.n4849 gnd.n1380 0.637812
R14307 gnd.n3188 gnd.n1383 0.637812
R14308 gnd.n4843 gnd.n1391 0.637812
R14309 gnd.n3258 gnd.n1394 0.637812
R14310 gnd.n4837 gnd.n1402 0.637812
R14311 gnd.n3329 gnd.n1405 0.637812
R14312 gnd.n3550 gnd.t185 0.637812
R14313 gnd.n3691 gnd.t21 0.637812
R14314 gnd.n3688 gnd.n2410 0.637812
R14315 gnd.n3709 gnd.n2402 0.637812
R14316 gnd.n3872 gnd.n2324 0.637812
R14317 gnd.n3880 gnd.n2318 0.637812
R14318 gnd.n3899 gnd.t0 0.637812
R14319 gnd.n3966 gnd.t165 0.637812
R14320 gnd.n4610 gnd.n1633 0.637812
R14321 gnd.n4609 gnd.n1636 0.637812
R14322 gnd.n4284 gnd.n1646 0.637812
R14323 gnd.n4603 gnd.n1649 0.637812
R14324 gnd.n4337 gnd.n4336 0.637812
R14325 gnd.n4348 gnd.n1825 0.637812
R14326 gnd.n4347 gnd.n4346 0.637812
R14327 gnd.n4359 gnd.n4358 0.637812
R14328 gnd.n1807 gnd.n1795 0.637812
R14329 gnd.n4369 gnd.n1797 0.637812
R14330 gnd.n4379 gnd.n1787 0.637812
R14331 gnd.n4378 gnd.n1778 0.637812
R14332 gnd.n4391 gnd.n4389 0.637812
R14333 gnd.n4321 gnd.n1769 0.637812
R14334 gnd.n4401 gnd.n1771 0.637812
R14335 gnd.n4412 gnd.n1761 0.637812
R14336 gnd.n4411 gnd.n1752 0.637812
R14337 gnd.n4423 gnd.n4422 0.637812
R14338 gnd.n4313 gnd.n1743 0.637812
R14339 gnd.n4433 gnd.n1745 0.637812
R14340 gnd.n4449 gnd.n1735 0.637812
R14341 gnd.n4448 gnd.n1725 0.637812
R14342 gnd.n4477 gnd.n4476 0.637812
R14343 gnd.n4439 gnd.n1716 0.637812
R14344 gnd.n4487 gnd.n1718 0.637812
R14345 gnd.n4469 gnd.n4468 0.637812
R14346 gnd.n4559 gnd.n1683 0.637812
R14347 gnd.n4562 gnd.n1686 0.637812
R14348 gnd.n7413 gnd.n313 0.637812
R14349 gnd.n4532 gnd.n4531 0.637812
R14350 gnd.n4547 gnd.n1699 0.637812
R14351 gnd.n4542 gnd.n4541 0.637812
R14352 gnd.n4521 gnd.n1704 0.637812
R14353 gnd.n4523 gnd.n332 0.637812
R14354 gnd.n7394 gnd.n7393 0.637812
R14355 gnd.n7398 gnd.n328 0.637812
R14356 gnd.n4515 gnd.n296 0.637812
R14357 gnd.n7422 gnd.n298 0.637812
R14358 gnd.n4511 gnd.n287 0.637812
R14359 gnd.n7430 gnd.n290 0.637812
R14360 gnd.n7380 gnd.n7379 0.637812
R14361 gnd.n7438 gnd.n281 0.637812
R14362 gnd.n7373 gnd.n7372 0.637812
R14363 gnd.n7721 gnd.n7720 0.63688
R14364 gnd gnd.n0 0.634843
R14365 gnd.n5307 gnd.n5306 0.573776
R14366 gnd.n5306 gnd.n5304 0.573776
R14367 gnd.n5304 gnd.n5302 0.573776
R14368 gnd.n5302 gnd.n5300 0.573776
R14369 gnd.n5300 gnd.n5298 0.573776
R14370 gnd.n5298 gnd.n5296 0.573776
R14371 gnd.n5296 gnd.n5294 0.573776
R14372 gnd.n5294 gnd.n5292 0.573776
R14373 gnd.n5292 gnd.n5290 0.573776
R14374 gnd.n5326 gnd.n5325 0.573776
R14375 gnd.n5325 gnd.n5323 0.573776
R14376 gnd.n5323 gnd.n5321 0.573776
R14377 gnd.n5321 gnd.n5319 0.573776
R14378 gnd.n5319 gnd.n5317 0.573776
R14379 gnd.n5317 gnd.n5315 0.573776
R14380 gnd.n5315 gnd.n5313 0.573776
R14381 gnd.n5313 gnd.n5311 0.573776
R14382 gnd.n5311 gnd.n5309 0.573776
R14383 gnd.n19 gnd.n17 0.573776
R14384 gnd.n21 gnd.n19 0.573776
R14385 gnd.n23 gnd.n21 0.573776
R14386 gnd.n25 gnd.n23 0.573776
R14387 gnd.n27 gnd.n25 0.573776
R14388 gnd.n29 gnd.n27 0.573776
R14389 gnd.n31 gnd.n29 0.573776
R14390 gnd.n33 gnd.n31 0.573776
R14391 gnd.n34 gnd.n33 0.573776
R14392 gnd.n38 gnd.n36 0.573776
R14393 gnd.n40 gnd.n38 0.573776
R14394 gnd.n42 gnd.n40 0.573776
R14395 gnd.n44 gnd.n42 0.573776
R14396 gnd.n46 gnd.n44 0.573776
R14397 gnd.n48 gnd.n46 0.573776
R14398 gnd.n50 gnd.n48 0.573776
R14399 gnd.n52 gnd.n50 0.573776
R14400 gnd.n53 gnd.n52 0.573776
R14401 gnd.n7418 gnd.n302 0.548625
R14402 gnd.n2851 gnd.n1225 0.548625
R14403 gnd.n3378 gnd.n3377 0.523366
R14404 gnd.n1887 gnd.n1610 0.523366
R14405 gnd.n4256 gnd.n4255 0.489829
R14406 gnd.n3235 gnd.n2559 0.489829
R14407 gnd.n6424 gnd.n5168 0.486781
R14408 gnd.n5629 gnd.n5525 0.48678
R14409 gnd.n5119 gnd.n994 0.480683
R14410 gnd.n5697 gnd.n5475 0.480683
R14411 gnd.n2940 gnd.n2938 0.477634
R14412 gnd.n2978 gnd.n2977 0.477634
R14413 gnd.n7569 gnd.n7568 0.477634
R14414 gnd.n7671 gnd.n7670 0.477634
R14415 gnd.n7663 gnd.n7662 0.465439
R14416 gnd.n7592 gnd.n7591 0.465439
R14417 gnd.n2176 gnd.n2170 0.465439
R14418 gnd.n2096 gnd.n2095 0.465439
R14419 gnd.n4833 gnd.n4832 0.465439
R14420 gnd.n3326 gnd.n3325 0.465439
R14421 gnd.n5031 gnd.n1087 0.465439
R14422 gnd.n2987 gnd.n1044 0.465439
R14423 gnd.n798 gnd.n793 0.425805
R14424 gnd.n7157 gnd.n7156 0.425805
R14425 gnd.n7369 gnd.n7368 0.425805
R14426 gnd.n2758 gnd.n2757 0.425805
R14427 gnd.n3242 gnd.n2644 0.388379
R14428 gnd.n6376 gnd.n6375 0.388379
R14429 gnd.n6344 gnd.n6343 0.388379
R14430 gnd.n6312 gnd.n6311 0.388379
R14431 gnd.n6281 gnd.n6280 0.388379
R14432 gnd.n6249 gnd.n6248 0.388379
R14433 gnd.n6217 gnd.n6216 0.388379
R14434 gnd.n6185 gnd.n6184 0.388379
R14435 gnd.n6154 gnd.n6153 0.388379
R14436 gnd.n7632 gnd.n7631 0.388379
R14437 gnd.n5072 gnd.n5071 0.388379
R14438 gnd.n1985 gnd.n1981 0.388379
R14439 gnd.n3376 gnd.n2569 0.377553
R14440 gnd.n1886 gnd.n1885 0.377553
R14441 gnd.n7721 gnd.n15 0.374463
R14442 gnd.n5195 gnd.t5 0.319156
R14443 gnd.n3065 gnd.t248 0.319156
R14444 gnd.t202 gnd.n1259 0.319156
R14445 gnd.n3097 gnd.t202 0.319156
R14446 gnd.n2716 gnd.t204 0.319156
R14447 gnd.n2563 gnd.t161 0.319156
R14448 gnd.n4796 gnd.n1497 0.319156
R14449 gnd.n2431 gnd.t48 0.319156
R14450 gnd.t62 gnd.n3905 0.319156
R14451 gnd.n4163 gnd.n4162 0.319156
R14452 gnd.n4250 gnd.t132 0.319156
R14453 gnd.n4449 gnd.t242 0.319156
R14454 gnd.n4495 gnd.t298 0.319156
R14455 gnd.t298 gnd.n310 0.319156
R14456 gnd.n7398 gnd.t313 0.319156
R14457 gnd.n5623 gnd.n5622 0.311721
R14458 gnd gnd.n7721 0.295112
R14459 gnd.n6481 gnd.n6480 0.268793
R14460 gnd.n3253 gnd.n3252 0.247451
R14461 gnd.n4279 gnd.n1837 0.247451
R14462 gnd.n6480 gnd.n6479 0.241354
R14463 gnd.n2136 gnd.n2135 0.229039
R14464 gnd.n2139 gnd.n2136 0.229039
R14465 gnd.n1461 gnd.n1456 0.229039
R14466 gnd.n3278 gnd.n1461 0.229039
R14467 gnd.n5348 gnd.n0 0.210825
R14468 gnd.n5752 gnd.n5493 0.206293
R14469 gnd.n6393 gnd.n6365 0.155672
R14470 gnd.n6386 gnd.n6365 0.155672
R14471 gnd.n6386 gnd.n6385 0.155672
R14472 gnd.n6385 gnd.n6369 0.155672
R14473 gnd.n6378 gnd.n6369 0.155672
R14474 gnd.n6378 gnd.n6377 0.155672
R14475 gnd.n6361 gnd.n6333 0.155672
R14476 gnd.n6354 gnd.n6333 0.155672
R14477 gnd.n6354 gnd.n6353 0.155672
R14478 gnd.n6353 gnd.n6337 0.155672
R14479 gnd.n6346 gnd.n6337 0.155672
R14480 gnd.n6346 gnd.n6345 0.155672
R14481 gnd.n6329 gnd.n6301 0.155672
R14482 gnd.n6322 gnd.n6301 0.155672
R14483 gnd.n6322 gnd.n6321 0.155672
R14484 gnd.n6321 gnd.n6305 0.155672
R14485 gnd.n6314 gnd.n6305 0.155672
R14486 gnd.n6314 gnd.n6313 0.155672
R14487 gnd.n6298 gnd.n6270 0.155672
R14488 gnd.n6291 gnd.n6270 0.155672
R14489 gnd.n6291 gnd.n6290 0.155672
R14490 gnd.n6290 gnd.n6274 0.155672
R14491 gnd.n6283 gnd.n6274 0.155672
R14492 gnd.n6283 gnd.n6282 0.155672
R14493 gnd.n6266 gnd.n6238 0.155672
R14494 gnd.n6259 gnd.n6238 0.155672
R14495 gnd.n6259 gnd.n6258 0.155672
R14496 gnd.n6258 gnd.n6242 0.155672
R14497 gnd.n6251 gnd.n6242 0.155672
R14498 gnd.n6251 gnd.n6250 0.155672
R14499 gnd.n6234 gnd.n6206 0.155672
R14500 gnd.n6227 gnd.n6206 0.155672
R14501 gnd.n6227 gnd.n6226 0.155672
R14502 gnd.n6226 gnd.n6210 0.155672
R14503 gnd.n6219 gnd.n6210 0.155672
R14504 gnd.n6219 gnd.n6218 0.155672
R14505 gnd.n6202 gnd.n6174 0.155672
R14506 gnd.n6195 gnd.n6174 0.155672
R14507 gnd.n6195 gnd.n6194 0.155672
R14508 gnd.n6194 gnd.n6178 0.155672
R14509 gnd.n6187 gnd.n6178 0.155672
R14510 gnd.n6187 gnd.n6186 0.155672
R14511 gnd.n6171 gnd.n6143 0.155672
R14512 gnd.n6164 gnd.n6143 0.155672
R14513 gnd.n6164 gnd.n6163 0.155672
R14514 gnd.n6163 gnd.n6147 0.155672
R14515 gnd.n6156 gnd.n6147 0.155672
R14516 gnd.n6156 gnd.n6155 0.155672
R14517 gnd.n5120 gnd.n5119 0.152939
R14518 gnd.n5121 gnd.n5120 0.152939
R14519 gnd.n5122 gnd.n5121 0.152939
R14520 gnd.n5123 gnd.n5122 0.152939
R14521 gnd.n5124 gnd.n5123 0.152939
R14522 gnd.n5125 gnd.n5124 0.152939
R14523 gnd.n5126 gnd.n5125 0.152939
R14524 gnd.n5127 gnd.n5126 0.152939
R14525 gnd.n5128 gnd.n5127 0.152939
R14526 gnd.n5129 gnd.n5128 0.152939
R14527 gnd.n5130 gnd.n5129 0.152939
R14528 gnd.n5131 gnd.n5130 0.152939
R14529 gnd.n5132 gnd.n5131 0.152939
R14530 gnd.n5133 gnd.n5132 0.152939
R14531 gnd.n6482 gnd.n5133 0.152939
R14532 gnd.n6482 gnd.n6481 0.152939
R14533 gnd.n5771 gnd.n5475 0.152939
R14534 gnd.n5772 gnd.n5771 0.152939
R14535 gnd.n5773 gnd.n5772 0.152939
R14536 gnd.n5773 gnd.n5454 0.152939
R14537 gnd.n5801 gnd.n5454 0.152939
R14538 gnd.n5802 gnd.n5801 0.152939
R14539 gnd.n5803 gnd.n5802 0.152939
R14540 gnd.n5804 gnd.n5803 0.152939
R14541 gnd.n5804 gnd.n5428 0.152939
R14542 gnd.n5835 gnd.n5428 0.152939
R14543 gnd.n5836 gnd.n5835 0.152939
R14544 gnd.n5837 gnd.n5836 0.152939
R14545 gnd.n5838 gnd.n5837 0.152939
R14546 gnd.n5839 gnd.n5838 0.152939
R14547 gnd.n5839 gnd.n5395 0.152939
R14548 gnd.n5896 gnd.n5395 0.152939
R14549 gnd.n5897 gnd.n5896 0.152939
R14550 gnd.n5898 gnd.n5897 0.152939
R14551 gnd.n5899 gnd.n5898 0.152939
R14552 gnd.n5899 gnd.n5368 0.152939
R14553 gnd.n5936 gnd.n5368 0.152939
R14554 gnd.n5937 gnd.n5936 0.152939
R14555 gnd.n5938 gnd.n5937 0.152939
R14556 gnd.n5939 gnd.n5938 0.152939
R14557 gnd.n5939 gnd.n5281 0.152939
R14558 gnd.n5981 gnd.n5281 0.152939
R14559 gnd.n5982 gnd.n5981 0.152939
R14560 gnd.n5983 gnd.n5982 0.152939
R14561 gnd.n5984 gnd.n5983 0.152939
R14562 gnd.n5984 gnd.n5253 0.152939
R14563 gnd.n6021 gnd.n5253 0.152939
R14564 gnd.n6022 gnd.n6021 0.152939
R14565 gnd.n6023 gnd.n6022 0.152939
R14566 gnd.n6024 gnd.n6023 0.152939
R14567 gnd.n6024 gnd.n5226 0.152939
R14568 gnd.n6067 gnd.n5226 0.152939
R14569 gnd.n6068 gnd.n6067 0.152939
R14570 gnd.n6069 gnd.n6068 0.152939
R14571 gnd.n6070 gnd.n6069 0.152939
R14572 gnd.n6070 gnd.n5199 0.152939
R14573 gnd.n6106 gnd.n5199 0.152939
R14574 gnd.n6107 gnd.n6106 0.152939
R14575 gnd.n6108 gnd.n6107 0.152939
R14576 gnd.n6110 gnd.n6108 0.152939
R14577 gnd.n6110 gnd.n6109 0.152939
R14578 gnd.n6109 gnd.n968 0.152939
R14579 gnd.n969 gnd.n968 0.152939
R14580 gnd.n970 gnd.n969 0.152939
R14581 gnd.n990 gnd.n970 0.152939
R14582 gnd.n991 gnd.n990 0.152939
R14583 gnd.n992 gnd.n991 0.152939
R14584 gnd.n993 gnd.n992 0.152939
R14585 gnd.n994 gnd.n993 0.152939
R14586 gnd.n5698 gnd.n5697 0.152939
R14587 gnd.n5699 gnd.n5698 0.152939
R14588 gnd.n5700 gnd.n5699 0.152939
R14589 gnd.n5701 gnd.n5700 0.152939
R14590 gnd.n5702 gnd.n5701 0.152939
R14591 gnd.n5703 gnd.n5702 0.152939
R14592 gnd.n5704 gnd.n5703 0.152939
R14593 gnd.n5705 gnd.n5704 0.152939
R14594 gnd.n5706 gnd.n5705 0.152939
R14595 gnd.n5707 gnd.n5706 0.152939
R14596 gnd.n5708 gnd.n5707 0.152939
R14597 gnd.n5709 gnd.n5708 0.152939
R14598 gnd.n5710 gnd.n5709 0.152939
R14599 gnd.n5711 gnd.n5710 0.152939
R14600 gnd.n5715 gnd.n5711 0.152939
R14601 gnd.n5715 gnd.n5493 0.152939
R14602 gnd.n6479 gnd.n5139 0.152939
R14603 gnd.n5141 gnd.n5139 0.152939
R14604 gnd.n5142 gnd.n5141 0.152939
R14605 gnd.n5143 gnd.n5142 0.152939
R14606 gnd.n5144 gnd.n5143 0.152939
R14607 gnd.n5145 gnd.n5144 0.152939
R14608 gnd.n5146 gnd.n5145 0.152939
R14609 gnd.n5147 gnd.n5146 0.152939
R14610 gnd.n5148 gnd.n5147 0.152939
R14611 gnd.n5149 gnd.n5148 0.152939
R14612 gnd.n5150 gnd.n5149 0.152939
R14613 gnd.n5151 gnd.n5150 0.152939
R14614 gnd.n5152 gnd.n5151 0.152939
R14615 gnd.n5153 gnd.n5152 0.152939
R14616 gnd.n5154 gnd.n5153 0.152939
R14617 gnd.n5155 gnd.n5154 0.152939
R14618 gnd.n5156 gnd.n5155 0.152939
R14619 gnd.n5157 gnd.n5156 0.152939
R14620 gnd.n5158 gnd.n5157 0.152939
R14621 gnd.n5159 gnd.n5158 0.152939
R14622 gnd.n5160 gnd.n5159 0.152939
R14623 gnd.n5161 gnd.n5160 0.152939
R14624 gnd.n5165 gnd.n5161 0.152939
R14625 gnd.n5166 gnd.n5165 0.152939
R14626 gnd.n5167 gnd.n5166 0.152939
R14627 gnd.n5168 gnd.n5167 0.152939
R14628 gnd.n5958 gnd.n5957 0.152939
R14629 gnd.n5959 gnd.n5958 0.152939
R14630 gnd.n5960 gnd.n5959 0.152939
R14631 gnd.n5961 gnd.n5960 0.152939
R14632 gnd.n5962 gnd.n5961 0.152939
R14633 gnd.n5963 gnd.n5962 0.152939
R14634 gnd.n5964 gnd.n5963 0.152939
R14635 gnd.n5965 gnd.n5964 0.152939
R14636 gnd.n5965 gnd.n5233 0.152939
R14637 gnd.n6042 gnd.n5233 0.152939
R14638 gnd.n6043 gnd.n6042 0.152939
R14639 gnd.n6044 gnd.n6043 0.152939
R14640 gnd.n6045 gnd.n6044 0.152939
R14641 gnd.n6046 gnd.n6045 0.152939
R14642 gnd.n6047 gnd.n6046 0.152939
R14643 gnd.n6048 gnd.n6047 0.152939
R14644 gnd.n6049 gnd.n6048 0.152939
R14645 gnd.n6050 gnd.n6049 0.152939
R14646 gnd.n6050 gnd.n5181 0.152939
R14647 gnd.n6126 gnd.n5181 0.152939
R14648 gnd.n6127 gnd.n6126 0.152939
R14649 gnd.n6128 gnd.n6127 0.152939
R14650 gnd.n6130 gnd.n6128 0.152939
R14651 gnd.n6130 gnd.n6129 0.152939
R14652 gnd.n6129 gnd.n5171 0.152939
R14653 gnd.n6422 gnd.n5171 0.152939
R14654 gnd.n6423 gnd.n6422 0.152939
R14655 gnd.n6424 gnd.n6423 0.152939
R14656 gnd.n5630 gnd.n5629 0.152939
R14657 gnd.n5631 gnd.n5630 0.152939
R14658 gnd.n5631 gnd.n5513 0.152939
R14659 gnd.n5645 gnd.n5513 0.152939
R14660 gnd.n5646 gnd.n5645 0.152939
R14661 gnd.n5647 gnd.n5646 0.152939
R14662 gnd.n5647 gnd.n5500 0.152939
R14663 gnd.n5661 gnd.n5500 0.152939
R14664 gnd.n5662 gnd.n5661 0.152939
R14665 gnd.n5663 gnd.n5662 0.152939
R14666 gnd.n5664 gnd.n5663 0.152939
R14667 gnd.n5665 gnd.n5664 0.152939
R14668 gnd.n5666 gnd.n5665 0.152939
R14669 gnd.n5667 gnd.n5666 0.152939
R14670 gnd.n5668 gnd.n5667 0.152939
R14671 gnd.n5669 gnd.n5668 0.152939
R14672 gnd.n5670 gnd.n5669 0.152939
R14673 gnd.n5671 gnd.n5670 0.152939
R14674 gnd.n5672 gnd.n5671 0.152939
R14675 gnd.n5672 gnd.n5435 0.152939
R14676 gnd.n5824 gnd.n5435 0.152939
R14677 gnd.n5825 gnd.n5824 0.152939
R14678 gnd.n5826 gnd.n5825 0.152939
R14679 gnd.n5827 gnd.n5826 0.152939
R14680 gnd.n5827 gnd.n5402 0.152939
R14681 gnd.n5871 gnd.n5402 0.152939
R14682 gnd.n5872 gnd.n5871 0.152939
R14683 gnd.n5873 gnd.n5872 0.152939
R14684 gnd.n5622 gnd.n5529 0.152939
R14685 gnd.n5532 gnd.n5529 0.152939
R14686 gnd.n5533 gnd.n5532 0.152939
R14687 gnd.n5534 gnd.n5533 0.152939
R14688 gnd.n5537 gnd.n5534 0.152939
R14689 gnd.n5538 gnd.n5537 0.152939
R14690 gnd.n5539 gnd.n5538 0.152939
R14691 gnd.n5540 gnd.n5539 0.152939
R14692 gnd.n5543 gnd.n5540 0.152939
R14693 gnd.n5544 gnd.n5543 0.152939
R14694 gnd.n5545 gnd.n5544 0.152939
R14695 gnd.n5546 gnd.n5545 0.152939
R14696 gnd.n5549 gnd.n5546 0.152939
R14697 gnd.n5550 gnd.n5549 0.152939
R14698 gnd.n5551 gnd.n5550 0.152939
R14699 gnd.n5552 gnd.n5551 0.152939
R14700 gnd.n5555 gnd.n5552 0.152939
R14701 gnd.n5556 gnd.n5555 0.152939
R14702 gnd.n5557 gnd.n5556 0.152939
R14703 gnd.n5558 gnd.n5557 0.152939
R14704 gnd.n5561 gnd.n5558 0.152939
R14705 gnd.n5562 gnd.n5561 0.152939
R14706 gnd.n5565 gnd.n5562 0.152939
R14707 gnd.n5566 gnd.n5565 0.152939
R14708 gnd.n5568 gnd.n5566 0.152939
R14709 gnd.n5568 gnd.n5525 0.152939
R14710 gnd.n6706 gnd.n793 0.152939
R14711 gnd.n6707 gnd.n6706 0.152939
R14712 gnd.n6708 gnd.n6707 0.152939
R14713 gnd.n6708 gnd.n787 0.152939
R14714 gnd.n6716 gnd.n787 0.152939
R14715 gnd.n6717 gnd.n6716 0.152939
R14716 gnd.n6718 gnd.n6717 0.152939
R14717 gnd.n6718 gnd.n781 0.152939
R14718 gnd.n6726 gnd.n781 0.152939
R14719 gnd.n6727 gnd.n6726 0.152939
R14720 gnd.n6728 gnd.n6727 0.152939
R14721 gnd.n6728 gnd.n775 0.152939
R14722 gnd.n6736 gnd.n775 0.152939
R14723 gnd.n6737 gnd.n6736 0.152939
R14724 gnd.n6738 gnd.n6737 0.152939
R14725 gnd.n6738 gnd.n769 0.152939
R14726 gnd.n6746 gnd.n769 0.152939
R14727 gnd.n6747 gnd.n6746 0.152939
R14728 gnd.n6748 gnd.n6747 0.152939
R14729 gnd.n6748 gnd.n763 0.152939
R14730 gnd.n6756 gnd.n763 0.152939
R14731 gnd.n6757 gnd.n6756 0.152939
R14732 gnd.n6758 gnd.n6757 0.152939
R14733 gnd.n6758 gnd.n757 0.152939
R14734 gnd.n6766 gnd.n757 0.152939
R14735 gnd.n6767 gnd.n6766 0.152939
R14736 gnd.n6768 gnd.n6767 0.152939
R14737 gnd.n6768 gnd.n751 0.152939
R14738 gnd.n6776 gnd.n751 0.152939
R14739 gnd.n6777 gnd.n6776 0.152939
R14740 gnd.n6778 gnd.n6777 0.152939
R14741 gnd.n6778 gnd.n745 0.152939
R14742 gnd.n6786 gnd.n745 0.152939
R14743 gnd.n6787 gnd.n6786 0.152939
R14744 gnd.n6788 gnd.n6787 0.152939
R14745 gnd.n6788 gnd.n739 0.152939
R14746 gnd.n6796 gnd.n739 0.152939
R14747 gnd.n6797 gnd.n6796 0.152939
R14748 gnd.n6798 gnd.n6797 0.152939
R14749 gnd.n6798 gnd.n733 0.152939
R14750 gnd.n6806 gnd.n733 0.152939
R14751 gnd.n6807 gnd.n6806 0.152939
R14752 gnd.n6808 gnd.n6807 0.152939
R14753 gnd.n6808 gnd.n727 0.152939
R14754 gnd.n6816 gnd.n727 0.152939
R14755 gnd.n6817 gnd.n6816 0.152939
R14756 gnd.n6818 gnd.n6817 0.152939
R14757 gnd.n6818 gnd.n721 0.152939
R14758 gnd.n6826 gnd.n721 0.152939
R14759 gnd.n6827 gnd.n6826 0.152939
R14760 gnd.n6828 gnd.n6827 0.152939
R14761 gnd.n6828 gnd.n715 0.152939
R14762 gnd.n6836 gnd.n715 0.152939
R14763 gnd.n6837 gnd.n6836 0.152939
R14764 gnd.n6838 gnd.n6837 0.152939
R14765 gnd.n6838 gnd.n709 0.152939
R14766 gnd.n6846 gnd.n709 0.152939
R14767 gnd.n6847 gnd.n6846 0.152939
R14768 gnd.n6848 gnd.n6847 0.152939
R14769 gnd.n6848 gnd.n703 0.152939
R14770 gnd.n6856 gnd.n703 0.152939
R14771 gnd.n6857 gnd.n6856 0.152939
R14772 gnd.n6858 gnd.n6857 0.152939
R14773 gnd.n6858 gnd.n697 0.152939
R14774 gnd.n6866 gnd.n697 0.152939
R14775 gnd.n6867 gnd.n6866 0.152939
R14776 gnd.n6868 gnd.n6867 0.152939
R14777 gnd.n6868 gnd.n691 0.152939
R14778 gnd.n6876 gnd.n691 0.152939
R14779 gnd.n6877 gnd.n6876 0.152939
R14780 gnd.n6878 gnd.n6877 0.152939
R14781 gnd.n6878 gnd.n685 0.152939
R14782 gnd.n6886 gnd.n685 0.152939
R14783 gnd.n6887 gnd.n6886 0.152939
R14784 gnd.n6888 gnd.n6887 0.152939
R14785 gnd.n6888 gnd.n679 0.152939
R14786 gnd.n6896 gnd.n679 0.152939
R14787 gnd.n6897 gnd.n6896 0.152939
R14788 gnd.n6898 gnd.n6897 0.152939
R14789 gnd.n6898 gnd.n673 0.152939
R14790 gnd.n6906 gnd.n673 0.152939
R14791 gnd.n6907 gnd.n6906 0.152939
R14792 gnd.n6908 gnd.n6907 0.152939
R14793 gnd.n6908 gnd.n667 0.152939
R14794 gnd.n6916 gnd.n667 0.152939
R14795 gnd.n6917 gnd.n6916 0.152939
R14796 gnd.n6918 gnd.n6917 0.152939
R14797 gnd.n6918 gnd.n661 0.152939
R14798 gnd.n6926 gnd.n661 0.152939
R14799 gnd.n6927 gnd.n6926 0.152939
R14800 gnd.n6928 gnd.n6927 0.152939
R14801 gnd.n6928 gnd.n655 0.152939
R14802 gnd.n6936 gnd.n655 0.152939
R14803 gnd.n6937 gnd.n6936 0.152939
R14804 gnd.n6938 gnd.n6937 0.152939
R14805 gnd.n6938 gnd.n649 0.152939
R14806 gnd.n6946 gnd.n649 0.152939
R14807 gnd.n6947 gnd.n6946 0.152939
R14808 gnd.n6948 gnd.n6947 0.152939
R14809 gnd.n6948 gnd.n643 0.152939
R14810 gnd.n6956 gnd.n643 0.152939
R14811 gnd.n6957 gnd.n6956 0.152939
R14812 gnd.n6958 gnd.n6957 0.152939
R14813 gnd.n6958 gnd.n637 0.152939
R14814 gnd.n6966 gnd.n637 0.152939
R14815 gnd.n6967 gnd.n6966 0.152939
R14816 gnd.n6968 gnd.n6967 0.152939
R14817 gnd.n6968 gnd.n631 0.152939
R14818 gnd.n6976 gnd.n631 0.152939
R14819 gnd.n6977 gnd.n6976 0.152939
R14820 gnd.n6978 gnd.n6977 0.152939
R14821 gnd.n6978 gnd.n625 0.152939
R14822 gnd.n6986 gnd.n625 0.152939
R14823 gnd.n6987 gnd.n6986 0.152939
R14824 gnd.n6988 gnd.n6987 0.152939
R14825 gnd.n6988 gnd.n619 0.152939
R14826 gnd.n6996 gnd.n619 0.152939
R14827 gnd.n6997 gnd.n6996 0.152939
R14828 gnd.n6998 gnd.n6997 0.152939
R14829 gnd.n6998 gnd.n613 0.152939
R14830 gnd.n7006 gnd.n613 0.152939
R14831 gnd.n7007 gnd.n7006 0.152939
R14832 gnd.n7008 gnd.n7007 0.152939
R14833 gnd.n7008 gnd.n607 0.152939
R14834 gnd.n7016 gnd.n607 0.152939
R14835 gnd.n7017 gnd.n7016 0.152939
R14836 gnd.n7018 gnd.n7017 0.152939
R14837 gnd.n7018 gnd.n601 0.152939
R14838 gnd.n7026 gnd.n601 0.152939
R14839 gnd.n7027 gnd.n7026 0.152939
R14840 gnd.n7028 gnd.n7027 0.152939
R14841 gnd.n7028 gnd.n595 0.152939
R14842 gnd.n7036 gnd.n595 0.152939
R14843 gnd.n7037 gnd.n7036 0.152939
R14844 gnd.n7038 gnd.n7037 0.152939
R14845 gnd.n7038 gnd.n589 0.152939
R14846 gnd.n7046 gnd.n589 0.152939
R14847 gnd.n7047 gnd.n7046 0.152939
R14848 gnd.n7048 gnd.n7047 0.152939
R14849 gnd.n7048 gnd.n583 0.152939
R14850 gnd.n7056 gnd.n583 0.152939
R14851 gnd.n7057 gnd.n7056 0.152939
R14852 gnd.n7058 gnd.n7057 0.152939
R14853 gnd.n7058 gnd.n577 0.152939
R14854 gnd.n7066 gnd.n577 0.152939
R14855 gnd.n7067 gnd.n7066 0.152939
R14856 gnd.n7068 gnd.n7067 0.152939
R14857 gnd.n7068 gnd.n571 0.152939
R14858 gnd.n7076 gnd.n571 0.152939
R14859 gnd.n7077 gnd.n7076 0.152939
R14860 gnd.n7078 gnd.n7077 0.152939
R14861 gnd.n7078 gnd.n565 0.152939
R14862 gnd.n7086 gnd.n565 0.152939
R14863 gnd.n7087 gnd.n7086 0.152939
R14864 gnd.n7088 gnd.n7087 0.152939
R14865 gnd.n7088 gnd.n559 0.152939
R14866 gnd.n7096 gnd.n559 0.152939
R14867 gnd.n7097 gnd.n7096 0.152939
R14868 gnd.n7098 gnd.n7097 0.152939
R14869 gnd.n7098 gnd.n553 0.152939
R14870 gnd.n7106 gnd.n553 0.152939
R14871 gnd.n7107 gnd.n7106 0.152939
R14872 gnd.n7108 gnd.n7107 0.152939
R14873 gnd.n7108 gnd.n547 0.152939
R14874 gnd.n7116 gnd.n547 0.152939
R14875 gnd.n7117 gnd.n7116 0.152939
R14876 gnd.n7118 gnd.n7117 0.152939
R14877 gnd.n7118 gnd.n541 0.152939
R14878 gnd.n7126 gnd.n541 0.152939
R14879 gnd.n7127 gnd.n7126 0.152939
R14880 gnd.n7128 gnd.n7127 0.152939
R14881 gnd.n7128 gnd.n535 0.152939
R14882 gnd.n7136 gnd.n535 0.152939
R14883 gnd.n7137 gnd.n7136 0.152939
R14884 gnd.n7138 gnd.n7137 0.152939
R14885 gnd.n7138 gnd.n529 0.152939
R14886 gnd.n7146 gnd.n529 0.152939
R14887 gnd.n7147 gnd.n7146 0.152939
R14888 gnd.n7148 gnd.n7147 0.152939
R14889 gnd.n7148 gnd.n523 0.152939
R14890 gnd.n7156 gnd.n523 0.152939
R14891 gnd.n7158 gnd.n7157 0.152939
R14892 gnd.n7158 gnd.n517 0.152939
R14893 gnd.n7166 gnd.n517 0.152939
R14894 gnd.n7167 gnd.n7166 0.152939
R14895 gnd.n7168 gnd.n7167 0.152939
R14896 gnd.n7168 gnd.n511 0.152939
R14897 gnd.n7176 gnd.n511 0.152939
R14898 gnd.n7177 gnd.n7176 0.152939
R14899 gnd.n7178 gnd.n7177 0.152939
R14900 gnd.n7178 gnd.n505 0.152939
R14901 gnd.n7186 gnd.n505 0.152939
R14902 gnd.n7187 gnd.n7186 0.152939
R14903 gnd.n7188 gnd.n7187 0.152939
R14904 gnd.n7188 gnd.n499 0.152939
R14905 gnd.n7196 gnd.n499 0.152939
R14906 gnd.n7197 gnd.n7196 0.152939
R14907 gnd.n7198 gnd.n7197 0.152939
R14908 gnd.n7198 gnd.n493 0.152939
R14909 gnd.n7206 gnd.n493 0.152939
R14910 gnd.n7207 gnd.n7206 0.152939
R14911 gnd.n7208 gnd.n7207 0.152939
R14912 gnd.n7208 gnd.n487 0.152939
R14913 gnd.n7216 gnd.n487 0.152939
R14914 gnd.n7217 gnd.n7216 0.152939
R14915 gnd.n7218 gnd.n7217 0.152939
R14916 gnd.n7218 gnd.n481 0.152939
R14917 gnd.n7226 gnd.n481 0.152939
R14918 gnd.n7227 gnd.n7226 0.152939
R14919 gnd.n7228 gnd.n7227 0.152939
R14920 gnd.n7228 gnd.n475 0.152939
R14921 gnd.n7236 gnd.n475 0.152939
R14922 gnd.n7237 gnd.n7236 0.152939
R14923 gnd.n7238 gnd.n7237 0.152939
R14924 gnd.n7238 gnd.n469 0.152939
R14925 gnd.n7246 gnd.n469 0.152939
R14926 gnd.n7247 gnd.n7246 0.152939
R14927 gnd.n7248 gnd.n7247 0.152939
R14928 gnd.n7248 gnd.n463 0.152939
R14929 gnd.n7256 gnd.n463 0.152939
R14930 gnd.n7257 gnd.n7256 0.152939
R14931 gnd.n7258 gnd.n7257 0.152939
R14932 gnd.n7258 gnd.n457 0.152939
R14933 gnd.n7266 gnd.n457 0.152939
R14934 gnd.n7267 gnd.n7266 0.152939
R14935 gnd.n7268 gnd.n7267 0.152939
R14936 gnd.n7268 gnd.n451 0.152939
R14937 gnd.n7276 gnd.n451 0.152939
R14938 gnd.n7277 gnd.n7276 0.152939
R14939 gnd.n7278 gnd.n7277 0.152939
R14940 gnd.n7278 gnd.n445 0.152939
R14941 gnd.n7286 gnd.n445 0.152939
R14942 gnd.n7287 gnd.n7286 0.152939
R14943 gnd.n7288 gnd.n7287 0.152939
R14944 gnd.n7288 gnd.n439 0.152939
R14945 gnd.n7296 gnd.n439 0.152939
R14946 gnd.n7297 gnd.n7296 0.152939
R14947 gnd.n7298 gnd.n7297 0.152939
R14948 gnd.n7298 gnd.n433 0.152939
R14949 gnd.n7306 gnd.n433 0.152939
R14950 gnd.n7307 gnd.n7306 0.152939
R14951 gnd.n7308 gnd.n7307 0.152939
R14952 gnd.n7308 gnd.n427 0.152939
R14953 gnd.n7316 gnd.n427 0.152939
R14954 gnd.n7317 gnd.n7316 0.152939
R14955 gnd.n7318 gnd.n7317 0.152939
R14956 gnd.n7318 gnd.n421 0.152939
R14957 gnd.n7326 gnd.n421 0.152939
R14958 gnd.n7327 gnd.n7326 0.152939
R14959 gnd.n7328 gnd.n7327 0.152939
R14960 gnd.n7328 gnd.n415 0.152939
R14961 gnd.n7336 gnd.n415 0.152939
R14962 gnd.n7337 gnd.n7336 0.152939
R14963 gnd.n7338 gnd.n7337 0.152939
R14964 gnd.n7338 gnd.n409 0.152939
R14965 gnd.n7346 gnd.n409 0.152939
R14966 gnd.n7347 gnd.n7346 0.152939
R14967 gnd.n7348 gnd.n7347 0.152939
R14968 gnd.n7348 gnd.n403 0.152939
R14969 gnd.n7356 gnd.n403 0.152939
R14970 gnd.n7357 gnd.n7356 0.152939
R14971 gnd.n7359 gnd.n7357 0.152939
R14972 gnd.n7359 gnd.n7358 0.152939
R14973 gnd.n7358 gnd.n397 0.152939
R14974 gnd.n7368 gnd.n397 0.152939
R14975 gnd.n340 gnd.n337 0.152939
R14976 gnd.n341 gnd.n340 0.152939
R14977 gnd.n342 gnd.n341 0.152939
R14978 gnd.n343 gnd.n342 0.152939
R14979 gnd.n396 gnd.n343 0.152939
R14980 gnd.n7369 gnd.n396 0.152939
R14981 gnd.n7419 gnd.n7418 0.152939
R14982 gnd.n7419 gnd.n284 0.152939
R14983 gnd.n7433 gnd.n284 0.152939
R14984 gnd.n7434 gnd.n7433 0.152939
R14985 gnd.n7435 gnd.n7434 0.152939
R14986 gnd.n7435 gnd.n269 0.152939
R14987 gnd.n7449 gnd.n269 0.152939
R14988 gnd.n7450 gnd.n7449 0.152939
R14989 gnd.n7451 gnd.n7450 0.152939
R14990 gnd.n7451 gnd.n253 0.152939
R14991 gnd.n7465 gnd.n253 0.152939
R14992 gnd.n7466 gnd.n7465 0.152939
R14993 gnd.n7467 gnd.n7466 0.152939
R14994 gnd.n7467 gnd.n239 0.152939
R14995 gnd.n7481 gnd.n239 0.152939
R14996 gnd.n7482 gnd.n7481 0.152939
R14997 gnd.n7483 gnd.n7482 0.152939
R14998 gnd.n7483 gnd.n223 0.152939
R14999 gnd.n7497 gnd.n223 0.152939
R15000 gnd.n7498 gnd.n7497 0.152939
R15001 gnd.n7499 gnd.n7498 0.152939
R15002 gnd.n7499 gnd.n206 0.152939
R15003 gnd.n7581 gnd.n206 0.152939
R15004 gnd.n7582 gnd.n7581 0.152939
R15005 gnd.n7583 gnd.n7582 0.152939
R15006 gnd.n7583 gnd.n129 0.152939
R15007 gnd.n7663 gnd.n129 0.152939
R15008 gnd.n7662 gnd.n130 0.152939
R15009 gnd.n132 gnd.n130 0.152939
R15010 gnd.n136 gnd.n132 0.152939
R15011 gnd.n137 gnd.n136 0.152939
R15012 gnd.n138 gnd.n137 0.152939
R15013 gnd.n139 gnd.n138 0.152939
R15014 gnd.n143 gnd.n139 0.152939
R15015 gnd.n144 gnd.n143 0.152939
R15016 gnd.n145 gnd.n144 0.152939
R15017 gnd.n146 gnd.n145 0.152939
R15018 gnd.n150 gnd.n146 0.152939
R15019 gnd.n151 gnd.n150 0.152939
R15020 gnd.n152 gnd.n151 0.152939
R15021 gnd.n153 gnd.n152 0.152939
R15022 gnd.n157 gnd.n153 0.152939
R15023 gnd.n158 gnd.n157 0.152939
R15024 gnd.n159 gnd.n158 0.152939
R15025 gnd.n160 gnd.n159 0.152939
R15026 gnd.n164 gnd.n160 0.152939
R15027 gnd.n165 gnd.n164 0.152939
R15028 gnd.n166 gnd.n165 0.152939
R15029 gnd.n167 gnd.n166 0.152939
R15030 gnd.n171 gnd.n167 0.152939
R15031 gnd.n172 gnd.n171 0.152939
R15032 gnd.n173 gnd.n172 0.152939
R15033 gnd.n174 gnd.n173 0.152939
R15034 gnd.n178 gnd.n174 0.152939
R15035 gnd.n179 gnd.n178 0.152939
R15036 gnd.n180 gnd.n179 0.152939
R15037 gnd.n181 gnd.n180 0.152939
R15038 gnd.n185 gnd.n181 0.152939
R15039 gnd.n186 gnd.n185 0.152939
R15040 gnd.n187 gnd.n186 0.152939
R15041 gnd.n188 gnd.n187 0.152939
R15042 gnd.n192 gnd.n188 0.152939
R15043 gnd.n193 gnd.n192 0.152939
R15044 gnd.n7593 gnd.n193 0.152939
R15045 gnd.n7593 gnd.n7592 0.152939
R15046 gnd.n2170 gnd.n1834 0.152939
R15047 gnd.n4287 gnd.n1834 0.152939
R15048 gnd.n4288 gnd.n4287 0.152939
R15049 gnd.n4289 gnd.n4288 0.152939
R15050 gnd.n4290 gnd.n4289 0.152939
R15051 gnd.n4291 gnd.n4290 0.152939
R15052 gnd.n4292 gnd.n4291 0.152939
R15053 gnd.n4293 gnd.n4292 0.152939
R15054 gnd.n4294 gnd.n4293 0.152939
R15055 gnd.n4295 gnd.n4294 0.152939
R15056 gnd.n4296 gnd.n4295 0.152939
R15057 gnd.n4297 gnd.n4296 0.152939
R15058 gnd.n4298 gnd.n4297 0.152939
R15059 gnd.n4299 gnd.n4298 0.152939
R15060 gnd.n4300 gnd.n4299 0.152939
R15061 gnd.n4301 gnd.n4300 0.152939
R15062 gnd.n4302 gnd.n4301 0.152939
R15063 gnd.n4303 gnd.n4302 0.152939
R15064 gnd.n4304 gnd.n4303 0.152939
R15065 gnd.n4305 gnd.n4304 0.152939
R15066 gnd.n4306 gnd.n4305 0.152939
R15067 gnd.n4307 gnd.n4306 0.152939
R15068 gnd.n4307 gnd.n1712 0.152939
R15069 gnd.n4490 gnd.n1712 0.152939
R15070 gnd.n4491 gnd.n4490 0.152939
R15071 gnd.n4492 gnd.n4491 0.152939
R15072 gnd.n4492 gnd.n1710 0.152939
R15073 gnd.n4498 gnd.n1710 0.152939
R15074 gnd.n4499 gnd.n4498 0.152939
R15075 gnd.n4500 gnd.n4499 0.152939
R15076 gnd.n4501 gnd.n4500 0.152939
R15077 gnd.n4502 gnd.n4501 0.152939
R15078 gnd.n4503 gnd.n4502 0.152939
R15079 gnd.n4504 gnd.n4503 0.152939
R15080 gnd.n4505 gnd.n4504 0.152939
R15081 gnd.n4506 gnd.n4505 0.152939
R15082 gnd.n4507 gnd.n4506 0.152939
R15083 gnd.n4508 gnd.n4507 0.152939
R15084 gnd.n4510 gnd.n4508 0.152939
R15085 gnd.n4510 gnd.n4509 0.152939
R15086 gnd.n4509 gnd.n347 0.152939
R15087 gnd.n348 gnd.n347 0.152939
R15088 gnd.n349 gnd.n348 0.152939
R15089 gnd.n350 gnd.n349 0.152939
R15090 gnd.n351 gnd.n350 0.152939
R15091 gnd.n352 gnd.n351 0.152939
R15092 gnd.n353 gnd.n352 0.152939
R15093 gnd.n354 gnd.n353 0.152939
R15094 gnd.n355 gnd.n354 0.152939
R15095 gnd.n356 gnd.n355 0.152939
R15096 gnd.n357 gnd.n356 0.152939
R15097 gnd.n358 gnd.n357 0.152939
R15098 gnd.n359 gnd.n358 0.152939
R15099 gnd.n360 gnd.n359 0.152939
R15100 gnd.n361 gnd.n360 0.152939
R15101 gnd.n362 gnd.n361 0.152939
R15102 gnd.n363 gnd.n362 0.152939
R15103 gnd.n364 gnd.n363 0.152939
R15104 gnd.n365 gnd.n364 0.152939
R15105 gnd.n366 gnd.n365 0.152939
R15106 gnd.n368 gnd.n366 0.152939
R15107 gnd.n368 gnd.n367 0.152939
R15108 gnd.n367 gnd.n199 0.152939
R15109 gnd.n7591 gnd.n199 0.152939
R15110 gnd.n2102 gnd.n2096 0.152939
R15111 gnd.n2103 gnd.n2102 0.152939
R15112 gnd.n2104 gnd.n2103 0.152939
R15113 gnd.n2104 gnd.n2091 0.152939
R15114 gnd.n2112 gnd.n2091 0.152939
R15115 gnd.n2113 gnd.n2112 0.152939
R15116 gnd.n2114 gnd.n2113 0.152939
R15117 gnd.n2114 gnd.n2087 0.152939
R15118 gnd.n2122 gnd.n2087 0.152939
R15119 gnd.n2123 gnd.n2122 0.152939
R15120 gnd.n2125 gnd.n2123 0.152939
R15121 gnd.n2125 gnd.n2124 0.152939
R15122 gnd.n2124 gnd.n2080 0.152939
R15123 gnd.n2134 gnd.n2080 0.152939
R15124 gnd.n2135 gnd.n2134 0.152939
R15125 gnd.n2142 gnd.n2139 0.152939
R15126 gnd.n2143 gnd.n2142 0.152939
R15127 gnd.n2144 gnd.n2143 0.152939
R15128 gnd.n2145 gnd.n2144 0.152939
R15129 gnd.n2148 gnd.n2145 0.152939
R15130 gnd.n2149 gnd.n2148 0.152939
R15131 gnd.n2150 gnd.n2149 0.152939
R15132 gnd.n2151 gnd.n2150 0.152939
R15133 gnd.n2154 gnd.n2151 0.152939
R15134 gnd.n2155 gnd.n2154 0.152939
R15135 gnd.n2156 gnd.n2155 0.152939
R15136 gnd.n2157 gnd.n2156 0.152939
R15137 gnd.n2160 gnd.n2157 0.152939
R15138 gnd.n2161 gnd.n2160 0.152939
R15139 gnd.n2162 gnd.n2161 0.152939
R15140 gnd.n2163 gnd.n2162 0.152939
R15141 gnd.n2169 gnd.n2163 0.152939
R15142 gnd.n2178 gnd.n2169 0.152939
R15143 gnd.n2178 gnd.n2177 0.152939
R15144 gnd.n2177 gnd.n2176 0.152939
R15145 gnd.n2095 gnd.n1641 0.152939
R15146 gnd.n1642 gnd.n1641 0.152939
R15147 gnd.n1643 gnd.n1642 0.152939
R15148 gnd.n1821 gnd.n1643 0.152939
R15149 gnd.n1822 gnd.n1821 0.152939
R15150 gnd.n1822 gnd.n1801 0.152939
R15151 gnd.n4362 gnd.n1801 0.152939
R15152 gnd.n4363 gnd.n4362 0.152939
R15153 gnd.n4364 gnd.n4363 0.152939
R15154 gnd.n4365 gnd.n4364 0.152939
R15155 gnd.n4365 gnd.n1775 0.152939
R15156 gnd.n4394 gnd.n1775 0.152939
R15157 gnd.n4395 gnd.n4394 0.152939
R15158 gnd.n4396 gnd.n4395 0.152939
R15159 gnd.n4397 gnd.n4396 0.152939
R15160 gnd.n4397 gnd.n1749 0.152939
R15161 gnd.n4426 gnd.n1749 0.152939
R15162 gnd.n4427 gnd.n4426 0.152939
R15163 gnd.n4428 gnd.n4427 0.152939
R15164 gnd.n4429 gnd.n4428 0.152939
R15165 gnd.n4429 gnd.n1722 0.152939
R15166 gnd.n4480 gnd.n1722 0.152939
R15167 gnd.n4481 gnd.n4480 0.152939
R15168 gnd.n4482 gnd.n4481 0.152939
R15169 gnd.n4483 gnd.n4482 0.152939
R15170 gnd.n4483 gnd.n301 0.152939
R15171 gnd.n7418 gnd.n301 0.152939
R15172 gnd.n2778 gnd.n2771 0.152939
R15173 gnd.n2781 gnd.n2778 0.152939
R15174 gnd.n2782 gnd.n2781 0.152939
R15175 gnd.n2783 gnd.n2782 0.152939
R15176 gnd.n2784 gnd.n2783 0.152939
R15177 gnd.n2787 gnd.n2784 0.152939
R15178 gnd.n2788 gnd.n2787 0.152939
R15179 gnd.n2789 gnd.n2788 0.152939
R15180 gnd.n2790 gnd.n2789 0.152939
R15181 gnd.n2793 gnd.n2790 0.152939
R15182 gnd.n2794 gnd.n2793 0.152939
R15183 gnd.n2795 gnd.n2794 0.152939
R15184 gnd.n2796 gnd.n2795 0.152939
R15185 gnd.n2799 gnd.n2796 0.152939
R15186 gnd.n2800 gnd.n2799 0.152939
R15187 gnd.n2801 gnd.n2800 0.152939
R15188 gnd.n2802 gnd.n2801 0.152939
R15189 gnd.n2803 gnd.n2802 0.152939
R15190 gnd.n2804 gnd.n2803 0.152939
R15191 gnd.n2804 gnd.n2685 0.152939
R15192 gnd.n3201 gnd.n2685 0.152939
R15193 gnd.n3202 gnd.n3201 0.152939
R15194 gnd.n3203 gnd.n3202 0.152939
R15195 gnd.n3203 gnd.n2681 0.152939
R15196 gnd.n3209 gnd.n2681 0.152939
R15197 gnd.n3210 gnd.n3209 0.152939
R15198 gnd.n3211 gnd.n3210 0.152939
R15199 gnd.n3211 gnd.n2677 0.152939
R15200 gnd.n3218 gnd.n2677 0.152939
R15201 gnd.n3219 gnd.n3218 0.152939
R15202 gnd.n3220 gnd.n3219 0.152939
R15203 gnd.n3221 gnd.n3220 0.152939
R15204 gnd.n3222 gnd.n3221 0.152939
R15205 gnd.n3222 gnd.n2552 0.152939
R15206 gnd.n3396 gnd.n2552 0.152939
R15207 gnd.n3397 gnd.n3396 0.152939
R15208 gnd.n3398 gnd.n3397 0.152939
R15209 gnd.n3399 gnd.n3398 0.152939
R15210 gnd.n3399 gnd.n2527 0.152939
R15211 gnd.n3426 gnd.n2527 0.152939
R15212 gnd.n3427 gnd.n3426 0.152939
R15213 gnd.n3428 gnd.n3427 0.152939
R15214 gnd.n3429 gnd.n3428 0.152939
R15215 gnd.n3430 gnd.n3429 0.152939
R15216 gnd.n3431 gnd.n3430 0.152939
R15217 gnd.n3431 gnd.n2492 0.152939
R15218 gnd.n3473 gnd.n2492 0.152939
R15219 gnd.n3474 gnd.n3473 0.152939
R15220 gnd.n3475 gnd.n3474 0.152939
R15221 gnd.n3476 gnd.n3475 0.152939
R15222 gnd.n3476 gnd.n2477 0.152939
R15223 gnd.n3595 gnd.n2477 0.152939
R15224 gnd.n3596 gnd.n3595 0.152939
R15225 gnd.n3597 gnd.n3596 0.152939
R15226 gnd.n3597 gnd.n2456 0.152939
R15227 gnd.n3622 gnd.n2456 0.152939
R15228 gnd.n3623 gnd.n3622 0.152939
R15229 gnd.n3624 gnd.n3623 0.152939
R15230 gnd.n3625 gnd.n3624 0.152939
R15231 gnd.n3625 gnd.n2423 0.152939
R15232 gnd.n3664 gnd.n2423 0.152939
R15233 gnd.n3665 gnd.n3664 0.152939
R15234 gnd.n3666 gnd.n3665 0.152939
R15235 gnd.n3667 gnd.n3666 0.152939
R15236 gnd.n3668 gnd.n3667 0.152939
R15237 gnd.n3669 gnd.n3668 0.152939
R15238 gnd.n3669 gnd.n2389 0.152939
R15239 gnd.n3747 gnd.n2389 0.152939
R15240 gnd.n3748 gnd.n3747 0.152939
R15241 gnd.n3749 gnd.n3748 0.152939
R15242 gnd.n3749 gnd.n2366 0.152939
R15243 gnd.n3790 gnd.n2366 0.152939
R15244 gnd.n3791 gnd.n3790 0.152939
R15245 gnd.n3792 gnd.n3791 0.152939
R15246 gnd.n3792 gnd.n2350 0.152939
R15247 gnd.n3838 gnd.n2350 0.152939
R15248 gnd.n3839 gnd.n3838 0.152939
R15249 gnd.n3840 gnd.n3839 0.152939
R15250 gnd.n3841 gnd.n3840 0.152939
R15251 gnd.n3841 gnd.n2321 0.152939
R15252 gnd.n3875 gnd.n2321 0.152939
R15253 gnd.n3876 gnd.n3875 0.152939
R15254 gnd.n3877 gnd.n3876 0.152939
R15255 gnd.n3877 gnd.n2284 0.152939
R15256 gnd.n3909 gnd.n2284 0.152939
R15257 gnd.n3910 gnd.n3909 0.152939
R15258 gnd.n3911 gnd.n3910 0.152939
R15259 gnd.n3912 gnd.n3911 0.152939
R15260 gnd.n3912 gnd.n2255 0.152939
R15261 gnd.n3961 gnd.n2255 0.152939
R15262 gnd.n3962 gnd.n3961 0.152939
R15263 gnd.n3963 gnd.n3962 0.152939
R15264 gnd.n3963 gnd.n2236 0.152939
R15265 gnd.n3987 gnd.n2236 0.152939
R15266 gnd.n3988 gnd.n3987 0.152939
R15267 gnd.n3989 gnd.n3988 0.152939
R15268 gnd.n3990 gnd.n3989 0.152939
R15269 gnd.n3990 gnd.n2035 0.152939
R15270 gnd.n4179 gnd.n2035 0.152939
R15271 gnd.n4180 gnd.n4179 0.152939
R15272 gnd.n4181 gnd.n4180 0.152939
R15273 gnd.n4181 gnd.n2023 0.152939
R15274 gnd.n4200 gnd.n2023 0.152939
R15275 gnd.n4201 gnd.n4200 0.152939
R15276 gnd.n4202 gnd.n4201 0.152939
R15277 gnd.n4202 gnd.n2011 0.152939
R15278 gnd.n4221 gnd.n2011 0.152939
R15279 gnd.n4222 gnd.n4221 0.152939
R15280 gnd.n4223 gnd.n4222 0.152939
R15281 gnd.n4223 gnd.n1999 0.152939
R15282 gnd.n4244 gnd.n1999 0.152939
R15283 gnd.n4245 gnd.n4244 0.152939
R15284 gnd.n4247 gnd.n4245 0.152939
R15285 gnd.n4247 gnd.n4246 0.152939
R15286 gnd.n4246 gnd.n1618 0.152939
R15287 gnd.n1619 gnd.n1618 0.152939
R15288 gnd.n1620 gnd.n1619 0.152939
R15289 gnd.n1626 gnd.n1620 0.152939
R15290 gnd.n1627 gnd.n1626 0.152939
R15291 gnd.n1628 gnd.n1627 0.152939
R15292 gnd.n1629 gnd.n1628 0.152939
R15293 gnd.n1815 gnd.n1629 0.152939
R15294 gnd.n1816 gnd.n1815 0.152939
R15295 gnd.n1817 gnd.n1816 0.152939
R15296 gnd.n1817 gnd.n1811 0.152939
R15297 gnd.n4351 gnd.n1811 0.152939
R15298 gnd.n4352 gnd.n4351 0.152939
R15299 gnd.n4353 gnd.n4352 0.152939
R15300 gnd.n4354 gnd.n4353 0.152939
R15301 gnd.n4354 gnd.n1784 0.152939
R15302 gnd.n4382 gnd.n1784 0.152939
R15303 gnd.n4383 gnd.n4382 0.152939
R15304 gnd.n4384 gnd.n4383 0.152939
R15305 gnd.n4385 gnd.n4384 0.152939
R15306 gnd.n4385 gnd.n1758 0.152939
R15307 gnd.n4415 gnd.n1758 0.152939
R15308 gnd.n4416 gnd.n4415 0.152939
R15309 gnd.n4417 gnd.n4416 0.152939
R15310 gnd.n4418 gnd.n4417 0.152939
R15311 gnd.n4418 gnd.n1731 0.152939
R15312 gnd.n4452 gnd.n1731 0.152939
R15313 gnd.n4453 gnd.n4452 0.152939
R15314 gnd.n4454 gnd.n4453 0.152939
R15315 gnd.n4455 gnd.n4454 0.152939
R15316 gnd.n4456 gnd.n4455 0.152939
R15317 gnd.n4459 gnd.n4456 0.152939
R15318 gnd.n4460 gnd.n4459 0.152939
R15319 gnd.n2938 gnd.n2911 0.152939
R15320 gnd.n2996 gnd.n2911 0.152939
R15321 gnd.n2997 gnd.n2996 0.152939
R15322 gnd.n2998 gnd.n2997 0.152939
R15323 gnd.n2998 gnd.n2909 0.152939
R15324 gnd.n3004 gnd.n2909 0.152939
R15325 gnd.n3005 gnd.n3004 0.152939
R15326 gnd.n3006 gnd.n3005 0.152939
R15327 gnd.n3006 gnd.n2907 0.152939
R15328 gnd.n3012 gnd.n2907 0.152939
R15329 gnd.n3013 gnd.n3012 0.152939
R15330 gnd.n3014 gnd.n3013 0.152939
R15331 gnd.n3014 gnd.n2905 0.152939
R15332 gnd.n3020 gnd.n2905 0.152939
R15333 gnd.n3021 gnd.n3020 0.152939
R15334 gnd.n3022 gnd.n3021 0.152939
R15335 gnd.n3022 gnd.n2903 0.152939
R15336 gnd.n3028 gnd.n2903 0.152939
R15337 gnd.n3029 gnd.n3028 0.152939
R15338 gnd.n3030 gnd.n3029 0.152939
R15339 gnd.n3030 gnd.n2862 0.152939
R15340 gnd.n3044 gnd.n2862 0.152939
R15341 gnd.n3045 gnd.n3044 0.152939
R15342 gnd.n3046 gnd.n3045 0.152939
R15343 gnd.n3046 gnd.n2745 0.152939
R15344 gnd.n3060 gnd.n2745 0.152939
R15345 gnd.n3061 gnd.n3060 0.152939
R15346 gnd.n3062 gnd.n3061 0.152939
R15347 gnd.n3062 gnd.n2739 0.152939
R15348 gnd.n3076 gnd.n2739 0.152939
R15349 gnd.n3077 gnd.n3076 0.152939
R15350 gnd.n2977 gnd.n2918 0.152939
R15351 gnd.n2919 gnd.n2918 0.152939
R15352 gnd.n2920 gnd.n2919 0.152939
R15353 gnd.n2921 gnd.n2920 0.152939
R15354 gnd.n2922 gnd.n2921 0.152939
R15355 gnd.n2923 gnd.n2922 0.152939
R15356 gnd.n2924 gnd.n2923 0.152939
R15357 gnd.n2925 gnd.n2924 0.152939
R15358 gnd.n2926 gnd.n2925 0.152939
R15359 gnd.n2927 gnd.n2926 0.152939
R15360 gnd.n2928 gnd.n2927 0.152939
R15361 gnd.n2929 gnd.n2928 0.152939
R15362 gnd.n2930 gnd.n2929 0.152939
R15363 gnd.n2931 gnd.n2930 0.152939
R15364 gnd.n2932 gnd.n2931 0.152939
R15365 gnd.n2942 gnd.n2932 0.152939
R15366 gnd.n2942 gnd.n2941 0.152939
R15367 gnd.n2941 gnd.n2940 0.152939
R15368 gnd.n2983 gnd.n2978 0.152939
R15369 gnd.n2983 gnd.n2982 0.152939
R15370 gnd.n2982 gnd.n2981 0.152939
R15371 gnd.n2981 gnd.n2979 0.152939
R15372 gnd.n2979 gnd.n1112 0.152939
R15373 gnd.n1113 gnd.n1112 0.152939
R15374 gnd.n1114 gnd.n1113 0.152939
R15375 gnd.n1130 gnd.n1114 0.152939
R15376 gnd.n1131 gnd.n1130 0.152939
R15377 gnd.n1132 gnd.n1131 0.152939
R15378 gnd.n1133 gnd.n1132 0.152939
R15379 gnd.n1151 gnd.n1133 0.152939
R15380 gnd.n1152 gnd.n1151 0.152939
R15381 gnd.n1153 gnd.n1152 0.152939
R15382 gnd.n1154 gnd.n1153 0.152939
R15383 gnd.n1170 gnd.n1154 0.152939
R15384 gnd.n1171 gnd.n1170 0.152939
R15385 gnd.n1172 gnd.n1171 0.152939
R15386 gnd.n1173 gnd.n1172 0.152939
R15387 gnd.n1192 gnd.n1173 0.152939
R15388 gnd.n1193 gnd.n1192 0.152939
R15389 gnd.n1194 gnd.n1193 0.152939
R15390 gnd.n1195 gnd.n1194 0.152939
R15391 gnd.n1213 gnd.n1195 0.152939
R15392 gnd.n1214 gnd.n1213 0.152939
R15393 gnd.n1215 gnd.n1214 0.152939
R15394 gnd.n1216 gnd.n1215 0.152939
R15395 gnd.n1233 gnd.n1216 0.152939
R15396 gnd.n1234 gnd.n1233 0.152939
R15397 gnd.n1235 gnd.n1234 0.152939
R15398 gnd.n1236 gnd.n1235 0.152939
R15399 gnd.n2735 gnd.n1236 0.152939
R15400 gnd.n2735 gnd.n1251 0.152939
R15401 gnd.n1252 gnd.n1251 0.152939
R15402 gnd.n1253 gnd.n1252 0.152939
R15403 gnd.n1269 gnd.n1253 0.152939
R15404 gnd.n1270 gnd.n1269 0.152939
R15405 gnd.n1271 gnd.n1270 0.152939
R15406 gnd.n1272 gnd.n1271 0.152939
R15407 gnd.n1290 gnd.n1272 0.152939
R15408 gnd.n1291 gnd.n1290 0.152939
R15409 gnd.n1292 gnd.n1291 0.152939
R15410 gnd.n1293 gnd.n1292 0.152939
R15411 gnd.n1311 gnd.n1293 0.152939
R15412 gnd.n1312 gnd.n1311 0.152939
R15413 gnd.n1313 gnd.n1312 0.152939
R15414 gnd.n1314 gnd.n1313 0.152939
R15415 gnd.n1332 gnd.n1314 0.152939
R15416 gnd.n1333 gnd.n1332 0.152939
R15417 gnd.n1334 gnd.n1333 0.152939
R15418 gnd.n1335 gnd.n1334 0.152939
R15419 gnd.n1353 gnd.n1335 0.152939
R15420 gnd.n1354 gnd.n1353 0.152939
R15421 gnd.n1355 gnd.n1354 0.152939
R15422 gnd.n1356 gnd.n1355 0.152939
R15423 gnd.n1374 gnd.n1356 0.152939
R15424 gnd.n1375 gnd.n1374 0.152939
R15425 gnd.n1376 gnd.n1375 0.152939
R15426 gnd.n1377 gnd.n1376 0.152939
R15427 gnd.n1396 gnd.n1377 0.152939
R15428 gnd.n1397 gnd.n1396 0.152939
R15429 gnd.n1398 gnd.n1397 0.152939
R15430 gnd.n1399 gnd.n1398 0.152939
R15431 gnd.n2569 gnd.n1399 0.152939
R15432 gnd.n1280 gnd.n1225 0.152939
R15433 gnd.n1281 gnd.n1280 0.152939
R15434 gnd.n1282 gnd.n1281 0.152939
R15435 gnd.n1283 gnd.n1282 0.152939
R15436 gnd.n1300 gnd.n1283 0.152939
R15437 gnd.n1301 gnd.n1300 0.152939
R15438 gnd.n1302 gnd.n1301 0.152939
R15439 gnd.n1303 gnd.n1302 0.152939
R15440 gnd.n1322 gnd.n1303 0.152939
R15441 gnd.n1323 gnd.n1322 0.152939
R15442 gnd.n1324 gnd.n1323 0.152939
R15443 gnd.n1325 gnd.n1324 0.152939
R15444 gnd.n1342 gnd.n1325 0.152939
R15445 gnd.n1343 gnd.n1342 0.152939
R15446 gnd.n1344 gnd.n1343 0.152939
R15447 gnd.n1345 gnd.n1344 0.152939
R15448 gnd.n1364 gnd.n1345 0.152939
R15449 gnd.n1365 gnd.n1364 0.152939
R15450 gnd.n1366 gnd.n1365 0.152939
R15451 gnd.n1367 gnd.n1366 0.152939
R15452 gnd.n1385 gnd.n1367 0.152939
R15453 gnd.n1386 gnd.n1385 0.152939
R15454 gnd.n1387 gnd.n1386 0.152939
R15455 gnd.n1388 gnd.n1387 0.152939
R15456 gnd.n1407 gnd.n1388 0.152939
R15457 gnd.n1408 gnd.n1407 0.152939
R15458 gnd.n4833 gnd.n1408 0.152939
R15459 gnd.n4832 gnd.n1409 0.152939
R15460 gnd.n1443 gnd.n1409 0.152939
R15461 gnd.n1444 gnd.n1443 0.152939
R15462 gnd.n1445 gnd.n1444 0.152939
R15463 gnd.n1446 gnd.n1445 0.152939
R15464 gnd.n1447 gnd.n1446 0.152939
R15465 gnd.n1448 gnd.n1447 0.152939
R15466 gnd.n1449 gnd.n1448 0.152939
R15467 gnd.n1450 gnd.n1449 0.152939
R15468 gnd.n1451 gnd.n1450 0.152939
R15469 gnd.n1452 gnd.n1451 0.152939
R15470 gnd.n1453 gnd.n1452 0.152939
R15471 gnd.n1454 gnd.n1453 0.152939
R15472 gnd.n1455 gnd.n1454 0.152939
R15473 gnd.n1456 gnd.n1455 0.152939
R15474 gnd.n3279 gnd.n3278 0.152939
R15475 gnd.n3280 gnd.n3279 0.152939
R15476 gnd.n3280 gnd.n3274 0.152939
R15477 gnd.n3288 gnd.n3274 0.152939
R15478 gnd.n3289 gnd.n3288 0.152939
R15479 gnd.n3290 gnd.n3289 0.152939
R15480 gnd.n3290 gnd.n3272 0.152939
R15481 gnd.n3298 gnd.n3272 0.152939
R15482 gnd.n3299 gnd.n3298 0.152939
R15483 gnd.n3300 gnd.n3299 0.152939
R15484 gnd.n3300 gnd.n3270 0.152939
R15485 gnd.n3308 gnd.n3270 0.152939
R15486 gnd.n3309 gnd.n3308 0.152939
R15487 gnd.n3310 gnd.n3309 0.152939
R15488 gnd.n3310 gnd.n3268 0.152939
R15489 gnd.n3318 gnd.n3268 0.152939
R15490 gnd.n3319 gnd.n3318 0.152939
R15491 gnd.n3320 gnd.n3319 0.152939
R15492 gnd.n3320 gnd.n3263 0.152939
R15493 gnd.n3325 gnd.n3263 0.152939
R15494 gnd.n5025 gnd.n1087 0.152939
R15495 gnd.n5025 gnd.n5024 0.152939
R15496 gnd.n5024 gnd.n5023 0.152939
R15497 gnd.n5023 gnd.n1090 0.152939
R15498 gnd.n2873 gnd.n1090 0.152939
R15499 gnd.n2874 gnd.n2873 0.152939
R15500 gnd.n2874 gnd.n2871 0.152939
R15501 gnd.n2880 gnd.n2871 0.152939
R15502 gnd.n2881 gnd.n2880 0.152939
R15503 gnd.n2882 gnd.n2881 0.152939
R15504 gnd.n2882 gnd.n2869 0.152939
R15505 gnd.n2888 gnd.n2869 0.152939
R15506 gnd.n2889 gnd.n2888 0.152939
R15507 gnd.n2890 gnd.n2889 0.152939
R15508 gnd.n2890 gnd.n2867 0.152939
R15509 gnd.n2896 gnd.n2867 0.152939
R15510 gnd.n2897 gnd.n2896 0.152939
R15511 gnd.n2898 gnd.n2897 0.152939
R15512 gnd.n2898 gnd.n2865 0.152939
R15513 gnd.n3036 gnd.n2865 0.152939
R15514 gnd.n3037 gnd.n3036 0.152939
R15515 gnd.n3038 gnd.n3037 0.152939
R15516 gnd.n3038 gnd.n2859 0.152939
R15517 gnd.n3052 gnd.n2859 0.152939
R15518 gnd.n3053 gnd.n3052 0.152939
R15519 gnd.n3054 gnd.n3053 0.152939
R15520 gnd.n3054 gnd.n2742 0.152939
R15521 gnd.n3068 gnd.n2742 0.152939
R15522 gnd.n3069 gnd.n3068 0.152939
R15523 gnd.n3070 gnd.n3069 0.152939
R15524 gnd.n3070 gnd.n2736 0.152939
R15525 gnd.n3084 gnd.n2736 0.152939
R15526 gnd.n3085 gnd.n3084 0.152939
R15527 gnd.n3086 gnd.n3085 0.152939
R15528 gnd.n3086 gnd.n2728 0.152939
R15529 gnd.n3100 gnd.n2728 0.152939
R15530 gnd.n3101 gnd.n3100 0.152939
R15531 gnd.n3102 gnd.n3101 0.152939
R15532 gnd.n3102 gnd.n2722 0.152939
R15533 gnd.n3116 gnd.n2722 0.152939
R15534 gnd.n3117 gnd.n3116 0.152939
R15535 gnd.n3118 gnd.n3117 0.152939
R15536 gnd.n3118 gnd.n2714 0.152939
R15537 gnd.n3132 gnd.n2714 0.152939
R15538 gnd.n3133 gnd.n3132 0.152939
R15539 gnd.n3134 gnd.n3133 0.152939
R15540 gnd.n3134 gnd.n2708 0.152939
R15541 gnd.n3148 gnd.n2708 0.152939
R15542 gnd.n3149 gnd.n3148 0.152939
R15543 gnd.n3150 gnd.n3149 0.152939
R15544 gnd.n3150 gnd.n2700 0.152939
R15545 gnd.n3164 gnd.n2700 0.152939
R15546 gnd.n3165 gnd.n3164 0.152939
R15547 gnd.n3167 gnd.n3165 0.152939
R15548 gnd.n3167 gnd.n3166 0.152939
R15549 gnd.n3166 gnd.n2695 0.152939
R15550 gnd.n2695 gnd.n2693 0.152939
R15551 gnd.n3183 gnd.n2693 0.152939
R15552 gnd.n3184 gnd.n3183 0.152939
R15553 gnd.n3185 gnd.n3184 0.152939
R15554 gnd.n3185 gnd.n2626 0.152939
R15555 gnd.n3261 gnd.n2626 0.152939
R15556 gnd.n3262 gnd.n3261 0.152939
R15557 gnd.n3326 gnd.n3262 0.152939
R15558 gnd.n1045 gnd.n1044 0.152939
R15559 gnd.n1046 gnd.n1045 0.152939
R15560 gnd.n1047 gnd.n1046 0.152939
R15561 gnd.n1048 gnd.n1047 0.152939
R15562 gnd.n1049 gnd.n1048 0.152939
R15563 gnd.n1050 gnd.n1049 0.152939
R15564 gnd.n1051 gnd.n1050 0.152939
R15565 gnd.n1052 gnd.n1051 0.152939
R15566 gnd.n1053 gnd.n1052 0.152939
R15567 gnd.n1054 gnd.n1053 0.152939
R15568 gnd.n1055 gnd.n1054 0.152939
R15569 gnd.n1056 gnd.n1055 0.152939
R15570 gnd.n1057 gnd.n1056 0.152939
R15571 gnd.n1058 gnd.n1057 0.152939
R15572 gnd.n1059 gnd.n1058 0.152939
R15573 gnd.n1060 gnd.n1059 0.152939
R15574 gnd.n1061 gnd.n1060 0.152939
R15575 gnd.n1064 gnd.n1061 0.152939
R15576 gnd.n1065 gnd.n1064 0.152939
R15577 gnd.n1066 gnd.n1065 0.152939
R15578 gnd.n1067 gnd.n1066 0.152939
R15579 gnd.n1068 gnd.n1067 0.152939
R15580 gnd.n1069 gnd.n1068 0.152939
R15581 gnd.n1070 gnd.n1069 0.152939
R15582 gnd.n1071 gnd.n1070 0.152939
R15583 gnd.n1072 gnd.n1071 0.152939
R15584 gnd.n1073 gnd.n1072 0.152939
R15585 gnd.n1074 gnd.n1073 0.152939
R15586 gnd.n1075 gnd.n1074 0.152939
R15587 gnd.n1076 gnd.n1075 0.152939
R15588 gnd.n1077 gnd.n1076 0.152939
R15589 gnd.n1078 gnd.n1077 0.152939
R15590 gnd.n1079 gnd.n1078 0.152939
R15591 gnd.n1080 gnd.n1079 0.152939
R15592 gnd.n1081 gnd.n1080 0.152939
R15593 gnd.n5033 gnd.n1081 0.152939
R15594 gnd.n5033 gnd.n5032 0.152939
R15595 gnd.n5032 gnd.n5031 0.152939
R15596 gnd.n2989 gnd.n2987 0.152939
R15597 gnd.n2989 gnd.n2988 0.152939
R15598 gnd.n2988 gnd.n1101 0.152939
R15599 gnd.n1102 gnd.n1101 0.152939
R15600 gnd.n1103 gnd.n1102 0.152939
R15601 gnd.n1121 gnd.n1103 0.152939
R15602 gnd.n1122 gnd.n1121 0.152939
R15603 gnd.n1123 gnd.n1122 0.152939
R15604 gnd.n1124 gnd.n1123 0.152939
R15605 gnd.n1141 gnd.n1124 0.152939
R15606 gnd.n1142 gnd.n1141 0.152939
R15607 gnd.n1143 gnd.n1142 0.152939
R15608 gnd.n1144 gnd.n1143 0.152939
R15609 gnd.n1161 gnd.n1144 0.152939
R15610 gnd.n1162 gnd.n1161 0.152939
R15611 gnd.n1163 gnd.n1162 0.152939
R15612 gnd.n1164 gnd.n1163 0.152939
R15613 gnd.n1181 gnd.n1164 0.152939
R15614 gnd.n1182 gnd.n1181 0.152939
R15615 gnd.n1183 gnd.n1182 0.152939
R15616 gnd.n1184 gnd.n1183 0.152939
R15617 gnd.n1203 gnd.n1184 0.152939
R15618 gnd.n1204 gnd.n1203 0.152939
R15619 gnd.n1205 gnd.n1204 0.152939
R15620 gnd.n1206 gnd.n1205 0.152939
R15621 gnd.n1224 gnd.n1206 0.152939
R15622 gnd.n1225 gnd.n1224 0.152939
R15623 gnd.n2759 gnd.n2758 0.152939
R15624 gnd.n2759 gnd.n2750 0.152939
R15625 gnd.n2765 gnd.n2750 0.152939
R15626 gnd.n2766 gnd.n2765 0.152939
R15627 gnd.n2767 gnd.n2766 0.152939
R15628 gnd.n2768 gnd.n2767 0.152939
R15629 gnd.n799 gnd.n798 0.152939
R15630 gnd.n800 gnd.n799 0.152939
R15631 gnd.n805 gnd.n800 0.152939
R15632 gnd.n806 gnd.n805 0.152939
R15633 gnd.n807 gnd.n806 0.152939
R15634 gnd.n808 gnd.n807 0.152939
R15635 gnd.n813 gnd.n808 0.152939
R15636 gnd.n814 gnd.n813 0.152939
R15637 gnd.n815 gnd.n814 0.152939
R15638 gnd.n816 gnd.n815 0.152939
R15639 gnd.n821 gnd.n816 0.152939
R15640 gnd.n822 gnd.n821 0.152939
R15641 gnd.n823 gnd.n822 0.152939
R15642 gnd.n824 gnd.n823 0.152939
R15643 gnd.n829 gnd.n824 0.152939
R15644 gnd.n830 gnd.n829 0.152939
R15645 gnd.n831 gnd.n830 0.152939
R15646 gnd.n832 gnd.n831 0.152939
R15647 gnd.n837 gnd.n832 0.152939
R15648 gnd.n838 gnd.n837 0.152939
R15649 gnd.n839 gnd.n838 0.152939
R15650 gnd.n840 gnd.n839 0.152939
R15651 gnd.n845 gnd.n840 0.152939
R15652 gnd.n846 gnd.n845 0.152939
R15653 gnd.n847 gnd.n846 0.152939
R15654 gnd.n848 gnd.n847 0.152939
R15655 gnd.n853 gnd.n848 0.152939
R15656 gnd.n854 gnd.n853 0.152939
R15657 gnd.n855 gnd.n854 0.152939
R15658 gnd.n856 gnd.n855 0.152939
R15659 gnd.n861 gnd.n856 0.152939
R15660 gnd.n862 gnd.n861 0.152939
R15661 gnd.n863 gnd.n862 0.152939
R15662 gnd.n864 gnd.n863 0.152939
R15663 gnd.n869 gnd.n864 0.152939
R15664 gnd.n870 gnd.n869 0.152939
R15665 gnd.n871 gnd.n870 0.152939
R15666 gnd.n872 gnd.n871 0.152939
R15667 gnd.n877 gnd.n872 0.152939
R15668 gnd.n878 gnd.n877 0.152939
R15669 gnd.n879 gnd.n878 0.152939
R15670 gnd.n880 gnd.n879 0.152939
R15671 gnd.n885 gnd.n880 0.152939
R15672 gnd.n886 gnd.n885 0.152939
R15673 gnd.n887 gnd.n886 0.152939
R15674 gnd.n888 gnd.n887 0.152939
R15675 gnd.n893 gnd.n888 0.152939
R15676 gnd.n894 gnd.n893 0.152939
R15677 gnd.n895 gnd.n894 0.152939
R15678 gnd.n896 gnd.n895 0.152939
R15679 gnd.n901 gnd.n896 0.152939
R15680 gnd.n902 gnd.n901 0.152939
R15681 gnd.n903 gnd.n902 0.152939
R15682 gnd.n904 gnd.n903 0.152939
R15683 gnd.n909 gnd.n904 0.152939
R15684 gnd.n910 gnd.n909 0.152939
R15685 gnd.n911 gnd.n910 0.152939
R15686 gnd.n912 gnd.n911 0.152939
R15687 gnd.n917 gnd.n912 0.152939
R15688 gnd.n918 gnd.n917 0.152939
R15689 gnd.n919 gnd.n918 0.152939
R15690 gnd.n920 gnd.n919 0.152939
R15691 gnd.n925 gnd.n920 0.152939
R15692 gnd.n926 gnd.n925 0.152939
R15693 gnd.n927 gnd.n926 0.152939
R15694 gnd.n928 gnd.n927 0.152939
R15695 gnd.n933 gnd.n928 0.152939
R15696 gnd.n934 gnd.n933 0.152939
R15697 gnd.n935 gnd.n934 0.152939
R15698 gnd.n936 gnd.n935 0.152939
R15699 gnd.n941 gnd.n936 0.152939
R15700 gnd.n942 gnd.n941 0.152939
R15701 gnd.n943 gnd.n942 0.152939
R15702 gnd.n944 gnd.n943 0.152939
R15703 gnd.n949 gnd.n944 0.152939
R15704 gnd.n950 gnd.n949 0.152939
R15705 gnd.n951 gnd.n950 0.152939
R15706 gnd.n952 gnd.n951 0.152939
R15707 gnd.n957 gnd.n952 0.152939
R15708 gnd.n958 gnd.n957 0.152939
R15709 gnd.n959 gnd.n958 0.152939
R15710 gnd.n960 gnd.n959 0.152939
R15711 gnd.n2754 gnd.n960 0.152939
R15712 gnd.n2757 gnd.n2754 0.152939
R15713 gnd.n4269 gnd.n4268 0.152939
R15714 gnd.n4268 gnd.n4267 0.152939
R15715 gnd.n4267 gnd.n1974 0.152939
R15716 gnd.n4263 gnd.n1974 0.152939
R15717 gnd.n4263 gnd.n4262 0.152939
R15718 gnd.n4262 gnd.n4261 0.152939
R15719 gnd.n4261 gnd.n1982 0.152939
R15720 gnd.n4257 gnd.n1982 0.152939
R15721 gnd.n4257 gnd.n4256 0.152939
R15722 gnd.n3386 gnd.n2559 0.152939
R15723 gnd.n3387 gnd.n3386 0.152939
R15724 gnd.n3389 gnd.n3387 0.152939
R15725 gnd.n3389 gnd.n3388 0.152939
R15726 gnd.n3388 gnd.n2534 0.152939
R15727 gnd.n3416 gnd.n2534 0.152939
R15728 gnd.n3417 gnd.n3416 0.152939
R15729 gnd.n3419 gnd.n3417 0.152939
R15730 gnd.n3419 gnd.n3418 0.152939
R15731 gnd.n3418 gnd.n2510 0.152939
R15732 gnd.n3451 gnd.n2510 0.152939
R15733 gnd.n3452 gnd.n3451 0.152939
R15734 gnd.n3456 gnd.n3452 0.152939
R15735 gnd.n3456 gnd.n3455 0.152939
R15736 gnd.n3455 gnd.n3454 0.152939
R15737 gnd.n3454 gnd.n2486 0.152939
R15738 gnd.n3553 gnd.n2486 0.152939
R15739 gnd.n3554 gnd.n3553 0.152939
R15740 gnd.n3556 gnd.n3554 0.152939
R15741 gnd.n3556 gnd.n3555 0.152939
R15742 gnd.n3555 gnd.n2463 0.152939
R15743 gnd.n3613 gnd.n2463 0.152939
R15744 gnd.n3614 gnd.n3613 0.152939
R15745 gnd.n3615 gnd.n3614 0.152939
R15746 gnd.n3615 gnd.n2442 0.152939
R15747 gnd.n3642 gnd.n2442 0.152939
R15748 gnd.n3643 gnd.n3642 0.152939
R15749 gnd.n3648 gnd.n3643 0.152939
R15750 gnd.n3648 gnd.n3647 0.152939
R15751 gnd.n3647 gnd.n3646 0.152939
R15752 gnd.n3646 gnd.n2407 0.152939
R15753 gnd.n3702 gnd.n2407 0.152939
R15754 gnd.n3703 gnd.n3702 0.152939
R15755 gnd.n3705 gnd.n3703 0.152939
R15756 gnd.n3705 gnd.n3704 0.152939
R15757 gnd.n3704 gnd.n2382 0.152939
R15758 gnd.n3756 gnd.n2382 0.152939
R15759 gnd.n3757 gnd.n3756 0.152939
R15760 gnd.n3770 gnd.n3757 0.152939
R15761 gnd.n3770 gnd.n3769 0.152939
R15762 gnd.n3769 gnd.n3768 0.152939
R15763 gnd.n3768 gnd.n3758 0.152939
R15764 gnd.n3764 gnd.n3758 0.152939
R15765 gnd.n3764 gnd.n3763 0.152939
R15766 gnd.n3763 gnd.n2336 0.152939
R15767 gnd.n3856 gnd.n2336 0.152939
R15768 gnd.n3857 gnd.n3856 0.152939
R15769 gnd.n3859 gnd.n3857 0.152939
R15770 gnd.n3859 gnd.n3858 0.152939
R15771 gnd.n3858 gnd.n2314 0.152939
R15772 gnd.n3885 gnd.n2314 0.152939
R15773 gnd.n3886 gnd.n3885 0.152939
R15774 gnd.n3887 gnd.n3886 0.152939
R15775 gnd.n3887 gnd.n2270 0.152939
R15776 gnd.n3929 gnd.n2270 0.152939
R15777 gnd.n3930 gnd.n3929 0.152939
R15778 gnd.n3947 gnd.n3930 0.152939
R15779 gnd.n3947 gnd.n3946 0.152939
R15780 gnd.n3946 gnd.n3945 0.152939
R15781 gnd.n3945 gnd.n3931 0.152939
R15782 gnd.n3941 gnd.n3931 0.152939
R15783 gnd.n3941 gnd.n3940 0.152939
R15784 gnd.n3940 gnd.n3939 0.152939
R15785 gnd.n3939 gnd.n2040 0.152939
R15786 gnd.n4168 gnd.n2040 0.152939
R15787 gnd.n4169 gnd.n4168 0.152939
R15788 gnd.n4170 gnd.n4169 0.152939
R15789 gnd.n4170 gnd.n2029 0.152939
R15790 gnd.n4189 gnd.n2029 0.152939
R15791 gnd.n4190 gnd.n4189 0.152939
R15792 gnd.n4191 gnd.n4190 0.152939
R15793 gnd.n4191 gnd.n2017 0.152939
R15794 gnd.n4210 gnd.n2017 0.152939
R15795 gnd.n4211 gnd.n4210 0.152939
R15796 gnd.n4212 gnd.n4211 0.152939
R15797 gnd.n4212 gnd.n2005 0.152939
R15798 gnd.n4231 gnd.n2005 0.152939
R15799 gnd.n4232 gnd.n4231 0.152939
R15800 gnd.n4234 gnd.n4232 0.152939
R15801 gnd.n4234 gnd.n4233 0.152939
R15802 gnd.n4233 gnd.n1994 0.152939
R15803 gnd.n4255 gnd.n1994 0.152939
R15804 gnd.n3247 gnd.n2631 0.152939
R15805 gnd.n3247 gnd.n3246 0.152939
R15806 gnd.n3246 gnd.n3245 0.152939
R15807 gnd.n3245 gnd.n2638 0.152939
R15808 gnd.n3241 gnd.n2638 0.152939
R15809 gnd.n3241 gnd.n3240 0.152939
R15810 gnd.n3240 gnd.n2645 0.152939
R15811 gnd.n3236 gnd.n2645 0.152939
R15812 gnd.n3236 gnd.n3235 0.152939
R15813 gnd.n3092 gnd.n2731 0.152939
R15814 gnd.n3093 gnd.n3092 0.152939
R15815 gnd.n3094 gnd.n3093 0.152939
R15816 gnd.n3094 gnd.n2725 0.152939
R15817 gnd.n3108 gnd.n2725 0.152939
R15818 gnd.n3109 gnd.n3108 0.152939
R15819 gnd.n3110 gnd.n3109 0.152939
R15820 gnd.n3110 gnd.n2718 0.152939
R15821 gnd.n3124 gnd.n2718 0.152939
R15822 gnd.n3125 gnd.n3124 0.152939
R15823 gnd.n3126 gnd.n3125 0.152939
R15824 gnd.n3126 gnd.n2711 0.152939
R15825 gnd.n3140 gnd.n2711 0.152939
R15826 gnd.n3141 gnd.n3140 0.152939
R15827 gnd.n3142 gnd.n3141 0.152939
R15828 gnd.n3142 gnd.n2704 0.152939
R15829 gnd.n3156 gnd.n2704 0.152939
R15830 gnd.n3157 gnd.n3156 0.152939
R15831 gnd.n3158 gnd.n3157 0.152939
R15832 gnd.n3158 gnd.n2697 0.152939
R15833 gnd.n3173 gnd.n2697 0.152939
R15834 gnd.n3174 gnd.n3173 0.152939
R15835 gnd.n3175 gnd.n3174 0.152939
R15836 gnd.n3175 gnd.n2691 0.152939
R15837 gnd.n3193 gnd.n2691 0.152939
R15838 gnd.n3193 gnd.n3192 0.152939
R15839 gnd.n3192 gnd.n3191 0.152939
R15840 gnd.n3191 gnd.n2630 0.152939
R15841 gnd.n3255 gnd.n2630 0.152939
R15842 gnd.n3255 gnd.n3254 0.152939
R15843 gnd.n3254 gnd.n3253 0.152939
R15844 gnd.n3380 gnd.n3378 0.152939
R15845 gnd.n3380 gnd.n3379 0.152939
R15846 gnd.n3379 gnd.n2543 0.152939
R15847 gnd.n3407 gnd.n2543 0.152939
R15848 gnd.n3408 gnd.n3407 0.152939
R15849 gnd.n3410 gnd.n3408 0.152939
R15850 gnd.n3410 gnd.n3409 0.152939
R15851 gnd.n3409 gnd.n2517 0.152939
R15852 gnd.n3443 gnd.n2517 0.152939
R15853 gnd.n3444 gnd.n3443 0.152939
R15854 gnd.n3445 gnd.n3444 0.152939
R15855 gnd.n3445 gnd.n2502 0.152939
R15856 gnd.n3463 gnd.n2502 0.152939
R15857 gnd.n3464 gnd.n3463 0.152939
R15858 gnd.n3466 gnd.n3464 0.152939
R15859 gnd.n3466 gnd.n3465 0.152939
R15860 gnd.n3465 gnd.n1531 0.152939
R15861 gnd.n4722 gnd.n1531 0.152939
R15862 gnd.n4722 gnd.n4721 0.152939
R15863 gnd.n4721 gnd.n4720 0.152939
R15864 gnd.n4720 gnd.n1532 0.152939
R15865 gnd.n4716 gnd.n1532 0.152939
R15866 gnd.n4716 gnd.n4715 0.152939
R15867 gnd.n4715 gnd.n4714 0.152939
R15868 gnd.n4714 gnd.n1537 0.152939
R15869 gnd.n4710 gnd.n1537 0.152939
R15870 gnd.n4710 gnd.n4709 0.152939
R15871 gnd.n4709 gnd.n4708 0.152939
R15872 gnd.n4708 gnd.n1542 0.152939
R15873 gnd.n4704 gnd.n1542 0.152939
R15874 gnd.n4704 gnd.n4703 0.152939
R15875 gnd.n4703 gnd.n4702 0.152939
R15876 gnd.n4702 gnd.n1547 0.152939
R15877 gnd.n4698 gnd.n1547 0.152939
R15878 gnd.n4698 gnd.n4697 0.152939
R15879 gnd.n4697 gnd.n4696 0.152939
R15880 gnd.n4696 gnd.n1552 0.152939
R15881 gnd.n4692 gnd.n1552 0.152939
R15882 gnd.n4692 gnd.n4691 0.152939
R15883 gnd.n4691 gnd.n4690 0.152939
R15884 gnd.n4690 gnd.n1557 0.152939
R15885 gnd.n4686 gnd.n1557 0.152939
R15886 gnd.n4686 gnd.n4685 0.152939
R15887 gnd.n4685 gnd.n4684 0.152939
R15888 gnd.n4684 gnd.n1562 0.152939
R15889 gnd.n4680 gnd.n1562 0.152939
R15890 gnd.n4680 gnd.n4679 0.152939
R15891 gnd.n4679 gnd.n4678 0.152939
R15892 gnd.n4678 gnd.n1567 0.152939
R15893 gnd.n4674 gnd.n1567 0.152939
R15894 gnd.n4674 gnd.n4673 0.152939
R15895 gnd.n4673 gnd.n4672 0.152939
R15896 gnd.n4672 gnd.n1572 0.152939
R15897 gnd.n4668 gnd.n1572 0.152939
R15898 gnd.n4668 gnd.n4667 0.152939
R15899 gnd.n4667 gnd.n4666 0.152939
R15900 gnd.n4666 gnd.n1577 0.152939
R15901 gnd.n4662 gnd.n1577 0.152939
R15902 gnd.n4662 gnd.n4661 0.152939
R15903 gnd.n4661 gnd.n4660 0.152939
R15904 gnd.n4660 gnd.n1582 0.152939
R15905 gnd.n4656 gnd.n1582 0.152939
R15906 gnd.n4656 gnd.n4655 0.152939
R15907 gnd.n4655 gnd.n4654 0.152939
R15908 gnd.n4654 gnd.n1587 0.152939
R15909 gnd.n4650 gnd.n1587 0.152939
R15910 gnd.n4650 gnd.n4649 0.152939
R15911 gnd.n4649 gnd.n4648 0.152939
R15912 gnd.n4648 gnd.n1592 0.152939
R15913 gnd.n4644 gnd.n1592 0.152939
R15914 gnd.n4644 gnd.n4643 0.152939
R15915 gnd.n4643 gnd.n4642 0.152939
R15916 gnd.n4642 gnd.n1597 0.152939
R15917 gnd.n4638 gnd.n1597 0.152939
R15918 gnd.n4638 gnd.n4637 0.152939
R15919 gnd.n4637 gnd.n4636 0.152939
R15920 gnd.n4636 gnd.n1602 0.152939
R15921 gnd.n4632 gnd.n1602 0.152939
R15922 gnd.n4632 gnd.n4631 0.152939
R15923 gnd.n4631 gnd.n4630 0.152939
R15924 gnd.n4630 gnd.n1607 0.152939
R15925 gnd.n1610 gnd.n1607 0.152939
R15926 gnd.n1885 gnd.n1879 0.152939
R15927 gnd.n1879 gnd.n1654 0.152939
R15928 gnd.n4600 gnd.n1654 0.152939
R15929 gnd.n4600 gnd.n4599 0.152939
R15930 gnd.n4599 gnd.n4598 0.152939
R15931 gnd.n4598 gnd.n1655 0.152939
R15932 gnd.n4594 gnd.n1655 0.152939
R15933 gnd.n4594 gnd.n4593 0.152939
R15934 gnd.n4593 gnd.n4592 0.152939
R15935 gnd.n4592 gnd.n1660 0.152939
R15936 gnd.n4588 gnd.n1660 0.152939
R15937 gnd.n4588 gnd.n4587 0.152939
R15938 gnd.n4587 gnd.n4586 0.152939
R15939 gnd.n4586 gnd.n1665 0.152939
R15940 gnd.n4582 gnd.n1665 0.152939
R15941 gnd.n4582 gnd.n4581 0.152939
R15942 gnd.n4581 gnd.n4580 0.152939
R15943 gnd.n4580 gnd.n1670 0.152939
R15944 gnd.n4576 gnd.n1670 0.152939
R15945 gnd.n4576 gnd.n4575 0.152939
R15946 gnd.n4575 gnd.n4574 0.152939
R15947 gnd.n4574 gnd.n1675 0.152939
R15948 gnd.n4570 gnd.n1675 0.152939
R15949 gnd.n4570 gnd.n4569 0.152939
R15950 gnd.n4569 gnd.n4568 0.152939
R15951 gnd.n4568 gnd.n1680 0.152939
R15952 gnd.n4564 gnd.n1680 0.152939
R15953 gnd.n4564 gnd.n318 0.152939
R15954 gnd.n7410 gnd.n318 0.152939
R15955 gnd.n7410 gnd.n7409 0.152939
R15956 gnd.n7409 gnd.n7408 0.152939
R15957 gnd.n7408 gnd.n319 0.152939
R15958 gnd.n7404 gnd.n319 0.152939
R15959 gnd.n7404 gnd.n7403 0.152939
R15960 gnd.n7403 gnd.n7402 0.152939
R15961 gnd.n7402 gnd.n324 0.152939
R15962 gnd.n324 gnd.n293 0.152939
R15963 gnd.n7425 gnd.n293 0.152939
R15964 gnd.n7426 gnd.n7425 0.152939
R15965 gnd.n7427 gnd.n7426 0.152939
R15966 gnd.n7427 gnd.n277 0.152939
R15967 gnd.n7441 gnd.n277 0.152939
R15968 gnd.n7442 gnd.n7441 0.152939
R15969 gnd.n7443 gnd.n7442 0.152939
R15970 gnd.n7443 gnd.n262 0.152939
R15971 gnd.n7457 gnd.n262 0.152939
R15972 gnd.n7458 gnd.n7457 0.152939
R15973 gnd.n7459 gnd.n7458 0.152939
R15974 gnd.n7459 gnd.n246 0.152939
R15975 gnd.n7473 gnd.n246 0.152939
R15976 gnd.n7474 gnd.n7473 0.152939
R15977 gnd.n7475 gnd.n7474 0.152939
R15978 gnd.n7475 gnd.n232 0.152939
R15979 gnd.n7489 gnd.n232 0.152939
R15980 gnd.n7490 gnd.n7489 0.152939
R15981 gnd.n7491 gnd.n7490 0.152939
R15982 gnd.n7491 gnd.n217 0.152939
R15983 gnd.n7505 gnd.n217 0.152939
R15984 gnd.n7506 gnd.n7505 0.152939
R15985 gnd.n7575 gnd.n7506 0.152939
R15986 gnd.n7575 gnd.n7574 0.152939
R15987 gnd.n7574 gnd.n7573 0.152939
R15988 gnd.n7573 gnd.n7507 0.152939
R15989 gnd.n7569 gnd.n7507 0.152939
R15990 gnd.n7568 gnd.n7509 0.152939
R15991 gnd.n7564 gnd.n7509 0.152939
R15992 gnd.n7564 gnd.n7563 0.152939
R15993 gnd.n7563 gnd.n7562 0.152939
R15994 gnd.n7562 gnd.n7515 0.152939
R15995 gnd.n7558 gnd.n7515 0.152939
R15996 gnd.n7558 gnd.n7557 0.152939
R15997 gnd.n7557 gnd.n7556 0.152939
R15998 gnd.n7556 gnd.n7523 0.152939
R15999 gnd.n7552 gnd.n7523 0.152939
R16000 gnd.n7552 gnd.n7551 0.152939
R16001 gnd.n7551 gnd.n7550 0.152939
R16002 gnd.n7550 gnd.n7531 0.152939
R16003 gnd.n7546 gnd.n7531 0.152939
R16004 gnd.n7546 gnd.n7545 0.152939
R16005 gnd.n7545 gnd.n7544 0.152939
R16006 gnd.n7544 gnd.n117 0.152939
R16007 gnd.n7670 gnd.n117 0.152939
R16008 gnd.n4280 gnd.n4279 0.152939
R16009 gnd.n4281 gnd.n4280 0.152939
R16010 gnd.n4281 gnd.n1830 0.152939
R16011 gnd.n4340 gnd.n1830 0.152939
R16012 gnd.n4341 gnd.n4340 0.152939
R16013 gnd.n4343 gnd.n4341 0.152939
R16014 gnd.n4343 gnd.n4342 0.152939
R16015 gnd.n4342 gnd.n1792 0.152939
R16016 gnd.n4372 gnd.n1792 0.152939
R16017 gnd.n4373 gnd.n4372 0.152939
R16018 gnd.n4375 gnd.n4373 0.152939
R16019 gnd.n4375 gnd.n4374 0.152939
R16020 gnd.n4374 gnd.n1766 0.152939
R16021 gnd.n4404 gnd.n1766 0.152939
R16022 gnd.n4405 gnd.n4404 0.152939
R16023 gnd.n4407 gnd.n4405 0.152939
R16024 gnd.n4407 gnd.n4406 0.152939
R16025 gnd.n4406 gnd.n1740 0.152939
R16026 gnd.n4436 gnd.n1740 0.152939
R16027 gnd.n4437 gnd.n4436 0.152939
R16028 gnd.n4445 gnd.n4437 0.152939
R16029 gnd.n4445 gnd.n4444 0.152939
R16030 gnd.n4444 gnd.n4443 0.152939
R16031 gnd.n4443 gnd.n4438 0.152939
R16032 gnd.n4438 gnd.n1693 0.152939
R16033 gnd.n4556 gnd.n1693 0.152939
R16034 gnd.n4556 gnd.n4555 0.152939
R16035 gnd.n4555 gnd.n4554 0.152939
R16036 gnd.n4554 gnd.n1694 0.152939
R16037 gnd.n4550 gnd.n1694 0.152939
R16038 gnd.n4550 gnd.n75 0.152939
R16039 gnd.n7719 gnd.n75 0.152939
R16040 gnd.n7719 gnd.n7718 0.152939
R16041 gnd.n7718 gnd.n77 0.152939
R16042 gnd.n7714 gnd.n77 0.152939
R16043 gnd.n7714 gnd.n7713 0.152939
R16044 gnd.n7713 gnd.n7712 0.152939
R16045 gnd.n7712 gnd.n82 0.152939
R16046 gnd.n7708 gnd.n82 0.152939
R16047 gnd.n7708 gnd.n7707 0.152939
R16048 gnd.n7707 gnd.n7706 0.152939
R16049 gnd.n7706 gnd.n87 0.152939
R16050 gnd.n7702 gnd.n87 0.152939
R16051 gnd.n7702 gnd.n7701 0.152939
R16052 gnd.n7701 gnd.n7700 0.152939
R16053 gnd.n7700 gnd.n92 0.152939
R16054 gnd.n7696 gnd.n92 0.152939
R16055 gnd.n7696 gnd.n7695 0.152939
R16056 gnd.n7695 gnd.n7694 0.152939
R16057 gnd.n7694 gnd.n97 0.152939
R16058 gnd.n7690 gnd.n97 0.152939
R16059 gnd.n7690 gnd.n7689 0.152939
R16060 gnd.n7689 gnd.n7688 0.152939
R16061 gnd.n7688 gnd.n102 0.152939
R16062 gnd.n7684 gnd.n102 0.152939
R16063 gnd.n7684 gnd.n7683 0.152939
R16064 gnd.n7683 gnd.n7682 0.152939
R16065 gnd.n7682 gnd.n107 0.152939
R16066 gnd.n7678 gnd.n107 0.152939
R16067 gnd.n7678 gnd.n7677 0.152939
R16068 gnd.n7677 gnd.n7676 0.152939
R16069 gnd.n7676 gnd.n112 0.152939
R16070 gnd.n7672 gnd.n112 0.152939
R16071 gnd.n7672 gnd.n7671 0.152939
R16072 gnd.n4269 gnd.n1837 0.151415
R16073 gnd.n3252 gnd.n2631 0.151415
R16074 gnd.n2851 gnd.n2771 0.14989
R16075 gnd.n4460 gnd.n302 0.14989
R16076 gnd.n3078 gnd.n3077 0.145814
R16077 gnd.n3078 gnd.n2731 0.145814
R16078 gnd.n5957 gnd.n5349 0.0767195
R16079 gnd.n5873 gnd.n5349 0.0767195
R16080 gnd.n3377 gnd.n3376 0.063
R16081 gnd.n1887 gnd.n1886 0.063
R16082 gnd.n6480 gnd.n5138 0.0477147
R16083 gnd.n5623 gnd.n5519 0.0442063
R16084 gnd.n5637 gnd.n5519 0.0442063
R16085 gnd.n5638 gnd.n5637 0.0442063
R16086 gnd.n5639 gnd.n5638 0.0442063
R16087 gnd.n5639 gnd.n5507 0.0442063
R16088 gnd.n5653 gnd.n5507 0.0442063
R16089 gnd.n5654 gnd.n5653 0.0442063
R16090 gnd.n5655 gnd.n5654 0.0442063
R16091 gnd.n5655 gnd.n5494 0.0442063
R16092 gnd.n5751 gnd.n5494 0.0442063
R16093 gnd.n5754 gnd.n5753 0.0344674
R16094 gnd.n4273 gnd.n1843 0.0344674
R16095 gnd.n3251 gnd.n2632 0.0344674
R16096 gnd.n5487 gnd.n5486 0.0269946
R16097 gnd.n5764 gnd.n5484 0.0269946
R16098 gnd.n5763 gnd.n5485 0.0269946
R16099 gnd.n5783 gnd.n5466 0.0269946
R16100 gnd.n5785 gnd.n5784 0.0269946
R16101 gnd.n5786 gnd.n5464 0.0269946
R16102 gnd.n5793 gnd.n5789 0.0269946
R16103 gnd.n5792 gnd.n5791 0.0269946
R16104 gnd.n5790 gnd.n5443 0.0269946
R16105 gnd.n5817 gnd.n5444 0.0269946
R16106 gnd.n5816 gnd.n5445 0.0269946
R16107 gnd.n5849 gnd.n5419 0.0269946
R16108 gnd.n5851 gnd.n5850 0.0269946
R16109 gnd.n5852 gnd.n5411 0.0269946
R16110 gnd.n5415 gnd.n5412 0.0269946
R16111 gnd.n5862 gnd.n5413 0.0269946
R16112 gnd.n5861 gnd.n5414 0.0269946
R16113 gnd.n5907 gnd.n5387 0.0269946
R16114 gnd.n5909 gnd.n5908 0.0269946
R16115 gnd.n5918 gnd.n5380 0.0269946
R16116 gnd.n5920 gnd.n5919 0.0269946
R16117 gnd.n5921 gnd.n5378 0.0269946
R16118 gnd.n5928 gnd.n5924 0.0269946
R16119 gnd.n5927 gnd.n5926 0.0269946
R16120 gnd.n5925 gnd.n5357 0.0269946
R16121 gnd.n5950 gnd.n5358 0.0269946
R16122 gnd.n5949 gnd.n5359 0.0269946
R16123 gnd.n5992 gnd.n5272 0.0269946
R16124 gnd.n5994 gnd.n5993 0.0269946
R16125 gnd.n6003 gnd.n5265 0.0269946
R16126 gnd.n6005 gnd.n6004 0.0269946
R16127 gnd.n6006 gnd.n5263 0.0269946
R16128 gnd.n6013 gnd.n6009 0.0269946
R16129 gnd.n6012 gnd.n6011 0.0269946
R16130 gnd.n6010 gnd.n5242 0.0269946
R16131 gnd.n6035 gnd.n5243 0.0269946
R16132 gnd.n6034 gnd.n5244 0.0269946
R16133 gnd.n6078 gnd.n5218 0.0269946
R16134 gnd.n6080 gnd.n6079 0.0269946
R16135 gnd.n6089 gnd.n5211 0.0269946
R16136 gnd.n6091 gnd.n6090 0.0269946
R16137 gnd.n6092 gnd.n5209 0.0269946
R16138 gnd.n6098 gnd.n6095 0.0269946
R16139 gnd.n6097 gnd.n6096 0.0269946
R16140 gnd.n6120 gnd.n5188 0.0269946
R16141 gnd.n6119 gnd.n5189 0.0269946
R16142 gnd.n6139 gnd.n5175 0.0269946
R16143 gnd.n6141 gnd.n6140 0.0269946
R16144 gnd.n6400 gnd.n981 0.0269946
R16145 gnd.n6402 gnd.n982 0.0269946
R16146 gnd.n6404 gnd.n6403 0.0269946
R16147 gnd.n6408 gnd.n6407 0.0269946
R16148 gnd.n1888 gnd.n1887 0.0246168
R16149 gnd.n3377 gnd.n2568 0.0246168
R16150 gnd.n5753 gnd.n5752 0.0202011
R16151 gnd.n1889 gnd.n1888 0.0174837
R16152 gnd.n1897 gnd.n1889 0.0174837
R16153 gnd.n1897 gnd.n1896 0.0174837
R16154 gnd.n1896 gnd.n1890 0.0174837
R16155 gnd.n1890 gnd.n1874 0.0174837
R16156 gnd.n1905 gnd.n1874 0.0174837
R16157 gnd.n1907 gnd.n1905 0.0174837
R16158 gnd.n1907 gnd.n1906 0.0174837
R16159 gnd.n1906 gnd.n1869 0.0174837
R16160 gnd.n1916 gnd.n1869 0.0174837
R16161 gnd.n1916 gnd.n1915 0.0174837
R16162 gnd.n1915 gnd.n1870 0.0174837
R16163 gnd.n1870 gnd.n1865 0.0174837
R16164 gnd.n1924 gnd.n1865 0.0174837
R16165 gnd.n1926 gnd.n1924 0.0174837
R16166 gnd.n1926 gnd.n1925 0.0174837
R16167 gnd.n1925 gnd.n1860 0.0174837
R16168 gnd.n1935 gnd.n1860 0.0174837
R16169 gnd.n1935 gnd.n1934 0.0174837
R16170 gnd.n1934 gnd.n1861 0.0174837
R16171 gnd.n1861 gnd.n1856 0.0174837
R16172 gnd.n1943 gnd.n1856 0.0174837
R16173 gnd.n1945 gnd.n1943 0.0174837
R16174 gnd.n1945 gnd.n1944 0.0174837
R16175 gnd.n1944 gnd.n1851 0.0174837
R16176 gnd.n1954 gnd.n1851 0.0174837
R16177 gnd.n1954 gnd.n1953 0.0174837
R16178 gnd.n1953 gnd.n1852 0.0174837
R16179 gnd.n1852 gnd.n1847 0.0174837
R16180 gnd.n1962 gnd.n1847 0.0174837
R16181 gnd.n1964 gnd.n1962 0.0174837
R16182 gnd.n1964 gnd.n1963 0.0174837
R16183 gnd.n1963 gnd.n1842 0.0174837
R16184 gnd.n4274 gnd.n1842 0.0174837
R16185 gnd.n4274 gnd.n4273 0.0174837
R16186 gnd.n2574 gnd.n2568 0.0174837
R16187 gnd.n3372 gnd.n2574 0.0174837
R16188 gnd.n3372 gnd.n3371 0.0174837
R16189 gnd.n3371 gnd.n2575 0.0174837
R16190 gnd.n3368 gnd.n2575 0.0174837
R16191 gnd.n3368 gnd.n3367 0.0174837
R16192 gnd.n3367 gnd.n2580 0.0174837
R16193 gnd.n3364 gnd.n2580 0.0174837
R16194 gnd.n3364 gnd.n3363 0.0174837
R16195 gnd.n3363 gnd.n2584 0.0174837
R16196 gnd.n3360 gnd.n2584 0.0174837
R16197 gnd.n3360 gnd.n3359 0.0174837
R16198 gnd.n3359 gnd.n2588 0.0174837
R16199 gnd.n3356 gnd.n2588 0.0174837
R16200 gnd.n3356 gnd.n3355 0.0174837
R16201 gnd.n3355 gnd.n2594 0.0174837
R16202 gnd.n3352 gnd.n2594 0.0174837
R16203 gnd.n3352 gnd.n3351 0.0174837
R16204 gnd.n3351 gnd.n2598 0.0174837
R16205 gnd.n3348 gnd.n2598 0.0174837
R16206 gnd.n3348 gnd.n3347 0.0174837
R16207 gnd.n3347 gnd.n2602 0.0174837
R16208 gnd.n3344 gnd.n2602 0.0174837
R16209 gnd.n3344 gnd.n3343 0.0174837
R16210 gnd.n3343 gnd.n2606 0.0174837
R16211 gnd.n3340 gnd.n2606 0.0174837
R16212 gnd.n3340 gnd.n3339 0.0174837
R16213 gnd.n3339 gnd.n2612 0.0174837
R16214 gnd.n3336 gnd.n2612 0.0174837
R16215 gnd.n3336 gnd.n3335 0.0174837
R16216 gnd.n3335 gnd.n2616 0.0174837
R16217 gnd.n2620 gnd.n2616 0.0174837
R16218 gnd.n2662 gnd.n2620 0.0174837
R16219 gnd.n2662 gnd.n2622 0.0174837
R16220 gnd.n2632 gnd.n2622 0.0174837
R16221 gnd.n5752 gnd.n5751 0.0148637
R16222 gnd.n6398 gnd.n6397 0.0144266
R16223 gnd.n6397 gnd.n980 0.0130679
R16224 gnd.n5754 gnd.n5487 0.00797283
R16225 gnd.n5486 gnd.n5484 0.00797283
R16226 gnd.n5764 gnd.n5763 0.00797283
R16227 gnd.n5485 gnd.n5466 0.00797283
R16228 gnd.n5784 gnd.n5783 0.00797283
R16229 gnd.n5786 gnd.n5785 0.00797283
R16230 gnd.n5789 gnd.n5464 0.00797283
R16231 gnd.n5793 gnd.n5792 0.00797283
R16232 gnd.n5791 gnd.n5790 0.00797283
R16233 gnd.n5444 gnd.n5443 0.00797283
R16234 gnd.n5817 gnd.n5816 0.00797283
R16235 gnd.n5445 gnd.n5419 0.00797283
R16236 gnd.n5850 gnd.n5849 0.00797283
R16237 gnd.n5852 gnd.n5851 0.00797283
R16238 gnd.n5415 gnd.n5411 0.00797283
R16239 gnd.n5413 gnd.n5412 0.00797283
R16240 gnd.n5862 gnd.n5861 0.00797283
R16241 gnd.n5414 gnd.n5387 0.00797283
R16242 gnd.n5909 gnd.n5907 0.00797283
R16243 gnd.n5908 gnd.n5380 0.00797283
R16244 gnd.n5919 gnd.n5918 0.00797283
R16245 gnd.n5921 gnd.n5920 0.00797283
R16246 gnd.n5924 gnd.n5378 0.00797283
R16247 gnd.n5928 gnd.n5927 0.00797283
R16248 gnd.n5926 gnd.n5925 0.00797283
R16249 gnd.n5358 gnd.n5357 0.00797283
R16250 gnd.n5950 gnd.n5949 0.00797283
R16251 gnd.n5359 gnd.n5272 0.00797283
R16252 gnd.n5994 gnd.n5992 0.00797283
R16253 gnd.n5993 gnd.n5265 0.00797283
R16254 gnd.n6004 gnd.n6003 0.00797283
R16255 gnd.n6006 gnd.n6005 0.00797283
R16256 gnd.n6009 gnd.n5263 0.00797283
R16257 gnd.n6013 gnd.n6012 0.00797283
R16258 gnd.n6011 gnd.n6010 0.00797283
R16259 gnd.n5243 gnd.n5242 0.00797283
R16260 gnd.n6035 gnd.n6034 0.00797283
R16261 gnd.n5244 gnd.n5218 0.00797283
R16262 gnd.n6080 gnd.n6078 0.00797283
R16263 gnd.n6079 gnd.n5211 0.00797283
R16264 gnd.n6090 gnd.n6089 0.00797283
R16265 gnd.n6092 gnd.n6091 0.00797283
R16266 gnd.n6095 gnd.n5209 0.00797283
R16267 gnd.n6098 gnd.n6097 0.00797283
R16268 gnd.n6096 gnd.n5188 0.00797283
R16269 gnd.n6120 gnd.n6119 0.00797283
R16270 gnd.n5189 gnd.n5175 0.00797283
R16271 gnd.n6140 gnd.n6139 0.00797283
R16272 gnd.n6398 gnd.n6141 0.00797283
R16273 gnd.n6400 gnd.n980 0.00797283
R16274 gnd.n6402 gnd.n981 0.00797283
R16275 gnd.n6403 gnd.n982 0.00797283
R16276 gnd.n6408 gnd.n6404 0.00797283
R16277 gnd.n6407 gnd.n5138 0.00797283
R16278 gnd.n4502 gnd.n319 0.00433921
R16279 gnd.n3084 gnd.n2735 0.00433921
R16280 gnd.n337 gnd.n302 0.00354878
R16281 gnd.n2851 gnd.n2768 0.00354878
R16282 gnd.n1843 gnd.n1837 0.000839674
R16283 gnd.n3252 gnd.n3251 0.000839674
R16284 a_n8300_8799.n225 a_n8300_8799.t145 485.149
R16285 a_n8300_8799.n244 a_n8300_8799.t38 485.149
R16286 a_n8300_8799.n264 a_n8300_8799.t120 485.149
R16287 a_n8300_8799.n164 a_n8300_8799.t103 485.149
R16288 a_n8300_8799.n183 a_n8300_8799.t119 485.149
R16289 a_n8300_8799.n203 a_n8300_8799.t121 485.149
R16290 a_n8300_8799.n56 a_n8300_8799.t85 485.135
R16291 a_n8300_8799.n237 a_n8300_8799.t61 464.166
R16292 a_n8300_8799.n219 a_n8300_8799.t140 464.166
R16293 a_n8300_8799.n236 a_n8300_8799.t102 464.166
R16294 a_n8300_8799.n235 a_n8300_8799.t99 464.166
R16295 a_n8300_8799.n220 a_n8300_8799.t39 464.166
R16296 a_n8300_8799.n234 a_n8300_8799.t107 464.166
R16297 a_n8300_8799.n233 a_n8300_8799.t106 464.166
R16298 a_n8300_8799.n221 a_n8300_8799.t41 464.166
R16299 a_n8300_8799.n232 a_n8300_8799.t40 464.166
R16300 a_n8300_8799.n231 a_n8300_8799.t128 464.166
R16301 a_n8300_8799.n222 a_n8300_8799.t56 464.166
R16302 a_n8300_8799.n230 a_n8300_8799.t45 464.166
R16303 a_n8300_8799.n229 a_n8300_8799.t132 464.166
R16304 a_n8300_8799.n223 a_n8300_8799.t84 464.166
R16305 a_n8300_8799.n228 a_n8300_8799.t60 464.166
R16306 a_n8300_8799.n227 a_n8300_8799.t152 464.166
R16307 a_n8300_8799.n224 a_n8300_8799.t101 464.166
R16308 a_n8300_8799.n226 a_n8300_8799.t63 464.166
R16309 a_n8300_8799.n71 a_n8300_8799.t96 485.135
R16310 a_n8300_8799.n256 a_n8300_8799.t72 464.166
R16311 a_n8300_8799.n238 a_n8300_8799.t154 464.166
R16312 a_n8300_8799.n255 a_n8300_8799.t117 464.166
R16313 a_n8300_8799.n254 a_n8300_8799.t116 464.166
R16314 a_n8300_8799.n239 a_n8300_8799.t50 464.166
R16315 a_n8300_8799.n253 a_n8300_8799.t124 464.166
R16316 a_n8300_8799.n252 a_n8300_8799.t123 464.166
R16317 a_n8300_8799.n240 a_n8300_8799.t52 464.166
R16318 a_n8300_8799.n251 a_n8300_8799.t51 464.166
R16319 a_n8300_8799.n250 a_n8300_8799.t144 464.166
R16320 a_n8300_8799.n241 a_n8300_8799.t69 464.166
R16321 a_n8300_8799.n249 a_n8300_8799.t55 464.166
R16322 a_n8300_8799.n248 a_n8300_8799.t146 464.166
R16323 a_n8300_8799.n242 a_n8300_8799.t97 464.166
R16324 a_n8300_8799.n247 a_n8300_8799.t73 464.166
R16325 a_n8300_8799.n246 a_n8300_8799.t43 464.166
R16326 a_n8300_8799.n243 a_n8300_8799.t118 464.166
R16327 a_n8300_8799.n245 a_n8300_8799.t74 464.166
R16328 a_n8300_8799.n86 a_n8300_8799.t127 485.135
R16329 a_n8300_8799.n276 a_n8300_8799.t58 464.166
R16330 a_n8300_8799.n258 a_n8300_8799.t105 464.166
R16331 a_n8300_8799.n275 a_n8300_8799.t44 464.166
R16332 a_n8300_8799.n274 a_n8300_8799.t64 464.166
R16333 a_n8300_8799.n259 a_n8300_8799.t149 464.166
R16334 a_n8300_8799.n273 a_n8300_8799.t115 464.166
R16335 a_n8300_8799.n272 a_n8300_8799.t143 464.166
R16336 a_n8300_8799.n260 a_n8300_8799.t95 464.166
R16337 a_n8300_8799.n271 a_n8300_8799.t122 464.166
R16338 a_n8300_8799.n270 a_n8300_8799.t54 464.166
R16339 a_n8300_8799.n261 a_n8300_8799.t139 464.166
R16340 a_n8300_8799.n269 a_n8300_8799.t78 464.166
R16341 a_n8300_8799.n268 a_n8300_8799.t133 464.166
R16342 a_n8300_8799.n262 a_n8300_8799.t62 464.166
R16343 a_n8300_8799.n267 a_n8300_8799.t110 464.166
R16344 a_n8300_8799.n266 a_n8300_8799.t49 464.166
R16345 a_n8300_8799.n263 a_n8300_8799.t92 464.166
R16346 a_n8300_8799.n265 a_n8300_8799.t71 464.166
R16347 a_n8300_8799.n165 a_n8300_8799.t142 464.166
R16348 a_n8300_8799.n166 a_n8300_8799.t65 464.166
R16349 a_n8300_8799.n167 a_n8300_8799.t98 464.166
R16350 a_n8300_8799.n168 a_n8300_8799.t135 464.166
R16351 a_n8300_8799.n163 a_n8300_8799.t137 464.166
R16352 a_n8300_8799.n169 a_n8300_8799.t83 464.166
R16353 a_n8300_8799.n170 a_n8300_8799.t114 464.166
R16354 a_n8300_8799.n171 a_n8300_8799.t134 464.166
R16355 a_n8300_8799.n172 a_n8300_8799.t81 464.166
R16356 a_n8300_8799.n162 a_n8300_8799.t82 464.166
R16357 a_n8300_8799.n173 a_n8300_8799.t111 464.166
R16358 a_n8300_8799.n161 a_n8300_8799.t67 464.166
R16359 a_n8300_8799.n174 a_n8300_8799.t68 464.166
R16360 a_n8300_8799.n175 a_n8300_8799.t108 464.166
R16361 a_n8300_8799.n176 a_n8300_8799.t36 464.166
R16362 a_n8300_8799.n177 a_n8300_8799.t66 464.166
R16363 a_n8300_8799.n160 a_n8300_8799.t88 464.166
R16364 a_n8300_8799.n178 a_n8300_8799.t136 464.166
R16365 a_n8300_8799.n184 a_n8300_8799.t155 464.166
R16366 a_n8300_8799.n185 a_n8300_8799.t75 464.166
R16367 a_n8300_8799.n186 a_n8300_8799.t112 464.166
R16368 a_n8300_8799.n187 a_n8300_8799.t150 464.166
R16369 a_n8300_8799.n182 a_n8300_8799.t153 464.166
R16370 a_n8300_8799.n188 a_n8300_8799.t93 464.166
R16371 a_n8300_8799.n189 a_n8300_8799.t131 464.166
R16372 a_n8300_8799.n190 a_n8300_8799.t148 464.166
R16373 a_n8300_8799.n191 a_n8300_8799.t89 464.166
R16374 a_n8300_8799.n181 a_n8300_8799.t90 464.166
R16375 a_n8300_8799.n192 a_n8300_8799.t129 464.166
R16376 a_n8300_8799.n180 a_n8300_8799.t79 464.166
R16377 a_n8300_8799.n193 a_n8300_8799.t80 464.166
R16378 a_n8300_8799.n194 a_n8300_8799.t125 464.166
R16379 a_n8300_8799.n195 a_n8300_8799.t46 464.166
R16380 a_n8300_8799.n196 a_n8300_8799.t76 464.166
R16381 a_n8300_8799.n179 a_n8300_8799.t100 464.166
R16382 a_n8300_8799.n197 a_n8300_8799.t151 464.166
R16383 a_n8300_8799.n204 a_n8300_8799.t70 464.166
R16384 a_n8300_8799.n205 a_n8300_8799.t91 464.166
R16385 a_n8300_8799.n206 a_n8300_8799.t48 464.166
R16386 a_n8300_8799.n207 a_n8300_8799.t109 464.166
R16387 a_n8300_8799.n202 a_n8300_8799.t86 464.166
R16388 a_n8300_8799.n208 a_n8300_8799.t130 464.166
R16389 a_n8300_8799.n209 a_n8300_8799.t77 464.166
R16390 a_n8300_8799.n210 a_n8300_8799.t138 464.166
R16391 a_n8300_8799.n211 a_n8300_8799.t53 464.166
R16392 a_n8300_8799.n201 a_n8300_8799.t37 464.166
R16393 a_n8300_8799.n212 a_n8300_8799.t94 464.166
R16394 a_n8300_8799.n200 a_n8300_8799.t141 464.166
R16395 a_n8300_8799.n213 a_n8300_8799.t113 464.166
R16396 a_n8300_8799.n214 a_n8300_8799.t147 464.166
R16397 a_n8300_8799.n215 a_n8300_8799.t87 464.166
R16398 a_n8300_8799.n216 a_n8300_8799.t42 464.166
R16399 a_n8300_8799.n199 a_n8300_8799.t104 464.166
R16400 a_n8300_8799.n217 a_n8300_8799.t57 464.166
R16401 a_n8300_8799.n41 a_n8300_8799.n70 71.7212
R16402 a_n8300_8799.n70 a_n8300_8799.n224 17.8606
R16403 a_n8300_8799.n69 a_n8300_8799.n41 76.9909
R16404 a_n8300_8799.n227 a_n8300_8799.n69 7.32118
R16405 a_n8300_8799.n68 a_n8300_8799.n40 78.3454
R16406 a_n8300_8799.n40 a_n8300_8799.n67 72.8951
R16407 a_n8300_8799.n66 a_n8300_8799.n42 70.1674
R16408 a_n8300_8799.n230 a_n8300_8799.n66 20.9683
R16409 a_n8300_8799.n42 a_n8300_8799.n65 72.3034
R16410 a_n8300_8799.n65 a_n8300_8799.n222 16.6962
R16411 a_n8300_8799.n64 a_n8300_8799.n43 77.6622
R16412 a_n8300_8799.n231 a_n8300_8799.n64 5.97853
R16413 a_n8300_8799.n63 a_n8300_8799.n43 77.6622
R16414 a_n8300_8799.n44 a_n8300_8799.n62 72.3034
R16415 a_n8300_8799.n61 a_n8300_8799.n44 70.1674
R16416 a_n8300_8799.n234 a_n8300_8799.n61 20.9683
R16417 a_n8300_8799.n46 a_n8300_8799.n60 72.8951
R16418 a_n8300_8799.n60 a_n8300_8799.n220 15.5127
R16419 a_n8300_8799.n59 a_n8300_8799.n46 78.3454
R16420 a_n8300_8799.n235 a_n8300_8799.n59 4.61226
R16421 a_n8300_8799.n58 a_n8300_8799.n45 76.9909
R16422 a_n8300_8799.n45 a_n8300_8799.n57 71.7212
R16423 a_n8300_8799.n237 a_n8300_8799.n56 20.9683
R16424 a_n8300_8799.n47 a_n8300_8799.n56 70.1674
R16425 a_n8300_8799.n33 a_n8300_8799.n85 71.7212
R16426 a_n8300_8799.n85 a_n8300_8799.n243 17.8606
R16427 a_n8300_8799.n84 a_n8300_8799.n33 76.9909
R16428 a_n8300_8799.n246 a_n8300_8799.n84 7.32118
R16429 a_n8300_8799.n83 a_n8300_8799.n32 78.3454
R16430 a_n8300_8799.n32 a_n8300_8799.n82 72.8951
R16431 a_n8300_8799.n81 a_n8300_8799.n34 70.1674
R16432 a_n8300_8799.n249 a_n8300_8799.n81 20.9683
R16433 a_n8300_8799.n34 a_n8300_8799.n80 72.3034
R16434 a_n8300_8799.n80 a_n8300_8799.n241 16.6962
R16435 a_n8300_8799.n79 a_n8300_8799.n35 77.6622
R16436 a_n8300_8799.n250 a_n8300_8799.n79 5.97853
R16437 a_n8300_8799.n78 a_n8300_8799.n35 77.6622
R16438 a_n8300_8799.n36 a_n8300_8799.n77 72.3034
R16439 a_n8300_8799.n76 a_n8300_8799.n36 70.1674
R16440 a_n8300_8799.n253 a_n8300_8799.n76 20.9683
R16441 a_n8300_8799.n38 a_n8300_8799.n75 72.8951
R16442 a_n8300_8799.n75 a_n8300_8799.n239 15.5127
R16443 a_n8300_8799.n74 a_n8300_8799.n38 78.3454
R16444 a_n8300_8799.n254 a_n8300_8799.n74 4.61226
R16445 a_n8300_8799.n73 a_n8300_8799.n37 76.9909
R16446 a_n8300_8799.n37 a_n8300_8799.n72 71.7212
R16447 a_n8300_8799.n256 a_n8300_8799.n71 20.9683
R16448 a_n8300_8799.n39 a_n8300_8799.n71 70.1674
R16449 a_n8300_8799.n25 a_n8300_8799.n100 71.7212
R16450 a_n8300_8799.n100 a_n8300_8799.n263 17.8606
R16451 a_n8300_8799.n99 a_n8300_8799.n25 76.9909
R16452 a_n8300_8799.n266 a_n8300_8799.n99 7.32118
R16453 a_n8300_8799.n98 a_n8300_8799.n24 78.3454
R16454 a_n8300_8799.n24 a_n8300_8799.n97 72.8951
R16455 a_n8300_8799.n96 a_n8300_8799.n26 70.1674
R16456 a_n8300_8799.n269 a_n8300_8799.n96 20.9683
R16457 a_n8300_8799.n26 a_n8300_8799.n95 72.3034
R16458 a_n8300_8799.n95 a_n8300_8799.n261 16.6962
R16459 a_n8300_8799.n94 a_n8300_8799.n27 77.6622
R16460 a_n8300_8799.n270 a_n8300_8799.n94 5.97853
R16461 a_n8300_8799.n93 a_n8300_8799.n27 77.6622
R16462 a_n8300_8799.n28 a_n8300_8799.n92 72.3034
R16463 a_n8300_8799.n91 a_n8300_8799.n28 70.1674
R16464 a_n8300_8799.n273 a_n8300_8799.n91 20.9683
R16465 a_n8300_8799.n30 a_n8300_8799.n90 72.8951
R16466 a_n8300_8799.n90 a_n8300_8799.n259 15.5127
R16467 a_n8300_8799.n89 a_n8300_8799.n30 78.3454
R16468 a_n8300_8799.n274 a_n8300_8799.n89 4.61226
R16469 a_n8300_8799.n88 a_n8300_8799.n29 76.9909
R16470 a_n8300_8799.n29 a_n8300_8799.n87 71.7212
R16471 a_n8300_8799.n276 a_n8300_8799.n86 20.9683
R16472 a_n8300_8799.n31 a_n8300_8799.n86 70.1674
R16473 a_n8300_8799.n17 a_n8300_8799.n115 70.1674
R16474 a_n8300_8799.n178 a_n8300_8799.n115 20.9683
R16475 a_n8300_8799.n114 a_n8300_8799.n17 71.7212
R16476 a_n8300_8799.n114 a_n8300_8799.n160 17.8606
R16477 a_n8300_8799.n16 a_n8300_8799.n113 76.9909
R16478 a_n8300_8799.n177 a_n8300_8799.n113 7.32118
R16479 a_n8300_8799.n112 a_n8300_8799.n16 78.3454
R16480 a_n8300_8799.n18 a_n8300_8799.n111 72.8951
R16481 a_n8300_8799.n110 a_n8300_8799.n18 70.1674
R16482 a_n8300_8799.n110 a_n8300_8799.n161 20.9683
R16483 a_n8300_8799.n19 a_n8300_8799.n109 72.3034
R16484 a_n8300_8799.n173 a_n8300_8799.n109 16.6962
R16485 a_n8300_8799.n108 a_n8300_8799.n19 77.6622
R16486 a_n8300_8799.n108 a_n8300_8799.n162 5.97853
R16487 a_n8300_8799.n20 a_n8300_8799.n107 77.6622
R16488 a_n8300_8799.n106 a_n8300_8799.n20 72.3034
R16489 a_n8300_8799.n21 a_n8300_8799.n105 70.1674
R16490 a_n8300_8799.n169 a_n8300_8799.n105 20.9683
R16491 a_n8300_8799.n104 a_n8300_8799.n21 72.8951
R16492 a_n8300_8799.n104 a_n8300_8799.n163 15.5127
R16493 a_n8300_8799.n22 a_n8300_8799.n103 78.3454
R16494 a_n8300_8799.n168 a_n8300_8799.n103 4.61226
R16495 a_n8300_8799.n102 a_n8300_8799.n22 76.9909
R16496 a_n8300_8799.n101 a_n8300_8799.n166 17.8606
R16497 a_n8300_8799.n101 a_n8300_8799.n23 71.7212
R16498 a_n8300_8799.n9 a_n8300_8799.n130 70.1674
R16499 a_n8300_8799.n197 a_n8300_8799.n130 20.9683
R16500 a_n8300_8799.n129 a_n8300_8799.n9 71.7212
R16501 a_n8300_8799.n129 a_n8300_8799.n179 17.8606
R16502 a_n8300_8799.n8 a_n8300_8799.n128 76.9909
R16503 a_n8300_8799.n196 a_n8300_8799.n128 7.32118
R16504 a_n8300_8799.n127 a_n8300_8799.n8 78.3454
R16505 a_n8300_8799.n10 a_n8300_8799.n126 72.8951
R16506 a_n8300_8799.n125 a_n8300_8799.n10 70.1674
R16507 a_n8300_8799.n125 a_n8300_8799.n180 20.9683
R16508 a_n8300_8799.n11 a_n8300_8799.n124 72.3034
R16509 a_n8300_8799.n192 a_n8300_8799.n124 16.6962
R16510 a_n8300_8799.n123 a_n8300_8799.n11 77.6622
R16511 a_n8300_8799.n123 a_n8300_8799.n181 5.97853
R16512 a_n8300_8799.n12 a_n8300_8799.n122 77.6622
R16513 a_n8300_8799.n121 a_n8300_8799.n12 72.3034
R16514 a_n8300_8799.n13 a_n8300_8799.n120 70.1674
R16515 a_n8300_8799.n188 a_n8300_8799.n120 20.9683
R16516 a_n8300_8799.n119 a_n8300_8799.n13 72.8951
R16517 a_n8300_8799.n119 a_n8300_8799.n182 15.5127
R16518 a_n8300_8799.n14 a_n8300_8799.n118 78.3454
R16519 a_n8300_8799.n187 a_n8300_8799.n118 4.61226
R16520 a_n8300_8799.n117 a_n8300_8799.n14 76.9909
R16521 a_n8300_8799.n116 a_n8300_8799.n185 17.8606
R16522 a_n8300_8799.n116 a_n8300_8799.n15 71.7212
R16523 a_n8300_8799.n1 a_n8300_8799.n145 70.1674
R16524 a_n8300_8799.n217 a_n8300_8799.n145 20.9683
R16525 a_n8300_8799.n144 a_n8300_8799.n1 71.7212
R16526 a_n8300_8799.n144 a_n8300_8799.n199 17.8606
R16527 a_n8300_8799.n0 a_n8300_8799.n143 76.9909
R16528 a_n8300_8799.n216 a_n8300_8799.n143 7.32118
R16529 a_n8300_8799.n142 a_n8300_8799.n0 78.3454
R16530 a_n8300_8799.n2 a_n8300_8799.n141 72.8951
R16531 a_n8300_8799.n140 a_n8300_8799.n2 70.1674
R16532 a_n8300_8799.n140 a_n8300_8799.n200 20.9683
R16533 a_n8300_8799.n3 a_n8300_8799.n139 72.3034
R16534 a_n8300_8799.n212 a_n8300_8799.n139 16.6962
R16535 a_n8300_8799.n138 a_n8300_8799.n3 77.6622
R16536 a_n8300_8799.n138 a_n8300_8799.n201 5.97853
R16537 a_n8300_8799.n4 a_n8300_8799.n137 77.6622
R16538 a_n8300_8799.n136 a_n8300_8799.n4 72.3034
R16539 a_n8300_8799.n5 a_n8300_8799.n135 70.1674
R16540 a_n8300_8799.n208 a_n8300_8799.n135 20.9683
R16541 a_n8300_8799.n134 a_n8300_8799.n5 72.8951
R16542 a_n8300_8799.n134 a_n8300_8799.n202 15.5127
R16543 a_n8300_8799.n6 a_n8300_8799.n133 78.3454
R16544 a_n8300_8799.n207 a_n8300_8799.n133 4.61226
R16545 a_n8300_8799.n132 a_n8300_8799.n6 76.9909
R16546 a_n8300_8799.n131 a_n8300_8799.n205 17.8606
R16547 a_n8300_8799.n131 a_n8300_8799.n7 71.7212
R16548 a_n8300_8799.n52 a_n8300_8799.n146 98.9633
R16549 a_n8300_8799.n55 a_n8300_8799.n283 98.9631
R16550 a_n8300_8799.n55 a_n8300_8799.n282 98.6055
R16551 a_n8300_8799.n54 a_n8300_8799.n281 98.6055
R16552 a_n8300_8799.n53 a_n8300_8799.n149 98.6055
R16553 a_n8300_8799.n53 a_n8300_8799.n148 98.6055
R16554 a_n8300_8799.n52 a_n8300_8799.n147 98.6055
R16555 a_n8300_8799.n284 a_n8300_8799.n55 98.6054
R16556 a_n8300_8799.n51 a_n8300_8799.n150 81.2902
R16557 a_n8300_8799.n49 a_n8300_8799.n156 81.2902
R16558 a_n8300_8799.n48 a_n8300_8799.n153 81.2902
R16559 a_n8300_8799.n50 a_n8300_8799.n158 80.9324
R16560 a_n8300_8799.n50 a_n8300_8799.n159 80.9324
R16561 a_n8300_8799.n51 a_n8300_8799.n152 80.9324
R16562 a_n8300_8799.n51 a_n8300_8799.n151 80.9324
R16563 a_n8300_8799.n49 a_n8300_8799.n157 80.9324
R16564 a_n8300_8799.n49 a_n8300_8799.n155 80.9324
R16565 a_n8300_8799.n48 a_n8300_8799.n154 80.9324
R16566 a_n8300_8799.n41 a_n8300_8799.n225 70.4033
R16567 a_n8300_8799.n33 a_n8300_8799.n244 70.4033
R16568 a_n8300_8799.n25 a_n8300_8799.n264 70.4033
R16569 a_n8300_8799.n164 a_n8300_8799.n23 70.4033
R16570 a_n8300_8799.n183 a_n8300_8799.n15 70.4033
R16571 a_n8300_8799.n203 a_n8300_8799.n7 70.4033
R16572 a_n8300_8799.n236 a_n8300_8799.n235 48.2005
R16573 a_n8300_8799.n61 a_n8300_8799.n233 20.9683
R16574 a_n8300_8799.n232 a_n8300_8799.n231 48.2005
R16575 a_n8300_8799.n66 a_n8300_8799.n229 20.9683
R16576 a_n8300_8799.n228 a_n8300_8799.n227 48.2005
R16577 a_n8300_8799.n255 a_n8300_8799.n254 48.2005
R16578 a_n8300_8799.n76 a_n8300_8799.n252 20.9683
R16579 a_n8300_8799.n251 a_n8300_8799.n250 48.2005
R16580 a_n8300_8799.n81 a_n8300_8799.n248 20.9683
R16581 a_n8300_8799.n247 a_n8300_8799.n246 48.2005
R16582 a_n8300_8799.n275 a_n8300_8799.n274 48.2005
R16583 a_n8300_8799.n91 a_n8300_8799.n272 20.9683
R16584 a_n8300_8799.n271 a_n8300_8799.n270 48.2005
R16585 a_n8300_8799.n96 a_n8300_8799.n268 20.9683
R16586 a_n8300_8799.n267 a_n8300_8799.n266 48.2005
R16587 a_n8300_8799.n168 a_n8300_8799.n167 48.2005
R16588 a_n8300_8799.n170 a_n8300_8799.n105 20.9683
R16589 a_n8300_8799.n172 a_n8300_8799.n162 48.2005
R16590 a_n8300_8799.n174 a_n8300_8799.n110 20.9683
R16591 a_n8300_8799.n177 a_n8300_8799.n176 48.2005
R16592 a_n8300_8799.t47 a_n8300_8799.n115 485.135
R16593 a_n8300_8799.n187 a_n8300_8799.n186 48.2005
R16594 a_n8300_8799.n189 a_n8300_8799.n120 20.9683
R16595 a_n8300_8799.n191 a_n8300_8799.n181 48.2005
R16596 a_n8300_8799.n193 a_n8300_8799.n125 20.9683
R16597 a_n8300_8799.n196 a_n8300_8799.n195 48.2005
R16598 a_n8300_8799.t59 a_n8300_8799.n130 485.135
R16599 a_n8300_8799.n207 a_n8300_8799.n206 48.2005
R16600 a_n8300_8799.n209 a_n8300_8799.n135 20.9683
R16601 a_n8300_8799.n211 a_n8300_8799.n201 48.2005
R16602 a_n8300_8799.n213 a_n8300_8799.n140 20.9683
R16603 a_n8300_8799.n216 a_n8300_8799.n215 48.2005
R16604 a_n8300_8799.t126 a_n8300_8799.n145 485.135
R16605 a_n8300_8799.n57 a_n8300_8799.n219 17.8606
R16606 a_n8300_8799.n226 a_n8300_8799.n70 25.894
R16607 a_n8300_8799.n72 a_n8300_8799.n238 17.8606
R16608 a_n8300_8799.n245 a_n8300_8799.n85 25.894
R16609 a_n8300_8799.n87 a_n8300_8799.n258 17.8606
R16610 a_n8300_8799.n265 a_n8300_8799.n100 25.894
R16611 a_n8300_8799.n178 a_n8300_8799.n114 25.894
R16612 a_n8300_8799.n197 a_n8300_8799.n129 25.894
R16613 a_n8300_8799.n217 a_n8300_8799.n144 25.894
R16614 a_n8300_8799.n68 a_n8300_8799.n223 43.3183
R16615 a_n8300_8799.n83 a_n8300_8799.n242 43.3183
R16616 a_n8300_8799.n98 a_n8300_8799.n262 43.3183
R16617 a_n8300_8799.n175 a_n8300_8799.n112 43.3183
R16618 a_n8300_8799.n194 a_n8300_8799.n127 43.3183
R16619 a_n8300_8799.n214 a_n8300_8799.n142 43.3183
R16620 a_n8300_8799.n62 a_n8300_8799.n221 16.6962
R16621 a_n8300_8799.n230 a_n8300_8799.n65 27.6507
R16622 a_n8300_8799.n77 a_n8300_8799.n240 16.6962
R16623 a_n8300_8799.n249 a_n8300_8799.n80 27.6507
R16624 a_n8300_8799.n92 a_n8300_8799.n260 16.6962
R16625 a_n8300_8799.n269 a_n8300_8799.n95 27.6507
R16626 a_n8300_8799.n171 a_n8300_8799.n106 16.6962
R16627 a_n8300_8799.n161 a_n8300_8799.n109 27.6507
R16628 a_n8300_8799.n190 a_n8300_8799.n121 16.6962
R16629 a_n8300_8799.n180 a_n8300_8799.n124 27.6507
R16630 a_n8300_8799.n210 a_n8300_8799.n136 16.6962
R16631 a_n8300_8799.n200 a_n8300_8799.n139 27.6507
R16632 a_n8300_8799.n63 a_n8300_8799.n221 41.7634
R16633 a_n8300_8799.n78 a_n8300_8799.n240 41.7634
R16634 a_n8300_8799.n93 a_n8300_8799.n260 41.7634
R16635 a_n8300_8799.n107 a_n8300_8799.n171 41.7634
R16636 a_n8300_8799.n122 a_n8300_8799.n190 41.7634
R16637 a_n8300_8799.n137 a_n8300_8799.n210 41.7634
R16638 a_n8300_8799.n234 a_n8300_8799.n60 29.3885
R16639 a_n8300_8799.n67 a_n8300_8799.n223 15.5127
R16640 a_n8300_8799.n253 a_n8300_8799.n75 29.3885
R16641 a_n8300_8799.n82 a_n8300_8799.n242 15.5127
R16642 a_n8300_8799.n273 a_n8300_8799.n90 29.3885
R16643 a_n8300_8799.n97 a_n8300_8799.n262 15.5127
R16644 a_n8300_8799.n169 a_n8300_8799.n104 29.3885
R16645 a_n8300_8799.n175 a_n8300_8799.n111 15.5127
R16646 a_n8300_8799.n188 a_n8300_8799.n119 29.3885
R16647 a_n8300_8799.n194 a_n8300_8799.n126 15.5127
R16648 a_n8300_8799.n208 a_n8300_8799.n134 29.3885
R16649 a_n8300_8799.n214 a_n8300_8799.n141 15.5127
R16650 a_n8300_8799.n58 a_n8300_8799.n219 40.1848
R16651 a_n8300_8799.n73 a_n8300_8799.n238 40.1848
R16652 a_n8300_8799.n88 a_n8300_8799.n258 40.1848
R16653 a_n8300_8799.n166 a_n8300_8799.n102 40.1848
R16654 a_n8300_8799.n185 a_n8300_8799.n117 40.1848
R16655 a_n8300_8799.n205 a_n8300_8799.n132 40.1848
R16656 a_n8300_8799.n50 a_n8300_8799.n49 31.9767
R16657 a_n8300_8799.n54 a_n8300_8799.n280 31.5713
R16658 a_n8300_8799.n226 a_n8300_8799.n225 20.9576
R16659 a_n8300_8799.n245 a_n8300_8799.n244 20.9576
R16660 a_n8300_8799.n265 a_n8300_8799.n264 20.9576
R16661 a_n8300_8799.n165 a_n8300_8799.n164 20.9576
R16662 a_n8300_8799.n184 a_n8300_8799.n183 20.9576
R16663 a_n8300_8799.n204 a_n8300_8799.n203 20.9576
R16664 a_n8300_8799.n280 a_n8300_8799.n53 19.0249
R16665 a_n8300_8799.n58 a_n8300_8799.n236 7.32118
R16666 a_n8300_8799.n69 a_n8300_8799.n224 40.1848
R16667 a_n8300_8799.n73 a_n8300_8799.n255 7.32118
R16668 a_n8300_8799.n84 a_n8300_8799.n243 40.1848
R16669 a_n8300_8799.n88 a_n8300_8799.n275 7.32118
R16670 a_n8300_8799.n99 a_n8300_8799.n263 40.1848
R16671 a_n8300_8799.n167 a_n8300_8799.n102 7.32118
R16672 a_n8300_8799.n160 a_n8300_8799.n113 40.1848
R16673 a_n8300_8799.n186 a_n8300_8799.n117 7.32118
R16674 a_n8300_8799.n179 a_n8300_8799.n128 40.1848
R16675 a_n8300_8799.n206 a_n8300_8799.n132 7.32118
R16676 a_n8300_8799.n199 a_n8300_8799.n143 40.1848
R16677 a_n8300_8799.n229 a_n8300_8799.n67 29.3885
R16678 a_n8300_8799.n248 a_n8300_8799.n82 29.3885
R16679 a_n8300_8799.n268 a_n8300_8799.n97 29.3885
R16680 a_n8300_8799.n111 a_n8300_8799.n174 29.3885
R16681 a_n8300_8799.n126 a_n8300_8799.n193 29.3885
R16682 a_n8300_8799.n141 a_n8300_8799.n213 29.3885
R16683 a_n8300_8799.n63 a_n8300_8799.n232 5.97853
R16684 a_n8300_8799.n64 a_n8300_8799.n222 41.7634
R16685 a_n8300_8799.n78 a_n8300_8799.n251 5.97853
R16686 a_n8300_8799.n79 a_n8300_8799.n241 41.7634
R16687 a_n8300_8799.n93 a_n8300_8799.n271 5.97853
R16688 a_n8300_8799.n94 a_n8300_8799.n261 41.7634
R16689 a_n8300_8799.n172 a_n8300_8799.n107 5.97853
R16690 a_n8300_8799.n173 a_n8300_8799.n108 41.7634
R16691 a_n8300_8799.n191 a_n8300_8799.n122 5.97853
R16692 a_n8300_8799.n192 a_n8300_8799.n123 41.7634
R16693 a_n8300_8799.n211 a_n8300_8799.n137 5.97853
R16694 a_n8300_8799.n212 a_n8300_8799.n138 41.7634
R16695 a_n8300_8799.n279 a_n8300_8799.n51 12.3339
R16696 a_n8300_8799.n280 a_n8300_8799.n279 11.4887
R16697 a_n8300_8799.n233 a_n8300_8799.n62 27.6507
R16698 a_n8300_8799.n252 a_n8300_8799.n77 27.6507
R16699 a_n8300_8799.n272 a_n8300_8799.n92 27.6507
R16700 a_n8300_8799.n170 a_n8300_8799.n106 27.6507
R16701 a_n8300_8799.n189 a_n8300_8799.n121 27.6507
R16702 a_n8300_8799.n209 a_n8300_8799.n136 27.6507
R16703 a_n8300_8799.n59 a_n8300_8799.n220 43.3183
R16704 a_n8300_8799.n68 a_n8300_8799.n228 4.61226
R16705 a_n8300_8799.n74 a_n8300_8799.n239 43.3183
R16706 a_n8300_8799.n83 a_n8300_8799.n247 4.61226
R16707 a_n8300_8799.n89 a_n8300_8799.n259 43.3183
R16708 a_n8300_8799.n98 a_n8300_8799.n267 4.61226
R16709 a_n8300_8799.n163 a_n8300_8799.n103 43.3183
R16710 a_n8300_8799.n176 a_n8300_8799.n112 4.61226
R16711 a_n8300_8799.n182 a_n8300_8799.n118 43.3183
R16712 a_n8300_8799.n195 a_n8300_8799.n127 4.61226
R16713 a_n8300_8799.n202 a_n8300_8799.n133 43.3183
R16714 a_n8300_8799.n215 a_n8300_8799.n142 4.61226
R16715 a_n8300_8799.n257 a_n8300_8799.n47 9.04406
R16716 a_n8300_8799.n198 a_n8300_8799.n17 9.04406
R16717 a_n8300_8799.n237 a_n8300_8799.n57 25.894
R16718 a_n8300_8799.n256 a_n8300_8799.n72 25.894
R16719 a_n8300_8799.n276 a_n8300_8799.n87 25.894
R16720 a_n8300_8799.n101 a_n8300_8799.n165 25.894
R16721 a_n8300_8799.n116 a_n8300_8799.n184 25.894
R16722 a_n8300_8799.n131 a_n8300_8799.n204 25.894
R16723 a_n8300_8799.n278 a_n8300_8799.n218 6.94254
R16724 a_n8300_8799.n278 a_n8300_8799.n277 6.64832
R16725 a_n8300_8799.n257 a_n8300_8799.n39 4.93611
R16726 a_n8300_8799.n277 a_n8300_8799.n31 4.93611
R16727 a_n8300_8799.n198 a_n8300_8799.n9 4.93611
R16728 a_n8300_8799.n218 a_n8300_8799.n1 4.93611
R16729 a_n8300_8799.n277 a_n8300_8799.n257 4.10845
R16730 a_n8300_8799.n218 a_n8300_8799.n198 4.10845
R16731 a_n8300_8799.n283 a_n8300_8799.t28 3.61217
R16732 a_n8300_8799.n283 a_n8300_8799.t15 3.61217
R16733 a_n8300_8799.n282 a_n8300_8799.t22 3.61217
R16734 a_n8300_8799.n282 a_n8300_8799.t26 3.61217
R16735 a_n8300_8799.n281 a_n8300_8799.t24 3.61217
R16736 a_n8300_8799.n281 a_n8300_8799.t20 3.61217
R16737 a_n8300_8799.n149 a_n8300_8799.t19 3.61217
R16738 a_n8300_8799.n149 a_n8300_8799.t14 3.61217
R16739 a_n8300_8799.n148 a_n8300_8799.t27 3.61217
R16740 a_n8300_8799.n148 a_n8300_8799.t25 3.61217
R16741 a_n8300_8799.n147 a_n8300_8799.t11 3.61217
R16742 a_n8300_8799.n147 a_n8300_8799.t21 3.61217
R16743 a_n8300_8799.n146 a_n8300_8799.t23 3.61217
R16744 a_n8300_8799.n146 a_n8300_8799.t13 3.61217
R16745 a_n8300_8799.t5 a_n8300_8799.n284 3.61217
R16746 a_n8300_8799.n284 a_n8300_8799.t12 3.61217
R16747 a_n8300_8799.n279 a_n8300_8799.n278 3.4105
R16748 a_n8300_8799.n158 a_n8300_8799.t34 2.82907
R16749 a_n8300_8799.n158 a_n8300_8799.t7 2.82907
R16750 a_n8300_8799.n159 a_n8300_8799.t29 2.82907
R16751 a_n8300_8799.n159 a_n8300_8799.t6 2.82907
R16752 a_n8300_8799.n152 a_n8300_8799.t2 2.82907
R16753 a_n8300_8799.n152 a_n8300_8799.t3 2.82907
R16754 a_n8300_8799.n151 a_n8300_8799.t35 2.82907
R16755 a_n8300_8799.n151 a_n8300_8799.t33 2.82907
R16756 a_n8300_8799.n150 a_n8300_8799.t18 2.82907
R16757 a_n8300_8799.n150 a_n8300_8799.t31 2.82907
R16758 a_n8300_8799.n156 a_n8300_8799.t30 2.82907
R16759 a_n8300_8799.n156 a_n8300_8799.t0 2.82907
R16760 a_n8300_8799.n157 a_n8300_8799.t4 2.82907
R16761 a_n8300_8799.n157 a_n8300_8799.t17 2.82907
R16762 a_n8300_8799.n155 a_n8300_8799.t1 2.82907
R16763 a_n8300_8799.n155 a_n8300_8799.t10 2.82907
R16764 a_n8300_8799.n154 a_n8300_8799.t32 2.82907
R16765 a_n8300_8799.n154 a_n8300_8799.t8 2.82907
R16766 a_n8300_8799.n153 a_n8300_8799.t9 2.82907
R16767 a_n8300_8799.n153 a_n8300_8799.t16 2.82907
R16768 a_n8300_8799.n41 a_n8300_8799.n40 1.13686
R16769 a_n8300_8799.n33 a_n8300_8799.n32 1.13686
R16770 a_n8300_8799.n25 a_n8300_8799.n24 1.13686
R16771 a_n8300_8799.n17 a_n8300_8799.n16 1.13686
R16772 a_n8300_8799.n9 a_n8300_8799.n8 1.13686
R16773 a_n8300_8799.n1 a_n8300_8799.n0 1.13686
R16774 a_n8300_8799.n51 a_n8300_8799.n50 1.07378
R16775 a_n8300_8799.n46 a_n8300_8799.n45 0.758076
R16776 a_n8300_8799.n46 a_n8300_8799.n44 0.758076
R16777 a_n8300_8799.n44 a_n8300_8799.n43 0.758076
R16778 a_n8300_8799.n43 a_n8300_8799.n42 0.758076
R16779 a_n8300_8799.n40 a_n8300_8799.n42 0.758076
R16780 a_n8300_8799.n38 a_n8300_8799.n37 0.758076
R16781 a_n8300_8799.n38 a_n8300_8799.n36 0.758076
R16782 a_n8300_8799.n36 a_n8300_8799.n35 0.758076
R16783 a_n8300_8799.n35 a_n8300_8799.n34 0.758076
R16784 a_n8300_8799.n32 a_n8300_8799.n34 0.758076
R16785 a_n8300_8799.n30 a_n8300_8799.n29 0.758076
R16786 a_n8300_8799.n30 a_n8300_8799.n28 0.758076
R16787 a_n8300_8799.n28 a_n8300_8799.n27 0.758076
R16788 a_n8300_8799.n27 a_n8300_8799.n26 0.758076
R16789 a_n8300_8799.n24 a_n8300_8799.n26 0.758076
R16790 a_n8300_8799.n21 a_n8300_8799.n22 0.758076
R16791 a_n8300_8799.n20 a_n8300_8799.n21 0.758076
R16792 a_n8300_8799.n19 a_n8300_8799.n20 0.758076
R16793 a_n8300_8799.n18 a_n8300_8799.n19 0.758076
R16794 a_n8300_8799.n16 a_n8300_8799.n18 0.758076
R16795 a_n8300_8799.n13 a_n8300_8799.n14 0.758076
R16796 a_n8300_8799.n12 a_n8300_8799.n13 0.758076
R16797 a_n8300_8799.n11 a_n8300_8799.n12 0.758076
R16798 a_n8300_8799.n10 a_n8300_8799.n11 0.758076
R16799 a_n8300_8799.n8 a_n8300_8799.n10 0.758076
R16800 a_n8300_8799.n5 a_n8300_8799.n6 0.758076
R16801 a_n8300_8799.n4 a_n8300_8799.n5 0.758076
R16802 a_n8300_8799.n3 a_n8300_8799.n4 0.758076
R16803 a_n8300_8799.n2 a_n8300_8799.n3 0.758076
R16804 a_n8300_8799.n0 a_n8300_8799.n2 0.758076
R16805 a_n8300_8799.n55 a_n8300_8799.n54 0.716017
R16806 a_n8300_8799.n53 a_n8300_8799.n52 0.716017
R16807 a_n8300_8799.n49 a_n8300_8799.n48 0.716017
R16808 a_n8300_8799.n6 a_n8300_8799.n7 0.568682
R16809 a_n8300_8799.n14 a_n8300_8799.n15 0.568682
R16810 a_n8300_8799.n22 a_n8300_8799.n23 0.568682
R16811 a_n8300_8799.n29 a_n8300_8799.n31 0.568682
R16812 a_n8300_8799.n37 a_n8300_8799.n39 0.568682
R16813 a_n8300_8799.n45 a_n8300_8799.n47 0.568682
R16814 vdd.n327 vdd.n291 756.745
R16815 vdd.n268 vdd.n232 756.745
R16816 vdd.n225 vdd.n189 756.745
R16817 vdd.n166 vdd.n130 756.745
R16818 vdd.n124 vdd.n88 756.745
R16819 vdd.n65 vdd.n29 756.745
R16820 vdd.n2108 vdd.n2072 756.745
R16821 vdd.n2167 vdd.n2131 756.745
R16822 vdd.n2006 vdd.n1970 756.745
R16823 vdd.n2065 vdd.n2029 756.745
R16824 vdd.n1905 vdd.n1869 756.745
R16825 vdd.n1964 vdd.n1928 756.745
R16826 vdd.n1253 vdd.t30 640.208
R16827 vdd.n981 vdd.t72 640.208
R16828 vdd.n1273 vdd.t45 640.208
R16829 vdd.n972 vdd.t96 640.208
R16830 vdd.n872 vdd.t52 640.208
R16831 vdd.n2704 vdd.t87 640.208
R16832 vdd.n832 vdd.t99 640.208
R16833 vdd.n2701 vdd.t76 640.208
R16834 vdd.n799 vdd.t26 640.208
R16835 vdd.n1043 vdd.t83 640.208
R16836 vdd.n1679 vdd.t62 592.009
R16837 vdd.n1717 vdd.t80 592.009
R16838 vdd.n1613 vdd.t93 592.009
R16839 vdd.n2269 vdd.t38 592.009
R16840 vdd.n1190 vdd.t69 592.009
R16841 vdd.n1150 vdd.t90 592.009
R16842 vdd.n426 vdd.t59 592.009
R16843 vdd.n440 vdd.t48 592.009
R16844 vdd.n452 vdd.t66 592.009
R16845 vdd.n768 vdd.t42 592.009
R16846 vdd.n3276 vdd.t56 592.009
R16847 vdd.n688 vdd.t34 592.009
R16848 vdd.n328 vdd.n327 585
R16849 vdd.n326 vdd.n293 585
R16850 vdd.n325 vdd.n324 585
R16851 vdd.n296 vdd.n294 585
R16852 vdd.n319 vdd.n318 585
R16853 vdd.n317 vdd.n316 585
R16854 vdd.n300 vdd.n299 585
R16855 vdd.n311 vdd.n310 585
R16856 vdd.n309 vdd.n308 585
R16857 vdd.n304 vdd.n303 585
R16858 vdd.n269 vdd.n268 585
R16859 vdd.n267 vdd.n234 585
R16860 vdd.n266 vdd.n265 585
R16861 vdd.n237 vdd.n235 585
R16862 vdd.n260 vdd.n259 585
R16863 vdd.n258 vdd.n257 585
R16864 vdd.n241 vdd.n240 585
R16865 vdd.n252 vdd.n251 585
R16866 vdd.n250 vdd.n249 585
R16867 vdd.n245 vdd.n244 585
R16868 vdd.n226 vdd.n225 585
R16869 vdd.n224 vdd.n191 585
R16870 vdd.n223 vdd.n222 585
R16871 vdd.n194 vdd.n192 585
R16872 vdd.n217 vdd.n216 585
R16873 vdd.n215 vdd.n214 585
R16874 vdd.n198 vdd.n197 585
R16875 vdd.n209 vdd.n208 585
R16876 vdd.n207 vdd.n206 585
R16877 vdd.n202 vdd.n201 585
R16878 vdd.n167 vdd.n166 585
R16879 vdd.n165 vdd.n132 585
R16880 vdd.n164 vdd.n163 585
R16881 vdd.n135 vdd.n133 585
R16882 vdd.n158 vdd.n157 585
R16883 vdd.n156 vdd.n155 585
R16884 vdd.n139 vdd.n138 585
R16885 vdd.n150 vdd.n149 585
R16886 vdd.n148 vdd.n147 585
R16887 vdd.n143 vdd.n142 585
R16888 vdd.n125 vdd.n124 585
R16889 vdd.n123 vdd.n90 585
R16890 vdd.n122 vdd.n121 585
R16891 vdd.n93 vdd.n91 585
R16892 vdd.n116 vdd.n115 585
R16893 vdd.n114 vdd.n113 585
R16894 vdd.n97 vdd.n96 585
R16895 vdd.n108 vdd.n107 585
R16896 vdd.n106 vdd.n105 585
R16897 vdd.n101 vdd.n100 585
R16898 vdd.n66 vdd.n65 585
R16899 vdd.n64 vdd.n31 585
R16900 vdd.n63 vdd.n62 585
R16901 vdd.n34 vdd.n32 585
R16902 vdd.n57 vdd.n56 585
R16903 vdd.n55 vdd.n54 585
R16904 vdd.n38 vdd.n37 585
R16905 vdd.n49 vdd.n48 585
R16906 vdd.n47 vdd.n46 585
R16907 vdd.n42 vdd.n41 585
R16908 vdd.n2109 vdd.n2108 585
R16909 vdd.n2107 vdd.n2074 585
R16910 vdd.n2106 vdd.n2105 585
R16911 vdd.n2077 vdd.n2075 585
R16912 vdd.n2100 vdd.n2099 585
R16913 vdd.n2098 vdd.n2097 585
R16914 vdd.n2081 vdd.n2080 585
R16915 vdd.n2092 vdd.n2091 585
R16916 vdd.n2090 vdd.n2089 585
R16917 vdd.n2085 vdd.n2084 585
R16918 vdd.n2168 vdd.n2167 585
R16919 vdd.n2166 vdd.n2133 585
R16920 vdd.n2165 vdd.n2164 585
R16921 vdd.n2136 vdd.n2134 585
R16922 vdd.n2159 vdd.n2158 585
R16923 vdd.n2157 vdd.n2156 585
R16924 vdd.n2140 vdd.n2139 585
R16925 vdd.n2151 vdd.n2150 585
R16926 vdd.n2149 vdd.n2148 585
R16927 vdd.n2144 vdd.n2143 585
R16928 vdd.n2007 vdd.n2006 585
R16929 vdd.n2005 vdd.n1972 585
R16930 vdd.n2004 vdd.n2003 585
R16931 vdd.n1975 vdd.n1973 585
R16932 vdd.n1998 vdd.n1997 585
R16933 vdd.n1996 vdd.n1995 585
R16934 vdd.n1979 vdd.n1978 585
R16935 vdd.n1990 vdd.n1989 585
R16936 vdd.n1988 vdd.n1987 585
R16937 vdd.n1983 vdd.n1982 585
R16938 vdd.n2066 vdd.n2065 585
R16939 vdd.n2064 vdd.n2031 585
R16940 vdd.n2063 vdd.n2062 585
R16941 vdd.n2034 vdd.n2032 585
R16942 vdd.n2057 vdd.n2056 585
R16943 vdd.n2055 vdd.n2054 585
R16944 vdd.n2038 vdd.n2037 585
R16945 vdd.n2049 vdd.n2048 585
R16946 vdd.n2047 vdd.n2046 585
R16947 vdd.n2042 vdd.n2041 585
R16948 vdd.n1906 vdd.n1905 585
R16949 vdd.n1904 vdd.n1871 585
R16950 vdd.n1903 vdd.n1902 585
R16951 vdd.n1874 vdd.n1872 585
R16952 vdd.n1897 vdd.n1896 585
R16953 vdd.n1895 vdd.n1894 585
R16954 vdd.n1878 vdd.n1877 585
R16955 vdd.n1889 vdd.n1888 585
R16956 vdd.n1887 vdd.n1886 585
R16957 vdd.n1882 vdd.n1881 585
R16958 vdd.n1965 vdd.n1964 585
R16959 vdd.n1963 vdd.n1930 585
R16960 vdd.n1962 vdd.n1961 585
R16961 vdd.n1933 vdd.n1931 585
R16962 vdd.n1956 vdd.n1955 585
R16963 vdd.n1954 vdd.n1953 585
R16964 vdd.n1937 vdd.n1936 585
R16965 vdd.n1948 vdd.n1947 585
R16966 vdd.n1946 vdd.n1945 585
R16967 vdd.n1941 vdd.n1940 585
R16968 vdd.n3448 vdd.n392 509.269
R16969 vdd.n3444 vdd.n393 509.269
R16970 vdd.n3316 vdd.n685 509.269
R16971 vdd.n3313 vdd.n684 509.269
R16972 vdd.n2264 vdd.n1437 509.269
R16973 vdd.n2267 vdd.n2266 509.269
R16974 vdd.n1586 vdd.n1550 509.269
R16975 vdd.n1782 vdd.n1551 509.269
R16976 vdd.n305 vdd.t161 329.043
R16977 vdd.n246 vdd.t246 329.043
R16978 vdd.n203 vdd.t297 329.043
R16979 vdd.n144 vdd.t230 329.043
R16980 vdd.n102 vdd.t198 329.043
R16981 vdd.n43 vdd.t187 329.043
R16982 vdd.n2086 vdd.t288 329.043
R16983 vdd.n2145 vdd.t222 329.043
R16984 vdd.n1984 vdd.t276 329.043
R16985 vdd.n2043 vdd.t199 329.043
R16986 vdd.n1883 vdd.t189 329.043
R16987 vdd.n1942 vdd.t197 329.043
R16988 vdd.n1679 vdd.t65 319.788
R16989 vdd.n1717 vdd.t82 319.788
R16990 vdd.n1613 vdd.t95 319.788
R16991 vdd.n2269 vdd.t40 319.788
R16992 vdd.n1190 vdd.t70 319.788
R16993 vdd.n1150 vdd.t91 319.788
R16994 vdd.n426 vdd.t60 319.788
R16995 vdd.n440 vdd.t50 319.788
R16996 vdd.n452 vdd.t67 319.788
R16997 vdd.n768 vdd.t44 319.788
R16998 vdd.n3276 vdd.t58 319.788
R16999 vdd.n688 vdd.t37 319.788
R17000 vdd.n1680 vdd.t64 303.69
R17001 vdd.n1718 vdd.t81 303.69
R17002 vdd.n1614 vdd.t94 303.69
R17003 vdd.n2270 vdd.t41 303.69
R17004 vdd.n1191 vdd.t71 303.69
R17005 vdd.n1151 vdd.t92 303.69
R17006 vdd.n427 vdd.t61 303.69
R17007 vdd.n441 vdd.t51 303.69
R17008 vdd.n453 vdd.t68 303.69
R17009 vdd.n769 vdd.t43 303.69
R17010 vdd.n3277 vdd.t57 303.69
R17011 vdd.n689 vdd.t36 303.69
R17012 vdd.n2936 vdd.n927 291.221
R17013 vdd.n3150 vdd.n809 291.221
R17014 vdd.n3087 vdd.n806 291.221
R17015 vdd.n2868 vdd.n2867 291.221
R17016 vdd.n2664 vdd.n969 291.221
R17017 vdd.n2595 vdd.n2594 291.221
R17018 vdd.n1309 vdd.n1308 291.221
R17019 vdd.n2415 vdd.n1075 291.221
R17020 vdd.n3066 vdd.n807 291.221
R17021 vdd.n3153 vdd.n3152 291.221
R17022 vdd.n2772 vdd.n2698 291.221
R17023 vdd.n2940 vdd.n931 291.221
R17024 vdd.n2592 vdd.n979 291.221
R17025 vdd.n977 vdd.n951 291.221
R17026 vdd.n1387 vdd.n1116 291.221
R17027 vdd.n2419 vdd.n1080 291.221
R17028 vdd.n3068 vdd.n807 185
R17029 vdd.n3151 vdd.n807 185
R17030 vdd.n3070 vdd.n3069 185
R17031 vdd.n3069 vdd.n805 185
R17032 vdd.n3071 vdd.n839 185
R17033 vdd.n3081 vdd.n839 185
R17034 vdd.n3072 vdd.n848 185
R17035 vdd.n848 vdd.n846 185
R17036 vdd.n3074 vdd.n3073 185
R17037 vdd.n3075 vdd.n3074 185
R17038 vdd.n3027 vdd.n847 185
R17039 vdd.n847 vdd.n843 185
R17040 vdd.n3026 vdd.n3025 185
R17041 vdd.n3025 vdd.n3024 185
R17042 vdd.n850 vdd.n849 185
R17043 vdd.n851 vdd.n850 185
R17044 vdd.n3017 vdd.n3016 185
R17045 vdd.n3018 vdd.n3017 185
R17046 vdd.n3015 vdd.n860 185
R17047 vdd.n860 vdd.n857 185
R17048 vdd.n3014 vdd.n3013 185
R17049 vdd.n3013 vdd.n3012 185
R17050 vdd.n862 vdd.n861 185
R17051 vdd.n870 vdd.n862 185
R17052 vdd.n3005 vdd.n3004 185
R17053 vdd.n3006 vdd.n3005 185
R17054 vdd.n3002 vdd.n871 185
R17055 vdd.n878 vdd.n871 185
R17056 vdd.n3001 vdd.n3000 185
R17057 vdd.n3000 vdd.n2999 185
R17058 vdd.n874 vdd.n873 185
R17059 vdd.n875 vdd.n874 185
R17060 vdd.n2992 vdd.n2991 185
R17061 vdd.n2993 vdd.n2992 185
R17062 vdd.n2990 vdd.n885 185
R17063 vdd.n885 vdd.n882 185
R17064 vdd.n2989 vdd.n2988 185
R17065 vdd.n2988 vdd.n2987 185
R17066 vdd.n887 vdd.n886 185
R17067 vdd.n895 vdd.n887 185
R17068 vdd.n2980 vdd.n2979 185
R17069 vdd.n2981 vdd.n2980 185
R17070 vdd.n2978 vdd.n896 185
R17071 vdd.n901 vdd.n896 185
R17072 vdd.n2977 vdd.n2976 185
R17073 vdd.n2976 vdd.n2975 185
R17074 vdd.n898 vdd.n897 185
R17075 vdd.n2847 vdd.n898 185
R17076 vdd.n2968 vdd.n2967 185
R17077 vdd.n2969 vdd.n2968 185
R17078 vdd.n2966 vdd.n908 185
R17079 vdd.n908 vdd.n905 185
R17080 vdd.n2965 vdd.n2964 185
R17081 vdd.n2964 vdd.n2963 185
R17082 vdd.n910 vdd.n909 185
R17083 vdd.n911 vdd.n910 185
R17084 vdd.n2956 vdd.n2955 185
R17085 vdd.n2957 vdd.n2956 185
R17086 vdd.n2954 vdd.n920 185
R17087 vdd.n920 vdd.n917 185
R17088 vdd.n2953 vdd.n2952 185
R17089 vdd.n2952 vdd.n2951 185
R17090 vdd.n922 vdd.n921 185
R17091 vdd.n2862 vdd.n922 185
R17092 vdd.n2944 vdd.n2943 185
R17093 vdd.n2945 vdd.n2944 185
R17094 vdd.n2942 vdd.n931 185
R17095 vdd.n931 vdd.n928 185
R17096 vdd.n2941 vdd.n2940 185
R17097 vdd.n933 vdd.n932 185
R17098 vdd.n2708 vdd.n2707 185
R17099 vdd.n2710 vdd.n2709 185
R17100 vdd.n2712 vdd.n2711 185
R17101 vdd.n2714 vdd.n2713 185
R17102 vdd.n2716 vdd.n2715 185
R17103 vdd.n2718 vdd.n2717 185
R17104 vdd.n2720 vdd.n2719 185
R17105 vdd.n2722 vdd.n2721 185
R17106 vdd.n2724 vdd.n2723 185
R17107 vdd.n2726 vdd.n2725 185
R17108 vdd.n2728 vdd.n2727 185
R17109 vdd.n2730 vdd.n2729 185
R17110 vdd.n2732 vdd.n2731 185
R17111 vdd.n2734 vdd.n2733 185
R17112 vdd.n2736 vdd.n2735 185
R17113 vdd.n2738 vdd.n2737 185
R17114 vdd.n2740 vdd.n2739 185
R17115 vdd.n2742 vdd.n2741 185
R17116 vdd.n2744 vdd.n2743 185
R17117 vdd.n2746 vdd.n2745 185
R17118 vdd.n2748 vdd.n2747 185
R17119 vdd.n2750 vdd.n2749 185
R17120 vdd.n2752 vdd.n2751 185
R17121 vdd.n2754 vdd.n2753 185
R17122 vdd.n2756 vdd.n2755 185
R17123 vdd.n2758 vdd.n2757 185
R17124 vdd.n2760 vdd.n2759 185
R17125 vdd.n2762 vdd.n2761 185
R17126 vdd.n2764 vdd.n2763 185
R17127 vdd.n2766 vdd.n2765 185
R17128 vdd.n2768 vdd.n2767 185
R17129 vdd.n2770 vdd.n2769 185
R17130 vdd.n2771 vdd.n2698 185
R17131 vdd.n2938 vdd.n2698 185
R17132 vdd.n3154 vdd.n3153 185
R17133 vdd.n3155 vdd.n798 185
R17134 vdd.n3157 vdd.n3156 185
R17135 vdd.n3159 vdd.n796 185
R17136 vdd.n3161 vdd.n3160 185
R17137 vdd.n3162 vdd.n795 185
R17138 vdd.n3164 vdd.n3163 185
R17139 vdd.n3166 vdd.n793 185
R17140 vdd.n3168 vdd.n3167 185
R17141 vdd.n3169 vdd.n792 185
R17142 vdd.n3171 vdd.n3170 185
R17143 vdd.n3173 vdd.n790 185
R17144 vdd.n3175 vdd.n3174 185
R17145 vdd.n3176 vdd.n789 185
R17146 vdd.n3178 vdd.n3177 185
R17147 vdd.n3180 vdd.n788 185
R17148 vdd.n3181 vdd.n786 185
R17149 vdd.n3184 vdd.n3183 185
R17150 vdd.n787 vdd.n785 185
R17151 vdd.n3040 vdd.n3039 185
R17152 vdd.n3042 vdd.n3041 185
R17153 vdd.n3044 vdd.n3036 185
R17154 vdd.n3046 vdd.n3045 185
R17155 vdd.n3047 vdd.n3035 185
R17156 vdd.n3049 vdd.n3048 185
R17157 vdd.n3051 vdd.n3033 185
R17158 vdd.n3053 vdd.n3052 185
R17159 vdd.n3054 vdd.n3032 185
R17160 vdd.n3056 vdd.n3055 185
R17161 vdd.n3058 vdd.n3030 185
R17162 vdd.n3060 vdd.n3059 185
R17163 vdd.n3061 vdd.n3029 185
R17164 vdd.n3063 vdd.n3062 185
R17165 vdd.n3065 vdd.n3028 185
R17166 vdd.n3067 vdd.n3066 185
R17167 vdd.n3066 vdd.n692 185
R17168 vdd.n3152 vdd.n802 185
R17169 vdd.n3152 vdd.n3151 185
R17170 vdd.n2775 vdd.n804 185
R17171 vdd.n805 vdd.n804 185
R17172 vdd.n2776 vdd.n838 185
R17173 vdd.n3081 vdd.n838 185
R17174 vdd.n2778 vdd.n2777 185
R17175 vdd.n2777 vdd.n846 185
R17176 vdd.n2779 vdd.n845 185
R17177 vdd.n3075 vdd.n845 185
R17178 vdd.n2781 vdd.n2780 185
R17179 vdd.n2780 vdd.n843 185
R17180 vdd.n2782 vdd.n853 185
R17181 vdd.n3024 vdd.n853 185
R17182 vdd.n2784 vdd.n2783 185
R17183 vdd.n2783 vdd.n851 185
R17184 vdd.n2785 vdd.n859 185
R17185 vdd.n3018 vdd.n859 185
R17186 vdd.n2787 vdd.n2786 185
R17187 vdd.n2786 vdd.n857 185
R17188 vdd.n2788 vdd.n864 185
R17189 vdd.n3012 vdd.n864 185
R17190 vdd.n2790 vdd.n2789 185
R17191 vdd.n2789 vdd.n870 185
R17192 vdd.n2791 vdd.n869 185
R17193 vdd.n3006 vdd.n869 185
R17194 vdd.n2793 vdd.n2792 185
R17195 vdd.n2792 vdd.n878 185
R17196 vdd.n2794 vdd.n877 185
R17197 vdd.n2999 vdd.n877 185
R17198 vdd.n2796 vdd.n2795 185
R17199 vdd.n2795 vdd.n875 185
R17200 vdd.n2797 vdd.n884 185
R17201 vdd.n2993 vdd.n884 185
R17202 vdd.n2799 vdd.n2798 185
R17203 vdd.n2798 vdd.n882 185
R17204 vdd.n2800 vdd.n889 185
R17205 vdd.n2987 vdd.n889 185
R17206 vdd.n2802 vdd.n2801 185
R17207 vdd.n2801 vdd.n895 185
R17208 vdd.n2803 vdd.n894 185
R17209 vdd.n2981 vdd.n894 185
R17210 vdd.n2805 vdd.n2804 185
R17211 vdd.n2804 vdd.n901 185
R17212 vdd.n2806 vdd.n900 185
R17213 vdd.n2975 vdd.n900 185
R17214 vdd.n2849 vdd.n2848 185
R17215 vdd.n2848 vdd.n2847 185
R17216 vdd.n2850 vdd.n907 185
R17217 vdd.n2969 vdd.n907 185
R17218 vdd.n2852 vdd.n2851 185
R17219 vdd.n2851 vdd.n905 185
R17220 vdd.n2853 vdd.n913 185
R17221 vdd.n2963 vdd.n913 185
R17222 vdd.n2855 vdd.n2854 185
R17223 vdd.n2854 vdd.n911 185
R17224 vdd.n2856 vdd.n919 185
R17225 vdd.n2957 vdd.n919 185
R17226 vdd.n2858 vdd.n2857 185
R17227 vdd.n2857 vdd.n917 185
R17228 vdd.n2859 vdd.n924 185
R17229 vdd.n2951 vdd.n924 185
R17230 vdd.n2861 vdd.n2860 185
R17231 vdd.n2862 vdd.n2861 185
R17232 vdd.n2774 vdd.n930 185
R17233 vdd.n2945 vdd.n930 185
R17234 vdd.n2773 vdd.n2772 185
R17235 vdd.n2772 vdd.n928 185
R17236 vdd.n2264 vdd.n2263 185
R17237 vdd.n2265 vdd.n2264 185
R17238 vdd.n1438 vdd.n1436 185
R17239 vdd.n2256 vdd.n1436 185
R17240 vdd.n2259 vdd.n2258 185
R17241 vdd.n2258 vdd.n2257 185
R17242 vdd.n1441 vdd.n1440 185
R17243 vdd.n1442 vdd.n1441 185
R17244 vdd.n2245 vdd.n2244 185
R17245 vdd.n2246 vdd.n2245 185
R17246 vdd.n1450 vdd.n1449 185
R17247 vdd.n2237 vdd.n1449 185
R17248 vdd.n2240 vdd.n2239 185
R17249 vdd.n2239 vdd.n2238 185
R17250 vdd.n1453 vdd.n1452 185
R17251 vdd.n1460 vdd.n1453 185
R17252 vdd.n2228 vdd.n2227 185
R17253 vdd.n2229 vdd.n2228 185
R17254 vdd.n1462 vdd.n1461 185
R17255 vdd.n1461 vdd.n1459 185
R17256 vdd.n2223 vdd.n2222 185
R17257 vdd.n2222 vdd.n2221 185
R17258 vdd.n1465 vdd.n1464 185
R17259 vdd.n1466 vdd.n1465 185
R17260 vdd.n2212 vdd.n2211 185
R17261 vdd.n2213 vdd.n2212 185
R17262 vdd.n1473 vdd.n1472 185
R17263 vdd.n2204 vdd.n1472 185
R17264 vdd.n2207 vdd.n2206 185
R17265 vdd.n2206 vdd.n2205 185
R17266 vdd.n1476 vdd.n1475 185
R17267 vdd.n1482 vdd.n1476 185
R17268 vdd.n2195 vdd.n2194 185
R17269 vdd.n2196 vdd.n2195 185
R17270 vdd.n1484 vdd.n1483 185
R17271 vdd.n2187 vdd.n1483 185
R17272 vdd.n2190 vdd.n2189 185
R17273 vdd.n2189 vdd.n2188 185
R17274 vdd.n1487 vdd.n1486 185
R17275 vdd.n1488 vdd.n1487 185
R17276 vdd.n2178 vdd.n2177 185
R17277 vdd.n2179 vdd.n2178 185
R17278 vdd.n1496 vdd.n1495 185
R17279 vdd.n1495 vdd.n1494 185
R17280 vdd.n1866 vdd.n1865 185
R17281 vdd.n1865 vdd.n1864 185
R17282 vdd.n1499 vdd.n1498 185
R17283 vdd.n1505 vdd.n1499 185
R17284 vdd.n1855 vdd.n1854 185
R17285 vdd.n1856 vdd.n1855 185
R17286 vdd.n1507 vdd.n1506 185
R17287 vdd.n1847 vdd.n1506 185
R17288 vdd.n1850 vdd.n1849 185
R17289 vdd.n1849 vdd.n1848 185
R17290 vdd.n1510 vdd.n1509 185
R17291 vdd.n1517 vdd.n1510 185
R17292 vdd.n1838 vdd.n1837 185
R17293 vdd.n1839 vdd.n1838 185
R17294 vdd.n1519 vdd.n1518 185
R17295 vdd.n1518 vdd.n1516 185
R17296 vdd.n1833 vdd.n1832 185
R17297 vdd.n1832 vdd.n1831 185
R17298 vdd.n1522 vdd.n1521 185
R17299 vdd.n1523 vdd.n1522 185
R17300 vdd.n1822 vdd.n1821 185
R17301 vdd.n1823 vdd.n1822 185
R17302 vdd.n1530 vdd.n1529 185
R17303 vdd.n1814 vdd.n1529 185
R17304 vdd.n1817 vdd.n1816 185
R17305 vdd.n1816 vdd.n1815 185
R17306 vdd.n1533 vdd.n1532 185
R17307 vdd.n1539 vdd.n1533 185
R17308 vdd.n1805 vdd.n1804 185
R17309 vdd.n1806 vdd.n1805 185
R17310 vdd.n1541 vdd.n1540 185
R17311 vdd.n1797 vdd.n1540 185
R17312 vdd.n1800 vdd.n1799 185
R17313 vdd.n1799 vdd.n1798 185
R17314 vdd.n1544 vdd.n1543 185
R17315 vdd.n1545 vdd.n1544 185
R17316 vdd.n1788 vdd.n1787 185
R17317 vdd.n1789 vdd.n1788 185
R17318 vdd.n1552 vdd.n1551 185
R17319 vdd.n1587 vdd.n1551 185
R17320 vdd.n1783 vdd.n1782 185
R17321 vdd.n1555 vdd.n1554 185
R17322 vdd.n1779 vdd.n1778 185
R17323 vdd.n1780 vdd.n1779 185
R17324 vdd.n1589 vdd.n1588 185
R17325 vdd.n1774 vdd.n1591 185
R17326 vdd.n1773 vdd.n1592 185
R17327 vdd.n1772 vdd.n1593 185
R17328 vdd.n1595 vdd.n1594 185
R17329 vdd.n1768 vdd.n1597 185
R17330 vdd.n1767 vdd.n1598 185
R17331 vdd.n1766 vdd.n1599 185
R17332 vdd.n1601 vdd.n1600 185
R17333 vdd.n1762 vdd.n1603 185
R17334 vdd.n1761 vdd.n1604 185
R17335 vdd.n1760 vdd.n1605 185
R17336 vdd.n1607 vdd.n1606 185
R17337 vdd.n1756 vdd.n1609 185
R17338 vdd.n1755 vdd.n1610 185
R17339 vdd.n1754 vdd.n1611 185
R17340 vdd.n1615 vdd.n1612 185
R17341 vdd.n1750 vdd.n1617 185
R17342 vdd.n1749 vdd.n1618 185
R17343 vdd.n1748 vdd.n1619 185
R17344 vdd.n1621 vdd.n1620 185
R17345 vdd.n1744 vdd.n1623 185
R17346 vdd.n1743 vdd.n1624 185
R17347 vdd.n1742 vdd.n1625 185
R17348 vdd.n1627 vdd.n1626 185
R17349 vdd.n1738 vdd.n1629 185
R17350 vdd.n1737 vdd.n1630 185
R17351 vdd.n1736 vdd.n1631 185
R17352 vdd.n1633 vdd.n1632 185
R17353 vdd.n1732 vdd.n1635 185
R17354 vdd.n1731 vdd.n1636 185
R17355 vdd.n1730 vdd.n1637 185
R17356 vdd.n1639 vdd.n1638 185
R17357 vdd.n1726 vdd.n1641 185
R17358 vdd.n1725 vdd.n1642 185
R17359 vdd.n1724 vdd.n1643 185
R17360 vdd.n1645 vdd.n1644 185
R17361 vdd.n1720 vdd.n1647 185
R17362 vdd.n1719 vdd.n1716 185
R17363 vdd.n1715 vdd.n1648 185
R17364 vdd.n1650 vdd.n1649 185
R17365 vdd.n1711 vdd.n1652 185
R17366 vdd.n1710 vdd.n1653 185
R17367 vdd.n1709 vdd.n1654 185
R17368 vdd.n1656 vdd.n1655 185
R17369 vdd.n1705 vdd.n1658 185
R17370 vdd.n1704 vdd.n1659 185
R17371 vdd.n1703 vdd.n1660 185
R17372 vdd.n1662 vdd.n1661 185
R17373 vdd.n1699 vdd.n1664 185
R17374 vdd.n1698 vdd.n1665 185
R17375 vdd.n1697 vdd.n1666 185
R17376 vdd.n1668 vdd.n1667 185
R17377 vdd.n1693 vdd.n1670 185
R17378 vdd.n1692 vdd.n1671 185
R17379 vdd.n1691 vdd.n1672 185
R17380 vdd.n1674 vdd.n1673 185
R17381 vdd.n1687 vdd.n1676 185
R17382 vdd.n1686 vdd.n1677 185
R17383 vdd.n1685 vdd.n1678 185
R17384 vdd.n1682 vdd.n1586 185
R17385 vdd.n1780 vdd.n1586 185
R17386 vdd.n2268 vdd.n2267 185
R17387 vdd.n2272 vdd.n1432 185
R17388 vdd.n1431 vdd.n1425 185
R17389 vdd.n1429 vdd.n1428 185
R17390 vdd.n1427 vdd.n1221 185
R17391 vdd.n2276 vdd.n1218 185
R17392 vdd.n2278 vdd.n2277 185
R17393 vdd.n2280 vdd.n1216 185
R17394 vdd.n2282 vdd.n2281 185
R17395 vdd.n2283 vdd.n1211 185
R17396 vdd.n2285 vdd.n2284 185
R17397 vdd.n2287 vdd.n1209 185
R17398 vdd.n2289 vdd.n2288 185
R17399 vdd.n2290 vdd.n1204 185
R17400 vdd.n2292 vdd.n2291 185
R17401 vdd.n2294 vdd.n1202 185
R17402 vdd.n2296 vdd.n2295 185
R17403 vdd.n2297 vdd.n1198 185
R17404 vdd.n2299 vdd.n2298 185
R17405 vdd.n2301 vdd.n1195 185
R17406 vdd.n2303 vdd.n2302 185
R17407 vdd.n1196 vdd.n1189 185
R17408 vdd.n2307 vdd.n1193 185
R17409 vdd.n2308 vdd.n1185 185
R17410 vdd.n2310 vdd.n2309 185
R17411 vdd.n2312 vdd.n1183 185
R17412 vdd.n2314 vdd.n2313 185
R17413 vdd.n2315 vdd.n1178 185
R17414 vdd.n2317 vdd.n2316 185
R17415 vdd.n2319 vdd.n1176 185
R17416 vdd.n2321 vdd.n2320 185
R17417 vdd.n2322 vdd.n1171 185
R17418 vdd.n2324 vdd.n2323 185
R17419 vdd.n2326 vdd.n1169 185
R17420 vdd.n2328 vdd.n2327 185
R17421 vdd.n2329 vdd.n1164 185
R17422 vdd.n2331 vdd.n2330 185
R17423 vdd.n2333 vdd.n1162 185
R17424 vdd.n2335 vdd.n2334 185
R17425 vdd.n2336 vdd.n1158 185
R17426 vdd.n2338 vdd.n2337 185
R17427 vdd.n2340 vdd.n1155 185
R17428 vdd.n2342 vdd.n2341 185
R17429 vdd.n1156 vdd.n1149 185
R17430 vdd.n2346 vdd.n1153 185
R17431 vdd.n2347 vdd.n1145 185
R17432 vdd.n2349 vdd.n2348 185
R17433 vdd.n2351 vdd.n1143 185
R17434 vdd.n2353 vdd.n2352 185
R17435 vdd.n2354 vdd.n1138 185
R17436 vdd.n2356 vdd.n2355 185
R17437 vdd.n2358 vdd.n1136 185
R17438 vdd.n2360 vdd.n2359 185
R17439 vdd.n2361 vdd.n1131 185
R17440 vdd.n2363 vdd.n2362 185
R17441 vdd.n2365 vdd.n1129 185
R17442 vdd.n2367 vdd.n2366 185
R17443 vdd.n2368 vdd.n1127 185
R17444 vdd.n2370 vdd.n2369 185
R17445 vdd.n2373 vdd.n2372 185
R17446 vdd.n2375 vdd.n2374 185
R17447 vdd.n2377 vdd.n1125 185
R17448 vdd.n2379 vdd.n2378 185
R17449 vdd.n1437 vdd.n1124 185
R17450 vdd.n2266 vdd.n1435 185
R17451 vdd.n2266 vdd.n2265 185
R17452 vdd.n1445 vdd.n1434 185
R17453 vdd.n2256 vdd.n1434 185
R17454 vdd.n2255 vdd.n2254 185
R17455 vdd.n2257 vdd.n2255 185
R17456 vdd.n1444 vdd.n1443 185
R17457 vdd.n1443 vdd.n1442 185
R17458 vdd.n2248 vdd.n2247 185
R17459 vdd.n2247 vdd.n2246 185
R17460 vdd.n1448 vdd.n1447 185
R17461 vdd.n2237 vdd.n1448 185
R17462 vdd.n2236 vdd.n2235 185
R17463 vdd.n2238 vdd.n2236 185
R17464 vdd.n1455 vdd.n1454 185
R17465 vdd.n1460 vdd.n1454 185
R17466 vdd.n2231 vdd.n2230 185
R17467 vdd.n2230 vdd.n2229 185
R17468 vdd.n1458 vdd.n1457 185
R17469 vdd.n1459 vdd.n1458 185
R17470 vdd.n2220 vdd.n2219 185
R17471 vdd.n2221 vdd.n2220 185
R17472 vdd.n1468 vdd.n1467 185
R17473 vdd.n1467 vdd.n1466 185
R17474 vdd.n2215 vdd.n2214 185
R17475 vdd.n2214 vdd.n2213 185
R17476 vdd.n1471 vdd.n1470 185
R17477 vdd.n2204 vdd.n1471 185
R17478 vdd.n2203 vdd.n2202 185
R17479 vdd.n2205 vdd.n2203 185
R17480 vdd.n1478 vdd.n1477 185
R17481 vdd.n1482 vdd.n1477 185
R17482 vdd.n2198 vdd.n2197 185
R17483 vdd.n2197 vdd.n2196 185
R17484 vdd.n1481 vdd.n1480 185
R17485 vdd.n2187 vdd.n1481 185
R17486 vdd.n2186 vdd.n2185 185
R17487 vdd.n2188 vdd.n2186 185
R17488 vdd.n1490 vdd.n1489 185
R17489 vdd.n1489 vdd.n1488 185
R17490 vdd.n2181 vdd.n2180 185
R17491 vdd.n2180 vdd.n2179 185
R17492 vdd.n1493 vdd.n1492 185
R17493 vdd.n1494 vdd.n1493 185
R17494 vdd.n1863 vdd.n1862 185
R17495 vdd.n1864 vdd.n1863 185
R17496 vdd.n1501 vdd.n1500 185
R17497 vdd.n1505 vdd.n1500 185
R17498 vdd.n1858 vdd.n1857 185
R17499 vdd.n1857 vdd.n1856 185
R17500 vdd.n1504 vdd.n1503 185
R17501 vdd.n1847 vdd.n1504 185
R17502 vdd.n1846 vdd.n1845 185
R17503 vdd.n1848 vdd.n1846 185
R17504 vdd.n1512 vdd.n1511 185
R17505 vdd.n1517 vdd.n1511 185
R17506 vdd.n1841 vdd.n1840 185
R17507 vdd.n1840 vdd.n1839 185
R17508 vdd.n1515 vdd.n1514 185
R17509 vdd.n1516 vdd.n1515 185
R17510 vdd.n1830 vdd.n1829 185
R17511 vdd.n1831 vdd.n1830 185
R17512 vdd.n1525 vdd.n1524 185
R17513 vdd.n1524 vdd.n1523 185
R17514 vdd.n1825 vdd.n1824 185
R17515 vdd.n1824 vdd.n1823 185
R17516 vdd.n1528 vdd.n1527 185
R17517 vdd.n1814 vdd.n1528 185
R17518 vdd.n1813 vdd.n1812 185
R17519 vdd.n1815 vdd.n1813 185
R17520 vdd.n1535 vdd.n1534 185
R17521 vdd.n1539 vdd.n1534 185
R17522 vdd.n1808 vdd.n1807 185
R17523 vdd.n1807 vdd.n1806 185
R17524 vdd.n1538 vdd.n1537 185
R17525 vdd.n1797 vdd.n1538 185
R17526 vdd.n1796 vdd.n1795 185
R17527 vdd.n1798 vdd.n1796 185
R17528 vdd.n1547 vdd.n1546 185
R17529 vdd.n1546 vdd.n1545 185
R17530 vdd.n1791 vdd.n1790 185
R17531 vdd.n1790 vdd.n1789 185
R17532 vdd.n1550 vdd.n1549 185
R17533 vdd.n1587 vdd.n1550 185
R17534 vdd.n971 vdd.n969 185
R17535 vdd.n2593 vdd.n969 185
R17536 vdd.n2515 vdd.n989 185
R17537 vdd.n989 vdd.n976 185
R17538 vdd.n2517 vdd.n2516 185
R17539 vdd.n2518 vdd.n2517 185
R17540 vdd.n2514 vdd.n988 185
R17541 vdd.n1338 vdd.n988 185
R17542 vdd.n2513 vdd.n2512 185
R17543 vdd.n2512 vdd.n2511 185
R17544 vdd.n991 vdd.n990 185
R17545 vdd.n992 vdd.n991 185
R17546 vdd.n2502 vdd.n2501 185
R17547 vdd.n2503 vdd.n2502 185
R17548 vdd.n2500 vdd.n1002 185
R17549 vdd.n1002 vdd.n999 185
R17550 vdd.n2499 vdd.n2498 185
R17551 vdd.n2498 vdd.n2497 185
R17552 vdd.n1004 vdd.n1003 185
R17553 vdd.n1005 vdd.n1004 185
R17554 vdd.n2490 vdd.n2489 185
R17555 vdd.n2491 vdd.n2490 185
R17556 vdd.n2488 vdd.n1013 185
R17557 vdd.n1018 vdd.n1013 185
R17558 vdd.n2487 vdd.n2486 185
R17559 vdd.n2486 vdd.n2485 185
R17560 vdd.n1015 vdd.n1014 185
R17561 vdd.n1024 vdd.n1015 185
R17562 vdd.n2478 vdd.n2477 185
R17563 vdd.n2479 vdd.n2478 185
R17564 vdd.n2476 vdd.n1025 185
R17565 vdd.n1359 vdd.n1025 185
R17566 vdd.n2475 vdd.n2474 185
R17567 vdd.n2474 vdd.n2473 185
R17568 vdd.n1027 vdd.n1026 185
R17569 vdd.n1028 vdd.n1027 185
R17570 vdd.n2466 vdd.n2465 185
R17571 vdd.n2467 vdd.n2466 185
R17572 vdd.n2464 vdd.n1037 185
R17573 vdd.n1037 vdd.n1034 185
R17574 vdd.n2463 vdd.n2462 185
R17575 vdd.n2462 vdd.n2461 185
R17576 vdd.n1039 vdd.n1038 185
R17577 vdd.n1048 vdd.n1039 185
R17578 vdd.n2453 vdd.n2452 185
R17579 vdd.n2454 vdd.n2453 185
R17580 vdd.n2451 vdd.n1049 185
R17581 vdd.n1055 vdd.n1049 185
R17582 vdd.n2450 vdd.n2449 185
R17583 vdd.n2449 vdd.n2448 185
R17584 vdd.n1051 vdd.n1050 185
R17585 vdd.n1052 vdd.n1051 185
R17586 vdd.n2441 vdd.n2440 185
R17587 vdd.n2442 vdd.n2441 185
R17588 vdd.n2439 vdd.n1062 185
R17589 vdd.n1062 vdd.n1059 185
R17590 vdd.n2438 vdd.n2437 185
R17591 vdd.n2437 vdd.n2436 185
R17592 vdd.n1064 vdd.n1063 185
R17593 vdd.n1065 vdd.n1064 185
R17594 vdd.n2429 vdd.n2428 185
R17595 vdd.n2430 vdd.n2429 185
R17596 vdd.n2427 vdd.n1073 185
R17597 vdd.n1079 vdd.n1073 185
R17598 vdd.n2426 vdd.n2425 185
R17599 vdd.n2425 vdd.n2424 185
R17600 vdd.n1075 vdd.n1074 185
R17601 vdd.n1076 vdd.n1075 185
R17602 vdd.n2415 vdd.n2414 185
R17603 vdd.n2413 vdd.n1118 185
R17604 vdd.n2412 vdd.n1117 185
R17605 vdd.n2417 vdd.n1117 185
R17606 vdd.n2411 vdd.n2410 185
R17607 vdd.n2409 vdd.n2408 185
R17608 vdd.n2407 vdd.n2406 185
R17609 vdd.n2405 vdd.n2404 185
R17610 vdd.n2403 vdd.n2402 185
R17611 vdd.n2401 vdd.n2400 185
R17612 vdd.n2399 vdd.n2398 185
R17613 vdd.n2397 vdd.n2396 185
R17614 vdd.n2395 vdd.n2394 185
R17615 vdd.n2393 vdd.n2392 185
R17616 vdd.n2391 vdd.n2390 185
R17617 vdd.n2389 vdd.n2388 185
R17618 vdd.n2387 vdd.n2386 185
R17619 vdd.n2385 vdd.n2384 185
R17620 vdd.n2383 vdd.n2382 185
R17621 vdd.n1275 vdd.n1119 185
R17622 vdd.n1277 vdd.n1276 185
R17623 vdd.n1279 vdd.n1278 185
R17624 vdd.n1281 vdd.n1280 185
R17625 vdd.n1283 vdd.n1282 185
R17626 vdd.n1285 vdd.n1284 185
R17627 vdd.n1287 vdd.n1286 185
R17628 vdd.n1289 vdd.n1288 185
R17629 vdd.n1291 vdd.n1290 185
R17630 vdd.n1293 vdd.n1292 185
R17631 vdd.n1295 vdd.n1294 185
R17632 vdd.n1297 vdd.n1296 185
R17633 vdd.n1299 vdd.n1298 185
R17634 vdd.n1301 vdd.n1300 185
R17635 vdd.n1304 vdd.n1303 185
R17636 vdd.n1306 vdd.n1305 185
R17637 vdd.n1308 vdd.n1307 185
R17638 vdd.n2596 vdd.n2595 185
R17639 vdd.n2598 vdd.n2597 185
R17640 vdd.n2600 vdd.n2599 185
R17641 vdd.n2603 vdd.n2602 185
R17642 vdd.n2605 vdd.n2604 185
R17643 vdd.n2607 vdd.n2606 185
R17644 vdd.n2609 vdd.n2608 185
R17645 vdd.n2611 vdd.n2610 185
R17646 vdd.n2613 vdd.n2612 185
R17647 vdd.n2615 vdd.n2614 185
R17648 vdd.n2617 vdd.n2616 185
R17649 vdd.n2619 vdd.n2618 185
R17650 vdd.n2621 vdd.n2620 185
R17651 vdd.n2623 vdd.n2622 185
R17652 vdd.n2625 vdd.n2624 185
R17653 vdd.n2627 vdd.n2626 185
R17654 vdd.n2629 vdd.n2628 185
R17655 vdd.n2631 vdd.n2630 185
R17656 vdd.n2633 vdd.n2632 185
R17657 vdd.n2635 vdd.n2634 185
R17658 vdd.n2637 vdd.n2636 185
R17659 vdd.n2639 vdd.n2638 185
R17660 vdd.n2641 vdd.n2640 185
R17661 vdd.n2643 vdd.n2642 185
R17662 vdd.n2645 vdd.n2644 185
R17663 vdd.n2647 vdd.n2646 185
R17664 vdd.n2649 vdd.n2648 185
R17665 vdd.n2651 vdd.n2650 185
R17666 vdd.n2653 vdd.n2652 185
R17667 vdd.n2655 vdd.n2654 185
R17668 vdd.n2657 vdd.n2656 185
R17669 vdd.n2659 vdd.n2658 185
R17670 vdd.n2661 vdd.n2660 185
R17671 vdd.n2662 vdd.n970 185
R17672 vdd.n2664 vdd.n2663 185
R17673 vdd.n2665 vdd.n2664 185
R17674 vdd.n2594 vdd.n974 185
R17675 vdd.n2594 vdd.n2593 185
R17676 vdd.n1336 vdd.n975 185
R17677 vdd.n976 vdd.n975 185
R17678 vdd.n1337 vdd.n986 185
R17679 vdd.n2518 vdd.n986 185
R17680 vdd.n1340 vdd.n1339 185
R17681 vdd.n1339 vdd.n1338 185
R17682 vdd.n1341 vdd.n993 185
R17683 vdd.n2511 vdd.n993 185
R17684 vdd.n1343 vdd.n1342 185
R17685 vdd.n1342 vdd.n992 185
R17686 vdd.n1344 vdd.n1000 185
R17687 vdd.n2503 vdd.n1000 185
R17688 vdd.n1346 vdd.n1345 185
R17689 vdd.n1345 vdd.n999 185
R17690 vdd.n1347 vdd.n1006 185
R17691 vdd.n2497 vdd.n1006 185
R17692 vdd.n1349 vdd.n1348 185
R17693 vdd.n1348 vdd.n1005 185
R17694 vdd.n1350 vdd.n1011 185
R17695 vdd.n2491 vdd.n1011 185
R17696 vdd.n1352 vdd.n1351 185
R17697 vdd.n1351 vdd.n1018 185
R17698 vdd.n1353 vdd.n1016 185
R17699 vdd.n2485 vdd.n1016 185
R17700 vdd.n1355 vdd.n1354 185
R17701 vdd.n1354 vdd.n1024 185
R17702 vdd.n1356 vdd.n1022 185
R17703 vdd.n2479 vdd.n1022 185
R17704 vdd.n1358 vdd.n1357 185
R17705 vdd.n1359 vdd.n1358 185
R17706 vdd.n1335 vdd.n1029 185
R17707 vdd.n2473 vdd.n1029 185
R17708 vdd.n1334 vdd.n1333 185
R17709 vdd.n1333 vdd.n1028 185
R17710 vdd.n1332 vdd.n1035 185
R17711 vdd.n2467 vdd.n1035 185
R17712 vdd.n1331 vdd.n1330 185
R17713 vdd.n1330 vdd.n1034 185
R17714 vdd.n1329 vdd.n1040 185
R17715 vdd.n2461 vdd.n1040 185
R17716 vdd.n1328 vdd.n1327 185
R17717 vdd.n1327 vdd.n1048 185
R17718 vdd.n1326 vdd.n1046 185
R17719 vdd.n2454 vdd.n1046 185
R17720 vdd.n1325 vdd.n1324 185
R17721 vdd.n1324 vdd.n1055 185
R17722 vdd.n1323 vdd.n1053 185
R17723 vdd.n2448 vdd.n1053 185
R17724 vdd.n1322 vdd.n1321 185
R17725 vdd.n1321 vdd.n1052 185
R17726 vdd.n1320 vdd.n1060 185
R17727 vdd.n2442 vdd.n1060 185
R17728 vdd.n1319 vdd.n1318 185
R17729 vdd.n1318 vdd.n1059 185
R17730 vdd.n1317 vdd.n1066 185
R17731 vdd.n2436 vdd.n1066 185
R17732 vdd.n1316 vdd.n1315 185
R17733 vdd.n1315 vdd.n1065 185
R17734 vdd.n1314 vdd.n1071 185
R17735 vdd.n2430 vdd.n1071 185
R17736 vdd.n1313 vdd.n1312 185
R17737 vdd.n1312 vdd.n1079 185
R17738 vdd.n1311 vdd.n1077 185
R17739 vdd.n2424 vdd.n1077 185
R17740 vdd.n1310 vdd.n1309 185
R17741 vdd.n1309 vdd.n1076 185
R17742 vdd.n3449 vdd.n3448 185
R17743 vdd.n3448 vdd.n3447 185
R17744 vdd.n3450 vdd.n387 185
R17745 vdd.n387 vdd.n386 185
R17746 vdd.n3452 vdd.n3451 185
R17747 vdd.n3453 vdd.n3452 185
R17748 vdd.n382 vdd.n381 185
R17749 vdd.n3454 vdd.n382 185
R17750 vdd.n3457 vdd.n3456 185
R17751 vdd.n3456 vdd.n3455 185
R17752 vdd.n3458 vdd.n376 185
R17753 vdd.n376 vdd.n375 185
R17754 vdd.n3460 vdd.n3459 185
R17755 vdd.n3461 vdd.n3460 185
R17756 vdd.n371 vdd.n370 185
R17757 vdd.n3462 vdd.n371 185
R17758 vdd.n3465 vdd.n3464 185
R17759 vdd.n3464 vdd.n3463 185
R17760 vdd.n3466 vdd.n365 185
R17761 vdd.n3423 vdd.n365 185
R17762 vdd.n3468 vdd.n3467 185
R17763 vdd.n3469 vdd.n3468 185
R17764 vdd.n360 vdd.n359 185
R17765 vdd.n3470 vdd.n360 185
R17766 vdd.n3473 vdd.n3472 185
R17767 vdd.n3472 vdd.n3471 185
R17768 vdd.n3474 vdd.n354 185
R17769 vdd.n361 vdd.n354 185
R17770 vdd.n3476 vdd.n3475 185
R17771 vdd.n3477 vdd.n3476 185
R17772 vdd.n350 vdd.n349 185
R17773 vdd.n3478 vdd.n350 185
R17774 vdd.n3481 vdd.n3480 185
R17775 vdd.n3480 vdd.n3479 185
R17776 vdd.n3482 vdd.n345 185
R17777 vdd.n345 vdd.n344 185
R17778 vdd.n3484 vdd.n3483 185
R17779 vdd.n3485 vdd.n3484 185
R17780 vdd.n339 vdd.n337 185
R17781 vdd.n3486 vdd.n339 185
R17782 vdd.n3489 vdd.n3488 185
R17783 vdd.n3488 vdd.n3487 185
R17784 vdd.n338 vdd.n336 185
R17785 vdd.n340 vdd.n338 185
R17786 vdd.n3399 vdd.n3398 185
R17787 vdd.n3400 vdd.n3399 185
R17788 vdd.n635 vdd.n634 185
R17789 vdd.n634 vdd.n633 185
R17790 vdd.n3394 vdd.n3393 185
R17791 vdd.n3393 vdd.n3392 185
R17792 vdd.n638 vdd.n637 185
R17793 vdd.n644 vdd.n638 185
R17794 vdd.n3380 vdd.n3379 185
R17795 vdd.n3381 vdd.n3380 185
R17796 vdd.n646 vdd.n645 185
R17797 vdd.n3372 vdd.n645 185
R17798 vdd.n3375 vdd.n3374 185
R17799 vdd.n3374 vdd.n3373 185
R17800 vdd.n649 vdd.n648 185
R17801 vdd.n656 vdd.n649 185
R17802 vdd.n3363 vdd.n3362 185
R17803 vdd.n3364 vdd.n3363 185
R17804 vdd.n658 vdd.n657 185
R17805 vdd.n657 vdd.n655 185
R17806 vdd.n3358 vdd.n3357 185
R17807 vdd.n3357 vdd.n3356 185
R17808 vdd.n661 vdd.n660 185
R17809 vdd.n662 vdd.n661 185
R17810 vdd.n3347 vdd.n3346 185
R17811 vdd.n3348 vdd.n3347 185
R17812 vdd.n669 vdd.n668 185
R17813 vdd.n3339 vdd.n668 185
R17814 vdd.n3342 vdd.n3341 185
R17815 vdd.n3341 vdd.n3340 185
R17816 vdd.n672 vdd.n671 185
R17817 vdd.n679 vdd.n672 185
R17818 vdd.n3330 vdd.n3329 185
R17819 vdd.n3331 vdd.n3330 185
R17820 vdd.n681 vdd.n680 185
R17821 vdd.n680 vdd.n678 185
R17822 vdd.n3325 vdd.n3324 185
R17823 vdd.n3324 vdd.n3323 185
R17824 vdd.n684 vdd.n683 185
R17825 vdd.n723 vdd.n684 185
R17826 vdd.n3313 vdd.n3312 185
R17827 vdd.n3311 vdd.n725 185
R17828 vdd.n3310 vdd.n724 185
R17829 vdd.n3315 vdd.n724 185
R17830 vdd.n729 vdd.n728 185
R17831 vdd.n733 vdd.n732 185
R17832 vdd.n3306 vdd.n734 185
R17833 vdd.n3305 vdd.n3304 185
R17834 vdd.n3303 vdd.n3302 185
R17835 vdd.n3301 vdd.n3300 185
R17836 vdd.n3299 vdd.n3298 185
R17837 vdd.n3297 vdd.n3296 185
R17838 vdd.n3295 vdd.n3294 185
R17839 vdd.n3293 vdd.n3292 185
R17840 vdd.n3291 vdd.n3290 185
R17841 vdd.n3289 vdd.n3288 185
R17842 vdd.n3287 vdd.n3286 185
R17843 vdd.n3285 vdd.n3284 185
R17844 vdd.n3283 vdd.n3282 185
R17845 vdd.n3281 vdd.n3280 185
R17846 vdd.n3279 vdd.n3278 185
R17847 vdd.n3270 vdd.n747 185
R17848 vdd.n3272 vdd.n3271 185
R17849 vdd.n3269 vdd.n3268 185
R17850 vdd.n3267 vdd.n3266 185
R17851 vdd.n3265 vdd.n3264 185
R17852 vdd.n3263 vdd.n3262 185
R17853 vdd.n3261 vdd.n3260 185
R17854 vdd.n3259 vdd.n3258 185
R17855 vdd.n3257 vdd.n3256 185
R17856 vdd.n3255 vdd.n3254 185
R17857 vdd.n3253 vdd.n3252 185
R17858 vdd.n3251 vdd.n3250 185
R17859 vdd.n3249 vdd.n3248 185
R17860 vdd.n3247 vdd.n3246 185
R17861 vdd.n3245 vdd.n3244 185
R17862 vdd.n3243 vdd.n3242 185
R17863 vdd.n3241 vdd.n3240 185
R17864 vdd.n3239 vdd.n3238 185
R17865 vdd.n3237 vdd.n3236 185
R17866 vdd.n3235 vdd.n3234 185
R17867 vdd.n3233 vdd.n3232 185
R17868 vdd.n3231 vdd.n3230 185
R17869 vdd.n3224 vdd.n767 185
R17870 vdd.n3226 vdd.n3225 185
R17871 vdd.n3223 vdd.n3222 185
R17872 vdd.n3221 vdd.n3220 185
R17873 vdd.n3219 vdd.n3218 185
R17874 vdd.n3217 vdd.n3216 185
R17875 vdd.n3215 vdd.n3214 185
R17876 vdd.n3213 vdd.n3212 185
R17877 vdd.n3211 vdd.n3210 185
R17878 vdd.n3209 vdd.n3208 185
R17879 vdd.n3207 vdd.n3206 185
R17880 vdd.n3205 vdd.n3204 185
R17881 vdd.n3203 vdd.n3202 185
R17882 vdd.n3201 vdd.n3200 185
R17883 vdd.n3199 vdd.n3198 185
R17884 vdd.n3197 vdd.n3196 185
R17885 vdd.n3195 vdd.n3194 185
R17886 vdd.n3193 vdd.n3192 185
R17887 vdd.n3191 vdd.n3190 185
R17888 vdd.n3189 vdd.n3188 185
R17889 vdd.n3187 vdd.n691 185
R17890 vdd.n3317 vdd.n3316 185
R17891 vdd.n3316 vdd.n3315 185
R17892 vdd.n3444 vdd.n3443 185
R17893 vdd.n618 vdd.n425 185
R17894 vdd.n617 vdd.n616 185
R17895 vdd.n615 vdd.n614 185
R17896 vdd.n613 vdd.n430 185
R17897 vdd.n609 vdd.n608 185
R17898 vdd.n607 vdd.n606 185
R17899 vdd.n605 vdd.n604 185
R17900 vdd.n603 vdd.n432 185
R17901 vdd.n599 vdd.n598 185
R17902 vdd.n597 vdd.n596 185
R17903 vdd.n595 vdd.n594 185
R17904 vdd.n593 vdd.n434 185
R17905 vdd.n589 vdd.n588 185
R17906 vdd.n587 vdd.n586 185
R17907 vdd.n585 vdd.n584 185
R17908 vdd.n583 vdd.n436 185
R17909 vdd.n579 vdd.n578 185
R17910 vdd.n577 vdd.n576 185
R17911 vdd.n575 vdd.n574 185
R17912 vdd.n573 vdd.n438 185
R17913 vdd.n569 vdd.n568 185
R17914 vdd.n567 vdd.n566 185
R17915 vdd.n565 vdd.n564 185
R17916 vdd.n563 vdd.n442 185
R17917 vdd.n559 vdd.n558 185
R17918 vdd.n557 vdd.n556 185
R17919 vdd.n555 vdd.n554 185
R17920 vdd.n553 vdd.n444 185
R17921 vdd.n549 vdd.n548 185
R17922 vdd.n547 vdd.n546 185
R17923 vdd.n545 vdd.n544 185
R17924 vdd.n543 vdd.n446 185
R17925 vdd.n539 vdd.n538 185
R17926 vdd.n537 vdd.n536 185
R17927 vdd.n535 vdd.n534 185
R17928 vdd.n533 vdd.n448 185
R17929 vdd.n529 vdd.n528 185
R17930 vdd.n527 vdd.n526 185
R17931 vdd.n525 vdd.n524 185
R17932 vdd.n523 vdd.n450 185
R17933 vdd.n519 vdd.n518 185
R17934 vdd.n517 vdd.n516 185
R17935 vdd.n515 vdd.n514 185
R17936 vdd.n513 vdd.n454 185
R17937 vdd.n509 vdd.n508 185
R17938 vdd.n507 vdd.n506 185
R17939 vdd.n505 vdd.n504 185
R17940 vdd.n503 vdd.n456 185
R17941 vdd.n499 vdd.n498 185
R17942 vdd.n497 vdd.n496 185
R17943 vdd.n495 vdd.n494 185
R17944 vdd.n493 vdd.n458 185
R17945 vdd.n489 vdd.n488 185
R17946 vdd.n487 vdd.n486 185
R17947 vdd.n485 vdd.n484 185
R17948 vdd.n483 vdd.n460 185
R17949 vdd.n479 vdd.n478 185
R17950 vdd.n477 vdd.n476 185
R17951 vdd.n475 vdd.n474 185
R17952 vdd.n473 vdd.n462 185
R17953 vdd.n469 vdd.n468 185
R17954 vdd.n467 vdd.n466 185
R17955 vdd.n465 vdd.n392 185
R17956 vdd.n3440 vdd.n393 185
R17957 vdd.n3447 vdd.n393 185
R17958 vdd.n3439 vdd.n3438 185
R17959 vdd.n3438 vdd.n386 185
R17960 vdd.n3437 vdd.n385 185
R17961 vdd.n3453 vdd.n385 185
R17962 vdd.n621 vdd.n384 185
R17963 vdd.n3454 vdd.n384 185
R17964 vdd.n3433 vdd.n383 185
R17965 vdd.n3455 vdd.n383 185
R17966 vdd.n3432 vdd.n3431 185
R17967 vdd.n3431 vdd.n375 185
R17968 vdd.n3430 vdd.n374 185
R17969 vdd.n3461 vdd.n374 185
R17970 vdd.n623 vdd.n373 185
R17971 vdd.n3462 vdd.n373 185
R17972 vdd.n3426 vdd.n372 185
R17973 vdd.n3463 vdd.n372 185
R17974 vdd.n3425 vdd.n3424 185
R17975 vdd.n3424 vdd.n3423 185
R17976 vdd.n3422 vdd.n364 185
R17977 vdd.n3469 vdd.n364 185
R17978 vdd.n625 vdd.n363 185
R17979 vdd.n3470 vdd.n363 185
R17980 vdd.n3418 vdd.n362 185
R17981 vdd.n3471 vdd.n362 185
R17982 vdd.n3417 vdd.n3416 185
R17983 vdd.n3416 vdd.n361 185
R17984 vdd.n3415 vdd.n353 185
R17985 vdd.n3477 vdd.n353 185
R17986 vdd.n627 vdd.n352 185
R17987 vdd.n3478 vdd.n352 185
R17988 vdd.n3411 vdd.n351 185
R17989 vdd.n3479 vdd.n351 185
R17990 vdd.n3410 vdd.n3409 185
R17991 vdd.n3409 vdd.n344 185
R17992 vdd.n3408 vdd.n343 185
R17993 vdd.n3485 vdd.n343 185
R17994 vdd.n629 vdd.n342 185
R17995 vdd.n3486 vdd.n342 185
R17996 vdd.n3404 vdd.n341 185
R17997 vdd.n3487 vdd.n341 185
R17998 vdd.n3403 vdd.n3402 185
R17999 vdd.n3402 vdd.n340 185
R18000 vdd.n3401 vdd.n631 185
R18001 vdd.n3401 vdd.n3400 185
R18002 vdd.n3389 vdd.n632 185
R18003 vdd.n633 vdd.n632 185
R18004 vdd.n3391 vdd.n3390 185
R18005 vdd.n3392 vdd.n3391 185
R18006 vdd.n640 vdd.n639 185
R18007 vdd.n644 vdd.n639 185
R18008 vdd.n3383 vdd.n3382 185
R18009 vdd.n3382 vdd.n3381 185
R18010 vdd.n643 vdd.n642 185
R18011 vdd.n3372 vdd.n643 185
R18012 vdd.n3371 vdd.n3370 185
R18013 vdd.n3373 vdd.n3371 185
R18014 vdd.n651 vdd.n650 185
R18015 vdd.n656 vdd.n650 185
R18016 vdd.n3366 vdd.n3365 185
R18017 vdd.n3365 vdd.n3364 185
R18018 vdd.n654 vdd.n653 185
R18019 vdd.n655 vdd.n654 185
R18020 vdd.n3355 vdd.n3354 185
R18021 vdd.n3356 vdd.n3355 185
R18022 vdd.n664 vdd.n663 185
R18023 vdd.n663 vdd.n662 185
R18024 vdd.n3350 vdd.n3349 185
R18025 vdd.n3349 vdd.n3348 185
R18026 vdd.n667 vdd.n666 185
R18027 vdd.n3339 vdd.n667 185
R18028 vdd.n3338 vdd.n3337 185
R18029 vdd.n3340 vdd.n3338 185
R18030 vdd.n674 vdd.n673 185
R18031 vdd.n679 vdd.n673 185
R18032 vdd.n3333 vdd.n3332 185
R18033 vdd.n3332 vdd.n3331 185
R18034 vdd.n677 vdd.n676 185
R18035 vdd.n678 vdd.n677 185
R18036 vdd.n3322 vdd.n3321 185
R18037 vdd.n3323 vdd.n3322 185
R18038 vdd.n686 vdd.n685 185
R18039 vdd.n723 vdd.n685 185
R18040 vdd.n2936 vdd.n2935 185
R18041 vdd.n2934 vdd.n2700 185
R18042 vdd.n2933 vdd.n2699 185
R18043 vdd.n2938 vdd.n2699 185
R18044 vdd.n2932 vdd.n2931 185
R18045 vdd.n2930 vdd.n2929 185
R18046 vdd.n2928 vdd.n2927 185
R18047 vdd.n2926 vdd.n2925 185
R18048 vdd.n2924 vdd.n2923 185
R18049 vdd.n2922 vdd.n2921 185
R18050 vdd.n2920 vdd.n2919 185
R18051 vdd.n2918 vdd.n2917 185
R18052 vdd.n2916 vdd.n2915 185
R18053 vdd.n2914 vdd.n2913 185
R18054 vdd.n2912 vdd.n2911 185
R18055 vdd.n2910 vdd.n2909 185
R18056 vdd.n2908 vdd.n2907 185
R18057 vdd.n2906 vdd.n2905 185
R18058 vdd.n2904 vdd.n2903 185
R18059 vdd.n2902 vdd.n2901 185
R18060 vdd.n2900 vdd.n2899 185
R18061 vdd.n2898 vdd.n2897 185
R18062 vdd.n2896 vdd.n2895 185
R18063 vdd.n2894 vdd.n2893 185
R18064 vdd.n2892 vdd.n2891 185
R18065 vdd.n2890 vdd.n2889 185
R18066 vdd.n2888 vdd.n2887 185
R18067 vdd.n2886 vdd.n2885 185
R18068 vdd.n2884 vdd.n2883 185
R18069 vdd.n2882 vdd.n2881 185
R18070 vdd.n2880 vdd.n2879 185
R18071 vdd.n2878 vdd.n2877 185
R18072 vdd.n2876 vdd.n2875 185
R18073 vdd.n2873 vdd.n2872 185
R18074 vdd.n2871 vdd.n2870 185
R18075 vdd.n2869 vdd.n2868 185
R18076 vdd.n3087 vdd.n3086 185
R18077 vdd.n3089 vdd.n834 185
R18078 vdd.n3091 vdd.n3090 185
R18079 vdd.n3093 vdd.n831 185
R18080 vdd.n3095 vdd.n3094 185
R18081 vdd.n3097 vdd.n829 185
R18082 vdd.n3099 vdd.n3098 185
R18083 vdd.n3100 vdd.n828 185
R18084 vdd.n3102 vdd.n3101 185
R18085 vdd.n3104 vdd.n826 185
R18086 vdd.n3106 vdd.n3105 185
R18087 vdd.n3107 vdd.n825 185
R18088 vdd.n3109 vdd.n3108 185
R18089 vdd.n3111 vdd.n823 185
R18090 vdd.n3113 vdd.n3112 185
R18091 vdd.n3114 vdd.n822 185
R18092 vdd.n3116 vdd.n3115 185
R18093 vdd.n3118 vdd.n731 185
R18094 vdd.n3120 vdd.n3119 185
R18095 vdd.n3122 vdd.n820 185
R18096 vdd.n3124 vdd.n3123 185
R18097 vdd.n3125 vdd.n819 185
R18098 vdd.n3127 vdd.n3126 185
R18099 vdd.n3129 vdd.n817 185
R18100 vdd.n3131 vdd.n3130 185
R18101 vdd.n3132 vdd.n816 185
R18102 vdd.n3134 vdd.n3133 185
R18103 vdd.n3136 vdd.n814 185
R18104 vdd.n3138 vdd.n3137 185
R18105 vdd.n3139 vdd.n813 185
R18106 vdd.n3141 vdd.n3140 185
R18107 vdd.n3143 vdd.n812 185
R18108 vdd.n3144 vdd.n811 185
R18109 vdd.n3147 vdd.n3146 185
R18110 vdd.n3148 vdd.n809 185
R18111 vdd.n809 vdd.n692 185
R18112 vdd.n3085 vdd.n806 185
R18113 vdd.n3151 vdd.n806 185
R18114 vdd.n3084 vdd.n3083 185
R18115 vdd.n3083 vdd.n805 185
R18116 vdd.n3082 vdd.n836 185
R18117 vdd.n3082 vdd.n3081 185
R18118 vdd.n2816 vdd.n837 185
R18119 vdd.n846 vdd.n837 185
R18120 vdd.n2817 vdd.n844 185
R18121 vdd.n3075 vdd.n844 185
R18122 vdd.n2819 vdd.n2818 185
R18123 vdd.n2818 vdd.n843 185
R18124 vdd.n2820 vdd.n852 185
R18125 vdd.n3024 vdd.n852 185
R18126 vdd.n2822 vdd.n2821 185
R18127 vdd.n2821 vdd.n851 185
R18128 vdd.n2823 vdd.n858 185
R18129 vdd.n3018 vdd.n858 185
R18130 vdd.n2825 vdd.n2824 185
R18131 vdd.n2824 vdd.n857 185
R18132 vdd.n2826 vdd.n863 185
R18133 vdd.n3012 vdd.n863 185
R18134 vdd.n2828 vdd.n2827 185
R18135 vdd.n2827 vdd.n870 185
R18136 vdd.n2829 vdd.n868 185
R18137 vdd.n3006 vdd.n868 185
R18138 vdd.n2831 vdd.n2830 185
R18139 vdd.n2830 vdd.n878 185
R18140 vdd.n2832 vdd.n876 185
R18141 vdd.n2999 vdd.n876 185
R18142 vdd.n2834 vdd.n2833 185
R18143 vdd.n2833 vdd.n875 185
R18144 vdd.n2835 vdd.n883 185
R18145 vdd.n2993 vdd.n883 185
R18146 vdd.n2837 vdd.n2836 185
R18147 vdd.n2836 vdd.n882 185
R18148 vdd.n2838 vdd.n888 185
R18149 vdd.n2987 vdd.n888 185
R18150 vdd.n2840 vdd.n2839 185
R18151 vdd.n2839 vdd.n895 185
R18152 vdd.n2841 vdd.n893 185
R18153 vdd.n2981 vdd.n893 185
R18154 vdd.n2843 vdd.n2842 185
R18155 vdd.n2842 vdd.n901 185
R18156 vdd.n2844 vdd.n899 185
R18157 vdd.n2975 vdd.n899 185
R18158 vdd.n2846 vdd.n2845 185
R18159 vdd.n2847 vdd.n2846 185
R18160 vdd.n2815 vdd.n906 185
R18161 vdd.n2969 vdd.n906 185
R18162 vdd.n2814 vdd.n2813 185
R18163 vdd.n2813 vdd.n905 185
R18164 vdd.n2812 vdd.n912 185
R18165 vdd.n2963 vdd.n912 185
R18166 vdd.n2811 vdd.n2810 185
R18167 vdd.n2810 vdd.n911 185
R18168 vdd.n2809 vdd.n918 185
R18169 vdd.n2957 vdd.n918 185
R18170 vdd.n2808 vdd.n2807 185
R18171 vdd.n2807 vdd.n917 185
R18172 vdd.n2703 vdd.n923 185
R18173 vdd.n2951 vdd.n923 185
R18174 vdd.n2864 vdd.n2863 185
R18175 vdd.n2863 vdd.n2862 185
R18176 vdd.n2865 vdd.n929 185
R18177 vdd.n2945 vdd.n929 185
R18178 vdd.n2867 vdd.n2866 185
R18179 vdd.n2867 vdd.n928 185
R18180 vdd.n927 vdd.n926 185
R18181 vdd.n928 vdd.n927 185
R18182 vdd.n2947 vdd.n2946 185
R18183 vdd.n2946 vdd.n2945 185
R18184 vdd.n2948 vdd.n925 185
R18185 vdd.n2862 vdd.n925 185
R18186 vdd.n2950 vdd.n2949 185
R18187 vdd.n2951 vdd.n2950 185
R18188 vdd.n916 vdd.n915 185
R18189 vdd.n917 vdd.n916 185
R18190 vdd.n2959 vdd.n2958 185
R18191 vdd.n2958 vdd.n2957 185
R18192 vdd.n2960 vdd.n914 185
R18193 vdd.n914 vdd.n911 185
R18194 vdd.n2962 vdd.n2961 185
R18195 vdd.n2963 vdd.n2962 185
R18196 vdd.n904 vdd.n903 185
R18197 vdd.n905 vdd.n904 185
R18198 vdd.n2971 vdd.n2970 185
R18199 vdd.n2970 vdd.n2969 185
R18200 vdd.n2972 vdd.n902 185
R18201 vdd.n2847 vdd.n902 185
R18202 vdd.n2974 vdd.n2973 185
R18203 vdd.n2975 vdd.n2974 185
R18204 vdd.n892 vdd.n891 185
R18205 vdd.n901 vdd.n892 185
R18206 vdd.n2983 vdd.n2982 185
R18207 vdd.n2982 vdd.n2981 185
R18208 vdd.n2984 vdd.n890 185
R18209 vdd.n895 vdd.n890 185
R18210 vdd.n2986 vdd.n2985 185
R18211 vdd.n2987 vdd.n2986 185
R18212 vdd.n881 vdd.n880 185
R18213 vdd.n882 vdd.n881 185
R18214 vdd.n2995 vdd.n2994 185
R18215 vdd.n2994 vdd.n2993 185
R18216 vdd.n2996 vdd.n879 185
R18217 vdd.n879 vdd.n875 185
R18218 vdd.n2998 vdd.n2997 185
R18219 vdd.n2999 vdd.n2998 185
R18220 vdd.n867 vdd.n866 185
R18221 vdd.n878 vdd.n867 185
R18222 vdd.n3008 vdd.n3007 185
R18223 vdd.n3007 vdd.n3006 185
R18224 vdd.n3009 vdd.n865 185
R18225 vdd.n870 vdd.n865 185
R18226 vdd.n3011 vdd.n3010 185
R18227 vdd.n3012 vdd.n3011 185
R18228 vdd.n856 vdd.n855 185
R18229 vdd.n857 vdd.n856 185
R18230 vdd.n3020 vdd.n3019 185
R18231 vdd.n3019 vdd.n3018 185
R18232 vdd.n3021 vdd.n854 185
R18233 vdd.n854 vdd.n851 185
R18234 vdd.n3023 vdd.n3022 185
R18235 vdd.n3024 vdd.n3023 185
R18236 vdd.n842 vdd.n841 185
R18237 vdd.n843 vdd.n842 185
R18238 vdd.n3077 vdd.n3076 185
R18239 vdd.n3076 vdd.n3075 185
R18240 vdd.n3078 vdd.n840 185
R18241 vdd.n846 vdd.n840 185
R18242 vdd.n3080 vdd.n3079 185
R18243 vdd.n3081 vdd.n3080 185
R18244 vdd.n810 vdd.n808 185
R18245 vdd.n808 vdd.n805 185
R18246 vdd.n3150 vdd.n3149 185
R18247 vdd.n3151 vdd.n3150 185
R18248 vdd.n2592 vdd.n2591 185
R18249 vdd.n2593 vdd.n2592 185
R18250 vdd.n980 vdd.n978 185
R18251 vdd.n978 vdd.n976 185
R18252 vdd.n2507 vdd.n987 185
R18253 vdd.n2518 vdd.n987 185
R18254 vdd.n2508 vdd.n996 185
R18255 vdd.n1338 vdd.n996 185
R18256 vdd.n2510 vdd.n2509 185
R18257 vdd.n2511 vdd.n2510 185
R18258 vdd.n2506 vdd.n995 185
R18259 vdd.n995 vdd.n992 185
R18260 vdd.n2505 vdd.n2504 185
R18261 vdd.n2504 vdd.n2503 185
R18262 vdd.n998 vdd.n997 185
R18263 vdd.n999 vdd.n998 185
R18264 vdd.n2496 vdd.n2495 185
R18265 vdd.n2497 vdd.n2496 185
R18266 vdd.n2494 vdd.n1008 185
R18267 vdd.n1008 vdd.n1005 185
R18268 vdd.n2493 vdd.n2492 185
R18269 vdd.n2492 vdd.n2491 185
R18270 vdd.n1010 vdd.n1009 185
R18271 vdd.n1018 vdd.n1010 185
R18272 vdd.n2484 vdd.n2483 185
R18273 vdd.n2485 vdd.n2484 185
R18274 vdd.n2482 vdd.n1019 185
R18275 vdd.n1024 vdd.n1019 185
R18276 vdd.n2481 vdd.n2480 185
R18277 vdd.n2480 vdd.n2479 185
R18278 vdd.n1021 vdd.n1020 185
R18279 vdd.n1359 vdd.n1021 185
R18280 vdd.n2472 vdd.n2471 185
R18281 vdd.n2473 vdd.n2472 185
R18282 vdd.n2470 vdd.n1031 185
R18283 vdd.n1031 vdd.n1028 185
R18284 vdd.n2469 vdd.n2468 185
R18285 vdd.n2468 vdd.n2467 185
R18286 vdd.n1033 vdd.n1032 185
R18287 vdd.n1034 vdd.n1033 185
R18288 vdd.n2460 vdd.n2459 185
R18289 vdd.n2461 vdd.n2460 185
R18290 vdd.n2457 vdd.n1042 185
R18291 vdd.n1048 vdd.n1042 185
R18292 vdd.n2456 vdd.n2455 185
R18293 vdd.n2455 vdd.n2454 185
R18294 vdd.n1045 vdd.n1044 185
R18295 vdd.n1055 vdd.n1045 185
R18296 vdd.n2447 vdd.n2446 185
R18297 vdd.n2448 vdd.n2447 185
R18298 vdd.n2445 vdd.n1056 185
R18299 vdd.n1056 vdd.n1052 185
R18300 vdd.n2444 vdd.n2443 185
R18301 vdd.n2443 vdd.n2442 185
R18302 vdd.n1058 vdd.n1057 185
R18303 vdd.n1059 vdd.n1058 185
R18304 vdd.n2435 vdd.n2434 185
R18305 vdd.n2436 vdd.n2435 185
R18306 vdd.n2433 vdd.n1068 185
R18307 vdd.n1068 vdd.n1065 185
R18308 vdd.n2432 vdd.n2431 185
R18309 vdd.n2431 vdd.n2430 185
R18310 vdd.n1070 vdd.n1069 185
R18311 vdd.n1079 vdd.n1070 185
R18312 vdd.n2423 vdd.n2422 185
R18313 vdd.n2424 vdd.n2423 185
R18314 vdd.n2421 vdd.n1080 185
R18315 vdd.n1080 vdd.n1076 185
R18316 vdd.n2523 vdd.n951 185
R18317 vdd.n2665 vdd.n951 185
R18318 vdd.n2525 vdd.n2524 185
R18319 vdd.n2527 vdd.n2526 185
R18320 vdd.n2529 vdd.n2528 185
R18321 vdd.n2531 vdd.n2530 185
R18322 vdd.n2533 vdd.n2532 185
R18323 vdd.n2535 vdd.n2534 185
R18324 vdd.n2537 vdd.n2536 185
R18325 vdd.n2539 vdd.n2538 185
R18326 vdd.n2541 vdd.n2540 185
R18327 vdd.n2543 vdd.n2542 185
R18328 vdd.n2545 vdd.n2544 185
R18329 vdd.n2547 vdd.n2546 185
R18330 vdd.n2549 vdd.n2548 185
R18331 vdd.n2551 vdd.n2550 185
R18332 vdd.n2553 vdd.n2552 185
R18333 vdd.n2555 vdd.n2554 185
R18334 vdd.n2557 vdd.n2556 185
R18335 vdd.n2559 vdd.n2558 185
R18336 vdd.n2561 vdd.n2560 185
R18337 vdd.n2563 vdd.n2562 185
R18338 vdd.n2565 vdd.n2564 185
R18339 vdd.n2567 vdd.n2566 185
R18340 vdd.n2569 vdd.n2568 185
R18341 vdd.n2571 vdd.n2570 185
R18342 vdd.n2573 vdd.n2572 185
R18343 vdd.n2575 vdd.n2574 185
R18344 vdd.n2577 vdd.n2576 185
R18345 vdd.n2579 vdd.n2578 185
R18346 vdd.n2581 vdd.n2580 185
R18347 vdd.n2583 vdd.n2582 185
R18348 vdd.n2585 vdd.n2584 185
R18349 vdd.n2587 vdd.n2586 185
R18350 vdd.n2589 vdd.n2588 185
R18351 vdd.n2590 vdd.n979 185
R18352 vdd.n2522 vdd.n977 185
R18353 vdd.n2593 vdd.n977 185
R18354 vdd.n2521 vdd.n2520 185
R18355 vdd.n2520 vdd.n976 185
R18356 vdd.n2519 vdd.n984 185
R18357 vdd.n2519 vdd.n2518 185
R18358 vdd.n1256 vdd.n985 185
R18359 vdd.n1338 vdd.n985 185
R18360 vdd.n1257 vdd.n994 185
R18361 vdd.n2511 vdd.n994 185
R18362 vdd.n1259 vdd.n1258 185
R18363 vdd.n1258 vdd.n992 185
R18364 vdd.n1260 vdd.n1001 185
R18365 vdd.n2503 vdd.n1001 185
R18366 vdd.n1262 vdd.n1261 185
R18367 vdd.n1261 vdd.n999 185
R18368 vdd.n1263 vdd.n1007 185
R18369 vdd.n2497 vdd.n1007 185
R18370 vdd.n1265 vdd.n1264 185
R18371 vdd.n1264 vdd.n1005 185
R18372 vdd.n1266 vdd.n1012 185
R18373 vdd.n2491 vdd.n1012 185
R18374 vdd.n1268 vdd.n1267 185
R18375 vdd.n1267 vdd.n1018 185
R18376 vdd.n1269 vdd.n1017 185
R18377 vdd.n2485 vdd.n1017 185
R18378 vdd.n1271 vdd.n1270 185
R18379 vdd.n1270 vdd.n1024 185
R18380 vdd.n1272 vdd.n1023 185
R18381 vdd.n2479 vdd.n1023 185
R18382 vdd.n1361 vdd.n1360 185
R18383 vdd.n1360 vdd.n1359 185
R18384 vdd.n1362 vdd.n1030 185
R18385 vdd.n2473 vdd.n1030 185
R18386 vdd.n1364 vdd.n1363 185
R18387 vdd.n1363 vdd.n1028 185
R18388 vdd.n1365 vdd.n1036 185
R18389 vdd.n2467 vdd.n1036 185
R18390 vdd.n1367 vdd.n1366 185
R18391 vdd.n1366 vdd.n1034 185
R18392 vdd.n1368 vdd.n1041 185
R18393 vdd.n2461 vdd.n1041 185
R18394 vdd.n1370 vdd.n1369 185
R18395 vdd.n1369 vdd.n1048 185
R18396 vdd.n1371 vdd.n1047 185
R18397 vdd.n2454 vdd.n1047 185
R18398 vdd.n1373 vdd.n1372 185
R18399 vdd.n1372 vdd.n1055 185
R18400 vdd.n1374 vdd.n1054 185
R18401 vdd.n2448 vdd.n1054 185
R18402 vdd.n1376 vdd.n1375 185
R18403 vdd.n1375 vdd.n1052 185
R18404 vdd.n1377 vdd.n1061 185
R18405 vdd.n2442 vdd.n1061 185
R18406 vdd.n1379 vdd.n1378 185
R18407 vdd.n1378 vdd.n1059 185
R18408 vdd.n1380 vdd.n1067 185
R18409 vdd.n2436 vdd.n1067 185
R18410 vdd.n1382 vdd.n1381 185
R18411 vdd.n1381 vdd.n1065 185
R18412 vdd.n1383 vdd.n1072 185
R18413 vdd.n2430 vdd.n1072 185
R18414 vdd.n1385 vdd.n1384 185
R18415 vdd.n1384 vdd.n1079 185
R18416 vdd.n1386 vdd.n1078 185
R18417 vdd.n2424 vdd.n1078 185
R18418 vdd.n1388 vdd.n1387 185
R18419 vdd.n1387 vdd.n1076 185
R18420 vdd.n2420 vdd.n2419 185
R18421 vdd.n1082 vdd.n1081 185
R18422 vdd.n1223 vdd.n1222 185
R18423 vdd.n1225 vdd.n1224 185
R18424 vdd.n1227 vdd.n1226 185
R18425 vdd.n1229 vdd.n1228 185
R18426 vdd.n1231 vdd.n1230 185
R18427 vdd.n1233 vdd.n1232 185
R18428 vdd.n1235 vdd.n1234 185
R18429 vdd.n1237 vdd.n1236 185
R18430 vdd.n1239 vdd.n1238 185
R18431 vdd.n1241 vdd.n1240 185
R18432 vdd.n1243 vdd.n1242 185
R18433 vdd.n1245 vdd.n1244 185
R18434 vdd.n1247 vdd.n1246 185
R18435 vdd.n1249 vdd.n1248 185
R18436 vdd.n1251 vdd.n1250 185
R18437 vdd.n1422 vdd.n1252 185
R18438 vdd.n1421 vdd.n1420 185
R18439 vdd.n1419 vdd.n1418 185
R18440 vdd.n1417 vdd.n1416 185
R18441 vdd.n1415 vdd.n1414 185
R18442 vdd.n1413 vdd.n1412 185
R18443 vdd.n1411 vdd.n1410 185
R18444 vdd.n1409 vdd.n1408 185
R18445 vdd.n1407 vdd.n1406 185
R18446 vdd.n1405 vdd.n1404 185
R18447 vdd.n1403 vdd.n1402 185
R18448 vdd.n1401 vdd.n1400 185
R18449 vdd.n1399 vdd.n1398 185
R18450 vdd.n1397 vdd.n1396 185
R18451 vdd.n1395 vdd.n1394 185
R18452 vdd.n1393 vdd.n1392 185
R18453 vdd.n1391 vdd.n1390 185
R18454 vdd.n1389 vdd.n1116 185
R18455 vdd.n2417 vdd.n1116 185
R18456 vdd.n2417 vdd.n1083 179.345
R18457 vdd.n3315 vdd.n692 179.345
R18458 vdd.n327 vdd.n326 171.744
R18459 vdd.n326 vdd.n325 171.744
R18460 vdd.n325 vdd.n294 171.744
R18461 vdd.n318 vdd.n294 171.744
R18462 vdd.n318 vdd.n317 171.744
R18463 vdd.n317 vdd.n299 171.744
R18464 vdd.n310 vdd.n299 171.744
R18465 vdd.n310 vdd.n309 171.744
R18466 vdd.n309 vdd.n303 171.744
R18467 vdd.n268 vdd.n267 171.744
R18468 vdd.n267 vdd.n266 171.744
R18469 vdd.n266 vdd.n235 171.744
R18470 vdd.n259 vdd.n235 171.744
R18471 vdd.n259 vdd.n258 171.744
R18472 vdd.n258 vdd.n240 171.744
R18473 vdd.n251 vdd.n240 171.744
R18474 vdd.n251 vdd.n250 171.744
R18475 vdd.n250 vdd.n244 171.744
R18476 vdd.n225 vdd.n224 171.744
R18477 vdd.n224 vdd.n223 171.744
R18478 vdd.n223 vdd.n192 171.744
R18479 vdd.n216 vdd.n192 171.744
R18480 vdd.n216 vdd.n215 171.744
R18481 vdd.n215 vdd.n197 171.744
R18482 vdd.n208 vdd.n197 171.744
R18483 vdd.n208 vdd.n207 171.744
R18484 vdd.n207 vdd.n201 171.744
R18485 vdd.n166 vdd.n165 171.744
R18486 vdd.n165 vdd.n164 171.744
R18487 vdd.n164 vdd.n133 171.744
R18488 vdd.n157 vdd.n133 171.744
R18489 vdd.n157 vdd.n156 171.744
R18490 vdd.n156 vdd.n138 171.744
R18491 vdd.n149 vdd.n138 171.744
R18492 vdd.n149 vdd.n148 171.744
R18493 vdd.n148 vdd.n142 171.744
R18494 vdd.n124 vdd.n123 171.744
R18495 vdd.n123 vdd.n122 171.744
R18496 vdd.n122 vdd.n91 171.744
R18497 vdd.n115 vdd.n91 171.744
R18498 vdd.n115 vdd.n114 171.744
R18499 vdd.n114 vdd.n96 171.744
R18500 vdd.n107 vdd.n96 171.744
R18501 vdd.n107 vdd.n106 171.744
R18502 vdd.n106 vdd.n100 171.744
R18503 vdd.n65 vdd.n64 171.744
R18504 vdd.n64 vdd.n63 171.744
R18505 vdd.n63 vdd.n32 171.744
R18506 vdd.n56 vdd.n32 171.744
R18507 vdd.n56 vdd.n55 171.744
R18508 vdd.n55 vdd.n37 171.744
R18509 vdd.n48 vdd.n37 171.744
R18510 vdd.n48 vdd.n47 171.744
R18511 vdd.n47 vdd.n41 171.744
R18512 vdd.n2108 vdd.n2107 171.744
R18513 vdd.n2107 vdd.n2106 171.744
R18514 vdd.n2106 vdd.n2075 171.744
R18515 vdd.n2099 vdd.n2075 171.744
R18516 vdd.n2099 vdd.n2098 171.744
R18517 vdd.n2098 vdd.n2080 171.744
R18518 vdd.n2091 vdd.n2080 171.744
R18519 vdd.n2091 vdd.n2090 171.744
R18520 vdd.n2090 vdd.n2084 171.744
R18521 vdd.n2167 vdd.n2166 171.744
R18522 vdd.n2166 vdd.n2165 171.744
R18523 vdd.n2165 vdd.n2134 171.744
R18524 vdd.n2158 vdd.n2134 171.744
R18525 vdd.n2158 vdd.n2157 171.744
R18526 vdd.n2157 vdd.n2139 171.744
R18527 vdd.n2150 vdd.n2139 171.744
R18528 vdd.n2150 vdd.n2149 171.744
R18529 vdd.n2149 vdd.n2143 171.744
R18530 vdd.n2006 vdd.n2005 171.744
R18531 vdd.n2005 vdd.n2004 171.744
R18532 vdd.n2004 vdd.n1973 171.744
R18533 vdd.n1997 vdd.n1973 171.744
R18534 vdd.n1997 vdd.n1996 171.744
R18535 vdd.n1996 vdd.n1978 171.744
R18536 vdd.n1989 vdd.n1978 171.744
R18537 vdd.n1989 vdd.n1988 171.744
R18538 vdd.n1988 vdd.n1982 171.744
R18539 vdd.n2065 vdd.n2064 171.744
R18540 vdd.n2064 vdd.n2063 171.744
R18541 vdd.n2063 vdd.n2032 171.744
R18542 vdd.n2056 vdd.n2032 171.744
R18543 vdd.n2056 vdd.n2055 171.744
R18544 vdd.n2055 vdd.n2037 171.744
R18545 vdd.n2048 vdd.n2037 171.744
R18546 vdd.n2048 vdd.n2047 171.744
R18547 vdd.n2047 vdd.n2041 171.744
R18548 vdd.n1905 vdd.n1904 171.744
R18549 vdd.n1904 vdd.n1903 171.744
R18550 vdd.n1903 vdd.n1872 171.744
R18551 vdd.n1896 vdd.n1872 171.744
R18552 vdd.n1896 vdd.n1895 171.744
R18553 vdd.n1895 vdd.n1877 171.744
R18554 vdd.n1888 vdd.n1877 171.744
R18555 vdd.n1888 vdd.n1887 171.744
R18556 vdd.n1887 vdd.n1881 171.744
R18557 vdd.n1964 vdd.n1963 171.744
R18558 vdd.n1963 vdd.n1962 171.744
R18559 vdd.n1962 vdd.n1931 171.744
R18560 vdd.n1955 vdd.n1931 171.744
R18561 vdd.n1955 vdd.n1954 171.744
R18562 vdd.n1954 vdd.n1936 171.744
R18563 vdd.n1947 vdd.n1936 171.744
R18564 vdd.n1947 vdd.n1946 171.744
R18565 vdd.n1946 vdd.n1940 171.744
R18566 vdd.n468 vdd.n467 146.341
R18567 vdd.n474 vdd.n473 146.341
R18568 vdd.n478 vdd.n477 146.341
R18569 vdd.n484 vdd.n483 146.341
R18570 vdd.n488 vdd.n487 146.341
R18571 vdd.n494 vdd.n493 146.341
R18572 vdd.n498 vdd.n497 146.341
R18573 vdd.n504 vdd.n503 146.341
R18574 vdd.n508 vdd.n507 146.341
R18575 vdd.n514 vdd.n513 146.341
R18576 vdd.n518 vdd.n517 146.341
R18577 vdd.n524 vdd.n523 146.341
R18578 vdd.n528 vdd.n527 146.341
R18579 vdd.n534 vdd.n533 146.341
R18580 vdd.n538 vdd.n537 146.341
R18581 vdd.n544 vdd.n543 146.341
R18582 vdd.n548 vdd.n547 146.341
R18583 vdd.n554 vdd.n553 146.341
R18584 vdd.n558 vdd.n557 146.341
R18585 vdd.n564 vdd.n563 146.341
R18586 vdd.n568 vdd.n567 146.341
R18587 vdd.n574 vdd.n573 146.341
R18588 vdd.n578 vdd.n577 146.341
R18589 vdd.n584 vdd.n583 146.341
R18590 vdd.n588 vdd.n587 146.341
R18591 vdd.n594 vdd.n593 146.341
R18592 vdd.n598 vdd.n597 146.341
R18593 vdd.n604 vdd.n603 146.341
R18594 vdd.n608 vdd.n607 146.341
R18595 vdd.n614 vdd.n613 146.341
R18596 vdd.n616 vdd.n425 146.341
R18597 vdd.n3322 vdd.n685 146.341
R18598 vdd.n3322 vdd.n677 146.341
R18599 vdd.n3332 vdd.n677 146.341
R18600 vdd.n3332 vdd.n673 146.341
R18601 vdd.n3338 vdd.n673 146.341
R18602 vdd.n3338 vdd.n667 146.341
R18603 vdd.n3349 vdd.n667 146.341
R18604 vdd.n3349 vdd.n663 146.341
R18605 vdd.n3355 vdd.n663 146.341
R18606 vdd.n3355 vdd.n654 146.341
R18607 vdd.n3365 vdd.n654 146.341
R18608 vdd.n3365 vdd.n650 146.341
R18609 vdd.n3371 vdd.n650 146.341
R18610 vdd.n3371 vdd.n643 146.341
R18611 vdd.n3382 vdd.n643 146.341
R18612 vdd.n3382 vdd.n639 146.341
R18613 vdd.n3391 vdd.n639 146.341
R18614 vdd.n3391 vdd.n632 146.341
R18615 vdd.n3401 vdd.n632 146.341
R18616 vdd.n3402 vdd.n3401 146.341
R18617 vdd.n3402 vdd.n341 146.341
R18618 vdd.n342 vdd.n341 146.341
R18619 vdd.n343 vdd.n342 146.341
R18620 vdd.n3409 vdd.n343 146.341
R18621 vdd.n3409 vdd.n351 146.341
R18622 vdd.n352 vdd.n351 146.341
R18623 vdd.n353 vdd.n352 146.341
R18624 vdd.n3416 vdd.n353 146.341
R18625 vdd.n3416 vdd.n362 146.341
R18626 vdd.n363 vdd.n362 146.341
R18627 vdd.n364 vdd.n363 146.341
R18628 vdd.n3424 vdd.n364 146.341
R18629 vdd.n3424 vdd.n372 146.341
R18630 vdd.n373 vdd.n372 146.341
R18631 vdd.n374 vdd.n373 146.341
R18632 vdd.n3431 vdd.n374 146.341
R18633 vdd.n3431 vdd.n383 146.341
R18634 vdd.n384 vdd.n383 146.341
R18635 vdd.n385 vdd.n384 146.341
R18636 vdd.n3438 vdd.n385 146.341
R18637 vdd.n3438 vdd.n393 146.341
R18638 vdd.n725 vdd.n724 146.341
R18639 vdd.n728 vdd.n724 146.341
R18640 vdd.n734 vdd.n733 146.341
R18641 vdd.n3304 vdd.n3303 146.341
R18642 vdd.n3300 vdd.n3299 146.341
R18643 vdd.n3296 vdd.n3295 146.341
R18644 vdd.n3292 vdd.n3291 146.341
R18645 vdd.n3288 vdd.n3287 146.341
R18646 vdd.n3284 vdd.n3283 146.341
R18647 vdd.n3280 vdd.n3279 146.341
R18648 vdd.n3271 vdd.n3270 146.341
R18649 vdd.n3268 vdd.n3267 146.341
R18650 vdd.n3264 vdd.n3263 146.341
R18651 vdd.n3260 vdd.n3259 146.341
R18652 vdd.n3256 vdd.n3255 146.341
R18653 vdd.n3252 vdd.n3251 146.341
R18654 vdd.n3248 vdd.n3247 146.341
R18655 vdd.n3244 vdd.n3243 146.341
R18656 vdd.n3240 vdd.n3239 146.341
R18657 vdd.n3236 vdd.n3235 146.341
R18658 vdd.n3232 vdd.n3231 146.341
R18659 vdd.n3225 vdd.n3224 146.341
R18660 vdd.n3222 vdd.n3221 146.341
R18661 vdd.n3218 vdd.n3217 146.341
R18662 vdd.n3214 vdd.n3213 146.341
R18663 vdd.n3210 vdd.n3209 146.341
R18664 vdd.n3206 vdd.n3205 146.341
R18665 vdd.n3202 vdd.n3201 146.341
R18666 vdd.n3198 vdd.n3197 146.341
R18667 vdd.n3194 vdd.n3193 146.341
R18668 vdd.n3190 vdd.n3189 146.341
R18669 vdd.n3316 vdd.n691 146.341
R18670 vdd.n3324 vdd.n684 146.341
R18671 vdd.n3324 vdd.n680 146.341
R18672 vdd.n3330 vdd.n680 146.341
R18673 vdd.n3330 vdd.n672 146.341
R18674 vdd.n3341 vdd.n672 146.341
R18675 vdd.n3341 vdd.n668 146.341
R18676 vdd.n3347 vdd.n668 146.341
R18677 vdd.n3347 vdd.n661 146.341
R18678 vdd.n3357 vdd.n661 146.341
R18679 vdd.n3357 vdd.n657 146.341
R18680 vdd.n3363 vdd.n657 146.341
R18681 vdd.n3363 vdd.n649 146.341
R18682 vdd.n3374 vdd.n649 146.341
R18683 vdd.n3374 vdd.n645 146.341
R18684 vdd.n3380 vdd.n645 146.341
R18685 vdd.n3380 vdd.n638 146.341
R18686 vdd.n3393 vdd.n638 146.341
R18687 vdd.n3393 vdd.n634 146.341
R18688 vdd.n3399 vdd.n634 146.341
R18689 vdd.n3399 vdd.n338 146.341
R18690 vdd.n3488 vdd.n338 146.341
R18691 vdd.n3488 vdd.n339 146.341
R18692 vdd.n3484 vdd.n339 146.341
R18693 vdd.n3484 vdd.n345 146.341
R18694 vdd.n3480 vdd.n345 146.341
R18695 vdd.n3480 vdd.n350 146.341
R18696 vdd.n3476 vdd.n350 146.341
R18697 vdd.n3476 vdd.n354 146.341
R18698 vdd.n3472 vdd.n354 146.341
R18699 vdd.n3472 vdd.n360 146.341
R18700 vdd.n3468 vdd.n360 146.341
R18701 vdd.n3468 vdd.n365 146.341
R18702 vdd.n3464 vdd.n365 146.341
R18703 vdd.n3464 vdd.n371 146.341
R18704 vdd.n3460 vdd.n371 146.341
R18705 vdd.n3460 vdd.n376 146.341
R18706 vdd.n3456 vdd.n376 146.341
R18707 vdd.n3456 vdd.n382 146.341
R18708 vdd.n3452 vdd.n382 146.341
R18709 vdd.n3452 vdd.n387 146.341
R18710 vdd.n3448 vdd.n387 146.341
R18711 vdd.n2378 vdd.n2377 146.341
R18712 vdd.n2375 vdd.n2372 146.341
R18713 vdd.n2370 vdd.n1127 146.341
R18714 vdd.n2366 vdd.n2365 146.341
R18715 vdd.n2363 vdd.n1131 146.341
R18716 vdd.n2359 vdd.n2358 146.341
R18717 vdd.n2356 vdd.n1138 146.341
R18718 vdd.n2352 vdd.n2351 146.341
R18719 vdd.n2349 vdd.n1145 146.341
R18720 vdd.n1156 vdd.n1153 146.341
R18721 vdd.n2341 vdd.n2340 146.341
R18722 vdd.n2338 vdd.n1158 146.341
R18723 vdd.n2334 vdd.n2333 146.341
R18724 vdd.n2331 vdd.n1164 146.341
R18725 vdd.n2327 vdd.n2326 146.341
R18726 vdd.n2324 vdd.n1171 146.341
R18727 vdd.n2320 vdd.n2319 146.341
R18728 vdd.n2317 vdd.n1178 146.341
R18729 vdd.n2313 vdd.n2312 146.341
R18730 vdd.n2310 vdd.n1185 146.341
R18731 vdd.n1196 vdd.n1193 146.341
R18732 vdd.n2302 vdd.n2301 146.341
R18733 vdd.n2299 vdd.n1198 146.341
R18734 vdd.n2295 vdd.n2294 146.341
R18735 vdd.n2292 vdd.n1204 146.341
R18736 vdd.n2288 vdd.n2287 146.341
R18737 vdd.n2285 vdd.n1211 146.341
R18738 vdd.n2281 vdd.n2280 146.341
R18739 vdd.n2278 vdd.n1218 146.341
R18740 vdd.n1429 vdd.n1427 146.341
R18741 vdd.n1432 vdd.n1431 146.341
R18742 vdd.n1790 vdd.n1550 146.341
R18743 vdd.n1790 vdd.n1546 146.341
R18744 vdd.n1796 vdd.n1546 146.341
R18745 vdd.n1796 vdd.n1538 146.341
R18746 vdd.n1807 vdd.n1538 146.341
R18747 vdd.n1807 vdd.n1534 146.341
R18748 vdd.n1813 vdd.n1534 146.341
R18749 vdd.n1813 vdd.n1528 146.341
R18750 vdd.n1824 vdd.n1528 146.341
R18751 vdd.n1824 vdd.n1524 146.341
R18752 vdd.n1830 vdd.n1524 146.341
R18753 vdd.n1830 vdd.n1515 146.341
R18754 vdd.n1840 vdd.n1515 146.341
R18755 vdd.n1840 vdd.n1511 146.341
R18756 vdd.n1846 vdd.n1511 146.341
R18757 vdd.n1846 vdd.n1504 146.341
R18758 vdd.n1857 vdd.n1504 146.341
R18759 vdd.n1857 vdd.n1500 146.341
R18760 vdd.n1863 vdd.n1500 146.341
R18761 vdd.n1863 vdd.n1493 146.341
R18762 vdd.n2180 vdd.n1493 146.341
R18763 vdd.n2180 vdd.n1489 146.341
R18764 vdd.n2186 vdd.n1489 146.341
R18765 vdd.n2186 vdd.n1481 146.341
R18766 vdd.n2197 vdd.n1481 146.341
R18767 vdd.n2197 vdd.n1477 146.341
R18768 vdd.n2203 vdd.n1477 146.341
R18769 vdd.n2203 vdd.n1471 146.341
R18770 vdd.n2214 vdd.n1471 146.341
R18771 vdd.n2214 vdd.n1467 146.341
R18772 vdd.n2220 vdd.n1467 146.341
R18773 vdd.n2220 vdd.n1458 146.341
R18774 vdd.n2230 vdd.n1458 146.341
R18775 vdd.n2230 vdd.n1454 146.341
R18776 vdd.n2236 vdd.n1454 146.341
R18777 vdd.n2236 vdd.n1448 146.341
R18778 vdd.n2247 vdd.n1448 146.341
R18779 vdd.n2247 vdd.n1443 146.341
R18780 vdd.n2255 vdd.n1443 146.341
R18781 vdd.n2255 vdd.n1434 146.341
R18782 vdd.n2266 vdd.n1434 146.341
R18783 vdd.n1779 vdd.n1555 146.341
R18784 vdd.n1779 vdd.n1588 146.341
R18785 vdd.n1592 vdd.n1591 146.341
R18786 vdd.n1594 vdd.n1593 146.341
R18787 vdd.n1598 vdd.n1597 146.341
R18788 vdd.n1600 vdd.n1599 146.341
R18789 vdd.n1604 vdd.n1603 146.341
R18790 vdd.n1606 vdd.n1605 146.341
R18791 vdd.n1610 vdd.n1609 146.341
R18792 vdd.n1612 vdd.n1611 146.341
R18793 vdd.n1618 vdd.n1617 146.341
R18794 vdd.n1620 vdd.n1619 146.341
R18795 vdd.n1624 vdd.n1623 146.341
R18796 vdd.n1626 vdd.n1625 146.341
R18797 vdd.n1630 vdd.n1629 146.341
R18798 vdd.n1632 vdd.n1631 146.341
R18799 vdd.n1636 vdd.n1635 146.341
R18800 vdd.n1638 vdd.n1637 146.341
R18801 vdd.n1642 vdd.n1641 146.341
R18802 vdd.n1644 vdd.n1643 146.341
R18803 vdd.n1716 vdd.n1647 146.341
R18804 vdd.n1649 vdd.n1648 146.341
R18805 vdd.n1653 vdd.n1652 146.341
R18806 vdd.n1655 vdd.n1654 146.341
R18807 vdd.n1659 vdd.n1658 146.341
R18808 vdd.n1661 vdd.n1660 146.341
R18809 vdd.n1665 vdd.n1664 146.341
R18810 vdd.n1667 vdd.n1666 146.341
R18811 vdd.n1671 vdd.n1670 146.341
R18812 vdd.n1673 vdd.n1672 146.341
R18813 vdd.n1677 vdd.n1676 146.341
R18814 vdd.n1678 vdd.n1586 146.341
R18815 vdd.n1788 vdd.n1551 146.341
R18816 vdd.n1788 vdd.n1544 146.341
R18817 vdd.n1799 vdd.n1544 146.341
R18818 vdd.n1799 vdd.n1540 146.341
R18819 vdd.n1805 vdd.n1540 146.341
R18820 vdd.n1805 vdd.n1533 146.341
R18821 vdd.n1816 vdd.n1533 146.341
R18822 vdd.n1816 vdd.n1529 146.341
R18823 vdd.n1822 vdd.n1529 146.341
R18824 vdd.n1822 vdd.n1522 146.341
R18825 vdd.n1832 vdd.n1522 146.341
R18826 vdd.n1832 vdd.n1518 146.341
R18827 vdd.n1838 vdd.n1518 146.341
R18828 vdd.n1838 vdd.n1510 146.341
R18829 vdd.n1849 vdd.n1510 146.341
R18830 vdd.n1849 vdd.n1506 146.341
R18831 vdd.n1855 vdd.n1506 146.341
R18832 vdd.n1855 vdd.n1499 146.341
R18833 vdd.n1865 vdd.n1499 146.341
R18834 vdd.n1865 vdd.n1495 146.341
R18835 vdd.n2178 vdd.n1495 146.341
R18836 vdd.n2178 vdd.n1487 146.341
R18837 vdd.n2189 vdd.n1487 146.341
R18838 vdd.n2189 vdd.n1483 146.341
R18839 vdd.n2195 vdd.n1483 146.341
R18840 vdd.n2195 vdd.n1476 146.341
R18841 vdd.n2206 vdd.n1476 146.341
R18842 vdd.n2206 vdd.n1472 146.341
R18843 vdd.n2212 vdd.n1472 146.341
R18844 vdd.n2212 vdd.n1465 146.341
R18845 vdd.n2222 vdd.n1465 146.341
R18846 vdd.n2222 vdd.n1461 146.341
R18847 vdd.n2228 vdd.n1461 146.341
R18848 vdd.n2228 vdd.n1453 146.341
R18849 vdd.n2239 vdd.n1453 146.341
R18850 vdd.n2239 vdd.n1449 146.341
R18851 vdd.n2245 vdd.n1449 146.341
R18852 vdd.n2245 vdd.n1441 146.341
R18853 vdd.n2258 vdd.n1441 146.341
R18854 vdd.n2258 vdd.n1436 146.341
R18855 vdd.n2264 vdd.n1436 146.341
R18856 vdd.n1253 vdd.t33 127.284
R18857 vdd.n981 vdd.t74 127.284
R18858 vdd.n1273 vdd.t47 127.284
R18859 vdd.n972 vdd.t97 127.284
R18860 vdd.n872 vdd.t54 127.284
R18861 vdd.n872 vdd.t55 127.284
R18862 vdd.n2704 vdd.t89 127.284
R18863 vdd.n832 vdd.t100 127.284
R18864 vdd.n2701 vdd.t79 127.284
R18865 vdd.n799 vdd.t28 127.284
R18866 vdd.n1043 vdd.t85 127.284
R18867 vdd.n1043 vdd.t86 127.284
R18868 vdd.n22 vdd.n20 117.314
R18869 vdd.n17 vdd.n15 117.314
R18870 vdd.n27 vdd.n26 116.927
R18871 vdd.n24 vdd.n23 116.927
R18872 vdd.n22 vdd.n21 116.927
R18873 vdd.n17 vdd.n16 116.927
R18874 vdd.n19 vdd.n18 116.927
R18875 vdd.n27 vdd.n25 116.927
R18876 vdd.n1254 vdd.t32 111.188
R18877 vdd.n982 vdd.t75 111.188
R18878 vdd.n1274 vdd.t46 111.188
R18879 vdd.n973 vdd.t98 111.188
R18880 vdd.n2705 vdd.t88 111.188
R18881 vdd.n833 vdd.t101 111.188
R18882 vdd.n2702 vdd.t78 111.188
R18883 vdd.n800 vdd.t29 111.188
R18884 vdd.n2946 vdd.n927 99.5127
R18885 vdd.n2946 vdd.n925 99.5127
R18886 vdd.n2950 vdd.n925 99.5127
R18887 vdd.n2950 vdd.n916 99.5127
R18888 vdd.n2958 vdd.n916 99.5127
R18889 vdd.n2958 vdd.n914 99.5127
R18890 vdd.n2962 vdd.n914 99.5127
R18891 vdd.n2962 vdd.n904 99.5127
R18892 vdd.n2970 vdd.n904 99.5127
R18893 vdd.n2970 vdd.n902 99.5127
R18894 vdd.n2974 vdd.n902 99.5127
R18895 vdd.n2974 vdd.n892 99.5127
R18896 vdd.n2982 vdd.n892 99.5127
R18897 vdd.n2982 vdd.n890 99.5127
R18898 vdd.n2986 vdd.n890 99.5127
R18899 vdd.n2986 vdd.n881 99.5127
R18900 vdd.n2994 vdd.n881 99.5127
R18901 vdd.n2994 vdd.n879 99.5127
R18902 vdd.n2998 vdd.n879 99.5127
R18903 vdd.n2998 vdd.n867 99.5127
R18904 vdd.n3007 vdd.n867 99.5127
R18905 vdd.n3007 vdd.n865 99.5127
R18906 vdd.n3011 vdd.n865 99.5127
R18907 vdd.n3011 vdd.n856 99.5127
R18908 vdd.n3019 vdd.n856 99.5127
R18909 vdd.n3019 vdd.n854 99.5127
R18910 vdd.n3023 vdd.n854 99.5127
R18911 vdd.n3023 vdd.n842 99.5127
R18912 vdd.n3076 vdd.n842 99.5127
R18913 vdd.n3076 vdd.n840 99.5127
R18914 vdd.n3080 vdd.n840 99.5127
R18915 vdd.n3080 vdd.n808 99.5127
R18916 vdd.n3150 vdd.n808 99.5127
R18917 vdd.n3146 vdd.n809 99.5127
R18918 vdd.n3144 vdd.n3143 99.5127
R18919 vdd.n3141 vdd.n813 99.5127
R18920 vdd.n3137 vdd.n3136 99.5127
R18921 vdd.n3134 vdd.n816 99.5127
R18922 vdd.n3130 vdd.n3129 99.5127
R18923 vdd.n3127 vdd.n819 99.5127
R18924 vdd.n3123 vdd.n3122 99.5127
R18925 vdd.n3120 vdd.n3118 99.5127
R18926 vdd.n3116 vdd.n822 99.5127
R18927 vdd.n3112 vdd.n3111 99.5127
R18928 vdd.n3109 vdd.n825 99.5127
R18929 vdd.n3105 vdd.n3104 99.5127
R18930 vdd.n3102 vdd.n828 99.5127
R18931 vdd.n3098 vdd.n3097 99.5127
R18932 vdd.n3095 vdd.n831 99.5127
R18933 vdd.n3090 vdd.n3089 99.5127
R18934 vdd.n2867 vdd.n929 99.5127
R18935 vdd.n2863 vdd.n929 99.5127
R18936 vdd.n2863 vdd.n923 99.5127
R18937 vdd.n2807 vdd.n923 99.5127
R18938 vdd.n2807 vdd.n918 99.5127
R18939 vdd.n2810 vdd.n918 99.5127
R18940 vdd.n2810 vdd.n912 99.5127
R18941 vdd.n2813 vdd.n912 99.5127
R18942 vdd.n2813 vdd.n906 99.5127
R18943 vdd.n2846 vdd.n906 99.5127
R18944 vdd.n2846 vdd.n899 99.5127
R18945 vdd.n2842 vdd.n899 99.5127
R18946 vdd.n2842 vdd.n893 99.5127
R18947 vdd.n2839 vdd.n893 99.5127
R18948 vdd.n2839 vdd.n888 99.5127
R18949 vdd.n2836 vdd.n888 99.5127
R18950 vdd.n2836 vdd.n883 99.5127
R18951 vdd.n2833 vdd.n883 99.5127
R18952 vdd.n2833 vdd.n876 99.5127
R18953 vdd.n2830 vdd.n876 99.5127
R18954 vdd.n2830 vdd.n868 99.5127
R18955 vdd.n2827 vdd.n868 99.5127
R18956 vdd.n2827 vdd.n863 99.5127
R18957 vdd.n2824 vdd.n863 99.5127
R18958 vdd.n2824 vdd.n858 99.5127
R18959 vdd.n2821 vdd.n858 99.5127
R18960 vdd.n2821 vdd.n852 99.5127
R18961 vdd.n2818 vdd.n852 99.5127
R18962 vdd.n2818 vdd.n844 99.5127
R18963 vdd.n844 vdd.n837 99.5127
R18964 vdd.n3082 vdd.n837 99.5127
R18965 vdd.n3083 vdd.n3082 99.5127
R18966 vdd.n3083 vdd.n806 99.5127
R18967 vdd.n2700 vdd.n2699 99.5127
R18968 vdd.n2931 vdd.n2699 99.5127
R18969 vdd.n2929 vdd.n2928 99.5127
R18970 vdd.n2925 vdd.n2924 99.5127
R18971 vdd.n2921 vdd.n2920 99.5127
R18972 vdd.n2917 vdd.n2916 99.5127
R18973 vdd.n2913 vdd.n2912 99.5127
R18974 vdd.n2909 vdd.n2908 99.5127
R18975 vdd.n2905 vdd.n2904 99.5127
R18976 vdd.n2901 vdd.n2900 99.5127
R18977 vdd.n2897 vdd.n2896 99.5127
R18978 vdd.n2893 vdd.n2892 99.5127
R18979 vdd.n2889 vdd.n2888 99.5127
R18980 vdd.n2885 vdd.n2884 99.5127
R18981 vdd.n2881 vdd.n2880 99.5127
R18982 vdd.n2877 vdd.n2876 99.5127
R18983 vdd.n2872 vdd.n2871 99.5127
R18984 vdd.n2664 vdd.n970 99.5127
R18985 vdd.n2660 vdd.n2659 99.5127
R18986 vdd.n2656 vdd.n2655 99.5127
R18987 vdd.n2652 vdd.n2651 99.5127
R18988 vdd.n2648 vdd.n2647 99.5127
R18989 vdd.n2644 vdd.n2643 99.5127
R18990 vdd.n2640 vdd.n2639 99.5127
R18991 vdd.n2636 vdd.n2635 99.5127
R18992 vdd.n2632 vdd.n2631 99.5127
R18993 vdd.n2628 vdd.n2627 99.5127
R18994 vdd.n2624 vdd.n2623 99.5127
R18995 vdd.n2620 vdd.n2619 99.5127
R18996 vdd.n2616 vdd.n2615 99.5127
R18997 vdd.n2612 vdd.n2611 99.5127
R18998 vdd.n2608 vdd.n2607 99.5127
R18999 vdd.n2604 vdd.n2603 99.5127
R19000 vdd.n2599 vdd.n2598 99.5127
R19001 vdd.n1309 vdd.n1077 99.5127
R19002 vdd.n1312 vdd.n1077 99.5127
R19003 vdd.n1312 vdd.n1071 99.5127
R19004 vdd.n1315 vdd.n1071 99.5127
R19005 vdd.n1315 vdd.n1066 99.5127
R19006 vdd.n1318 vdd.n1066 99.5127
R19007 vdd.n1318 vdd.n1060 99.5127
R19008 vdd.n1321 vdd.n1060 99.5127
R19009 vdd.n1321 vdd.n1053 99.5127
R19010 vdd.n1324 vdd.n1053 99.5127
R19011 vdd.n1324 vdd.n1046 99.5127
R19012 vdd.n1327 vdd.n1046 99.5127
R19013 vdd.n1327 vdd.n1040 99.5127
R19014 vdd.n1330 vdd.n1040 99.5127
R19015 vdd.n1330 vdd.n1035 99.5127
R19016 vdd.n1333 vdd.n1035 99.5127
R19017 vdd.n1333 vdd.n1029 99.5127
R19018 vdd.n1358 vdd.n1029 99.5127
R19019 vdd.n1358 vdd.n1022 99.5127
R19020 vdd.n1354 vdd.n1022 99.5127
R19021 vdd.n1354 vdd.n1016 99.5127
R19022 vdd.n1351 vdd.n1016 99.5127
R19023 vdd.n1351 vdd.n1011 99.5127
R19024 vdd.n1348 vdd.n1011 99.5127
R19025 vdd.n1348 vdd.n1006 99.5127
R19026 vdd.n1345 vdd.n1006 99.5127
R19027 vdd.n1345 vdd.n1000 99.5127
R19028 vdd.n1342 vdd.n1000 99.5127
R19029 vdd.n1342 vdd.n993 99.5127
R19030 vdd.n1339 vdd.n993 99.5127
R19031 vdd.n1339 vdd.n986 99.5127
R19032 vdd.n986 vdd.n975 99.5127
R19033 vdd.n2594 vdd.n975 99.5127
R19034 vdd.n1118 vdd.n1117 99.5127
R19035 vdd.n2410 vdd.n1117 99.5127
R19036 vdd.n2408 vdd.n2407 99.5127
R19037 vdd.n2404 vdd.n2403 99.5127
R19038 vdd.n2400 vdd.n2399 99.5127
R19039 vdd.n2396 vdd.n2395 99.5127
R19040 vdd.n2392 vdd.n2391 99.5127
R19041 vdd.n2388 vdd.n2387 99.5127
R19042 vdd.n2384 vdd.n2383 99.5127
R19043 vdd.n1276 vdd.n1275 99.5127
R19044 vdd.n1280 vdd.n1279 99.5127
R19045 vdd.n1284 vdd.n1283 99.5127
R19046 vdd.n1288 vdd.n1287 99.5127
R19047 vdd.n1292 vdd.n1291 99.5127
R19048 vdd.n1296 vdd.n1295 99.5127
R19049 vdd.n1300 vdd.n1299 99.5127
R19050 vdd.n1305 vdd.n1304 99.5127
R19051 vdd.n2425 vdd.n1075 99.5127
R19052 vdd.n2425 vdd.n1073 99.5127
R19053 vdd.n2429 vdd.n1073 99.5127
R19054 vdd.n2429 vdd.n1064 99.5127
R19055 vdd.n2437 vdd.n1064 99.5127
R19056 vdd.n2437 vdd.n1062 99.5127
R19057 vdd.n2441 vdd.n1062 99.5127
R19058 vdd.n2441 vdd.n1051 99.5127
R19059 vdd.n2449 vdd.n1051 99.5127
R19060 vdd.n2449 vdd.n1049 99.5127
R19061 vdd.n2453 vdd.n1049 99.5127
R19062 vdd.n2453 vdd.n1039 99.5127
R19063 vdd.n2462 vdd.n1039 99.5127
R19064 vdd.n2462 vdd.n1037 99.5127
R19065 vdd.n2466 vdd.n1037 99.5127
R19066 vdd.n2466 vdd.n1027 99.5127
R19067 vdd.n2474 vdd.n1027 99.5127
R19068 vdd.n2474 vdd.n1025 99.5127
R19069 vdd.n2478 vdd.n1025 99.5127
R19070 vdd.n2478 vdd.n1015 99.5127
R19071 vdd.n2486 vdd.n1015 99.5127
R19072 vdd.n2486 vdd.n1013 99.5127
R19073 vdd.n2490 vdd.n1013 99.5127
R19074 vdd.n2490 vdd.n1004 99.5127
R19075 vdd.n2498 vdd.n1004 99.5127
R19076 vdd.n2498 vdd.n1002 99.5127
R19077 vdd.n2502 vdd.n1002 99.5127
R19078 vdd.n2502 vdd.n991 99.5127
R19079 vdd.n2512 vdd.n991 99.5127
R19080 vdd.n2512 vdd.n988 99.5127
R19081 vdd.n2517 vdd.n988 99.5127
R19082 vdd.n2517 vdd.n989 99.5127
R19083 vdd.n989 vdd.n969 99.5127
R19084 vdd.n3066 vdd.n3065 99.5127
R19085 vdd.n3063 vdd.n3029 99.5127
R19086 vdd.n3059 vdd.n3058 99.5127
R19087 vdd.n3056 vdd.n3032 99.5127
R19088 vdd.n3052 vdd.n3051 99.5127
R19089 vdd.n3049 vdd.n3035 99.5127
R19090 vdd.n3045 vdd.n3044 99.5127
R19091 vdd.n3042 vdd.n3039 99.5127
R19092 vdd.n3183 vdd.n787 99.5127
R19093 vdd.n3181 vdd.n3180 99.5127
R19094 vdd.n3178 vdd.n789 99.5127
R19095 vdd.n3174 vdd.n3173 99.5127
R19096 vdd.n3171 vdd.n792 99.5127
R19097 vdd.n3167 vdd.n3166 99.5127
R19098 vdd.n3164 vdd.n795 99.5127
R19099 vdd.n3160 vdd.n3159 99.5127
R19100 vdd.n3157 vdd.n798 99.5127
R19101 vdd.n2772 vdd.n930 99.5127
R19102 vdd.n2861 vdd.n930 99.5127
R19103 vdd.n2861 vdd.n924 99.5127
R19104 vdd.n2857 vdd.n924 99.5127
R19105 vdd.n2857 vdd.n919 99.5127
R19106 vdd.n2854 vdd.n919 99.5127
R19107 vdd.n2854 vdd.n913 99.5127
R19108 vdd.n2851 vdd.n913 99.5127
R19109 vdd.n2851 vdd.n907 99.5127
R19110 vdd.n2848 vdd.n907 99.5127
R19111 vdd.n2848 vdd.n900 99.5127
R19112 vdd.n2804 vdd.n900 99.5127
R19113 vdd.n2804 vdd.n894 99.5127
R19114 vdd.n2801 vdd.n894 99.5127
R19115 vdd.n2801 vdd.n889 99.5127
R19116 vdd.n2798 vdd.n889 99.5127
R19117 vdd.n2798 vdd.n884 99.5127
R19118 vdd.n2795 vdd.n884 99.5127
R19119 vdd.n2795 vdd.n877 99.5127
R19120 vdd.n2792 vdd.n877 99.5127
R19121 vdd.n2792 vdd.n869 99.5127
R19122 vdd.n2789 vdd.n869 99.5127
R19123 vdd.n2789 vdd.n864 99.5127
R19124 vdd.n2786 vdd.n864 99.5127
R19125 vdd.n2786 vdd.n859 99.5127
R19126 vdd.n2783 vdd.n859 99.5127
R19127 vdd.n2783 vdd.n853 99.5127
R19128 vdd.n2780 vdd.n853 99.5127
R19129 vdd.n2780 vdd.n845 99.5127
R19130 vdd.n2777 vdd.n845 99.5127
R19131 vdd.n2777 vdd.n838 99.5127
R19132 vdd.n838 vdd.n804 99.5127
R19133 vdd.n3152 vdd.n804 99.5127
R19134 vdd.n2707 vdd.n933 99.5127
R19135 vdd.n2711 vdd.n2710 99.5127
R19136 vdd.n2715 vdd.n2714 99.5127
R19137 vdd.n2719 vdd.n2718 99.5127
R19138 vdd.n2723 vdd.n2722 99.5127
R19139 vdd.n2727 vdd.n2726 99.5127
R19140 vdd.n2731 vdd.n2730 99.5127
R19141 vdd.n2735 vdd.n2734 99.5127
R19142 vdd.n2739 vdd.n2738 99.5127
R19143 vdd.n2743 vdd.n2742 99.5127
R19144 vdd.n2747 vdd.n2746 99.5127
R19145 vdd.n2751 vdd.n2750 99.5127
R19146 vdd.n2755 vdd.n2754 99.5127
R19147 vdd.n2759 vdd.n2758 99.5127
R19148 vdd.n2763 vdd.n2762 99.5127
R19149 vdd.n2767 vdd.n2766 99.5127
R19150 vdd.n2769 vdd.n2698 99.5127
R19151 vdd.n2944 vdd.n931 99.5127
R19152 vdd.n2944 vdd.n922 99.5127
R19153 vdd.n2952 vdd.n922 99.5127
R19154 vdd.n2952 vdd.n920 99.5127
R19155 vdd.n2956 vdd.n920 99.5127
R19156 vdd.n2956 vdd.n910 99.5127
R19157 vdd.n2964 vdd.n910 99.5127
R19158 vdd.n2964 vdd.n908 99.5127
R19159 vdd.n2968 vdd.n908 99.5127
R19160 vdd.n2968 vdd.n898 99.5127
R19161 vdd.n2976 vdd.n898 99.5127
R19162 vdd.n2976 vdd.n896 99.5127
R19163 vdd.n2980 vdd.n896 99.5127
R19164 vdd.n2980 vdd.n887 99.5127
R19165 vdd.n2988 vdd.n887 99.5127
R19166 vdd.n2988 vdd.n885 99.5127
R19167 vdd.n2992 vdd.n885 99.5127
R19168 vdd.n2992 vdd.n874 99.5127
R19169 vdd.n3000 vdd.n874 99.5127
R19170 vdd.n3000 vdd.n871 99.5127
R19171 vdd.n3005 vdd.n871 99.5127
R19172 vdd.n3005 vdd.n862 99.5127
R19173 vdd.n3013 vdd.n862 99.5127
R19174 vdd.n3013 vdd.n860 99.5127
R19175 vdd.n3017 vdd.n860 99.5127
R19176 vdd.n3017 vdd.n850 99.5127
R19177 vdd.n3025 vdd.n850 99.5127
R19178 vdd.n3025 vdd.n847 99.5127
R19179 vdd.n3074 vdd.n847 99.5127
R19180 vdd.n3074 vdd.n848 99.5127
R19181 vdd.n848 vdd.n839 99.5127
R19182 vdd.n3069 vdd.n839 99.5127
R19183 vdd.n3069 vdd.n807 99.5127
R19184 vdd.n2588 vdd.n2587 99.5127
R19185 vdd.n2584 vdd.n2583 99.5127
R19186 vdd.n2580 vdd.n2579 99.5127
R19187 vdd.n2576 vdd.n2575 99.5127
R19188 vdd.n2572 vdd.n2571 99.5127
R19189 vdd.n2568 vdd.n2567 99.5127
R19190 vdd.n2564 vdd.n2563 99.5127
R19191 vdd.n2560 vdd.n2559 99.5127
R19192 vdd.n2556 vdd.n2555 99.5127
R19193 vdd.n2552 vdd.n2551 99.5127
R19194 vdd.n2548 vdd.n2547 99.5127
R19195 vdd.n2544 vdd.n2543 99.5127
R19196 vdd.n2540 vdd.n2539 99.5127
R19197 vdd.n2536 vdd.n2535 99.5127
R19198 vdd.n2532 vdd.n2531 99.5127
R19199 vdd.n2528 vdd.n2527 99.5127
R19200 vdd.n2524 vdd.n951 99.5127
R19201 vdd.n1387 vdd.n1078 99.5127
R19202 vdd.n1384 vdd.n1078 99.5127
R19203 vdd.n1384 vdd.n1072 99.5127
R19204 vdd.n1381 vdd.n1072 99.5127
R19205 vdd.n1381 vdd.n1067 99.5127
R19206 vdd.n1378 vdd.n1067 99.5127
R19207 vdd.n1378 vdd.n1061 99.5127
R19208 vdd.n1375 vdd.n1061 99.5127
R19209 vdd.n1375 vdd.n1054 99.5127
R19210 vdd.n1372 vdd.n1054 99.5127
R19211 vdd.n1372 vdd.n1047 99.5127
R19212 vdd.n1369 vdd.n1047 99.5127
R19213 vdd.n1369 vdd.n1041 99.5127
R19214 vdd.n1366 vdd.n1041 99.5127
R19215 vdd.n1366 vdd.n1036 99.5127
R19216 vdd.n1363 vdd.n1036 99.5127
R19217 vdd.n1363 vdd.n1030 99.5127
R19218 vdd.n1360 vdd.n1030 99.5127
R19219 vdd.n1360 vdd.n1023 99.5127
R19220 vdd.n1270 vdd.n1023 99.5127
R19221 vdd.n1270 vdd.n1017 99.5127
R19222 vdd.n1267 vdd.n1017 99.5127
R19223 vdd.n1267 vdd.n1012 99.5127
R19224 vdd.n1264 vdd.n1012 99.5127
R19225 vdd.n1264 vdd.n1007 99.5127
R19226 vdd.n1261 vdd.n1007 99.5127
R19227 vdd.n1261 vdd.n1001 99.5127
R19228 vdd.n1258 vdd.n1001 99.5127
R19229 vdd.n1258 vdd.n994 99.5127
R19230 vdd.n994 vdd.n985 99.5127
R19231 vdd.n2519 vdd.n985 99.5127
R19232 vdd.n2520 vdd.n2519 99.5127
R19233 vdd.n2520 vdd.n977 99.5127
R19234 vdd.n1222 vdd.n1082 99.5127
R19235 vdd.n1226 vdd.n1225 99.5127
R19236 vdd.n1230 vdd.n1229 99.5127
R19237 vdd.n1234 vdd.n1233 99.5127
R19238 vdd.n1238 vdd.n1237 99.5127
R19239 vdd.n1242 vdd.n1241 99.5127
R19240 vdd.n1246 vdd.n1245 99.5127
R19241 vdd.n1250 vdd.n1249 99.5127
R19242 vdd.n1420 vdd.n1252 99.5127
R19243 vdd.n1418 vdd.n1417 99.5127
R19244 vdd.n1414 vdd.n1413 99.5127
R19245 vdd.n1410 vdd.n1409 99.5127
R19246 vdd.n1406 vdd.n1405 99.5127
R19247 vdd.n1402 vdd.n1401 99.5127
R19248 vdd.n1398 vdd.n1397 99.5127
R19249 vdd.n1394 vdd.n1393 99.5127
R19250 vdd.n1390 vdd.n1116 99.5127
R19251 vdd.n2423 vdd.n1080 99.5127
R19252 vdd.n2423 vdd.n1070 99.5127
R19253 vdd.n2431 vdd.n1070 99.5127
R19254 vdd.n2431 vdd.n1068 99.5127
R19255 vdd.n2435 vdd.n1068 99.5127
R19256 vdd.n2435 vdd.n1058 99.5127
R19257 vdd.n2443 vdd.n1058 99.5127
R19258 vdd.n2443 vdd.n1056 99.5127
R19259 vdd.n2447 vdd.n1056 99.5127
R19260 vdd.n2447 vdd.n1045 99.5127
R19261 vdd.n2455 vdd.n1045 99.5127
R19262 vdd.n2455 vdd.n1042 99.5127
R19263 vdd.n2460 vdd.n1042 99.5127
R19264 vdd.n2460 vdd.n1033 99.5127
R19265 vdd.n2468 vdd.n1033 99.5127
R19266 vdd.n2468 vdd.n1031 99.5127
R19267 vdd.n2472 vdd.n1031 99.5127
R19268 vdd.n2472 vdd.n1021 99.5127
R19269 vdd.n2480 vdd.n1021 99.5127
R19270 vdd.n2480 vdd.n1019 99.5127
R19271 vdd.n2484 vdd.n1019 99.5127
R19272 vdd.n2484 vdd.n1010 99.5127
R19273 vdd.n2492 vdd.n1010 99.5127
R19274 vdd.n2492 vdd.n1008 99.5127
R19275 vdd.n2496 vdd.n1008 99.5127
R19276 vdd.n2496 vdd.n998 99.5127
R19277 vdd.n2504 vdd.n998 99.5127
R19278 vdd.n2504 vdd.n995 99.5127
R19279 vdd.n2510 vdd.n995 99.5127
R19280 vdd.n2510 vdd.n996 99.5127
R19281 vdd.n996 vdd.n987 99.5127
R19282 vdd.n987 vdd.n978 99.5127
R19283 vdd.n2592 vdd.n978 99.5127
R19284 vdd.n9 vdd.n7 98.9633
R19285 vdd.n2 vdd.n0 98.9633
R19286 vdd.n9 vdd.n8 98.6055
R19287 vdd.n11 vdd.n10 98.6055
R19288 vdd.n13 vdd.n12 98.6055
R19289 vdd.n6 vdd.n5 98.6055
R19290 vdd.n4 vdd.n3 98.6055
R19291 vdd.n2 vdd.n1 98.6055
R19292 vdd.t161 vdd.n303 85.8723
R19293 vdd.t246 vdd.n244 85.8723
R19294 vdd.t297 vdd.n201 85.8723
R19295 vdd.t230 vdd.n142 85.8723
R19296 vdd.t198 vdd.n100 85.8723
R19297 vdd.t187 vdd.n41 85.8723
R19298 vdd.t288 vdd.n2084 85.8723
R19299 vdd.t222 vdd.n2143 85.8723
R19300 vdd.t276 vdd.n1982 85.8723
R19301 vdd.t199 vdd.n2041 85.8723
R19302 vdd.t189 vdd.n1881 85.8723
R19303 vdd.t197 vdd.n1940 85.8723
R19304 vdd.n3003 vdd.n872 78.546
R19305 vdd.n2458 vdd.n1043 78.546
R19306 vdd.n290 vdd.n289 75.1835
R19307 vdd.n288 vdd.n287 75.1835
R19308 vdd.n286 vdd.n285 75.1835
R19309 vdd.n284 vdd.n283 75.1835
R19310 vdd.n282 vdd.n281 75.1835
R19311 vdd.n280 vdd.n279 75.1835
R19312 vdd.n278 vdd.n277 75.1835
R19313 vdd.n276 vdd.n275 75.1835
R19314 vdd.n274 vdd.n273 75.1835
R19315 vdd.n188 vdd.n187 75.1835
R19316 vdd.n186 vdd.n185 75.1835
R19317 vdd.n184 vdd.n183 75.1835
R19318 vdd.n182 vdd.n181 75.1835
R19319 vdd.n180 vdd.n179 75.1835
R19320 vdd.n178 vdd.n177 75.1835
R19321 vdd.n176 vdd.n175 75.1835
R19322 vdd.n174 vdd.n173 75.1835
R19323 vdd.n172 vdd.n171 75.1835
R19324 vdd.n87 vdd.n86 75.1835
R19325 vdd.n85 vdd.n84 75.1835
R19326 vdd.n83 vdd.n82 75.1835
R19327 vdd.n81 vdd.n80 75.1835
R19328 vdd.n79 vdd.n78 75.1835
R19329 vdd.n77 vdd.n76 75.1835
R19330 vdd.n75 vdd.n74 75.1835
R19331 vdd.n73 vdd.n72 75.1835
R19332 vdd.n71 vdd.n70 75.1835
R19333 vdd.n2114 vdd.n2113 75.1835
R19334 vdd.n2116 vdd.n2115 75.1835
R19335 vdd.n2118 vdd.n2117 75.1835
R19336 vdd.n2120 vdd.n2119 75.1835
R19337 vdd.n2122 vdd.n2121 75.1835
R19338 vdd.n2124 vdd.n2123 75.1835
R19339 vdd.n2126 vdd.n2125 75.1835
R19340 vdd.n2128 vdd.n2127 75.1835
R19341 vdd.n2130 vdd.n2129 75.1835
R19342 vdd.n2012 vdd.n2011 75.1835
R19343 vdd.n2014 vdd.n2013 75.1835
R19344 vdd.n2016 vdd.n2015 75.1835
R19345 vdd.n2018 vdd.n2017 75.1835
R19346 vdd.n2020 vdd.n2019 75.1835
R19347 vdd.n2022 vdd.n2021 75.1835
R19348 vdd.n2024 vdd.n2023 75.1835
R19349 vdd.n2026 vdd.n2025 75.1835
R19350 vdd.n2028 vdd.n2027 75.1835
R19351 vdd.n1911 vdd.n1910 75.1835
R19352 vdd.n1913 vdd.n1912 75.1835
R19353 vdd.n1915 vdd.n1914 75.1835
R19354 vdd.n1917 vdd.n1916 75.1835
R19355 vdd.n1919 vdd.n1918 75.1835
R19356 vdd.n1921 vdd.n1920 75.1835
R19357 vdd.n1923 vdd.n1922 75.1835
R19358 vdd.n1925 vdd.n1924 75.1835
R19359 vdd.n1927 vdd.n1926 75.1835
R19360 vdd.n2939 vdd.n2938 72.8958
R19361 vdd.n2938 vdd.n2682 72.8958
R19362 vdd.n2938 vdd.n2683 72.8958
R19363 vdd.n2938 vdd.n2684 72.8958
R19364 vdd.n2938 vdd.n2685 72.8958
R19365 vdd.n2938 vdd.n2686 72.8958
R19366 vdd.n2938 vdd.n2687 72.8958
R19367 vdd.n2938 vdd.n2688 72.8958
R19368 vdd.n2938 vdd.n2689 72.8958
R19369 vdd.n2938 vdd.n2690 72.8958
R19370 vdd.n2938 vdd.n2691 72.8958
R19371 vdd.n2938 vdd.n2692 72.8958
R19372 vdd.n2938 vdd.n2693 72.8958
R19373 vdd.n2938 vdd.n2694 72.8958
R19374 vdd.n2938 vdd.n2695 72.8958
R19375 vdd.n2938 vdd.n2696 72.8958
R19376 vdd.n2938 vdd.n2697 72.8958
R19377 vdd.n803 vdd.n692 72.8958
R19378 vdd.n3158 vdd.n692 72.8958
R19379 vdd.n797 vdd.n692 72.8958
R19380 vdd.n3165 vdd.n692 72.8958
R19381 vdd.n794 vdd.n692 72.8958
R19382 vdd.n3172 vdd.n692 72.8958
R19383 vdd.n791 vdd.n692 72.8958
R19384 vdd.n3179 vdd.n692 72.8958
R19385 vdd.n3182 vdd.n692 72.8958
R19386 vdd.n3038 vdd.n692 72.8958
R19387 vdd.n3043 vdd.n692 72.8958
R19388 vdd.n3037 vdd.n692 72.8958
R19389 vdd.n3050 vdd.n692 72.8958
R19390 vdd.n3034 vdd.n692 72.8958
R19391 vdd.n3057 vdd.n692 72.8958
R19392 vdd.n3031 vdd.n692 72.8958
R19393 vdd.n3064 vdd.n692 72.8958
R19394 vdd.n2417 vdd.n2416 72.8958
R19395 vdd.n2417 vdd.n1084 72.8958
R19396 vdd.n2417 vdd.n1085 72.8958
R19397 vdd.n2417 vdd.n1086 72.8958
R19398 vdd.n2417 vdd.n1087 72.8958
R19399 vdd.n2417 vdd.n1088 72.8958
R19400 vdd.n2417 vdd.n1089 72.8958
R19401 vdd.n2417 vdd.n1090 72.8958
R19402 vdd.n2417 vdd.n1091 72.8958
R19403 vdd.n2417 vdd.n1092 72.8958
R19404 vdd.n2417 vdd.n1093 72.8958
R19405 vdd.n2417 vdd.n1094 72.8958
R19406 vdd.n2417 vdd.n1095 72.8958
R19407 vdd.n2417 vdd.n1096 72.8958
R19408 vdd.n2417 vdd.n1097 72.8958
R19409 vdd.n2417 vdd.n1098 72.8958
R19410 vdd.n2417 vdd.n1099 72.8958
R19411 vdd.n2665 vdd.n952 72.8958
R19412 vdd.n2665 vdd.n953 72.8958
R19413 vdd.n2665 vdd.n954 72.8958
R19414 vdd.n2665 vdd.n955 72.8958
R19415 vdd.n2665 vdd.n956 72.8958
R19416 vdd.n2665 vdd.n957 72.8958
R19417 vdd.n2665 vdd.n958 72.8958
R19418 vdd.n2665 vdd.n959 72.8958
R19419 vdd.n2665 vdd.n960 72.8958
R19420 vdd.n2665 vdd.n961 72.8958
R19421 vdd.n2665 vdd.n962 72.8958
R19422 vdd.n2665 vdd.n963 72.8958
R19423 vdd.n2665 vdd.n964 72.8958
R19424 vdd.n2665 vdd.n965 72.8958
R19425 vdd.n2665 vdd.n966 72.8958
R19426 vdd.n2665 vdd.n967 72.8958
R19427 vdd.n2665 vdd.n968 72.8958
R19428 vdd.n2938 vdd.n2937 72.8958
R19429 vdd.n2938 vdd.n2666 72.8958
R19430 vdd.n2938 vdd.n2667 72.8958
R19431 vdd.n2938 vdd.n2668 72.8958
R19432 vdd.n2938 vdd.n2669 72.8958
R19433 vdd.n2938 vdd.n2670 72.8958
R19434 vdd.n2938 vdd.n2671 72.8958
R19435 vdd.n2938 vdd.n2672 72.8958
R19436 vdd.n2938 vdd.n2673 72.8958
R19437 vdd.n2938 vdd.n2674 72.8958
R19438 vdd.n2938 vdd.n2675 72.8958
R19439 vdd.n2938 vdd.n2676 72.8958
R19440 vdd.n2938 vdd.n2677 72.8958
R19441 vdd.n2938 vdd.n2678 72.8958
R19442 vdd.n2938 vdd.n2679 72.8958
R19443 vdd.n2938 vdd.n2680 72.8958
R19444 vdd.n2938 vdd.n2681 72.8958
R19445 vdd.n3088 vdd.n692 72.8958
R19446 vdd.n835 vdd.n692 72.8958
R19447 vdd.n3096 vdd.n692 72.8958
R19448 vdd.n830 vdd.n692 72.8958
R19449 vdd.n3103 vdd.n692 72.8958
R19450 vdd.n827 vdd.n692 72.8958
R19451 vdd.n3110 vdd.n692 72.8958
R19452 vdd.n824 vdd.n692 72.8958
R19453 vdd.n3117 vdd.n692 72.8958
R19454 vdd.n3121 vdd.n692 72.8958
R19455 vdd.n821 vdd.n692 72.8958
R19456 vdd.n3128 vdd.n692 72.8958
R19457 vdd.n818 vdd.n692 72.8958
R19458 vdd.n3135 vdd.n692 72.8958
R19459 vdd.n815 vdd.n692 72.8958
R19460 vdd.n3142 vdd.n692 72.8958
R19461 vdd.n3145 vdd.n692 72.8958
R19462 vdd.n2665 vdd.n950 72.8958
R19463 vdd.n2665 vdd.n949 72.8958
R19464 vdd.n2665 vdd.n948 72.8958
R19465 vdd.n2665 vdd.n947 72.8958
R19466 vdd.n2665 vdd.n946 72.8958
R19467 vdd.n2665 vdd.n945 72.8958
R19468 vdd.n2665 vdd.n944 72.8958
R19469 vdd.n2665 vdd.n943 72.8958
R19470 vdd.n2665 vdd.n942 72.8958
R19471 vdd.n2665 vdd.n941 72.8958
R19472 vdd.n2665 vdd.n940 72.8958
R19473 vdd.n2665 vdd.n939 72.8958
R19474 vdd.n2665 vdd.n938 72.8958
R19475 vdd.n2665 vdd.n937 72.8958
R19476 vdd.n2665 vdd.n936 72.8958
R19477 vdd.n2665 vdd.n935 72.8958
R19478 vdd.n2665 vdd.n934 72.8958
R19479 vdd.n2418 vdd.n2417 72.8958
R19480 vdd.n2417 vdd.n1100 72.8958
R19481 vdd.n2417 vdd.n1101 72.8958
R19482 vdd.n2417 vdd.n1102 72.8958
R19483 vdd.n2417 vdd.n1103 72.8958
R19484 vdd.n2417 vdd.n1104 72.8958
R19485 vdd.n2417 vdd.n1105 72.8958
R19486 vdd.n2417 vdd.n1106 72.8958
R19487 vdd.n2417 vdd.n1107 72.8958
R19488 vdd.n2417 vdd.n1108 72.8958
R19489 vdd.n2417 vdd.n1109 72.8958
R19490 vdd.n2417 vdd.n1110 72.8958
R19491 vdd.n2417 vdd.n1111 72.8958
R19492 vdd.n2417 vdd.n1112 72.8958
R19493 vdd.n2417 vdd.n1113 72.8958
R19494 vdd.n2417 vdd.n1114 72.8958
R19495 vdd.n2417 vdd.n1115 72.8958
R19496 vdd.n1781 vdd.n1780 66.2847
R19497 vdd.n1780 vdd.n1556 66.2847
R19498 vdd.n1780 vdd.n1557 66.2847
R19499 vdd.n1780 vdd.n1558 66.2847
R19500 vdd.n1780 vdd.n1559 66.2847
R19501 vdd.n1780 vdd.n1560 66.2847
R19502 vdd.n1780 vdd.n1561 66.2847
R19503 vdd.n1780 vdd.n1562 66.2847
R19504 vdd.n1780 vdd.n1563 66.2847
R19505 vdd.n1780 vdd.n1564 66.2847
R19506 vdd.n1780 vdd.n1565 66.2847
R19507 vdd.n1780 vdd.n1566 66.2847
R19508 vdd.n1780 vdd.n1567 66.2847
R19509 vdd.n1780 vdd.n1568 66.2847
R19510 vdd.n1780 vdd.n1569 66.2847
R19511 vdd.n1780 vdd.n1570 66.2847
R19512 vdd.n1780 vdd.n1571 66.2847
R19513 vdd.n1780 vdd.n1572 66.2847
R19514 vdd.n1780 vdd.n1573 66.2847
R19515 vdd.n1780 vdd.n1574 66.2847
R19516 vdd.n1780 vdd.n1575 66.2847
R19517 vdd.n1780 vdd.n1576 66.2847
R19518 vdd.n1780 vdd.n1577 66.2847
R19519 vdd.n1780 vdd.n1578 66.2847
R19520 vdd.n1780 vdd.n1579 66.2847
R19521 vdd.n1780 vdd.n1580 66.2847
R19522 vdd.n1780 vdd.n1581 66.2847
R19523 vdd.n1780 vdd.n1582 66.2847
R19524 vdd.n1780 vdd.n1583 66.2847
R19525 vdd.n1780 vdd.n1584 66.2847
R19526 vdd.n1780 vdd.n1585 66.2847
R19527 vdd.n1433 vdd.n1083 66.2847
R19528 vdd.n1430 vdd.n1083 66.2847
R19529 vdd.n1426 vdd.n1083 66.2847
R19530 vdd.n2279 vdd.n1083 66.2847
R19531 vdd.n1217 vdd.n1083 66.2847
R19532 vdd.n2286 vdd.n1083 66.2847
R19533 vdd.n1210 vdd.n1083 66.2847
R19534 vdd.n2293 vdd.n1083 66.2847
R19535 vdd.n1203 vdd.n1083 66.2847
R19536 vdd.n2300 vdd.n1083 66.2847
R19537 vdd.n1197 vdd.n1083 66.2847
R19538 vdd.n1192 vdd.n1083 66.2847
R19539 vdd.n2311 vdd.n1083 66.2847
R19540 vdd.n1184 vdd.n1083 66.2847
R19541 vdd.n2318 vdd.n1083 66.2847
R19542 vdd.n1177 vdd.n1083 66.2847
R19543 vdd.n2325 vdd.n1083 66.2847
R19544 vdd.n1170 vdd.n1083 66.2847
R19545 vdd.n2332 vdd.n1083 66.2847
R19546 vdd.n1163 vdd.n1083 66.2847
R19547 vdd.n2339 vdd.n1083 66.2847
R19548 vdd.n1157 vdd.n1083 66.2847
R19549 vdd.n1152 vdd.n1083 66.2847
R19550 vdd.n2350 vdd.n1083 66.2847
R19551 vdd.n1144 vdd.n1083 66.2847
R19552 vdd.n2357 vdd.n1083 66.2847
R19553 vdd.n1137 vdd.n1083 66.2847
R19554 vdd.n2364 vdd.n1083 66.2847
R19555 vdd.n1130 vdd.n1083 66.2847
R19556 vdd.n2371 vdd.n1083 66.2847
R19557 vdd.n2376 vdd.n1083 66.2847
R19558 vdd.n1126 vdd.n1083 66.2847
R19559 vdd.n3315 vdd.n3314 66.2847
R19560 vdd.n3315 vdd.n693 66.2847
R19561 vdd.n3315 vdd.n694 66.2847
R19562 vdd.n3315 vdd.n695 66.2847
R19563 vdd.n3315 vdd.n696 66.2847
R19564 vdd.n3315 vdd.n697 66.2847
R19565 vdd.n3315 vdd.n698 66.2847
R19566 vdd.n3315 vdd.n699 66.2847
R19567 vdd.n3315 vdd.n700 66.2847
R19568 vdd.n3315 vdd.n701 66.2847
R19569 vdd.n3315 vdd.n702 66.2847
R19570 vdd.n3315 vdd.n703 66.2847
R19571 vdd.n3315 vdd.n704 66.2847
R19572 vdd.n3315 vdd.n705 66.2847
R19573 vdd.n3315 vdd.n706 66.2847
R19574 vdd.n3315 vdd.n707 66.2847
R19575 vdd.n3315 vdd.n708 66.2847
R19576 vdd.n3315 vdd.n709 66.2847
R19577 vdd.n3315 vdd.n710 66.2847
R19578 vdd.n3315 vdd.n711 66.2847
R19579 vdd.n3315 vdd.n712 66.2847
R19580 vdd.n3315 vdd.n713 66.2847
R19581 vdd.n3315 vdd.n714 66.2847
R19582 vdd.n3315 vdd.n715 66.2847
R19583 vdd.n3315 vdd.n716 66.2847
R19584 vdd.n3315 vdd.n717 66.2847
R19585 vdd.n3315 vdd.n718 66.2847
R19586 vdd.n3315 vdd.n719 66.2847
R19587 vdd.n3315 vdd.n720 66.2847
R19588 vdd.n3315 vdd.n721 66.2847
R19589 vdd.n3315 vdd.n722 66.2847
R19590 vdd.n3446 vdd.n3445 66.2847
R19591 vdd.n3446 vdd.n424 66.2847
R19592 vdd.n3446 vdd.n423 66.2847
R19593 vdd.n3446 vdd.n422 66.2847
R19594 vdd.n3446 vdd.n421 66.2847
R19595 vdd.n3446 vdd.n420 66.2847
R19596 vdd.n3446 vdd.n419 66.2847
R19597 vdd.n3446 vdd.n418 66.2847
R19598 vdd.n3446 vdd.n417 66.2847
R19599 vdd.n3446 vdd.n416 66.2847
R19600 vdd.n3446 vdd.n415 66.2847
R19601 vdd.n3446 vdd.n414 66.2847
R19602 vdd.n3446 vdd.n413 66.2847
R19603 vdd.n3446 vdd.n412 66.2847
R19604 vdd.n3446 vdd.n411 66.2847
R19605 vdd.n3446 vdd.n410 66.2847
R19606 vdd.n3446 vdd.n409 66.2847
R19607 vdd.n3446 vdd.n408 66.2847
R19608 vdd.n3446 vdd.n407 66.2847
R19609 vdd.n3446 vdd.n406 66.2847
R19610 vdd.n3446 vdd.n405 66.2847
R19611 vdd.n3446 vdd.n404 66.2847
R19612 vdd.n3446 vdd.n403 66.2847
R19613 vdd.n3446 vdd.n402 66.2847
R19614 vdd.n3446 vdd.n401 66.2847
R19615 vdd.n3446 vdd.n400 66.2847
R19616 vdd.n3446 vdd.n399 66.2847
R19617 vdd.n3446 vdd.n398 66.2847
R19618 vdd.n3446 vdd.n397 66.2847
R19619 vdd.n3446 vdd.n396 66.2847
R19620 vdd.n3446 vdd.n395 66.2847
R19621 vdd.n3446 vdd.n394 66.2847
R19622 vdd.n467 vdd.n394 52.4337
R19623 vdd.n473 vdd.n395 52.4337
R19624 vdd.n477 vdd.n396 52.4337
R19625 vdd.n483 vdd.n397 52.4337
R19626 vdd.n487 vdd.n398 52.4337
R19627 vdd.n493 vdd.n399 52.4337
R19628 vdd.n497 vdd.n400 52.4337
R19629 vdd.n503 vdd.n401 52.4337
R19630 vdd.n507 vdd.n402 52.4337
R19631 vdd.n513 vdd.n403 52.4337
R19632 vdd.n517 vdd.n404 52.4337
R19633 vdd.n523 vdd.n405 52.4337
R19634 vdd.n527 vdd.n406 52.4337
R19635 vdd.n533 vdd.n407 52.4337
R19636 vdd.n537 vdd.n408 52.4337
R19637 vdd.n543 vdd.n409 52.4337
R19638 vdd.n547 vdd.n410 52.4337
R19639 vdd.n553 vdd.n411 52.4337
R19640 vdd.n557 vdd.n412 52.4337
R19641 vdd.n563 vdd.n413 52.4337
R19642 vdd.n567 vdd.n414 52.4337
R19643 vdd.n573 vdd.n415 52.4337
R19644 vdd.n577 vdd.n416 52.4337
R19645 vdd.n583 vdd.n417 52.4337
R19646 vdd.n587 vdd.n418 52.4337
R19647 vdd.n593 vdd.n419 52.4337
R19648 vdd.n597 vdd.n420 52.4337
R19649 vdd.n603 vdd.n421 52.4337
R19650 vdd.n607 vdd.n422 52.4337
R19651 vdd.n613 vdd.n423 52.4337
R19652 vdd.n616 vdd.n424 52.4337
R19653 vdd.n3445 vdd.n3444 52.4337
R19654 vdd.n3314 vdd.n3313 52.4337
R19655 vdd.n728 vdd.n693 52.4337
R19656 vdd.n734 vdd.n694 52.4337
R19657 vdd.n3303 vdd.n695 52.4337
R19658 vdd.n3299 vdd.n696 52.4337
R19659 vdd.n3295 vdd.n697 52.4337
R19660 vdd.n3291 vdd.n698 52.4337
R19661 vdd.n3287 vdd.n699 52.4337
R19662 vdd.n3283 vdd.n700 52.4337
R19663 vdd.n3279 vdd.n701 52.4337
R19664 vdd.n3271 vdd.n702 52.4337
R19665 vdd.n3267 vdd.n703 52.4337
R19666 vdd.n3263 vdd.n704 52.4337
R19667 vdd.n3259 vdd.n705 52.4337
R19668 vdd.n3255 vdd.n706 52.4337
R19669 vdd.n3251 vdd.n707 52.4337
R19670 vdd.n3247 vdd.n708 52.4337
R19671 vdd.n3243 vdd.n709 52.4337
R19672 vdd.n3239 vdd.n710 52.4337
R19673 vdd.n3235 vdd.n711 52.4337
R19674 vdd.n3231 vdd.n712 52.4337
R19675 vdd.n3225 vdd.n713 52.4337
R19676 vdd.n3221 vdd.n714 52.4337
R19677 vdd.n3217 vdd.n715 52.4337
R19678 vdd.n3213 vdd.n716 52.4337
R19679 vdd.n3209 vdd.n717 52.4337
R19680 vdd.n3205 vdd.n718 52.4337
R19681 vdd.n3201 vdd.n719 52.4337
R19682 vdd.n3197 vdd.n720 52.4337
R19683 vdd.n3193 vdd.n721 52.4337
R19684 vdd.n3189 vdd.n722 52.4337
R19685 vdd.n2378 vdd.n1126 52.4337
R19686 vdd.n2376 vdd.n2375 52.4337
R19687 vdd.n2371 vdd.n2370 52.4337
R19688 vdd.n2366 vdd.n1130 52.4337
R19689 vdd.n2364 vdd.n2363 52.4337
R19690 vdd.n2359 vdd.n1137 52.4337
R19691 vdd.n2357 vdd.n2356 52.4337
R19692 vdd.n2352 vdd.n1144 52.4337
R19693 vdd.n2350 vdd.n2349 52.4337
R19694 vdd.n1153 vdd.n1152 52.4337
R19695 vdd.n2341 vdd.n1157 52.4337
R19696 vdd.n2339 vdd.n2338 52.4337
R19697 vdd.n2334 vdd.n1163 52.4337
R19698 vdd.n2332 vdd.n2331 52.4337
R19699 vdd.n2327 vdd.n1170 52.4337
R19700 vdd.n2325 vdd.n2324 52.4337
R19701 vdd.n2320 vdd.n1177 52.4337
R19702 vdd.n2318 vdd.n2317 52.4337
R19703 vdd.n2313 vdd.n1184 52.4337
R19704 vdd.n2311 vdd.n2310 52.4337
R19705 vdd.n1193 vdd.n1192 52.4337
R19706 vdd.n2302 vdd.n1197 52.4337
R19707 vdd.n2300 vdd.n2299 52.4337
R19708 vdd.n2295 vdd.n1203 52.4337
R19709 vdd.n2293 vdd.n2292 52.4337
R19710 vdd.n2288 vdd.n1210 52.4337
R19711 vdd.n2286 vdd.n2285 52.4337
R19712 vdd.n2281 vdd.n1217 52.4337
R19713 vdd.n2279 vdd.n2278 52.4337
R19714 vdd.n1427 vdd.n1426 52.4337
R19715 vdd.n1431 vdd.n1430 52.4337
R19716 vdd.n2267 vdd.n1433 52.4337
R19717 vdd.n1782 vdd.n1781 52.4337
R19718 vdd.n1588 vdd.n1556 52.4337
R19719 vdd.n1592 vdd.n1557 52.4337
R19720 vdd.n1594 vdd.n1558 52.4337
R19721 vdd.n1598 vdd.n1559 52.4337
R19722 vdd.n1600 vdd.n1560 52.4337
R19723 vdd.n1604 vdd.n1561 52.4337
R19724 vdd.n1606 vdd.n1562 52.4337
R19725 vdd.n1610 vdd.n1563 52.4337
R19726 vdd.n1612 vdd.n1564 52.4337
R19727 vdd.n1618 vdd.n1565 52.4337
R19728 vdd.n1620 vdd.n1566 52.4337
R19729 vdd.n1624 vdd.n1567 52.4337
R19730 vdd.n1626 vdd.n1568 52.4337
R19731 vdd.n1630 vdd.n1569 52.4337
R19732 vdd.n1632 vdd.n1570 52.4337
R19733 vdd.n1636 vdd.n1571 52.4337
R19734 vdd.n1638 vdd.n1572 52.4337
R19735 vdd.n1642 vdd.n1573 52.4337
R19736 vdd.n1644 vdd.n1574 52.4337
R19737 vdd.n1716 vdd.n1575 52.4337
R19738 vdd.n1649 vdd.n1576 52.4337
R19739 vdd.n1653 vdd.n1577 52.4337
R19740 vdd.n1655 vdd.n1578 52.4337
R19741 vdd.n1659 vdd.n1579 52.4337
R19742 vdd.n1661 vdd.n1580 52.4337
R19743 vdd.n1665 vdd.n1581 52.4337
R19744 vdd.n1667 vdd.n1582 52.4337
R19745 vdd.n1671 vdd.n1583 52.4337
R19746 vdd.n1673 vdd.n1584 52.4337
R19747 vdd.n1677 vdd.n1585 52.4337
R19748 vdd.n1781 vdd.n1555 52.4337
R19749 vdd.n1591 vdd.n1556 52.4337
R19750 vdd.n1593 vdd.n1557 52.4337
R19751 vdd.n1597 vdd.n1558 52.4337
R19752 vdd.n1599 vdd.n1559 52.4337
R19753 vdd.n1603 vdd.n1560 52.4337
R19754 vdd.n1605 vdd.n1561 52.4337
R19755 vdd.n1609 vdd.n1562 52.4337
R19756 vdd.n1611 vdd.n1563 52.4337
R19757 vdd.n1617 vdd.n1564 52.4337
R19758 vdd.n1619 vdd.n1565 52.4337
R19759 vdd.n1623 vdd.n1566 52.4337
R19760 vdd.n1625 vdd.n1567 52.4337
R19761 vdd.n1629 vdd.n1568 52.4337
R19762 vdd.n1631 vdd.n1569 52.4337
R19763 vdd.n1635 vdd.n1570 52.4337
R19764 vdd.n1637 vdd.n1571 52.4337
R19765 vdd.n1641 vdd.n1572 52.4337
R19766 vdd.n1643 vdd.n1573 52.4337
R19767 vdd.n1647 vdd.n1574 52.4337
R19768 vdd.n1648 vdd.n1575 52.4337
R19769 vdd.n1652 vdd.n1576 52.4337
R19770 vdd.n1654 vdd.n1577 52.4337
R19771 vdd.n1658 vdd.n1578 52.4337
R19772 vdd.n1660 vdd.n1579 52.4337
R19773 vdd.n1664 vdd.n1580 52.4337
R19774 vdd.n1666 vdd.n1581 52.4337
R19775 vdd.n1670 vdd.n1582 52.4337
R19776 vdd.n1672 vdd.n1583 52.4337
R19777 vdd.n1676 vdd.n1584 52.4337
R19778 vdd.n1678 vdd.n1585 52.4337
R19779 vdd.n1433 vdd.n1432 52.4337
R19780 vdd.n1430 vdd.n1429 52.4337
R19781 vdd.n1426 vdd.n1218 52.4337
R19782 vdd.n2280 vdd.n2279 52.4337
R19783 vdd.n1217 vdd.n1211 52.4337
R19784 vdd.n2287 vdd.n2286 52.4337
R19785 vdd.n1210 vdd.n1204 52.4337
R19786 vdd.n2294 vdd.n2293 52.4337
R19787 vdd.n1203 vdd.n1198 52.4337
R19788 vdd.n2301 vdd.n2300 52.4337
R19789 vdd.n1197 vdd.n1196 52.4337
R19790 vdd.n1192 vdd.n1185 52.4337
R19791 vdd.n2312 vdd.n2311 52.4337
R19792 vdd.n1184 vdd.n1178 52.4337
R19793 vdd.n2319 vdd.n2318 52.4337
R19794 vdd.n1177 vdd.n1171 52.4337
R19795 vdd.n2326 vdd.n2325 52.4337
R19796 vdd.n1170 vdd.n1164 52.4337
R19797 vdd.n2333 vdd.n2332 52.4337
R19798 vdd.n1163 vdd.n1158 52.4337
R19799 vdd.n2340 vdd.n2339 52.4337
R19800 vdd.n1157 vdd.n1156 52.4337
R19801 vdd.n1152 vdd.n1145 52.4337
R19802 vdd.n2351 vdd.n2350 52.4337
R19803 vdd.n1144 vdd.n1138 52.4337
R19804 vdd.n2358 vdd.n2357 52.4337
R19805 vdd.n1137 vdd.n1131 52.4337
R19806 vdd.n2365 vdd.n2364 52.4337
R19807 vdd.n1130 vdd.n1127 52.4337
R19808 vdd.n2372 vdd.n2371 52.4337
R19809 vdd.n2377 vdd.n2376 52.4337
R19810 vdd.n1437 vdd.n1126 52.4337
R19811 vdd.n3314 vdd.n725 52.4337
R19812 vdd.n733 vdd.n693 52.4337
R19813 vdd.n3304 vdd.n694 52.4337
R19814 vdd.n3300 vdd.n695 52.4337
R19815 vdd.n3296 vdd.n696 52.4337
R19816 vdd.n3292 vdd.n697 52.4337
R19817 vdd.n3288 vdd.n698 52.4337
R19818 vdd.n3284 vdd.n699 52.4337
R19819 vdd.n3280 vdd.n700 52.4337
R19820 vdd.n3270 vdd.n701 52.4337
R19821 vdd.n3268 vdd.n702 52.4337
R19822 vdd.n3264 vdd.n703 52.4337
R19823 vdd.n3260 vdd.n704 52.4337
R19824 vdd.n3256 vdd.n705 52.4337
R19825 vdd.n3252 vdd.n706 52.4337
R19826 vdd.n3248 vdd.n707 52.4337
R19827 vdd.n3244 vdd.n708 52.4337
R19828 vdd.n3240 vdd.n709 52.4337
R19829 vdd.n3236 vdd.n710 52.4337
R19830 vdd.n3232 vdd.n711 52.4337
R19831 vdd.n3224 vdd.n712 52.4337
R19832 vdd.n3222 vdd.n713 52.4337
R19833 vdd.n3218 vdd.n714 52.4337
R19834 vdd.n3214 vdd.n715 52.4337
R19835 vdd.n3210 vdd.n716 52.4337
R19836 vdd.n3206 vdd.n717 52.4337
R19837 vdd.n3202 vdd.n718 52.4337
R19838 vdd.n3198 vdd.n719 52.4337
R19839 vdd.n3194 vdd.n720 52.4337
R19840 vdd.n3190 vdd.n721 52.4337
R19841 vdd.n722 vdd.n691 52.4337
R19842 vdd.n3445 vdd.n425 52.4337
R19843 vdd.n614 vdd.n424 52.4337
R19844 vdd.n608 vdd.n423 52.4337
R19845 vdd.n604 vdd.n422 52.4337
R19846 vdd.n598 vdd.n421 52.4337
R19847 vdd.n594 vdd.n420 52.4337
R19848 vdd.n588 vdd.n419 52.4337
R19849 vdd.n584 vdd.n418 52.4337
R19850 vdd.n578 vdd.n417 52.4337
R19851 vdd.n574 vdd.n416 52.4337
R19852 vdd.n568 vdd.n415 52.4337
R19853 vdd.n564 vdd.n414 52.4337
R19854 vdd.n558 vdd.n413 52.4337
R19855 vdd.n554 vdd.n412 52.4337
R19856 vdd.n548 vdd.n411 52.4337
R19857 vdd.n544 vdd.n410 52.4337
R19858 vdd.n538 vdd.n409 52.4337
R19859 vdd.n534 vdd.n408 52.4337
R19860 vdd.n528 vdd.n407 52.4337
R19861 vdd.n524 vdd.n406 52.4337
R19862 vdd.n518 vdd.n405 52.4337
R19863 vdd.n514 vdd.n404 52.4337
R19864 vdd.n508 vdd.n403 52.4337
R19865 vdd.n504 vdd.n402 52.4337
R19866 vdd.n498 vdd.n401 52.4337
R19867 vdd.n494 vdd.n400 52.4337
R19868 vdd.n488 vdd.n399 52.4337
R19869 vdd.n484 vdd.n398 52.4337
R19870 vdd.n478 vdd.n397 52.4337
R19871 vdd.n474 vdd.n396 52.4337
R19872 vdd.n468 vdd.n395 52.4337
R19873 vdd.n394 vdd.n392 52.4337
R19874 vdd.t130 vdd.t136 51.4683
R19875 vdd.n274 vdd.n272 42.0461
R19876 vdd.n172 vdd.n170 42.0461
R19877 vdd.n71 vdd.n69 42.0461
R19878 vdd.n2114 vdd.n2112 42.0461
R19879 vdd.n2012 vdd.n2010 42.0461
R19880 vdd.n1911 vdd.n1909 42.0461
R19881 vdd.n332 vdd.n331 41.6884
R19882 vdd.n230 vdd.n229 41.6884
R19883 vdd.n129 vdd.n128 41.6884
R19884 vdd.n2172 vdd.n2171 41.6884
R19885 vdd.n2070 vdd.n2069 41.6884
R19886 vdd.n1969 vdd.n1968 41.6884
R19887 vdd.n1681 vdd.n1680 41.1157
R19888 vdd.n1719 vdd.n1718 41.1157
R19889 vdd.n1615 vdd.n1614 41.1157
R19890 vdd.n428 vdd.n427 41.1157
R19891 vdd.n566 vdd.n441 41.1157
R19892 vdd.n454 vdd.n453 41.1157
R19893 vdd.n3145 vdd.n3144 39.2114
R19894 vdd.n3142 vdd.n3141 39.2114
R19895 vdd.n3137 vdd.n815 39.2114
R19896 vdd.n3135 vdd.n3134 39.2114
R19897 vdd.n3130 vdd.n818 39.2114
R19898 vdd.n3128 vdd.n3127 39.2114
R19899 vdd.n3123 vdd.n821 39.2114
R19900 vdd.n3121 vdd.n3120 39.2114
R19901 vdd.n3117 vdd.n3116 39.2114
R19902 vdd.n3112 vdd.n824 39.2114
R19903 vdd.n3110 vdd.n3109 39.2114
R19904 vdd.n3105 vdd.n827 39.2114
R19905 vdd.n3103 vdd.n3102 39.2114
R19906 vdd.n3098 vdd.n830 39.2114
R19907 vdd.n3096 vdd.n3095 39.2114
R19908 vdd.n3090 vdd.n835 39.2114
R19909 vdd.n3088 vdd.n3087 39.2114
R19910 vdd.n2937 vdd.n2936 39.2114
R19911 vdd.n2931 vdd.n2666 39.2114
R19912 vdd.n2928 vdd.n2667 39.2114
R19913 vdd.n2924 vdd.n2668 39.2114
R19914 vdd.n2920 vdd.n2669 39.2114
R19915 vdd.n2916 vdd.n2670 39.2114
R19916 vdd.n2912 vdd.n2671 39.2114
R19917 vdd.n2908 vdd.n2672 39.2114
R19918 vdd.n2904 vdd.n2673 39.2114
R19919 vdd.n2900 vdd.n2674 39.2114
R19920 vdd.n2896 vdd.n2675 39.2114
R19921 vdd.n2892 vdd.n2676 39.2114
R19922 vdd.n2888 vdd.n2677 39.2114
R19923 vdd.n2884 vdd.n2678 39.2114
R19924 vdd.n2880 vdd.n2679 39.2114
R19925 vdd.n2876 vdd.n2680 39.2114
R19926 vdd.n2871 vdd.n2681 39.2114
R19927 vdd.n2660 vdd.n968 39.2114
R19928 vdd.n2656 vdd.n967 39.2114
R19929 vdd.n2652 vdd.n966 39.2114
R19930 vdd.n2648 vdd.n965 39.2114
R19931 vdd.n2644 vdd.n964 39.2114
R19932 vdd.n2640 vdd.n963 39.2114
R19933 vdd.n2636 vdd.n962 39.2114
R19934 vdd.n2632 vdd.n961 39.2114
R19935 vdd.n2628 vdd.n960 39.2114
R19936 vdd.n2624 vdd.n959 39.2114
R19937 vdd.n2620 vdd.n958 39.2114
R19938 vdd.n2616 vdd.n957 39.2114
R19939 vdd.n2612 vdd.n956 39.2114
R19940 vdd.n2608 vdd.n955 39.2114
R19941 vdd.n2604 vdd.n954 39.2114
R19942 vdd.n2599 vdd.n953 39.2114
R19943 vdd.n2595 vdd.n952 39.2114
R19944 vdd.n2416 vdd.n2415 39.2114
R19945 vdd.n2410 vdd.n1084 39.2114
R19946 vdd.n2407 vdd.n1085 39.2114
R19947 vdd.n2403 vdd.n1086 39.2114
R19948 vdd.n2399 vdd.n1087 39.2114
R19949 vdd.n2395 vdd.n1088 39.2114
R19950 vdd.n2391 vdd.n1089 39.2114
R19951 vdd.n2387 vdd.n1090 39.2114
R19952 vdd.n2383 vdd.n1091 39.2114
R19953 vdd.n1276 vdd.n1092 39.2114
R19954 vdd.n1280 vdd.n1093 39.2114
R19955 vdd.n1284 vdd.n1094 39.2114
R19956 vdd.n1288 vdd.n1095 39.2114
R19957 vdd.n1292 vdd.n1096 39.2114
R19958 vdd.n1296 vdd.n1097 39.2114
R19959 vdd.n1300 vdd.n1098 39.2114
R19960 vdd.n1305 vdd.n1099 39.2114
R19961 vdd.n3064 vdd.n3063 39.2114
R19962 vdd.n3059 vdd.n3031 39.2114
R19963 vdd.n3057 vdd.n3056 39.2114
R19964 vdd.n3052 vdd.n3034 39.2114
R19965 vdd.n3050 vdd.n3049 39.2114
R19966 vdd.n3045 vdd.n3037 39.2114
R19967 vdd.n3043 vdd.n3042 39.2114
R19968 vdd.n3038 vdd.n787 39.2114
R19969 vdd.n3182 vdd.n3181 39.2114
R19970 vdd.n3179 vdd.n3178 39.2114
R19971 vdd.n3174 vdd.n791 39.2114
R19972 vdd.n3172 vdd.n3171 39.2114
R19973 vdd.n3167 vdd.n794 39.2114
R19974 vdd.n3165 vdd.n3164 39.2114
R19975 vdd.n3160 vdd.n797 39.2114
R19976 vdd.n3158 vdd.n3157 39.2114
R19977 vdd.n3153 vdd.n803 39.2114
R19978 vdd.n2940 vdd.n2939 39.2114
R19979 vdd.n2707 vdd.n2682 39.2114
R19980 vdd.n2711 vdd.n2683 39.2114
R19981 vdd.n2715 vdd.n2684 39.2114
R19982 vdd.n2719 vdd.n2685 39.2114
R19983 vdd.n2723 vdd.n2686 39.2114
R19984 vdd.n2727 vdd.n2687 39.2114
R19985 vdd.n2731 vdd.n2688 39.2114
R19986 vdd.n2735 vdd.n2689 39.2114
R19987 vdd.n2739 vdd.n2690 39.2114
R19988 vdd.n2743 vdd.n2691 39.2114
R19989 vdd.n2747 vdd.n2692 39.2114
R19990 vdd.n2751 vdd.n2693 39.2114
R19991 vdd.n2755 vdd.n2694 39.2114
R19992 vdd.n2759 vdd.n2695 39.2114
R19993 vdd.n2763 vdd.n2696 39.2114
R19994 vdd.n2767 vdd.n2697 39.2114
R19995 vdd.n2939 vdd.n933 39.2114
R19996 vdd.n2710 vdd.n2682 39.2114
R19997 vdd.n2714 vdd.n2683 39.2114
R19998 vdd.n2718 vdd.n2684 39.2114
R19999 vdd.n2722 vdd.n2685 39.2114
R20000 vdd.n2726 vdd.n2686 39.2114
R20001 vdd.n2730 vdd.n2687 39.2114
R20002 vdd.n2734 vdd.n2688 39.2114
R20003 vdd.n2738 vdd.n2689 39.2114
R20004 vdd.n2742 vdd.n2690 39.2114
R20005 vdd.n2746 vdd.n2691 39.2114
R20006 vdd.n2750 vdd.n2692 39.2114
R20007 vdd.n2754 vdd.n2693 39.2114
R20008 vdd.n2758 vdd.n2694 39.2114
R20009 vdd.n2762 vdd.n2695 39.2114
R20010 vdd.n2766 vdd.n2696 39.2114
R20011 vdd.n2769 vdd.n2697 39.2114
R20012 vdd.n803 vdd.n798 39.2114
R20013 vdd.n3159 vdd.n3158 39.2114
R20014 vdd.n797 vdd.n795 39.2114
R20015 vdd.n3166 vdd.n3165 39.2114
R20016 vdd.n794 vdd.n792 39.2114
R20017 vdd.n3173 vdd.n3172 39.2114
R20018 vdd.n791 vdd.n789 39.2114
R20019 vdd.n3180 vdd.n3179 39.2114
R20020 vdd.n3183 vdd.n3182 39.2114
R20021 vdd.n3039 vdd.n3038 39.2114
R20022 vdd.n3044 vdd.n3043 39.2114
R20023 vdd.n3037 vdd.n3035 39.2114
R20024 vdd.n3051 vdd.n3050 39.2114
R20025 vdd.n3034 vdd.n3032 39.2114
R20026 vdd.n3058 vdd.n3057 39.2114
R20027 vdd.n3031 vdd.n3029 39.2114
R20028 vdd.n3065 vdd.n3064 39.2114
R20029 vdd.n2416 vdd.n1118 39.2114
R20030 vdd.n2408 vdd.n1084 39.2114
R20031 vdd.n2404 vdd.n1085 39.2114
R20032 vdd.n2400 vdd.n1086 39.2114
R20033 vdd.n2396 vdd.n1087 39.2114
R20034 vdd.n2392 vdd.n1088 39.2114
R20035 vdd.n2388 vdd.n1089 39.2114
R20036 vdd.n2384 vdd.n1090 39.2114
R20037 vdd.n1275 vdd.n1091 39.2114
R20038 vdd.n1279 vdd.n1092 39.2114
R20039 vdd.n1283 vdd.n1093 39.2114
R20040 vdd.n1287 vdd.n1094 39.2114
R20041 vdd.n1291 vdd.n1095 39.2114
R20042 vdd.n1295 vdd.n1096 39.2114
R20043 vdd.n1299 vdd.n1097 39.2114
R20044 vdd.n1304 vdd.n1098 39.2114
R20045 vdd.n1308 vdd.n1099 39.2114
R20046 vdd.n2598 vdd.n952 39.2114
R20047 vdd.n2603 vdd.n953 39.2114
R20048 vdd.n2607 vdd.n954 39.2114
R20049 vdd.n2611 vdd.n955 39.2114
R20050 vdd.n2615 vdd.n956 39.2114
R20051 vdd.n2619 vdd.n957 39.2114
R20052 vdd.n2623 vdd.n958 39.2114
R20053 vdd.n2627 vdd.n959 39.2114
R20054 vdd.n2631 vdd.n960 39.2114
R20055 vdd.n2635 vdd.n961 39.2114
R20056 vdd.n2639 vdd.n962 39.2114
R20057 vdd.n2643 vdd.n963 39.2114
R20058 vdd.n2647 vdd.n964 39.2114
R20059 vdd.n2651 vdd.n965 39.2114
R20060 vdd.n2655 vdd.n966 39.2114
R20061 vdd.n2659 vdd.n967 39.2114
R20062 vdd.n970 vdd.n968 39.2114
R20063 vdd.n2937 vdd.n2700 39.2114
R20064 vdd.n2929 vdd.n2666 39.2114
R20065 vdd.n2925 vdd.n2667 39.2114
R20066 vdd.n2921 vdd.n2668 39.2114
R20067 vdd.n2917 vdd.n2669 39.2114
R20068 vdd.n2913 vdd.n2670 39.2114
R20069 vdd.n2909 vdd.n2671 39.2114
R20070 vdd.n2905 vdd.n2672 39.2114
R20071 vdd.n2901 vdd.n2673 39.2114
R20072 vdd.n2897 vdd.n2674 39.2114
R20073 vdd.n2893 vdd.n2675 39.2114
R20074 vdd.n2889 vdd.n2676 39.2114
R20075 vdd.n2885 vdd.n2677 39.2114
R20076 vdd.n2881 vdd.n2678 39.2114
R20077 vdd.n2877 vdd.n2679 39.2114
R20078 vdd.n2872 vdd.n2680 39.2114
R20079 vdd.n2868 vdd.n2681 39.2114
R20080 vdd.n3089 vdd.n3088 39.2114
R20081 vdd.n835 vdd.n831 39.2114
R20082 vdd.n3097 vdd.n3096 39.2114
R20083 vdd.n830 vdd.n828 39.2114
R20084 vdd.n3104 vdd.n3103 39.2114
R20085 vdd.n827 vdd.n825 39.2114
R20086 vdd.n3111 vdd.n3110 39.2114
R20087 vdd.n824 vdd.n822 39.2114
R20088 vdd.n3118 vdd.n3117 39.2114
R20089 vdd.n3122 vdd.n3121 39.2114
R20090 vdd.n821 vdd.n819 39.2114
R20091 vdd.n3129 vdd.n3128 39.2114
R20092 vdd.n818 vdd.n816 39.2114
R20093 vdd.n3136 vdd.n3135 39.2114
R20094 vdd.n815 vdd.n813 39.2114
R20095 vdd.n3143 vdd.n3142 39.2114
R20096 vdd.n3146 vdd.n3145 39.2114
R20097 vdd.n979 vdd.n934 39.2114
R20098 vdd.n2587 vdd.n935 39.2114
R20099 vdd.n2583 vdd.n936 39.2114
R20100 vdd.n2579 vdd.n937 39.2114
R20101 vdd.n2575 vdd.n938 39.2114
R20102 vdd.n2571 vdd.n939 39.2114
R20103 vdd.n2567 vdd.n940 39.2114
R20104 vdd.n2563 vdd.n941 39.2114
R20105 vdd.n2559 vdd.n942 39.2114
R20106 vdd.n2555 vdd.n943 39.2114
R20107 vdd.n2551 vdd.n944 39.2114
R20108 vdd.n2547 vdd.n945 39.2114
R20109 vdd.n2543 vdd.n946 39.2114
R20110 vdd.n2539 vdd.n947 39.2114
R20111 vdd.n2535 vdd.n948 39.2114
R20112 vdd.n2531 vdd.n949 39.2114
R20113 vdd.n2527 vdd.n950 39.2114
R20114 vdd.n2419 vdd.n2418 39.2114
R20115 vdd.n1222 vdd.n1100 39.2114
R20116 vdd.n1226 vdd.n1101 39.2114
R20117 vdd.n1230 vdd.n1102 39.2114
R20118 vdd.n1234 vdd.n1103 39.2114
R20119 vdd.n1238 vdd.n1104 39.2114
R20120 vdd.n1242 vdd.n1105 39.2114
R20121 vdd.n1246 vdd.n1106 39.2114
R20122 vdd.n1250 vdd.n1107 39.2114
R20123 vdd.n1420 vdd.n1108 39.2114
R20124 vdd.n1417 vdd.n1109 39.2114
R20125 vdd.n1413 vdd.n1110 39.2114
R20126 vdd.n1409 vdd.n1111 39.2114
R20127 vdd.n1405 vdd.n1112 39.2114
R20128 vdd.n1401 vdd.n1113 39.2114
R20129 vdd.n1397 vdd.n1114 39.2114
R20130 vdd.n1393 vdd.n1115 39.2114
R20131 vdd.n2524 vdd.n950 39.2114
R20132 vdd.n2528 vdd.n949 39.2114
R20133 vdd.n2532 vdd.n948 39.2114
R20134 vdd.n2536 vdd.n947 39.2114
R20135 vdd.n2540 vdd.n946 39.2114
R20136 vdd.n2544 vdd.n945 39.2114
R20137 vdd.n2548 vdd.n944 39.2114
R20138 vdd.n2552 vdd.n943 39.2114
R20139 vdd.n2556 vdd.n942 39.2114
R20140 vdd.n2560 vdd.n941 39.2114
R20141 vdd.n2564 vdd.n940 39.2114
R20142 vdd.n2568 vdd.n939 39.2114
R20143 vdd.n2572 vdd.n938 39.2114
R20144 vdd.n2576 vdd.n937 39.2114
R20145 vdd.n2580 vdd.n936 39.2114
R20146 vdd.n2584 vdd.n935 39.2114
R20147 vdd.n2588 vdd.n934 39.2114
R20148 vdd.n2418 vdd.n1082 39.2114
R20149 vdd.n1225 vdd.n1100 39.2114
R20150 vdd.n1229 vdd.n1101 39.2114
R20151 vdd.n1233 vdd.n1102 39.2114
R20152 vdd.n1237 vdd.n1103 39.2114
R20153 vdd.n1241 vdd.n1104 39.2114
R20154 vdd.n1245 vdd.n1105 39.2114
R20155 vdd.n1249 vdd.n1106 39.2114
R20156 vdd.n1252 vdd.n1107 39.2114
R20157 vdd.n1418 vdd.n1108 39.2114
R20158 vdd.n1414 vdd.n1109 39.2114
R20159 vdd.n1410 vdd.n1110 39.2114
R20160 vdd.n1406 vdd.n1111 39.2114
R20161 vdd.n1402 vdd.n1112 39.2114
R20162 vdd.n1398 vdd.n1113 39.2114
R20163 vdd.n1394 vdd.n1114 39.2114
R20164 vdd.n1390 vdd.n1115 39.2114
R20165 vdd.n2271 vdd.n2270 37.2369
R20166 vdd.n2307 vdd.n1191 37.2369
R20167 vdd.n2346 vdd.n1151 37.2369
R20168 vdd.n3230 vdd.n769 37.2369
R20169 vdd.n3278 vdd.n3277 37.2369
R20170 vdd.n690 vdd.n689 37.2369
R20171 vdd.n2414 vdd.n1074 31.0639
R20172 vdd.n2663 vdd.n971 31.0639
R20173 vdd.n2596 vdd.n974 31.0639
R20174 vdd.n1310 vdd.n1307 31.0639
R20175 vdd.n2869 vdd.n2866 31.0639
R20176 vdd.n3086 vdd.n3085 31.0639
R20177 vdd.n2935 vdd.n926 31.0639
R20178 vdd.n3149 vdd.n3148 31.0639
R20179 vdd.n3068 vdd.n3067 31.0639
R20180 vdd.n3154 vdd.n802 31.0639
R20181 vdd.n2773 vdd.n2771 31.0639
R20182 vdd.n2942 vdd.n2941 31.0639
R20183 vdd.n2421 vdd.n2420 31.0639
R20184 vdd.n2591 vdd.n2590 31.0639
R20185 vdd.n2523 vdd.n2522 31.0639
R20186 vdd.n1389 vdd.n1388 31.0639
R20187 vdd.n1255 vdd.n1254 30.449
R20188 vdd.n983 vdd.n982 30.449
R20189 vdd.n1302 vdd.n1274 30.449
R20190 vdd.n2601 vdd.n973 30.449
R20191 vdd.n2706 vdd.n2705 30.449
R20192 vdd.n3092 vdd.n833 30.449
R20193 vdd.n2874 vdd.n2702 30.449
R20194 vdd.n801 vdd.n800 30.449
R20195 vdd.n1780 vdd.n1587 22.2201
R20196 vdd.n2265 vdd.n1083 22.2201
R20197 vdd.n3315 vdd.n723 22.2201
R20198 vdd.n3447 vdd.n3446 22.2201
R20199 vdd.n1791 vdd.n1549 19.3944
R20200 vdd.n1791 vdd.n1547 19.3944
R20201 vdd.n1795 vdd.n1547 19.3944
R20202 vdd.n1795 vdd.n1537 19.3944
R20203 vdd.n1808 vdd.n1537 19.3944
R20204 vdd.n1808 vdd.n1535 19.3944
R20205 vdd.n1812 vdd.n1535 19.3944
R20206 vdd.n1812 vdd.n1527 19.3944
R20207 vdd.n1825 vdd.n1527 19.3944
R20208 vdd.n1825 vdd.n1525 19.3944
R20209 vdd.n1829 vdd.n1525 19.3944
R20210 vdd.n1829 vdd.n1514 19.3944
R20211 vdd.n1841 vdd.n1514 19.3944
R20212 vdd.n1841 vdd.n1512 19.3944
R20213 vdd.n1845 vdd.n1512 19.3944
R20214 vdd.n1845 vdd.n1503 19.3944
R20215 vdd.n1858 vdd.n1503 19.3944
R20216 vdd.n1858 vdd.n1501 19.3944
R20217 vdd.n1862 vdd.n1501 19.3944
R20218 vdd.n1862 vdd.n1492 19.3944
R20219 vdd.n2181 vdd.n1492 19.3944
R20220 vdd.n2181 vdd.n1490 19.3944
R20221 vdd.n2185 vdd.n1490 19.3944
R20222 vdd.n2185 vdd.n1480 19.3944
R20223 vdd.n2198 vdd.n1480 19.3944
R20224 vdd.n2198 vdd.n1478 19.3944
R20225 vdd.n2202 vdd.n1478 19.3944
R20226 vdd.n2202 vdd.n1470 19.3944
R20227 vdd.n2215 vdd.n1470 19.3944
R20228 vdd.n2215 vdd.n1468 19.3944
R20229 vdd.n2219 vdd.n1468 19.3944
R20230 vdd.n2219 vdd.n1457 19.3944
R20231 vdd.n2231 vdd.n1457 19.3944
R20232 vdd.n2231 vdd.n1455 19.3944
R20233 vdd.n2235 vdd.n1455 19.3944
R20234 vdd.n2235 vdd.n1447 19.3944
R20235 vdd.n2248 vdd.n1447 19.3944
R20236 vdd.n2248 vdd.n1444 19.3944
R20237 vdd.n2254 vdd.n1444 19.3944
R20238 vdd.n2254 vdd.n1445 19.3944
R20239 vdd.n1445 vdd.n1435 19.3944
R20240 vdd.n1715 vdd.n1650 19.3944
R20241 vdd.n1711 vdd.n1650 19.3944
R20242 vdd.n1711 vdd.n1710 19.3944
R20243 vdd.n1710 vdd.n1709 19.3944
R20244 vdd.n1709 vdd.n1656 19.3944
R20245 vdd.n1705 vdd.n1656 19.3944
R20246 vdd.n1705 vdd.n1704 19.3944
R20247 vdd.n1704 vdd.n1703 19.3944
R20248 vdd.n1703 vdd.n1662 19.3944
R20249 vdd.n1699 vdd.n1662 19.3944
R20250 vdd.n1699 vdd.n1698 19.3944
R20251 vdd.n1698 vdd.n1697 19.3944
R20252 vdd.n1697 vdd.n1668 19.3944
R20253 vdd.n1693 vdd.n1668 19.3944
R20254 vdd.n1693 vdd.n1692 19.3944
R20255 vdd.n1692 vdd.n1691 19.3944
R20256 vdd.n1691 vdd.n1674 19.3944
R20257 vdd.n1687 vdd.n1674 19.3944
R20258 vdd.n1687 vdd.n1686 19.3944
R20259 vdd.n1686 vdd.n1685 19.3944
R20260 vdd.n1750 vdd.n1749 19.3944
R20261 vdd.n1749 vdd.n1748 19.3944
R20262 vdd.n1748 vdd.n1621 19.3944
R20263 vdd.n1744 vdd.n1621 19.3944
R20264 vdd.n1744 vdd.n1743 19.3944
R20265 vdd.n1743 vdd.n1742 19.3944
R20266 vdd.n1742 vdd.n1627 19.3944
R20267 vdd.n1738 vdd.n1627 19.3944
R20268 vdd.n1738 vdd.n1737 19.3944
R20269 vdd.n1737 vdd.n1736 19.3944
R20270 vdd.n1736 vdd.n1633 19.3944
R20271 vdd.n1732 vdd.n1633 19.3944
R20272 vdd.n1732 vdd.n1731 19.3944
R20273 vdd.n1731 vdd.n1730 19.3944
R20274 vdd.n1730 vdd.n1639 19.3944
R20275 vdd.n1726 vdd.n1639 19.3944
R20276 vdd.n1726 vdd.n1725 19.3944
R20277 vdd.n1725 vdd.n1724 19.3944
R20278 vdd.n1724 vdd.n1645 19.3944
R20279 vdd.n1720 vdd.n1645 19.3944
R20280 vdd.n1783 vdd.n1554 19.3944
R20281 vdd.n1778 vdd.n1554 19.3944
R20282 vdd.n1778 vdd.n1589 19.3944
R20283 vdd.n1774 vdd.n1589 19.3944
R20284 vdd.n1774 vdd.n1773 19.3944
R20285 vdd.n1773 vdd.n1772 19.3944
R20286 vdd.n1772 vdd.n1595 19.3944
R20287 vdd.n1768 vdd.n1595 19.3944
R20288 vdd.n1768 vdd.n1767 19.3944
R20289 vdd.n1767 vdd.n1766 19.3944
R20290 vdd.n1766 vdd.n1601 19.3944
R20291 vdd.n1762 vdd.n1601 19.3944
R20292 vdd.n1762 vdd.n1761 19.3944
R20293 vdd.n1761 vdd.n1760 19.3944
R20294 vdd.n1760 vdd.n1607 19.3944
R20295 vdd.n1756 vdd.n1607 19.3944
R20296 vdd.n1756 vdd.n1755 19.3944
R20297 vdd.n1755 vdd.n1754 19.3944
R20298 vdd.n2303 vdd.n1189 19.3944
R20299 vdd.n2303 vdd.n1195 19.3944
R20300 vdd.n2298 vdd.n1195 19.3944
R20301 vdd.n2298 vdd.n2297 19.3944
R20302 vdd.n2297 vdd.n2296 19.3944
R20303 vdd.n2296 vdd.n1202 19.3944
R20304 vdd.n2291 vdd.n1202 19.3944
R20305 vdd.n2291 vdd.n2290 19.3944
R20306 vdd.n2290 vdd.n2289 19.3944
R20307 vdd.n2289 vdd.n1209 19.3944
R20308 vdd.n2284 vdd.n1209 19.3944
R20309 vdd.n2284 vdd.n2283 19.3944
R20310 vdd.n2283 vdd.n2282 19.3944
R20311 vdd.n2282 vdd.n1216 19.3944
R20312 vdd.n2277 vdd.n1216 19.3944
R20313 vdd.n2277 vdd.n2276 19.3944
R20314 vdd.n1428 vdd.n1221 19.3944
R20315 vdd.n2272 vdd.n1425 19.3944
R20316 vdd.n2342 vdd.n1149 19.3944
R20317 vdd.n2342 vdd.n1155 19.3944
R20318 vdd.n2337 vdd.n1155 19.3944
R20319 vdd.n2337 vdd.n2336 19.3944
R20320 vdd.n2336 vdd.n2335 19.3944
R20321 vdd.n2335 vdd.n1162 19.3944
R20322 vdd.n2330 vdd.n1162 19.3944
R20323 vdd.n2330 vdd.n2329 19.3944
R20324 vdd.n2329 vdd.n2328 19.3944
R20325 vdd.n2328 vdd.n1169 19.3944
R20326 vdd.n2323 vdd.n1169 19.3944
R20327 vdd.n2323 vdd.n2322 19.3944
R20328 vdd.n2322 vdd.n2321 19.3944
R20329 vdd.n2321 vdd.n1176 19.3944
R20330 vdd.n2316 vdd.n1176 19.3944
R20331 vdd.n2316 vdd.n2315 19.3944
R20332 vdd.n2315 vdd.n2314 19.3944
R20333 vdd.n2314 vdd.n1183 19.3944
R20334 vdd.n2309 vdd.n1183 19.3944
R20335 vdd.n2309 vdd.n2308 19.3944
R20336 vdd.n2379 vdd.n1124 19.3944
R20337 vdd.n2379 vdd.n1125 19.3944
R20338 vdd.n2374 vdd.n2373 19.3944
R20339 vdd.n2369 vdd.n2368 19.3944
R20340 vdd.n2368 vdd.n2367 19.3944
R20341 vdd.n2367 vdd.n1129 19.3944
R20342 vdd.n2362 vdd.n1129 19.3944
R20343 vdd.n2362 vdd.n2361 19.3944
R20344 vdd.n2361 vdd.n2360 19.3944
R20345 vdd.n2360 vdd.n1136 19.3944
R20346 vdd.n2355 vdd.n1136 19.3944
R20347 vdd.n2355 vdd.n2354 19.3944
R20348 vdd.n2354 vdd.n2353 19.3944
R20349 vdd.n2353 vdd.n1143 19.3944
R20350 vdd.n2348 vdd.n1143 19.3944
R20351 vdd.n2348 vdd.n2347 19.3944
R20352 vdd.n1787 vdd.n1552 19.3944
R20353 vdd.n1787 vdd.n1543 19.3944
R20354 vdd.n1800 vdd.n1543 19.3944
R20355 vdd.n1800 vdd.n1541 19.3944
R20356 vdd.n1804 vdd.n1541 19.3944
R20357 vdd.n1804 vdd.n1532 19.3944
R20358 vdd.n1817 vdd.n1532 19.3944
R20359 vdd.n1817 vdd.n1530 19.3944
R20360 vdd.n1821 vdd.n1530 19.3944
R20361 vdd.n1821 vdd.n1521 19.3944
R20362 vdd.n1833 vdd.n1521 19.3944
R20363 vdd.n1833 vdd.n1519 19.3944
R20364 vdd.n1837 vdd.n1519 19.3944
R20365 vdd.n1837 vdd.n1509 19.3944
R20366 vdd.n1850 vdd.n1509 19.3944
R20367 vdd.n1850 vdd.n1507 19.3944
R20368 vdd.n1854 vdd.n1507 19.3944
R20369 vdd.n1854 vdd.n1498 19.3944
R20370 vdd.n1866 vdd.n1498 19.3944
R20371 vdd.n1866 vdd.n1496 19.3944
R20372 vdd.n2177 vdd.n1496 19.3944
R20373 vdd.n2177 vdd.n1486 19.3944
R20374 vdd.n2190 vdd.n1486 19.3944
R20375 vdd.n2190 vdd.n1484 19.3944
R20376 vdd.n2194 vdd.n1484 19.3944
R20377 vdd.n2194 vdd.n1475 19.3944
R20378 vdd.n2207 vdd.n1475 19.3944
R20379 vdd.n2207 vdd.n1473 19.3944
R20380 vdd.n2211 vdd.n1473 19.3944
R20381 vdd.n2211 vdd.n1464 19.3944
R20382 vdd.n2223 vdd.n1464 19.3944
R20383 vdd.n2223 vdd.n1462 19.3944
R20384 vdd.n2227 vdd.n1462 19.3944
R20385 vdd.n2227 vdd.n1452 19.3944
R20386 vdd.n2240 vdd.n1452 19.3944
R20387 vdd.n2240 vdd.n1450 19.3944
R20388 vdd.n2244 vdd.n1450 19.3944
R20389 vdd.n2244 vdd.n1440 19.3944
R20390 vdd.n2259 vdd.n1440 19.3944
R20391 vdd.n2259 vdd.n1438 19.3944
R20392 vdd.n2263 vdd.n1438 19.3944
R20393 vdd.n3321 vdd.n686 19.3944
R20394 vdd.n3321 vdd.n676 19.3944
R20395 vdd.n3333 vdd.n676 19.3944
R20396 vdd.n3333 vdd.n674 19.3944
R20397 vdd.n3337 vdd.n674 19.3944
R20398 vdd.n3337 vdd.n666 19.3944
R20399 vdd.n3350 vdd.n666 19.3944
R20400 vdd.n3350 vdd.n664 19.3944
R20401 vdd.n3354 vdd.n664 19.3944
R20402 vdd.n3354 vdd.n653 19.3944
R20403 vdd.n3366 vdd.n653 19.3944
R20404 vdd.n3366 vdd.n651 19.3944
R20405 vdd.n3370 vdd.n651 19.3944
R20406 vdd.n3370 vdd.n642 19.3944
R20407 vdd.n3383 vdd.n642 19.3944
R20408 vdd.n3383 vdd.n640 19.3944
R20409 vdd.n3390 vdd.n640 19.3944
R20410 vdd.n3390 vdd.n3389 19.3944
R20411 vdd.n3389 vdd.n631 19.3944
R20412 vdd.n3403 vdd.n631 19.3944
R20413 vdd.n3404 vdd.n3403 19.3944
R20414 vdd.n3404 vdd.n629 19.3944
R20415 vdd.n3408 vdd.n629 19.3944
R20416 vdd.n3410 vdd.n3408 19.3944
R20417 vdd.n3411 vdd.n3410 19.3944
R20418 vdd.n3411 vdd.n627 19.3944
R20419 vdd.n3415 vdd.n627 19.3944
R20420 vdd.n3417 vdd.n3415 19.3944
R20421 vdd.n3418 vdd.n3417 19.3944
R20422 vdd.n3418 vdd.n625 19.3944
R20423 vdd.n3422 vdd.n625 19.3944
R20424 vdd.n3425 vdd.n3422 19.3944
R20425 vdd.n3426 vdd.n3425 19.3944
R20426 vdd.n3426 vdd.n623 19.3944
R20427 vdd.n3430 vdd.n623 19.3944
R20428 vdd.n3432 vdd.n3430 19.3944
R20429 vdd.n3433 vdd.n3432 19.3944
R20430 vdd.n3433 vdd.n621 19.3944
R20431 vdd.n3437 vdd.n621 19.3944
R20432 vdd.n3439 vdd.n3437 19.3944
R20433 vdd.n3440 vdd.n3439 19.3944
R20434 vdd.n569 vdd.n438 19.3944
R20435 vdd.n575 vdd.n438 19.3944
R20436 vdd.n576 vdd.n575 19.3944
R20437 vdd.n579 vdd.n576 19.3944
R20438 vdd.n579 vdd.n436 19.3944
R20439 vdd.n585 vdd.n436 19.3944
R20440 vdd.n586 vdd.n585 19.3944
R20441 vdd.n589 vdd.n586 19.3944
R20442 vdd.n589 vdd.n434 19.3944
R20443 vdd.n595 vdd.n434 19.3944
R20444 vdd.n596 vdd.n595 19.3944
R20445 vdd.n599 vdd.n596 19.3944
R20446 vdd.n599 vdd.n432 19.3944
R20447 vdd.n605 vdd.n432 19.3944
R20448 vdd.n606 vdd.n605 19.3944
R20449 vdd.n609 vdd.n606 19.3944
R20450 vdd.n609 vdd.n430 19.3944
R20451 vdd.n615 vdd.n430 19.3944
R20452 vdd.n617 vdd.n615 19.3944
R20453 vdd.n618 vdd.n617 19.3944
R20454 vdd.n516 vdd.n515 19.3944
R20455 vdd.n519 vdd.n516 19.3944
R20456 vdd.n519 vdd.n450 19.3944
R20457 vdd.n525 vdd.n450 19.3944
R20458 vdd.n526 vdd.n525 19.3944
R20459 vdd.n529 vdd.n526 19.3944
R20460 vdd.n529 vdd.n448 19.3944
R20461 vdd.n535 vdd.n448 19.3944
R20462 vdd.n536 vdd.n535 19.3944
R20463 vdd.n539 vdd.n536 19.3944
R20464 vdd.n539 vdd.n446 19.3944
R20465 vdd.n545 vdd.n446 19.3944
R20466 vdd.n546 vdd.n545 19.3944
R20467 vdd.n549 vdd.n546 19.3944
R20468 vdd.n549 vdd.n444 19.3944
R20469 vdd.n555 vdd.n444 19.3944
R20470 vdd.n556 vdd.n555 19.3944
R20471 vdd.n559 vdd.n556 19.3944
R20472 vdd.n559 vdd.n442 19.3944
R20473 vdd.n565 vdd.n442 19.3944
R20474 vdd.n466 vdd.n465 19.3944
R20475 vdd.n469 vdd.n466 19.3944
R20476 vdd.n469 vdd.n462 19.3944
R20477 vdd.n475 vdd.n462 19.3944
R20478 vdd.n476 vdd.n475 19.3944
R20479 vdd.n479 vdd.n476 19.3944
R20480 vdd.n479 vdd.n460 19.3944
R20481 vdd.n485 vdd.n460 19.3944
R20482 vdd.n486 vdd.n485 19.3944
R20483 vdd.n489 vdd.n486 19.3944
R20484 vdd.n489 vdd.n458 19.3944
R20485 vdd.n495 vdd.n458 19.3944
R20486 vdd.n496 vdd.n495 19.3944
R20487 vdd.n499 vdd.n496 19.3944
R20488 vdd.n499 vdd.n456 19.3944
R20489 vdd.n505 vdd.n456 19.3944
R20490 vdd.n506 vdd.n505 19.3944
R20491 vdd.n509 vdd.n506 19.3944
R20492 vdd.n3325 vdd.n683 19.3944
R20493 vdd.n3325 vdd.n681 19.3944
R20494 vdd.n3329 vdd.n681 19.3944
R20495 vdd.n3329 vdd.n671 19.3944
R20496 vdd.n3342 vdd.n671 19.3944
R20497 vdd.n3342 vdd.n669 19.3944
R20498 vdd.n3346 vdd.n669 19.3944
R20499 vdd.n3346 vdd.n660 19.3944
R20500 vdd.n3358 vdd.n660 19.3944
R20501 vdd.n3358 vdd.n658 19.3944
R20502 vdd.n3362 vdd.n658 19.3944
R20503 vdd.n3362 vdd.n648 19.3944
R20504 vdd.n3375 vdd.n648 19.3944
R20505 vdd.n3375 vdd.n646 19.3944
R20506 vdd.n3379 vdd.n646 19.3944
R20507 vdd.n3379 vdd.n637 19.3944
R20508 vdd.n3394 vdd.n637 19.3944
R20509 vdd.n3394 vdd.n635 19.3944
R20510 vdd.n3398 vdd.n635 19.3944
R20511 vdd.n3398 vdd.n336 19.3944
R20512 vdd.n3489 vdd.n336 19.3944
R20513 vdd.n3489 vdd.n337 19.3944
R20514 vdd.n3483 vdd.n337 19.3944
R20515 vdd.n3483 vdd.n3482 19.3944
R20516 vdd.n3482 vdd.n3481 19.3944
R20517 vdd.n3481 vdd.n349 19.3944
R20518 vdd.n3475 vdd.n349 19.3944
R20519 vdd.n3475 vdd.n3474 19.3944
R20520 vdd.n3474 vdd.n3473 19.3944
R20521 vdd.n3473 vdd.n359 19.3944
R20522 vdd.n3467 vdd.n359 19.3944
R20523 vdd.n3467 vdd.n3466 19.3944
R20524 vdd.n3466 vdd.n3465 19.3944
R20525 vdd.n3465 vdd.n370 19.3944
R20526 vdd.n3459 vdd.n370 19.3944
R20527 vdd.n3459 vdd.n3458 19.3944
R20528 vdd.n3458 vdd.n3457 19.3944
R20529 vdd.n3457 vdd.n381 19.3944
R20530 vdd.n3451 vdd.n381 19.3944
R20531 vdd.n3451 vdd.n3450 19.3944
R20532 vdd.n3450 vdd.n3449 19.3944
R20533 vdd.n3272 vdd.n747 19.3944
R20534 vdd.n3272 vdd.n3269 19.3944
R20535 vdd.n3269 vdd.n3266 19.3944
R20536 vdd.n3266 vdd.n3265 19.3944
R20537 vdd.n3265 vdd.n3262 19.3944
R20538 vdd.n3262 vdd.n3261 19.3944
R20539 vdd.n3261 vdd.n3258 19.3944
R20540 vdd.n3258 vdd.n3257 19.3944
R20541 vdd.n3257 vdd.n3254 19.3944
R20542 vdd.n3254 vdd.n3253 19.3944
R20543 vdd.n3253 vdd.n3250 19.3944
R20544 vdd.n3250 vdd.n3249 19.3944
R20545 vdd.n3249 vdd.n3246 19.3944
R20546 vdd.n3246 vdd.n3245 19.3944
R20547 vdd.n3245 vdd.n3242 19.3944
R20548 vdd.n3242 vdd.n3241 19.3944
R20549 vdd.n3241 vdd.n3238 19.3944
R20550 vdd.n3238 vdd.n3237 19.3944
R20551 vdd.n3237 vdd.n3234 19.3944
R20552 vdd.n3234 vdd.n3233 19.3944
R20553 vdd.n3312 vdd.n3311 19.3944
R20554 vdd.n3311 vdd.n3310 19.3944
R20555 vdd.n732 vdd.n729 19.3944
R20556 vdd.n3306 vdd.n3305 19.3944
R20557 vdd.n3305 vdd.n3302 19.3944
R20558 vdd.n3302 vdd.n3301 19.3944
R20559 vdd.n3301 vdd.n3298 19.3944
R20560 vdd.n3298 vdd.n3297 19.3944
R20561 vdd.n3297 vdd.n3294 19.3944
R20562 vdd.n3294 vdd.n3293 19.3944
R20563 vdd.n3293 vdd.n3290 19.3944
R20564 vdd.n3290 vdd.n3289 19.3944
R20565 vdd.n3289 vdd.n3286 19.3944
R20566 vdd.n3286 vdd.n3285 19.3944
R20567 vdd.n3285 vdd.n3282 19.3944
R20568 vdd.n3282 vdd.n3281 19.3944
R20569 vdd.n3226 vdd.n767 19.3944
R20570 vdd.n3226 vdd.n3223 19.3944
R20571 vdd.n3223 vdd.n3220 19.3944
R20572 vdd.n3220 vdd.n3219 19.3944
R20573 vdd.n3219 vdd.n3216 19.3944
R20574 vdd.n3216 vdd.n3215 19.3944
R20575 vdd.n3215 vdd.n3212 19.3944
R20576 vdd.n3212 vdd.n3211 19.3944
R20577 vdd.n3211 vdd.n3208 19.3944
R20578 vdd.n3208 vdd.n3207 19.3944
R20579 vdd.n3207 vdd.n3204 19.3944
R20580 vdd.n3204 vdd.n3203 19.3944
R20581 vdd.n3203 vdd.n3200 19.3944
R20582 vdd.n3200 vdd.n3199 19.3944
R20583 vdd.n3199 vdd.n3196 19.3944
R20584 vdd.n3196 vdd.n3195 19.3944
R20585 vdd.n3192 vdd.n3191 19.3944
R20586 vdd.n3188 vdd.n3187 19.3944
R20587 vdd.n1719 vdd.n1715 19.0066
R20588 vdd.n2307 vdd.n1189 19.0066
R20589 vdd.n569 vdd.n566 19.0066
R20590 vdd.n3230 vdd.n767 19.0066
R20591 vdd.n1254 vdd.n1253 16.0975
R20592 vdd.n982 vdd.n981 16.0975
R20593 vdd.n1680 vdd.n1679 16.0975
R20594 vdd.n1718 vdd.n1717 16.0975
R20595 vdd.n1614 vdd.n1613 16.0975
R20596 vdd.n2270 vdd.n2269 16.0975
R20597 vdd.n1191 vdd.n1190 16.0975
R20598 vdd.n1151 vdd.n1150 16.0975
R20599 vdd.n1274 vdd.n1273 16.0975
R20600 vdd.n973 vdd.n972 16.0975
R20601 vdd.n2705 vdd.n2704 16.0975
R20602 vdd.n427 vdd.n426 16.0975
R20603 vdd.n441 vdd.n440 16.0975
R20604 vdd.n453 vdd.n452 16.0975
R20605 vdd.n769 vdd.n768 16.0975
R20606 vdd.n3277 vdd.n3276 16.0975
R20607 vdd.n833 vdd.n832 16.0975
R20608 vdd.n2702 vdd.n2701 16.0975
R20609 vdd.n689 vdd.n688 16.0975
R20610 vdd.n800 vdd.n799 16.0975
R20611 vdd.t136 vdd.n2665 15.4182
R20612 vdd.n2938 vdd.t130 15.4182
R20613 vdd.n28 vdd.n27 14.8572
R20614 vdd.n2417 vdd.n1076 14.0578
R20615 vdd.n3151 vdd.n692 14.0578
R20616 vdd.n328 vdd.n293 13.1884
R20617 vdd.n269 vdd.n234 13.1884
R20618 vdd.n226 vdd.n191 13.1884
R20619 vdd.n167 vdd.n132 13.1884
R20620 vdd.n125 vdd.n90 13.1884
R20621 vdd.n66 vdd.n31 13.1884
R20622 vdd.n2109 vdd.n2074 13.1884
R20623 vdd.n2168 vdd.n2133 13.1884
R20624 vdd.n2007 vdd.n1972 13.1884
R20625 vdd.n2066 vdd.n2031 13.1884
R20626 vdd.n1906 vdd.n1871 13.1884
R20627 vdd.n1965 vdd.n1930 13.1884
R20628 vdd.n1750 vdd.n1615 12.9944
R20629 vdd.n1754 vdd.n1615 12.9944
R20630 vdd.n2346 vdd.n1149 12.9944
R20631 vdd.n2347 vdd.n2346 12.9944
R20632 vdd.n515 vdd.n454 12.9944
R20633 vdd.n509 vdd.n454 12.9944
R20634 vdd.n3278 vdd.n747 12.9944
R20635 vdd.n3281 vdd.n3278 12.9944
R20636 vdd.n329 vdd.n291 12.8005
R20637 vdd.n324 vdd.n295 12.8005
R20638 vdd.n270 vdd.n232 12.8005
R20639 vdd.n265 vdd.n236 12.8005
R20640 vdd.n227 vdd.n189 12.8005
R20641 vdd.n222 vdd.n193 12.8005
R20642 vdd.n168 vdd.n130 12.8005
R20643 vdd.n163 vdd.n134 12.8005
R20644 vdd.n126 vdd.n88 12.8005
R20645 vdd.n121 vdd.n92 12.8005
R20646 vdd.n67 vdd.n29 12.8005
R20647 vdd.n62 vdd.n33 12.8005
R20648 vdd.n2110 vdd.n2072 12.8005
R20649 vdd.n2105 vdd.n2076 12.8005
R20650 vdd.n2169 vdd.n2131 12.8005
R20651 vdd.n2164 vdd.n2135 12.8005
R20652 vdd.n2008 vdd.n1970 12.8005
R20653 vdd.n2003 vdd.n1974 12.8005
R20654 vdd.n2067 vdd.n2029 12.8005
R20655 vdd.n2062 vdd.n2033 12.8005
R20656 vdd.n1907 vdd.n1869 12.8005
R20657 vdd.n1902 vdd.n1873 12.8005
R20658 vdd.n1966 vdd.n1928 12.8005
R20659 vdd.n1961 vdd.n1932 12.8005
R20660 vdd.n323 vdd.n296 12.0247
R20661 vdd.n264 vdd.n237 12.0247
R20662 vdd.n221 vdd.n194 12.0247
R20663 vdd.n162 vdd.n135 12.0247
R20664 vdd.n120 vdd.n93 12.0247
R20665 vdd.n61 vdd.n34 12.0247
R20666 vdd.n2104 vdd.n2077 12.0247
R20667 vdd.n2163 vdd.n2136 12.0247
R20668 vdd.n2002 vdd.n1975 12.0247
R20669 vdd.n2061 vdd.n2034 12.0247
R20670 vdd.n1901 vdd.n1874 12.0247
R20671 vdd.n1960 vdd.n1933 12.0247
R20672 vdd.n1789 vdd.n1545 11.337
R20673 vdd.n1798 vdd.n1545 11.337
R20674 vdd.n1798 vdd.n1797 11.337
R20675 vdd.n1806 vdd.n1539 11.337
R20676 vdd.n1815 vdd.n1814 11.337
R20677 vdd.n1831 vdd.n1523 11.337
R20678 vdd.n1839 vdd.n1516 11.337
R20679 vdd.n1848 vdd.n1847 11.337
R20680 vdd.n1856 vdd.n1505 11.337
R20681 vdd.n2179 vdd.n1494 11.337
R20682 vdd.n2188 vdd.n1488 11.337
R20683 vdd.n2196 vdd.n1482 11.337
R20684 vdd.n2205 vdd.n2204 11.337
R20685 vdd.n2221 vdd.n1466 11.337
R20686 vdd.n2229 vdd.n1459 11.337
R20687 vdd.n2238 vdd.n2237 11.337
R20688 vdd.n2246 vdd.n1442 11.337
R20689 vdd.n2257 vdd.n1442 11.337
R20690 vdd.n2257 vdd.n2256 11.337
R20691 vdd.n3323 vdd.n678 11.337
R20692 vdd.n3331 vdd.n678 11.337
R20693 vdd.n3331 vdd.n679 11.337
R20694 vdd.n3340 vdd.n3339 11.337
R20695 vdd.n3356 vdd.n662 11.337
R20696 vdd.n3364 vdd.n655 11.337
R20697 vdd.n3373 vdd.n3372 11.337
R20698 vdd.n3381 vdd.n644 11.337
R20699 vdd.n3400 vdd.n633 11.337
R20700 vdd.n3487 vdd.n340 11.337
R20701 vdd.n3485 vdd.n344 11.337
R20702 vdd.n3479 vdd.n3478 11.337
R20703 vdd.n3471 vdd.n361 11.337
R20704 vdd.n3470 vdd.n3469 11.337
R20705 vdd.n3463 vdd.n3462 11.337
R20706 vdd.n3461 vdd.n375 11.337
R20707 vdd.n3455 vdd.n3454 11.337
R20708 vdd.n3454 vdd.n3453 11.337
R20709 vdd.n3453 vdd.n386 11.337
R20710 vdd.n320 vdd.n319 11.249
R20711 vdd.n261 vdd.n260 11.249
R20712 vdd.n218 vdd.n217 11.249
R20713 vdd.n159 vdd.n158 11.249
R20714 vdd.n117 vdd.n116 11.249
R20715 vdd.n58 vdd.n57 11.249
R20716 vdd.n2101 vdd.n2100 11.249
R20717 vdd.n2160 vdd.n2159 11.249
R20718 vdd.n1999 vdd.n1998 11.249
R20719 vdd.n2058 vdd.n2057 11.249
R20720 vdd.n1898 vdd.n1897 11.249
R20721 vdd.n1957 vdd.n1956 11.249
R20722 vdd.n1587 vdd.t63 11.2237
R20723 vdd.n3447 vdd.t49 11.2237
R20724 vdd.t220 vdd.n1460 10.7702
R20725 vdd.n3348 vdd.t142 10.7702
R20726 vdd.n305 vdd.n304 10.7238
R20727 vdd.n246 vdd.n245 10.7238
R20728 vdd.n203 vdd.n202 10.7238
R20729 vdd.n144 vdd.n143 10.7238
R20730 vdd.n102 vdd.n101 10.7238
R20731 vdd.n43 vdd.n42 10.7238
R20732 vdd.n2086 vdd.n2085 10.7238
R20733 vdd.n2145 vdd.n2144 10.7238
R20734 vdd.n1984 vdd.n1983 10.7238
R20735 vdd.n2043 vdd.n2042 10.7238
R20736 vdd.n1883 vdd.n1882 10.7238
R20737 vdd.n1942 vdd.n1941 10.7238
R20738 vdd.n2593 vdd.t120 10.6568
R20739 vdd.t102 vdd.n928 10.6568
R20740 vdd.n2426 vdd.n1074 10.6151
R20741 vdd.n2427 vdd.n2426 10.6151
R20742 vdd.n2428 vdd.n2427 10.6151
R20743 vdd.n2428 vdd.n1063 10.6151
R20744 vdd.n2438 vdd.n1063 10.6151
R20745 vdd.n2439 vdd.n2438 10.6151
R20746 vdd.n2440 vdd.n2439 10.6151
R20747 vdd.n2440 vdd.n1050 10.6151
R20748 vdd.n2450 vdd.n1050 10.6151
R20749 vdd.n2451 vdd.n2450 10.6151
R20750 vdd.n2452 vdd.n2451 10.6151
R20751 vdd.n2452 vdd.n1038 10.6151
R20752 vdd.n2463 vdd.n1038 10.6151
R20753 vdd.n2464 vdd.n2463 10.6151
R20754 vdd.n2465 vdd.n2464 10.6151
R20755 vdd.n2465 vdd.n1026 10.6151
R20756 vdd.n2475 vdd.n1026 10.6151
R20757 vdd.n2476 vdd.n2475 10.6151
R20758 vdd.n2477 vdd.n2476 10.6151
R20759 vdd.n2477 vdd.n1014 10.6151
R20760 vdd.n2487 vdd.n1014 10.6151
R20761 vdd.n2488 vdd.n2487 10.6151
R20762 vdd.n2489 vdd.n2488 10.6151
R20763 vdd.n2489 vdd.n1003 10.6151
R20764 vdd.n2499 vdd.n1003 10.6151
R20765 vdd.n2500 vdd.n2499 10.6151
R20766 vdd.n2501 vdd.n2500 10.6151
R20767 vdd.n2501 vdd.n990 10.6151
R20768 vdd.n2513 vdd.n990 10.6151
R20769 vdd.n2514 vdd.n2513 10.6151
R20770 vdd.n2516 vdd.n2514 10.6151
R20771 vdd.n2516 vdd.n2515 10.6151
R20772 vdd.n2515 vdd.n971 10.6151
R20773 vdd.n2663 vdd.n2662 10.6151
R20774 vdd.n2662 vdd.n2661 10.6151
R20775 vdd.n2661 vdd.n2658 10.6151
R20776 vdd.n2658 vdd.n2657 10.6151
R20777 vdd.n2657 vdd.n2654 10.6151
R20778 vdd.n2654 vdd.n2653 10.6151
R20779 vdd.n2653 vdd.n2650 10.6151
R20780 vdd.n2650 vdd.n2649 10.6151
R20781 vdd.n2649 vdd.n2646 10.6151
R20782 vdd.n2646 vdd.n2645 10.6151
R20783 vdd.n2645 vdd.n2642 10.6151
R20784 vdd.n2642 vdd.n2641 10.6151
R20785 vdd.n2641 vdd.n2638 10.6151
R20786 vdd.n2638 vdd.n2637 10.6151
R20787 vdd.n2637 vdd.n2634 10.6151
R20788 vdd.n2634 vdd.n2633 10.6151
R20789 vdd.n2633 vdd.n2630 10.6151
R20790 vdd.n2630 vdd.n2629 10.6151
R20791 vdd.n2629 vdd.n2626 10.6151
R20792 vdd.n2626 vdd.n2625 10.6151
R20793 vdd.n2625 vdd.n2622 10.6151
R20794 vdd.n2622 vdd.n2621 10.6151
R20795 vdd.n2621 vdd.n2618 10.6151
R20796 vdd.n2618 vdd.n2617 10.6151
R20797 vdd.n2617 vdd.n2614 10.6151
R20798 vdd.n2614 vdd.n2613 10.6151
R20799 vdd.n2613 vdd.n2610 10.6151
R20800 vdd.n2610 vdd.n2609 10.6151
R20801 vdd.n2609 vdd.n2606 10.6151
R20802 vdd.n2606 vdd.n2605 10.6151
R20803 vdd.n2605 vdd.n2602 10.6151
R20804 vdd.n2600 vdd.n2597 10.6151
R20805 vdd.n2597 vdd.n2596 10.6151
R20806 vdd.n1311 vdd.n1310 10.6151
R20807 vdd.n1313 vdd.n1311 10.6151
R20808 vdd.n1314 vdd.n1313 10.6151
R20809 vdd.n1316 vdd.n1314 10.6151
R20810 vdd.n1317 vdd.n1316 10.6151
R20811 vdd.n1319 vdd.n1317 10.6151
R20812 vdd.n1320 vdd.n1319 10.6151
R20813 vdd.n1322 vdd.n1320 10.6151
R20814 vdd.n1323 vdd.n1322 10.6151
R20815 vdd.n1325 vdd.n1323 10.6151
R20816 vdd.n1326 vdd.n1325 10.6151
R20817 vdd.n1328 vdd.n1326 10.6151
R20818 vdd.n1329 vdd.n1328 10.6151
R20819 vdd.n1331 vdd.n1329 10.6151
R20820 vdd.n1332 vdd.n1331 10.6151
R20821 vdd.n1334 vdd.n1332 10.6151
R20822 vdd.n1335 vdd.n1334 10.6151
R20823 vdd.n1357 vdd.n1335 10.6151
R20824 vdd.n1357 vdd.n1356 10.6151
R20825 vdd.n1356 vdd.n1355 10.6151
R20826 vdd.n1355 vdd.n1353 10.6151
R20827 vdd.n1353 vdd.n1352 10.6151
R20828 vdd.n1352 vdd.n1350 10.6151
R20829 vdd.n1350 vdd.n1349 10.6151
R20830 vdd.n1349 vdd.n1347 10.6151
R20831 vdd.n1347 vdd.n1346 10.6151
R20832 vdd.n1346 vdd.n1344 10.6151
R20833 vdd.n1344 vdd.n1343 10.6151
R20834 vdd.n1343 vdd.n1341 10.6151
R20835 vdd.n1341 vdd.n1340 10.6151
R20836 vdd.n1340 vdd.n1337 10.6151
R20837 vdd.n1337 vdd.n1336 10.6151
R20838 vdd.n1336 vdd.n974 10.6151
R20839 vdd.n2414 vdd.n2413 10.6151
R20840 vdd.n2413 vdd.n2412 10.6151
R20841 vdd.n2412 vdd.n2411 10.6151
R20842 vdd.n2411 vdd.n2409 10.6151
R20843 vdd.n2409 vdd.n2406 10.6151
R20844 vdd.n2406 vdd.n2405 10.6151
R20845 vdd.n2405 vdd.n2402 10.6151
R20846 vdd.n2402 vdd.n2401 10.6151
R20847 vdd.n2401 vdd.n2398 10.6151
R20848 vdd.n2398 vdd.n2397 10.6151
R20849 vdd.n2397 vdd.n2394 10.6151
R20850 vdd.n2394 vdd.n2393 10.6151
R20851 vdd.n2393 vdd.n2390 10.6151
R20852 vdd.n2390 vdd.n2389 10.6151
R20853 vdd.n2389 vdd.n2386 10.6151
R20854 vdd.n2386 vdd.n2385 10.6151
R20855 vdd.n2385 vdd.n2382 10.6151
R20856 vdd.n2382 vdd.n1119 10.6151
R20857 vdd.n1277 vdd.n1119 10.6151
R20858 vdd.n1278 vdd.n1277 10.6151
R20859 vdd.n1281 vdd.n1278 10.6151
R20860 vdd.n1282 vdd.n1281 10.6151
R20861 vdd.n1285 vdd.n1282 10.6151
R20862 vdd.n1286 vdd.n1285 10.6151
R20863 vdd.n1289 vdd.n1286 10.6151
R20864 vdd.n1290 vdd.n1289 10.6151
R20865 vdd.n1293 vdd.n1290 10.6151
R20866 vdd.n1294 vdd.n1293 10.6151
R20867 vdd.n1297 vdd.n1294 10.6151
R20868 vdd.n1298 vdd.n1297 10.6151
R20869 vdd.n1301 vdd.n1298 10.6151
R20870 vdd.n1306 vdd.n1303 10.6151
R20871 vdd.n1307 vdd.n1306 10.6151
R20872 vdd.n2866 vdd.n2865 10.6151
R20873 vdd.n2865 vdd.n2864 10.6151
R20874 vdd.n2864 vdd.n2703 10.6151
R20875 vdd.n2808 vdd.n2703 10.6151
R20876 vdd.n2809 vdd.n2808 10.6151
R20877 vdd.n2811 vdd.n2809 10.6151
R20878 vdd.n2812 vdd.n2811 10.6151
R20879 vdd.n2814 vdd.n2812 10.6151
R20880 vdd.n2815 vdd.n2814 10.6151
R20881 vdd.n2845 vdd.n2815 10.6151
R20882 vdd.n2845 vdd.n2844 10.6151
R20883 vdd.n2844 vdd.n2843 10.6151
R20884 vdd.n2843 vdd.n2841 10.6151
R20885 vdd.n2841 vdd.n2840 10.6151
R20886 vdd.n2840 vdd.n2838 10.6151
R20887 vdd.n2838 vdd.n2837 10.6151
R20888 vdd.n2837 vdd.n2835 10.6151
R20889 vdd.n2835 vdd.n2834 10.6151
R20890 vdd.n2834 vdd.n2832 10.6151
R20891 vdd.n2832 vdd.n2831 10.6151
R20892 vdd.n2831 vdd.n2829 10.6151
R20893 vdd.n2829 vdd.n2828 10.6151
R20894 vdd.n2828 vdd.n2826 10.6151
R20895 vdd.n2826 vdd.n2825 10.6151
R20896 vdd.n2825 vdd.n2823 10.6151
R20897 vdd.n2823 vdd.n2822 10.6151
R20898 vdd.n2822 vdd.n2820 10.6151
R20899 vdd.n2820 vdd.n2819 10.6151
R20900 vdd.n2819 vdd.n2817 10.6151
R20901 vdd.n2817 vdd.n2816 10.6151
R20902 vdd.n2816 vdd.n836 10.6151
R20903 vdd.n3084 vdd.n836 10.6151
R20904 vdd.n3085 vdd.n3084 10.6151
R20905 vdd.n2935 vdd.n2934 10.6151
R20906 vdd.n2934 vdd.n2933 10.6151
R20907 vdd.n2933 vdd.n2932 10.6151
R20908 vdd.n2932 vdd.n2930 10.6151
R20909 vdd.n2930 vdd.n2927 10.6151
R20910 vdd.n2927 vdd.n2926 10.6151
R20911 vdd.n2926 vdd.n2923 10.6151
R20912 vdd.n2923 vdd.n2922 10.6151
R20913 vdd.n2922 vdd.n2919 10.6151
R20914 vdd.n2919 vdd.n2918 10.6151
R20915 vdd.n2918 vdd.n2915 10.6151
R20916 vdd.n2915 vdd.n2914 10.6151
R20917 vdd.n2914 vdd.n2911 10.6151
R20918 vdd.n2911 vdd.n2910 10.6151
R20919 vdd.n2910 vdd.n2907 10.6151
R20920 vdd.n2907 vdd.n2906 10.6151
R20921 vdd.n2906 vdd.n2903 10.6151
R20922 vdd.n2903 vdd.n2902 10.6151
R20923 vdd.n2902 vdd.n2899 10.6151
R20924 vdd.n2899 vdd.n2898 10.6151
R20925 vdd.n2898 vdd.n2895 10.6151
R20926 vdd.n2895 vdd.n2894 10.6151
R20927 vdd.n2894 vdd.n2891 10.6151
R20928 vdd.n2891 vdd.n2890 10.6151
R20929 vdd.n2890 vdd.n2887 10.6151
R20930 vdd.n2887 vdd.n2886 10.6151
R20931 vdd.n2886 vdd.n2883 10.6151
R20932 vdd.n2883 vdd.n2882 10.6151
R20933 vdd.n2882 vdd.n2879 10.6151
R20934 vdd.n2879 vdd.n2878 10.6151
R20935 vdd.n2878 vdd.n2875 10.6151
R20936 vdd.n2873 vdd.n2870 10.6151
R20937 vdd.n2870 vdd.n2869 10.6151
R20938 vdd.n2947 vdd.n926 10.6151
R20939 vdd.n2948 vdd.n2947 10.6151
R20940 vdd.n2949 vdd.n2948 10.6151
R20941 vdd.n2949 vdd.n915 10.6151
R20942 vdd.n2959 vdd.n915 10.6151
R20943 vdd.n2960 vdd.n2959 10.6151
R20944 vdd.n2961 vdd.n2960 10.6151
R20945 vdd.n2961 vdd.n903 10.6151
R20946 vdd.n2971 vdd.n903 10.6151
R20947 vdd.n2972 vdd.n2971 10.6151
R20948 vdd.n2973 vdd.n2972 10.6151
R20949 vdd.n2973 vdd.n891 10.6151
R20950 vdd.n2983 vdd.n891 10.6151
R20951 vdd.n2984 vdd.n2983 10.6151
R20952 vdd.n2985 vdd.n2984 10.6151
R20953 vdd.n2985 vdd.n880 10.6151
R20954 vdd.n2995 vdd.n880 10.6151
R20955 vdd.n2996 vdd.n2995 10.6151
R20956 vdd.n2997 vdd.n2996 10.6151
R20957 vdd.n2997 vdd.n866 10.6151
R20958 vdd.n3008 vdd.n866 10.6151
R20959 vdd.n3009 vdd.n3008 10.6151
R20960 vdd.n3010 vdd.n3009 10.6151
R20961 vdd.n3010 vdd.n855 10.6151
R20962 vdd.n3020 vdd.n855 10.6151
R20963 vdd.n3021 vdd.n3020 10.6151
R20964 vdd.n3022 vdd.n3021 10.6151
R20965 vdd.n3022 vdd.n841 10.6151
R20966 vdd.n3077 vdd.n841 10.6151
R20967 vdd.n3078 vdd.n3077 10.6151
R20968 vdd.n3079 vdd.n3078 10.6151
R20969 vdd.n3079 vdd.n810 10.6151
R20970 vdd.n3149 vdd.n810 10.6151
R20971 vdd.n3148 vdd.n3147 10.6151
R20972 vdd.n3147 vdd.n811 10.6151
R20973 vdd.n812 vdd.n811 10.6151
R20974 vdd.n3140 vdd.n812 10.6151
R20975 vdd.n3140 vdd.n3139 10.6151
R20976 vdd.n3139 vdd.n3138 10.6151
R20977 vdd.n3138 vdd.n814 10.6151
R20978 vdd.n3133 vdd.n814 10.6151
R20979 vdd.n3133 vdd.n3132 10.6151
R20980 vdd.n3132 vdd.n3131 10.6151
R20981 vdd.n3131 vdd.n817 10.6151
R20982 vdd.n3126 vdd.n817 10.6151
R20983 vdd.n3126 vdd.n3125 10.6151
R20984 vdd.n3125 vdd.n3124 10.6151
R20985 vdd.n3124 vdd.n820 10.6151
R20986 vdd.n3119 vdd.n820 10.6151
R20987 vdd.n3119 vdd.n731 10.6151
R20988 vdd.n3115 vdd.n731 10.6151
R20989 vdd.n3115 vdd.n3114 10.6151
R20990 vdd.n3114 vdd.n3113 10.6151
R20991 vdd.n3113 vdd.n823 10.6151
R20992 vdd.n3108 vdd.n823 10.6151
R20993 vdd.n3108 vdd.n3107 10.6151
R20994 vdd.n3107 vdd.n3106 10.6151
R20995 vdd.n3106 vdd.n826 10.6151
R20996 vdd.n3101 vdd.n826 10.6151
R20997 vdd.n3101 vdd.n3100 10.6151
R20998 vdd.n3100 vdd.n3099 10.6151
R20999 vdd.n3099 vdd.n829 10.6151
R21000 vdd.n3094 vdd.n829 10.6151
R21001 vdd.n3094 vdd.n3093 10.6151
R21002 vdd.n3091 vdd.n834 10.6151
R21003 vdd.n3086 vdd.n834 10.6151
R21004 vdd.n3067 vdd.n3028 10.6151
R21005 vdd.n3062 vdd.n3028 10.6151
R21006 vdd.n3062 vdd.n3061 10.6151
R21007 vdd.n3061 vdd.n3060 10.6151
R21008 vdd.n3060 vdd.n3030 10.6151
R21009 vdd.n3055 vdd.n3030 10.6151
R21010 vdd.n3055 vdd.n3054 10.6151
R21011 vdd.n3054 vdd.n3053 10.6151
R21012 vdd.n3053 vdd.n3033 10.6151
R21013 vdd.n3048 vdd.n3033 10.6151
R21014 vdd.n3048 vdd.n3047 10.6151
R21015 vdd.n3047 vdd.n3046 10.6151
R21016 vdd.n3046 vdd.n3036 10.6151
R21017 vdd.n3041 vdd.n3036 10.6151
R21018 vdd.n3041 vdd.n3040 10.6151
R21019 vdd.n3040 vdd.n785 10.6151
R21020 vdd.n3184 vdd.n785 10.6151
R21021 vdd.n3184 vdd.n786 10.6151
R21022 vdd.n788 vdd.n786 10.6151
R21023 vdd.n3177 vdd.n788 10.6151
R21024 vdd.n3177 vdd.n3176 10.6151
R21025 vdd.n3176 vdd.n3175 10.6151
R21026 vdd.n3175 vdd.n790 10.6151
R21027 vdd.n3170 vdd.n790 10.6151
R21028 vdd.n3170 vdd.n3169 10.6151
R21029 vdd.n3169 vdd.n3168 10.6151
R21030 vdd.n3168 vdd.n793 10.6151
R21031 vdd.n3163 vdd.n793 10.6151
R21032 vdd.n3163 vdd.n3162 10.6151
R21033 vdd.n3162 vdd.n3161 10.6151
R21034 vdd.n3161 vdd.n796 10.6151
R21035 vdd.n3156 vdd.n3155 10.6151
R21036 vdd.n3155 vdd.n3154 10.6151
R21037 vdd.n2774 vdd.n2773 10.6151
R21038 vdd.n2860 vdd.n2774 10.6151
R21039 vdd.n2860 vdd.n2859 10.6151
R21040 vdd.n2859 vdd.n2858 10.6151
R21041 vdd.n2858 vdd.n2856 10.6151
R21042 vdd.n2856 vdd.n2855 10.6151
R21043 vdd.n2855 vdd.n2853 10.6151
R21044 vdd.n2853 vdd.n2852 10.6151
R21045 vdd.n2852 vdd.n2850 10.6151
R21046 vdd.n2850 vdd.n2849 10.6151
R21047 vdd.n2849 vdd.n2806 10.6151
R21048 vdd.n2806 vdd.n2805 10.6151
R21049 vdd.n2805 vdd.n2803 10.6151
R21050 vdd.n2803 vdd.n2802 10.6151
R21051 vdd.n2802 vdd.n2800 10.6151
R21052 vdd.n2800 vdd.n2799 10.6151
R21053 vdd.n2799 vdd.n2797 10.6151
R21054 vdd.n2797 vdd.n2796 10.6151
R21055 vdd.n2796 vdd.n2794 10.6151
R21056 vdd.n2794 vdd.n2793 10.6151
R21057 vdd.n2793 vdd.n2791 10.6151
R21058 vdd.n2791 vdd.n2790 10.6151
R21059 vdd.n2790 vdd.n2788 10.6151
R21060 vdd.n2788 vdd.n2787 10.6151
R21061 vdd.n2787 vdd.n2785 10.6151
R21062 vdd.n2785 vdd.n2784 10.6151
R21063 vdd.n2784 vdd.n2782 10.6151
R21064 vdd.n2782 vdd.n2781 10.6151
R21065 vdd.n2781 vdd.n2779 10.6151
R21066 vdd.n2779 vdd.n2778 10.6151
R21067 vdd.n2778 vdd.n2776 10.6151
R21068 vdd.n2776 vdd.n2775 10.6151
R21069 vdd.n2775 vdd.n802 10.6151
R21070 vdd.n2941 vdd.n932 10.6151
R21071 vdd.n2708 vdd.n932 10.6151
R21072 vdd.n2709 vdd.n2708 10.6151
R21073 vdd.n2712 vdd.n2709 10.6151
R21074 vdd.n2713 vdd.n2712 10.6151
R21075 vdd.n2716 vdd.n2713 10.6151
R21076 vdd.n2717 vdd.n2716 10.6151
R21077 vdd.n2720 vdd.n2717 10.6151
R21078 vdd.n2721 vdd.n2720 10.6151
R21079 vdd.n2724 vdd.n2721 10.6151
R21080 vdd.n2725 vdd.n2724 10.6151
R21081 vdd.n2728 vdd.n2725 10.6151
R21082 vdd.n2729 vdd.n2728 10.6151
R21083 vdd.n2732 vdd.n2729 10.6151
R21084 vdd.n2733 vdd.n2732 10.6151
R21085 vdd.n2736 vdd.n2733 10.6151
R21086 vdd.n2737 vdd.n2736 10.6151
R21087 vdd.n2740 vdd.n2737 10.6151
R21088 vdd.n2741 vdd.n2740 10.6151
R21089 vdd.n2744 vdd.n2741 10.6151
R21090 vdd.n2745 vdd.n2744 10.6151
R21091 vdd.n2748 vdd.n2745 10.6151
R21092 vdd.n2749 vdd.n2748 10.6151
R21093 vdd.n2752 vdd.n2749 10.6151
R21094 vdd.n2753 vdd.n2752 10.6151
R21095 vdd.n2756 vdd.n2753 10.6151
R21096 vdd.n2757 vdd.n2756 10.6151
R21097 vdd.n2760 vdd.n2757 10.6151
R21098 vdd.n2761 vdd.n2760 10.6151
R21099 vdd.n2764 vdd.n2761 10.6151
R21100 vdd.n2765 vdd.n2764 10.6151
R21101 vdd.n2770 vdd.n2768 10.6151
R21102 vdd.n2771 vdd.n2770 10.6151
R21103 vdd.n2943 vdd.n2942 10.6151
R21104 vdd.n2943 vdd.n921 10.6151
R21105 vdd.n2953 vdd.n921 10.6151
R21106 vdd.n2954 vdd.n2953 10.6151
R21107 vdd.n2955 vdd.n2954 10.6151
R21108 vdd.n2955 vdd.n909 10.6151
R21109 vdd.n2965 vdd.n909 10.6151
R21110 vdd.n2966 vdd.n2965 10.6151
R21111 vdd.n2967 vdd.n2966 10.6151
R21112 vdd.n2967 vdd.n897 10.6151
R21113 vdd.n2977 vdd.n897 10.6151
R21114 vdd.n2978 vdd.n2977 10.6151
R21115 vdd.n2979 vdd.n2978 10.6151
R21116 vdd.n2979 vdd.n886 10.6151
R21117 vdd.n2989 vdd.n886 10.6151
R21118 vdd.n2990 vdd.n2989 10.6151
R21119 vdd.n2991 vdd.n2990 10.6151
R21120 vdd.n2991 vdd.n873 10.6151
R21121 vdd.n3001 vdd.n873 10.6151
R21122 vdd.n3002 vdd.n3001 10.6151
R21123 vdd.n3004 vdd.n861 10.6151
R21124 vdd.n3014 vdd.n861 10.6151
R21125 vdd.n3015 vdd.n3014 10.6151
R21126 vdd.n3016 vdd.n3015 10.6151
R21127 vdd.n3016 vdd.n849 10.6151
R21128 vdd.n3026 vdd.n849 10.6151
R21129 vdd.n3027 vdd.n3026 10.6151
R21130 vdd.n3073 vdd.n3027 10.6151
R21131 vdd.n3073 vdd.n3072 10.6151
R21132 vdd.n3072 vdd.n3071 10.6151
R21133 vdd.n3071 vdd.n3070 10.6151
R21134 vdd.n3070 vdd.n3068 10.6151
R21135 vdd.n2422 vdd.n2421 10.6151
R21136 vdd.n2422 vdd.n1069 10.6151
R21137 vdd.n2432 vdd.n1069 10.6151
R21138 vdd.n2433 vdd.n2432 10.6151
R21139 vdd.n2434 vdd.n2433 10.6151
R21140 vdd.n2434 vdd.n1057 10.6151
R21141 vdd.n2444 vdd.n1057 10.6151
R21142 vdd.n2445 vdd.n2444 10.6151
R21143 vdd.n2446 vdd.n2445 10.6151
R21144 vdd.n2446 vdd.n1044 10.6151
R21145 vdd.n2456 vdd.n1044 10.6151
R21146 vdd.n2457 vdd.n2456 10.6151
R21147 vdd.n2459 vdd.n1032 10.6151
R21148 vdd.n2469 vdd.n1032 10.6151
R21149 vdd.n2470 vdd.n2469 10.6151
R21150 vdd.n2471 vdd.n2470 10.6151
R21151 vdd.n2471 vdd.n1020 10.6151
R21152 vdd.n2481 vdd.n1020 10.6151
R21153 vdd.n2482 vdd.n2481 10.6151
R21154 vdd.n2483 vdd.n2482 10.6151
R21155 vdd.n2483 vdd.n1009 10.6151
R21156 vdd.n2493 vdd.n1009 10.6151
R21157 vdd.n2494 vdd.n2493 10.6151
R21158 vdd.n2495 vdd.n2494 10.6151
R21159 vdd.n2495 vdd.n997 10.6151
R21160 vdd.n2505 vdd.n997 10.6151
R21161 vdd.n2506 vdd.n2505 10.6151
R21162 vdd.n2509 vdd.n2506 10.6151
R21163 vdd.n2509 vdd.n2508 10.6151
R21164 vdd.n2508 vdd.n2507 10.6151
R21165 vdd.n2507 vdd.n980 10.6151
R21166 vdd.n2591 vdd.n980 10.6151
R21167 vdd.n2590 vdd.n2589 10.6151
R21168 vdd.n2589 vdd.n2586 10.6151
R21169 vdd.n2586 vdd.n2585 10.6151
R21170 vdd.n2585 vdd.n2582 10.6151
R21171 vdd.n2582 vdd.n2581 10.6151
R21172 vdd.n2581 vdd.n2578 10.6151
R21173 vdd.n2578 vdd.n2577 10.6151
R21174 vdd.n2577 vdd.n2574 10.6151
R21175 vdd.n2574 vdd.n2573 10.6151
R21176 vdd.n2573 vdd.n2570 10.6151
R21177 vdd.n2570 vdd.n2569 10.6151
R21178 vdd.n2569 vdd.n2566 10.6151
R21179 vdd.n2566 vdd.n2565 10.6151
R21180 vdd.n2565 vdd.n2562 10.6151
R21181 vdd.n2562 vdd.n2561 10.6151
R21182 vdd.n2561 vdd.n2558 10.6151
R21183 vdd.n2558 vdd.n2557 10.6151
R21184 vdd.n2557 vdd.n2554 10.6151
R21185 vdd.n2554 vdd.n2553 10.6151
R21186 vdd.n2553 vdd.n2550 10.6151
R21187 vdd.n2550 vdd.n2549 10.6151
R21188 vdd.n2549 vdd.n2546 10.6151
R21189 vdd.n2546 vdd.n2545 10.6151
R21190 vdd.n2545 vdd.n2542 10.6151
R21191 vdd.n2542 vdd.n2541 10.6151
R21192 vdd.n2541 vdd.n2538 10.6151
R21193 vdd.n2538 vdd.n2537 10.6151
R21194 vdd.n2537 vdd.n2534 10.6151
R21195 vdd.n2534 vdd.n2533 10.6151
R21196 vdd.n2533 vdd.n2530 10.6151
R21197 vdd.n2530 vdd.n2529 10.6151
R21198 vdd.n2526 vdd.n2525 10.6151
R21199 vdd.n2525 vdd.n2523 10.6151
R21200 vdd.n1388 vdd.n1386 10.6151
R21201 vdd.n1386 vdd.n1385 10.6151
R21202 vdd.n1385 vdd.n1383 10.6151
R21203 vdd.n1383 vdd.n1382 10.6151
R21204 vdd.n1382 vdd.n1380 10.6151
R21205 vdd.n1380 vdd.n1379 10.6151
R21206 vdd.n1379 vdd.n1377 10.6151
R21207 vdd.n1377 vdd.n1376 10.6151
R21208 vdd.n1376 vdd.n1374 10.6151
R21209 vdd.n1374 vdd.n1373 10.6151
R21210 vdd.n1373 vdd.n1371 10.6151
R21211 vdd.n1371 vdd.n1370 10.6151
R21212 vdd.n1370 vdd.n1368 10.6151
R21213 vdd.n1368 vdd.n1367 10.6151
R21214 vdd.n1367 vdd.n1365 10.6151
R21215 vdd.n1365 vdd.n1364 10.6151
R21216 vdd.n1364 vdd.n1362 10.6151
R21217 vdd.n1362 vdd.n1361 10.6151
R21218 vdd.n1361 vdd.n1272 10.6151
R21219 vdd.n1272 vdd.n1271 10.6151
R21220 vdd.n1271 vdd.n1269 10.6151
R21221 vdd.n1269 vdd.n1268 10.6151
R21222 vdd.n1268 vdd.n1266 10.6151
R21223 vdd.n1266 vdd.n1265 10.6151
R21224 vdd.n1265 vdd.n1263 10.6151
R21225 vdd.n1263 vdd.n1262 10.6151
R21226 vdd.n1262 vdd.n1260 10.6151
R21227 vdd.n1260 vdd.n1259 10.6151
R21228 vdd.n1259 vdd.n1257 10.6151
R21229 vdd.n1257 vdd.n1256 10.6151
R21230 vdd.n1256 vdd.n984 10.6151
R21231 vdd.n2521 vdd.n984 10.6151
R21232 vdd.n2522 vdd.n2521 10.6151
R21233 vdd.n2420 vdd.n1081 10.6151
R21234 vdd.n1223 vdd.n1081 10.6151
R21235 vdd.n1224 vdd.n1223 10.6151
R21236 vdd.n1227 vdd.n1224 10.6151
R21237 vdd.n1228 vdd.n1227 10.6151
R21238 vdd.n1231 vdd.n1228 10.6151
R21239 vdd.n1232 vdd.n1231 10.6151
R21240 vdd.n1235 vdd.n1232 10.6151
R21241 vdd.n1236 vdd.n1235 10.6151
R21242 vdd.n1239 vdd.n1236 10.6151
R21243 vdd.n1240 vdd.n1239 10.6151
R21244 vdd.n1243 vdd.n1240 10.6151
R21245 vdd.n1244 vdd.n1243 10.6151
R21246 vdd.n1247 vdd.n1244 10.6151
R21247 vdd.n1248 vdd.n1247 10.6151
R21248 vdd.n1251 vdd.n1248 10.6151
R21249 vdd.n1422 vdd.n1251 10.6151
R21250 vdd.n1422 vdd.n1421 10.6151
R21251 vdd.n1421 vdd.n1419 10.6151
R21252 vdd.n1419 vdd.n1416 10.6151
R21253 vdd.n1416 vdd.n1415 10.6151
R21254 vdd.n1415 vdd.n1412 10.6151
R21255 vdd.n1412 vdd.n1411 10.6151
R21256 vdd.n1411 vdd.n1408 10.6151
R21257 vdd.n1408 vdd.n1407 10.6151
R21258 vdd.n1407 vdd.n1404 10.6151
R21259 vdd.n1404 vdd.n1403 10.6151
R21260 vdd.n1403 vdd.n1400 10.6151
R21261 vdd.n1400 vdd.n1399 10.6151
R21262 vdd.n1399 vdd.n1396 10.6151
R21263 vdd.n1396 vdd.n1395 10.6151
R21264 vdd.n1392 vdd.n1391 10.6151
R21265 vdd.n1391 vdd.n1389 10.6151
R21266 vdd.n2213 vdd.t156 10.5435
R21267 vdd.n656 vdd.t152 10.5435
R21268 vdd.n316 vdd.n298 10.4732
R21269 vdd.n257 vdd.n239 10.4732
R21270 vdd.n214 vdd.n196 10.4732
R21271 vdd.n155 vdd.n137 10.4732
R21272 vdd.n113 vdd.n95 10.4732
R21273 vdd.n54 vdd.n36 10.4732
R21274 vdd.n2097 vdd.n2079 10.4732
R21275 vdd.n2156 vdd.n2138 10.4732
R21276 vdd.n1995 vdd.n1977 10.4732
R21277 vdd.n2054 vdd.n2036 10.4732
R21278 vdd.n1894 vdd.n1876 10.4732
R21279 vdd.n1953 vdd.n1935 10.4732
R21280 vdd.t183 vdd.n2187 10.3167
R21281 vdd.n3392 vdd.t231 10.3167
R21282 vdd.n1864 vdd.t154 10.09
R21283 vdd.n3486 vdd.t170 10.09
R21284 vdd.t144 vdd.n1517 9.86327
R21285 vdd.n3477 vdd.t228 9.86327
R21286 vdd.n2382 vdd.n2381 9.78206
R21287 vdd.n3308 vdd.n731 9.78206
R21288 vdd.n3185 vdd.n3184 9.78206
R21289 vdd.n2274 vdd.n1422 9.78206
R21290 vdd.n315 vdd.n300 9.69747
R21291 vdd.n256 vdd.n241 9.69747
R21292 vdd.n213 vdd.n198 9.69747
R21293 vdd.n154 vdd.n139 9.69747
R21294 vdd.n112 vdd.n97 9.69747
R21295 vdd.n53 vdd.n38 9.69747
R21296 vdd.n2096 vdd.n2081 9.69747
R21297 vdd.n2155 vdd.n2140 9.69747
R21298 vdd.n1994 vdd.n1979 9.69747
R21299 vdd.n2053 vdd.n2038 9.69747
R21300 vdd.n1893 vdd.n1878 9.69747
R21301 vdd.n1952 vdd.n1937 9.69747
R21302 vdd.n1823 vdd.t236 9.63654
R21303 vdd.n3423 vdd.t200 9.63654
R21304 vdd.n331 vdd.n330 9.45567
R21305 vdd.n272 vdd.n271 9.45567
R21306 vdd.n229 vdd.n228 9.45567
R21307 vdd.n170 vdd.n169 9.45567
R21308 vdd.n128 vdd.n127 9.45567
R21309 vdd.n69 vdd.n68 9.45567
R21310 vdd.n2112 vdd.n2111 9.45567
R21311 vdd.n2171 vdd.n2170 9.45567
R21312 vdd.n2010 vdd.n2009 9.45567
R21313 vdd.n2069 vdd.n2068 9.45567
R21314 vdd.n1909 vdd.n1908 9.45567
R21315 vdd.n1968 vdd.n1967 9.45567
R21316 vdd.n1797 vdd.t196 9.40981
R21317 vdd.n3455 vdd.t160 9.40981
R21318 vdd.n2344 vdd.n1149 9.3005
R21319 vdd.n2343 vdd.n2342 9.3005
R21320 vdd.n1155 vdd.n1154 9.3005
R21321 vdd.n2337 vdd.n1159 9.3005
R21322 vdd.n2336 vdd.n1160 9.3005
R21323 vdd.n2335 vdd.n1161 9.3005
R21324 vdd.n1165 vdd.n1162 9.3005
R21325 vdd.n2330 vdd.n1166 9.3005
R21326 vdd.n2329 vdd.n1167 9.3005
R21327 vdd.n2328 vdd.n1168 9.3005
R21328 vdd.n1172 vdd.n1169 9.3005
R21329 vdd.n2323 vdd.n1173 9.3005
R21330 vdd.n2322 vdd.n1174 9.3005
R21331 vdd.n2321 vdd.n1175 9.3005
R21332 vdd.n1179 vdd.n1176 9.3005
R21333 vdd.n2316 vdd.n1180 9.3005
R21334 vdd.n2315 vdd.n1181 9.3005
R21335 vdd.n2314 vdd.n1182 9.3005
R21336 vdd.n1186 vdd.n1183 9.3005
R21337 vdd.n2309 vdd.n1187 9.3005
R21338 vdd.n2308 vdd.n1188 9.3005
R21339 vdd.n2307 vdd.n2306 9.3005
R21340 vdd.n2305 vdd.n1189 9.3005
R21341 vdd.n2304 vdd.n2303 9.3005
R21342 vdd.n1195 vdd.n1194 9.3005
R21343 vdd.n2298 vdd.n1199 9.3005
R21344 vdd.n2297 vdd.n1200 9.3005
R21345 vdd.n2296 vdd.n1201 9.3005
R21346 vdd.n1205 vdd.n1202 9.3005
R21347 vdd.n2291 vdd.n1206 9.3005
R21348 vdd.n2290 vdd.n1207 9.3005
R21349 vdd.n2289 vdd.n1208 9.3005
R21350 vdd.n1212 vdd.n1209 9.3005
R21351 vdd.n2284 vdd.n1213 9.3005
R21352 vdd.n2283 vdd.n1214 9.3005
R21353 vdd.n2282 vdd.n1215 9.3005
R21354 vdd.n1219 vdd.n1216 9.3005
R21355 vdd.n2277 vdd.n1220 9.3005
R21356 vdd.n2346 vdd.n2345 9.3005
R21357 vdd.n2368 vdd.n1120 9.3005
R21358 vdd.n2367 vdd.n1128 9.3005
R21359 vdd.n1132 vdd.n1129 9.3005
R21360 vdd.n2362 vdd.n1133 9.3005
R21361 vdd.n2361 vdd.n1134 9.3005
R21362 vdd.n2360 vdd.n1135 9.3005
R21363 vdd.n1139 vdd.n1136 9.3005
R21364 vdd.n2355 vdd.n1140 9.3005
R21365 vdd.n2354 vdd.n1141 9.3005
R21366 vdd.n2353 vdd.n1142 9.3005
R21367 vdd.n1146 vdd.n1143 9.3005
R21368 vdd.n2348 vdd.n1147 9.3005
R21369 vdd.n2347 vdd.n1148 9.3005
R21370 vdd.n2380 vdd.n2379 9.3005
R21371 vdd.n1124 vdd.n1123 9.3005
R21372 vdd.n2177 vdd.n2176 9.3005
R21373 vdd.n1486 vdd.n1485 9.3005
R21374 vdd.n2191 vdd.n2190 9.3005
R21375 vdd.n2192 vdd.n1484 9.3005
R21376 vdd.n2194 vdd.n2193 9.3005
R21377 vdd.n1475 vdd.n1474 9.3005
R21378 vdd.n2208 vdd.n2207 9.3005
R21379 vdd.n2209 vdd.n1473 9.3005
R21380 vdd.n2211 vdd.n2210 9.3005
R21381 vdd.n1464 vdd.n1463 9.3005
R21382 vdd.n2224 vdd.n2223 9.3005
R21383 vdd.n2225 vdd.n1462 9.3005
R21384 vdd.n2227 vdd.n2226 9.3005
R21385 vdd.n1452 vdd.n1451 9.3005
R21386 vdd.n2241 vdd.n2240 9.3005
R21387 vdd.n2242 vdd.n1450 9.3005
R21388 vdd.n2244 vdd.n2243 9.3005
R21389 vdd.n1440 vdd.n1439 9.3005
R21390 vdd.n2260 vdd.n2259 9.3005
R21391 vdd.n2261 vdd.n1438 9.3005
R21392 vdd.n2263 vdd.n2262 9.3005
R21393 vdd.n307 vdd.n306 9.3005
R21394 vdd.n302 vdd.n301 9.3005
R21395 vdd.n313 vdd.n312 9.3005
R21396 vdd.n315 vdd.n314 9.3005
R21397 vdd.n298 vdd.n297 9.3005
R21398 vdd.n321 vdd.n320 9.3005
R21399 vdd.n323 vdd.n322 9.3005
R21400 vdd.n295 vdd.n292 9.3005
R21401 vdd.n330 vdd.n329 9.3005
R21402 vdd.n248 vdd.n247 9.3005
R21403 vdd.n243 vdd.n242 9.3005
R21404 vdd.n254 vdd.n253 9.3005
R21405 vdd.n256 vdd.n255 9.3005
R21406 vdd.n239 vdd.n238 9.3005
R21407 vdd.n262 vdd.n261 9.3005
R21408 vdd.n264 vdd.n263 9.3005
R21409 vdd.n236 vdd.n233 9.3005
R21410 vdd.n271 vdd.n270 9.3005
R21411 vdd.n205 vdd.n204 9.3005
R21412 vdd.n200 vdd.n199 9.3005
R21413 vdd.n211 vdd.n210 9.3005
R21414 vdd.n213 vdd.n212 9.3005
R21415 vdd.n196 vdd.n195 9.3005
R21416 vdd.n219 vdd.n218 9.3005
R21417 vdd.n221 vdd.n220 9.3005
R21418 vdd.n193 vdd.n190 9.3005
R21419 vdd.n228 vdd.n227 9.3005
R21420 vdd.n146 vdd.n145 9.3005
R21421 vdd.n141 vdd.n140 9.3005
R21422 vdd.n152 vdd.n151 9.3005
R21423 vdd.n154 vdd.n153 9.3005
R21424 vdd.n137 vdd.n136 9.3005
R21425 vdd.n160 vdd.n159 9.3005
R21426 vdd.n162 vdd.n161 9.3005
R21427 vdd.n134 vdd.n131 9.3005
R21428 vdd.n169 vdd.n168 9.3005
R21429 vdd.n104 vdd.n103 9.3005
R21430 vdd.n99 vdd.n98 9.3005
R21431 vdd.n110 vdd.n109 9.3005
R21432 vdd.n112 vdd.n111 9.3005
R21433 vdd.n95 vdd.n94 9.3005
R21434 vdd.n118 vdd.n117 9.3005
R21435 vdd.n120 vdd.n119 9.3005
R21436 vdd.n92 vdd.n89 9.3005
R21437 vdd.n127 vdd.n126 9.3005
R21438 vdd.n45 vdd.n44 9.3005
R21439 vdd.n40 vdd.n39 9.3005
R21440 vdd.n51 vdd.n50 9.3005
R21441 vdd.n53 vdd.n52 9.3005
R21442 vdd.n36 vdd.n35 9.3005
R21443 vdd.n59 vdd.n58 9.3005
R21444 vdd.n61 vdd.n60 9.3005
R21445 vdd.n33 vdd.n30 9.3005
R21446 vdd.n68 vdd.n67 9.3005
R21447 vdd.n3230 vdd.n3229 9.3005
R21448 vdd.n3233 vdd.n766 9.3005
R21449 vdd.n3234 vdd.n765 9.3005
R21450 vdd.n3237 vdd.n764 9.3005
R21451 vdd.n3238 vdd.n763 9.3005
R21452 vdd.n3241 vdd.n762 9.3005
R21453 vdd.n3242 vdd.n761 9.3005
R21454 vdd.n3245 vdd.n760 9.3005
R21455 vdd.n3246 vdd.n759 9.3005
R21456 vdd.n3249 vdd.n758 9.3005
R21457 vdd.n3250 vdd.n757 9.3005
R21458 vdd.n3253 vdd.n756 9.3005
R21459 vdd.n3254 vdd.n755 9.3005
R21460 vdd.n3257 vdd.n754 9.3005
R21461 vdd.n3258 vdd.n753 9.3005
R21462 vdd.n3261 vdd.n752 9.3005
R21463 vdd.n3262 vdd.n751 9.3005
R21464 vdd.n3265 vdd.n750 9.3005
R21465 vdd.n3266 vdd.n749 9.3005
R21466 vdd.n3269 vdd.n748 9.3005
R21467 vdd.n3273 vdd.n3272 9.3005
R21468 vdd.n3274 vdd.n747 9.3005
R21469 vdd.n3278 vdd.n3275 9.3005
R21470 vdd.n3281 vdd.n746 9.3005
R21471 vdd.n3282 vdd.n745 9.3005
R21472 vdd.n3285 vdd.n744 9.3005
R21473 vdd.n3286 vdd.n743 9.3005
R21474 vdd.n3289 vdd.n742 9.3005
R21475 vdd.n3290 vdd.n741 9.3005
R21476 vdd.n3293 vdd.n740 9.3005
R21477 vdd.n3294 vdd.n739 9.3005
R21478 vdd.n3297 vdd.n738 9.3005
R21479 vdd.n3298 vdd.n737 9.3005
R21480 vdd.n3301 vdd.n736 9.3005
R21481 vdd.n3302 vdd.n735 9.3005
R21482 vdd.n3305 vdd.n730 9.3005
R21483 vdd.n3311 vdd.n727 9.3005
R21484 vdd.n3312 vdd.n726 9.3005
R21485 vdd.n3326 vdd.n3325 9.3005
R21486 vdd.n3327 vdd.n681 9.3005
R21487 vdd.n3329 vdd.n3328 9.3005
R21488 vdd.n671 vdd.n670 9.3005
R21489 vdd.n3343 vdd.n3342 9.3005
R21490 vdd.n3344 vdd.n669 9.3005
R21491 vdd.n3346 vdd.n3345 9.3005
R21492 vdd.n660 vdd.n659 9.3005
R21493 vdd.n3359 vdd.n3358 9.3005
R21494 vdd.n3360 vdd.n658 9.3005
R21495 vdd.n3362 vdd.n3361 9.3005
R21496 vdd.n648 vdd.n647 9.3005
R21497 vdd.n3376 vdd.n3375 9.3005
R21498 vdd.n3377 vdd.n646 9.3005
R21499 vdd.n3379 vdd.n3378 9.3005
R21500 vdd.n637 vdd.n636 9.3005
R21501 vdd.n3395 vdd.n3394 9.3005
R21502 vdd.n3396 vdd.n635 9.3005
R21503 vdd.n3398 vdd.n3397 9.3005
R21504 vdd.n336 vdd.n334 9.3005
R21505 vdd.n683 vdd.n682 9.3005
R21506 vdd.n3490 vdd.n3489 9.3005
R21507 vdd.n337 vdd.n335 9.3005
R21508 vdd.n3483 vdd.n346 9.3005
R21509 vdd.n3482 vdd.n347 9.3005
R21510 vdd.n3481 vdd.n348 9.3005
R21511 vdd.n355 vdd.n349 9.3005
R21512 vdd.n3475 vdd.n356 9.3005
R21513 vdd.n3474 vdd.n357 9.3005
R21514 vdd.n3473 vdd.n358 9.3005
R21515 vdd.n366 vdd.n359 9.3005
R21516 vdd.n3467 vdd.n367 9.3005
R21517 vdd.n3466 vdd.n368 9.3005
R21518 vdd.n3465 vdd.n369 9.3005
R21519 vdd.n377 vdd.n370 9.3005
R21520 vdd.n3459 vdd.n378 9.3005
R21521 vdd.n3458 vdd.n379 9.3005
R21522 vdd.n3457 vdd.n380 9.3005
R21523 vdd.n388 vdd.n381 9.3005
R21524 vdd.n3451 vdd.n389 9.3005
R21525 vdd.n3450 vdd.n390 9.3005
R21526 vdd.n3449 vdd.n391 9.3005
R21527 vdd.n466 vdd.n463 9.3005
R21528 vdd.n470 vdd.n469 9.3005
R21529 vdd.n471 vdd.n462 9.3005
R21530 vdd.n475 vdd.n472 9.3005
R21531 vdd.n476 vdd.n461 9.3005
R21532 vdd.n480 vdd.n479 9.3005
R21533 vdd.n481 vdd.n460 9.3005
R21534 vdd.n485 vdd.n482 9.3005
R21535 vdd.n486 vdd.n459 9.3005
R21536 vdd.n490 vdd.n489 9.3005
R21537 vdd.n491 vdd.n458 9.3005
R21538 vdd.n495 vdd.n492 9.3005
R21539 vdd.n496 vdd.n457 9.3005
R21540 vdd.n500 vdd.n499 9.3005
R21541 vdd.n501 vdd.n456 9.3005
R21542 vdd.n505 vdd.n502 9.3005
R21543 vdd.n506 vdd.n455 9.3005
R21544 vdd.n510 vdd.n509 9.3005
R21545 vdd.n511 vdd.n454 9.3005
R21546 vdd.n515 vdd.n512 9.3005
R21547 vdd.n516 vdd.n451 9.3005
R21548 vdd.n520 vdd.n519 9.3005
R21549 vdd.n521 vdd.n450 9.3005
R21550 vdd.n525 vdd.n522 9.3005
R21551 vdd.n526 vdd.n449 9.3005
R21552 vdd.n530 vdd.n529 9.3005
R21553 vdd.n531 vdd.n448 9.3005
R21554 vdd.n535 vdd.n532 9.3005
R21555 vdd.n536 vdd.n447 9.3005
R21556 vdd.n540 vdd.n539 9.3005
R21557 vdd.n541 vdd.n446 9.3005
R21558 vdd.n545 vdd.n542 9.3005
R21559 vdd.n546 vdd.n445 9.3005
R21560 vdd.n550 vdd.n549 9.3005
R21561 vdd.n551 vdd.n444 9.3005
R21562 vdd.n555 vdd.n552 9.3005
R21563 vdd.n556 vdd.n443 9.3005
R21564 vdd.n560 vdd.n559 9.3005
R21565 vdd.n561 vdd.n442 9.3005
R21566 vdd.n565 vdd.n562 9.3005
R21567 vdd.n566 vdd.n439 9.3005
R21568 vdd.n570 vdd.n569 9.3005
R21569 vdd.n571 vdd.n438 9.3005
R21570 vdd.n575 vdd.n572 9.3005
R21571 vdd.n576 vdd.n437 9.3005
R21572 vdd.n580 vdd.n579 9.3005
R21573 vdd.n581 vdd.n436 9.3005
R21574 vdd.n585 vdd.n582 9.3005
R21575 vdd.n586 vdd.n435 9.3005
R21576 vdd.n590 vdd.n589 9.3005
R21577 vdd.n591 vdd.n434 9.3005
R21578 vdd.n595 vdd.n592 9.3005
R21579 vdd.n596 vdd.n433 9.3005
R21580 vdd.n600 vdd.n599 9.3005
R21581 vdd.n601 vdd.n432 9.3005
R21582 vdd.n605 vdd.n602 9.3005
R21583 vdd.n606 vdd.n431 9.3005
R21584 vdd.n610 vdd.n609 9.3005
R21585 vdd.n611 vdd.n430 9.3005
R21586 vdd.n615 vdd.n612 9.3005
R21587 vdd.n617 vdd.n429 9.3005
R21588 vdd.n619 vdd.n618 9.3005
R21589 vdd.n3443 vdd.n3442 9.3005
R21590 vdd.n465 vdd.n464 9.3005
R21591 vdd.n3321 vdd.n3320 9.3005
R21592 vdd.n676 vdd.n675 9.3005
R21593 vdd.n3334 vdd.n3333 9.3005
R21594 vdd.n3335 vdd.n674 9.3005
R21595 vdd.n3337 vdd.n3336 9.3005
R21596 vdd.n666 vdd.n665 9.3005
R21597 vdd.n3351 vdd.n3350 9.3005
R21598 vdd.n3352 vdd.n664 9.3005
R21599 vdd.n3354 vdd.n3353 9.3005
R21600 vdd.n653 vdd.n652 9.3005
R21601 vdd.n3367 vdd.n3366 9.3005
R21602 vdd.n3368 vdd.n651 9.3005
R21603 vdd.n3370 vdd.n3369 9.3005
R21604 vdd.n642 vdd.n641 9.3005
R21605 vdd.n3384 vdd.n3383 9.3005
R21606 vdd.n3385 vdd.n640 9.3005
R21607 vdd.n3390 vdd.n3386 9.3005
R21608 vdd.n3389 vdd.n3388 9.3005
R21609 vdd.n3387 vdd.n631 9.3005
R21610 vdd.n3403 vdd.n630 9.3005
R21611 vdd.n3405 vdd.n3404 9.3005
R21612 vdd.n3406 vdd.n629 9.3005
R21613 vdd.n3408 vdd.n3407 9.3005
R21614 vdd.n3410 vdd.n628 9.3005
R21615 vdd.n3412 vdd.n3411 9.3005
R21616 vdd.n3413 vdd.n627 9.3005
R21617 vdd.n3415 vdd.n3414 9.3005
R21618 vdd.n3417 vdd.n626 9.3005
R21619 vdd.n3419 vdd.n3418 9.3005
R21620 vdd.n3420 vdd.n625 9.3005
R21621 vdd.n3422 vdd.n3421 9.3005
R21622 vdd.n3425 vdd.n624 9.3005
R21623 vdd.n3427 vdd.n3426 9.3005
R21624 vdd.n3428 vdd.n623 9.3005
R21625 vdd.n3430 vdd.n3429 9.3005
R21626 vdd.n3432 vdd.n622 9.3005
R21627 vdd.n3434 vdd.n3433 9.3005
R21628 vdd.n3435 vdd.n621 9.3005
R21629 vdd.n3437 vdd.n3436 9.3005
R21630 vdd.n3439 vdd.n620 9.3005
R21631 vdd.n3441 vdd.n3440 9.3005
R21632 vdd.n3319 vdd.n686 9.3005
R21633 vdd.n3318 vdd.n3317 9.3005
R21634 vdd.n3187 vdd.n687 9.3005
R21635 vdd.n3196 vdd.n783 9.3005
R21636 vdd.n3199 vdd.n782 9.3005
R21637 vdd.n3200 vdd.n781 9.3005
R21638 vdd.n3203 vdd.n780 9.3005
R21639 vdd.n3204 vdd.n779 9.3005
R21640 vdd.n3207 vdd.n778 9.3005
R21641 vdd.n3208 vdd.n777 9.3005
R21642 vdd.n3211 vdd.n776 9.3005
R21643 vdd.n3212 vdd.n775 9.3005
R21644 vdd.n3215 vdd.n774 9.3005
R21645 vdd.n3216 vdd.n773 9.3005
R21646 vdd.n3219 vdd.n772 9.3005
R21647 vdd.n3220 vdd.n771 9.3005
R21648 vdd.n3223 vdd.n770 9.3005
R21649 vdd.n3227 vdd.n3226 9.3005
R21650 vdd.n3228 vdd.n767 9.3005
R21651 vdd.n2273 vdd.n2272 9.3005
R21652 vdd.n2268 vdd.n1424 9.3005
R21653 vdd.n1792 vdd.n1791 9.3005
R21654 vdd.n1793 vdd.n1547 9.3005
R21655 vdd.n1795 vdd.n1794 9.3005
R21656 vdd.n1537 vdd.n1536 9.3005
R21657 vdd.n1809 vdd.n1808 9.3005
R21658 vdd.n1810 vdd.n1535 9.3005
R21659 vdd.n1812 vdd.n1811 9.3005
R21660 vdd.n1527 vdd.n1526 9.3005
R21661 vdd.n1826 vdd.n1825 9.3005
R21662 vdd.n1827 vdd.n1525 9.3005
R21663 vdd.n1829 vdd.n1828 9.3005
R21664 vdd.n1514 vdd.n1513 9.3005
R21665 vdd.n1842 vdd.n1841 9.3005
R21666 vdd.n1843 vdd.n1512 9.3005
R21667 vdd.n1845 vdd.n1844 9.3005
R21668 vdd.n1503 vdd.n1502 9.3005
R21669 vdd.n1859 vdd.n1858 9.3005
R21670 vdd.n1860 vdd.n1501 9.3005
R21671 vdd.n1862 vdd.n1861 9.3005
R21672 vdd.n1492 vdd.n1491 9.3005
R21673 vdd.n2182 vdd.n2181 9.3005
R21674 vdd.n2183 vdd.n1490 9.3005
R21675 vdd.n2185 vdd.n2184 9.3005
R21676 vdd.n1480 vdd.n1479 9.3005
R21677 vdd.n2199 vdd.n2198 9.3005
R21678 vdd.n2200 vdd.n1478 9.3005
R21679 vdd.n2202 vdd.n2201 9.3005
R21680 vdd.n1470 vdd.n1469 9.3005
R21681 vdd.n2216 vdd.n2215 9.3005
R21682 vdd.n2217 vdd.n1468 9.3005
R21683 vdd.n2219 vdd.n2218 9.3005
R21684 vdd.n1457 vdd.n1456 9.3005
R21685 vdd.n2232 vdd.n2231 9.3005
R21686 vdd.n2233 vdd.n1455 9.3005
R21687 vdd.n2235 vdd.n2234 9.3005
R21688 vdd.n1447 vdd.n1446 9.3005
R21689 vdd.n2249 vdd.n2248 9.3005
R21690 vdd.n2250 vdd.n1444 9.3005
R21691 vdd.n2254 vdd.n2253 9.3005
R21692 vdd.n2252 vdd.n1445 9.3005
R21693 vdd.n2251 vdd.n1435 9.3005
R21694 vdd.n1549 vdd.n1548 9.3005
R21695 vdd.n1685 vdd.n1684 9.3005
R21696 vdd.n1686 vdd.n1675 9.3005
R21697 vdd.n1688 vdd.n1687 9.3005
R21698 vdd.n1689 vdd.n1674 9.3005
R21699 vdd.n1691 vdd.n1690 9.3005
R21700 vdd.n1692 vdd.n1669 9.3005
R21701 vdd.n1694 vdd.n1693 9.3005
R21702 vdd.n1695 vdd.n1668 9.3005
R21703 vdd.n1697 vdd.n1696 9.3005
R21704 vdd.n1698 vdd.n1663 9.3005
R21705 vdd.n1700 vdd.n1699 9.3005
R21706 vdd.n1701 vdd.n1662 9.3005
R21707 vdd.n1703 vdd.n1702 9.3005
R21708 vdd.n1704 vdd.n1657 9.3005
R21709 vdd.n1706 vdd.n1705 9.3005
R21710 vdd.n1707 vdd.n1656 9.3005
R21711 vdd.n1709 vdd.n1708 9.3005
R21712 vdd.n1710 vdd.n1651 9.3005
R21713 vdd.n1712 vdd.n1711 9.3005
R21714 vdd.n1713 vdd.n1650 9.3005
R21715 vdd.n1715 vdd.n1714 9.3005
R21716 vdd.n1719 vdd.n1646 9.3005
R21717 vdd.n1721 vdd.n1720 9.3005
R21718 vdd.n1722 vdd.n1645 9.3005
R21719 vdd.n1724 vdd.n1723 9.3005
R21720 vdd.n1725 vdd.n1640 9.3005
R21721 vdd.n1727 vdd.n1726 9.3005
R21722 vdd.n1728 vdd.n1639 9.3005
R21723 vdd.n1730 vdd.n1729 9.3005
R21724 vdd.n1731 vdd.n1634 9.3005
R21725 vdd.n1733 vdd.n1732 9.3005
R21726 vdd.n1734 vdd.n1633 9.3005
R21727 vdd.n1736 vdd.n1735 9.3005
R21728 vdd.n1737 vdd.n1628 9.3005
R21729 vdd.n1739 vdd.n1738 9.3005
R21730 vdd.n1740 vdd.n1627 9.3005
R21731 vdd.n1742 vdd.n1741 9.3005
R21732 vdd.n1743 vdd.n1622 9.3005
R21733 vdd.n1745 vdd.n1744 9.3005
R21734 vdd.n1746 vdd.n1621 9.3005
R21735 vdd.n1748 vdd.n1747 9.3005
R21736 vdd.n1749 vdd.n1616 9.3005
R21737 vdd.n1751 vdd.n1750 9.3005
R21738 vdd.n1752 vdd.n1615 9.3005
R21739 vdd.n1754 vdd.n1753 9.3005
R21740 vdd.n1755 vdd.n1608 9.3005
R21741 vdd.n1757 vdd.n1756 9.3005
R21742 vdd.n1758 vdd.n1607 9.3005
R21743 vdd.n1760 vdd.n1759 9.3005
R21744 vdd.n1761 vdd.n1602 9.3005
R21745 vdd.n1763 vdd.n1762 9.3005
R21746 vdd.n1764 vdd.n1601 9.3005
R21747 vdd.n1766 vdd.n1765 9.3005
R21748 vdd.n1767 vdd.n1596 9.3005
R21749 vdd.n1769 vdd.n1768 9.3005
R21750 vdd.n1770 vdd.n1595 9.3005
R21751 vdd.n1772 vdd.n1771 9.3005
R21752 vdd.n1773 vdd.n1590 9.3005
R21753 vdd.n1775 vdd.n1774 9.3005
R21754 vdd.n1776 vdd.n1589 9.3005
R21755 vdd.n1778 vdd.n1777 9.3005
R21756 vdd.n1554 vdd.n1553 9.3005
R21757 vdd.n1784 vdd.n1783 9.3005
R21758 vdd.n1683 vdd.n1682 9.3005
R21759 vdd.n1787 vdd.n1786 9.3005
R21760 vdd.n1543 vdd.n1542 9.3005
R21761 vdd.n1801 vdd.n1800 9.3005
R21762 vdd.n1802 vdd.n1541 9.3005
R21763 vdd.n1804 vdd.n1803 9.3005
R21764 vdd.n1532 vdd.n1531 9.3005
R21765 vdd.n1818 vdd.n1817 9.3005
R21766 vdd.n1819 vdd.n1530 9.3005
R21767 vdd.n1821 vdd.n1820 9.3005
R21768 vdd.n1521 vdd.n1520 9.3005
R21769 vdd.n1834 vdd.n1833 9.3005
R21770 vdd.n1835 vdd.n1519 9.3005
R21771 vdd.n1837 vdd.n1836 9.3005
R21772 vdd.n1509 vdd.n1508 9.3005
R21773 vdd.n1851 vdd.n1850 9.3005
R21774 vdd.n1852 vdd.n1507 9.3005
R21775 vdd.n1854 vdd.n1853 9.3005
R21776 vdd.n1498 vdd.n1497 9.3005
R21777 vdd.n1867 vdd.n1866 9.3005
R21778 vdd.n1868 vdd.n1496 9.3005
R21779 vdd.n1785 vdd.n1552 9.3005
R21780 vdd.n2088 vdd.n2087 9.3005
R21781 vdd.n2083 vdd.n2082 9.3005
R21782 vdd.n2094 vdd.n2093 9.3005
R21783 vdd.n2096 vdd.n2095 9.3005
R21784 vdd.n2079 vdd.n2078 9.3005
R21785 vdd.n2102 vdd.n2101 9.3005
R21786 vdd.n2104 vdd.n2103 9.3005
R21787 vdd.n2076 vdd.n2073 9.3005
R21788 vdd.n2111 vdd.n2110 9.3005
R21789 vdd.n2147 vdd.n2146 9.3005
R21790 vdd.n2142 vdd.n2141 9.3005
R21791 vdd.n2153 vdd.n2152 9.3005
R21792 vdd.n2155 vdd.n2154 9.3005
R21793 vdd.n2138 vdd.n2137 9.3005
R21794 vdd.n2161 vdd.n2160 9.3005
R21795 vdd.n2163 vdd.n2162 9.3005
R21796 vdd.n2135 vdd.n2132 9.3005
R21797 vdd.n2170 vdd.n2169 9.3005
R21798 vdd.n1986 vdd.n1985 9.3005
R21799 vdd.n1981 vdd.n1980 9.3005
R21800 vdd.n1992 vdd.n1991 9.3005
R21801 vdd.n1994 vdd.n1993 9.3005
R21802 vdd.n1977 vdd.n1976 9.3005
R21803 vdd.n2000 vdd.n1999 9.3005
R21804 vdd.n2002 vdd.n2001 9.3005
R21805 vdd.n1974 vdd.n1971 9.3005
R21806 vdd.n2009 vdd.n2008 9.3005
R21807 vdd.n2045 vdd.n2044 9.3005
R21808 vdd.n2040 vdd.n2039 9.3005
R21809 vdd.n2051 vdd.n2050 9.3005
R21810 vdd.n2053 vdd.n2052 9.3005
R21811 vdd.n2036 vdd.n2035 9.3005
R21812 vdd.n2059 vdd.n2058 9.3005
R21813 vdd.n2061 vdd.n2060 9.3005
R21814 vdd.n2033 vdd.n2030 9.3005
R21815 vdd.n2068 vdd.n2067 9.3005
R21816 vdd.n1885 vdd.n1884 9.3005
R21817 vdd.n1880 vdd.n1879 9.3005
R21818 vdd.n1891 vdd.n1890 9.3005
R21819 vdd.n1893 vdd.n1892 9.3005
R21820 vdd.n1876 vdd.n1875 9.3005
R21821 vdd.n1899 vdd.n1898 9.3005
R21822 vdd.n1901 vdd.n1900 9.3005
R21823 vdd.n1873 vdd.n1870 9.3005
R21824 vdd.n1908 vdd.n1907 9.3005
R21825 vdd.n1944 vdd.n1943 9.3005
R21826 vdd.n1939 vdd.n1938 9.3005
R21827 vdd.n1950 vdd.n1949 9.3005
R21828 vdd.n1952 vdd.n1951 9.3005
R21829 vdd.n1935 vdd.n1934 9.3005
R21830 vdd.n1958 vdd.n1957 9.3005
R21831 vdd.n1960 vdd.n1959 9.3005
R21832 vdd.n1932 vdd.n1929 9.3005
R21833 vdd.n1967 vdd.n1966 9.3005
R21834 vdd.n1823 vdd.t210 9.18308
R21835 vdd.n3423 vdd.t146 9.18308
R21836 vdd.n1517 vdd.t181 8.95635
R21837 vdd.n2265 vdd.t39 8.95635
R21838 vdd.n723 vdd.t35 8.95635
R21839 vdd.t158 vdd.n3477 8.95635
R21840 vdd.n312 vdd.n311 8.92171
R21841 vdd.n253 vdd.n252 8.92171
R21842 vdd.n210 vdd.n209 8.92171
R21843 vdd.n151 vdd.n150 8.92171
R21844 vdd.n109 vdd.n108 8.92171
R21845 vdd.n50 vdd.n49 8.92171
R21846 vdd.n2093 vdd.n2092 8.92171
R21847 vdd.n2152 vdd.n2151 8.92171
R21848 vdd.n1991 vdd.n1990 8.92171
R21849 vdd.n2050 vdd.n2049 8.92171
R21850 vdd.n1890 vdd.n1889 8.92171
R21851 vdd.n1949 vdd.n1948 8.92171
R21852 vdd.n231 vdd.n129 8.81535
R21853 vdd.n2071 vdd.n1969 8.81535
R21854 vdd.n1864 vdd.t240 8.72962
R21855 vdd.t162 vdd.n3486 8.72962
R21856 vdd.n2187 vdd.t167 8.50289
R21857 vdd.n3392 vdd.t164 8.50289
R21858 vdd.n28 vdd.n14 8.42249
R21859 vdd.n2213 vdd.t243 8.27616
R21860 vdd.t204 vdd.n656 8.27616
R21861 vdd.n3492 vdd.n3491 8.16225
R21862 vdd.n2175 vdd.n2174 8.16225
R21863 vdd.n308 vdd.n302 8.14595
R21864 vdd.n249 vdd.n243 8.14595
R21865 vdd.n206 vdd.n200 8.14595
R21866 vdd.n147 vdd.n141 8.14595
R21867 vdd.n105 vdd.n99 8.14595
R21868 vdd.n46 vdd.n40 8.14595
R21869 vdd.n2089 vdd.n2083 8.14595
R21870 vdd.n2148 vdd.n2142 8.14595
R21871 vdd.n1987 vdd.n1981 8.14595
R21872 vdd.n2046 vdd.n2040 8.14595
R21873 vdd.n1886 vdd.n1880 8.14595
R21874 vdd.n1945 vdd.n1939 8.14595
R21875 vdd.n1460 vdd.t148 8.04943
R21876 vdd.n3348 vdd.t262 8.04943
R21877 vdd.n2424 vdd.n1076 7.70933
R21878 vdd.n2424 vdd.n1079 7.70933
R21879 vdd.n2430 vdd.n1065 7.70933
R21880 vdd.n2436 vdd.n1065 7.70933
R21881 vdd.n2436 vdd.n1059 7.70933
R21882 vdd.n2442 vdd.n1059 7.70933
R21883 vdd.n2448 vdd.n1052 7.70933
R21884 vdd.n2448 vdd.n1055 7.70933
R21885 vdd.n2454 vdd.n1048 7.70933
R21886 vdd.n2461 vdd.n1034 7.70933
R21887 vdd.n2467 vdd.n1034 7.70933
R21888 vdd.n2473 vdd.n1028 7.70933
R21889 vdd.n2479 vdd.n1024 7.70933
R21890 vdd.n2485 vdd.n1018 7.70933
R21891 vdd.n2497 vdd.n1005 7.70933
R21892 vdd.n2503 vdd.n999 7.70933
R21893 vdd.n2503 vdd.n992 7.70933
R21894 vdd.n2511 vdd.n992 7.70933
R21895 vdd.n2593 vdd.n976 7.70933
R21896 vdd.n2945 vdd.n928 7.70933
R21897 vdd.n2957 vdd.n917 7.70933
R21898 vdd.n2957 vdd.n911 7.70933
R21899 vdd.n2963 vdd.n911 7.70933
R21900 vdd.n2969 vdd.n905 7.70933
R21901 vdd.n2975 vdd.n901 7.70933
R21902 vdd.n2981 vdd.n895 7.70933
R21903 vdd.n2993 vdd.n882 7.70933
R21904 vdd.n2999 vdd.n875 7.70933
R21905 vdd.n2999 vdd.n878 7.70933
R21906 vdd.n3006 vdd.n870 7.70933
R21907 vdd.n3012 vdd.n857 7.70933
R21908 vdd.n3018 vdd.n857 7.70933
R21909 vdd.n3024 vdd.n851 7.70933
R21910 vdd.n3024 vdd.n843 7.70933
R21911 vdd.n3075 vdd.n843 7.70933
R21912 vdd.n3075 vdd.n846 7.70933
R21913 vdd.n3081 vdd.n805 7.70933
R21914 vdd.n3151 vdd.n805 7.70933
R21915 vdd.n3004 vdd.n3003 7.49318
R21916 vdd.n2458 vdd.n2457 7.49318
R21917 vdd.n307 vdd.n304 7.3702
R21918 vdd.n248 vdd.n245 7.3702
R21919 vdd.n205 vdd.n202 7.3702
R21920 vdd.n146 vdd.n143 7.3702
R21921 vdd.n104 vdd.n101 7.3702
R21922 vdd.n45 vdd.n42 7.3702
R21923 vdd.n2088 vdd.n2085 7.3702
R21924 vdd.n2147 vdd.n2144 7.3702
R21925 vdd.n1986 vdd.n1983 7.3702
R21926 vdd.n2045 vdd.n2042 7.3702
R21927 vdd.n1885 vdd.n1882 7.3702
R21928 vdd.n1944 vdd.n1941 7.3702
R21929 vdd.n2442 vdd.t18 7.36923
R21930 vdd.t114 vdd.n851 7.36923
R21931 vdd.n2518 vdd.t118 7.25587
R21932 vdd.n2862 vdd.t106 7.25587
R21933 vdd.n2246 vdd.t188 7.1425
R21934 vdd.n679 vdd.t186 7.1425
R21935 vdd.n1720 vdd.n1719 6.98232
R21936 vdd.n2308 vdd.n2307 6.98232
R21937 vdd.n566 vdd.n565 6.98232
R21938 vdd.n3233 vdd.n3230 6.98232
R21939 vdd.t256 vdd.n1459 6.91577
R21940 vdd.n3356 vdd.t202 6.91577
R21941 vdd.n2205 vdd.t208 6.68904
R21942 vdd.n3372 vdd.t191 6.68904
R21943 vdd.t238 vdd.n1488 6.46231
R21944 vdd.n3400 vdd.t194 6.46231
R21945 vdd.n3492 vdd.n333 6.38151
R21946 vdd.n2174 vdd.n2173 6.38151
R21947 vdd.n1856 vdd.t179 6.23558
R21948 vdd.t253 vdd.n344 6.23558
R21949 vdd.t150 vdd.n1516 6.00885
R21950 vdd.n3471 vdd.t213 6.00885
R21951 vdd.t128 vdd.n1005 5.89549
R21952 vdd.n2969 vdd.t110 5.89549
R21953 vdd.n308 vdd.n307 5.81868
R21954 vdd.n249 vdd.n248 5.81868
R21955 vdd.n206 vdd.n205 5.81868
R21956 vdd.n147 vdd.n146 5.81868
R21957 vdd.n105 vdd.n104 5.81868
R21958 vdd.n46 vdd.n45 5.81868
R21959 vdd.n2089 vdd.n2088 5.81868
R21960 vdd.n2148 vdd.n2147 5.81868
R21961 vdd.n1987 vdd.n1986 5.81868
R21962 vdd.n2046 vdd.n2045 5.81868
R21963 vdd.n1886 vdd.n1885 5.81868
R21964 vdd.n1945 vdd.n1944 5.81868
R21965 vdd.n1815 vdd.t140 5.78212
R21966 vdd.n3462 vdd.t259 5.78212
R21967 vdd.n2601 vdd.n2600 5.77611
R21968 vdd.n1303 vdd.n1302 5.77611
R21969 vdd.n2874 vdd.n2873 5.77611
R21970 vdd.n3092 vdd.n3091 5.77611
R21971 vdd.n3156 vdd.n801 5.77611
R21972 vdd.n2768 vdd.n2706 5.77611
R21973 vdd.n2526 vdd.n983 5.77611
R21974 vdd.n1392 vdd.n1255 5.77611
R21975 vdd.n1682 vdd.n1681 5.62474
R21976 vdd.n2271 vdd.n2268 5.62474
R21977 vdd.n3443 vdd.n428 5.62474
R21978 vdd.n3317 vdd.n690 5.62474
R21979 vdd.n1539 vdd.t140 5.55539
R21980 vdd.t124 vdd.n1028 5.55539
R21981 vdd.n2473 vdd.t19 5.55539
R21982 vdd.t25 vdd.n882 5.55539
R21983 vdd.n2993 vdd.t21 5.55539
R21984 vdd.t259 vdd.n3461 5.55539
R21985 vdd.n1048 vdd.t84 5.44203
R21986 vdd.n3006 vdd.t53 5.44203
R21987 vdd.n1831 vdd.t150 5.32866
R21988 vdd.n2430 vdd.t31 5.32866
R21989 vdd.n1338 vdd.t73 5.32866
R21990 vdd.n2951 vdd.t77 5.32866
R21991 vdd.n846 vdd.t27 5.32866
R21992 vdd.t213 vdd.n3470 5.32866
R21993 vdd.n1847 vdd.t179 5.10193
R21994 vdd.n3479 vdd.t253 5.10193
R21995 vdd.n311 vdd.n302 5.04292
R21996 vdd.n252 vdd.n243 5.04292
R21997 vdd.n209 vdd.n200 5.04292
R21998 vdd.n150 vdd.n141 5.04292
R21999 vdd.n108 vdd.n99 5.04292
R22000 vdd.n49 vdd.n40 5.04292
R22001 vdd.n2092 vdd.n2083 5.04292
R22002 vdd.n2151 vdd.n2142 5.04292
R22003 vdd.n1990 vdd.n1981 5.04292
R22004 vdd.n2049 vdd.n2040 5.04292
R22005 vdd.n1889 vdd.n1880 5.04292
R22006 vdd.n1948 vdd.n1939 5.04292
R22007 vdd.n2479 vdd.t112 4.98857
R22008 vdd.n895 vdd.t125 4.98857
R22009 vdd.n2179 vdd.t238 4.8752
R22010 vdd.t108 vdd.t134 4.8752
R22011 vdd.t20 vdd.t104 4.8752
R22012 vdd.t138 vdd.t127 4.8752
R22013 vdd.t23 vdd.t1 4.8752
R22014 vdd.t194 vdd.n340 4.8752
R22015 vdd.n2602 vdd.n2601 4.83952
R22016 vdd.n1302 vdd.n1301 4.83952
R22017 vdd.n2875 vdd.n2874 4.83952
R22018 vdd.n3093 vdd.n3092 4.83952
R22019 vdd.n801 vdd.n796 4.83952
R22020 vdd.n2765 vdd.n2706 4.83952
R22021 vdd.n2529 vdd.n983 4.83952
R22022 vdd.n1395 vdd.n1255 4.83952
R22023 vdd.n2276 vdd.n2275 4.74817
R22024 vdd.n1428 vdd.n1423 4.74817
R22025 vdd.n1125 vdd.n1122 4.74817
R22026 vdd.n2369 vdd.n1121 4.74817
R22027 vdd.n2374 vdd.n1122 4.74817
R22028 vdd.n2373 vdd.n1121 4.74817
R22029 vdd.n3310 vdd.n3309 4.74817
R22030 vdd.n3307 vdd.n3306 4.74817
R22031 vdd.n3307 vdd.n732 4.74817
R22032 vdd.n3309 vdd.n729 4.74817
R22033 vdd.n3192 vdd.n784 4.74817
R22034 vdd.n3188 vdd.n3186 4.74817
R22035 vdd.n3191 vdd.n3186 4.74817
R22036 vdd.n3195 vdd.n784 4.74817
R22037 vdd.n2275 vdd.n1221 4.74817
R22038 vdd.n1425 vdd.n1423 4.74817
R22039 vdd.n333 vdd.n332 4.7074
R22040 vdd.n231 vdd.n230 4.7074
R22041 vdd.n2173 vdd.n2172 4.7074
R22042 vdd.n2071 vdd.n2070 4.7074
R22043 vdd.n1482 vdd.t208 4.64847
R22044 vdd.n2454 vdd.t122 4.64847
R22045 vdd.n1018 vdd.t117 4.64847
R22046 vdd.n2975 vdd.t109 4.64847
R22047 vdd.n870 vdd.t0 4.64847
R22048 vdd.n3381 vdd.t191 4.64847
R22049 vdd.n2221 vdd.t256 4.42174
R22050 vdd.t202 vdd.n655 4.42174
R22051 vdd.n312 vdd.n300 4.26717
R22052 vdd.n253 vdd.n241 4.26717
R22053 vdd.n210 vdd.n198 4.26717
R22054 vdd.n151 vdd.n139 4.26717
R22055 vdd.n109 vdd.n97 4.26717
R22056 vdd.n50 vdd.n38 4.26717
R22057 vdd.n2093 vdd.n2081 4.26717
R22058 vdd.n2152 vdd.n2140 4.26717
R22059 vdd.n1991 vdd.n1979 4.26717
R22060 vdd.n2050 vdd.n2038 4.26717
R22061 vdd.n1890 vdd.n1878 4.26717
R22062 vdd.n1949 vdd.n1937 4.26717
R22063 vdd.n2237 vdd.t188 4.19501
R22064 vdd.n3340 vdd.t186 4.19501
R22065 vdd.n333 vdd.n231 4.10845
R22066 vdd.n2173 vdd.n2071 4.10845
R22067 vdd.n289 vdd.t224 4.06363
R22068 vdd.n289 vdd.t272 4.06363
R22069 vdd.n287 vdd.t275 4.06363
R22070 vdd.n287 vdd.t147 4.06363
R22071 vdd.n285 vdd.t178 4.06363
R22072 vdd.n285 vdd.t247 4.06363
R22073 vdd.n283 vdd.t279 4.06363
R22074 vdd.n283 vdd.t290 4.06363
R22075 vdd.n281 vdd.t295 4.06363
R22076 vdd.n281 vdd.t185 4.06363
R22077 vdd.n279 vdd.t218 4.06363
R22078 vdd.n279 vdd.t294 4.06363
R22079 vdd.n277 vdd.t296 4.06363
R22080 vdd.n277 vdd.t217 4.06363
R22081 vdd.n275 vdd.t223 4.06363
R22082 vdd.n275 vdd.t226 4.06363
R22083 vdd.n273 vdd.t274 4.06363
R22084 vdd.n273 vdd.t169 4.06363
R22085 vdd.n187 vdd.t201 4.06363
R22086 vdd.n187 vdd.t260 4.06363
R22087 vdd.n185 vdd.t261 4.06363
R22088 vdd.n185 vdd.t292 4.06363
R22089 vdd.n183 vdd.t159 4.06363
R22090 vdd.n183 vdd.t229 4.06363
R22091 vdd.n181 vdd.t266 4.06363
R22092 vdd.n181 vdd.t280 4.06363
R22093 vdd.n179 vdd.t284 4.06363
R22094 vdd.n179 vdd.t163 4.06363
R22095 vdd.n177 vdd.t193 4.06363
R22096 vdd.n177 vdd.t283 4.06363
R22097 vdd.n175 vdd.t285 4.06363
R22098 vdd.n175 vdd.t192 4.06363
R22099 vdd.n173 vdd.t203 4.06363
R22100 vdd.n173 vdd.t205 4.06363
R22101 vdd.n171 vdd.t263 4.06363
R22102 vdd.n171 vdd.t143 4.06363
R22103 vdd.n86 vdd.t235 4.06363
R22104 vdd.n86 vdd.t264 4.06363
R22105 vdd.n84 vdd.t214 4.06363
R22106 vdd.n84 vdd.t286 4.06363
R22107 vdd.n82 vdd.t177 4.06363
R22108 vdd.n82 vdd.t273 4.06363
R22109 vdd.n80 vdd.t171 4.06363
R22110 vdd.n80 vdd.t254 4.06363
R22111 vdd.n78 vdd.t195 4.06363
R22112 vdd.n78 vdd.t281 4.06363
R22113 vdd.n76 vdd.t165 4.06363
R22114 vdd.n76 vdd.t232 4.06363
R22115 vdd.n74 vdd.t153 4.06363
R22116 vdd.n74 vdd.t206 4.06363
R22117 vdd.n72 vdd.t291 4.06363
R22118 vdd.n72 vdd.t271 4.06363
R22119 vdd.n70 vdd.t277 4.06363
R22120 vdd.n70 vdd.t219 4.06363
R22121 vdd.n2113 vdd.t242 4.06363
R22122 vdd.n2113 vdd.t174 4.06363
R22123 vdd.n2115 vdd.t299 4.06363
R22124 vdd.n2115 vdd.t269 4.06363
R22125 vdd.n2117 vdd.t267 4.06363
R22126 vdd.n2117 vdd.t216 4.06363
R22127 vdd.n2119 vdd.t212 4.06363
R22128 vdd.n2119 vdd.t268 4.06363
R22129 vdd.n2121 vdd.t250 4.06363
R22130 vdd.n2121 vdd.t249 4.06363
R22131 vdd.n2123 vdd.t207 4.06363
R22132 vdd.n2123 vdd.t176 4.06363
R22133 vdd.n2125 vdd.t173 4.06363
R22134 vdd.n2125 vdd.t248 4.06363
R22135 vdd.n2127 vdd.t227 4.06363
R22136 vdd.n2127 vdd.t175 4.06363
R22137 vdd.n2129 vdd.t166 4.06363
R22138 vdd.n2129 vdd.t270 4.06363
R22139 vdd.n2011 vdd.t225 4.06363
R22140 vdd.n2011 vdd.t149 4.06363
R22141 vdd.n2013 vdd.t289 4.06363
R22142 vdd.n2013 vdd.t257 4.06363
R22143 vdd.n2015 vdd.t251 4.06363
R22144 vdd.n2015 vdd.t190 4.06363
R22145 vdd.n2017 vdd.t184 4.06363
R22146 vdd.n2017 vdd.t252 4.06363
R22147 vdd.n2019 vdd.t241 4.06363
R22148 vdd.n2019 vdd.t239 4.06363
R22149 vdd.n2021 vdd.t180 4.06363
R22150 vdd.n2021 vdd.t155 4.06363
R22151 vdd.n2023 vdd.t145 4.06363
R22152 vdd.n2023 vdd.t234 4.06363
R22153 vdd.n2025 vdd.t211 4.06363
R22154 vdd.n2025 vdd.t151 4.06363
R22155 vdd.n2027 vdd.t141 4.06363
R22156 vdd.n2027 vdd.t258 4.06363
R22157 vdd.n1910 vdd.t221 4.06363
R22158 vdd.n1910 vdd.t278 4.06363
R22159 vdd.n1912 vdd.t244 4.06363
R22160 vdd.n1912 vdd.t293 4.06363
R22161 vdd.n1914 vdd.t209 4.06363
R22162 vdd.n1914 vdd.t157 4.06363
R22163 vdd.n1916 vdd.t233 4.06363
R22164 vdd.n1916 vdd.t168 4.06363
R22165 vdd.n1918 vdd.t282 4.06363
R22166 vdd.n1918 vdd.t298 4.06363
R22167 vdd.n1920 vdd.t255 4.06363
R22168 vdd.n1920 vdd.t172 4.06363
R22169 vdd.n1922 vdd.t245 4.06363
R22170 vdd.n1922 vdd.t182 4.06363
R22171 vdd.n1924 vdd.t287 4.06363
R22172 vdd.n1924 vdd.t215 4.06363
R22173 vdd.n1926 vdd.t265 4.06363
R22174 vdd.n1926 vdd.t237 4.06363
R22175 vdd.n26 vdd.t13 3.9605
R22176 vdd.n26 vdd.t11 3.9605
R22177 vdd.n23 vdd.t6 3.9605
R22178 vdd.n23 vdd.t2 3.9605
R22179 vdd.n21 vdd.t8 3.9605
R22180 vdd.n21 vdd.t12 3.9605
R22181 vdd.n20 vdd.t7 3.9605
R22182 vdd.n20 vdd.t10 3.9605
R22183 vdd.n15 vdd.t3 3.9605
R22184 vdd.n15 vdd.t4 3.9605
R22185 vdd.n16 vdd.t16 3.9605
R22186 vdd.n16 vdd.t5 3.9605
R22187 vdd.n18 vdd.t15 3.9605
R22188 vdd.n18 vdd.t9 3.9605
R22189 vdd.n25 vdd.t14 3.9605
R22190 vdd.n25 vdd.t17 3.9605
R22191 vdd.n2511 vdd.t132 3.85492
R22192 vdd.n1338 vdd.t132 3.85492
R22193 vdd.n2951 vdd.t115 3.85492
R22194 vdd.t115 vdd.n917 3.85492
R22195 vdd.n7 vdd.t24 3.61217
R22196 vdd.n7 vdd.t126 3.61217
R22197 vdd.n8 vdd.t139 3.61217
R22198 vdd.n8 vdd.t111 3.61217
R22199 vdd.n10 vdd.t107 3.61217
R22200 vdd.n10 vdd.t116 3.61217
R22201 vdd.n12 vdd.t131 3.61217
R22202 vdd.n12 vdd.t103 3.61217
R22203 vdd.n5 vdd.t121 3.61217
R22204 vdd.n5 vdd.t137 3.61217
R22205 vdd.n3 vdd.t133 3.61217
R22206 vdd.n3 vdd.t119 3.61217
R22207 vdd.n1 vdd.t129 3.61217
R22208 vdd.n1 vdd.t105 3.61217
R22209 vdd.n0 vdd.t113 3.61217
R22210 vdd.n0 vdd.t135 3.61217
R22211 vdd.n316 vdd.n315 3.49141
R22212 vdd.n257 vdd.n256 3.49141
R22213 vdd.n214 vdd.n213 3.49141
R22214 vdd.n155 vdd.n154 3.49141
R22215 vdd.n113 vdd.n112 3.49141
R22216 vdd.n54 vdd.n53 3.49141
R22217 vdd.n2097 vdd.n2096 3.49141
R22218 vdd.n2156 vdd.n2155 3.49141
R22219 vdd.n1995 vdd.n1994 3.49141
R22220 vdd.n2054 vdd.n2053 3.49141
R22221 vdd.n1894 vdd.n1893 3.49141
R22222 vdd.n1953 vdd.n1952 3.49141
R22223 vdd.n2665 vdd.t120 3.40145
R22224 vdd.n2938 vdd.t102 3.40145
R22225 vdd.n2238 vdd.t148 3.28809
R22226 vdd.n3339 vdd.t262 3.28809
R22227 vdd.n3003 vdd.n3002 3.12245
R22228 vdd.n2459 vdd.n2458 3.12245
R22229 vdd.t243 vdd.n1466 3.06136
R22230 vdd.n1055 vdd.t122 3.06136
R22231 vdd.n2491 vdd.t117 3.06136
R22232 vdd.n2847 vdd.t109 3.06136
R22233 vdd.n3012 vdd.t0 3.06136
R22234 vdd.n3364 vdd.t204 3.06136
R22235 vdd.n2196 vdd.t167 2.83463
R22236 vdd.n644 vdd.t164 2.83463
R22237 vdd.n1359 vdd.t112 2.72126
R22238 vdd.n2987 vdd.t125 2.72126
R22239 vdd.n319 vdd.n298 2.71565
R22240 vdd.n260 vdd.n239 2.71565
R22241 vdd.n217 vdd.n196 2.71565
R22242 vdd.n158 vdd.n137 2.71565
R22243 vdd.n116 vdd.n95 2.71565
R22244 vdd.n57 vdd.n36 2.71565
R22245 vdd.n2100 vdd.n2079 2.71565
R22246 vdd.n2159 vdd.n2138 2.71565
R22247 vdd.n1998 vdd.n1977 2.71565
R22248 vdd.n2057 vdd.n2036 2.71565
R22249 vdd.n1897 vdd.n1876 2.71565
R22250 vdd.n1956 vdd.n1935 2.71565
R22251 vdd.t240 vdd.n1494 2.6079
R22252 vdd.n3487 vdd.t162 2.6079
R22253 vdd.t104 vdd.n999 2.49453
R22254 vdd.n2963 vdd.t138 2.49453
R22255 vdd.n306 vdd.n305 2.4129
R22256 vdd.n247 vdd.n246 2.4129
R22257 vdd.n204 vdd.n203 2.4129
R22258 vdd.n145 vdd.n144 2.4129
R22259 vdd.n103 vdd.n102 2.4129
R22260 vdd.n44 vdd.n43 2.4129
R22261 vdd.n2087 vdd.n2086 2.4129
R22262 vdd.n2146 vdd.n2145 2.4129
R22263 vdd.n1985 vdd.n1984 2.4129
R22264 vdd.n2044 vdd.n2043 2.4129
R22265 vdd.n1884 vdd.n1883 2.4129
R22266 vdd.n1943 vdd.n1942 2.4129
R22267 vdd.n1848 vdd.t181 2.38117
R22268 vdd.n2256 vdd.t39 2.38117
R22269 vdd.n1079 vdd.t31 2.38117
R22270 vdd.n2518 vdd.t73 2.38117
R22271 vdd.n2862 vdd.t77 2.38117
R22272 vdd.n3081 vdd.t27 2.38117
R22273 vdd.n3323 vdd.t35 2.38117
R22274 vdd.n3478 vdd.t158 2.38117
R22275 vdd.n2381 vdd.n1122 2.27742
R22276 vdd.n2381 vdd.n1121 2.27742
R22277 vdd.n3308 vdd.n3307 2.27742
R22278 vdd.n3309 vdd.n3308 2.27742
R22279 vdd.n3186 vdd.n3185 2.27742
R22280 vdd.n3185 vdd.n784 2.27742
R22281 vdd.n2275 vdd.n2274 2.27742
R22282 vdd.n2274 vdd.n1423 2.27742
R22283 vdd.t210 vdd.n1523 2.15444
R22284 vdd.n2467 vdd.t124 2.15444
R22285 vdd.n1359 vdd.t19 2.15444
R22286 vdd.n2987 vdd.t25 2.15444
R22287 vdd.t21 vdd.n875 2.15444
R22288 vdd.n3469 vdd.t146 2.15444
R22289 vdd.n320 vdd.n296 1.93989
R22290 vdd.n261 vdd.n237 1.93989
R22291 vdd.n218 vdd.n194 1.93989
R22292 vdd.n159 vdd.n135 1.93989
R22293 vdd.n117 vdd.n93 1.93989
R22294 vdd.n58 vdd.n34 1.93989
R22295 vdd.n2101 vdd.n2077 1.93989
R22296 vdd.n2160 vdd.n2136 1.93989
R22297 vdd.n1999 vdd.n1975 1.93989
R22298 vdd.n2058 vdd.n2034 1.93989
R22299 vdd.n1898 vdd.n1874 1.93989
R22300 vdd.n1957 vdd.n1933 1.93989
R22301 vdd.n1806 vdd.t196 1.92771
R22302 vdd.t160 vdd.n375 1.92771
R22303 vdd.n2491 vdd.t128 1.81434
R22304 vdd.n2847 vdd.t110 1.81434
R22305 vdd.n1814 vdd.t236 1.70098
R22306 vdd.n3463 vdd.t200 1.70098
R22307 vdd.n2485 vdd.t134 1.58761
R22308 vdd.n901 vdd.t23 1.58761
R22309 vdd.n1839 vdd.t144 1.47425
R22310 vdd.n361 vdd.t228 1.47425
R22311 vdd.n1505 vdd.t154 1.24752
R22312 vdd.n2461 vdd.t22 1.24752
R22313 vdd.n1024 vdd.t108 1.24752
R22314 vdd.n2981 vdd.t1 1.24752
R22315 vdd.n878 vdd.t123 1.24752
R22316 vdd.t170 vdd.n3485 1.24752
R22317 vdd.n331 vdd.n291 1.16414
R22318 vdd.n324 vdd.n323 1.16414
R22319 vdd.n272 vdd.n232 1.16414
R22320 vdd.n265 vdd.n264 1.16414
R22321 vdd.n229 vdd.n189 1.16414
R22322 vdd.n222 vdd.n221 1.16414
R22323 vdd.n170 vdd.n130 1.16414
R22324 vdd.n163 vdd.n162 1.16414
R22325 vdd.n128 vdd.n88 1.16414
R22326 vdd.n121 vdd.n120 1.16414
R22327 vdd.n69 vdd.n29 1.16414
R22328 vdd.n62 vdd.n61 1.16414
R22329 vdd.n2112 vdd.n2072 1.16414
R22330 vdd.n2105 vdd.n2104 1.16414
R22331 vdd.n2171 vdd.n2131 1.16414
R22332 vdd.n2164 vdd.n2163 1.16414
R22333 vdd.n2010 vdd.n1970 1.16414
R22334 vdd.n2003 vdd.n2002 1.16414
R22335 vdd.n2069 vdd.n2029 1.16414
R22336 vdd.n2062 vdd.n2061 1.16414
R22337 vdd.n1909 vdd.n1869 1.16414
R22338 vdd.n1902 vdd.n1901 1.16414
R22339 vdd.n1968 vdd.n1928 1.16414
R22340 vdd.n1961 vdd.n1960 1.16414
R22341 vdd.n2188 vdd.t183 1.02079
R22342 vdd.t84 vdd.t22 1.02079
R22343 vdd.t123 vdd.t53 1.02079
R22344 vdd.t231 vdd.n633 1.02079
R22345 vdd.n2174 vdd.n28 1.00834
R22346 vdd vdd.n3492 1.0005
R22347 vdd.n1685 vdd.n1681 0.970197
R22348 vdd.n2272 vdd.n2271 0.970197
R22349 vdd.n618 vdd.n428 0.970197
R22350 vdd.n3187 vdd.n690 0.970197
R22351 vdd.n2204 vdd.t156 0.794056
R22352 vdd.n3373 vdd.t152 0.794056
R22353 vdd.n2229 vdd.t220 0.567326
R22354 vdd.t142 vdd.n662 0.567326
R22355 vdd.n2262 vdd.n1123 0.530988
R22356 vdd.n726 vdd.n682 0.530988
R22357 vdd.n464 vdd.n391 0.530988
R22358 vdd.n3442 vdd.n3441 0.530988
R22359 vdd.n3319 vdd.n3318 0.530988
R22360 vdd.n2251 vdd.n1424 0.530988
R22361 vdd.n1683 vdd.n1548 0.530988
R22362 vdd.n1785 vdd.n1784 0.530988
R22363 vdd.n4 vdd.n2 0.459552
R22364 vdd.n11 vdd.n9 0.459552
R22365 vdd.t118 vdd.n976 0.453961
R22366 vdd.n2945 vdd.t106 0.453961
R22367 vdd.n329 vdd.n328 0.388379
R22368 vdd.n295 vdd.n293 0.388379
R22369 vdd.n270 vdd.n269 0.388379
R22370 vdd.n236 vdd.n234 0.388379
R22371 vdd.n227 vdd.n226 0.388379
R22372 vdd.n193 vdd.n191 0.388379
R22373 vdd.n168 vdd.n167 0.388379
R22374 vdd.n134 vdd.n132 0.388379
R22375 vdd.n126 vdd.n125 0.388379
R22376 vdd.n92 vdd.n90 0.388379
R22377 vdd.n67 vdd.n66 0.388379
R22378 vdd.n33 vdd.n31 0.388379
R22379 vdd.n2110 vdd.n2109 0.388379
R22380 vdd.n2076 vdd.n2074 0.388379
R22381 vdd.n2169 vdd.n2168 0.388379
R22382 vdd.n2135 vdd.n2133 0.388379
R22383 vdd.n2008 vdd.n2007 0.388379
R22384 vdd.n1974 vdd.n1972 0.388379
R22385 vdd.n2067 vdd.n2066 0.388379
R22386 vdd.n2033 vdd.n2031 0.388379
R22387 vdd.n1907 vdd.n1906 0.388379
R22388 vdd.n1873 vdd.n1871 0.388379
R22389 vdd.n1966 vdd.n1965 0.388379
R22390 vdd.n1932 vdd.n1930 0.388379
R22391 vdd.n19 vdd.n17 0.387128
R22392 vdd.n24 vdd.n22 0.387128
R22393 vdd.n6 vdd.n4 0.358259
R22394 vdd.n13 vdd.n11 0.358259
R22395 vdd.n276 vdd.n274 0.358259
R22396 vdd.n278 vdd.n276 0.358259
R22397 vdd.n280 vdd.n278 0.358259
R22398 vdd.n282 vdd.n280 0.358259
R22399 vdd.n284 vdd.n282 0.358259
R22400 vdd.n286 vdd.n284 0.358259
R22401 vdd.n288 vdd.n286 0.358259
R22402 vdd.n290 vdd.n288 0.358259
R22403 vdd.n332 vdd.n290 0.358259
R22404 vdd.n174 vdd.n172 0.358259
R22405 vdd.n176 vdd.n174 0.358259
R22406 vdd.n178 vdd.n176 0.358259
R22407 vdd.n180 vdd.n178 0.358259
R22408 vdd.n182 vdd.n180 0.358259
R22409 vdd.n184 vdd.n182 0.358259
R22410 vdd.n186 vdd.n184 0.358259
R22411 vdd.n188 vdd.n186 0.358259
R22412 vdd.n230 vdd.n188 0.358259
R22413 vdd.n73 vdd.n71 0.358259
R22414 vdd.n75 vdd.n73 0.358259
R22415 vdd.n77 vdd.n75 0.358259
R22416 vdd.n79 vdd.n77 0.358259
R22417 vdd.n81 vdd.n79 0.358259
R22418 vdd.n83 vdd.n81 0.358259
R22419 vdd.n85 vdd.n83 0.358259
R22420 vdd.n87 vdd.n85 0.358259
R22421 vdd.n129 vdd.n87 0.358259
R22422 vdd.n2172 vdd.n2130 0.358259
R22423 vdd.n2130 vdd.n2128 0.358259
R22424 vdd.n2128 vdd.n2126 0.358259
R22425 vdd.n2126 vdd.n2124 0.358259
R22426 vdd.n2124 vdd.n2122 0.358259
R22427 vdd.n2122 vdd.n2120 0.358259
R22428 vdd.n2120 vdd.n2118 0.358259
R22429 vdd.n2118 vdd.n2116 0.358259
R22430 vdd.n2116 vdd.n2114 0.358259
R22431 vdd.n2070 vdd.n2028 0.358259
R22432 vdd.n2028 vdd.n2026 0.358259
R22433 vdd.n2026 vdd.n2024 0.358259
R22434 vdd.n2024 vdd.n2022 0.358259
R22435 vdd.n2022 vdd.n2020 0.358259
R22436 vdd.n2020 vdd.n2018 0.358259
R22437 vdd.n2018 vdd.n2016 0.358259
R22438 vdd.n2016 vdd.n2014 0.358259
R22439 vdd.n2014 vdd.n2012 0.358259
R22440 vdd.n1969 vdd.n1927 0.358259
R22441 vdd.n1927 vdd.n1925 0.358259
R22442 vdd.n1925 vdd.n1923 0.358259
R22443 vdd.n1923 vdd.n1921 0.358259
R22444 vdd.n1921 vdd.n1919 0.358259
R22445 vdd.n1919 vdd.n1917 0.358259
R22446 vdd.n1917 vdd.n1915 0.358259
R22447 vdd.n1915 vdd.n1913 0.358259
R22448 vdd.n1913 vdd.n1911 0.358259
R22449 vdd.t18 vdd.n1052 0.340595
R22450 vdd.n2497 vdd.t20 0.340595
R22451 vdd.t127 vdd.n905 0.340595
R22452 vdd.n3018 vdd.t114 0.340595
R22453 vdd.n14 vdd.n6 0.334552
R22454 vdd.n14 vdd.n13 0.334552
R22455 vdd.n27 vdd.n19 0.21707
R22456 vdd.n27 vdd.n24 0.21707
R22457 vdd.n330 vdd.n292 0.155672
R22458 vdd.n322 vdd.n292 0.155672
R22459 vdd.n322 vdd.n321 0.155672
R22460 vdd.n321 vdd.n297 0.155672
R22461 vdd.n314 vdd.n297 0.155672
R22462 vdd.n314 vdd.n313 0.155672
R22463 vdd.n313 vdd.n301 0.155672
R22464 vdd.n306 vdd.n301 0.155672
R22465 vdd.n271 vdd.n233 0.155672
R22466 vdd.n263 vdd.n233 0.155672
R22467 vdd.n263 vdd.n262 0.155672
R22468 vdd.n262 vdd.n238 0.155672
R22469 vdd.n255 vdd.n238 0.155672
R22470 vdd.n255 vdd.n254 0.155672
R22471 vdd.n254 vdd.n242 0.155672
R22472 vdd.n247 vdd.n242 0.155672
R22473 vdd.n228 vdd.n190 0.155672
R22474 vdd.n220 vdd.n190 0.155672
R22475 vdd.n220 vdd.n219 0.155672
R22476 vdd.n219 vdd.n195 0.155672
R22477 vdd.n212 vdd.n195 0.155672
R22478 vdd.n212 vdd.n211 0.155672
R22479 vdd.n211 vdd.n199 0.155672
R22480 vdd.n204 vdd.n199 0.155672
R22481 vdd.n169 vdd.n131 0.155672
R22482 vdd.n161 vdd.n131 0.155672
R22483 vdd.n161 vdd.n160 0.155672
R22484 vdd.n160 vdd.n136 0.155672
R22485 vdd.n153 vdd.n136 0.155672
R22486 vdd.n153 vdd.n152 0.155672
R22487 vdd.n152 vdd.n140 0.155672
R22488 vdd.n145 vdd.n140 0.155672
R22489 vdd.n127 vdd.n89 0.155672
R22490 vdd.n119 vdd.n89 0.155672
R22491 vdd.n119 vdd.n118 0.155672
R22492 vdd.n118 vdd.n94 0.155672
R22493 vdd.n111 vdd.n94 0.155672
R22494 vdd.n111 vdd.n110 0.155672
R22495 vdd.n110 vdd.n98 0.155672
R22496 vdd.n103 vdd.n98 0.155672
R22497 vdd.n68 vdd.n30 0.155672
R22498 vdd.n60 vdd.n30 0.155672
R22499 vdd.n60 vdd.n59 0.155672
R22500 vdd.n59 vdd.n35 0.155672
R22501 vdd.n52 vdd.n35 0.155672
R22502 vdd.n52 vdd.n51 0.155672
R22503 vdd.n51 vdd.n39 0.155672
R22504 vdd.n44 vdd.n39 0.155672
R22505 vdd.n2111 vdd.n2073 0.155672
R22506 vdd.n2103 vdd.n2073 0.155672
R22507 vdd.n2103 vdd.n2102 0.155672
R22508 vdd.n2102 vdd.n2078 0.155672
R22509 vdd.n2095 vdd.n2078 0.155672
R22510 vdd.n2095 vdd.n2094 0.155672
R22511 vdd.n2094 vdd.n2082 0.155672
R22512 vdd.n2087 vdd.n2082 0.155672
R22513 vdd.n2170 vdd.n2132 0.155672
R22514 vdd.n2162 vdd.n2132 0.155672
R22515 vdd.n2162 vdd.n2161 0.155672
R22516 vdd.n2161 vdd.n2137 0.155672
R22517 vdd.n2154 vdd.n2137 0.155672
R22518 vdd.n2154 vdd.n2153 0.155672
R22519 vdd.n2153 vdd.n2141 0.155672
R22520 vdd.n2146 vdd.n2141 0.155672
R22521 vdd.n2009 vdd.n1971 0.155672
R22522 vdd.n2001 vdd.n1971 0.155672
R22523 vdd.n2001 vdd.n2000 0.155672
R22524 vdd.n2000 vdd.n1976 0.155672
R22525 vdd.n1993 vdd.n1976 0.155672
R22526 vdd.n1993 vdd.n1992 0.155672
R22527 vdd.n1992 vdd.n1980 0.155672
R22528 vdd.n1985 vdd.n1980 0.155672
R22529 vdd.n2068 vdd.n2030 0.155672
R22530 vdd.n2060 vdd.n2030 0.155672
R22531 vdd.n2060 vdd.n2059 0.155672
R22532 vdd.n2059 vdd.n2035 0.155672
R22533 vdd.n2052 vdd.n2035 0.155672
R22534 vdd.n2052 vdd.n2051 0.155672
R22535 vdd.n2051 vdd.n2039 0.155672
R22536 vdd.n2044 vdd.n2039 0.155672
R22537 vdd.n1908 vdd.n1870 0.155672
R22538 vdd.n1900 vdd.n1870 0.155672
R22539 vdd.n1900 vdd.n1899 0.155672
R22540 vdd.n1899 vdd.n1875 0.155672
R22541 vdd.n1892 vdd.n1875 0.155672
R22542 vdd.n1892 vdd.n1891 0.155672
R22543 vdd.n1891 vdd.n1879 0.155672
R22544 vdd.n1884 vdd.n1879 0.155672
R22545 vdd.n1967 vdd.n1929 0.155672
R22546 vdd.n1959 vdd.n1929 0.155672
R22547 vdd.n1959 vdd.n1958 0.155672
R22548 vdd.n1958 vdd.n1934 0.155672
R22549 vdd.n1951 vdd.n1934 0.155672
R22550 vdd.n1951 vdd.n1950 0.155672
R22551 vdd.n1950 vdd.n1938 0.155672
R22552 vdd.n1943 vdd.n1938 0.155672
R22553 vdd.n1128 vdd.n1120 0.152939
R22554 vdd.n1132 vdd.n1128 0.152939
R22555 vdd.n1133 vdd.n1132 0.152939
R22556 vdd.n1134 vdd.n1133 0.152939
R22557 vdd.n1135 vdd.n1134 0.152939
R22558 vdd.n1139 vdd.n1135 0.152939
R22559 vdd.n1140 vdd.n1139 0.152939
R22560 vdd.n1141 vdd.n1140 0.152939
R22561 vdd.n1142 vdd.n1141 0.152939
R22562 vdd.n1146 vdd.n1142 0.152939
R22563 vdd.n1147 vdd.n1146 0.152939
R22564 vdd.n1148 vdd.n1147 0.152939
R22565 vdd.n2345 vdd.n1148 0.152939
R22566 vdd.n2345 vdd.n2344 0.152939
R22567 vdd.n2344 vdd.n2343 0.152939
R22568 vdd.n2343 vdd.n1154 0.152939
R22569 vdd.n1159 vdd.n1154 0.152939
R22570 vdd.n1160 vdd.n1159 0.152939
R22571 vdd.n1161 vdd.n1160 0.152939
R22572 vdd.n1165 vdd.n1161 0.152939
R22573 vdd.n1166 vdd.n1165 0.152939
R22574 vdd.n1167 vdd.n1166 0.152939
R22575 vdd.n1168 vdd.n1167 0.152939
R22576 vdd.n1172 vdd.n1168 0.152939
R22577 vdd.n1173 vdd.n1172 0.152939
R22578 vdd.n1174 vdd.n1173 0.152939
R22579 vdd.n1175 vdd.n1174 0.152939
R22580 vdd.n1179 vdd.n1175 0.152939
R22581 vdd.n1180 vdd.n1179 0.152939
R22582 vdd.n1181 vdd.n1180 0.152939
R22583 vdd.n1182 vdd.n1181 0.152939
R22584 vdd.n1186 vdd.n1182 0.152939
R22585 vdd.n1187 vdd.n1186 0.152939
R22586 vdd.n1188 vdd.n1187 0.152939
R22587 vdd.n2306 vdd.n1188 0.152939
R22588 vdd.n2306 vdd.n2305 0.152939
R22589 vdd.n2305 vdd.n2304 0.152939
R22590 vdd.n2304 vdd.n1194 0.152939
R22591 vdd.n1199 vdd.n1194 0.152939
R22592 vdd.n1200 vdd.n1199 0.152939
R22593 vdd.n1201 vdd.n1200 0.152939
R22594 vdd.n1205 vdd.n1201 0.152939
R22595 vdd.n1206 vdd.n1205 0.152939
R22596 vdd.n1207 vdd.n1206 0.152939
R22597 vdd.n1208 vdd.n1207 0.152939
R22598 vdd.n1212 vdd.n1208 0.152939
R22599 vdd.n1213 vdd.n1212 0.152939
R22600 vdd.n1214 vdd.n1213 0.152939
R22601 vdd.n1215 vdd.n1214 0.152939
R22602 vdd.n1219 vdd.n1215 0.152939
R22603 vdd.n1220 vdd.n1219 0.152939
R22604 vdd.n2380 vdd.n1123 0.152939
R22605 vdd.n2176 vdd.n1485 0.152939
R22606 vdd.n2191 vdd.n1485 0.152939
R22607 vdd.n2192 vdd.n2191 0.152939
R22608 vdd.n2193 vdd.n2192 0.152939
R22609 vdd.n2193 vdd.n1474 0.152939
R22610 vdd.n2208 vdd.n1474 0.152939
R22611 vdd.n2209 vdd.n2208 0.152939
R22612 vdd.n2210 vdd.n2209 0.152939
R22613 vdd.n2210 vdd.n1463 0.152939
R22614 vdd.n2224 vdd.n1463 0.152939
R22615 vdd.n2225 vdd.n2224 0.152939
R22616 vdd.n2226 vdd.n2225 0.152939
R22617 vdd.n2226 vdd.n1451 0.152939
R22618 vdd.n2241 vdd.n1451 0.152939
R22619 vdd.n2242 vdd.n2241 0.152939
R22620 vdd.n2243 vdd.n2242 0.152939
R22621 vdd.n2243 vdd.n1439 0.152939
R22622 vdd.n2260 vdd.n1439 0.152939
R22623 vdd.n2261 vdd.n2260 0.152939
R22624 vdd.n2262 vdd.n2261 0.152939
R22625 vdd.n735 vdd.n730 0.152939
R22626 vdd.n736 vdd.n735 0.152939
R22627 vdd.n737 vdd.n736 0.152939
R22628 vdd.n738 vdd.n737 0.152939
R22629 vdd.n739 vdd.n738 0.152939
R22630 vdd.n740 vdd.n739 0.152939
R22631 vdd.n741 vdd.n740 0.152939
R22632 vdd.n742 vdd.n741 0.152939
R22633 vdd.n743 vdd.n742 0.152939
R22634 vdd.n744 vdd.n743 0.152939
R22635 vdd.n745 vdd.n744 0.152939
R22636 vdd.n746 vdd.n745 0.152939
R22637 vdd.n3275 vdd.n746 0.152939
R22638 vdd.n3275 vdd.n3274 0.152939
R22639 vdd.n3274 vdd.n3273 0.152939
R22640 vdd.n3273 vdd.n748 0.152939
R22641 vdd.n749 vdd.n748 0.152939
R22642 vdd.n750 vdd.n749 0.152939
R22643 vdd.n751 vdd.n750 0.152939
R22644 vdd.n752 vdd.n751 0.152939
R22645 vdd.n753 vdd.n752 0.152939
R22646 vdd.n754 vdd.n753 0.152939
R22647 vdd.n755 vdd.n754 0.152939
R22648 vdd.n756 vdd.n755 0.152939
R22649 vdd.n757 vdd.n756 0.152939
R22650 vdd.n758 vdd.n757 0.152939
R22651 vdd.n759 vdd.n758 0.152939
R22652 vdd.n760 vdd.n759 0.152939
R22653 vdd.n761 vdd.n760 0.152939
R22654 vdd.n762 vdd.n761 0.152939
R22655 vdd.n763 vdd.n762 0.152939
R22656 vdd.n764 vdd.n763 0.152939
R22657 vdd.n765 vdd.n764 0.152939
R22658 vdd.n766 vdd.n765 0.152939
R22659 vdd.n3229 vdd.n766 0.152939
R22660 vdd.n3229 vdd.n3228 0.152939
R22661 vdd.n3228 vdd.n3227 0.152939
R22662 vdd.n3227 vdd.n770 0.152939
R22663 vdd.n771 vdd.n770 0.152939
R22664 vdd.n772 vdd.n771 0.152939
R22665 vdd.n773 vdd.n772 0.152939
R22666 vdd.n774 vdd.n773 0.152939
R22667 vdd.n775 vdd.n774 0.152939
R22668 vdd.n776 vdd.n775 0.152939
R22669 vdd.n777 vdd.n776 0.152939
R22670 vdd.n778 vdd.n777 0.152939
R22671 vdd.n779 vdd.n778 0.152939
R22672 vdd.n780 vdd.n779 0.152939
R22673 vdd.n781 vdd.n780 0.152939
R22674 vdd.n782 vdd.n781 0.152939
R22675 vdd.n783 vdd.n782 0.152939
R22676 vdd.n727 vdd.n726 0.152939
R22677 vdd.n3326 vdd.n682 0.152939
R22678 vdd.n3327 vdd.n3326 0.152939
R22679 vdd.n3328 vdd.n3327 0.152939
R22680 vdd.n3328 vdd.n670 0.152939
R22681 vdd.n3343 vdd.n670 0.152939
R22682 vdd.n3344 vdd.n3343 0.152939
R22683 vdd.n3345 vdd.n3344 0.152939
R22684 vdd.n3345 vdd.n659 0.152939
R22685 vdd.n3359 vdd.n659 0.152939
R22686 vdd.n3360 vdd.n3359 0.152939
R22687 vdd.n3361 vdd.n3360 0.152939
R22688 vdd.n3361 vdd.n647 0.152939
R22689 vdd.n3376 vdd.n647 0.152939
R22690 vdd.n3377 vdd.n3376 0.152939
R22691 vdd.n3378 vdd.n3377 0.152939
R22692 vdd.n3378 vdd.n636 0.152939
R22693 vdd.n3395 vdd.n636 0.152939
R22694 vdd.n3396 vdd.n3395 0.152939
R22695 vdd.n3397 vdd.n3396 0.152939
R22696 vdd.n3397 vdd.n334 0.152939
R22697 vdd.n3490 vdd.n335 0.152939
R22698 vdd.n346 vdd.n335 0.152939
R22699 vdd.n347 vdd.n346 0.152939
R22700 vdd.n348 vdd.n347 0.152939
R22701 vdd.n355 vdd.n348 0.152939
R22702 vdd.n356 vdd.n355 0.152939
R22703 vdd.n357 vdd.n356 0.152939
R22704 vdd.n358 vdd.n357 0.152939
R22705 vdd.n366 vdd.n358 0.152939
R22706 vdd.n367 vdd.n366 0.152939
R22707 vdd.n368 vdd.n367 0.152939
R22708 vdd.n369 vdd.n368 0.152939
R22709 vdd.n377 vdd.n369 0.152939
R22710 vdd.n378 vdd.n377 0.152939
R22711 vdd.n379 vdd.n378 0.152939
R22712 vdd.n380 vdd.n379 0.152939
R22713 vdd.n388 vdd.n380 0.152939
R22714 vdd.n389 vdd.n388 0.152939
R22715 vdd.n390 vdd.n389 0.152939
R22716 vdd.n391 vdd.n390 0.152939
R22717 vdd.n464 vdd.n463 0.152939
R22718 vdd.n470 vdd.n463 0.152939
R22719 vdd.n471 vdd.n470 0.152939
R22720 vdd.n472 vdd.n471 0.152939
R22721 vdd.n472 vdd.n461 0.152939
R22722 vdd.n480 vdd.n461 0.152939
R22723 vdd.n481 vdd.n480 0.152939
R22724 vdd.n482 vdd.n481 0.152939
R22725 vdd.n482 vdd.n459 0.152939
R22726 vdd.n490 vdd.n459 0.152939
R22727 vdd.n491 vdd.n490 0.152939
R22728 vdd.n492 vdd.n491 0.152939
R22729 vdd.n492 vdd.n457 0.152939
R22730 vdd.n500 vdd.n457 0.152939
R22731 vdd.n501 vdd.n500 0.152939
R22732 vdd.n502 vdd.n501 0.152939
R22733 vdd.n502 vdd.n455 0.152939
R22734 vdd.n510 vdd.n455 0.152939
R22735 vdd.n511 vdd.n510 0.152939
R22736 vdd.n512 vdd.n511 0.152939
R22737 vdd.n512 vdd.n451 0.152939
R22738 vdd.n520 vdd.n451 0.152939
R22739 vdd.n521 vdd.n520 0.152939
R22740 vdd.n522 vdd.n521 0.152939
R22741 vdd.n522 vdd.n449 0.152939
R22742 vdd.n530 vdd.n449 0.152939
R22743 vdd.n531 vdd.n530 0.152939
R22744 vdd.n532 vdd.n531 0.152939
R22745 vdd.n532 vdd.n447 0.152939
R22746 vdd.n540 vdd.n447 0.152939
R22747 vdd.n541 vdd.n540 0.152939
R22748 vdd.n542 vdd.n541 0.152939
R22749 vdd.n542 vdd.n445 0.152939
R22750 vdd.n550 vdd.n445 0.152939
R22751 vdd.n551 vdd.n550 0.152939
R22752 vdd.n552 vdd.n551 0.152939
R22753 vdd.n552 vdd.n443 0.152939
R22754 vdd.n560 vdd.n443 0.152939
R22755 vdd.n561 vdd.n560 0.152939
R22756 vdd.n562 vdd.n561 0.152939
R22757 vdd.n562 vdd.n439 0.152939
R22758 vdd.n570 vdd.n439 0.152939
R22759 vdd.n571 vdd.n570 0.152939
R22760 vdd.n572 vdd.n571 0.152939
R22761 vdd.n572 vdd.n437 0.152939
R22762 vdd.n580 vdd.n437 0.152939
R22763 vdd.n581 vdd.n580 0.152939
R22764 vdd.n582 vdd.n581 0.152939
R22765 vdd.n582 vdd.n435 0.152939
R22766 vdd.n590 vdd.n435 0.152939
R22767 vdd.n591 vdd.n590 0.152939
R22768 vdd.n592 vdd.n591 0.152939
R22769 vdd.n592 vdd.n433 0.152939
R22770 vdd.n600 vdd.n433 0.152939
R22771 vdd.n601 vdd.n600 0.152939
R22772 vdd.n602 vdd.n601 0.152939
R22773 vdd.n602 vdd.n431 0.152939
R22774 vdd.n610 vdd.n431 0.152939
R22775 vdd.n611 vdd.n610 0.152939
R22776 vdd.n612 vdd.n611 0.152939
R22777 vdd.n612 vdd.n429 0.152939
R22778 vdd.n619 vdd.n429 0.152939
R22779 vdd.n3442 vdd.n619 0.152939
R22780 vdd.n3320 vdd.n3319 0.152939
R22781 vdd.n3320 vdd.n675 0.152939
R22782 vdd.n3334 vdd.n675 0.152939
R22783 vdd.n3335 vdd.n3334 0.152939
R22784 vdd.n3336 vdd.n3335 0.152939
R22785 vdd.n3336 vdd.n665 0.152939
R22786 vdd.n3351 vdd.n665 0.152939
R22787 vdd.n3352 vdd.n3351 0.152939
R22788 vdd.n3353 vdd.n3352 0.152939
R22789 vdd.n3353 vdd.n652 0.152939
R22790 vdd.n3367 vdd.n652 0.152939
R22791 vdd.n3368 vdd.n3367 0.152939
R22792 vdd.n3369 vdd.n3368 0.152939
R22793 vdd.n3369 vdd.n641 0.152939
R22794 vdd.n3384 vdd.n641 0.152939
R22795 vdd.n3385 vdd.n3384 0.152939
R22796 vdd.n3386 vdd.n3385 0.152939
R22797 vdd.n3388 vdd.n3386 0.152939
R22798 vdd.n3388 vdd.n3387 0.152939
R22799 vdd.n3387 vdd.n630 0.152939
R22800 vdd.n3405 vdd.n630 0.152939
R22801 vdd.n3406 vdd.n3405 0.152939
R22802 vdd.n3407 vdd.n3406 0.152939
R22803 vdd.n3407 vdd.n628 0.152939
R22804 vdd.n3412 vdd.n628 0.152939
R22805 vdd.n3413 vdd.n3412 0.152939
R22806 vdd.n3414 vdd.n3413 0.152939
R22807 vdd.n3414 vdd.n626 0.152939
R22808 vdd.n3419 vdd.n626 0.152939
R22809 vdd.n3420 vdd.n3419 0.152939
R22810 vdd.n3421 vdd.n3420 0.152939
R22811 vdd.n3421 vdd.n624 0.152939
R22812 vdd.n3427 vdd.n624 0.152939
R22813 vdd.n3428 vdd.n3427 0.152939
R22814 vdd.n3429 vdd.n3428 0.152939
R22815 vdd.n3429 vdd.n622 0.152939
R22816 vdd.n3434 vdd.n622 0.152939
R22817 vdd.n3435 vdd.n3434 0.152939
R22818 vdd.n3436 vdd.n3435 0.152939
R22819 vdd.n3436 vdd.n620 0.152939
R22820 vdd.n3441 vdd.n620 0.152939
R22821 vdd.n3318 vdd.n687 0.152939
R22822 vdd.n2273 vdd.n1424 0.152939
R22823 vdd.n1792 vdd.n1548 0.152939
R22824 vdd.n1793 vdd.n1792 0.152939
R22825 vdd.n1794 vdd.n1793 0.152939
R22826 vdd.n1794 vdd.n1536 0.152939
R22827 vdd.n1809 vdd.n1536 0.152939
R22828 vdd.n1810 vdd.n1809 0.152939
R22829 vdd.n1811 vdd.n1810 0.152939
R22830 vdd.n1811 vdd.n1526 0.152939
R22831 vdd.n1826 vdd.n1526 0.152939
R22832 vdd.n1827 vdd.n1826 0.152939
R22833 vdd.n1828 vdd.n1827 0.152939
R22834 vdd.n1828 vdd.n1513 0.152939
R22835 vdd.n1842 vdd.n1513 0.152939
R22836 vdd.n1843 vdd.n1842 0.152939
R22837 vdd.n1844 vdd.n1843 0.152939
R22838 vdd.n1844 vdd.n1502 0.152939
R22839 vdd.n1859 vdd.n1502 0.152939
R22840 vdd.n1860 vdd.n1859 0.152939
R22841 vdd.n1861 vdd.n1860 0.152939
R22842 vdd.n1861 vdd.n1491 0.152939
R22843 vdd.n2182 vdd.n1491 0.152939
R22844 vdd.n2183 vdd.n2182 0.152939
R22845 vdd.n2184 vdd.n2183 0.152939
R22846 vdd.n2184 vdd.n1479 0.152939
R22847 vdd.n2199 vdd.n1479 0.152939
R22848 vdd.n2200 vdd.n2199 0.152939
R22849 vdd.n2201 vdd.n2200 0.152939
R22850 vdd.n2201 vdd.n1469 0.152939
R22851 vdd.n2216 vdd.n1469 0.152939
R22852 vdd.n2217 vdd.n2216 0.152939
R22853 vdd.n2218 vdd.n2217 0.152939
R22854 vdd.n2218 vdd.n1456 0.152939
R22855 vdd.n2232 vdd.n1456 0.152939
R22856 vdd.n2233 vdd.n2232 0.152939
R22857 vdd.n2234 vdd.n2233 0.152939
R22858 vdd.n2234 vdd.n1446 0.152939
R22859 vdd.n2249 vdd.n1446 0.152939
R22860 vdd.n2250 vdd.n2249 0.152939
R22861 vdd.n2253 vdd.n2250 0.152939
R22862 vdd.n2253 vdd.n2252 0.152939
R22863 vdd.n2252 vdd.n2251 0.152939
R22864 vdd.n1784 vdd.n1553 0.152939
R22865 vdd.n1777 vdd.n1553 0.152939
R22866 vdd.n1777 vdd.n1776 0.152939
R22867 vdd.n1776 vdd.n1775 0.152939
R22868 vdd.n1775 vdd.n1590 0.152939
R22869 vdd.n1771 vdd.n1590 0.152939
R22870 vdd.n1771 vdd.n1770 0.152939
R22871 vdd.n1770 vdd.n1769 0.152939
R22872 vdd.n1769 vdd.n1596 0.152939
R22873 vdd.n1765 vdd.n1596 0.152939
R22874 vdd.n1765 vdd.n1764 0.152939
R22875 vdd.n1764 vdd.n1763 0.152939
R22876 vdd.n1763 vdd.n1602 0.152939
R22877 vdd.n1759 vdd.n1602 0.152939
R22878 vdd.n1759 vdd.n1758 0.152939
R22879 vdd.n1758 vdd.n1757 0.152939
R22880 vdd.n1757 vdd.n1608 0.152939
R22881 vdd.n1753 vdd.n1608 0.152939
R22882 vdd.n1753 vdd.n1752 0.152939
R22883 vdd.n1752 vdd.n1751 0.152939
R22884 vdd.n1751 vdd.n1616 0.152939
R22885 vdd.n1747 vdd.n1616 0.152939
R22886 vdd.n1747 vdd.n1746 0.152939
R22887 vdd.n1746 vdd.n1745 0.152939
R22888 vdd.n1745 vdd.n1622 0.152939
R22889 vdd.n1741 vdd.n1622 0.152939
R22890 vdd.n1741 vdd.n1740 0.152939
R22891 vdd.n1740 vdd.n1739 0.152939
R22892 vdd.n1739 vdd.n1628 0.152939
R22893 vdd.n1735 vdd.n1628 0.152939
R22894 vdd.n1735 vdd.n1734 0.152939
R22895 vdd.n1734 vdd.n1733 0.152939
R22896 vdd.n1733 vdd.n1634 0.152939
R22897 vdd.n1729 vdd.n1634 0.152939
R22898 vdd.n1729 vdd.n1728 0.152939
R22899 vdd.n1728 vdd.n1727 0.152939
R22900 vdd.n1727 vdd.n1640 0.152939
R22901 vdd.n1723 vdd.n1640 0.152939
R22902 vdd.n1723 vdd.n1722 0.152939
R22903 vdd.n1722 vdd.n1721 0.152939
R22904 vdd.n1721 vdd.n1646 0.152939
R22905 vdd.n1714 vdd.n1646 0.152939
R22906 vdd.n1714 vdd.n1713 0.152939
R22907 vdd.n1713 vdd.n1712 0.152939
R22908 vdd.n1712 vdd.n1651 0.152939
R22909 vdd.n1708 vdd.n1651 0.152939
R22910 vdd.n1708 vdd.n1707 0.152939
R22911 vdd.n1707 vdd.n1706 0.152939
R22912 vdd.n1706 vdd.n1657 0.152939
R22913 vdd.n1702 vdd.n1657 0.152939
R22914 vdd.n1702 vdd.n1701 0.152939
R22915 vdd.n1701 vdd.n1700 0.152939
R22916 vdd.n1700 vdd.n1663 0.152939
R22917 vdd.n1696 vdd.n1663 0.152939
R22918 vdd.n1696 vdd.n1695 0.152939
R22919 vdd.n1695 vdd.n1694 0.152939
R22920 vdd.n1694 vdd.n1669 0.152939
R22921 vdd.n1690 vdd.n1669 0.152939
R22922 vdd.n1690 vdd.n1689 0.152939
R22923 vdd.n1689 vdd.n1688 0.152939
R22924 vdd.n1688 vdd.n1675 0.152939
R22925 vdd.n1684 vdd.n1675 0.152939
R22926 vdd.n1684 vdd.n1683 0.152939
R22927 vdd.n1786 vdd.n1785 0.152939
R22928 vdd.n1786 vdd.n1542 0.152939
R22929 vdd.n1801 vdd.n1542 0.152939
R22930 vdd.n1802 vdd.n1801 0.152939
R22931 vdd.n1803 vdd.n1802 0.152939
R22932 vdd.n1803 vdd.n1531 0.152939
R22933 vdd.n1818 vdd.n1531 0.152939
R22934 vdd.n1819 vdd.n1818 0.152939
R22935 vdd.n1820 vdd.n1819 0.152939
R22936 vdd.n1820 vdd.n1520 0.152939
R22937 vdd.n1834 vdd.n1520 0.152939
R22938 vdd.n1835 vdd.n1834 0.152939
R22939 vdd.n1836 vdd.n1835 0.152939
R22940 vdd.n1836 vdd.n1508 0.152939
R22941 vdd.n1851 vdd.n1508 0.152939
R22942 vdd.n1852 vdd.n1851 0.152939
R22943 vdd.n1853 vdd.n1852 0.152939
R22944 vdd.n1853 vdd.n1497 0.152939
R22945 vdd.n1867 vdd.n1497 0.152939
R22946 vdd.n1868 vdd.n1867 0.152939
R22947 vdd.n1789 vdd.t63 0.113865
R22948 vdd.t49 vdd.n386 0.113865
R22949 vdd.n2381 vdd.n2380 0.110256
R22950 vdd.n3308 vdd.n727 0.110256
R22951 vdd.n3185 vdd.n687 0.110256
R22952 vdd.n2274 vdd.n2273 0.110256
R22953 vdd.n2176 vdd.n2175 0.0695946
R22954 vdd.n3491 vdd.n334 0.0695946
R22955 vdd.n3491 vdd.n3490 0.0695946
R22956 vdd.n2175 vdd.n1868 0.0695946
R22957 vdd.n2381 vdd.n1120 0.0431829
R22958 vdd.n2274 vdd.n1220 0.0431829
R22959 vdd.n3308 vdd.n730 0.0431829
R22960 vdd.n3185 vdd.n783 0.0431829
R22961 vdd vdd.n28 0.00833333
R22962 a_n2318_13878.n59 a_n2318_13878.t82 533.335
R22963 a_n2318_13878.n75 a_n2318_13878.t63 512.366
R22964 a_n2318_13878.n70 a_n2318_13878.t67 512.366
R22965 a_n2318_13878.n74 a_n2318_13878.t57 512.366
R22966 a_n2318_13878.n73 a_n2318_13878.t72 512.366
R22967 a_n2318_13878.n71 a_n2318_13878.t79 512.366
R22968 a_n2318_13878.n72 a_n2318_13878.t80 512.366
R22969 a_n2318_13878.n53 a_n2318_13878.t35 533.335
R22970 a_n2318_13878.n89 a_n2318_13878.t43 512.366
R22971 a_n2318_13878.n68 a_n2318_13878.t21 512.366
R22972 a_n2318_13878.n88 a_n2318_13878.t33 512.366
R22973 a_n2318_13878.n87 a_n2318_13878.t25 512.366
R22974 a_n2318_13878.n69 a_n2318_13878.t45 512.366
R22975 a_n2318_13878.n86 a_n2318_13878.t27 512.366
R22976 a_n2318_13878.n37 a_n2318_13878.t23 533.335
R22977 a_n2318_13878.n112 a_n2318_13878.t31 512.366
R22978 a_n2318_13878.n113 a_n2318_13878.t19 512.366
R22979 a_n2318_13878.n114 a_n2318_13878.t29 512.366
R22980 a_n2318_13878.n115 a_n2318_13878.t17 512.366
R22981 a_n2318_13878.n66 a_n2318_13878.t37 512.366
R22982 a_n2318_13878.n116 a_n2318_13878.t41 512.366
R22983 a_n2318_13878.n30 a_n2318_13878.t78 533.335
R22984 a_n2318_13878.n107 a_n2318_13878.t56 512.366
R22985 a_n2318_13878.n108 a_n2318_13878.t75 512.366
R22986 a_n2318_13878.n109 a_n2318_13878.t76 512.366
R22987 a_n2318_13878.n110 a_n2318_13878.t53 512.366
R22988 a_n2318_13878.n67 a_n2318_13878.t62 512.366
R22989 a_n2318_13878.n111 a_n2318_13878.t70 512.366
R22990 a_n2318_13878.n99 a_n2318_13878.t69 512.366
R22991 a_n2318_13878.n98 a_n2318_13878.t60 512.366
R22992 a_n2318_13878.n97 a_n2318_13878.t52 512.366
R22993 a_n2318_13878.n101 a_n2318_13878.t77 512.366
R22994 a_n2318_13878.n100 a_n2318_13878.t66 512.366
R22995 a_n2318_13878.n96 a_n2318_13878.t65 512.366
R22996 a_n2318_13878.n103 a_n2318_13878.t73 512.366
R22997 a_n2318_13878.n102 a_n2318_13878.t58 512.366
R22998 a_n2318_13878.n95 a_n2318_13878.t59 512.366
R22999 a_n2318_13878.n105 a_n2318_13878.t61 512.366
R23000 a_n2318_13878.n104 a_n2318_13878.t71 512.366
R23001 a_n2318_13878.n94 a_n2318_13878.t83 512.366
R23002 a_n2318_13878.n64 a_n2318_13878.n1 70.1674
R23003 a_n2318_13878.n58 a_n2318_13878.n5 70.1674
R23004 a_n2318_13878.n16 a_n2318_13878.n43 70.1674
R23005 a_n2318_13878.n19 a_n2318_13878.n36 70.1674
R23006 a_n2318_13878.n111 a_n2318_13878.n36 20.9683
R23007 a_n2318_13878.n35 a_n2318_13878.n20 72.3034
R23008 a_n2318_13878.n35 a_n2318_13878.n67 16.6962
R23009 a_n2318_13878.n20 a_n2318_13878.n34 77.6622
R23010 a_n2318_13878.n110 a_n2318_13878.n34 5.97853
R23011 a_n2318_13878.n33 a_n2318_13878.n21 77.6622
R23012 a_n2318_13878.n21 a_n2318_13878.n32 72.3034
R23013 a_n2318_13878.n107 a_n2318_13878.n30 20.9683
R23014 a_n2318_13878.n31 a_n2318_13878.n30 70.1674
R23015 a_n2318_13878.n116 a_n2318_13878.n43 20.9683
R23016 a_n2318_13878.n42 a_n2318_13878.n17 72.3034
R23017 a_n2318_13878.n42 a_n2318_13878.n66 16.6962
R23018 a_n2318_13878.n17 a_n2318_13878.n41 77.6622
R23019 a_n2318_13878.n115 a_n2318_13878.n41 5.97853
R23020 a_n2318_13878.n40 a_n2318_13878.n18 77.6622
R23021 a_n2318_13878.n18 a_n2318_13878.n39 72.3034
R23022 a_n2318_13878.n112 a_n2318_13878.n37 20.9683
R23023 a_n2318_13878.n38 a_n2318_13878.n37 70.1674
R23024 a_n2318_13878.n8 a_n2318_13878.n52 70.1674
R23025 a_n2318_13878.n10 a_n2318_13878.n49 70.1674
R23026 a_n2318_13878.n12 a_n2318_13878.n47 70.1674
R23027 a_n2318_13878.n14 a_n2318_13878.n45 70.1674
R23028 a_n2318_13878.n45 a_n2318_13878.n94 20.9683
R23029 a_n2318_13878.n44 a_n2318_13878.n15 75.0448
R23030 a_n2318_13878.n104 a_n2318_13878.n44 11.2134
R23031 a_n2318_13878.n15 a_n2318_13878.n105 161.3
R23032 a_n2318_13878.n47 a_n2318_13878.n95 20.9683
R23033 a_n2318_13878.n46 a_n2318_13878.n13 75.0448
R23034 a_n2318_13878.n102 a_n2318_13878.n46 11.2134
R23035 a_n2318_13878.n13 a_n2318_13878.n103 161.3
R23036 a_n2318_13878.n49 a_n2318_13878.n96 20.9683
R23037 a_n2318_13878.n48 a_n2318_13878.n11 75.0448
R23038 a_n2318_13878.n100 a_n2318_13878.n48 11.2134
R23039 a_n2318_13878.n11 a_n2318_13878.n101 161.3
R23040 a_n2318_13878.n52 a_n2318_13878.n97 20.9683
R23041 a_n2318_13878.n50 a_n2318_13878.n9 75.0448
R23042 a_n2318_13878.n98 a_n2318_13878.n50 11.2134
R23043 a_n2318_13878.n9 a_n2318_13878.n99 161.3
R23044 a_n2318_13878.n86 a_n2318_13878.n58 20.9683
R23045 a_n2318_13878.n6 a_n2318_13878.n57 72.3034
R23046 a_n2318_13878.n57 a_n2318_13878.n69 16.6962
R23047 a_n2318_13878.n56 a_n2318_13878.n6 77.6622
R23048 a_n2318_13878.n87 a_n2318_13878.n56 5.97853
R23049 a_n2318_13878.n55 a_n2318_13878.n4 77.6622
R23050 a_n2318_13878.n4 a_n2318_13878.n54 72.3034
R23051 a_n2318_13878.n89 a_n2318_13878.n53 20.9683
R23052 a_n2318_13878.n7 a_n2318_13878.n53 70.1674
R23053 a_n2318_13878.n72 a_n2318_13878.n64 20.9683
R23054 a_n2318_13878.n2 a_n2318_13878.n63 72.3034
R23055 a_n2318_13878.n63 a_n2318_13878.n71 16.6962
R23056 a_n2318_13878.n62 a_n2318_13878.n2 77.6622
R23057 a_n2318_13878.n73 a_n2318_13878.n62 5.97853
R23058 a_n2318_13878.n61 a_n2318_13878.n0 77.6622
R23059 a_n2318_13878.n0 a_n2318_13878.n60 72.3034
R23060 a_n2318_13878.n75 a_n2318_13878.n59 20.9683
R23061 a_n2318_13878.n3 a_n2318_13878.n59 70.1674
R23062 a_n2318_13878.n25 a_n2318_13878.n84 81.2902
R23063 a_n2318_13878.n23 a_n2318_13878.n79 81.2902
R23064 a_n2318_13878.n22 a_n2318_13878.n76 81.2902
R23065 a_n2318_13878.n25 a_n2318_13878.n85 80.9324
R23066 a_n2318_13878.n25 a_n2318_13878.n83 80.9324
R23067 a_n2318_13878.n24 a_n2318_13878.n82 80.9324
R23068 a_n2318_13878.n24 a_n2318_13878.n81 80.9324
R23069 a_n2318_13878.n23 a_n2318_13878.n80 80.9324
R23070 a_n2318_13878.n23 a_n2318_13878.n78 80.9324
R23071 a_n2318_13878.n22 a_n2318_13878.n77 80.9324
R23072 a_n2318_13878.n29 a_n2318_13878.t24 74.6477
R23073 a_n2318_13878.n26 a_n2318_13878.t40 74.6477
R23074 a_n2318_13878.n27 a_n2318_13878.t36 74.2899
R23075 a_n2318_13878.n28 a_n2318_13878.t48 74.2897
R23076 a_n2318_13878.n28 a_n2318_13878.n118 70.6783
R23077 a_n2318_13878.n29 a_n2318_13878.n65 70.6783
R23078 a_n2318_13878.n26 a_n2318_13878.n90 70.6783
R23079 a_n2318_13878.n26 a_n2318_13878.n91 70.6783
R23080 a_n2318_13878.n27 a_n2318_13878.n92 70.6783
R23081 a_n2318_13878.n119 a_n2318_13878.n29 70.6782
R23082 a_n2318_13878.n74 a_n2318_13878.n73 48.2005
R23083 a_n2318_13878.n64 a_n2318_13878.t54 533.335
R23084 a_n2318_13878.n88 a_n2318_13878.n87 48.2005
R23085 a_n2318_13878.n58 a_n2318_13878.t39 533.335
R23086 a_n2318_13878.n115 a_n2318_13878.n114 48.2005
R23087 a_n2318_13878.t47 a_n2318_13878.n43 533.335
R23088 a_n2318_13878.n110 a_n2318_13878.n109 48.2005
R23089 a_n2318_13878.t55 a_n2318_13878.n36 533.335
R23090 a_n2318_13878.n99 a_n2318_13878.n98 48.2005
R23091 a_n2318_13878.t74 a_n2318_13878.n52 533.335
R23092 a_n2318_13878.n101 a_n2318_13878.n100 48.2005
R23093 a_n2318_13878.t81 a_n2318_13878.n49 533.335
R23094 a_n2318_13878.n103 a_n2318_13878.n102 48.2005
R23095 a_n2318_13878.t68 a_n2318_13878.n47 533.335
R23096 a_n2318_13878.n105 a_n2318_13878.n104 48.2005
R23097 a_n2318_13878.t64 a_n2318_13878.n45 533.335
R23098 a_n2318_13878.n60 a_n2318_13878.n70 16.6962
R23099 a_n2318_13878.n72 a_n2318_13878.n63 27.6507
R23100 a_n2318_13878.n54 a_n2318_13878.n68 16.6962
R23101 a_n2318_13878.n86 a_n2318_13878.n57 27.6507
R23102 a_n2318_13878.n113 a_n2318_13878.n39 16.6962
R23103 a_n2318_13878.n116 a_n2318_13878.n42 27.6507
R23104 a_n2318_13878.n108 a_n2318_13878.n32 16.6962
R23105 a_n2318_13878.n111 a_n2318_13878.n35 27.6507
R23106 a_n2318_13878.n61 a_n2318_13878.n70 41.7634
R23107 a_n2318_13878.n55 a_n2318_13878.n68 41.7634
R23108 a_n2318_13878.n113 a_n2318_13878.n40 41.7634
R23109 a_n2318_13878.n108 a_n2318_13878.n33 41.7634
R23110 a_n2318_13878.n24 a_n2318_13878.n23 31.238
R23111 a_n2318_13878.n50 a_n2318_13878.n97 35.3134
R23112 a_n2318_13878.n48 a_n2318_13878.n96 35.3134
R23113 a_n2318_13878.n46 a_n2318_13878.n95 35.3134
R23114 a_n2318_13878.n44 a_n2318_13878.n94 35.3134
R23115 a_n2318_13878.n5 a_n2318_13878.n25 23.891
R23116 a_n2318_13878.n31 a_n2318_13878.n106 12.705
R23117 a_n2318_13878.n1 a_n2318_13878.n51 12.5005
R23118 a_n2318_13878.n61 a_n2318_13878.n74 5.97853
R23119 a_n2318_13878.n62 a_n2318_13878.n71 41.7634
R23120 a_n2318_13878.n55 a_n2318_13878.n88 5.97853
R23121 a_n2318_13878.n56 a_n2318_13878.n69 41.7634
R23122 a_n2318_13878.n114 a_n2318_13878.n40 5.97853
R23123 a_n2318_13878.n66 a_n2318_13878.n41 41.7634
R23124 a_n2318_13878.n109 a_n2318_13878.n33 5.97853
R23125 a_n2318_13878.n67 a_n2318_13878.n34 41.7634
R23126 a_n2318_13878.n93 a_n2318_13878.n7 11.1956
R23127 a_n2318_13878.n75 a_n2318_13878.n60 27.6507
R23128 a_n2318_13878.n89 a_n2318_13878.n54 27.6507
R23129 a_n2318_13878.n39 a_n2318_13878.n112 27.6507
R23130 a_n2318_13878.n32 a_n2318_13878.n107 27.6507
R23131 a_n2318_13878.n28 a_n2318_13878.n117 9.85898
R23132 a_n2318_13878.n8 a_n2318_13878.n51 8.73345
R23133 a_n2318_13878.n106 a_n2318_13878.n15 8.73345
R23134 a_n2318_13878.n117 a_n2318_13878.n16 7.36035
R23135 a_n2318_13878.n93 a_n2318_13878.n27 6.01559
R23136 a_n2318_13878.n117 a_n2318_13878.n51 5.3452
R23137 a_n2318_13878.n38 a_n2318_13878.n19 4.01186
R23138 a_n2318_13878.n5 a_n2318_13878.n3 3.76565
R23139 a_n2318_13878.n118 a_n2318_13878.t38 3.61217
R23140 a_n2318_13878.n118 a_n2318_13878.t42 3.61217
R23141 a_n2318_13878.n65 a_n2318_13878.t32 3.61217
R23142 a_n2318_13878.n65 a_n2318_13878.t20 3.61217
R23143 a_n2318_13878.n90 a_n2318_13878.t46 3.61217
R23144 a_n2318_13878.n90 a_n2318_13878.t28 3.61217
R23145 a_n2318_13878.n91 a_n2318_13878.t34 3.61217
R23146 a_n2318_13878.n91 a_n2318_13878.t26 3.61217
R23147 a_n2318_13878.n92 a_n2318_13878.t44 3.61217
R23148 a_n2318_13878.n92 a_n2318_13878.t22 3.61217
R23149 a_n2318_13878.n119 a_n2318_13878.t30 3.61217
R23150 a_n2318_13878.t18 a_n2318_13878.n119 3.61217
R23151 a_n2318_13878.n84 a_n2318_13878.t4 2.82907
R23152 a_n2318_13878.n84 a_n2318_13878.t2 2.82907
R23153 a_n2318_13878.n85 a_n2318_13878.t7 2.82907
R23154 a_n2318_13878.n85 a_n2318_13878.t16 2.82907
R23155 a_n2318_13878.n83 a_n2318_13878.t3 2.82907
R23156 a_n2318_13878.n83 a_n2318_13878.t1 2.82907
R23157 a_n2318_13878.n82 a_n2318_13878.t51 2.82907
R23158 a_n2318_13878.n82 a_n2318_13878.t50 2.82907
R23159 a_n2318_13878.n81 a_n2318_13878.t15 2.82907
R23160 a_n2318_13878.n81 a_n2318_13878.t6 2.82907
R23161 a_n2318_13878.n79 a_n2318_13878.t10 2.82907
R23162 a_n2318_13878.n79 a_n2318_13878.t5 2.82907
R23163 a_n2318_13878.n80 a_n2318_13878.t14 2.82907
R23164 a_n2318_13878.n80 a_n2318_13878.t49 2.82907
R23165 a_n2318_13878.n78 a_n2318_13878.t13 2.82907
R23166 a_n2318_13878.n78 a_n2318_13878.t0 2.82907
R23167 a_n2318_13878.n77 a_n2318_13878.t9 2.82907
R23168 a_n2318_13878.n77 a_n2318_13878.t8 2.82907
R23169 a_n2318_13878.n76 a_n2318_13878.t12 2.82907
R23170 a_n2318_13878.n76 a_n2318_13878.t11 2.82907
R23171 a_n2318_13878.n106 a_n2318_13878.n93 1.30542
R23172 a_n2318_13878.n29 a_n2318_13878.n28 1.07378
R23173 a_n2318_13878.n27 a_n2318_13878.n26 1.07378
R23174 a_n2318_13878.n25 a_n2318_13878.n24 1.07378
R23175 a_n2318_13878.n12 a_n2318_13878.n11 1.04595
R23176 a_n2318_13878.n6 a_n2318_13878.n5 0.966409
R23177 a_n2318_13878.n21 a_n2318_13878.n20 0.758076
R23178 a_n2318_13878.n20 a_n2318_13878.n19 0.758076
R23179 a_n2318_13878.n18 a_n2318_13878.n17 0.758076
R23180 a_n2318_13878.n17 a_n2318_13878.n16 0.758076
R23181 a_n2318_13878.n15 a_n2318_13878.n14 0.758076
R23182 a_n2318_13878.n13 a_n2318_13878.n12 0.758076
R23183 a_n2318_13878.n11 a_n2318_13878.n10 0.758076
R23184 a_n2318_13878.n9 a_n2318_13878.n8 0.758076
R23185 a_n2318_13878.n6 a_n2318_13878.n4 0.758076
R23186 a_n2318_13878.n2 a_n2318_13878.n0 0.758076
R23187 a_n2318_13878.n2 a_n2318_13878.n1 0.758076
R23188 a_n2318_13878.n23 a_n2318_13878.n22 0.716017
R23189 a_n2318_13878.n14 a_n2318_13878.n13 0.67853
R23190 a_n2318_13878.n10 a_n2318_13878.n9 0.67853
R23191 a_n2318_13878.n0 a_n2318_13878.n3 0.568682
R23192 a_n2318_13878.n4 a_n2318_13878.n7 0.568682
R23193 a_n2318_13878.n38 a_n2318_13878.n18 0.568682
R23194 a_n2318_13878.n31 a_n2318_13878.n21 0.568682
R23195 a_n2140_13878.n2 a_n2140_13878.n0 98.9633
R23196 a_n2140_13878.n5 a_n2140_13878.n3 98.7517
R23197 a_n2140_13878.n2 a_n2140_13878.n1 98.6055
R23198 a_n2140_13878.n9 a_n2140_13878.n8 98.6055
R23199 a_n2140_13878.n7 a_n2140_13878.n6 98.6055
R23200 a_n2140_13878.n5 a_n2140_13878.n4 98.6055
R23201 a_n2140_13878.n21 a_n2140_13878.n20 98.6054
R23202 a_n2140_13878.n19 a_n2140_13878.n18 98.6054
R23203 a_n2140_13878.n11 a_n2140_13878.t1 74.6477
R23204 a_n2140_13878.n16 a_n2140_13878.t2 74.2899
R23205 a_n2140_13878.n13 a_n2140_13878.t3 74.2899
R23206 a_n2140_13878.n12 a_n2140_13878.t0 74.2899
R23207 a_n2140_13878.n15 a_n2140_13878.n14 70.6783
R23208 a_n2140_13878.n11 a_n2140_13878.n10 70.6783
R23209 a_n2140_13878.n17 a_n2140_13878.n9 14.2849
R23210 a_n2140_13878.n19 a_n2140_13878.n17 11.9339
R23211 a_n2140_13878.n17 a_n2140_13878.n16 6.95632
R23212 a_n2140_13878.n18 a_n2140_13878.t14 3.61217
R23213 a_n2140_13878.n18 a_n2140_13878.t15 3.61217
R23214 a_n2140_13878.n1 a_n2140_13878.t8 3.61217
R23215 a_n2140_13878.n1 a_n2140_13878.t16 3.61217
R23216 a_n2140_13878.n0 a_n2140_13878.t19 3.61217
R23217 a_n2140_13878.n0 a_n2140_13878.t23 3.61217
R23218 a_n2140_13878.n14 a_n2140_13878.t6 3.61217
R23219 a_n2140_13878.n14 a_n2140_13878.t7 3.61217
R23220 a_n2140_13878.n10 a_n2140_13878.t4 3.61217
R23221 a_n2140_13878.n10 a_n2140_13878.t5 3.61217
R23222 a_n2140_13878.n8 a_n2140_13878.t17 3.61217
R23223 a_n2140_13878.n8 a_n2140_13878.t9 3.61217
R23224 a_n2140_13878.n6 a_n2140_13878.t20 3.61217
R23225 a_n2140_13878.n6 a_n2140_13878.t11 3.61217
R23226 a_n2140_13878.n4 a_n2140_13878.t10 3.61217
R23227 a_n2140_13878.n4 a_n2140_13878.t12 3.61217
R23228 a_n2140_13878.n3 a_n2140_13878.t18 3.61217
R23229 a_n2140_13878.n3 a_n2140_13878.t13 3.61217
R23230 a_n2140_13878.n21 a_n2140_13878.t21 3.61217
R23231 a_n2140_13878.t22 a_n2140_13878.n21 3.61217
R23232 a_n2140_13878.n12 a_n2140_13878.n11 0.358259
R23233 a_n2140_13878.n15 a_n2140_13878.n13 0.358259
R23234 a_n2140_13878.n16 a_n2140_13878.n15 0.358259
R23235 a_n2140_13878.n20 a_n2140_13878.n2 0.358259
R23236 a_n2140_13878.n20 a_n2140_13878.n19 0.358259
R23237 a_n2140_13878.n7 a_n2140_13878.n5 0.146627
R23238 a_n2140_13878.n9 a_n2140_13878.n7 0.146627
R23239 a_n2140_13878.n13 a_n2140_13878.n12 0.101793
R23240 outputibias.n27 outputibias.n1 289.615
R23241 outputibias.n58 outputibias.n32 289.615
R23242 outputibias.n90 outputibias.n64 289.615
R23243 outputibias.n122 outputibias.n96 289.615
R23244 outputibias.n28 outputibias.n27 185
R23245 outputibias.n26 outputibias.n25 185
R23246 outputibias.n5 outputibias.n4 185
R23247 outputibias.n20 outputibias.n19 185
R23248 outputibias.n18 outputibias.n17 185
R23249 outputibias.n9 outputibias.n8 185
R23250 outputibias.n12 outputibias.n11 185
R23251 outputibias.n59 outputibias.n58 185
R23252 outputibias.n57 outputibias.n56 185
R23253 outputibias.n36 outputibias.n35 185
R23254 outputibias.n51 outputibias.n50 185
R23255 outputibias.n49 outputibias.n48 185
R23256 outputibias.n40 outputibias.n39 185
R23257 outputibias.n43 outputibias.n42 185
R23258 outputibias.n91 outputibias.n90 185
R23259 outputibias.n89 outputibias.n88 185
R23260 outputibias.n68 outputibias.n67 185
R23261 outputibias.n83 outputibias.n82 185
R23262 outputibias.n81 outputibias.n80 185
R23263 outputibias.n72 outputibias.n71 185
R23264 outputibias.n75 outputibias.n74 185
R23265 outputibias.n123 outputibias.n122 185
R23266 outputibias.n121 outputibias.n120 185
R23267 outputibias.n100 outputibias.n99 185
R23268 outputibias.n115 outputibias.n114 185
R23269 outputibias.n113 outputibias.n112 185
R23270 outputibias.n104 outputibias.n103 185
R23271 outputibias.n107 outputibias.n106 185
R23272 outputibias.n0 outputibias.t9 178.945
R23273 outputibias.n133 outputibias.t10 177.018
R23274 outputibias.n132 outputibias.t11 177.018
R23275 outputibias.n0 outputibias.t8 177.018
R23276 outputibias.t7 outputibias.n10 147.661
R23277 outputibias.t1 outputibias.n41 147.661
R23278 outputibias.t3 outputibias.n73 147.661
R23279 outputibias.t5 outputibias.n105 147.661
R23280 outputibias.n128 outputibias.t6 132.363
R23281 outputibias.n128 outputibias.t0 130.436
R23282 outputibias.n129 outputibias.t2 130.436
R23283 outputibias.n130 outputibias.t4 130.436
R23284 outputibias.n27 outputibias.n26 104.615
R23285 outputibias.n26 outputibias.n4 104.615
R23286 outputibias.n19 outputibias.n4 104.615
R23287 outputibias.n19 outputibias.n18 104.615
R23288 outputibias.n18 outputibias.n8 104.615
R23289 outputibias.n11 outputibias.n8 104.615
R23290 outputibias.n58 outputibias.n57 104.615
R23291 outputibias.n57 outputibias.n35 104.615
R23292 outputibias.n50 outputibias.n35 104.615
R23293 outputibias.n50 outputibias.n49 104.615
R23294 outputibias.n49 outputibias.n39 104.615
R23295 outputibias.n42 outputibias.n39 104.615
R23296 outputibias.n90 outputibias.n89 104.615
R23297 outputibias.n89 outputibias.n67 104.615
R23298 outputibias.n82 outputibias.n67 104.615
R23299 outputibias.n82 outputibias.n81 104.615
R23300 outputibias.n81 outputibias.n71 104.615
R23301 outputibias.n74 outputibias.n71 104.615
R23302 outputibias.n122 outputibias.n121 104.615
R23303 outputibias.n121 outputibias.n99 104.615
R23304 outputibias.n114 outputibias.n99 104.615
R23305 outputibias.n114 outputibias.n113 104.615
R23306 outputibias.n113 outputibias.n103 104.615
R23307 outputibias.n106 outputibias.n103 104.615
R23308 outputibias.n63 outputibias.n31 95.6354
R23309 outputibias.n63 outputibias.n62 94.6732
R23310 outputibias.n95 outputibias.n94 94.6732
R23311 outputibias.n127 outputibias.n126 94.6732
R23312 outputibias.n11 outputibias.t7 52.3082
R23313 outputibias.n42 outputibias.t1 52.3082
R23314 outputibias.n74 outputibias.t3 52.3082
R23315 outputibias.n106 outputibias.t5 52.3082
R23316 outputibias.n12 outputibias.n10 15.6674
R23317 outputibias.n43 outputibias.n41 15.6674
R23318 outputibias.n75 outputibias.n73 15.6674
R23319 outputibias.n107 outputibias.n105 15.6674
R23320 outputibias.n13 outputibias.n9 12.8005
R23321 outputibias.n44 outputibias.n40 12.8005
R23322 outputibias.n76 outputibias.n72 12.8005
R23323 outputibias.n108 outputibias.n104 12.8005
R23324 outputibias.n17 outputibias.n16 12.0247
R23325 outputibias.n48 outputibias.n47 12.0247
R23326 outputibias.n80 outputibias.n79 12.0247
R23327 outputibias.n112 outputibias.n111 12.0247
R23328 outputibias.n20 outputibias.n7 11.249
R23329 outputibias.n51 outputibias.n38 11.249
R23330 outputibias.n83 outputibias.n70 11.249
R23331 outputibias.n115 outputibias.n102 11.249
R23332 outputibias.n21 outputibias.n5 10.4732
R23333 outputibias.n52 outputibias.n36 10.4732
R23334 outputibias.n84 outputibias.n68 10.4732
R23335 outputibias.n116 outputibias.n100 10.4732
R23336 outputibias.n25 outputibias.n24 9.69747
R23337 outputibias.n56 outputibias.n55 9.69747
R23338 outputibias.n88 outputibias.n87 9.69747
R23339 outputibias.n120 outputibias.n119 9.69747
R23340 outputibias.n31 outputibias.n30 9.45567
R23341 outputibias.n62 outputibias.n61 9.45567
R23342 outputibias.n94 outputibias.n93 9.45567
R23343 outputibias.n126 outputibias.n125 9.45567
R23344 outputibias.n30 outputibias.n29 9.3005
R23345 outputibias.n3 outputibias.n2 9.3005
R23346 outputibias.n24 outputibias.n23 9.3005
R23347 outputibias.n22 outputibias.n21 9.3005
R23348 outputibias.n7 outputibias.n6 9.3005
R23349 outputibias.n16 outputibias.n15 9.3005
R23350 outputibias.n14 outputibias.n13 9.3005
R23351 outputibias.n61 outputibias.n60 9.3005
R23352 outputibias.n34 outputibias.n33 9.3005
R23353 outputibias.n55 outputibias.n54 9.3005
R23354 outputibias.n53 outputibias.n52 9.3005
R23355 outputibias.n38 outputibias.n37 9.3005
R23356 outputibias.n47 outputibias.n46 9.3005
R23357 outputibias.n45 outputibias.n44 9.3005
R23358 outputibias.n93 outputibias.n92 9.3005
R23359 outputibias.n66 outputibias.n65 9.3005
R23360 outputibias.n87 outputibias.n86 9.3005
R23361 outputibias.n85 outputibias.n84 9.3005
R23362 outputibias.n70 outputibias.n69 9.3005
R23363 outputibias.n79 outputibias.n78 9.3005
R23364 outputibias.n77 outputibias.n76 9.3005
R23365 outputibias.n125 outputibias.n124 9.3005
R23366 outputibias.n98 outputibias.n97 9.3005
R23367 outputibias.n119 outputibias.n118 9.3005
R23368 outputibias.n117 outputibias.n116 9.3005
R23369 outputibias.n102 outputibias.n101 9.3005
R23370 outputibias.n111 outputibias.n110 9.3005
R23371 outputibias.n109 outputibias.n108 9.3005
R23372 outputibias.n28 outputibias.n3 8.92171
R23373 outputibias.n59 outputibias.n34 8.92171
R23374 outputibias.n91 outputibias.n66 8.92171
R23375 outputibias.n123 outputibias.n98 8.92171
R23376 outputibias.n29 outputibias.n1 8.14595
R23377 outputibias.n60 outputibias.n32 8.14595
R23378 outputibias.n92 outputibias.n64 8.14595
R23379 outputibias.n124 outputibias.n96 8.14595
R23380 outputibias.n31 outputibias.n1 5.81868
R23381 outputibias.n62 outputibias.n32 5.81868
R23382 outputibias.n94 outputibias.n64 5.81868
R23383 outputibias.n126 outputibias.n96 5.81868
R23384 outputibias.n131 outputibias.n130 5.20947
R23385 outputibias.n29 outputibias.n28 5.04292
R23386 outputibias.n60 outputibias.n59 5.04292
R23387 outputibias.n92 outputibias.n91 5.04292
R23388 outputibias.n124 outputibias.n123 5.04292
R23389 outputibias.n131 outputibias.n127 4.42209
R23390 outputibias.n14 outputibias.n10 4.38594
R23391 outputibias.n45 outputibias.n41 4.38594
R23392 outputibias.n77 outputibias.n73 4.38594
R23393 outputibias.n109 outputibias.n105 4.38594
R23394 outputibias.n132 outputibias.n131 4.28454
R23395 outputibias.n25 outputibias.n3 4.26717
R23396 outputibias.n56 outputibias.n34 4.26717
R23397 outputibias.n88 outputibias.n66 4.26717
R23398 outputibias.n120 outputibias.n98 4.26717
R23399 outputibias.n24 outputibias.n5 3.49141
R23400 outputibias.n55 outputibias.n36 3.49141
R23401 outputibias.n87 outputibias.n68 3.49141
R23402 outputibias.n119 outputibias.n100 3.49141
R23403 outputibias.n21 outputibias.n20 2.71565
R23404 outputibias.n52 outputibias.n51 2.71565
R23405 outputibias.n84 outputibias.n83 2.71565
R23406 outputibias.n116 outputibias.n115 2.71565
R23407 outputibias.n17 outputibias.n7 1.93989
R23408 outputibias.n48 outputibias.n38 1.93989
R23409 outputibias.n80 outputibias.n70 1.93989
R23410 outputibias.n112 outputibias.n102 1.93989
R23411 outputibias.n130 outputibias.n129 1.9266
R23412 outputibias.n129 outputibias.n128 1.9266
R23413 outputibias.n133 outputibias.n132 1.92658
R23414 outputibias.n134 outputibias.n133 1.29913
R23415 outputibias.n16 outputibias.n9 1.16414
R23416 outputibias.n47 outputibias.n40 1.16414
R23417 outputibias.n79 outputibias.n72 1.16414
R23418 outputibias.n111 outputibias.n104 1.16414
R23419 outputibias.n127 outputibias.n95 0.962709
R23420 outputibias.n95 outputibias.n63 0.962709
R23421 outputibias.n13 outputibias.n12 0.388379
R23422 outputibias.n44 outputibias.n43 0.388379
R23423 outputibias.n76 outputibias.n75 0.388379
R23424 outputibias.n108 outputibias.n107 0.388379
R23425 outputibias.n134 outputibias.n0 0.337251
R23426 outputibias outputibias.n134 0.302375
R23427 outputibias.n30 outputibias.n2 0.155672
R23428 outputibias.n23 outputibias.n2 0.155672
R23429 outputibias.n23 outputibias.n22 0.155672
R23430 outputibias.n22 outputibias.n6 0.155672
R23431 outputibias.n15 outputibias.n6 0.155672
R23432 outputibias.n15 outputibias.n14 0.155672
R23433 outputibias.n61 outputibias.n33 0.155672
R23434 outputibias.n54 outputibias.n33 0.155672
R23435 outputibias.n54 outputibias.n53 0.155672
R23436 outputibias.n53 outputibias.n37 0.155672
R23437 outputibias.n46 outputibias.n37 0.155672
R23438 outputibias.n46 outputibias.n45 0.155672
R23439 outputibias.n93 outputibias.n65 0.155672
R23440 outputibias.n86 outputibias.n65 0.155672
R23441 outputibias.n86 outputibias.n85 0.155672
R23442 outputibias.n85 outputibias.n69 0.155672
R23443 outputibias.n78 outputibias.n69 0.155672
R23444 outputibias.n78 outputibias.n77 0.155672
R23445 outputibias.n125 outputibias.n97 0.155672
R23446 outputibias.n118 outputibias.n97 0.155672
R23447 outputibias.n118 outputibias.n117 0.155672
R23448 outputibias.n117 outputibias.n101 0.155672
R23449 outputibias.n110 outputibias.n101 0.155672
R23450 outputibias.n110 outputibias.n109 0.155672
R23451 a_n2318_8322.n9 a_n2318_8322.t7 74.6477
R23452 a_n2318_8322.t26 a_n2318_8322.n22 74.6477
R23453 a_n2318_8322.n1 a_n2318_8322.t25 74.6474
R23454 a_n2318_8322.n16 a_n2318_8322.t12 74.2899
R23455 a_n2318_8322.n6 a_n2318_8322.t15 74.2899
R23456 a_n2318_8322.n10 a_n2318_8322.t5 74.2899
R23457 a_n2318_8322.n11 a_n2318_8322.t8 74.2899
R23458 a_n2318_8322.n14 a_n2318_8322.t9 74.2899
R23459 a_n2318_8322.n22 a_n2318_8322.n21 70.6783
R23460 a_n2318_8322.n20 a_n2318_8322.n19 70.6783
R23461 a_n2318_8322.n18 a_n2318_8322.n17 70.6783
R23462 a_n2318_8322.n1 a_n2318_8322.n0 70.6783
R23463 a_n2318_8322.n3 a_n2318_8322.n2 70.6783
R23464 a_n2318_8322.n5 a_n2318_8322.n4 70.6783
R23465 a_n2318_8322.n9 a_n2318_8322.n8 70.6783
R23466 a_n2318_8322.n13 a_n2318_8322.n12 70.6783
R23467 a_n2318_8322.n16 a_n2318_8322.n15 23.4712
R23468 a_n2318_8322.n7 a_n2318_8322.t3 10.0266
R23469 a_n2318_8322.n15 a_n2318_8322.n14 6.95632
R23470 a_n2318_8322.n7 a_n2318_8322.n6 6.19447
R23471 a_n2318_8322.n15 a_n2318_8322.n7 5.3452
R23472 a_n2318_8322.n21 a_n2318_8322.t14 3.61217
R23473 a_n2318_8322.n21 a_n2318_8322.t13 3.61217
R23474 a_n2318_8322.n19 a_n2318_8322.t23 3.61217
R23475 a_n2318_8322.n19 a_n2318_8322.t18 3.61217
R23476 a_n2318_8322.n17 a_n2318_8322.t21 3.61217
R23477 a_n2318_8322.n17 a_n2318_8322.t20 3.61217
R23478 a_n2318_8322.n0 a_n2318_8322.t22 3.61217
R23479 a_n2318_8322.n0 a_n2318_8322.t19 3.61217
R23480 a_n2318_8322.n2 a_n2318_8322.t16 3.61217
R23481 a_n2318_8322.n2 a_n2318_8322.t27 3.61217
R23482 a_n2318_8322.n4 a_n2318_8322.t24 3.61217
R23483 a_n2318_8322.n4 a_n2318_8322.t17 3.61217
R23484 a_n2318_8322.n8 a_n2318_8322.t11 3.61217
R23485 a_n2318_8322.n8 a_n2318_8322.t10 3.61217
R23486 a_n2318_8322.n12 a_n2318_8322.t6 3.61217
R23487 a_n2318_8322.n12 a_n2318_8322.t4 3.61217
R23488 a_n2318_8322.n6 a_n2318_8322.n5 0.358259
R23489 a_n2318_8322.n5 a_n2318_8322.n3 0.358259
R23490 a_n2318_8322.n3 a_n2318_8322.n1 0.358259
R23491 a_n2318_8322.n14 a_n2318_8322.n13 0.358259
R23492 a_n2318_8322.n13 a_n2318_8322.n11 0.358259
R23493 a_n2318_8322.n10 a_n2318_8322.n9 0.358259
R23494 a_n2318_8322.n18 a_n2318_8322.n16 0.358259
R23495 a_n2318_8322.n20 a_n2318_8322.n18 0.358259
R23496 a_n2318_8322.n22 a_n2318_8322.n20 0.358259
R23497 a_n2318_8322.n11 a_n2318_8322.n10 0.101793
R23498 a_n2318_8322.t2 a_n2318_8322.t1 0.0788333
R23499 a_n2318_8322.t0 a_n2318_8322.t2 0.0631667
R23500 a_n2318_8322.t3 a_n2318_8322.t0 0.0471944
R23501 a_n2318_8322.t3 a_n2318_8322.t1 0.0453889
R23502 output.n41 output.n15 289.615
R23503 output.n72 output.n46 289.615
R23504 output.n104 output.n78 289.615
R23505 output.n136 output.n110 289.615
R23506 output.n77 output.n45 197.26
R23507 output.n77 output.n76 196.298
R23508 output.n109 output.n108 196.298
R23509 output.n141 output.n140 196.298
R23510 output.n42 output.n41 185
R23511 output.n40 output.n39 185
R23512 output.n19 output.n18 185
R23513 output.n34 output.n33 185
R23514 output.n32 output.n31 185
R23515 output.n23 output.n22 185
R23516 output.n26 output.n25 185
R23517 output.n73 output.n72 185
R23518 output.n71 output.n70 185
R23519 output.n50 output.n49 185
R23520 output.n65 output.n64 185
R23521 output.n63 output.n62 185
R23522 output.n54 output.n53 185
R23523 output.n57 output.n56 185
R23524 output.n105 output.n104 185
R23525 output.n103 output.n102 185
R23526 output.n82 output.n81 185
R23527 output.n97 output.n96 185
R23528 output.n95 output.n94 185
R23529 output.n86 output.n85 185
R23530 output.n89 output.n88 185
R23531 output.n137 output.n136 185
R23532 output.n135 output.n134 185
R23533 output.n114 output.n113 185
R23534 output.n129 output.n128 185
R23535 output.n127 output.n126 185
R23536 output.n118 output.n117 185
R23537 output.n121 output.n120 185
R23538 output.t18 output.n24 147.661
R23539 output.t19 output.n55 147.661
R23540 output.t17 output.n87 147.661
R23541 output.t16 output.n119 147.661
R23542 output.n41 output.n40 104.615
R23543 output.n40 output.n18 104.615
R23544 output.n33 output.n18 104.615
R23545 output.n33 output.n32 104.615
R23546 output.n32 output.n22 104.615
R23547 output.n25 output.n22 104.615
R23548 output.n72 output.n71 104.615
R23549 output.n71 output.n49 104.615
R23550 output.n64 output.n49 104.615
R23551 output.n64 output.n63 104.615
R23552 output.n63 output.n53 104.615
R23553 output.n56 output.n53 104.615
R23554 output.n104 output.n103 104.615
R23555 output.n103 output.n81 104.615
R23556 output.n96 output.n81 104.615
R23557 output.n96 output.n95 104.615
R23558 output.n95 output.n85 104.615
R23559 output.n88 output.n85 104.615
R23560 output.n136 output.n135 104.615
R23561 output.n135 output.n113 104.615
R23562 output.n128 output.n113 104.615
R23563 output.n128 output.n127 104.615
R23564 output.n127 output.n117 104.615
R23565 output.n120 output.n117 104.615
R23566 output.n1 output.t10 77.056
R23567 output.n14 output.t11 76.6694
R23568 output.n1 output.n0 72.7095
R23569 output.n3 output.n2 72.7095
R23570 output.n5 output.n4 72.7095
R23571 output.n7 output.n6 72.7095
R23572 output.n9 output.n8 72.7095
R23573 output.n11 output.n10 72.7095
R23574 output.n13 output.n12 72.7095
R23575 output.n25 output.t18 52.3082
R23576 output.n56 output.t19 52.3082
R23577 output.n88 output.t17 52.3082
R23578 output.n120 output.t16 52.3082
R23579 output.n26 output.n24 15.6674
R23580 output.n57 output.n55 15.6674
R23581 output.n89 output.n87 15.6674
R23582 output.n121 output.n119 15.6674
R23583 output.n27 output.n23 12.8005
R23584 output.n58 output.n54 12.8005
R23585 output.n90 output.n86 12.8005
R23586 output.n122 output.n118 12.8005
R23587 output.n31 output.n30 12.0247
R23588 output.n62 output.n61 12.0247
R23589 output.n94 output.n93 12.0247
R23590 output.n126 output.n125 12.0247
R23591 output.n34 output.n21 11.249
R23592 output.n65 output.n52 11.249
R23593 output.n97 output.n84 11.249
R23594 output.n129 output.n116 11.249
R23595 output.n35 output.n19 10.4732
R23596 output.n66 output.n50 10.4732
R23597 output.n98 output.n82 10.4732
R23598 output.n130 output.n114 10.4732
R23599 output.n39 output.n38 9.69747
R23600 output.n70 output.n69 9.69747
R23601 output.n102 output.n101 9.69747
R23602 output.n134 output.n133 9.69747
R23603 output.n45 output.n44 9.45567
R23604 output.n76 output.n75 9.45567
R23605 output.n108 output.n107 9.45567
R23606 output.n140 output.n139 9.45567
R23607 output.n44 output.n43 9.3005
R23608 output.n17 output.n16 9.3005
R23609 output.n38 output.n37 9.3005
R23610 output.n36 output.n35 9.3005
R23611 output.n21 output.n20 9.3005
R23612 output.n30 output.n29 9.3005
R23613 output.n28 output.n27 9.3005
R23614 output.n75 output.n74 9.3005
R23615 output.n48 output.n47 9.3005
R23616 output.n69 output.n68 9.3005
R23617 output.n67 output.n66 9.3005
R23618 output.n52 output.n51 9.3005
R23619 output.n61 output.n60 9.3005
R23620 output.n59 output.n58 9.3005
R23621 output.n107 output.n106 9.3005
R23622 output.n80 output.n79 9.3005
R23623 output.n101 output.n100 9.3005
R23624 output.n99 output.n98 9.3005
R23625 output.n84 output.n83 9.3005
R23626 output.n93 output.n92 9.3005
R23627 output.n91 output.n90 9.3005
R23628 output.n139 output.n138 9.3005
R23629 output.n112 output.n111 9.3005
R23630 output.n133 output.n132 9.3005
R23631 output.n131 output.n130 9.3005
R23632 output.n116 output.n115 9.3005
R23633 output.n125 output.n124 9.3005
R23634 output.n123 output.n122 9.3005
R23635 output.n42 output.n17 8.92171
R23636 output.n73 output.n48 8.92171
R23637 output.n105 output.n80 8.92171
R23638 output.n137 output.n112 8.92171
R23639 output output.n141 8.15037
R23640 output.n43 output.n15 8.14595
R23641 output.n74 output.n46 8.14595
R23642 output.n106 output.n78 8.14595
R23643 output.n138 output.n110 8.14595
R23644 output.n45 output.n15 5.81868
R23645 output.n76 output.n46 5.81868
R23646 output.n108 output.n78 5.81868
R23647 output.n140 output.n110 5.81868
R23648 output.n43 output.n42 5.04292
R23649 output.n74 output.n73 5.04292
R23650 output.n106 output.n105 5.04292
R23651 output.n138 output.n137 5.04292
R23652 output.n28 output.n24 4.38594
R23653 output.n59 output.n55 4.38594
R23654 output.n91 output.n87 4.38594
R23655 output.n123 output.n119 4.38594
R23656 output.n39 output.n17 4.26717
R23657 output.n70 output.n48 4.26717
R23658 output.n102 output.n80 4.26717
R23659 output.n134 output.n112 4.26717
R23660 output.n0 output.t4 3.9605
R23661 output.n0 output.t2 3.9605
R23662 output.n2 output.t9 3.9605
R23663 output.n2 output.t12 3.9605
R23664 output.n4 output.t14 3.9605
R23665 output.n4 output.t6 3.9605
R23666 output.n6 output.t8 3.9605
R23667 output.n6 output.t15 3.9605
R23668 output.n8 output.t0 3.9605
R23669 output.n8 output.t5 3.9605
R23670 output.n10 output.t7 3.9605
R23671 output.n10 output.t13 3.9605
R23672 output.n12 output.t3 3.9605
R23673 output.n12 output.t1 3.9605
R23674 output.n38 output.n19 3.49141
R23675 output.n69 output.n50 3.49141
R23676 output.n101 output.n82 3.49141
R23677 output.n133 output.n114 3.49141
R23678 output.n35 output.n34 2.71565
R23679 output.n66 output.n65 2.71565
R23680 output.n98 output.n97 2.71565
R23681 output.n130 output.n129 2.71565
R23682 output.n31 output.n21 1.93989
R23683 output.n62 output.n52 1.93989
R23684 output.n94 output.n84 1.93989
R23685 output.n126 output.n116 1.93989
R23686 output.n30 output.n23 1.16414
R23687 output.n61 output.n54 1.16414
R23688 output.n93 output.n86 1.16414
R23689 output.n125 output.n118 1.16414
R23690 output.n141 output.n109 0.962709
R23691 output.n109 output.n77 0.962709
R23692 output.n27 output.n26 0.388379
R23693 output.n58 output.n57 0.388379
R23694 output.n90 output.n89 0.388379
R23695 output.n122 output.n121 0.388379
R23696 output.n14 output.n13 0.387128
R23697 output.n13 output.n11 0.387128
R23698 output.n11 output.n9 0.387128
R23699 output.n9 output.n7 0.387128
R23700 output.n7 output.n5 0.387128
R23701 output.n5 output.n3 0.387128
R23702 output.n3 output.n1 0.387128
R23703 output.n44 output.n16 0.155672
R23704 output.n37 output.n16 0.155672
R23705 output.n37 output.n36 0.155672
R23706 output.n36 output.n20 0.155672
R23707 output.n29 output.n20 0.155672
R23708 output.n29 output.n28 0.155672
R23709 output.n75 output.n47 0.155672
R23710 output.n68 output.n47 0.155672
R23711 output.n68 output.n67 0.155672
R23712 output.n67 output.n51 0.155672
R23713 output.n60 output.n51 0.155672
R23714 output.n60 output.n59 0.155672
R23715 output.n107 output.n79 0.155672
R23716 output.n100 output.n79 0.155672
R23717 output.n100 output.n99 0.155672
R23718 output.n99 output.n83 0.155672
R23719 output.n92 output.n83 0.155672
R23720 output.n92 output.n91 0.155672
R23721 output.n139 output.n111 0.155672
R23722 output.n132 output.n111 0.155672
R23723 output.n132 output.n131 0.155672
R23724 output.n131 output.n115 0.155672
R23725 output.n124 output.n115 0.155672
R23726 output.n124 output.n123 0.155672
R23727 output output.n14 0.126227
R23728 plus.n34 plus.t22 436.949
R23729 plus.n8 plus.t12 436.949
R23730 plus.n35 plus.t5 415.966
R23731 plus.n33 plus.t19 415.966
R23732 plus.n41 plus.t23 415.966
R23733 plus.n42 plus.t11 415.966
R23734 plus.n46 plus.t6 415.966
R23735 plus.n47 plus.t10 415.966
R23736 plus.n29 plus.t18 415.966
R23737 plus.n53 plus.t8 415.966
R23738 plus.n54 plus.t15 415.966
R23739 plus.n26 plus.t24 415.966
R23740 plus.n25 plus.t20 415.966
R23741 plus.n1 plus.t7 415.966
R23742 plus.n19 plus.t17 415.966
R23743 plus.n18 plus.t13 415.966
R23744 plus.n4 plus.t21 415.966
R23745 plus.n13 plus.t16 415.966
R23746 plus.n11 plus.t9 415.966
R23747 plus.n7 plus.t14 415.966
R23748 plus.n58 plus.t0 243.97
R23749 plus.n58 plus.n57 223.454
R23750 plus.n60 plus.n59 223.454
R23751 plus.n55 plus.n54 161.3
R23752 plus.n53 plus.n28 161.3
R23753 plus.n52 plus.n51 161.3
R23754 plus.n50 plus.n29 161.3
R23755 plus.n49 plus.n48 161.3
R23756 plus.n47 plus.n30 161.3
R23757 plus.n46 plus.n45 161.3
R23758 plus.n44 plus.n31 161.3
R23759 plus.n43 plus.n42 161.3
R23760 plus.n41 plus.n32 161.3
R23761 plus.n40 plus.n39 161.3
R23762 plus.n38 plus.n33 161.3
R23763 plus.n37 plus.n36 161.3
R23764 plus.n10 plus.n9 161.3
R23765 plus.n11 plus.n6 161.3
R23766 plus.n12 plus.n5 161.3
R23767 plus.n14 plus.n13 161.3
R23768 plus.n15 plus.n4 161.3
R23769 plus.n17 plus.n16 161.3
R23770 plus.n18 plus.n3 161.3
R23771 plus.n19 plus.n2 161.3
R23772 plus.n21 plus.n20 161.3
R23773 plus.n22 plus.n1 161.3
R23774 plus.n24 plus.n23 161.3
R23775 plus.n25 plus.n0 161.3
R23776 plus.n27 plus.n26 161.3
R23777 plus.n37 plus.n34 70.4033
R23778 plus.n9 plus.n8 70.4033
R23779 plus.n42 plus.n41 48.2005
R23780 plus.n47 plus.n46 48.2005
R23781 plus.n54 plus.n53 48.2005
R23782 plus.n26 plus.n25 48.2005
R23783 plus.n19 plus.n18 48.2005
R23784 plus.n13 plus.n4 48.2005
R23785 plus.n40 plus.n33 47.4702
R23786 plus.n48 plus.n29 47.4702
R23787 plus.n20 plus.n1 47.4702
R23788 plus.n12 plus.n11 47.4702
R23789 plus.n56 plus.n55 29.8622
R23790 plus.n36 plus.n33 25.5611
R23791 plus.n52 plus.n29 25.5611
R23792 plus.n24 plus.n1 25.5611
R23793 plus.n11 plus.n10 25.5611
R23794 plus.n42 plus.n31 24.1005
R23795 plus.n46 plus.n31 24.1005
R23796 plus.n18 plus.n17 24.1005
R23797 plus.n17 plus.n4 24.1005
R23798 plus.n36 plus.n35 22.6399
R23799 plus.n53 plus.n52 22.6399
R23800 plus.n25 plus.n24 22.6399
R23801 plus.n10 plus.n7 22.6399
R23802 plus.n35 plus.n34 20.9576
R23803 plus.n8 plus.n7 20.9576
R23804 plus.n57 plus.t3 19.8005
R23805 plus.n57 plus.t2 19.8005
R23806 plus.n59 plus.t4 19.8005
R23807 plus.n59 plus.t1 19.8005
R23808 plus plus.n61 14.6396
R23809 plus.n56 plus.n27 11.7903
R23810 plus.n61 plus.n60 5.40567
R23811 plus.n61 plus.n56 1.188
R23812 plus.n41 plus.n40 0.730803
R23813 plus.n48 plus.n47 0.730803
R23814 plus.n20 plus.n19 0.730803
R23815 plus.n13 plus.n12 0.730803
R23816 plus.n60 plus.n58 0.716017
R23817 plus.n38 plus.n37 0.189894
R23818 plus.n39 plus.n38 0.189894
R23819 plus.n39 plus.n32 0.189894
R23820 plus.n43 plus.n32 0.189894
R23821 plus.n44 plus.n43 0.189894
R23822 plus.n45 plus.n44 0.189894
R23823 plus.n45 plus.n30 0.189894
R23824 plus.n49 plus.n30 0.189894
R23825 plus.n50 plus.n49 0.189894
R23826 plus.n51 plus.n50 0.189894
R23827 plus.n51 plus.n28 0.189894
R23828 plus.n55 plus.n28 0.189894
R23829 plus.n27 plus.n0 0.189894
R23830 plus.n23 plus.n0 0.189894
R23831 plus.n23 plus.n22 0.189894
R23832 plus.n22 plus.n21 0.189894
R23833 plus.n21 plus.n2 0.189894
R23834 plus.n3 plus.n2 0.189894
R23835 plus.n16 plus.n3 0.189894
R23836 plus.n16 plus.n15 0.189894
R23837 plus.n15 plus.n14 0.189894
R23838 plus.n14 plus.n5 0.189894
R23839 plus.n6 plus.n5 0.189894
R23840 plus.n9 plus.n6 0.189894
R23841 a_n2903_n3924.n12 a_n2903_n3924.t26 214.994
R23842 a_n2903_n3924.n1 a_n2903_n3924.t35 214.733
R23843 a_n2903_n3924.n13 a_n2903_n3924.t34 214.321
R23844 a_n2903_n3924.n14 a_n2903_n3924.t40 214.321
R23845 a_n2903_n3924.n15 a_n2903_n3924.t28 214.321
R23846 a_n2903_n3924.n16 a_n2903_n3924.t29 214.321
R23847 a_n2903_n3924.n17 a_n2903_n3924.t41 214.321
R23848 a_n2903_n3924.n12 a_n2903_n3924.t27 214.321
R23849 a_n2903_n3924.n0 a_n2903_n3924.t8 55.8337
R23850 a_n2903_n3924.n2 a_n2903_n3924.t2 55.8337
R23851 a_n2903_n3924.n11 a_n2903_n3924.t43 55.8337
R23852 a_n2903_n3924.n41 a_n2903_n3924.t15 55.8335
R23853 a_n2903_n3924.n39 a_n2903_n3924.t5 55.8335
R23854 a_n2903_n3924.n30 a_n2903_n3924.t38 55.8335
R23855 a_n2903_n3924.n29 a_n2903_n3924.t18 55.8335
R23856 a_n2903_n3924.n20 a_n2903_n3924.t6 55.8335
R23857 a_n2903_n3924.n43 a_n2903_n3924.n42 53.0052
R23858 a_n2903_n3924.n45 a_n2903_n3924.n44 53.0052
R23859 a_n2903_n3924.n47 a_n2903_n3924.n46 53.0052
R23860 a_n2903_n3924.n4 a_n2903_n3924.n3 53.0052
R23861 a_n2903_n3924.n6 a_n2903_n3924.n5 53.0052
R23862 a_n2903_n3924.n8 a_n2903_n3924.n7 53.0052
R23863 a_n2903_n3924.n10 a_n2903_n3924.n9 53.0052
R23864 a_n2903_n3924.n38 a_n2903_n3924.n37 53.0051
R23865 a_n2903_n3924.n36 a_n2903_n3924.n35 53.0051
R23866 a_n2903_n3924.n34 a_n2903_n3924.n33 53.0051
R23867 a_n2903_n3924.n32 a_n2903_n3924.n31 53.0051
R23868 a_n2903_n3924.n28 a_n2903_n3924.n27 53.0051
R23869 a_n2903_n3924.n26 a_n2903_n3924.n25 53.0051
R23870 a_n2903_n3924.n24 a_n2903_n3924.n23 53.0051
R23871 a_n2903_n3924.n22 a_n2903_n3924.n21 53.0051
R23872 a_n2903_n3924.n49 a_n2903_n3924.n48 53.0051
R23873 a_n2903_n3924.n19 a_n2903_n3924.n11 12.1555
R23874 a_n2903_n3924.n41 a_n2903_n3924.n40 12.1555
R23875 a_n2903_n3924.n20 a_n2903_n3924.n19 5.07593
R23876 a_n2903_n3924.n40 a_n2903_n3924.n39 5.07593
R23877 a_n2903_n3924.n42 a_n2903_n3924.t12 2.82907
R23878 a_n2903_n3924.n42 a_n2903_n3924.t22 2.82907
R23879 a_n2903_n3924.n44 a_n2903_n3924.t24 2.82907
R23880 a_n2903_n3924.n44 a_n2903_n3924.t20 2.82907
R23881 a_n2903_n3924.n46 a_n2903_n3924.t7 2.82907
R23882 a_n2903_n3924.n46 a_n2903_n3924.t19 2.82907
R23883 a_n2903_n3924.n3 a_n2903_n3924.t44 2.82907
R23884 a_n2903_n3924.n3 a_n2903_n3924.t4 2.82907
R23885 a_n2903_n3924.n5 a_n2903_n3924.t1 2.82907
R23886 a_n2903_n3924.n5 a_n2903_n3924.t31 2.82907
R23887 a_n2903_n3924.n7 a_n2903_n3924.t46 2.82907
R23888 a_n2903_n3924.n7 a_n2903_n3924.t3 2.82907
R23889 a_n2903_n3924.n9 a_n2903_n3924.t30 2.82907
R23890 a_n2903_n3924.n9 a_n2903_n3924.t47 2.82907
R23891 a_n2903_n3924.n37 a_n2903_n3924.t45 2.82907
R23892 a_n2903_n3924.n37 a_n2903_n3924.t36 2.82907
R23893 a_n2903_n3924.n35 a_n2903_n3924.t0 2.82907
R23894 a_n2903_n3924.n35 a_n2903_n3924.t42 2.82907
R23895 a_n2903_n3924.n33 a_n2903_n3924.t32 2.82907
R23896 a_n2903_n3924.n33 a_n2903_n3924.t39 2.82907
R23897 a_n2903_n3924.n31 a_n2903_n3924.t37 2.82907
R23898 a_n2903_n3924.n31 a_n2903_n3924.t33 2.82907
R23899 a_n2903_n3924.n27 a_n2903_n3924.t21 2.82907
R23900 a_n2903_n3924.n27 a_n2903_n3924.t16 2.82907
R23901 a_n2903_n3924.n25 a_n2903_n3924.t9 2.82907
R23902 a_n2903_n3924.n25 a_n2903_n3924.t14 2.82907
R23903 a_n2903_n3924.n23 a_n2903_n3924.t13 2.82907
R23904 a_n2903_n3924.n23 a_n2903_n3924.t17 2.82907
R23905 a_n2903_n3924.n21 a_n2903_n3924.t10 2.82907
R23906 a_n2903_n3924.n21 a_n2903_n3924.t23 2.82907
R23907 a_n2903_n3924.t25 a_n2903_n3924.n49 2.82907
R23908 a_n2903_n3924.n49 a_n2903_n3924.t11 2.82907
R23909 a_n2903_n3924.n40 a_n2903_n3924.n1 1.95694
R23910 a_n2903_n3924.n19 a_n2903_n3924.n18 1.95694
R23911 a_n2903_n3924.n17 a_n2903_n3924.n16 0.672012
R23912 a_n2903_n3924.n16 a_n2903_n3924.n15 0.672012
R23913 a_n2903_n3924.n15 a_n2903_n3924.n14 0.672012
R23914 a_n2903_n3924.n14 a_n2903_n3924.n13 0.672012
R23915 a_n2903_n3924.n18 a_n2903_n3924.n17 0.40239
R23916 a_n2903_n3924.n22 a_n2903_n3924.n20 0.358259
R23917 a_n2903_n3924.n24 a_n2903_n3924.n22 0.358259
R23918 a_n2903_n3924.n26 a_n2903_n3924.n24 0.358259
R23919 a_n2903_n3924.n28 a_n2903_n3924.n26 0.358259
R23920 a_n2903_n3924.n29 a_n2903_n3924.n28 0.358259
R23921 a_n2903_n3924.n32 a_n2903_n3924.n30 0.358259
R23922 a_n2903_n3924.n34 a_n2903_n3924.n32 0.358259
R23923 a_n2903_n3924.n36 a_n2903_n3924.n34 0.358259
R23924 a_n2903_n3924.n38 a_n2903_n3924.n36 0.358259
R23925 a_n2903_n3924.n39 a_n2903_n3924.n38 0.358259
R23926 a_n2903_n3924.n11 a_n2903_n3924.n10 0.358259
R23927 a_n2903_n3924.n10 a_n2903_n3924.n8 0.358259
R23928 a_n2903_n3924.n8 a_n2903_n3924.n6 0.358259
R23929 a_n2903_n3924.n6 a_n2903_n3924.n4 0.358259
R23930 a_n2903_n3924.n4 a_n2903_n3924.n2 0.358259
R23931 a_n2903_n3924.n48 a_n2903_n3924.n0 0.358259
R23932 a_n2903_n3924.n48 a_n2903_n3924.n47 0.358259
R23933 a_n2903_n3924.n47 a_n2903_n3924.n45 0.358259
R23934 a_n2903_n3924.n45 a_n2903_n3924.n43 0.358259
R23935 a_n2903_n3924.n43 a_n2903_n3924.n41 0.358259
R23936 a_n2903_n3924.n18 a_n2903_n3924.n12 0.270122
R23937 a_n2903_n3924.n13 a_n2903_n3924.n1 0.259948
R23938 a_n2903_n3924.n30 a_n2903_n3924.n29 0.235414
R23939 a_n2903_n3924.n2 a_n2903_n3924.n0 0.235414
R23940 minus.n36 minus.t23 436.949
R23941 minus.n6 minus.t11 436.949
R23942 minus.n54 minus.t18 415.966
R23943 minus.n53 minus.t13 415.966
R23944 minus.n29 minus.t20 415.966
R23945 minus.n47 minus.t10 415.966
R23946 minus.n46 minus.t5 415.966
R23947 minus.n32 minus.t14 415.966
R23948 minus.n41 minus.t9 415.966
R23949 minus.n39 minus.t22 415.966
R23950 minus.n35 minus.t7 415.966
R23951 minus.n7 minus.t15 415.966
R23952 minus.n5 minus.t8 415.966
R23953 minus.n13 minus.t12 415.966
R23954 minus.n14 minus.t21 415.966
R23955 minus.n18 minus.t16 415.966
R23956 minus.n19 minus.t19 415.966
R23957 minus.n1 minus.t6 415.966
R23958 minus.n25 minus.t17 415.966
R23959 minus.n26 minus.t24 415.966
R23960 minus.n60 minus.t1 243.255
R23961 minus.n59 minus.n57 224.169
R23962 minus.n59 minus.n58 223.454
R23963 minus.n38 minus.n37 161.3
R23964 minus.n39 minus.n34 161.3
R23965 minus.n40 minus.n33 161.3
R23966 minus.n42 minus.n41 161.3
R23967 minus.n43 minus.n32 161.3
R23968 minus.n45 minus.n44 161.3
R23969 minus.n46 minus.n31 161.3
R23970 minus.n47 minus.n30 161.3
R23971 minus.n49 minus.n48 161.3
R23972 minus.n50 minus.n29 161.3
R23973 minus.n52 minus.n51 161.3
R23974 minus.n53 minus.n28 161.3
R23975 minus.n55 minus.n54 161.3
R23976 minus.n27 minus.n26 161.3
R23977 minus.n25 minus.n0 161.3
R23978 minus.n24 minus.n23 161.3
R23979 minus.n22 minus.n1 161.3
R23980 minus.n21 minus.n20 161.3
R23981 minus.n19 minus.n2 161.3
R23982 minus.n18 minus.n17 161.3
R23983 minus.n16 minus.n3 161.3
R23984 minus.n15 minus.n14 161.3
R23985 minus.n13 minus.n4 161.3
R23986 minus.n12 minus.n11 161.3
R23987 minus.n10 minus.n5 161.3
R23988 minus.n9 minus.n8 161.3
R23989 minus.n37 minus.n36 70.4033
R23990 minus.n9 minus.n6 70.4033
R23991 minus.n54 minus.n53 48.2005
R23992 minus.n47 minus.n46 48.2005
R23993 minus.n41 minus.n32 48.2005
R23994 minus.n14 minus.n13 48.2005
R23995 minus.n19 minus.n18 48.2005
R23996 minus.n26 minus.n25 48.2005
R23997 minus.n48 minus.n29 47.4702
R23998 minus.n40 minus.n39 47.4702
R23999 minus.n12 minus.n5 47.4702
R24000 minus.n20 minus.n1 47.4702
R24001 minus.n56 minus.n55 30.0782
R24002 minus.n52 minus.n29 25.5611
R24003 minus.n39 minus.n38 25.5611
R24004 minus.n8 minus.n5 25.5611
R24005 minus.n24 minus.n1 25.5611
R24006 minus.n46 minus.n45 24.1005
R24007 minus.n45 minus.n32 24.1005
R24008 minus.n14 minus.n3 24.1005
R24009 minus.n18 minus.n3 24.1005
R24010 minus.n53 minus.n52 22.6399
R24011 minus.n38 minus.n35 22.6399
R24012 minus.n8 minus.n7 22.6399
R24013 minus.n25 minus.n24 22.6399
R24014 minus.n36 minus.n35 20.9576
R24015 minus.n7 minus.n6 20.9576
R24016 minus.n58 minus.t0 19.8005
R24017 minus.n58 minus.t4 19.8005
R24018 minus.n57 minus.t2 19.8005
R24019 minus.n57 minus.t3 19.8005
R24020 minus minus.n61 12.0099
R24021 minus.n56 minus.n27 12.0062
R24022 minus.n61 minus.n60 4.80222
R24023 minus.n61 minus.n56 0.972091
R24024 minus.n48 minus.n47 0.730803
R24025 minus.n41 minus.n40 0.730803
R24026 minus.n13 minus.n12 0.730803
R24027 minus.n20 minus.n19 0.730803
R24028 minus.n60 minus.n59 0.716017
R24029 minus.n55 minus.n28 0.189894
R24030 minus.n51 minus.n28 0.189894
R24031 minus.n51 minus.n50 0.189894
R24032 minus.n50 minus.n49 0.189894
R24033 minus.n49 minus.n30 0.189894
R24034 minus.n31 minus.n30 0.189894
R24035 minus.n44 minus.n31 0.189894
R24036 minus.n44 minus.n43 0.189894
R24037 minus.n43 minus.n42 0.189894
R24038 minus.n42 minus.n33 0.189894
R24039 minus.n34 minus.n33 0.189894
R24040 minus.n37 minus.n34 0.189894
R24041 minus.n10 minus.n9 0.189894
R24042 minus.n11 minus.n10 0.189894
R24043 minus.n11 minus.n4 0.189894
R24044 minus.n15 minus.n4 0.189894
R24045 minus.n16 minus.n15 0.189894
R24046 minus.n17 minus.n16 0.189894
R24047 minus.n17 minus.n2 0.189894
R24048 minus.n21 minus.n2 0.189894
R24049 minus.n22 minus.n21 0.189894
R24050 minus.n23 minus.n22 0.189894
R24051 minus.n23 minus.n0 0.189894
R24052 minus.n27 minus.n0 0.189894
R24053 diffpairibias.n0 diffpairibias.t18 436.822
R24054 diffpairibias.n21 diffpairibias.t19 435.479
R24055 diffpairibias.n20 diffpairibias.t16 435.479
R24056 diffpairibias.n19 diffpairibias.t17 435.479
R24057 diffpairibias.n18 diffpairibias.t21 435.479
R24058 diffpairibias.n0 diffpairibias.t22 435.479
R24059 diffpairibias.n1 diffpairibias.t20 435.479
R24060 diffpairibias.n2 diffpairibias.t23 435.479
R24061 diffpairibias.n10 diffpairibias.t0 377.536
R24062 diffpairibias.n10 diffpairibias.t8 376.193
R24063 diffpairibias.n11 diffpairibias.t10 376.193
R24064 diffpairibias.n12 diffpairibias.t6 376.193
R24065 diffpairibias.n13 diffpairibias.t2 376.193
R24066 diffpairibias.n14 diffpairibias.t12 376.193
R24067 diffpairibias.n15 diffpairibias.t4 376.193
R24068 diffpairibias.n16 diffpairibias.t14 376.193
R24069 diffpairibias.n3 diffpairibias.t1 113.368
R24070 diffpairibias.n3 diffpairibias.t9 112.698
R24071 diffpairibias.n4 diffpairibias.t11 112.698
R24072 diffpairibias.n5 diffpairibias.t7 112.698
R24073 diffpairibias.n6 diffpairibias.t3 112.698
R24074 diffpairibias.n7 diffpairibias.t13 112.698
R24075 diffpairibias.n8 diffpairibias.t5 112.698
R24076 diffpairibias.n9 diffpairibias.t15 112.698
R24077 diffpairibias.n17 diffpairibias.n16 4.77242
R24078 diffpairibias.n17 diffpairibias.n9 4.30807
R24079 diffpairibias.n18 diffpairibias.n17 4.13945
R24080 diffpairibias.n16 diffpairibias.n15 1.34352
R24081 diffpairibias.n15 diffpairibias.n14 1.34352
R24082 diffpairibias.n14 diffpairibias.n13 1.34352
R24083 diffpairibias.n13 diffpairibias.n12 1.34352
R24084 diffpairibias.n12 diffpairibias.n11 1.34352
R24085 diffpairibias.n11 diffpairibias.n10 1.34352
R24086 diffpairibias.n2 diffpairibias.n1 1.34352
R24087 diffpairibias.n1 diffpairibias.n0 1.34352
R24088 diffpairibias.n19 diffpairibias.n18 1.34352
R24089 diffpairibias.n20 diffpairibias.n19 1.34352
R24090 diffpairibias.n21 diffpairibias.n20 1.34352
R24091 diffpairibias.n22 diffpairibias.n21 0.862419
R24092 diffpairibias diffpairibias.n22 0.684875
R24093 diffpairibias.n9 diffpairibias.n8 0.672012
R24094 diffpairibias.n8 diffpairibias.n7 0.672012
R24095 diffpairibias.n7 diffpairibias.n6 0.672012
R24096 diffpairibias.n6 diffpairibias.n5 0.672012
R24097 diffpairibias.n5 diffpairibias.n4 0.672012
R24098 diffpairibias.n4 diffpairibias.n3 0.672012
R24099 diffpairibias.n22 diffpairibias.n2 0.190907
C0 plus commonsourceibias 0.272687f
C1 output outputibias 2.34152f
C2 vdd output 7.23429f
C3 CSoutput output 6.13571f
C4 CSoutput outputibias 0.032386f
C5 vdd CSoutput 0.140911p
C6 commonsourceibias output 0.006808f
C7 minus diffpairibias 2.77e-19
C8 CSoutput minus 3.14657f
C9 vdd plus 0.090721f
C10 plus diffpairibias 2.54e-19
C11 commonsourceibias outputibias 0.003832f
C12 vdd commonsourceibias 0.004218f
C13 CSoutput plus 0.861832f
C14 commonsourceibias diffpairibias 0.052851f
C15 CSoutput commonsourceibias 44.9728f
C16 minus plus 9.21705f
C17 minus commonsourceibias 0.31863f
C18 diffpairibias gnd 48.968338f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.1814p
C22 plus gnd 31.923103f
C23 minus gnd 27.60523f
C24 CSoutput gnd 0.11419p
C25 vdd gnd 0.474282p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.031174f
C74 minus.t6 gnd 0.314946f
C75 minus.n1 gnd 0.145609f
C76 minus.n2 gnd 0.031174f
C77 minus.n3 gnd 0.007074f
C78 minus.n4 gnd 0.031174f
C79 minus.t8 gnd 0.314946f
C80 minus.n5 gnd 0.145609f
C81 minus.t11 gnd 0.321783f
C82 minus.n6 gnd 0.135744f
C83 minus.t15 gnd 0.314946f
C84 minus.n7 gnd 0.145321f
C85 minus.n8 gnd 0.007074f
C86 minus.n9 gnd 0.102316f
C87 minus.n10 gnd 0.031174f
C88 minus.n11 gnd 0.031174f
C89 minus.n12 gnd 0.007074f
C90 minus.t12 gnd 0.314946f
C91 minus.n13 gnd 0.142438f
C92 minus.t21 gnd 0.314946f
C93 minus.n14 gnd 0.145513f
C94 minus.n15 gnd 0.031174f
C95 minus.n16 gnd 0.031174f
C96 minus.n17 gnd 0.031174f
C97 minus.t16 gnd 0.314946f
C98 minus.n18 gnd 0.145513f
C99 minus.t19 gnd 0.314946f
C100 minus.n19 gnd 0.142438f
C101 minus.n20 gnd 0.007074f
C102 minus.n21 gnd 0.031174f
C103 minus.n22 gnd 0.031174f
C104 minus.n23 gnd 0.031174f
C105 minus.n24 gnd 0.007074f
C106 minus.t17 gnd 0.314946f
C107 minus.n25 gnd 0.145321f
C108 minus.t24 gnd 0.314946f
C109 minus.n26 gnd 0.142342f
C110 minus.n27 gnd 0.354613f
C111 minus.n28 gnd 0.031174f
C112 minus.t18 gnd 0.314946f
C113 minus.t13 gnd 0.314946f
C114 minus.t20 gnd 0.314946f
C115 minus.n29 gnd 0.145609f
C116 minus.n30 gnd 0.031174f
C117 minus.t10 gnd 0.314946f
C118 minus.t5 gnd 0.314946f
C119 minus.n31 gnd 0.031174f
C120 minus.t14 gnd 0.314946f
C121 minus.n32 gnd 0.145513f
C122 minus.n33 gnd 0.031174f
C123 minus.t9 gnd 0.314946f
C124 minus.t22 gnd 0.314946f
C125 minus.n34 gnd 0.031174f
C126 minus.t7 gnd 0.314946f
C127 minus.n35 gnd 0.145321f
C128 minus.t23 gnd 0.321783f
C129 minus.n36 gnd 0.135744f
C130 minus.n37 gnd 0.102316f
C131 minus.n38 gnd 0.007074f
C132 minus.n39 gnd 0.145609f
C133 minus.n40 gnd 0.007074f
C134 minus.n41 gnd 0.142438f
C135 minus.n42 gnd 0.031174f
C136 minus.n43 gnd 0.031174f
C137 minus.n44 gnd 0.031174f
C138 minus.n45 gnd 0.007074f
C139 minus.n46 gnd 0.145513f
C140 minus.n47 gnd 0.142438f
C141 minus.n48 gnd 0.007074f
C142 minus.n49 gnd 0.031174f
C143 minus.n50 gnd 0.031174f
C144 minus.n51 gnd 0.031174f
C145 minus.n52 gnd 0.007074f
C146 minus.n53 gnd 0.145321f
C147 minus.n54 gnd 0.142342f
C148 minus.n55 gnd 0.89555f
C149 minus.n56 gnd 1.36609f
C150 minus.t2 gnd 0.00961f
C151 minus.t3 gnd 0.00961f
C152 minus.n57 gnd 0.0316f
C153 minus.t0 gnd 0.00961f
C154 minus.t4 gnd 0.00961f
C155 minus.n58 gnd 0.031167f
C156 minus.n59 gnd 0.265994f
C157 minus.t1 gnd 0.053488f
C158 minus.n60 gnd 0.145151f
C159 minus.n61 gnd 2.29369f
C160 a_n2903_n3924.t11 gnd 0.102414f
C161 a_n2903_n3924.t8 gnd 1.06441f
C162 a_n2903_n3924.n0 gnd 0.361252f
C163 a_n2903_n3924.t35 gnd 1.32447f
C164 a_n2903_n3924.n1 gnd 1.52483f
C165 a_n2903_n3924.t2 gnd 1.06441f
C166 a_n2903_n3924.n2 gnd 0.361252f
C167 a_n2903_n3924.t44 gnd 0.102414f
C168 a_n2903_n3924.t4 gnd 0.102414f
C169 a_n2903_n3924.n3 gnd 0.836435f
C170 a_n2903_n3924.n4 gnd 0.33923f
C171 a_n2903_n3924.t1 gnd 0.102414f
C172 a_n2903_n3924.t31 gnd 0.102414f
C173 a_n2903_n3924.n5 gnd 0.836435f
C174 a_n2903_n3924.n6 gnd 0.33923f
C175 a_n2903_n3924.t46 gnd 0.102414f
C176 a_n2903_n3924.t3 gnd 0.102414f
C177 a_n2903_n3924.n7 gnd 0.836435f
C178 a_n2903_n3924.n8 gnd 0.33923f
C179 a_n2903_n3924.t30 gnd 0.102414f
C180 a_n2903_n3924.t47 gnd 0.102414f
C181 a_n2903_n3924.n9 gnd 0.836435f
C182 a_n2903_n3924.n10 gnd 0.33923f
C183 a_n2903_n3924.t43 gnd 1.06441f
C184 a_n2903_n3924.n11 gnd 0.918548f
C185 a_n2903_n3924.t26 gnd 1.32439f
C186 a_n2903_n3924.t27 gnd 1.32251f
C187 a_n2903_n3924.n12 gnd 1.32305f
C188 a_n2903_n3924.t34 gnd 1.32251f
C189 a_n2903_n3924.n13 gnd 0.715276f
C190 a_n2903_n3924.t40 gnd 1.32251f
C191 a_n2903_n3924.n14 gnd 0.931464f
C192 a_n2903_n3924.t28 gnd 1.32251f
C193 a_n2903_n3924.n15 gnd 0.931464f
C194 a_n2903_n3924.t29 gnd 1.32251f
C195 a_n2903_n3924.n16 gnd 0.931464f
C196 a_n2903_n3924.t41 gnd 1.32251f
C197 a_n2903_n3924.n17 gnd 0.790007f
C198 a_n2903_n3924.n18 gnd 0.50344f
C199 a_n2903_n3924.n19 gnd 0.956044f
C200 a_n2903_n3924.t6 gnd 1.06441f
C201 a_n2903_n3924.n20 gnd 0.583868f
C202 a_n2903_n3924.t10 gnd 0.102414f
C203 a_n2903_n3924.t23 gnd 0.102414f
C204 a_n2903_n3924.n21 gnd 0.836434f
C205 a_n2903_n3924.n22 gnd 0.339231f
C206 a_n2903_n3924.t13 gnd 0.102414f
C207 a_n2903_n3924.t17 gnd 0.102414f
C208 a_n2903_n3924.n23 gnd 0.836434f
C209 a_n2903_n3924.n24 gnd 0.339231f
C210 a_n2903_n3924.t9 gnd 0.102414f
C211 a_n2903_n3924.t14 gnd 0.102414f
C212 a_n2903_n3924.n25 gnd 0.836434f
C213 a_n2903_n3924.n26 gnd 0.339231f
C214 a_n2903_n3924.t21 gnd 0.102414f
C215 a_n2903_n3924.t16 gnd 0.102414f
C216 a_n2903_n3924.n27 gnd 0.836434f
C217 a_n2903_n3924.n28 gnd 0.339231f
C218 a_n2903_n3924.t18 gnd 1.06441f
C219 a_n2903_n3924.n29 gnd 0.361256f
C220 a_n2903_n3924.t38 gnd 1.06441f
C221 a_n2903_n3924.n30 gnd 0.361256f
C222 a_n2903_n3924.t37 gnd 0.102414f
C223 a_n2903_n3924.t33 gnd 0.102414f
C224 a_n2903_n3924.n31 gnd 0.836434f
C225 a_n2903_n3924.n32 gnd 0.339231f
C226 a_n2903_n3924.t32 gnd 0.102414f
C227 a_n2903_n3924.t39 gnd 0.102414f
C228 a_n2903_n3924.n33 gnd 0.836434f
C229 a_n2903_n3924.n34 gnd 0.339231f
C230 a_n2903_n3924.t0 gnd 0.102414f
C231 a_n2903_n3924.t42 gnd 0.102414f
C232 a_n2903_n3924.n35 gnd 0.836434f
C233 a_n2903_n3924.n36 gnd 0.339231f
C234 a_n2903_n3924.t45 gnd 0.102414f
C235 a_n2903_n3924.t36 gnd 0.102414f
C236 a_n2903_n3924.n37 gnd 0.836434f
C237 a_n2903_n3924.n38 gnd 0.339231f
C238 a_n2903_n3924.t5 gnd 1.06441f
C239 a_n2903_n3924.n39 gnd 0.583868f
C240 a_n2903_n3924.n40 gnd 0.956044f
C241 a_n2903_n3924.t15 gnd 1.06441f
C242 a_n2903_n3924.n41 gnd 0.918552f
C243 a_n2903_n3924.t12 gnd 0.102414f
C244 a_n2903_n3924.t22 gnd 0.102414f
C245 a_n2903_n3924.n42 gnd 0.836435f
C246 a_n2903_n3924.n43 gnd 0.33923f
C247 a_n2903_n3924.t24 gnd 0.102414f
C248 a_n2903_n3924.t20 gnd 0.102414f
C249 a_n2903_n3924.n44 gnd 0.836435f
C250 a_n2903_n3924.n45 gnd 0.33923f
C251 a_n2903_n3924.t7 gnd 0.102414f
C252 a_n2903_n3924.t19 gnd 0.102414f
C253 a_n2903_n3924.n46 gnd 0.836435f
C254 a_n2903_n3924.n47 gnd 0.33923f
C255 a_n2903_n3924.n48 gnd 0.339229f
C256 a_n2903_n3924.n49 gnd 0.836436f
C257 a_n2903_n3924.t25 gnd 0.102414f
C258 plus.n0 gnd 0.022616f
C259 plus.t24 gnd 0.228486f
C260 plus.t20 gnd 0.228486f
C261 plus.t7 gnd 0.228486f
C262 plus.n1 gnd 0.105636f
C263 plus.n2 gnd 0.022616f
C264 plus.t17 gnd 0.228486f
C265 plus.n3 gnd 0.022616f
C266 plus.t13 gnd 0.228486f
C267 plus.t21 gnd 0.228486f
C268 plus.n4 gnd 0.105567f
C269 plus.n5 gnd 0.022616f
C270 plus.t16 gnd 0.228486f
C271 plus.n6 gnd 0.022616f
C272 plus.t9 gnd 0.228486f
C273 plus.t14 gnd 0.228486f
C274 plus.n7 gnd 0.105427f
C275 plus.t12 gnd 0.233447f
C276 plus.n8 gnd 0.098479f
C277 plus.n9 gnd 0.074228f
C278 plus.n10 gnd 0.005132f
C279 plus.n11 gnd 0.105636f
C280 plus.n12 gnd 0.005132f
C281 plus.n13 gnd 0.103336f
C282 plus.n14 gnd 0.022616f
C283 plus.n15 gnd 0.022616f
C284 plus.n16 gnd 0.022616f
C285 plus.n17 gnd 0.005132f
C286 plus.n18 gnd 0.105567f
C287 plus.n19 gnd 0.103336f
C288 plus.n20 gnd 0.005132f
C289 plus.n21 gnd 0.022616f
C290 plus.n22 gnd 0.022616f
C291 plus.n23 gnd 0.022616f
C292 plus.n24 gnd 0.005132f
C293 plus.n25 gnd 0.105427f
C294 plus.n26 gnd 0.103266f
C295 plus.n27 gnd 0.251429f
C296 plus.n28 gnd 0.022616f
C297 plus.t18 gnd 0.228486f
C298 plus.n29 gnd 0.105636f
C299 plus.n30 gnd 0.022616f
C300 plus.n31 gnd 0.005132f
C301 plus.t6 gnd 0.228486f
C302 plus.n32 gnd 0.022616f
C303 plus.t19 gnd 0.228486f
C304 plus.n33 gnd 0.105636f
C305 plus.t22 gnd 0.233447f
C306 plus.n34 gnd 0.098479f
C307 plus.t5 gnd 0.228486f
C308 plus.n35 gnd 0.105427f
C309 plus.n36 gnd 0.005132f
C310 plus.n37 gnd 0.074228f
C311 plus.n38 gnd 0.022616f
C312 plus.n39 gnd 0.022616f
C313 plus.n40 gnd 0.005132f
C314 plus.t23 gnd 0.228486f
C315 plus.n41 gnd 0.103336f
C316 plus.t11 gnd 0.228486f
C317 plus.n42 gnd 0.105567f
C318 plus.n43 gnd 0.022616f
C319 plus.n44 gnd 0.022616f
C320 plus.n45 gnd 0.022616f
C321 plus.n46 gnd 0.105567f
C322 plus.t10 gnd 0.228486f
C323 plus.n47 gnd 0.103336f
C324 plus.n48 gnd 0.005132f
C325 plus.n49 gnd 0.022616f
C326 plus.n50 gnd 0.022616f
C327 plus.n51 gnd 0.022616f
C328 plus.n52 gnd 0.005132f
C329 plus.t8 gnd 0.228486f
C330 plus.n53 gnd 0.105427f
C331 plus.t15 gnd 0.228486f
C332 plus.n54 gnd 0.103266f
C333 plus.n55 gnd 0.640615f
C334 plus.n56 gnd 0.982144f
C335 plus.t0 gnd 0.039042f
C336 plus.t3 gnd 0.006972f
C337 plus.t2 gnd 0.006972f
C338 plus.n57 gnd 0.022611f
C339 plus.n58 gnd 0.17553f
C340 plus.t4 gnd 0.006972f
C341 plus.t1 gnd 0.006972f
C342 plus.n59 gnd 0.022611f
C343 plus.n60 gnd 0.131756f
C344 plus.n61 gnd 2.69131f
C345 output.t10 gnd 0.464308f
C346 output.t4 gnd 0.044422f
C347 output.t2 gnd 0.044422f
C348 output.n0 gnd 0.364624f
C349 output.n1 gnd 0.614102f
C350 output.t9 gnd 0.044422f
C351 output.t12 gnd 0.044422f
C352 output.n2 gnd 0.364624f
C353 output.n3 gnd 0.350265f
C354 output.t14 gnd 0.044422f
C355 output.t6 gnd 0.044422f
C356 output.n4 gnd 0.364624f
C357 output.n5 gnd 0.350265f
C358 output.t8 gnd 0.044422f
C359 output.t15 gnd 0.044422f
C360 output.n6 gnd 0.364624f
C361 output.n7 gnd 0.350265f
C362 output.t0 gnd 0.044422f
C363 output.t5 gnd 0.044422f
C364 output.n8 gnd 0.364624f
C365 output.n9 gnd 0.350265f
C366 output.t7 gnd 0.044422f
C367 output.t13 gnd 0.044422f
C368 output.n10 gnd 0.364624f
C369 output.n11 gnd 0.350265f
C370 output.t3 gnd 0.044422f
C371 output.t1 gnd 0.044422f
C372 output.n12 gnd 0.364624f
C373 output.n13 gnd 0.350265f
C374 output.t11 gnd 0.462979f
C375 output.n14 gnd 0.28994f
C376 output.n15 gnd 0.015803f
C377 output.n16 gnd 0.011243f
C378 output.n17 gnd 0.006041f
C379 output.n18 gnd 0.01428f
C380 output.n19 gnd 0.006397f
C381 output.n20 gnd 0.011243f
C382 output.n21 gnd 0.006041f
C383 output.n22 gnd 0.01428f
C384 output.n23 gnd 0.006397f
C385 output.n24 gnd 0.048111f
C386 output.t18 gnd 0.023274f
C387 output.n25 gnd 0.01071f
C388 output.n26 gnd 0.008435f
C389 output.n27 gnd 0.006041f
C390 output.n28 gnd 0.267512f
C391 output.n29 gnd 0.011243f
C392 output.n30 gnd 0.006041f
C393 output.n31 gnd 0.006397f
C394 output.n32 gnd 0.01428f
C395 output.n33 gnd 0.01428f
C396 output.n34 gnd 0.006397f
C397 output.n35 gnd 0.006041f
C398 output.n36 gnd 0.011243f
C399 output.n37 gnd 0.011243f
C400 output.n38 gnd 0.006041f
C401 output.n39 gnd 0.006397f
C402 output.n40 gnd 0.01428f
C403 output.n41 gnd 0.030913f
C404 output.n42 gnd 0.006397f
C405 output.n43 gnd 0.006041f
C406 output.n44 gnd 0.025987f
C407 output.n45 gnd 0.097665f
C408 output.n46 gnd 0.015803f
C409 output.n47 gnd 0.011243f
C410 output.n48 gnd 0.006041f
C411 output.n49 gnd 0.01428f
C412 output.n50 gnd 0.006397f
C413 output.n51 gnd 0.011243f
C414 output.n52 gnd 0.006041f
C415 output.n53 gnd 0.01428f
C416 output.n54 gnd 0.006397f
C417 output.n55 gnd 0.048111f
C418 output.t19 gnd 0.023274f
C419 output.n56 gnd 0.01071f
C420 output.n57 gnd 0.008435f
C421 output.n58 gnd 0.006041f
C422 output.n59 gnd 0.267512f
C423 output.n60 gnd 0.011243f
C424 output.n61 gnd 0.006041f
C425 output.n62 gnd 0.006397f
C426 output.n63 gnd 0.01428f
C427 output.n64 gnd 0.01428f
C428 output.n65 gnd 0.006397f
C429 output.n66 gnd 0.006041f
C430 output.n67 gnd 0.011243f
C431 output.n68 gnd 0.011243f
C432 output.n69 gnd 0.006041f
C433 output.n70 gnd 0.006397f
C434 output.n71 gnd 0.01428f
C435 output.n72 gnd 0.030913f
C436 output.n73 gnd 0.006397f
C437 output.n74 gnd 0.006041f
C438 output.n75 gnd 0.025987f
C439 output.n76 gnd 0.09306f
C440 output.n77 gnd 1.65264f
C441 output.n78 gnd 0.015803f
C442 output.n79 gnd 0.011243f
C443 output.n80 gnd 0.006041f
C444 output.n81 gnd 0.01428f
C445 output.n82 gnd 0.006397f
C446 output.n83 gnd 0.011243f
C447 output.n84 gnd 0.006041f
C448 output.n85 gnd 0.01428f
C449 output.n86 gnd 0.006397f
C450 output.n87 gnd 0.048111f
C451 output.t17 gnd 0.023274f
C452 output.n88 gnd 0.01071f
C453 output.n89 gnd 0.008435f
C454 output.n90 gnd 0.006041f
C455 output.n91 gnd 0.267512f
C456 output.n92 gnd 0.011243f
C457 output.n93 gnd 0.006041f
C458 output.n94 gnd 0.006397f
C459 output.n95 gnd 0.01428f
C460 output.n96 gnd 0.01428f
C461 output.n97 gnd 0.006397f
C462 output.n98 gnd 0.006041f
C463 output.n99 gnd 0.011243f
C464 output.n100 gnd 0.011243f
C465 output.n101 gnd 0.006041f
C466 output.n102 gnd 0.006397f
C467 output.n103 gnd 0.01428f
C468 output.n104 gnd 0.030913f
C469 output.n105 gnd 0.006397f
C470 output.n106 gnd 0.006041f
C471 output.n107 gnd 0.025987f
C472 output.n108 gnd 0.09306f
C473 output.n109 gnd 0.713089f
C474 output.n110 gnd 0.015803f
C475 output.n111 gnd 0.011243f
C476 output.n112 gnd 0.006041f
C477 output.n113 gnd 0.01428f
C478 output.n114 gnd 0.006397f
C479 output.n115 gnd 0.011243f
C480 output.n116 gnd 0.006041f
C481 output.n117 gnd 0.01428f
C482 output.n118 gnd 0.006397f
C483 output.n119 gnd 0.048111f
C484 output.t16 gnd 0.023274f
C485 output.n120 gnd 0.01071f
C486 output.n121 gnd 0.008435f
C487 output.n122 gnd 0.006041f
C488 output.n123 gnd 0.267512f
C489 output.n124 gnd 0.011243f
C490 output.n125 gnd 0.006041f
C491 output.n126 gnd 0.006397f
C492 output.n127 gnd 0.01428f
C493 output.n128 gnd 0.01428f
C494 output.n129 gnd 0.006397f
C495 output.n130 gnd 0.006041f
C496 output.n131 gnd 0.011243f
C497 output.n132 gnd 0.011243f
C498 output.n133 gnd 0.006041f
C499 output.n134 gnd 0.006397f
C500 output.n135 gnd 0.01428f
C501 output.n136 gnd 0.030913f
C502 output.n137 gnd 0.006397f
C503 output.n138 gnd 0.006041f
C504 output.n139 gnd 0.025987f
C505 output.n140 gnd 0.09306f
C506 output.n141 gnd 1.67353f
C507 a_n2318_8322.t1 gnd 39.602997f
C508 a_n2318_8322.t3 gnd 29.1868f
C509 a_n2318_8322.t2 gnd 19.7318f
C510 a_n2318_8322.t0 gnd 39.602997f
C511 a_n2318_8322.t25 gnd 0.896865f
C512 a_n2318_8322.t22 gnd 0.095784f
C513 a_n2318_8322.t19 gnd 0.095784f
C514 a_n2318_8322.n0 gnd 0.674698f
C515 a_n2318_8322.n1 gnd 0.753878f
C516 a_n2318_8322.t16 gnd 0.095784f
C517 a_n2318_8322.t27 gnd 0.095784f
C518 a_n2318_8322.n2 gnd 0.674698f
C519 a_n2318_8322.n3 gnd 0.383035f
C520 a_n2318_8322.t24 gnd 0.095784f
C521 a_n2318_8322.t17 gnd 0.095784f
C522 a_n2318_8322.n4 gnd 0.674698f
C523 a_n2318_8322.n5 gnd 0.383035f
C524 a_n2318_8322.t15 gnd 0.895082f
C525 a_n2318_8322.n6 gnd 0.881139f
C526 a_n2318_8322.n7 gnd 3.71089f
C527 a_n2318_8322.t7 gnd 0.896867f
C528 a_n2318_8322.t11 gnd 0.095784f
C529 a_n2318_8322.t10 gnd 0.095784f
C530 a_n2318_8322.n8 gnd 0.674698f
C531 a_n2318_8322.n9 gnd 0.753876f
C532 a_n2318_8322.t5 gnd 0.895082f
C533 a_n2318_8322.n10 gnd 0.379361f
C534 a_n2318_8322.t8 gnd 0.895082f
C535 a_n2318_8322.n11 gnd 0.379361f
C536 a_n2318_8322.t6 gnd 0.095784f
C537 a_n2318_8322.t4 gnd 0.095784f
C538 a_n2318_8322.n12 gnd 0.674698f
C539 a_n2318_8322.n13 gnd 0.383035f
C540 a_n2318_8322.t9 gnd 0.895082f
C541 a_n2318_8322.n14 gnd 1.07426f
C542 a_n2318_8322.n15 gnd 1.82616f
C543 a_n2318_8322.t12 gnd 0.895082f
C544 a_n2318_8322.n16 gnd 1.55131f
C545 a_n2318_8322.t21 gnd 0.095784f
C546 a_n2318_8322.t20 gnd 0.095784f
C547 a_n2318_8322.n17 gnd 0.674698f
C548 a_n2318_8322.n18 gnd 0.383035f
C549 a_n2318_8322.t23 gnd 0.095784f
C550 a_n2318_8322.t18 gnd 0.095784f
C551 a_n2318_8322.n19 gnd 0.674698f
C552 a_n2318_8322.n20 gnd 0.383035f
C553 a_n2318_8322.t14 gnd 0.095784f
C554 a_n2318_8322.t13 gnd 0.095784f
C555 a_n2318_8322.n21 gnd 0.674698f
C556 a_n2318_8322.n22 gnd 0.753876f
C557 a_n2318_8322.t26 gnd 0.896867f
C558 outputibias.t8 gnd 0.11477f
C559 outputibias.t9 gnd 0.115567f
C560 outputibias.n0 gnd 0.130108f
C561 outputibias.n1 gnd 0.001372f
C562 outputibias.n2 gnd 9.76e-19
C563 outputibias.n3 gnd 5.24e-19
C564 outputibias.n4 gnd 0.001239f
C565 outputibias.n5 gnd 5.55e-19
C566 outputibias.n6 gnd 9.76e-19
C567 outputibias.n7 gnd 5.24e-19
C568 outputibias.n8 gnd 0.001239f
C569 outputibias.n9 gnd 5.55e-19
C570 outputibias.n10 gnd 0.004176f
C571 outputibias.t7 gnd 0.00202f
C572 outputibias.n11 gnd 9.3e-19
C573 outputibias.n12 gnd 7.32e-19
C574 outputibias.n13 gnd 5.24e-19
C575 outputibias.n14 gnd 0.02322f
C576 outputibias.n15 gnd 9.76e-19
C577 outputibias.n16 gnd 5.24e-19
C578 outputibias.n17 gnd 5.55e-19
C579 outputibias.n18 gnd 0.001239f
C580 outputibias.n19 gnd 0.001239f
C581 outputibias.n20 gnd 5.55e-19
C582 outputibias.n21 gnd 5.24e-19
C583 outputibias.n22 gnd 9.76e-19
C584 outputibias.n23 gnd 9.76e-19
C585 outputibias.n24 gnd 5.24e-19
C586 outputibias.n25 gnd 5.55e-19
C587 outputibias.n26 gnd 0.001239f
C588 outputibias.n27 gnd 0.002683f
C589 outputibias.n28 gnd 5.55e-19
C590 outputibias.n29 gnd 5.24e-19
C591 outputibias.n30 gnd 0.002256f
C592 outputibias.n31 gnd 0.005781f
C593 outputibias.n32 gnd 0.001372f
C594 outputibias.n33 gnd 9.76e-19
C595 outputibias.n34 gnd 5.24e-19
C596 outputibias.n35 gnd 0.001239f
C597 outputibias.n36 gnd 5.55e-19
C598 outputibias.n37 gnd 9.76e-19
C599 outputibias.n38 gnd 5.24e-19
C600 outputibias.n39 gnd 0.001239f
C601 outputibias.n40 gnd 5.55e-19
C602 outputibias.n41 gnd 0.004176f
C603 outputibias.t1 gnd 0.00202f
C604 outputibias.n42 gnd 9.3e-19
C605 outputibias.n43 gnd 7.32e-19
C606 outputibias.n44 gnd 5.24e-19
C607 outputibias.n45 gnd 0.02322f
C608 outputibias.n46 gnd 9.76e-19
C609 outputibias.n47 gnd 5.24e-19
C610 outputibias.n48 gnd 5.55e-19
C611 outputibias.n49 gnd 0.001239f
C612 outputibias.n50 gnd 0.001239f
C613 outputibias.n51 gnd 5.55e-19
C614 outputibias.n52 gnd 5.24e-19
C615 outputibias.n53 gnd 9.76e-19
C616 outputibias.n54 gnd 9.76e-19
C617 outputibias.n55 gnd 5.24e-19
C618 outputibias.n56 gnd 5.55e-19
C619 outputibias.n57 gnd 0.001239f
C620 outputibias.n58 gnd 0.002683f
C621 outputibias.n59 gnd 5.55e-19
C622 outputibias.n60 gnd 5.24e-19
C623 outputibias.n61 gnd 0.002256f
C624 outputibias.n62 gnd 0.005197f
C625 outputibias.n63 gnd 0.121892f
C626 outputibias.n64 gnd 0.001372f
C627 outputibias.n65 gnd 9.76e-19
C628 outputibias.n66 gnd 5.24e-19
C629 outputibias.n67 gnd 0.001239f
C630 outputibias.n68 gnd 5.55e-19
C631 outputibias.n69 gnd 9.76e-19
C632 outputibias.n70 gnd 5.24e-19
C633 outputibias.n71 gnd 0.001239f
C634 outputibias.n72 gnd 5.55e-19
C635 outputibias.n73 gnd 0.004176f
C636 outputibias.t3 gnd 0.00202f
C637 outputibias.n74 gnd 9.3e-19
C638 outputibias.n75 gnd 7.32e-19
C639 outputibias.n76 gnd 5.24e-19
C640 outputibias.n77 gnd 0.02322f
C641 outputibias.n78 gnd 9.76e-19
C642 outputibias.n79 gnd 5.24e-19
C643 outputibias.n80 gnd 5.55e-19
C644 outputibias.n81 gnd 0.001239f
C645 outputibias.n82 gnd 0.001239f
C646 outputibias.n83 gnd 5.55e-19
C647 outputibias.n84 gnd 5.24e-19
C648 outputibias.n85 gnd 9.76e-19
C649 outputibias.n86 gnd 9.76e-19
C650 outputibias.n87 gnd 5.24e-19
C651 outputibias.n88 gnd 5.55e-19
C652 outputibias.n89 gnd 0.001239f
C653 outputibias.n90 gnd 0.002683f
C654 outputibias.n91 gnd 5.55e-19
C655 outputibias.n92 gnd 5.24e-19
C656 outputibias.n93 gnd 0.002256f
C657 outputibias.n94 gnd 0.005197f
C658 outputibias.n95 gnd 0.064513f
C659 outputibias.n96 gnd 0.001372f
C660 outputibias.n97 gnd 9.76e-19
C661 outputibias.n98 gnd 5.24e-19
C662 outputibias.n99 gnd 0.001239f
C663 outputibias.n100 gnd 5.55e-19
C664 outputibias.n101 gnd 9.76e-19
C665 outputibias.n102 gnd 5.24e-19
C666 outputibias.n103 gnd 0.001239f
C667 outputibias.n104 gnd 5.55e-19
C668 outputibias.n105 gnd 0.004176f
C669 outputibias.t5 gnd 0.00202f
C670 outputibias.n106 gnd 9.3e-19
C671 outputibias.n107 gnd 7.32e-19
C672 outputibias.n108 gnd 5.24e-19
C673 outputibias.n109 gnd 0.02322f
C674 outputibias.n110 gnd 9.76e-19
C675 outputibias.n111 gnd 5.24e-19
C676 outputibias.n112 gnd 5.55e-19
C677 outputibias.n113 gnd 0.001239f
C678 outputibias.n114 gnd 0.001239f
C679 outputibias.n115 gnd 5.55e-19
C680 outputibias.n116 gnd 5.24e-19
C681 outputibias.n117 gnd 9.76e-19
C682 outputibias.n118 gnd 9.76e-19
C683 outputibias.n119 gnd 5.24e-19
C684 outputibias.n120 gnd 5.55e-19
C685 outputibias.n121 gnd 0.001239f
C686 outputibias.n122 gnd 0.002683f
C687 outputibias.n123 gnd 5.55e-19
C688 outputibias.n124 gnd 5.24e-19
C689 outputibias.n125 gnd 0.002256f
C690 outputibias.n126 gnd 0.005197f
C691 outputibias.n127 gnd 0.084814f
C692 outputibias.t4 gnd 0.108319f
C693 outputibias.t2 gnd 0.108319f
C694 outputibias.t0 gnd 0.108319f
C695 outputibias.t6 gnd 0.109238f
C696 outputibias.n128 gnd 0.134674f
C697 outputibias.n129 gnd 0.07244f
C698 outputibias.n130 gnd 0.079818f
C699 outputibias.n131 gnd 0.164901f
C700 outputibias.t11 gnd 0.11477f
C701 outputibias.n132 gnd 0.067481f
C702 outputibias.t10 gnd 0.11477f
C703 outputibias.n133 gnd 0.065115f
C704 outputibias.n134 gnd 0.029159f
C705 a_n2140_13878.t21 gnd 0.186452f
C706 a_n2140_13878.t19 gnd 0.186452f
C707 a_n2140_13878.t23 gnd 0.186452f
C708 a_n2140_13878.n0 gnd 1.47058f
C709 a_n2140_13878.t8 gnd 0.186452f
C710 a_n2140_13878.t16 gnd 0.186452f
C711 a_n2140_13878.n1 gnd 1.46815f
C712 a_n2140_13878.n2 gnd 1.31969f
C713 a_n2140_13878.t18 gnd 0.186452f
C714 a_n2140_13878.t13 gnd 0.186452f
C715 a_n2140_13878.n3 gnd 1.46971f
C716 a_n2140_13878.t10 gnd 0.186452f
C717 a_n2140_13878.t12 gnd 0.186452f
C718 a_n2140_13878.n4 gnd 1.46815f
C719 a_n2140_13878.n5 gnd 2.05145f
C720 a_n2140_13878.t20 gnd 0.186452f
C721 a_n2140_13878.t11 gnd 0.186452f
C722 a_n2140_13878.n6 gnd 1.46815f
C723 a_n2140_13878.n7 gnd 1.00065f
C724 a_n2140_13878.t17 gnd 0.186452f
C725 a_n2140_13878.t9 gnd 0.186452f
C726 a_n2140_13878.n8 gnd 1.46815f
C727 a_n2140_13878.n9 gnd 4.05307f
C728 a_n2140_13878.t1 gnd 1.74584f
C729 a_n2140_13878.t4 gnd 0.186452f
C730 a_n2140_13878.t5 gnd 0.186452f
C731 a_n2140_13878.n10 gnd 1.31337f
C732 a_n2140_13878.n11 gnd 1.4675f
C733 a_n2140_13878.t0 gnd 1.74237f
C734 a_n2140_13878.n12 gnd 0.738464f
C735 a_n2140_13878.t3 gnd 1.74237f
C736 a_n2140_13878.n13 gnd 0.738464f
C737 a_n2140_13878.t6 gnd 0.186452f
C738 a_n2140_13878.t7 gnd 0.186452f
C739 a_n2140_13878.n14 gnd 1.31337f
C740 a_n2140_13878.n15 gnd 0.745616f
C741 a_n2140_13878.t2 gnd 1.74237f
C742 a_n2140_13878.n16 gnd 2.09116f
C743 a_n2140_13878.n17 gnd 2.85337f
C744 a_n2140_13878.t14 gnd 0.186452f
C745 a_n2140_13878.t15 gnd 0.186452f
C746 a_n2140_13878.n18 gnd 1.46815f
C747 a_n2140_13878.n19 gnd 2.01216f
C748 a_n2140_13878.n20 gnd 0.650496f
C749 a_n2140_13878.n21 gnd 1.46815f
C750 a_n2140_13878.t22 gnd 0.186452f
C751 a_n2318_13878.n0 gnd 0.217886f
C752 a_n2318_13878.n1 gnd 0.753716f
C753 a_n2318_13878.n2 gnd 0.217886f
C754 a_n2318_13878.n3 gnd 0.42604f
C755 a_n2318_13878.n4 gnd 0.217886f
C756 a_n2318_13878.n5 gnd 3.16141f
C757 a_n2318_13878.n6 gnd 0.217886f
C758 a_n2318_13878.n7 gnd 0.674574f
C759 a_n2318_13878.n8 gnd 0.674551f
C760 a_n2318_13878.n9 gnd 0.206738f
C761 a_n2318_13878.n10 gnd 0.152266f
C762 a_n2318_13878.n11 gnd 0.239314f
C763 a_n2318_13878.n12 gnd 0.184843f
C764 a_n2318_13878.n13 gnd 0.206738f
C765 a_n2318_13878.n14 gnd 0.152266f
C766 a_n2318_13878.n15 gnd 0.729022f
C767 a_n2318_13878.n16 gnd 0.51701f
C768 a_n2318_13878.n17 gnd 0.217886f
C769 a_n2318_13878.n18 gnd 0.217886f
C770 a_n2318_13878.n19 gnd 0.447806f
C771 a_n2318_13878.n20 gnd 0.217886f
C772 a_n2318_13878.n21 gnd 0.217886f
C773 a_n2318_13878.n22 gnd 0.733554f
C774 a_n2318_13878.n23 gnd 2.98994f
C775 a_n2318_13878.n24 gnd 2.92523f
C776 a_n2318_13878.n25 gnd 3.7969f
C777 a_n2318_13878.n26 gnd 1.79383f
C778 a_n2318_13878.n27 gnd 1.91464f
C779 a_n2318_13878.n28 gnd 2.09784f
C780 a_n2318_13878.n29 gnd 1.79383f
C781 a_n2318_13878.n30 gnd 0.287827f
C782 a_n2318_13878.n31 gnd 0.766802f
C783 a_n2318_13878.n32 gnd 0.004897f
C784 a_n2318_13878.n33 gnd 0.010591f
C785 a_n2318_13878.n34 gnd 0.010591f
C786 a_n2318_13878.n35 gnd 0.004897f
C787 a_n2318_13878.n36 gnd 0.287827f
C788 a_n2318_13878.n37 gnd 0.287827f
C789 a_n2318_13878.n38 gnd 0.447806f
C790 a_n2318_13878.n39 gnd 0.004897f
C791 a_n2318_13878.n40 gnd 0.010591f
C792 a_n2318_13878.n41 gnd 0.010591f
C793 a_n2318_13878.n42 gnd 0.004897f
C794 a_n2318_13878.n43 gnd 0.287827f
C795 a_n2318_13878.n44 gnd 0.008436f
C796 a_n2318_13878.n45 gnd 0.287827f
C797 a_n2318_13878.n46 gnd 0.008436f
C798 a_n2318_13878.n47 gnd 0.287827f
C799 a_n2318_13878.n48 gnd 0.008436f
C800 a_n2318_13878.n49 gnd 0.287827f
C801 a_n2318_13878.n50 gnd 0.008436f
C802 a_n2318_13878.n51 gnd 1.46328f
C803 a_n2318_13878.n52 gnd 0.287827f
C804 a_n2318_13878.n53 gnd 0.287827f
C805 a_n2318_13878.n54 gnd 0.004897f
C806 a_n2318_13878.n55 gnd 0.010591f
C807 a_n2318_13878.n56 gnd 0.010591f
C808 a_n2318_13878.n57 gnd 0.004897f
C809 a_n2318_13878.n58 gnd 0.287827f
C810 a_n2318_13878.n59 gnd 0.287827f
C811 a_n2318_13878.n60 gnd 0.004897f
C812 a_n2318_13878.n61 gnd 0.010591f
C813 a_n2318_13878.n62 gnd 0.010591f
C814 a_n2318_13878.n63 gnd 0.004897f
C815 a_n2318_13878.n64 gnd 0.287827f
C816 a_n2318_13878.t30 gnd 0.151128f
C817 a_n2318_13878.t24 gnd 1.41509f
C818 a_n2318_13878.t32 gnd 0.151128f
C819 a_n2318_13878.t20 gnd 0.151128f
C820 a_n2318_13878.n65 gnd 1.06455f
C821 a_n2318_13878.t37 gnd 0.702974f
C822 a_n2318_13878.n66 gnd 0.307084f
C823 a_n2318_13878.t29 gnd 0.702974f
C824 a_n2318_13878.t23 gnd 0.714753f
C825 a_n2318_13878.t31 gnd 0.702974f
C826 a_n2318_13878.t62 gnd 0.702974f
C827 a_n2318_13878.n67 gnd 0.307084f
C828 a_n2318_13878.t76 gnd 0.702974f
C829 a_n2318_13878.t78 gnd 0.714753f
C830 a_n2318_13878.t56 gnd 0.702974f
C831 a_n2318_13878.t35 gnd 0.714753f
C832 a_n2318_13878.t43 gnd 0.702974f
C833 a_n2318_13878.t21 gnd 0.702974f
C834 a_n2318_13878.n68 gnd 0.307084f
C835 a_n2318_13878.t33 gnd 0.702974f
C836 a_n2318_13878.t25 gnd 0.702974f
C837 a_n2318_13878.t45 gnd 0.702974f
C838 a_n2318_13878.n69 gnd 0.307084f
C839 a_n2318_13878.t27 gnd 0.702974f
C840 a_n2318_13878.t39 gnd 0.714753f
C841 a_n2318_13878.t82 gnd 0.714753f
C842 a_n2318_13878.t63 gnd 0.702974f
C843 a_n2318_13878.t67 gnd 0.702974f
C844 a_n2318_13878.n70 gnd 0.307084f
C845 a_n2318_13878.t57 gnd 0.702974f
C846 a_n2318_13878.t72 gnd 0.702974f
C847 a_n2318_13878.t79 gnd 0.702974f
C848 a_n2318_13878.n71 gnd 0.307084f
C849 a_n2318_13878.t80 gnd 0.702974f
C850 a_n2318_13878.t54 gnd 0.714753f
C851 a_n2318_13878.n72 gnd 0.309588f
C852 a_n2318_13878.n73 gnd 0.30246f
C853 a_n2318_13878.n74 gnd 0.30246f
C854 a_n2318_13878.n75 gnd 0.309588f
C855 a_n2318_13878.t12 gnd 0.117544f
C856 a_n2318_13878.t11 gnd 0.117544f
C857 a_n2318_13878.n76 gnd 1.04031f
C858 a_n2318_13878.t9 gnd 0.117544f
C859 a_n2318_13878.t8 gnd 0.117544f
C860 a_n2318_13878.n77 gnd 1.03866f
C861 a_n2318_13878.t13 gnd 0.117544f
C862 a_n2318_13878.t0 gnd 0.117544f
C863 a_n2318_13878.n78 gnd 1.03866f
C864 a_n2318_13878.t10 gnd 0.117544f
C865 a_n2318_13878.t5 gnd 0.117544f
C866 a_n2318_13878.n79 gnd 1.04031f
C867 a_n2318_13878.t14 gnd 0.117544f
C868 a_n2318_13878.t49 gnd 0.117544f
C869 a_n2318_13878.n80 gnd 1.03866f
C870 a_n2318_13878.t15 gnd 0.117544f
C871 a_n2318_13878.t6 gnd 0.117544f
C872 a_n2318_13878.n81 gnd 1.03866f
C873 a_n2318_13878.t51 gnd 0.117544f
C874 a_n2318_13878.t50 gnd 0.117544f
C875 a_n2318_13878.n82 gnd 1.03866f
C876 a_n2318_13878.t3 gnd 0.117544f
C877 a_n2318_13878.t1 gnd 0.117544f
C878 a_n2318_13878.n83 gnd 1.03866f
C879 a_n2318_13878.t4 gnd 0.117544f
C880 a_n2318_13878.t2 gnd 0.117544f
C881 a_n2318_13878.n84 gnd 1.04032f
C882 a_n2318_13878.t7 gnd 0.117544f
C883 a_n2318_13878.t16 gnd 0.117544f
C884 a_n2318_13878.n85 gnd 1.03866f
C885 a_n2318_13878.n86 gnd 0.309588f
C886 a_n2318_13878.n87 gnd 0.30246f
C887 a_n2318_13878.n88 gnd 0.30246f
C888 a_n2318_13878.n89 gnd 0.309588f
C889 a_n2318_13878.t40 gnd 1.41509f
C890 a_n2318_13878.t46 gnd 0.151128f
C891 a_n2318_13878.t28 gnd 0.151128f
C892 a_n2318_13878.n90 gnd 1.06455f
C893 a_n2318_13878.t34 gnd 0.151128f
C894 a_n2318_13878.t26 gnd 0.151128f
C895 a_n2318_13878.n91 gnd 1.06455f
C896 a_n2318_13878.t44 gnd 0.151128f
C897 a_n2318_13878.t22 gnd 0.151128f
C898 a_n2318_13878.n92 gnd 1.06455f
C899 a_n2318_13878.t36 gnd 1.41227f
C900 a_n2318_13878.n93 gnd 0.867362f
C901 a_n2318_13878.t61 gnd 0.702974f
C902 a_n2318_13878.t71 gnd 0.702974f
C903 a_n2318_13878.t83 gnd 0.702974f
C904 a_n2318_13878.n94 gnd 0.309072f
C905 a_n2318_13878.t73 gnd 0.702974f
C906 a_n2318_13878.t58 gnd 0.702974f
C907 a_n2318_13878.t59 gnd 0.702974f
C908 a_n2318_13878.n95 gnd 0.309072f
C909 a_n2318_13878.t77 gnd 0.702974f
C910 a_n2318_13878.t66 gnd 0.702974f
C911 a_n2318_13878.t65 gnd 0.702974f
C912 a_n2318_13878.n96 gnd 0.309072f
C913 a_n2318_13878.t69 gnd 0.702974f
C914 a_n2318_13878.t60 gnd 0.702974f
C915 a_n2318_13878.t52 gnd 0.702974f
C916 a_n2318_13878.n97 gnd 0.309072f
C917 a_n2318_13878.t74 gnd 0.714753f
C918 a_n2318_13878.n98 gnd 0.305147f
C919 a_n2318_13878.n99 gnd 0.299606f
C920 a_n2318_13878.t81 gnd 0.714753f
C921 a_n2318_13878.n100 gnd 0.305147f
C922 a_n2318_13878.n101 gnd 0.299606f
C923 a_n2318_13878.t68 gnd 0.714753f
C924 a_n2318_13878.n102 gnd 0.305147f
C925 a_n2318_13878.n103 gnd 0.299606f
C926 a_n2318_13878.t64 gnd 0.714753f
C927 a_n2318_13878.n104 gnd 0.305147f
C928 a_n2318_13878.n105 gnd 0.299606f
C929 a_n2318_13878.n106 gnd 1.12829f
C930 a_n2318_13878.n107 gnd 0.309588f
C931 a_n2318_13878.t75 gnd 0.702974f
C932 a_n2318_13878.n108 gnd 0.307084f
C933 a_n2318_13878.n109 gnd 0.30246f
C934 a_n2318_13878.t53 gnd 0.702974f
C935 a_n2318_13878.n110 gnd 0.30246f
C936 a_n2318_13878.t70 gnd 0.702974f
C937 a_n2318_13878.n111 gnd 0.309588f
C938 a_n2318_13878.t55 gnd 0.714753f
C939 a_n2318_13878.n112 gnd 0.309588f
C940 a_n2318_13878.t19 gnd 0.702974f
C941 a_n2318_13878.n113 gnd 0.307084f
C942 a_n2318_13878.n114 gnd 0.30246f
C943 a_n2318_13878.t17 gnd 0.702974f
C944 a_n2318_13878.n115 gnd 0.30246f
C945 a_n2318_13878.t41 gnd 0.702974f
C946 a_n2318_13878.n116 gnd 0.309588f
C947 a_n2318_13878.t47 gnd 0.714753f
C948 a_n2318_13878.n117 gnd 1.20932f
C949 a_n2318_13878.t48 gnd 1.41226f
C950 a_n2318_13878.t38 gnd 0.151128f
C951 a_n2318_13878.t42 gnd 0.151128f
C952 a_n2318_13878.n118 gnd 1.06455f
C953 a_n2318_13878.n119 gnd 1.06455f
C954 a_n2318_13878.t18 gnd 0.151128f
C955 vdd.t113 gnd 0.039229f
C956 vdd.t135 gnd 0.039229f
C957 vdd.n0 gnd 0.309405f
C958 vdd.t129 gnd 0.039229f
C959 vdd.t105 gnd 0.039229f
C960 vdd.n1 gnd 0.308894f
C961 vdd.n2 gnd 0.284859f
C962 vdd.t133 gnd 0.039229f
C963 vdd.t119 gnd 0.039229f
C964 vdd.n3 gnd 0.308894f
C965 vdd.n4 gnd 0.144064f
C966 vdd.t121 gnd 0.039229f
C967 vdd.t137 gnd 0.039229f
C968 vdd.n5 gnd 0.308894f
C969 vdd.n6 gnd 0.135177f
C970 vdd.t24 gnd 0.039229f
C971 vdd.t126 gnd 0.039229f
C972 vdd.n7 gnd 0.309405f
C973 vdd.t139 gnd 0.039229f
C974 vdd.t111 gnd 0.039229f
C975 vdd.n8 gnd 0.308894f
C976 vdd.n9 gnd 0.284859f
C977 vdd.t107 gnd 0.039229f
C978 vdd.t116 gnd 0.039229f
C979 vdd.n10 gnd 0.308894f
C980 vdd.n11 gnd 0.144064f
C981 vdd.t131 gnd 0.039229f
C982 vdd.t103 gnd 0.039229f
C983 vdd.n12 gnd 0.308894f
C984 vdd.n13 gnd 0.135177f
C985 vdd.n14 gnd 0.095568f
C986 vdd.t3 gnd 0.021794f
C987 vdd.t4 gnd 0.021794f
C988 vdd.n15 gnd 0.200603f
C989 vdd.t16 gnd 0.021794f
C990 vdd.t5 gnd 0.021794f
C991 vdd.n16 gnd 0.200016f
C992 vdd.n17 gnd 0.34809f
C993 vdd.t15 gnd 0.021794f
C994 vdd.t9 gnd 0.021794f
C995 vdd.n18 gnd 0.200016f
C996 vdd.n19 gnd 0.14401f
C997 vdd.t7 gnd 0.021794f
C998 vdd.t10 gnd 0.021794f
C999 vdd.n20 gnd 0.200603f
C1000 vdd.t8 gnd 0.021794f
C1001 vdd.t12 gnd 0.021794f
C1002 vdd.n21 gnd 0.200016f
C1003 vdd.n22 gnd 0.34809f
C1004 vdd.t6 gnd 0.021794f
C1005 vdd.t2 gnd 0.021794f
C1006 vdd.n23 gnd 0.200016f
C1007 vdd.n24 gnd 0.14401f
C1008 vdd.t14 gnd 0.021794f
C1009 vdd.t17 gnd 0.021794f
C1010 vdd.n25 gnd 0.200016f
C1011 vdd.t13 gnd 0.021794f
C1012 vdd.t11 gnd 0.021794f
C1013 vdd.n26 gnd 0.200016f
C1014 vdd.n27 gnd 23.282999f
C1015 vdd.n28 gnd 8.88987f
C1016 vdd.n29 gnd 0.005944f
C1017 vdd.n30 gnd 0.005516f
C1018 vdd.n31 gnd 0.003051f
C1019 vdd.n32 gnd 0.007006f
C1020 vdd.n33 gnd 0.002964f
C1021 vdd.n34 gnd 0.003138f
C1022 vdd.n35 gnd 0.005516f
C1023 vdd.n36 gnd 0.002964f
C1024 vdd.n37 gnd 0.007006f
C1025 vdd.n38 gnd 0.003138f
C1026 vdd.n39 gnd 0.005516f
C1027 vdd.n40 gnd 0.002964f
C1028 vdd.n41 gnd 0.005254f
C1029 vdd.n42 gnd 0.00527f
C1030 vdd.t187 gnd 0.015051f
C1031 vdd.n43 gnd 0.033489f
C1032 vdd.n44 gnd 0.174283f
C1033 vdd.n45 gnd 0.002964f
C1034 vdd.n46 gnd 0.003138f
C1035 vdd.n47 gnd 0.007006f
C1036 vdd.n48 gnd 0.007006f
C1037 vdd.n49 gnd 0.003138f
C1038 vdd.n50 gnd 0.002964f
C1039 vdd.n51 gnd 0.005516f
C1040 vdd.n52 gnd 0.005516f
C1041 vdd.n53 gnd 0.002964f
C1042 vdd.n54 gnd 0.003138f
C1043 vdd.n55 gnd 0.007006f
C1044 vdd.n56 gnd 0.007006f
C1045 vdd.n57 gnd 0.003138f
C1046 vdd.n58 gnd 0.002964f
C1047 vdd.n59 gnd 0.005516f
C1048 vdd.n60 gnd 0.005516f
C1049 vdd.n61 gnd 0.002964f
C1050 vdd.n62 gnd 0.003138f
C1051 vdd.n63 gnd 0.007006f
C1052 vdd.n64 gnd 0.007006f
C1053 vdd.n65 gnd 0.016563f
C1054 vdd.n66 gnd 0.003051f
C1055 vdd.n67 gnd 0.002964f
C1056 vdd.n68 gnd 0.014257f
C1057 vdd.n69 gnd 0.009953f
C1058 vdd.t277 gnd 0.03487f
C1059 vdd.t219 gnd 0.03487f
C1060 vdd.n70 gnd 0.239652f
C1061 vdd.n71 gnd 0.188449f
C1062 vdd.t291 gnd 0.03487f
C1063 vdd.t271 gnd 0.03487f
C1064 vdd.n72 gnd 0.239652f
C1065 vdd.n73 gnd 0.152078f
C1066 vdd.t153 gnd 0.03487f
C1067 vdd.t206 gnd 0.03487f
C1068 vdd.n74 gnd 0.239652f
C1069 vdd.n75 gnd 0.152078f
C1070 vdd.t165 gnd 0.03487f
C1071 vdd.t232 gnd 0.03487f
C1072 vdd.n76 gnd 0.239652f
C1073 vdd.n77 gnd 0.152078f
C1074 vdd.t195 gnd 0.03487f
C1075 vdd.t281 gnd 0.03487f
C1076 vdd.n78 gnd 0.239652f
C1077 vdd.n79 gnd 0.152078f
C1078 vdd.t171 gnd 0.03487f
C1079 vdd.t254 gnd 0.03487f
C1080 vdd.n80 gnd 0.239652f
C1081 vdd.n81 gnd 0.152078f
C1082 vdd.t177 gnd 0.03487f
C1083 vdd.t273 gnd 0.03487f
C1084 vdd.n82 gnd 0.239652f
C1085 vdd.n83 gnd 0.152078f
C1086 vdd.t214 gnd 0.03487f
C1087 vdd.t286 gnd 0.03487f
C1088 vdd.n84 gnd 0.239652f
C1089 vdd.n85 gnd 0.152078f
C1090 vdd.t235 gnd 0.03487f
C1091 vdd.t264 gnd 0.03487f
C1092 vdd.n86 gnd 0.239652f
C1093 vdd.n87 gnd 0.152078f
C1094 vdd.n88 gnd 0.005944f
C1095 vdd.n89 gnd 0.005516f
C1096 vdd.n90 gnd 0.003051f
C1097 vdd.n91 gnd 0.007006f
C1098 vdd.n92 gnd 0.002964f
C1099 vdd.n93 gnd 0.003138f
C1100 vdd.n94 gnd 0.005516f
C1101 vdd.n95 gnd 0.002964f
C1102 vdd.n96 gnd 0.007006f
C1103 vdd.n97 gnd 0.003138f
C1104 vdd.n98 gnd 0.005516f
C1105 vdd.n99 gnd 0.002964f
C1106 vdd.n100 gnd 0.005254f
C1107 vdd.n101 gnd 0.00527f
C1108 vdd.t198 gnd 0.015051f
C1109 vdd.n102 gnd 0.033489f
C1110 vdd.n103 gnd 0.174283f
C1111 vdd.n104 gnd 0.002964f
C1112 vdd.n105 gnd 0.003138f
C1113 vdd.n106 gnd 0.007006f
C1114 vdd.n107 gnd 0.007006f
C1115 vdd.n108 gnd 0.003138f
C1116 vdd.n109 gnd 0.002964f
C1117 vdd.n110 gnd 0.005516f
C1118 vdd.n111 gnd 0.005516f
C1119 vdd.n112 gnd 0.002964f
C1120 vdd.n113 gnd 0.003138f
C1121 vdd.n114 gnd 0.007006f
C1122 vdd.n115 gnd 0.007006f
C1123 vdd.n116 gnd 0.003138f
C1124 vdd.n117 gnd 0.002964f
C1125 vdd.n118 gnd 0.005516f
C1126 vdd.n119 gnd 0.005516f
C1127 vdd.n120 gnd 0.002964f
C1128 vdd.n121 gnd 0.003138f
C1129 vdd.n122 gnd 0.007006f
C1130 vdd.n123 gnd 0.007006f
C1131 vdd.n124 gnd 0.016563f
C1132 vdd.n125 gnd 0.003051f
C1133 vdd.n126 gnd 0.002964f
C1134 vdd.n127 gnd 0.014257f
C1135 vdd.n128 gnd 0.009641f
C1136 vdd.n129 gnd 0.113146f
C1137 vdd.n130 gnd 0.005944f
C1138 vdd.n131 gnd 0.005516f
C1139 vdd.n132 gnd 0.003051f
C1140 vdd.n133 gnd 0.007006f
C1141 vdd.n134 gnd 0.002964f
C1142 vdd.n135 gnd 0.003138f
C1143 vdd.n136 gnd 0.005516f
C1144 vdd.n137 gnd 0.002964f
C1145 vdd.n138 gnd 0.007006f
C1146 vdd.n139 gnd 0.003138f
C1147 vdd.n140 gnd 0.005516f
C1148 vdd.n141 gnd 0.002964f
C1149 vdd.n142 gnd 0.005254f
C1150 vdd.n143 gnd 0.00527f
C1151 vdd.t230 gnd 0.015051f
C1152 vdd.n144 gnd 0.033489f
C1153 vdd.n145 gnd 0.174283f
C1154 vdd.n146 gnd 0.002964f
C1155 vdd.n147 gnd 0.003138f
C1156 vdd.n148 gnd 0.007006f
C1157 vdd.n149 gnd 0.007006f
C1158 vdd.n150 gnd 0.003138f
C1159 vdd.n151 gnd 0.002964f
C1160 vdd.n152 gnd 0.005516f
C1161 vdd.n153 gnd 0.005516f
C1162 vdd.n154 gnd 0.002964f
C1163 vdd.n155 gnd 0.003138f
C1164 vdd.n156 gnd 0.007006f
C1165 vdd.n157 gnd 0.007006f
C1166 vdd.n158 gnd 0.003138f
C1167 vdd.n159 gnd 0.002964f
C1168 vdd.n160 gnd 0.005516f
C1169 vdd.n161 gnd 0.005516f
C1170 vdd.n162 gnd 0.002964f
C1171 vdd.n163 gnd 0.003138f
C1172 vdd.n164 gnd 0.007006f
C1173 vdd.n165 gnd 0.007006f
C1174 vdd.n166 gnd 0.016563f
C1175 vdd.n167 gnd 0.003051f
C1176 vdd.n168 gnd 0.002964f
C1177 vdd.n169 gnd 0.014257f
C1178 vdd.n170 gnd 0.009953f
C1179 vdd.t263 gnd 0.03487f
C1180 vdd.t143 gnd 0.03487f
C1181 vdd.n171 gnd 0.239652f
C1182 vdd.n172 gnd 0.188449f
C1183 vdd.t203 gnd 0.03487f
C1184 vdd.t205 gnd 0.03487f
C1185 vdd.n173 gnd 0.239652f
C1186 vdd.n174 gnd 0.152078f
C1187 vdd.t285 gnd 0.03487f
C1188 vdd.t192 gnd 0.03487f
C1189 vdd.n175 gnd 0.239652f
C1190 vdd.n176 gnd 0.152078f
C1191 vdd.t193 gnd 0.03487f
C1192 vdd.t283 gnd 0.03487f
C1193 vdd.n177 gnd 0.239652f
C1194 vdd.n178 gnd 0.152078f
C1195 vdd.t284 gnd 0.03487f
C1196 vdd.t163 gnd 0.03487f
C1197 vdd.n179 gnd 0.239652f
C1198 vdd.n180 gnd 0.152078f
C1199 vdd.t266 gnd 0.03487f
C1200 vdd.t280 gnd 0.03487f
C1201 vdd.n181 gnd 0.239652f
C1202 vdd.n182 gnd 0.152078f
C1203 vdd.t159 gnd 0.03487f
C1204 vdd.t229 gnd 0.03487f
C1205 vdd.n183 gnd 0.239652f
C1206 vdd.n184 gnd 0.152078f
C1207 vdd.t261 gnd 0.03487f
C1208 vdd.t292 gnd 0.03487f
C1209 vdd.n185 gnd 0.239652f
C1210 vdd.n186 gnd 0.152078f
C1211 vdd.t201 gnd 0.03487f
C1212 vdd.t260 gnd 0.03487f
C1213 vdd.n187 gnd 0.239652f
C1214 vdd.n188 gnd 0.152078f
C1215 vdd.n189 gnd 0.005944f
C1216 vdd.n190 gnd 0.005516f
C1217 vdd.n191 gnd 0.003051f
C1218 vdd.n192 gnd 0.007006f
C1219 vdd.n193 gnd 0.002964f
C1220 vdd.n194 gnd 0.003138f
C1221 vdd.n195 gnd 0.005516f
C1222 vdd.n196 gnd 0.002964f
C1223 vdd.n197 gnd 0.007006f
C1224 vdd.n198 gnd 0.003138f
C1225 vdd.n199 gnd 0.005516f
C1226 vdd.n200 gnd 0.002964f
C1227 vdd.n201 gnd 0.005254f
C1228 vdd.n202 gnd 0.00527f
C1229 vdd.t297 gnd 0.015051f
C1230 vdd.n203 gnd 0.033489f
C1231 vdd.n204 gnd 0.174283f
C1232 vdd.n205 gnd 0.002964f
C1233 vdd.n206 gnd 0.003138f
C1234 vdd.n207 gnd 0.007006f
C1235 vdd.n208 gnd 0.007006f
C1236 vdd.n209 gnd 0.003138f
C1237 vdd.n210 gnd 0.002964f
C1238 vdd.n211 gnd 0.005516f
C1239 vdd.n212 gnd 0.005516f
C1240 vdd.n213 gnd 0.002964f
C1241 vdd.n214 gnd 0.003138f
C1242 vdd.n215 gnd 0.007006f
C1243 vdd.n216 gnd 0.007006f
C1244 vdd.n217 gnd 0.003138f
C1245 vdd.n218 gnd 0.002964f
C1246 vdd.n219 gnd 0.005516f
C1247 vdd.n220 gnd 0.005516f
C1248 vdd.n221 gnd 0.002964f
C1249 vdd.n222 gnd 0.003138f
C1250 vdd.n223 gnd 0.007006f
C1251 vdd.n224 gnd 0.007006f
C1252 vdd.n225 gnd 0.016563f
C1253 vdd.n226 gnd 0.003051f
C1254 vdd.n227 gnd 0.002964f
C1255 vdd.n228 gnd 0.014257f
C1256 vdd.n229 gnd 0.009641f
C1257 vdd.n230 gnd 0.067311f
C1258 vdd.n231 gnd 0.242538f
C1259 vdd.n232 gnd 0.005944f
C1260 vdd.n233 gnd 0.005516f
C1261 vdd.n234 gnd 0.003051f
C1262 vdd.n235 gnd 0.007006f
C1263 vdd.n236 gnd 0.002964f
C1264 vdd.n237 gnd 0.003138f
C1265 vdd.n238 gnd 0.005516f
C1266 vdd.n239 gnd 0.002964f
C1267 vdd.n240 gnd 0.007006f
C1268 vdd.n241 gnd 0.003138f
C1269 vdd.n242 gnd 0.005516f
C1270 vdd.n243 gnd 0.002964f
C1271 vdd.n244 gnd 0.005254f
C1272 vdd.n245 gnd 0.00527f
C1273 vdd.t246 gnd 0.015051f
C1274 vdd.n246 gnd 0.033489f
C1275 vdd.n247 gnd 0.174283f
C1276 vdd.n248 gnd 0.002964f
C1277 vdd.n249 gnd 0.003138f
C1278 vdd.n250 gnd 0.007006f
C1279 vdd.n251 gnd 0.007006f
C1280 vdd.n252 gnd 0.003138f
C1281 vdd.n253 gnd 0.002964f
C1282 vdd.n254 gnd 0.005516f
C1283 vdd.n255 gnd 0.005516f
C1284 vdd.n256 gnd 0.002964f
C1285 vdd.n257 gnd 0.003138f
C1286 vdd.n258 gnd 0.007006f
C1287 vdd.n259 gnd 0.007006f
C1288 vdd.n260 gnd 0.003138f
C1289 vdd.n261 gnd 0.002964f
C1290 vdd.n262 gnd 0.005516f
C1291 vdd.n263 gnd 0.005516f
C1292 vdd.n264 gnd 0.002964f
C1293 vdd.n265 gnd 0.003138f
C1294 vdd.n266 gnd 0.007006f
C1295 vdd.n267 gnd 0.007006f
C1296 vdd.n268 gnd 0.016563f
C1297 vdd.n269 gnd 0.003051f
C1298 vdd.n270 gnd 0.002964f
C1299 vdd.n271 gnd 0.014257f
C1300 vdd.n272 gnd 0.009953f
C1301 vdd.t274 gnd 0.03487f
C1302 vdd.t169 gnd 0.03487f
C1303 vdd.n273 gnd 0.239652f
C1304 vdd.n274 gnd 0.188449f
C1305 vdd.t223 gnd 0.03487f
C1306 vdd.t226 gnd 0.03487f
C1307 vdd.n275 gnd 0.239652f
C1308 vdd.n276 gnd 0.152078f
C1309 vdd.t296 gnd 0.03487f
C1310 vdd.t217 gnd 0.03487f
C1311 vdd.n277 gnd 0.239652f
C1312 vdd.n278 gnd 0.152078f
C1313 vdd.t218 gnd 0.03487f
C1314 vdd.t294 gnd 0.03487f
C1315 vdd.n279 gnd 0.239652f
C1316 vdd.n280 gnd 0.152078f
C1317 vdd.t295 gnd 0.03487f
C1318 vdd.t185 gnd 0.03487f
C1319 vdd.n281 gnd 0.239652f
C1320 vdd.n282 gnd 0.152078f
C1321 vdd.t279 gnd 0.03487f
C1322 vdd.t290 gnd 0.03487f
C1323 vdd.n283 gnd 0.239652f
C1324 vdd.n284 gnd 0.152078f
C1325 vdd.t178 gnd 0.03487f
C1326 vdd.t247 gnd 0.03487f
C1327 vdd.n285 gnd 0.239652f
C1328 vdd.n286 gnd 0.152078f
C1329 vdd.t275 gnd 0.03487f
C1330 vdd.t147 gnd 0.03487f
C1331 vdd.n287 gnd 0.239652f
C1332 vdd.n288 gnd 0.152078f
C1333 vdd.t224 gnd 0.03487f
C1334 vdd.t272 gnd 0.03487f
C1335 vdd.n289 gnd 0.239652f
C1336 vdd.n290 gnd 0.152078f
C1337 vdd.n291 gnd 0.005944f
C1338 vdd.n292 gnd 0.005516f
C1339 vdd.n293 gnd 0.003051f
C1340 vdd.n294 gnd 0.007006f
C1341 vdd.n295 gnd 0.002964f
C1342 vdd.n296 gnd 0.003138f
C1343 vdd.n297 gnd 0.005516f
C1344 vdd.n298 gnd 0.002964f
C1345 vdd.n299 gnd 0.007006f
C1346 vdd.n300 gnd 0.003138f
C1347 vdd.n301 gnd 0.005516f
C1348 vdd.n302 gnd 0.002964f
C1349 vdd.n303 gnd 0.005254f
C1350 vdd.n304 gnd 0.00527f
C1351 vdd.t161 gnd 0.015051f
C1352 vdd.n305 gnd 0.033489f
C1353 vdd.n306 gnd 0.174283f
C1354 vdd.n307 gnd 0.002964f
C1355 vdd.n308 gnd 0.003138f
C1356 vdd.n309 gnd 0.007006f
C1357 vdd.n310 gnd 0.007006f
C1358 vdd.n311 gnd 0.003138f
C1359 vdd.n312 gnd 0.002964f
C1360 vdd.n313 gnd 0.005516f
C1361 vdd.n314 gnd 0.005516f
C1362 vdd.n315 gnd 0.002964f
C1363 vdd.n316 gnd 0.003138f
C1364 vdd.n317 gnd 0.007006f
C1365 vdd.n318 gnd 0.007006f
C1366 vdd.n319 gnd 0.003138f
C1367 vdd.n320 gnd 0.002964f
C1368 vdd.n321 gnd 0.005516f
C1369 vdd.n322 gnd 0.005516f
C1370 vdd.n323 gnd 0.002964f
C1371 vdd.n324 gnd 0.003138f
C1372 vdd.n325 gnd 0.007006f
C1373 vdd.n326 gnd 0.007006f
C1374 vdd.n327 gnd 0.016563f
C1375 vdd.n328 gnd 0.003051f
C1376 vdd.n329 gnd 0.002964f
C1377 vdd.n330 gnd 0.014257f
C1378 vdd.n331 gnd 0.009641f
C1379 vdd.n332 gnd 0.067311f
C1380 vdd.n333 gnd 0.277654f
C1381 vdd.n334 gnd 0.008324f
C1382 vdd.n335 gnd 0.010831f
C1383 vdd.n336 gnd 0.008718f
C1384 vdd.n337 gnd 0.008718f
C1385 vdd.n338 gnd 0.010831f
C1386 vdd.n339 gnd 0.010831f
C1387 vdd.n340 gnd 0.791407f
C1388 vdd.n341 gnd 0.010831f
C1389 vdd.n342 gnd 0.010831f
C1390 vdd.n343 gnd 0.010831f
C1391 vdd.n344 gnd 0.857819f
C1392 vdd.n345 gnd 0.010831f
C1393 vdd.n346 gnd 0.010831f
C1394 vdd.n347 gnd 0.010831f
C1395 vdd.n348 gnd 0.010831f
C1396 vdd.n349 gnd 0.008718f
C1397 vdd.n350 gnd 0.010831f
C1398 vdd.t253 gnd 0.553432f
C1399 vdd.n351 gnd 0.010831f
C1400 vdd.n352 gnd 0.010831f
C1401 vdd.n353 gnd 0.010831f
C1402 vdd.t228 gnd 0.553432f
C1403 vdd.n354 gnd 0.010831f
C1404 vdd.n355 gnd 0.010831f
C1405 vdd.n356 gnd 0.010831f
C1406 vdd.n357 gnd 0.010831f
C1407 vdd.n358 gnd 0.010831f
C1408 vdd.n359 gnd 0.008718f
C1409 vdd.n360 gnd 0.010831f
C1410 vdd.n361 gnd 0.625378f
C1411 vdd.n362 gnd 0.010831f
C1412 vdd.n363 gnd 0.010831f
C1413 vdd.n364 gnd 0.010831f
C1414 vdd.t146 gnd 0.553432f
C1415 vdd.n365 gnd 0.010831f
C1416 vdd.n366 gnd 0.010831f
C1417 vdd.n367 gnd 0.010831f
C1418 vdd.n368 gnd 0.010831f
C1419 vdd.n369 gnd 0.010831f
C1420 vdd.n370 gnd 0.008718f
C1421 vdd.n371 gnd 0.010831f
C1422 vdd.t200 gnd 0.553432f
C1423 vdd.n372 gnd 0.010831f
C1424 vdd.n373 gnd 0.010831f
C1425 vdd.n374 gnd 0.010831f
C1426 vdd.n375 gnd 0.647515f
C1427 vdd.n376 gnd 0.010831f
C1428 vdd.n377 gnd 0.010831f
C1429 vdd.n378 gnd 0.010831f
C1430 vdd.n379 gnd 0.010831f
C1431 vdd.n380 gnd 0.010831f
C1432 vdd.n381 gnd 0.008718f
C1433 vdd.n382 gnd 0.010831f
C1434 vdd.t160 gnd 0.553432f
C1435 vdd.n383 gnd 0.010831f
C1436 vdd.n384 gnd 0.010831f
C1437 vdd.n385 gnd 0.010831f
C1438 vdd.n386 gnd 0.558966f
C1439 vdd.n387 gnd 0.010831f
C1440 vdd.n388 gnd 0.010831f
C1441 vdd.n389 gnd 0.010831f
C1442 vdd.n390 gnd 0.010831f
C1443 vdd.n391 gnd 0.026201f
C1444 vdd.n392 gnd 0.026762f
C1445 vdd.t49 gnd 0.553432f
C1446 vdd.n393 gnd 0.026201f
C1447 vdd.n425 gnd 0.010831f
C1448 vdd.t61 gnd 0.133248f
C1449 vdd.t60 gnd 0.142406f
C1450 vdd.t59 gnd 0.17402f
C1451 vdd.n426 gnd 0.223069f
C1452 vdd.n427 gnd 0.18829f
C1453 vdd.n428 gnd 0.014297f
C1454 vdd.n429 gnd 0.010831f
C1455 vdd.n430 gnd 0.008718f
C1456 vdd.n431 gnd 0.010831f
C1457 vdd.n432 gnd 0.008718f
C1458 vdd.n433 gnd 0.010831f
C1459 vdd.n434 gnd 0.008718f
C1460 vdd.n435 gnd 0.010831f
C1461 vdd.n436 gnd 0.008718f
C1462 vdd.n437 gnd 0.010831f
C1463 vdd.n438 gnd 0.008718f
C1464 vdd.n439 gnd 0.010831f
C1465 vdd.t51 gnd 0.133248f
C1466 vdd.t50 gnd 0.142406f
C1467 vdd.t48 gnd 0.17402f
C1468 vdd.n440 gnd 0.223069f
C1469 vdd.n441 gnd 0.18829f
C1470 vdd.n442 gnd 0.008718f
C1471 vdd.n443 gnd 0.010831f
C1472 vdd.n444 gnd 0.008718f
C1473 vdd.n445 gnd 0.010831f
C1474 vdd.n446 gnd 0.008718f
C1475 vdd.n447 gnd 0.010831f
C1476 vdd.n448 gnd 0.008718f
C1477 vdd.n449 gnd 0.010831f
C1478 vdd.n450 gnd 0.008718f
C1479 vdd.n451 gnd 0.010831f
C1480 vdd.t68 gnd 0.133248f
C1481 vdd.t67 gnd 0.142406f
C1482 vdd.t66 gnd 0.17402f
C1483 vdd.n452 gnd 0.223069f
C1484 vdd.n453 gnd 0.18829f
C1485 vdd.n454 gnd 0.018655f
C1486 vdd.n455 gnd 0.010831f
C1487 vdd.n456 gnd 0.008718f
C1488 vdd.n457 gnd 0.010831f
C1489 vdd.n458 gnd 0.008718f
C1490 vdd.n459 gnd 0.010831f
C1491 vdd.n460 gnd 0.008718f
C1492 vdd.n461 gnd 0.010831f
C1493 vdd.n462 gnd 0.008718f
C1494 vdd.n463 gnd 0.010831f
C1495 vdd.n464 gnd 0.026762f
C1496 vdd.n465 gnd 0.007236f
C1497 vdd.n466 gnd 0.008718f
C1498 vdd.n467 gnd 0.010831f
C1499 vdd.n468 gnd 0.010831f
C1500 vdd.n469 gnd 0.008718f
C1501 vdd.n470 gnd 0.010831f
C1502 vdd.n471 gnd 0.010831f
C1503 vdd.n472 gnd 0.010831f
C1504 vdd.n473 gnd 0.010831f
C1505 vdd.n474 gnd 0.010831f
C1506 vdd.n475 gnd 0.008718f
C1507 vdd.n476 gnd 0.008718f
C1508 vdd.n477 gnd 0.010831f
C1509 vdd.n478 gnd 0.010831f
C1510 vdd.n479 gnd 0.008718f
C1511 vdd.n480 gnd 0.010831f
C1512 vdd.n481 gnd 0.010831f
C1513 vdd.n482 gnd 0.010831f
C1514 vdd.n483 gnd 0.010831f
C1515 vdd.n484 gnd 0.010831f
C1516 vdd.n485 gnd 0.008718f
C1517 vdd.n486 gnd 0.008718f
C1518 vdd.n487 gnd 0.010831f
C1519 vdd.n488 gnd 0.010831f
C1520 vdd.n489 gnd 0.008718f
C1521 vdd.n490 gnd 0.010831f
C1522 vdd.n491 gnd 0.010831f
C1523 vdd.n492 gnd 0.010831f
C1524 vdd.n493 gnd 0.010831f
C1525 vdd.n494 gnd 0.010831f
C1526 vdd.n495 gnd 0.008718f
C1527 vdd.n496 gnd 0.008718f
C1528 vdd.n497 gnd 0.010831f
C1529 vdd.n498 gnd 0.010831f
C1530 vdd.n499 gnd 0.008718f
C1531 vdd.n500 gnd 0.010831f
C1532 vdd.n501 gnd 0.010831f
C1533 vdd.n502 gnd 0.010831f
C1534 vdd.n503 gnd 0.010831f
C1535 vdd.n504 gnd 0.010831f
C1536 vdd.n505 gnd 0.008718f
C1537 vdd.n506 gnd 0.008718f
C1538 vdd.n507 gnd 0.010831f
C1539 vdd.n508 gnd 0.010831f
C1540 vdd.n509 gnd 0.007279f
C1541 vdd.n510 gnd 0.010831f
C1542 vdd.n511 gnd 0.010831f
C1543 vdd.n512 gnd 0.010831f
C1544 vdd.n513 gnd 0.010831f
C1545 vdd.n514 gnd 0.010831f
C1546 vdd.n515 gnd 0.007279f
C1547 vdd.n516 gnd 0.008718f
C1548 vdd.n517 gnd 0.010831f
C1549 vdd.n518 gnd 0.010831f
C1550 vdd.n519 gnd 0.008718f
C1551 vdd.n520 gnd 0.010831f
C1552 vdd.n521 gnd 0.010831f
C1553 vdd.n522 gnd 0.010831f
C1554 vdd.n523 gnd 0.010831f
C1555 vdd.n524 gnd 0.010831f
C1556 vdd.n525 gnd 0.008718f
C1557 vdd.n526 gnd 0.008718f
C1558 vdd.n527 gnd 0.010831f
C1559 vdd.n528 gnd 0.010831f
C1560 vdd.n529 gnd 0.008718f
C1561 vdd.n530 gnd 0.010831f
C1562 vdd.n531 gnd 0.010831f
C1563 vdd.n532 gnd 0.010831f
C1564 vdd.n533 gnd 0.010831f
C1565 vdd.n534 gnd 0.010831f
C1566 vdd.n535 gnd 0.008718f
C1567 vdd.n536 gnd 0.008718f
C1568 vdd.n537 gnd 0.010831f
C1569 vdd.n538 gnd 0.010831f
C1570 vdd.n539 gnd 0.008718f
C1571 vdd.n540 gnd 0.010831f
C1572 vdd.n541 gnd 0.010831f
C1573 vdd.n542 gnd 0.010831f
C1574 vdd.n543 gnd 0.010831f
C1575 vdd.n544 gnd 0.010831f
C1576 vdd.n545 gnd 0.008718f
C1577 vdd.n546 gnd 0.008718f
C1578 vdd.n547 gnd 0.010831f
C1579 vdd.n548 gnd 0.010831f
C1580 vdd.n549 gnd 0.008718f
C1581 vdd.n550 gnd 0.010831f
C1582 vdd.n551 gnd 0.010831f
C1583 vdd.n552 gnd 0.010831f
C1584 vdd.n553 gnd 0.010831f
C1585 vdd.n554 gnd 0.010831f
C1586 vdd.n555 gnd 0.008718f
C1587 vdd.n556 gnd 0.008718f
C1588 vdd.n557 gnd 0.010831f
C1589 vdd.n558 gnd 0.010831f
C1590 vdd.n559 gnd 0.008718f
C1591 vdd.n560 gnd 0.010831f
C1592 vdd.n561 gnd 0.010831f
C1593 vdd.n562 gnd 0.010831f
C1594 vdd.n563 gnd 0.010831f
C1595 vdd.n564 gnd 0.010831f
C1596 vdd.n565 gnd 0.005928f
C1597 vdd.n566 gnd 0.018655f
C1598 vdd.n567 gnd 0.010831f
C1599 vdd.n568 gnd 0.010831f
C1600 vdd.n569 gnd 0.00863f
C1601 vdd.n570 gnd 0.010831f
C1602 vdd.n571 gnd 0.010831f
C1603 vdd.n572 gnd 0.010831f
C1604 vdd.n573 gnd 0.010831f
C1605 vdd.n574 gnd 0.010831f
C1606 vdd.n575 gnd 0.008718f
C1607 vdd.n576 gnd 0.008718f
C1608 vdd.n577 gnd 0.010831f
C1609 vdd.n578 gnd 0.010831f
C1610 vdd.n579 gnd 0.008718f
C1611 vdd.n580 gnd 0.010831f
C1612 vdd.n581 gnd 0.010831f
C1613 vdd.n582 gnd 0.010831f
C1614 vdd.n583 gnd 0.010831f
C1615 vdd.n584 gnd 0.010831f
C1616 vdd.n585 gnd 0.008718f
C1617 vdd.n586 gnd 0.008718f
C1618 vdd.n587 gnd 0.010831f
C1619 vdd.n588 gnd 0.010831f
C1620 vdd.n589 gnd 0.008718f
C1621 vdd.n590 gnd 0.010831f
C1622 vdd.n591 gnd 0.010831f
C1623 vdd.n592 gnd 0.010831f
C1624 vdd.n593 gnd 0.010831f
C1625 vdd.n594 gnd 0.010831f
C1626 vdd.n595 gnd 0.008718f
C1627 vdd.n596 gnd 0.008718f
C1628 vdd.n597 gnd 0.010831f
C1629 vdd.n598 gnd 0.010831f
C1630 vdd.n599 gnd 0.008718f
C1631 vdd.n600 gnd 0.010831f
C1632 vdd.n601 gnd 0.010831f
C1633 vdd.n602 gnd 0.010831f
C1634 vdd.n603 gnd 0.010831f
C1635 vdd.n604 gnd 0.010831f
C1636 vdd.n605 gnd 0.008718f
C1637 vdd.n606 gnd 0.008718f
C1638 vdd.n607 gnd 0.010831f
C1639 vdd.n608 gnd 0.010831f
C1640 vdd.n609 gnd 0.008718f
C1641 vdd.n610 gnd 0.010831f
C1642 vdd.n611 gnd 0.010831f
C1643 vdd.n612 gnd 0.010831f
C1644 vdd.n613 gnd 0.010831f
C1645 vdd.n614 gnd 0.010831f
C1646 vdd.n615 gnd 0.008718f
C1647 vdd.n616 gnd 0.010831f
C1648 vdd.n617 gnd 0.008718f
C1649 vdd.n618 gnd 0.004577f
C1650 vdd.n619 gnd 0.010831f
C1651 vdd.n620 gnd 0.010831f
C1652 vdd.n621 gnd 0.008718f
C1653 vdd.n622 gnd 0.010831f
C1654 vdd.n623 gnd 0.008718f
C1655 vdd.n624 gnd 0.010831f
C1656 vdd.n625 gnd 0.008718f
C1657 vdd.n626 gnd 0.010831f
C1658 vdd.n627 gnd 0.008718f
C1659 vdd.n628 gnd 0.010831f
C1660 vdd.n629 gnd 0.008718f
C1661 vdd.n630 gnd 0.010831f
C1662 vdd.n631 gnd 0.008718f
C1663 vdd.n632 gnd 0.010831f
C1664 vdd.n633 gnd 0.60324f
C1665 vdd.t194 gnd 0.553432f
C1666 vdd.n634 gnd 0.010831f
C1667 vdd.n635 gnd 0.008718f
C1668 vdd.n636 gnd 0.010831f
C1669 vdd.n637 gnd 0.008718f
C1670 vdd.n638 gnd 0.010831f
C1671 vdd.t164 gnd 0.553432f
C1672 vdd.n639 gnd 0.010831f
C1673 vdd.n640 gnd 0.008718f
C1674 vdd.n641 gnd 0.010831f
C1675 vdd.n642 gnd 0.008718f
C1676 vdd.n643 gnd 0.010831f
C1677 vdd.t191 gnd 0.553432f
C1678 vdd.n644 gnd 0.691789f
C1679 vdd.n645 gnd 0.010831f
C1680 vdd.n646 gnd 0.008718f
C1681 vdd.n647 gnd 0.010831f
C1682 vdd.n648 gnd 0.008718f
C1683 vdd.n649 gnd 0.010831f
C1684 vdd.t152 gnd 0.553432f
C1685 vdd.n650 gnd 0.010831f
C1686 vdd.n651 gnd 0.008718f
C1687 vdd.n652 gnd 0.010831f
C1688 vdd.n653 gnd 0.008718f
C1689 vdd.n654 gnd 0.010831f
C1690 vdd.n655 gnd 0.76927f
C1691 vdd.n656 gnd 0.918696f
C1692 vdd.t204 gnd 0.553432f
C1693 vdd.n657 gnd 0.010831f
C1694 vdd.n658 gnd 0.008718f
C1695 vdd.n659 gnd 0.010831f
C1696 vdd.n660 gnd 0.008718f
C1697 vdd.n661 gnd 0.010831f
C1698 vdd.n662 gnd 0.581103f
C1699 vdd.n663 gnd 0.010831f
C1700 vdd.n664 gnd 0.008718f
C1701 vdd.n665 gnd 0.010831f
C1702 vdd.n666 gnd 0.008718f
C1703 vdd.n667 gnd 0.010831f
C1704 vdd.t262 gnd 0.553432f
C1705 vdd.t142 gnd 0.553432f
C1706 vdd.n668 gnd 0.010831f
C1707 vdd.n669 gnd 0.008718f
C1708 vdd.n670 gnd 0.010831f
C1709 vdd.n671 gnd 0.008718f
C1710 vdd.n672 gnd 0.010831f
C1711 vdd.t186 gnd 0.553432f
C1712 vdd.n673 gnd 0.010831f
C1713 vdd.n674 gnd 0.008718f
C1714 vdd.n675 gnd 0.010831f
C1715 vdd.n676 gnd 0.008718f
C1716 vdd.n677 gnd 0.010831f
C1717 vdd.n678 gnd 1.10686f
C1718 vdd.n679 gnd 0.902093f
C1719 vdd.n680 gnd 0.010831f
C1720 vdd.n681 gnd 0.008718f
C1721 vdd.n682 gnd 0.026201f
C1722 vdd.n683 gnd 0.007236f
C1723 vdd.n684 gnd 0.026201f
C1724 vdd.t35 gnd 0.553432f
C1725 vdd.n685 gnd 0.026201f
C1726 vdd.n686 gnd 0.007236f
C1727 vdd.n687 gnd 0.009315f
C1728 vdd.t36 gnd 0.133248f
C1729 vdd.t37 gnd 0.142406f
C1730 vdd.t34 gnd 0.17402f
C1731 vdd.n688 gnd 0.223069f
C1732 vdd.n689 gnd 0.187419f
C1733 vdd.n690 gnd 0.013425f
C1734 vdd.n691 gnd 0.010831f
C1735 vdd.n692 gnd 9.44154f
C1736 vdd.n723 gnd 1.52194f
C1737 vdd.n724 gnd 0.010831f
C1738 vdd.n725 gnd 0.010831f
C1739 vdd.n726 gnd 0.026762f
C1740 vdd.n727 gnd 0.009315f
C1741 vdd.n728 gnd 0.010831f
C1742 vdd.n729 gnd 0.008718f
C1743 vdd.n730 gnd 0.006932f
C1744 vdd.n731 gnd 0.025294f
C1745 vdd.n732 gnd 0.008718f
C1746 vdd.n733 gnd 0.010831f
C1747 vdd.n734 gnd 0.010831f
C1748 vdd.n735 gnd 0.010831f
C1749 vdd.n736 gnd 0.010831f
C1750 vdd.n737 gnd 0.010831f
C1751 vdd.n738 gnd 0.010831f
C1752 vdd.n739 gnd 0.010831f
C1753 vdd.n740 gnd 0.010831f
C1754 vdd.n741 gnd 0.010831f
C1755 vdd.n742 gnd 0.010831f
C1756 vdd.n743 gnd 0.010831f
C1757 vdd.n744 gnd 0.010831f
C1758 vdd.n745 gnd 0.010831f
C1759 vdd.n746 gnd 0.010831f
C1760 vdd.n747 gnd 0.007279f
C1761 vdd.n748 gnd 0.010831f
C1762 vdd.n749 gnd 0.010831f
C1763 vdd.n750 gnd 0.010831f
C1764 vdd.n751 gnd 0.010831f
C1765 vdd.n752 gnd 0.010831f
C1766 vdd.n753 gnd 0.010831f
C1767 vdd.n754 gnd 0.010831f
C1768 vdd.n755 gnd 0.010831f
C1769 vdd.n756 gnd 0.010831f
C1770 vdd.n757 gnd 0.010831f
C1771 vdd.n758 gnd 0.010831f
C1772 vdd.n759 gnd 0.010831f
C1773 vdd.n760 gnd 0.010831f
C1774 vdd.n761 gnd 0.010831f
C1775 vdd.n762 gnd 0.010831f
C1776 vdd.n763 gnd 0.010831f
C1777 vdd.n764 gnd 0.010831f
C1778 vdd.n765 gnd 0.010831f
C1779 vdd.n766 gnd 0.010831f
C1780 vdd.n767 gnd 0.00863f
C1781 vdd.t43 gnd 0.133248f
C1782 vdd.t44 gnd 0.142406f
C1783 vdd.t42 gnd 0.17402f
C1784 vdd.n768 gnd 0.223069f
C1785 vdd.n769 gnd 0.187419f
C1786 vdd.n770 gnd 0.010831f
C1787 vdd.n771 gnd 0.010831f
C1788 vdd.n772 gnd 0.010831f
C1789 vdd.n773 gnd 0.010831f
C1790 vdd.n774 gnd 0.010831f
C1791 vdd.n775 gnd 0.010831f
C1792 vdd.n776 gnd 0.010831f
C1793 vdd.n777 gnd 0.010831f
C1794 vdd.n778 gnd 0.010831f
C1795 vdd.n779 gnd 0.010831f
C1796 vdd.n780 gnd 0.010831f
C1797 vdd.n781 gnd 0.010831f
C1798 vdd.n782 gnd 0.010831f
C1799 vdd.n783 gnd 0.006932f
C1800 vdd.n785 gnd 0.007365f
C1801 vdd.n786 gnd 0.007365f
C1802 vdd.n787 gnd 0.007365f
C1803 vdd.n788 gnd 0.007365f
C1804 vdd.n789 gnd 0.007365f
C1805 vdd.n790 gnd 0.007365f
C1806 vdd.n792 gnd 0.007365f
C1807 vdd.n793 gnd 0.007365f
C1808 vdd.n795 gnd 0.007365f
C1809 vdd.n796 gnd 0.005361f
C1810 vdd.n798 gnd 0.007365f
C1811 vdd.t29 gnd 0.297618f
C1812 vdd.t28 gnd 0.304649f
C1813 vdd.t26 gnd 0.194297f
C1814 vdd.n799 gnd 0.105007f
C1815 vdd.n800 gnd 0.059563f
C1816 vdd.n801 gnd 0.010526f
C1817 vdd.n802 gnd 0.017048f
C1818 vdd.n804 gnd 0.007365f
C1819 vdd.n805 gnd 0.752667f
C1820 vdd.n806 gnd 0.016133f
C1821 vdd.n807 gnd 0.016133f
C1822 vdd.n808 gnd 0.007365f
C1823 vdd.n809 gnd 0.017226f
C1824 vdd.n810 gnd 0.007365f
C1825 vdd.n811 gnd 0.007365f
C1826 vdd.n812 gnd 0.007365f
C1827 vdd.n813 gnd 0.007365f
C1828 vdd.n814 gnd 0.007365f
C1829 vdd.n816 gnd 0.007365f
C1830 vdd.n817 gnd 0.007365f
C1831 vdd.n819 gnd 0.007365f
C1832 vdd.n820 gnd 0.007365f
C1833 vdd.n822 gnd 0.007365f
C1834 vdd.n823 gnd 0.007365f
C1835 vdd.n825 gnd 0.007365f
C1836 vdd.n826 gnd 0.007365f
C1837 vdd.n828 gnd 0.007365f
C1838 vdd.n829 gnd 0.007365f
C1839 vdd.n831 gnd 0.007365f
C1840 vdd.t101 gnd 0.297618f
C1841 vdd.t100 gnd 0.304649f
C1842 vdd.t99 gnd 0.194297f
C1843 vdd.n832 gnd 0.105007f
C1844 vdd.n833 gnd 0.059563f
C1845 vdd.n834 gnd 0.007365f
C1846 vdd.n836 gnd 0.007365f
C1847 vdd.n837 gnd 0.007365f
C1848 vdd.t27 gnd 0.376333f
C1849 vdd.n838 gnd 0.007365f
C1850 vdd.n839 gnd 0.007365f
C1851 vdd.n840 gnd 0.007365f
C1852 vdd.n841 gnd 0.007365f
C1853 vdd.n842 gnd 0.007365f
C1854 vdd.n843 gnd 0.752667f
C1855 vdd.n844 gnd 0.007365f
C1856 vdd.n845 gnd 0.007365f
C1857 vdd.n846 gnd 0.636446f
C1858 vdd.n847 gnd 0.007365f
C1859 vdd.n848 gnd 0.007365f
C1860 vdd.n849 gnd 0.007365f
C1861 vdd.n850 gnd 0.007365f
C1862 vdd.n851 gnd 0.736064f
C1863 vdd.n852 gnd 0.007365f
C1864 vdd.n853 gnd 0.007365f
C1865 vdd.n854 gnd 0.007365f
C1866 vdd.n855 gnd 0.007365f
C1867 vdd.n856 gnd 0.007365f
C1868 vdd.n857 gnd 0.752667f
C1869 vdd.n858 gnd 0.007365f
C1870 vdd.n859 gnd 0.007365f
C1871 vdd.t114 gnd 0.376333f
C1872 vdd.n860 gnd 0.007365f
C1873 vdd.n861 gnd 0.007365f
C1874 vdd.n862 gnd 0.007365f
C1875 vdd.t0 gnd 0.376333f
C1876 vdd.n863 gnd 0.007365f
C1877 vdd.n864 gnd 0.007365f
C1878 vdd.n865 gnd 0.007365f
C1879 vdd.n866 gnd 0.007365f
C1880 vdd.n867 gnd 0.007365f
C1881 vdd.t53 gnd 0.315456f
C1882 vdd.n868 gnd 0.007365f
C1883 vdd.n869 gnd 0.007365f
C1884 vdd.n870 gnd 0.60324f
C1885 vdd.n871 gnd 0.007365f
C1886 vdd.t54 gnd 0.304649f
C1887 vdd.t52 gnd 0.194297f
C1888 vdd.t55 gnd 0.304649f
C1889 vdd.n872 gnd 0.171225f
C1890 vdd.n873 gnd 0.007365f
C1891 vdd.n874 gnd 0.007365f
C1892 vdd.n875 gnd 0.481485f
C1893 vdd.n876 gnd 0.007365f
C1894 vdd.n877 gnd 0.007365f
C1895 vdd.t123 gnd 0.110686f
C1896 vdd.n878 gnd 0.437211f
C1897 vdd.n879 gnd 0.007365f
C1898 vdd.n880 gnd 0.007365f
C1899 vdd.n881 gnd 0.007365f
C1900 vdd.n882 gnd 0.647515f
C1901 vdd.n883 gnd 0.007365f
C1902 vdd.n884 gnd 0.007365f
C1903 vdd.t21 gnd 0.376333f
C1904 vdd.n885 gnd 0.007365f
C1905 vdd.n886 gnd 0.007365f
C1906 vdd.n887 gnd 0.007365f
C1907 vdd.t125 gnd 0.376333f
C1908 vdd.n888 gnd 0.007365f
C1909 vdd.n889 gnd 0.007365f
C1910 vdd.t25 gnd 0.376333f
C1911 vdd.n890 gnd 0.007365f
C1912 vdd.n891 gnd 0.007365f
C1913 vdd.n892 gnd 0.007365f
C1914 vdd.t1 gnd 0.298853f
C1915 vdd.n893 gnd 0.007365f
C1916 vdd.n894 gnd 0.007365f
C1917 vdd.n895 gnd 0.619843f
C1918 vdd.n896 gnd 0.007365f
C1919 vdd.n897 gnd 0.007365f
C1920 vdd.n898 gnd 0.007365f
C1921 vdd.t109 gnd 0.376333f
C1922 vdd.n899 gnd 0.007365f
C1923 vdd.n900 gnd 0.007365f
C1924 vdd.t23 gnd 0.315456f
C1925 vdd.n901 gnd 0.453814f
C1926 vdd.n902 gnd 0.007365f
C1927 vdd.n903 gnd 0.007365f
C1928 vdd.n904 gnd 0.007365f
C1929 vdd.n905 gnd 0.392936f
C1930 vdd.n906 gnd 0.007365f
C1931 vdd.n907 gnd 0.007365f
C1932 vdd.t110 gnd 0.376333f
C1933 vdd.n908 gnd 0.007365f
C1934 vdd.n909 gnd 0.007365f
C1935 vdd.n910 gnd 0.007365f
C1936 vdd.n911 gnd 0.752667f
C1937 vdd.n912 gnd 0.007365f
C1938 vdd.n913 gnd 0.007365f
C1939 vdd.t127 gnd 0.254579f
C1940 vdd.t138 gnd 0.35973f
C1941 vdd.n914 gnd 0.007365f
C1942 vdd.n915 gnd 0.007365f
C1943 vdd.n916 gnd 0.007365f
C1944 vdd.n917 gnd 0.5645f
C1945 vdd.n918 gnd 0.007365f
C1946 vdd.n919 gnd 0.007365f
C1947 vdd.n920 gnd 0.007365f
C1948 vdd.n921 gnd 0.007365f
C1949 vdd.n922 gnd 0.007365f
C1950 vdd.t77 gnd 0.376333f
C1951 vdd.n923 gnd 0.007365f
C1952 vdd.n924 gnd 0.007365f
C1953 vdd.t115 gnd 0.376333f
C1954 vdd.n925 gnd 0.007365f
C1955 vdd.n926 gnd 0.016133f
C1956 vdd.n927 gnd 0.016133f
C1957 vdd.n928 gnd 0.896559f
C1958 vdd.n929 gnd 0.007365f
C1959 vdd.n930 gnd 0.007365f
C1960 vdd.t106 gnd 0.376333f
C1961 vdd.n931 gnd 0.016133f
C1962 vdd.n932 gnd 0.007365f
C1963 vdd.n933 gnd 0.007365f
C1964 vdd.t120 gnd 0.686255f
C1965 vdd.n951 gnd 0.017226f
C1966 vdd.n969 gnd 0.016133f
C1967 vdd.n970 gnd 0.007365f
C1968 vdd.n971 gnd 0.016133f
C1969 vdd.t98 gnd 0.297618f
C1970 vdd.t97 gnd 0.304649f
C1971 vdd.t96 gnd 0.194297f
C1972 vdd.n972 gnd 0.105007f
C1973 vdd.n973 gnd 0.059563f
C1974 vdd.n974 gnd 0.017048f
C1975 vdd.n975 gnd 0.007365f
C1976 vdd.n976 gnd 0.398471f
C1977 vdd.n977 gnd 0.016133f
C1978 vdd.n978 gnd 0.007365f
C1979 vdd.n979 gnd 0.017226f
C1980 vdd.n980 gnd 0.007365f
C1981 vdd.t75 gnd 0.297618f
C1982 vdd.t74 gnd 0.304649f
C1983 vdd.t72 gnd 0.194297f
C1984 vdd.n981 gnd 0.105007f
C1985 vdd.n982 gnd 0.059563f
C1986 vdd.n983 gnd 0.010526f
C1987 vdd.n984 gnd 0.007365f
C1988 vdd.n985 gnd 0.007365f
C1989 vdd.t73 gnd 0.376333f
C1990 vdd.n986 gnd 0.007365f
C1991 vdd.t118 gnd 0.376333f
C1992 vdd.n987 gnd 0.007365f
C1993 vdd.n988 gnd 0.007365f
C1994 vdd.n989 gnd 0.007365f
C1995 vdd.n990 gnd 0.007365f
C1996 vdd.n991 gnd 0.007365f
C1997 vdd.n992 gnd 0.752667f
C1998 vdd.n993 gnd 0.007365f
C1999 vdd.n994 gnd 0.007365f
C2000 vdd.t132 gnd 0.376333f
C2001 vdd.n995 gnd 0.007365f
C2002 vdd.n996 gnd 0.007365f
C2003 vdd.n997 gnd 0.007365f
C2004 vdd.n998 gnd 0.007365f
C2005 vdd.n999 gnd 0.498088f
C2006 vdd.n1000 gnd 0.007365f
C2007 vdd.n1001 gnd 0.007365f
C2008 vdd.n1002 gnd 0.007365f
C2009 vdd.n1003 gnd 0.007365f
C2010 vdd.n1004 gnd 0.007365f
C2011 vdd.n1005 gnd 0.664118f
C2012 vdd.n1006 gnd 0.007365f
C2013 vdd.n1007 gnd 0.007365f
C2014 vdd.t104 gnd 0.35973f
C2015 vdd.t20 gnd 0.254579f
C2016 vdd.n1008 gnd 0.007365f
C2017 vdd.n1009 gnd 0.007365f
C2018 vdd.n1010 gnd 0.007365f
C2019 vdd.t117 gnd 0.376333f
C2020 vdd.n1011 gnd 0.007365f
C2021 vdd.n1012 gnd 0.007365f
C2022 vdd.t128 gnd 0.376333f
C2023 vdd.n1013 gnd 0.007365f
C2024 vdd.n1014 gnd 0.007365f
C2025 vdd.n1015 gnd 0.007365f
C2026 vdd.t134 gnd 0.315456f
C2027 vdd.n1016 gnd 0.007365f
C2028 vdd.n1017 gnd 0.007365f
C2029 vdd.n1018 gnd 0.60324f
C2030 vdd.n1019 gnd 0.007365f
C2031 vdd.n1020 gnd 0.007365f
C2032 vdd.n1021 gnd 0.007365f
C2033 vdd.t112 gnd 0.376333f
C2034 vdd.n1022 gnd 0.007365f
C2035 vdd.n1023 gnd 0.007365f
C2036 vdd.t108 gnd 0.298853f
C2037 vdd.n1024 gnd 0.437211f
C2038 vdd.n1025 gnd 0.007365f
C2039 vdd.n1026 gnd 0.007365f
C2040 vdd.n1027 gnd 0.007365f
C2041 vdd.n1028 gnd 0.647515f
C2042 vdd.n1029 gnd 0.007365f
C2043 vdd.n1030 gnd 0.007365f
C2044 vdd.t19 gnd 0.376333f
C2045 vdd.n1031 gnd 0.007365f
C2046 vdd.n1032 gnd 0.007365f
C2047 vdd.n1033 gnd 0.007365f
C2048 vdd.n1034 gnd 0.752667f
C2049 vdd.n1035 gnd 0.007365f
C2050 vdd.n1036 gnd 0.007365f
C2051 vdd.t124 gnd 0.376333f
C2052 vdd.n1037 gnd 0.007365f
C2053 vdd.n1038 gnd 0.007365f
C2054 vdd.n1039 gnd 0.007365f
C2055 vdd.t22 gnd 0.110686f
C2056 vdd.n1040 gnd 0.007365f
C2057 vdd.n1041 gnd 0.007365f
C2058 vdd.n1042 gnd 0.007365f
C2059 vdd.t85 gnd 0.304649f
C2060 vdd.t83 gnd 0.194297f
C2061 vdd.t86 gnd 0.304649f
C2062 vdd.n1043 gnd 0.171225f
C2063 vdd.n1044 gnd 0.007365f
C2064 vdd.n1045 gnd 0.007365f
C2065 vdd.t122 gnd 0.376333f
C2066 vdd.n1046 gnd 0.007365f
C2067 vdd.n1047 gnd 0.007365f
C2068 vdd.t84 gnd 0.315456f
C2069 vdd.n1048 gnd 0.641981f
C2070 vdd.n1049 gnd 0.007365f
C2071 vdd.n1050 gnd 0.007365f
C2072 vdd.n1051 gnd 0.007365f
C2073 vdd.n1052 gnd 0.392936f
C2074 vdd.n1053 gnd 0.007365f
C2075 vdd.n1054 gnd 0.007365f
C2076 vdd.n1055 gnd 0.52576f
C2077 vdd.n1056 gnd 0.007365f
C2078 vdd.n1057 gnd 0.007365f
C2079 vdd.n1058 gnd 0.007365f
C2080 vdd.n1059 gnd 0.752667f
C2081 vdd.n1060 gnd 0.007365f
C2082 vdd.n1061 gnd 0.007365f
C2083 vdd.t18 gnd 0.376333f
C2084 vdd.n1062 gnd 0.007365f
C2085 vdd.n1063 gnd 0.007365f
C2086 vdd.n1064 gnd 0.007365f
C2087 vdd.n1065 gnd 0.752667f
C2088 vdd.n1066 gnd 0.007365f
C2089 vdd.n1067 gnd 0.007365f
C2090 vdd.n1068 gnd 0.007365f
C2091 vdd.n1069 gnd 0.007365f
C2092 vdd.n1070 gnd 0.007365f
C2093 vdd.t31 gnd 0.376333f
C2094 vdd.n1071 gnd 0.007365f
C2095 vdd.n1072 gnd 0.007365f
C2096 vdd.n1073 gnd 0.007365f
C2097 vdd.n1074 gnd 0.016133f
C2098 vdd.n1075 gnd 0.016133f
C2099 vdd.n1076 gnd 1.06259f
C2100 vdd.n1077 gnd 0.007365f
C2101 vdd.n1078 gnd 0.007365f
C2102 vdd.n1079 gnd 0.492554f
C2103 vdd.n1080 gnd 0.016133f
C2104 vdd.n1081 gnd 0.007365f
C2105 vdd.n1082 gnd 0.007365f
C2106 vdd.n1083 gnd 9.84001f
C2107 vdd.n1116 gnd 0.017226f
C2108 vdd.n1117 gnd 0.007365f
C2109 vdd.n1118 gnd 0.007365f
C2110 vdd.n1119 gnd 0.007365f
C2111 vdd.n1120 gnd 0.006932f
C2112 vdd.n1123 gnd 0.026762f
C2113 vdd.n1124 gnd 0.007236f
C2114 vdd.n1125 gnd 0.008718f
C2115 vdd.n1127 gnd 0.010831f
C2116 vdd.n1128 gnd 0.010831f
C2117 vdd.n1129 gnd 0.008718f
C2118 vdd.n1131 gnd 0.010831f
C2119 vdd.n1132 gnd 0.010831f
C2120 vdd.n1133 gnd 0.010831f
C2121 vdd.n1134 gnd 0.010831f
C2122 vdd.n1135 gnd 0.010831f
C2123 vdd.n1136 gnd 0.008718f
C2124 vdd.n1138 gnd 0.010831f
C2125 vdd.n1139 gnd 0.010831f
C2126 vdd.n1140 gnd 0.010831f
C2127 vdd.n1141 gnd 0.010831f
C2128 vdd.n1142 gnd 0.010831f
C2129 vdd.n1143 gnd 0.008718f
C2130 vdd.n1145 gnd 0.010831f
C2131 vdd.n1146 gnd 0.010831f
C2132 vdd.n1147 gnd 0.010831f
C2133 vdd.n1148 gnd 0.010831f
C2134 vdd.n1149 gnd 0.007279f
C2135 vdd.t92 gnd 0.133248f
C2136 vdd.t91 gnd 0.142406f
C2137 vdd.t90 gnd 0.17402f
C2138 vdd.n1150 gnd 0.223069f
C2139 vdd.n1151 gnd 0.187419f
C2140 vdd.n1153 gnd 0.010831f
C2141 vdd.n1154 gnd 0.010831f
C2142 vdd.n1155 gnd 0.008718f
C2143 vdd.n1156 gnd 0.010831f
C2144 vdd.n1158 gnd 0.010831f
C2145 vdd.n1159 gnd 0.010831f
C2146 vdd.n1160 gnd 0.010831f
C2147 vdd.n1161 gnd 0.010831f
C2148 vdd.n1162 gnd 0.008718f
C2149 vdd.n1164 gnd 0.010831f
C2150 vdd.n1165 gnd 0.010831f
C2151 vdd.n1166 gnd 0.010831f
C2152 vdd.n1167 gnd 0.010831f
C2153 vdd.n1168 gnd 0.010831f
C2154 vdd.n1169 gnd 0.008718f
C2155 vdd.n1171 gnd 0.010831f
C2156 vdd.n1172 gnd 0.010831f
C2157 vdd.n1173 gnd 0.010831f
C2158 vdd.n1174 gnd 0.010831f
C2159 vdd.n1175 gnd 0.010831f
C2160 vdd.n1176 gnd 0.008718f
C2161 vdd.n1178 gnd 0.010831f
C2162 vdd.n1179 gnd 0.010831f
C2163 vdd.n1180 gnd 0.010831f
C2164 vdd.n1181 gnd 0.010831f
C2165 vdd.n1182 gnd 0.010831f
C2166 vdd.n1183 gnd 0.008718f
C2167 vdd.n1185 gnd 0.010831f
C2168 vdd.n1186 gnd 0.010831f
C2169 vdd.n1187 gnd 0.010831f
C2170 vdd.n1188 gnd 0.010831f
C2171 vdd.n1189 gnd 0.00863f
C2172 vdd.t71 gnd 0.133248f
C2173 vdd.t70 gnd 0.142406f
C2174 vdd.t69 gnd 0.17402f
C2175 vdd.n1190 gnd 0.223069f
C2176 vdd.n1191 gnd 0.187419f
C2177 vdd.n1193 gnd 0.010831f
C2178 vdd.n1194 gnd 0.010831f
C2179 vdd.n1195 gnd 0.008718f
C2180 vdd.n1196 gnd 0.010831f
C2181 vdd.n1198 gnd 0.010831f
C2182 vdd.n1199 gnd 0.010831f
C2183 vdd.n1200 gnd 0.010831f
C2184 vdd.n1201 gnd 0.010831f
C2185 vdd.n1202 gnd 0.008718f
C2186 vdd.n1204 gnd 0.010831f
C2187 vdd.n1205 gnd 0.010831f
C2188 vdd.n1206 gnd 0.010831f
C2189 vdd.n1207 gnd 0.010831f
C2190 vdd.n1208 gnd 0.010831f
C2191 vdd.n1209 gnd 0.008718f
C2192 vdd.n1211 gnd 0.010831f
C2193 vdd.n1212 gnd 0.010831f
C2194 vdd.n1213 gnd 0.010831f
C2195 vdd.n1214 gnd 0.010831f
C2196 vdd.n1215 gnd 0.010831f
C2197 vdd.n1216 gnd 0.008718f
C2198 vdd.n1218 gnd 0.010831f
C2199 vdd.n1219 gnd 0.010831f
C2200 vdd.n1220 gnd 0.006932f
C2201 vdd.n1221 gnd 0.008718f
C2202 vdd.n1222 gnd 0.007365f
C2203 vdd.n1223 gnd 0.007365f
C2204 vdd.n1224 gnd 0.007365f
C2205 vdd.n1225 gnd 0.007365f
C2206 vdd.n1226 gnd 0.007365f
C2207 vdd.n1227 gnd 0.007365f
C2208 vdd.n1228 gnd 0.007365f
C2209 vdd.n1229 gnd 0.007365f
C2210 vdd.n1230 gnd 0.007365f
C2211 vdd.n1231 gnd 0.007365f
C2212 vdd.n1232 gnd 0.007365f
C2213 vdd.n1233 gnd 0.007365f
C2214 vdd.n1234 gnd 0.007365f
C2215 vdd.n1235 gnd 0.007365f
C2216 vdd.n1236 gnd 0.007365f
C2217 vdd.n1237 gnd 0.007365f
C2218 vdd.n1238 gnd 0.007365f
C2219 vdd.n1239 gnd 0.007365f
C2220 vdd.n1240 gnd 0.007365f
C2221 vdd.n1241 gnd 0.007365f
C2222 vdd.n1242 gnd 0.007365f
C2223 vdd.n1243 gnd 0.007365f
C2224 vdd.n1244 gnd 0.007365f
C2225 vdd.n1245 gnd 0.007365f
C2226 vdd.n1246 gnd 0.007365f
C2227 vdd.n1247 gnd 0.007365f
C2228 vdd.n1248 gnd 0.007365f
C2229 vdd.n1249 gnd 0.007365f
C2230 vdd.n1250 gnd 0.007365f
C2231 vdd.n1251 gnd 0.007365f
C2232 vdd.n1252 gnd 0.007365f
C2233 vdd.t32 gnd 0.297618f
C2234 vdd.t33 gnd 0.304649f
C2235 vdd.t30 gnd 0.194297f
C2236 vdd.n1253 gnd 0.105007f
C2237 vdd.n1254 gnd 0.059563f
C2238 vdd.n1255 gnd 0.010526f
C2239 vdd.n1256 gnd 0.007365f
C2240 vdd.n1257 gnd 0.007365f
C2241 vdd.n1258 gnd 0.007365f
C2242 vdd.n1259 gnd 0.007365f
C2243 vdd.n1260 gnd 0.007365f
C2244 vdd.n1261 gnd 0.007365f
C2245 vdd.n1262 gnd 0.007365f
C2246 vdd.n1263 gnd 0.007365f
C2247 vdd.n1264 gnd 0.007365f
C2248 vdd.n1265 gnd 0.007365f
C2249 vdd.n1266 gnd 0.007365f
C2250 vdd.n1267 gnd 0.007365f
C2251 vdd.n1268 gnd 0.007365f
C2252 vdd.n1269 gnd 0.007365f
C2253 vdd.n1270 gnd 0.007365f
C2254 vdd.n1271 gnd 0.007365f
C2255 vdd.n1272 gnd 0.007365f
C2256 vdd.t46 gnd 0.297618f
C2257 vdd.t47 gnd 0.304649f
C2258 vdd.t45 gnd 0.194297f
C2259 vdd.n1273 gnd 0.105007f
C2260 vdd.n1274 gnd 0.059563f
C2261 vdd.n1275 gnd 0.007365f
C2262 vdd.n1276 gnd 0.007365f
C2263 vdd.n1277 gnd 0.007365f
C2264 vdd.n1278 gnd 0.007365f
C2265 vdd.n1279 gnd 0.007365f
C2266 vdd.n1280 gnd 0.007365f
C2267 vdd.n1281 gnd 0.007365f
C2268 vdd.n1282 gnd 0.007365f
C2269 vdd.n1283 gnd 0.007365f
C2270 vdd.n1284 gnd 0.007365f
C2271 vdd.n1285 gnd 0.007365f
C2272 vdd.n1286 gnd 0.007365f
C2273 vdd.n1287 gnd 0.007365f
C2274 vdd.n1288 gnd 0.007365f
C2275 vdd.n1289 gnd 0.007365f
C2276 vdd.n1290 gnd 0.007365f
C2277 vdd.n1291 gnd 0.007365f
C2278 vdd.n1292 gnd 0.007365f
C2279 vdd.n1293 gnd 0.007365f
C2280 vdd.n1294 gnd 0.007365f
C2281 vdd.n1295 gnd 0.007365f
C2282 vdd.n1296 gnd 0.007365f
C2283 vdd.n1297 gnd 0.007365f
C2284 vdd.n1298 gnd 0.007365f
C2285 vdd.n1299 gnd 0.007365f
C2286 vdd.n1300 gnd 0.007365f
C2287 vdd.n1301 gnd 0.005361f
C2288 vdd.n1302 gnd 0.010526f
C2289 vdd.n1303 gnd 0.005686f
C2290 vdd.n1304 gnd 0.007365f
C2291 vdd.n1305 gnd 0.007365f
C2292 vdd.n1306 gnd 0.007365f
C2293 vdd.n1307 gnd 0.017226f
C2294 vdd.n1308 gnd 0.017226f
C2295 vdd.n1309 gnd 0.016133f
C2296 vdd.n1310 gnd 0.016133f
C2297 vdd.n1311 gnd 0.007365f
C2298 vdd.n1312 gnd 0.007365f
C2299 vdd.n1313 gnd 0.007365f
C2300 vdd.n1314 gnd 0.007365f
C2301 vdd.n1315 gnd 0.007365f
C2302 vdd.n1316 gnd 0.007365f
C2303 vdd.n1317 gnd 0.007365f
C2304 vdd.n1318 gnd 0.007365f
C2305 vdd.n1319 gnd 0.007365f
C2306 vdd.n1320 gnd 0.007365f
C2307 vdd.n1321 gnd 0.007365f
C2308 vdd.n1322 gnd 0.007365f
C2309 vdd.n1323 gnd 0.007365f
C2310 vdd.n1324 gnd 0.007365f
C2311 vdd.n1325 gnd 0.007365f
C2312 vdd.n1326 gnd 0.007365f
C2313 vdd.n1327 gnd 0.007365f
C2314 vdd.n1328 gnd 0.007365f
C2315 vdd.n1329 gnd 0.007365f
C2316 vdd.n1330 gnd 0.007365f
C2317 vdd.n1331 gnd 0.007365f
C2318 vdd.n1332 gnd 0.007365f
C2319 vdd.n1333 gnd 0.007365f
C2320 vdd.n1334 gnd 0.007365f
C2321 vdd.n1335 gnd 0.007365f
C2322 vdd.n1336 gnd 0.007365f
C2323 vdd.n1337 gnd 0.007365f
C2324 vdd.n1338 gnd 0.44828f
C2325 vdd.n1339 gnd 0.007365f
C2326 vdd.n1340 gnd 0.007365f
C2327 vdd.n1341 gnd 0.007365f
C2328 vdd.n1342 gnd 0.007365f
C2329 vdd.n1343 gnd 0.007365f
C2330 vdd.n1344 gnd 0.007365f
C2331 vdd.n1345 gnd 0.007365f
C2332 vdd.n1346 gnd 0.007365f
C2333 vdd.n1347 gnd 0.007365f
C2334 vdd.n1348 gnd 0.007365f
C2335 vdd.n1349 gnd 0.007365f
C2336 vdd.n1350 gnd 0.007365f
C2337 vdd.n1351 gnd 0.007365f
C2338 vdd.n1352 gnd 0.007365f
C2339 vdd.n1353 gnd 0.007365f
C2340 vdd.n1354 gnd 0.007365f
C2341 vdd.n1355 gnd 0.007365f
C2342 vdd.n1356 gnd 0.007365f
C2343 vdd.n1357 gnd 0.007365f
C2344 vdd.n1358 gnd 0.007365f
C2345 vdd.n1359 gnd 0.237976f
C2346 vdd.n1360 gnd 0.007365f
C2347 vdd.n1361 gnd 0.007365f
C2348 vdd.n1362 gnd 0.007365f
C2349 vdd.n1363 gnd 0.007365f
C2350 vdd.n1364 gnd 0.007365f
C2351 vdd.n1365 gnd 0.007365f
C2352 vdd.n1366 gnd 0.007365f
C2353 vdd.n1367 gnd 0.007365f
C2354 vdd.n1368 gnd 0.007365f
C2355 vdd.n1369 gnd 0.007365f
C2356 vdd.n1370 gnd 0.007365f
C2357 vdd.n1371 gnd 0.007365f
C2358 vdd.n1372 gnd 0.007365f
C2359 vdd.n1373 gnd 0.007365f
C2360 vdd.n1374 gnd 0.007365f
C2361 vdd.n1375 gnd 0.007365f
C2362 vdd.n1376 gnd 0.007365f
C2363 vdd.n1377 gnd 0.007365f
C2364 vdd.n1378 gnd 0.007365f
C2365 vdd.n1379 gnd 0.007365f
C2366 vdd.n1380 gnd 0.007365f
C2367 vdd.n1381 gnd 0.007365f
C2368 vdd.n1382 gnd 0.007365f
C2369 vdd.n1383 gnd 0.007365f
C2370 vdd.n1384 gnd 0.007365f
C2371 vdd.n1385 gnd 0.007365f
C2372 vdd.n1386 gnd 0.007365f
C2373 vdd.n1387 gnd 0.016133f
C2374 vdd.n1388 gnd 0.016133f
C2375 vdd.n1389 gnd 0.017226f
C2376 vdd.n1390 gnd 0.007365f
C2377 vdd.n1391 gnd 0.007365f
C2378 vdd.n1392 gnd 0.005686f
C2379 vdd.n1393 gnd 0.007365f
C2380 vdd.n1394 gnd 0.007365f
C2381 vdd.n1395 gnd 0.005361f
C2382 vdd.n1396 gnd 0.007365f
C2383 vdd.n1397 gnd 0.007365f
C2384 vdd.n1398 gnd 0.007365f
C2385 vdd.n1399 gnd 0.007365f
C2386 vdd.n1400 gnd 0.007365f
C2387 vdd.n1401 gnd 0.007365f
C2388 vdd.n1402 gnd 0.007365f
C2389 vdd.n1403 gnd 0.007365f
C2390 vdd.n1404 gnd 0.007365f
C2391 vdd.n1405 gnd 0.007365f
C2392 vdd.n1406 gnd 0.007365f
C2393 vdd.n1407 gnd 0.007365f
C2394 vdd.n1408 gnd 0.007365f
C2395 vdd.n1409 gnd 0.007365f
C2396 vdd.n1410 gnd 0.007365f
C2397 vdd.n1411 gnd 0.007365f
C2398 vdd.n1412 gnd 0.007365f
C2399 vdd.n1413 gnd 0.007365f
C2400 vdd.n1414 gnd 0.007365f
C2401 vdd.n1415 gnd 0.007365f
C2402 vdd.n1416 gnd 0.007365f
C2403 vdd.n1417 gnd 0.007365f
C2404 vdd.n1418 gnd 0.007365f
C2405 vdd.n1419 gnd 0.007365f
C2406 vdd.n1420 gnd 0.007365f
C2407 vdd.n1421 gnd 0.007365f
C2408 vdd.n1422 gnd 0.029519f
C2409 vdd.n1424 gnd 0.026762f
C2410 vdd.n1425 gnd 0.008718f
C2411 vdd.n1427 gnd 0.010831f
C2412 vdd.n1428 gnd 0.008718f
C2413 vdd.n1429 gnd 0.010831f
C2414 vdd.n1431 gnd 0.010831f
C2415 vdd.n1432 gnd 0.010831f
C2416 vdd.n1434 gnd 0.010831f
C2417 vdd.n1435 gnd 0.007236f
C2418 vdd.t39 gnd 0.553432f
C2419 vdd.n1436 gnd 0.010831f
C2420 vdd.n1437 gnd 0.026762f
C2421 vdd.n1438 gnd 0.008718f
C2422 vdd.n1439 gnd 0.010831f
C2423 vdd.n1440 gnd 0.008718f
C2424 vdd.n1441 gnd 0.010831f
C2425 vdd.n1442 gnd 1.10686f
C2426 vdd.n1443 gnd 0.010831f
C2427 vdd.n1444 gnd 0.008718f
C2428 vdd.n1445 gnd 0.008718f
C2429 vdd.n1446 gnd 0.010831f
C2430 vdd.n1447 gnd 0.008718f
C2431 vdd.n1448 gnd 0.010831f
C2432 vdd.t188 gnd 0.553432f
C2433 vdd.n1449 gnd 0.010831f
C2434 vdd.n1450 gnd 0.008718f
C2435 vdd.n1451 gnd 0.010831f
C2436 vdd.n1452 gnd 0.008718f
C2437 vdd.n1453 gnd 0.010831f
C2438 vdd.t148 gnd 0.553432f
C2439 vdd.n1454 gnd 0.010831f
C2440 vdd.n1455 gnd 0.008718f
C2441 vdd.n1456 gnd 0.010831f
C2442 vdd.n1457 gnd 0.008718f
C2443 vdd.n1458 gnd 0.010831f
C2444 vdd.n1459 gnd 0.891025f
C2445 vdd.n1460 gnd 0.918696f
C2446 vdd.t220 gnd 0.553432f
C2447 vdd.n1461 gnd 0.010831f
C2448 vdd.n1462 gnd 0.008718f
C2449 vdd.n1463 gnd 0.010831f
C2450 vdd.n1464 gnd 0.008718f
C2451 vdd.n1465 gnd 0.010831f
C2452 vdd.n1466 gnd 0.702858f
C2453 vdd.n1467 gnd 0.010831f
C2454 vdd.n1468 gnd 0.008718f
C2455 vdd.n1469 gnd 0.010831f
C2456 vdd.n1470 gnd 0.008718f
C2457 vdd.n1471 gnd 0.010831f
C2458 vdd.t156 gnd 0.553432f
C2459 vdd.t243 gnd 0.553432f
C2460 vdd.n1472 gnd 0.010831f
C2461 vdd.n1473 gnd 0.008718f
C2462 vdd.n1474 gnd 0.010831f
C2463 vdd.n1475 gnd 0.008718f
C2464 vdd.n1476 gnd 0.010831f
C2465 vdd.t208 gnd 0.553432f
C2466 vdd.n1477 gnd 0.010831f
C2467 vdd.n1478 gnd 0.008718f
C2468 vdd.n1479 gnd 0.010831f
C2469 vdd.n1480 gnd 0.008718f
C2470 vdd.n1481 gnd 0.010831f
C2471 vdd.t167 gnd 0.553432f
C2472 vdd.n1482 gnd 0.780339f
C2473 vdd.n1483 gnd 0.010831f
C2474 vdd.n1484 gnd 0.008718f
C2475 vdd.n1485 gnd 0.010831f
C2476 vdd.n1486 gnd 0.008718f
C2477 vdd.n1487 gnd 0.010831f
C2478 vdd.n1488 gnd 0.868888f
C2479 vdd.n1489 gnd 0.010831f
C2480 vdd.n1490 gnd 0.008718f
C2481 vdd.n1491 gnd 0.010831f
C2482 vdd.n1492 gnd 0.008718f
C2483 vdd.n1493 gnd 0.010831f
C2484 vdd.n1494 gnd 0.680721f
C2485 vdd.t238 gnd 0.553432f
C2486 vdd.n1495 gnd 0.010831f
C2487 vdd.n1496 gnd 0.008718f
C2488 vdd.n1497 gnd 0.010831f
C2489 vdd.n1498 gnd 0.008718f
C2490 vdd.n1499 gnd 0.010831f
C2491 vdd.t154 gnd 0.553432f
C2492 vdd.n1500 gnd 0.010831f
C2493 vdd.n1501 gnd 0.008718f
C2494 vdd.n1502 gnd 0.010831f
C2495 vdd.n1503 gnd 0.008718f
C2496 vdd.n1504 gnd 0.010831f
C2497 vdd.t179 gnd 0.553432f
C2498 vdd.n1505 gnd 0.614309f
C2499 vdd.n1506 gnd 0.010831f
C2500 vdd.n1507 gnd 0.008718f
C2501 vdd.n1508 gnd 0.010831f
C2502 vdd.n1509 gnd 0.008718f
C2503 vdd.n1510 gnd 0.010831f
C2504 vdd.t181 gnd 0.553432f
C2505 vdd.n1511 gnd 0.010831f
C2506 vdd.n1512 gnd 0.008718f
C2507 vdd.n1513 gnd 0.010831f
C2508 vdd.n1514 gnd 0.008718f
C2509 vdd.n1515 gnd 0.010831f
C2510 vdd.n1516 gnd 0.84675f
C2511 vdd.n1517 gnd 0.918696f
C2512 vdd.t144 gnd 0.553432f
C2513 vdd.n1518 gnd 0.010831f
C2514 vdd.n1519 gnd 0.008718f
C2515 vdd.n1520 gnd 0.010831f
C2516 vdd.n1521 gnd 0.008718f
C2517 vdd.n1522 gnd 0.010831f
C2518 vdd.n1523 gnd 0.658584f
C2519 vdd.n1524 gnd 0.010831f
C2520 vdd.n1525 gnd 0.008718f
C2521 vdd.n1526 gnd 0.010831f
C2522 vdd.n1527 gnd 0.008718f
C2523 vdd.n1528 gnd 0.010831f
C2524 vdd.t236 gnd 0.553432f
C2525 vdd.t210 gnd 0.553432f
C2526 vdd.n1529 gnd 0.010831f
C2527 vdd.n1530 gnd 0.008718f
C2528 vdd.n1531 gnd 0.010831f
C2529 vdd.n1532 gnd 0.008718f
C2530 vdd.n1533 gnd 0.010831f
C2531 vdd.t140 gnd 0.553432f
C2532 vdd.n1534 gnd 0.010831f
C2533 vdd.n1535 gnd 0.008718f
C2534 vdd.n1536 gnd 0.010831f
C2535 vdd.n1537 gnd 0.008718f
C2536 vdd.n1538 gnd 0.010831f
C2537 vdd.t196 gnd 0.553432f
C2538 vdd.n1539 gnd 0.824613f
C2539 vdd.n1540 gnd 0.010831f
C2540 vdd.n1541 gnd 0.008718f
C2541 vdd.n1542 gnd 0.010831f
C2542 vdd.n1543 gnd 0.008718f
C2543 vdd.n1544 gnd 0.010831f
C2544 vdd.n1545 gnd 1.10686f
C2545 vdd.n1546 gnd 0.010831f
C2546 vdd.n1547 gnd 0.008718f
C2547 vdd.n1548 gnd 0.026201f
C2548 vdd.n1549 gnd 0.007236f
C2549 vdd.n1550 gnd 0.026201f
C2550 vdd.t63 gnd 0.553432f
C2551 vdd.n1551 gnd 0.026201f
C2552 vdd.n1552 gnd 0.007236f
C2553 vdd.n1553 gnd 0.010831f
C2554 vdd.n1554 gnd 0.008718f
C2555 vdd.n1555 gnd 0.010831f
C2556 vdd.n1586 gnd 0.026762f
C2557 vdd.n1587 gnd 1.63262f
C2558 vdd.n1588 gnd 0.010831f
C2559 vdd.n1589 gnd 0.008718f
C2560 vdd.n1590 gnd 0.010831f
C2561 vdd.n1591 gnd 0.010831f
C2562 vdd.n1592 gnd 0.010831f
C2563 vdd.n1593 gnd 0.010831f
C2564 vdd.n1594 gnd 0.010831f
C2565 vdd.n1595 gnd 0.008718f
C2566 vdd.n1596 gnd 0.010831f
C2567 vdd.n1597 gnd 0.010831f
C2568 vdd.n1598 gnd 0.010831f
C2569 vdd.n1599 gnd 0.010831f
C2570 vdd.n1600 gnd 0.010831f
C2571 vdd.n1601 gnd 0.008718f
C2572 vdd.n1602 gnd 0.010831f
C2573 vdd.n1603 gnd 0.010831f
C2574 vdd.n1604 gnd 0.010831f
C2575 vdd.n1605 gnd 0.010831f
C2576 vdd.n1606 gnd 0.010831f
C2577 vdd.n1607 gnd 0.008718f
C2578 vdd.n1608 gnd 0.010831f
C2579 vdd.n1609 gnd 0.010831f
C2580 vdd.n1610 gnd 0.010831f
C2581 vdd.n1611 gnd 0.010831f
C2582 vdd.n1612 gnd 0.010831f
C2583 vdd.t94 gnd 0.133248f
C2584 vdd.t95 gnd 0.142406f
C2585 vdd.t93 gnd 0.17402f
C2586 vdd.n1613 gnd 0.223069f
C2587 vdd.n1614 gnd 0.18829f
C2588 vdd.n1615 gnd 0.018655f
C2589 vdd.n1616 gnd 0.010831f
C2590 vdd.n1617 gnd 0.010831f
C2591 vdd.n1618 gnd 0.010831f
C2592 vdd.n1619 gnd 0.010831f
C2593 vdd.n1620 gnd 0.010831f
C2594 vdd.n1621 gnd 0.008718f
C2595 vdd.n1622 gnd 0.010831f
C2596 vdd.n1623 gnd 0.010831f
C2597 vdd.n1624 gnd 0.010831f
C2598 vdd.n1625 gnd 0.010831f
C2599 vdd.n1626 gnd 0.010831f
C2600 vdd.n1627 gnd 0.008718f
C2601 vdd.n1628 gnd 0.010831f
C2602 vdd.n1629 gnd 0.010831f
C2603 vdd.n1630 gnd 0.010831f
C2604 vdd.n1631 gnd 0.010831f
C2605 vdd.n1632 gnd 0.010831f
C2606 vdd.n1633 gnd 0.008718f
C2607 vdd.n1634 gnd 0.010831f
C2608 vdd.n1635 gnd 0.010831f
C2609 vdd.n1636 gnd 0.010831f
C2610 vdd.n1637 gnd 0.010831f
C2611 vdd.n1638 gnd 0.010831f
C2612 vdd.n1639 gnd 0.008718f
C2613 vdd.n1640 gnd 0.010831f
C2614 vdd.n1641 gnd 0.010831f
C2615 vdd.n1642 gnd 0.010831f
C2616 vdd.n1643 gnd 0.010831f
C2617 vdd.n1644 gnd 0.010831f
C2618 vdd.n1645 gnd 0.008718f
C2619 vdd.n1646 gnd 0.010831f
C2620 vdd.n1647 gnd 0.010831f
C2621 vdd.n1648 gnd 0.010831f
C2622 vdd.n1649 gnd 0.010831f
C2623 vdd.n1650 gnd 0.008718f
C2624 vdd.n1651 gnd 0.010831f
C2625 vdd.n1652 gnd 0.010831f
C2626 vdd.n1653 gnd 0.010831f
C2627 vdd.n1654 gnd 0.010831f
C2628 vdd.n1655 gnd 0.010831f
C2629 vdd.n1656 gnd 0.008718f
C2630 vdd.n1657 gnd 0.010831f
C2631 vdd.n1658 gnd 0.010831f
C2632 vdd.n1659 gnd 0.010831f
C2633 vdd.n1660 gnd 0.010831f
C2634 vdd.n1661 gnd 0.010831f
C2635 vdd.n1662 gnd 0.008718f
C2636 vdd.n1663 gnd 0.010831f
C2637 vdd.n1664 gnd 0.010831f
C2638 vdd.n1665 gnd 0.010831f
C2639 vdd.n1666 gnd 0.010831f
C2640 vdd.n1667 gnd 0.010831f
C2641 vdd.n1668 gnd 0.008718f
C2642 vdd.n1669 gnd 0.010831f
C2643 vdd.n1670 gnd 0.010831f
C2644 vdd.n1671 gnd 0.010831f
C2645 vdd.n1672 gnd 0.010831f
C2646 vdd.n1673 gnd 0.010831f
C2647 vdd.n1674 gnd 0.008718f
C2648 vdd.n1675 gnd 0.010831f
C2649 vdd.n1676 gnd 0.010831f
C2650 vdd.n1677 gnd 0.010831f
C2651 vdd.n1678 gnd 0.010831f
C2652 vdd.t64 gnd 0.133248f
C2653 vdd.t65 gnd 0.142406f
C2654 vdd.t62 gnd 0.17402f
C2655 vdd.n1679 gnd 0.223069f
C2656 vdd.n1680 gnd 0.18829f
C2657 vdd.n1681 gnd 0.014297f
C2658 vdd.n1682 gnd 0.004141f
C2659 vdd.n1683 gnd 0.026762f
C2660 vdd.n1684 gnd 0.010831f
C2661 vdd.n1685 gnd 0.004577f
C2662 vdd.n1686 gnd 0.008718f
C2663 vdd.n1687 gnd 0.008718f
C2664 vdd.n1688 gnd 0.010831f
C2665 vdd.n1689 gnd 0.010831f
C2666 vdd.n1690 gnd 0.010831f
C2667 vdd.n1691 gnd 0.008718f
C2668 vdd.n1692 gnd 0.008718f
C2669 vdd.n1693 gnd 0.008718f
C2670 vdd.n1694 gnd 0.010831f
C2671 vdd.n1695 gnd 0.010831f
C2672 vdd.n1696 gnd 0.010831f
C2673 vdd.n1697 gnd 0.008718f
C2674 vdd.n1698 gnd 0.008718f
C2675 vdd.n1699 gnd 0.008718f
C2676 vdd.n1700 gnd 0.010831f
C2677 vdd.n1701 gnd 0.010831f
C2678 vdd.n1702 gnd 0.010831f
C2679 vdd.n1703 gnd 0.008718f
C2680 vdd.n1704 gnd 0.008718f
C2681 vdd.n1705 gnd 0.008718f
C2682 vdd.n1706 gnd 0.010831f
C2683 vdd.n1707 gnd 0.010831f
C2684 vdd.n1708 gnd 0.010831f
C2685 vdd.n1709 gnd 0.008718f
C2686 vdd.n1710 gnd 0.008718f
C2687 vdd.n1711 gnd 0.008718f
C2688 vdd.n1712 gnd 0.010831f
C2689 vdd.n1713 gnd 0.010831f
C2690 vdd.n1714 gnd 0.010831f
C2691 vdd.n1715 gnd 0.00863f
C2692 vdd.n1716 gnd 0.010831f
C2693 vdd.t81 gnd 0.133248f
C2694 vdd.t82 gnd 0.142406f
C2695 vdd.t80 gnd 0.17402f
C2696 vdd.n1717 gnd 0.223069f
C2697 vdd.n1718 gnd 0.18829f
C2698 vdd.n1719 gnd 0.018655f
C2699 vdd.n1720 gnd 0.005928f
C2700 vdd.n1721 gnd 0.010831f
C2701 vdd.n1722 gnd 0.010831f
C2702 vdd.n1723 gnd 0.010831f
C2703 vdd.n1724 gnd 0.008718f
C2704 vdd.n1725 gnd 0.008718f
C2705 vdd.n1726 gnd 0.008718f
C2706 vdd.n1727 gnd 0.010831f
C2707 vdd.n1728 gnd 0.010831f
C2708 vdd.n1729 gnd 0.010831f
C2709 vdd.n1730 gnd 0.008718f
C2710 vdd.n1731 gnd 0.008718f
C2711 vdd.n1732 gnd 0.008718f
C2712 vdd.n1733 gnd 0.010831f
C2713 vdd.n1734 gnd 0.010831f
C2714 vdd.n1735 gnd 0.010831f
C2715 vdd.n1736 gnd 0.008718f
C2716 vdd.n1737 gnd 0.008718f
C2717 vdd.n1738 gnd 0.008718f
C2718 vdd.n1739 gnd 0.010831f
C2719 vdd.n1740 gnd 0.010831f
C2720 vdd.n1741 gnd 0.010831f
C2721 vdd.n1742 gnd 0.008718f
C2722 vdd.n1743 gnd 0.008718f
C2723 vdd.n1744 gnd 0.008718f
C2724 vdd.n1745 gnd 0.010831f
C2725 vdd.n1746 gnd 0.010831f
C2726 vdd.n1747 gnd 0.010831f
C2727 vdd.n1748 gnd 0.008718f
C2728 vdd.n1749 gnd 0.008718f
C2729 vdd.n1750 gnd 0.007279f
C2730 vdd.n1751 gnd 0.010831f
C2731 vdd.n1752 gnd 0.010831f
C2732 vdd.n1753 gnd 0.010831f
C2733 vdd.n1754 gnd 0.007279f
C2734 vdd.n1755 gnd 0.008718f
C2735 vdd.n1756 gnd 0.008718f
C2736 vdd.n1757 gnd 0.010831f
C2737 vdd.n1758 gnd 0.010831f
C2738 vdd.n1759 gnd 0.010831f
C2739 vdd.n1760 gnd 0.008718f
C2740 vdd.n1761 gnd 0.008718f
C2741 vdd.n1762 gnd 0.008718f
C2742 vdd.n1763 gnd 0.010831f
C2743 vdd.n1764 gnd 0.010831f
C2744 vdd.n1765 gnd 0.010831f
C2745 vdd.n1766 gnd 0.008718f
C2746 vdd.n1767 gnd 0.008718f
C2747 vdd.n1768 gnd 0.008718f
C2748 vdd.n1769 gnd 0.010831f
C2749 vdd.n1770 gnd 0.010831f
C2750 vdd.n1771 gnd 0.010831f
C2751 vdd.n1772 gnd 0.008718f
C2752 vdd.n1773 gnd 0.008718f
C2753 vdd.n1774 gnd 0.008718f
C2754 vdd.n1775 gnd 0.010831f
C2755 vdd.n1776 gnd 0.010831f
C2756 vdd.n1777 gnd 0.010831f
C2757 vdd.n1778 gnd 0.008718f
C2758 vdd.n1779 gnd 0.010831f
C2759 vdd.n1780 gnd 2.62327f
C2760 vdd.n1782 gnd 0.026762f
C2761 vdd.n1783 gnd 0.007236f
C2762 vdd.n1784 gnd 0.026762f
C2763 vdd.n1785 gnd 0.026201f
C2764 vdd.n1786 gnd 0.010831f
C2765 vdd.n1787 gnd 0.008718f
C2766 vdd.n1788 gnd 0.010831f
C2767 vdd.n1789 gnd 0.558966f
C2768 vdd.n1790 gnd 0.010831f
C2769 vdd.n1791 gnd 0.008718f
C2770 vdd.n1792 gnd 0.010831f
C2771 vdd.n1793 gnd 0.010831f
C2772 vdd.n1794 gnd 0.010831f
C2773 vdd.n1795 gnd 0.008718f
C2774 vdd.n1796 gnd 0.010831f
C2775 vdd.n1797 gnd 1.01278f
C2776 vdd.n1798 gnd 1.10686f
C2777 vdd.n1799 gnd 0.010831f
C2778 vdd.n1800 gnd 0.008718f
C2779 vdd.n1801 gnd 0.010831f
C2780 vdd.n1802 gnd 0.010831f
C2781 vdd.n1803 gnd 0.010831f
C2782 vdd.n1804 gnd 0.008718f
C2783 vdd.n1805 gnd 0.010831f
C2784 vdd.n1806 gnd 0.647515f
C2785 vdd.n1807 gnd 0.010831f
C2786 vdd.n1808 gnd 0.008718f
C2787 vdd.n1809 gnd 0.010831f
C2788 vdd.n1810 gnd 0.010831f
C2789 vdd.n1811 gnd 0.010831f
C2790 vdd.n1812 gnd 0.008718f
C2791 vdd.n1813 gnd 0.010831f
C2792 vdd.n1814 gnd 0.636446f
C2793 vdd.n1815 gnd 0.835682f
C2794 vdd.n1816 gnd 0.010831f
C2795 vdd.n1817 gnd 0.008718f
C2796 vdd.n1818 gnd 0.010831f
C2797 vdd.n1819 gnd 0.010831f
C2798 vdd.n1820 gnd 0.010831f
C2799 vdd.n1821 gnd 0.008718f
C2800 vdd.n1822 gnd 0.010831f
C2801 vdd.n1823 gnd 0.918696f
C2802 vdd.n1824 gnd 0.010831f
C2803 vdd.n1825 gnd 0.008718f
C2804 vdd.n1826 gnd 0.010831f
C2805 vdd.n1827 gnd 0.010831f
C2806 vdd.n1828 gnd 0.010831f
C2807 vdd.n1829 gnd 0.008718f
C2808 vdd.n1830 gnd 0.010831f
C2809 vdd.t150 gnd 0.553432f
C2810 vdd.n1831 gnd 0.813544f
C2811 vdd.n1832 gnd 0.010831f
C2812 vdd.n1833 gnd 0.008718f
C2813 vdd.n1834 gnd 0.010831f
C2814 vdd.n1835 gnd 0.010831f
C2815 vdd.n1836 gnd 0.010831f
C2816 vdd.n1837 gnd 0.008718f
C2817 vdd.n1838 gnd 0.010831f
C2818 vdd.n1839 gnd 0.625378f
C2819 vdd.n1840 gnd 0.010831f
C2820 vdd.n1841 gnd 0.008718f
C2821 vdd.n1842 gnd 0.010831f
C2822 vdd.n1843 gnd 0.010831f
C2823 vdd.n1844 gnd 0.010831f
C2824 vdd.n1845 gnd 0.008718f
C2825 vdd.n1846 gnd 0.010831f
C2826 vdd.n1847 gnd 0.802476f
C2827 vdd.n1848 gnd 0.669652f
C2828 vdd.n1849 gnd 0.010831f
C2829 vdd.n1850 gnd 0.008718f
C2830 vdd.n1851 gnd 0.010831f
C2831 vdd.n1852 gnd 0.010831f
C2832 vdd.n1853 gnd 0.010831f
C2833 vdd.n1854 gnd 0.008718f
C2834 vdd.n1855 gnd 0.010831f
C2835 vdd.n1856 gnd 0.857819f
C2836 vdd.n1857 gnd 0.010831f
C2837 vdd.n1858 gnd 0.008718f
C2838 vdd.n1859 gnd 0.010831f
C2839 vdd.n1860 gnd 0.010831f
C2840 vdd.n1861 gnd 0.010831f
C2841 vdd.n1862 gnd 0.008718f
C2842 vdd.n1863 gnd 0.010831f
C2843 vdd.t240 gnd 0.553432f
C2844 vdd.n1864 gnd 0.918696f
C2845 vdd.n1865 gnd 0.010831f
C2846 vdd.n1866 gnd 0.008718f
C2847 vdd.n1867 gnd 0.010831f
C2848 vdd.n1868 gnd 0.008324f
C2849 vdd.n1869 gnd 0.005944f
C2850 vdd.n1870 gnd 0.005516f
C2851 vdd.n1871 gnd 0.003051f
C2852 vdd.n1872 gnd 0.007006f
C2853 vdd.n1873 gnd 0.002964f
C2854 vdd.n1874 gnd 0.003138f
C2855 vdd.n1875 gnd 0.005516f
C2856 vdd.n1876 gnd 0.002964f
C2857 vdd.n1877 gnd 0.007006f
C2858 vdd.n1878 gnd 0.003138f
C2859 vdd.n1879 gnd 0.005516f
C2860 vdd.n1880 gnd 0.002964f
C2861 vdd.n1881 gnd 0.005254f
C2862 vdd.n1882 gnd 0.00527f
C2863 vdd.t189 gnd 0.015051f
C2864 vdd.n1883 gnd 0.033489f
C2865 vdd.n1884 gnd 0.174283f
C2866 vdd.n1885 gnd 0.002964f
C2867 vdd.n1886 gnd 0.003138f
C2868 vdd.n1887 gnd 0.007006f
C2869 vdd.n1888 gnd 0.007006f
C2870 vdd.n1889 gnd 0.003138f
C2871 vdd.n1890 gnd 0.002964f
C2872 vdd.n1891 gnd 0.005516f
C2873 vdd.n1892 gnd 0.005516f
C2874 vdd.n1893 gnd 0.002964f
C2875 vdd.n1894 gnd 0.003138f
C2876 vdd.n1895 gnd 0.007006f
C2877 vdd.n1896 gnd 0.007006f
C2878 vdd.n1897 gnd 0.003138f
C2879 vdd.n1898 gnd 0.002964f
C2880 vdd.n1899 gnd 0.005516f
C2881 vdd.n1900 gnd 0.005516f
C2882 vdd.n1901 gnd 0.002964f
C2883 vdd.n1902 gnd 0.003138f
C2884 vdd.n1903 gnd 0.007006f
C2885 vdd.n1904 gnd 0.007006f
C2886 vdd.n1905 gnd 0.016563f
C2887 vdd.n1906 gnd 0.003051f
C2888 vdd.n1907 gnd 0.002964f
C2889 vdd.n1908 gnd 0.014257f
C2890 vdd.n1909 gnd 0.009953f
C2891 vdd.t221 gnd 0.03487f
C2892 vdd.t278 gnd 0.03487f
C2893 vdd.n1910 gnd 0.239652f
C2894 vdd.n1911 gnd 0.188449f
C2895 vdd.t244 gnd 0.03487f
C2896 vdd.t293 gnd 0.03487f
C2897 vdd.n1912 gnd 0.239652f
C2898 vdd.n1913 gnd 0.152078f
C2899 vdd.t209 gnd 0.03487f
C2900 vdd.t157 gnd 0.03487f
C2901 vdd.n1914 gnd 0.239652f
C2902 vdd.n1915 gnd 0.152078f
C2903 vdd.t233 gnd 0.03487f
C2904 vdd.t168 gnd 0.03487f
C2905 vdd.n1916 gnd 0.239652f
C2906 vdd.n1917 gnd 0.152078f
C2907 vdd.t282 gnd 0.03487f
C2908 vdd.t298 gnd 0.03487f
C2909 vdd.n1918 gnd 0.239652f
C2910 vdd.n1919 gnd 0.152078f
C2911 vdd.t255 gnd 0.03487f
C2912 vdd.t172 gnd 0.03487f
C2913 vdd.n1920 gnd 0.239652f
C2914 vdd.n1921 gnd 0.152078f
C2915 vdd.t245 gnd 0.03487f
C2916 vdd.t182 gnd 0.03487f
C2917 vdd.n1922 gnd 0.239652f
C2918 vdd.n1923 gnd 0.152078f
C2919 vdd.t287 gnd 0.03487f
C2920 vdd.t215 gnd 0.03487f
C2921 vdd.n1924 gnd 0.239652f
C2922 vdd.n1925 gnd 0.152078f
C2923 vdd.t265 gnd 0.03487f
C2924 vdd.t237 gnd 0.03487f
C2925 vdd.n1926 gnd 0.239652f
C2926 vdd.n1927 gnd 0.152078f
C2927 vdd.n1928 gnd 0.005944f
C2928 vdd.n1929 gnd 0.005516f
C2929 vdd.n1930 gnd 0.003051f
C2930 vdd.n1931 gnd 0.007006f
C2931 vdd.n1932 gnd 0.002964f
C2932 vdd.n1933 gnd 0.003138f
C2933 vdd.n1934 gnd 0.005516f
C2934 vdd.n1935 gnd 0.002964f
C2935 vdd.n1936 gnd 0.007006f
C2936 vdd.n1937 gnd 0.003138f
C2937 vdd.n1938 gnd 0.005516f
C2938 vdd.n1939 gnd 0.002964f
C2939 vdd.n1940 gnd 0.005254f
C2940 vdd.n1941 gnd 0.00527f
C2941 vdd.t197 gnd 0.015051f
C2942 vdd.n1942 gnd 0.033489f
C2943 vdd.n1943 gnd 0.174283f
C2944 vdd.n1944 gnd 0.002964f
C2945 vdd.n1945 gnd 0.003138f
C2946 vdd.n1946 gnd 0.007006f
C2947 vdd.n1947 gnd 0.007006f
C2948 vdd.n1948 gnd 0.003138f
C2949 vdd.n1949 gnd 0.002964f
C2950 vdd.n1950 gnd 0.005516f
C2951 vdd.n1951 gnd 0.005516f
C2952 vdd.n1952 gnd 0.002964f
C2953 vdd.n1953 gnd 0.003138f
C2954 vdd.n1954 gnd 0.007006f
C2955 vdd.n1955 gnd 0.007006f
C2956 vdd.n1956 gnd 0.003138f
C2957 vdd.n1957 gnd 0.002964f
C2958 vdd.n1958 gnd 0.005516f
C2959 vdd.n1959 gnd 0.005516f
C2960 vdd.n1960 gnd 0.002964f
C2961 vdd.n1961 gnd 0.003138f
C2962 vdd.n1962 gnd 0.007006f
C2963 vdd.n1963 gnd 0.007006f
C2964 vdd.n1964 gnd 0.016563f
C2965 vdd.n1965 gnd 0.003051f
C2966 vdd.n1966 gnd 0.002964f
C2967 vdd.n1967 gnd 0.014257f
C2968 vdd.n1968 gnd 0.009641f
C2969 vdd.n1969 gnd 0.113146f
C2970 vdd.n1970 gnd 0.005944f
C2971 vdd.n1971 gnd 0.005516f
C2972 vdd.n1972 gnd 0.003051f
C2973 vdd.n1973 gnd 0.007006f
C2974 vdd.n1974 gnd 0.002964f
C2975 vdd.n1975 gnd 0.003138f
C2976 vdd.n1976 gnd 0.005516f
C2977 vdd.n1977 gnd 0.002964f
C2978 vdd.n1978 gnd 0.007006f
C2979 vdd.n1979 gnd 0.003138f
C2980 vdd.n1980 gnd 0.005516f
C2981 vdd.n1981 gnd 0.002964f
C2982 vdd.n1982 gnd 0.005254f
C2983 vdd.n1983 gnd 0.00527f
C2984 vdd.t276 gnd 0.015051f
C2985 vdd.n1984 gnd 0.033489f
C2986 vdd.n1985 gnd 0.174283f
C2987 vdd.n1986 gnd 0.002964f
C2988 vdd.n1987 gnd 0.003138f
C2989 vdd.n1988 gnd 0.007006f
C2990 vdd.n1989 gnd 0.007006f
C2991 vdd.n1990 gnd 0.003138f
C2992 vdd.n1991 gnd 0.002964f
C2993 vdd.n1992 gnd 0.005516f
C2994 vdd.n1993 gnd 0.005516f
C2995 vdd.n1994 gnd 0.002964f
C2996 vdd.n1995 gnd 0.003138f
C2997 vdd.n1996 gnd 0.007006f
C2998 vdd.n1997 gnd 0.007006f
C2999 vdd.n1998 gnd 0.003138f
C3000 vdd.n1999 gnd 0.002964f
C3001 vdd.n2000 gnd 0.005516f
C3002 vdd.n2001 gnd 0.005516f
C3003 vdd.n2002 gnd 0.002964f
C3004 vdd.n2003 gnd 0.003138f
C3005 vdd.n2004 gnd 0.007006f
C3006 vdd.n2005 gnd 0.007006f
C3007 vdd.n2006 gnd 0.016563f
C3008 vdd.n2007 gnd 0.003051f
C3009 vdd.n2008 gnd 0.002964f
C3010 vdd.n2009 gnd 0.014257f
C3011 vdd.n2010 gnd 0.009953f
C3012 vdd.t225 gnd 0.03487f
C3013 vdd.t149 gnd 0.03487f
C3014 vdd.n2011 gnd 0.239652f
C3015 vdd.n2012 gnd 0.188449f
C3016 vdd.t289 gnd 0.03487f
C3017 vdd.t257 gnd 0.03487f
C3018 vdd.n2013 gnd 0.239652f
C3019 vdd.n2014 gnd 0.152078f
C3020 vdd.t251 gnd 0.03487f
C3021 vdd.t190 gnd 0.03487f
C3022 vdd.n2015 gnd 0.239652f
C3023 vdd.n2016 gnd 0.152078f
C3024 vdd.t184 gnd 0.03487f
C3025 vdd.t252 gnd 0.03487f
C3026 vdd.n2017 gnd 0.239652f
C3027 vdd.n2018 gnd 0.152078f
C3028 vdd.t241 gnd 0.03487f
C3029 vdd.t239 gnd 0.03487f
C3030 vdd.n2019 gnd 0.239652f
C3031 vdd.n2020 gnd 0.152078f
C3032 vdd.t180 gnd 0.03487f
C3033 vdd.t155 gnd 0.03487f
C3034 vdd.n2021 gnd 0.239652f
C3035 vdd.n2022 gnd 0.152078f
C3036 vdd.t145 gnd 0.03487f
C3037 vdd.t234 gnd 0.03487f
C3038 vdd.n2023 gnd 0.239652f
C3039 vdd.n2024 gnd 0.152078f
C3040 vdd.t211 gnd 0.03487f
C3041 vdd.t151 gnd 0.03487f
C3042 vdd.n2025 gnd 0.239652f
C3043 vdd.n2026 gnd 0.152078f
C3044 vdd.t141 gnd 0.03487f
C3045 vdd.t258 gnd 0.03487f
C3046 vdd.n2027 gnd 0.239652f
C3047 vdd.n2028 gnd 0.152078f
C3048 vdd.n2029 gnd 0.005944f
C3049 vdd.n2030 gnd 0.005516f
C3050 vdd.n2031 gnd 0.003051f
C3051 vdd.n2032 gnd 0.007006f
C3052 vdd.n2033 gnd 0.002964f
C3053 vdd.n2034 gnd 0.003138f
C3054 vdd.n2035 gnd 0.005516f
C3055 vdd.n2036 gnd 0.002964f
C3056 vdd.n2037 gnd 0.007006f
C3057 vdd.n2038 gnd 0.003138f
C3058 vdd.n2039 gnd 0.005516f
C3059 vdd.n2040 gnd 0.002964f
C3060 vdd.n2041 gnd 0.005254f
C3061 vdd.n2042 gnd 0.00527f
C3062 vdd.t199 gnd 0.015051f
C3063 vdd.n2043 gnd 0.033489f
C3064 vdd.n2044 gnd 0.174283f
C3065 vdd.n2045 gnd 0.002964f
C3066 vdd.n2046 gnd 0.003138f
C3067 vdd.n2047 gnd 0.007006f
C3068 vdd.n2048 gnd 0.007006f
C3069 vdd.n2049 gnd 0.003138f
C3070 vdd.n2050 gnd 0.002964f
C3071 vdd.n2051 gnd 0.005516f
C3072 vdd.n2052 gnd 0.005516f
C3073 vdd.n2053 gnd 0.002964f
C3074 vdd.n2054 gnd 0.003138f
C3075 vdd.n2055 gnd 0.007006f
C3076 vdd.n2056 gnd 0.007006f
C3077 vdd.n2057 gnd 0.003138f
C3078 vdd.n2058 gnd 0.002964f
C3079 vdd.n2059 gnd 0.005516f
C3080 vdd.n2060 gnd 0.005516f
C3081 vdd.n2061 gnd 0.002964f
C3082 vdd.n2062 gnd 0.003138f
C3083 vdd.n2063 gnd 0.007006f
C3084 vdd.n2064 gnd 0.007006f
C3085 vdd.n2065 gnd 0.016563f
C3086 vdd.n2066 gnd 0.003051f
C3087 vdd.n2067 gnd 0.002964f
C3088 vdd.n2068 gnd 0.014257f
C3089 vdd.n2069 gnd 0.009641f
C3090 vdd.n2070 gnd 0.067311f
C3091 vdd.n2071 gnd 0.242538f
C3092 vdd.n2072 gnd 0.005944f
C3093 vdd.n2073 gnd 0.005516f
C3094 vdd.n2074 gnd 0.003051f
C3095 vdd.n2075 gnd 0.007006f
C3096 vdd.n2076 gnd 0.002964f
C3097 vdd.n2077 gnd 0.003138f
C3098 vdd.n2078 gnd 0.005516f
C3099 vdd.n2079 gnd 0.002964f
C3100 vdd.n2080 gnd 0.007006f
C3101 vdd.n2081 gnd 0.003138f
C3102 vdd.n2082 gnd 0.005516f
C3103 vdd.n2083 gnd 0.002964f
C3104 vdd.n2084 gnd 0.005254f
C3105 vdd.n2085 gnd 0.00527f
C3106 vdd.t288 gnd 0.015051f
C3107 vdd.n2086 gnd 0.033489f
C3108 vdd.n2087 gnd 0.174283f
C3109 vdd.n2088 gnd 0.002964f
C3110 vdd.n2089 gnd 0.003138f
C3111 vdd.n2090 gnd 0.007006f
C3112 vdd.n2091 gnd 0.007006f
C3113 vdd.n2092 gnd 0.003138f
C3114 vdd.n2093 gnd 0.002964f
C3115 vdd.n2094 gnd 0.005516f
C3116 vdd.n2095 gnd 0.005516f
C3117 vdd.n2096 gnd 0.002964f
C3118 vdd.n2097 gnd 0.003138f
C3119 vdd.n2098 gnd 0.007006f
C3120 vdd.n2099 gnd 0.007006f
C3121 vdd.n2100 gnd 0.003138f
C3122 vdd.n2101 gnd 0.002964f
C3123 vdd.n2102 gnd 0.005516f
C3124 vdd.n2103 gnd 0.005516f
C3125 vdd.n2104 gnd 0.002964f
C3126 vdd.n2105 gnd 0.003138f
C3127 vdd.n2106 gnd 0.007006f
C3128 vdd.n2107 gnd 0.007006f
C3129 vdd.n2108 gnd 0.016563f
C3130 vdd.n2109 gnd 0.003051f
C3131 vdd.n2110 gnd 0.002964f
C3132 vdd.n2111 gnd 0.014257f
C3133 vdd.n2112 gnd 0.009953f
C3134 vdd.t242 gnd 0.03487f
C3135 vdd.t174 gnd 0.03487f
C3136 vdd.n2113 gnd 0.239652f
C3137 vdd.n2114 gnd 0.188449f
C3138 vdd.t299 gnd 0.03487f
C3139 vdd.t269 gnd 0.03487f
C3140 vdd.n2115 gnd 0.239652f
C3141 vdd.n2116 gnd 0.152078f
C3142 vdd.t267 gnd 0.03487f
C3143 vdd.t216 gnd 0.03487f
C3144 vdd.n2117 gnd 0.239652f
C3145 vdd.n2118 gnd 0.152078f
C3146 vdd.t212 gnd 0.03487f
C3147 vdd.t268 gnd 0.03487f
C3148 vdd.n2119 gnd 0.239652f
C3149 vdd.n2120 gnd 0.152078f
C3150 vdd.t250 gnd 0.03487f
C3151 vdd.t249 gnd 0.03487f
C3152 vdd.n2121 gnd 0.239652f
C3153 vdd.n2122 gnd 0.152078f
C3154 vdd.t207 gnd 0.03487f
C3155 vdd.t176 gnd 0.03487f
C3156 vdd.n2123 gnd 0.239652f
C3157 vdd.n2124 gnd 0.152078f
C3158 vdd.t173 gnd 0.03487f
C3159 vdd.t248 gnd 0.03487f
C3160 vdd.n2125 gnd 0.239652f
C3161 vdd.n2126 gnd 0.152078f
C3162 vdd.t227 gnd 0.03487f
C3163 vdd.t175 gnd 0.03487f
C3164 vdd.n2127 gnd 0.239652f
C3165 vdd.n2128 gnd 0.152078f
C3166 vdd.t166 gnd 0.03487f
C3167 vdd.t270 gnd 0.03487f
C3168 vdd.n2129 gnd 0.239652f
C3169 vdd.n2130 gnd 0.152078f
C3170 vdd.n2131 gnd 0.005944f
C3171 vdd.n2132 gnd 0.005516f
C3172 vdd.n2133 gnd 0.003051f
C3173 vdd.n2134 gnd 0.007006f
C3174 vdd.n2135 gnd 0.002964f
C3175 vdd.n2136 gnd 0.003138f
C3176 vdd.n2137 gnd 0.005516f
C3177 vdd.n2138 gnd 0.002964f
C3178 vdd.n2139 gnd 0.007006f
C3179 vdd.n2140 gnd 0.003138f
C3180 vdd.n2141 gnd 0.005516f
C3181 vdd.n2142 gnd 0.002964f
C3182 vdd.n2143 gnd 0.005254f
C3183 vdd.n2144 gnd 0.00527f
C3184 vdd.t222 gnd 0.015051f
C3185 vdd.n2145 gnd 0.033489f
C3186 vdd.n2146 gnd 0.174283f
C3187 vdd.n2147 gnd 0.002964f
C3188 vdd.n2148 gnd 0.003138f
C3189 vdd.n2149 gnd 0.007006f
C3190 vdd.n2150 gnd 0.007006f
C3191 vdd.n2151 gnd 0.003138f
C3192 vdd.n2152 gnd 0.002964f
C3193 vdd.n2153 gnd 0.005516f
C3194 vdd.n2154 gnd 0.005516f
C3195 vdd.n2155 gnd 0.002964f
C3196 vdd.n2156 gnd 0.003138f
C3197 vdd.n2157 gnd 0.007006f
C3198 vdd.n2158 gnd 0.007006f
C3199 vdd.n2159 gnd 0.003138f
C3200 vdd.n2160 gnd 0.002964f
C3201 vdd.n2161 gnd 0.005516f
C3202 vdd.n2162 gnd 0.005516f
C3203 vdd.n2163 gnd 0.002964f
C3204 vdd.n2164 gnd 0.003138f
C3205 vdd.n2165 gnd 0.007006f
C3206 vdd.n2166 gnd 0.007006f
C3207 vdd.n2167 gnd 0.016563f
C3208 vdd.n2168 gnd 0.003051f
C3209 vdd.n2169 gnd 0.002964f
C3210 vdd.n2170 gnd 0.014257f
C3211 vdd.n2171 gnd 0.009641f
C3212 vdd.n2172 gnd 0.067311f
C3213 vdd.n2173 gnd 0.277654f
C3214 vdd.n2174 gnd 2.91269f
C3215 vdd.n2175 gnd 0.638846f
C3216 vdd.n2176 gnd 0.008324f
C3217 vdd.n2177 gnd 0.008718f
C3218 vdd.n2178 gnd 0.010831f
C3219 vdd.n2179 gnd 0.791407f
C3220 vdd.n2180 gnd 0.010831f
C3221 vdd.n2181 gnd 0.008718f
C3222 vdd.n2182 gnd 0.010831f
C3223 vdd.n2183 gnd 0.010831f
C3224 vdd.n2184 gnd 0.010831f
C3225 vdd.n2185 gnd 0.008718f
C3226 vdd.n2186 gnd 0.010831f
C3227 vdd.n2187 gnd 0.918696f
C3228 vdd.t183 gnd 0.553432f
C3229 vdd.n2188 gnd 0.60324f
C3230 vdd.n2189 gnd 0.010831f
C3231 vdd.n2190 gnd 0.008718f
C3232 vdd.n2191 gnd 0.010831f
C3233 vdd.n2192 gnd 0.010831f
C3234 vdd.n2193 gnd 0.010831f
C3235 vdd.n2194 gnd 0.008718f
C3236 vdd.n2195 gnd 0.010831f
C3237 vdd.n2196 gnd 0.691789f
C3238 vdd.n2197 gnd 0.010831f
C3239 vdd.n2198 gnd 0.008718f
C3240 vdd.n2199 gnd 0.010831f
C3241 vdd.n2200 gnd 0.010831f
C3242 vdd.n2201 gnd 0.010831f
C3243 vdd.n2202 gnd 0.008718f
C3244 vdd.n2203 gnd 0.010831f
C3245 vdd.n2204 gnd 0.592172f
C3246 vdd.n2205 gnd 0.879956f
C3247 vdd.n2206 gnd 0.010831f
C3248 vdd.n2207 gnd 0.008718f
C3249 vdd.n2208 gnd 0.010831f
C3250 vdd.n2209 gnd 0.010831f
C3251 vdd.n2210 gnd 0.010831f
C3252 vdd.n2211 gnd 0.008718f
C3253 vdd.n2212 gnd 0.010831f
C3254 vdd.n2213 gnd 0.918696f
C3255 vdd.n2214 gnd 0.010831f
C3256 vdd.n2215 gnd 0.008718f
C3257 vdd.n2216 gnd 0.010831f
C3258 vdd.n2217 gnd 0.010831f
C3259 vdd.n2218 gnd 0.010831f
C3260 vdd.n2219 gnd 0.008718f
C3261 vdd.n2220 gnd 0.010831f
C3262 vdd.t256 gnd 0.553432f
C3263 vdd.n2221 gnd 0.76927f
C3264 vdd.n2222 gnd 0.010831f
C3265 vdd.n2223 gnd 0.008718f
C3266 vdd.n2224 gnd 0.010831f
C3267 vdd.n2225 gnd 0.010831f
C3268 vdd.n2226 gnd 0.010831f
C3269 vdd.n2227 gnd 0.008718f
C3270 vdd.n2228 gnd 0.010831f
C3271 vdd.n2229 gnd 0.581103f
C3272 vdd.n2230 gnd 0.010831f
C3273 vdd.n2231 gnd 0.008718f
C3274 vdd.n2232 gnd 0.010831f
C3275 vdd.n2233 gnd 0.010831f
C3276 vdd.n2234 gnd 0.010831f
C3277 vdd.n2235 gnd 0.008718f
C3278 vdd.n2236 gnd 0.010831f
C3279 vdd.n2237 gnd 0.758201f
C3280 vdd.n2238 gnd 0.713927f
C3281 vdd.n2239 gnd 0.010831f
C3282 vdd.n2240 gnd 0.008718f
C3283 vdd.n2241 gnd 0.010831f
C3284 vdd.n2242 gnd 0.010831f
C3285 vdd.n2243 gnd 0.010831f
C3286 vdd.n2244 gnd 0.008718f
C3287 vdd.n2245 gnd 0.010831f
C3288 vdd.n2246 gnd 0.902093f
C3289 vdd.n2247 gnd 0.010831f
C3290 vdd.n2248 gnd 0.008718f
C3291 vdd.n2249 gnd 0.010831f
C3292 vdd.n2250 gnd 0.010831f
C3293 vdd.n2251 gnd 0.026201f
C3294 vdd.n2252 gnd 0.010831f
C3295 vdd.n2253 gnd 0.010831f
C3296 vdd.n2254 gnd 0.008718f
C3297 vdd.n2255 gnd 0.010831f
C3298 vdd.n2256 gnd 0.669652f
C3299 vdd.n2257 gnd 1.10686f
C3300 vdd.n2258 gnd 0.010831f
C3301 vdd.n2259 gnd 0.008718f
C3302 vdd.n2260 gnd 0.010831f
C3303 vdd.n2261 gnd 0.010831f
C3304 vdd.n2262 gnd 0.026201f
C3305 vdd.n2263 gnd 0.007236f
C3306 vdd.n2264 gnd 0.026201f
C3307 vdd.n2265 gnd 1.52194f
C3308 vdd.n2266 gnd 0.026201f
C3309 vdd.n2267 gnd 0.026762f
C3310 vdd.n2268 gnd 0.004141f
C3311 vdd.t41 gnd 0.133248f
C3312 vdd.t40 gnd 0.142406f
C3313 vdd.t38 gnd 0.17402f
C3314 vdd.n2269 gnd 0.223069f
C3315 vdd.n2270 gnd 0.187419f
C3316 vdd.n2271 gnd 0.013425f
C3317 vdd.n2272 gnd 0.004577f
C3318 vdd.n2273 gnd 0.009315f
C3319 vdd.n2274 gnd 0.819089f
C3320 vdd.n2276 gnd 0.008718f
C3321 vdd.n2277 gnd 0.008718f
C3322 vdd.n2278 gnd 0.010831f
C3323 vdd.n2280 gnd 0.010831f
C3324 vdd.n2281 gnd 0.010831f
C3325 vdd.n2282 gnd 0.008718f
C3326 vdd.n2283 gnd 0.008718f
C3327 vdd.n2284 gnd 0.008718f
C3328 vdd.n2285 gnd 0.010831f
C3329 vdd.n2287 gnd 0.010831f
C3330 vdd.n2288 gnd 0.010831f
C3331 vdd.n2289 gnd 0.008718f
C3332 vdd.n2290 gnd 0.008718f
C3333 vdd.n2291 gnd 0.008718f
C3334 vdd.n2292 gnd 0.010831f
C3335 vdd.n2294 gnd 0.010831f
C3336 vdd.n2295 gnd 0.010831f
C3337 vdd.n2296 gnd 0.008718f
C3338 vdd.n2297 gnd 0.008718f
C3339 vdd.n2298 gnd 0.008718f
C3340 vdd.n2299 gnd 0.010831f
C3341 vdd.n2301 gnd 0.010831f
C3342 vdd.n2302 gnd 0.010831f
C3343 vdd.n2303 gnd 0.008718f
C3344 vdd.n2304 gnd 0.010831f
C3345 vdd.n2305 gnd 0.010831f
C3346 vdd.n2306 gnd 0.010831f
C3347 vdd.n2307 gnd 0.017784f
C3348 vdd.n2308 gnd 0.005928f
C3349 vdd.n2309 gnd 0.008718f
C3350 vdd.n2310 gnd 0.010831f
C3351 vdd.n2312 gnd 0.010831f
C3352 vdd.n2313 gnd 0.010831f
C3353 vdd.n2314 gnd 0.008718f
C3354 vdd.n2315 gnd 0.008718f
C3355 vdd.n2316 gnd 0.008718f
C3356 vdd.n2317 gnd 0.010831f
C3357 vdd.n2319 gnd 0.010831f
C3358 vdd.n2320 gnd 0.010831f
C3359 vdd.n2321 gnd 0.008718f
C3360 vdd.n2322 gnd 0.008718f
C3361 vdd.n2323 gnd 0.008718f
C3362 vdd.n2324 gnd 0.010831f
C3363 vdd.n2326 gnd 0.010831f
C3364 vdd.n2327 gnd 0.010831f
C3365 vdd.n2328 gnd 0.008718f
C3366 vdd.n2329 gnd 0.008718f
C3367 vdd.n2330 gnd 0.008718f
C3368 vdd.n2331 gnd 0.010831f
C3369 vdd.n2333 gnd 0.010831f
C3370 vdd.n2334 gnd 0.010831f
C3371 vdd.n2335 gnd 0.008718f
C3372 vdd.n2336 gnd 0.008718f
C3373 vdd.n2337 gnd 0.008718f
C3374 vdd.n2338 gnd 0.010831f
C3375 vdd.n2340 gnd 0.010831f
C3376 vdd.n2341 gnd 0.010831f
C3377 vdd.n2342 gnd 0.008718f
C3378 vdd.n2343 gnd 0.010831f
C3379 vdd.n2344 gnd 0.010831f
C3380 vdd.n2345 gnd 0.010831f
C3381 vdd.n2346 gnd 0.017784f
C3382 vdd.n2347 gnd 0.007279f
C3383 vdd.n2348 gnd 0.008718f
C3384 vdd.n2349 gnd 0.010831f
C3385 vdd.n2351 gnd 0.010831f
C3386 vdd.n2352 gnd 0.010831f
C3387 vdd.n2353 gnd 0.008718f
C3388 vdd.n2354 gnd 0.008718f
C3389 vdd.n2355 gnd 0.008718f
C3390 vdd.n2356 gnd 0.010831f
C3391 vdd.n2358 gnd 0.010831f
C3392 vdd.n2359 gnd 0.010831f
C3393 vdd.n2360 gnd 0.008718f
C3394 vdd.n2361 gnd 0.008718f
C3395 vdd.n2362 gnd 0.008718f
C3396 vdd.n2363 gnd 0.010831f
C3397 vdd.n2365 gnd 0.010831f
C3398 vdd.n2366 gnd 0.010831f
C3399 vdd.n2367 gnd 0.008718f
C3400 vdd.n2368 gnd 0.008718f
C3401 vdd.n2369 gnd 0.008718f
C3402 vdd.n2370 gnd 0.010831f
C3403 vdd.n2372 gnd 0.010831f
C3404 vdd.n2373 gnd 0.008718f
C3405 vdd.n2374 gnd 0.008718f
C3406 vdd.n2375 gnd 0.010831f
C3407 vdd.n2377 gnd 0.010831f
C3408 vdd.n2378 gnd 0.010831f
C3409 vdd.n2379 gnd 0.008718f
C3410 vdd.n2380 gnd 0.009315f
C3411 vdd.n2381 gnd 0.819089f
C3412 vdd.n2382 gnd 0.029519f
C3413 vdd.n2383 gnd 0.007365f
C3414 vdd.n2384 gnd 0.007365f
C3415 vdd.n2385 gnd 0.007365f
C3416 vdd.n2386 gnd 0.007365f
C3417 vdd.n2387 gnd 0.007365f
C3418 vdd.n2388 gnd 0.007365f
C3419 vdd.n2389 gnd 0.007365f
C3420 vdd.n2390 gnd 0.007365f
C3421 vdd.n2391 gnd 0.007365f
C3422 vdd.n2392 gnd 0.007365f
C3423 vdd.n2393 gnd 0.007365f
C3424 vdd.n2394 gnd 0.007365f
C3425 vdd.n2395 gnd 0.007365f
C3426 vdd.n2396 gnd 0.007365f
C3427 vdd.n2397 gnd 0.007365f
C3428 vdd.n2398 gnd 0.007365f
C3429 vdd.n2399 gnd 0.007365f
C3430 vdd.n2400 gnd 0.007365f
C3431 vdd.n2401 gnd 0.007365f
C3432 vdd.n2402 gnd 0.007365f
C3433 vdd.n2403 gnd 0.007365f
C3434 vdd.n2404 gnd 0.007365f
C3435 vdd.n2405 gnd 0.007365f
C3436 vdd.n2406 gnd 0.007365f
C3437 vdd.n2407 gnd 0.007365f
C3438 vdd.n2408 gnd 0.007365f
C3439 vdd.n2409 gnd 0.007365f
C3440 vdd.n2410 gnd 0.007365f
C3441 vdd.n2411 gnd 0.007365f
C3442 vdd.n2412 gnd 0.007365f
C3443 vdd.n2413 gnd 0.007365f
C3444 vdd.n2414 gnd 0.017226f
C3445 vdd.n2415 gnd 0.017226f
C3446 vdd.n2417 gnd 9.44154f
C3447 vdd.n2419 gnd 0.017226f
C3448 vdd.n2420 gnd 0.017226f
C3449 vdd.n2421 gnd 0.016133f
C3450 vdd.n2422 gnd 0.007365f
C3451 vdd.n2423 gnd 0.007365f
C3452 vdd.n2424 gnd 0.752667f
C3453 vdd.n2425 gnd 0.007365f
C3454 vdd.n2426 gnd 0.007365f
C3455 vdd.n2427 gnd 0.007365f
C3456 vdd.n2428 gnd 0.007365f
C3457 vdd.n2429 gnd 0.007365f
C3458 vdd.n2430 gnd 0.636446f
C3459 vdd.n2431 gnd 0.007365f
C3460 vdd.n2432 gnd 0.007365f
C3461 vdd.n2433 gnd 0.007365f
C3462 vdd.n2434 gnd 0.007365f
C3463 vdd.n2435 gnd 0.007365f
C3464 vdd.n2436 gnd 0.752667f
C3465 vdd.n2437 gnd 0.007365f
C3466 vdd.n2438 gnd 0.007365f
C3467 vdd.n2439 gnd 0.007365f
C3468 vdd.n2440 gnd 0.007365f
C3469 vdd.n2441 gnd 0.007365f
C3470 vdd.n2442 gnd 0.736064f
C3471 vdd.n2443 gnd 0.007365f
C3472 vdd.n2444 gnd 0.007365f
C3473 vdd.n2445 gnd 0.007365f
C3474 vdd.n2446 gnd 0.007365f
C3475 vdd.n2447 gnd 0.007365f
C3476 vdd.n2448 gnd 0.752667f
C3477 vdd.n2449 gnd 0.007365f
C3478 vdd.n2450 gnd 0.007365f
C3479 vdd.n2451 gnd 0.007365f
C3480 vdd.n2452 gnd 0.007365f
C3481 vdd.n2453 gnd 0.007365f
C3482 vdd.n2454 gnd 0.60324f
C3483 vdd.n2455 gnd 0.007365f
C3484 vdd.n2456 gnd 0.007365f
C3485 vdd.n2457 gnd 0.006282f
C3486 vdd.n2458 gnd 0.021336f
C3487 vdd.n2459 gnd 0.004766f
C3488 vdd.n2460 gnd 0.007365f
C3489 vdd.n2461 gnd 0.437211f
C3490 vdd.n2462 gnd 0.007365f
C3491 vdd.n2463 gnd 0.007365f
C3492 vdd.n2464 gnd 0.007365f
C3493 vdd.n2465 gnd 0.007365f
C3494 vdd.n2466 gnd 0.007365f
C3495 vdd.n2467 gnd 0.481485f
C3496 vdd.n2468 gnd 0.007365f
C3497 vdd.n2469 gnd 0.007365f
C3498 vdd.n2470 gnd 0.007365f
C3499 vdd.n2471 gnd 0.007365f
C3500 vdd.n2472 gnd 0.007365f
C3501 vdd.n2473 gnd 0.647515f
C3502 vdd.n2474 gnd 0.007365f
C3503 vdd.n2475 gnd 0.007365f
C3504 vdd.n2476 gnd 0.007365f
C3505 vdd.n2477 gnd 0.007365f
C3506 vdd.n2478 gnd 0.007365f
C3507 vdd.n2479 gnd 0.619843f
C3508 vdd.n2480 gnd 0.007365f
C3509 vdd.n2481 gnd 0.007365f
C3510 vdd.n2482 gnd 0.007365f
C3511 vdd.n2483 gnd 0.007365f
C3512 vdd.n2484 gnd 0.007365f
C3513 vdd.n2485 gnd 0.453814f
C3514 vdd.n2486 gnd 0.007365f
C3515 vdd.n2487 gnd 0.007365f
C3516 vdd.n2488 gnd 0.007365f
C3517 vdd.n2489 gnd 0.007365f
C3518 vdd.n2490 gnd 0.007365f
C3519 vdd.n2491 gnd 0.237976f
C3520 vdd.n2492 gnd 0.007365f
C3521 vdd.n2493 gnd 0.007365f
C3522 vdd.n2494 gnd 0.007365f
C3523 vdd.n2495 gnd 0.007365f
C3524 vdd.n2496 gnd 0.007365f
C3525 vdd.n2497 gnd 0.392936f
C3526 vdd.n2498 gnd 0.007365f
C3527 vdd.n2499 gnd 0.007365f
C3528 vdd.n2500 gnd 0.007365f
C3529 vdd.n2501 gnd 0.007365f
C3530 vdd.n2502 gnd 0.007365f
C3531 vdd.n2503 gnd 0.752667f
C3532 vdd.n2504 gnd 0.007365f
C3533 vdd.n2505 gnd 0.007365f
C3534 vdd.n2506 gnd 0.007365f
C3535 vdd.n2507 gnd 0.007365f
C3536 vdd.n2508 gnd 0.007365f
C3537 vdd.n2509 gnd 0.007365f
C3538 vdd.n2510 gnd 0.007365f
C3539 vdd.n2511 gnd 0.5645f
C3540 vdd.n2512 gnd 0.007365f
C3541 vdd.n2513 gnd 0.007365f
C3542 vdd.n2514 gnd 0.007365f
C3543 vdd.n2515 gnd 0.007365f
C3544 vdd.n2516 gnd 0.007365f
C3545 vdd.n2517 gnd 0.007365f
C3546 vdd.n2518 gnd 0.470417f
C3547 vdd.n2519 gnd 0.007365f
C3548 vdd.n2520 gnd 0.007365f
C3549 vdd.n2521 gnd 0.007365f
C3550 vdd.n2522 gnd 0.017048f
C3551 vdd.n2523 gnd 0.016311f
C3552 vdd.n2524 gnd 0.007365f
C3553 vdd.n2525 gnd 0.007365f
C3554 vdd.n2526 gnd 0.005686f
C3555 vdd.n2527 gnd 0.007365f
C3556 vdd.n2528 gnd 0.007365f
C3557 vdd.n2529 gnd 0.005361f
C3558 vdd.n2530 gnd 0.007365f
C3559 vdd.n2531 gnd 0.007365f
C3560 vdd.n2532 gnd 0.007365f
C3561 vdd.n2533 gnd 0.007365f
C3562 vdd.n2534 gnd 0.007365f
C3563 vdd.n2535 gnd 0.007365f
C3564 vdd.n2536 gnd 0.007365f
C3565 vdd.n2537 gnd 0.007365f
C3566 vdd.n2538 gnd 0.007365f
C3567 vdd.n2539 gnd 0.007365f
C3568 vdd.n2540 gnd 0.007365f
C3569 vdd.n2541 gnd 0.007365f
C3570 vdd.n2542 gnd 0.007365f
C3571 vdd.n2543 gnd 0.007365f
C3572 vdd.n2544 gnd 0.007365f
C3573 vdd.n2545 gnd 0.007365f
C3574 vdd.n2546 gnd 0.007365f
C3575 vdd.n2547 gnd 0.007365f
C3576 vdd.n2548 gnd 0.007365f
C3577 vdd.n2549 gnd 0.007365f
C3578 vdd.n2550 gnd 0.007365f
C3579 vdd.n2551 gnd 0.007365f
C3580 vdd.n2552 gnd 0.007365f
C3581 vdd.n2553 gnd 0.007365f
C3582 vdd.n2554 gnd 0.007365f
C3583 vdd.n2555 gnd 0.007365f
C3584 vdd.n2556 gnd 0.007365f
C3585 vdd.n2557 gnd 0.007365f
C3586 vdd.n2558 gnd 0.007365f
C3587 vdd.n2559 gnd 0.007365f
C3588 vdd.n2560 gnd 0.007365f
C3589 vdd.n2561 gnd 0.007365f
C3590 vdd.n2562 gnd 0.007365f
C3591 vdd.n2563 gnd 0.007365f
C3592 vdd.n2564 gnd 0.007365f
C3593 vdd.n2565 gnd 0.007365f
C3594 vdd.n2566 gnd 0.007365f
C3595 vdd.n2567 gnd 0.007365f
C3596 vdd.n2568 gnd 0.007365f
C3597 vdd.n2569 gnd 0.007365f
C3598 vdd.n2570 gnd 0.007365f
C3599 vdd.n2571 gnd 0.007365f
C3600 vdd.n2572 gnd 0.007365f
C3601 vdd.n2573 gnd 0.007365f
C3602 vdd.n2574 gnd 0.007365f
C3603 vdd.n2575 gnd 0.007365f
C3604 vdd.n2576 gnd 0.007365f
C3605 vdd.n2577 gnd 0.007365f
C3606 vdd.n2578 gnd 0.007365f
C3607 vdd.n2579 gnd 0.007365f
C3608 vdd.n2580 gnd 0.007365f
C3609 vdd.n2581 gnd 0.007365f
C3610 vdd.n2582 gnd 0.007365f
C3611 vdd.n2583 gnd 0.007365f
C3612 vdd.n2584 gnd 0.007365f
C3613 vdd.n2585 gnd 0.007365f
C3614 vdd.n2586 gnd 0.007365f
C3615 vdd.n2587 gnd 0.007365f
C3616 vdd.n2588 gnd 0.007365f
C3617 vdd.n2589 gnd 0.007365f
C3618 vdd.n2590 gnd 0.017226f
C3619 vdd.n2591 gnd 0.016133f
C3620 vdd.n2592 gnd 0.016133f
C3621 vdd.n2593 gnd 0.896559f
C3622 vdd.n2594 gnd 0.016133f
C3623 vdd.n2595 gnd 0.017226f
C3624 vdd.n2596 gnd 0.016311f
C3625 vdd.n2597 gnd 0.007365f
C3626 vdd.n2598 gnd 0.007365f
C3627 vdd.n2599 gnd 0.007365f
C3628 vdd.n2600 gnd 0.005686f
C3629 vdd.n2601 gnd 0.010526f
C3630 vdd.n2602 gnd 0.005361f
C3631 vdd.n2603 gnd 0.007365f
C3632 vdd.n2604 gnd 0.007365f
C3633 vdd.n2605 gnd 0.007365f
C3634 vdd.n2606 gnd 0.007365f
C3635 vdd.n2607 gnd 0.007365f
C3636 vdd.n2608 gnd 0.007365f
C3637 vdd.n2609 gnd 0.007365f
C3638 vdd.n2610 gnd 0.007365f
C3639 vdd.n2611 gnd 0.007365f
C3640 vdd.n2612 gnd 0.007365f
C3641 vdd.n2613 gnd 0.007365f
C3642 vdd.n2614 gnd 0.007365f
C3643 vdd.n2615 gnd 0.007365f
C3644 vdd.n2616 gnd 0.007365f
C3645 vdd.n2617 gnd 0.007365f
C3646 vdd.n2618 gnd 0.007365f
C3647 vdd.n2619 gnd 0.007365f
C3648 vdd.n2620 gnd 0.007365f
C3649 vdd.n2621 gnd 0.007365f
C3650 vdd.n2622 gnd 0.007365f
C3651 vdd.n2623 gnd 0.007365f
C3652 vdd.n2624 gnd 0.007365f
C3653 vdd.n2625 gnd 0.007365f
C3654 vdd.n2626 gnd 0.007365f
C3655 vdd.n2627 gnd 0.007365f
C3656 vdd.n2628 gnd 0.007365f
C3657 vdd.n2629 gnd 0.007365f
C3658 vdd.n2630 gnd 0.007365f
C3659 vdd.n2631 gnd 0.007365f
C3660 vdd.n2632 gnd 0.007365f
C3661 vdd.n2633 gnd 0.007365f
C3662 vdd.n2634 gnd 0.007365f
C3663 vdd.n2635 gnd 0.007365f
C3664 vdd.n2636 gnd 0.007365f
C3665 vdd.n2637 gnd 0.007365f
C3666 vdd.n2638 gnd 0.007365f
C3667 vdd.n2639 gnd 0.007365f
C3668 vdd.n2640 gnd 0.007365f
C3669 vdd.n2641 gnd 0.007365f
C3670 vdd.n2642 gnd 0.007365f
C3671 vdd.n2643 gnd 0.007365f
C3672 vdd.n2644 gnd 0.007365f
C3673 vdd.n2645 gnd 0.007365f
C3674 vdd.n2646 gnd 0.007365f
C3675 vdd.n2647 gnd 0.007365f
C3676 vdd.n2648 gnd 0.007365f
C3677 vdd.n2649 gnd 0.007365f
C3678 vdd.n2650 gnd 0.007365f
C3679 vdd.n2651 gnd 0.007365f
C3680 vdd.n2652 gnd 0.007365f
C3681 vdd.n2653 gnd 0.007365f
C3682 vdd.n2654 gnd 0.007365f
C3683 vdd.n2655 gnd 0.007365f
C3684 vdd.n2656 gnd 0.007365f
C3685 vdd.n2657 gnd 0.007365f
C3686 vdd.n2658 gnd 0.007365f
C3687 vdd.n2659 gnd 0.007365f
C3688 vdd.n2660 gnd 0.007365f
C3689 vdd.n2661 gnd 0.007365f
C3690 vdd.n2662 gnd 0.007365f
C3691 vdd.n2663 gnd 0.017226f
C3692 vdd.n2664 gnd 0.017226f
C3693 vdd.n2665 gnd 0.918696f
C3694 vdd.t136 gnd 3.26525f
C3695 vdd.t130 gnd 3.26525f
C3696 vdd.n2698 gnd 0.017226f
C3697 vdd.t102 gnd 0.686255f
C3698 vdd.n2699 gnd 0.007365f
C3699 vdd.n2700 gnd 0.007365f
C3700 vdd.t78 gnd 0.297618f
C3701 vdd.t79 gnd 0.304649f
C3702 vdd.t76 gnd 0.194297f
C3703 vdd.n2701 gnd 0.105007f
C3704 vdd.n2702 gnd 0.059563f
C3705 vdd.n2703 gnd 0.007365f
C3706 vdd.t88 gnd 0.297618f
C3707 vdd.t89 gnd 0.304649f
C3708 vdd.t87 gnd 0.194297f
C3709 vdd.n2704 gnd 0.105007f
C3710 vdd.n2705 gnd 0.059563f
C3711 vdd.n2706 gnd 0.010526f
C3712 vdd.n2707 gnd 0.007365f
C3713 vdd.n2708 gnd 0.007365f
C3714 vdd.n2709 gnd 0.007365f
C3715 vdd.n2710 gnd 0.007365f
C3716 vdd.n2711 gnd 0.007365f
C3717 vdd.n2712 gnd 0.007365f
C3718 vdd.n2713 gnd 0.007365f
C3719 vdd.n2714 gnd 0.007365f
C3720 vdd.n2715 gnd 0.007365f
C3721 vdd.n2716 gnd 0.007365f
C3722 vdd.n2717 gnd 0.007365f
C3723 vdd.n2718 gnd 0.007365f
C3724 vdd.n2719 gnd 0.007365f
C3725 vdd.n2720 gnd 0.007365f
C3726 vdd.n2721 gnd 0.007365f
C3727 vdd.n2722 gnd 0.007365f
C3728 vdd.n2723 gnd 0.007365f
C3729 vdd.n2724 gnd 0.007365f
C3730 vdd.n2725 gnd 0.007365f
C3731 vdd.n2726 gnd 0.007365f
C3732 vdd.n2727 gnd 0.007365f
C3733 vdd.n2728 gnd 0.007365f
C3734 vdd.n2729 gnd 0.007365f
C3735 vdd.n2730 gnd 0.007365f
C3736 vdd.n2731 gnd 0.007365f
C3737 vdd.n2732 gnd 0.007365f
C3738 vdd.n2733 gnd 0.007365f
C3739 vdd.n2734 gnd 0.007365f
C3740 vdd.n2735 gnd 0.007365f
C3741 vdd.n2736 gnd 0.007365f
C3742 vdd.n2737 gnd 0.007365f
C3743 vdd.n2738 gnd 0.007365f
C3744 vdd.n2739 gnd 0.007365f
C3745 vdd.n2740 gnd 0.007365f
C3746 vdd.n2741 gnd 0.007365f
C3747 vdd.n2742 gnd 0.007365f
C3748 vdd.n2743 gnd 0.007365f
C3749 vdd.n2744 gnd 0.007365f
C3750 vdd.n2745 gnd 0.007365f
C3751 vdd.n2746 gnd 0.007365f
C3752 vdd.n2747 gnd 0.007365f
C3753 vdd.n2748 gnd 0.007365f
C3754 vdd.n2749 gnd 0.007365f
C3755 vdd.n2750 gnd 0.007365f
C3756 vdd.n2751 gnd 0.007365f
C3757 vdd.n2752 gnd 0.007365f
C3758 vdd.n2753 gnd 0.007365f
C3759 vdd.n2754 gnd 0.007365f
C3760 vdd.n2755 gnd 0.007365f
C3761 vdd.n2756 gnd 0.007365f
C3762 vdd.n2757 gnd 0.007365f
C3763 vdd.n2758 gnd 0.007365f
C3764 vdd.n2759 gnd 0.007365f
C3765 vdd.n2760 gnd 0.007365f
C3766 vdd.n2761 gnd 0.007365f
C3767 vdd.n2762 gnd 0.007365f
C3768 vdd.n2763 gnd 0.007365f
C3769 vdd.n2764 gnd 0.007365f
C3770 vdd.n2765 gnd 0.005361f
C3771 vdd.n2766 gnd 0.007365f
C3772 vdd.n2767 gnd 0.007365f
C3773 vdd.n2768 gnd 0.005686f
C3774 vdd.n2769 gnd 0.007365f
C3775 vdd.n2770 gnd 0.007365f
C3776 vdd.n2771 gnd 0.017226f
C3777 vdd.n2772 gnd 0.016133f
C3778 vdd.n2773 gnd 0.016133f
C3779 vdd.n2774 gnd 0.007365f
C3780 vdd.n2775 gnd 0.007365f
C3781 vdd.n2776 gnd 0.007365f
C3782 vdd.n2777 gnd 0.007365f
C3783 vdd.n2778 gnd 0.007365f
C3784 vdd.n2779 gnd 0.007365f
C3785 vdd.n2780 gnd 0.007365f
C3786 vdd.n2781 gnd 0.007365f
C3787 vdd.n2782 gnd 0.007365f
C3788 vdd.n2783 gnd 0.007365f
C3789 vdd.n2784 gnd 0.007365f
C3790 vdd.n2785 gnd 0.007365f
C3791 vdd.n2786 gnd 0.007365f
C3792 vdd.n2787 gnd 0.007365f
C3793 vdd.n2788 gnd 0.007365f
C3794 vdd.n2789 gnd 0.007365f
C3795 vdd.n2790 gnd 0.007365f
C3796 vdd.n2791 gnd 0.007365f
C3797 vdd.n2792 gnd 0.007365f
C3798 vdd.n2793 gnd 0.007365f
C3799 vdd.n2794 gnd 0.007365f
C3800 vdd.n2795 gnd 0.007365f
C3801 vdd.n2796 gnd 0.007365f
C3802 vdd.n2797 gnd 0.007365f
C3803 vdd.n2798 gnd 0.007365f
C3804 vdd.n2799 gnd 0.007365f
C3805 vdd.n2800 gnd 0.007365f
C3806 vdd.n2801 gnd 0.007365f
C3807 vdd.n2802 gnd 0.007365f
C3808 vdd.n2803 gnd 0.007365f
C3809 vdd.n2804 gnd 0.007365f
C3810 vdd.n2805 gnd 0.007365f
C3811 vdd.n2806 gnd 0.007365f
C3812 vdd.n2807 gnd 0.007365f
C3813 vdd.n2808 gnd 0.007365f
C3814 vdd.n2809 gnd 0.007365f
C3815 vdd.n2810 gnd 0.007365f
C3816 vdd.n2811 gnd 0.007365f
C3817 vdd.n2812 gnd 0.007365f
C3818 vdd.n2813 gnd 0.007365f
C3819 vdd.n2814 gnd 0.007365f
C3820 vdd.n2815 gnd 0.007365f
C3821 vdd.n2816 gnd 0.007365f
C3822 vdd.n2817 gnd 0.007365f
C3823 vdd.n2818 gnd 0.007365f
C3824 vdd.n2819 gnd 0.007365f
C3825 vdd.n2820 gnd 0.007365f
C3826 vdd.n2821 gnd 0.007365f
C3827 vdd.n2822 gnd 0.007365f
C3828 vdd.n2823 gnd 0.007365f
C3829 vdd.n2824 gnd 0.007365f
C3830 vdd.n2825 gnd 0.007365f
C3831 vdd.n2826 gnd 0.007365f
C3832 vdd.n2827 gnd 0.007365f
C3833 vdd.n2828 gnd 0.007365f
C3834 vdd.n2829 gnd 0.007365f
C3835 vdd.n2830 gnd 0.007365f
C3836 vdd.n2831 gnd 0.007365f
C3837 vdd.n2832 gnd 0.007365f
C3838 vdd.n2833 gnd 0.007365f
C3839 vdd.n2834 gnd 0.007365f
C3840 vdd.n2835 gnd 0.007365f
C3841 vdd.n2836 gnd 0.007365f
C3842 vdd.n2837 gnd 0.007365f
C3843 vdd.n2838 gnd 0.007365f
C3844 vdd.n2839 gnd 0.007365f
C3845 vdd.n2840 gnd 0.007365f
C3846 vdd.n2841 gnd 0.007365f
C3847 vdd.n2842 gnd 0.007365f
C3848 vdd.n2843 gnd 0.007365f
C3849 vdd.n2844 gnd 0.007365f
C3850 vdd.n2845 gnd 0.007365f
C3851 vdd.n2846 gnd 0.007365f
C3852 vdd.n2847 gnd 0.237976f
C3853 vdd.n2848 gnd 0.007365f
C3854 vdd.n2849 gnd 0.007365f
C3855 vdd.n2850 gnd 0.007365f
C3856 vdd.n2851 gnd 0.007365f
C3857 vdd.n2852 gnd 0.007365f
C3858 vdd.n2853 gnd 0.007365f
C3859 vdd.n2854 gnd 0.007365f
C3860 vdd.n2855 gnd 0.007365f
C3861 vdd.n2856 gnd 0.007365f
C3862 vdd.n2857 gnd 0.007365f
C3863 vdd.n2858 gnd 0.007365f
C3864 vdd.n2859 gnd 0.007365f
C3865 vdd.n2860 gnd 0.007365f
C3866 vdd.n2861 gnd 0.007365f
C3867 vdd.n2862 gnd 0.470417f
C3868 vdd.n2863 gnd 0.007365f
C3869 vdd.n2864 gnd 0.007365f
C3870 vdd.n2865 gnd 0.007365f
C3871 vdd.n2866 gnd 0.016133f
C3872 vdd.n2867 gnd 0.016133f
C3873 vdd.n2868 gnd 0.017226f
C3874 vdd.n2869 gnd 0.017226f
C3875 vdd.n2870 gnd 0.007365f
C3876 vdd.n2871 gnd 0.007365f
C3877 vdd.n2872 gnd 0.007365f
C3878 vdd.n2873 gnd 0.005686f
C3879 vdd.n2874 gnd 0.010526f
C3880 vdd.n2875 gnd 0.005361f
C3881 vdd.n2876 gnd 0.007365f
C3882 vdd.n2877 gnd 0.007365f
C3883 vdd.n2878 gnd 0.007365f
C3884 vdd.n2879 gnd 0.007365f
C3885 vdd.n2880 gnd 0.007365f
C3886 vdd.n2881 gnd 0.007365f
C3887 vdd.n2882 gnd 0.007365f
C3888 vdd.n2883 gnd 0.007365f
C3889 vdd.n2884 gnd 0.007365f
C3890 vdd.n2885 gnd 0.007365f
C3891 vdd.n2886 gnd 0.007365f
C3892 vdd.n2887 gnd 0.007365f
C3893 vdd.n2888 gnd 0.007365f
C3894 vdd.n2889 gnd 0.007365f
C3895 vdd.n2890 gnd 0.007365f
C3896 vdd.n2891 gnd 0.007365f
C3897 vdd.n2892 gnd 0.007365f
C3898 vdd.n2893 gnd 0.007365f
C3899 vdd.n2894 gnd 0.007365f
C3900 vdd.n2895 gnd 0.007365f
C3901 vdd.n2896 gnd 0.007365f
C3902 vdd.n2897 gnd 0.007365f
C3903 vdd.n2898 gnd 0.007365f
C3904 vdd.n2899 gnd 0.007365f
C3905 vdd.n2900 gnd 0.007365f
C3906 vdd.n2901 gnd 0.007365f
C3907 vdd.n2902 gnd 0.007365f
C3908 vdd.n2903 gnd 0.007365f
C3909 vdd.n2904 gnd 0.007365f
C3910 vdd.n2905 gnd 0.007365f
C3911 vdd.n2906 gnd 0.007365f
C3912 vdd.n2907 gnd 0.007365f
C3913 vdd.n2908 gnd 0.007365f
C3914 vdd.n2909 gnd 0.007365f
C3915 vdd.n2910 gnd 0.007365f
C3916 vdd.n2911 gnd 0.007365f
C3917 vdd.n2912 gnd 0.007365f
C3918 vdd.n2913 gnd 0.007365f
C3919 vdd.n2914 gnd 0.007365f
C3920 vdd.n2915 gnd 0.007365f
C3921 vdd.n2916 gnd 0.007365f
C3922 vdd.n2917 gnd 0.007365f
C3923 vdd.n2918 gnd 0.007365f
C3924 vdd.n2919 gnd 0.007365f
C3925 vdd.n2920 gnd 0.007365f
C3926 vdd.n2921 gnd 0.007365f
C3927 vdd.n2922 gnd 0.007365f
C3928 vdd.n2923 gnd 0.007365f
C3929 vdd.n2924 gnd 0.007365f
C3930 vdd.n2925 gnd 0.007365f
C3931 vdd.n2926 gnd 0.007365f
C3932 vdd.n2927 gnd 0.007365f
C3933 vdd.n2928 gnd 0.007365f
C3934 vdd.n2929 gnd 0.007365f
C3935 vdd.n2930 gnd 0.007365f
C3936 vdd.n2931 gnd 0.007365f
C3937 vdd.n2932 gnd 0.007365f
C3938 vdd.n2933 gnd 0.007365f
C3939 vdd.n2934 gnd 0.007365f
C3940 vdd.n2935 gnd 0.017226f
C3941 vdd.n2936 gnd 0.017226f
C3942 vdd.n2938 gnd 0.918696f
C3943 vdd.n2940 gnd 0.017226f
C3944 vdd.n2941 gnd 0.017226f
C3945 vdd.n2942 gnd 0.016133f
C3946 vdd.n2943 gnd 0.007365f
C3947 vdd.n2944 gnd 0.007365f
C3948 vdd.n2945 gnd 0.398471f
C3949 vdd.n2946 gnd 0.007365f
C3950 vdd.n2947 gnd 0.007365f
C3951 vdd.n2948 gnd 0.007365f
C3952 vdd.n2949 gnd 0.007365f
C3953 vdd.n2950 gnd 0.007365f
C3954 vdd.n2951 gnd 0.44828f
C3955 vdd.n2952 gnd 0.007365f
C3956 vdd.n2953 gnd 0.007365f
C3957 vdd.n2954 gnd 0.007365f
C3958 vdd.n2955 gnd 0.007365f
C3959 vdd.n2956 gnd 0.007365f
C3960 vdd.n2957 gnd 0.752667f
C3961 vdd.n2958 gnd 0.007365f
C3962 vdd.n2959 gnd 0.007365f
C3963 vdd.n2960 gnd 0.007365f
C3964 vdd.n2961 gnd 0.007365f
C3965 vdd.n2962 gnd 0.007365f
C3966 vdd.n2963 gnd 0.498088f
C3967 vdd.n2964 gnd 0.007365f
C3968 vdd.n2965 gnd 0.007365f
C3969 vdd.n2966 gnd 0.007365f
C3970 vdd.n2967 gnd 0.007365f
C3971 vdd.n2968 gnd 0.007365f
C3972 vdd.n2969 gnd 0.664118f
C3973 vdd.n2970 gnd 0.007365f
C3974 vdd.n2971 gnd 0.007365f
C3975 vdd.n2972 gnd 0.007365f
C3976 vdd.n2973 gnd 0.007365f
C3977 vdd.n2974 gnd 0.007365f
C3978 vdd.n2975 gnd 0.60324f
C3979 vdd.n2976 gnd 0.007365f
C3980 vdd.n2977 gnd 0.007365f
C3981 vdd.n2978 gnd 0.007365f
C3982 vdd.n2979 gnd 0.007365f
C3983 vdd.n2980 gnd 0.007365f
C3984 vdd.n2981 gnd 0.437211f
C3985 vdd.n2982 gnd 0.007365f
C3986 vdd.n2983 gnd 0.007365f
C3987 vdd.n2984 gnd 0.007365f
C3988 vdd.n2985 gnd 0.007365f
C3989 vdd.n2986 gnd 0.007365f
C3990 vdd.n2987 gnd 0.237976f
C3991 vdd.n2988 gnd 0.007365f
C3992 vdd.n2989 gnd 0.007365f
C3993 vdd.n2990 gnd 0.007365f
C3994 vdd.n2991 gnd 0.007365f
C3995 vdd.n2992 gnd 0.007365f
C3996 vdd.n2993 gnd 0.647515f
C3997 vdd.n2994 gnd 0.007365f
C3998 vdd.n2995 gnd 0.007365f
C3999 vdd.n2996 gnd 0.007365f
C4000 vdd.n2997 gnd 0.007365f
C4001 vdd.n2998 gnd 0.007365f
C4002 vdd.n2999 gnd 0.752667f
C4003 vdd.n3000 gnd 0.007365f
C4004 vdd.n3001 gnd 0.007365f
C4005 vdd.n3002 gnd 0.004766f
C4006 vdd.n3003 gnd 0.021336f
C4007 vdd.n3004 gnd 0.006282f
C4008 vdd.n3005 gnd 0.007365f
C4009 vdd.n3006 gnd 0.641981f
C4010 vdd.n3007 gnd 0.007365f
C4011 vdd.n3008 gnd 0.007365f
C4012 vdd.n3009 gnd 0.007365f
C4013 vdd.n3010 gnd 0.007365f
C4014 vdd.n3011 gnd 0.007365f
C4015 vdd.n3012 gnd 0.52576f
C4016 vdd.n3013 gnd 0.007365f
C4017 vdd.n3014 gnd 0.007365f
C4018 vdd.n3015 gnd 0.007365f
C4019 vdd.n3016 gnd 0.007365f
C4020 vdd.n3017 gnd 0.007365f
C4021 vdd.n3018 gnd 0.392936f
C4022 vdd.n3019 gnd 0.007365f
C4023 vdd.n3020 gnd 0.007365f
C4024 vdd.n3021 gnd 0.007365f
C4025 vdd.n3022 gnd 0.007365f
C4026 vdd.n3023 gnd 0.007365f
C4027 vdd.n3024 gnd 0.752667f
C4028 vdd.n3025 gnd 0.007365f
C4029 vdd.n3026 gnd 0.007365f
C4030 vdd.n3027 gnd 0.007365f
C4031 vdd.n3028 gnd 0.007365f
C4032 vdd.n3029 gnd 0.007365f
C4033 vdd.n3030 gnd 0.007365f
C4034 vdd.n3032 gnd 0.007365f
C4035 vdd.n3033 gnd 0.007365f
C4036 vdd.n3035 gnd 0.007365f
C4037 vdd.n3036 gnd 0.007365f
C4038 vdd.n3039 gnd 0.007365f
C4039 vdd.n3040 gnd 0.007365f
C4040 vdd.n3041 gnd 0.007365f
C4041 vdd.n3042 gnd 0.007365f
C4042 vdd.n3044 gnd 0.007365f
C4043 vdd.n3045 gnd 0.007365f
C4044 vdd.n3046 gnd 0.007365f
C4045 vdd.n3047 gnd 0.007365f
C4046 vdd.n3048 gnd 0.007365f
C4047 vdd.n3049 gnd 0.007365f
C4048 vdd.n3051 gnd 0.007365f
C4049 vdd.n3052 gnd 0.007365f
C4050 vdd.n3053 gnd 0.007365f
C4051 vdd.n3054 gnd 0.007365f
C4052 vdd.n3055 gnd 0.007365f
C4053 vdd.n3056 gnd 0.007365f
C4054 vdd.n3058 gnd 0.007365f
C4055 vdd.n3059 gnd 0.007365f
C4056 vdd.n3060 gnd 0.007365f
C4057 vdd.n3061 gnd 0.007365f
C4058 vdd.n3062 gnd 0.007365f
C4059 vdd.n3063 gnd 0.007365f
C4060 vdd.n3065 gnd 0.007365f
C4061 vdd.n3066 gnd 0.017226f
C4062 vdd.n3067 gnd 0.017226f
C4063 vdd.n3068 gnd 0.016133f
C4064 vdd.n3069 gnd 0.007365f
C4065 vdd.n3070 gnd 0.007365f
C4066 vdd.n3071 gnd 0.007365f
C4067 vdd.n3072 gnd 0.007365f
C4068 vdd.n3073 gnd 0.007365f
C4069 vdd.n3074 gnd 0.007365f
C4070 vdd.n3075 gnd 0.752667f
C4071 vdd.n3076 gnd 0.007365f
C4072 vdd.n3077 gnd 0.007365f
C4073 vdd.n3078 gnd 0.007365f
C4074 vdd.n3079 gnd 0.007365f
C4075 vdd.n3080 gnd 0.007365f
C4076 vdd.n3081 gnd 0.492554f
C4077 vdd.n3082 gnd 0.007365f
C4078 vdd.n3083 gnd 0.007365f
C4079 vdd.n3084 gnd 0.007365f
C4080 vdd.n3085 gnd 0.017048f
C4081 vdd.n3086 gnd 0.016311f
C4082 vdd.n3087 gnd 0.017226f
C4083 vdd.n3089 gnd 0.007365f
C4084 vdd.n3090 gnd 0.007365f
C4085 vdd.n3091 gnd 0.005686f
C4086 vdd.n3092 gnd 0.010526f
C4087 vdd.n3093 gnd 0.005361f
C4088 vdd.n3094 gnd 0.007365f
C4089 vdd.n3095 gnd 0.007365f
C4090 vdd.n3097 gnd 0.007365f
C4091 vdd.n3098 gnd 0.007365f
C4092 vdd.n3099 gnd 0.007365f
C4093 vdd.n3100 gnd 0.007365f
C4094 vdd.n3101 gnd 0.007365f
C4095 vdd.n3102 gnd 0.007365f
C4096 vdd.n3104 gnd 0.007365f
C4097 vdd.n3105 gnd 0.007365f
C4098 vdd.n3106 gnd 0.007365f
C4099 vdd.n3107 gnd 0.007365f
C4100 vdd.n3108 gnd 0.007365f
C4101 vdd.n3109 gnd 0.007365f
C4102 vdd.n3111 gnd 0.007365f
C4103 vdd.n3112 gnd 0.007365f
C4104 vdd.n3113 gnd 0.007365f
C4105 vdd.n3114 gnd 0.007365f
C4106 vdd.n3115 gnd 0.007365f
C4107 vdd.n3116 gnd 0.007365f
C4108 vdd.n3118 gnd 0.007365f
C4109 vdd.n3119 gnd 0.007365f
C4110 vdd.n3120 gnd 0.007365f
C4111 vdd.n3122 gnd 0.007365f
C4112 vdd.n3123 gnd 0.007365f
C4113 vdd.n3124 gnd 0.007365f
C4114 vdd.n3125 gnd 0.007365f
C4115 vdd.n3126 gnd 0.007365f
C4116 vdd.n3127 gnd 0.007365f
C4117 vdd.n3129 gnd 0.007365f
C4118 vdd.n3130 gnd 0.007365f
C4119 vdd.n3131 gnd 0.007365f
C4120 vdd.n3132 gnd 0.007365f
C4121 vdd.n3133 gnd 0.007365f
C4122 vdd.n3134 gnd 0.007365f
C4123 vdd.n3136 gnd 0.007365f
C4124 vdd.n3137 gnd 0.007365f
C4125 vdd.n3138 gnd 0.007365f
C4126 vdd.n3139 gnd 0.007365f
C4127 vdd.n3140 gnd 0.007365f
C4128 vdd.n3141 gnd 0.007365f
C4129 vdd.n3143 gnd 0.007365f
C4130 vdd.n3144 gnd 0.007365f
C4131 vdd.n3146 gnd 0.007365f
C4132 vdd.n3147 gnd 0.007365f
C4133 vdd.n3148 gnd 0.017226f
C4134 vdd.n3149 gnd 0.016133f
C4135 vdd.n3150 gnd 0.016133f
C4136 vdd.n3151 gnd 1.06259f
C4137 vdd.n3152 gnd 0.016133f
C4138 vdd.n3153 gnd 0.017226f
C4139 vdd.n3154 gnd 0.016311f
C4140 vdd.n3155 gnd 0.007365f
C4141 vdd.n3156 gnd 0.005686f
C4142 vdd.n3157 gnd 0.007365f
C4143 vdd.n3159 gnd 0.007365f
C4144 vdd.n3160 gnd 0.007365f
C4145 vdd.n3161 gnd 0.007365f
C4146 vdd.n3162 gnd 0.007365f
C4147 vdd.n3163 gnd 0.007365f
C4148 vdd.n3164 gnd 0.007365f
C4149 vdd.n3166 gnd 0.007365f
C4150 vdd.n3167 gnd 0.007365f
C4151 vdd.n3168 gnd 0.007365f
C4152 vdd.n3169 gnd 0.007365f
C4153 vdd.n3170 gnd 0.007365f
C4154 vdd.n3171 gnd 0.007365f
C4155 vdd.n3173 gnd 0.007365f
C4156 vdd.n3174 gnd 0.007365f
C4157 vdd.n3175 gnd 0.007365f
C4158 vdd.n3176 gnd 0.007365f
C4159 vdd.n3177 gnd 0.007365f
C4160 vdd.n3178 gnd 0.007365f
C4161 vdd.n3180 gnd 0.007365f
C4162 vdd.n3181 gnd 0.007365f
C4163 vdd.n3183 gnd 0.007365f
C4164 vdd.n3184 gnd 0.025294f
C4165 vdd.n3185 gnd 0.823313f
C4166 vdd.n3187 gnd 0.004577f
C4167 vdd.n3188 gnd 0.008718f
C4168 vdd.n3189 gnd 0.010831f
C4169 vdd.n3190 gnd 0.010831f
C4170 vdd.n3191 gnd 0.008718f
C4171 vdd.n3192 gnd 0.008718f
C4172 vdd.n3193 gnd 0.010831f
C4173 vdd.n3194 gnd 0.010831f
C4174 vdd.n3195 gnd 0.008718f
C4175 vdd.n3196 gnd 0.008718f
C4176 vdd.n3197 gnd 0.010831f
C4177 vdd.n3198 gnd 0.010831f
C4178 vdd.n3199 gnd 0.008718f
C4179 vdd.n3200 gnd 0.008718f
C4180 vdd.n3201 gnd 0.010831f
C4181 vdd.n3202 gnd 0.010831f
C4182 vdd.n3203 gnd 0.008718f
C4183 vdd.n3204 gnd 0.008718f
C4184 vdd.n3205 gnd 0.010831f
C4185 vdd.n3206 gnd 0.010831f
C4186 vdd.n3207 gnd 0.008718f
C4187 vdd.n3208 gnd 0.008718f
C4188 vdd.n3209 gnd 0.010831f
C4189 vdd.n3210 gnd 0.010831f
C4190 vdd.n3211 gnd 0.008718f
C4191 vdd.n3212 gnd 0.008718f
C4192 vdd.n3213 gnd 0.010831f
C4193 vdd.n3214 gnd 0.010831f
C4194 vdd.n3215 gnd 0.008718f
C4195 vdd.n3216 gnd 0.008718f
C4196 vdd.n3217 gnd 0.010831f
C4197 vdd.n3218 gnd 0.010831f
C4198 vdd.n3219 gnd 0.008718f
C4199 vdd.n3220 gnd 0.008718f
C4200 vdd.n3221 gnd 0.010831f
C4201 vdd.n3222 gnd 0.010831f
C4202 vdd.n3223 gnd 0.008718f
C4203 vdd.n3224 gnd 0.010831f
C4204 vdd.n3225 gnd 0.010831f
C4205 vdd.n3226 gnd 0.008718f
C4206 vdd.n3227 gnd 0.010831f
C4207 vdd.n3228 gnd 0.010831f
C4208 vdd.n3229 gnd 0.010831f
C4209 vdd.n3230 gnd 0.017784f
C4210 vdd.n3231 gnd 0.010831f
C4211 vdd.n3232 gnd 0.010831f
C4212 vdd.n3233 gnd 0.005928f
C4213 vdd.n3234 gnd 0.008718f
C4214 vdd.n3235 gnd 0.010831f
C4215 vdd.n3236 gnd 0.010831f
C4216 vdd.n3237 gnd 0.008718f
C4217 vdd.n3238 gnd 0.008718f
C4218 vdd.n3239 gnd 0.010831f
C4219 vdd.n3240 gnd 0.010831f
C4220 vdd.n3241 gnd 0.008718f
C4221 vdd.n3242 gnd 0.008718f
C4222 vdd.n3243 gnd 0.010831f
C4223 vdd.n3244 gnd 0.010831f
C4224 vdd.n3245 gnd 0.008718f
C4225 vdd.n3246 gnd 0.008718f
C4226 vdd.n3247 gnd 0.010831f
C4227 vdd.n3248 gnd 0.010831f
C4228 vdd.n3249 gnd 0.008718f
C4229 vdd.n3250 gnd 0.008718f
C4230 vdd.n3251 gnd 0.010831f
C4231 vdd.n3252 gnd 0.010831f
C4232 vdd.n3253 gnd 0.008718f
C4233 vdd.n3254 gnd 0.008718f
C4234 vdd.n3255 gnd 0.010831f
C4235 vdd.n3256 gnd 0.010831f
C4236 vdd.n3257 gnd 0.008718f
C4237 vdd.n3258 gnd 0.008718f
C4238 vdd.n3259 gnd 0.010831f
C4239 vdd.n3260 gnd 0.010831f
C4240 vdd.n3261 gnd 0.008718f
C4241 vdd.n3262 gnd 0.008718f
C4242 vdd.n3263 gnd 0.010831f
C4243 vdd.n3264 gnd 0.010831f
C4244 vdd.n3265 gnd 0.008718f
C4245 vdd.n3266 gnd 0.008718f
C4246 vdd.n3267 gnd 0.010831f
C4247 vdd.n3268 gnd 0.010831f
C4248 vdd.n3269 gnd 0.008718f
C4249 vdd.n3270 gnd 0.010831f
C4250 vdd.n3271 gnd 0.010831f
C4251 vdd.n3272 gnd 0.008718f
C4252 vdd.n3273 gnd 0.010831f
C4253 vdd.n3274 gnd 0.010831f
C4254 vdd.n3275 gnd 0.010831f
C4255 vdd.t57 gnd 0.133248f
C4256 vdd.t58 gnd 0.142406f
C4257 vdd.t56 gnd 0.17402f
C4258 vdd.n3276 gnd 0.223069f
C4259 vdd.n3277 gnd 0.187419f
C4260 vdd.n3278 gnd 0.017784f
C4261 vdd.n3279 gnd 0.010831f
C4262 vdd.n3280 gnd 0.010831f
C4263 vdd.n3281 gnd 0.007279f
C4264 vdd.n3282 gnd 0.008718f
C4265 vdd.n3283 gnd 0.010831f
C4266 vdd.n3284 gnd 0.010831f
C4267 vdd.n3285 gnd 0.008718f
C4268 vdd.n3286 gnd 0.008718f
C4269 vdd.n3287 gnd 0.010831f
C4270 vdd.n3288 gnd 0.010831f
C4271 vdd.n3289 gnd 0.008718f
C4272 vdd.n3290 gnd 0.008718f
C4273 vdd.n3291 gnd 0.010831f
C4274 vdd.n3292 gnd 0.010831f
C4275 vdd.n3293 gnd 0.008718f
C4276 vdd.n3294 gnd 0.008718f
C4277 vdd.n3295 gnd 0.010831f
C4278 vdd.n3296 gnd 0.010831f
C4279 vdd.n3297 gnd 0.008718f
C4280 vdd.n3298 gnd 0.008718f
C4281 vdd.n3299 gnd 0.010831f
C4282 vdd.n3300 gnd 0.010831f
C4283 vdd.n3301 gnd 0.008718f
C4284 vdd.n3302 gnd 0.008718f
C4285 vdd.n3303 gnd 0.010831f
C4286 vdd.n3304 gnd 0.010831f
C4287 vdd.n3305 gnd 0.008718f
C4288 vdd.n3306 gnd 0.008718f
C4289 vdd.n3308 gnd 0.823313f
C4290 vdd.n3310 gnd 0.008718f
C4291 vdd.n3311 gnd 0.008718f
C4292 vdd.n3312 gnd 0.007236f
C4293 vdd.n3313 gnd 0.026762f
C4294 vdd.n3315 gnd 9.84001f
C4295 vdd.n3316 gnd 0.026762f
C4296 vdd.n3317 gnd 0.004141f
C4297 vdd.n3318 gnd 0.026762f
C4298 vdd.n3319 gnd 0.026201f
C4299 vdd.n3320 gnd 0.010831f
C4300 vdd.n3321 gnd 0.008718f
C4301 vdd.n3322 gnd 0.010831f
C4302 vdd.n3323 gnd 0.669652f
C4303 vdd.n3324 gnd 0.010831f
C4304 vdd.n3325 gnd 0.008718f
C4305 vdd.n3326 gnd 0.010831f
C4306 vdd.n3327 gnd 0.010831f
C4307 vdd.n3328 gnd 0.010831f
C4308 vdd.n3329 gnd 0.008718f
C4309 vdd.n3330 gnd 0.010831f
C4310 vdd.n3331 gnd 1.10686f
C4311 vdd.n3332 gnd 0.010831f
C4312 vdd.n3333 gnd 0.008718f
C4313 vdd.n3334 gnd 0.010831f
C4314 vdd.n3335 gnd 0.010831f
C4315 vdd.n3336 gnd 0.010831f
C4316 vdd.n3337 gnd 0.008718f
C4317 vdd.n3338 gnd 0.010831f
C4318 vdd.n3339 gnd 0.713927f
C4319 vdd.n3340 gnd 0.758201f
C4320 vdd.n3341 gnd 0.010831f
C4321 vdd.n3342 gnd 0.008718f
C4322 vdd.n3343 gnd 0.010831f
C4323 vdd.n3344 gnd 0.010831f
C4324 vdd.n3345 gnd 0.010831f
C4325 vdd.n3346 gnd 0.008718f
C4326 vdd.n3347 gnd 0.010831f
C4327 vdd.n3348 gnd 0.918696f
C4328 vdd.n3349 gnd 0.010831f
C4329 vdd.n3350 gnd 0.008718f
C4330 vdd.n3351 gnd 0.010831f
C4331 vdd.n3352 gnd 0.010831f
C4332 vdd.n3353 gnd 0.010831f
C4333 vdd.n3354 gnd 0.008718f
C4334 vdd.n3355 gnd 0.010831f
C4335 vdd.t202 gnd 0.553432f
C4336 vdd.n3356 gnd 0.891025f
C4337 vdd.n3357 gnd 0.010831f
C4338 vdd.n3358 gnd 0.008718f
C4339 vdd.n3359 gnd 0.010831f
C4340 vdd.n3360 gnd 0.010831f
C4341 vdd.n3361 gnd 0.010831f
C4342 vdd.n3362 gnd 0.008718f
C4343 vdd.n3363 gnd 0.010831f
C4344 vdd.n3364 gnd 0.702858f
C4345 vdd.n3365 gnd 0.010831f
C4346 vdd.n3366 gnd 0.008718f
C4347 vdd.n3367 gnd 0.010831f
C4348 vdd.n3368 gnd 0.010831f
C4349 vdd.n3369 gnd 0.010831f
C4350 vdd.n3370 gnd 0.008718f
C4351 vdd.n3371 gnd 0.010831f
C4352 vdd.n3372 gnd 0.879956f
C4353 vdd.n3373 gnd 0.592172f
C4354 vdd.n3374 gnd 0.010831f
C4355 vdd.n3375 gnd 0.008718f
C4356 vdd.n3376 gnd 0.010831f
C4357 vdd.n3377 gnd 0.010831f
C4358 vdd.n3378 gnd 0.010831f
C4359 vdd.n3379 gnd 0.008718f
C4360 vdd.n3380 gnd 0.010831f
C4361 vdd.n3381 gnd 0.780339f
C4362 vdd.n3382 gnd 0.010831f
C4363 vdd.n3383 gnd 0.008718f
C4364 vdd.n3384 gnd 0.010831f
C4365 vdd.n3385 gnd 0.010831f
C4366 vdd.n3386 gnd 0.010831f
C4367 vdd.n3387 gnd 0.010831f
C4368 vdd.n3388 gnd 0.010831f
C4369 vdd.n3389 gnd 0.008718f
C4370 vdd.n3390 gnd 0.008718f
C4371 vdd.n3391 gnd 0.010831f
C4372 vdd.t231 gnd 0.553432f
C4373 vdd.n3392 gnd 0.918696f
C4374 vdd.n3393 gnd 0.010831f
C4375 vdd.n3394 gnd 0.008718f
C4376 vdd.n3395 gnd 0.010831f
C4377 vdd.n3396 gnd 0.010831f
C4378 vdd.n3397 gnd 0.010831f
C4379 vdd.n3398 gnd 0.008718f
C4380 vdd.n3399 gnd 0.010831f
C4381 vdd.n3400 gnd 0.868888f
C4382 vdd.n3401 gnd 0.010831f
C4383 vdd.n3402 gnd 0.010831f
C4384 vdd.n3403 gnd 0.008718f
C4385 vdd.n3404 gnd 0.008718f
C4386 vdd.n3405 gnd 0.010831f
C4387 vdd.n3406 gnd 0.010831f
C4388 vdd.n3407 gnd 0.010831f
C4389 vdd.n3408 gnd 0.008718f
C4390 vdd.n3409 gnd 0.010831f
C4391 vdd.n3410 gnd 0.008718f
C4392 vdd.n3411 gnd 0.008718f
C4393 vdd.n3412 gnd 0.010831f
C4394 vdd.n3413 gnd 0.010831f
C4395 vdd.n3414 gnd 0.010831f
C4396 vdd.n3415 gnd 0.008718f
C4397 vdd.n3416 gnd 0.010831f
C4398 vdd.n3417 gnd 0.008718f
C4399 vdd.n3418 gnd 0.008718f
C4400 vdd.n3419 gnd 0.010831f
C4401 vdd.n3420 gnd 0.010831f
C4402 vdd.n3421 gnd 0.010831f
C4403 vdd.n3422 gnd 0.008718f
C4404 vdd.n3423 gnd 0.918696f
C4405 vdd.n3424 gnd 0.010831f
C4406 vdd.n3425 gnd 0.008718f
C4407 vdd.n3426 gnd 0.008718f
C4408 vdd.n3427 gnd 0.010831f
C4409 vdd.n3428 gnd 0.010831f
C4410 vdd.n3429 gnd 0.010831f
C4411 vdd.n3430 gnd 0.008718f
C4412 vdd.n3431 gnd 0.010831f
C4413 vdd.n3432 gnd 0.008718f
C4414 vdd.n3433 gnd 0.008718f
C4415 vdd.n3434 gnd 0.010831f
C4416 vdd.n3435 gnd 0.010831f
C4417 vdd.n3436 gnd 0.010831f
C4418 vdd.n3437 gnd 0.008718f
C4419 vdd.n3438 gnd 0.010831f
C4420 vdd.n3439 gnd 0.008718f
C4421 vdd.n3440 gnd 0.007236f
C4422 vdd.n3441 gnd 0.026201f
C4423 vdd.n3442 gnd 0.026762f
C4424 vdd.n3443 gnd 0.004141f
C4425 vdd.n3444 gnd 0.026762f
C4426 vdd.n3446 gnd 2.62327f
C4427 vdd.n3447 gnd 1.63262f
C4428 vdd.n3448 gnd 0.026201f
C4429 vdd.n3449 gnd 0.007236f
C4430 vdd.n3450 gnd 0.008718f
C4431 vdd.n3451 gnd 0.008718f
C4432 vdd.n3452 gnd 0.010831f
C4433 vdd.n3453 gnd 1.10686f
C4434 vdd.n3454 gnd 1.10686f
C4435 vdd.n3455 gnd 1.01278f
C4436 vdd.n3456 gnd 0.010831f
C4437 vdd.n3457 gnd 0.008718f
C4438 vdd.n3458 gnd 0.008718f
C4439 vdd.n3459 gnd 0.008718f
C4440 vdd.n3460 gnd 0.010831f
C4441 vdd.n3461 gnd 0.824613f
C4442 vdd.t259 gnd 0.553432f
C4443 vdd.n3462 gnd 0.835682f
C4444 vdd.n3463 gnd 0.636446f
C4445 vdd.n3464 gnd 0.010831f
C4446 vdd.n3465 gnd 0.008718f
C4447 vdd.n3466 gnd 0.008718f
C4448 vdd.n3467 gnd 0.008718f
C4449 vdd.n3468 gnd 0.010831f
C4450 vdd.n3469 gnd 0.658584f
C4451 vdd.n3470 gnd 0.813544f
C4452 vdd.t213 gnd 0.553432f
C4453 vdd.n3471 gnd 0.84675f
C4454 vdd.n3472 gnd 0.010831f
C4455 vdd.n3473 gnd 0.008718f
C4456 vdd.n3474 gnd 0.008718f
C4457 vdd.n3475 gnd 0.008718f
C4458 vdd.n3476 gnd 0.010831f
C4459 vdd.n3477 gnd 0.918696f
C4460 vdd.t158 gnd 0.553432f
C4461 vdd.n3478 gnd 0.669652f
C4462 vdd.n3479 gnd 0.802476f
C4463 vdd.n3480 gnd 0.010831f
C4464 vdd.n3481 gnd 0.008718f
C4465 vdd.n3482 gnd 0.008718f
C4466 vdd.n3483 gnd 0.008718f
C4467 vdd.n3484 gnd 0.010831f
C4468 vdd.n3485 gnd 0.614309f
C4469 vdd.t170 gnd 0.553432f
C4470 vdd.n3486 gnd 0.918696f
C4471 vdd.t162 gnd 0.553432f
C4472 vdd.n3487 gnd 0.680721f
C4473 vdd.n3488 gnd 0.010831f
C4474 vdd.n3489 gnd 0.008718f
C4475 vdd.n3490 gnd 0.008324f
C4476 vdd.n3491 gnd 0.638845f
C4477 vdd.n3492 gnd 2.90073f
C4478 a_n8300_8799.n0 gnd 0.209735f
C4479 a_n8300_8799.n1 gnd 0.287993f
C4480 a_n8300_8799.n2 gnd 0.209735f
C4481 a_n8300_8799.n3 gnd 0.209735f
C4482 a_n8300_8799.n4 gnd 0.209735f
C4483 a_n8300_8799.n5 gnd 0.209735f
C4484 a_n8300_8799.n6 gnd 0.209735f
C4485 a_n8300_8799.n7 gnd 0.218086f
C4486 a_n8300_8799.n8 gnd 0.209735f
C4487 a_n8300_8799.n9 gnd 0.287993f
C4488 a_n8300_8799.n10 gnd 0.209735f
C4489 a_n8300_8799.n11 gnd 0.209735f
C4490 a_n8300_8799.n12 gnd 0.209735f
C4491 a_n8300_8799.n13 gnd 0.209735f
C4492 a_n8300_8799.n14 gnd 0.209735f
C4493 a_n8300_8799.n15 gnd 0.218086f
C4494 a_n8300_8799.n16 gnd 0.209735f
C4495 a_n8300_8799.n17 gnd 0.454587f
C4496 a_n8300_8799.n18 gnd 0.209735f
C4497 a_n8300_8799.n19 gnd 0.209735f
C4498 a_n8300_8799.n20 gnd 0.209735f
C4499 a_n8300_8799.n21 gnd 0.209735f
C4500 a_n8300_8799.n22 gnd 0.209735f
C4501 a_n8300_8799.n23 gnd 0.218086f
C4502 a_n8300_8799.n24 gnd 0.209735f
C4503 a_n8300_8799.n25 gnd 0.322954f
C4504 a_n8300_8799.n26 gnd 0.209735f
C4505 a_n8300_8799.n27 gnd 0.209735f
C4506 a_n8300_8799.n28 gnd 0.209735f
C4507 a_n8300_8799.n29 gnd 0.209735f
C4508 a_n8300_8799.n30 gnd 0.209735f
C4509 a_n8300_8799.n31 gnd 0.183126f
C4510 a_n8300_8799.n32 gnd 0.209735f
C4511 a_n8300_8799.n33 gnd 0.322954f
C4512 a_n8300_8799.n34 gnd 0.209735f
C4513 a_n8300_8799.n35 gnd 0.209735f
C4514 a_n8300_8799.n36 gnd 0.209735f
C4515 a_n8300_8799.n37 gnd 0.209735f
C4516 a_n8300_8799.n38 gnd 0.209735f
C4517 a_n8300_8799.n39 gnd 0.183126f
C4518 a_n8300_8799.n40 gnd 0.209735f
C4519 a_n8300_8799.n41 gnd 0.322954f
C4520 a_n8300_8799.n42 gnd 0.209735f
C4521 a_n8300_8799.n43 gnd 0.209735f
C4522 a_n8300_8799.n44 gnd 0.209735f
C4523 a_n8300_8799.n45 gnd 0.209735f
C4524 a_n8300_8799.n46 gnd 0.209735f
C4525 a_n8300_8799.n47 gnd 0.349719f
C4526 a_n8300_8799.n48 gnd 0.706113f
C4527 a_n8300_8799.n49 gnd 2.92842f
C4528 a_n8300_8799.n50 gnd 2.87118f
C4529 a_n8300_8799.n51 gnd 1.40945f
C4530 a_n8300_8799.n52 gnd 1.02965f
C4531 a_n8300_8799.n53 gnd 2.58843f
C4532 a_n8300_8799.n54 gnd 3.19734f
C4533 a_n8300_8799.n55 gnd 1.53719f
C4534 a_n8300_8799.n56 gnd 0.252501f
C4535 a_n8300_8799.n57 gnd 0.003691f
C4536 a_n8300_8799.n58 gnd 0.009731f
C4537 a_n8300_8799.n59 gnd 0.010632f
C4538 a_n8300_8799.n60 gnd 0.005618f
C4539 a_n8300_8799.n62 gnd 0.004714f
C4540 a_n8300_8799.n63 gnd 0.010195f
C4541 a_n8300_8799.n64 gnd 0.010195f
C4542 a_n8300_8799.n65 gnd 0.004714f
C4543 a_n8300_8799.n67 gnd 0.005618f
C4544 a_n8300_8799.n68 gnd 0.010632f
C4545 a_n8300_8799.n69 gnd 0.009731f
C4546 a_n8300_8799.n70 gnd 0.003691f
C4547 a_n8300_8799.n71 gnd 0.252501f
C4548 a_n8300_8799.n72 gnd 0.003691f
C4549 a_n8300_8799.n73 gnd 0.009731f
C4550 a_n8300_8799.n74 gnd 0.010632f
C4551 a_n8300_8799.n75 gnd 0.005618f
C4552 a_n8300_8799.n77 gnd 0.004714f
C4553 a_n8300_8799.n78 gnd 0.010195f
C4554 a_n8300_8799.n79 gnd 0.010195f
C4555 a_n8300_8799.n80 gnd 0.004714f
C4556 a_n8300_8799.n82 gnd 0.005618f
C4557 a_n8300_8799.n83 gnd 0.010632f
C4558 a_n8300_8799.n84 gnd 0.009731f
C4559 a_n8300_8799.n85 gnd 0.003691f
C4560 a_n8300_8799.n86 gnd 0.252501f
C4561 a_n8300_8799.n87 gnd 0.003691f
C4562 a_n8300_8799.n88 gnd 0.009731f
C4563 a_n8300_8799.n89 gnd 0.010632f
C4564 a_n8300_8799.n90 gnd 0.005618f
C4565 a_n8300_8799.n92 gnd 0.004714f
C4566 a_n8300_8799.n93 gnd 0.010195f
C4567 a_n8300_8799.n94 gnd 0.010195f
C4568 a_n8300_8799.n95 gnd 0.004714f
C4569 a_n8300_8799.n97 gnd 0.005618f
C4570 a_n8300_8799.n98 gnd 0.010632f
C4571 a_n8300_8799.n99 gnd 0.009731f
C4572 a_n8300_8799.n100 gnd 0.003691f
C4573 a_n8300_8799.n101 gnd 0.003691f
C4574 a_n8300_8799.n102 gnd 0.009731f
C4575 a_n8300_8799.n103 gnd 0.010632f
C4576 a_n8300_8799.n104 gnd 0.005618f
C4577 a_n8300_8799.n106 gnd 0.004714f
C4578 a_n8300_8799.n107 gnd 0.010195f
C4579 a_n8300_8799.n108 gnd 0.010195f
C4580 a_n8300_8799.n109 gnd 0.004714f
C4581 a_n8300_8799.n111 gnd 0.005618f
C4582 a_n8300_8799.n112 gnd 0.010632f
C4583 a_n8300_8799.n113 gnd 0.009731f
C4584 a_n8300_8799.n114 gnd 0.003691f
C4585 a_n8300_8799.n115 gnd 0.252501f
C4586 a_n8300_8799.n116 gnd 0.003691f
C4587 a_n8300_8799.n117 gnd 0.009731f
C4588 a_n8300_8799.n118 gnd 0.010632f
C4589 a_n8300_8799.n119 gnd 0.005618f
C4590 a_n8300_8799.n121 gnd 0.004714f
C4591 a_n8300_8799.n122 gnd 0.010195f
C4592 a_n8300_8799.n123 gnd 0.010195f
C4593 a_n8300_8799.n124 gnd 0.004714f
C4594 a_n8300_8799.n126 gnd 0.005618f
C4595 a_n8300_8799.n127 gnd 0.010632f
C4596 a_n8300_8799.n128 gnd 0.009731f
C4597 a_n8300_8799.n129 gnd 0.003691f
C4598 a_n8300_8799.n130 gnd 0.252501f
C4599 a_n8300_8799.n131 gnd 0.003691f
C4600 a_n8300_8799.n132 gnd 0.009731f
C4601 a_n8300_8799.n133 gnd 0.010632f
C4602 a_n8300_8799.n134 gnd 0.005618f
C4603 a_n8300_8799.n136 gnd 0.004714f
C4604 a_n8300_8799.n137 gnd 0.010195f
C4605 a_n8300_8799.n138 gnd 0.010195f
C4606 a_n8300_8799.n139 gnd 0.004714f
C4607 a_n8300_8799.n141 gnd 0.005618f
C4608 a_n8300_8799.n142 gnd 0.010632f
C4609 a_n8300_8799.n143 gnd 0.009731f
C4610 a_n8300_8799.n144 gnd 0.003691f
C4611 a_n8300_8799.n145 gnd 0.252501f
C4612 a_n8300_8799.t12 gnd 0.145474f
C4613 a_n8300_8799.t23 gnd 0.145474f
C4614 a_n8300_8799.t13 gnd 0.145474f
C4615 a_n8300_8799.n146 gnd 1.14738f
C4616 a_n8300_8799.t11 gnd 0.145474f
C4617 a_n8300_8799.t21 gnd 0.145474f
C4618 a_n8300_8799.n147 gnd 1.14549f
C4619 a_n8300_8799.t27 gnd 0.145474f
C4620 a_n8300_8799.t25 gnd 0.145474f
C4621 a_n8300_8799.n148 gnd 1.14549f
C4622 a_n8300_8799.t19 gnd 0.145474f
C4623 a_n8300_8799.t14 gnd 0.145474f
C4624 a_n8300_8799.n149 gnd 1.14549f
C4625 a_n8300_8799.t18 gnd 0.113147f
C4626 a_n8300_8799.t31 gnd 0.113147f
C4627 a_n8300_8799.n150 gnd 1.0014f
C4628 a_n8300_8799.t35 gnd 0.113147f
C4629 a_n8300_8799.t33 gnd 0.113147f
C4630 a_n8300_8799.n151 gnd 0.999805f
C4631 a_n8300_8799.t2 gnd 0.113147f
C4632 a_n8300_8799.t3 gnd 0.113147f
C4633 a_n8300_8799.n152 gnd 0.999805f
C4634 a_n8300_8799.t9 gnd 0.113147f
C4635 a_n8300_8799.t16 gnd 0.113147f
C4636 a_n8300_8799.n153 gnd 1.0014f
C4637 a_n8300_8799.t32 gnd 0.113147f
C4638 a_n8300_8799.t8 gnd 0.113147f
C4639 a_n8300_8799.n154 gnd 0.999804f
C4640 a_n8300_8799.t1 gnd 0.113147f
C4641 a_n8300_8799.t10 gnd 0.113147f
C4642 a_n8300_8799.n155 gnd 0.999804f
C4643 a_n8300_8799.t30 gnd 0.113147f
C4644 a_n8300_8799.t0 gnd 0.113147f
C4645 a_n8300_8799.n156 gnd 1.0014f
C4646 a_n8300_8799.t4 gnd 0.113147f
C4647 a_n8300_8799.t17 gnd 0.113147f
C4648 a_n8300_8799.n157 gnd 0.999804f
C4649 a_n8300_8799.t34 gnd 0.113147f
C4650 a_n8300_8799.t7 gnd 0.113147f
C4651 a_n8300_8799.n158 gnd 0.999805f
C4652 a_n8300_8799.t29 gnd 0.113147f
C4653 a_n8300_8799.t6 gnd 0.113147f
C4654 a_n8300_8799.n159 gnd 0.999805f
C4655 a_n8300_8799.t88 gnd 0.603205f
C4656 a_n8300_8799.n160 gnd 0.27157f
C4657 a_n8300_8799.t36 gnd 0.603205f
C4658 a_n8300_8799.t67 gnd 0.603205f
C4659 a_n8300_8799.n161 gnd 0.273516f
C4660 a_n8300_8799.t68 gnd 0.603205f
C4661 a_n8300_8799.t82 gnd 0.603205f
C4662 a_n8300_8799.n162 gnd 0.266655f
C4663 a_n8300_8799.t134 gnd 0.603205f
C4664 a_n8300_8799.t137 gnd 0.603205f
C4665 a_n8300_8799.n163 gnd 0.270669f
C4666 a_n8300_8799.t98 gnd 0.603205f
C4667 a_n8300_8799.t142 gnd 0.603205f
C4668 a_n8300_8799.t103 gnd 0.614621f
C4669 a_n8300_8799.n164 gnd 0.252868f
C4670 a_n8300_8799.n165 gnd 0.273892f
C4671 a_n8300_8799.t65 gnd 0.603205f
C4672 a_n8300_8799.n166 gnd 0.27157f
C4673 a_n8300_8799.n167 gnd 0.267301f
C4674 a_n8300_8799.t135 gnd 0.603205f
C4675 a_n8300_8799.n168 gnd 0.266008f
C4676 a_n8300_8799.t83 gnd 0.603205f
C4677 a_n8300_8799.n169 gnd 0.273259f
C4678 a_n8300_8799.t114 gnd 0.603205f
C4679 a_n8300_8799.n170 gnd 0.273516f
C4680 a_n8300_8799.n171 gnd 0.271106f
C4681 a_n8300_8799.t81 gnd 0.603205f
C4682 a_n8300_8799.n172 gnd 0.266655f
C4683 a_n8300_8799.t111 gnd 0.603205f
C4684 a_n8300_8799.n173 gnd 0.271106f
C4685 a_n8300_8799.n174 gnd 0.273259f
C4686 a_n8300_8799.t108 gnd 0.603205f
C4687 a_n8300_8799.n175 gnd 0.270669f
C4688 a_n8300_8799.n176 gnd 0.266008f
C4689 a_n8300_8799.t66 gnd 0.603205f
C4690 a_n8300_8799.n177 gnd 0.267301f
C4691 a_n8300_8799.t136 gnd 0.603205f
C4692 a_n8300_8799.n178 gnd 0.273892f
C4693 a_n8300_8799.t47 gnd 0.614611f
C4694 a_n8300_8799.t100 gnd 0.603205f
C4695 a_n8300_8799.n179 gnd 0.27157f
C4696 a_n8300_8799.t46 gnd 0.603205f
C4697 a_n8300_8799.t79 gnd 0.603205f
C4698 a_n8300_8799.n180 gnd 0.273516f
C4699 a_n8300_8799.t80 gnd 0.603205f
C4700 a_n8300_8799.t90 gnd 0.603205f
C4701 a_n8300_8799.n181 gnd 0.266655f
C4702 a_n8300_8799.t148 gnd 0.603205f
C4703 a_n8300_8799.t153 gnd 0.603205f
C4704 a_n8300_8799.n182 gnd 0.270669f
C4705 a_n8300_8799.t112 gnd 0.603205f
C4706 a_n8300_8799.t155 gnd 0.603205f
C4707 a_n8300_8799.t119 gnd 0.614621f
C4708 a_n8300_8799.n183 gnd 0.252868f
C4709 a_n8300_8799.n184 gnd 0.273892f
C4710 a_n8300_8799.t75 gnd 0.603205f
C4711 a_n8300_8799.n185 gnd 0.27157f
C4712 a_n8300_8799.n186 gnd 0.267301f
C4713 a_n8300_8799.t150 gnd 0.603205f
C4714 a_n8300_8799.n187 gnd 0.266008f
C4715 a_n8300_8799.t93 gnd 0.603205f
C4716 a_n8300_8799.n188 gnd 0.273259f
C4717 a_n8300_8799.t131 gnd 0.603205f
C4718 a_n8300_8799.n189 gnd 0.273516f
C4719 a_n8300_8799.n190 gnd 0.271106f
C4720 a_n8300_8799.t89 gnd 0.603205f
C4721 a_n8300_8799.n191 gnd 0.266655f
C4722 a_n8300_8799.t129 gnd 0.603205f
C4723 a_n8300_8799.n192 gnd 0.271106f
C4724 a_n8300_8799.n193 gnd 0.273259f
C4725 a_n8300_8799.t125 gnd 0.603205f
C4726 a_n8300_8799.n194 gnd 0.270669f
C4727 a_n8300_8799.n195 gnd 0.266008f
C4728 a_n8300_8799.t76 gnd 0.603205f
C4729 a_n8300_8799.n196 gnd 0.267301f
C4730 a_n8300_8799.t151 gnd 0.603205f
C4731 a_n8300_8799.n197 gnd 0.273892f
C4732 a_n8300_8799.t59 gnd 0.614611f
C4733 a_n8300_8799.n198 gnd 0.906834f
C4734 a_n8300_8799.t104 gnd 0.603205f
C4735 a_n8300_8799.n199 gnd 0.27157f
C4736 a_n8300_8799.t87 gnd 0.603205f
C4737 a_n8300_8799.t141 gnd 0.603205f
C4738 a_n8300_8799.n200 gnd 0.273516f
C4739 a_n8300_8799.t113 gnd 0.603205f
C4740 a_n8300_8799.t37 gnd 0.603205f
C4741 a_n8300_8799.n201 gnd 0.266655f
C4742 a_n8300_8799.t138 gnd 0.603205f
C4743 a_n8300_8799.t86 gnd 0.603205f
C4744 a_n8300_8799.n202 gnd 0.270669f
C4745 a_n8300_8799.t48 gnd 0.603205f
C4746 a_n8300_8799.t70 gnd 0.603205f
C4747 a_n8300_8799.t121 gnd 0.614621f
C4748 a_n8300_8799.n203 gnd 0.252868f
C4749 a_n8300_8799.n204 gnd 0.273892f
C4750 a_n8300_8799.t91 gnd 0.603205f
C4751 a_n8300_8799.n205 gnd 0.27157f
C4752 a_n8300_8799.n206 gnd 0.267301f
C4753 a_n8300_8799.t109 gnd 0.603205f
C4754 a_n8300_8799.n207 gnd 0.266008f
C4755 a_n8300_8799.t130 gnd 0.603205f
C4756 a_n8300_8799.n208 gnd 0.273259f
C4757 a_n8300_8799.t77 gnd 0.603205f
C4758 a_n8300_8799.n209 gnd 0.273516f
C4759 a_n8300_8799.n210 gnd 0.271106f
C4760 a_n8300_8799.t53 gnd 0.603205f
C4761 a_n8300_8799.n211 gnd 0.266655f
C4762 a_n8300_8799.t94 gnd 0.603205f
C4763 a_n8300_8799.n212 gnd 0.271106f
C4764 a_n8300_8799.n213 gnd 0.273259f
C4765 a_n8300_8799.t147 gnd 0.603205f
C4766 a_n8300_8799.n214 gnd 0.270669f
C4767 a_n8300_8799.n215 gnd 0.266008f
C4768 a_n8300_8799.t42 gnd 0.603205f
C4769 a_n8300_8799.n216 gnd 0.267301f
C4770 a_n8300_8799.t57 gnd 0.603205f
C4771 a_n8300_8799.n217 gnd 0.273892f
C4772 a_n8300_8799.t126 gnd 0.614611f
C4773 a_n8300_8799.n218 gnd 1.55651f
C4774 a_n8300_8799.t85 gnd 0.614611f
C4775 a_n8300_8799.t61 gnd 0.603205f
C4776 a_n8300_8799.t140 gnd 0.603205f
C4777 a_n8300_8799.n219 gnd 0.27157f
C4778 a_n8300_8799.t102 gnd 0.603205f
C4779 a_n8300_8799.t99 gnd 0.603205f
C4780 a_n8300_8799.t39 gnd 0.603205f
C4781 a_n8300_8799.n220 gnd 0.270669f
C4782 a_n8300_8799.t107 gnd 0.603205f
C4783 a_n8300_8799.t106 gnd 0.603205f
C4784 a_n8300_8799.t41 gnd 0.603205f
C4785 a_n8300_8799.n221 gnd 0.271106f
C4786 a_n8300_8799.t40 gnd 0.603205f
C4787 a_n8300_8799.t128 gnd 0.603205f
C4788 a_n8300_8799.t56 gnd 0.603205f
C4789 a_n8300_8799.n222 gnd 0.271106f
C4790 a_n8300_8799.t45 gnd 0.603205f
C4791 a_n8300_8799.t132 gnd 0.603205f
C4792 a_n8300_8799.t84 gnd 0.603205f
C4793 a_n8300_8799.n223 gnd 0.270669f
C4794 a_n8300_8799.t60 gnd 0.603205f
C4795 a_n8300_8799.t152 gnd 0.603205f
C4796 a_n8300_8799.t101 gnd 0.603205f
C4797 a_n8300_8799.n224 gnd 0.27157f
C4798 a_n8300_8799.t145 gnd 0.614621f
C4799 a_n8300_8799.n225 gnd 0.252868f
C4800 a_n8300_8799.t63 gnd 0.603205f
C4801 a_n8300_8799.n226 gnd 0.273892f
C4802 a_n8300_8799.n227 gnd 0.267301f
C4803 a_n8300_8799.n228 gnd 0.266008f
C4804 a_n8300_8799.n229 gnd 0.273259f
C4805 a_n8300_8799.n230 gnd 0.273516f
C4806 a_n8300_8799.n231 gnd 0.266655f
C4807 a_n8300_8799.n232 gnd 0.266655f
C4808 a_n8300_8799.n233 gnd 0.273516f
C4809 a_n8300_8799.n234 gnd 0.273259f
C4810 a_n8300_8799.n235 gnd 0.266008f
C4811 a_n8300_8799.n236 gnd 0.267301f
C4812 a_n8300_8799.n237 gnd 0.273892f
C4813 a_n8300_8799.t96 gnd 0.614611f
C4814 a_n8300_8799.t72 gnd 0.603205f
C4815 a_n8300_8799.t154 gnd 0.603205f
C4816 a_n8300_8799.n238 gnd 0.27157f
C4817 a_n8300_8799.t117 gnd 0.603205f
C4818 a_n8300_8799.t116 gnd 0.603205f
C4819 a_n8300_8799.t50 gnd 0.603205f
C4820 a_n8300_8799.n239 gnd 0.270669f
C4821 a_n8300_8799.t124 gnd 0.603205f
C4822 a_n8300_8799.t123 gnd 0.603205f
C4823 a_n8300_8799.t52 gnd 0.603205f
C4824 a_n8300_8799.n240 gnd 0.271106f
C4825 a_n8300_8799.t51 gnd 0.603205f
C4826 a_n8300_8799.t144 gnd 0.603205f
C4827 a_n8300_8799.t69 gnd 0.603205f
C4828 a_n8300_8799.n241 gnd 0.271106f
C4829 a_n8300_8799.t55 gnd 0.603205f
C4830 a_n8300_8799.t146 gnd 0.603205f
C4831 a_n8300_8799.t97 gnd 0.603205f
C4832 a_n8300_8799.n242 gnd 0.270669f
C4833 a_n8300_8799.t73 gnd 0.603205f
C4834 a_n8300_8799.t43 gnd 0.603205f
C4835 a_n8300_8799.t118 gnd 0.603205f
C4836 a_n8300_8799.n243 gnd 0.27157f
C4837 a_n8300_8799.t38 gnd 0.614621f
C4838 a_n8300_8799.n244 gnd 0.252868f
C4839 a_n8300_8799.t74 gnd 0.603205f
C4840 a_n8300_8799.n245 gnd 0.273892f
C4841 a_n8300_8799.n246 gnd 0.267301f
C4842 a_n8300_8799.n247 gnd 0.266008f
C4843 a_n8300_8799.n248 gnd 0.273259f
C4844 a_n8300_8799.n249 gnd 0.273516f
C4845 a_n8300_8799.n250 gnd 0.266655f
C4846 a_n8300_8799.n251 gnd 0.266655f
C4847 a_n8300_8799.n252 gnd 0.273516f
C4848 a_n8300_8799.n253 gnd 0.273259f
C4849 a_n8300_8799.n254 gnd 0.266008f
C4850 a_n8300_8799.n255 gnd 0.267301f
C4851 a_n8300_8799.n256 gnd 0.273892f
C4852 a_n8300_8799.n257 gnd 0.906834f
C4853 a_n8300_8799.t127 gnd 0.614611f
C4854 a_n8300_8799.t58 gnd 0.603205f
C4855 a_n8300_8799.t105 gnd 0.603205f
C4856 a_n8300_8799.n258 gnd 0.27157f
C4857 a_n8300_8799.t44 gnd 0.603205f
C4858 a_n8300_8799.t64 gnd 0.603205f
C4859 a_n8300_8799.t149 gnd 0.603205f
C4860 a_n8300_8799.n259 gnd 0.270669f
C4861 a_n8300_8799.t115 gnd 0.603205f
C4862 a_n8300_8799.t143 gnd 0.603205f
C4863 a_n8300_8799.t95 gnd 0.603205f
C4864 a_n8300_8799.n260 gnd 0.271106f
C4865 a_n8300_8799.t122 gnd 0.603205f
C4866 a_n8300_8799.t54 gnd 0.603205f
C4867 a_n8300_8799.t139 gnd 0.603205f
C4868 a_n8300_8799.n261 gnd 0.271106f
C4869 a_n8300_8799.t78 gnd 0.603205f
C4870 a_n8300_8799.t133 gnd 0.603205f
C4871 a_n8300_8799.t62 gnd 0.603205f
C4872 a_n8300_8799.n262 gnd 0.270669f
C4873 a_n8300_8799.t110 gnd 0.603205f
C4874 a_n8300_8799.t49 gnd 0.603205f
C4875 a_n8300_8799.t92 gnd 0.603205f
C4876 a_n8300_8799.n263 gnd 0.27157f
C4877 a_n8300_8799.t120 gnd 0.614621f
C4878 a_n8300_8799.n264 gnd 0.252868f
C4879 a_n8300_8799.t71 gnd 0.603205f
C4880 a_n8300_8799.n265 gnd 0.273892f
C4881 a_n8300_8799.n266 gnd 0.267301f
C4882 a_n8300_8799.n267 gnd 0.266008f
C4883 a_n8300_8799.n268 gnd 0.273259f
C4884 a_n8300_8799.n269 gnd 0.273516f
C4885 a_n8300_8799.n270 gnd 0.266655f
C4886 a_n8300_8799.n271 gnd 0.266655f
C4887 a_n8300_8799.n272 gnd 0.273516f
C4888 a_n8300_8799.n273 gnd 0.273259f
C4889 a_n8300_8799.n274 gnd 0.266008f
C4890 a_n8300_8799.n275 gnd 0.267301f
C4891 a_n8300_8799.n276 gnd 0.273892f
C4892 a_n8300_8799.n277 gnd 1.25096f
C4893 a_n8300_8799.n278 gnd 14.1132f
C4894 a_n8300_8799.n279 gnd 4.41458f
C4895 a_n8300_8799.n280 gnd 6.40591f
C4896 a_n8300_8799.t24 gnd 0.145474f
C4897 a_n8300_8799.t20 gnd 0.145474f
C4898 a_n8300_8799.n281 gnd 1.14549f
C4899 a_n8300_8799.t22 gnd 0.145474f
C4900 a_n8300_8799.t26 gnd 0.145474f
C4901 a_n8300_8799.n282 gnd 1.14549f
C4902 a_n8300_8799.t28 gnd 0.145474f
C4903 a_n8300_8799.t15 gnd 0.145474f
C4904 a_n8300_8799.n283 gnd 1.14738f
C4905 a_n8300_8799.n284 gnd 1.14549f
C4906 a_n8300_8799.t5 gnd 0.145474f
C4907 CSoutput.n0 gnd 0.048434f
C4908 CSoutput.t218 gnd 0.320378f
C4909 CSoutput.n1 gnd 0.144666f
C4910 CSoutput.n2 gnd 0.048434f
C4911 CSoutput.t216 gnd 0.320378f
C4912 CSoutput.n3 gnd 0.038387f
C4913 CSoutput.n4 gnd 0.048434f
C4914 CSoutput.t209 gnd 0.320378f
C4915 CSoutput.n5 gnd 0.033102f
C4916 CSoutput.n6 gnd 0.048434f
C4917 CSoutput.t213 gnd 0.320378f
C4918 CSoutput.t202 gnd 0.320378f
C4919 CSoutput.n7 gnd 0.14309f
C4920 CSoutput.n8 gnd 0.048434f
C4921 CSoutput.t201 gnd 0.320378f
C4922 CSoutput.n9 gnd 0.031561f
C4923 CSoutput.n10 gnd 0.048434f
C4924 CSoutput.t210 gnd 0.320378f
C4925 CSoutput.t215 gnd 0.320378f
C4926 CSoutput.n11 gnd 0.14309f
C4927 CSoutput.n12 gnd 0.048434f
C4928 CSoutput.t221 gnd 0.320378f
C4929 CSoutput.n13 gnd 0.033102f
C4930 CSoutput.n14 gnd 0.048434f
C4931 CSoutput.t203 gnd 0.320378f
C4932 CSoutput.t212 gnd 0.320378f
C4933 CSoutput.n15 gnd 0.14309f
C4934 CSoutput.n16 gnd 0.048434f
C4935 CSoutput.t219 gnd 0.320378f
C4936 CSoutput.n17 gnd 0.035354f
C4937 CSoutput.t206 gnd 0.38286f
C4938 CSoutput.t217 gnd 0.320378f
C4939 CSoutput.n18 gnd 0.18267f
C4940 CSoutput.n19 gnd 0.177253f
C4941 CSoutput.n20 gnd 0.205635f
C4942 CSoutput.n21 gnd 0.048434f
C4943 CSoutput.n22 gnd 0.040423f
C4944 CSoutput.n23 gnd 0.14309f
C4945 CSoutput.n24 gnd 0.038967f
C4946 CSoutput.n25 gnd 0.038387f
C4947 CSoutput.n26 gnd 0.048434f
C4948 CSoutput.n27 gnd 0.048434f
C4949 CSoutput.n28 gnd 0.040112f
C4950 CSoutput.n29 gnd 0.034056f
C4951 CSoutput.n30 gnd 0.146275f
C4952 CSoutput.n31 gnd 0.034525f
C4953 CSoutput.n32 gnd 0.048434f
C4954 CSoutput.n33 gnd 0.048434f
C4955 CSoutput.n34 gnd 0.048434f
C4956 CSoutput.n35 gnd 0.039685f
C4957 CSoutput.n36 gnd 0.14309f
C4958 CSoutput.n37 gnd 0.037953f
C4959 CSoutput.n38 gnd 0.039401f
C4960 CSoutput.n39 gnd 0.048434f
C4961 CSoutput.n40 gnd 0.048434f
C4962 CSoutput.n41 gnd 0.040415f
C4963 CSoutput.n42 gnd 0.036939f
C4964 CSoutput.n43 gnd 0.14309f
C4965 CSoutput.n44 gnd 0.037876f
C4966 CSoutput.n45 gnd 0.048434f
C4967 CSoutput.n46 gnd 0.048434f
C4968 CSoutput.n47 gnd 0.048434f
C4969 CSoutput.n48 gnd 0.037876f
C4970 CSoutput.n49 gnd 0.14309f
C4971 CSoutput.n50 gnd 0.036939f
C4972 CSoutput.n51 gnd 0.040415f
C4973 CSoutput.n52 gnd 0.048434f
C4974 CSoutput.n53 gnd 0.048434f
C4975 CSoutput.n54 gnd 0.039401f
C4976 CSoutput.n55 gnd 0.037953f
C4977 CSoutput.n56 gnd 0.14309f
C4978 CSoutput.n57 gnd 0.039685f
C4979 CSoutput.n58 gnd 0.048434f
C4980 CSoutput.n59 gnd 0.048434f
C4981 CSoutput.n60 gnd 0.048434f
C4982 CSoutput.n61 gnd 0.034525f
C4983 CSoutput.n62 gnd 0.146275f
C4984 CSoutput.n63 gnd 0.034056f
C4985 CSoutput.t205 gnd 0.320378f
C4986 CSoutput.n64 gnd 0.14309f
C4987 CSoutput.n65 gnd 0.040112f
C4988 CSoutput.n66 gnd 0.048434f
C4989 CSoutput.n67 gnd 0.048434f
C4990 CSoutput.n68 gnd 0.048434f
C4991 CSoutput.n69 gnd 0.038967f
C4992 CSoutput.n70 gnd 0.14309f
C4993 CSoutput.n71 gnd 0.040423f
C4994 CSoutput.n72 gnd 0.035354f
C4995 CSoutput.n73 gnd 0.048434f
C4996 CSoutput.n74 gnd 0.048434f
C4997 CSoutput.n75 gnd 0.036665f
C4998 CSoutput.n76 gnd 0.021775f
C4999 CSoutput.t208 gnd 0.359967f
C5000 CSoutput.n77 gnd 0.178817f
C5001 CSoutput.n78 gnd 0.765143f
C5002 CSoutput.t62 gnd 0.060414f
C5003 CSoutput.t9 gnd 0.060414f
C5004 CSoutput.n79 gnd 0.467746f
C5005 CSoutput.t194 gnd 0.060414f
C5006 CSoutput.t60 gnd 0.060414f
C5007 CSoutput.n80 gnd 0.466912f
C5008 CSoutput.n81 gnd 0.473915f
C5009 CSoutput.t196 gnd 0.060414f
C5010 CSoutput.t186 gnd 0.060414f
C5011 CSoutput.n82 gnd 0.466912f
C5012 CSoutput.n83 gnd 0.233525f
C5013 CSoutput.t56 gnd 0.060414f
C5014 CSoutput.t89 gnd 0.060414f
C5015 CSoutput.n84 gnd 0.466912f
C5016 CSoutput.n85 gnd 0.233525f
C5017 CSoutput.t0 gnd 0.060414f
C5018 CSoutput.t65 gnd 0.060414f
C5019 CSoutput.n86 gnd 0.466912f
C5020 CSoutput.n87 gnd 0.233525f
C5021 CSoutput.t68 gnd 0.060414f
C5022 CSoutput.t180 gnd 0.060414f
C5023 CSoutput.n88 gnd 0.466912f
C5024 CSoutput.n89 gnd 0.233525f
C5025 CSoutput.t50 gnd 0.060414f
C5026 CSoutput.t72 gnd 0.060414f
C5027 CSoutput.n90 gnd 0.466912f
C5028 CSoutput.n91 gnd 0.233525f
C5029 CSoutput.t73 gnd 0.060414f
C5030 CSoutput.t71 gnd 0.060414f
C5031 CSoutput.n92 gnd 0.466912f
C5032 CSoutput.n93 gnd 0.233525f
C5033 CSoutput.t99 gnd 0.060414f
C5034 CSoutput.t43 gnd 0.060414f
C5035 CSoutput.n94 gnd 0.466912f
C5036 CSoutput.n95 gnd 0.233525f
C5037 CSoutput.t187 gnd 0.060414f
C5038 CSoutput.t4 gnd 0.060414f
C5039 CSoutput.n96 gnd 0.466912f
C5040 CSoutput.n97 gnd 0.428232f
C5041 CSoutput.t190 gnd 0.060414f
C5042 CSoutput.t10 gnd 0.060414f
C5043 CSoutput.n98 gnd 0.467746f
C5044 CSoutput.t24 gnd 0.060414f
C5045 CSoutput.t18 gnd 0.060414f
C5046 CSoutput.n99 gnd 0.466912f
C5047 CSoutput.n100 gnd 0.473915f
C5048 CSoutput.t192 gnd 0.060414f
C5049 CSoutput.t61 gnd 0.060414f
C5050 CSoutput.n101 gnd 0.466912f
C5051 CSoutput.n102 gnd 0.233525f
C5052 CSoutput.t69 gnd 0.060414f
C5053 CSoutput.t91 gnd 0.060414f
C5054 CSoutput.n103 gnd 0.466912f
C5055 CSoutput.n104 gnd 0.233525f
C5056 CSoutput.t41 gnd 0.060414f
C5057 CSoutput.t83 gnd 0.060414f
C5058 CSoutput.n105 gnd 0.466912f
C5059 CSoutput.n106 gnd 0.233525f
C5060 CSoutput.t31 gnd 0.060414f
C5061 CSoutput.t193 gnd 0.060414f
C5062 CSoutput.n107 gnd 0.466912f
C5063 CSoutput.n108 gnd 0.233525f
C5064 CSoutput.t16 gnd 0.060414f
C5065 CSoutput.t64 gnd 0.060414f
C5066 CSoutput.n109 gnd 0.466912f
C5067 CSoutput.n110 gnd 0.233525f
C5068 CSoutput.t79 gnd 0.060414f
C5069 CSoutput.t199 gnd 0.060414f
C5070 CSoutput.n111 gnd 0.466912f
C5071 CSoutput.n112 gnd 0.233525f
C5072 CSoutput.t52 gnd 0.060414f
C5073 CSoutput.t21 gnd 0.060414f
C5074 CSoutput.n113 gnd 0.466912f
C5075 CSoutput.n114 gnd 0.233525f
C5076 CSoutput.t14 gnd 0.060414f
C5077 CSoutput.t49 gnd 0.060414f
C5078 CSoutput.n115 gnd 0.466912f
C5079 CSoutput.n116 gnd 0.348245f
C5080 CSoutput.n117 gnd 0.439135f
C5081 CSoutput.t3 gnd 0.060414f
C5082 CSoutput.t80 gnd 0.060414f
C5083 CSoutput.n118 gnd 0.467746f
C5084 CSoutput.t19 gnd 0.060414f
C5085 CSoutput.t37 gnd 0.060414f
C5086 CSoutput.n119 gnd 0.466912f
C5087 CSoutput.n120 gnd 0.473915f
C5088 CSoutput.t181 gnd 0.060414f
C5089 CSoutput.t48 gnd 0.060414f
C5090 CSoutput.n121 gnd 0.466912f
C5091 CSoutput.n122 gnd 0.233525f
C5092 CSoutput.t183 gnd 0.060414f
C5093 CSoutput.t184 gnd 0.060414f
C5094 CSoutput.n123 gnd 0.466912f
C5095 CSoutput.n124 gnd 0.233525f
C5096 CSoutput.t93 gnd 0.060414f
C5097 CSoutput.t182 gnd 0.060414f
C5098 CSoutput.n125 gnd 0.466912f
C5099 CSoutput.n126 gnd 0.233525f
C5100 CSoutput.t63 gnd 0.060414f
C5101 CSoutput.t92 gnd 0.060414f
C5102 CSoutput.n127 gnd 0.466912f
C5103 CSoutput.n128 gnd 0.233525f
C5104 CSoutput.t94 gnd 0.060414f
C5105 CSoutput.t32 gnd 0.060414f
C5106 CSoutput.n129 gnd 0.466912f
C5107 CSoutput.n130 gnd 0.233525f
C5108 CSoutput.t40 gnd 0.060414f
C5109 CSoutput.t45 gnd 0.060414f
C5110 CSoutput.n131 gnd 0.466912f
C5111 CSoutput.n132 gnd 0.233525f
C5112 CSoutput.t8 gnd 0.060414f
C5113 CSoutput.t5 gnd 0.060414f
C5114 CSoutput.n133 gnd 0.466912f
C5115 CSoutput.n134 gnd 0.233525f
C5116 CSoutput.t28 gnd 0.060414f
C5117 CSoutput.t78 gnd 0.060414f
C5118 CSoutput.n135 gnd 0.466912f
C5119 CSoutput.n136 gnd 0.348245f
C5120 CSoutput.n137 gnd 0.49084f
C5121 CSoutput.n138 gnd 9.77039f
C5122 CSoutput.n140 gnd 0.856782f
C5123 CSoutput.n141 gnd 0.642586f
C5124 CSoutput.n142 gnd 0.856782f
C5125 CSoutput.n143 gnd 0.856782f
C5126 CSoutput.n144 gnd 2.30672f
C5127 CSoutput.n145 gnd 0.856782f
C5128 CSoutput.n146 gnd 0.856782f
C5129 CSoutput.t211 gnd 1.07098f
C5130 CSoutput.n147 gnd 0.856782f
C5131 CSoutput.n148 gnd 0.856782f
C5132 CSoutput.n152 gnd 0.856782f
C5133 CSoutput.n156 gnd 0.856782f
C5134 CSoutput.n157 gnd 0.856782f
C5135 CSoutput.n159 gnd 0.856782f
C5136 CSoutput.n164 gnd 0.856782f
C5137 CSoutput.n166 gnd 0.856782f
C5138 CSoutput.n167 gnd 0.856782f
C5139 CSoutput.n169 gnd 0.856782f
C5140 CSoutput.n170 gnd 0.856782f
C5141 CSoutput.n172 gnd 0.856782f
C5142 CSoutput.t204 gnd 14.3167f
C5143 CSoutput.n174 gnd 0.856782f
C5144 CSoutput.n175 gnd 0.642586f
C5145 CSoutput.n176 gnd 0.856782f
C5146 CSoutput.n177 gnd 0.856782f
C5147 CSoutput.n178 gnd 2.30672f
C5148 CSoutput.n179 gnd 0.856782f
C5149 CSoutput.n180 gnd 0.856782f
C5150 CSoutput.t220 gnd 1.07098f
C5151 CSoutput.n181 gnd 0.856782f
C5152 CSoutput.n182 gnd 0.856782f
C5153 CSoutput.n186 gnd 0.856782f
C5154 CSoutput.n190 gnd 0.856782f
C5155 CSoutput.n191 gnd 0.856782f
C5156 CSoutput.n193 gnd 0.856782f
C5157 CSoutput.n198 gnd 0.856782f
C5158 CSoutput.n200 gnd 0.856782f
C5159 CSoutput.n201 gnd 0.856782f
C5160 CSoutput.n203 gnd 0.856782f
C5161 CSoutput.n204 gnd 0.856782f
C5162 CSoutput.n206 gnd 0.856782f
C5163 CSoutput.n207 gnd 0.642586f
C5164 CSoutput.n209 gnd 0.856782f
C5165 CSoutput.n210 gnd 0.642586f
C5166 CSoutput.n211 gnd 0.856782f
C5167 CSoutput.n212 gnd 0.856782f
C5168 CSoutput.n213 gnd 2.30672f
C5169 CSoutput.n214 gnd 0.856782f
C5170 CSoutput.n215 gnd 0.856782f
C5171 CSoutput.t214 gnd 1.07098f
C5172 CSoutput.n216 gnd 0.856782f
C5173 CSoutput.n217 gnd 2.30672f
C5174 CSoutput.n219 gnd 0.856782f
C5175 CSoutput.n220 gnd 0.856782f
C5176 CSoutput.n222 gnd 0.856782f
C5177 CSoutput.n223 gnd 0.856782f
C5178 CSoutput.t200 gnd 14.0834f
C5179 CSoutput.t207 gnd 14.3167f
C5180 CSoutput.n229 gnd 2.68785f
C5181 CSoutput.n230 gnd 10.9493f
C5182 CSoutput.n231 gnd 11.4075f
C5183 CSoutput.n236 gnd 2.91167f
C5184 CSoutput.n242 gnd 0.856782f
C5185 CSoutput.n244 gnd 0.856782f
C5186 CSoutput.n246 gnd 0.856782f
C5187 CSoutput.n248 gnd 0.856782f
C5188 CSoutput.n250 gnd 0.856782f
C5189 CSoutput.n256 gnd 0.856782f
C5190 CSoutput.n263 gnd 1.57187f
C5191 CSoutput.n264 gnd 1.57186f
C5192 CSoutput.n265 gnd 0.856782f
C5193 CSoutput.n266 gnd 0.856782f
C5194 CSoutput.n268 gnd 0.642586f
C5195 CSoutput.n269 gnd 0.550318f
C5196 CSoutput.n271 gnd 0.642586f
C5197 CSoutput.n272 gnd 0.550318f
C5198 CSoutput.n273 gnd 0.642586f
C5199 CSoutput.n275 gnd 0.856782f
C5200 CSoutput.n277 gnd 2.30672f
C5201 CSoutput.n278 gnd 2.68785f
C5202 CSoutput.n279 gnd 10.0706f
C5203 CSoutput.n281 gnd 0.642586f
C5204 CSoutput.n282 gnd 1.65341f
C5205 CSoutput.n283 gnd 0.642586f
C5206 CSoutput.n285 gnd 0.856782f
C5207 CSoutput.n287 gnd 2.30672f
C5208 CSoutput.n288 gnd 5.02441f
C5209 CSoutput.t39 gnd 0.060414f
C5210 CSoutput.t81 gnd 0.060414f
C5211 CSoutput.n289 gnd 0.467746f
C5212 CSoutput.t70 gnd 0.060414f
C5213 CSoutput.t2 gnd 0.060414f
C5214 CSoutput.n290 gnd 0.466912f
C5215 CSoutput.n291 gnd 0.473915f
C5216 CSoutput.t11 gnd 0.060414f
C5217 CSoutput.t197 gnd 0.060414f
C5218 CSoutput.n292 gnd 0.466912f
C5219 CSoutput.n293 gnd 0.233525f
C5220 CSoutput.t51 gnd 0.060414f
C5221 CSoutput.t55 gnd 0.060414f
C5222 CSoutput.n294 gnd 0.466912f
C5223 CSoutput.n295 gnd 0.233525f
C5224 CSoutput.t36 gnd 0.060414f
C5225 CSoutput.t33 gnd 0.060414f
C5226 CSoutput.n296 gnd 0.466912f
C5227 CSoutput.n297 gnd 0.233525f
C5228 CSoutput.t47 gnd 0.060414f
C5229 CSoutput.t44 gnd 0.060414f
C5230 CSoutput.n298 gnd 0.466912f
C5231 CSoutput.n299 gnd 0.233525f
C5232 CSoutput.t97 gnd 0.060414f
C5233 CSoutput.t195 gnd 0.060414f
C5234 CSoutput.n300 gnd 0.466912f
C5235 CSoutput.n301 gnd 0.233525f
C5236 CSoutput.t86 gnd 0.060414f
C5237 CSoutput.t34 gnd 0.060414f
C5238 CSoutput.n302 gnd 0.466912f
C5239 CSoutput.n303 gnd 0.233525f
C5240 CSoutput.t27 gnd 0.060414f
C5241 CSoutput.t15 gnd 0.060414f
C5242 CSoutput.n304 gnd 0.466912f
C5243 CSoutput.n305 gnd 0.233525f
C5244 CSoutput.t54 gnd 0.060414f
C5245 CSoutput.t58 gnd 0.060414f
C5246 CSoutput.n306 gnd 0.466912f
C5247 CSoutput.n307 gnd 0.428232f
C5248 CSoutput.t17 gnd 0.060414f
C5249 CSoutput.t85 gnd 0.060414f
C5250 CSoutput.n308 gnd 0.467746f
C5251 CSoutput.t59 gnd 0.060414f
C5252 CSoutput.t23 gnd 0.060414f
C5253 CSoutput.n309 gnd 0.466912f
C5254 CSoutput.n310 gnd 0.473915f
C5255 CSoutput.t1 gnd 0.060414f
C5256 CSoutput.t42 gnd 0.060414f
C5257 CSoutput.n311 gnd 0.466912f
C5258 CSoutput.n312 gnd 0.233525f
C5259 CSoutput.t38 gnd 0.060414f
C5260 CSoutput.t198 gnd 0.060414f
C5261 CSoutput.n313 gnd 0.466912f
C5262 CSoutput.n314 gnd 0.233525f
C5263 CSoutput.t66 gnd 0.060414f
C5264 CSoutput.t26 gnd 0.060414f
C5265 CSoutput.n315 gnd 0.466912f
C5266 CSoutput.n316 gnd 0.233525f
C5267 CSoutput.t67 gnd 0.060414f
C5268 CSoutput.t96 gnd 0.060414f
C5269 CSoutput.n317 gnd 0.466912f
C5270 CSoutput.n318 gnd 0.233525f
C5271 CSoutput.t25 gnd 0.060414f
C5272 CSoutput.t77 gnd 0.060414f
C5273 CSoutput.n319 gnd 0.466912f
C5274 CSoutput.n320 gnd 0.233525f
C5275 CSoutput.t90 gnd 0.060414f
C5276 CSoutput.t20 gnd 0.060414f
C5277 CSoutput.n321 gnd 0.466912f
C5278 CSoutput.n322 gnd 0.233525f
C5279 CSoutput.t29 gnd 0.060414f
C5280 CSoutput.t35 gnd 0.060414f
C5281 CSoutput.n323 gnd 0.466912f
C5282 CSoutput.n324 gnd 0.233525f
C5283 CSoutput.t57 gnd 0.060414f
C5284 CSoutput.t53 gnd 0.060414f
C5285 CSoutput.n325 gnd 0.466912f
C5286 CSoutput.n326 gnd 0.348245f
C5287 CSoutput.n327 gnd 0.439135f
C5288 CSoutput.t98 gnd 0.060414f
C5289 CSoutput.t46 gnd 0.060414f
C5290 CSoutput.n328 gnd 0.467746f
C5291 CSoutput.t191 gnd 0.060414f
C5292 CSoutput.t6 gnd 0.060414f
C5293 CSoutput.n329 gnd 0.466912f
C5294 CSoutput.n330 gnd 0.473915f
C5295 CSoutput.t12 gnd 0.060414f
C5296 CSoutput.t188 gnd 0.060414f
C5297 CSoutput.n331 gnd 0.466912f
C5298 CSoutput.n332 gnd 0.233525f
C5299 CSoutput.t7 gnd 0.060414f
C5300 CSoutput.t22 gnd 0.060414f
C5301 CSoutput.n333 gnd 0.466912f
C5302 CSoutput.n334 gnd 0.233525f
C5303 CSoutput.t76 gnd 0.060414f
C5304 CSoutput.t82 gnd 0.060414f
C5305 CSoutput.n335 gnd 0.466912f
C5306 CSoutput.n336 gnd 0.233525f
C5307 CSoutput.t30 gnd 0.060414f
C5308 CSoutput.t88 gnd 0.060414f
C5309 CSoutput.n337 gnd 0.466912f
C5310 CSoutput.n338 gnd 0.233525f
C5311 CSoutput.t75 gnd 0.060414f
C5312 CSoutput.t189 gnd 0.060414f
C5313 CSoutput.n339 gnd 0.466912f
C5314 CSoutput.n340 gnd 0.233525f
C5315 CSoutput.t95 gnd 0.060414f
C5316 CSoutput.t74 gnd 0.060414f
C5317 CSoutput.n341 gnd 0.466912f
C5318 CSoutput.n342 gnd 0.233525f
C5319 CSoutput.t84 gnd 0.060414f
C5320 CSoutput.t13 gnd 0.060414f
C5321 CSoutput.n343 gnd 0.466912f
C5322 CSoutput.n344 gnd 0.233525f
C5323 CSoutput.t185 gnd 0.060414f
C5324 CSoutput.t87 gnd 0.060414f
C5325 CSoutput.n345 gnd 0.46691f
C5326 CSoutput.n346 gnd 0.348247f
C5327 CSoutput.n347 gnd 0.49084f
C5328 CSoutput.n348 gnd 13.6516f
C5329 CSoutput.t159 gnd 0.052862f
C5330 CSoutput.t140 gnd 0.052862f
C5331 CSoutput.n349 gnd 0.468673f
C5332 CSoutput.t144 gnd 0.052862f
C5333 CSoutput.t146 gnd 0.052862f
C5334 CSoutput.n350 gnd 0.46711f
C5335 CSoutput.n351 gnd 0.435259f
C5336 CSoutput.t131 gnd 0.052862f
C5337 CSoutput.t175 gnd 0.052862f
C5338 CSoutput.n352 gnd 0.46711f
C5339 CSoutput.n353 gnd 0.214562f
C5340 CSoutput.t111 gnd 0.052862f
C5341 CSoutput.t160 gnd 0.052862f
C5342 CSoutput.n354 gnd 0.46711f
C5343 CSoutput.n355 gnd 0.214562f
C5344 CSoutput.t102 gnd 0.052862f
C5345 CSoutput.t126 gnd 0.052862f
C5346 CSoutput.n356 gnd 0.46711f
C5347 CSoutput.n357 gnd 0.214562f
C5348 CSoutput.t105 gnd 0.052862f
C5349 CSoutput.t116 gnd 0.052862f
C5350 CSoutput.n358 gnd 0.46711f
C5351 CSoutput.n359 gnd 0.214562f
C5352 CSoutput.t154 gnd 0.052862f
C5353 CSoutput.t137 gnd 0.052862f
C5354 CSoutput.n360 gnd 0.46711f
C5355 CSoutput.n361 gnd 0.214562f
C5356 CSoutput.t141 gnd 0.052862f
C5357 CSoutput.t101 gnd 0.052862f
C5358 CSoutput.n362 gnd 0.46711f
C5359 CSoutput.n363 gnd 0.214562f
C5360 CSoutput.t127 gnd 0.052862f
C5361 CSoutput.t149 gnd 0.052862f
C5362 CSoutput.n364 gnd 0.46711f
C5363 CSoutput.n365 gnd 0.214562f
C5364 CSoutput.t110 gnd 0.052862f
C5365 CSoutput.t156 gnd 0.052862f
C5366 CSoutput.n366 gnd 0.46711f
C5367 CSoutput.n367 gnd 0.395696f
C5368 CSoutput.t118 gnd 0.052862f
C5369 CSoutput.t155 gnd 0.052862f
C5370 CSoutput.n368 gnd 0.468673f
C5371 CSoutput.t113 gnd 0.052862f
C5372 CSoutput.t151 gnd 0.052862f
C5373 CSoutput.n369 gnd 0.46711f
C5374 CSoutput.n370 gnd 0.435259f
C5375 CSoutput.t103 gnd 0.052862f
C5376 CSoutput.t128 gnd 0.052862f
C5377 CSoutput.n371 gnd 0.46711f
C5378 CSoutput.n372 gnd 0.214562f
C5379 CSoutput.t170 gnd 0.052862f
C5380 CSoutput.t119 gnd 0.052862f
C5381 CSoutput.n373 gnd 0.46711f
C5382 CSoutput.n374 gnd 0.214562f
C5383 CSoutput.t122 gnd 0.052862f
C5384 CSoutput.t163 gnd 0.052862f
C5385 CSoutput.n375 gnd 0.46711f
C5386 CSoutput.n376 gnd 0.214562f
C5387 CSoutput.t142 gnd 0.052862f
C5388 CSoutput.t145 gnd 0.052862f
C5389 CSoutput.n377 gnd 0.46711f
C5390 CSoutput.n378 gnd 0.214562f
C5391 CSoutput.t115 gnd 0.052862f
C5392 CSoutput.t150 gnd 0.052862f
C5393 CSoutput.n379 gnd 0.46711f
C5394 CSoutput.n380 gnd 0.214562f
C5395 CSoutput.t109 gnd 0.052862f
C5396 CSoutput.t121 gnd 0.052862f
C5397 CSoutput.n381 gnd 0.46711f
C5398 CSoutput.n382 gnd 0.214562f
C5399 CSoutput.t100 gnd 0.052862f
C5400 CSoutput.t178 gnd 0.052862f
C5401 CSoutput.n383 gnd 0.46711f
C5402 CSoutput.n384 gnd 0.214562f
C5403 CSoutput.t168 gnd 0.052862f
C5404 CSoutput.t117 gnd 0.052862f
C5405 CSoutput.n385 gnd 0.46711f
C5406 CSoutput.n386 gnd 0.325752f
C5407 CSoutput.n387 gnd 0.605271f
C5408 CSoutput.n388 gnd 14.1857f
C5409 CSoutput.t167 gnd 0.052862f
C5410 CSoutput.t135 gnd 0.052862f
C5411 CSoutput.n389 gnd 0.468673f
C5412 CSoutput.t107 gnd 0.052862f
C5413 CSoutput.t108 gnd 0.052862f
C5414 CSoutput.n390 gnd 0.46711f
C5415 CSoutput.n391 gnd 0.435259f
C5416 CSoutput.t114 gnd 0.052862f
C5417 CSoutput.t174 gnd 0.052862f
C5418 CSoutput.n392 gnd 0.46711f
C5419 CSoutput.n393 gnd 0.214562f
C5420 CSoutput.t136 gnd 0.052862f
C5421 CSoutput.t164 gnd 0.052862f
C5422 CSoutput.n394 gnd 0.46711f
C5423 CSoutput.n395 gnd 0.214562f
C5424 CSoutput.t172 gnd 0.052862f
C5425 CSoutput.t124 gnd 0.052862f
C5426 CSoutput.n396 gnd 0.46711f
C5427 CSoutput.n397 gnd 0.214562f
C5428 CSoutput.t132 gnd 0.052862f
C5429 CSoutput.t157 gnd 0.052862f
C5430 CSoutput.n398 gnd 0.46711f
C5431 CSoutput.n399 gnd 0.214562f
C5432 CSoutput.t165 gnd 0.052862f
C5433 CSoutput.t177 gnd 0.052862f
C5434 CSoutput.n400 gnd 0.46711f
C5435 CSoutput.n401 gnd 0.214562f
C5436 CSoutput.t123 gnd 0.052862f
C5437 CSoutput.t162 gnd 0.052862f
C5438 CSoutput.n402 gnd 0.46711f
C5439 CSoutput.n403 gnd 0.214562f
C5440 CSoutput.t112 gnd 0.052862f
C5441 CSoutput.t173 gnd 0.052862f
C5442 CSoutput.n404 gnd 0.46711f
C5443 CSoutput.n405 gnd 0.214562f
C5444 CSoutput.t130 gnd 0.052862f
C5445 CSoutput.t147 gnd 0.052862f
C5446 CSoutput.n406 gnd 0.46711f
C5447 CSoutput.n407 gnd 0.395696f
C5448 CSoutput.t134 gnd 0.052862f
C5449 CSoutput.t133 gnd 0.052862f
C5450 CSoutput.n408 gnd 0.468673f
C5451 CSoutput.t143 gnd 0.052862f
C5452 CSoutput.t166 gnd 0.052862f
C5453 CSoutput.n409 gnd 0.46711f
C5454 CSoutput.n410 gnd 0.435259f
C5455 CSoutput.t169 gnd 0.052862f
C5456 CSoutput.t125 gnd 0.052862f
C5457 CSoutput.n411 gnd 0.46711f
C5458 CSoutput.n412 gnd 0.214562f
C5459 CSoutput.t153 gnd 0.052862f
C5460 CSoutput.t176 gnd 0.052862f
C5461 CSoutput.n413 gnd 0.46711f
C5462 CSoutput.n414 gnd 0.214562f
C5463 CSoutput.t138 gnd 0.052862f
C5464 CSoutput.t161 gnd 0.052862f
C5465 CSoutput.n415 gnd 0.46711f
C5466 CSoutput.n416 gnd 0.214562f
C5467 CSoutput.t106 gnd 0.052862f
C5468 CSoutput.t148 gnd 0.052862f
C5469 CSoutput.n417 gnd 0.46711f
C5470 CSoutput.n418 gnd 0.214562f
C5471 CSoutput.t179 gnd 0.052862f
C5472 CSoutput.t129 gnd 0.052862f
C5473 CSoutput.n419 gnd 0.46711f
C5474 CSoutput.n420 gnd 0.214562f
C5475 CSoutput.t158 gnd 0.052862f
C5476 CSoutput.t120 gnd 0.052862f
C5477 CSoutput.n421 gnd 0.46711f
C5478 CSoutput.n422 gnd 0.214562f
C5479 CSoutput.t171 gnd 0.052862f
C5480 CSoutput.t139 gnd 0.052862f
C5481 CSoutput.n423 gnd 0.46711f
C5482 CSoutput.n424 gnd 0.214562f
C5483 CSoutput.t104 gnd 0.052862f
C5484 CSoutput.t152 gnd 0.052862f
C5485 CSoutput.n425 gnd 0.46711f
C5486 CSoutput.n426 gnd 0.325752f
C5487 CSoutput.n427 gnd 0.605271f
C5488 CSoutput.n428 gnd 8.51017f
C5489 CSoutput.n429 gnd 15.605599f
C5490 commonsourceibias.n0 gnd 0.010705f
C5491 commonsourceibias.t117 gnd 0.162096f
C5492 commonsourceibias.t135 gnd 0.149881f
C5493 commonsourceibias.n1 gnd 0.007808f
C5494 commonsourceibias.n2 gnd 0.008022f
C5495 commonsourceibias.t92 gnd 0.149881f
C5496 commonsourceibias.n3 gnd 0.010321f
C5497 commonsourceibias.n4 gnd 0.008022f
C5498 commonsourceibias.t90 gnd 0.149881f
C5499 commonsourceibias.n5 gnd 0.059802f
C5500 commonsourceibias.t127 gnd 0.149881f
C5501 commonsourceibias.n6 gnd 0.007564f
C5502 commonsourceibias.n7 gnd 0.008022f
C5503 commonsourceibias.t145 gnd 0.149881f
C5504 commonsourceibias.n8 gnd 0.010168f
C5505 commonsourceibias.n9 gnd 0.008022f
C5506 commonsourceibias.t83 gnd 0.149881f
C5507 commonsourceibias.n10 gnd 0.059802f
C5508 commonsourceibias.t116 gnd 0.149881f
C5509 commonsourceibias.n11 gnd 0.007348f
C5510 commonsourceibias.n12 gnd 0.008022f
C5511 commonsourceibias.t110 gnd 0.149881f
C5512 commonsourceibias.n13 gnd 0.009997f
C5513 commonsourceibias.n14 gnd 0.010705f
C5514 commonsourceibias.t22 gnd 0.162096f
C5515 commonsourceibias.t74 gnd 0.149881f
C5516 commonsourceibias.n15 gnd 0.007808f
C5517 commonsourceibias.n16 gnd 0.008022f
C5518 commonsourceibias.t4 gnd 0.149881f
C5519 commonsourceibias.n17 gnd 0.010321f
C5520 commonsourceibias.n18 gnd 0.008022f
C5521 commonsourceibias.t20 gnd 0.149881f
C5522 commonsourceibias.n19 gnd 0.059802f
C5523 commonsourceibias.t28 gnd 0.149881f
C5524 commonsourceibias.n20 gnd 0.007564f
C5525 commonsourceibias.n21 gnd 0.008022f
C5526 commonsourceibias.t40 gnd 0.149881f
C5527 commonsourceibias.n22 gnd 0.010168f
C5528 commonsourceibias.n23 gnd 0.008022f
C5529 commonsourceibias.t10 gnd 0.149881f
C5530 commonsourceibias.n24 gnd 0.059802f
C5531 commonsourceibias.t16 gnd 0.149881f
C5532 commonsourceibias.n25 gnd 0.007348f
C5533 commonsourceibias.n26 gnd 0.008022f
C5534 commonsourceibias.t24 gnd 0.149881f
C5535 commonsourceibias.n27 gnd 0.009997f
C5536 commonsourceibias.n28 gnd 0.008022f
C5537 commonsourceibias.t68 gnd 0.149881f
C5538 commonsourceibias.n29 gnd 0.059802f
C5539 commonsourceibias.t50 gnd 0.149881f
C5540 commonsourceibias.n30 gnd 0.007159f
C5541 commonsourceibias.n31 gnd 0.008022f
C5542 commonsourceibias.t12 gnd 0.149881f
C5543 commonsourceibias.n32 gnd 0.009806f
C5544 commonsourceibias.n33 gnd 0.008022f
C5545 commonsourceibias.t38 gnd 0.149881f
C5546 commonsourceibias.n34 gnd 0.059802f
C5547 commonsourceibias.t42 gnd 0.149881f
C5548 commonsourceibias.n35 gnd 0.006995f
C5549 commonsourceibias.n36 gnd 0.008022f
C5550 commonsourceibias.t76 gnd 0.149881f
C5551 commonsourceibias.n37 gnd 0.009595f
C5552 commonsourceibias.n38 gnd 0.008022f
C5553 commonsourceibias.t0 gnd 0.149881f
C5554 commonsourceibias.n39 gnd 0.059802f
C5555 commonsourceibias.t54 gnd 0.149881f
C5556 commonsourceibias.n40 gnd 0.006855f
C5557 commonsourceibias.n41 gnd 0.008022f
C5558 commonsourceibias.t66 gnd 0.149881f
C5559 commonsourceibias.n42 gnd 0.00936f
C5560 commonsourceibias.t46 gnd 0.16664f
C5561 commonsourceibias.t72 gnd 0.149881f
C5562 commonsourceibias.n43 gnd 0.065328f
C5563 commonsourceibias.n44 gnd 0.07169f
C5564 commonsourceibias.n45 gnd 0.033265f
C5565 commonsourceibias.n46 gnd 0.008022f
C5566 commonsourceibias.n47 gnd 0.007808f
C5567 commonsourceibias.n48 gnd 0.01119f
C5568 commonsourceibias.n49 gnd 0.059802f
C5569 commonsourceibias.n50 gnd 0.011182f
C5570 commonsourceibias.n51 gnd 0.008022f
C5571 commonsourceibias.n52 gnd 0.008022f
C5572 commonsourceibias.n53 gnd 0.008022f
C5573 commonsourceibias.n54 gnd 0.010321f
C5574 commonsourceibias.n55 gnd 0.059802f
C5575 commonsourceibias.n56 gnd 0.010563f
C5576 commonsourceibias.n57 gnd 0.010263f
C5577 commonsourceibias.n58 gnd 0.008022f
C5578 commonsourceibias.n59 gnd 0.008022f
C5579 commonsourceibias.n60 gnd 0.008022f
C5580 commonsourceibias.n61 gnd 0.007564f
C5581 commonsourceibias.n62 gnd 0.0112f
C5582 commonsourceibias.n63 gnd 0.059802f
C5583 commonsourceibias.n64 gnd 0.011196f
C5584 commonsourceibias.n65 gnd 0.008022f
C5585 commonsourceibias.n66 gnd 0.008022f
C5586 commonsourceibias.n67 gnd 0.008022f
C5587 commonsourceibias.n68 gnd 0.010168f
C5588 commonsourceibias.n69 gnd 0.059802f
C5589 commonsourceibias.n70 gnd 0.010488f
C5590 commonsourceibias.n71 gnd 0.010338f
C5591 commonsourceibias.n72 gnd 0.008022f
C5592 commonsourceibias.n73 gnd 0.008022f
C5593 commonsourceibias.n74 gnd 0.008022f
C5594 commonsourceibias.n75 gnd 0.007348f
C5595 commonsourceibias.n76 gnd 0.011204f
C5596 commonsourceibias.n77 gnd 0.059802f
C5597 commonsourceibias.n78 gnd 0.011203f
C5598 commonsourceibias.n79 gnd 0.008022f
C5599 commonsourceibias.n80 gnd 0.008022f
C5600 commonsourceibias.n81 gnd 0.008022f
C5601 commonsourceibias.n82 gnd 0.009997f
C5602 commonsourceibias.n83 gnd 0.059802f
C5603 commonsourceibias.n84 gnd 0.010413f
C5604 commonsourceibias.n85 gnd 0.010413f
C5605 commonsourceibias.n86 gnd 0.008022f
C5606 commonsourceibias.n87 gnd 0.008022f
C5607 commonsourceibias.n88 gnd 0.008022f
C5608 commonsourceibias.n89 gnd 0.007159f
C5609 commonsourceibias.n90 gnd 0.011203f
C5610 commonsourceibias.n91 gnd 0.059802f
C5611 commonsourceibias.n92 gnd 0.011204f
C5612 commonsourceibias.n93 gnd 0.008022f
C5613 commonsourceibias.n94 gnd 0.008022f
C5614 commonsourceibias.n95 gnd 0.008022f
C5615 commonsourceibias.n96 gnd 0.009806f
C5616 commonsourceibias.n97 gnd 0.059802f
C5617 commonsourceibias.n98 gnd 0.010338f
C5618 commonsourceibias.n99 gnd 0.010488f
C5619 commonsourceibias.n100 gnd 0.008022f
C5620 commonsourceibias.n101 gnd 0.008022f
C5621 commonsourceibias.n102 gnd 0.008022f
C5622 commonsourceibias.n103 gnd 0.006995f
C5623 commonsourceibias.n104 gnd 0.011196f
C5624 commonsourceibias.n105 gnd 0.059802f
C5625 commonsourceibias.n106 gnd 0.0112f
C5626 commonsourceibias.n107 gnd 0.008022f
C5627 commonsourceibias.n108 gnd 0.008022f
C5628 commonsourceibias.n109 gnd 0.008022f
C5629 commonsourceibias.n110 gnd 0.009595f
C5630 commonsourceibias.n111 gnd 0.059802f
C5631 commonsourceibias.n112 gnd 0.010263f
C5632 commonsourceibias.n113 gnd 0.010563f
C5633 commonsourceibias.n114 gnd 0.008022f
C5634 commonsourceibias.n115 gnd 0.008022f
C5635 commonsourceibias.n116 gnd 0.008022f
C5636 commonsourceibias.n117 gnd 0.006855f
C5637 commonsourceibias.n118 gnd 0.011182f
C5638 commonsourceibias.n119 gnd 0.059802f
C5639 commonsourceibias.n120 gnd 0.01119f
C5640 commonsourceibias.n121 gnd 0.008022f
C5641 commonsourceibias.n122 gnd 0.008022f
C5642 commonsourceibias.n123 gnd 0.008022f
C5643 commonsourceibias.n124 gnd 0.00936f
C5644 commonsourceibias.n125 gnd 0.059802f
C5645 commonsourceibias.n126 gnd 0.009843f
C5646 commonsourceibias.n127 gnd 0.071758f
C5647 commonsourceibias.n128 gnd 0.079928f
C5648 commonsourceibias.t23 gnd 0.017311f
C5649 commonsourceibias.t75 gnd 0.017311f
C5650 commonsourceibias.n129 gnd 0.152968f
C5651 commonsourceibias.n130 gnd 0.132319f
C5652 commonsourceibias.t5 gnd 0.017311f
C5653 commonsourceibias.t21 gnd 0.017311f
C5654 commonsourceibias.n131 gnd 0.152968f
C5655 commonsourceibias.n132 gnd 0.070264f
C5656 commonsourceibias.t29 gnd 0.017311f
C5657 commonsourceibias.t41 gnd 0.017311f
C5658 commonsourceibias.n133 gnd 0.152968f
C5659 commonsourceibias.n134 gnd 0.070264f
C5660 commonsourceibias.t11 gnd 0.017311f
C5661 commonsourceibias.t17 gnd 0.017311f
C5662 commonsourceibias.n135 gnd 0.152968f
C5663 commonsourceibias.n136 gnd 0.070264f
C5664 commonsourceibias.t25 gnd 0.017311f
C5665 commonsourceibias.t69 gnd 0.017311f
C5666 commonsourceibias.n137 gnd 0.152968f
C5667 commonsourceibias.n138 gnd 0.058702f
C5668 commonsourceibias.t73 gnd 0.017311f
C5669 commonsourceibias.t47 gnd 0.017311f
C5670 commonsourceibias.n139 gnd 0.15348f
C5671 commonsourceibias.t55 gnd 0.017311f
C5672 commonsourceibias.t67 gnd 0.017311f
C5673 commonsourceibias.n140 gnd 0.152968f
C5674 commonsourceibias.n141 gnd 0.142538f
C5675 commonsourceibias.t77 gnd 0.017311f
C5676 commonsourceibias.t1 gnd 0.017311f
C5677 commonsourceibias.n142 gnd 0.152968f
C5678 commonsourceibias.n143 gnd 0.070264f
C5679 commonsourceibias.t39 gnd 0.017311f
C5680 commonsourceibias.t43 gnd 0.017311f
C5681 commonsourceibias.n144 gnd 0.152968f
C5682 commonsourceibias.n145 gnd 0.070264f
C5683 commonsourceibias.t51 gnd 0.017311f
C5684 commonsourceibias.t13 gnd 0.017311f
C5685 commonsourceibias.n146 gnd 0.152968f
C5686 commonsourceibias.n147 gnd 0.058702f
C5687 commonsourceibias.n148 gnd 0.071082f
C5688 commonsourceibias.n149 gnd 0.05192f
C5689 commonsourceibias.t131 gnd 0.149881f
C5690 commonsourceibias.n150 gnd 0.059802f
C5691 commonsourceibias.t107 gnd 0.149881f
C5692 commonsourceibias.n151 gnd 0.059802f
C5693 commonsourceibias.n152 gnd 0.008022f
C5694 commonsourceibias.t103 gnd 0.149881f
C5695 commonsourceibias.n153 gnd 0.059802f
C5696 commonsourceibias.n154 gnd 0.008022f
C5697 commonsourceibias.t121 gnd 0.149881f
C5698 commonsourceibias.n155 gnd 0.059802f
C5699 commonsourceibias.n156 gnd 0.008022f
C5700 commonsourceibias.t138 gnd 0.149881f
C5701 commonsourceibias.n157 gnd 0.006995f
C5702 commonsourceibias.n158 gnd 0.008022f
C5703 commonsourceibias.t95 gnd 0.149881f
C5704 commonsourceibias.n159 gnd 0.009595f
C5705 commonsourceibias.n160 gnd 0.008022f
C5706 commonsourceibias.t111 gnd 0.149881f
C5707 commonsourceibias.n161 gnd 0.059802f
C5708 commonsourceibias.t130 gnd 0.149881f
C5709 commonsourceibias.n162 gnd 0.006855f
C5710 commonsourceibias.n163 gnd 0.008022f
C5711 commonsourceibias.t87 gnd 0.149881f
C5712 commonsourceibias.n164 gnd 0.00936f
C5713 commonsourceibias.t119 gnd 0.16664f
C5714 commonsourceibias.t84 gnd 0.149881f
C5715 commonsourceibias.n165 gnd 0.065328f
C5716 commonsourceibias.n166 gnd 0.07169f
C5717 commonsourceibias.n167 gnd 0.033265f
C5718 commonsourceibias.n168 gnd 0.008022f
C5719 commonsourceibias.n169 gnd 0.007808f
C5720 commonsourceibias.n170 gnd 0.01119f
C5721 commonsourceibias.n171 gnd 0.059802f
C5722 commonsourceibias.n172 gnd 0.011182f
C5723 commonsourceibias.n173 gnd 0.008022f
C5724 commonsourceibias.n174 gnd 0.008022f
C5725 commonsourceibias.n175 gnd 0.008022f
C5726 commonsourceibias.n176 gnd 0.010321f
C5727 commonsourceibias.n177 gnd 0.059802f
C5728 commonsourceibias.n178 gnd 0.010563f
C5729 commonsourceibias.n179 gnd 0.010263f
C5730 commonsourceibias.n180 gnd 0.008022f
C5731 commonsourceibias.n181 gnd 0.008022f
C5732 commonsourceibias.n182 gnd 0.008022f
C5733 commonsourceibias.n183 gnd 0.007564f
C5734 commonsourceibias.n184 gnd 0.0112f
C5735 commonsourceibias.n185 gnd 0.059802f
C5736 commonsourceibias.n186 gnd 0.011196f
C5737 commonsourceibias.n187 gnd 0.008022f
C5738 commonsourceibias.n188 gnd 0.008022f
C5739 commonsourceibias.n189 gnd 0.008022f
C5740 commonsourceibias.n190 gnd 0.010168f
C5741 commonsourceibias.n191 gnd 0.059802f
C5742 commonsourceibias.n192 gnd 0.010488f
C5743 commonsourceibias.n193 gnd 0.010338f
C5744 commonsourceibias.n194 gnd 0.008022f
C5745 commonsourceibias.n195 gnd 0.008022f
C5746 commonsourceibias.n196 gnd 0.009806f
C5747 commonsourceibias.n197 gnd 0.007348f
C5748 commonsourceibias.n198 gnd 0.011204f
C5749 commonsourceibias.n199 gnd 0.008022f
C5750 commonsourceibias.n200 gnd 0.008022f
C5751 commonsourceibias.n201 gnd 0.011203f
C5752 commonsourceibias.n202 gnd 0.007159f
C5753 commonsourceibias.n203 gnd 0.009997f
C5754 commonsourceibias.n204 gnd 0.008022f
C5755 commonsourceibias.n205 gnd 0.007008f
C5756 commonsourceibias.n206 gnd 0.010413f
C5757 commonsourceibias.n207 gnd 0.010413f
C5758 commonsourceibias.n208 gnd 0.007008f
C5759 commonsourceibias.n209 gnd 0.008022f
C5760 commonsourceibias.n210 gnd 0.008022f
C5761 commonsourceibias.n211 gnd 0.007159f
C5762 commonsourceibias.n212 gnd 0.011203f
C5763 commonsourceibias.n213 gnd 0.059802f
C5764 commonsourceibias.n214 gnd 0.011204f
C5765 commonsourceibias.n215 gnd 0.008022f
C5766 commonsourceibias.n216 gnd 0.008022f
C5767 commonsourceibias.n217 gnd 0.008022f
C5768 commonsourceibias.n218 gnd 0.009806f
C5769 commonsourceibias.n219 gnd 0.059802f
C5770 commonsourceibias.n220 gnd 0.010338f
C5771 commonsourceibias.n221 gnd 0.010488f
C5772 commonsourceibias.n222 gnd 0.008022f
C5773 commonsourceibias.n223 gnd 0.008022f
C5774 commonsourceibias.n224 gnd 0.008022f
C5775 commonsourceibias.n225 gnd 0.006995f
C5776 commonsourceibias.n226 gnd 0.011196f
C5777 commonsourceibias.n227 gnd 0.059802f
C5778 commonsourceibias.n228 gnd 0.0112f
C5779 commonsourceibias.n229 gnd 0.008022f
C5780 commonsourceibias.n230 gnd 0.008022f
C5781 commonsourceibias.n231 gnd 0.008022f
C5782 commonsourceibias.n232 gnd 0.009595f
C5783 commonsourceibias.n233 gnd 0.059802f
C5784 commonsourceibias.n234 gnd 0.010263f
C5785 commonsourceibias.n235 gnd 0.010563f
C5786 commonsourceibias.n236 gnd 0.008022f
C5787 commonsourceibias.n237 gnd 0.008022f
C5788 commonsourceibias.n238 gnd 0.008022f
C5789 commonsourceibias.n239 gnd 0.006855f
C5790 commonsourceibias.n240 gnd 0.011182f
C5791 commonsourceibias.n241 gnd 0.059802f
C5792 commonsourceibias.n242 gnd 0.01119f
C5793 commonsourceibias.n243 gnd 0.008022f
C5794 commonsourceibias.n244 gnd 0.008022f
C5795 commonsourceibias.n245 gnd 0.008022f
C5796 commonsourceibias.n246 gnd 0.00936f
C5797 commonsourceibias.n247 gnd 0.059802f
C5798 commonsourceibias.n248 gnd 0.009843f
C5799 commonsourceibias.n249 gnd 0.071758f
C5800 commonsourceibias.n250 gnd 0.046883f
C5801 commonsourceibias.n251 gnd 0.010705f
C5802 commonsourceibias.t120 gnd 0.149881f
C5803 commonsourceibias.n252 gnd 0.007808f
C5804 commonsourceibias.n253 gnd 0.008022f
C5805 commonsourceibias.t81 gnd 0.149881f
C5806 commonsourceibias.n254 gnd 0.010321f
C5807 commonsourceibias.n255 gnd 0.008022f
C5808 commonsourceibias.t159 gnd 0.149881f
C5809 commonsourceibias.n256 gnd 0.059802f
C5810 commonsourceibias.t109 gnd 0.149881f
C5811 commonsourceibias.n257 gnd 0.007564f
C5812 commonsourceibias.n258 gnd 0.008022f
C5813 commonsourceibias.t129 gnd 0.149881f
C5814 commonsourceibias.n259 gnd 0.010168f
C5815 commonsourceibias.n260 gnd 0.008022f
C5816 commonsourceibias.t151 gnd 0.149881f
C5817 commonsourceibias.n261 gnd 0.059802f
C5818 commonsourceibias.t100 gnd 0.149881f
C5819 commonsourceibias.n262 gnd 0.007348f
C5820 commonsourceibias.n263 gnd 0.008022f
C5821 commonsourceibias.t96 gnd 0.149881f
C5822 commonsourceibias.n264 gnd 0.009997f
C5823 commonsourceibias.n265 gnd 0.008022f
C5824 commonsourceibias.t113 gnd 0.149881f
C5825 commonsourceibias.n266 gnd 0.059802f
C5826 commonsourceibias.t94 gnd 0.149881f
C5827 commonsourceibias.n267 gnd 0.007159f
C5828 commonsourceibias.n268 gnd 0.008022f
C5829 commonsourceibias.t91 gnd 0.149881f
C5830 commonsourceibias.n269 gnd 0.009806f
C5831 commonsourceibias.n270 gnd 0.008022f
C5832 commonsourceibias.t104 gnd 0.149881f
C5833 commonsourceibias.n271 gnd 0.059802f
C5834 commonsourceibias.t122 gnd 0.149881f
C5835 commonsourceibias.n272 gnd 0.006995f
C5836 commonsourceibias.n273 gnd 0.008022f
C5837 commonsourceibias.t85 gnd 0.149881f
C5838 commonsourceibias.n274 gnd 0.009595f
C5839 commonsourceibias.n275 gnd 0.008022f
C5840 commonsourceibias.t97 gnd 0.149881f
C5841 commonsourceibias.n276 gnd 0.059802f
C5842 commonsourceibias.t112 gnd 0.149881f
C5843 commonsourceibias.n277 gnd 0.006855f
C5844 commonsourceibias.n278 gnd 0.008022f
C5845 commonsourceibias.t157 gnd 0.149881f
C5846 commonsourceibias.n279 gnd 0.00936f
C5847 commonsourceibias.t102 gnd 0.16664f
C5848 commonsourceibias.t152 gnd 0.149881f
C5849 commonsourceibias.n280 gnd 0.065328f
C5850 commonsourceibias.n281 gnd 0.07169f
C5851 commonsourceibias.n282 gnd 0.033265f
C5852 commonsourceibias.n283 gnd 0.008022f
C5853 commonsourceibias.n284 gnd 0.007808f
C5854 commonsourceibias.n285 gnd 0.01119f
C5855 commonsourceibias.n286 gnd 0.059802f
C5856 commonsourceibias.n287 gnd 0.011182f
C5857 commonsourceibias.n288 gnd 0.008022f
C5858 commonsourceibias.n289 gnd 0.008022f
C5859 commonsourceibias.n290 gnd 0.008022f
C5860 commonsourceibias.n291 gnd 0.010321f
C5861 commonsourceibias.n292 gnd 0.059802f
C5862 commonsourceibias.n293 gnd 0.010563f
C5863 commonsourceibias.n294 gnd 0.010263f
C5864 commonsourceibias.n295 gnd 0.008022f
C5865 commonsourceibias.n296 gnd 0.008022f
C5866 commonsourceibias.n297 gnd 0.008022f
C5867 commonsourceibias.n298 gnd 0.007564f
C5868 commonsourceibias.n299 gnd 0.0112f
C5869 commonsourceibias.n300 gnd 0.059802f
C5870 commonsourceibias.n301 gnd 0.011196f
C5871 commonsourceibias.n302 gnd 0.008022f
C5872 commonsourceibias.n303 gnd 0.008022f
C5873 commonsourceibias.n304 gnd 0.008022f
C5874 commonsourceibias.n305 gnd 0.010168f
C5875 commonsourceibias.n306 gnd 0.059802f
C5876 commonsourceibias.n307 gnd 0.010488f
C5877 commonsourceibias.n308 gnd 0.010338f
C5878 commonsourceibias.n309 gnd 0.008022f
C5879 commonsourceibias.n310 gnd 0.008022f
C5880 commonsourceibias.n311 gnd 0.008022f
C5881 commonsourceibias.n312 gnd 0.007348f
C5882 commonsourceibias.n313 gnd 0.011204f
C5883 commonsourceibias.n314 gnd 0.059802f
C5884 commonsourceibias.n315 gnd 0.011203f
C5885 commonsourceibias.n316 gnd 0.008022f
C5886 commonsourceibias.n317 gnd 0.008022f
C5887 commonsourceibias.n318 gnd 0.008022f
C5888 commonsourceibias.n319 gnd 0.009997f
C5889 commonsourceibias.n320 gnd 0.059802f
C5890 commonsourceibias.n321 gnd 0.010413f
C5891 commonsourceibias.n322 gnd 0.010413f
C5892 commonsourceibias.n323 gnd 0.008022f
C5893 commonsourceibias.n324 gnd 0.008022f
C5894 commonsourceibias.n325 gnd 0.008022f
C5895 commonsourceibias.n326 gnd 0.007159f
C5896 commonsourceibias.n327 gnd 0.011203f
C5897 commonsourceibias.n328 gnd 0.059802f
C5898 commonsourceibias.n329 gnd 0.011204f
C5899 commonsourceibias.n330 gnd 0.008022f
C5900 commonsourceibias.n331 gnd 0.008022f
C5901 commonsourceibias.n332 gnd 0.008022f
C5902 commonsourceibias.n333 gnd 0.009806f
C5903 commonsourceibias.n334 gnd 0.059802f
C5904 commonsourceibias.n335 gnd 0.010338f
C5905 commonsourceibias.n336 gnd 0.010488f
C5906 commonsourceibias.n337 gnd 0.008022f
C5907 commonsourceibias.n338 gnd 0.008022f
C5908 commonsourceibias.n339 gnd 0.008022f
C5909 commonsourceibias.n340 gnd 0.006995f
C5910 commonsourceibias.n341 gnd 0.011196f
C5911 commonsourceibias.n342 gnd 0.059802f
C5912 commonsourceibias.n343 gnd 0.0112f
C5913 commonsourceibias.n344 gnd 0.008022f
C5914 commonsourceibias.n345 gnd 0.008022f
C5915 commonsourceibias.n346 gnd 0.008022f
C5916 commonsourceibias.n347 gnd 0.009595f
C5917 commonsourceibias.n348 gnd 0.059802f
C5918 commonsourceibias.n349 gnd 0.010263f
C5919 commonsourceibias.n350 gnd 0.010563f
C5920 commonsourceibias.n351 gnd 0.008022f
C5921 commonsourceibias.n352 gnd 0.008022f
C5922 commonsourceibias.n353 gnd 0.008022f
C5923 commonsourceibias.n354 gnd 0.006855f
C5924 commonsourceibias.n355 gnd 0.011182f
C5925 commonsourceibias.n356 gnd 0.059802f
C5926 commonsourceibias.n357 gnd 0.01119f
C5927 commonsourceibias.n358 gnd 0.008022f
C5928 commonsourceibias.n359 gnd 0.008022f
C5929 commonsourceibias.n360 gnd 0.008022f
C5930 commonsourceibias.n361 gnd 0.00936f
C5931 commonsourceibias.n362 gnd 0.059802f
C5932 commonsourceibias.n363 gnd 0.009843f
C5933 commonsourceibias.t101 gnd 0.162096f
C5934 commonsourceibias.n364 gnd 0.071758f
C5935 commonsourceibias.n365 gnd 0.024957f
C5936 commonsourceibias.n366 gnd 0.404135f
C5937 commonsourceibias.n367 gnd 0.010705f
C5938 commonsourceibias.t140 gnd 0.162096f
C5939 commonsourceibias.t153 gnd 0.149881f
C5940 commonsourceibias.n368 gnd 0.007808f
C5941 commonsourceibias.n369 gnd 0.008022f
C5942 commonsourceibias.t86 gnd 0.149881f
C5943 commonsourceibias.n370 gnd 0.010321f
C5944 commonsourceibias.n371 gnd 0.008022f
C5945 commonsourceibias.t146 gnd 0.149881f
C5946 commonsourceibias.n372 gnd 0.007564f
C5947 commonsourceibias.n373 gnd 0.008022f
C5948 commonsourceibias.t80 gnd 0.149881f
C5949 commonsourceibias.n374 gnd 0.010168f
C5950 commonsourceibias.n375 gnd 0.008022f
C5951 commonsourceibias.t139 gnd 0.149881f
C5952 commonsourceibias.n376 gnd 0.007348f
C5953 commonsourceibias.n377 gnd 0.008022f
C5954 commonsourceibias.t133 gnd 0.149881f
C5955 commonsourceibias.n378 gnd 0.009997f
C5956 commonsourceibias.t37 gnd 0.017311f
C5957 commonsourceibias.t15 gnd 0.017311f
C5958 commonsourceibias.n379 gnd 0.15348f
C5959 commonsourceibias.t7 gnd 0.017311f
C5960 commonsourceibias.t35 gnd 0.017311f
C5961 commonsourceibias.n380 gnd 0.152968f
C5962 commonsourceibias.n381 gnd 0.142538f
C5963 commonsourceibias.t49 gnd 0.017311f
C5964 commonsourceibias.t65 gnd 0.017311f
C5965 commonsourceibias.n382 gnd 0.152968f
C5966 commonsourceibias.n383 gnd 0.070264f
C5967 commonsourceibias.t61 gnd 0.017311f
C5968 commonsourceibias.t3 gnd 0.017311f
C5969 commonsourceibias.n384 gnd 0.152968f
C5970 commonsourceibias.n385 gnd 0.070264f
C5971 commonsourceibias.t33 gnd 0.017311f
C5972 commonsourceibias.t63 gnd 0.017311f
C5973 commonsourceibias.n386 gnd 0.152968f
C5974 commonsourceibias.n387 gnd 0.058702f
C5975 commonsourceibias.n388 gnd 0.010705f
C5976 commonsourceibias.t30 gnd 0.149881f
C5977 commonsourceibias.n389 gnd 0.007808f
C5978 commonsourceibias.n390 gnd 0.008022f
C5979 commonsourceibias.t44 gnd 0.149881f
C5980 commonsourceibias.n391 gnd 0.010321f
C5981 commonsourceibias.n392 gnd 0.008022f
C5982 commonsourceibias.t18 gnd 0.149881f
C5983 commonsourceibias.n393 gnd 0.007564f
C5984 commonsourceibias.n394 gnd 0.008022f
C5985 commonsourceibias.t58 gnd 0.149881f
C5986 commonsourceibias.n395 gnd 0.010168f
C5987 commonsourceibias.n396 gnd 0.008022f
C5988 commonsourceibias.t8 gnd 0.149881f
C5989 commonsourceibias.n397 gnd 0.007348f
C5990 commonsourceibias.n398 gnd 0.008022f
C5991 commonsourceibias.t56 gnd 0.149881f
C5992 commonsourceibias.n399 gnd 0.009997f
C5993 commonsourceibias.n400 gnd 0.008022f
C5994 commonsourceibias.t62 gnd 0.149881f
C5995 commonsourceibias.n401 gnd 0.007159f
C5996 commonsourceibias.n402 gnd 0.008022f
C5997 commonsourceibias.t32 gnd 0.149881f
C5998 commonsourceibias.n403 gnd 0.009806f
C5999 commonsourceibias.n404 gnd 0.008022f
C6000 commonsourceibias.t60 gnd 0.149881f
C6001 commonsourceibias.n405 gnd 0.006995f
C6002 commonsourceibias.n406 gnd 0.008022f
C6003 commonsourceibias.t64 gnd 0.149881f
C6004 commonsourceibias.n407 gnd 0.009595f
C6005 commonsourceibias.n408 gnd 0.008022f
C6006 commonsourceibias.t34 gnd 0.149881f
C6007 commonsourceibias.n409 gnd 0.006855f
C6008 commonsourceibias.n410 gnd 0.008022f
C6009 commonsourceibias.t6 gnd 0.149881f
C6010 commonsourceibias.n411 gnd 0.00936f
C6011 commonsourceibias.t36 gnd 0.16664f
C6012 commonsourceibias.t14 gnd 0.149881f
C6013 commonsourceibias.n412 gnd 0.065328f
C6014 commonsourceibias.n413 gnd 0.07169f
C6015 commonsourceibias.n414 gnd 0.033265f
C6016 commonsourceibias.n415 gnd 0.008022f
C6017 commonsourceibias.n416 gnd 0.007808f
C6018 commonsourceibias.n417 gnd 0.01119f
C6019 commonsourceibias.n418 gnd 0.059802f
C6020 commonsourceibias.n419 gnd 0.011182f
C6021 commonsourceibias.n420 gnd 0.008022f
C6022 commonsourceibias.n421 gnd 0.008022f
C6023 commonsourceibias.n422 gnd 0.008022f
C6024 commonsourceibias.n423 gnd 0.010321f
C6025 commonsourceibias.n424 gnd 0.059802f
C6026 commonsourceibias.n425 gnd 0.010563f
C6027 commonsourceibias.t48 gnd 0.149881f
C6028 commonsourceibias.n426 gnd 0.059802f
C6029 commonsourceibias.n427 gnd 0.010263f
C6030 commonsourceibias.n428 gnd 0.008022f
C6031 commonsourceibias.n429 gnd 0.008022f
C6032 commonsourceibias.n430 gnd 0.008022f
C6033 commonsourceibias.n431 gnd 0.007564f
C6034 commonsourceibias.n432 gnd 0.0112f
C6035 commonsourceibias.n433 gnd 0.059802f
C6036 commonsourceibias.n434 gnd 0.011196f
C6037 commonsourceibias.n435 gnd 0.008022f
C6038 commonsourceibias.n436 gnd 0.008022f
C6039 commonsourceibias.n437 gnd 0.008022f
C6040 commonsourceibias.n438 gnd 0.010168f
C6041 commonsourceibias.n439 gnd 0.059802f
C6042 commonsourceibias.n440 gnd 0.010488f
C6043 commonsourceibias.t2 gnd 0.149881f
C6044 commonsourceibias.n441 gnd 0.059802f
C6045 commonsourceibias.n442 gnd 0.010338f
C6046 commonsourceibias.n443 gnd 0.008022f
C6047 commonsourceibias.n444 gnd 0.008022f
C6048 commonsourceibias.n445 gnd 0.008022f
C6049 commonsourceibias.n446 gnd 0.007348f
C6050 commonsourceibias.n447 gnd 0.011204f
C6051 commonsourceibias.n448 gnd 0.059802f
C6052 commonsourceibias.n449 gnd 0.011203f
C6053 commonsourceibias.n450 gnd 0.008022f
C6054 commonsourceibias.n451 gnd 0.008022f
C6055 commonsourceibias.n452 gnd 0.008022f
C6056 commonsourceibias.n453 gnd 0.009997f
C6057 commonsourceibias.n454 gnd 0.059802f
C6058 commonsourceibias.n455 gnd 0.010413f
C6059 commonsourceibias.t26 gnd 0.149881f
C6060 commonsourceibias.n456 gnd 0.059802f
C6061 commonsourceibias.n457 gnd 0.010413f
C6062 commonsourceibias.n458 gnd 0.008022f
C6063 commonsourceibias.n459 gnd 0.008022f
C6064 commonsourceibias.n460 gnd 0.008022f
C6065 commonsourceibias.n461 gnd 0.007159f
C6066 commonsourceibias.n462 gnd 0.011203f
C6067 commonsourceibias.n463 gnd 0.059802f
C6068 commonsourceibias.n464 gnd 0.011204f
C6069 commonsourceibias.n465 gnd 0.008022f
C6070 commonsourceibias.n466 gnd 0.008022f
C6071 commonsourceibias.n467 gnd 0.008022f
C6072 commonsourceibias.n468 gnd 0.009806f
C6073 commonsourceibias.n469 gnd 0.059802f
C6074 commonsourceibias.n470 gnd 0.010338f
C6075 commonsourceibias.t70 gnd 0.149881f
C6076 commonsourceibias.n471 gnd 0.059802f
C6077 commonsourceibias.n472 gnd 0.010488f
C6078 commonsourceibias.n473 gnd 0.008022f
C6079 commonsourceibias.n474 gnd 0.008022f
C6080 commonsourceibias.n475 gnd 0.008022f
C6081 commonsourceibias.n476 gnd 0.006995f
C6082 commonsourceibias.n477 gnd 0.011196f
C6083 commonsourceibias.n478 gnd 0.059802f
C6084 commonsourceibias.n479 gnd 0.0112f
C6085 commonsourceibias.n480 gnd 0.008022f
C6086 commonsourceibias.n481 gnd 0.008022f
C6087 commonsourceibias.n482 gnd 0.008022f
C6088 commonsourceibias.n483 gnd 0.009595f
C6089 commonsourceibias.n484 gnd 0.059802f
C6090 commonsourceibias.n485 gnd 0.010263f
C6091 commonsourceibias.t78 gnd 0.149881f
C6092 commonsourceibias.n486 gnd 0.059802f
C6093 commonsourceibias.n487 gnd 0.010563f
C6094 commonsourceibias.n488 gnd 0.008022f
C6095 commonsourceibias.n489 gnd 0.008022f
C6096 commonsourceibias.n490 gnd 0.008022f
C6097 commonsourceibias.n491 gnd 0.006855f
C6098 commonsourceibias.n492 gnd 0.011182f
C6099 commonsourceibias.n493 gnd 0.059802f
C6100 commonsourceibias.n494 gnd 0.01119f
C6101 commonsourceibias.n495 gnd 0.008022f
C6102 commonsourceibias.n496 gnd 0.008022f
C6103 commonsourceibias.n497 gnd 0.008022f
C6104 commonsourceibias.n498 gnd 0.00936f
C6105 commonsourceibias.n499 gnd 0.059802f
C6106 commonsourceibias.n500 gnd 0.009843f
C6107 commonsourceibias.t52 gnd 0.162096f
C6108 commonsourceibias.n501 gnd 0.071758f
C6109 commonsourceibias.n502 gnd 0.079928f
C6110 commonsourceibias.t31 gnd 0.017311f
C6111 commonsourceibias.t53 gnd 0.017311f
C6112 commonsourceibias.n503 gnd 0.152968f
C6113 commonsourceibias.n504 gnd 0.132319f
C6114 commonsourceibias.t79 gnd 0.017311f
C6115 commonsourceibias.t45 gnd 0.017311f
C6116 commonsourceibias.n505 gnd 0.152968f
C6117 commonsourceibias.n506 gnd 0.070264f
C6118 commonsourceibias.t59 gnd 0.017311f
C6119 commonsourceibias.t19 gnd 0.017311f
C6120 commonsourceibias.n507 gnd 0.152968f
C6121 commonsourceibias.n508 gnd 0.070264f
C6122 commonsourceibias.t9 gnd 0.017311f
C6123 commonsourceibias.t71 gnd 0.017311f
C6124 commonsourceibias.n509 gnd 0.152968f
C6125 commonsourceibias.n510 gnd 0.070264f
C6126 commonsourceibias.t27 gnd 0.017311f
C6127 commonsourceibias.t57 gnd 0.017311f
C6128 commonsourceibias.n511 gnd 0.152968f
C6129 commonsourceibias.n512 gnd 0.058702f
C6130 commonsourceibias.n513 gnd 0.071082f
C6131 commonsourceibias.n514 gnd 0.05192f
C6132 commonsourceibias.t98 gnd 0.149881f
C6133 commonsourceibias.n515 gnd 0.059802f
C6134 commonsourceibias.n516 gnd 0.008022f
C6135 commonsourceibias.t125 gnd 0.149881f
C6136 commonsourceibias.n517 gnd 0.059802f
C6137 commonsourceibias.n518 gnd 0.008022f
C6138 commonsourceibias.t142 gnd 0.149881f
C6139 commonsourceibias.n519 gnd 0.059802f
C6140 commonsourceibias.n520 gnd 0.008022f
C6141 commonsourceibias.t155 gnd 0.149881f
C6142 commonsourceibias.n521 gnd 0.006995f
C6143 commonsourceibias.n522 gnd 0.008022f
C6144 commonsourceibias.t114 gnd 0.149881f
C6145 commonsourceibias.n523 gnd 0.009595f
C6146 commonsourceibias.n524 gnd 0.008022f
C6147 commonsourceibias.t148 gnd 0.149881f
C6148 commonsourceibias.n525 gnd 0.006855f
C6149 commonsourceibias.n526 gnd 0.008022f
C6150 commonsourceibias.t82 gnd 0.149881f
C6151 commonsourceibias.n527 gnd 0.00936f
C6152 commonsourceibias.t126 gnd 0.16664f
C6153 commonsourceibias.t89 gnd 0.149881f
C6154 commonsourceibias.n528 gnd 0.065328f
C6155 commonsourceibias.n529 gnd 0.07169f
C6156 commonsourceibias.n530 gnd 0.033265f
C6157 commonsourceibias.n531 gnd 0.008022f
C6158 commonsourceibias.n532 gnd 0.007808f
C6159 commonsourceibias.n533 gnd 0.01119f
C6160 commonsourceibias.n534 gnd 0.059802f
C6161 commonsourceibias.n535 gnd 0.011182f
C6162 commonsourceibias.n536 gnd 0.008022f
C6163 commonsourceibias.n537 gnd 0.008022f
C6164 commonsourceibias.n538 gnd 0.008022f
C6165 commonsourceibias.n539 gnd 0.010321f
C6166 commonsourceibias.n540 gnd 0.059802f
C6167 commonsourceibias.n541 gnd 0.010563f
C6168 commonsourceibias.t134 gnd 0.149881f
C6169 commonsourceibias.n542 gnd 0.059802f
C6170 commonsourceibias.n543 gnd 0.010263f
C6171 commonsourceibias.n544 gnd 0.008022f
C6172 commonsourceibias.n545 gnd 0.008022f
C6173 commonsourceibias.n546 gnd 0.008022f
C6174 commonsourceibias.n547 gnd 0.007564f
C6175 commonsourceibias.n548 gnd 0.0112f
C6176 commonsourceibias.n549 gnd 0.059802f
C6177 commonsourceibias.n550 gnd 0.011196f
C6178 commonsourceibias.n551 gnd 0.008022f
C6179 commonsourceibias.n552 gnd 0.008022f
C6180 commonsourceibias.n553 gnd 0.008022f
C6181 commonsourceibias.n554 gnd 0.010168f
C6182 commonsourceibias.n555 gnd 0.059802f
C6183 commonsourceibias.n556 gnd 0.010488f
C6184 commonsourceibias.n557 gnd 0.010338f
C6185 commonsourceibias.n558 gnd 0.008022f
C6186 commonsourceibias.n559 gnd 0.008022f
C6187 commonsourceibias.n560 gnd 0.009806f
C6188 commonsourceibias.n561 gnd 0.007348f
C6189 commonsourceibias.n562 gnd 0.011204f
C6190 commonsourceibias.n563 gnd 0.008022f
C6191 commonsourceibias.n564 gnd 0.008022f
C6192 commonsourceibias.n565 gnd 0.011203f
C6193 commonsourceibias.n566 gnd 0.007159f
C6194 commonsourceibias.n567 gnd 0.009997f
C6195 commonsourceibias.n568 gnd 0.008022f
C6196 commonsourceibias.n569 gnd 0.007008f
C6197 commonsourceibias.n570 gnd 0.010413f
C6198 commonsourceibias.t149 gnd 0.149881f
C6199 commonsourceibias.n571 gnd 0.059802f
C6200 commonsourceibias.n572 gnd 0.010413f
C6201 commonsourceibias.n573 gnd 0.007008f
C6202 commonsourceibias.n574 gnd 0.008022f
C6203 commonsourceibias.n575 gnd 0.008022f
C6204 commonsourceibias.n576 gnd 0.007159f
C6205 commonsourceibias.n577 gnd 0.011203f
C6206 commonsourceibias.n578 gnd 0.059802f
C6207 commonsourceibias.n579 gnd 0.011204f
C6208 commonsourceibias.n580 gnd 0.008022f
C6209 commonsourceibias.n581 gnd 0.008022f
C6210 commonsourceibias.n582 gnd 0.008022f
C6211 commonsourceibias.n583 gnd 0.009806f
C6212 commonsourceibias.n584 gnd 0.059802f
C6213 commonsourceibias.n585 gnd 0.010338f
C6214 commonsourceibias.t156 gnd 0.149881f
C6215 commonsourceibias.n586 gnd 0.059802f
C6216 commonsourceibias.n587 gnd 0.010488f
C6217 commonsourceibias.n588 gnd 0.008022f
C6218 commonsourceibias.n589 gnd 0.008022f
C6219 commonsourceibias.n590 gnd 0.008022f
C6220 commonsourceibias.n591 gnd 0.006995f
C6221 commonsourceibias.n592 gnd 0.011196f
C6222 commonsourceibias.n593 gnd 0.059802f
C6223 commonsourceibias.n594 gnd 0.0112f
C6224 commonsourceibias.n595 gnd 0.008022f
C6225 commonsourceibias.n596 gnd 0.008022f
C6226 commonsourceibias.n597 gnd 0.008022f
C6227 commonsourceibias.n598 gnd 0.009595f
C6228 commonsourceibias.n599 gnd 0.059802f
C6229 commonsourceibias.n600 gnd 0.010263f
C6230 commonsourceibias.t105 gnd 0.149881f
C6231 commonsourceibias.n601 gnd 0.059802f
C6232 commonsourceibias.n602 gnd 0.010563f
C6233 commonsourceibias.n603 gnd 0.008022f
C6234 commonsourceibias.n604 gnd 0.008022f
C6235 commonsourceibias.n605 gnd 0.008022f
C6236 commonsourceibias.n606 gnd 0.006855f
C6237 commonsourceibias.n607 gnd 0.011182f
C6238 commonsourceibias.n608 gnd 0.059802f
C6239 commonsourceibias.n609 gnd 0.01119f
C6240 commonsourceibias.n610 gnd 0.008022f
C6241 commonsourceibias.n611 gnd 0.008022f
C6242 commonsourceibias.n612 gnd 0.008022f
C6243 commonsourceibias.n613 gnd 0.00936f
C6244 commonsourceibias.n614 gnd 0.059802f
C6245 commonsourceibias.n615 gnd 0.009843f
C6246 commonsourceibias.n616 gnd 0.071758f
C6247 commonsourceibias.n617 gnd 0.046883f
C6248 commonsourceibias.n618 gnd 0.010705f
C6249 commonsourceibias.t141 gnd 0.149881f
C6250 commonsourceibias.n619 gnd 0.007808f
C6251 commonsourceibias.n620 gnd 0.008022f
C6252 commonsourceibias.t154 gnd 0.149881f
C6253 commonsourceibias.n621 gnd 0.010321f
C6254 commonsourceibias.n622 gnd 0.008022f
C6255 commonsourceibias.t132 gnd 0.149881f
C6256 commonsourceibias.n623 gnd 0.007564f
C6257 commonsourceibias.n624 gnd 0.008022f
C6258 commonsourceibias.t147 gnd 0.149881f
C6259 commonsourceibias.n625 gnd 0.010168f
C6260 commonsourceibias.n626 gnd 0.008022f
C6261 commonsourceibias.t123 gnd 0.149881f
C6262 commonsourceibias.n627 gnd 0.007348f
C6263 commonsourceibias.n628 gnd 0.008022f
C6264 commonsourceibias.t115 gnd 0.149881f
C6265 commonsourceibias.n629 gnd 0.009997f
C6266 commonsourceibias.n630 gnd 0.008022f
C6267 commonsourceibias.t88 gnd 0.149881f
C6268 commonsourceibias.n631 gnd 0.007159f
C6269 commonsourceibias.n632 gnd 0.008022f
C6270 commonsourceibias.t106 gnd 0.149881f
C6271 commonsourceibias.n633 gnd 0.009806f
C6272 commonsourceibias.n634 gnd 0.008022f
C6273 commonsourceibias.t143 gnd 0.149881f
C6274 commonsourceibias.n635 gnd 0.006995f
C6275 commonsourceibias.n636 gnd 0.008022f
C6276 commonsourceibias.t99 gnd 0.149881f
C6277 commonsourceibias.n637 gnd 0.009595f
C6278 commonsourceibias.n638 gnd 0.008022f
C6279 commonsourceibias.t136 gnd 0.149881f
C6280 commonsourceibias.n639 gnd 0.006855f
C6281 commonsourceibias.n640 gnd 0.008022f
C6282 commonsourceibias.t150 gnd 0.149881f
C6283 commonsourceibias.n641 gnd 0.00936f
C6284 commonsourceibias.t108 gnd 0.16664f
C6285 commonsourceibias.t158 gnd 0.149881f
C6286 commonsourceibias.n642 gnd 0.065328f
C6287 commonsourceibias.n643 gnd 0.07169f
C6288 commonsourceibias.n644 gnd 0.033265f
C6289 commonsourceibias.n645 gnd 0.008022f
C6290 commonsourceibias.n646 gnd 0.007808f
C6291 commonsourceibias.n647 gnd 0.01119f
C6292 commonsourceibias.n648 gnd 0.059802f
C6293 commonsourceibias.n649 gnd 0.011182f
C6294 commonsourceibias.n650 gnd 0.008022f
C6295 commonsourceibias.n651 gnd 0.008022f
C6296 commonsourceibias.n652 gnd 0.008022f
C6297 commonsourceibias.n653 gnd 0.010321f
C6298 commonsourceibias.n654 gnd 0.059802f
C6299 commonsourceibias.n655 gnd 0.010563f
C6300 commonsourceibias.t118 gnd 0.149881f
C6301 commonsourceibias.n656 gnd 0.059802f
C6302 commonsourceibias.n657 gnd 0.010263f
C6303 commonsourceibias.n658 gnd 0.008022f
C6304 commonsourceibias.n659 gnd 0.008022f
C6305 commonsourceibias.n660 gnd 0.008022f
C6306 commonsourceibias.n661 gnd 0.007564f
C6307 commonsourceibias.n662 gnd 0.0112f
C6308 commonsourceibias.n663 gnd 0.059802f
C6309 commonsourceibias.n664 gnd 0.011196f
C6310 commonsourceibias.n665 gnd 0.008022f
C6311 commonsourceibias.n666 gnd 0.008022f
C6312 commonsourceibias.n667 gnd 0.008022f
C6313 commonsourceibias.n668 gnd 0.010168f
C6314 commonsourceibias.n669 gnd 0.059802f
C6315 commonsourceibias.n670 gnd 0.010488f
C6316 commonsourceibias.t128 gnd 0.149881f
C6317 commonsourceibias.n671 gnd 0.059802f
C6318 commonsourceibias.n672 gnd 0.010338f
C6319 commonsourceibias.n673 gnd 0.008022f
C6320 commonsourceibias.n674 gnd 0.008022f
C6321 commonsourceibias.n675 gnd 0.008022f
C6322 commonsourceibias.n676 gnd 0.007348f
C6323 commonsourceibias.n677 gnd 0.011204f
C6324 commonsourceibias.n678 gnd 0.059802f
C6325 commonsourceibias.n679 gnd 0.011203f
C6326 commonsourceibias.n680 gnd 0.008022f
C6327 commonsourceibias.n681 gnd 0.008022f
C6328 commonsourceibias.n682 gnd 0.008022f
C6329 commonsourceibias.n683 gnd 0.009997f
C6330 commonsourceibias.n684 gnd 0.059802f
C6331 commonsourceibias.n685 gnd 0.010413f
C6332 commonsourceibias.t137 gnd 0.149881f
C6333 commonsourceibias.n686 gnd 0.059802f
C6334 commonsourceibias.n687 gnd 0.010413f
C6335 commonsourceibias.n688 gnd 0.008022f
C6336 commonsourceibias.n689 gnd 0.008022f
C6337 commonsourceibias.n690 gnd 0.008022f
C6338 commonsourceibias.n691 gnd 0.007159f
C6339 commonsourceibias.n692 gnd 0.011203f
C6340 commonsourceibias.n693 gnd 0.059802f
C6341 commonsourceibias.n694 gnd 0.011204f
C6342 commonsourceibias.n695 gnd 0.008022f
C6343 commonsourceibias.n696 gnd 0.008022f
C6344 commonsourceibias.n697 gnd 0.008022f
C6345 commonsourceibias.n698 gnd 0.009806f
C6346 commonsourceibias.n699 gnd 0.059802f
C6347 commonsourceibias.n700 gnd 0.010338f
C6348 commonsourceibias.t144 gnd 0.149881f
C6349 commonsourceibias.n701 gnd 0.059802f
C6350 commonsourceibias.n702 gnd 0.010488f
C6351 commonsourceibias.n703 gnd 0.008022f
C6352 commonsourceibias.n704 gnd 0.008022f
C6353 commonsourceibias.n705 gnd 0.008022f
C6354 commonsourceibias.n706 gnd 0.006995f
C6355 commonsourceibias.n707 gnd 0.011196f
C6356 commonsourceibias.n708 gnd 0.059802f
C6357 commonsourceibias.n709 gnd 0.0112f
C6358 commonsourceibias.n710 gnd 0.008022f
C6359 commonsourceibias.n711 gnd 0.008022f
C6360 commonsourceibias.n712 gnd 0.008022f
C6361 commonsourceibias.n713 gnd 0.009595f
C6362 commonsourceibias.n714 gnd 0.059802f
C6363 commonsourceibias.n715 gnd 0.010263f
C6364 commonsourceibias.t93 gnd 0.149881f
C6365 commonsourceibias.n716 gnd 0.059802f
C6366 commonsourceibias.n717 gnd 0.010563f
C6367 commonsourceibias.n718 gnd 0.008022f
C6368 commonsourceibias.n719 gnd 0.008022f
C6369 commonsourceibias.n720 gnd 0.008022f
C6370 commonsourceibias.n721 gnd 0.006855f
C6371 commonsourceibias.n722 gnd 0.011182f
C6372 commonsourceibias.n723 gnd 0.059802f
C6373 commonsourceibias.n724 gnd 0.01119f
C6374 commonsourceibias.n725 gnd 0.008022f
C6375 commonsourceibias.n726 gnd 0.008022f
C6376 commonsourceibias.n727 gnd 0.008022f
C6377 commonsourceibias.n728 gnd 0.00936f
C6378 commonsourceibias.n729 gnd 0.059802f
C6379 commonsourceibias.n730 gnd 0.009843f
C6380 commonsourceibias.t124 gnd 0.162096f
C6381 commonsourceibias.n731 gnd 0.071758f
C6382 commonsourceibias.n732 gnd 0.024957f
C6383 commonsourceibias.n733 gnd 0.221543f
C6384 commonsourceibias.n734 gnd 4.49224f
.ends

