* NGSPICE file created from opamp158.ext - technology: sky130A

.subckt opamp158 gnd CSoutput output vdd plus minus commonsourceibias outputibias
+ diffpairibias
X0 a_n2472_13878.t24 a_n2848_n452.t52 a_n2848_n452.t53 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 CSoutput.t71 a_n6972_8799.t44 vdd.t16 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X2 a_n2472_13878.t3 a_n2848_n452.t64 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X3 vdd.t130 a_n6972_8799.t45 CSoutput.t70 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X4 commonsourceibias.t39 commonsourceibias.t38 gnd.t351 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X5 gnd.t350 commonsourceibias.t80 CSoutput.t91 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X6 vdd.t103 vdd.t101 vdd.t102 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X7 gnd.t118 gnd.t116 gnd.t117 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X8 a_n6972_8799.t43 plus.t5 a_n3106_n452.t29 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X9 outputibias.t7 outputibias.t6 gnd.t160 gnd.t159 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X10 CSoutput.t69 a_n6972_8799.t46 vdd.t140 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X11 gnd.t338 commonsourceibias.t81 CSoutput.t15 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 a_n3106_n452.t28 plus.t6 a_n6972_8799.t41 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X13 CSoutput.t128 a_n2650_8322.t5 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X14 gnd.t349 commonsourceibias.t36 commonsourceibias.t37 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X15 gnd.t348 commonsourceibias.t82 CSoutput.t107 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X16 a_n2650_8322.t33 a_n2848_n452.t65 a_n6972_8799.t29 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 gnd.t347 commonsourceibias.t83 CSoutput.t109 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X18 gnd.t346 commonsourceibias.t84 CSoutput.t72 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X19 output.t19 CSoutput.t129 vdd.t113 gnd.t151 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X20 CSoutput.t68 a_n6972_8799.t47 vdd.t148 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X21 vdd.t118 a_n6972_8799.t48 CSoutput.t67 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X22 gnd.t345 commonsourceibias.t85 CSoutput.t94 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X23 outputibias.t5 outputibias.t4 gnd.t158 gnd.t157 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X24 a_n6972_8799.t27 a_n2848_n452.t66 a_n2650_8322.t32 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X25 a_n2848_n452.t11 minus.t5 a_n3106_n452.t41 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X26 a_n6972_8799.t39 plus.t7 a_n3106_n452.t27 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X27 gnd.t344 commonsourceibias.t78 commonsourceibias.t79 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 plus.t4 gnd.t113 gnd.t115 gnd.t114 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X29 a_n2848_n452.t10 minus.t6 a_n3106_n452.t40 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X30 a_n6972_8799.t36 a_n2848_n452.t67 a_n2650_8322.t31 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X31 CSoutput.t0 commonsourceibias.t86 gnd.t343 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 gnd.t342 commonsourceibias.t76 commonsourceibias.t77 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X33 CSoutput.t66 a_n6972_8799.t49 vdd.t112 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X34 CSoutput.t4 commonsourceibias.t87 gnd.t341 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X35 a_n3106_n452.t26 plus.t8 a_n6972_8799.t7 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X36 vdd.t114 CSoutput.t130 output.t18 gnd.t150 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X37 vdd.t100 vdd.t98 vdd.t99 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X38 a_n3106_n452.t43 minus.t7 a_n2848_n452.t13 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X39 CSoutput.t95 commonsourceibias.t88 gnd.t337 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X40 a_n3106_n452.t35 diffpairibias.t16 gnd.t162 gnd.t161 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X41 CSoutput.t105 commonsourceibias.t89 gnd.t340 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X42 CSoutput.t65 a_n6972_8799.t50 vdd.t141 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X43 CSoutput.t84 commonsourceibias.t90 gnd.t339 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X44 vdd.t97 vdd.t95 vdd.t96 vdd.t45 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X45 output.t17 CSoutput.t131 vdd.t115 gnd.t149 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X46 outputibias.t3 outputibias.t2 gnd.t10 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X47 gnd.t336 commonsourceibias.t34 commonsourceibias.t35 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X48 a_n2472_13878.t23 a_n2848_n452.t58 a_n2848_n452.t59 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X49 a_n2848_n452.t37 a_n2848_n452.t36 a_n2472_13878.t22 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X50 CSoutput.t92 commonsourceibias.t91 gnd.t335 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 commonsourceibias.t33 commonsourceibias.t32 gnd.t334 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X52 CSoutput.t64 a_n6972_8799.t51 vdd.t11 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X53 gnd.t112 gnd.t110 gnd.t111 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X54 CSoutput.t132 a_n2650_8322.t4 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X55 vdd.t94 vdd.t92 vdd.t93 vdd.t75 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X56 vdd.t206 a_n6972_8799.t52 CSoutput.t63 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X57 a_n3106_n452.t25 plus.t9 a_n6972_8799.t4 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X58 a_n3106_n452.t24 plus.t10 a_n6972_8799.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X59 a_n3106_n452.t39 minus.t8 a_n2848_n452.t9 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X60 diffpairibias.t15 diffpairibias.t14 gnd.t153 gnd.t152 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X61 a_n2848_n452.t27 a_n2848_n452.t26 a_n2472_13878.t21 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X62 a_n6972_8799.t22 a_n2848_n452.t68 a_n2650_8322.t30 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X63 vdd.t125 a_n6972_8799.t53 CSoutput.t62 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X64 a_n2848_n452.t29 a_n2848_n452.t28 a_n2472_13878.t20 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X65 CSoutput.t61 a_n6972_8799.t54 vdd.t131 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X66 gnd.t109 gnd.t107 gnd.t108 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X67 a_n6972_8799.t21 a_n2848_n452.t69 a_n2650_8322.t29 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X68 gnd.t333 commonsourceibias.t92 CSoutput.t16 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X69 gnd.t332 commonsourceibias.t93 CSoutput.t5 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X70 diffpairibias.t13 diffpairibias.t12 gnd.t355 gnd.t354 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X71 CSoutput.t60 a_n6972_8799.t55 vdd.t9 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X72 output.t16 CSoutput.t133 vdd.t26 gnd.t148 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X73 gnd.t324 commonsourceibias.t94 CSoutput.t108 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X74 commonsourceibias.t31 commonsourceibias.t30 gnd.t331 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X75 a_n2650_8322.t28 a_n2848_n452.t70 a_n6972_8799.t25 vdd.t198 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X76 gnd.t323 commonsourceibias.t95 CSoutput.t110 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X77 a_n3106_n452.t42 minus.t9 a_n2848_n452.t12 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X78 commonsourceibias.t29 commonsourceibias.t28 gnd.t330 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X79 a_n3106_n452.t23 plus.t11 a_n6972_8799.t11 gnd.t173 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X80 output.t15 CSoutput.t134 vdd.t27 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X81 gnd.t329 commonsourceibias.t96 CSoutput.t77 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X82 a_n6972_8799.t42 plus.t12 a_n3106_n452.t22 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X83 commonsourceibias.t17 commonsourceibias.t16 gnd.t328 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X84 CSoutput.t73 commonsourceibias.t97 gnd.t327 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 CSoutput.t135 a_n2650_8322.t3 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X86 a_n3106_n452.t53 diffpairibias.t17 gnd.t191 gnd.t190 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X87 gnd.t326 commonsourceibias.t14 commonsourceibias.t15 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X88 vdd.t108 a_n6972_8799.t56 CSoutput.t59 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X89 a_n6972_8799.t20 a_n2848_n452.t71 a_n2650_8322.t27 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X90 a_n2848_n452.t55 a_n2848_n452.t54 a_n2472_13878.t19 vdd.t197 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X91 a_n3106_n452.t21 plus.t13 a_n6972_8799.t38 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X92 a_n2848_n452.t25 a_n2848_n452.t24 a_n2472_13878.t18 vdd.t153 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X93 gnd.t325 commonsourceibias.t12 commonsourceibias.t13 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X94 commonsourceibias.t11 commonsourceibias.t10 gnd.t322 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X95 CSoutput.t58 a_n6972_8799.t57 vdd.t17 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X96 vdd.t202 a_n6972_8799.t58 CSoutput.t57 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X97 CSoutput.t119 commonsourceibias.t98 gnd.t321 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 a_n2848_n452.t15 minus.t10 a_n3106_n452.t46 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X99 CSoutput.t112 commonsourceibias.t99 gnd.t320 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 vdd.t132 CSoutput.t136 output.t14 gnd.t146 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X101 CSoutput.t56 a_n6972_8799.t59 vdd.t146 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X102 vdd.t91 vdd.t89 vdd.t90 vdd.t79 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X103 CSoutput.t81 commonsourceibias.t100 gnd.t319 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X104 vdd.t88 vdd.t85 vdd.t87 vdd.t86 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X105 CSoutput.t6 commonsourceibias.t101 gnd.t318 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X106 gnd.t317 commonsourceibias.t102 CSoutput.t96 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X107 commonsourceibias.t25 commonsourceibias.t24 gnd.t316 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 CSoutput.t85 commonsourceibias.t103 gnd.t315 gnd.t314 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 vdd.t84 vdd.t82 vdd.t83 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X110 a_n2650_8322.t13 a_n2848_n452.t72 vdd.t192 vdd.t191 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X111 vdd.t194 a_n2848_n452.t73 a_n2650_8322.t12 vdd.t193 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X112 a_n2848_n452.t41 a_n2848_n452.t40 a_n2472_13878.t17 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X113 gnd.t313 commonsourceibias.t104 CSoutput.t78 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X114 a_n3106_n452.t2 diffpairibias.t18 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X115 gnd.t106 gnd.t104 minus.t4 gnd.t105 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X116 gnd.t103 gnd.t101 gnd.t102 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X117 commonsourceibias.t23 commonsourceibias.t22 gnd.t312 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X118 vdd.t196 a_n2848_n452.t74 a_n2472_13878.t0 vdd.t195 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X119 commonsourceibias.t21 commonsourceibias.t20 gnd.t311 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X120 vdd.t81 vdd.t78 vdd.t80 vdd.t79 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X121 gnd.t310 commonsourceibias.t44 commonsourceibias.t45 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X122 gnd.t309 commonsourceibias.t42 commonsourceibias.t43 gnd.t308 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X123 gnd.t307 commonsourceibias.t105 CSoutput.t74 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 gnd.t100 gnd.t98 plus.t3 gnd.t99 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X125 outputibias.t1 outputibias.t0 gnd.t353 gnd.t352 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X126 a_n6972_8799.t34 a_n2848_n452.t75 a_n2650_8322.t26 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X127 a_n2650_8322.t11 a_n2848_n452.t76 vdd.t190 vdd.t189 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X128 vdd.t77 vdd.t74 vdd.t76 vdd.t75 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X129 gnd.t306 commonsourceibias.t106 CSoutput.t120 gnd.t305 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 a_n2848_n452.t21 minus.t11 a_n3106_n452.t52 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X131 a_n6972_8799.t14 plus.t14 a_n3106_n452.t20 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X132 gnd.t304 commonsourceibias.t107 CSoutput.t113 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X133 commonsourceibias.t41 commonsourceibias.t40 gnd.t303 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X134 vdd.t7 a_n6972_8799.t60 CSoutput.t55 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X135 a_n2848_n452.t61 a_n2848_n452.t60 a_n2472_13878.t16 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X136 a_n6972_8799.t5 plus.t15 a_n3106_n452.t19 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X137 a_n2848_n452.t20 minus.t12 a_n3106_n452.t51 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X138 gnd.t302 commonsourceibias.t108 CSoutput.t86 gnd.t262 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X139 diffpairibias.t11 diffpairibias.t10 gnd.t168 gnd.t167 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X140 CSoutput.t54 a_n6972_8799.t61 vdd.t1 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X141 a_n6972_8799.t30 a_n2848_n452.t77 a_n2650_8322.t25 vdd.t188 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X142 gnd.t301 commonsourceibias.t109 CSoutput.t124 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X143 a_n2472_13878.t15 a_n2848_n452.t56 a_n2848_n452.t57 vdd.t187 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X144 output.t3 outputibias.t8 gnd.t135 gnd.t134 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X145 CSoutput.t114 commonsourceibias.t110 gnd.t300 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 gnd.t299 commonsourceibias.t111 CSoutput.t97 gnd.t298 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X147 a_n3106_n452.t50 minus.t13 a_n2848_n452.t19 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X148 commonsourceibias.t19 commonsourceibias.t18 gnd.t297 gnd.t296 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X149 a_n2472_13878.t14 a_n2848_n452.t48 a_n2848_n452.t49 vdd.t186 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X150 CSoutput.t53 a_n6972_8799.t62 vdd.t127 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X151 vdd.t185 a_n2848_n452.t78 a_n2650_8322.t10 vdd.t184 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X152 gnd.t295 commonsourceibias.t112 CSoutput.t87 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X153 CSoutput.t125 commonsourceibias.t113 gnd.t294 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X154 a_n2848_n452.t51 a_n2848_n452.t50 a_n2472_13878.t13 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X155 vdd.t13 a_n6972_8799.t63 CSoutput.t52 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X156 vdd.t73 vdd.t71 vdd.t72 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X157 a_n3106_n452.t18 plus.t16 a_n6972_8799.t12 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X158 a_n2848_n452.t18 minus.t14 a_n3106_n452.t49 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X159 gnd.t97 gnd.t94 gnd.t96 gnd.t95 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X160 a_n3106_n452.t3 diffpairibias.t19 gnd.t6 gnd.t5 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X161 CSoutput.t115 commonsourceibias.t114 gnd.t293 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X162 CSoutput.t98 commonsourceibias.t115 gnd.t292 gnd.t291 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X163 a_n6972_8799.t1 plus.t17 a_n3106_n452.t17 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X164 CSoutput.t1 commonsourceibias.t116 gnd.t290 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 vdd.t133 CSoutput.t137 output.t13 gnd.t145 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X166 a_n3106_n452.t30 diffpairibias.t20 gnd.t122 gnd.t121 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X167 CSoutput.t7 commonsourceibias.t117 gnd.t289 gnd.t288 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X168 gnd.t287 commonsourceibias.t118 CSoutput.t99 gnd.t286 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X169 gnd.t285 commonsourceibias.t119 CSoutput.t106 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 CSoutput.t88 commonsourceibias.t120 gnd.t284 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X171 commonsourceibias.t27 commonsourceibias.t26 gnd.t283 gnd.t282 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X172 a_n2472_13878.t12 a_n2848_n452.t30 a_n2848_n452.t31 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X173 a_n6972_8799.t2 plus.t18 a_n3106_n452.t16 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X174 gnd.t93 gnd.t91 gnd.t92 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X175 vdd.t70 vdd.t68 vdd.t69 vdd.t41 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X176 a_n2650_8322.t24 a_n2848_n452.t79 a_n6972_8799.t31 vdd.t183 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X177 gnd.t281 commonsourceibias.t121 CSoutput.t93 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X178 gnd.t90 gnd.t87 gnd.t89 gnd.t88 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X179 CSoutput.t51 a_n6972_8799.t64 vdd.t203 vdd.t15 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X180 minus.t3 gnd.t84 gnd.t86 gnd.t85 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X181 a_n2472_13878.t26 a_n2848_n452.t80 vdd.t182 vdd.t181 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 CSoutput.t17 commonsourceibias.t122 gnd.t280 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 gnd.t83 gnd.t81 gnd.t82 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X184 diffpairibias.t9 diffpairibias.t8 gnd.t178 gnd.t177 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X185 vdd.t180 a_n2848_n452.t81 a_n2472_13878.t25 vdd.t179 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X186 a_n2848_n452.t17 minus.t15 a_n3106_n452.t48 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X187 vdd.t147 a_n6972_8799.t65 CSoutput.t50 vdd.t12 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X188 CSoutput.t49 a_n6972_8799.t66 vdd.t205 vdd.t126 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 a_n3106_n452.t15 plus.t19 a_n6972_8799.t16 gnd.t182 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X190 CSoutput.t8 commonsourceibias.t123 gnd.t279 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X191 gnd.t278 commonsourceibias.t124 CSoutput.t111 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X192 a_n2472_13878.t11 a_n2848_n452.t46 a_n2848_n452.t47 vdd.t178 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X193 gnd.t277 commonsourceibias.t48 commonsourceibias.t49 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X194 gnd.t276 commonsourceibias.t125 CSoutput.t79 gnd.t262 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X195 gnd.t275 commonsourceibias.t126 CSoutput.t76 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X196 a_n2650_8322.t23 a_n2848_n452.t82 a_n6972_8799.t18 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X197 gnd.t274 commonsourceibias.t127 CSoutput.t75 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 a_n3106_n452.t47 minus.t16 a_n2848_n452.t16 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X199 a_n2472_13878.t10 a_n2848_n452.t22 a_n2848_n452.t23 vdd.t177 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X200 vdd.t135 a_n6972_8799.t67 CSoutput.t48 vdd.t117 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X201 CSoutput.t47 a_n6972_8799.t68 vdd.t123 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 CSoutput.t121 commonsourceibias.t128 gnd.t273 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X203 vdd.t104 CSoutput.t138 output.t12 gnd.t144 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X204 diffpairibias.t7 diffpairibias.t6 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X205 vdd.t173 a_n2848_n452.t83 a_n2650_8322.t9 vdd.t172 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X206 gnd.t272 commonsourceibias.t46 commonsourceibias.t47 gnd.t271 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X207 CSoutput.t116 commonsourceibias.t129 gnd.t270 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X208 a_n3106_n452.t33 minus.t17 a_n2848_n452.t6 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X209 a_n3106_n452.t14 plus.t20 a_n6972_8799.t3 gnd.t120 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X210 gnd.t80 gnd.t78 gnd.t79 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X211 gnd.t269 commonsourceibias.t130 CSoutput.t82 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X212 CSoutput.t18 commonsourceibias.t131 gnd.t261 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X213 a_n3106_n452.t36 minus.t18 a_n2848_n452.t8 gnd.t166 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X214 a_n2472_13878.t2 a_n2848_n452.t84 vdd.t176 vdd.t175 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X215 vdd.t3 a_n6972_8799.t69 CSoutput.t46 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X216 gnd.t268 commonsourceibias.t2 commonsourceibias.t3 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X217 gnd.t77 gnd.t74 gnd.t76 gnd.t75 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X218 a_n2650_8322.t22 a_n2848_n452.t85 a_n6972_8799.t17 vdd.t174 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X219 vdd.t171 a_n2848_n452.t86 a_n2650_8322.t8 vdd.t170 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X220 minus.t2 gnd.t71 gnd.t73 gnd.t72 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X221 CSoutput.t100 commonsourceibias.t132 gnd.t267 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X222 CSoutput.t139 a_n2650_8322.t2 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X223 a_n3106_n452.t38 diffpairibias.t21 gnd.t176 gnd.t175 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X224 CSoutput.t45 a_n6972_8799.t70 vdd.t128 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 vdd.t67 vdd.t65 vdd.t66 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X226 vdd.t64 vdd.t61 vdd.t63 vdd.t62 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X227 a_n6972_8799.t37 plus.t21 a_n3106_n452.t13 gnd.t181 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X228 a_n2848_n452.t7 minus.t19 a_n3106_n452.t34 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X229 CSoutput.t89 commonsourceibias.t133 gnd.t260 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X230 vdd.t116 a_n6972_8799.t71 CSoutput.t44 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X231 vdd.t22 a_n6972_8799.t72 CSoutput.t43 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X232 vdd.t60 vdd.t58 vdd.t59 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X233 a_n3106_n452.t44 minus.t20 a_n2848_n452.t14 gnd.t173 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X234 gnd.t266 commonsourceibias.t134 CSoutput.t126 gnd.t265 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 CSoutput.t117 commonsourceibias.t135 gnd.t264 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X236 vdd.t105 CSoutput.t140 output.t11 gnd.t143 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X237 gnd.t263 commonsourceibias.t0 commonsourceibias.t1 gnd.t262 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X238 gnd.t259 commonsourceibias.t8 commonsourceibias.t9 gnd.t258 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X239 gnd.t257 commonsourceibias.t136 CSoutput.t127 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X240 CSoutput.t101 commonsourceibias.t137 gnd.t249 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X241 output.t10 CSoutput.t141 vdd.t136 gnd.t142 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X242 vdd.t57 vdd.t54 vdd.t56 vdd.t55 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X243 a_n3106_n452.t31 minus.t21 a_n2848_n452.t4 gnd.t130 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X244 gnd.t70 gnd.t68 gnd.t69 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X245 CSoutput.t42 a_n6972_8799.t73 vdd.t138 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X246 a_n2472_13878.t9 a_n2848_n452.t32 a_n2848_n452.t33 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X247 a_n3106_n452.t0 minus.t22 a_n2848_n452.t0 gnd.t0 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X248 gnd.t67 gnd.t64 gnd.t66 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X249 vdd.t53 vdd.t51 vdd.t52 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X250 a_n2650_8322.t21 a_n2848_n452.t87 a_n6972_8799.t32 vdd.t169 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X251 gnd.t63 gnd.t61 gnd.t62 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X252 CSoutput.t103 commonsourceibias.t138 gnd.t256 gnd.t255 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X253 CSoutput.t142 a_n2650_8322.t1 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X254 diffpairibias.t5 diffpairibias.t4 gnd.t124 gnd.t123 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X255 CSoutput.t41 a_n6972_8799.t74 vdd.t134 vdd.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 commonsourceibias.t7 commonsourceibias.t6 gnd.t254 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X257 vdd.t25 a_n6972_8799.t75 CSoutput.t40 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X258 CSoutput.t102 commonsourceibias.t139 gnd.t253 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X259 gnd.t252 commonsourceibias.t140 CSoutput.t104 gnd.t251 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X260 vdd.t14 a_n6972_8799.t76 CSoutput.t39 vdd.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X261 a_n2650_8322.t7 a_n2848_n452.t88 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X262 gnd.t60 gnd.t57 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X263 gnd.t250 commonsourceibias.t141 CSoutput.t90 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 gnd.t248 commonsourceibias.t4 commonsourceibias.t5 gnd.t247 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X265 a_n3106_n452.t5 minus.t23 a_n2848_n452.t3 gnd.t8 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X266 vdd.t166 a_n2848_n452.t89 a_n2472_13878.t4 vdd.t165 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X267 gnd.t56 gnd.t54 gnd.t55 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X268 output.t2 outputibias.t9 gnd.t129 gnd.t128 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X269 CSoutput.t14 commonsourceibias.t142 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X270 CSoutput.t38 a_n6972_8799.t77 vdd.t19 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X271 vdd.t50 vdd.t48 vdd.t49 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X272 CSoutput.t37 a_n6972_8799.t78 vdd.t20 vdd.t10 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 output.t9 CSoutput.t143 vdd.t137 gnd.t141 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X274 vdd.t129 a_n6972_8799.t79 CSoutput.t36 vdd.t24 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 vdd.t120 a_n6972_8799.t80 CSoutput.t35 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 gnd.t53 gnd.t51 plus.t2 gnd.t52 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X277 CSoutput.t9 commonsourceibias.t143 gnd.t244 gnd.t243 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X278 gnd.t50 gnd.t47 gnd.t49 gnd.t48 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X279 CSoutput.t80 commonsourceibias.t144 gnd.t242 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X280 gnd.t241 commonsourceibias.t145 CSoutput.t122 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 vdd.t109 CSoutput.t144 output.t8 gnd.t140 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X282 gnd.t46 gnd.t43 gnd.t45 gnd.t44 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X283 output.t1 outputibias.t10 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X284 gnd.t240 commonsourceibias.t68 commonsourceibias.t69 gnd.t239 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X285 a_n6972_8799.t26 a_n2848_n452.t90 a_n2650_8322.t20 vdd.t164 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X286 a_n2650_8322.t19 a_n2848_n452.t91 a_n6972_8799.t23 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X287 a_n2472_13878.t1 a_n2848_n452.t92 vdd.t163 vdd.t162 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X288 vdd.t47 vdd.t44 vdd.t46 vdd.t45 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X289 vdd.t110 CSoutput.t145 output.t7 gnd.t139 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X290 output.t0 outputibias.t11 gnd.t132 gnd.t131 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X291 vdd.t207 a_n6972_8799.t81 CSoutput.t34 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X292 CSoutput.t33 a_n6972_8799.t82 vdd.t107 vdd.t106 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X293 vdd.t43 vdd.t40 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X294 vdd.t39 vdd.t36 vdd.t38 vdd.t37 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X295 a_n3106_n452.t12 plus.t22 a_n6972_8799.t8 gnd.t165 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X296 a_n2650_8322.t18 a_n2848_n452.t93 a_n6972_8799.t28 vdd.t161 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X297 a_n6972_8799.t35 a_n2848_n452.t94 a_n2650_8322.t17 vdd.t160 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X298 vdd.t35 vdd.t32 vdd.t34 vdd.t33 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X299 gnd.t42 gnd.t40 minus.t1 gnd.t41 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X300 a_n2848_n452.t5 minus.t24 a_n3106_n452.t32 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X301 a_n6972_8799.t40 plus.t23 a_n3106_n452.t11 gnd.t187 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X302 gnd.t39 gnd.t36 gnd.t38 gnd.t37 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X303 CSoutput.t118 commonsourceibias.t146 gnd.t238 gnd.t237 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X304 vdd.t31 vdd.t28 vdd.t30 vdd.t29 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X305 a_n2848_n452.t2 minus.t25 a_n3106_n452.t4 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X306 a_n2472_13878.t8 a_n2848_n452.t34 a_n2848_n452.t35 vdd.t159 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X307 output.t6 CSoutput.t146 vdd.t111 gnd.t138 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X308 commonsourceibias.t67 commonsourceibias.t66 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X309 vdd.t122 a_n6972_8799.t83 CSoutput.t32 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X310 gnd.t234 commonsourceibias.t147 CSoutput.t23 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X311 gnd.t233 commonsourceibias.t64 commonsourceibias.t65 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X312 CSoutput.t83 commonsourceibias.t148 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X313 gnd.t230 commonsourceibias.t149 CSoutput.t19 gnd.t229 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X314 gnd.t35 gnd.t32 gnd.t34 gnd.t33 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X315 a_n3106_n452.t54 minus.t26 a_n2848_n452.t62 gnd.t174 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X316 gnd.t228 commonsourceibias.t150 CSoutput.t11 gnd.t227 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 output.t5 CSoutput.t147 vdd.t4 gnd.t137 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X318 a_n3106_n452.t37 diffpairibias.t22 gnd.t171 gnd.t170 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X319 a_n6972_8799.t24 a_n2848_n452.t95 a_n2650_8322.t16 vdd.t158 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X320 a_n2848_n452.t39 a_n2848_n452.t38 a_n2472_13878.t7 vdd.t157 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X321 gnd.t226 commonsourceibias.t151 CSoutput.t10 gnd.t225 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 commonsourceibias.t51 commonsourceibias.t50 gnd.t224 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X323 CSoutput.t31 a_n6972_8799.t84 vdd.t23 vdd.t8 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X324 vdd.t144 a_n6972_8799.t85 CSoutput.t30 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X325 gnd.t223 commonsourceibias.t152 CSoutput.t2 gnd.t222 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X326 a_n6972_8799.t9 plus.t24 a_n3106_n452.t10 gnd.t169 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X327 gnd.t31 gnd.t28 gnd.t30 gnd.t29 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X328 CSoutput.t29 a_n6972_8799.t86 vdd.t145 vdd.t18 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X329 vdd.t119 a_n6972_8799.t87 CSoutput.t28 vdd.t6 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X330 diffpairibias.t3 diffpairibias.t2 gnd.t164 gnd.t163 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X331 a_n2650_8322.t15 a_n2848_n452.t96 a_n6972_8799.t19 vdd.t156 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X332 gnd.t16 gnd.t14 plus.t1 gnd.t15 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X333 a_n2848_n452.t1 minus.t27 a_n3106_n452.t1 gnd.t1 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X334 vdd.t143 a_n6972_8799.t88 CSoutput.t27 vdd.t124 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X335 gnd.t221 commonsourceibias.t153 CSoutput.t20 gnd.t220 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 commonsourceibias.t55 commonsourceibias.t54 gnd.t219 gnd.t218 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X337 CSoutput.t148 a_n2650_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X338 diffpairibias.t1 diffpairibias.t0 gnd.t155 gnd.t154 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X339 CSoutput.t21 commonsourceibias.t154 gnd.t217 gnd.t216 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X340 gnd.t27 gnd.t24 gnd.t26 gnd.t25 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X341 vdd.t155 a_n2848_n452.t97 a_n2472_13878.t27 vdd.t154 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X342 gnd.t23 gnd.t20 gnd.t22 gnd.t21 sky130_fd_pr__nfet_01v8 ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X343 commonsourceibias.t53 commonsourceibias.t52 gnd.t215 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X344 vdd.t204 a_n6972_8799.t89 CSoutput.t26 vdd.t21 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X345 plus.t0 gnd.t17 gnd.t19 gnd.t18 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X346 CSoutput.t22 commonsourceibias.t155 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X347 gnd.t212 commonsourceibias.t156 CSoutput.t123 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X348 CSoutput.t3 commonsourceibias.t157 gnd.t211 gnd.t210 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X349 vdd.t201 a_n6972_8799.t90 CSoutput.t25 vdd.t121 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X350 CSoutput.t24 a_n6972_8799.t91 vdd.t142 vdd.t139 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X351 CSoutput.t12 commonsourceibias.t158 gnd.t209 gnd.t208 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X352 commonsourceibias.t75 commonsourceibias.t74 gnd.t207 gnd.t206 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X353 gnd.t13 gnd.t11 minus.t0 gnd.t12 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X354 a_n6972_8799.t6 plus.t25 a_n3106_n452.t9 gnd.t133 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X355 vdd.t5 CSoutput.t149 output.t4 gnd.t136 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X356 gnd.t205 commonsourceibias.t72 commonsourceibias.t73 gnd.t204 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X357 a_n2650_8322.t14 a_n2848_n452.t98 a_n6972_8799.t33 vdd.t153 sky130_fd_pr__pfet_01v8 ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X358 CSoutput.t13 commonsourceibias.t159 gnd.t203 gnd.t202 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 a_n6972_8799.t13 plus.t26 a_n3106_n452.t8 gnd.t179 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X360 a_n2848_n452.t63 minus.t28 a_n3106_n452.t55 gnd.t180 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X361 gnd.t201 commonsourceibias.t70 commonsourceibias.t71 gnd.t200 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 commonsourceibias.t63 commonsourceibias.t62 gnd.t199 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X363 a_n2650_8322.t6 a_n2848_n452.t99 vdd.t152 vdd.t151 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X364 a_n2472_13878.t6 a_n2848_n452.t42 a_n2848_n452.t43 vdd.t150 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X365 gnd.t197 commonsourceibias.t60 commonsourceibias.t61 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X366 a_n3106_n452.t7 plus.t27 a_n6972_8799.t15 gnd.t183 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X367 commonsourceibias.t59 commonsourceibias.t58 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X368 a_n2848_n452.t45 a_n2848_n452.t44 a_n2472_13878.t5 vdd.t149 sky130_fd_pr__pfet_01v8 ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X369 a_n3106_n452.t6 plus.t28 a_n6972_8799.t10 gnd.t172 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X370 gnd.t193 commonsourceibias.t56 commonsourceibias.t57 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 a_n3106_n452.t45 diffpairibias.t23 gnd.t185 gnd.t184 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
R0 a_n2848_n452.n88 a_n2848_n452.t98 512.366
R1 a_n2848_n452.n87 a_n2848_n452.t77 512.366
R2 a_n2848_n452.n80 a_n2848_n452.t82 512.366
R3 a_n2848_n452.n86 a_n2848_n452.t71 512.366
R4 a_n2848_n452.n85 a_n2848_n452.t87 512.366
R5 a_n2848_n452.n81 a_n2848_n452.t95 512.366
R6 a_n2848_n452.n84 a_n2848_n452.t96 512.366
R7 a_n2848_n452.n83 a_n2848_n452.t66 512.366
R8 a_n2848_n452.n82 a_n2848_n452.t79 512.366
R9 a_n2848_n452.n61 a_n2848_n452.t42 533.335
R10 a_n2848_n452.n89 a_n2848_n452.t60 512.366
R11 a_n2848_n452.n90 a_n2848_n452.t34 512.366
R12 a_n2848_n452.n92 a_n2848_n452.t54 512.366
R13 a_n2848_n452.n109 a_n2848_n452.t28 512.366
R14 a_n2848_n452.n108 a_n2848_n452.t30 512.366
R15 a_n2848_n452.n79 a_n2848_n452.t40 512.366
R16 a_n2848_n452.n107 a_n2848_n452.t46 512.366
R17 a_n2848_n452.n106 a_n2848_n452.t38 512.366
R18 a_n2848_n452.n69 a_n2848_n452.t32 512.366
R19 a_n2848_n452.n136 a_n2848_n452.t24 512.366
R20 a_n2848_n452.n137 a_n2848_n452.t52 512.366
R21 a_n2848_n452.n76 a_n2848_n452.t44 512.366
R22 a_n2848_n452.n138 a_n2848_n452.t56 512.366
R23 a_n2848_n452.n139 a_n2848_n452.t36 512.366
R24 a_n2848_n452.n140 a_n2848_n452.t58 512.366
R25 a_n2848_n452.n141 a_n2848_n452.t50 512.366
R26 a_n2848_n452.n75 a_n2848_n452.t48 512.366
R27 a_n2848_n452.n142 a_n2848_n452.t26 512.366
R28 a_n2848_n452.n129 a_n2848_n452.t70 512.366
R29 a_n2848_n452.n130 a_n2848_n452.t94 512.366
R30 a_n2848_n452.n78 a_n2848_n452.t93 512.366
R31 a_n2848_n452.n131 a_n2848_n452.t68 512.366
R32 a_n2848_n452.n132 a_n2848_n452.t91 512.366
R33 a_n2848_n452.n133 a_n2848_n452.t90 512.366
R34 a_n2848_n452.n134 a_n2848_n452.t65 512.366
R35 a_n2848_n452.n77 a_n2848_n452.t75 512.366
R36 a_n2848_n452.n135 a_n2848_n452.t85 512.366
R37 a_n2848_n452.n121 a_n2848_n452.t84 512.366
R38 a_n2848_n452.n120 a_n2848_n452.t74 512.366
R39 a_n2848_n452.n119 a_n2848_n452.t64 512.366
R40 a_n2848_n452.n123 a_n2848_n452.t92 512.366
R41 a_n2848_n452.n122 a_n2848_n452.t81 512.366
R42 a_n2848_n452.n118 a_n2848_n452.t80 512.366
R43 a_n2848_n452.n125 a_n2848_n452.t88 512.366
R44 a_n2848_n452.n124 a_n2848_n452.t73 512.366
R45 a_n2848_n452.n117 a_n2848_n452.t72 512.366
R46 a_n2848_n452.n127 a_n2848_n452.t76 512.366
R47 a_n2848_n452.n126 a_n2848_n452.t86 512.366
R48 a_n2848_n452.n116 a_n2848_n452.t99 512.366
R49 a_n2848_n452.n6 a_n2848_n452.n68 70.1674
R50 a_n2848_n452.n10 a_n2848_n452.n70 70.1674
R51 a_n2848_n452.n22 a_n2848_n452.n47 70.1674
R52 a_n2848_n452.n26 a_n2848_n452.n40 70.1674
R53 a_n2848_n452.n135 a_n2848_n452.n40 20.9683
R54 a_n2848_n452.n39 a_n2848_n452.n26 74.73
R55 a_n2848_n452.n39 a_n2848_n452.n77 11.843
R56 a_n2848_n452.n25 a_n2848_n452.n38 80.4688
R57 a_n2848_n452.n134 a_n2848_n452.n38 0.365327
R58 a_n2848_n452.n37 a_n2848_n452.n25 75.0448
R59 a_n2848_n452.n27 a_n2848_n452.n36 70.1674
R60 a_n2848_n452.n131 a_n2848_n452.n36 20.9683
R61 a_n2848_n452.n35 a_n2848_n452.n27 70.3058
R62 a_n2848_n452.n35 a_n2848_n452.n78 20.6913
R63 a_n2848_n452.n28 a_n2848_n452.n34 75.3623
R64 a_n2848_n452.n130 a_n2848_n452.n34 10.5784
R65 a_n2848_n452.n129 a_n2848_n452.n28 161.3
R66 a_n2848_n452.n142 a_n2848_n452.n47 20.9683
R67 a_n2848_n452.n46 a_n2848_n452.n22 74.73
R68 a_n2848_n452.n46 a_n2848_n452.n75 11.843
R69 a_n2848_n452.n21 a_n2848_n452.n45 80.4688
R70 a_n2848_n452.n141 a_n2848_n452.n45 0.365327
R71 a_n2848_n452.n44 a_n2848_n452.n21 75.0448
R72 a_n2848_n452.n23 a_n2848_n452.n43 70.1674
R73 a_n2848_n452.n138 a_n2848_n452.n43 20.9683
R74 a_n2848_n452.n42 a_n2848_n452.n23 70.3058
R75 a_n2848_n452.n42 a_n2848_n452.n76 20.6913
R76 a_n2848_n452.n24 a_n2848_n452.n41 75.3623
R77 a_n2848_n452.n137 a_n2848_n452.n41 10.5784
R78 a_n2848_n452.n136 a_n2848_n452.n24 161.3
R79 a_n2848_n452.n13 a_n2848_n452.n56 70.1674
R80 a_n2848_n452.n15 a_n2848_n452.n53 70.1674
R81 a_n2848_n452.n17 a_n2848_n452.n51 70.1674
R82 a_n2848_n452.n19 a_n2848_n452.n49 70.1674
R83 a_n2848_n452.n49 a_n2848_n452.n116 20.9683
R84 a_n2848_n452.n48 a_n2848_n452.n20 75.0448
R85 a_n2848_n452.n126 a_n2848_n452.n48 11.2134
R86 a_n2848_n452.n20 a_n2848_n452.n127 161.3
R87 a_n2848_n452.n51 a_n2848_n452.n117 20.9683
R88 a_n2848_n452.n50 a_n2848_n452.n18 75.0448
R89 a_n2848_n452.n124 a_n2848_n452.n50 11.2134
R90 a_n2848_n452.n18 a_n2848_n452.n125 161.3
R91 a_n2848_n452.n53 a_n2848_n452.n118 20.9683
R92 a_n2848_n452.n52 a_n2848_n452.n16 75.0448
R93 a_n2848_n452.n122 a_n2848_n452.n52 11.2134
R94 a_n2848_n452.n16 a_n2848_n452.n123 161.3
R95 a_n2848_n452.n56 a_n2848_n452.n119 20.9683
R96 a_n2848_n452.n54 a_n2848_n452.n14 75.0448
R97 a_n2848_n452.n120 a_n2848_n452.n54 11.2134
R98 a_n2848_n452.n14 a_n2848_n452.n121 161.3
R99 a_n2848_n452.n105 a_n2848_n452.n10 161.3
R100 a_n2848_n452.n59 a_n2848_n452.n11 70.1674
R101 a_n2848_n452.n107 a_n2848_n452.n59 20.9683
R102 a_n2848_n452.n11 a_n2848_n452.n58 70.3058
R103 a_n2848_n452.n58 a_n2848_n452.n79 20.6913
R104 a_n2848_n452.n57 a_n2848_n452.n12 75.3623
R105 a_n2848_n452.n108 a_n2848_n452.n57 10.5784
R106 a_n2848_n452.n12 a_n2848_n452.n109 161.3
R107 a_n2848_n452.n70 a_n2848_n452.n92 20.9683
R108 a_n2848_n452.n61 a_n2848_n452.n9 70.1674
R109 a_n2848_n452.n61 a_n2848_n452.n89 20.9683
R110 a_n2848_n452.n10 a_n2848_n452.n60 74.73
R111 a_n2848_n452.n90 a_n2848_n452.n60 11.843
R112 a_n2848_n452.n91 a_n2848_n452.n10 161.3
R113 a_n2848_n452.n68 a_n2848_n452.n82 20.9683
R114 a_n2848_n452.n67 a_n2848_n452.n6 74.73
R115 a_n2848_n452.n83 a_n2848_n452.n67 11.843
R116 a_n2848_n452.n66 a_n2848_n452.n5 80.4688
R117 a_n2848_n452.n66 a_n2848_n452.n84 0.365327
R118 a_n2848_n452.n5 a_n2848_n452.n65 75.0448
R119 a_n2848_n452.n64 a_n2848_n452.n7 70.1674
R120 a_n2848_n452.n86 a_n2848_n452.n64 20.9683
R121 a_n2848_n452.n7 a_n2848_n452.n63 70.3058
R122 a_n2848_n452.n63 a_n2848_n452.n80 20.6913
R123 a_n2848_n452.n62 a_n2848_n452.n8 75.3623
R124 a_n2848_n452.n87 a_n2848_n452.n62 10.5784
R125 a_n2848_n452.n8 a_n2848_n452.n88 161.3
R126 a_n2848_n452.n3 a_n2848_n452.n102 81.4626
R127 a_n2848_n452.n4 a_n2848_n452.n96 81.4626
R128 a_n2848_n452.n0 a_n2848_n452.n93 81.4626
R129 a_n2848_n452.n3 a_n2848_n452.n103 80.9324
R130 a_n2848_n452.n2 a_n2848_n452.n104 80.9324
R131 a_n2848_n452.n2 a_n2848_n452.n101 80.9324
R132 a_n2848_n452.n2 a_n2848_n452.n100 80.9324
R133 a_n2848_n452.n1 a_n2848_n452.n99 80.9324
R134 a_n2848_n452.n4 a_n2848_n452.n97 80.9324
R135 a_n2848_n452.n0 a_n2848_n452.n98 80.9324
R136 a_n2848_n452.n0 a_n2848_n452.n95 80.9324
R137 a_n2848_n452.n0 a_n2848_n452.n94 80.9324
R138 a_n2848_n452.n31 a_n2848_n452.t25 74.6477
R139 a_n2848_n452.n29 a_n2848_n452.t43 74.6477
R140 a_n2848_n452.n114 a_n2848_n452.t29 74.2899
R141 a_n2848_n452.t23 a_n2848_n452.n33 74.2898
R142 a_n2848_n452.n33 a_n2848_n452.n74 70.6783
R143 a_n2848_n452.n32 a_n2848_n452.n73 70.6783
R144 a_n2848_n452.n32 a_n2848_n452.n72 70.6783
R145 a_n2848_n452.n31 a_n2848_n452.n71 70.6783
R146 a_n2848_n452.n29 a_n2848_n452.n110 70.6783
R147 a_n2848_n452.n29 a_n2848_n452.n111 70.6783
R148 a_n2848_n452.n30 a_n2848_n452.n112 70.6783
R149 a_n2848_n452.n30 a_n2848_n452.n113 70.6783
R150 a_n2848_n452.n88 a_n2848_n452.n87 48.2005
R151 a_n2848_n452.n64 a_n2848_n452.n85 20.9683
R152 a_n2848_n452.n84 a_n2848_n452.n81 48.2005
R153 a_n2848_n452.t69 a_n2848_n452.n68 533.335
R154 a_n2848_n452.n109 a_n2848_n452.n108 48.2005
R155 a_n2848_n452.n59 a_n2848_n452.n106 20.9683
R156 a_n2848_n452.n70 a_n2848_n452.n69 20.9683
R157 a_n2848_n452.n137 a_n2848_n452.n136 48.2005
R158 a_n2848_n452.n139 a_n2848_n452.n43 20.9683
R159 a_n2848_n452.n141 a_n2848_n452.n140 48.2005
R160 a_n2848_n452.t22 a_n2848_n452.n47 533.335
R161 a_n2848_n452.n130 a_n2848_n452.n129 48.2005
R162 a_n2848_n452.n132 a_n2848_n452.n36 20.9683
R163 a_n2848_n452.n134 a_n2848_n452.n133 48.2005
R164 a_n2848_n452.t67 a_n2848_n452.n40 533.335
R165 a_n2848_n452.n121 a_n2848_n452.n120 48.2005
R166 a_n2848_n452.t89 a_n2848_n452.n56 533.335
R167 a_n2848_n452.n123 a_n2848_n452.n122 48.2005
R168 a_n2848_n452.t97 a_n2848_n452.n53 533.335
R169 a_n2848_n452.n125 a_n2848_n452.n124 48.2005
R170 a_n2848_n452.t83 a_n2848_n452.n51 533.335
R171 a_n2848_n452.n127 a_n2848_n452.n126 48.2005
R172 a_n2848_n452.t78 a_n2848_n452.n49 533.335
R173 a_n2848_n452.n86 a_n2848_n452.n63 21.4216
R174 a_n2848_n452.n91 a_n2848_n452.n90 47.4702
R175 a_n2848_n452.n107 a_n2848_n452.n58 21.4216
R176 a_n2848_n452.n138 a_n2848_n452.n42 21.4216
R177 a_n2848_n452.n131 a_n2848_n452.n35 21.4216
R178 a_n2848_n452.n1 a_n2848_n452.n0 33.585
R179 a_n2848_n452.n67 a_n2848_n452.n82 34.4824
R180 a_n2848_n452.n60 a_n2848_n452.n89 34.4824
R181 a_n2848_n452.n142 a_n2848_n452.n46 34.4824
R182 a_n2848_n452.n135 a_n2848_n452.n39 34.4824
R183 a_n2848_n452.n85 a_n2848_n452.n65 35.3134
R184 a_n2848_n452.n65 a_n2848_n452.n81 11.2134
R185 a_n2848_n452.n106 a_n2848_n452.n105 24.1005
R186 a_n2848_n452.n105 a_n2848_n452.n69 24.1005
R187 a_n2848_n452.n139 a_n2848_n452.n44 35.3134
R188 a_n2848_n452.n140 a_n2848_n452.n44 11.2134
R189 a_n2848_n452.n132 a_n2848_n452.n37 35.3134
R190 a_n2848_n452.n133 a_n2848_n452.n37 11.2134
R191 a_n2848_n452.n54 a_n2848_n452.n119 35.3134
R192 a_n2848_n452.n52 a_n2848_n452.n118 35.3134
R193 a_n2848_n452.n50 a_n2848_n452.n117 35.3134
R194 a_n2848_n452.n48 a_n2848_n452.n116 35.3134
R195 a_n2848_n452.n10 a_n2848_n452.n2 23.891
R196 a_n2848_n452.n62 a_n2848_n452.n80 36.139
R197 a_n2848_n452.n57 a_n2848_n452.n79 36.139
R198 a_n2848_n452.n76 a_n2848_n452.n41 36.139
R199 a_n2848_n452.n78 a_n2848_n452.n34 36.139
R200 a_n2848_n452.n28 a_n2848_n452.n128 13.3641
R201 a_n2848_n452.n6 a_n2848_n452.n55 13.1596
R202 a_n2848_n452.n115 a_n2848_n452.n12 11.8547
R203 a_n2848_n452.n33 a_n2848_n452.n143 10.2167
R204 a_n2848_n452.n13 a_n2848_n452.n55 9.99103
R205 a_n2848_n452.n128 a_n2848_n452.n20 9.99103
R206 a_n2848_n452.n143 a_n2848_n452.n22 8.01944
R207 a_n2848_n452.n115 a_n2848_n452.n114 6.37334
R208 a_n2848_n452.n143 a_n2848_n452.n55 5.3452
R209 a_n2848_n452.n24 a_n2848_n452.n26 4.07247
R210 a_n2848_n452.n9 a_n2848_n452.n8 4.07247
R211 a_n2848_n452.n74 a_n2848_n452.t49 3.61217
R212 a_n2848_n452.n74 a_n2848_n452.t27 3.61217
R213 a_n2848_n452.n73 a_n2848_n452.t59 3.61217
R214 a_n2848_n452.n73 a_n2848_n452.t51 3.61217
R215 a_n2848_n452.n72 a_n2848_n452.t57 3.61217
R216 a_n2848_n452.n72 a_n2848_n452.t37 3.61217
R217 a_n2848_n452.n71 a_n2848_n452.t53 3.61217
R218 a_n2848_n452.n71 a_n2848_n452.t45 3.61217
R219 a_n2848_n452.n110 a_n2848_n452.t35 3.61217
R220 a_n2848_n452.n110 a_n2848_n452.t61 3.61217
R221 a_n2848_n452.n111 a_n2848_n452.t33 3.61217
R222 a_n2848_n452.n111 a_n2848_n452.t55 3.61217
R223 a_n2848_n452.n112 a_n2848_n452.t47 3.61217
R224 a_n2848_n452.n112 a_n2848_n452.t39 3.61217
R225 a_n2848_n452.n113 a_n2848_n452.t31 3.61217
R226 a_n2848_n452.n113 a_n2848_n452.t41 3.61217
R227 a_n2848_n452.n102 a_n2848_n452.t3 2.82907
R228 a_n2848_n452.n102 a_n2848_n452.t63 2.82907
R229 a_n2848_n452.n103 a_n2848_n452.t16 2.82907
R230 a_n2848_n452.n103 a_n2848_n452.t17 2.82907
R231 a_n2848_n452.n104 a_n2848_n452.t13 2.82907
R232 a_n2848_n452.n104 a_n2848_n452.t10 2.82907
R233 a_n2848_n452.n101 a_n2848_n452.t0 2.82907
R234 a_n2848_n452.n101 a_n2848_n452.t7 2.82907
R235 a_n2848_n452.n100 a_n2848_n452.t8 2.82907
R236 a_n2848_n452.n100 a_n2848_n452.t2 2.82907
R237 a_n2848_n452.n99 a_n2848_n452.t9 2.82907
R238 a_n2848_n452.n99 a_n2848_n452.t20 2.82907
R239 a_n2848_n452.n96 a_n2848_n452.t19 2.82907
R240 a_n2848_n452.n96 a_n2848_n452.t15 2.82907
R241 a_n2848_n452.n97 a_n2848_n452.t6 2.82907
R242 a_n2848_n452.n97 a_n2848_n452.t21 2.82907
R243 a_n2848_n452.n98 a_n2848_n452.t4 2.82907
R244 a_n2848_n452.n98 a_n2848_n452.t5 2.82907
R245 a_n2848_n452.n95 a_n2848_n452.t62 2.82907
R246 a_n2848_n452.n95 a_n2848_n452.t1 2.82907
R247 a_n2848_n452.n94 a_n2848_n452.t12 2.82907
R248 a_n2848_n452.n94 a_n2848_n452.t11 2.82907
R249 a_n2848_n452.n93 a_n2848_n452.t14 2.82907
R250 a_n2848_n452.n93 a_n2848_n452.t18 2.82907
R251 a_n2848_n452.n128 a_n2848_n452.n115 1.30542
R252 a_n2848_n452.n17 a_n2848_n452.n16 1.04595
R253 a_n2848_n452.n66 a_n2848_n452.n83 47.835
R254 a_n2848_n452.n92 a_n2848_n452.n91 0.730803
R255 a_n2848_n452.n75 a_n2848_n452.n45 47.835
R256 a_n2848_n452.n77 a_n2848_n452.n38 47.835
R257 a_n2848_n452.n0 a_n2848_n452.n4 1.59102
R258 a_n2848_n452.n26 a_n2848_n452.n25 1.13686
R259 a_n2848_n452.n22 a_n2848_n452.n21 1.13686
R260 a_n2848_n452.n6 a_n2848_n452.n5 1.13686
R261 a_n2848_n452.n10 a_n2848_n452.n11 1.09898
R262 a_n2848_n452.n2 a_n2848_n452.n3 1.06084
R263 a_n2848_n452.n2 a_n2848_n452.n1 1.06084
R264 a_n2848_n452.n27 a_n2848_n452.n28 0.758076
R265 a_n2848_n452.n25 a_n2848_n452.n27 0.758076
R266 a_n2848_n452.n23 a_n2848_n452.n24 0.758076
R267 a_n2848_n452.n21 a_n2848_n452.n23 0.758076
R268 a_n2848_n452.n20 a_n2848_n452.n19 0.758076
R269 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R270 a_n2848_n452.n16 a_n2848_n452.n15 0.758076
R271 a_n2848_n452.n14 a_n2848_n452.n13 0.758076
R272 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R273 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R274 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R275 a_n2848_n452.n5 a_n2848_n452.n7 0.758076
R276 a_n2848_n452.n33 a_n2848_n452.n32 0.716017
R277 a_n2848_n452.n32 a_n2848_n452.n31 0.716017
R278 a_n2848_n452.n30 a_n2848_n452.n29 0.716017
R279 a_n2848_n452.n114 a_n2848_n452.n30 0.716017
R280 a_n2848_n452.n19 a_n2848_n452.n18 0.67853
R281 a_n2848_n452.n15 a_n2848_n452.n14 0.67853
R282 a_n2472_13878.n25 a_n2472_13878.n24 98.9632
R283 a_n2472_13878.n2 a_n2472_13878.n0 98.7517
R284 a_n2472_13878.n20 a_n2472_13878.n19 98.6055
R285 a_n2472_13878.n22 a_n2472_13878.n21 98.6055
R286 a_n2472_13878.n24 a_n2472_13878.n23 98.6055
R287 a_n2472_13878.n8 a_n2472_13878.n7 98.6055
R288 a_n2472_13878.n6 a_n2472_13878.n5 98.6055
R289 a_n2472_13878.n4 a_n2472_13878.n3 98.6055
R290 a_n2472_13878.n2 a_n2472_13878.n1 98.6055
R291 a_n2472_13878.n18 a_n2472_13878.n17 98.6054
R292 a_n2472_13878.n10 a_n2472_13878.t1 74.6477
R293 a_n2472_13878.n15 a_n2472_13878.t4 74.2899
R294 a_n2472_13878.n12 a_n2472_13878.t2 74.2899
R295 a_n2472_13878.n11 a_n2472_13878.t27 74.2899
R296 a_n2472_13878.n14 a_n2472_13878.n13 70.6783
R297 a_n2472_13878.n10 a_n2472_13878.n9 70.6783
R298 a_n2472_13878.n16 a_n2472_13878.n8 15.0004
R299 a_n2472_13878.n18 a_n2472_13878.n16 12.2917
R300 a_n2472_13878.n16 a_n2472_13878.n15 7.67184
R301 a_n2472_13878.n17 a_n2472_13878.t21 3.61217
R302 a_n2472_13878.n17 a_n2472_13878.t10 3.61217
R303 a_n2472_13878.n19 a_n2472_13878.t13 3.61217
R304 a_n2472_13878.n19 a_n2472_13878.t14 3.61217
R305 a_n2472_13878.n21 a_n2472_13878.t22 3.61217
R306 a_n2472_13878.n21 a_n2472_13878.t23 3.61217
R307 a_n2472_13878.n23 a_n2472_13878.t5 3.61217
R308 a_n2472_13878.n23 a_n2472_13878.t15 3.61217
R309 a_n2472_13878.n13 a_n2472_13878.t0 3.61217
R310 a_n2472_13878.n13 a_n2472_13878.t3 3.61217
R311 a_n2472_13878.n9 a_n2472_13878.t25 3.61217
R312 a_n2472_13878.n9 a_n2472_13878.t26 3.61217
R313 a_n2472_13878.n7 a_n2472_13878.t16 3.61217
R314 a_n2472_13878.n7 a_n2472_13878.t6 3.61217
R315 a_n2472_13878.n5 a_n2472_13878.t19 3.61217
R316 a_n2472_13878.n5 a_n2472_13878.t8 3.61217
R317 a_n2472_13878.n3 a_n2472_13878.t7 3.61217
R318 a_n2472_13878.n3 a_n2472_13878.t9 3.61217
R319 a_n2472_13878.n1 a_n2472_13878.t17 3.61217
R320 a_n2472_13878.n1 a_n2472_13878.t11 3.61217
R321 a_n2472_13878.n0 a_n2472_13878.t20 3.61217
R322 a_n2472_13878.n0 a_n2472_13878.t12 3.61217
R323 a_n2472_13878.n25 a_n2472_13878.t18 3.61217
R324 a_n2472_13878.t24 a_n2472_13878.n25 3.61217
R325 a_n2472_13878.n11 a_n2472_13878.n10 0.358259
R326 a_n2472_13878.n14 a_n2472_13878.n12 0.358259
R327 a_n2472_13878.n15 a_n2472_13878.n14 0.358259
R328 a_n2472_13878.n24 a_n2472_13878.n22 0.358259
R329 a_n2472_13878.n22 a_n2472_13878.n20 0.358259
R330 a_n2472_13878.n20 a_n2472_13878.n18 0.358259
R331 a_n2472_13878.n4 a_n2472_13878.n2 0.146627
R332 a_n2472_13878.n6 a_n2472_13878.n4 0.146627
R333 a_n2472_13878.n8 a_n2472_13878.n6 0.146627
R334 a_n2472_13878.n12 a_n2472_13878.n11 0.101793
R335 vdd.n291 vdd.n255 756.745
R336 vdd.n244 vdd.n208 756.745
R337 vdd.n201 vdd.n165 756.745
R338 vdd.n154 vdd.n118 756.745
R339 vdd.n112 vdd.n76 756.745
R340 vdd.n65 vdd.n29 756.745
R341 vdd.n1186 vdd.n1150 756.745
R342 vdd.n1233 vdd.n1197 756.745
R343 vdd.n1096 vdd.n1060 756.745
R344 vdd.n1143 vdd.n1107 756.745
R345 vdd.n1007 vdd.n971 756.745
R346 vdd.n1054 vdd.n1018 756.745
R347 vdd.n926 vdd.t44 640.208
R348 vdd.n787 vdd.t74 640.208
R349 vdd.n920 vdd.t95 640.208
R350 vdd.n778 vdd.t92 640.208
R351 vdd.n675 vdd.t54 640.208
R352 vdd.n2375 vdd.t89 640.208
R353 vdd.n622 vdd.t68 640.208
R354 vdd.n2444 vdd.t78 640.208
R355 vdd.n589 vdd.t40 640.208
R356 vdd.n848 vdd.t85 640.208
R357 vdd.n1400 vdd.t32 592.009
R358 vdd.n1438 vdd.t48 592.009
R359 vdd.n1334 vdd.t65 592.009
R360 vdd.n1814 vdd.t61 592.009
R361 vdd.n1664 vdd.t71 592.009
R362 vdd.n1624 vdd.t82 592.009
R363 vdd.n3090 vdd.t28 592.009
R364 vdd.n405 vdd.t98 592.009
R365 vdd.n365 vdd.t101 592.009
R366 vdd.n557 vdd.t36 592.009
R367 vdd.n2986 vdd.t51 592.009
R368 vdd.n2893 vdd.t58 592.009
R369 vdd.n292 vdd.n291 585
R370 vdd.n290 vdd.n257 585
R371 vdd.n289 vdd.n288 585
R372 vdd.n260 vdd.n258 585
R373 vdd.n283 vdd.n282 585
R374 vdd.n281 vdd.n280 585
R375 vdd.n264 vdd.n263 585
R376 vdd.n275 vdd.n274 585
R377 vdd.n273 vdd.n272 585
R378 vdd.n268 vdd.n267 585
R379 vdd.n245 vdd.n244 585
R380 vdd.n243 vdd.n210 585
R381 vdd.n242 vdd.n241 585
R382 vdd.n213 vdd.n211 585
R383 vdd.n236 vdd.n235 585
R384 vdd.n234 vdd.n233 585
R385 vdd.n217 vdd.n216 585
R386 vdd.n228 vdd.n227 585
R387 vdd.n226 vdd.n225 585
R388 vdd.n221 vdd.n220 585
R389 vdd.n202 vdd.n201 585
R390 vdd.n200 vdd.n167 585
R391 vdd.n199 vdd.n198 585
R392 vdd.n170 vdd.n168 585
R393 vdd.n193 vdd.n192 585
R394 vdd.n191 vdd.n190 585
R395 vdd.n174 vdd.n173 585
R396 vdd.n185 vdd.n184 585
R397 vdd.n183 vdd.n182 585
R398 vdd.n178 vdd.n177 585
R399 vdd.n155 vdd.n154 585
R400 vdd.n153 vdd.n120 585
R401 vdd.n152 vdd.n151 585
R402 vdd.n123 vdd.n121 585
R403 vdd.n146 vdd.n145 585
R404 vdd.n144 vdd.n143 585
R405 vdd.n127 vdd.n126 585
R406 vdd.n138 vdd.n137 585
R407 vdd.n136 vdd.n135 585
R408 vdd.n131 vdd.n130 585
R409 vdd.n113 vdd.n112 585
R410 vdd.n111 vdd.n78 585
R411 vdd.n110 vdd.n109 585
R412 vdd.n81 vdd.n79 585
R413 vdd.n104 vdd.n103 585
R414 vdd.n102 vdd.n101 585
R415 vdd.n85 vdd.n84 585
R416 vdd.n96 vdd.n95 585
R417 vdd.n94 vdd.n93 585
R418 vdd.n89 vdd.n88 585
R419 vdd.n66 vdd.n65 585
R420 vdd.n64 vdd.n31 585
R421 vdd.n63 vdd.n62 585
R422 vdd.n34 vdd.n32 585
R423 vdd.n57 vdd.n56 585
R424 vdd.n55 vdd.n54 585
R425 vdd.n38 vdd.n37 585
R426 vdd.n49 vdd.n48 585
R427 vdd.n47 vdd.n46 585
R428 vdd.n42 vdd.n41 585
R429 vdd.n1187 vdd.n1186 585
R430 vdd.n1185 vdd.n1152 585
R431 vdd.n1184 vdd.n1183 585
R432 vdd.n1155 vdd.n1153 585
R433 vdd.n1178 vdd.n1177 585
R434 vdd.n1176 vdd.n1175 585
R435 vdd.n1159 vdd.n1158 585
R436 vdd.n1170 vdd.n1169 585
R437 vdd.n1168 vdd.n1167 585
R438 vdd.n1163 vdd.n1162 585
R439 vdd.n1234 vdd.n1233 585
R440 vdd.n1232 vdd.n1199 585
R441 vdd.n1231 vdd.n1230 585
R442 vdd.n1202 vdd.n1200 585
R443 vdd.n1225 vdd.n1224 585
R444 vdd.n1223 vdd.n1222 585
R445 vdd.n1206 vdd.n1205 585
R446 vdd.n1217 vdd.n1216 585
R447 vdd.n1215 vdd.n1214 585
R448 vdd.n1210 vdd.n1209 585
R449 vdd.n1097 vdd.n1096 585
R450 vdd.n1095 vdd.n1062 585
R451 vdd.n1094 vdd.n1093 585
R452 vdd.n1065 vdd.n1063 585
R453 vdd.n1088 vdd.n1087 585
R454 vdd.n1086 vdd.n1085 585
R455 vdd.n1069 vdd.n1068 585
R456 vdd.n1080 vdd.n1079 585
R457 vdd.n1078 vdd.n1077 585
R458 vdd.n1073 vdd.n1072 585
R459 vdd.n1144 vdd.n1143 585
R460 vdd.n1142 vdd.n1109 585
R461 vdd.n1141 vdd.n1140 585
R462 vdd.n1112 vdd.n1110 585
R463 vdd.n1135 vdd.n1134 585
R464 vdd.n1133 vdd.n1132 585
R465 vdd.n1116 vdd.n1115 585
R466 vdd.n1127 vdd.n1126 585
R467 vdd.n1125 vdd.n1124 585
R468 vdd.n1120 vdd.n1119 585
R469 vdd.n1008 vdd.n1007 585
R470 vdd.n1006 vdd.n973 585
R471 vdd.n1005 vdd.n1004 585
R472 vdd.n976 vdd.n974 585
R473 vdd.n999 vdd.n998 585
R474 vdd.n997 vdd.n996 585
R475 vdd.n980 vdd.n979 585
R476 vdd.n991 vdd.n990 585
R477 vdd.n989 vdd.n988 585
R478 vdd.n984 vdd.n983 585
R479 vdd.n1055 vdd.n1054 585
R480 vdd.n1053 vdd.n1020 585
R481 vdd.n1052 vdd.n1051 585
R482 vdd.n1023 vdd.n1021 585
R483 vdd.n1046 vdd.n1045 585
R484 vdd.n1044 vdd.n1043 585
R485 vdd.n1027 vdd.n1026 585
R486 vdd.n1038 vdd.n1037 585
R487 vdd.n1036 vdd.n1035 585
R488 vdd.n1031 vdd.n1030 585
R489 vdd.n3206 vdd.n330 515.122
R490 vdd.n3088 vdd.n328 515.122
R491 vdd.n515 vdd.n478 515.122
R492 vdd.n3024 vdd.n479 515.122
R493 vdd.n1809 vdd.n945 515.122
R494 vdd.n1812 vdd.n1811 515.122
R495 vdd.n1307 vdd.n1271 515.122
R496 vdd.n1503 vdd.n1272 515.122
R497 vdd.n269 vdd.t9 329.043
R498 vdd.n222 vdd.t3 329.043
R499 vdd.n179 vdd.t146 329.043
R500 vdd.n132 vdd.t14 329.043
R501 vdd.n90 vdd.t23 329.043
R502 vdd.n43 vdd.t108 329.043
R503 vdd.n1164 vdd.t16 329.043
R504 vdd.n1211 vdd.t122 329.043
R505 vdd.n1074 vdd.t112 329.043
R506 vdd.n1121 vdd.t201 329.043
R507 vdd.n985 vdd.t203 329.043
R508 vdd.n1032 vdd.t144 329.043
R509 vdd.n1400 vdd.t35 319.788
R510 vdd.n1438 vdd.t50 319.788
R511 vdd.n1334 vdd.t67 319.788
R512 vdd.n1814 vdd.t63 319.788
R513 vdd.n1664 vdd.t72 319.788
R514 vdd.n1624 vdd.t83 319.788
R515 vdd.n3090 vdd.t30 319.788
R516 vdd.n405 vdd.t99 319.788
R517 vdd.n365 vdd.t102 319.788
R518 vdd.n557 vdd.t39 319.788
R519 vdd.n2986 vdd.t53 319.788
R520 vdd.n2893 vdd.t60 319.788
R521 vdd.n1401 vdd.t34 303.69
R522 vdd.n1439 vdd.t49 303.69
R523 vdd.n1335 vdd.t66 303.69
R524 vdd.n1815 vdd.t64 303.69
R525 vdd.n1665 vdd.t73 303.69
R526 vdd.n1625 vdd.t84 303.69
R527 vdd.n3091 vdd.t31 303.69
R528 vdd.n406 vdd.t100 303.69
R529 vdd.n366 vdd.t103 303.69
R530 vdd.n558 vdd.t38 303.69
R531 vdd.n2987 vdd.t52 303.69
R532 vdd.n2894 vdd.t59 303.69
R533 vdd.n2630 vdd.n737 285.366
R534 vdd.n2854 vdd.n599 285.366
R535 vdd.n2791 vdd.n596 285.366
R536 vdd.n2509 vdd.n734 285.366
R537 vdd.n2339 vdd.n775 285.366
R538 vdd.n2270 vdd.n2269 285.366
R539 vdd.n2010 vdd.n901 285.366
R540 vdd.n2080 vdd.n903 285.366
R541 vdd.n2770 vdd.n597 285.366
R542 vdd.n2857 vdd.n2856 285.366
R543 vdd.n2623 vdd.n735 285.366
R544 vdd.n2632 vdd.n733 285.366
R545 vdd.n2267 vdd.n785 285.366
R546 vdd.n783 vdd.n757 285.366
R547 vdd.n1896 vdd.n902 285.366
R548 vdd.n2082 vdd.n899 285.366
R549 vdd.n943 vdd.n900 216.982
R550 vdd.n3022 vdd.n484 216.982
R551 vdd.n2772 vdd.n597 185
R552 vdd.n2855 vdd.n597 185
R553 vdd.n2774 vdd.n2773 185
R554 vdd.n2773 vdd.n595 185
R555 vdd.n2775 vdd.n629 185
R556 vdd.n2785 vdd.n629 185
R557 vdd.n2776 vdd.n638 185
R558 vdd.n638 vdd.n636 185
R559 vdd.n2778 vdd.n2777 185
R560 vdd.n2779 vdd.n2778 185
R561 vdd.n2731 vdd.n637 185
R562 vdd.n637 vdd.n633 185
R563 vdd.n2730 vdd.n2729 185
R564 vdd.n2729 vdd.n2728 185
R565 vdd.n640 vdd.n639 185
R566 vdd.n641 vdd.n640 185
R567 vdd.n2721 vdd.n2720 185
R568 vdd.n2722 vdd.n2721 185
R569 vdd.n2719 vdd.n649 185
R570 vdd.n654 vdd.n649 185
R571 vdd.n2718 vdd.n2717 185
R572 vdd.n2717 vdd.n2716 185
R573 vdd.n651 vdd.n650 185
R574 vdd.n660 vdd.n651 185
R575 vdd.n2709 vdd.n2708 185
R576 vdd.n2710 vdd.n2709 185
R577 vdd.n2707 vdd.n661 185
R578 vdd.n667 vdd.n661 185
R579 vdd.n2706 vdd.n2705 185
R580 vdd.n2705 vdd.n2704 185
R581 vdd.n663 vdd.n662 185
R582 vdd.n664 vdd.n663 185
R583 vdd.n2697 vdd.n2696 185
R584 vdd.n2698 vdd.n2697 185
R585 vdd.n2695 vdd.n674 185
R586 vdd.n674 vdd.n671 185
R587 vdd.n2693 vdd.n2692 185
R588 vdd.n2692 vdd.n2691 185
R589 vdd.n677 vdd.n676 185
R590 vdd.n678 vdd.n677 185
R591 vdd.n2684 vdd.n2683 185
R592 vdd.n2685 vdd.n2684 185
R593 vdd.n2682 vdd.n686 185
R594 vdd.n691 vdd.n686 185
R595 vdd.n2681 vdd.n2680 185
R596 vdd.n2680 vdd.n2679 185
R597 vdd.n688 vdd.n687 185
R598 vdd.n2591 vdd.n688 185
R599 vdd.n2672 vdd.n2671 185
R600 vdd.n2673 vdd.n2672 185
R601 vdd.n2670 vdd.n698 185
R602 vdd.n698 vdd.n695 185
R603 vdd.n2669 vdd.n2668 185
R604 vdd.n2668 vdd.n2667 185
R605 vdd.n700 vdd.n699 185
R606 vdd.n701 vdd.n700 185
R607 vdd.n2660 vdd.n2659 185
R608 vdd.n2661 vdd.n2660 185
R609 vdd.n2658 vdd.n709 185
R610 vdd.n2603 vdd.n709 185
R611 vdd.n2657 vdd.n2656 185
R612 vdd.n2656 vdd.n2655 185
R613 vdd.n711 vdd.n710 185
R614 vdd.n720 vdd.n711 185
R615 vdd.n2648 vdd.n2647 185
R616 vdd.n2649 vdd.n2648 185
R617 vdd.n2646 vdd.n721 185
R618 vdd.n721 vdd.n717 185
R619 vdd.n2645 vdd.n2644 185
R620 vdd.n2644 vdd.n2643 185
R621 vdd.n723 vdd.n722 185
R622 vdd.n2615 vdd.n723 185
R623 vdd.n2636 vdd.n2635 185
R624 vdd.n2637 vdd.n2636 185
R625 vdd.n2634 vdd.n731 185
R626 vdd.n736 vdd.n731 185
R627 vdd.n2633 vdd.n2632 185
R628 vdd.n2632 vdd.n2631 185
R629 vdd.n733 vdd.n732 185
R630 vdd.n2379 vdd.n2378 185
R631 vdd.n2381 vdd.n2380 185
R632 vdd.n2383 vdd.n2382 185
R633 vdd.n2385 vdd.n2384 185
R634 vdd.n2387 vdd.n2386 185
R635 vdd.n2389 vdd.n2388 185
R636 vdd.n2391 vdd.n2390 185
R637 vdd.n2393 vdd.n2392 185
R638 vdd.n2395 vdd.n2394 185
R639 vdd.n2397 vdd.n2396 185
R640 vdd.n2399 vdd.n2398 185
R641 vdd.n2401 vdd.n2400 185
R642 vdd.n2403 vdd.n2402 185
R643 vdd.n2405 vdd.n2404 185
R644 vdd.n2407 vdd.n2406 185
R645 vdd.n2409 vdd.n2408 185
R646 vdd.n2411 vdd.n2410 185
R647 vdd.n2413 vdd.n2412 185
R648 vdd.n2415 vdd.n2414 185
R649 vdd.n2417 vdd.n2416 185
R650 vdd.n2419 vdd.n2418 185
R651 vdd.n2421 vdd.n2420 185
R652 vdd.n2423 vdd.n2422 185
R653 vdd.n2425 vdd.n2424 185
R654 vdd.n2427 vdd.n2426 185
R655 vdd.n2429 vdd.n2428 185
R656 vdd.n2431 vdd.n2430 185
R657 vdd.n2433 vdd.n2432 185
R658 vdd.n2435 vdd.n2434 185
R659 vdd.n2437 vdd.n2436 185
R660 vdd.n2439 vdd.n2438 185
R661 vdd.n2441 vdd.n2440 185
R662 vdd.n2442 vdd.n2374 185
R663 vdd.n2623 vdd.n2622 185
R664 vdd.n2624 vdd.n2623 185
R665 vdd.n2858 vdd.n2857 185
R666 vdd.n2859 vdd.n588 185
R667 vdd.n2861 vdd.n2860 185
R668 vdd.n2863 vdd.n586 185
R669 vdd.n2865 vdd.n2864 185
R670 vdd.n2866 vdd.n585 185
R671 vdd.n2868 vdd.n2867 185
R672 vdd.n2870 vdd.n583 185
R673 vdd.n2872 vdd.n2871 185
R674 vdd.n2873 vdd.n582 185
R675 vdd.n2875 vdd.n2874 185
R676 vdd.n2877 vdd.n580 185
R677 vdd.n2879 vdd.n2878 185
R678 vdd.n2880 vdd.n579 185
R679 vdd.n2882 vdd.n2881 185
R680 vdd.n2884 vdd.n578 185
R681 vdd.n2885 vdd.n576 185
R682 vdd.n2888 vdd.n2887 185
R683 vdd.n577 vdd.n575 185
R684 vdd.n2744 vdd.n2743 185
R685 vdd.n2746 vdd.n2745 185
R686 vdd.n2748 vdd.n2740 185
R687 vdd.n2750 vdd.n2749 185
R688 vdd.n2751 vdd.n2739 185
R689 vdd.n2753 vdd.n2752 185
R690 vdd.n2755 vdd.n2737 185
R691 vdd.n2757 vdd.n2756 185
R692 vdd.n2758 vdd.n2736 185
R693 vdd.n2760 vdd.n2759 185
R694 vdd.n2762 vdd.n2734 185
R695 vdd.n2764 vdd.n2763 185
R696 vdd.n2765 vdd.n2733 185
R697 vdd.n2767 vdd.n2766 185
R698 vdd.n2769 vdd.n2732 185
R699 vdd.n2771 vdd.n2770 185
R700 vdd.n2770 vdd.n484 185
R701 vdd.n2856 vdd.n592 185
R702 vdd.n2856 vdd.n2855 185
R703 vdd.n2522 vdd.n594 185
R704 vdd.n595 vdd.n594 185
R705 vdd.n2523 vdd.n628 185
R706 vdd.n2785 vdd.n628 185
R707 vdd.n2525 vdd.n2524 185
R708 vdd.n2524 vdd.n636 185
R709 vdd.n2526 vdd.n635 185
R710 vdd.n2779 vdd.n635 185
R711 vdd.n2528 vdd.n2527 185
R712 vdd.n2527 vdd.n633 185
R713 vdd.n2529 vdd.n643 185
R714 vdd.n2728 vdd.n643 185
R715 vdd.n2531 vdd.n2530 185
R716 vdd.n2530 vdd.n641 185
R717 vdd.n2532 vdd.n648 185
R718 vdd.n2722 vdd.n648 185
R719 vdd.n2534 vdd.n2533 185
R720 vdd.n2533 vdd.n654 185
R721 vdd.n2535 vdd.n653 185
R722 vdd.n2716 vdd.n653 185
R723 vdd.n2537 vdd.n2536 185
R724 vdd.n2536 vdd.n660 185
R725 vdd.n2538 vdd.n659 185
R726 vdd.n2710 vdd.n659 185
R727 vdd.n2540 vdd.n2539 185
R728 vdd.n2539 vdd.n667 185
R729 vdd.n2541 vdd.n666 185
R730 vdd.n2704 vdd.n666 185
R731 vdd.n2543 vdd.n2542 185
R732 vdd.n2542 vdd.n664 185
R733 vdd.n2544 vdd.n673 185
R734 vdd.n2698 vdd.n673 185
R735 vdd.n2546 vdd.n2545 185
R736 vdd.n2545 vdd.n671 185
R737 vdd.n2547 vdd.n680 185
R738 vdd.n2691 vdd.n680 185
R739 vdd.n2549 vdd.n2548 185
R740 vdd.n2548 vdd.n678 185
R741 vdd.n2550 vdd.n685 185
R742 vdd.n2685 vdd.n685 185
R743 vdd.n2552 vdd.n2551 185
R744 vdd.n2551 vdd.n691 185
R745 vdd.n2553 vdd.n690 185
R746 vdd.n2679 vdd.n690 185
R747 vdd.n2593 vdd.n2592 185
R748 vdd.n2592 vdd.n2591 185
R749 vdd.n2594 vdd.n697 185
R750 vdd.n2673 vdd.n697 185
R751 vdd.n2596 vdd.n2595 185
R752 vdd.n2595 vdd.n695 185
R753 vdd.n2597 vdd.n703 185
R754 vdd.n2667 vdd.n703 185
R755 vdd.n2599 vdd.n2598 185
R756 vdd.n2598 vdd.n701 185
R757 vdd.n2600 vdd.n708 185
R758 vdd.n2661 vdd.n708 185
R759 vdd.n2602 vdd.n2601 185
R760 vdd.n2603 vdd.n2602 185
R761 vdd.n2521 vdd.n713 185
R762 vdd.n2655 vdd.n713 185
R763 vdd.n2520 vdd.n2519 185
R764 vdd.n2519 vdd.n720 185
R765 vdd.n2518 vdd.n719 185
R766 vdd.n2649 vdd.n719 185
R767 vdd.n2517 vdd.n2516 185
R768 vdd.n2516 vdd.n717 185
R769 vdd.n2443 vdd.n725 185
R770 vdd.n2643 vdd.n725 185
R771 vdd.n2617 vdd.n2616 185
R772 vdd.n2616 vdd.n2615 185
R773 vdd.n2618 vdd.n730 185
R774 vdd.n2637 vdd.n730 185
R775 vdd.n2620 vdd.n2619 185
R776 vdd.n2619 vdd.n736 185
R777 vdd.n2621 vdd.n735 185
R778 vdd.n2631 vdd.n735 185
R779 vdd.n1809 vdd.n1808 185
R780 vdd.n1810 vdd.n1809 185
R781 vdd.n946 vdd.n944 185
R782 vdd.n1588 vdd.n944 185
R783 vdd.n1591 vdd.n1590 185
R784 vdd.n1590 vdd.n1589 185
R785 vdd.n949 vdd.n948 185
R786 vdd.n950 vdd.n949 185
R787 vdd.n1577 vdd.n1576 185
R788 vdd.n1578 vdd.n1577 185
R789 vdd.n958 vdd.n957 185
R790 vdd.n1569 vdd.n957 185
R791 vdd.n1572 vdd.n1571 185
R792 vdd.n1571 vdd.n1570 185
R793 vdd.n961 vdd.n960 185
R794 vdd.n968 vdd.n961 185
R795 vdd.n1560 vdd.n1559 185
R796 vdd.n1561 vdd.n1560 185
R797 vdd.n970 vdd.n969 185
R798 vdd.n969 vdd.n967 185
R799 vdd.n1555 vdd.n1554 185
R800 vdd.n1554 vdd.n1553 185
R801 vdd.n1243 vdd.n1242 185
R802 vdd.n1244 vdd.n1243 185
R803 vdd.n1544 vdd.n1543 185
R804 vdd.n1545 vdd.n1544 185
R805 vdd.n1251 vdd.n1250 185
R806 vdd.n1535 vdd.n1250 185
R807 vdd.n1538 vdd.n1537 185
R808 vdd.n1537 vdd.n1536 185
R809 vdd.n1254 vdd.n1253 185
R810 vdd.n1260 vdd.n1254 185
R811 vdd.n1526 vdd.n1525 185
R812 vdd.n1527 vdd.n1526 185
R813 vdd.n1262 vdd.n1261 185
R814 vdd.n1518 vdd.n1261 185
R815 vdd.n1521 vdd.n1520 185
R816 vdd.n1520 vdd.n1519 185
R817 vdd.n1265 vdd.n1264 185
R818 vdd.n1266 vdd.n1265 185
R819 vdd.n1509 vdd.n1508 185
R820 vdd.n1510 vdd.n1509 185
R821 vdd.n1273 vdd.n1272 185
R822 vdd.n1308 vdd.n1272 185
R823 vdd.n1504 vdd.n1503 185
R824 vdd.n1276 vdd.n1275 185
R825 vdd.n1500 vdd.n1499 185
R826 vdd.n1501 vdd.n1500 185
R827 vdd.n1310 vdd.n1309 185
R828 vdd.n1495 vdd.n1312 185
R829 vdd.n1494 vdd.n1313 185
R830 vdd.n1493 vdd.n1314 185
R831 vdd.n1316 vdd.n1315 185
R832 vdd.n1489 vdd.n1318 185
R833 vdd.n1488 vdd.n1319 185
R834 vdd.n1487 vdd.n1320 185
R835 vdd.n1322 vdd.n1321 185
R836 vdd.n1483 vdd.n1324 185
R837 vdd.n1482 vdd.n1325 185
R838 vdd.n1481 vdd.n1326 185
R839 vdd.n1328 vdd.n1327 185
R840 vdd.n1477 vdd.n1330 185
R841 vdd.n1476 vdd.n1331 185
R842 vdd.n1475 vdd.n1332 185
R843 vdd.n1336 vdd.n1333 185
R844 vdd.n1471 vdd.n1338 185
R845 vdd.n1470 vdd.n1339 185
R846 vdd.n1469 vdd.n1340 185
R847 vdd.n1342 vdd.n1341 185
R848 vdd.n1465 vdd.n1344 185
R849 vdd.n1464 vdd.n1345 185
R850 vdd.n1463 vdd.n1346 185
R851 vdd.n1348 vdd.n1347 185
R852 vdd.n1459 vdd.n1350 185
R853 vdd.n1458 vdd.n1351 185
R854 vdd.n1457 vdd.n1352 185
R855 vdd.n1354 vdd.n1353 185
R856 vdd.n1453 vdd.n1356 185
R857 vdd.n1452 vdd.n1357 185
R858 vdd.n1451 vdd.n1358 185
R859 vdd.n1360 vdd.n1359 185
R860 vdd.n1447 vdd.n1362 185
R861 vdd.n1446 vdd.n1363 185
R862 vdd.n1445 vdd.n1364 185
R863 vdd.n1366 vdd.n1365 185
R864 vdd.n1441 vdd.n1368 185
R865 vdd.n1440 vdd.n1437 185
R866 vdd.n1436 vdd.n1369 185
R867 vdd.n1371 vdd.n1370 185
R868 vdd.n1432 vdd.n1373 185
R869 vdd.n1431 vdd.n1374 185
R870 vdd.n1430 vdd.n1375 185
R871 vdd.n1377 vdd.n1376 185
R872 vdd.n1426 vdd.n1379 185
R873 vdd.n1425 vdd.n1380 185
R874 vdd.n1424 vdd.n1381 185
R875 vdd.n1383 vdd.n1382 185
R876 vdd.n1420 vdd.n1385 185
R877 vdd.n1419 vdd.n1386 185
R878 vdd.n1418 vdd.n1387 185
R879 vdd.n1389 vdd.n1388 185
R880 vdd.n1414 vdd.n1391 185
R881 vdd.n1413 vdd.n1392 185
R882 vdd.n1412 vdd.n1393 185
R883 vdd.n1395 vdd.n1394 185
R884 vdd.n1408 vdd.n1397 185
R885 vdd.n1407 vdd.n1398 185
R886 vdd.n1406 vdd.n1399 185
R887 vdd.n1403 vdd.n1307 185
R888 vdd.n1501 vdd.n1307 185
R889 vdd.n1813 vdd.n1812 185
R890 vdd.n1817 vdd.n939 185
R891 vdd.n1693 vdd.n938 185
R892 vdd.n1696 vdd.n1695 185
R893 vdd.n1698 vdd.n1697 185
R894 vdd.n1701 vdd.n1700 185
R895 vdd.n1703 vdd.n1702 185
R896 vdd.n1705 vdd.n1691 185
R897 vdd.n1707 vdd.n1706 185
R898 vdd.n1708 vdd.n1685 185
R899 vdd.n1710 vdd.n1709 185
R900 vdd.n1712 vdd.n1683 185
R901 vdd.n1714 vdd.n1713 185
R902 vdd.n1715 vdd.n1678 185
R903 vdd.n1717 vdd.n1716 185
R904 vdd.n1719 vdd.n1676 185
R905 vdd.n1721 vdd.n1720 185
R906 vdd.n1722 vdd.n1672 185
R907 vdd.n1724 vdd.n1723 185
R908 vdd.n1726 vdd.n1669 185
R909 vdd.n1728 vdd.n1727 185
R910 vdd.n1670 vdd.n1663 185
R911 vdd.n1732 vdd.n1667 185
R912 vdd.n1733 vdd.n1659 185
R913 vdd.n1735 vdd.n1734 185
R914 vdd.n1737 vdd.n1657 185
R915 vdd.n1739 vdd.n1738 185
R916 vdd.n1740 vdd.n1652 185
R917 vdd.n1742 vdd.n1741 185
R918 vdd.n1744 vdd.n1650 185
R919 vdd.n1746 vdd.n1745 185
R920 vdd.n1747 vdd.n1645 185
R921 vdd.n1749 vdd.n1748 185
R922 vdd.n1751 vdd.n1643 185
R923 vdd.n1753 vdd.n1752 185
R924 vdd.n1754 vdd.n1638 185
R925 vdd.n1756 vdd.n1755 185
R926 vdd.n1758 vdd.n1636 185
R927 vdd.n1760 vdd.n1759 185
R928 vdd.n1761 vdd.n1632 185
R929 vdd.n1763 vdd.n1762 185
R930 vdd.n1765 vdd.n1629 185
R931 vdd.n1767 vdd.n1766 185
R932 vdd.n1630 vdd.n1623 185
R933 vdd.n1771 vdd.n1627 185
R934 vdd.n1772 vdd.n1619 185
R935 vdd.n1774 vdd.n1773 185
R936 vdd.n1776 vdd.n1617 185
R937 vdd.n1778 vdd.n1777 185
R938 vdd.n1779 vdd.n1612 185
R939 vdd.n1781 vdd.n1780 185
R940 vdd.n1783 vdd.n1610 185
R941 vdd.n1785 vdd.n1784 185
R942 vdd.n1786 vdd.n1605 185
R943 vdd.n1788 vdd.n1787 185
R944 vdd.n1790 vdd.n1604 185
R945 vdd.n1791 vdd.n1601 185
R946 vdd.n1794 vdd.n1793 185
R947 vdd.n1603 vdd.n1599 185
R948 vdd.n1798 vdd.n1597 185
R949 vdd.n1800 vdd.n1799 185
R950 vdd.n1802 vdd.n1595 185
R951 vdd.n1804 vdd.n1803 185
R952 vdd.n1805 vdd.n945 185
R953 vdd.n1811 vdd.n942 185
R954 vdd.n1811 vdd.n1810 185
R955 vdd.n953 vdd.n941 185
R956 vdd.n1588 vdd.n941 185
R957 vdd.n1587 vdd.n1586 185
R958 vdd.n1589 vdd.n1587 185
R959 vdd.n952 vdd.n951 185
R960 vdd.n951 vdd.n950 185
R961 vdd.n1580 vdd.n1579 185
R962 vdd.n1579 vdd.n1578 185
R963 vdd.n956 vdd.n955 185
R964 vdd.n1569 vdd.n956 185
R965 vdd.n1568 vdd.n1567 185
R966 vdd.n1570 vdd.n1568 185
R967 vdd.n963 vdd.n962 185
R968 vdd.n968 vdd.n962 185
R969 vdd.n1563 vdd.n1562 185
R970 vdd.n1562 vdd.n1561 185
R971 vdd.n966 vdd.n965 185
R972 vdd.n967 vdd.n966 185
R973 vdd.n1552 vdd.n1551 185
R974 vdd.n1553 vdd.n1552 185
R975 vdd.n1246 vdd.n1245 185
R976 vdd.n1245 vdd.n1244 185
R977 vdd.n1547 vdd.n1546 185
R978 vdd.n1546 vdd.n1545 185
R979 vdd.n1249 vdd.n1248 185
R980 vdd.n1535 vdd.n1249 185
R981 vdd.n1534 vdd.n1533 185
R982 vdd.n1536 vdd.n1534 185
R983 vdd.n1256 vdd.n1255 185
R984 vdd.n1260 vdd.n1255 185
R985 vdd.n1529 vdd.n1528 185
R986 vdd.n1528 vdd.n1527 185
R987 vdd.n1259 vdd.n1258 185
R988 vdd.n1518 vdd.n1259 185
R989 vdd.n1517 vdd.n1516 185
R990 vdd.n1519 vdd.n1517 185
R991 vdd.n1268 vdd.n1267 185
R992 vdd.n1267 vdd.n1266 185
R993 vdd.n1512 vdd.n1511 185
R994 vdd.n1511 vdd.n1510 185
R995 vdd.n1271 vdd.n1270 185
R996 vdd.n1308 vdd.n1271 185
R997 vdd.n777 vdd.n775 185
R998 vdd.n2268 vdd.n775 185
R999 vdd.n2190 vdd.n795 185
R1000 vdd.n795 vdd.n782 185
R1001 vdd.n2192 vdd.n2191 185
R1002 vdd.n2193 vdd.n2192 185
R1003 vdd.n2189 vdd.n794 185
R1004 vdd.n1948 vdd.n794 185
R1005 vdd.n2188 vdd.n2187 185
R1006 vdd.n2187 vdd.n2186 185
R1007 vdd.n797 vdd.n796 185
R1008 vdd.n798 vdd.n797 185
R1009 vdd.n2177 vdd.n2176 185
R1010 vdd.n2178 vdd.n2177 185
R1011 vdd.n2175 vdd.n808 185
R1012 vdd.n808 vdd.n805 185
R1013 vdd.n2174 vdd.n2173 185
R1014 vdd.n2173 vdd.n2172 185
R1015 vdd.n810 vdd.n809 185
R1016 vdd.n1960 vdd.n810 185
R1017 vdd.n2165 vdd.n2164 185
R1018 vdd.n2166 vdd.n2165 185
R1019 vdd.n2163 vdd.n818 185
R1020 vdd.n823 vdd.n818 185
R1021 vdd.n2162 vdd.n2161 185
R1022 vdd.n2161 vdd.n2160 185
R1023 vdd.n820 vdd.n819 185
R1024 vdd.n829 vdd.n820 185
R1025 vdd.n2153 vdd.n2152 185
R1026 vdd.n2154 vdd.n2153 185
R1027 vdd.n2151 vdd.n830 185
R1028 vdd.n1972 vdd.n830 185
R1029 vdd.n2150 vdd.n2149 185
R1030 vdd.n2149 vdd.n2148 185
R1031 vdd.n832 vdd.n831 185
R1032 vdd.n833 vdd.n832 185
R1033 vdd.n2141 vdd.n2140 185
R1034 vdd.n2142 vdd.n2141 185
R1035 vdd.n2139 vdd.n842 185
R1036 vdd.n842 vdd.n839 185
R1037 vdd.n2138 vdd.n2137 185
R1038 vdd.n2137 vdd.n2136 185
R1039 vdd.n844 vdd.n843 185
R1040 vdd.n853 vdd.n844 185
R1041 vdd.n2128 vdd.n2127 185
R1042 vdd.n2129 vdd.n2128 185
R1043 vdd.n2126 vdd.n854 185
R1044 vdd.n860 vdd.n854 185
R1045 vdd.n2125 vdd.n2124 185
R1046 vdd.n2124 vdd.n2123 185
R1047 vdd.n856 vdd.n855 185
R1048 vdd.n857 vdd.n856 185
R1049 vdd.n2116 vdd.n2115 185
R1050 vdd.n2117 vdd.n2116 185
R1051 vdd.n2114 vdd.n867 185
R1052 vdd.n867 vdd.n864 185
R1053 vdd.n2113 vdd.n2112 185
R1054 vdd.n2112 vdd.n2111 185
R1055 vdd.n869 vdd.n868 185
R1056 vdd.n870 vdd.n869 185
R1057 vdd.n2104 vdd.n2103 185
R1058 vdd.n2105 vdd.n2104 185
R1059 vdd.n2102 vdd.n879 185
R1060 vdd.n879 vdd.n876 185
R1061 vdd.n2101 vdd.n2100 185
R1062 vdd.n2100 vdd.n2099 185
R1063 vdd.n881 vdd.n880 185
R1064 vdd.n882 vdd.n881 185
R1065 vdd.n2092 vdd.n2091 185
R1066 vdd.n2093 vdd.n2092 185
R1067 vdd.n2090 vdd.n891 185
R1068 vdd.n891 vdd.n888 185
R1069 vdd.n2089 vdd.n2088 185
R1070 vdd.n2088 vdd.n2087 185
R1071 vdd.n893 vdd.n892 185
R1072 vdd.n894 vdd.n893 185
R1073 vdd.n2080 vdd.n2079 185
R1074 vdd.n2081 vdd.n2080 185
R1075 vdd.n2078 vdd.n903 185
R1076 vdd.n2077 vdd.n2076 185
R1077 vdd.n2074 vdd.n904 185
R1078 vdd.n2074 vdd.n900 185
R1079 vdd.n2073 vdd.n2072 185
R1080 vdd.n2071 vdd.n2070 185
R1081 vdd.n2069 vdd.n906 185
R1082 vdd.n2067 vdd.n2066 185
R1083 vdd.n2065 vdd.n907 185
R1084 vdd.n2064 vdd.n2063 185
R1085 vdd.n2061 vdd.n908 185
R1086 vdd.n2059 vdd.n2058 185
R1087 vdd.n2057 vdd.n909 185
R1088 vdd.n2056 vdd.n2055 185
R1089 vdd.n2053 vdd.n910 185
R1090 vdd.n2051 vdd.n2050 185
R1091 vdd.n2049 vdd.n911 185
R1092 vdd.n2048 vdd.n2047 185
R1093 vdd.n2045 vdd.n912 185
R1094 vdd.n2043 vdd.n2042 185
R1095 vdd.n2041 vdd.n913 185
R1096 vdd.n2040 vdd.n2039 185
R1097 vdd.n2037 vdd.n914 185
R1098 vdd.n2035 vdd.n2034 185
R1099 vdd.n2033 vdd.n915 185
R1100 vdd.n2032 vdd.n2031 185
R1101 vdd.n2029 vdd.n916 185
R1102 vdd.n2027 vdd.n2026 185
R1103 vdd.n2025 vdd.n917 185
R1104 vdd.n2024 vdd.n2023 185
R1105 vdd.n2021 vdd.n918 185
R1106 vdd.n2019 vdd.n2018 185
R1107 vdd.n2017 vdd.n919 185
R1108 vdd.n2015 vdd.n2014 185
R1109 vdd.n2012 vdd.n922 185
R1110 vdd.n2010 vdd.n2009 185
R1111 vdd.n2271 vdd.n2270 185
R1112 vdd.n2273 vdd.n2272 185
R1113 vdd.n2275 vdd.n2274 185
R1114 vdd.n2278 vdd.n2277 185
R1115 vdd.n2280 vdd.n2279 185
R1116 vdd.n2282 vdd.n2281 185
R1117 vdd.n2284 vdd.n2283 185
R1118 vdd.n2286 vdd.n2285 185
R1119 vdd.n2288 vdd.n2287 185
R1120 vdd.n2290 vdd.n2289 185
R1121 vdd.n2292 vdd.n2291 185
R1122 vdd.n2294 vdd.n2293 185
R1123 vdd.n2296 vdd.n2295 185
R1124 vdd.n2298 vdd.n2297 185
R1125 vdd.n2300 vdd.n2299 185
R1126 vdd.n2302 vdd.n2301 185
R1127 vdd.n2304 vdd.n2303 185
R1128 vdd.n2306 vdd.n2305 185
R1129 vdd.n2308 vdd.n2307 185
R1130 vdd.n2310 vdd.n2309 185
R1131 vdd.n2312 vdd.n2311 185
R1132 vdd.n2314 vdd.n2313 185
R1133 vdd.n2316 vdd.n2315 185
R1134 vdd.n2318 vdd.n2317 185
R1135 vdd.n2320 vdd.n2319 185
R1136 vdd.n2322 vdd.n2321 185
R1137 vdd.n2324 vdd.n2323 185
R1138 vdd.n2326 vdd.n2325 185
R1139 vdd.n2328 vdd.n2327 185
R1140 vdd.n2330 vdd.n2329 185
R1141 vdd.n2332 vdd.n2331 185
R1142 vdd.n2334 vdd.n2333 185
R1143 vdd.n2336 vdd.n2335 185
R1144 vdd.n2337 vdd.n776 185
R1145 vdd.n2339 vdd.n2338 185
R1146 vdd.n2340 vdd.n2339 185
R1147 vdd.n2269 vdd.n780 185
R1148 vdd.n2269 vdd.n2268 185
R1149 vdd.n1946 vdd.n781 185
R1150 vdd.n782 vdd.n781 185
R1151 vdd.n1947 vdd.n792 185
R1152 vdd.n2193 vdd.n792 185
R1153 vdd.n1950 vdd.n1949 185
R1154 vdd.n1949 vdd.n1948 185
R1155 vdd.n1951 vdd.n799 185
R1156 vdd.n2186 vdd.n799 185
R1157 vdd.n1953 vdd.n1952 185
R1158 vdd.n1952 vdd.n798 185
R1159 vdd.n1954 vdd.n806 185
R1160 vdd.n2178 vdd.n806 185
R1161 vdd.n1956 vdd.n1955 185
R1162 vdd.n1955 vdd.n805 185
R1163 vdd.n1957 vdd.n811 185
R1164 vdd.n2172 vdd.n811 185
R1165 vdd.n1959 vdd.n1958 185
R1166 vdd.n1960 vdd.n1959 185
R1167 vdd.n1945 vdd.n816 185
R1168 vdd.n2166 vdd.n816 185
R1169 vdd.n1944 vdd.n1943 185
R1170 vdd.n1943 vdd.n823 185
R1171 vdd.n1942 vdd.n821 185
R1172 vdd.n2160 vdd.n821 185
R1173 vdd.n1941 vdd.n1940 185
R1174 vdd.n1940 vdd.n829 185
R1175 vdd.n923 vdd.n827 185
R1176 vdd.n2154 vdd.n827 185
R1177 vdd.n1974 vdd.n1973 185
R1178 vdd.n1973 vdd.n1972 185
R1179 vdd.n1975 vdd.n834 185
R1180 vdd.n2148 vdd.n834 185
R1181 vdd.n1977 vdd.n1976 185
R1182 vdd.n1976 vdd.n833 185
R1183 vdd.n1978 vdd.n840 185
R1184 vdd.n2142 vdd.n840 185
R1185 vdd.n1980 vdd.n1979 185
R1186 vdd.n1979 vdd.n839 185
R1187 vdd.n1981 vdd.n845 185
R1188 vdd.n2136 vdd.n845 185
R1189 vdd.n1983 vdd.n1982 185
R1190 vdd.n1982 vdd.n853 185
R1191 vdd.n1984 vdd.n851 185
R1192 vdd.n2129 vdd.n851 185
R1193 vdd.n1986 vdd.n1985 185
R1194 vdd.n1985 vdd.n860 185
R1195 vdd.n1987 vdd.n858 185
R1196 vdd.n2123 vdd.n858 185
R1197 vdd.n1989 vdd.n1988 185
R1198 vdd.n1988 vdd.n857 185
R1199 vdd.n1990 vdd.n865 185
R1200 vdd.n2117 vdd.n865 185
R1201 vdd.n1992 vdd.n1991 185
R1202 vdd.n1991 vdd.n864 185
R1203 vdd.n1993 vdd.n871 185
R1204 vdd.n2111 vdd.n871 185
R1205 vdd.n1995 vdd.n1994 185
R1206 vdd.n1994 vdd.n870 185
R1207 vdd.n1996 vdd.n877 185
R1208 vdd.n2105 vdd.n877 185
R1209 vdd.n1998 vdd.n1997 185
R1210 vdd.n1997 vdd.n876 185
R1211 vdd.n1999 vdd.n883 185
R1212 vdd.n2099 vdd.n883 185
R1213 vdd.n2001 vdd.n2000 185
R1214 vdd.n2000 vdd.n882 185
R1215 vdd.n2002 vdd.n889 185
R1216 vdd.n2093 vdd.n889 185
R1217 vdd.n2004 vdd.n2003 185
R1218 vdd.n2003 vdd.n888 185
R1219 vdd.n2005 vdd.n895 185
R1220 vdd.n2087 vdd.n895 185
R1221 vdd.n2007 vdd.n2006 185
R1222 vdd.n2006 vdd.n894 185
R1223 vdd.n2008 vdd.n901 185
R1224 vdd.n2081 vdd.n901 185
R1225 vdd.n3206 vdd.n3205 185
R1226 vdd.n3207 vdd.n3206 185
R1227 vdd.n325 vdd.n324 185
R1228 vdd.n3208 vdd.n325 185
R1229 vdd.n3211 vdd.n3210 185
R1230 vdd.n3210 vdd.n3209 185
R1231 vdd.n3212 vdd.n319 185
R1232 vdd.n319 vdd.n318 185
R1233 vdd.n3214 vdd.n3213 185
R1234 vdd.n3215 vdd.n3214 185
R1235 vdd.n314 vdd.n313 185
R1236 vdd.n3216 vdd.n314 185
R1237 vdd.n3219 vdd.n3218 185
R1238 vdd.n3218 vdd.n3217 185
R1239 vdd.n3220 vdd.n309 185
R1240 vdd.n309 vdd.n308 185
R1241 vdd.n3222 vdd.n3221 185
R1242 vdd.n3223 vdd.n3222 185
R1243 vdd.n303 vdd.n301 185
R1244 vdd.n3224 vdd.n303 185
R1245 vdd.n3227 vdd.n3226 185
R1246 vdd.n3226 vdd.n3225 185
R1247 vdd.n302 vdd.n300 185
R1248 vdd.n304 vdd.n302 185
R1249 vdd.n3063 vdd.n3062 185
R1250 vdd.n3064 vdd.n3063 185
R1251 vdd.n458 vdd.n457 185
R1252 vdd.n457 vdd.n456 185
R1253 vdd.n3058 vdd.n3057 185
R1254 vdd.n3057 vdd.n3056 185
R1255 vdd.n461 vdd.n460 185
R1256 vdd.n467 vdd.n461 185
R1257 vdd.n3047 vdd.n3046 185
R1258 vdd.n3048 vdd.n3047 185
R1259 vdd.n469 vdd.n468 185
R1260 vdd.n3039 vdd.n468 185
R1261 vdd.n3042 vdd.n3041 185
R1262 vdd.n3041 vdd.n3040 185
R1263 vdd.n472 vdd.n471 185
R1264 vdd.n473 vdd.n472 185
R1265 vdd.n3030 vdd.n3029 185
R1266 vdd.n3031 vdd.n3030 185
R1267 vdd.n480 vdd.n479 185
R1268 vdd.n516 vdd.n479 185
R1269 vdd.n3025 vdd.n3024 185
R1270 vdd.n483 vdd.n482 185
R1271 vdd.n3021 vdd.n3020 185
R1272 vdd.n3022 vdd.n3021 185
R1273 vdd.n518 vdd.n517 185
R1274 vdd.n522 vdd.n521 185
R1275 vdd.n3016 vdd.n523 185
R1276 vdd.n3015 vdd.n3014 185
R1277 vdd.n3013 vdd.n3012 185
R1278 vdd.n3011 vdd.n3010 185
R1279 vdd.n3009 vdd.n3008 185
R1280 vdd.n3007 vdd.n3006 185
R1281 vdd.n3005 vdd.n3004 185
R1282 vdd.n3003 vdd.n3002 185
R1283 vdd.n3001 vdd.n3000 185
R1284 vdd.n2999 vdd.n2998 185
R1285 vdd.n2997 vdd.n2996 185
R1286 vdd.n2995 vdd.n2994 185
R1287 vdd.n2993 vdd.n2992 185
R1288 vdd.n2991 vdd.n2990 185
R1289 vdd.n2989 vdd.n2988 185
R1290 vdd.n2980 vdd.n536 185
R1291 vdd.n2982 vdd.n2981 185
R1292 vdd.n2979 vdd.n2978 185
R1293 vdd.n2977 vdd.n2976 185
R1294 vdd.n2975 vdd.n2974 185
R1295 vdd.n2973 vdd.n2972 185
R1296 vdd.n2971 vdd.n2970 185
R1297 vdd.n2969 vdd.n2968 185
R1298 vdd.n2967 vdd.n2966 185
R1299 vdd.n2965 vdd.n2964 185
R1300 vdd.n2963 vdd.n2962 185
R1301 vdd.n2961 vdd.n2960 185
R1302 vdd.n2959 vdd.n2958 185
R1303 vdd.n2957 vdd.n2956 185
R1304 vdd.n2955 vdd.n2954 185
R1305 vdd.n2953 vdd.n2952 185
R1306 vdd.n2951 vdd.n2950 185
R1307 vdd.n2949 vdd.n2948 185
R1308 vdd.n2947 vdd.n2946 185
R1309 vdd.n2945 vdd.n2944 185
R1310 vdd.n2943 vdd.n2942 185
R1311 vdd.n2941 vdd.n2940 185
R1312 vdd.n2934 vdd.n556 185
R1313 vdd.n2936 vdd.n2935 185
R1314 vdd.n2933 vdd.n2932 185
R1315 vdd.n2931 vdd.n2930 185
R1316 vdd.n2929 vdd.n2928 185
R1317 vdd.n2927 vdd.n2926 185
R1318 vdd.n2925 vdd.n2924 185
R1319 vdd.n2923 vdd.n2922 185
R1320 vdd.n2921 vdd.n2920 185
R1321 vdd.n2919 vdd.n2918 185
R1322 vdd.n2917 vdd.n2916 185
R1323 vdd.n2915 vdd.n2914 185
R1324 vdd.n2913 vdd.n2912 185
R1325 vdd.n2911 vdd.n2910 185
R1326 vdd.n2909 vdd.n2908 185
R1327 vdd.n2907 vdd.n2906 185
R1328 vdd.n2905 vdd.n2904 185
R1329 vdd.n2903 vdd.n2902 185
R1330 vdd.n2901 vdd.n2900 185
R1331 vdd.n2899 vdd.n2898 185
R1332 vdd.n2897 vdd.n2896 185
R1333 vdd.n2892 vdd.n515 185
R1334 vdd.n3022 vdd.n515 185
R1335 vdd.n3089 vdd.n3088 185
R1336 vdd.n3093 vdd.n440 185
R1337 vdd.n3095 vdd.n3094 185
R1338 vdd.n3097 vdd.n438 185
R1339 vdd.n3099 vdd.n3098 185
R1340 vdd.n3100 vdd.n433 185
R1341 vdd.n3102 vdd.n3101 185
R1342 vdd.n3104 vdd.n431 185
R1343 vdd.n3106 vdd.n3105 185
R1344 vdd.n3107 vdd.n426 185
R1345 vdd.n3109 vdd.n3108 185
R1346 vdd.n3111 vdd.n424 185
R1347 vdd.n3113 vdd.n3112 185
R1348 vdd.n3114 vdd.n419 185
R1349 vdd.n3116 vdd.n3115 185
R1350 vdd.n3118 vdd.n417 185
R1351 vdd.n3120 vdd.n3119 185
R1352 vdd.n3121 vdd.n413 185
R1353 vdd.n3123 vdd.n3122 185
R1354 vdd.n3125 vdd.n410 185
R1355 vdd.n3127 vdd.n3126 185
R1356 vdd.n411 vdd.n404 185
R1357 vdd.n3131 vdd.n408 185
R1358 vdd.n3132 vdd.n400 185
R1359 vdd.n3134 vdd.n3133 185
R1360 vdd.n3136 vdd.n398 185
R1361 vdd.n3138 vdd.n3137 185
R1362 vdd.n3139 vdd.n393 185
R1363 vdd.n3141 vdd.n3140 185
R1364 vdd.n3143 vdd.n391 185
R1365 vdd.n3145 vdd.n3144 185
R1366 vdd.n3146 vdd.n386 185
R1367 vdd.n3148 vdd.n3147 185
R1368 vdd.n3150 vdd.n384 185
R1369 vdd.n3152 vdd.n3151 185
R1370 vdd.n3153 vdd.n379 185
R1371 vdd.n3155 vdd.n3154 185
R1372 vdd.n3157 vdd.n377 185
R1373 vdd.n3159 vdd.n3158 185
R1374 vdd.n3160 vdd.n373 185
R1375 vdd.n3162 vdd.n3161 185
R1376 vdd.n3164 vdd.n370 185
R1377 vdd.n3166 vdd.n3165 185
R1378 vdd.n371 vdd.n364 185
R1379 vdd.n3170 vdd.n368 185
R1380 vdd.n3171 vdd.n360 185
R1381 vdd.n3173 vdd.n3172 185
R1382 vdd.n3175 vdd.n358 185
R1383 vdd.n3177 vdd.n3176 185
R1384 vdd.n3178 vdd.n353 185
R1385 vdd.n3180 vdd.n3179 185
R1386 vdd.n3182 vdd.n351 185
R1387 vdd.n3184 vdd.n3183 185
R1388 vdd.n3185 vdd.n346 185
R1389 vdd.n3187 vdd.n3186 185
R1390 vdd.n3189 vdd.n344 185
R1391 vdd.n3191 vdd.n3190 185
R1392 vdd.n3192 vdd.n338 185
R1393 vdd.n3194 vdd.n3193 185
R1394 vdd.n3196 vdd.n337 185
R1395 vdd.n3197 vdd.n336 185
R1396 vdd.n3200 vdd.n3199 185
R1397 vdd.n3201 vdd.n334 185
R1398 vdd.n3202 vdd.n330 185
R1399 vdd.n3084 vdd.n328 185
R1400 vdd.n3207 vdd.n328 185
R1401 vdd.n3083 vdd.n327 185
R1402 vdd.n3208 vdd.n327 185
R1403 vdd.n3082 vdd.n326 185
R1404 vdd.n3209 vdd.n326 185
R1405 vdd.n446 vdd.n445 185
R1406 vdd.n445 vdd.n318 185
R1407 vdd.n3078 vdd.n317 185
R1408 vdd.n3215 vdd.n317 185
R1409 vdd.n3077 vdd.n316 185
R1410 vdd.n3216 vdd.n316 185
R1411 vdd.n3076 vdd.n315 185
R1412 vdd.n3217 vdd.n315 185
R1413 vdd.n449 vdd.n448 185
R1414 vdd.n448 vdd.n308 185
R1415 vdd.n3072 vdd.n307 185
R1416 vdd.n3223 vdd.n307 185
R1417 vdd.n3071 vdd.n306 185
R1418 vdd.n3224 vdd.n306 185
R1419 vdd.n3070 vdd.n305 185
R1420 vdd.n3225 vdd.n305 185
R1421 vdd.n455 vdd.n451 185
R1422 vdd.n455 vdd.n304 185
R1423 vdd.n3066 vdd.n3065 185
R1424 vdd.n3065 vdd.n3064 185
R1425 vdd.n454 vdd.n453 185
R1426 vdd.n456 vdd.n454 185
R1427 vdd.n3055 vdd.n3054 185
R1428 vdd.n3056 vdd.n3055 185
R1429 vdd.n463 vdd.n462 185
R1430 vdd.n467 vdd.n462 185
R1431 vdd.n3050 vdd.n3049 185
R1432 vdd.n3049 vdd.n3048 185
R1433 vdd.n466 vdd.n465 185
R1434 vdd.n3039 vdd.n466 185
R1435 vdd.n3038 vdd.n3037 185
R1436 vdd.n3040 vdd.n3038 185
R1437 vdd.n475 vdd.n474 185
R1438 vdd.n474 vdd.n473 185
R1439 vdd.n3033 vdd.n3032 185
R1440 vdd.n3032 vdd.n3031 185
R1441 vdd.n478 vdd.n477 185
R1442 vdd.n516 vdd.n478 185
R1443 vdd.n2628 vdd.n737 185
R1444 vdd.n2627 vdd.n2626 185
R1445 vdd.n739 vdd.n738 185
R1446 vdd.n2624 vdd.n739 185
R1447 vdd.n2447 vdd.n2446 185
R1448 vdd.n2449 vdd.n2448 185
R1449 vdd.n2451 vdd.n2450 185
R1450 vdd.n2453 vdd.n2452 185
R1451 vdd.n2455 vdd.n2454 185
R1452 vdd.n2457 vdd.n2456 185
R1453 vdd.n2459 vdd.n2458 185
R1454 vdd.n2461 vdd.n2460 185
R1455 vdd.n2463 vdd.n2462 185
R1456 vdd.n2465 vdd.n2464 185
R1457 vdd.n2467 vdd.n2466 185
R1458 vdd.n2469 vdd.n2468 185
R1459 vdd.n2471 vdd.n2470 185
R1460 vdd.n2473 vdd.n2472 185
R1461 vdd.n2475 vdd.n2474 185
R1462 vdd.n2477 vdd.n2476 185
R1463 vdd.n2479 vdd.n2478 185
R1464 vdd.n2481 vdd.n2480 185
R1465 vdd.n2483 vdd.n2482 185
R1466 vdd.n2485 vdd.n2484 185
R1467 vdd.n2487 vdd.n2486 185
R1468 vdd.n2489 vdd.n2488 185
R1469 vdd.n2491 vdd.n2490 185
R1470 vdd.n2493 vdd.n2492 185
R1471 vdd.n2495 vdd.n2494 185
R1472 vdd.n2497 vdd.n2496 185
R1473 vdd.n2499 vdd.n2498 185
R1474 vdd.n2501 vdd.n2500 185
R1475 vdd.n2503 vdd.n2502 185
R1476 vdd.n2506 vdd.n2505 185
R1477 vdd.n2508 vdd.n2507 185
R1478 vdd.n2510 vdd.n2509 185
R1479 vdd.n2791 vdd.n2790 185
R1480 vdd.n2793 vdd.n624 185
R1481 vdd.n2795 vdd.n2794 185
R1482 vdd.n2797 vdd.n621 185
R1483 vdd.n2799 vdd.n2798 185
R1484 vdd.n2801 vdd.n619 185
R1485 vdd.n2803 vdd.n2802 185
R1486 vdd.n2804 vdd.n618 185
R1487 vdd.n2806 vdd.n2805 185
R1488 vdd.n2808 vdd.n616 185
R1489 vdd.n2810 vdd.n2809 185
R1490 vdd.n2811 vdd.n615 185
R1491 vdd.n2813 vdd.n2812 185
R1492 vdd.n2815 vdd.n613 185
R1493 vdd.n2817 vdd.n2816 185
R1494 vdd.n2818 vdd.n612 185
R1495 vdd.n2820 vdd.n2819 185
R1496 vdd.n2822 vdd.n520 185
R1497 vdd.n2824 vdd.n2823 185
R1498 vdd.n2826 vdd.n610 185
R1499 vdd.n2828 vdd.n2827 185
R1500 vdd.n2829 vdd.n609 185
R1501 vdd.n2831 vdd.n2830 185
R1502 vdd.n2833 vdd.n607 185
R1503 vdd.n2835 vdd.n2834 185
R1504 vdd.n2836 vdd.n606 185
R1505 vdd.n2838 vdd.n2837 185
R1506 vdd.n2840 vdd.n604 185
R1507 vdd.n2842 vdd.n2841 185
R1508 vdd.n2843 vdd.n603 185
R1509 vdd.n2845 vdd.n2844 185
R1510 vdd.n2847 vdd.n602 185
R1511 vdd.n2848 vdd.n601 185
R1512 vdd.n2851 vdd.n2850 185
R1513 vdd.n2852 vdd.n599 185
R1514 vdd.n599 vdd.n484 185
R1515 vdd.n2789 vdd.n596 185
R1516 vdd.n2855 vdd.n596 185
R1517 vdd.n2788 vdd.n2787 185
R1518 vdd.n2787 vdd.n595 185
R1519 vdd.n2786 vdd.n626 185
R1520 vdd.n2786 vdd.n2785 185
R1521 vdd.n2560 vdd.n627 185
R1522 vdd.n636 vdd.n627 185
R1523 vdd.n2561 vdd.n634 185
R1524 vdd.n2779 vdd.n634 185
R1525 vdd.n2563 vdd.n2562 185
R1526 vdd.n2562 vdd.n633 185
R1527 vdd.n2564 vdd.n642 185
R1528 vdd.n2728 vdd.n642 185
R1529 vdd.n2566 vdd.n2565 185
R1530 vdd.n2565 vdd.n641 185
R1531 vdd.n2567 vdd.n647 185
R1532 vdd.n2722 vdd.n647 185
R1533 vdd.n2569 vdd.n2568 185
R1534 vdd.n2568 vdd.n654 185
R1535 vdd.n2570 vdd.n652 185
R1536 vdd.n2716 vdd.n652 185
R1537 vdd.n2572 vdd.n2571 185
R1538 vdd.n2571 vdd.n660 185
R1539 vdd.n2573 vdd.n658 185
R1540 vdd.n2710 vdd.n658 185
R1541 vdd.n2575 vdd.n2574 185
R1542 vdd.n2574 vdd.n667 185
R1543 vdd.n2576 vdd.n665 185
R1544 vdd.n2704 vdd.n665 185
R1545 vdd.n2578 vdd.n2577 185
R1546 vdd.n2577 vdd.n664 185
R1547 vdd.n2579 vdd.n672 185
R1548 vdd.n2698 vdd.n672 185
R1549 vdd.n2581 vdd.n2580 185
R1550 vdd.n2580 vdd.n671 185
R1551 vdd.n2582 vdd.n679 185
R1552 vdd.n2691 vdd.n679 185
R1553 vdd.n2584 vdd.n2583 185
R1554 vdd.n2583 vdd.n678 185
R1555 vdd.n2585 vdd.n684 185
R1556 vdd.n2685 vdd.n684 185
R1557 vdd.n2587 vdd.n2586 185
R1558 vdd.n2586 vdd.n691 185
R1559 vdd.n2588 vdd.n689 185
R1560 vdd.n2679 vdd.n689 185
R1561 vdd.n2590 vdd.n2589 185
R1562 vdd.n2591 vdd.n2590 185
R1563 vdd.n2559 vdd.n696 185
R1564 vdd.n2673 vdd.n696 185
R1565 vdd.n2558 vdd.n2557 185
R1566 vdd.n2557 vdd.n695 185
R1567 vdd.n2556 vdd.n702 185
R1568 vdd.n2667 vdd.n702 185
R1569 vdd.n2555 vdd.n2554 185
R1570 vdd.n2554 vdd.n701 185
R1571 vdd.n2515 vdd.n707 185
R1572 vdd.n2661 vdd.n707 185
R1573 vdd.n2605 vdd.n2604 185
R1574 vdd.n2604 vdd.n2603 185
R1575 vdd.n2606 vdd.n712 185
R1576 vdd.n2655 vdd.n712 185
R1577 vdd.n2608 vdd.n2607 185
R1578 vdd.n2607 vdd.n720 185
R1579 vdd.n2609 vdd.n718 185
R1580 vdd.n2649 vdd.n718 185
R1581 vdd.n2611 vdd.n2610 185
R1582 vdd.n2610 vdd.n717 185
R1583 vdd.n2612 vdd.n724 185
R1584 vdd.n2643 vdd.n724 185
R1585 vdd.n2614 vdd.n2613 185
R1586 vdd.n2615 vdd.n2614 185
R1587 vdd.n2514 vdd.n729 185
R1588 vdd.n2637 vdd.n729 185
R1589 vdd.n2513 vdd.n2512 185
R1590 vdd.n2512 vdd.n736 185
R1591 vdd.n2511 vdd.n734 185
R1592 vdd.n2631 vdd.n734 185
R1593 vdd.n2630 vdd.n2629 185
R1594 vdd.n2631 vdd.n2630 185
R1595 vdd.n728 vdd.n727 185
R1596 vdd.n736 vdd.n728 185
R1597 vdd.n2639 vdd.n2638 185
R1598 vdd.n2638 vdd.n2637 185
R1599 vdd.n2640 vdd.n726 185
R1600 vdd.n2615 vdd.n726 185
R1601 vdd.n2642 vdd.n2641 185
R1602 vdd.n2643 vdd.n2642 185
R1603 vdd.n716 vdd.n715 185
R1604 vdd.n717 vdd.n716 185
R1605 vdd.n2651 vdd.n2650 185
R1606 vdd.n2650 vdd.n2649 185
R1607 vdd.n2652 vdd.n714 185
R1608 vdd.n720 vdd.n714 185
R1609 vdd.n2654 vdd.n2653 185
R1610 vdd.n2655 vdd.n2654 185
R1611 vdd.n706 vdd.n705 185
R1612 vdd.n2603 vdd.n706 185
R1613 vdd.n2663 vdd.n2662 185
R1614 vdd.n2662 vdd.n2661 185
R1615 vdd.n2664 vdd.n704 185
R1616 vdd.n704 vdd.n701 185
R1617 vdd.n2666 vdd.n2665 185
R1618 vdd.n2667 vdd.n2666 185
R1619 vdd.n694 vdd.n693 185
R1620 vdd.n695 vdd.n694 185
R1621 vdd.n2675 vdd.n2674 185
R1622 vdd.n2674 vdd.n2673 185
R1623 vdd.n2676 vdd.n692 185
R1624 vdd.n2591 vdd.n692 185
R1625 vdd.n2678 vdd.n2677 185
R1626 vdd.n2679 vdd.n2678 185
R1627 vdd.n683 vdd.n682 185
R1628 vdd.n691 vdd.n683 185
R1629 vdd.n2687 vdd.n2686 185
R1630 vdd.n2686 vdd.n2685 185
R1631 vdd.n2688 vdd.n681 185
R1632 vdd.n681 vdd.n678 185
R1633 vdd.n2690 vdd.n2689 185
R1634 vdd.n2691 vdd.n2690 185
R1635 vdd.n670 vdd.n669 185
R1636 vdd.n671 vdd.n670 185
R1637 vdd.n2700 vdd.n2699 185
R1638 vdd.n2699 vdd.n2698 185
R1639 vdd.n2701 vdd.n668 185
R1640 vdd.n668 vdd.n664 185
R1641 vdd.n2703 vdd.n2702 185
R1642 vdd.n2704 vdd.n2703 185
R1643 vdd.n657 vdd.n656 185
R1644 vdd.n667 vdd.n657 185
R1645 vdd.n2712 vdd.n2711 185
R1646 vdd.n2711 vdd.n2710 185
R1647 vdd.n2713 vdd.n655 185
R1648 vdd.n660 vdd.n655 185
R1649 vdd.n2715 vdd.n2714 185
R1650 vdd.n2716 vdd.n2715 185
R1651 vdd.n646 vdd.n645 185
R1652 vdd.n654 vdd.n646 185
R1653 vdd.n2724 vdd.n2723 185
R1654 vdd.n2723 vdd.n2722 185
R1655 vdd.n2725 vdd.n644 185
R1656 vdd.n644 vdd.n641 185
R1657 vdd.n2727 vdd.n2726 185
R1658 vdd.n2728 vdd.n2727 185
R1659 vdd.n632 vdd.n631 185
R1660 vdd.n633 vdd.n632 185
R1661 vdd.n2781 vdd.n2780 185
R1662 vdd.n2780 vdd.n2779 185
R1663 vdd.n2782 vdd.n630 185
R1664 vdd.n636 vdd.n630 185
R1665 vdd.n2784 vdd.n2783 185
R1666 vdd.n2785 vdd.n2784 185
R1667 vdd.n600 vdd.n598 185
R1668 vdd.n598 vdd.n595 185
R1669 vdd.n2854 vdd.n2853 185
R1670 vdd.n2855 vdd.n2854 185
R1671 vdd.n2267 vdd.n2266 185
R1672 vdd.n2268 vdd.n2267 185
R1673 vdd.n786 vdd.n784 185
R1674 vdd.n784 vdd.n782 185
R1675 vdd.n2182 vdd.n793 185
R1676 vdd.n2193 vdd.n793 185
R1677 vdd.n2183 vdd.n802 185
R1678 vdd.n1948 vdd.n802 185
R1679 vdd.n2185 vdd.n2184 185
R1680 vdd.n2186 vdd.n2185 185
R1681 vdd.n2181 vdd.n801 185
R1682 vdd.n801 vdd.n798 185
R1683 vdd.n2180 vdd.n2179 185
R1684 vdd.n2179 vdd.n2178 185
R1685 vdd.n804 vdd.n803 185
R1686 vdd.n805 vdd.n804 185
R1687 vdd.n2171 vdd.n2170 185
R1688 vdd.n2172 vdd.n2171 185
R1689 vdd.n2169 vdd.n813 185
R1690 vdd.n1960 vdd.n813 185
R1691 vdd.n2168 vdd.n2167 185
R1692 vdd.n2167 vdd.n2166 185
R1693 vdd.n815 vdd.n814 185
R1694 vdd.n823 vdd.n815 185
R1695 vdd.n2159 vdd.n2158 185
R1696 vdd.n2160 vdd.n2159 185
R1697 vdd.n2157 vdd.n824 185
R1698 vdd.n829 vdd.n824 185
R1699 vdd.n2156 vdd.n2155 185
R1700 vdd.n2155 vdd.n2154 185
R1701 vdd.n826 vdd.n825 185
R1702 vdd.n1972 vdd.n826 185
R1703 vdd.n2147 vdd.n2146 185
R1704 vdd.n2148 vdd.n2147 185
R1705 vdd.n2145 vdd.n836 185
R1706 vdd.n836 vdd.n833 185
R1707 vdd.n2144 vdd.n2143 185
R1708 vdd.n2143 vdd.n2142 185
R1709 vdd.n838 vdd.n837 185
R1710 vdd.n839 vdd.n838 185
R1711 vdd.n2135 vdd.n2134 185
R1712 vdd.n2136 vdd.n2135 185
R1713 vdd.n2132 vdd.n847 185
R1714 vdd.n853 vdd.n847 185
R1715 vdd.n2131 vdd.n2130 185
R1716 vdd.n2130 vdd.n2129 185
R1717 vdd.n850 vdd.n849 185
R1718 vdd.n860 vdd.n850 185
R1719 vdd.n2122 vdd.n2121 185
R1720 vdd.n2123 vdd.n2122 185
R1721 vdd.n2120 vdd.n861 185
R1722 vdd.n861 vdd.n857 185
R1723 vdd.n2119 vdd.n2118 185
R1724 vdd.n2118 vdd.n2117 185
R1725 vdd.n863 vdd.n862 185
R1726 vdd.n864 vdd.n863 185
R1727 vdd.n2110 vdd.n2109 185
R1728 vdd.n2111 vdd.n2110 185
R1729 vdd.n2108 vdd.n873 185
R1730 vdd.n873 vdd.n870 185
R1731 vdd.n2107 vdd.n2106 185
R1732 vdd.n2106 vdd.n2105 185
R1733 vdd.n875 vdd.n874 185
R1734 vdd.n876 vdd.n875 185
R1735 vdd.n2098 vdd.n2097 185
R1736 vdd.n2099 vdd.n2098 185
R1737 vdd.n2096 vdd.n885 185
R1738 vdd.n885 vdd.n882 185
R1739 vdd.n2095 vdd.n2094 185
R1740 vdd.n2094 vdd.n2093 185
R1741 vdd.n887 vdd.n886 185
R1742 vdd.n888 vdd.n887 185
R1743 vdd.n2086 vdd.n2085 185
R1744 vdd.n2087 vdd.n2086 185
R1745 vdd.n2084 vdd.n897 185
R1746 vdd.n897 vdd.n894 185
R1747 vdd.n2083 vdd.n2082 185
R1748 vdd.n2082 vdd.n2081 185
R1749 vdd.n2198 vdd.n757 185
R1750 vdd.n2340 vdd.n757 185
R1751 vdd.n2200 vdd.n2199 185
R1752 vdd.n2202 vdd.n2201 185
R1753 vdd.n2204 vdd.n2203 185
R1754 vdd.n2206 vdd.n2205 185
R1755 vdd.n2208 vdd.n2207 185
R1756 vdd.n2210 vdd.n2209 185
R1757 vdd.n2212 vdd.n2211 185
R1758 vdd.n2214 vdd.n2213 185
R1759 vdd.n2216 vdd.n2215 185
R1760 vdd.n2218 vdd.n2217 185
R1761 vdd.n2220 vdd.n2219 185
R1762 vdd.n2222 vdd.n2221 185
R1763 vdd.n2224 vdd.n2223 185
R1764 vdd.n2226 vdd.n2225 185
R1765 vdd.n2228 vdd.n2227 185
R1766 vdd.n2230 vdd.n2229 185
R1767 vdd.n2232 vdd.n2231 185
R1768 vdd.n2234 vdd.n2233 185
R1769 vdd.n2236 vdd.n2235 185
R1770 vdd.n2238 vdd.n2237 185
R1771 vdd.n2240 vdd.n2239 185
R1772 vdd.n2242 vdd.n2241 185
R1773 vdd.n2244 vdd.n2243 185
R1774 vdd.n2246 vdd.n2245 185
R1775 vdd.n2248 vdd.n2247 185
R1776 vdd.n2250 vdd.n2249 185
R1777 vdd.n2252 vdd.n2251 185
R1778 vdd.n2254 vdd.n2253 185
R1779 vdd.n2256 vdd.n2255 185
R1780 vdd.n2258 vdd.n2257 185
R1781 vdd.n2260 vdd.n2259 185
R1782 vdd.n2262 vdd.n2261 185
R1783 vdd.n2264 vdd.n2263 185
R1784 vdd.n2265 vdd.n785 185
R1785 vdd.n2197 vdd.n783 185
R1786 vdd.n2268 vdd.n783 185
R1787 vdd.n2196 vdd.n2195 185
R1788 vdd.n2195 vdd.n782 185
R1789 vdd.n2194 vdd.n790 185
R1790 vdd.n2194 vdd.n2193 185
R1791 vdd.n1932 vdd.n791 185
R1792 vdd.n1948 vdd.n791 185
R1793 vdd.n1933 vdd.n800 185
R1794 vdd.n2186 vdd.n800 185
R1795 vdd.n1935 vdd.n1934 185
R1796 vdd.n1934 vdd.n798 185
R1797 vdd.n1936 vdd.n807 185
R1798 vdd.n2178 vdd.n807 185
R1799 vdd.n1938 vdd.n1937 185
R1800 vdd.n1937 vdd.n805 185
R1801 vdd.n1939 vdd.n812 185
R1802 vdd.n2172 vdd.n812 185
R1803 vdd.n1962 vdd.n1961 185
R1804 vdd.n1961 vdd.n1960 185
R1805 vdd.n1963 vdd.n817 185
R1806 vdd.n2166 vdd.n817 185
R1807 vdd.n1965 vdd.n1964 185
R1808 vdd.n1964 vdd.n823 185
R1809 vdd.n1966 vdd.n822 185
R1810 vdd.n2160 vdd.n822 185
R1811 vdd.n1968 vdd.n1967 185
R1812 vdd.n1967 vdd.n829 185
R1813 vdd.n1969 vdd.n828 185
R1814 vdd.n2154 vdd.n828 185
R1815 vdd.n1971 vdd.n1970 185
R1816 vdd.n1972 vdd.n1971 185
R1817 vdd.n1931 vdd.n835 185
R1818 vdd.n2148 vdd.n835 185
R1819 vdd.n1930 vdd.n1929 185
R1820 vdd.n1929 vdd.n833 185
R1821 vdd.n1928 vdd.n841 185
R1822 vdd.n2142 vdd.n841 185
R1823 vdd.n1927 vdd.n1926 185
R1824 vdd.n1926 vdd.n839 185
R1825 vdd.n1925 vdd.n846 185
R1826 vdd.n2136 vdd.n846 185
R1827 vdd.n1924 vdd.n1923 185
R1828 vdd.n1923 vdd.n853 185
R1829 vdd.n1922 vdd.n852 185
R1830 vdd.n2129 vdd.n852 185
R1831 vdd.n1921 vdd.n1920 185
R1832 vdd.n1920 vdd.n860 185
R1833 vdd.n1919 vdd.n859 185
R1834 vdd.n2123 vdd.n859 185
R1835 vdd.n1918 vdd.n1917 185
R1836 vdd.n1917 vdd.n857 185
R1837 vdd.n1916 vdd.n866 185
R1838 vdd.n2117 vdd.n866 185
R1839 vdd.n1915 vdd.n1914 185
R1840 vdd.n1914 vdd.n864 185
R1841 vdd.n1913 vdd.n872 185
R1842 vdd.n2111 vdd.n872 185
R1843 vdd.n1912 vdd.n1911 185
R1844 vdd.n1911 vdd.n870 185
R1845 vdd.n1910 vdd.n878 185
R1846 vdd.n2105 vdd.n878 185
R1847 vdd.n1909 vdd.n1908 185
R1848 vdd.n1908 vdd.n876 185
R1849 vdd.n1907 vdd.n884 185
R1850 vdd.n2099 vdd.n884 185
R1851 vdd.n1906 vdd.n1905 185
R1852 vdd.n1905 vdd.n882 185
R1853 vdd.n1904 vdd.n890 185
R1854 vdd.n2093 vdd.n890 185
R1855 vdd.n1903 vdd.n1902 185
R1856 vdd.n1902 vdd.n888 185
R1857 vdd.n1901 vdd.n896 185
R1858 vdd.n2087 vdd.n896 185
R1859 vdd.n1900 vdd.n1899 185
R1860 vdd.n1899 vdd.n894 185
R1861 vdd.n1898 vdd.n902 185
R1862 vdd.n2081 vdd.n902 185
R1863 vdd.n899 vdd.n898 185
R1864 vdd.n1830 vdd.n1828 185
R1865 vdd.n1833 vdd.n1832 185
R1866 vdd.n1834 vdd.n1827 185
R1867 vdd.n1836 vdd.n1835 185
R1868 vdd.n1838 vdd.n1826 185
R1869 vdd.n1841 vdd.n1840 185
R1870 vdd.n1842 vdd.n1825 185
R1871 vdd.n1844 vdd.n1843 185
R1872 vdd.n1846 vdd.n1824 185
R1873 vdd.n1849 vdd.n1848 185
R1874 vdd.n1850 vdd.n1823 185
R1875 vdd.n1852 vdd.n1851 185
R1876 vdd.n1854 vdd.n1822 185
R1877 vdd.n1857 vdd.n1856 185
R1878 vdd.n1858 vdd.n1821 185
R1879 vdd.n1860 vdd.n1859 185
R1880 vdd.n1862 vdd.n1820 185
R1881 vdd.n1865 vdd.n1864 185
R1882 vdd.n1866 vdd.n933 185
R1883 vdd.n1868 vdd.n1867 185
R1884 vdd.n1870 vdd.n932 185
R1885 vdd.n1873 vdd.n1872 185
R1886 vdd.n1874 vdd.n931 185
R1887 vdd.n1876 vdd.n1875 185
R1888 vdd.n1878 vdd.n930 185
R1889 vdd.n1881 vdd.n1880 185
R1890 vdd.n1882 vdd.n929 185
R1891 vdd.n1884 vdd.n1883 185
R1892 vdd.n1886 vdd.n928 185
R1893 vdd.n1889 vdd.n1888 185
R1894 vdd.n1890 vdd.n925 185
R1895 vdd.n1893 vdd.n1892 185
R1896 vdd.n1895 vdd.n924 185
R1897 vdd.n1897 vdd.n1896 185
R1898 vdd.n1896 vdd.n900 185
R1899 vdd.n291 vdd.n290 171.744
R1900 vdd.n290 vdd.n289 171.744
R1901 vdd.n289 vdd.n258 171.744
R1902 vdd.n282 vdd.n258 171.744
R1903 vdd.n282 vdd.n281 171.744
R1904 vdd.n281 vdd.n263 171.744
R1905 vdd.n274 vdd.n263 171.744
R1906 vdd.n274 vdd.n273 171.744
R1907 vdd.n273 vdd.n267 171.744
R1908 vdd.n244 vdd.n243 171.744
R1909 vdd.n243 vdd.n242 171.744
R1910 vdd.n242 vdd.n211 171.744
R1911 vdd.n235 vdd.n211 171.744
R1912 vdd.n235 vdd.n234 171.744
R1913 vdd.n234 vdd.n216 171.744
R1914 vdd.n227 vdd.n216 171.744
R1915 vdd.n227 vdd.n226 171.744
R1916 vdd.n226 vdd.n220 171.744
R1917 vdd.n201 vdd.n200 171.744
R1918 vdd.n200 vdd.n199 171.744
R1919 vdd.n199 vdd.n168 171.744
R1920 vdd.n192 vdd.n168 171.744
R1921 vdd.n192 vdd.n191 171.744
R1922 vdd.n191 vdd.n173 171.744
R1923 vdd.n184 vdd.n173 171.744
R1924 vdd.n184 vdd.n183 171.744
R1925 vdd.n183 vdd.n177 171.744
R1926 vdd.n154 vdd.n153 171.744
R1927 vdd.n153 vdd.n152 171.744
R1928 vdd.n152 vdd.n121 171.744
R1929 vdd.n145 vdd.n121 171.744
R1930 vdd.n145 vdd.n144 171.744
R1931 vdd.n144 vdd.n126 171.744
R1932 vdd.n137 vdd.n126 171.744
R1933 vdd.n137 vdd.n136 171.744
R1934 vdd.n136 vdd.n130 171.744
R1935 vdd.n112 vdd.n111 171.744
R1936 vdd.n111 vdd.n110 171.744
R1937 vdd.n110 vdd.n79 171.744
R1938 vdd.n103 vdd.n79 171.744
R1939 vdd.n103 vdd.n102 171.744
R1940 vdd.n102 vdd.n84 171.744
R1941 vdd.n95 vdd.n84 171.744
R1942 vdd.n95 vdd.n94 171.744
R1943 vdd.n94 vdd.n88 171.744
R1944 vdd.n65 vdd.n64 171.744
R1945 vdd.n64 vdd.n63 171.744
R1946 vdd.n63 vdd.n32 171.744
R1947 vdd.n56 vdd.n32 171.744
R1948 vdd.n56 vdd.n55 171.744
R1949 vdd.n55 vdd.n37 171.744
R1950 vdd.n48 vdd.n37 171.744
R1951 vdd.n48 vdd.n47 171.744
R1952 vdd.n47 vdd.n41 171.744
R1953 vdd.n1186 vdd.n1185 171.744
R1954 vdd.n1185 vdd.n1184 171.744
R1955 vdd.n1184 vdd.n1153 171.744
R1956 vdd.n1177 vdd.n1153 171.744
R1957 vdd.n1177 vdd.n1176 171.744
R1958 vdd.n1176 vdd.n1158 171.744
R1959 vdd.n1169 vdd.n1158 171.744
R1960 vdd.n1169 vdd.n1168 171.744
R1961 vdd.n1168 vdd.n1162 171.744
R1962 vdd.n1233 vdd.n1232 171.744
R1963 vdd.n1232 vdd.n1231 171.744
R1964 vdd.n1231 vdd.n1200 171.744
R1965 vdd.n1224 vdd.n1200 171.744
R1966 vdd.n1224 vdd.n1223 171.744
R1967 vdd.n1223 vdd.n1205 171.744
R1968 vdd.n1216 vdd.n1205 171.744
R1969 vdd.n1216 vdd.n1215 171.744
R1970 vdd.n1215 vdd.n1209 171.744
R1971 vdd.n1096 vdd.n1095 171.744
R1972 vdd.n1095 vdd.n1094 171.744
R1973 vdd.n1094 vdd.n1063 171.744
R1974 vdd.n1087 vdd.n1063 171.744
R1975 vdd.n1087 vdd.n1086 171.744
R1976 vdd.n1086 vdd.n1068 171.744
R1977 vdd.n1079 vdd.n1068 171.744
R1978 vdd.n1079 vdd.n1078 171.744
R1979 vdd.n1078 vdd.n1072 171.744
R1980 vdd.n1143 vdd.n1142 171.744
R1981 vdd.n1142 vdd.n1141 171.744
R1982 vdd.n1141 vdd.n1110 171.744
R1983 vdd.n1134 vdd.n1110 171.744
R1984 vdd.n1134 vdd.n1133 171.744
R1985 vdd.n1133 vdd.n1115 171.744
R1986 vdd.n1126 vdd.n1115 171.744
R1987 vdd.n1126 vdd.n1125 171.744
R1988 vdd.n1125 vdd.n1119 171.744
R1989 vdd.n1007 vdd.n1006 171.744
R1990 vdd.n1006 vdd.n1005 171.744
R1991 vdd.n1005 vdd.n974 171.744
R1992 vdd.n998 vdd.n974 171.744
R1993 vdd.n998 vdd.n997 171.744
R1994 vdd.n997 vdd.n979 171.744
R1995 vdd.n990 vdd.n979 171.744
R1996 vdd.n990 vdd.n989 171.744
R1997 vdd.n989 vdd.n983 171.744
R1998 vdd.n1054 vdd.n1053 171.744
R1999 vdd.n1053 vdd.n1052 171.744
R2000 vdd.n1052 vdd.n1021 171.744
R2001 vdd.n1045 vdd.n1021 171.744
R2002 vdd.n1045 vdd.n1044 171.744
R2003 vdd.n1044 vdd.n1026 171.744
R2004 vdd.n1037 vdd.n1026 171.744
R2005 vdd.n1037 vdd.n1036 171.744
R2006 vdd.n1036 vdd.n1030 171.744
R2007 vdd.n3199 vdd.n334 146.341
R2008 vdd.n3197 vdd.n3196 146.341
R2009 vdd.n3194 vdd.n338 146.341
R2010 vdd.n3190 vdd.n3189 146.341
R2011 vdd.n3187 vdd.n346 146.341
R2012 vdd.n3183 vdd.n3182 146.341
R2013 vdd.n3180 vdd.n353 146.341
R2014 vdd.n3176 vdd.n3175 146.341
R2015 vdd.n3173 vdd.n360 146.341
R2016 vdd.n371 vdd.n368 146.341
R2017 vdd.n3165 vdd.n3164 146.341
R2018 vdd.n3162 vdd.n373 146.341
R2019 vdd.n3158 vdd.n3157 146.341
R2020 vdd.n3155 vdd.n379 146.341
R2021 vdd.n3151 vdd.n3150 146.341
R2022 vdd.n3148 vdd.n386 146.341
R2023 vdd.n3144 vdd.n3143 146.341
R2024 vdd.n3141 vdd.n393 146.341
R2025 vdd.n3137 vdd.n3136 146.341
R2026 vdd.n3134 vdd.n400 146.341
R2027 vdd.n411 vdd.n408 146.341
R2028 vdd.n3126 vdd.n3125 146.341
R2029 vdd.n3123 vdd.n413 146.341
R2030 vdd.n3119 vdd.n3118 146.341
R2031 vdd.n3116 vdd.n419 146.341
R2032 vdd.n3112 vdd.n3111 146.341
R2033 vdd.n3109 vdd.n426 146.341
R2034 vdd.n3105 vdd.n3104 146.341
R2035 vdd.n3102 vdd.n433 146.341
R2036 vdd.n3098 vdd.n3097 146.341
R2037 vdd.n3095 vdd.n440 146.341
R2038 vdd.n3032 vdd.n478 146.341
R2039 vdd.n3032 vdd.n474 146.341
R2040 vdd.n3038 vdd.n474 146.341
R2041 vdd.n3038 vdd.n466 146.341
R2042 vdd.n3049 vdd.n466 146.341
R2043 vdd.n3049 vdd.n462 146.341
R2044 vdd.n3055 vdd.n462 146.341
R2045 vdd.n3055 vdd.n454 146.341
R2046 vdd.n3065 vdd.n454 146.341
R2047 vdd.n3065 vdd.n455 146.341
R2048 vdd.n455 vdd.n305 146.341
R2049 vdd.n306 vdd.n305 146.341
R2050 vdd.n307 vdd.n306 146.341
R2051 vdd.n448 vdd.n307 146.341
R2052 vdd.n448 vdd.n315 146.341
R2053 vdd.n316 vdd.n315 146.341
R2054 vdd.n317 vdd.n316 146.341
R2055 vdd.n445 vdd.n317 146.341
R2056 vdd.n445 vdd.n326 146.341
R2057 vdd.n327 vdd.n326 146.341
R2058 vdd.n328 vdd.n327 146.341
R2059 vdd.n3021 vdd.n483 146.341
R2060 vdd.n3021 vdd.n517 146.341
R2061 vdd.n523 vdd.n522 146.341
R2062 vdd.n3014 vdd.n3013 146.341
R2063 vdd.n3010 vdd.n3009 146.341
R2064 vdd.n3006 vdd.n3005 146.341
R2065 vdd.n3002 vdd.n3001 146.341
R2066 vdd.n2998 vdd.n2997 146.341
R2067 vdd.n2994 vdd.n2993 146.341
R2068 vdd.n2990 vdd.n2989 146.341
R2069 vdd.n2981 vdd.n2980 146.341
R2070 vdd.n2978 vdd.n2977 146.341
R2071 vdd.n2974 vdd.n2973 146.341
R2072 vdd.n2970 vdd.n2969 146.341
R2073 vdd.n2966 vdd.n2965 146.341
R2074 vdd.n2962 vdd.n2961 146.341
R2075 vdd.n2958 vdd.n2957 146.341
R2076 vdd.n2954 vdd.n2953 146.341
R2077 vdd.n2950 vdd.n2949 146.341
R2078 vdd.n2946 vdd.n2945 146.341
R2079 vdd.n2942 vdd.n2941 146.341
R2080 vdd.n2935 vdd.n2934 146.341
R2081 vdd.n2932 vdd.n2931 146.341
R2082 vdd.n2928 vdd.n2927 146.341
R2083 vdd.n2924 vdd.n2923 146.341
R2084 vdd.n2920 vdd.n2919 146.341
R2085 vdd.n2916 vdd.n2915 146.341
R2086 vdd.n2912 vdd.n2911 146.341
R2087 vdd.n2908 vdd.n2907 146.341
R2088 vdd.n2904 vdd.n2903 146.341
R2089 vdd.n2900 vdd.n2899 146.341
R2090 vdd.n2896 vdd.n515 146.341
R2091 vdd.n3030 vdd.n479 146.341
R2092 vdd.n3030 vdd.n472 146.341
R2093 vdd.n3041 vdd.n472 146.341
R2094 vdd.n3041 vdd.n468 146.341
R2095 vdd.n3047 vdd.n468 146.341
R2096 vdd.n3047 vdd.n461 146.341
R2097 vdd.n3057 vdd.n461 146.341
R2098 vdd.n3057 vdd.n457 146.341
R2099 vdd.n3063 vdd.n457 146.341
R2100 vdd.n3063 vdd.n302 146.341
R2101 vdd.n3226 vdd.n302 146.341
R2102 vdd.n3226 vdd.n303 146.341
R2103 vdd.n3222 vdd.n303 146.341
R2104 vdd.n3222 vdd.n309 146.341
R2105 vdd.n3218 vdd.n309 146.341
R2106 vdd.n3218 vdd.n314 146.341
R2107 vdd.n3214 vdd.n314 146.341
R2108 vdd.n3214 vdd.n319 146.341
R2109 vdd.n3210 vdd.n319 146.341
R2110 vdd.n3210 vdd.n325 146.341
R2111 vdd.n3206 vdd.n325 146.341
R2112 vdd.n1803 vdd.n1802 146.341
R2113 vdd.n1800 vdd.n1597 146.341
R2114 vdd.n1793 vdd.n1603 146.341
R2115 vdd.n1791 vdd.n1790 146.341
R2116 vdd.n1788 vdd.n1605 146.341
R2117 vdd.n1784 vdd.n1783 146.341
R2118 vdd.n1781 vdd.n1612 146.341
R2119 vdd.n1777 vdd.n1776 146.341
R2120 vdd.n1774 vdd.n1619 146.341
R2121 vdd.n1630 vdd.n1627 146.341
R2122 vdd.n1766 vdd.n1765 146.341
R2123 vdd.n1763 vdd.n1632 146.341
R2124 vdd.n1759 vdd.n1758 146.341
R2125 vdd.n1756 vdd.n1638 146.341
R2126 vdd.n1752 vdd.n1751 146.341
R2127 vdd.n1749 vdd.n1645 146.341
R2128 vdd.n1745 vdd.n1744 146.341
R2129 vdd.n1742 vdd.n1652 146.341
R2130 vdd.n1738 vdd.n1737 146.341
R2131 vdd.n1735 vdd.n1659 146.341
R2132 vdd.n1670 vdd.n1667 146.341
R2133 vdd.n1727 vdd.n1726 146.341
R2134 vdd.n1724 vdd.n1672 146.341
R2135 vdd.n1720 vdd.n1719 146.341
R2136 vdd.n1717 vdd.n1678 146.341
R2137 vdd.n1713 vdd.n1712 146.341
R2138 vdd.n1710 vdd.n1685 146.341
R2139 vdd.n1706 vdd.n1705 146.341
R2140 vdd.n1703 vdd.n1700 146.341
R2141 vdd.n1698 vdd.n1695 146.341
R2142 vdd.n1693 vdd.n939 146.341
R2143 vdd.n1511 vdd.n1271 146.341
R2144 vdd.n1511 vdd.n1267 146.341
R2145 vdd.n1517 vdd.n1267 146.341
R2146 vdd.n1517 vdd.n1259 146.341
R2147 vdd.n1528 vdd.n1259 146.341
R2148 vdd.n1528 vdd.n1255 146.341
R2149 vdd.n1534 vdd.n1255 146.341
R2150 vdd.n1534 vdd.n1249 146.341
R2151 vdd.n1546 vdd.n1249 146.341
R2152 vdd.n1546 vdd.n1245 146.341
R2153 vdd.n1552 vdd.n1245 146.341
R2154 vdd.n1552 vdd.n966 146.341
R2155 vdd.n1562 vdd.n966 146.341
R2156 vdd.n1562 vdd.n962 146.341
R2157 vdd.n1568 vdd.n962 146.341
R2158 vdd.n1568 vdd.n956 146.341
R2159 vdd.n1579 vdd.n956 146.341
R2160 vdd.n1579 vdd.n951 146.341
R2161 vdd.n1587 vdd.n951 146.341
R2162 vdd.n1587 vdd.n941 146.341
R2163 vdd.n1811 vdd.n941 146.341
R2164 vdd.n1500 vdd.n1276 146.341
R2165 vdd.n1500 vdd.n1309 146.341
R2166 vdd.n1313 vdd.n1312 146.341
R2167 vdd.n1315 vdd.n1314 146.341
R2168 vdd.n1319 vdd.n1318 146.341
R2169 vdd.n1321 vdd.n1320 146.341
R2170 vdd.n1325 vdd.n1324 146.341
R2171 vdd.n1327 vdd.n1326 146.341
R2172 vdd.n1331 vdd.n1330 146.341
R2173 vdd.n1333 vdd.n1332 146.341
R2174 vdd.n1339 vdd.n1338 146.341
R2175 vdd.n1341 vdd.n1340 146.341
R2176 vdd.n1345 vdd.n1344 146.341
R2177 vdd.n1347 vdd.n1346 146.341
R2178 vdd.n1351 vdd.n1350 146.341
R2179 vdd.n1353 vdd.n1352 146.341
R2180 vdd.n1357 vdd.n1356 146.341
R2181 vdd.n1359 vdd.n1358 146.341
R2182 vdd.n1363 vdd.n1362 146.341
R2183 vdd.n1365 vdd.n1364 146.341
R2184 vdd.n1437 vdd.n1368 146.341
R2185 vdd.n1370 vdd.n1369 146.341
R2186 vdd.n1374 vdd.n1373 146.341
R2187 vdd.n1376 vdd.n1375 146.341
R2188 vdd.n1380 vdd.n1379 146.341
R2189 vdd.n1382 vdd.n1381 146.341
R2190 vdd.n1386 vdd.n1385 146.341
R2191 vdd.n1388 vdd.n1387 146.341
R2192 vdd.n1392 vdd.n1391 146.341
R2193 vdd.n1394 vdd.n1393 146.341
R2194 vdd.n1398 vdd.n1397 146.341
R2195 vdd.n1399 vdd.n1307 146.341
R2196 vdd.n1509 vdd.n1272 146.341
R2197 vdd.n1509 vdd.n1265 146.341
R2198 vdd.n1520 vdd.n1265 146.341
R2199 vdd.n1520 vdd.n1261 146.341
R2200 vdd.n1526 vdd.n1261 146.341
R2201 vdd.n1526 vdd.n1254 146.341
R2202 vdd.n1537 vdd.n1254 146.341
R2203 vdd.n1537 vdd.n1250 146.341
R2204 vdd.n1544 vdd.n1250 146.341
R2205 vdd.n1544 vdd.n1243 146.341
R2206 vdd.n1554 vdd.n1243 146.341
R2207 vdd.n1554 vdd.n969 146.341
R2208 vdd.n1560 vdd.n969 146.341
R2209 vdd.n1560 vdd.n961 146.341
R2210 vdd.n1571 vdd.n961 146.341
R2211 vdd.n1571 vdd.n957 146.341
R2212 vdd.n1577 vdd.n957 146.341
R2213 vdd.n1577 vdd.n949 146.341
R2214 vdd.n1590 vdd.n949 146.341
R2215 vdd.n1590 vdd.n944 146.341
R2216 vdd.n1809 vdd.n944 146.341
R2217 vdd.n926 vdd.t47 127.284
R2218 vdd.n787 vdd.t76 127.284
R2219 vdd.n920 vdd.t97 127.284
R2220 vdd.n778 vdd.t93 127.284
R2221 vdd.n675 vdd.t56 127.284
R2222 vdd.n675 vdd.t57 127.284
R2223 vdd.n2375 vdd.t91 127.284
R2224 vdd.n622 vdd.t69 127.284
R2225 vdd.n2444 vdd.t81 127.284
R2226 vdd.n589 vdd.t42 127.284
R2227 vdd.n848 vdd.t87 127.284
R2228 vdd.n848 vdd.t88 127.284
R2229 vdd.n22 vdd.n20 117.314
R2230 vdd.n17 vdd.n15 117.314
R2231 vdd.n27 vdd.n26 116.927
R2232 vdd.n24 vdd.n23 116.927
R2233 vdd.n22 vdd.n21 116.927
R2234 vdd.n17 vdd.n16 116.927
R2235 vdd.n19 vdd.n18 116.927
R2236 vdd.n27 vdd.n25 116.927
R2237 vdd.n927 vdd.t46 111.188
R2238 vdd.n788 vdd.t77 111.188
R2239 vdd.n921 vdd.t96 111.188
R2240 vdd.n779 vdd.t94 111.188
R2241 vdd.n2376 vdd.t90 111.188
R2242 vdd.n623 vdd.t70 111.188
R2243 vdd.n2445 vdd.t80 111.188
R2244 vdd.n590 vdd.t43 111.188
R2245 vdd.n2630 vdd.n728 99.5127
R2246 vdd.n2638 vdd.n728 99.5127
R2247 vdd.n2638 vdd.n726 99.5127
R2248 vdd.n2642 vdd.n726 99.5127
R2249 vdd.n2642 vdd.n716 99.5127
R2250 vdd.n2650 vdd.n716 99.5127
R2251 vdd.n2650 vdd.n714 99.5127
R2252 vdd.n2654 vdd.n714 99.5127
R2253 vdd.n2654 vdd.n706 99.5127
R2254 vdd.n2662 vdd.n706 99.5127
R2255 vdd.n2662 vdd.n704 99.5127
R2256 vdd.n2666 vdd.n704 99.5127
R2257 vdd.n2666 vdd.n694 99.5127
R2258 vdd.n2674 vdd.n694 99.5127
R2259 vdd.n2674 vdd.n692 99.5127
R2260 vdd.n2678 vdd.n692 99.5127
R2261 vdd.n2678 vdd.n683 99.5127
R2262 vdd.n2686 vdd.n683 99.5127
R2263 vdd.n2686 vdd.n681 99.5127
R2264 vdd.n2690 vdd.n681 99.5127
R2265 vdd.n2690 vdd.n670 99.5127
R2266 vdd.n2699 vdd.n670 99.5127
R2267 vdd.n2699 vdd.n668 99.5127
R2268 vdd.n2703 vdd.n668 99.5127
R2269 vdd.n2703 vdd.n657 99.5127
R2270 vdd.n2711 vdd.n657 99.5127
R2271 vdd.n2711 vdd.n655 99.5127
R2272 vdd.n2715 vdd.n655 99.5127
R2273 vdd.n2715 vdd.n646 99.5127
R2274 vdd.n2723 vdd.n646 99.5127
R2275 vdd.n2723 vdd.n644 99.5127
R2276 vdd.n2727 vdd.n644 99.5127
R2277 vdd.n2727 vdd.n632 99.5127
R2278 vdd.n2780 vdd.n632 99.5127
R2279 vdd.n2780 vdd.n630 99.5127
R2280 vdd.n2784 vdd.n630 99.5127
R2281 vdd.n2784 vdd.n598 99.5127
R2282 vdd.n2854 vdd.n598 99.5127
R2283 vdd.n2850 vdd.n599 99.5127
R2284 vdd.n2848 vdd.n2847 99.5127
R2285 vdd.n2845 vdd.n603 99.5127
R2286 vdd.n2841 vdd.n2840 99.5127
R2287 vdd.n2838 vdd.n606 99.5127
R2288 vdd.n2834 vdd.n2833 99.5127
R2289 vdd.n2831 vdd.n609 99.5127
R2290 vdd.n2827 vdd.n2826 99.5127
R2291 vdd.n2824 vdd.n2822 99.5127
R2292 vdd.n2820 vdd.n612 99.5127
R2293 vdd.n2816 vdd.n2815 99.5127
R2294 vdd.n2813 vdd.n615 99.5127
R2295 vdd.n2809 vdd.n2808 99.5127
R2296 vdd.n2806 vdd.n618 99.5127
R2297 vdd.n2802 vdd.n2801 99.5127
R2298 vdd.n2799 vdd.n621 99.5127
R2299 vdd.n2794 vdd.n2793 99.5127
R2300 vdd.n2512 vdd.n734 99.5127
R2301 vdd.n2512 vdd.n729 99.5127
R2302 vdd.n2614 vdd.n729 99.5127
R2303 vdd.n2614 vdd.n724 99.5127
R2304 vdd.n2610 vdd.n724 99.5127
R2305 vdd.n2610 vdd.n718 99.5127
R2306 vdd.n2607 vdd.n718 99.5127
R2307 vdd.n2607 vdd.n712 99.5127
R2308 vdd.n2604 vdd.n712 99.5127
R2309 vdd.n2604 vdd.n707 99.5127
R2310 vdd.n2554 vdd.n707 99.5127
R2311 vdd.n2554 vdd.n702 99.5127
R2312 vdd.n2557 vdd.n702 99.5127
R2313 vdd.n2557 vdd.n696 99.5127
R2314 vdd.n2590 vdd.n696 99.5127
R2315 vdd.n2590 vdd.n689 99.5127
R2316 vdd.n2586 vdd.n689 99.5127
R2317 vdd.n2586 vdd.n684 99.5127
R2318 vdd.n2583 vdd.n684 99.5127
R2319 vdd.n2583 vdd.n679 99.5127
R2320 vdd.n2580 vdd.n679 99.5127
R2321 vdd.n2580 vdd.n672 99.5127
R2322 vdd.n2577 vdd.n672 99.5127
R2323 vdd.n2577 vdd.n665 99.5127
R2324 vdd.n2574 vdd.n665 99.5127
R2325 vdd.n2574 vdd.n658 99.5127
R2326 vdd.n2571 vdd.n658 99.5127
R2327 vdd.n2571 vdd.n652 99.5127
R2328 vdd.n2568 vdd.n652 99.5127
R2329 vdd.n2568 vdd.n647 99.5127
R2330 vdd.n2565 vdd.n647 99.5127
R2331 vdd.n2565 vdd.n642 99.5127
R2332 vdd.n2562 vdd.n642 99.5127
R2333 vdd.n2562 vdd.n634 99.5127
R2334 vdd.n634 vdd.n627 99.5127
R2335 vdd.n2786 vdd.n627 99.5127
R2336 vdd.n2787 vdd.n2786 99.5127
R2337 vdd.n2787 vdd.n596 99.5127
R2338 vdd.n2626 vdd.n739 99.5127
R2339 vdd.n2446 vdd.n739 99.5127
R2340 vdd.n2450 vdd.n2449 99.5127
R2341 vdd.n2454 vdd.n2453 99.5127
R2342 vdd.n2458 vdd.n2457 99.5127
R2343 vdd.n2462 vdd.n2461 99.5127
R2344 vdd.n2466 vdd.n2465 99.5127
R2345 vdd.n2470 vdd.n2469 99.5127
R2346 vdd.n2474 vdd.n2473 99.5127
R2347 vdd.n2478 vdd.n2477 99.5127
R2348 vdd.n2482 vdd.n2481 99.5127
R2349 vdd.n2486 vdd.n2485 99.5127
R2350 vdd.n2490 vdd.n2489 99.5127
R2351 vdd.n2494 vdd.n2493 99.5127
R2352 vdd.n2498 vdd.n2497 99.5127
R2353 vdd.n2502 vdd.n2501 99.5127
R2354 vdd.n2507 vdd.n2506 99.5127
R2355 vdd.n2339 vdd.n776 99.5127
R2356 vdd.n2335 vdd.n2334 99.5127
R2357 vdd.n2331 vdd.n2330 99.5127
R2358 vdd.n2327 vdd.n2326 99.5127
R2359 vdd.n2323 vdd.n2322 99.5127
R2360 vdd.n2319 vdd.n2318 99.5127
R2361 vdd.n2315 vdd.n2314 99.5127
R2362 vdd.n2311 vdd.n2310 99.5127
R2363 vdd.n2307 vdd.n2306 99.5127
R2364 vdd.n2303 vdd.n2302 99.5127
R2365 vdd.n2299 vdd.n2298 99.5127
R2366 vdd.n2295 vdd.n2294 99.5127
R2367 vdd.n2291 vdd.n2290 99.5127
R2368 vdd.n2287 vdd.n2286 99.5127
R2369 vdd.n2283 vdd.n2282 99.5127
R2370 vdd.n2279 vdd.n2278 99.5127
R2371 vdd.n2274 vdd.n2273 99.5127
R2372 vdd.n2006 vdd.n901 99.5127
R2373 vdd.n2006 vdd.n895 99.5127
R2374 vdd.n2003 vdd.n895 99.5127
R2375 vdd.n2003 vdd.n889 99.5127
R2376 vdd.n2000 vdd.n889 99.5127
R2377 vdd.n2000 vdd.n883 99.5127
R2378 vdd.n1997 vdd.n883 99.5127
R2379 vdd.n1997 vdd.n877 99.5127
R2380 vdd.n1994 vdd.n877 99.5127
R2381 vdd.n1994 vdd.n871 99.5127
R2382 vdd.n1991 vdd.n871 99.5127
R2383 vdd.n1991 vdd.n865 99.5127
R2384 vdd.n1988 vdd.n865 99.5127
R2385 vdd.n1988 vdd.n858 99.5127
R2386 vdd.n1985 vdd.n858 99.5127
R2387 vdd.n1985 vdd.n851 99.5127
R2388 vdd.n1982 vdd.n851 99.5127
R2389 vdd.n1982 vdd.n845 99.5127
R2390 vdd.n1979 vdd.n845 99.5127
R2391 vdd.n1979 vdd.n840 99.5127
R2392 vdd.n1976 vdd.n840 99.5127
R2393 vdd.n1976 vdd.n834 99.5127
R2394 vdd.n1973 vdd.n834 99.5127
R2395 vdd.n1973 vdd.n827 99.5127
R2396 vdd.n1940 vdd.n827 99.5127
R2397 vdd.n1940 vdd.n821 99.5127
R2398 vdd.n1943 vdd.n821 99.5127
R2399 vdd.n1943 vdd.n816 99.5127
R2400 vdd.n1959 vdd.n816 99.5127
R2401 vdd.n1959 vdd.n811 99.5127
R2402 vdd.n1955 vdd.n811 99.5127
R2403 vdd.n1955 vdd.n806 99.5127
R2404 vdd.n1952 vdd.n806 99.5127
R2405 vdd.n1952 vdd.n799 99.5127
R2406 vdd.n1949 vdd.n799 99.5127
R2407 vdd.n1949 vdd.n792 99.5127
R2408 vdd.n792 vdd.n781 99.5127
R2409 vdd.n2269 vdd.n781 99.5127
R2410 vdd.n2076 vdd.n2074 99.5127
R2411 vdd.n2074 vdd.n2073 99.5127
R2412 vdd.n2070 vdd.n2069 99.5127
R2413 vdd.n2067 vdd.n907 99.5127
R2414 vdd.n2063 vdd.n2061 99.5127
R2415 vdd.n2059 vdd.n909 99.5127
R2416 vdd.n2055 vdd.n2053 99.5127
R2417 vdd.n2051 vdd.n911 99.5127
R2418 vdd.n2047 vdd.n2045 99.5127
R2419 vdd.n2043 vdd.n913 99.5127
R2420 vdd.n2039 vdd.n2037 99.5127
R2421 vdd.n2035 vdd.n915 99.5127
R2422 vdd.n2031 vdd.n2029 99.5127
R2423 vdd.n2027 vdd.n917 99.5127
R2424 vdd.n2023 vdd.n2021 99.5127
R2425 vdd.n2019 vdd.n919 99.5127
R2426 vdd.n2014 vdd.n2012 99.5127
R2427 vdd.n2080 vdd.n893 99.5127
R2428 vdd.n2088 vdd.n893 99.5127
R2429 vdd.n2088 vdd.n891 99.5127
R2430 vdd.n2092 vdd.n891 99.5127
R2431 vdd.n2092 vdd.n881 99.5127
R2432 vdd.n2100 vdd.n881 99.5127
R2433 vdd.n2100 vdd.n879 99.5127
R2434 vdd.n2104 vdd.n879 99.5127
R2435 vdd.n2104 vdd.n869 99.5127
R2436 vdd.n2112 vdd.n869 99.5127
R2437 vdd.n2112 vdd.n867 99.5127
R2438 vdd.n2116 vdd.n867 99.5127
R2439 vdd.n2116 vdd.n856 99.5127
R2440 vdd.n2124 vdd.n856 99.5127
R2441 vdd.n2124 vdd.n854 99.5127
R2442 vdd.n2128 vdd.n854 99.5127
R2443 vdd.n2128 vdd.n844 99.5127
R2444 vdd.n2137 vdd.n844 99.5127
R2445 vdd.n2137 vdd.n842 99.5127
R2446 vdd.n2141 vdd.n842 99.5127
R2447 vdd.n2141 vdd.n832 99.5127
R2448 vdd.n2149 vdd.n832 99.5127
R2449 vdd.n2149 vdd.n830 99.5127
R2450 vdd.n2153 vdd.n830 99.5127
R2451 vdd.n2153 vdd.n820 99.5127
R2452 vdd.n2161 vdd.n820 99.5127
R2453 vdd.n2161 vdd.n818 99.5127
R2454 vdd.n2165 vdd.n818 99.5127
R2455 vdd.n2165 vdd.n810 99.5127
R2456 vdd.n2173 vdd.n810 99.5127
R2457 vdd.n2173 vdd.n808 99.5127
R2458 vdd.n2177 vdd.n808 99.5127
R2459 vdd.n2177 vdd.n797 99.5127
R2460 vdd.n2187 vdd.n797 99.5127
R2461 vdd.n2187 vdd.n794 99.5127
R2462 vdd.n2192 vdd.n794 99.5127
R2463 vdd.n2192 vdd.n795 99.5127
R2464 vdd.n795 vdd.n775 99.5127
R2465 vdd.n2770 vdd.n2769 99.5127
R2466 vdd.n2767 vdd.n2733 99.5127
R2467 vdd.n2763 vdd.n2762 99.5127
R2468 vdd.n2760 vdd.n2736 99.5127
R2469 vdd.n2756 vdd.n2755 99.5127
R2470 vdd.n2753 vdd.n2739 99.5127
R2471 vdd.n2749 vdd.n2748 99.5127
R2472 vdd.n2746 vdd.n2743 99.5127
R2473 vdd.n2887 vdd.n577 99.5127
R2474 vdd.n2885 vdd.n2884 99.5127
R2475 vdd.n2882 vdd.n579 99.5127
R2476 vdd.n2878 vdd.n2877 99.5127
R2477 vdd.n2875 vdd.n582 99.5127
R2478 vdd.n2871 vdd.n2870 99.5127
R2479 vdd.n2868 vdd.n585 99.5127
R2480 vdd.n2864 vdd.n2863 99.5127
R2481 vdd.n2861 vdd.n588 99.5127
R2482 vdd.n2619 vdd.n735 99.5127
R2483 vdd.n2619 vdd.n730 99.5127
R2484 vdd.n2616 vdd.n730 99.5127
R2485 vdd.n2616 vdd.n725 99.5127
R2486 vdd.n2516 vdd.n725 99.5127
R2487 vdd.n2516 vdd.n719 99.5127
R2488 vdd.n2519 vdd.n719 99.5127
R2489 vdd.n2519 vdd.n713 99.5127
R2490 vdd.n2602 vdd.n713 99.5127
R2491 vdd.n2602 vdd.n708 99.5127
R2492 vdd.n2598 vdd.n708 99.5127
R2493 vdd.n2598 vdd.n703 99.5127
R2494 vdd.n2595 vdd.n703 99.5127
R2495 vdd.n2595 vdd.n697 99.5127
R2496 vdd.n2592 vdd.n697 99.5127
R2497 vdd.n2592 vdd.n690 99.5127
R2498 vdd.n2551 vdd.n690 99.5127
R2499 vdd.n2551 vdd.n685 99.5127
R2500 vdd.n2548 vdd.n685 99.5127
R2501 vdd.n2548 vdd.n680 99.5127
R2502 vdd.n2545 vdd.n680 99.5127
R2503 vdd.n2545 vdd.n673 99.5127
R2504 vdd.n2542 vdd.n673 99.5127
R2505 vdd.n2542 vdd.n666 99.5127
R2506 vdd.n2539 vdd.n666 99.5127
R2507 vdd.n2539 vdd.n659 99.5127
R2508 vdd.n2536 vdd.n659 99.5127
R2509 vdd.n2536 vdd.n653 99.5127
R2510 vdd.n2533 vdd.n653 99.5127
R2511 vdd.n2533 vdd.n648 99.5127
R2512 vdd.n2530 vdd.n648 99.5127
R2513 vdd.n2530 vdd.n643 99.5127
R2514 vdd.n2527 vdd.n643 99.5127
R2515 vdd.n2527 vdd.n635 99.5127
R2516 vdd.n2524 vdd.n635 99.5127
R2517 vdd.n2524 vdd.n628 99.5127
R2518 vdd.n628 vdd.n594 99.5127
R2519 vdd.n2856 vdd.n594 99.5127
R2520 vdd.n2380 vdd.n2379 99.5127
R2521 vdd.n2384 vdd.n2383 99.5127
R2522 vdd.n2388 vdd.n2387 99.5127
R2523 vdd.n2392 vdd.n2391 99.5127
R2524 vdd.n2396 vdd.n2395 99.5127
R2525 vdd.n2400 vdd.n2399 99.5127
R2526 vdd.n2404 vdd.n2403 99.5127
R2527 vdd.n2408 vdd.n2407 99.5127
R2528 vdd.n2412 vdd.n2411 99.5127
R2529 vdd.n2416 vdd.n2415 99.5127
R2530 vdd.n2420 vdd.n2419 99.5127
R2531 vdd.n2424 vdd.n2423 99.5127
R2532 vdd.n2428 vdd.n2427 99.5127
R2533 vdd.n2432 vdd.n2431 99.5127
R2534 vdd.n2436 vdd.n2435 99.5127
R2535 vdd.n2440 vdd.n2439 99.5127
R2536 vdd.n2623 vdd.n2374 99.5127
R2537 vdd.n2632 vdd.n731 99.5127
R2538 vdd.n2636 vdd.n731 99.5127
R2539 vdd.n2636 vdd.n723 99.5127
R2540 vdd.n2644 vdd.n723 99.5127
R2541 vdd.n2644 vdd.n721 99.5127
R2542 vdd.n2648 vdd.n721 99.5127
R2543 vdd.n2648 vdd.n711 99.5127
R2544 vdd.n2656 vdd.n711 99.5127
R2545 vdd.n2656 vdd.n709 99.5127
R2546 vdd.n2660 vdd.n709 99.5127
R2547 vdd.n2660 vdd.n700 99.5127
R2548 vdd.n2668 vdd.n700 99.5127
R2549 vdd.n2668 vdd.n698 99.5127
R2550 vdd.n2672 vdd.n698 99.5127
R2551 vdd.n2672 vdd.n688 99.5127
R2552 vdd.n2680 vdd.n688 99.5127
R2553 vdd.n2680 vdd.n686 99.5127
R2554 vdd.n2684 vdd.n686 99.5127
R2555 vdd.n2684 vdd.n677 99.5127
R2556 vdd.n2692 vdd.n677 99.5127
R2557 vdd.n2692 vdd.n674 99.5127
R2558 vdd.n2697 vdd.n674 99.5127
R2559 vdd.n2697 vdd.n663 99.5127
R2560 vdd.n2705 vdd.n663 99.5127
R2561 vdd.n2705 vdd.n661 99.5127
R2562 vdd.n2709 vdd.n661 99.5127
R2563 vdd.n2709 vdd.n651 99.5127
R2564 vdd.n2717 vdd.n651 99.5127
R2565 vdd.n2717 vdd.n649 99.5127
R2566 vdd.n2721 vdd.n649 99.5127
R2567 vdd.n2721 vdd.n640 99.5127
R2568 vdd.n2729 vdd.n640 99.5127
R2569 vdd.n2729 vdd.n637 99.5127
R2570 vdd.n2778 vdd.n637 99.5127
R2571 vdd.n2778 vdd.n638 99.5127
R2572 vdd.n638 vdd.n629 99.5127
R2573 vdd.n2773 vdd.n629 99.5127
R2574 vdd.n2773 vdd.n597 99.5127
R2575 vdd.n2263 vdd.n2262 99.5127
R2576 vdd.n2259 vdd.n2258 99.5127
R2577 vdd.n2255 vdd.n2254 99.5127
R2578 vdd.n2251 vdd.n2250 99.5127
R2579 vdd.n2247 vdd.n2246 99.5127
R2580 vdd.n2243 vdd.n2242 99.5127
R2581 vdd.n2239 vdd.n2238 99.5127
R2582 vdd.n2235 vdd.n2234 99.5127
R2583 vdd.n2231 vdd.n2230 99.5127
R2584 vdd.n2227 vdd.n2226 99.5127
R2585 vdd.n2223 vdd.n2222 99.5127
R2586 vdd.n2219 vdd.n2218 99.5127
R2587 vdd.n2215 vdd.n2214 99.5127
R2588 vdd.n2211 vdd.n2210 99.5127
R2589 vdd.n2207 vdd.n2206 99.5127
R2590 vdd.n2203 vdd.n2202 99.5127
R2591 vdd.n2199 vdd.n757 99.5127
R2592 vdd.n1899 vdd.n902 99.5127
R2593 vdd.n1899 vdd.n896 99.5127
R2594 vdd.n1902 vdd.n896 99.5127
R2595 vdd.n1902 vdd.n890 99.5127
R2596 vdd.n1905 vdd.n890 99.5127
R2597 vdd.n1905 vdd.n884 99.5127
R2598 vdd.n1908 vdd.n884 99.5127
R2599 vdd.n1908 vdd.n878 99.5127
R2600 vdd.n1911 vdd.n878 99.5127
R2601 vdd.n1911 vdd.n872 99.5127
R2602 vdd.n1914 vdd.n872 99.5127
R2603 vdd.n1914 vdd.n866 99.5127
R2604 vdd.n1917 vdd.n866 99.5127
R2605 vdd.n1917 vdd.n859 99.5127
R2606 vdd.n1920 vdd.n859 99.5127
R2607 vdd.n1920 vdd.n852 99.5127
R2608 vdd.n1923 vdd.n852 99.5127
R2609 vdd.n1923 vdd.n846 99.5127
R2610 vdd.n1926 vdd.n846 99.5127
R2611 vdd.n1926 vdd.n841 99.5127
R2612 vdd.n1929 vdd.n841 99.5127
R2613 vdd.n1929 vdd.n835 99.5127
R2614 vdd.n1971 vdd.n835 99.5127
R2615 vdd.n1971 vdd.n828 99.5127
R2616 vdd.n1967 vdd.n828 99.5127
R2617 vdd.n1967 vdd.n822 99.5127
R2618 vdd.n1964 vdd.n822 99.5127
R2619 vdd.n1964 vdd.n817 99.5127
R2620 vdd.n1961 vdd.n817 99.5127
R2621 vdd.n1961 vdd.n812 99.5127
R2622 vdd.n1937 vdd.n812 99.5127
R2623 vdd.n1937 vdd.n807 99.5127
R2624 vdd.n1934 vdd.n807 99.5127
R2625 vdd.n1934 vdd.n800 99.5127
R2626 vdd.n800 vdd.n791 99.5127
R2627 vdd.n2194 vdd.n791 99.5127
R2628 vdd.n2195 vdd.n2194 99.5127
R2629 vdd.n2195 vdd.n783 99.5127
R2630 vdd.n1832 vdd.n1830 99.5127
R2631 vdd.n1836 vdd.n1827 99.5127
R2632 vdd.n1840 vdd.n1838 99.5127
R2633 vdd.n1844 vdd.n1825 99.5127
R2634 vdd.n1848 vdd.n1846 99.5127
R2635 vdd.n1852 vdd.n1823 99.5127
R2636 vdd.n1856 vdd.n1854 99.5127
R2637 vdd.n1860 vdd.n1821 99.5127
R2638 vdd.n1864 vdd.n1862 99.5127
R2639 vdd.n1868 vdd.n933 99.5127
R2640 vdd.n1872 vdd.n1870 99.5127
R2641 vdd.n1876 vdd.n931 99.5127
R2642 vdd.n1880 vdd.n1878 99.5127
R2643 vdd.n1884 vdd.n929 99.5127
R2644 vdd.n1888 vdd.n1886 99.5127
R2645 vdd.n1893 vdd.n925 99.5127
R2646 vdd.n1896 vdd.n1895 99.5127
R2647 vdd.n2082 vdd.n897 99.5127
R2648 vdd.n2086 vdd.n897 99.5127
R2649 vdd.n2086 vdd.n887 99.5127
R2650 vdd.n2094 vdd.n887 99.5127
R2651 vdd.n2094 vdd.n885 99.5127
R2652 vdd.n2098 vdd.n885 99.5127
R2653 vdd.n2098 vdd.n875 99.5127
R2654 vdd.n2106 vdd.n875 99.5127
R2655 vdd.n2106 vdd.n873 99.5127
R2656 vdd.n2110 vdd.n873 99.5127
R2657 vdd.n2110 vdd.n863 99.5127
R2658 vdd.n2118 vdd.n863 99.5127
R2659 vdd.n2118 vdd.n861 99.5127
R2660 vdd.n2122 vdd.n861 99.5127
R2661 vdd.n2122 vdd.n850 99.5127
R2662 vdd.n2130 vdd.n850 99.5127
R2663 vdd.n2130 vdd.n847 99.5127
R2664 vdd.n2135 vdd.n847 99.5127
R2665 vdd.n2135 vdd.n838 99.5127
R2666 vdd.n2143 vdd.n838 99.5127
R2667 vdd.n2143 vdd.n836 99.5127
R2668 vdd.n2147 vdd.n836 99.5127
R2669 vdd.n2147 vdd.n826 99.5127
R2670 vdd.n2155 vdd.n826 99.5127
R2671 vdd.n2155 vdd.n824 99.5127
R2672 vdd.n2159 vdd.n824 99.5127
R2673 vdd.n2159 vdd.n815 99.5127
R2674 vdd.n2167 vdd.n815 99.5127
R2675 vdd.n2167 vdd.n813 99.5127
R2676 vdd.n2171 vdd.n813 99.5127
R2677 vdd.n2171 vdd.n804 99.5127
R2678 vdd.n2179 vdd.n804 99.5127
R2679 vdd.n2179 vdd.n801 99.5127
R2680 vdd.n2185 vdd.n801 99.5127
R2681 vdd.n2185 vdd.n802 99.5127
R2682 vdd.n802 vdd.n793 99.5127
R2683 vdd.n793 vdd.n784 99.5127
R2684 vdd.n2267 vdd.n784 99.5127
R2685 vdd.n9 vdd.n7 98.9633
R2686 vdd.n2 vdd.n0 98.9633
R2687 vdd.n9 vdd.n8 98.6055
R2688 vdd.n11 vdd.n10 98.6055
R2689 vdd.n13 vdd.n12 98.6055
R2690 vdd.n6 vdd.n5 98.6055
R2691 vdd.n4 vdd.n3 98.6055
R2692 vdd.n2 vdd.n1 98.6055
R2693 vdd.t9 vdd.n267 85.8723
R2694 vdd.t3 vdd.n220 85.8723
R2695 vdd.t146 vdd.n177 85.8723
R2696 vdd.t14 vdd.n130 85.8723
R2697 vdd.t23 vdd.n88 85.8723
R2698 vdd.t108 vdd.n41 85.8723
R2699 vdd.t16 vdd.n1162 85.8723
R2700 vdd.t122 vdd.n1209 85.8723
R2701 vdd.t112 vdd.n1072 85.8723
R2702 vdd.t201 vdd.n1119 85.8723
R2703 vdd.t203 vdd.n983 85.8723
R2704 vdd.t144 vdd.n1030 85.8723
R2705 vdd.n2694 vdd.n675 78.546
R2706 vdd.n2133 vdd.n848 78.546
R2707 vdd.n254 vdd.n253 75.1835
R2708 vdd.n252 vdd.n251 75.1835
R2709 vdd.n250 vdd.n249 75.1835
R2710 vdd.n164 vdd.n163 75.1835
R2711 vdd.n162 vdd.n161 75.1835
R2712 vdd.n160 vdd.n159 75.1835
R2713 vdd.n75 vdd.n74 75.1835
R2714 vdd.n73 vdd.n72 75.1835
R2715 vdd.n71 vdd.n70 75.1835
R2716 vdd.n1192 vdd.n1191 75.1835
R2717 vdd.n1194 vdd.n1193 75.1835
R2718 vdd.n1196 vdd.n1195 75.1835
R2719 vdd.n1102 vdd.n1101 75.1835
R2720 vdd.n1104 vdd.n1103 75.1835
R2721 vdd.n1106 vdd.n1105 75.1835
R2722 vdd.n1013 vdd.n1012 75.1835
R2723 vdd.n1015 vdd.n1014 75.1835
R2724 vdd.n1017 vdd.n1016 75.1835
R2725 vdd.n2624 vdd.n2357 72.8958
R2726 vdd.n2624 vdd.n2358 72.8958
R2727 vdd.n2624 vdd.n2359 72.8958
R2728 vdd.n2624 vdd.n2360 72.8958
R2729 vdd.n2624 vdd.n2361 72.8958
R2730 vdd.n2624 vdd.n2362 72.8958
R2731 vdd.n2624 vdd.n2363 72.8958
R2732 vdd.n2624 vdd.n2364 72.8958
R2733 vdd.n2624 vdd.n2365 72.8958
R2734 vdd.n2624 vdd.n2366 72.8958
R2735 vdd.n2624 vdd.n2367 72.8958
R2736 vdd.n2624 vdd.n2368 72.8958
R2737 vdd.n2624 vdd.n2369 72.8958
R2738 vdd.n2624 vdd.n2370 72.8958
R2739 vdd.n2624 vdd.n2371 72.8958
R2740 vdd.n2624 vdd.n2372 72.8958
R2741 vdd.n2624 vdd.n2373 72.8958
R2742 vdd.n593 vdd.n484 72.8958
R2743 vdd.n2862 vdd.n484 72.8958
R2744 vdd.n587 vdd.n484 72.8958
R2745 vdd.n2869 vdd.n484 72.8958
R2746 vdd.n584 vdd.n484 72.8958
R2747 vdd.n2876 vdd.n484 72.8958
R2748 vdd.n581 vdd.n484 72.8958
R2749 vdd.n2883 vdd.n484 72.8958
R2750 vdd.n2886 vdd.n484 72.8958
R2751 vdd.n2742 vdd.n484 72.8958
R2752 vdd.n2747 vdd.n484 72.8958
R2753 vdd.n2741 vdd.n484 72.8958
R2754 vdd.n2754 vdd.n484 72.8958
R2755 vdd.n2738 vdd.n484 72.8958
R2756 vdd.n2761 vdd.n484 72.8958
R2757 vdd.n2735 vdd.n484 72.8958
R2758 vdd.n2768 vdd.n484 72.8958
R2759 vdd.n2075 vdd.n900 72.8958
R2760 vdd.n905 vdd.n900 72.8958
R2761 vdd.n2068 vdd.n900 72.8958
R2762 vdd.n2062 vdd.n900 72.8958
R2763 vdd.n2060 vdd.n900 72.8958
R2764 vdd.n2054 vdd.n900 72.8958
R2765 vdd.n2052 vdd.n900 72.8958
R2766 vdd.n2046 vdd.n900 72.8958
R2767 vdd.n2044 vdd.n900 72.8958
R2768 vdd.n2038 vdd.n900 72.8958
R2769 vdd.n2036 vdd.n900 72.8958
R2770 vdd.n2030 vdd.n900 72.8958
R2771 vdd.n2028 vdd.n900 72.8958
R2772 vdd.n2022 vdd.n900 72.8958
R2773 vdd.n2020 vdd.n900 72.8958
R2774 vdd.n2013 vdd.n900 72.8958
R2775 vdd.n2011 vdd.n900 72.8958
R2776 vdd.n2340 vdd.n758 72.8958
R2777 vdd.n2340 vdd.n759 72.8958
R2778 vdd.n2340 vdd.n760 72.8958
R2779 vdd.n2340 vdd.n761 72.8958
R2780 vdd.n2340 vdd.n762 72.8958
R2781 vdd.n2340 vdd.n763 72.8958
R2782 vdd.n2340 vdd.n764 72.8958
R2783 vdd.n2340 vdd.n765 72.8958
R2784 vdd.n2340 vdd.n766 72.8958
R2785 vdd.n2340 vdd.n767 72.8958
R2786 vdd.n2340 vdd.n768 72.8958
R2787 vdd.n2340 vdd.n769 72.8958
R2788 vdd.n2340 vdd.n770 72.8958
R2789 vdd.n2340 vdd.n771 72.8958
R2790 vdd.n2340 vdd.n772 72.8958
R2791 vdd.n2340 vdd.n773 72.8958
R2792 vdd.n2340 vdd.n774 72.8958
R2793 vdd.n2625 vdd.n2624 72.8958
R2794 vdd.n2624 vdd.n2341 72.8958
R2795 vdd.n2624 vdd.n2342 72.8958
R2796 vdd.n2624 vdd.n2343 72.8958
R2797 vdd.n2624 vdd.n2344 72.8958
R2798 vdd.n2624 vdd.n2345 72.8958
R2799 vdd.n2624 vdd.n2346 72.8958
R2800 vdd.n2624 vdd.n2347 72.8958
R2801 vdd.n2624 vdd.n2348 72.8958
R2802 vdd.n2624 vdd.n2349 72.8958
R2803 vdd.n2624 vdd.n2350 72.8958
R2804 vdd.n2624 vdd.n2351 72.8958
R2805 vdd.n2624 vdd.n2352 72.8958
R2806 vdd.n2624 vdd.n2353 72.8958
R2807 vdd.n2624 vdd.n2354 72.8958
R2808 vdd.n2624 vdd.n2355 72.8958
R2809 vdd.n2624 vdd.n2356 72.8958
R2810 vdd.n2792 vdd.n484 72.8958
R2811 vdd.n625 vdd.n484 72.8958
R2812 vdd.n2800 vdd.n484 72.8958
R2813 vdd.n620 vdd.n484 72.8958
R2814 vdd.n2807 vdd.n484 72.8958
R2815 vdd.n617 vdd.n484 72.8958
R2816 vdd.n2814 vdd.n484 72.8958
R2817 vdd.n614 vdd.n484 72.8958
R2818 vdd.n2821 vdd.n484 72.8958
R2819 vdd.n2825 vdd.n484 72.8958
R2820 vdd.n611 vdd.n484 72.8958
R2821 vdd.n2832 vdd.n484 72.8958
R2822 vdd.n608 vdd.n484 72.8958
R2823 vdd.n2839 vdd.n484 72.8958
R2824 vdd.n605 vdd.n484 72.8958
R2825 vdd.n2846 vdd.n484 72.8958
R2826 vdd.n2849 vdd.n484 72.8958
R2827 vdd.n2340 vdd.n756 72.8958
R2828 vdd.n2340 vdd.n755 72.8958
R2829 vdd.n2340 vdd.n754 72.8958
R2830 vdd.n2340 vdd.n753 72.8958
R2831 vdd.n2340 vdd.n752 72.8958
R2832 vdd.n2340 vdd.n751 72.8958
R2833 vdd.n2340 vdd.n750 72.8958
R2834 vdd.n2340 vdd.n749 72.8958
R2835 vdd.n2340 vdd.n748 72.8958
R2836 vdd.n2340 vdd.n747 72.8958
R2837 vdd.n2340 vdd.n746 72.8958
R2838 vdd.n2340 vdd.n745 72.8958
R2839 vdd.n2340 vdd.n744 72.8958
R2840 vdd.n2340 vdd.n743 72.8958
R2841 vdd.n2340 vdd.n742 72.8958
R2842 vdd.n2340 vdd.n741 72.8958
R2843 vdd.n2340 vdd.n740 72.8958
R2844 vdd.n1829 vdd.n900 72.8958
R2845 vdd.n1831 vdd.n900 72.8958
R2846 vdd.n1837 vdd.n900 72.8958
R2847 vdd.n1839 vdd.n900 72.8958
R2848 vdd.n1845 vdd.n900 72.8958
R2849 vdd.n1847 vdd.n900 72.8958
R2850 vdd.n1853 vdd.n900 72.8958
R2851 vdd.n1855 vdd.n900 72.8958
R2852 vdd.n1861 vdd.n900 72.8958
R2853 vdd.n1863 vdd.n900 72.8958
R2854 vdd.n1869 vdd.n900 72.8958
R2855 vdd.n1871 vdd.n900 72.8958
R2856 vdd.n1877 vdd.n900 72.8958
R2857 vdd.n1879 vdd.n900 72.8958
R2858 vdd.n1885 vdd.n900 72.8958
R2859 vdd.n1887 vdd.n900 72.8958
R2860 vdd.n1894 vdd.n900 72.8958
R2861 vdd.n1502 vdd.n1501 66.2847
R2862 vdd.n1501 vdd.n1277 66.2847
R2863 vdd.n1501 vdd.n1278 66.2847
R2864 vdd.n1501 vdd.n1279 66.2847
R2865 vdd.n1501 vdd.n1280 66.2847
R2866 vdd.n1501 vdd.n1281 66.2847
R2867 vdd.n1501 vdd.n1282 66.2847
R2868 vdd.n1501 vdd.n1283 66.2847
R2869 vdd.n1501 vdd.n1284 66.2847
R2870 vdd.n1501 vdd.n1285 66.2847
R2871 vdd.n1501 vdd.n1286 66.2847
R2872 vdd.n1501 vdd.n1287 66.2847
R2873 vdd.n1501 vdd.n1288 66.2847
R2874 vdd.n1501 vdd.n1289 66.2847
R2875 vdd.n1501 vdd.n1290 66.2847
R2876 vdd.n1501 vdd.n1291 66.2847
R2877 vdd.n1501 vdd.n1292 66.2847
R2878 vdd.n1501 vdd.n1293 66.2847
R2879 vdd.n1501 vdd.n1294 66.2847
R2880 vdd.n1501 vdd.n1295 66.2847
R2881 vdd.n1501 vdd.n1296 66.2847
R2882 vdd.n1501 vdd.n1297 66.2847
R2883 vdd.n1501 vdd.n1298 66.2847
R2884 vdd.n1501 vdd.n1299 66.2847
R2885 vdd.n1501 vdd.n1300 66.2847
R2886 vdd.n1501 vdd.n1301 66.2847
R2887 vdd.n1501 vdd.n1302 66.2847
R2888 vdd.n1501 vdd.n1303 66.2847
R2889 vdd.n1501 vdd.n1304 66.2847
R2890 vdd.n1501 vdd.n1305 66.2847
R2891 vdd.n1501 vdd.n1306 66.2847
R2892 vdd.n943 vdd.n940 66.2847
R2893 vdd.n1694 vdd.n943 66.2847
R2894 vdd.n1699 vdd.n943 66.2847
R2895 vdd.n1704 vdd.n943 66.2847
R2896 vdd.n1692 vdd.n943 66.2847
R2897 vdd.n1711 vdd.n943 66.2847
R2898 vdd.n1684 vdd.n943 66.2847
R2899 vdd.n1718 vdd.n943 66.2847
R2900 vdd.n1677 vdd.n943 66.2847
R2901 vdd.n1725 vdd.n943 66.2847
R2902 vdd.n1671 vdd.n943 66.2847
R2903 vdd.n1666 vdd.n943 66.2847
R2904 vdd.n1736 vdd.n943 66.2847
R2905 vdd.n1658 vdd.n943 66.2847
R2906 vdd.n1743 vdd.n943 66.2847
R2907 vdd.n1651 vdd.n943 66.2847
R2908 vdd.n1750 vdd.n943 66.2847
R2909 vdd.n1644 vdd.n943 66.2847
R2910 vdd.n1757 vdd.n943 66.2847
R2911 vdd.n1637 vdd.n943 66.2847
R2912 vdd.n1764 vdd.n943 66.2847
R2913 vdd.n1631 vdd.n943 66.2847
R2914 vdd.n1626 vdd.n943 66.2847
R2915 vdd.n1775 vdd.n943 66.2847
R2916 vdd.n1618 vdd.n943 66.2847
R2917 vdd.n1782 vdd.n943 66.2847
R2918 vdd.n1611 vdd.n943 66.2847
R2919 vdd.n1789 vdd.n943 66.2847
R2920 vdd.n1792 vdd.n943 66.2847
R2921 vdd.n1602 vdd.n943 66.2847
R2922 vdd.n1801 vdd.n943 66.2847
R2923 vdd.n1596 vdd.n943 66.2847
R2924 vdd.n3023 vdd.n3022 66.2847
R2925 vdd.n3022 vdd.n485 66.2847
R2926 vdd.n3022 vdd.n486 66.2847
R2927 vdd.n3022 vdd.n487 66.2847
R2928 vdd.n3022 vdd.n488 66.2847
R2929 vdd.n3022 vdd.n489 66.2847
R2930 vdd.n3022 vdd.n490 66.2847
R2931 vdd.n3022 vdd.n491 66.2847
R2932 vdd.n3022 vdd.n492 66.2847
R2933 vdd.n3022 vdd.n493 66.2847
R2934 vdd.n3022 vdd.n494 66.2847
R2935 vdd.n3022 vdd.n495 66.2847
R2936 vdd.n3022 vdd.n496 66.2847
R2937 vdd.n3022 vdd.n497 66.2847
R2938 vdd.n3022 vdd.n498 66.2847
R2939 vdd.n3022 vdd.n499 66.2847
R2940 vdd.n3022 vdd.n500 66.2847
R2941 vdd.n3022 vdd.n501 66.2847
R2942 vdd.n3022 vdd.n502 66.2847
R2943 vdd.n3022 vdd.n503 66.2847
R2944 vdd.n3022 vdd.n504 66.2847
R2945 vdd.n3022 vdd.n505 66.2847
R2946 vdd.n3022 vdd.n506 66.2847
R2947 vdd.n3022 vdd.n507 66.2847
R2948 vdd.n3022 vdd.n508 66.2847
R2949 vdd.n3022 vdd.n509 66.2847
R2950 vdd.n3022 vdd.n510 66.2847
R2951 vdd.n3022 vdd.n511 66.2847
R2952 vdd.n3022 vdd.n512 66.2847
R2953 vdd.n3022 vdd.n513 66.2847
R2954 vdd.n3022 vdd.n514 66.2847
R2955 vdd.n3087 vdd.n329 66.2847
R2956 vdd.n3096 vdd.n329 66.2847
R2957 vdd.n439 vdd.n329 66.2847
R2958 vdd.n3103 vdd.n329 66.2847
R2959 vdd.n432 vdd.n329 66.2847
R2960 vdd.n3110 vdd.n329 66.2847
R2961 vdd.n425 vdd.n329 66.2847
R2962 vdd.n3117 vdd.n329 66.2847
R2963 vdd.n418 vdd.n329 66.2847
R2964 vdd.n3124 vdd.n329 66.2847
R2965 vdd.n412 vdd.n329 66.2847
R2966 vdd.n407 vdd.n329 66.2847
R2967 vdd.n3135 vdd.n329 66.2847
R2968 vdd.n399 vdd.n329 66.2847
R2969 vdd.n3142 vdd.n329 66.2847
R2970 vdd.n392 vdd.n329 66.2847
R2971 vdd.n3149 vdd.n329 66.2847
R2972 vdd.n385 vdd.n329 66.2847
R2973 vdd.n3156 vdd.n329 66.2847
R2974 vdd.n378 vdd.n329 66.2847
R2975 vdd.n3163 vdd.n329 66.2847
R2976 vdd.n372 vdd.n329 66.2847
R2977 vdd.n367 vdd.n329 66.2847
R2978 vdd.n3174 vdd.n329 66.2847
R2979 vdd.n359 vdd.n329 66.2847
R2980 vdd.n3181 vdd.n329 66.2847
R2981 vdd.n352 vdd.n329 66.2847
R2982 vdd.n3188 vdd.n329 66.2847
R2983 vdd.n345 vdd.n329 66.2847
R2984 vdd.n3195 vdd.n329 66.2847
R2985 vdd.n3198 vdd.n329 66.2847
R2986 vdd.n333 vdd.n329 66.2847
R2987 vdd.n334 vdd.n333 52.4337
R2988 vdd.n3198 vdd.n3197 52.4337
R2989 vdd.n3195 vdd.n3194 52.4337
R2990 vdd.n3190 vdd.n345 52.4337
R2991 vdd.n3188 vdd.n3187 52.4337
R2992 vdd.n3183 vdd.n352 52.4337
R2993 vdd.n3181 vdd.n3180 52.4337
R2994 vdd.n3176 vdd.n359 52.4337
R2995 vdd.n3174 vdd.n3173 52.4337
R2996 vdd.n368 vdd.n367 52.4337
R2997 vdd.n3165 vdd.n372 52.4337
R2998 vdd.n3163 vdd.n3162 52.4337
R2999 vdd.n3158 vdd.n378 52.4337
R3000 vdd.n3156 vdd.n3155 52.4337
R3001 vdd.n3151 vdd.n385 52.4337
R3002 vdd.n3149 vdd.n3148 52.4337
R3003 vdd.n3144 vdd.n392 52.4337
R3004 vdd.n3142 vdd.n3141 52.4337
R3005 vdd.n3137 vdd.n399 52.4337
R3006 vdd.n3135 vdd.n3134 52.4337
R3007 vdd.n408 vdd.n407 52.4337
R3008 vdd.n3126 vdd.n412 52.4337
R3009 vdd.n3124 vdd.n3123 52.4337
R3010 vdd.n3119 vdd.n418 52.4337
R3011 vdd.n3117 vdd.n3116 52.4337
R3012 vdd.n3112 vdd.n425 52.4337
R3013 vdd.n3110 vdd.n3109 52.4337
R3014 vdd.n3105 vdd.n432 52.4337
R3015 vdd.n3103 vdd.n3102 52.4337
R3016 vdd.n3098 vdd.n439 52.4337
R3017 vdd.n3096 vdd.n3095 52.4337
R3018 vdd.n3088 vdd.n3087 52.4337
R3019 vdd.n3024 vdd.n3023 52.4337
R3020 vdd.n517 vdd.n485 52.4337
R3021 vdd.n523 vdd.n486 52.4337
R3022 vdd.n3013 vdd.n487 52.4337
R3023 vdd.n3009 vdd.n488 52.4337
R3024 vdd.n3005 vdd.n489 52.4337
R3025 vdd.n3001 vdd.n490 52.4337
R3026 vdd.n2997 vdd.n491 52.4337
R3027 vdd.n2993 vdd.n492 52.4337
R3028 vdd.n2989 vdd.n493 52.4337
R3029 vdd.n2981 vdd.n494 52.4337
R3030 vdd.n2977 vdd.n495 52.4337
R3031 vdd.n2973 vdd.n496 52.4337
R3032 vdd.n2969 vdd.n497 52.4337
R3033 vdd.n2965 vdd.n498 52.4337
R3034 vdd.n2961 vdd.n499 52.4337
R3035 vdd.n2957 vdd.n500 52.4337
R3036 vdd.n2953 vdd.n501 52.4337
R3037 vdd.n2949 vdd.n502 52.4337
R3038 vdd.n2945 vdd.n503 52.4337
R3039 vdd.n2941 vdd.n504 52.4337
R3040 vdd.n2935 vdd.n505 52.4337
R3041 vdd.n2931 vdd.n506 52.4337
R3042 vdd.n2927 vdd.n507 52.4337
R3043 vdd.n2923 vdd.n508 52.4337
R3044 vdd.n2919 vdd.n509 52.4337
R3045 vdd.n2915 vdd.n510 52.4337
R3046 vdd.n2911 vdd.n511 52.4337
R3047 vdd.n2907 vdd.n512 52.4337
R3048 vdd.n2903 vdd.n513 52.4337
R3049 vdd.n2899 vdd.n514 52.4337
R3050 vdd.n1803 vdd.n1596 52.4337
R3051 vdd.n1801 vdd.n1800 52.4337
R3052 vdd.n1603 vdd.n1602 52.4337
R3053 vdd.n1792 vdd.n1791 52.4337
R3054 vdd.n1789 vdd.n1788 52.4337
R3055 vdd.n1784 vdd.n1611 52.4337
R3056 vdd.n1782 vdd.n1781 52.4337
R3057 vdd.n1777 vdd.n1618 52.4337
R3058 vdd.n1775 vdd.n1774 52.4337
R3059 vdd.n1627 vdd.n1626 52.4337
R3060 vdd.n1766 vdd.n1631 52.4337
R3061 vdd.n1764 vdd.n1763 52.4337
R3062 vdd.n1759 vdd.n1637 52.4337
R3063 vdd.n1757 vdd.n1756 52.4337
R3064 vdd.n1752 vdd.n1644 52.4337
R3065 vdd.n1750 vdd.n1749 52.4337
R3066 vdd.n1745 vdd.n1651 52.4337
R3067 vdd.n1743 vdd.n1742 52.4337
R3068 vdd.n1738 vdd.n1658 52.4337
R3069 vdd.n1736 vdd.n1735 52.4337
R3070 vdd.n1667 vdd.n1666 52.4337
R3071 vdd.n1727 vdd.n1671 52.4337
R3072 vdd.n1725 vdd.n1724 52.4337
R3073 vdd.n1720 vdd.n1677 52.4337
R3074 vdd.n1718 vdd.n1717 52.4337
R3075 vdd.n1713 vdd.n1684 52.4337
R3076 vdd.n1711 vdd.n1710 52.4337
R3077 vdd.n1706 vdd.n1692 52.4337
R3078 vdd.n1704 vdd.n1703 52.4337
R3079 vdd.n1699 vdd.n1698 52.4337
R3080 vdd.n1694 vdd.n1693 52.4337
R3081 vdd.n1812 vdd.n940 52.4337
R3082 vdd.n1503 vdd.n1502 52.4337
R3083 vdd.n1309 vdd.n1277 52.4337
R3084 vdd.n1313 vdd.n1278 52.4337
R3085 vdd.n1315 vdd.n1279 52.4337
R3086 vdd.n1319 vdd.n1280 52.4337
R3087 vdd.n1321 vdd.n1281 52.4337
R3088 vdd.n1325 vdd.n1282 52.4337
R3089 vdd.n1327 vdd.n1283 52.4337
R3090 vdd.n1331 vdd.n1284 52.4337
R3091 vdd.n1333 vdd.n1285 52.4337
R3092 vdd.n1339 vdd.n1286 52.4337
R3093 vdd.n1341 vdd.n1287 52.4337
R3094 vdd.n1345 vdd.n1288 52.4337
R3095 vdd.n1347 vdd.n1289 52.4337
R3096 vdd.n1351 vdd.n1290 52.4337
R3097 vdd.n1353 vdd.n1291 52.4337
R3098 vdd.n1357 vdd.n1292 52.4337
R3099 vdd.n1359 vdd.n1293 52.4337
R3100 vdd.n1363 vdd.n1294 52.4337
R3101 vdd.n1365 vdd.n1295 52.4337
R3102 vdd.n1437 vdd.n1296 52.4337
R3103 vdd.n1370 vdd.n1297 52.4337
R3104 vdd.n1374 vdd.n1298 52.4337
R3105 vdd.n1376 vdd.n1299 52.4337
R3106 vdd.n1380 vdd.n1300 52.4337
R3107 vdd.n1382 vdd.n1301 52.4337
R3108 vdd.n1386 vdd.n1302 52.4337
R3109 vdd.n1388 vdd.n1303 52.4337
R3110 vdd.n1392 vdd.n1304 52.4337
R3111 vdd.n1394 vdd.n1305 52.4337
R3112 vdd.n1398 vdd.n1306 52.4337
R3113 vdd.n1502 vdd.n1276 52.4337
R3114 vdd.n1312 vdd.n1277 52.4337
R3115 vdd.n1314 vdd.n1278 52.4337
R3116 vdd.n1318 vdd.n1279 52.4337
R3117 vdd.n1320 vdd.n1280 52.4337
R3118 vdd.n1324 vdd.n1281 52.4337
R3119 vdd.n1326 vdd.n1282 52.4337
R3120 vdd.n1330 vdd.n1283 52.4337
R3121 vdd.n1332 vdd.n1284 52.4337
R3122 vdd.n1338 vdd.n1285 52.4337
R3123 vdd.n1340 vdd.n1286 52.4337
R3124 vdd.n1344 vdd.n1287 52.4337
R3125 vdd.n1346 vdd.n1288 52.4337
R3126 vdd.n1350 vdd.n1289 52.4337
R3127 vdd.n1352 vdd.n1290 52.4337
R3128 vdd.n1356 vdd.n1291 52.4337
R3129 vdd.n1358 vdd.n1292 52.4337
R3130 vdd.n1362 vdd.n1293 52.4337
R3131 vdd.n1364 vdd.n1294 52.4337
R3132 vdd.n1368 vdd.n1295 52.4337
R3133 vdd.n1369 vdd.n1296 52.4337
R3134 vdd.n1373 vdd.n1297 52.4337
R3135 vdd.n1375 vdd.n1298 52.4337
R3136 vdd.n1379 vdd.n1299 52.4337
R3137 vdd.n1381 vdd.n1300 52.4337
R3138 vdd.n1385 vdd.n1301 52.4337
R3139 vdd.n1387 vdd.n1302 52.4337
R3140 vdd.n1391 vdd.n1303 52.4337
R3141 vdd.n1393 vdd.n1304 52.4337
R3142 vdd.n1397 vdd.n1305 52.4337
R3143 vdd.n1399 vdd.n1306 52.4337
R3144 vdd.n940 vdd.n939 52.4337
R3145 vdd.n1695 vdd.n1694 52.4337
R3146 vdd.n1700 vdd.n1699 52.4337
R3147 vdd.n1705 vdd.n1704 52.4337
R3148 vdd.n1692 vdd.n1685 52.4337
R3149 vdd.n1712 vdd.n1711 52.4337
R3150 vdd.n1684 vdd.n1678 52.4337
R3151 vdd.n1719 vdd.n1718 52.4337
R3152 vdd.n1677 vdd.n1672 52.4337
R3153 vdd.n1726 vdd.n1725 52.4337
R3154 vdd.n1671 vdd.n1670 52.4337
R3155 vdd.n1666 vdd.n1659 52.4337
R3156 vdd.n1737 vdd.n1736 52.4337
R3157 vdd.n1658 vdd.n1652 52.4337
R3158 vdd.n1744 vdd.n1743 52.4337
R3159 vdd.n1651 vdd.n1645 52.4337
R3160 vdd.n1751 vdd.n1750 52.4337
R3161 vdd.n1644 vdd.n1638 52.4337
R3162 vdd.n1758 vdd.n1757 52.4337
R3163 vdd.n1637 vdd.n1632 52.4337
R3164 vdd.n1765 vdd.n1764 52.4337
R3165 vdd.n1631 vdd.n1630 52.4337
R3166 vdd.n1626 vdd.n1619 52.4337
R3167 vdd.n1776 vdd.n1775 52.4337
R3168 vdd.n1618 vdd.n1612 52.4337
R3169 vdd.n1783 vdd.n1782 52.4337
R3170 vdd.n1611 vdd.n1605 52.4337
R3171 vdd.n1790 vdd.n1789 52.4337
R3172 vdd.n1793 vdd.n1792 52.4337
R3173 vdd.n1602 vdd.n1597 52.4337
R3174 vdd.n1802 vdd.n1801 52.4337
R3175 vdd.n1596 vdd.n945 52.4337
R3176 vdd.n3023 vdd.n483 52.4337
R3177 vdd.n522 vdd.n485 52.4337
R3178 vdd.n3014 vdd.n486 52.4337
R3179 vdd.n3010 vdd.n487 52.4337
R3180 vdd.n3006 vdd.n488 52.4337
R3181 vdd.n3002 vdd.n489 52.4337
R3182 vdd.n2998 vdd.n490 52.4337
R3183 vdd.n2994 vdd.n491 52.4337
R3184 vdd.n2990 vdd.n492 52.4337
R3185 vdd.n2980 vdd.n493 52.4337
R3186 vdd.n2978 vdd.n494 52.4337
R3187 vdd.n2974 vdd.n495 52.4337
R3188 vdd.n2970 vdd.n496 52.4337
R3189 vdd.n2966 vdd.n497 52.4337
R3190 vdd.n2962 vdd.n498 52.4337
R3191 vdd.n2958 vdd.n499 52.4337
R3192 vdd.n2954 vdd.n500 52.4337
R3193 vdd.n2950 vdd.n501 52.4337
R3194 vdd.n2946 vdd.n502 52.4337
R3195 vdd.n2942 vdd.n503 52.4337
R3196 vdd.n2934 vdd.n504 52.4337
R3197 vdd.n2932 vdd.n505 52.4337
R3198 vdd.n2928 vdd.n506 52.4337
R3199 vdd.n2924 vdd.n507 52.4337
R3200 vdd.n2920 vdd.n508 52.4337
R3201 vdd.n2916 vdd.n509 52.4337
R3202 vdd.n2912 vdd.n510 52.4337
R3203 vdd.n2908 vdd.n511 52.4337
R3204 vdd.n2904 vdd.n512 52.4337
R3205 vdd.n2900 vdd.n513 52.4337
R3206 vdd.n2896 vdd.n514 52.4337
R3207 vdd.n3087 vdd.n440 52.4337
R3208 vdd.n3097 vdd.n3096 52.4337
R3209 vdd.n439 vdd.n433 52.4337
R3210 vdd.n3104 vdd.n3103 52.4337
R3211 vdd.n432 vdd.n426 52.4337
R3212 vdd.n3111 vdd.n3110 52.4337
R3213 vdd.n425 vdd.n419 52.4337
R3214 vdd.n3118 vdd.n3117 52.4337
R3215 vdd.n418 vdd.n413 52.4337
R3216 vdd.n3125 vdd.n3124 52.4337
R3217 vdd.n412 vdd.n411 52.4337
R3218 vdd.n407 vdd.n400 52.4337
R3219 vdd.n3136 vdd.n3135 52.4337
R3220 vdd.n399 vdd.n393 52.4337
R3221 vdd.n3143 vdd.n3142 52.4337
R3222 vdd.n392 vdd.n386 52.4337
R3223 vdd.n3150 vdd.n3149 52.4337
R3224 vdd.n385 vdd.n379 52.4337
R3225 vdd.n3157 vdd.n3156 52.4337
R3226 vdd.n378 vdd.n373 52.4337
R3227 vdd.n3164 vdd.n3163 52.4337
R3228 vdd.n372 vdd.n371 52.4337
R3229 vdd.n367 vdd.n360 52.4337
R3230 vdd.n3175 vdd.n3174 52.4337
R3231 vdd.n359 vdd.n353 52.4337
R3232 vdd.n3182 vdd.n3181 52.4337
R3233 vdd.n352 vdd.n346 52.4337
R3234 vdd.n3189 vdd.n3188 52.4337
R3235 vdd.n345 vdd.n338 52.4337
R3236 vdd.n3196 vdd.n3195 52.4337
R3237 vdd.n3199 vdd.n3198 52.4337
R3238 vdd.n333 vdd.n330 52.4337
R3239 vdd.t162 vdd.t172 51.4683
R3240 vdd.n250 vdd.n248 42.0461
R3241 vdd.n160 vdd.n158 42.0461
R3242 vdd.n71 vdd.n69 42.0461
R3243 vdd.n1192 vdd.n1190 42.0461
R3244 vdd.n1102 vdd.n1100 42.0461
R3245 vdd.n1013 vdd.n1011 42.0461
R3246 vdd.n296 vdd.n295 41.6884
R3247 vdd.n206 vdd.n205 41.6884
R3248 vdd.n117 vdd.n116 41.6884
R3249 vdd.n1238 vdd.n1237 41.6884
R3250 vdd.n1148 vdd.n1147 41.6884
R3251 vdd.n1059 vdd.n1058 41.6884
R3252 vdd.n1402 vdd.n1401 41.1157
R3253 vdd.n1440 vdd.n1439 41.1157
R3254 vdd.n1336 vdd.n1335 41.1157
R3255 vdd.n3092 vdd.n3091 41.1157
R3256 vdd.n3131 vdd.n406 41.1157
R3257 vdd.n3170 vdd.n366 41.1157
R3258 vdd.n2849 vdd.n2848 39.2114
R3259 vdd.n2846 vdd.n2845 39.2114
R3260 vdd.n2841 vdd.n605 39.2114
R3261 vdd.n2839 vdd.n2838 39.2114
R3262 vdd.n2834 vdd.n608 39.2114
R3263 vdd.n2832 vdd.n2831 39.2114
R3264 vdd.n2827 vdd.n611 39.2114
R3265 vdd.n2825 vdd.n2824 39.2114
R3266 vdd.n2821 vdd.n2820 39.2114
R3267 vdd.n2816 vdd.n614 39.2114
R3268 vdd.n2814 vdd.n2813 39.2114
R3269 vdd.n2809 vdd.n617 39.2114
R3270 vdd.n2807 vdd.n2806 39.2114
R3271 vdd.n2802 vdd.n620 39.2114
R3272 vdd.n2800 vdd.n2799 39.2114
R3273 vdd.n2794 vdd.n625 39.2114
R3274 vdd.n2792 vdd.n2791 39.2114
R3275 vdd.n2625 vdd.n737 39.2114
R3276 vdd.n2446 vdd.n2341 39.2114
R3277 vdd.n2450 vdd.n2342 39.2114
R3278 vdd.n2454 vdd.n2343 39.2114
R3279 vdd.n2458 vdd.n2344 39.2114
R3280 vdd.n2462 vdd.n2345 39.2114
R3281 vdd.n2466 vdd.n2346 39.2114
R3282 vdd.n2470 vdd.n2347 39.2114
R3283 vdd.n2474 vdd.n2348 39.2114
R3284 vdd.n2478 vdd.n2349 39.2114
R3285 vdd.n2482 vdd.n2350 39.2114
R3286 vdd.n2486 vdd.n2351 39.2114
R3287 vdd.n2490 vdd.n2352 39.2114
R3288 vdd.n2494 vdd.n2353 39.2114
R3289 vdd.n2498 vdd.n2354 39.2114
R3290 vdd.n2502 vdd.n2355 39.2114
R3291 vdd.n2507 vdd.n2356 39.2114
R3292 vdd.n2335 vdd.n774 39.2114
R3293 vdd.n2331 vdd.n773 39.2114
R3294 vdd.n2327 vdd.n772 39.2114
R3295 vdd.n2323 vdd.n771 39.2114
R3296 vdd.n2319 vdd.n770 39.2114
R3297 vdd.n2315 vdd.n769 39.2114
R3298 vdd.n2311 vdd.n768 39.2114
R3299 vdd.n2307 vdd.n767 39.2114
R3300 vdd.n2303 vdd.n766 39.2114
R3301 vdd.n2299 vdd.n765 39.2114
R3302 vdd.n2295 vdd.n764 39.2114
R3303 vdd.n2291 vdd.n763 39.2114
R3304 vdd.n2287 vdd.n762 39.2114
R3305 vdd.n2283 vdd.n761 39.2114
R3306 vdd.n2279 vdd.n760 39.2114
R3307 vdd.n2274 vdd.n759 39.2114
R3308 vdd.n2270 vdd.n758 39.2114
R3309 vdd.n2075 vdd.n903 39.2114
R3310 vdd.n2073 vdd.n905 39.2114
R3311 vdd.n2069 vdd.n2068 39.2114
R3312 vdd.n2062 vdd.n907 39.2114
R3313 vdd.n2061 vdd.n2060 39.2114
R3314 vdd.n2054 vdd.n909 39.2114
R3315 vdd.n2053 vdd.n2052 39.2114
R3316 vdd.n2046 vdd.n911 39.2114
R3317 vdd.n2045 vdd.n2044 39.2114
R3318 vdd.n2038 vdd.n913 39.2114
R3319 vdd.n2037 vdd.n2036 39.2114
R3320 vdd.n2030 vdd.n915 39.2114
R3321 vdd.n2029 vdd.n2028 39.2114
R3322 vdd.n2022 vdd.n917 39.2114
R3323 vdd.n2021 vdd.n2020 39.2114
R3324 vdd.n2013 vdd.n919 39.2114
R3325 vdd.n2012 vdd.n2011 39.2114
R3326 vdd.n2768 vdd.n2767 39.2114
R3327 vdd.n2763 vdd.n2735 39.2114
R3328 vdd.n2761 vdd.n2760 39.2114
R3329 vdd.n2756 vdd.n2738 39.2114
R3330 vdd.n2754 vdd.n2753 39.2114
R3331 vdd.n2749 vdd.n2741 39.2114
R3332 vdd.n2747 vdd.n2746 39.2114
R3333 vdd.n2742 vdd.n577 39.2114
R3334 vdd.n2886 vdd.n2885 39.2114
R3335 vdd.n2883 vdd.n2882 39.2114
R3336 vdd.n2878 vdd.n581 39.2114
R3337 vdd.n2876 vdd.n2875 39.2114
R3338 vdd.n2871 vdd.n584 39.2114
R3339 vdd.n2869 vdd.n2868 39.2114
R3340 vdd.n2864 vdd.n587 39.2114
R3341 vdd.n2862 vdd.n2861 39.2114
R3342 vdd.n2857 vdd.n593 39.2114
R3343 vdd.n2357 vdd.n733 39.2114
R3344 vdd.n2380 vdd.n2358 39.2114
R3345 vdd.n2384 vdd.n2359 39.2114
R3346 vdd.n2388 vdd.n2360 39.2114
R3347 vdd.n2392 vdd.n2361 39.2114
R3348 vdd.n2396 vdd.n2362 39.2114
R3349 vdd.n2400 vdd.n2363 39.2114
R3350 vdd.n2404 vdd.n2364 39.2114
R3351 vdd.n2408 vdd.n2365 39.2114
R3352 vdd.n2412 vdd.n2366 39.2114
R3353 vdd.n2416 vdd.n2367 39.2114
R3354 vdd.n2420 vdd.n2368 39.2114
R3355 vdd.n2424 vdd.n2369 39.2114
R3356 vdd.n2428 vdd.n2370 39.2114
R3357 vdd.n2432 vdd.n2371 39.2114
R3358 vdd.n2436 vdd.n2372 39.2114
R3359 vdd.n2440 vdd.n2373 39.2114
R3360 vdd.n2379 vdd.n2357 39.2114
R3361 vdd.n2383 vdd.n2358 39.2114
R3362 vdd.n2387 vdd.n2359 39.2114
R3363 vdd.n2391 vdd.n2360 39.2114
R3364 vdd.n2395 vdd.n2361 39.2114
R3365 vdd.n2399 vdd.n2362 39.2114
R3366 vdd.n2403 vdd.n2363 39.2114
R3367 vdd.n2407 vdd.n2364 39.2114
R3368 vdd.n2411 vdd.n2365 39.2114
R3369 vdd.n2415 vdd.n2366 39.2114
R3370 vdd.n2419 vdd.n2367 39.2114
R3371 vdd.n2423 vdd.n2368 39.2114
R3372 vdd.n2427 vdd.n2369 39.2114
R3373 vdd.n2431 vdd.n2370 39.2114
R3374 vdd.n2435 vdd.n2371 39.2114
R3375 vdd.n2439 vdd.n2372 39.2114
R3376 vdd.n2374 vdd.n2373 39.2114
R3377 vdd.n593 vdd.n588 39.2114
R3378 vdd.n2863 vdd.n2862 39.2114
R3379 vdd.n587 vdd.n585 39.2114
R3380 vdd.n2870 vdd.n2869 39.2114
R3381 vdd.n584 vdd.n582 39.2114
R3382 vdd.n2877 vdd.n2876 39.2114
R3383 vdd.n581 vdd.n579 39.2114
R3384 vdd.n2884 vdd.n2883 39.2114
R3385 vdd.n2887 vdd.n2886 39.2114
R3386 vdd.n2743 vdd.n2742 39.2114
R3387 vdd.n2748 vdd.n2747 39.2114
R3388 vdd.n2741 vdd.n2739 39.2114
R3389 vdd.n2755 vdd.n2754 39.2114
R3390 vdd.n2738 vdd.n2736 39.2114
R3391 vdd.n2762 vdd.n2761 39.2114
R3392 vdd.n2735 vdd.n2733 39.2114
R3393 vdd.n2769 vdd.n2768 39.2114
R3394 vdd.n2076 vdd.n2075 39.2114
R3395 vdd.n2070 vdd.n905 39.2114
R3396 vdd.n2068 vdd.n2067 39.2114
R3397 vdd.n2063 vdd.n2062 39.2114
R3398 vdd.n2060 vdd.n2059 39.2114
R3399 vdd.n2055 vdd.n2054 39.2114
R3400 vdd.n2052 vdd.n2051 39.2114
R3401 vdd.n2047 vdd.n2046 39.2114
R3402 vdd.n2044 vdd.n2043 39.2114
R3403 vdd.n2039 vdd.n2038 39.2114
R3404 vdd.n2036 vdd.n2035 39.2114
R3405 vdd.n2031 vdd.n2030 39.2114
R3406 vdd.n2028 vdd.n2027 39.2114
R3407 vdd.n2023 vdd.n2022 39.2114
R3408 vdd.n2020 vdd.n2019 39.2114
R3409 vdd.n2014 vdd.n2013 39.2114
R3410 vdd.n2011 vdd.n2010 39.2114
R3411 vdd.n2273 vdd.n758 39.2114
R3412 vdd.n2278 vdd.n759 39.2114
R3413 vdd.n2282 vdd.n760 39.2114
R3414 vdd.n2286 vdd.n761 39.2114
R3415 vdd.n2290 vdd.n762 39.2114
R3416 vdd.n2294 vdd.n763 39.2114
R3417 vdd.n2298 vdd.n764 39.2114
R3418 vdd.n2302 vdd.n765 39.2114
R3419 vdd.n2306 vdd.n766 39.2114
R3420 vdd.n2310 vdd.n767 39.2114
R3421 vdd.n2314 vdd.n768 39.2114
R3422 vdd.n2318 vdd.n769 39.2114
R3423 vdd.n2322 vdd.n770 39.2114
R3424 vdd.n2326 vdd.n771 39.2114
R3425 vdd.n2330 vdd.n772 39.2114
R3426 vdd.n2334 vdd.n773 39.2114
R3427 vdd.n776 vdd.n774 39.2114
R3428 vdd.n2626 vdd.n2625 39.2114
R3429 vdd.n2449 vdd.n2341 39.2114
R3430 vdd.n2453 vdd.n2342 39.2114
R3431 vdd.n2457 vdd.n2343 39.2114
R3432 vdd.n2461 vdd.n2344 39.2114
R3433 vdd.n2465 vdd.n2345 39.2114
R3434 vdd.n2469 vdd.n2346 39.2114
R3435 vdd.n2473 vdd.n2347 39.2114
R3436 vdd.n2477 vdd.n2348 39.2114
R3437 vdd.n2481 vdd.n2349 39.2114
R3438 vdd.n2485 vdd.n2350 39.2114
R3439 vdd.n2489 vdd.n2351 39.2114
R3440 vdd.n2493 vdd.n2352 39.2114
R3441 vdd.n2497 vdd.n2353 39.2114
R3442 vdd.n2501 vdd.n2354 39.2114
R3443 vdd.n2506 vdd.n2355 39.2114
R3444 vdd.n2509 vdd.n2356 39.2114
R3445 vdd.n2793 vdd.n2792 39.2114
R3446 vdd.n625 vdd.n621 39.2114
R3447 vdd.n2801 vdd.n2800 39.2114
R3448 vdd.n620 vdd.n618 39.2114
R3449 vdd.n2808 vdd.n2807 39.2114
R3450 vdd.n617 vdd.n615 39.2114
R3451 vdd.n2815 vdd.n2814 39.2114
R3452 vdd.n614 vdd.n612 39.2114
R3453 vdd.n2822 vdd.n2821 39.2114
R3454 vdd.n2826 vdd.n2825 39.2114
R3455 vdd.n611 vdd.n609 39.2114
R3456 vdd.n2833 vdd.n2832 39.2114
R3457 vdd.n608 vdd.n606 39.2114
R3458 vdd.n2840 vdd.n2839 39.2114
R3459 vdd.n605 vdd.n603 39.2114
R3460 vdd.n2847 vdd.n2846 39.2114
R3461 vdd.n2850 vdd.n2849 39.2114
R3462 vdd.n785 vdd.n740 39.2114
R3463 vdd.n2262 vdd.n741 39.2114
R3464 vdd.n2258 vdd.n742 39.2114
R3465 vdd.n2254 vdd.n743 39.2114
R3466 vdd.n2250 vdd.n744 39.2114
R3467 vdd.n2246 vdd.n745 39.2114
R3468 vdd.n2242 vdd.n746 39.2114
R3469 vdd.n2238 vdd.n747 39.2114
R3470 vdd.n2234 vdd.n748 39.2114
R3471 vdd.n2230 vdd.n749 39.2114
R3472 vdd.n2226 vdd.n750 39.2114
R3473 vdd.n2222 vdd.n751 39.2114
R3474 vdd.n2218 vdd.n752 39.2114
R3475 vdd.n2214 vdd.n753 39.2114
R3476 vdd.n2210 vdd.n754 39.2114
R3477 vdd.n2206 vdd.n755 39.2114
R3478 vdd.n2202 vdd.n756 39.2114
R3479 vdd.n1829 vdd.n899 39.2114
R3480 vdd.n1832 vdd.n1831 39.2114
R3481 vdd.n1837 vdd.n1836 39.2114
R3482 vdd.n1840 vdd.n1839 39.2114
R3483 vdd.n1845 vdd.n1844 39.2114
R3484 vdd.n1848 vdd.n1847 39.2114
R3485 vdd.n1853 vdd.n1852 39.2114
R3486 vdd.n1856 vdd.n1855 39.2114
R3487 vdd.n1861 vdd.n1860 39.2114
R3488 vdd.n1864 vdd.n1863 39.2114
R3489 vdd.n1869 vdd.n1868 39.2114
R3490 vdd.n1872 vdd.n1871 39.2114
R3491 vdd.n1877 vdd.n1876 39.2114
R3492 vdd.n1880 vdd.n1879 39.2114
R3493 vdd.n1885 vdd.n1884 39.2114
R3494 vdd.n1888 vdd.n1887 39.2114
R3495 vdd.n1894 vdd.n1893 39.2114
R3496 vdd.n2199 vdd.n756 39.2114
R3497 vdd.n2203 vdd.n755 39.2114
R3498 vdd.n2207 vdd.n754 39.2114
R3499 vdd.n2211 vdd.n753 39.2114
R3500 vdd.n2215 vdd.n752 39.2114
R3501 vdd.n2219 vdd.n751 39.2114
R3502 vdd.n2223 vdd.n750 39.2114
R3503 vdd.n2227 vdd.n749 39.2114
R3504 vdd.n2231 vdd.n748 39.2114
R3505 vdd.n2235 vdd.n747 39.2114
R3506 vdd.n2239 vdd.n746 39.2114
R3507 vdd.n2243 vdd.n745 39.2114
R3508 vdd.n2247 vdd.n744 39.2114
R3509 vdd.n2251 vdd.n743 39.2114
R3510 vdd.n2255 vdd.n742 39.2114
R3511 vdd.n2259 vdd.n741 39.2114
R3512 vdd.n2263 vdd.n740 39.2114
R3513 vdd.n1830 vdd.n1829 39.2114
R3514 vdd.n1831 vdd.n1827 39.2114
R3515 vdd.n1838 vdd.n1837 39.2114
R3516 vdd.n1839 vdd.n1825 39.2114
R3517 vdd.n1846 vdd.n1845 39.2114
R3518 vdd.n1847 vdd.n1823 39.2114
R3519 vdd.n1854 vdd.n1853 39.2114
R3520 vdd.n1855 vdd.n1821 39.2114
R3521 vdd.n1862 vdd.n1861 39.2114
R3522 vdd.n1863 vdd.n933 39.2114
R3523 vdd.n1870 vdd.n1869 39.2114
R3524 vdd.n1871 vdd.n931 39.2114
R3525 vdd.n1878 vdd.n1877 39.2114
R3526 vdd.n1879 vdd.n929 39.2114
R3527 vdd.n1886 vdd.n1885 39.2114
R3528 vdd.n1887 vdd.n925 39.2114
R3529 vdd.n1895 vdd.n1894 39.2114
R3530 vdd.n1816 vdd.n1815 37.2369
R3531 vdd.n1732 vdd.n1665 37.2369
R3532 vdd.n1771 vdd.n1625 37.2369
R3533 vdd.n2940 vdd.n558 37.2369
R3534 vdd.n2988 vdd.n2987 37.2369
R3535 vdd.n2895 vdd.n2894 37.2369
R3536 vdd.n1891 vdd.n927 30.449
R3537 vdd.n789 vdd.n788 30.449
R3538 vdd.n2016 vdd.n921 30.449
R3539 vdd.n2276 vdd.n779 30.449
R3540 vdd.n2377 vdd.n2376 30.449
R3541 vdd.n2796 vdd.n623 30.449
R3542 vdd.n2504 vdd.n2445 30.449
R3543 vdd.n591 vdd.n590 30.449
R3544 vdd.n2079 vdd.n2078 30.4395
R3545 vdd.n2338 vdd.n777 30.4395
R3546 vdd.n2271 vdd.n780 30.4395
R3547 vdd.n2009 vdd.n2008 30.4395
R3548 vdd.n2511 vdd.n2510 30.4395
R3549 vdd.n2790 vdd.n2789 30.4395
R3550 vdd.n2629 vdd.n2628 30.4395
R3551 vdd.n2853 vdd.n2852 30.4395
R3552 vdd.n2772 vdd.n2771 30.4395
R3553 vdd.n2858 vdd.n592 30.4395
R3554 vdd.n2622 vdd.n2621 30.4395
R3555 vdd.n2633 vdd.n732 30.4395
R3556 vdd.n2083 vdd.n898 30.4395
R3557 vdd.n2266 vdd.n2265 30.4395
R3558 vdd.n2198 vdd.n2197 30.4395
R3559 vdd.n1898 vdd.n1897 30.4395
R3560 vdd.n1501 vdd.n1308 22.6735
R3561 vdd.n1810 vdd.n943 22.6735
R3562 vdd.n3022 vdd.n516 22.6735
R3563 vdd.n3207 vdd.n329 22.6735
R3564 vdd.n1512 vdd.n1270 19.3944
R3565 vdd.n1512 vdd.n1268 19.3944
R3566 vdd.n1516 vdd.n1268 19.3944
R3567 vdd.n1516 vdd.n1258 19.3944
R3568 vdd.n1529 vdd.n1258 19.3944
R3569 vdd.n1529 vdd.n1256 19.3944
R3570 vdd.n1533 vdd.n1256 19.3944
R3571 vdd.n1533 vdd.n1248 19.3944
R3572 vdd.n1547 vdd.n1248 19.3944
R3573 vdd.n1547 vdd.n1246 19.3944
R3574 vdd.n1551 vdd.n1246 19.3944
R3575 vdd.n1551 vdd.n965 19.3944
R3576 vdd.n1563 vdd.n965 19.3944
R3577 vdd.n1563 vdd.n963 19.3944
R3578 vdd.n1567 vdd.n963 19.3944
R3579 vdd.n1567 vdd.n955 19.3944
R3580 vdd.n1580 vdd.n955 19.3944
R3581 vdd.n1580 vdd.n952 19.3944
R3582 vdd.n1586 vdd.n952 19.3944
R3583 vdd.n1586 vdd.n953 19.3944
R3584 vdd.n953 vdd.n942 19.3944
R3585 vdd.n1436 vdd.n1371 19.3944
R3586 vdd.n1432 vdd.n1371 19.3944
R3587 vdd.n1432 vdd.n1431 19.3944
R3588 vdd.n1431 vdd.n1430 19.3944
R3589 vdd.n1430 vdd.n1377 19.3944
R3590 vdd.n1426 vdd.n1377 19.3944
R3591 vdd.n1426 vdd.n1425 19.3944
R3592 vdd.n1425 vdd.n1424 19.3944
R3593 vdd.n1424 vdd.n1383 19.3944
R3594 vdd.n1420 vdd.n1383 19.3944
R3595 vdd.n1420 vdd.n1419 19.3944
R3596 vdd.n1419 vdd.n1418 19.3944
R3597 vdd.n1418 vdd.n1389 19.3944
R3598 vdd.n1414 vdd.n1389 19.3944
R3599 vdd.n1414 vdd.n1413 19.3944
R3600 vdd.n1413 vdd.n1412 19.3944
R3601 vdd.n1412 vdd.n1395 19.3944
R3602 vdd.n1408 vdd.n1395 19.3944
R3603 vdd.n1408 vdd.n1407 19.3944
R3604 vdd.n1407 vdd.n1406 19.3944
R3605 vdd.n1471 vdd.n1470 19.3944
R3606 vdd.n1470 vdd.n1469 19.3944
R3607 vdd.n1469 vdd.n1342 19.3944
R3608 vdd.n1465 vdd.n1342 19.3944
R3609 vdd.n1465 vdd.n1464 19.3944
R3610 vdd.n1464 vdd.n1463 19.3944
R3611 vdd.n1463 vdd.n1348 19.3944
R3612 vdd.n1459 vdd.n1348 19.3944
R3613 vdd.n1459 vdd.n1458 19.3944
R3614 vdd.n1458 vdd.n1457 19.3944
R3615 vdd.n1457 vdd.n1354 19.3944
R3616 vdd.n1453 vdd.n1354 19.3944
R3617 vdd.n1453 vdd.n1452 19.3944
R3618 vdd.n1452 vdd.n1451 19.3944
R3619 vdd.n1451 vdd.n1360 19.3944
R3620 vdd.n1447 vdd.n1360 19.3944
R3621 vdd.n1447 vdd.n1446 19.3944
R3622 vdd.n1446 vdd.n1445 19.3944
R3623 vdd.n1445 vdd.n1366 19.3944
R3624 vdd.n1441 vdd.n1366 19.3944
R3625 vdd.n1504 vdd.n1275 19.3944
R3626 vdd.n1499 vdd.n1275 19.3944
R3627 vdd.n1499 vdd.n1310 19.3944
R3628 vdd.n1495 vdd.n1310 19.3944
R3629 vdd.n1495 vdd.n1494 19.3944
R3630 vdd.n1494 vdd.n1493 19.3944
R3631 vdd.n1493 vdd.n1316 19.3944
R3632 vdd.n1489 vdd.n1316 19.3944
R3633 vdd.n1489 vdd.n1488 19.3944
R3634 vdd.n1488 vdd.n1487 19.3944
R3635 vdd.n1487 vdd.n1322 19.3944
R3636 vdd.n1483 vdd.n1322 19.3944
R3637 vdd.n1483 vdd.n1482 19.3944
R3638 vdd.n1482 vdd.n1481 19.3944
R3639 vdd.n1481 vdd.n1328 19.3944
R3640 vdd.n1477 vdd.n1328 19.3944
R3641 vdd.n1477 vdd.n1476 19.3944
R3642 vdd.n1476 vdd.n1475 19.3944
R3643 vdd.n1728 vdd.n1663 19.3944
R3644 vdd.n1728 vdd.n1669 19.3944
R3645 vdd.n1723 vdd.n1669 19.3944
R3646 vdd.n1723 vdd.n1722 19.3944
R3647 vdd.n1722 vdd.n1721 19.3944
R3648 vdd.n1721 vdd.n1676 19.3944
R3649 vdd.n1716 vdd.n1676 19.3944
R3650 vdd.n1716 vdd.n1715 19.3944
R3651 vdd.n1715 vdd.n1714 19.3944
R3652 vdd.n1714 vdd.n1683 19.3944
R3653 vdd.n1709 vdd.n1683 19.3944
R3654 vdd.n1709 vdd.n1708 19.3944
R3655 vdd.n1708 vdd.n1707 19.3944
R3656 vdd.n1707 vdd.n1691 19.3944
R3657 vdd.n1702 vdd.n1691 19.3944
R3658 vdd.n1702 vdd.n1701 19.3944
R3659 vdd.n1697 vdd.n1696 19.3944
R3660 vdd.n1817 vdd.n938 19.3944
R3661 vdd.n1767 vdd.n1623 19.3944
R3662 vdd.n1767 vdd.n1629 19.3944
R3663 vdd.n1762 vdd.n1629 19.3944
R3664 vdd.n1762 vdd.n1761 19.3944
R3665 vdd.n1761 vdd.n1760 19.3944
R3666 vdd.n1760 vdd.n1636 19.3944
R3667 vdd.n1755 vdd.n1636 19.3944
R3668 vdd.n1755 vdd.n1754 19.3944
R3669 vdd.n1754 vdd.n1753 19.3944
R3670 vdd.n1753 vdd.n1643 19.3944
R3671 vdd.n1748 vdd.n1643 19.3944
R3672 vdd.n1748 vdd.n1747 19.3944
R3673 vdd.n1747 vdd.n1746 19.3944
R3674 vdd.n1746 vdd.n1650 19.3944
R3675 vdd.n1741 vdd.n1650 19.3944
R3676 vdd.n1741 vdd.n1740 19.3944
R3677 vdd.n1740 vdd.n1739 19.3944
R3678 vdd.n1739 vdd.n1657 19.3944
R3679 vdd.n1734 vdd.n1657 19.3944
R3680 vdd.n1734 vdd.n1733 19.3944
R3681 vdd.n1805 vdd.n1804 19.3944
R3682 vdd.n1804 vdd.n1595 19.3944
R3683 vdd.n1799 vdd.n1798 19.3944
R3684 vdd.n1794 vdd.n1599 19.3944
R3685 vdd.n1794 vdd.n1601 19.3944
R3686 vdd.n1604 vdd.n1601 19.3944
R3687 vdd.n1787 vdd.n1604 19.3944
R3688 vdd.n1787 vdd.n1786 19.3944
R3689 vdd.n1786 vdd.n1785 19.3944
R3690 vdd.n1785 vdd.n1610 19.3944
R3691 vdd.n1780 vdd.n1610 19.3944
R3692 vdd.n1780 vdd.n1779 19.3944
R3693 vdd.n1779 vdd.n1778 19.3944
R3694 vdd.n1778 vdd.n1617 19.3944
R3695 vdd.n1773 vdd.n1617 19.3944
R3696 vdd.n1773 vdd.n1772 19.3944
R3697 vdd.n1508 vdd.n1273 19.3944
R3698 vdd.n1508 vdd.n1264 19.3944
R3699 vdd.n1521 vdd.n1264 19.3944
R3700 vdd.n1521 vdd.n1262 19.3944
R3701 vdd.n1525 vdd.n1262 19.3944
R3702 vdd.n1525 vdd.n1253 19.3944
R3703 vdd.n1538 vdd.n1253 19.3944
R3704 vdd.n1538 vdd.n1251 19.3944
R3705 vdd.n1543 vdd.n1251 19.3944
R3706 vdd.n1543 vdd.n1242 19.3944
R3707 vdd.n1555 vdd.n1242 19.3944
R3708 vdd.n1555 vdd.n970 19.3944
R3709 vdd.n1559 vdd.n970 19.3944
R3710 vdd.n1559 vdd.n960 19.3944
R3711 vdd.n1572 vdd.n960 19.3944
R3712 vdd.n1572 vdd.n958 19.3944
R3713 vdd.n1576 vdd.n958 19.3944
R3714 vdd.n1576 vdd.n948 19.3944
R3715 vdd.n1591 vdd.n948 19.3944
R3716 vdd.n1591 vdd.n946 19.3944
R3717 vdd.n1808 vdd.n946 19.3944
R3718 vdd.n3033 vdd.n477 19.3944
R3719 vdd.n3033 vdd.n475 19.3944
R3720 vdd.n3037 vdd.n475 19.3944
R3721 vdd.n3037 vdd.n465 19.3944
R3722 vdd.n3050 vdd.n465 19.3944
R3723 vdd.n3050 vdd.n463 19.3944
R3724 vdd.n3054 vdd.n463 19.3944
R3725 vdd.n3054 vdd.n453 19.3944
R3726 vdd.n3066 vdd.n453 19.3944
R3727 vdd.n3066 vdd.n451 19.3944
R3728 vdd.n3070 vdd.n451 19.3944
R3729 vdd.n3071 vdd.n3070 19.3944
R3730 vdd.n3072 vdd.n3071 19.3944
R3731 vdd.n3072 vdd.n449 19.3944
R3732 vdd.n3076 vdd.n449 19.3944
R3733 vdd.n3077 vdd.n3076 19.3944
R3734 vdd.n3078 vdd.n3077 19.3944
R3735 vdd.n3078 vdd.n446 19.3944
R3736 vdd.n3082 vdd.n446 19.3944
R3737 vdd.n3083 vdd.n3082 19.3944
R3738 vdd.n3084 vdd.n3083 19.3944
R3739 vdd.n3127 vdd.n404 19.3944
R3740 vdd.n3127 vdd.n410 19.3944
R3741 vdd.n3122 vdd.n410 19.3944
R3742 vdd.n3122 vdd.n3121 19.3944
R3743 vdd.n3121 vdd.n3120 19.3944
R3744 vdd.n3120 vdd.n417 19.3944
R3745 vdd.n3115 vdd.n417 19.3944
R3746 vdd.n3115 vdd.n3114 19.3944
R3747 vdd.n3114 vdd.n3113 19.3944
R3748 vdd.n3113 vdd.n424 19.3944
R3749 vdd.n3108 vdd.n424 19.3944
R3750 vdd.n3108 vdd.n3107 19.3944
R3751 vdd.n3107 vdd.n3106 19.3944
R3752 vdd.n3106 vdd.n431 19.3944
R3753 vdd.n3101 vdd.n431 19.3944
R3754 vdd.n3101 vdd.n3100 19.3944
R3755 vdd.n3100 vdd.n3099 19.3944
R3756 vdd.n3099 vdd.n438 19.3944
R3757 vdd.n3094 vdd.n438 19.3944
R3758 vdd.n3094 vdd.n3093 19.3944
R3759 vdd.n3166 vdd.n364 19.3944
R3760 vdd.n3166 vdd.n370 19.3944
R3761 vdd.n3161 vdd.n370 19.3944
R3762 vdd.n3161 vdd.n3160 19.3944
R3763 vdd.n3160 vdd.n3159 19.3944
R3764 vdd.n3159 vdd.n377 19.3944
R3765 vdd.n3154 vdd.n377 19.3944
R3766 vdd.n3154 vdd.n3153 19.3944
R3767 vdd.n3153 vdd.n3152 19.3944
R3768 vdd.n3152 vdd.n384 19.3944
R3769 vdd.n3147 vdd.n384 19.3944
R3770 vdd.n3147 vdd.n3146 19.3944
R3771 vdd.n3146 vdd.n3145 19.3944
R3772 vdd.n3145 vdd.n391 19.3944
R3773 vdd.n3140 vdd.n391 19.3944
R3774 vdd.n3140 vdd.n3139 19.3944
R3775 vdd.n3139 vdd.n3138 19.3944
R3776 vdd.n3138 vdd.n398 19.3944
R3777 vdd.n3133 vdd.n398 19.3944
R3778 vdd.n3133 vdd.n3132 19.3944
R3779 vdd.n3202 vdd.n3201 19.3944
R3780 vdd.n3201 vdd.n3200 19.3944
R3781 vdd.n3200 vdd.n336 19.3944
R3782 vdd.n337 vdd.n336 19.3944
R3783 vdd.n3193 vdd.n337 19.3944
R3784 vdd.n3193 vdd.n3192 19.3944
R3785 vdd.n3192 vdd.n3191 19.3944
R3786 vdd.n3191 vdd.n344 19.3944
R3787 vdd.n3186 vdd.n344 19.3944
R3788 vdd.n3186 vdd.n3185 19.3944
R3789 vdd.n3185 vdd.n3184 19.3944
R3790 vdd.n3184 vdd.n351 19.3944
R3791 vdd.n3179 vdd.n351 19.3944
R3792 vdd.n3179 vdd.n3178 19.3944
R3793 vdd.n3178 vdd.n3177 19.3944
R3794 vdd.n3177 vdd.n358 19.3944
R3795 vdd.n3172 vdd.n358 19.3944
R3796 vdd.n3172 vdd.n3171 19.3944
R3797 vdd.n3029 vdd.n480 19.3944
R3798 vdd.n3029 vdd.n471 19.3944
R3799 vdd.n3042 vdd.n471 19.3944
R3800 vdd.n3042 vdd.n469 19.3944
R3801 vdd.n3046 vdd.n469 19.3944
R3802 vdd.n3046 vdd.n460 19.3944
R3803 vdd.n3058 vdd.n460 19.3944
R3804 vdd.n3058 vdd.n458 19.3944
R3805 vdd.n3062 vdd.n458 19.3944
R3806 vdd.n3062 vdd.n300 19.3944
R3807 vdd.n3227 vdd.n300 19.3944
R3808 vdd.n3227 vdd.n301 19.3944
R3809 vdd.n3221 vdd.n301 19.3944
R3810 vdd.n3221 vdd.n3220 19.3944
R3811 vdd.n3220 vdd.n3219 19.3944
R3812 vdd.n3219 vdd.n313 19.3944
R3813 vdd.n3213 vdd.n313 19.3944
R3814 vdd.n3213 vdd.n3212 19.3944
R3815 vdd.n3212 vdd.n3211 19.3944
R3816 vdd.n3211 vdd.n324 19.3944
R3817 vdd.n3205 vdd.n324 19.3944
R3818 vdd.n2982 vdd.n536 19.3944
R3819 vdd.n2982 vdd.n2979 19.3944
R3820 vdd.n2979 vdd.n2976 19.3944
R3821 vdd.n2976 vdd.n2975 19.3944
R3822 vdd.n2975 vdd.n2972 19.3944
R3823 vdd.n2972 vdd.n2971 19.3944
R3824 vdd.n2971 vdd.n2968 19.3944
R3825 vdd.n2968 vdd.n2967 19.3944
R3826 vdd.n2967 vdd.n2964 19.3944
R3827 vdd.n2964 vdd.n2963 19.3944
R3828 vdd.n2963 vdd.n2960 19.3944
R3829 vdd.n2960 vdd.n2959 19.3944
R3830 vdd.n2959 vdd.n2956 19.3944
R3831 vdd.n2956 vdd.n2955 19.3944
R3832 vdd.n2955 vdd.n2952 19.3944
R3833 vdd.n2952 vdd.n2951 19.3944
R3834 vdd.n2951 vdd.n2948 19.3944
R3835 vdd.n2948 vdd.n2947 19.3944
R3836 vdd.n2947 vdd.n2944 19.3944
R3837 vdd.n2944 vdd.n2943 19.3944
R3838 vdd.n3025 vdd.n482 19.3944
R3839 vdd.n3020 vdd.n482 19.3944
R3840 vdd.n521 vdd.n518 19.3944
R3841 vdd.n3016 vdd.n3015 19.3944
R3842 vdd.n3015 vdd.n3012 19.3944
R3843 vdd.n3012 vdd.n3011 19.3944
R3844 vdd.n3011 vdd.n3008 19.3944
R3845 vdd.n3008 vdd.n3007 19.3944
R3846 vdd.n3007 vdd.n3004 19.3944
R3847 vdd.n3004 vdd.n3003 19.3944
R3848 vdd.n3003 vdd.n3000 19.3944
R3849 vdd.n3000 vdd.n2999 19.3944
R3850 vdd.n2999 vdd.n2996 19.3944
R3851 vdd.n2996 vdd.n2995 19.3944
R3852 vdd.n2995 vdd.n2992 19.3944
R3853 vdd.n2992 vdd.n2991 19.3944
R3854 vdd.n2936 vdd.n556 19.3944
R3855 vdd.n2936 vdd.n2933 19.3944
R3856 vdd.n2933 vdd.n2930 19.3944
R3857 vdd.n2930 vdd.n2929 19.3944
R3858 vdd.n2929 vdd.n2926 19.3944
R3859 vdd.n2926 vdd.n2925 19.3944
R3860 vdd.n2925 vdd.n2922 19.3944
R3861 vdd.n2922 vdd.n2921 19.3944
R3862 vdd.n2921 vdd.n2918 19.3944
R3863 vdd.n2918 vdd.n2917 19.3944
R3864 vdd.n2917 vdd.n2914 19.3944
R3865 vdd.n2914 vdd.n2913 19.3944
R3866 vdd.n2913 vdd.n2910 19.3944
R3867 vdd.n2910 vdd.n2909 19.3944
R3868 vdd.n2909 vdd.n2906 19.3944
R3869 vdd.n2906 vdd.n2905 19.3944
R3870 vdd.n2902 vdd.n2901 19.3944
R3871 vdd.n2898 vdd.n2897 19.3944
R3872 vdd.n1440 vdd.n1436 19.0066
R3873 vdd.n1732 vdd.n1663 19.0066
R3874 vdd.n3131 vdd.n404 19.0066
R3875 vdd.n2940 vdd.n556 19.0066
R3876 vdd.n927 vdd.n926 16.0975
R3877 vdd.n788 vdd.n787 16.0975
R3878 vdd.n1401 vdd.n1400 16.0975
R3879 vdd.n1439 vdd.n1438 16.0975
R3880 vdd.n1335 vdd.n1334 16.0975
R3881 vdd.n1815 vdd.n1814 16.0975
R3882 vdd.n1665 vdd.n1664 16.0975
R3883 vdd.n1625 vdd.n1624 16.0975
R3884 vdd.n921 vdd.n920 16.0975
R3885 vdd.n779 vdd.n778 16.0975
R3886 vdd.n2376 vdd.n2375 16.0975
R3887 vdd.n3091 vdd.n3090 16.0975
R3888 vdd.n406 vdd.n405 16.0975
R3889 vdd.n366 vdd.n365 16.0975
R3890 vdd.n558 vdd.n557 16.0975
R3891 vdd.n2987 vdd.n2986 16.0975
R3892 vdd.n623 vdd.n622 16.0975
R3893 vdd.n2445 vdd.n2444 16.0975
R3894 vdd.n2894 vdd.n2893 16.0975
R3895 vdd.n590 vdd.n589 16.0975
R3896 vdd.t172 vdd.n2340 15.4182
R3897 vdd.n2624 vdd.t162 15.4182
R3898 vdd.n28 vdd.n27 14.8572
R3899 vdd.n2081 vdd.n900 13.6043
R3900 vdd.n2855 vdd.n484 13.6043
R3901 vdd.n292 vdd.n257 13.1884
R3902 vdd.n245 vdd.n210 13.1884
R3903 vdd.n202 vdd.n167 13.1884
R3904 vdd.n155 vdd.n120 13.1884
R3905 vdd.n113 vdd.n78 13.1884
R3906 vdd.n66 vdd.n31 13.1884
R3907 vdd.n1187 vdd.n1152 13.1884
R3908 vdd.n1234 vdd.n1199 13.1884
R3909 vdd.n1097 vdd.n1062 13.1884
R3910 vdd.n1144 vdd.n1109 13.1884
R3911 vdd.n1008 vdd.n973 13.1884
R3912 vdd.n1055 vdd.n1020 13.1884
R3913 vdd.n1471 vdd.n1336 12.9944
R3914 vdd.n1475 vdd.n1336 12.9944
R3915 vdd.n1771 vdd.n1623 12.9944
R3916 vdd.n1772 vdd.n1771 12.9944
R3917 vdd.n3170 vdd.n364 12.9944
R3918 vdd.n3171 vdd.n3170 12.9944
R3919 vdd.n2988 vdd.n536 12.9944
R3920 vdd.n2991 vdd.n2988 12.9944
R3921 vdd.n293 vdd.n255 12.8005
R3922 vdd.n288 vdd.n259 12.8005
R3923 vdd.n246 vdd.n208 12.8005
R3924 vdd.n241 vdd.n212 12.8005
R3925 vdd.n203 vdd.n165 12.8005
R3926 vdd.n198 vdd.n169 12.8005
R3927 vdd.n156 vdd.n118 12.8005
R3928 vdd.n151 vdd.n122 12.8005
R3929 vdd.n114 vdd.n76 12.8005
R3930 vdd.n109 vdd.n80 12.8005
R3931 vdd.n67 vdd.n29 12.8005
R3932 vdd.n62 vdd.n33 12.8005
R3933 vdd.n1188 vdd.n1150 12.8005
R3934 vdd.n1183 vdd.n1154 12.8005
R3935 vdd.n1235 vdd.n1197 12.8005
R3936 vdd.n1230 vdd.n1201 12.8005
R3937 vdd.n1098 vdd.n1060 12.8005
R3938 vdd.n1093 vdd.n1064 12.8005
R3939 vdd.n1145 vdd.n1107 12.8005
R3940 vdd.n1140 vdd.n1111 12.8005
R3941 vdd.n1009 vdd.n971 12.8005
R3942 vdd.n1004 vdd.n975 12.8005
R3943 vdd.n1056 vdd.n1018 12.8005
R3944 vdd.n1051 vdd.n1022 12.8005
R3945 vdd.n287 vdd.n260 12.0247
R3946 vdd.n240 vdd.n213 12.0247
R3947 vdd.n197 vdd.n170 12.0247
R3948 vdd.n150 vdd.n123 12.0247
R3949 vdd.n108 vdd.n81 12.0247
R3950 vdd.n61 vdd.n34 12.0247
R3951 vdd.n1182 vdd.n1155 12.0247
R3952 vdd.n1229 vdd.n1202 12.0247
R3953 vdd.n1092 vdd.n1065 12.0247
R3954 vdd.n1139 vdd.n1112 12.0247
R3955 vdd.n1003 vdd.n976 12.0247
R3956 vdd.n1050 vdd.n1023 12.0247
R3957 vdd.n1510 vdd.n1266 11.337
R3958 vdd.n1519 vdd.n1266 11.337
R3959 vdd.n1519 vdd.n1518 11.337
R3960 vdd.n1527 vdd.n1260 11.337
R3961 vdd.n1536 vdd.n1535 11.337
R3962 vdd.n1553 vdd.n1244 11.337
R3963 vdd.n1561 vdd.n967 11.337
R3964 vdd.n1570 vdd.n1569 11.337
R3965 vdd.n1578 vdd.n950 11.337
R3966 vdd.n1589 vdd.n950 11.337
R3967 vdd.n1589 vdd.n1588 11.337
R3968 vdd.n3031 vdd.n473 11.337
R3969 vdd.n3040 vdd.n473 11.337
R3970 vdd.n3040 vdd.n3039 11.337
R3971 vdd.n3048 vdd.n467 11.337
R3972 vdd.n3064 vdd.n456 11.337
R3973 vdd.n3225 vdd.n304 11.337
R3974 vdd.n3223 vdd.n308 11.337
R3975 vdd.n3217 vdd.n3216 11.337
R3976 vdd.n3215 vdd.n318 11.337
R3977 vdd.n3209 vdd.n318 11.337
R3978 vdd.n3209 vdd.n3208 11.337
R3979 vdd.n284 vdd.n283 11.249
R3980 vdd.n237 vdd.n236 11.249
R3981 vdd.n194 vdd.n193 11.249
R3982 vdd.n147 vdd.n146 11.249
R3983 vdd.n105 vdd.n104 11.249
R3984 vdd.n58 vdd.n57 11.249
R3985 vdd.n1179 vdd.n1178 11.249
R3986 vdd.n1226 vdd.n1225 11.249
R3987 vdd.n1089 vdd.n1088 11.249
R3988 vdd.n1136 vdd.n1135 11.249
R3989 vdd.n1000 vdd.n999 11.249
R3990 vdd.n1047 vdd.n1046 11.249
R3991 vdd.n1308 vdd.t33 10.7702
R3992 vdd.t29 vdd.n3207 10.7702
R3993 vdd.n269 vdd.n268 10.7238
R3994 vdd.n222 vdd.n221 10.7238
R3995 vdd.n179 vdd.n178 10.7238
R3996 vdd.n132 vdd.n131 10.7238
R3997 vdd.n90 vdd.n89 10.7238
R3998 vdd.n43 vdd.n42 10.7238
R3999 vdd.n1164 vdd.n1163 10.7238
R4000 vdd.n1211 vdd.n1210 10.7238
R4001 vdd.n1074 vdd.n1073 10.7238
R4002 vdd.n1121 vdd.n1120 10.7238
R4003 vdd.n985 vdd.n984 10.7238
R4004 vdd.n1032 vdd.n1031 10.7238
R4005 vdd.n2079 vdd.n892 10.6151
R4006 vdd.n2089 vdd.n892 10.6151
R4007 vdd.n2090 vdd.n2089 10.6151
R4008 vdd.n2091 vdd.n2090 10.6151
R4009 vdd.n2091 vdd.n880 10.6151
R4010 vdd.n2101 vdd.n880 10.6151
R4011 vdd.n2102 vdd.n2101 10.6151
R4012 vdd.n2103 vdd.n2102 10.6151
R4013 vdd.n2103 vdd.n868 10.6151
R4014 vdd.n2113 vdd.n868 10.6151
R4015 vdd.n2114 vdd.n2113 10.6151
R4016 vdd.n2115 vdd.n2114 10.6151
R4017 vdd.n2115 vdd.n855 10.6151
R4018 vdd.n2125 vdd.n855 10.6151
R4019 vdd.n2126 vdd.n2125 10.6151
R4020 vdd.n2127 vdd.n2126 10.6151
R4021 vdd.n2127 vdd.n843 10.6151
R4022 vdd.n2138 vdd.n843 10.6151
R4023 vdd.n2139 vdd.n2138 10.6151
R4024 vdd.n2140 vdd.n2139 10.6151
R4025 vdd.n2140 vdd.n831 10.6151
R4026 vdd.n2150 vdd.n831 10.6151
R4027 vdd.n2151 vdd.n2150 10.6151
R4028 vdd.n2152 vdd.n2151 10.6151
R4029 vdd.n2152 vdd.n819 10.6151
R4030 vdd.n2162 vdd.n819 10.6151
R4031 vdd.n2163 vdd.n2162 10.6151
R4032 vdd.n2164 vdd.n2163 10.6151
R4033 vdd.n2164 vdd.n809 10.6151
R4034 vdd.n2174 vdd.n809 10.6151
R4035 vdd.n2175 vdd.n2174 10.6151
R4036 vdd.n2176 vdd.n2175 10.6151
R4037 vdd.n2176 vdd.n796 10.6151
R4038 vdd.n2188 vdd.n796 10.6151
R4039 vdd.n2189 vdd.n2188 10.6151
R4040 vdd.n2191 vdd.n2189 10.6151
R4041 vdd.n2191 vdd.n2190 10.6151
R4042 vdd.n2190 vdd.n777 10.6151
R4043 vdd.n2338 vdd.n2337 10.6151
R4044 vdd.n2337 vdd.n2336 10.6151
R4045 vdd.n2336 vdd.n2333 10.6151
R4046 vdd.n2333 vdd.n2332 10.6151
R4047 vdd.n2332 vdd.n2329 10.6151
R4048 vdd.n2329 vdd.n2328 10.6151
R4049 vdd.n2328 vdd.n2325 10.6151
R4050 vdd.n2325 vdd.n2324 10.6151
R4051 vdd.n2324 vdd.n2321 10.6151
R4052 vdd.n2321 vdd.n2320 10.6151
R4053 vdd.n2320 vdd.n2317 10.6151
R4054 vdd.n2317 vdd.n2316 10.6151
R4055 vdd.n2316 vdd.n2313 10.6151
R4056 vdd.n2313 vdd.n2312 10.6151
R4057 vdd.n2312 vdd.n2309 10.6151
R4058 vdd.n2309 vdd.n2308 10.6151
R4059 vdd.n2308 vdd.n2305 10.6151
R4060 vdd.n2305 vdd.n2304 10.6151
R4061 vdd.n2304 vdd.n2301 10.6151
R4062 vdd.n2301 vdd.n2300 10.6151
R4063 vdd.n2300 vdd.n2297 10.6151
R4064 vdd.n2297 vdd.n2296 10.6151
R4065 vdd.n2296 vdd.n2293 10.6151
R4066 vdd.n2293 vdd.n2292 10.6151
R4067 vdd.n2292 vdd.n2289 10.6151
R4068 vdd.n2289 vdd.n2288 10.6151
R4069 vdd.n2288 vdd.n2285 10.6151
R4070 vdd.n2285 vdd.n2284 10.6151
R4071 vdd.n2284 vdd.n2281 10.6151
R4072 vdd.n2281 vdd.n2280 10.6151
R4073 vdd.n2280 vdd.n2277 10.6151
R4074 vdd.n2275 vdd.n2272 10.6151
R4075 vdd.n2272 vdd.n2271 10.6151
R4076 vdd.n2008 vdd.n2007 10.6151
R4077 vdd.n2007 vdd.n2005 10.6151
R4078 vdd.n2005 vdd.n2004 10.6151
R4079 vdd.n2004 vdd.n2002 10.6151
R4080 vdd.n2002 vdd.n2001 10.6151
R4081 vdd.n2001 vdd.n1999 10.6151
R4082 vdd.n1999 vdd.n1998 10.6151
R4083 vdd.n1998 vdd.n1996 10.6151
R4084 vdd.n1996 vdd.n1995 10.6151
R4085 vdd.n1995 vdd.n1993 10.6151
R4086 vdd.n1993 vdd.n1992 10.6151
R4087 vdd.n1992 vdd.n1990 10.6151
R4088 vdd.n1990 vdd.n1989 10.6151
R4089 vdd.n1989 vdd.n1987 10.6151
R4090 vdd.n1987 vdd.n1986 10.6151
R4091 vdd.n1986 vdd.n1984 10.6151
R4092 vdd.n1984 vdd.n1983 10.6151
R4093 vdd.n1983 vdd.n1981 10.6151
R4094 vdd.n1981 vdd.n1980 10.6151
R4095 vdd.n1980 vdd.n1978 10.6151
R4096 vdd.n1978 vdd.n1977 10.6151
R4097 vdd.n1977 vdd.n1975 10.6151
R4098 vdd.n1975 vdd.n1974 10.6151
R4099 vdd.n1974 vdd.n923 10.6151
R4100 vdd.n1941 vdd.n923 10.6151
R4101 vdd.n1942 vdd.n1941 10.6151
R4102 vdd.n1944 vdd.n1942 10.6151
R4103 vdd.n1945 vdd.n1944 10.6151
R4104 vdd.n1958 vdd.n1945 10.6151
R4105 vdd.n1958 vdd.n1957 10.6151
R4106 vdd.n1957 vdd.n1956 10.6151
R4107 vdd.n1956 vdd.n1954 10.6151
R4108 vdd.n1954 vdd.n1953 10.6151
R4109 vdd.n1953 vdd.n1951 10.6151
R4110 vdd.n1951 vdd.n1950 10.6151
R4111 vdd.n1950 vdd.n1947 10.6151
R4112 vdd.n1947 vdd.n1946 10.6151
R4113 vdd.n1946 vdd.n780 10.6151
R4114 vdd.n2078 vdd.n2077 10.6151
R4115 vdd.n2077 vdd.n904 10.6151
R4116 vdd.n2072 vdd.n904 10.6151
R4117 vdd.n2072 vdd.n2071 10.6151
R4118 vdd.n2071 vdd.n906 10.6151
R4119 vdd.n2066 vdd.n906 10.6151
R4120 vdd.n2066 vdd.n2065 10.6151
R4121 vdd.n2065 vdd.n2064 10.6151
R4122 vdd.n2064 vdd.n908 10.6151
R4123 vdd.n2058 vdd.n908 10.6151
R4124 vdd.n2058 vdd.n2057 10.6151
R4125 vdd.n2057 vdd.n2056 10.6151
R4126 vdd.n2056 vdd.n910 10.6151
R4127 vdd.n2050 vdd.n910 10.6151
R4128 vdd.n2050 vdd.n2049 10.6151
R4129 vdd.n2049 vdd.n2048 10.6151
R4130 vdd.n2048 vdd.n912 10.6151
R4131 vdd.n2042 vdd.n912 10.6151
R4132 vdd.n2042 vdd.n2041 10.6151
R4133 vdd.n2041 vdd.n2040 10.6151
R4134 vdd.n2040 vdd.n914 10.6151
R4135 vdd.n2034 vdd.n914 10.6151
R4136 vdd.n2034 vdd.n2033 10.6151
R4137 vdd.n2033 vdd.n2032 10.6151
R4138 vdd.n2032 vdd.n916 10.6151
R4139 vdd.n2026 vdd.n916 10.6151
R4140 vdd.n2026 vdd.n2025 10.6151
R4141 vdd.n2025 vdd.n2024 10.6151
R4142 vdd.n2024 vdd.n918 10.6151
R4143 vdd.n2018 vdd.n918 10.6151
R4144 vdd.n2018 vdd.n2017 10.6151
R4145 vdd.n2015 vdd.n922 10.6151
R4146 vdd.n2009 vdd.n922 10.6151
R4147 vdd.n2513 vdd.n2511 10.6151
R4148 vdd.n2514 vdd.n2513 10.6151
R4149 vdd.n2613 vdd.n2514 10.6151
R4150 vdd.n2613 vdd.n2612 10.6151
R4151 vdd.n2612 vdd.n2611 10.6151
R4152 vdd.n2611 vdd.n2609 10.6151
R4153 vdd.n2609 vdd.n2608 10.6151
R4154 vdd.n2608 vdd.n2606 10.6151
R4155 vdd.n2606 vdd.n2605 10.6151
R4156 vdd.n2605 vdd.n2515 10.6151
R4157 vdd.n2555 vdd.n2515 10.6151
R4158 vdd.n2556 vdd.n2555 10.6151
R4159 vdd.n2558 vdd.n2556 10.6151
R4160 vdd.n2559 vdd.n2558 10.6151
R4161 vdd.n2589 vdd.n2559 10.6151
R4162 vdd.n2589 vdd.n2588 10.6151
R4163 vdd.n2588 vdd.n2587 10.6151
R4164 vdd.n2587 vdd.n2585 10.6151
R4165 vdd.n2585 vdd.n2584 10.6151
R4166 vdd.n2584 vdd.n2582 10.6151
R4167 vdd.n2582 vdd.n2581 10.6151
R4168 vdd.n2581 vdd.n2579 10.6151
R4169 vdd.n2579 vdd.n2578 10.6151
R4170 vdd.n2578 vdd.n2576 10.6151
R4171 vdd.n2576 vdd.n2575 10.6151
R4172 vdd.n2575 vdd.n2573 10.6151
R4173 vdd.n2573 vdd.n2572 10.6151
R4174 vdd.n2572 vdd.n2570 10.6151
R4175 vdd.n2570 vdd.n2569 10.6151
R4176 vdd.n2569 vdd.n2567 10.6151
R4177 vdd.n2567 vdd.n2566 10.6151
R4178 vdd.n2566 vdd.n2564 10.6151
R4179 vdd.n2564 vdd.n2563 10.6151
R4180 vdd.n2563 vdd.n2561 10.6151
R4181 vdd.n2561 vdd.n2560 10.6151
R4182 vdd.n2560 vdd.n626 10.6151
R4183 vdd.n2788 vdd.n626 10.6151
R4184 vdd.n2789 vdd.n2788 10.6151
R4185 vdd.n2628 vdd.n2627 10.6151
R4186 vdd.n2627 vdd.n738 10.6151
R4187 vdd.n2447 vdd.n738 10.6151
R4188 vdd.n2448 vdd.n2447 10.6151
R4189 vdd.n2451 vdd.n2448 10.6151
R4190 vdd.n2452 vdd.n2451 10.6151
R4191 vdd.n2455 vdd.n2452 10.6151
R4192 vdd.n2456 vdd.n2455 10.6151
R4193 vdd.n2459 vdd.n2456 10.6151
R4194 vdd.n2460 vdd.n2459 10.6151
R4195 vdd.n2463 vdd.n2460 10.6151
R4196 vdd.n2464 vdd.n2463 10.6151
R4197 vdd.n2467 vdd.n2464 10.6151
R4198 vdd.n2468 vdd.n2467 10.6151
R4199 vdd.n2471 vdd.n2468 10.6151
R4200 vdd.n2472 vdd.n2471 10.6151
R4201 vdd.n2475 vdd.n2472 10.6151
R4202 vdd.n2476 vdd.n2475 10.6151
R4203 vdd.n2479 vdd.n2476 10.6151
R4204 vdd.n2480 vdd.n2479 10.6151
R4205 vdd.n2483 vdd.n2480 10.6151
R4206 vdd.n2484 vdd.n2483 10.6151
R4207 vdd.n2487 vdd.n2484 10.6151
R4208 vdd.n2488 vdd.n2487 10.6151
R4209 vdd.n2491 vdd.n2488 10.6151
R4210 vdd.n2492 vdd.n2491 10.6151
R4211 vdd.n2495 vdd.n2492 10.6151
R4212 vdd.n2496 vdd.n2495 10.6151
R4213 vdd.n2499 vdd.n2496 10.6151
R4214 vdd.n2500 vdd.n2499 10.6151
R4215 vdd.n2503 vdd.n2500 10.6151
R4216 vdd.n2508 vdd.n2505 10.6151
R4217 vdd.n2510 vdd.n2508 10.6151
R4218 vdd.n2629 vdd.n727 10.6151
R4219 vdd.n2639 vdd.n727 10.6151
R4220 vdd.n2640 vdd.n2639 10.6151
R4221 vdd.n2641 vdd.n2640 10.6151
R4222 vdd.n2641 vdd.n715 10.6151
R4223 vdd.n2651 vdd.n715 10.6151
R4224 vdd.n2652 vdd.n2651 10.6151
R4225 vdd.n2653 vdd.n2652 10.6151
R4226 vdd.n2653 vdd.n705 10.6151
R4227 vdd.n2663 vdd.n705 10.6151
R4228 vdd.n2664 vdd.n2663 10.6151
R4229 vdd.n2665 vdd.n2664 10.6151
R4230 vdd.n2665 vdd.n693 10.6151
R4231 vdd.n2675 vdd.n693 10.6151
R4232 vdd.n2676 vdd.n2675 10.6151
R4233 vdd.n2677 vdd.n2676 10.6151
R4234 vdd.n2677 vdd.n682 10.6151
R4235 vdd.n2687 vdd.n682 10.6151
R4236 vdd.n2688 vdd.n2687 10.6151
R4237 vdd.n2689 vdd.n2688 10.6151
R4238 vdd.n2689 vdd.n669 10.6151
R4239 vdd.n2700 vdd.n669 10.6151
R4240 vdd.n2701 vdd.n2700 10.6151
R4241 vdd.n2702 vdd.n2701 10.6151
R4242 vdd.n2702 vdd.n656 10.6151
R4243 vdd.n2712 vdd.n656 10.6151
R4244 vdd.n2713 vdd.n2712 10.6151
R4245 vdd.n2714 vdd.n2713 10.6151
R4246 vdd.n2714 vdd.n645 10.6151
R4247 vdd.n2724 vdd.n645 10.6151
R4248 vdd.n2725 vdd.n2724 10.6151
R4249 vdd.n2726 vdd.n2725 10.6151
R4250 vdd.n2726 vdd.n631 10.6151
R4251 vdd.n2781 vdd.n631 10.6151
R4252 vdd.n2782 vdd.n2781 10.6151
R4253 vdd.n2783 vdd.n2782 10.6151
R4254 vdd.n2783 vdd.n600 10.6151
R4255 vdd.n2853 vdd.n600 10.6151
R4256 vdd.n2852 vdd.n2851 10.6151
R4257 vdd.n2851 vdd.n601 10.6151
R4258 vdd.n602 vdd.n601 10.6151
R4259 vdd.n2844 vdd.n602 10.6151
R4260 vdd.n2844 vdd.n2843 10.6151
R4261 vdd.n2843 vdd.n2842 10.6151
R4262 vdd.n2842 vdd.n604 10.6151
R4263 vdd.n2837 vdd.n604 10.6151
R4264 vdd.n2837 vdd.n2836 10.6151
R4265 vdd.n2836 vdd.n2835 10.6151
R4266 vdd.n2835 vdd.n607 10.6151
R4267 vdd.n2830 vdd.n607 10.6151
R4268 vdd.n2830 vdd.n2829 10.6151
R4269 vdd.n2829 vdd.n2828 10.6151
R4270 vdd.n2828 vdd.n610 10.6151
R4271 vdd.n2823 vdd.n610 10.6151
R4272 vdd.n2823 vdd.n520 10.6151
R4273 vdd.n2819 vdd.n520 10.6151
R4274 vdd.n2819 vdd.n2818 10.6151
R4275 vdd.n2818 vdd.n2817 10.6151
R4276 vdd.n2817 vdd.n613 10.6151
R4277 vdd.n2812 vdd.n613 10.6151
R4278 vdd.n2812 vdd.n2811 10.6151
R4279 vdd.n2811 vdd.n2810 10.6151
R4280 vdd.n2810 vdd.n616 10.6151
R4281 vdd.n2805 vdd.n616 10.6151
R4282 vdd.n2805 vdd.n2804 10.6151
R4283 vdd.n2804 vdd.n2803 10.6151
R4284 vdd.n2803 vdd.n619 10.6151
R4285 vdd.n2798 vdd.n619 10.6151
R4286 vdd.n2798 vdd.n2797 10.6151
R4287 vdd.n2795 vdd.n624 10.6151
R4288 vdd.n2790 vdd.n624 10.6151
R4289 vdd.n2771 vdd.n2732 10.6151
R4290 vdd.n2766 vdd.n2732 10.6151
R4291 vdd.n2766 vdd.n2765 10.6151
R4292 vdd.n2765 vdd.n2764 10.6151
R4293 vdd.n2764 vdd.n2734 10.6151
R4294 vdd.n2759 vdd.n2734 10.6151
R4295 vdd.n2759 vdd.n2758 10.6151
R4296 vdd.n2758 vdd.n2757 10.6151
R4297 vdd.n2757 vdd.n2737 10.6151
R4298 vdd.n2752 vdd.n2737 10.6151
R4299 vdd.n2752 vdd.n2751 10.6151
R4300 vdd.n2751 vdd.n2750 10.6151
R4301 vdd.n2750 vdd.n2740 10.6151
R4302 vdd.n2745 vdd.n2740 10.6151
R4303 vdd.n2745 vdd.n2744 10.6151
R4304 vdd.n2744 vdd.n575 10.6151
R4305 vdd.n2888 vdd.n575 10.6151
R4306 vdd.n2888 vdd.n576 10.6151
R4307 vdd.n578 vdd.n576 10.6151
R4308 vdd.n2881 vdd.n578 10.6151
R4309 vdd.n2881 vdd.n2880 10.6151
R4310 vdd.n2880 vdd.n2879 10.6151
R4311 vdd.n2879 vdd.n580 10.6151
R4312 vdd.n2874 vdd.n580 10.6151
R4313 vdd.n2874 vdd.n2873 10.6151
R4314 vdd.n2873 vdd.n2872 10.6151
R4315 vdd.n2872 vdd.n583 10.6151
R4316 vdd.n2867 vdd.n583 10.6151
R4317 vdd.n2867 vdd.n2866 10.6151
R4318 vdd.n2866 vdd.n2865 10.6151
R4319 vdd.n2865 vdd.n586 10.6151
R4320 vdd.n2860 vdd.n2859 10.6151
R4321 vdd.n2859 vdd.n2858 10.6151
R4322 vdd.n2621 vdd.n2620 10.6151
R4323 vdd.n2620 vdd.n2618 10.6151
R4324 vdd.n2618 vdd.n2617 10.6151
R4325 vdd.n2617 vdd.n2443 10.6151
R4326 vdd.n2517 vdd.n2443 10.6151
R4327 vdd.n2518 vdd.n2517 10.6151
R4328 vdd.n2520 vdd.n2518 10.6151
R4329 vdd.n2521 vdd.n2520 10.6151
R4330 vdd.n2601 vdd.n2521 10.6151
R4331 vdd.n2601 vdd.n2600 10.6151
R4332 vdd.n2600 vdd.n2599 10.6151
R4333 vdd.n2599 vdd.n2597 10.6151
R4334 vdd.n2597 vdd.n2596 10.6151
R4335 vdd.n2596 vdd.n2594 10.6151
R4336 vdd.n2594 vdd.n2593 10.6151
R4337 vdd.n2593 vdd.n2553 10.6151
R4338 vdd.n2553 vdd.n2552 10.6151
R4339 vdd.n2552 vdd.n2550 10.6151
R4340 vdd.n2550 vdd.n2549 10.6151
R4341 vdd.n2549 vdd.n2547 10.6151
R4342 vdd.n2547 vdd.n2546 10.6151
R4343 vdd.n2546 vdd.n2544 10.6151
R4344 vdd.n2544 vdd.n2543 10.6151
R4345 vdd.n2543 vdd.n2541 10.6151
R4346 vdd.n2541 vdd.n2540 10.6151
R4347 vdd.n2540 vdd.n2538 10.6151
R4348 vdd.n2538 vdd.n2537 10.6151
R4349 vdd.n2537 vdd.n2535 10.6151
R4350 vdd.n2535 vdd.n2534 10.6151
R4351 vdd.n2534 vdd.n2532 10.6151
R4352 vdd.n2532 vdd.n2531 10.6151
R4353 vdd.n2531 vdd.n2529 10.6151
R4354 vdd.n2529 vdd.n2528 10.6151
R4355 vdd.n2528 vdd.n2526 10.6151
R4356 vdd.n2526 vdd.n2525 10.6151
R4357 vdd.n2525 vdd.n2523 10.6151
R4358 vdd.n2523 vdd.n2522 10.6151
R4359 vdd.n2522 vdd.n592 10.6151
R4360 vdd.n2378 vdd.n732 10.6151
R4361 vdd.n2381 vdd.n2378 10.6151
R4362 vdd.n2382 vdd.n2381 10.6151
R4363 vdd.n2385 vdd.n2382 10.6151
R4364 vdd.n2386 vdd.n2385 10.6151
R4365 vdd.n2389 vdd.n2386 10.6151
R4366 vdd.n2390 vdd.n2389 10.6151
R4367 vdd.n2393 vdd.n2390 10.6151
R4368 vdd.n2394 vdd.n2393 10.6151
R4369 vdd.n2397 vdd.n2394 10.6151
R4370 vdd.n2398 vdd.n2397 10.6151
R4371 vdd.n2401 vdd.n2398 10.6151
R4372 vdd.n2402 vdd.n2401 10.6151
R4373 vdd.n2405 vdd.n2402 10.6151
R4374 vdd.n2406 vdd.n2405 10.6151
R4375 vdd.n2409 vdd.n2406 10.6151
R4376 vdd.n2410 vdd.n2409 10.6151
R4377 vdd.n2413 vdd.n2410 10.6151
R4378 vdd.n2414 vdd.n2413 10.6151
R4379 vdd.n2417 vdd.n2414 10.6151
R4380 vdd.n2418 vdd.n2417 10.6151
R4381 vdd.n2421 vdd.n2418 10.6151
R4382 vdd.n2422 vdd.n2421 10.6151
R4383 vdd.n2425 vdd.n2422 10.6151
R4384 vdd.n2426 vdd.n2425 10.6151
R4385 vdd.n2429 vdd.n2426 10.6151
R4386 vdd.n2430 vdd.n2429 10.6151
R4387 vdd.n2433 vdd.n2430 10.6151
R4388 vdd.n2434 vdd.n2433 10.6151
R4389 vdd.n2437 vdd.n2434 10.6151
R4390 vdd.n2438 vdd.n2437 10.6151
R4391 vdd.n2442 vdd.n2441 10.6151
R4392 vdd.n2622 vdd.n2442 10.6151
R4393 vdd.n2634 vdd.n2633 10.6151
R4394 vdd.n2635 vdd.n2634 10.6151
R4395 vdd.n2635 vdd.n722 10.6151
R4396 vdd.n2645 vdd.n722 10.6151
R4397 vdd.n2646 vdd.n2645 10.6151
R4398 vdd.n2647 vdd.n2646 10.6151
R4399 vdd.n2647 vdd.n710 10.6151
R4400 vdd.n2657 vdd.n710 10.6151
R4401 vdd.n2658 vdd.n2657 10.6151
R4402 vdd.n2659 vdd.n2658 10.6151
R4403 vdd.n2659 vdd.n699 10.6151
R4404 vdd.n2669 vdd.n699 10.6151
R4405 vdd.n2670 vdd.n2669 10.6151
R4406 vdd.n2671 vdd.n2670 10.6151
R4407 vdd.n2671 vdd.n687 10.6151
R4408 vdd.n2681 vdd.n687 10.6151
R4409 vdd.n2682 vdd.n2681 10.6151
R4410 vdd.n2683 vdd.n2682 10.6151
R4411 vdd.n2683 vdd.n676 10.6151
R4412 vdd.n2693 vdd.n676 10.6151
R4413 vdd.n2696 vdd.n2695 10.6151
R4414 vdd.n2696 vdd.n662 10.6151
R4415 vdd.n2706 vdd.n662 10.6151
R4416 vdd.n2707 vdd.n2706 10.6151
R4417 vdd.n2708 vdd.n2707 10.6151
R4418 vdd.n2708 vdd.n650 10.6151
R4419 vdd.n2718 vdd.n650 10.6151
R4420 vdd.n2719 vdd.n2718 10.6151
R4421 vdd.n2720 vdd.n2719 10.6151
R4422 vdd.n2720 vdd.n639 10.6151
R4423 vdd.n2730 vdd.n639 10.6151
R4424 vdd.n2731 vdd.n2730 10.6151
R4425 vdd.n2777 vdd.n2731 10.6151
R4426 vdd.n2777 vdd.n2776 10.6151
R4427 vdd.n2776 vdd.n2775 10.6151
R4428 vdd.n2775 vdd.n2774 10.6151
R4429 vdd.n2774 vdd.n2772 10.6151
R4430 vdd.n2084 vdd.n2083 10.6151
R4431 vdd.n2085 vdd.n2084 10.6151
R4432 vdd.n2085 vdd.n886 10.6151
R4433 vdd.n2095 vdd.n886 10.6151
R4434 vdd.n2096 vdd.n2095 10.6151
R4435 vdd.n2097 vdd.n2096 10.6151
R4436 vdd.n2097 vdd.n874 10.6151
R4437 vdd.n2107 vdd.n874 10.6151
R4438 vdd.n2108 vdd.n2107 10.6151
R4439 vdd.n2109 vdd.n2108 10.6151
R4440 vdd.n2109 vdd.n862 10.6151
R4441 vdd.n2119 vdd.n862 10.6151
R4442 vdd.n2120 vdd.n2119 10.6151
R4443 vdd.n2121 vdd.n2120 10.6151
R4444 vdd.n2121 vdd.n849 10.6151
R4445 vdd.n2131 vdd.n849 10.6151
R4446 vdd.n2132 vdd.n2131 10.6151
R4447 vdd.n2134 vdd.n837 10.6151
R4448 vdd.n2144 vdd.n837 10.6151
R4449 vdd.n2145 vdd.n2144 10.6151
R4450 vdd.n2146 vdd.n2145 10.6151
R4451 vdd.n2146 vdd.n825 10.6151
R4452 vdd.n2156 vdd.n825 10.6151
R4453 vdd.n2157 vdd.n2156 10.6151
R4454 vdd.n2158 vdd.n2157 10.6151
R4455 vdd.n2158 vdd.n814 10.6151
R4456 vdd.n2168 vdd.n814 10.6151
R4457 vdd.n2169 vdd.n2168 10.6151
R4458 vdd.n2170 vdd.n2169 10.6151
R4459 vdd.n2170 vdd.n803 10.6151
R4460 vdd.n2180 vdd.n803 10.6151
R4461 vdd.n2181 vdd.n2180 10.6151
R4462 vdd.n2184 vdd.n2181 10.6151
R4463 vdd.n2184 vdd.n2183 10.6151
R4464 vdd.n2183 vdd.n2182 10.6151
R4465 vdd.n2182 vdd.n786 10.6151
R4466 vdd.n2266 vdd.n786 10.6151
R4467 vdd.n2265 vdd.n2264 10.6151
R4468 vdd.n2264 vdd.n2261 10.6151
R4469 vdd.n2261 vdd.n2260 10.6151
R4470 vdd.n2260 vdd.n2257 10.6151
R4471 vdd.n2257 vdd.n2256 10.6151
R4472 vdd.n2256 vdd.n2253 10.6151
R4473 vdd.n2253 vdd.n2252 10.6151
R4474 vdd.n2252 vdd.n2249 10.6151
R4475 vdd.n2249 vdd.n2248 10.6151
R4476 vdd.n2248 vdd.n2245 10.6151
R4477 vdd.n2245 vdd.n2244 10.6151
R4478 vdd.n2244 vdd.n2241 10.6151
R4479 vdd.n2241 vdd.n2240 10.6151
R4480 vdd.n2240 vdd.n2237 10.6151
R4481 vdd.n2237 vdd.n2236 10.6151
R4482 vdd.n2236 vdd.n2233 10.6151
R4483 vdd.n2233 vdd.n2232 10.6151
R4484 vdd.n2232 vdd.n2229 10.6151
R4485 vdd.n2229 vdd.n2228 10.6151
R4486 vdd.n2228 vdd.n2225 10.6151
R4487 vdd.n2225 vdd.n2224 10.6151
R4488 vdd.n2224 vdd.n2221 10.6151
R4489 vdd.n2221 vdd.n2220 10.6151
R4490 vdd.n2220 vdd.n2217 10.6151
R4491 vdd.n2217 vdd.n2216 10.6151
R4492 vdd.n2216 vdd.n2213 10.6151
R4493 vdd.n2213 vdd.n2212 10.6151
R4494 vdd.n2212 vdd.n2209 10.6151
R4495 vdd.n2209 vdd.n2208 10.6151
R4496 vdd.n2208 vdd.n2205 10.6151
R4497 vdd.n2205 vdd.n2204 10.6151
R4498 vdd.n2201 vdd.n2200 10.6151
R4499 vdd.n2200 vdd.n2198 10.6151
R4500 vdd.n1900 vdd.n1898 10.6151
R4501 vdd.n1901 vdd.n1900 10.6151
R4502 vdd.n1903 vdd.n1901 10.6151
R4503 vdd.n1904 vdd.n1903 10.6151
R4504 vdd.n1906 vdd.n1904 10.6151
R4505 vdd.n1907 vdd.n1906 10.6151
R4506 vdd.n1909 vdd.n1907 10.6151
R4507 vdd.n1910 vdd.n1909 10.6151
R4508 vdd.n1912 vdd.n1910 10.6151
R4509 vdd.n1913 vdd.n1912 10.6151
R4510 vdd.n1915 vdd.n1913 10.6151
R4511 vdd.n1916 vdd.n1915 10.6151
R4512 vdd.n1918 vdd.n1916 10.6151
R4513 vdd.n1919 vdd.n1918 10.6151
R4514 vdd.n1921 vdd.n1919 10.6151
R4515 vdd.n1922 vdd.n1921 10.6151
R4516 vdd.n1924 vdd.n1922 10.6151
R4517 vdd.n1925 vdd.n1924 10.6151
R4518 vdd.n1927 vdd.n1925 10.6151
R4519 vdd.n1928 vdd.n1927 10.6151
R4520 vdd.n1930 vdd.n1928 10.6151
R4521 vdd.n1931 vdd.n1930 10.6151
R4522 vdd.n1970 vdd.n1931 10.6151
R4523 vdd.n1970 vdd.n1969 10.6151
R4524 vdd.n1969 vdd.n1968 10.6151
R4525 vdd.n1968 vdd.n1966 10.6151
R4526 vdd.n1966 vdd.n1965 10.6151
R4527 vdd.n1965 vdd.n1963 10.6151
R4528 vdd.n1963 vdd.n1962 10.6151
R4529 vdd.n1962 vdd.n1939 10.6151
R4530 vdd.n1939 vdd.n1938 10.6151
R4531 vdd.n1938 vdd.n1936 10.6151
R4532 vdd.n1936 vdd.n1935 10.6151
R4533 vdd.n1935 vdd.n1933 10.6151
R4534 vdd.n1933 vdd.n1932 10.6151
R4535 vdd.n1932 vdd.n790 10.6151
R4536 vdd.n2196 vdd.n790 10.6151
R4537 vdd.n2197 vdd.n2196 10.6151
R4538 vdd.n1828 vdd.n898 10.6151
R4539 vdd.n1833 vdd.n1828 10.6151
R4540 vdd.n1834 vdd.n1833 10.6151
R4541 vdd.n1835 vdd.n1834 10.6151
R4542 vdd.n1835 vdd.n1826 10.6151
R4543 vdd.n1841 vdd.n1826 10.6151
R4544 vdd.n1842 vdd.n1841 10.6151
R4545 vdd.n1843 vdd.n1842 10.6151
R4546 vdd.n1843 vdd.n1824 10.6151
R4547 vdd.n1849 vdd.n1824 10.6151
R4548 vdd.n1850 vdd.n1849 10.6151
R4549 vdd.n1851 vdd.n1850 10.6151
R4550 vdd.n1851 vdd.n1822 10.6151
R4551 vdd.n1857 vdd.n1822 10.6151
R4552 vdd.n1858 vdd.n1857 10.6151
R4553 vdd.n1859 vdd.n1858 10.6151
R4554 vdd.n1859 vdd.n1820 10.6151
R4555 vdd.n1865 vdd.n1820 10.6151
R4556 vdd.n1866 vdd.n1865 10.6151
R4557 vdd.n1867 vdd.n1866 10.6151
R4558 vdd.n1867 vdd.n932 10.6151
R4559 vdd.n1873 vdd.n932 10.6151
R4560 vdd.n1874 vdd.n1873 10.6151
R4561 vdd.n1875 vdd.n1874 10.6151
R4562 vdd.n1875 vdd.n930 10.6151
R4563 vdd.n1881 vdd.n930 10.6151
R4564 vdd.n1882 vdd.n1881 10.6151
R4565 vdd.n1883 vdd.n1882 10.6151
R4566 vdd.n1883 vdd.n928 10.6151
R4567 vdd.n1889 vdd.n928 10.6151
R4568 vdd.n1890 vdd.n1889 10.6151
R4569 vdd.n1892 vdd.n924 10.6151
R4570 vdd.n1897 vdd.n924 10.6151
R4571 vdd.n280 vdd.n262 10.4732
R4572 vdd.n233 vdd.n215 10.4732
R4573 vdd.n190 vdd.n172 10.4732
R4574 vdd.n143 vdd.n125 10.4732
R4575 vdd.n101 vdd.n83 10.4732
R4576 vdd.n54 vdd.n36 10.4732
R4577 vdd.n1175 vdd.n1157 10.4732
R4578 vdd.n1222 vdd.n1204 10.4732
R4579 vdd.n1085 vdd.n1067 10.4732
R4580 vdd.n1132 vdd.n1114 10.4732
R4581 vdd.n996 vdd.n978 10.4732
R4582 vdd.n1043 vdd.n1025 10.4732
R4583 vdd.t0 vdd.n968 10.3167
R4584 vdd.n3056 vdd.t24 10.3167
R4585 vdd.n2268 vdd.t191 10.2034
R4586 vdd.n2631 vdd.t179 10.2034
R4587 vdd.n1545 vdd.t12 10.09
R4588 vdd.n3224 vdd.t10 10.09
R4589 vdd.n1796 vdd.n912 9.88581
R4590 vdd.n3018 vdd.n520 9.88581
R4591 vdd.n2889 vdd.n2888 9.88581
R4592 vdd.n1820 vdd.n1819 9.88581
R4593 vdd.n279 vdd.n264 9.69747
R4594 vdd.n232 vdd.n217 9.69747
R4595 vdd.n189 vdd.n174 9.69747
R4596 vdd.n142 vdd.n127 9.69747
R4597 vdd.n100 vdd.n85 9.69747
R4598 vdd.n53 vdd.n38 9.69747
R4599 vdd.n1174 vdd.n1159 9.69747
R4600 vdd.n1221 vdd.n1206 9.69747
R4601 vdd.n1084 vdd.n1069 9.69747
R4602 vdd.n1131 vdd.n1116 9.69747
R4603 vdd.n995 vdd.n980 9.69747
R4604 vdd.n1042 vdd.n1027 9.69747
R4605 vdd.n295 vdd.n294 9.45567
R4606 vdd.n248 vdd.n247 9.45567
R4607 vdd.n205 vdd.n204 9.45567
R4608 vdd.n158 vdd.n157 9.45567
R4609 vdd.n116 vdd.n115 9.45567
R4610 vdd.n69 vdd.n68 9.45567
R4611 vdd.n1190 vdd.n1189 9.45567
R4612 vdd.n1237 vdd.n1236 9.45567
R4613 vdd.n1100 vdd.n1099 9.45567
R4614 vdd.n1147 vdd.n1146 9.45567
R4615 vdd.n1011 vdd.n1010 9.45567
R4616 vdd.n1058 vdd.n1057 9.45567
R4617 vdd.n1769 vdd.n1623 9.3005
R4618 vdd.n1768 vdd.n1767 9.3005
R4619 vdd.n1629 vdd.n1628 9.3005
R4620 vdd.n1762 vdd.n1633 9.3005
R4621 vdd.n1761 vdd.n1634 9.3005
R4622 vdd.n1760 vdd.n1635 9.3005
R4623 vdd.n1639 vdd.n1636 9.3005
R4624 vdd.n1755 vdd.n1640 9.3005
R4625 vdd.n1754 vdd.n1641 9.3005
R4626 vdd.n1753 vdd.n1642 9.3005
R4627 vdd.n1646 vdd.n1643 9.3005
R4628 vdd.n1748 vdd.n1647 9.3005
R4629 vdd.n1747 vdd.n1648 9.3005
R4630 vdd.n1746 vdd.n1649 9.3005
R4631 vdd.n1653 vdd.n1650 9.3005
R4632 vdd.n1741 vdd.n1654 9.3005
R4633 vdd.n1740 vdd.n1655 9.3005
R4634 vdd.n1739 vdd.n1656 9.3005
R4635 vdd.n1660 vdd.n1657 9.3005
R4636 vdd.n1734 vdd.n1661 9.3005
R4637 vdd.n1733 vdd.n1662 9.3005
R4638 vdd.n1732 vdd.n1731 9.3005
R4639 vdd.n1730 vdd.n1663 9.3005
R4640 vdd.n1729 vdd.n1728 9.3005
R4641 vdd.n1669 vdd.n1668 9.3005
R4642 vdd.n1723 vdd.n1673 9.3005
R4643 vdd.n1722 vdd.n1674 9.3005
R4644 vdd.n1721 vdd.n1675 9.3005
R4645 vdd.n1679 vdd.n1676 9.3005
R4646 vdd.n1716 vdd.n1680 9.3005
R4647 vdd.n1715 vdd.n1681 9.3005
R4648 vdd.n1714 vdd.n1682 9.3005
R4649 vdd.n1686 vdd.n1683 9.3005
R4650 vdd.n1709 vdd.n1687 9.3005
R4651 vdd.n1708 vdd.n1688 9.3005
R4652 vdd.n1707 vdd.n1689 9.3005
R4653 vdd.n1691 vdd.n1690 9.3005
R4654 vdd.n1702 vdd.n934 9.3005
R4655 vdd.n1771 vdd.n1770 9.3005
R4656 vdd.n1795 vdd.n1794 9.3005
R4657 vdd.n1601 vdd.n1600 9.3005
R4658 vdd.n1606 vdd.n1604 9.3005
R4659 vdd.n1787 vdd.n1607 9.3005
R4660 vdd.n1786 vdd.n1608 9.3005
R4661 vdd.n1785 vdd.n1609 9.3005
R4662 vdd.n1613 vdd.n1610 9.3005
R4663 vdd.n1780 vdd.n1614 9.3005
R4664 vdd.n1779 vdd.n1615 9.3005
R4665 vdd.n1778 vdd.n1616 9.3005
R4666 vdd.n1620 vdd.n1617 9.3005
R4667 vdd.n1773 vdd.n1621 9.3005
R4668 vdd.n1772 vdd.n1622 9.3005
R4669 vdd.n1804 vdd.n1594 9.3005
R4670 vdd.n1806 vdd.n1805 9.3005
R4671 vdd.n1556 vdd.n1555 9.3005
R4672 vdd.n1557 vdd.n970 9.3005
R4673 vdd.n1559 vdd.n1558 9.3005
R4674 vdd.n960 vdd.n959 9.3005
R4675 vdd.n1573 vdd.n1572 9.3005
R4676 vdd.n1574 vdd.n958 9.3005
R4677 vdd.n1576 vdd.n1575 9.3005
R4678 vdd.n948 vdd.n947 9.3005
R4679 vdd.n1592 vdd.n1591 9.3005
R4680 vdd.n1593 vdd.n946 9.3005
R4681 vdd.n1808 vdd.n1807 9.3005
R4682 vdd.n271 vdd.n270 9.3005
R4683 vdd.n266 vdd.n265 9.3005
R4684 vdd.n277 vdd.n276 9.3005
R4685 vdd.n279 vdd.n278 9.3005
R4686 vdd.n262 vdd.n261 9.3005
R4687 vdd.n285 vdd.n284 9.3005
R4688 vdd.n287 vdd.n286 9.3005
R4689 vdd.n259 vdd.n256 9.3005
R4690 vdd.n294 vdd.n293 9.3005
R4691 vdd.n224 vdd.n223 9.3005
R4692 vdd.n219 vdd.n218 9.3005
R4693 vdd.n230 vdd.n229 9.3005
R4694 vdd.n232 vdd.n231 9.3005
R4695 vdd.n215 vdd.n214 9.3005
R4696 vdd.n238 vdd.n237 9.3005
R4697 vdd.n240 vdd.n239 9.3005
R4698 vdd.n212 vdd.n209 9.3005
R4699 vdd.n247 vdd.n246 9.3005
R4700 vdd.n181 vdd.n180 9.3005
R4701 vdd.n176 vdd.n175 9.3005
R4702 vdd.n187 vdd.n186 9.3005
R4703 vdd.n189 vdd.n188 9.3005
R4704 vdd.n172 vdd.n171 9.3005
R4705 vdd.n195 vdd.n194 9.3005
R4706 vdd.n197 vdd.n196 9.3005
R4707 vdd.n169 vdd.n166 9.3005
R4708 vdd.n204 vdd.n203 9.3005
R4709 vdd.n134 vdd.n133 9.3005
R4710 vdd.n129 vdd.n128 9.3005
R4711 vdd.n140 vdd.n139 9.3005
R4712 vdd.n142 vdd.n141 9.3005
R4713 vdd.n125 vdd.n124 9.3005
R4714 vdd.n148 vdd.n147 9.3005
R4715 vdd.n150 vdd.n149 9.3005
R4716 vdd.n122 vdd.n119 9.3005
R4717 vdd.n157 vdd.n156 9.3005
R4718 vdd.n92 vdd.n91 9.3005
R4719 vdd.n87 vdd.n86 9.3005
R4720 vdd.n98 vdd.n97 9.3005
R4721 vdd.n100 vdd.n99 9.3005
R4722 vdd.n83 vdd.n82 9.3005
R4723 vdd.n106 vdd.n105 9.3005
R4724 vdd.n108 vdd.n107 9.3005
R4725 vdd.n80 vdd.n77 9.3005
R4726 vdd.n115 vdd.n114 9.3005
R4727 vdd.n45 vdd.n44 9.3005
R4728 vdd.n40 vdd.n39 9.3005
R4729 vdd.n51 vdd.n50 9.3005
R4730 vdd.n53 vdd.n52 9.3005
R4731 vdd.n36 vdd.n35 9.3005
R4732 vdd.n59 vdd.n58 9.3005
R4733 vdd.n61 vdd.n60 9.3005
R4734 vdd.n33 vdd.n30 9.3005
R4735 vdd.n68 vdd.n67 9.3005
R4736 vdd.n2940 vdd.n2939 9.3005
R4737 vdd.n2943 vdd.n555 9.3005
R4738 vdd.n2944 vdd.n554 9.3005
R4739 vdd.n2947 vdd.n553 9.3005
R4740 vdd.n2948 vdd.n552 9.3005
R4741 vdd.n2951 vdd.n551 9.3005
R4742 vdd.n2952 vdd.n550 9.3005
R4743 vdd.n2955 vdd.n549 9.3005
R4744 vdd.n2956 vdd.n548 9.3005
R4745 vdd.n2959 vdd.n547 9.3005
R4746 vdd.n2960 vdd.n546 9.3005
R4747 vdd.n2963 vdd.n545 9.3005
R4748 vdd.n2964 vdd.n544 9.3005
R4749 vdd.n2967 vdd.n543 9.3005
R4750 vdd.n2968 vdd.n542 9.3005
R4751 vdd.n2971 vdd.n541 9.3005
R4752 vdd.n2972 vdd.n540 9.3005
R4753 vdd.n2975 vdd.n539 9.3005
R4754 vdd.n2976 vdd.n538 9.3005
R4755 vdd.n2979 vdd.n537 9.3005
R4756 vdd.n2983 vdd.n2982 9.3005
R4757 vdd.n2984 vdd.n536 9.3005
R4758 vdd.n2988 vdd.n2985 9.3005
R4759 vdd.n2991 vdd.n535 9.3005
R4760 vdd.n2992 vdd.n534 9.3005
R4761 vdd.n2995 vdd.n533 9.3005
R4762 vdd.n2996 vdd.n532 9.3005
R4763 vdd.n2999 vdd.n531 9.3005
R4764 vdd.n3000 vdd.n530 9.3005
R4765 vdd.n3003 vdd.n529 9.3005
R4766 vdd.n3004 vdd.n528 9.3005
R4767 vdd.n3007 vdd.n527 9.3005
R4768 vdd.n3008 vdd.n526 9.3005
R4769 vdd.n3011 vdd.n525 9.3005
R4770 vdd.n3012 vdd.n524 9.3005
R4771 vdd.n3015 vdd.n519 9.3005
R4772 vdd.n482 vdd.n481 9.3005
R4773 vdd.n3026 vdd.n3025 9.3005
R4774 vdd.n3029 vdd.n3028 9.3005
R4775 vdd.n471 vdd.n470 9.3005
R4776 vdd.n3043 vdd.n3042 9.3005
R4777 vdd.n3044 vdd.n469 9.3005
R4778 vdd.n3046 vdd.n3045 9.3005
R4779 vdd.n460 vdd.n459 9.3005
R4780 vdd.n3059 vdd.n3058 9.3005
R4781 vdd.n3060 vdd.n458 9.3005
R4782 vdd.n3062 vdd.n3061 9.3005
R4783 vdd.n300 vdd.n298 9.3005
R4784 vdd.n3027 vdd.n480 9.3005
R4785 vdd.n3228 vdd.n3227 9.3005
R4786 vdd.n301 vdd.n299 9.3005
R4787 vdd.n3221 vdd.n310 9.3005
R4788 vdd.n3220 vdd.n311 9.3005
R4789 vdd.n3219 vdd.n312 9.3005
R4790 vdd.n320 vdd.n313 9.3005
R4791 vdd.n3213 vdd.n321 9.3005
R4792 vdd.n3212 vdd.n322 9.3005
R4793 vdd.n3211 vdd.n323 9.3005
R4794 vdd.n331 vdd.n324 9.3005
R4795 vdd.n3205 vdd.n3204 9.3005
R4796 vdd.n3201 vdd.n332 9.3005
R4797 vdd.n3200 vdd.n335 9.3005
R4798 vdd.n339 vdd.n336 9.3005
R4799 vdd.n340 vdd.n337 9.3005
R4800 vdd.n3193 vdd.n341 9.3005
R4801 vdd.n3192 vdd.n342 9.3005
R4802 vdd.n3191 vdd.n343 9.3005
R4803 vdd.n347 vdd.n344 9.3005
R4804 vdd.n3186 vdd.n348 9.3005
R4805 vdd.n3185 vdd.n349 9.3005
R4806 vdd.n3184 vdd.n350 9.3005
R4807 vdd.n354 vdd.n351 9.3005
R4808 vdd.n3179 vdd.n355 9.3005
R4809 vdd.n3178 vdd.n356 9.3005
R4810 vdd.n3177 vdd.n357 9.3005
R4811 vdd.n361 vdd.n358 9.3005
R4812 vdd.n3172 vdd.n362 9.3005
R4813 vdd.n3171 vdd.n363 9.3005
R4814 vdd.n3170 vdd.n3169 9.3005
R4815 vdd.n3168 vdd.n364 9.3005
R4816 vdd.n3167 vdd.n3166 9.3005
R4817 vdd.n370 vdd.n369 9.3005
R4818 vdd.n3161 vdd.n374 9.3005
R4819 vdd.n3160 vdd.n375 9.3005
R4820 vdd.n3159 vdd.n376 9.3005
R4821 vdd.n380 vdd.n377 9.3005
R4822 vdd.n3154 vdd.n381 9.3005
R4823 vdd.n3153 vdd.n382 9.3005
R4824 vdd.n3152 vdd.n383 9.3005
R4825 vdd.n387 vdd.n384 9.3005
R4826 vdd.n3147 vdd.n388 9.3005
R4827 vdd.n3146 vdd.n389 9.3005
R4828 vdd.n3145 vdd.n390 9.3005
R4829 vdd.n394 vdd.n391 9.3005
R4830 vdd.n3140 vdd.n395 9.3005
R4831 vdd.n3139 vdd.n396 9.3005
R4832 vdd.n3138 vdd.n397 9.3005
R4833 vdd.n401 vdd.n398 9.3005
R4834 vdd.n3133 vdd.n402 9.3005
R4835 vdd.n3132 vdd.n403 9.3005
R4836 vdd.n3131 vdd.n3130 9.3005
R4837 vdd.n3129 vdd.n404 9.3005
R4838 vdd.n3128 vdd.n3127 9.3005
R4839 vdd.n410 vdd.n409 9.3005
R4840 vdd.n3122 vdd.n414 9.3005
R4841 vdd.n3121 vdd.n415 9.3005
R4842 vdd.n3120 vdd.n416 9.3005
R4843 vdd.n420 vdd.n417 9.3005
R4844 vdd.n3115 vdd.n421 9.3005
R4845 vdd.n3114 vdd.n422 9.3005
R4846 vdd.n3113 vdd.n423 9.3005
R4847 vdd.n427 vdd.n424 9.3005
R4848 vdd.n3108 vdd.n428 9.3005
R4849 vdd.n3107 vdd.n429 9.3005
R4850 vdd.n3106 vdd.n430 9.3005
R4851 vdd.n434 vdd.n431 9.3005
R4852 vdd.n3101 vdd.n435 9.3005
R4853 vdd.n3100 vdd.n436 9.3005
R4854 vdd.n3099 vdd.n437 9.3005
R4855 vdd.n441 vdd.n438 9.3005
R4856 vdd.n3094 vdd.n442 9.3005
R4857 vdd.n3093 vdd.n443 9.3005
R4858 vdd.n3089 vdd.n3086 9.3005
R4859 vdd.n3203 vdd.n3202 9.3005
R4860 vdd.n3034 vdd.n3033 9.3005
R4861 vdd.n3035 vdd.n475 9.3005
R4862 vdd.n3037 vdd.n3036 9.3005
R4863 vdd.n465 vdd.n464 9.3005
R4864 vdd.n3051 vdd.n3050 9.3005
R4865 vdd.n3052 vdd.n463 9.3005
R4866 vdd.n3054 vdd.n3053 9.3005
R4867 vdd.n453 vdd.n452 9.3005
R4868 vdd.n3067 vdd.n3066 9.3005
R4869 vdd.n3068 vdd.n451 9.3005
R4870 vdd.n3070 vdd.n3069 9.3005
R4871 vdd.n3071 vdd.n450 9.3005
R4872 vdd.n3073 vdd.n3072 9.3005
R4873 vdd.n3074 vdd.n449 9.3005
R4874 vdd.n3076 vdd.n3075 9.3005
R4875 vdd.n3077 vdd.n447 9.3005
R4876 vdd.n3079 vdd.n3078 9.3005
R4877 vdd.n3080 vdd.n446 9.3005
R4878 vdd.n3082 vdd.n3081 9.3005
R4879 vdd.n3083 vdd.n444 9.3005
R4880 vdd.n3085 vdd.n3084 9.3005
R4881 vdd.n477 vdd.n476 9.3005
R4882 vdd.n2892 vdd.n2891 9.3005
R4883 vdd.n2897 vdd.n2890 9.3005
R4884 vdd.n2906 vdd.n572 9.3005
R4885 vdd.n2909 vdd.n571 9.3005
R4886 vdd.n2910 vdd.n570 9.3005
R4887 vdd.n2913 vdd.n569 9.3005
R4888 vdd.n2914 vdd.n568 9.3005
R4889 vdd.n2917 vdd.n567 9.3005
R4890 vdd.n2918 vdd.n566 9.3005
R4891 vdd.n2921 vdd.n565 9.3005
R4892 vdd.n2922 vdd.n564 9.3005
R4893 vdd.n2925 vdd.n563 9.3005
R4894 vdd.n2926 vdd.n562 9.3005
R4895 vdd.n2929 vdd.n561 9.3005
R4896 vdd.n2930 vdd.n560 9.3005
R4897 vdd.n2933 vdd.n559 9.3005
R4898 vdd.n2937 vdd.n2936 9.3005
R4899 vdd.n2938 vdd.n556 9.3005
R4900 vdd.n1818 vdd.n1817 9.3005
R4901 vdd.n1813 vdd.n937 9.3005
R4902 vdd.n1513 vdd.n1512 9.3005
R4903 vdd.n1514 vdd.n1268 9.3005
R4904 vdd.n1516 vdd.n1515 9.3005
R4905 vdd.n1258 vdd.n1257 9.3005
R4906 vdd.n1530 vdd.n1529 9.3005
R4907 vdd.n1531 vdd.n1256 9.3005
R4908 vdd.n1533 vdd.n1532 9.3005
R4909 vdd.n1248 vdd.n1247 9.3005
R4910 vdd.n1548 vdd.n1547 9.3005
R4911 vdd.n1549 vdd.n1246 9.3005
R4912 vdd.n1551 vdd.n1550 9.3005
R4913 vdd.n965 vdd.n964 9.3005
R4914 vdd.n1564 vdd.n1563 9.3005
R4915 vdd.n1565 vdd.n963 9.3005
R4916 vdd.n1567 vdd.n1566 9.3005
R4917 vdd.n955 vdd.n954 9.3005
R4918 vdd.n1581 vdd.n1580 9.3005
R4919 vdd.n1582 vdd.n952 9.3005
R4920 vdd.n1586 vdd.n1585 9.3005
R4921 vdd.n1584 vdd.n953 9.3005
R4922 vdd.n1583 vdd.n942 9.3005
R4923 vdd.n1270 vdd.n1269 9.3005
R4924 vdd.n1406 vdd.n1405 9.3005
R4925 vdd.n1407 vdd.n1396 9.3005
R4926 vdd.n1409 vdd.n1408 9.3005
R4927 vdd.n1410 vdd.n1395 9.3005
R4928 vdd.n1412 vdd.n1411 9.3005
R4929 vdd.n1413 vdd.n1390 9.3005
R4930 vdd.n1415 vdd.n1414 9.3005
R4931 vdd.n1416 vdd.n1389 9.3005
R4932 vdd.n1418 vdd.n1417 9.3005
R4933 vdd.n1419 vdd.n1384 9.3005
R4934 vdd.n1421 vdd.n1420 9.3005
R4935 vdd.n1422 vdd.n1383 9.3005
R4936 vdd.n1424 vdd.n1423 9.3005
R4937 vdd.n1425 vdd.n1378 9.3005
R4938 vdd.n1427 vdd.n1426 9.3005
R4939 vdd.n1428 vdd.n1377 9.3005
R4940 vdd.n1430 vdd.n1429 9.3005
R4941 vdd.n1431 vdd.n1372 9.3005
R4942 vdd.n1433 vdd.n1432 9.3005
R4943 vdd.n1434 vdd.n1371 9.3005
R4944 vdd.n1436 vdd.n1435 9.3005
R4945 vdd.n1440 vdd.n1367 9.3005
R4946 vdd.n1442 vdd.n1441 9.3005
R4947 vdd.n1443 vdd.n1366 9.3005
R4948 vdd.n1445 vdd.n1444 9.3005
R4949 vdd.n1446 vdd.n1361 9.3005
R4950 vdd.n1448 vdd.n1447 9.3005
R4951 vdd.n1449 vdd.n1360 9.3005
R4952 vdd.n1451 vdd.n1450 9.3005
R4953 vdd.n1452 vdd.n1355 9.3005
R4954 vdd.n1454 vdd.n1453 9.3005
R4955 vdd.n1455 vdd.n1354 9.3005
R4956 vdd.n1457 vdd.n1456 9.3005
R4957 vdd.n1458 vdd.n1349 9.3005
R4958 vdd.n1460 vdd.n1459 9.3005
R4959 vdd.n1461 vdd.n1348 9.3005
R4960 vdd.n1463 vdd.n1462 9.3005
R4961 vdd.n1464 vdd.n1343 9.3005
R4962 vdd.n1466 vdd.n1465 9.3005
R4963 vdd.n1467 vdd.n1342 9.3005
R4964 vdd.n1469 vdd.n1468 9.3005
R4965 vdd.n1470 vdd.n1337 9.3005
R4966 vdd.n1472 vdd.n1471 9.3005
R4967 vdd.n1473 vdd.n1336 9.3005
R4968 vdd.n1475 vdd.n1474 9.3005
R4969 vdd.n1476 vdd.n1329 9.3005
R4970 vdd.n1478 vdd.n1477 9.3005
R4971 vdd.n1479 vdd.n1328 9.3005
R4972 vdd.n1481 vdd.n1480 9.3005
R4973 vdd.n1482 vdd.n1323 9.3005
R4974 vdd.n1484 vdd.n1483 9.3005
R4975 vdd.n1485 vdd.n1322 9.3005
R4976 vdd.n1487 vdd.n1486 9.3005
R4977 vdd.n1488 vdd.n1317 9.3005
R4978 vdd.n1490 vdd.n1489 9.3005
R4979 vdd.n1491 vdd.n1316 9.3005
R4980 vdd.n1493 vdd.n1492 9.3005
R4981 vdd.n1494 vdd.n1311 9.3005
R4982 vdd.n1496 vdd.n1495 9.3005
R4983 vdd.n1497 vdd.n1310 9.3005
R4984 vdd.n1499 vdd.n1498 9.3005
R4985 vdd.n1275 vdd.n1274 9.3005
R4986 vdd.n1505 vdd.n1504 9.3005
R4987 vdd.n1404 vdd.n1403 9.3005
R4988 vdd.n1508 vdd.n1507 9.3005
R4989 vdd.n1264 vdd.n1263 9.3005
R4990 vdd.n1522 vdd.n1521 9.3005
R4991 vdd.n1523 vdd.n1262 9.3005
R4992 vdd.n1525 vdd.n1524 9.3005
R4993 vdd.n1253 vdd.n1252 9.3005
R4994 vdd.n1539 vdd.n1538 9.3005
R4995 vdd.n1540 vdd.n1251 9.3005
R4996 vdd.n1543 vdd.n1542 9.3005
R4997 vdd.n1541 vdd.n1242 9.3005
R4998 vdd.n1506 vdd.n1273 9.3005
R4999 vdd.n1166 vdd.n1165 9.3005
R5000 vdd.n1161 vdd.n1160 9.3005
R5001 vdd.n1172 vdd.n1171 9.3005
R5002 vdd.n1174 vdd.n1173 9.3005
R5003 vdd.n1157 vdd.n1156 9.3005
R5004 vdd.n1180 vdd.n1179 9.3005
R5005 vdd.n1182 vdd.n1181 9.3005
R5006 vdd.n1154 vdd.n1151 9.3005
R5007 vdd.n1189 vdd.n1188 9.3005
R5008 vdd.n1213 vdd.n1212 9.3005
R5009 vdd.n1208 vdd.n1207 9.3005
R5010 vdd.n1219 vdd.n1218 9.3005
R5011 vdd.n1221 vdd.n1220 9.3005
R5012 vdd.n1204 vdd.n1203 9.3005
R5013 vdd.n1227 vdd.n1226 9.3005
R5014 vdd.n1229 vdd.n1228 9.3005
R5015 vdd.n1201 vdd.n1198 9.3005
R5016 vdd.n1236 vdd.n1235 9.3005
R5017 vdd.n1076 vdd.n1075 9.3005
R5018 vdd.n1071 vdd.n1070 9.3005
R5019 vdd.n1082 vdd.n1081 9.3005
R5020 vdd.n1084 vdd.n1083 9.3005
R5021 vdd.n1067 vdd.n1066 9.3005
R5022 vdd.n1090 vdd.n1089 9.3005
R5023 vdd.n1092 vdd.n1091 9.3005
R5024 vdd.n1064 vdd.n1061 9.3005
R5025 vdd.n1099 vdd.n1098 9.3005
R5026 vdd.n1123 vdd.n1122 9.3005
R5027 vdd.n1118 vdd.n1117 9.3005
R5028 vdd.n1129 vdd.n1128 9.3005
R5029 vdd.n1131 vdd.n1130 9.3005
R5030 vdd.n1114 vdd.n1113 9.3005
R5031 vdd.n1137 vdd.n1136 9.3005
R5032 vdd.n1139 vdd.n1138 9.3005
R5033 vdd.n1111 vdd.n1108 9.3005
R5034 vdd.n1146 vdd.n1145 9.3005
R5035 vdd.n987 vdd.n986 9.3005
R5036 vdd.n982 vdd.n981 9.3005
R5037 vdd.n993 vdd.n992 9.3005
R5038 vdd.n995 vdd.n994 9.3005
R5039 vdd.n978 vdd.n977 9.3005
R5040 vdd.n1001 vdd.n1000 9.3005
R5041 vdd.n1003 vdd.n1002 9.3005
R5042 vdd.n975 vdd.n972 9.3005
R5043 vdd.n1010 vdd.n1009 9.3005
R5044 vdd.n1034 vdd.n1033 9.3005
R5045 vdd.n1029 vdd.n1028 9.3005
R5046 vdd.n1040 vdd.n1039 9.3005
R5047 vdd.n1042 vdd.n1041 9.3005
R5048 vdd.n1025 vdd.n1024 9.3005
R5049 vdd.n1048 vdd.n1047 9.3005
R5050 vdd.n1050 vdd.n1049 9.3005
R5051 vdd.n1022 vdd.n1019 9.3005
R5052 vdd.n1057 vdd.n1056 9.3005
R5053 vdd.n1518 vdd.t121 8.95635
R5054 vdd.t8 vdd.n3215 8.95635
R5055 vdd.n276 vdd.n275 8.92171
R5056 vdd.n229 vdd.n228 8.92171
R5057 vdd.n186 vdd.n185 8.92171
R5058 vdd.n139 vdd.n138 8.92171
R5059 vdd.n97 vdd.n96 8.92171
R5060 vdd.n50 vdd.n49 8.92171
R5061 vdd.n1171 vdd.n1170 8.92171
R5062 vdd.n1218 vdd.n1217 8.92171
R5063 vdd.n1081 vdd.n1080 8.92171
R5064 vdd.n1128 vdd.n1127 8.92171
R5065 vdd.n992 vdd.n991 8.92171
R5066 vdd.n1039 vdd.n1038 8.92171
R5067 vdd.n207 vdd.n117 8.81535
R5068 vdd.n1149 vdd.n1059 8.81535
R5069 vdd.n1545 vdd.t106 8.72962
R5070 vdd.t117 vdd.n3224 8.72962
R5071 vdd.n968 vdd.t21 8.50289
R5072 vdd.n1810 vdd.t62 8.50289
R5073 vdd.n516 vdd.t37 8.50289
R5074 vdd.n3056 vdd.t139 8.50289
R5075 vdd.n28 vdd.n14 8.42249
R5076 vdd.n3230 vdd.n3229 8.16225
R5077 vdd.n1241 vdd.n1240 8.16225
R5078 vdd.n272 vdd.n266 8.14595
R5079 vdd.n225 vdd.n219 8.14595
R5080 vdd.n182 vdd.n176 8.14595
R5081 vdd.n135 vdd.n129 8.14595
R5082 vdd.n93 vdd.n87 8.14595
R5083 vdd.n46 vdd.n40 8.14595
R5084 vdd.n1167 vdd.n1161 8.14595
R5085 vdd.n1214 vdd.n1208 8.14595
R5086 vdd.n1077 vdd.n1071 8.14595
R5087 vdd.n1124 vdd.n1118 8.14595
R5088 vdd.n988 vdd.n982 8.14595
R5089 vdd.n1035 vdd.n1029 8.14595
R5090 vdd.n2081 vdd.n894 7.70933
R5091 vdd.n2087 vdd.n894 7.70933
R5092 vdd.n2093 vdd.n888 7.70933
R5093 vdd.n2093 vdd.n882 7.70933
R5094 vdd.n2099 vdd.n882 7.70933
R5095 vdd.n2099 vdd.n876 7.70933
R5096 vdd.n2105 vdd.n876 7.70933
R5097 vdd.n2111 vdd.n870 7.70933
R5098 vdd.n2117 vdd.n864 7.70933
R5099 vdd.n2123 vdd.n857 7.70933
R5100 vdd.n2123 vdd.n860 7.70933
R5101 vdd.n2129 vdd.n853 7.70933
R5102 vdd.n2136 vdd.n839 7.70933
R5103 vdd.n2142 vdd.n839 7.70933
R5104 vdd.n2148 vdd.n833 7.70933
R5105 vdd.n2154 vdd.n829 7.70933
R5106 vdd.n2160 vdd.n823 7.70933
R5107 vdd.n2178 vdd.n805 7.70933
R5108 vdd.n2178 vdd.n798 7.70933
R5109 vdd.n2186 vdd.n798 7.70933
R5110 vdd.n2268 vdd.n782 7.70933
R5111 vdd.n2631 vdd.n736 7.70933
R5112 vdd.n2643 vdd.n717 7.70933
R5113 vdd.n2649 vdd.n717 7.70933
R5114 vdd.n2649 vdd.n720 7.70933
R5115 vdd.n2667 vdd.n701 7.70933
R5116 vdd.n2673 vdd.n695 7.70933
R5117 vdd.n2679 vdd.n691 7.70933
R5118 vdd.n2685 vdd.n678 7.70933
R5119 vdd.n2691 vdd.n678 7.70933
R5120 vdd.n2698 vdd.n671 7.70933
R5121 vdd.n2704 vdd.n664 7.70933
R5122 vdd.n2704 vdd.n667 7.70933
R5123 vdd.n2710 vdd.n660 7.70933
R5124 vdd.n2716 vdd.n654 7.70933
R5125 vdd.n2722 vdd.n641 7.70933
R5126 vdd.n2728 vdd.n641 7.70933
R5127 vdd.n2728 vdd.n633 7.70933
R5128 vdd.n2779 vdd.n633 7.70933
R5129 vdd.n2779 vdd.n636 7.70933
R5130 vdd.n2785 vdd.n595 7.70933
R5131 vdd.n2855 vdd.n595 7.70933
R5132 vdd.t198 vdd.n870 7.59597
R5133 vdd.n1960 vdd.t150 7.59597
R5134 vdd.n2603 vdd.t153 7.59597
R5135 vdd.n654 vdd.t177 7.59597
R5136 vdd.n271 vdd.n268 7.3702
R5137 vdd.n224 vdd.n221 7.3702
R5138 vdd.n181 vdd.n178 7.3702
R5139 vdd.n134 vdd.n131 7.3702
R5140 vdd.n92 vdd.n89 7.3702
R5141 vdd.n45 vdd.n42 7.3702
R5142 vdd.n1166 vdd.n1163 7.3702
R5143 vdd.n1213 vdd.n1210 7.3702
R5144 vdd.n1076 vdd.n1073 7.3702
R5145 vdd.n1123 vdd.n1120 7.3702
R5146 vdd.n987 vdd.n984 7.3702
R5147 vdd.n1034 vdd.n1031 7.3702
R5148 vdd.n1441 vdd.n1440 6.98232
R5149 vdd.n1733 vdd.n1732 6.98232
R5150 vdd.n3132 vdd.n3131 6.98232
R5151 vdd.n2943 vdd.n2940 6.98232
R5152 vdd.n2117 vdd.t161 6.91577
R5153 vdd.n2710 vdd.t186 6.91577
R5154 vdd.n2695 vdd.n2694 6.86879
R5155 vdd.n2133 vdd.n2132 6.86879
R5156 vdd.n2193 vdd.t193 6.80241
R5157 vdd.n2637 vdd.t181 6.80241
R5158 vdd.n1578 vdd.t15 6.68904
R5159 vdd.n3039 vdd.t2 6.68904
R5160 vdd.t6 vdd.n967 6.46231
R5161 vdd.n3064 vdd.t18 6.46231
R5162 vdd.n1960 vdd.t151 6.34895
R5163 vdd.n2603 vdd.t195 6.34895
R5164 vdd.n1536 vdd.t126 6.23558
R5165 vdd.t124 vdd.n308 6.23558
R5166 vdd.n3230 vdd.n297 6.22547
R5167 vdd.n1240 vdd.n1239 6.22547
R5168 vdd.t164 vdd.n833 6.00885
R5169 vdd.n691 vdd.t169 6.00885
R5170 vdd.n272 vdd.n271 5.81868
R5171 vdd.n225 vdd.n224 5.81868
R5172 vdd.n182 vdd.n181 5.81868
R5173 vdd.n135 vdd.n134 5.81868
R5174 vdd.n93 vdd.n92 5.81868
R5175 vdd.n46 vdd.n45 5.81868
R5176 vdd.n1167 vdd.n1166 5.81868
R5177 vdd.n1214 vdd.n1213 5.81868
R5178 vdd.n1077 vdd.n1076 5.81868
R5179 vdd.n1124 vdd.n1123 5.81868
R5180 vdd.n988 vdd.n987 5.81868
R5181 vdd.n1035 vdd.n1034 5.81868
R5182 vdd.n2276 vdd.n2275 5.77611
R5183 vdd.n2016 vdd.n2015 5.77611
R5184 vdd.n2505 vdd.n2504 5.77611
R5185 vdd.n2796 vdd.n2795 5.77611
R5186 vdd.n2860 vdd.n591 5.77611
R5187 vdd.n2441 vdd.n2377 5.77611
R5188 vdd.n2201 vdd.n789 5.77611
R5189 vdd.n1892 vdd.n1891 5.77611
R5190 vdd.n1403 vdd.n1402 5.62474
R5191 vdd.n1816 vdd.n1813 5.62474
R5192 vdd.n3092 vdd.n3089 5.62474
R5193 vdd.n2895 vdd.n2892 5.62474
R5194 vdd.n2154 vdd.t189 5.44203
R5195 vdd.n2673 vdd.t165 5.44203
R5196 vdd.n1260 vdd.t126 5.10193
R5197 vdd.n2129 vdd.t178 5.10193
R5198 vdd.n2148 vdd.t197 5.10193
R5199 vdd.n2679 vdd.t187 5.10193
R5200 vdd.n2698 vdd.t156 5.10193
R5201 vdd.n3217 vdd.t124 5.10193
R5202 vdd.n275 vdd.n266 5.04292
R5203 vdd.n228 vdd.n219 5.04292
R5204 vdd.n185 vdd.n176 5.04292
R5205 vdd.n138 vdd.n129 5.04292
R5206 vdd.n96 vdd.n87 5.04292
R5207 vdd.n49 vdd.n40 5.04292
R5208 vdd.n1170 vdd.n1161 5.04292
R5209 vdd.n1217 vdd.n1208 5.04292
R5210 vdd.n1080 vdd.n1071 5.04292
R5211 vdd.n1127 vdd.n1118 5.04292
R5212 vdd.n991 vdd.n982 5.04292
R5213 vdd.n1038 vdd.n1029 5.04292
R5214 vdd.n853 vdd.t86 4.98857
R5215 vdd.t55 vdd.n671 4.98857
R5216 vdd.n1553 vdd.t6 4.8752
R5217 vdd.t45 vdd.n888 4.8752
R5218 vdd.t159 vdd.t170 4.8752
R5219 vdd.n1948 vdd.t75 4.8752
R5220 vdd.n2615 vdd.t79 4.8752
R5221 vdd.t199 vdd.t149 4.8752
R5222 vdd.n636 vdd.t41 4.8752
R5223 vdd.t18 vdd.n304 4.8752
R5224 vdd.n2277 vdd.n2276 4.83952
R5225 vdd.n2017 vdd.n2016 4.83952
R5226 vdd.n2504 vdd.n2503 4.83952
R5227 vdd.n2797 vdd.n2796 4.83952
R5228 vdd.n591 vdd.n586 4.83952
R5229 vdd.n2438 vdd.n2377 4.83952
R5230 vdd.n2204 vdd.n789 4.83952
R5231 vdd.n1891 vdd.n1890 4.83952
R5232 vdd.n2172 vdd.t184 4.76184
R5233 vdd.n2655 vdd.t175 4.76184
R5234 vdd.n1701 vdd.n935 4.74817
R5235 vdd.n1696 vdd.n936 4.74817
R5236 vdd.n1598 vdd.n1595 4.74817
R5237 vdd.n1797 vdd.n1599 4.74817
R5238 vdd.n1799 vdd.n1598 4.74817
R5239 vdd.n1798 vdd.n1797 4.74817
R5240 vdd.n3020 vdd.n3019 4.74817
R5241 vdd.n3017 vdd.n3016 4.74817
R5242 vdd.n3017 vdd.n521 4.74817
R5243 vdd.n3019 vdd.n518 4.74817
R5244 vdd.n2902 vdd.n573 4.74817
R5245 vdd.n2898 vdd.n574 4.74817
R5246 vdd.n2901 vdd.n574 4.74817
R5247 vdd.n2905 vdd.n573 4.74817
R5248 vdd.n1697 vdd.n935 4.74817
R5249 vdd.n938 vdd.n936 4.74817
R5250 vdd.n297 vdd.n296 4.7074
R5251 vdd.n207 vdd.n206 4.7074
R5252 vdd.n1239 vdd.n1238 4.7074
R5253 vdd.n1149 vdd.n1148 4.7074
R5254 vdd.n1569 vdd.t15 4.64847
R5255 vdd.n3048 vdd.t2 4.64847
R5256 vdd.n1948 vdd.t167 4.30838
R5257 vdd.n2615 vdd.t154 4.30838
R5258 vdd.n276 vdd.n264 4.26717
R5259 vdd.n229 vdd.n217 4.26717
R5260 vdd.n186 vdd.n174 4.26717
R5261 vdd.n139 vdd.n127 4.26717
R5262 vdd.n97 vdd.n85 4.26717
R5263 vdd.n50 vdd.n38 4.26717
R5264 vdd.n1171 vdd.n1159 4.26717
R5265 vdd.n1218 vdd.n1206 4.26717
R5266 vdd.n1081 vdd.n1069 4.26717
R5267 vdd.n1128 vdd.n1116 4.26717
R5268 vdd.n992 vdd.n980 4.26717
R5269 vdd.n1039 vdd.n1027 4.26717
R5270 vdd.t160 vdd.n864 4.19501
R5271 vdd.n823 vdd.t174 4.19501
R5272 vdd.t188 vdd.n701 4.19501
R5273 vdd.n660 vdd.t183 4.19501
R5274 vdd.n297 vdd.n207 4.10845
R5275 vdd.n1239 vdd.n1149 4.10845
R5276 vdd.n253 vdd.t148 4.06363
R5277 vdd.n253 vdd.t207 4.06363
R5278 vdd.n251 vdd.t128 4.06363
R5279 vdd.n251 vdd.t118 4.06363
R5280 vdd.n249 vdd.t140 4.06363
R5281 vdd.n249 vdd.t116 4.06363
R5282 vdd.n163 vdd.t11 4.06363
R5283 vdd.n163 vdd.t143 4.06363
R5284 vdd.n161 vdd.t19 4.06363
R5285 vdd.n161 vdd.t206 4.06363
R5286 vdd.n159 vdd.t141 4.06363
R5287 vdd.n159 vdd.t129 4.06363
R5288 vdd.n74 vdd.t20 4.06363
R5289 vdd.n74 vdd.t125 4.06363
R5290 vdd.n72 vdd.t145 4.06363
R5291 vdd.n72 vdd.t135 4.06363
R5292 vdd.n70 vdd.t142 4.06363
R5293 vdd.n70 vdd.t25 4.06363
R5294 vdd.n1191 vdd.t17 4.06363
R5295 vdd.n1191 vdd.t22 4.06363
R5296 vdd.n1193 vdd.t138 4.06363
R5297 vdd.n1193 vdd.t202 4.06363
R5298 vdd.n1195 vdd.t127 4.06363
R5299 vdd.n1195 vdd.t13 4.06363
R5300 vdd.n1101 vdd.t1 4.06363
R5301 vdd.n1101 vdd.t120 4.06363
R5302 vdd.n1103 vdd.t107 4.06363
R5303 vdd.n1103 vdd.t7 4.06363
R5304 vdd.n1105 vdd.t205 4.06363
R5305 vdd.n1105 vdd.t147 4.06363
R5306 vdd.n1012 vdd.t134 4.06363
R5307 vdd.n1012 vdd.t204 4.06363
R5308 vdd.n1014 vdd.t123 4.06363
R5309 vdd.n1014 vdd.t119 4.06363
R5310 vdd.n1016 vdd.t131 4.06363
R5311 vdd.n1016 vdd.t130 4.06363
R5312 vdd.n26 vdd.t113 3.9605
R5313 vdd.n26 vdd.t114 3.9605
R5314 vdd.n23 vdd.t115 3.9605
R5315 vdd.n23 vdd.t5 3.9605
R5316 vdd.n21 vdd.t4 3.9605
R5317 vdd.n21 vdd.t105 3.9605
R5318 vdd.n20 vdd.t27 3.9605
R5319 vdd.n20 vdd.t110 3.9605
R5320 vdd.n15 vdd.t111 3.9605
R5321 vdd.n15 vdd.t132 3.9605
R5322 vdd.n16 vdd.t26 3.9605
R5323 vdd.n16 vdd.t109 3.9605
R5324 vdd.n18 vdd.t136 3.9605
R5325 vdd.n18 vdd.t133 3.9605
R5326 vdd.n25 vdd.t137 3.9605
R5327 vdd.n25 vdd.t104 3.9605
R5328 vdd.n2694 vdd.n2693 3.74684
R5329 vdd.n2134 vdd.n2133 3.74684
R5330 vdd.n7 vdd.t200 3.61217
R5331 vdd.n7 vdd.t166 3.61217
R5332 vdd.n8 vdd.t176 3.61217
R5333 vdd.n8 vdd.t196 3.61217
R5334 vdd.n10 vdd.t182 3.61217
R5335 vdd.n10 vdd.t155 3.61217
R5336 vdd.n12 vdd.t163 3.61217
R5337 vdd.n12 vdd.t180 3.61217
R5338 vdd.n5 vdd.t192 3.61217
R5339 vdd.n5 vdd.t173 3.61217
R5340 vdd.n3 vdd.t168 3.61217
R5341 vdd.n3 vdd.t194 3.61217
R5342 vdd.n1 vdd.t152 3.61217
R5343 vdd.n1 vdd.t185 3.61217
R5344 vdd.n0 vdd.t190 3.61217
R5345 vdd.n0 vdd.t171 3.61217
R5346 vdd.n2111 vdd.t160 3.51482
R5347 vdd.n2166 vdd.t174 3.51482
R5348 vdd.n2661 vdd.t188 3.51482
R5349 vdd.n2716 vdd.t183 3.51482
R5350 vdd.n280 vdd.n279 3.49141
R5351 vdd.n233 vdd.n232 3.49141
R5352 vdd.n190 vdd.n189 3.49141
R5353 vdd.n143 vdd.n142 3.49141
R5354 vdd.n101 vdd.n100 3.49141
R5355 vdd.n54 vdd.n53 3.49141
R5356 vdd.n1175 vdd.n1174 3.49141
R5357 vdd.n1222 vdd.n1221 3.49141
R5358 vdd.n1085 vdd.n1084 3.49141
R5359 vdd.n1132 vdd.n1131 3.49141
R5360 vdd.n996 vdd.n995 3.49141
R5361 vdd.n1043 vdd.n1042 3.49141
R5362 vdd.n2186 vdd.t167 3.40145
R5363 vdd.n2340 vdd.t191 3.40145
R5364 vdd.n2624 vdd.t179 3.40145
R5365 vdd.n2643 vdd.t154 3.40145
R5366 vdd.t184 vdd.n805 2.94799
R5367 vdd.n720 vdd.t175 2.94799
R5368 vdd.n1570 vdd.t21 2.83463
R5369 vdd.n1588 vdd.t62 2.83463
R5370 vdd.n2087 vdd.t45 2.83463
R5371 vdd.n2193 vdd.t75 2.83463
R5372 vdd.n2637 vdd.t79 2.83463
R5373 vdd.n2785 vdd.t41 2.83463
R5374 vdd.n3031 vdd.t37 2.83463
R5375 vdd.n467 vdd.t139 2.83463
R5376 vdd.n283 vdd.n262 2.71565
R5377 vdd.n236 vdd.n215 2.71565
R5378 vdd.n193 vdd.n172 2.71565
R5379 vdd.n146 vdd.n125 2.71565
R5380 vdd.n104 vdd.n83 2.71565
R5381 vdd.n57 vdd.n36 2.71565
R5382 vdd.n1178 vdd.n1157 2.71565
R5383 vdd.n1225 vdd.n1204 2.71565
R5384 vdd.n1088 vdd.n1067 2.71565
R5385 vdd.n1135 vdd.n1114 2.71565
R5386 vdd.n999 vdd.n978 2.71565
R5387 vdd.n1046 vdd.n1025 2.71565
R5388 vdd.t106 vdd.n1244 2.6079
R5389 vdd.n860 vdd.t178 2.6079
R5390 vdd.n1972 vdd.t197 2.6079
R5391 vdd.n2591 vdd.t187 2.6079
R5392 vdd.t156 vdd.n664 2.6079
R5393 vdd.n3225 vdd.t117 2.6079
R5394 vdd.n270 vdd.n269 2.4129
R5395 vdd.n223 vdd.n222 2.4129
R5396 vdd.n180 vdd.n179 2.4129
R5397 vdd.n133 vdd.n132 2.4129
R5398 vdd.n91 vdd.n90 2.4129
R5399 vdd.n44 vdd.n43 2.4129
R5400 vdd.n1165 vdd.n1164 2.4129
R5401 vdd.n1212 vdd.n1211 2.4129
R5402 vdd.n1075 vdd.n1074 2.4129
R5403 vdd.n1122 vdd.n1121 2.4129
R5404 vdd.n986 vdd.n985 2.4129
R5405 vdd.n1033 vdd.n1032 2.4129
R5406 vdd.n1527 vdd.t121 2.38117
R5407 vdd.n3216 vdd.t8 2.38117
R5408 vdd.n1796 vdd.n1598 2.27742
R5409 vdd.n1797 vdd.n1796 2.27742
R5410 vdd.n3018 vdd.n3017 2.27742
R5411 vdd.n3019 vdd.n3018 2.27742
R5412 vdd.n2889 vdd.n574 2.27742
R5413 vdd.n2889 vdd.n573 2.27742
R5414 vdd.n1819 vdd.n935 2.27742
R5415 vdd.n1819 vdd.n936 2.27742
R5416 vdd.n1972 vdd.t189 2.2678
R5417 vdd.n2591 vdd.t165 2.2678
R5418 vdd.n2160 vdd.t170 2.04107
R5419 vdd.n2667 vdd.t199 2.04107
R5420 vdd.n284 vdd.n260 1.93989
R5421 vdd.n237 vdd.n213 1.93989
R5422 vdd.n194 vdd.n170 1.93989
R5423 vdd.n147 vdd.n123 1.93989
R5424 vdd.n105 vdd.n81 1.93989
R5425 vdd.n58 vdd.n34 1.93989
R5426 vdd.n1179 vdd.n1155 1.93989
R5427 vdd.n1226 vdd.n1202 1.93989
R5428 vdd.n1089 vdd.n1065 1.93989
R5429 vdd.n1136 vdd.n1112 1.93989
R5430 vdd.n1000 vdd.n976 1.93989
R5431 vdd.n1047 vdd.n1023 1.93989
R5432 vdd.n2136 vdd.t157 1.70098
R5433 vdd.n2142 vdd.t164 1.70098
R5434 vdd.n2685 vdd.t169 1.70098
R5435 vdd.n2691 vdd.t158 1.70098
R5436 vdd.n2166 vdd.t151 1.36088
R5437 vdd.n2661 vdd.t195 1.36088
R5438 vdd.n1535 vdd.t12 1.24752
R5439 vdd.t10 vdd.n3223 1.24752
R5440 vdd.n295 vdd.n255 1.16414
R5441 vdd.n288 vdd.n287 1.16414
R5442 vdd.n248 vdd.n208 1.16414
R5443 vdd.n241 vdd.n240 1.16414
R5444 vdd.n205 vdd.n165 1.16414
R5445 vdd.n198 vdd.n197 1.16414
R5446 vdd.n158 vdd.n118 1.16414
R5447 vdd.n151 vdd.n150 1.16414
R5448 vdd.n116 vdd.n76 1.16414
R5449 vdd.n109 vdd.n108 1.16414
R5450 vdd.n69 vdd.n29 1.16414
R5451 vdd.n62 vdd.n61 1.16414
R5452 vdd.n1190 vdd.n1150 1.16414
R5453 vdd.n1183 vdd.n1182 1.16414
R5454 vdd.n1237 vdd.n1197 1.16414
R5455 vdd.n1230 vdd.n1229 1.16414
R5456 vdd.n1100 vdd.n1060 1.16414
R5457 vdd.n1093 vdd.n1092 1.16414
R5458 vdd.n1147 vdd.n1107 1.16414
R5459 vdd.n1140 vdd.n1139 1.16414
R5460 vdd.n1011 vdd.n971 1.16414
R5461 vdd.n1004 vdd.n1003 1.16414
R5462 vdd.n1058 vdd.n1018 1.16414
R5463 vdd.n1051 vdd.n1050 1.16414
R5464 vdd.n1561 vdd.t0 1.02079
R5465 vdd.t86 vdd.t157 1.02079
R5466 vdd.t158 vdd.t55 1.02079
R5467 vdd.t24 vdd.n456 1.02079
R5468 vdd.n1406 vdd.n1402 0.970197
R5469 vdd.n1817 vdd.n1816 0.970197
R5470 vdd.n3093 vdd.n3092 0.970197
R5471 vdd.n2897 vdd.n2895 0.970197
R5472 vdd.n1240 vdd.n28 0.956323
R5473 vdd vdd.n3230 0.94849
R5474 vdd.t193 vdd.n782 0.907421
R5475 vdd.n736 vdd.t181 0.907421
R5476 vdd.t161 vdd.n857 0.794056
R5477 vdd.n829 vdd.t159 0.794056
R5478 vdd.t149 vdd.n695 0.794056
R5479 vdd.n667 vdd.t186 0.794056
R5480 vdd.n1510 vdd.t33 0.567326
R5481 vdd.n3208 vdd.t29 0.567326
R5482 vdd.n1807 vdd.n1806 0.537085
R5483 vdd.n3027 vdd.n3026 0.537085
R5484 vdd.n3204 vdd.n3203 0.537085
R5485 vdd.n3086 vdd.n3085 0.537085
R5486 vdd.n2891 vdd.n476 0.537085
R5487 vdd.n1583 vdd.n937 0.537085
R5488 vdd.n1404 vdd.n1269 0.537085
R5489 vdd.n1506 vdd.n1505 0.537085
R5490 vdd.n4 vdd.n2 0.459552
R5491 vdd.n11 vdd.n9 0.459552
R5492 vdd.n293 vdd.n292 0.388379
R5493 vdd.n259 vdd.n257 0.388379
R5494 vdd.n246 vdd.n245 0.388379
R5495 vdd.n212 vdd.n210 0.388379
R5496 vdd.n203 vdd.n202 0.388379
R5497 vdd.n169 vdd.n167 0.388379
R5498 vdd.n156 vdd.n155 0.388379
R5499 vdd.n122 vdd.n120 0.388379
R5500 vdd.n114 vdd.n113 0.388379
R5501 vdd.n80 vdd.n78 0.388379
R5502 vdd.n67 vdd.n66 0.388379
R5503 vdd.n33 vdd.n31 0.388379
R5504 vdd.n1188 vdd.n1187 0.388379
R5505 vdd.n1154 vdd.n1152 0.388379
R5506 vdd.n1235 vdd.n1234 0.388379
R5507 vdd.n1201 vdd.n1199 0.388379
R5508 vdd.n1098 vdd.n1097 0.388379
R5509 vdd.n1064 vdd.n1062 0.388379
R5510 vdd.n1145 vdd.n1144 0.388379
R5511 vdd.n1111 vdd.n1109 0.388379
R5512 vdd.n1009 vdd.n1008 0.388379
R5513 vdd.n975 vdd.n973 0.388379
R5514 vdd.n1056 vdd.n1055 0.388379
R5515 vdd.n1022 vdd.n1020 0.388379
R5516 vdd.n19 vdd.n17 0.387128
R5517 vdd.n24 vdd.n22 0.387128
R5518 vdd.n6 vdd.n4 0.358259
R5519 vdd.n13 vdd.n11 0.358259
R5520 vdd.n252 vdd.n250 0.358259
R5521 vdd.n254 vdd.n252 0.358259
R5522 vdd.n296 vdd.n254 0.358259
R5523 vdd.n162 vdd.n160 0.358259
R5524 vdd.n164 vdd.n162 0.358259
R5525 vdd.n206 vdd.n164 0.358259
R5526 vdd.n73 vdd.n71 0.358259
R5527 vdd.n75 vdd.n73 0.358259
R5528 vdd.n117 vdd.n75 0.358259
R5529 vdd.n1238 vdd.n1196 0.358259
R5530 vdd.n1196 vdd.n1194 0.358259
R5531 vdd.n1194 vdd.n1192 0.358259
R5532 vdd.n1148 vdd.n1106 0.358259
R5533 vdd.n1106 vdd.n1104 0.358259
R5534 vdd.n1104 vdd.n1102 0.358259
R5535 vdd.n1059 vdd.n1017 0.358259
R5536 vdd.n1017 vdd.n1015 0.358259
R5537 vdd.n1015 vdd.n1013 0.358259
R5538 vdd.n14 vdd.n6 0.334552
R5539 vdd.n14 vdd.n13 0.334552
R5540 vdd.n27 vdd.n19 0.21707
R5541 vdd.n27 vdd.n24 0.21707
R5542 vdd.n294 vdd.n256 0.155672
R5543 vdd.n286 vdd.n256 0.155672
R5544 vdd.n286 vdd.n285 0.155672
R5545 vdd.n285 vdd.n261 0.155672
R5546 vdd.n278 vdd.n261 0.155672
R5547 vdd.n278 vdd.n277 0.155672
R5548 vdd.n277 vdd.n265 0.155672
R5549 vdd.n270 vdd.n265 0.155672
R5550 vdd.n247 vdd.n209 0.155672
R5551 vdd.n239 vdd.n209 0.155672
R5552 vdd.n239 vdd.n238 0.155672
R5553 vdd.n238 vdd.n214 0.155672
R5554 vdd.n231 vdd.n214 0.155672
R5555 vdd.n231 vdd.n230 0.155672
R5556 vdd.n230 vdd.n218 0.155672
R5557 vdd.n223 vdd.n218 0.155672
R5558 vdd.n204 vdd.n166 0.155672
R5559 vdd.n196 vdd.n166 0.155672
R5560 vdd.n196 vdd.n195 0.155672
R5561 vdd.n195 vdd.n171 0.155672
R5562 vdd.n188 vdd.n171 0.155672
R5563 vdd.n188 vdd.n187 0.155672
R5564 vdd.n187 vdd.n175 0.155672
R5565 vdd.n180 vdd.n175 0.155672
R5566 vdd.n157 vdd.n119 0.155672
R5567 vdd.n149 vdd.n119 0.155672
R5568 vdd.n149 vdd.n148 0.155672
R5569 vdd.n148 vdd.n124 0.155672
R5570 vdd.n141 vdd.n124 0.155672
R5571 vdd.n141 vdd.n140 0.155672
R5572 vdd.n140 vdd.n128 0.155672
R5573 vdd.n133 vdd.n128 0.155672
R5574 vdd.n115 vdd.n77 0.155672
R5575 vdd.n107 vdd.n77 0.155672
R5576 vdd.n107 vdd.n106 0.155672
R5577 vdd.n106 vdd.n82 0.155672
R5578 vdd.n99 vdd.n82 0.155672
R5579 vdd.n99 vdd.n98 0.155672
R5580 vdd.n98 vdd.n86 0.155672
R5581 vdd.n91 vdd.n86 0.155672
R5582 vdd.n68 vdd.n30 0.155672
R5583 vdd.n60 vdd.n30 0.155672
R5584 vdd.n60 vdd.n59 0.155672
R5585 vdd.n59 vdd.n35 0.155672
R5586 vdd.n52 vdd.n35 0.155672
R5587 vdd.n52 vdd.n51 0.155672
R5588 vdd.n51 vdd.n39 0.155672
R5589 vdd.n44 vdd.n39 0.155672
R5590 vdd.n1189 vdd.n1151 0.155672
R5591 vdd.n1181 vdd.n1151 0.155672
R5592 vdd.n1181 vdd.n1180 0.155672
R5593 vdd.n1180 vdd.n1156 0.155672
R5594 vdd.n1173 vdd.n1156 0.155672
R5595 vdd.n1173 vdd.n1172 0.155672
R5596 vdd.n1172 vdd.n1160 0.155672
R5597 vdd.n1165 vdd.n1160 0.155672
R5598 vdd.n1236 vdd.n1198 0.155672
R5599 vdd.n1228 vdd.n1198 0.155672
R5600 vdd.n1228 vdd.n1227 0.155672
R5601 vdd.n1227 vdd.n1203 0.155672
R5602 vdd.n1220 vdd.n1203 0.155672
R5603 vdd.n1220 vdd.n1219 0.155672
R5604 vdd.n1219 vdd.n1207 0.155672
R5605 vdd.n1212 vdd.n1207 0.155672
R5606 vdd.n1099 vdd.n1061 0.155672
R5607 vdd.n1091 vdd.n1061 0.155672
R5608 vdd.n1091 vdd.n1090 0.155672
R5609 vdd.n1090 vdd.n1066 0.155672
R5610 vdd.n1083 vdd.n1066 0.155672
R5611 vdd.n1083 vdd.n1082 0.155672
R5612 vdd.n1082 vdd.n1070 0.155672
R5613 vdd.n1075 vdd.n1070 0.155672
R5614 vdd.n1146 vdd.n1108 0.155672
R5615 vdd.n1138 vdd.n1108 0.155672
R5616 vdd.n1138 vdd.n1137 0.155672
R5617 vdd.n1137 vdd.n1113 0.155672
R5618 vdd.n1130 vdd.n1113 0.155672
R5619 vdd.n1130 vdd.n1129 0.155672
R5620 vdd.n1129 vdd.n1117 0.155672
R5621 vdd.n1122 vdd.n1117 0.155672
R5622 vdd.n1010 vdd.n972 0.155672
R5623 vdd.n1002 vdd.n972 0.155672
R5624 vdd.n1002 vdd.n1001 0.155672
R5625 vdd.n1001 vdd.n977 0.155672
R5626 vdd.n994 vdd.n977 0.155672
R5627 vdd.n994 vdd.n993 0.155672
R5628 vdd.n993 vdd.n981 0.155672
R5629 vdd.n986 vdd.n981 0.155672
R5630 vdd.n1057 vdd.n1019 0.155672
R5631 vdd.n1049 vdd.n1019 0.155672
R5632 vdd.n1049 vdd.n1048 0.155672
R5633 vdd.n1048 vdd.n1024 0.155672
R5634 vdd.n1041 vdd.n1024 0.155672
R5635 vdd.n1041 vdd.n1040 0.155672
R5636 vdd.n1040 vdd.n1028 0.155672
R5637 vdd.n1033 vdd.n1028 0.155672
R5638 vdd.n1795 vdd.n1600 0.152939
R5639 vdd.n1606 vdd.n1600 0.152939
R5640 vdd.n1607 vdd.n1606 0.152939
R5641 vdd.n1608 vdd.n1607 0.152939
R5642 vdd.n1609 vdd.n1608 0.152939
R5643 vdd.n1613 vdd.n1609 0.152939
R5644 vdd.n1614 vdd.n1613 0.152939
R5645 vdd.n1615 vdd.n1614 0.152939
R5646 vdd.n1616 vdd.n1615 0.152939
R5647 vdd.n1620 vdd.n1616 0.152939
R5648 vdd.n1621 vdd.n1620 0.152939
R5649 vdd.n1622 vdd.n1621 0.152939
R5650 vdd.n1770 vdd.n1622 0.152939
R5651 vdd.n1770 vdd.n1769 0.152939
R5652 vdd.n1769 vdd.n1768 0.152939
R5653 vdd.n1768 vdd.n1628 0.152939
R5654 vdd.n1633 vdd.n1628 0.152939
R5655 vdd.n1634 vdd.n1633 0.152939
R5656 vdd.n1635 vdd.n1634 0.152939
R5657 vdd.n1639 vdd.n1635 0.152939
R5658 vdd.n1640 vdd.n1639 0.152939
R5659 vdd.n1641 vdd.n1640 0.152939
R5660 vdd.n1642 vdd.n1641 0.152939
R5661 vdd.n1646 vdd.n1642 0.152939
R5662 vdd.n1647 vdd.n1646 0.152939
R5663 vdd.n1648 vdd.n1647 0.152939
R5664 vdd.n1649 vdd.n1648 0.152939
R5665 vdd.n1653 vdd.n1649 0.152939
R5666 vdd.n1654 vdd.n1653 0.152939
R5667 vdd.n1655 vdd.n1654 0.152939
R5668 vdd.n1656 vdd.n1655 0.152939
R5669 vdd.n1660 vdd.n1656 0.152939
R5670 vdd.n1661 vdd.n1660 0.152939
R5671 vdd.n1662 vdd.n1661 0.152939
R5672 vdd.n1731 vdd.n1662 0.152939
R5673 vdd.n1731 vdd.n1730 0.152939
R5674 vdd.n1730 vdd.n1729 0.152939
R5675 vdd.n1729 vdd.n1668 0.152939
R5676 vdd.n1673 vdd.n1668 0.152939
R5677 vdd.n1674 vdd.n1673 0.152939
R5678 vdd.n1675 vdd.n1674 0.152939
R5679 vdd.n1679 vdd.n1675 0.152939
R5680 vdd.n1680 vdd.n1679 0.152939
R5681 vdd.n1681 vdd.n1680 0.152939
R5682 vdd.n1682 vdd.n1681 0.152939
R5683 vdd.n1686 vdd.n1682 0.152939
R5684 vdd.n1687 vdd.n1686 0.152939
R5685 vdd.n1688 vdd.n1687 0.152939
R5686 vdd.n1689 vdd.n1688 0.152939
R5687 vdd.n1690 vdd.n1689 0.152939
R5688 vdd.n1690 vdd.n934 0.152939
R5689 vdd.n1806 vdd.n1594 0.152939
R5690 vdd.n1557 vdd.n1556 0.152939
R5691 vdd.n1558 vdd.n1557 0.152939
R5692 vdd.n1558 vdd.n959 0.152939
R5693 vdd.n1573 vdd.n959 0.152939
R5694 vdd.n1574 vdd.n1573 0.152939
R5695 vdd.n1575 vdd.n1574 0.152939
R5696 vdd.n1575 vdd.n947 0.152939
R5697 vdd.n1592 vdd.n947 0.152939
R5698 vdd.n1593 vdd.n1592 0.152939
R5699 vdd.n1807 vdd.n1593 0.152939
R5700 vdd.n524 vdd.n519 0.152939
R5701 vdd.n525 vdd.n524 0.152939
R5702 vdd.n526 vdd.n525 0.152939
R5703 vdd.n527 vdd.n526 0.152939
R5704 vdd.n528 vdd.n527 0.152939
R5705 vdd.n529 vdd.n528 0.152939
R5706 vdd.n530 vdd.n529 0.152939
R5707 vdd.n531 vdd.n530 0.152939
R5708 vdd.n532 vdd.n531 0.152939
R5709 vdd.n533 vdd.n532 0.152939
R5710 vdd.n534 vdd.n533 0.152939
R5711 vdd.n535 vdd.n534 0.152939
R5712 vdd.n2985 vdd.n535 0.152939
R5713 vdd.n2985 vdd.n2984 0.152939
R5714 vdd.n2984 vdd.n2983 0.152939
R5715 vdd.n2983 vdd.n537 0.152939
R5716 vdd.n538 vdd.n537 0.152939
R5717 vdd.n539 vdd.n538 0.152939
R5718 vdd.n540 vdd.n539 0.152939
R5719 vdd.n541 vdd.n540 0.152939
R5720 vdd.n542 vdd.n541 0.152939
R5721 vdd.n543 vdd.n542 0.152939
R5722 vdd.n544 vdd.n543 0.152939
R5723 vdd.n545 vdd.n544 0.152939
R5724 vdd.n546 vdd.n545 0.152939
R5725 vdd.n547 vdd.n546 0.152939
R5726 vdd.n548 vdd.n547 0.152939
R5727 vdd.n549 vdd.n548 0.152939
R5728 vdd.n550 vdd.n549 0.152939
R5729 vdd.n551 vdd.n550 0.152939
R5730 vdd.n552 vdd.n551 0.152939
R5731 vdd.n553 vdd.n552 0.152939
R5732 vdd.n554 vdd.n553 0.152939
R5733 vdd.n555 vdd.n554 0.152939
R5734 vdd.n2939 vdd.n555 0.152939
R5735 vdd.n2939 vdd.n2938 0.152939
R5736 vdd.n2938 vdd.n2937 0.152939
R5737 vdd.n2937 vdd.n559 0.152939
R5738 vdd.n560 vdd.n559 0.152939
R5739 vdd.n561 vdd.n560 0.152939
R5740 vdd.n562 vdd.n561 0.152939
R5741 vdd.n563 vdd.n562 0.152939
R5742 vdd.n564 vdd.n563 0.152939
R5743 vdd.n565 vdd.n564 0.152939
R5744 vdd.n566 vdd.n565 0.152939
R5745 vdd.n567 vdd.n566 0.152939
R5746 vdd.n568 vdd.n567 0.152939
R5747 vdd.n569 vdd.n568 0.152939
R5748 vdd.n570 vdd.n569 0.152939
R5749 vdd.n571 vdd.n570 0.152939
R5750 vdd.n572 vdd.n571 0.152939
R5751 vdd.n3026 vdd.n481 0.152939
R5752 vdd.n3028 vdd.n3027 0.152939
R5753 vdd.n3028 vdd.n470 0.152939
R5754 vdd.n3043 vdd.n470 0.152939
R5755 vdd.n3044 vdd.n3043 0.152939
R5756 vdd.n3045 vdd.n3044 0.152939
R5757 vdd.n3045 vdd.n459 0.152939
R5758 vdd.n3059 vdd.n459 0.152939
R5759 vdd.n3060 vdd.n3059 0.152939
R5760 vdd.n3061 vdd.n3060 0.152939
R5761 vdd.n3061 vdd.n298 0.152939
R5762 vdd.n3228 vdd.n299 0.152939
R5763 vdd.n310 vdd.n299 0.152939
R5764 vdd.n311 vdd.n310 0.152939
R5765 vdd.n312 vdd.n311 0.152939
R5766 vdd.n320 vdd.n312 0.152939
R5767 vdd.n321 vdd.n320 0.152939
R5768 vdd.n322 vdd.n321 0.152939
R5769 vdd.n323 vdd.n322 0.152939
R5770 vdd.n331 vdd.n323 0.152939
R5771 vdd.n3204 vdd.n331 0.152939
R5772 vdd.n3203 vdd.n332 0.152939
R5773 vdd.n335 vdd.n332 0.152939
R5774 vdd.n339 vdd.n335 0.152939
R5775 vdd.n340 vdd.n339 0.152939
R5776 vdd.n341 vdd.n340 0.152939
R5777 vdd.n342 vdd.n341 0.152939
R5778 vdd.n343 vdd.n342 0.152939
R5779 vdd.n347 vdd.n343 0.152939
R5780 vdd.n348 vdd.n347 0.152939
R5781 vdd.n349 vdd.n348 0.152939
R5782 vdd.n350 vdd.n349 0.152939
R5783 vdd.n354 vdd.n350 0.152939
R5784 vdd.n355 vdd.n354 0.152939
R5785 vdd.n356 vdd.n355 0.152939
R5786 vdd.n357 vdd.n356 0.152939
R5787 vdd.n361 vdd.n357 0.152939
R5788 vdd.n362 vdd.n361 0.152939
R5789 vdd.n363 vdd.n362 0.152939
R5790 vdd.n3169 vdd.n363 0.152939
R5791 vdd.n3169 vdd.n3168 0.152939
R5792 vdd.n3168 vdd.n3167 0.152939
R5793 vdd.n3167 vdd.n369 0.152939
R5794 vdd.n374 vdd.n369 0.152939
R5795 vdd.n375 vdd.n374 0.152939
R5796 vdd.n376 vdd.n375 0.152939
R5797 vdd.n380 vdd.n376 0.152939
R5798 vdd.n381 vdd.n380 0.152939
R5799 vdd.n382 vdd.n381 0.152939
R5800 vdd.n383 vdd.n382 0.152939
R5801 vdd.n387 vdd.n383 0.152939
R5802 vdd.n388 vdd.n387 0.152939
R5803 vdd.n389 vdd.n388 0.152939
R5804 vdd.n390 vdd.n389 0.152939
R5805 vdd.n394 vdd.n390 0.152939
R5806 vdd.n395 vdd.n394 0.152939
R5807 vdd.n396 vdd.n395 0.152939
R5808 vdd.n397 vdd.n396 0.152939
R5809 vdd.n401 vdd.n397 0.152939
R5810 vdd.n402 vdd.n401 0.152939
R5811 vdd.n403 vdd.n402 0.152939
R5812 vdd.n3130 vdd.n403 0.152939
R5813 vdd.n3130 vdd.n3129 0.152939
R5814 vdd.n3129 vdd.n3128 0.152939
R5815 vdd.n3128 vdd.n409 0.152939
R5816 vdd.n414 vdd.n409 0.152939
R5817 vdd.n415 vdd.n414 0.152939
R5818 vdd.n416 vdd.n415 0.152939
R5819 vdd.n420 vdd.n416 0.152939
R5820 vdd.n421 vdd.n420 0.152939
R5821 vdd.n422 vdd.n421 0.152939
R5822 vdd.n423 vdd.n422 0.152939
R5823 vdd.n427 vdd.n423 0.152939
R5824 vdd.n428 vdd.n427 0.152939
R5825 vdd.n429 vdd.n428 0.152939
R5826 vdd.n430 vdd.n429 0.152939
R5827 vdd.n434 vdd.n430 0.152939
R5828 vdd.n435 vdd.n434 0.152939
R5829 vdd.n436 vdd.n435 0.152939
R5830 vdd.n437 vdd.n436 0.152939
R5831 vdd.n441 vdd.n437 0.152939
R5832 vdd.n442 vdd.n441 0.152939
R5833 vdd.n443 vdd.n442 0.152939
R5834 vdd.n3086 vdd.n443 0.152939
R5835 vdd.n3034 vdd.n476 0.152939
R5836 vdd.n3035 vdd.n3034 0.152939
R5837 vdd.n3036 vdd.n3035 0.152939
R5838 vdd.n3036 vdd.n464 0.152939
R5839 vdd.n3051 vdd.n464 0.152939
R5840 vdd.n3052 vdd.n3051 0.152939
R5841 vdd.n3053 vdd.n3052 0.152939
R5842 vdd.n3053 vdd.n452 0.152939
R5843 vdd.n3067 vdd.n452 0.152939
R5844 vdd.n3068 vdd.n3067 0.152939
R5845 vdd.n3069 vdd.n3068 0.152939
R5846 vdd.n3069 vdd.n450 0.152939
R5847 vdd.n3073 vdd.n450 0.152939
R5848 vdd.n3074 vdd.n3073 0.152939
R5849 vdd.n3075 vdd.n3074 0.152939
R5850 vdd.n3075 vdd.n447 0.152939
R5851 vdd.n3079 vdd.n447 0.152939
R5852 vdd.n3080 vdd.n3079 0.152939
R5853 vdd.n3081 vdd.n3080 0.152939
R5854 vdd.n3081 vdd.n444 0.152939
R5855 vdd.n3085 vdd.n444 0.152939
R5856 vdd.n2891 vdd.n2890 0.152939
R5857 vdd.n1818 vdd.n937 0.152939
R5858 vdd.n1513 vdd.n1269 0.152939
R5859 vdd.n1514 vdd.n1513 0.152939
R5860 vdd.n1515 vdd.n1514 0.152939
R5861 vdd.n1515 vdd.n1257 0.152939
R5862 vdd.n1530 vdd.n1257 0.152939
R5863 vdd.n1531 vdd.n1530 0.152939
R5864 vdd.n1532 vdd.n1531 0.152939
R5865 vdd.n1532 vdd.n1247 0.152939
R5866 vdd.n1548 vdd.n1247 0.152939
R5867 vdd.n1549 vdd.n1548 0.152939
R5868 vdd.n1550 vdd.n1549 0.152939
R5869 vdd.n1550 vdd.n964 0.152939
R5870 vdd.n1564 vdd.n964 0.152939
R5871 vdd.n1565 vdd.n1564 0.152939
R5872 vdd.n1566 vdd.n1565 0.152939
R5873 vdd.n1566 vdd.n954 0.152939
R5874 vdd.n1581 vdd.n954 0.152939
R5875 vdd.n1582 vdd.n1581 0.152939
R5876 vdd.n1585 vdd.n1582 0.152939
R5877 vdd.n1585 vdd.n1584 0.152939
R5878 vdd.n1584 vdd.n1583 0.152939
R5879 vdd.n1505 vdd.n1274 0.152939
R5880 vdd.n1498 vdd.n1274 0.152939
R5881 vdd.n1498 vdd.n1497 0.152939
R5882 vdd.n1497 vdd.n1496 0.152939
R5883 vdd.n1496 vdd.n1311 0.152939
R5884 vdd.n1492 vdd.n1311 0.152939
R5885 vdd.n1492 vdd.n1491 0.152939
R5886 vdd.n1491 vdd.n1490 0.152939
R5887 vdd.n1490 vdd.n1317 0.152939
R5888 vdd.n1486 vdd.n1317 0.152939
R5889 vdd.n1486 vdd.n1485 0.152939
R5890 vdd.n1485 vdd.n1484 0.152939
R5891 vdd.n1484 vdd.n1323 0.152939
R5892 vdd.n1480 vdd.n1323 0.152939
R5893 vdd.n1480 vdd.n1479 0.152939
R5894 vdd.n1479 vdd.n1478 0.152939
R5895 vdd.n1478 vdd.n1329 0.152939
R5896 vdd.n1474 vdd.n1329 0.152939
R5897 vdd.n1474 vdd.n1473 0.152939
R5898 vdd.n1473 vdd.n1472 0.152939
R5899 vdd.n1472 vdd.n1337 0.152939
R5900 vdd.n1468 vdd.n1337 0.152939
R5901 vdd.n1468 vdd.n1467 0.152939
R5902 vdd.n1467 vdd.n1466 0.152939
R5903 vdd.n1466 vdd.n1343 0.152939
R5904 vdd.n1462 vdd.n1343 0.152939
R5905 vdd.n1462 vdd.n1461 0.152939
R5906 vdd.n1461 vdd.n1460 0.152939
R5907 vdd.n1460 vdd.n1349 0.152939
R5908 vdd.n1456 vdd.n1349 0.152939
R5909 vdd.n1456 vdd.n1455 0.152939
R5910 vdd.n1455 vdd.n1454 0.152939
R5911 vdd.n1454 vdd.n1355 0.152939
R5912 vdd.n1450 vdd.n1355 0.152939
R5913 vdd.n1450 vdd.n1449 0.152939
R5914 vdd.n1449 vdd.n1448 0.152939
R5915 vdd.n1448 vdd.n1361 0.152939
R5916 vdd.n1444 vdd.n1361 0.152939
R5917 vdd.n1444 vdd.n1443 0.152939
R5918 vdd.n1443 vdd.n1442 0.152939
R5919 vdd.n1442 vdd.n1367 0.152939
R5920 vdd.n1435 vdd.n1367 0.152939
R5921 vdd.n1435 vdd.n1434 0.152939
R5922 vdd.n1434 vdd.n1433 0.152939
R5923 vdd.n1433 vdd.n1372 0.152939
R5924 vdd.n1429 vdd.n1372 0.152939
R5925 vdd.n1429 vdd.n1428 0.152939
R5926 vdd.n1428 vdd.n1427 0.152939
R5927 vdd.n1427 vdd.n1378 0.152939
R5928 vdd.n1423 vdd.n1378 0.152939
R5929 vdd.n1423 vdd.n1422 0.152939
R5930 vdd.n1422 vdd.n1421 0.152939
R5931 vdd.n1421 vdd.n1384 0.152939
R5932 vdd.n1417 vdd.n1384 0.152939
R5933 vdd.n1417 vdd.n1416 0.152939
R5934 vdd.n1416 vdd.n1415 0.152939
R5935 vdd.n1415 vdd.n1390 0.152939
R5936 vdd.n1411 vdd.n1390 0.152939
R5937 vdd.n1411 vdd.n1410 0.152939
R5938 vdd.n1410 vdd.n1409 0.152939
R5939 vdd.n1409 vdd.n1396 0.152939
R5940 vdd.n1405 vdd.n1396 0.152939
R5941 vdd.n1405 vdd.n1404 0.152939
R5942 vdd.n1507 vdd.n1506 0.152939
R5943 vdd.n1507 vdd.n1263 0.152939
R5944 vdd.n1522 vdd.n1263 0.152939
R5945 vdd.n1523 vdd.n1522 0.152939
R5946 vdd.n1524 vdd.n1523 0.152939
R5947 vdd.n1524 vdd.n1252 0.152939
R5948 vdd.n1539 vdd.n1252 0.152939
R5949 vdd.n1540 vdd.n1539 0.152939
R5950 vdd.n1542 vdd.n1540 0.152939
R5951 vdd.n1542 vdd.n1541 0.152939
R5952 vdd.n2105 vdd.t198 0.113865
R5953 vdd.n2172 vdd.t150 0.113865
R5954 vdd.n2655 vdd.t153 0.113865
R5955 vdd.n2722 vdd.t177 0.113865
R5956 vdd.n1796 vdd.n1594 0.110256
R5957 vdd.n3018 vdd.n481 0.110256
R5958 vdd.n2890 vdd.n2889 0.110256
R5959 vdd.n1819 vdd.n1818 0.110256
R5960 vdd.n1556 vdd.n1241 0.0695946
R5961 vdd.n3229 vdd.n298 0.0695946
R5962 vdd.n3229 vdd.n3228 0.0695946
R5963 vdd.n1541 vdd.n1241 0.0695946
R5964 vdd.n1796 vdd.n1795 0.0431829
R5965 vdd.n1819 vdd.n934 0.0431829
R5966 vdd.n3018 vdd.n519 0.0431829
R5967 vdd.n2889 vdd.n572 0.0431829
R5968 vdd vdd.n28 0.00833333
R5969 a_n6972_8799.n98 a_n6972_8799.t55 485.149
R5970 a_n6972_8799.n105 a_n6972_8799.t59 485.149
R5971 a_n6972_8799.n113 a_n6972_8799.t84 485.149
R5972 a_n6972_8799.n74 a_n6972_8799.t83 485.149
R5973 a_n6972_8799.n81 a_n6972_8799.t90 485.149
R5974 a_n6972_8799.n89 a_n6972_8799.t85 485.149
R5975 a_n6972_8799.n26 a_n6972_8799.t69 485.135
R5976 a_n6972_8799.n102 a_n6972_8799.t46 464.166
R5977 a_n6972_8799.n96 a_n6972_8799.t71 464.166
R5978 a_n6972_8799.n101 a_n6972_8799.t70 464.166
R5979 a_n6972_8799.n100 a_n6972_8799.t48 464.166
R5980 a_n6972_8799.n97 a_n6972_8799.t47 464.166
R5981 a_n6972_8799.n99 a_n6972_8799.t81 464.166
R5982 a_n6972_8799.n31 a_n6972_8799.t76 485.135
R5983 a_n6972_8799.n109 a_n6972_8799.t50 464.166
R5984 a_n6972_8799.n103 a_n6972_8799.t79 464.166
R5985 a_n6972_8799.n108 a_n6972_8799.t77 464.166
R5986 a_n6972_8799.n107 a_n6972_8799.t52 464.166
R5987 a_n6972_8799.n104 a_n6972_8799.t51 464.166
R5988 a_n6972_8799.n106 a_n6972_8799.t88 464.166
R5989 a_n6972_8799.n36 a_n6972_8799.t56 485.135
R5990 a_n6972_8799.n117 a_n6972_8799.t91 464.166
R5991 a_n6972_8799.n111 a_n6972_8799.t75 464.166
R5992 a_n6972_8799.n116 a_n6972_8799.t86 464.166
R5993 a_n6972_8799.n115 a_n6972_8799.t67 464.166
R5994 a_n6972_8799.n112 a_n6972_8799.t78 464.166
R5995 a_n6972_8799.n114 a_n6972_8799.t53 464.166
R5996 a_n6972_8799.n75 a_n6972_8799.t62 464.166
R5997 a_n6972_8799.n76 a_n6972_8799.t63 464.166
R5998 a_n6972_8799.n77 a_n6972_8799.t73 464.166
R5999 a_n6972_8799.n78 a_n6972_8799.t58 464.166
R6000 a_n6972_8799.n73 a_n6972_8799.t57 464.166
R6001 a_n6972_8799.n79 a_n6972_8799.t72 464.166
R6002 a_n6972_8799.n82 a_n6972_8799.t66 464.166
R6003 a_n6972_8799.n83 a_n6972_8799.t65 464.166
R6004 a_n6972_8799.n84 a_n6972_8799.t82 464.166
R6005 a_n6972_8799.n85 a_n6972_8799.t60 464.166
R6006 a_n6972_8799.n80 a_n6972_8799.t61 464.166
R6007 a_n6972_8799.n86 a_n6972_8799.t80 464.166
R6008 a_n6972_8799.n90 a_n6972_8799.t54 464.166
R6009 a_n6972_8799.n91 a_n6972_8799.t45 464.166
R6010 a_n6972_8799.n92 a_n6972_8799.t68 464.166
R6011 a_n6972_8799.n93 a_n6972_8799.t87 464.166
R6012 a_n6972_8799.n88 a_n6972_8799.t74 464.166
R6013 a_n6972_8799.n94 a_n6972_8799.t89 464.166
R6014 a_n6972_8799.n20 a_n6972_8799.n30 72.3034
R6015 a_n6972_8799.n30 a_n6972_8799.n97 16.6962
R6016 a_n6972_8799.n29 a_n6972_8799.n20 77.6622
R6017 a_n6972_8799.n100 a_n6972_8799.n29 5.97853
R6018 a_n6972_8799.n28 a_n6972_8799.n19 77.6622
R6019 a_n6972_8799.n19 a_n6972_8799.n27 72.3034
R6020 a_n6972_8799.n102 a_n6972_8799.n26 20.9683
R6021 a_n6972_8799.n21 a_n6972_8799.n26 70.1674
R6022 a_n6972_8799.n17 a_n6972_8799.n35 72.3034
R6023 a_n6972_8799.n35 a_n6972_8799.n104 16.6962
R6024 a_n6972_8799.n34 a_n6972_8799.n17 77.6622
R6025 a_n6972_8799.n107 a_n6972_8799.n34 5.97853
R6026 a_n6972_8799.n33 a_n6972_8799.n16 77.6622
R6027 a_n6972_8799.n16 a_n6972_8799.n32 72.3034
R6028 a_n6972_8799.n109 a_n6972_8799.n31 20.9683
R6029 a_n6972_8799.n18 a_n6972_8799.n31 70.1674
R6030 a_n6972_8799.n14 a_n6972_8799.n40 72.3034
R6031 a_n6972_8799.n40 a_n6972_8799.n112 16.6962
R6032 a_n6972_8799.n39 a_n6972_8799.n14 77.6622
R6033 a_n6972_8799.n115 a_n6972_8799.n39 5.97853
R6034 a_n6972_8799.n38 a_n6972_8799.n13 77.6622
R6035 a_n6972_8799.n13 a_n6972_8799.n37 72.3034
R6036 a_n6972_8799.n117 a_n6972_8799.n36 20.9683
R6037 a_n6972_8799.n15 a_n6972_8799.n36 70.1674
R6038 a_n6972_8799.n11 a_n6972_8799.n45 70.1674
R6039 a_n6972_8799.n79 a_n6972_8799.n45 20.9683
R6040 a_n6972_8799.n44 a_n6972_8799.n11 72.3034
R6041 a_n6972_8799.n44 a_n6972_8799.n73 16.6962
R6042 a_n6972_8799.n10 a_n6972_8799.n43 77.6622
R6043 a_n6972_8799.n78 a_n6972_8799.n43 5.97853
R6044 a_n6972_8799.n42 a_n6972_8799.n10 77.6622
R6045 a_n6972_8799.n41 a_n6972_8799.n76 16.6962
R6046 a_n6972_8799.n41 a_n6972_8799.n12 72.3034
R6047 a_n6972_8799.n8 a_n6972_8799.n50 70.1674
R6048 a_n6972_8799.n86 a_n6972_8799.n50 20.9683
R6049 a_n6972_8799.n49 a_n6972_8799.n8 72.3034
R6050 a_n6972_8799.n49 a_n6972_8799.n80 16.6962
R6051 a_n6972_8799.n7 a_n6972_8799.n48 77.6622
R6052 a_n6972_8799.n85 a_n6972_8799.n48 5.97853
R6053 a_n6972_8799.n47 a_n6972_8799.n7 77.6622
R6054 a_n6972_8799.n46 a_n6972_8799.n83 16.6962
R6055 a_n6972_8799.n46 a_n6972_8799.n9 72.3034
R6056 a_n6972_8799.n5 a_n6972_8799.n55 70.1674
R6057 a_n6972_8799.n94 a_n6972_8799.n55 20.9683
R6058 a_n6972_8799.n54 a_n6972_8799.n5 72.3034
R6059 a_n6972_8799.n54 a_n6972_8799.n88 16.6962
R6060 a_n6972_8799.n4 a_n6972_8799.n53 77.6622
R6061 a_n6972_8799.n93 a_n6972_8799.n53 5.97853
R6062 a_n6972_8799.n52 a_n6972_8799.n4 77.6622
R6063 a_n6972_8799.n51 a_n6972_8799.n91 16.6962
R6064 a_n6972_8799.n51 a_n6972_8799.n6 72.3034
R6065 a_n6972_8799.n22 a_n6972_8799.n56 98.9633
R6066 a_n6972_8799.n126 a_n6972_8799.n25 98.9632
R6067 a_n6972_8799.n25 a_n6972_8799.n125 98.6055
R6068 a_n6972_8799.n25 a_n6972_8799.n124 98.6055
R6069 a_n6972_8799.n24 a_n6972_8799.n123 98.6055
R6070 a_n6972_8799.n24 a_n6972_8799.n122 98.6055
R6071 a_n6972_8799.n23 a_n6972_8799.n60 98.6055
R6072 a_n6972_8799.n23 a_n6972_8799.n59 98.6055
R6073 a_n6972_8799.n22 a_n6972_8799.n58 98.6055
R6074 a_n6972_8799.n22 a_n6972_8799.n57 98.6055
R6075 a_n6972_8799.n1 a_n6972_8799.n61 81.4626
R6076 a_n6972_8799.n3 a_n6972_8799.n67 81.4626
R6077 a_n6972_8799.n0 a_n6972_8799.n64 81.4626
R6078 a_n6972_8799.n2 a_n6972_8799.n70 80.9324
R6079 a_n6972_8799.n2 a_n6972_8799.n71 80.9324
R6080 a_n6972_8799.n1 a_n6972_8799.n72 80.9324
R6081 a_n6972_8799.n1 a_n6972_8799.n63 80.9324
R6082 a_n6972_8799.n1 a_n6972_8799.n62 80.9324
R6083 a_n6972_8799.n3 a_n6972_8799.n68 80.9324
R6084 a_n6972_8799.n0 a_n6972_8799.n69 80.9324
R6085 a_n6972_8799.n0 a_n6972_8799.n66 80.9324
R6086 a_n6972_8799.n0 a_n6972_8799.n65 80.9324
R6087 a_n6972_8799.n20 a_n6972_8799.n98 70.4033
R6088 a_n6972_8799.n17 a_n6972_8799.n105 70.4033
R6089 a_n6972_8799.n14 a_n6972_8799.n113 70.4033
R6090 a_n6972_8799.n74 a_n6972_8799.n12 70.4033
R6091 a_n6972_8799.n81 a_n6972_8799.n9 70.4033
R6092 a_n6972_8799.n89 a_n6972_8799.n6 70.4033
R6093 a_n6972_8799.n101 a_n6972_8799.n100 48.2005
R6094 a_n6972_8799.n108 a_n6972_8799.n107 48.2005
R6095 a_n6972_8799.n116 a_n6972_8799.n115 48.2005
R6096 a_n6972_8799.n78 a_n6972_8799.n77 48.2005
R6097 a_n6972_8799.t44 a_n6972_8799.n45 485.135
R6098 a_n6972_8799.n85 a_n6972_8799.n84 48.2005
R6099 a_n6972_8799.t49 a_n6972_8799.n50 485.135
R6100 a_n6972_8799.n93 a_n6972_8799.n92 48.2005
R6101 a_n6972_8799.t64 a_n6972_8799.n55 485.135
R6102 a_n6972_8799.n27 a_n6972_8799.n96 16.6962
R6103 a_n6972_8799.n99 a_n6972_8799.n30 27.6507
R6104 a_n6972_8799.n32 a_n6972_8799.n103 16.6962
R6105 a_n6972_8799.n106 a_n6972_8799.n35 27.6507
R6106 a_n6972_8799.n37 a_n6972_8799.n111 16.6962
R6107 a_n6972_8799.n114 a_n6972_8799.n40 27.6507
R6108 a_n6972_8799.n79 a_n6972_8799.n44 27.6507
R6109 a_n6972_8799.n86 a_n6972_8799.n49 27.6507
R6110 a_n6972_8799.n94 a_n6972_8799.n54 27.6507
R6111 a_n6972_8799.n28 a_n6972_8799.n96 41.7634
R6112 a_n6972_8799.n33 a_n6972_8799.n103 41.7634
R6113 a_n6972_8799.n38 a_n6972_8799.n111 41.7634
R6114 a_n6972_8799.n76 a_n6972_8799.n42 41.7634
R6115 a_n6972_8799.n83 a_n6972_8799.n47 41.7634
R6116 a_n6972_8799.n91 a_n6972_8799.n52 41.7634
R6117 a_n6972_8799.n2 a_n6972_8799.n0 34.3237
R6118 a_n6972_8799.n24 a_n6972_8799.n121 33.3407
R6119 a_n6972_8799.n99 a_n6972_8799.n98 20.9576
R6120 a_n6972_8799.n106 a_n6972_8799.n105 20.9576
R6121 a_n6972_8799.n114 a_n6972_8799.n113 20.9576
R6122 a_n6972_8799.n75 a_n6972_8799.n74 20.9576
R6123 a_n6972_8799.n82 a_n6972_8799.n81 20.9576
R6124 a_n6972_8799.n90 a_n6972_8799.n89 20.9576
R6125 a_n6972_8799.n121 a_n6972_8799.n23 19.402
R6126 a_n6972_8799.n28 a_n6972_8799.n101 5.97853
R6127 a_n6972_8799.n29 a_n6972_8799.n97 41.7634
R6128 a_n6972_8799.n33 a_n6972_8799.n108 5.97853
R6129 a_n6972_8799.n34 a_n6972_8799.n104 41.7634
R6130 a_n6972_8799.n38 a_n6972_8799.n116 5.97853
R6131 a_n6972_8799.n39 a_n6972_8799.n112 41.7634
R6132 a_n6972_8799.n77 a_n6972_8799.n42 5.97853
R6133 a_n6972_8799.n73 a_n6972_8799.n43 41.7634
R6134 a_n6972_8799.n84 a_n6972_8799.n47 5.97853
R6135 a_n6972_8799.n80 a_n6972_8799.n48 41.7634
R6136 a_n6972_8799.n92 a_n6972_8799.n52 5.97853
R6137 a_n6972_8799.n88 a_n6972_8799.n53 41.7634
R6138 a_n6972_8799.n120 a_n6972_8799.n1 12.3339
R6139 a_n6972_8799.n121 a_n6972_8799.n120 11.4887
R6140 a_n6972_8799.n102 a_n6972_8799.n27 27.6507
R6141 a_n6972_8799.n109 a_n6972_8799.n32 27.6507
R6142 a_n6972_8799.n117 a_n6972_8799.n37 27.6507
R6143 a_n6972_8799.n41 a_n6972_8799.n75 27.6507
R6144 a_n6972_8799.n46 a_n6972_8799.n82 27.6507
R6145 a_n6972_8799.n51 a_n6972_8799.n90 27.6507
R6146 a_n6972_8799.n110 a_n6972_8799.n21 9.05164
R6147 a_n6972_8799.n87 a_n6972_8799.n11 9.05164
R6148 a_n6972_8799.n119 a_n6972_8799.n95 7.14777
R6149 a_n6972_8799.n119 a_n6972_8799.n118 6.65114
R6150 a_n6972_8799.n110 a_n6972_8799.n18 4.94368
R6151 a_n6972_8799.n118 a_n6972_8799.n15 4.94368
R6152 a_n6972_8799.n87 a_n6972_8799.n8 4.94368
R6153 a_n6972_8799.n95 a_n6972_8799.n5 4.94368
R6154 a_n6972_8799.n118 a_n6972_8799.n110 4.10845
R6155 a_n6972_8799.n95 a_n6972_8799.n87 4.10845
R6156 a_n6972_8799.n125 a_n6972_8799.t29 3.61217
R6157 a_n6972_8799.n125 a_n6972_8799.t34 3.61217
R6158 a_n6972_8799.n124 a_n6972_8799.t23 3.61217
R6159 a_n6972_8799.n124 a_n6972_8799.t26 3.61217
R6160 a_n6972_8799.n123 a_n6972_8799.t28 3.61217
R6161 a_n6972_8799.n123 a_n6972_8799.t22 3.61217
R6162 a_n6972_8799.n122 a_n6972_8799.t25 3.61217
R6163 a_n6972_8799.n122 a_n6972_8799.t35 3.61217
R6164 a_n6972_8799.n60 a_n6972_8799.t31 3.61217
R6165 a_n6972_8799.n60 a_n6972_8799.t21 3.61217
R6166 a_n6972_8799.n59 a_n6972_8799.t19 3.61217
R6167 a_n6972_8799.n59 a_n6972_8799.t27 3.61217
R6168 a_n6972_8799.n58 a_n6972_8799.t32 3.61217
R6169 a_n6972_8799.n58 a_n6972_8799.t24 3.61217
R6170 a_n6972_8799.n57 a_n6972_8799.t18 3.61217
R6171 a_n6972_8799.n57 a_n6972_8799.t20 3.61217
R6172 a_n6972_8799.n56 a_n6972_8799.t33 3.61217
R6173 a_n6972_8799.n56 a_n6972_8799.t30 3.61217
R6174 a_n6972_8799.t17 a_n6972_8799.n126 3.61217
R6175 a_n6972_8799.n126 a_n6972_8799.t36 3.61217
R6176 a_n6972_8799.n120 a_n6972_8799.n119 3.4105
R6177 a_n6972_8799.n70 a_n6972_8799.t10 2.82907
R6178 a_n6972_8799.n70 a_n6972_8799.t9 2.82907
R6179 a_n6972_8799.n71 a_n6972_8799.t0 2.82907
R6180 a_n6972_8799.n71 a_n6972_8799.t13 2.82907
R6181 a_n6972_8799.n72 a_n6972_8799.t38 2.82907
R6182 a_n6972_8799.n72 a_n6972_8799.t5 2.82907
R6183 a_n6972_8799.n63 a_n6972_8799.t12 2.82907
R6184 a_n6972_8799.n63 a_n6972_8799.t1 2.82907
R6185 a_n6972_8799.n62 a_n6972_8799.t8 2.82907
R6186 a_n6972_8799.n62 a_n6972_8799.t37 2.82907
R6187 a_n6972_8799.n61 a_n6972_8799.t11 2.82907
R6188 a_n6972_8799.n61 a_n6972_8799.t43 2.82907
R6189 a_n6972_8799.n67 a_n6972_8799.t4 2.82907
R6190 a_n6972_8799.n67 a_n6972_8799.t14 2.82907
R6191 a_n6972_8799.n68 a_n6972_8799.t15 2.82907
R6192 a_n6972_8799.n68 a_n6972_8799.t6 2.82907
R6193 a_n6972_8799.n69 a_n6972_8799.t16 2.82907
R6194 a_n6972_8799.n69 a_n6972_8799.t2 2.82907
R6195 a_n6972_8799.n66 a_n6972_8799.t7 2.82907
R6196 a_n6972_8799.n66 a_n6972_8799.t39 2.82907
R6197 a_n6972_8799.n65 a_n6972_8799.t41 2.82907
R6198 a_n6972_8799.n65 a_n6972_8799.t42 2.82907
R6199 a_n6972_8799.n64 a_n6972_8799.t3 2.82907
R6200 a_n6972_8799.n64 a_n6972_8799.t40 2.82907
R6201 a_n6972_8799.n1 a_n6972_8799.n2 2.12119
R6202 a_n6972_8799.n0 a_n6972_8799.n3 1.59102
R6203 a_n6972_8799.n20 a_n6972_8799.n19 1.13686
R6204 a_n6972_8799.n17 a_n6972_8799.n16 1.13686
R6205 a_n6972_8799.n14 a_n6972_8799.n13 1.13686
R6206 a_n6972_8799.n11 a_n6972_8799.n10 1.13686
R6207 a_n6972_8799.n8 a_n6972_8799.n7 1.13686
R6208 a_n6972_8799.n5 a_n6972_8799.n4 1.13686
R6209 a_n6972_8799.n25 a_n6972_8799.n24 1.07378
R6210 a_n6972_8799.n23 a_n6972_8799.n22 1.07378
R6211 a_n6972_8799.n4 a_n6972_8799.n6 0.568682
R6212 a_n6972_8799.n7 a_n6972_8799.n9 0.568682
R6213 a_n6972_8799.n10 a_n6972_8799.n12 0.568682
R6214 a_n6972_8799.n13 a_n6972_8799.n15 0.568682
R6215 a_n6972_8799.n16 a_n6972_8799.n18 0.568682
R6216 a_n6972_8799.n19 a_n6972_8799.n21 0.568682
R6217 CSoutput.n19 CSoutput.t134 184.661
R6218 CSoutput.n78 CSoutput.n77 165.8
R6219 CSoutput.n76 CSoutput.n0 165.8
R6220 CSoutput.n75 CSoutput.n74 165.8
R6221 CSoutput.n73 CSoutput.n72 165.8
R6222 CSoutput.n71 CSoutput.n2 165.8
R6223 CSoutput.n69 CSoutput.n68 165.8
R6224 CSoutput.n67 CSoutput.n3 165.8
R6225 CSoutput.n66 CSoutput.n65 165.8
R6226 CSoutput.n63 CSoutput.n4 165.8
R6227 CSoutput.n61 CSoutput.n60 165.8
R6228 CSoutput.n59 CSoutput.n5 165.8
R6229 CSoutput.n58 CSoutput.n57 165.8
R6230 CSoutput.n55 CSoutput.n6 165.8
R6231 CSoutput.n54 CSoutput.n53 165.8
R6232 CSoutput.n52 CSoutput.n51 165.8
R6233 CSoutput.n50 CSoutput.n8 165.8
R6234 CSoutput.n48 CSoutput.n47 165.8
R6235 CSoutput.n46 CSoutput.n9 165.8
R6236 CSoutput.n45 CSoutput.n44 165.8
R6237 CSoutput.n42 CSoutput.n10 165.8
R6238 CSoutput.n41 CSoutput.n40 165.8
R6239 CSoutput.n39 CSoutput.n38 165.8
R6240 CSoutput.n37 CSoutput.n12 165.8
R6241 CSoutput.n35 CSoutput.n34 165.8
R6242 CSoutput.n33 CSoutput.n13 165.8
R6243 CSoutput.n32 CSoutput.n31 165.8
R6244 CSoutput.n29 CSoutput.n14 165.8
R6245 CSoutput.n28 CSoutput.n27 165.8
R6246 CSoutput.n26 CSoutput.n25 165.8
R6247 CSoutput.n24 CSoutput.n16 165.8
R6248 CSoutput.n22 CSoutput.n21 165.8
R6249 CSoutput.n20 CSoutput.n17 165.8
R6250 CSoutput.n77 CSoutput.t136 162.194
R6251 CSoutput.n18 CSoutput.t145 120.501
R6252 CSoutput.n23 CSoutput.t147 120.501
R6253 CSoutput.n15 CSoutput.t140 120.501
R6254 CSoutput.n30 CSoutput.t131 120.501
R6255 CSoutput.n36 CSoutput.t149 120.501
R6256 CSoutput.n11 CSoutput.t143 120.501
R6257 CSoutput.n43 CSoutput.t138 120.501
R6258 CSoutput.n49 CSoutput.t129 120.501
R6259 CSoutput.n7 CSoutput.t130 120.501
R6260 CSoutput.n56 CSoutput.t141 120.501
R6261 CSoutput.n62 CSoutput.t137 120.501
R6262 CSoutput.n64 CSoutput.t133 120.501
R6263 CSoutput.n70 CSoutput.t144 120.501
R6264 CSoutput.n1 CSoutput.t146 120.501
R6265 CSoutput.n270 CSoutput.n268 103.469
R6266 CSoutput.n262 CSoutput.n260 103.469
R6267 CSoutput.n255 CSoutput.n253 103.469
R6268 CSoutput.n96 CSoutput.n94 103.469
R6269 CSoutput.n88 CSoutput.n86 103.469
R6270 CSoutput.n81 CSoutput.n79 103.469
R6271 CSoutput.n272 CSoutput.n271 103.111
R6272 CSoutput.n270 CSoutput.n269 103.111
R6273 CSoutput.n266 CSoutput.n265 103.111
R6274 CSoutput.n264 CSoutput.n263 103.111
R6275 CSoutput.n262 CSoutput.n261 103.111
R6276 CSoutput.n259 CSoutput.n258 103.111
R6277 CSoutput.n257 CSoutput.n256 103.111
R6278 CSoutput.n255 CSoutput.n254 103.111
R6279 CSoutput.n96 CSoutput.n95 103.111
R6280 CSoutput.n98 CSoutput.n97 103.111
R6281 CSoutput.n100 CSoutput.n99 103.111
R6282 CSoutput.n88 CSoutput.n87 103.111
R6283 CSoutput.n90 CSoutput.n89 103.111
R6284 CSoutput.n92 CSoutput.n91 103.111
R6285 CSoutput.n81 CSoutput.n80 103.111
R6286 CSoutput.n83 CSoutput.n82 103.111
R6287 CSoutput.n85 CSoutput.n84 103.111
R6288 CSoutput.n274 CSoutput.n273 103.111
R6289 CSoutput.n298 CSoutput.n296 81.5057
R6290 CSoutput.n279 CSoutput.n277 81.5057
R6291 CSoutput.n338 CSoutput.n336 81.5057
R6292 CSoutput.n319 CSoutput.n317 81.5057
R6293 CSoutput.n314 CSoutput.n313 80.9324
R6294 CSoutput.n312 CSoutput.n311 80.9324
R6295 CSoutput.n310 CSoutput.n309 80.9324
R6296 CSoutput.n308 CSoutput.n307 80.9324
R6297 CSoutput.n306 CSoutput.n305 80.9324
R6298 CSoutput.n304 CSoutput.n303 80.9324
R6299 CSoutput.n302 CSoutput.n301 80.9324
R6300 CSoutput.n300 CSoutput.n299 80.9324
R6301 CSoutput.n298 CSoutput.n297 80.9324
R6302 CSoutput.n295 CSoutput.n294 80.9324
R6303 CSoutput.n293 CSoutput.n292 80.9324
R6304 CSoutput.n291 CSoutput.n290 80.9324
R6305 CSoutput.n289 CSoutput.n288 80.9324
R6306 CSoutput.n287 CSoutput.n286 80.9324
R6307 CSoutput.n285 CSoutput.n284 80.9324
R6308 CSoutput.n283 CSoutput.n282 80.9324
R6309 CSoutput.n281 CSoutput.n280 80.9324
R6310 CSoutput.n279 CSoutput.n278 80.9324
R6311 CSoutput.n338 CSoutput.n337 80.9324
R6312 CSoutput.n340 CSoutput.n339 80.9324
R6313 CSoutput.n342 CSoutput.n341 80.9324
R6314 CSoutput.n344 CSoutput.n343 80.9324
R6315 CSoutput.n346 CSoutput.n345 80.9324
R6316 CSoutput.n348 CSoutput.n347 80.9324
R6317 CSoutput.n350 CSoutput.n349 80.9324
R6318 CSoutput.n352 CSoutput.n351 80.9324
R6319 CSoutput.n354 CSoutput.n353 80.9324
R6320 CSoutput.n319 CSoutput.n318 80.9324
R6321 CSoutput.n321 CSoutput.n320 80.9324
R6322 CSoutput.n323 CSoutput.n322 80.9324
R6323 CSoutput.n325 CSoutput.n324 80.9324
R6324 CSoutput.n327 CSoutput.n326 80.9324
R6325 CSoutput.n329 CSoutput.n328 80.9324
R6326 CSoutput.n331 CSoutput.n330 80.9324
R6327 CSoutput.n333 CSoutput.n332 80.9324
R6328 CSoutput.n335 CSoutput.n334 80.9324
R6329 CSoutput.n25 CSoutput.n24 48.1486
R6330 CSoutput.n69 CSoutput.n3 48.1486
R6331 CSoutput.n38 CSoutput.n37 48.1486
R6332 CSoutput.n42 CSoutput.n41 48.1486
R6333 CSoutput.n51 CSoutput.n50 48.1486
R6334 CSoutput.n55 CSoutput.n54 48.1486
R6335 CSoutput.n22 CSoutput.n17 46.462
R6336 CSoutput.n72 CSoutput.n71 46.462
R6337 CSoutput.n20 CSoutput.n19 44.9055
R6338 CSoutput.n29 CSoutput.n28 43.7635
R6339 CSoutput.n65 CSoutput.n63 43.7635
R6340 CSoutput.n35 CSoutput.n13 41.7396
R6341 CSoutput.n57 CSoutput.n5 41.7396
R6342 CSoutput.n44 CSoutput.n9 37.0171
R6343 CSoutput.n48 CSoutput.n9 37.0171
R6344 CSoutput.n76 CSoutput.n75 34.9932
R6345 CSoutput.n31 CSoutput.n13 32.2947
R6346 CSoutput.n61 CSoutput.n5 32.2947
R6347 CSoutput.n30 CSoutput.n29 29.6014
R6348 CSoutput.n63 CSoutput.n62 29.6014
R6349 CSoutput.n19 CSoutput.n18 28.4085
R6350 CSoutput.n18 CSoutput.n17 25.1176
R6351 CSoutput.n72 CSoutput.n1 25.1176
R6352 CSoutput.n43 CSoutput.n42 22.0922
R6353 CSoutput.n50 CSoutput.n49 22.0922
R6354 CSoutput.n77 CSoutput.n76 21.8586
R6355 CSoutput.n37 CSoutput.n36 18.9681
R6356 CSoutput.n56 CSoutput.n55 18.9681
R6357 CSoutput.n25 CSoutput.n15 17.6292
R6358 CSoutput.n64 CSoutput.n3 17.6292
R6359 CSoutput.n24 CSoutput.n23 15.844
R6360 CSoutput.n70 CSoutput.n69 15.844
R6361 CSoutput.n38 CSoutput.n11 14.5051
R6362 CSoutput.n54 CSoutput.n7 14.5051
R6363 CSoutput.n357 CSoutput.n78 11.6139
R6364 CSoutput.n41 CSoutput.n11 11.3811
R6365 CSoutput.n51 CSoutput.n7 11.3811
R6366 CSoutput.n23 CSoutput.n22 10.0422
R6367 CSoutput.n71 CSoutput.n70 10.0422
R6368 CSoutput.n267 CSoutput.n259 9.25285
R6369 CSoutput.n93 CSoutput.n85 9.25285
R6370 CSoutput.n316 CSoutput.n276 9.05363
R6371 CSoutput.n315 CSoutput.n295 8.97993
R6372 CSoutput.n355 CSoutput.n335 8.97993
R6373 CSoutput.n28 CSoutput.n15 8.25698
R6374 CSoutput.n65 CSoutput.n64 8.25698
R6375 CSoutput.n316 CSoutput.n315 7.89345
R6376 CSoutput.n356 CSoutput.n355 7.89345
R6377 CSoutput.n276 CSoutput.n275 7.12641
R6378 CSoutput.n102 CSoutput.n101 7.12641
R6379 CSoutput.n36 CSoutput.n35 6.91809
R6380 CSoutput.n57 CSoutput.n56 6.91809
R6381 CSoutput.n357 CSoutput.n102 5.46119
R6382 CSoutput.n315 CSoutput.n314 5.25266
R6383 CSoutput.n355 CSoutput.n354 5.25266
R6384 CSoutput.n275 CSoutput.n274 5.1449
R6385 CSoutput.n267 CSoutput.n266 5.1449
R6386 CSoutput.n101 CSoutput.n100 5.1449
R6387 CSoutput.n93 CSoutput.n92 5.1449
R6388 CSoutput.n193 CSoutput.n146 4.5005
R6389 CSoutput.n162 CSoutput.n146 4.5005
R6390 CSoutput.n157 CSoutput.n141 4.5005
R6391 CSoutput.n157 CSoutput.n143 4.5005
R6392 CSoutput.n157 CSoutput.n140 4.5005
R6393 CSoutput.n157 CSoutput.n144 4.5005
R6394 CSoutput.n157 CSoutput.n139 4.5005
R6395 CSoutput.n157 CSoutput.t148 4.5005
R6396 CSoutput.n157 CSoutput.n138 4.5005
R6397 CSoutput.n157 CSoutput.n145 4.5005
R6398 CSoutput.n157 CSoutput.n146 4.5005
R6399 CSoutput.n155 CSoutput.n141 4.5005
R6400 CSoutput.n155 CSoutput.n143 4.5005
R6401 CSoutput.n155 CSoutput.n140 4.5005
R6402 CSoutput.n155 CSoutput.n144 4.5005
R6403 CSoutput.n155 CSoutput.n139 4.5005
R6404 CSoutput.n155 CSoutput.t148 4.5005
R6405 CSoutput.n155 CSoutput.n138 4.5005
R6406 CSoutput.n155 CSoutput.n145 4.5005
R6407 CSoutput.n155 CSoutput.n146 4.5005
R6408 CSoutput.n154 CSoutput.n141 4.5005
R6409 CSoutput.n154 CSoutput.n143 4.5005
R6410 CSoutput.n154 CSoutput.n140 4.5005
R6411 CSoutput.n154 CSoutput.n144 4.5005
R6412 CSoutput.n154 CSoutput.n139 4.5005
R6413 CSoutput.n154 CSoutput.t148 4.5005
R6414 CSoutput.n154 CSoutput.n138 4.5005
R6415 CSoutput.n154 CSoutput.n145 4.5005
R6416 CSoutput.n154 CSoutput.n146 4.5005
R6417 CSoutput.n239 CSoutput.n141 4.5005
R6418 CSoutput.n239 CSoutput.n143 4.5005
R6419 CSoutput.n239 CSoutput.n140 4.5005
R6420 CSoutput.n239 CSoutput.n144 4.5005
R6421 CSoutput.n239 CSoutput.n139 4.5005
R6422 CSoutput.n239 CSoutput.t148 4.5005
R6423 CSoutput.n239 CSoutput.n138 4.5005
R6424 CSoutput.n239 CSoutput.n145 4.5005
R6425 CSoutput.n239 CSoutput.n146 4.5005
R6426 CSoutput.n237 CSoutput.n141 4.5005
R6427 CSoutput.n237 CSoutput.n143 4.5005
R6428 CSoutput.n237 CSoutput.n140 4.5005
R6429 CSoutput.n237 CSoutput.n144 4.5005
R6430 CSoutput.n237 CSoutput.n139 4.5005
R6431 CSoutput.n237 CSoutput.t148 4.5005
R6432 CSoutput.n237 CSoutput.n138 4.5005
R6433 CSoutput.n237 CSoutput.n145 4.5005
R6434 CSoutput.n235 CSoutput.n141 4.5005
R6435 CSoutput.n235 CSoutput.n143 4.5005
R6436 CSoutput.n235 CSoutput.n140 4.5005
R6437 CSoutput.n235 CSoutput.n144 4.5005
R6438 CSoutput.n235 CSoutput.n139 4.5005
R6439 CSoutput.n235 CSoutput.t148 4.5005
R6440 CSoutput.n235 CSoutput.n138 4.5005
R6441 CSoutput.n235 CSoutput.n145 4.5005
R6442 CSoutput.n165 CSoutput.n141 4.5005
R6443 CSoutput.n165 CSoutput.n143 4.5005
R6444 CSoutput.n165 CSoutput.n140 4.5005
R6445 CSoutput.n165 CSoutput.n144 4.5005
R6446 CSoutput.n165 CSoutput.n139 4.5005
R6447 CSoutput.n165 CSoutput.t148 4.5005
R6448 CSoutput.n165 CSoutput.n138 4.5005
R6449 CSoutput.n165 CSoutput.n145 4.5005
R6450 CSoutput.n165 CSoutput.n146 4.5005
R6451 CSoutput.n164 CSoutput.n141 4.5005
R6452 CSoutput.n164 CSoutput.n143 4.5005
R6453 CSoutput.n164 CSoutput.n140 4.5005
R6454 CSoutput.n164 CSoutput.n144 4.5005
R6455 CSoutput.n164 CSoutput.n139 4.5005
R6456 CSoutput.n164 CSoutput.t148 4.5005
R6457 CSoutput.n164 CSoutput.n138 4.5005
R6458 CSoutput.n164 CSoutput.n145 4.5005
R6459 CSoutput.n164 CSoutput.n146 4.5005
R6460 CSoutput.n168 CSoutput.n141 4.5005
R6461 CSoutput.n168 CSoutput.n143 4.5005
R6462 CSoutput.n168 CSoutput.n140 4.5005
R6463 CSoutput.n168 CSoutput.n144 4.5005
R6464 CSoutput.n168 CSoutput.n139 4.5005
R6465 CSoutput.n168 CSoutput.t148 4.5005
R6466 CSoutput.n168 CSoutput.n138 4.5005
R6467 CSoutput.n168 CSoutput.n145 4.5005
R6468 CSoutput.n168 CSoutput.n146 4.5005
R6469 CSoutput.n167 CSoutput.n141 4.5005
R6470 CSoutput.n167 CSoutput.n143 4.5005
R6471 CSoutput.n167 CSoutput.n140 4.5005
R6472 CSoutput.n167 CSoutput.n144 4.5005
R6473 CSoutput.n167 CSoutput.n139 4.5005
R6474 CSoutput.n167 CSoutput.t148 4.5005
R6475 CSoutput.n167 CSoutput.n138 4.5005
R6476 CSoutput.n167 CSoutput.n145 4.5005
R6477 CSoutput.n167 CSoutput.n146 4.5005
R6478 CSoutput.n150 CSoutput.n141 4.5005
R6479 CSoutput.n150 CSoutput.n143 4.5005
R6480 CSoutput.n150 CSoutput.n140 4.5005
R6481 CSoutput.n150 CSoutput.n144 4.5005
R6482 CSoutput.n150 CSoutput.n139 4.5005
R6483 CSoutput.n150 CSoutput.t148 4.5005
R6484 CSoutput.n150 CSoutput.n138 4.5005
R6485 CSoutput.n150 CSoutput.n145 4.5005
R6486 CSoutput.n150 CSoutput.n146 4.5005
R6487 CSoutput.n242 CSoutput.n141 4.5005
R6488 CSoutput.n242 CSoutput.n143 4.5005
R6489 CSoutput.n242 CSoutput.n140 4.5005
R6490 CSoutput.n242 CSoutput.n144 4.5005
R6491 CSoutput.n242 CSoutput.n139 4.5005
R6492 CSoutput.n242 CSoutput.t148 4.5005
R6493 CSoutput.n242 CSoutput.n138 4.5005
R6494 CSoutput.n242 CSoutput.n145 4.5005
R6495 CSoutput.n242 CSoutput.n146 4.5005
R6496 CSoutput.n229 CSoutput.n200 4.5005
R6497 CSoutput.n229 CSoutput.n206 4.5005
R6498 CSoutput.n187 CSoutput.n176 4.5005
R6499 CSoutput.n187 CSoutput.n178 4.5005
R6500 CSoutput.n187 CSoutput.n175 4.5005
R6501 CSoutput.n187 CSoutput.n179 4.5005
R6502 CSoutput.n187 CSoutput.n174 4.5005
R6503 CSoutput.n187 CSoutput.t142 4.5005
R6504 CSoutput.n187 CSoutput.n173 4.5005
R6505 CSoutput.n187 CSoutput.n180 4.5005
R6506 CSoutput.n229 CSoutput.n187 4.5005
R6507 CSoutput.n208 CSoutput.n176 4.5005
R6508 CSoutput.n208 CSoutput.n178 4.5005
R6509 CSoutput.n208 CSoutput.n175 4.5005
R6510 CSoutput.n208 CSoutput.n179 4.5005
R6511 CSoutput.n208 CSoutput.n174 4.5005
R6512 CSoutput.n208 CSoutput.t142 4.5005
R6513 CSoutput.n208 CSoutput.n173 4.5005
R6514 CSoutput.n208 CSoutput.n180 4.5005
R6515 CSoutput.n229 CSoutput.n208 4.5005
R6516 CSoutput.n186 CSoutput.n176 4.5005
R6517 CSoutput.n186 CSoutput.n178 4.5005
R6518 CSoutput.n186 CSoutput.n175 4.5005
R6519 CSoutput.n186 CSoutput.n179 4.5005
R6520 CSoutput.n186 CSoutput.n174 4.5005
R6521 CSoutput.n186 CSoutput.t142 4.5005
R6522 CSoutput.n186 CSoutput.n173 4.5005
R6523 CSoutput.n186 CSoutput.n180 4.5005
R6524 CSoutput.n229 CSoutput.n186 4.5005
R6525 CSoutput.n210 CSoutput.n176 4.5005
R6526 CSoutput.n210 CSoutput.n178 4.5005
R6527 CSoutput.n210 CSoutput.n175 4.5005
R6528 CSoutput.n210 CSoutput.n179 4.5005
R6529 CSoutput.n210 CSoutput.n174 4.5005
R6530 CSoutput.n210 CSoutput.t142 4.5005
R6531 CSoutput.n210 CSoutput.n173 4.5005
R6532 CSoutput.n210 CSoutput.n180 4.5005
R6533 CSoutput.n229 CSoutput.n210 4.5005
R6534 CSoutput.n176 CSoutput.n171 4.5005
R6535 CSoutput.n178 CSoutput.n171 4.5005
R6536 CSoutput.n175 CSoutput.n171 4.5005
R6537 CSoutput.n179 CSoutput.n171 4.5005
R6538 CSoutput.n174 CSoutput.n171 4.5005
R6539 CSoutput.t142 CSoutput.n171 4.5005
R6540 CSoutput.n173 CSoutput.n171 4.5005
R6541 CSoutput.n180 CSoutput.n171 4.5005
R6542 CSoutput.n232 CSoutput.n176 4.5005
R6543 CSoutput.n232 CSoutput.n178 4.5005
R6544 CSoutput.n232 CSoutput.n175 4.5005
R6545 CSoutput.n232 CSoutput.n179 4.5005
R6546 CSoutput.n232 CSoutput.n174 4.5005
R6547 CSoutput.n232 CSoutput.t142 4.5005
R6548 CSoutput.n232 CSoutput.n173 4.5005
R6549 CSoutput.n232 CSoutput.n180 4.5005
R6550 CSoutput.n230 CSoutput.n176 4.5005
R6551 CSoutput.n230 CSoutput.n178 4.5005
R6552 CSoutput.n230 CSoutput.n175 4.5005
R6553 CSoutput.n230 CSoutput.n179 4.5005
R6554 CSoutput.n230 CSoutput.n174 4.5005
R6555 CSoutput.n230 CSoutput.t142 4.5005
R6556 CSoutput.n230 CSoutput.n173 4.5005
R6557 CSoutput.n230 CSoutput.n180 4.5005
R6558 CSoutput.n230 CSoutput.n229 4.5005
R6559 CSoutput.n212 CSoutput.n176 4.5005
R6560 CSoutput.n212 CSoutput.n178 4.5005
R6561 CSoutput.n212 CSoutput.n175 4.5005
R6562 CSoutput.n212 CSoutput.n179 4.5005
R6563 CSoutput.n212 CSoutput.n174 4.5005
R6564 CSoutput.n212 CSoutput.t142 4.5005
R6565 CSoutput.n212 CSoutput.n173 4.5005
R6566 CSoutput.n212 CSoutput.n180 4.5005
R6567 CSoutput.n229 CSoutput.n212 4.5005
R6568 CSoutput.n184 CSoutput.n176 4.5005
R6569 CSoutput.n184 CSoutput.n178 4.5005
R6570 CSoutput.n184 CSoutput.n175 4.5005
R6571 CSoutput.n184 CSoutput.n179 4.5005
R6572 CSoutput.n184 CSoutput.n174 4.5005
R6573 CSoutput.n184 CSoutput.t142 4.5005
R6574 CSoutput.n184 CSoutput.n173 4.5005
R6575 CSoutput.n184 CSoutput.n180 4.5005
R6576 CSoutput.n229 CSoutput.n184 4.5005
R6577 CSoutput.n214 CSoutput.n176 4.5005
R6578 CSoutput.n214 CSoutput.n178 4.5005
R6579 CSoutput.n214 CSoutput.n175 4.5005
R6580 CSoutput.n214 CSoutput.n179 4.5005
R6581 CSoutput.n214 CSoutput.n174 4.5005
R6582 CSoutput.n214 CSoutput.t142 4.5005
R6583 CSoutput.n214 CSoutput.n173 4.5005
R6584 CSoutput.n214 CSoutput.n180 4.5005
R6585 CSoutput.n229 CSoutput.n214 4.5005
R6586 CSoutput.n183 CSoutput.n176 4.5005
R6587 CSoutput.n183 CSoutput.n178 4.5005
R6588 CSoutput.n183 CSoutput.n175 4.5005
R6589 CSoutput.n183 CSoutput.n179 4.5005
R6590 CSoutput.n183 CSoutput.n174 4.5005
R6591 CSoutput.n183 CSoutput.t142 4.5005
R6592 CSoutput.n183 CSoutput.n173 4.5005
R6593 CSoutput.n183 CSoutput.n180 4.5005
R6594 CSoutput.n229 CSoutput.n183 4.5005
R6595 CSoutput.n228 CSoutput.n176 4.5005
R6596 CSoutput.n228 CSoutput.n178 4.5005
R6597 CSoutput.n228 CSoutput.n175 4.5005
R6598 CSoutput.n228 CSoutput.n179 4.5005
R6599 CSoutput.n228 CSoutput.n174 4.5005
R6600 CSoutput.n228 CSoutput.t142 4.5005
R6601 CSoutput.n228 CSoutput.n173 4.5005
R6602 CSoutput.n228 CSoutput.n180 4.5005
R6603 CSoutput.n229 CSoutput.n228 4.5005
R6604 CSoutput.n227 CSoutput.n112 4.5005
R6605 CSoutput.n128 CSoutput.n112 4.5005
R6606 CSoutput.n123 CSoutput.n107 4.5005
R6607 CSoutput.n123 CSoutput.n109 4.5005
R6608 CSoutput.n123 CSoutput.n106 4.5005
R6609 CSoutput.n123 CSoutput.n110 4.5005
R6610 CSoutput.n123 CSoutput.n105 4.5005
R6611 CSoutput.n123 CSoutput.t139 4.5005
R6612 CSoutput.n123 CSoutput.n104 4.5005
R6613 CSoutput.n123 CSoutput.n111 4.5005
R6614 CSoutput.n123 CSoutput.n112 4.5005
R6615 CSoutput.n121 CSoutput.n107 4.5005
R6616 CSoutput.n121 CSoutput.n109 4.5005
R6617 CSoutput.n121 CSoutput.n106 4.5005
R6618 CSoutput.n121 CSoutput.n110 4.5005
R6619 CSoutput.n121 CSoutput.n105 4.5005
R6620 CSoutput.n121 CSoutput.t139 4.5005
R6621 CSoutput.n121 CSoutput.n104 4.5005
R6622 CSoutput.n121 CSoutput.n111 4.5005
R6623 CSoutput.n121 CSoutput.n112 4.5005
R6624 CSoutput.n120 CSoutput.n107 4.5005
R6625 CSoutput.n120 CSoutput.n109 4.5005
R6626 CSoutput.n120 CSoutput.n106 4.5005
R6627 CSoutput.n120 CSoutput.n110 4.5005
R6628 CSoutput.n120 CSoutput.n105 4.5005
R6629 CSoutput.n120 CSoutput.t139 4.5005
R6630 CSoutput.n120 CSoutput.n104 4.5005
R6631 CSoutput.n120 CSoutput.n111 4.5005
R6632 CSoutput.n120 CSoutput.n112 4.5005
R6633 CSoutput.n249 CSoutput.n107 4.5005
R6634 CSoutput.n249 CSoutput.n109 4.5005
R6635 CSoutput.n249 CSoutput.n106 4.5005
R6636 CSoutput.n249 CSoutput.n110 4.5005
R6637 CSoutput.n249 CSoutput.n105 4.5005
R6638 CSoutput.n249 CSoutput.t139 4.5005
R6639 CSoutput.n249 CSoutput.n104 4.5005
R6640 CSoutput.n249 CSoutput.n111 4.5005
R6641 CSoutput.n249 CSoutput.n112 4.5005
R6642 CSoutput.n247 CSoutput.n107 4.5005
R6643 CSoutput.n247 CSoutput.n109 4.5005
R6644 CSoutput.n247 CSoutput.n106 4.5005
R6645 CSoutput.n247 CSoutput.n110 4.5005
R6646 CSoutput.n247 CSoutput.n105 4.5005
R6647 CSoutput.n247 CSoutput.t139 4.5005
R6648 CSoutput.n247 CSoutput.n104 4.5005
R6649 CSoutput.n247 CSoutput.n111 4.5005
R6650 CSoutput.n245 CSoutput.n107 4.5005
R6651 CSoutput.n245 CSoutput.n109 4.5005
R6652 CSoutput.n245 CSoutput.n106 4.5005
R6653 CSoutput.n245 CSoutput.n110 4.5005
R6654 CSoutput.n245 CSoutput.n105 4.5005
R6655 CSoutput.n245 CSoutput.t139 4.5005
R6656 CSoutput.n245 CSoutput.n104 4.5005
R6657 CSoutput.n245 CSoutput.n111 4.5005
R6658 CSoutput.n131 CSoutput.n107 4.5005
R6659 CSoutput.n131 CSoutput.n109 4.5005
R6660 CSoutput.n131 CSoutput.n106 4.5005
R6661 CSoutput.n131 CSoutput.n110 4.5005
R6662 CSoutput.n131 CSoutput.n105 4.5005
R6663 CSoutput.n131 CSoutput.t139 4.5005
R6664 CSoutput.n131 CSoutput.n104 4.5005
R6665 CSoutput.n131 CSoutput.n111 4.5005
R6666 CSoutput.n131 CSoutput.n112 4.5005
R6667 CSoutput.n130 CSoutput.n107 4.5005
R6668 CSoutput.n130 CSoutput.n109 4.5005
R6669 CSoutput.n130 CSoutput.n106 4.5005
R6670 CSoutput.n130 CSoutput.n110 4.5005
R6671 CSoutput.n130 CSoutput.n105 4.5005
R6672 CSoutput.n130 CSoutput.t139 4.5005
R6673 CSoutput.n130 CSoutput.n104 4.5005
R6674 CSoutput.n130 CSoutput.n111 4.5005
R6675 CSoutput.n130 CSoutput.n112 4.5005
R6676 CSoutput.n134 CSoutput.n107 4.5005
R6677 CSoutput.n134 CSoutput.n109 4.5005
R6678 CSoutput.n134 CSoutput.n106 4.5005
R6679 CSoutput.n134 CSoutput.n110 4.5005
R6680 CSoutput.n134 CSoutput.n105 4.5005
R6681 CSoutput.n134 CSoutput.t139 4.5005
R6682 CSoutput.n134 CSoutput.n104 4.5005
R6683 CSoutput.n134 CSoutput.n111 4.5005
R6684 CSoutput.n134 CSoutput.n112 4.5005
R6685 CSoutput.n133 CSoutput.n107 4.5005
R6686 CSoutput.n133 CSoutput.n109 4.5005
R6687 CSoutput.n133 CSoutput.n106 4.5005
R6688 CSoutput.n133 CSoutput.n110 4.5005
R6689 CSoutput.n133 CSoutput.n105 4.5005
R6690 CSoutput.n133 CSoutput.t139 4.5005
R6691 CSoutput.n133 CSoutput.n104 4.5005
R6692 CSoutput.n133 CSoutput.n111 4.5005
R6693 CSoutput.n133 CSoutput.n112 4.5005
R6694 CSoutput.n116 CSoutput.n107 4.5005
R6695 CSoutput.n116 CSoutput.n109 4.5005
R6696 CSoutput.n116 CSoutput.n106 4.5005
R6697 CSoutput.n116 CSoutput.n110 4.5005
R6698 CSoutput.n116 CSoutput.n105 4.5005
R6699 CSoutput.n116 CSoutput.t139 4.5005
R6700 CSoutput.n116 CSoutput.n104 4.5005
R6701 CSoutput.n116 CSoutput.n111 4.5005
R6702 CSoutput.n116 CSoutput.n112 4.5005
R6703 CSoutput.n252 CSoutput.n107 4.5005
R6704 CSoutput.n252 CSoutput.n109 4.5005
R6705 CSoutput.n252 CSoutput.n106 4.5005
R6706 CSoutput.n252 CSoutput.n110 4.5005
R6707 CSoutput.n252 CSoutput.n105 4.5005
R6708 CSoutput.n252 CSoutput.t139 4.5005
R6709 CSoutput.n252 CSoutput.n104 4.5005
R6710 CSoutput.n252 CSoutput.n111 4.5005
R6711 CSoutput.n252 CSoutput.n112 4.5005
R6712 CSoutput.n275 CSoutput.n267 4.10845
R6713 CSoutput.n101 CSoutput.n93 4.10845
R6714 CSoutput.n273 CSoutput.t34 4.06363
R6715 CSoutput.n273 CSoutput.t60 4.06363
R6716 CSoutput.n271 CSoutput.t67 4.06363
R6717 CSoutput.n271 CSoutput.t68 4.06363
R6718 CSoutput.n269 CSoutput.t44 4.06363
R6719 CSoutput.n269 CSoutput.t45 4.06363
R6720 CSoutput.n268 CSoutput.t46 4.06363
R6721 CSoutput.n268 CSoutput.t69 4.06363
R6722 CSoutput.n265 CSoutput.t27 4.06363
R6723 CSoutput.n265 CSoutput.t56 4.06363
R6724 CSoutput.n263 CSoutput.t63 4.06363
R6725 CSoutput.n263 CSoutput.t64 4.06363
R6726 CSoutput.n261 CSoutput.t36 4.06363
R6727 CSoutput.n261 CSoutput.t38 4.06363
R6728 CSoutput.n260 CSoutput.t39 4.06363
R6729 CSoutput.n260 CSoutput.t65 4.06363
R6730 CSoutput.n258 CSoutput.t62 4.06363
R6731 CSoutput.n258 CSoutput.t31 4.06363
R6732 CSoutput.n256 CSoutput.t48 4.06363
R6733 CSoutput.n256 CSoutput.t37 4.06363
R6734 CSoutput.n254 CSoutput.t40 4.06363
R6735 CSoutput.n254 CSoutput.t29 4.06363
R6736 CSoutput.n253 CSoutput.t59 4.06363
R6737 CSoutput.n253 CSoutput.t24 4.06363
R6738 CSoutput.n94 CSoutput.t43 4.06363
R6739 CSoutput.n94 CSoutput.t71 4.06363
R6740 CSoutput.n95 CSoutput.t57 4.06363
R6741 CSoutput.n95 CSoutput.t58 4.06363
R6742 CSoutput.n97 CSoutput.t52 4.06363
R6743 CSoutput.n97 CSoutput.t42 4.06363
R6744 CSoutput.n99 CSoutput.t32 4.06363
R6745 CSoutput.n99 CSoutput.t53 4.06363
R6746 CSoutput.n86 CSoutput.t35 4.06363
R6747 CSoutput.n86 CSoutput.t66 4.06363
R6748 CSoutput.n87 CSoutput.t55 4.06363
R6749 CSoutput.n87 CSoutput.t54 4.06363
R6750 CSoutput.n89 CSoutput.t50 4.06363
R6751 CSoutput.n89 CSoutput.t33 4.06363
R6752 CSoutput.n91 CSoutput.t25 4.06363
R6753 CSoutput.n91 CSoutput.t49 4.06363
R6754 CSoutput.n79 CSoutput.t26 4.06363
R6755 CSoutput.n79 CSoutput.t51 4.06363
R6756 CSoutput.n80 CSoutput.t28 4.06363
R6757 CSoutput.n80 CSoutput.t41 4.06363
R6758 CSoutput.n82 CSoutput.t70 4.06363
R6759 CSoutput.n82 CSoutput.t47 4.06363
R6760 CSoutput.n84 CSoutput.t30 4.06363
R6761 CSoutput.n84 CSoutput.t61 4.06363
R6762 CSoutput.n44 CSoutput.n43 3.79402
R6763 CSoutput.n49 CSoutput.n48 3.79402
R6764 CSoutput.n357 CSoutput.n356 3.57343
R6765 CSoutput.n356 CSoutput.n316 3.42304
R6766 CSoutput.n313 CSoutput.t2 2.82907
R6767 CSoutput.n313 CSoutput.t6 2.82907
R6768 CSoutput.n311 CSoutput.t87 2.82907
R6769 CSoutput.n311 CSoutput.t22 2.82907
R6770 CSoutput.n309 CSoutput.t94 2.82907
R6771 CSoutput.n309 CSoutput.t73 2.82907
R6772 CSoutput.n307 CSoutput.t78 2.82907
R6773 CSoutput.n307 CSoutput.t17 2.82907
R6774 CSoutput.n305 CSoutput.t108 2.82907
R6775 CSoutput.n305 CSoutput.t92 2.82907
R6776 CSoutput.n303 CSoutput.t77 2.82907
R6777 CSoutput.n303 CSoutput.t125 2.82907
R6778 CSoutput.n301 CSoutput.t10 2.82907
R6779 CSoutput.n301 CSoutput.t81 2.82907
R6780 CSoutput.n299 CSoutput.t124 2.82907
R6781 CSoutput.n299 CSoutput.t116 2.82907
R6782 CSoutput.n297 CSoutput.t15 2.82907
R6783 CSoutput.n297 CSoutput.t13 2.82907
R6784 CSoutput.n296 CSoutput.t96 2.82907
R6785 CSoutput.n296 CSoutput.t88 2.82907
R6786 CSoutput.n294 CSoutput.t109 2.82907
R6787 CSoutput.n294 CSoutput.t7 2.82907
R6788 CSoutput.n292 CSoutput.t82 2.82907
R6789 CSoutput.n292 CSoutput.t4 2.82907
R6790 CSoutput.n290 CSoutput.t110 2.82907
R6791 CSoutput.n290 CSoutput.t114 2.82907
R6792 CSoutput.n288 CSoutput.t93 2.82907
R6793 CSoutput.n288 CSoutput.t103 2.82907
R6794 CSoutput.n286 CSoutput.t120 2.82907
R6795 CSoutput.n286 CSoutput.t85 2.82907
R6796 CSoutput.n284 CSoutput.t97 2.82907
R6797 CSoutput.n284 CSoutput.t18 2.82907
R6798 CSoutput.n282 CSoutput.t72 2.82907
R6799 CSoutput.n282 CSoutput.t98 2.82907
R6800 CSoutput.n280 CSoutput.t75 2.82907
R6801 CSoutput.n280 CSoutput.t9 2.82907
R6802 CSoutput.n278 CSoutput.t16 2.82907
R6803 CSoutput.n278 CSoutput.t84 2.82907
R6804 CSoutput.n277 CSoutput.t99 2.82907
R6805 CSoutput.n277 CSoutput.t117 2.82907
R6806 CSoutput.n336 CSoutput.t90 2.82907
R6807 CSoutput.n336 CSoutput.t8 2.82907
R6808 CSoutput.n337 CSoutput.t5 2.82907
R6809 CSoutput.n337 CSoutput.t21 2.82907
R6810 CSoutput.n339 CSoutput.t23 2.82907
R6811 CSoutput.n339 CSoutput.t100 2.82907
R6812 CSoutput.n341 CSoutput.t111 2.82907
R6813 CSoutput.n341 CSoutput.t80 2.82907
R6814 CSoutput.n343 CSoutput.t127 2.82907
R6815 CSoutput.n343 CSoutput.t1 2.82907
R6816 CSoutput.n345 CSoutput.t113 2.82907
R6817 CSoutput.n345 CSoutput.t95 2.82907
R6818 CSoutput.n347 CSoutput.t122 2.82907
R6819 CSoutput.n347 CSoutput.t121 2.82907
R6820 CSoutput.n349 CSoutput.t106 2.82907
R6821 CSoutput.n349 CSoutput.t112 2.82907
R6822 CSoutput.n351 CSoutput.t11 2.82907
R6823 CSoutput.n351 CSoutput.t101 2.82907
R6824 CSoutput.n353 CSoutput.t86 2.82907
R6825 CSoutput.n353 CSoutput.t12 2.82907
R6826 CSoutput.n317 CSoutput.t20 2.82907
R6827 CSoutput.n317 CSoutput.t102 2.82907
R6828 CSoutput.n318 CSoutput.t74 2.82907
R6829 CSoutput.n318 CSoutput.t0 2.82907
R6830 CSoutput.n320 CSoutput.t91 2.82907
R6831 CSoutput.n320 CSoutput.t118 2.82907
R6832 CSoutput.n322 CSoutput.t104 2.82907
R6833 CSoutput.n322 CSoutput.t3 2.82907
R6834 CSoutput.n324 CSoutput.t19 2.82907
R6835 CSoutput.n324 CSoutput.t89 2.82907
R6836 CSoutput.n326 CSoutput.t76 2.82907
R6837 CSoutput.n326 CSoutput.t119 2.82907
R6838 CSoutput.n328 CSoutput.t123 2.82907
R6839 CSoutput.n328 CSoutput.t14 2.82907
R6840 CSoutput.n330 CSoutput.t126 2.82907
R6841 CSoutput.n330 CSoutput.t115 2.82907
R6842 CSoutput.n332 CSoutput.t107 2.82907
R6843 CSoutput.n332 CSoutput.t83 2.82907
R6844 CSoutput.n334 CSoutput.t79 2.82907
R6845 CSoutput.n334 CSoutput.t105 2.82907
R6846 CSoutput.n75 CSoutput.n1 2.45513
R6847 CSoutput.n276 CSoutput.n102 2.36742
R6848 CSoutput.n193 CSoutput.n191 2.251
R6849 CSoutput.n193 CSoutput.n190 2.251
R6850 CSoutput.n193 CSoutput.n189 2.251
R6851 CSoutput.n193 CSoutput.n188 2.251
R6852 CSoutput.n162 CSoutput.n161 2.251
R6853 CSoutput.n162 CSoutput.n160 2.251
R6854 CSoutput.n162 CSoutput.n159 2.251
R6855 CSoutput.n162 CSoutput.n158 2.251
R6856 CSoutput.n235 CSoutput.n234 2.251
R6857 CSoutput.n200 CSoutput.n198 2.251
R6858 CSoutput.n200 CSoutput.n197 2.251
R6859 CSoutput.n200 CSoutput.n196 2.251
R6860 CSoutput.n218 CSoutput.n200 2.251
R6861 CSoutput.n206 CSoutput.n205 2.251
R6862 CSoutput.n206 CSoutput.n204 2.251
R6863 CSoutput.n206 CSoutput.n203 2.251
R6864 CSoutput.n206 CSoutput.n202 2.251
R6865 CSoutput.n232 CSoutput.n172 2.251
R6866 CSoutput.n227 CSoutput.n225 2.251
R6867 CSoutput.n227 CSoutput.n224 2.251
R6868 CSoutput.n227 CSoutput.n223 2.251
R6869 CSoutput.n227 CSoutput.n222 2.251
R6870 CSoutput.n128 CSoutput.n127 2.251
R6871 CSoutput.n128 CSoutput.n126 2.251
R6872 CSoutput.n128 CSoutput.n125 2.251
R6873 CSoutput.n128 CSoutput.n124 2.251
R6874 CSoutput.n245 CSoutput.n244 2.251
R6875 CSoutput.n162 CSoutput.n142 2.2505
R6876 CSoutput.n157 CSoutput.n142 2.2505
R6877 CSoutput.n155 CSoutput.n142 2.2505
R6878 CSoutput.n154 CSoutput.n142 2.2505
R6879 CSoutput.n239 CSoutput.n142 2.2505
R6880 CSoutput.n237 CSoutput.n142 2.2505
R6881 CSoutput.n235 CSoutput.n142 2.2505
R6882 CSoutput.n165 CSoutput.n142 2.2505
R6883 CSoutput.n164 CSoutput.n142 2.2505
R6884 CSoutput.n168 CSoutput.n142 2.2505
R6885 CSoutput.n167 CSoutput.n142 2.2505
R6886 CSoutput.n150 CSoutput.n142 2.2505
R6887 CSoutput.n242 CSoutput.n142 2.2505
R6888 CSoutput.n242 CSoutput.n241 2.2505
R6889 CSoutput.n206 CSoutput.n177 2.2505
R6890 CSoutput.n187 CSoutput.n177 2.2505
R6891 CSoutput.n208 CSoutput.n177 2.2505
R6892 CSoutput.n186 CSoutput.n177 2.2505
R6893 CSoutput.n210 CSoutput.n177 2.2505
R6894 CSoutput.n177 CSoutput.n171 2.2505
R6895 CSoutput.n232 CSoutput.n177 2.2505
R6896 CSoutput.n230 CSoutput.n177 2.2505
R6897 CSoutput.n212 CSoutput.n177 2.2505
R6898 CSoutput.n184 CSoutput.n177 2.2505
R6899 CSoutput.n214 CSoutput.n177 2.2505
R6900 CSoutput.n183 CSoutput.n177 2.2505
R6901 CSoutput.n228 CSoutput.n177 2.2505
R6902 CSoutput.n228 CSoutput.n181 2.2505
R6903 CSoutput.n128 CSoutput.n108 2.2505
R6904 CSoutput.n123 CSoutput.n108 2.2505
R6905 CSoutput.n121 CSoutput.n108 2.2505
R6906 CSoutput.n120 CSoutput.n108 2.2505
R6907 CSoutput.n249 CSoutput.n108 2.2505
R6908 CSoutput.n247 CSoutput.n108 2.2505
R6909 CSoutput.n245 CSoutput.n108 2.2505
R6910 CSoutput.n131 CSoutput.n108 2.2505
R6911 CSoutput.n130 CSoutput.n108 2.2505
R6912 CSoutput.n134 CSoutput.n108 2.2505
R6913 CSoutput.n133 CSoutput.n108 2.2505
R6914 CSoutput.n116 CSoutput.n108 2.2505
R6915 CSoutput.n252 CSoutput.n108 2.2505
R6916 CSoutput.n252 CSoutput.n251 2.2505
R6917 CSoutput.n170 CSoutput.n163 2.25024
R6918 CSoutput.n170 CSoutput.n156 2.25024
R6919 CSoutput.n238 CSoutput.n170 2.25024
R6920 CSoutput.n170 CSoutput.n166 2.25024
R6921 CSoutput.n170 CSoutput.n169 2.25024
R6922 CSoutput.n170 CSoutput.n137 2.25024
R6923 CSoutput.n220 CSoutput.n217 2.25024
R6924 CSoutput.n220 CSoutput.n216 2.25024
R6925 CSoutput.n220 CSoutput.n215 2.25024
R6926 CSoutput.n220 CSoutput.n182 2.25024
R6927 CSoutput.n220 CSoutput.n219 2.25024
R6928 CSoutput.n221 CSoutput.n220 2.25024
R6929 CSoutput.n136 CSoutput.n129 2.25024
R6930 CSoutput.n136 CSoutput.n122 2.25024
R6931 CSoutput.n248 CSoutput.n136 2.25024
R6932 CSoutput.n136 CSoutput.n132 2.25024
R6933 CSoutput.n136 CSoutput.n135 2.25024
R6934 CSoutput.n136 CSoutput.n103 2.25024
R6935 CSoutput.n237 CSoutput.n147 1.50111
R6936 CSoutput.n185 CSoutput.n171 1.50111
R6937 CSoutput.n247 CSoutput.n113 1.50111
R6938 CSoutput.n193 CSoutput.n192 1.501
R6939 CSoutput.n200 CSoutput.n199 1.501
R6940 CSoutput.n227 CSoutput.n226 1.501
R6941 CSoutput.n241 CSoutput.n152 1.12536
R6942 CSoutput.n241 CSoutput.n153 1.12536
R6943 CSoutput.n241 CSoutput.n240 1.12536
R6944 CSoutput.n201 CSoutput.n181 1.12536
R6945 CSoutput.n207 CSoutput.n181 1.12536
R6946 CSoutput.n209 CSoutput.n181 1.12536
R6947 CSoutput.n251 CSoutput.n118 1.12536
R6948 CSoutput.n251 CSoutput.n119 1.12536
R6949 CSoutput.n251 CSoutput.n250 1.12536
R6950 CSoutput.n241 CSoutput.n148 1.12536
R6951 CSoutput.n241 CSoutput.n149 1.12536
R6952 CSoutput.n241 CSoutput.n151 1.12536
R6953 CSoutput.n231 CSoutput.n181 1.12536
R6954 CSoutput.n211 CSoutput.n181 1.12536
R6955 CSoutput.n213 CSoutput.n181 1.12536
R6956 CSoutput.n251 CSoutput.n114 1.12536
R6957 CSoutput.n251 CSoutput.n115 1.12536
R6958 CSoutput.n251 CSoutput.n117 1.12536
R6959 CSoutput.n31 CSoutput.n30 0.669944
R6960 CSoutput.n62 CSoutput.n61 0.669944
R6961 CSoutput.n300 CSoutput.n298 0.573776
R6962 CSoutput.n302 CSoutput.n300 0.573776
R6963 CSoutput.n304 CSoutput.n302 0.573776
R6964 CSoutput.n306 CSoutput.n304 0.573776
R6965 CSoutput.n308 CSoutput.n306 0.573776
R6966 CSoutput.n310 CSoutput.n308 0.573776
R6967 CSoutput.n312 CSoutput.n310 0.573776
R6968 CSoutput.n314 CSoutput.n312 0.573776
R6969 CSoutput.n281 CSoutput.n279 0.573776
R6970 CSoutput.n283 CSoutput.n281 0.573776
R6971 CSoutput.n285 CSoutput.n283 0.573776
R6972 CSoutput.n287 CSoutput.n285 0.573776
R6973 CSoutput.n289 CSoutput.n287 0.573776
R6974 CSoutput.n291 CSoutput.n289 0.573776
R6975 CSoutput.n293 CSoutput.n291 0.573776
R6976 CSoutput.n295 CSoutput.n293 0.573776
R6977 CSoutput.n354 CSoutput.n352 0.573776
R6978 CSoutput.n352 CSoutput.n350 0.573776
R6979 CSoutput.n350 CSoutput.n348 0.573776
R6980 CSoutput.n348 CSoutput.n346 0.573776
R6981 CSoutput.n346 CSoutput.n344 0.573776
R6982 CSoutput.n344 CSoutput.n342 0.573776
R6983 CSoutput.n342 CSoutput.n340 0.573776
R6984 CSoutput.n340 CSoutput.n338 0.573776
R6985 CSoutput.n335 CSoutput.n333 0.573776
R6986 CSoutput.n333 CSoutput.n331 0.573776
R6987 CSoutput.n331 CSoutput.n329 0.573776
R6988 CSoutput.n329 CSoutput.n327 0.573776
R6989 CSoutput.n327 CSoutput.n325 0.573776
R6990 CSoutput.n325 CSoutput.n323 0.573776
R6991 CSoutput.n323 CSoutput.n321 0.573776
R6992 CSoutput.n321 CSoutput.n319 0.573776
R6993 CSoutput.n357 CSoutput.n252 0.53442
R6994 CSoutput.n272 CSoutput.n270 0.358259
R6995 CSoutput.n274 CSoutput.n272 0.358259
R6996 CSoutput.n264 CSoutput.n262 0.358259
R6997 CSoutput.n266 CSoutput.n264 0.358259
R6998 CSoutput.n257 CSoutput.n255 0.358259
R6999 CSoutput.n259 CSoutput.n257 0.358259
R7000 CSoutput.n100 CSoutput.n98 0.358259
R7001 CSoutput.n98 CSoutput.n96 0.358259
R7002 CSoutput.n92 CSoutput.n90 0.358259
R7003 CSoutput.n90 CSoutput.n88 0.358259
R7004 CSoutput.n85 CSoutput.n83 0.358259
R7005 CSoutput.n83 CSoutput.n81 0.358259
R7006 CSoutput.n21 CSoutput.n20 0.169105
R7007 CSoutput.n21 CSoutput.n16 0.169105
R7008 CSoutput.n26 CSoutput.n16 0.169105
R7009 CSoutput.n27 CSoutput.n26 0.169105
R7010 CSoutput.n27 CSoutput.n14 0.169105
R7011 CSoutput.n32 CSoutput.n14 0.169105
R7012 CSoutput.n33 CSoutput.n32 0.169105
R7013 CSoutput.n34 CSoutput.n33 0.169105
R7014 CSoutput.n34 CSoutput.n12 0.169105
R7015 CSoutput.n39 CSoutput.n12 0.169105
R7016 CSoutput.n40 CSoutput.n39 0.169105
R7017 CSoutput.n40 CSoutput.n10 0.169105
R7018 CSoutput.n45 CSoutput.n10 0.169105
R7019 CSoutput.n46 CSoutput.n45 0.169105
R7020 CSoutput.n47 CSoutput.n46 0.169105
R7021 CSoutput.n47 CSoutput.n8 0.169105
R7022 CSoutput.n52 CSoutput.n8 0.169105
R7023 CSoutput.n53 CSoutput.n52 0.169105
R7024 CSoutput.n53 CSoutput.n6 0.169105
R7025 CSoutput.n58 CSoutput.n6 0.169105
R7026 CSoutput.n59 CSoutput.n58 0.169105
R7027 CSoutput.n60 CSoutput.n59 0.169105
R7028 CSoutput.n60 CSoutput.n4 0.169105
R7029 CSoutput.n66 CSoutput.n4 0.169105
R7030 CSoutput.n67 CSoutput.n66 0.169105
R7031 CSoutput.n68 CSoutput.n67 0.169105
R7032 CSoutput.n68 CSoutput.n2 0.169105
R7033 CSoutput.n73 CSoutput.n2 0.169105
R7034 CSoutput.n74 CSoutput.n73 0.169105
R7035 CSoutput.n74 CSoutput.n0 0.169105
R7036 CSoutput.n78 CSoutput.n0 0.169105
R7037 CSoutput.n195 CSoutput.n194 0.0910737
R7038 CSoutput.n246 CSoutput.n243 0.0723685
R7039 CSoutput.n200 CSoutput.n195 0.0522944
R7040 CSoutput.n243 CSoutput.n242 0.0499135
R7041 CSoutput.n194 CSoutput.n193 0.0499135
R7042 CSoutput.n228 CSoutput.n227 0.0464294
R7043 CSoutput.n236 CSoutput.n233 0.0391444
R7044 CSoutput.n195 CSoutput.t128 0.023435
R7045 CSoutput.n243 CSoutput.t132 0.02262
R7046 CSoutput.n194 CSoutput.t135 0.02262
R7047 CSoutput CSoutput.n357 0.0052
R7048 CSoutput.n165 CSoutput.n148 0.00365111
R7049 CSoutput.n168 CSoutput.n149 0.00365111
R7050 CSoutput.n151 CSoutput.n150 0.00365111
R7051 CSoutput.n193 CSoutput.n152 0.00365111
R7052 CSoutput.n157 CSoutput.n153 0.00365111
R7053 CSoutput.n240 CSoutput.n154 0.00365111
R7054 CSoutput.n231 CSoutput.n230 0.00365111
R7055 CSoutput.n211 CSoutput.n184 0.00365111
R7056 CSoutput.n213 CSoutput.n183 0.00365111
R7057 CSoutput.n201 CSoutput.n200 0.00365111
R7058 CSoutput.n207 CSoutput.n187 0.00365111
R7059 CSoutput.n209 CSoutput.n186 0.00365111
R7060 CSoutput.n131 CSoutput.n114 0.00365111
R7061 CSoutput.n134 CSoutput.n115 0.00365111
R7062 CSoutput.n117 CSoutput.n116 0.00365111
R7063 CSoutput.n227 CSoutput.n118 0.00365111
R7064 CSoutput.n123 CSoutput.n119 0.00365111
R7065 CSoutput.n250 CSoutput.n120 0.00365111
R7066 CSoutput.n162 CSoutput.n152 0.00340054
R7067 CSoutput.n155 CSoutput.n153 0.00340054
R7068 CSoutput.n240 CSoutput.n239 0.00340054
R7069 CSoutput.n235 CSoutput.n148 0.00340054
R7070 CSoutput.n164 CSoutput.n149 0.00340054
R7071 CSoutput.n167 CSoutput.n151 0.00340054
R7072 CSoutput.n206 CSoutput.n201 0.00340054
R7073 CSoutput.n208 CSoutput.n207 0.00340054
R7074 CSoutput.n210 CSoutput.n209 0.00340054
R7075 CSoutput.n232 CSoutput.n231 0.00340054
R7076 CSoutput.n212 CSoutput.n211 0.00340054
R7077 CSoutput.n214 CSoutput.n213 0.00340054
R7078 CSoutput.n128 CSoutput.n118 0.00340054
R7079 CSoutput.n121 CSoutput.n119 0.00340054
R7080 CSoutput.n250 CSoutput.n249 0.00340054
R7081 CSoutput.n245 CSoutput.n114 0.00340054
R7082 CSoutput.n130 CSoutput.n115 0.00340054
R7083 CSoutput.n133 CSoutput.n117 0.00340054
R7084 CSoutput.n163 CSoutput.n157 0.00252698
R7085 CSoutput.n156 CSoutput.n154 0.00252698
R7086 CSoutput.n238 CSoutput.n237 0.00252698
R7087 CSoutput.n166 CSoutput.n164 0.00252698
R7088 CSoutput.n169 CSoutput.n167 0.00252698
R7089 CSoutput.n242 CSoutput.n137 0.00252698
R7090 CSoutput.n163 CSoutput.n162 0.00252698
R7091 CSoutput.n156 CSoutput.n155 0.00252698
R7092 CSoutput.n239 CSoutput.n238 0.00252698
R7093 CSoutput.n166 CSoutput.n165 0.00252698
R7094 CSoutput.n169 CSoutput.n168 0.00252698
R7095 CSoutput.n150 CSoutput.n137 0.00252698
R7096 CSoutput.n217 CSoutput.n187 0.00252698
R7097 CSoutput.n216 CSoutput.n186 0.00252698
R7098 CSoutput.n215 CSoutput.n171 0.00252698
R7099 CSoutput.n212 CSoutput.n182 0.00252698
R7100 CSoutput.n219 CSoutput.n214 0.00252698
R7101 CSoutput.n228 CSoutput.n221 0.00252698
R7102 CSoutput.n217 CSoutput.n206 0.00252698
R7103 CSoutput.n216 CSoutput.n208 0.00252698
R7104 CSoutput.n215 CSoutput.n210 0.00252698
R7105 CSoutput.n230 CSoutput.n182 0.00252698
R7106 CSoutput.n219 CSoutput.n184 0.00252698
R7107 CSoutput.n221 CSoutput.n183 0.00252698
R7108 CSoutput.n129 CSoutput.n123 0.00252698
R7109 CSoutput.n122 CSoutput.n120 0.00252698
R7110 CSoutput.n248 CSoutput.n247 0.00252698
R7111 CSoutput.n132 CSoutput.n130 0.00252698
R7112 CSoutput.n135 CSoutput.n133 0.00252698
R7113 CSoutput.n252 CSoutput.n103 0.00252698
R7114 CSoutput.n129 CSoutput.n128 0.00252698
R7115 CSoutput.n122 CSoutput.n121 0.00252698
R7116 CSoutput.n249 CSoutput.n248 0.00252698
R7117 CSoutput.n132 CSoutput.n131 0.00252698
R7118 CSoutput.n135 CSoutput.n134 0.00252698
R7119 CSoutput.n116 CSoutput.n103 0.00252698
R7120 CSoutput.n237 CSoutput.n236 0.0020275
R7121 CSoutput.n236 CSoutput.n235 0.0020275
R7122 CSoutput.n233 CSoutput.n171 0.0020275
R7123 CSoutput.n233 CSoutput.n232 0.0020275
R7124 CSoutput.n247 CSoutput.n246 0.0020275
R7125 CSoutput.n246 CSoutput.n245 0.0020275
R7126 CSoutput.n147 CSoutput.n146 0.00166668
R7127 CSoutput.n229 CSoutput.n185 0.00166668
R7128 CSoutput.n113 CSoutput.n112 0.00166668
R7129 CSoutput.n251 CSoutput.n113 0.00133328
R7130 CSoutput.n185 CSoutput.n181 0.00133328
R7131 CSoutput.n241 CSoutput.n147 0.00133328
R7132 CSoutput.n244 CSoutput.n136 0.001
R7133 CSoutput.n222 CSoutput.n136 0.001
R7134 CSoutput.n124 CSoutput.n104 0.001
R7135 CSoutput.n223 CSoutput.n104 0.001
R7136 CSoutput.n125 CSoutput.n105 0.001
R7137 CSoutput.n224 CSoutput.n105 0.001
R7138 CSoutput.n126 CSoutput.n106 0.001
R7139 CSoutput.n225 CSoutput.n106 0.001
R7140 CSoutput.n127 CSoutput.n107 0.001
R7141 CSoutput.n226 CSoutput.n107 0.001
R7142 CSoutput.n220 CSoutput.n172 0.001
R7143 CSoutput.n220 CSoutput.n218 0.001
R7144 CSoutput.n202 CSoutput.n173 0.001
R7145 CSoutput.n196 CSoutput.n173 0.001
R7146 CSoutput.n203 CSoutput.n174 0.001
R7147 CSoutput.n197 CSoutput.n174 0.001
R7148 CSoutput.n204 CSoutput.n175 0.001
R7149 CSoutput.n198 CSoutput.n175 0.001
R7150 CSoutput.n205 CSoutput.n176 0.001
R7151 CSoutput.n199 CSoutput.n176 0.001
R7152 CSoutput.n234 CSoutput.n170 0.001
R7153 CSoutput.n188 CSoutput.n170 0.001
R7154 CSoutput.n158 CSoutput.n138 0.001
R7155 CSoutput.n189 CSoutput.n138 0.001
R7156 CSoutput.n159 CSoutput.n139 0.001
R7157 CSoutput.n190 CSoutput.n139 0.001
R7158 CSoutput.n160 CSoutput.n140 0.001
R7159 CSoutput.n191 CSoutput.n140 0.001
R7160 CSoutput.n161 CSoutput.n141 0.001
R7161 CSoutput.n192 CSoutput.n141 0.001
R7162 CSoutput.n192 CSoutput.n142 0.001
R7163 CSoutput.n191 CSoutput.n143 0.001
R7164 CSoutput.n190 CSoutput.n144 0.001
R7165 CSoutput.n189 CSoutput.t148 0.001
R7166 CSoutput.n188 CSoutput.n145 0.001
R7167 CSoutput.n161 CSoutput.n143 0.001
R7168 CSoutput.n160 CSoutput.n144 0.001
R7169 CSoutput.n159 CSoutput.t148 0.001
R7170 CSoutput.n158 CSoutput.n145 0.001
R7171 CSoutput.n234 CSoutput.n146 0.001
R7172 CSoutput.n199 CSoutput.n177 0.001
R7173 CSoutput.n198 CSoutput.n178 0.001
R7174 CSoutput.n197 CSoutput.n179 0.001
R7175 CSoutput.n196 CSoutput.t142 0.001
R7176 CSoutput.n218 CSoutput.n180 0.001
R7177 CSoutput.n205 CSoutput.n178 0.001
R7178 CSoutput.n204 CSoutput.n179 0.001
R7179 CSoutput.n203 CSoutput.t142 0.001
R7180 CSoutput.n202 CSoutput.n180 0.001
R7181 CSoutput.n229 CSoutput.n172 0.001
R7182 CSoutput.n226 CSoutput.n108 0.001
R7183 CSoutput.n225 CSoutput.n109 0.001
R7184 CSoutput.n224 CSoutput.n110 0.001
R7185 CSoutput.n223 CSoutput.t139 0.001
R7186 CSoutput.n222 CSoutput.n111 0.001
R7187 CSoutput.n127 CSoutput.n109 0.001
R7188 CSoutput.n126 CSoutput.n110 0.001
R7189 CSoutput.n125 CSoutput.t139 0.001
R7190 CSoutput.n124 CSoutput.n111 0.001
R7191 CSoutput.n244 CSoutput.n112 0.001
R7192 commonsourceibias.n281 commonsourceibias.t101 222.032
R7193 commonsourceibias.n44 commonsourceibias.t32 222.032
R7194 commonsourceibias.n166 commonsourceibias.t117 222.032
R7195 commonsourceibias.n643 commonsourceibias.t108 222.032
R7196 commonsourceibias.n413 commonsourceibias.t0 222.032
R7197 commonsourceibias.n529 commonsourceibias.t125 222.032
R7198 commonsourceibias.n364 commonsourceibias.t102 207.983
R7199 commonsourceibias.n127 commonsourceibias.t12 207.983
R7200 commonsourceibias.n249 commonsourceibias.t118 207.983
R7201 commonsourceibias.n731 commonsourceibias.t123 207.983
R7202 commonsourceibias.n501 commonsourceibias.t58 207.983
R7203 commonsourceibias.n616 commonsourceibias.t139 207.983
R7204 commonsourceibias.n280 commonsourceibias.t152 168.701
R7205 commonsourceibias.n286 commonsourceibias.t155 168.701
R7206 commonsourceibias.n292 commonsourceibias.t112 168.701
R7207 commonsourceibias.n276 commonsourceibias.t97 168.701
R7208 commonsourceibias.n300 commonsourceibias.t85 168.701
R7209 commonsourceibias.n306 commonsourceibias.t122 168.701
R7210 commonsourceibias.n271 commonsourceibias.t104 168.701
R7211 commonsourceibias.n314 commonsourceibias.t91 168.701
R7212 commonsourceibias.n320 commonsourceibias.t94 168.701
R7213 commonsourceibias.n266 commonsourceibias.t113 168.701
R7214 commonsourceibias.n328 commonsourceibias.t96 168.701
R7215 commonsourceibias.n334 commonsourceibias.t100 168.701
R7216 commonsourceibias.n261 commonsourceibias.t151 168.701
R7217 commonsourceibias.n342 commonsourceibias.t129 168.701
R7218 commonsourceibias.n348 commonsourceibias.t109 168.701
R7219 commonsourceibias.n256 commonsourceibias.t159 168.701
R7220 commonsourceibias.n356 commonsourceibias.t81 168.701
R7221 commonsourceibias.n362 commonsourceibias.t120 168.701
R7222 commonsourceibias.n125 commonsourceibias.t66 168.701
R7223 commonsourceibias.n119 commonsourceibias.t42 168.701
R7224 commonsourceibias.n19 commonsourceibias.t10 168.701
R7225 commonsourceibias.n111 commonsourceibias.t46 168.701
R7226 commonsourceibias.n105 commonsourceibias.t16 168.701
R7227 commonsourceibias.n24 commonsourceibias.t36 168.701
R7228 commonsourceibias.n97 commonsourceibias.t22 168.701
R7229 commonsourceibias.n91 commonsourceibias.t14 168.701
R7230 commonsourceibias.n29 commonsourceibias.t54 168.701
R7231 commonsourceibias.n83 commonsourceibias.t76 168.701
R7232 commonsourceibias.n77 commonsourceibias.t38 168.701
R7233 commonsourceibias.n34 commonsourceibias.t8 168.701
R7234 commonsourceibias.n69 commonsourceibias.t28 168.701
R7235 commonsourceibias.n63 commonsourceibias.t68 168.701
R7236 commonsourceibias.n39 commonsourceibias.t18 168.701
R7237 commonsourceibias.n55 commonsourceibias.t60 168.701
R7238 commonsourceibias.n49 commonsourceibias.t52 168.701
R7239 commonsourceibias.n43 commonsourceibias.t64 168.701
R7240 commonsourceibias.n247 commonsourceibias.t135 168.701
R7241 commonsourceibias.n241 commonsourceibias.t92 168.701
R7242 commonsourceibias.n5 commonsourceibias.t90 168.701
R7243 commonsourceibias.n233 commonsourceibias.t127 168.701
R7244 commonsourceibias.n227 commonsourceibias.t143 168.701
R7245 commonsourceibias.n10 commonsourceibias.t84 168.701
R7246 commonsourceibias.n219 commonsourceibias.t115 168.701
R7247 commonsourceibias.n213 commonsourceibias.t111 168.701
R7248 commonsourceibias.n150 commonsourceibias.t131 168.701
R7249 commonsourceibias.n151 commonsourceibias.t106 168.701
R7250 commonsourceibias.n153 commonsourceibias.t103 168.701
R7251 commonsourceibias.n155 commonsourceibias.t121 168.701
R7252 commonsourceibias.n191 commonsourceibias.t138 168.701
R7253 commonsourceibias.n185 commonsourceibias.t95 168.701
R7254 commonsourceibias.n161 commonsourceibias.t110 168.701
R7255 commonsourceibias.n177 commonsourceibias.t130 168.701
R7256 commonsourceibias.n171 commonsourceibias.t87 168.701
R7257 commonsourceibias.n165 commonsourceibias.t83 168.701
R7258 commonsourceibias.n642 commonsourceibias.t158 168.701
R7259 commonsourceibias.n648 commonsourceibias.t150 168.701
R7260 commonsourceibias.n654 commonsourceibias.t137 168.701
R7261 commonsourceibias.n656 commonsourceibias.t119 168.701
R7262 commonsourceibias.n663 commonsourceibias.t99 168.701
R7263 commonsourceibias.n669 commonsourceibias.t145 168.701
R7264 commonsourceibias.n671 commonsourceibias.t128 168.701
R7265 commonsourceibias.n678 commonsourceibias.t107 168.701
R7266 commonsourceibias.n684 commonsourceibias.t88 168.701
R7267 commonsourceibias.n686 commonsourceibias.t136 168.701
R7268 commonsourceibias.n693 commonsourceibias.t116 168.701
R7269 commonsourceibias.n699 commonsourceibias.t124 168.701
R7270 commonsourceibias.n701 commonsourceibias.t144 168.701
R7271 commonsourceibias.n708 commonsourceibias.t147 168.701
R7272 commonsourceibias.n714 commonsourceibias.t132 168.701
R7273 commonsourceibias.n716 commonsourceibias.t93 168.701
R7274 commonsourceibias.n723 commonsourceibias.t154 168.701
R7275 commonsourceibias.n729 commonsourceibias.t141 168.701
R7276 commonsourceibias.n412 commonsourceibias.t20 168.701
R7277 commonsourceibias.n418 commonsourceibias.t44 168.701
R7278 commonsourceibias.n424 commonsourceibias.t6 168.701
R7279 commonsourceibias.n426 commonsourceibias.t34 168.701
R7280 commonsourceibias.n433 commonsourceibias.t26 168.701
R7281 commonsourceibias.n439 commonsourceibias.t72 168.701
R7282 commonsourceibias.n441 commonsourceibias.t40 168.701
R7283 commonsourceibias.n448 commonsourceibias.t4 168.701
R7284 commonsourceibias.n454 commonsourceibias.t74 168.701
R7285 commonsourceibias.n456 commonsourceibias.t2 168.701
R7286 commonsourceibias.n463 commonsourceibias.t62 168.701
R7287 commonsourceibias.n469 commonsourceibias.t78 168.701
R7288 commonsourceibias.n471 commonsourceibias.t50 168.701
R7289 commonsourceibias.n478 commonsourceibias.t70 168.701
R7290 commonsourceibias.n484 commonsourceibias.t24 168.701
R7291 commonsourceibias.n486 commonsourceibias.t56 168.701
R7292 commonsourceibias.n493 commonsourceibias.t30 168.701
R7293 commonsourceibias.n499 commonsourceibias.t48 168.701
R7294 commonsourceibias.n614 commonsourceibias.t153 168.701
R7295 commonsourceibias.n608 commonsourceibias.t86 168.701
R7296 commonsourceibias.n601 commonsourceibias.t105 168.701
R7297 commonsourceibias.n599 commonsourceibias.t146 168.701
R7298 commonsourceibias.n593 commonsourceibias.t80 168.701
R7299 commonsourceibias.n586 commonsourceibias.t157 168.701
R7300 commonsourceibias.n584 commonsourceibias.t140 168.701
R7301 commonsourceibias.n578 commonsourceibias.t133 168.701
R7302 commonsourceibias.n571 commonsourceibias.t149 168.701
R7303 commonsourceibias.n528 commonsourceibias.t89 168.701
R7304 commonsourceibias.n534 commonsourceibias.t82 168.701
R7305 commonsourceibias.n540 commonsourceibias.t148 168.701
R7306 commonsourceibias.n542 commonsourceibias.t134 168.701
R7307 commonsourceibias.n549 commonsourceibias.t114 168.701
R7308 commonsourceibias.n555 commonsourceibias.t156 168.701
R7309 commonsourceibias.n519 commonsourceibias.t142 168.701
R7310 commonsourceibias.n517 commonsourceibias.t126 168.701
R7311 commonsourceibias.n515 commonsourceibias.t98 168.701
R7312 commonsourceibias.n363 commonsourceibias.n251 161.3
R7313 commonsourceibias.n361 commonsourceibias.n360 161.3
R7314 commonsourceibias.n359 commonsourceibias.n252 161.3
R7315 commonsourceibias.n358 commonsourceibias.n357 161.3
R7316 commonsourceibias.n355 commonsourceibias.n253 161.3
R7317 commonsourceibias.n354 commonsourceibias.n353 161.3
R7318 commonsourceibias.n352 commonsourceibias.n254 161.3
R7319 commonsourceibias.n351 commonsourceibias.n350 161.3
R7320 commonsourceibias.n349 commonsourceibias.n255 161.3
R7321 commonsourceibias.n347 commonsourceibias.n346 161.3
R7322 commonsourceibias.n345 commonsourceibias.n257 161.3
R7323 commonsourceibias.n344 commonsourceibias.n343 161.3
R7324 commonsourceibias.n341 commonsourceibias.n258 161.3
R7325 commonsourceibias.n340 commonsourceibias.n339 161.3
R7326 commonsourceibias.n338 commonsourceibias.n259 161.3
R7327 commonsourceibias.n337 commonsourceibias.n336 161.3
R7328 commonsourceibias.n335 commonsourceibias.n260 161.3
R7329 commonsourceibias.n333 commonsourceibias.n332 161.3
R7330 commonsourceibias.n331 commonsourceibias.n262 161.3
R7331 commonsourceibias.n330 commonsourceibias.n329 161.3
R7332 commonsourceibias.n327 commonsourceibias.n263 161.3
R7333 commonsourceibias.n326 commonsourceibias.n325 161.3
R7334 commonsourceibias.n324 commonsourceibias.n264 161.3
R7335 commonsourceibias.n323 commonsourceibias.n322 161.3
R7336 commonsourceibias.n321 commonsourceibias.n265 161.3
R7337 commonsourceibias.n319 commonsourceibias.n318 161.3
R7338 commonsourceibias.n317 commonsourceibias.n267 161.3
R7339 commonsourceibias.n316 commonsourceibias.n315 161.3
R7340 commonsourceibias.n313 commonsourceibias.n268 161.3
R7341 commonsourceibias.n312 commonsourceibias.n311 161.3
R7342 commonsourceibias.n310 commonsourceibias.n269 161.3
R7343 commonsourceibias.n309 commonsourceibias.n308 161.3
R7344 commonsourceibias.n307 commonsourceibias.n270 161.3
R7345 commonsourceibias.n305 commonsourceibias.n304 161.3
R7346 commonsourceibias.n303 commonsourceibias.n272 161.3
R7347 commonsourceibias.n302 commonsourceibias.n301 161.3
R7348 commonsourceibias.n299 commonsourceibias.n273 161.3
R7349 commonsourceibias.n298 commonsourceibias.n297 161.3
R7350 commonsourceibias.n296 commonsourceibias.n274 161.3
R7351 commonsourceibias.n295 commonsourceibias.n294 161.3
R7352 commonsourceibias.n293 commonsourceibias.n275 161.3
R7353 commonsourceibias.n291 commonsourceibias.n290 161.3
R7354 commonsourceibias.n289 commonsourceibias.n277 161.3
R7355 commonsourceibias.n288 commonsourceibias.n287 161.3
R7356 commonsourceibias.n285 commonsourceibias.n278 161.3
R7357 commonsourceibias.n284 commonsourceibias.n283 161.3
R7358 commonsourceibias.n282 commonsourceibias.n279 161.3
R7359 commonsourceibias.n45 commonsourceibias.n42 161.3
R7360 commonsourceibias.n47 commonsourceibias.n46 161.3
R7361 commonsourceibias.n48 commonsourceibias.n41 161.3
R7362 commonsourceibias.n51 commonsourceibias.n50 161.3
R7363 commonsourceibias.n52 commonsourceibias.n40 161.3
R7364 commonsourceibias.n54 commonsourceibias.n53 161.3
R7365 commonsourceibias.n56 commonsourceibias.n38 161.3
R7366 commonsourceibias.n58 commonsourceibias.n57 161.3
R7367 commonsourceibias.n59 commonsourceibias.n37 161.3
R7368 commonsourceibias.n61 commonsourceibias.n60 161.3
R7369 commonsourceibias.n62 commonsourceibias.n36 161.3
R7370 commonsourceibias.n65 commonsourceibias.n64 161.3
R7371 commonsourceibias.n66 commonsourceibias.n35 161.3
R7372 commonsourceibias.n68 commonsourceibias.n67 161.3
R7373 commonsourceibias.n70 commonsourceibias.n33 161.3
R7374 commonsourceibias.n72 commonsourceibias.n71 161.3
R7375 commonsourceibias.n73 commonsourceibias.n32 161.3
R7376 commonsourceibias.n75 commonsourceibias.n74 161.3
R7377 commonsourceibias.n76 commonsourceibias.n31 161.3
R7378 commonsourceibias.n79 commonsourceibias.n78 161.3
R7379 commonsourceibias.n80 commonsourceibias.n30 161.3
R7380 commonsourceibias.n82 commonsourceibias.n81 161.3
R7381 commonsourceibias.n84 commonsourceibias.n28 161.3
R7382 commonsourceibias.n86 commonsourceibias.n85 161.3
R7383 commonsourceibias.n87 commonsourceibias.n27 161.3
R7384 commonsourceibias.n89 commonsourceibias.n88 161.3
R7385 commonsourceibias.n90 commonsourceibias.n26 161.3
R7386 commonsourceibias.n93 commonsourceibias.n92 161.3
R7387 commonsourceibias.n94 commonsourceibias.n25 161.3
R7388 commonsourceibias.n96 commonsourceibias.n95 161.3
R7389 commonsourceibias.n98 commonsourceibias.n23 161.3
R7390 commonsourceibias.n100 commonsourceibias.n99 161.3
R7391 commonsourceibias.n101 commonsourceibias.n22 161.3
R7392 commonsourceibias.n103 commonsourceibias.n102 161.3
R7393 commonsourceibias.n104 commonsourceibias.n21 161.3
R7394 commonsourceibias.n107 commonsourceibias.n106 161.3
R7395 commonsourceibias.n108 commonsourceibias.n20 161.3
R7396 commonsourceibias.n110 commonsourceibias.n109 161.3
R7397 commonsourceibias.n112 commonsourceibias.n18 161.3
R7398 commonsourceibias.n114 commonsourceibias.n113 161.3
R7399 commonsourceibias.n115 commonsourceibias.n17 161.3
R7400 commonsourceibias.n117 commonsourceibias.n116 161.3
R7401 commonsourceibias.n118 commonsourceibias.n16 161.3
R7402 commonsourceibias.n121 commonsourceibias.n120 161.3
R7403 commonsourceibias.n122 commonsourceibias.n15 161.3
R7404 commonsourceibias.n124 commonsourceibias.n123 161.3
R7405 commonsourceibias.n126 commonsourceibias.n14 161.3
R7406 commonsourceibias.n167 commonsourceibias.n164 161.3
R7407 commonsourceibias.n169 commonsourceibias.n168 161.3
R7408 commonsourceibias.n170 commonsourceibias.n163 161.3
R7409 commonsourceibias.n173 commonsourceibias.n172 161.3
R7410 commonsourceibias.n174 commonsourceibias.n162 161.3
R7411 commonsourceibias.n176 commonsourceibias.n175 161.3
R7412 commonsourceibias.n178 commonsourceibias.n160 161.3
R7413 commonsourceibias.n180 commonsourceibias.n179 161.3
R7414 commonsourceibias.n181 commonsourceibias.n159 161.3
R7415 commonsourceibias.n183 commonsourceibias.n182 161.3
R7416 commonsourceibias.n184 commonsourceibias.n158 161.3
R7417 commonsourceibias.n187 commonsourceibias.n186 161.3
R7418 commonsourceibias.n188 commonsourceibias.n157 161.3
R7419 commonsourceibias.n190 commonsourceibias.n189 161.3
R7420 commonsourceibias.n192 commonsourceibias.n156 161.3
R7421 commonsourceibias.n194 commonsourceibias.n193 161.3
R7422 commonsourceibias.n196 commonsourceibias.n195 161.3
R7423 commonsourceibias.n197 commonsourceibias.n154 161.3
R7424 commonsourceibias.n199 commonsourceibias.n198 161.3
R7425 commonsourceibias.n201 commonsourceibias.n200 161.3
R7426 commonsourceibias.n202 commonsourceibias.n152 161.3
R7427 commonsourceibias.n204 commonsourceibias.n203 161.3
R7428 commonsourceibias.n206 commonsourceibias.n205 161.3
R7429 commonsourceibias.n208 commonsourceibias.n207 161.3
R7430 commonsourceibias.n209 commonsourceibias.n13 161.3
R7431 commonsourceibias.n211 commonsourceibias.n210 161.3
R7432 commonsourceibias.n212 commonsourceibias.n12 161.3
R7433 commonsourceibias.n215 commonsourceibias.n214 161.3
R7434 commonsourceibias.n216 commonsourceibias.n11 161.3
R7435 commonsourceibias.n218 commonsourceibias.n217 161.3
R7436 commonsourceibias.n220 commonsourceibias.n9 161.3
R7437 commonsourceibias.n222 commonsourceibias.n221 161.3
R7438 commonsourceibias.n223 commonsourceibias.n8 161.3
R7439 commonsourceibias.n225 commonsourceibias.n224 161.3
R7440 commonsourceibias.n226 commonsourceibias.n7 161.3
R7441 commonsourceibias.n229 commonsourceibias.n228 161.3
R7442 commonsourceibias.n230 commonsourceibias.n6 161.3
R7443 commonsourceibias.n232 commonsourceibias.n231 161.3
R7444 commonsourceibias.n234 commonsourceibias.n4 161.3
R7445 commonsourceibias.n236 commonsourceibias.n235 161.3
R7446 commonsourceibias.n237 commonsourceibias.n3 161.3
R7447 commonsourceibias.n239 commonsourceibias.n238 161.3
R7448 commonsourceibias.n240 commonsourceibias.n2 161.3
R7449 commonsourceibias.n243 commonsourceibias.n242 161.3
R7450 commonsourceibias.n244 commonsourceibias.n1 161.3
R7451 commonsourceibias.n246 commonsourceibias.n245 161.3
R7452 commonsourceibias.n248 commonsourceibias.n0 161.3
R7453 commonsourceibias.n730 commonsourceibias.n618 161.3
R7454 commonsourceibias.n728 commonsourceibias.n727 161.3
R7455 commonsourceibias.n726 commonsourceibias.n619 161.3
R7456 commonsourceibias.n725 commonsourceibias.n724 161.3
R7457 commonsourceibias.n722 commonsourceibias.n620 161.3
R7458 commonsourceibias.n721 commonsourceibias.n720 161.3
R7459 commonsourceibias.n719 commonsourceibias.n621 161.3
R7460 commonsourceibias.n718 commonsourceibias.n717 161.3
R7461 commonsourceibias.n715 commonsourceibias.n622 161.3
R7462 commonsourceibias.n713 commonsourceibias.n712 161.3
R7463 commonsourceibias.n711 commonsourceibias.n623 161.3
R7464 commonsourceibias.n710 commonsourceibias.n709 161.3
R7465 commonsourceibias.n707 commonsourceibias.n624 161.3
R7466 commonsourceibias.n706 commonsourceibias.n705 161.3
R7467 commonsourceibias.n704 commonsourceibias.n625 161.3
R7468 commonsourceibias.n703 commonsourceibias.n702 161.3
R7469 commonsourceibias.n700 commonsourceibias.n626 161.3
R7470 commonsourceibias.n698 commonsourceibias.n697 161.3
R7471 commonsourceibias.n696 commonsourceibias.n627 161.3
R7472 commonsourceibias.n695 commonsourceibias.n694 161.3
R7473 commonsourceibias.n692 commonsourceibias.n628 161.3
R7474 commonsourceibias.n691 commonsourceibias.n690 161.3
R7475 commonsourceibias.n689 commonsourceibias.n629 161.3
R7476 commonsourceibias.n688 commonsourceibias.n687 161.3
R7477 commonsourceibias.n685 commonsourceibias.n630 161.3
R7478 commonsourceibias.n683 commonsourceibias.n682 161.3
R7479 commonsourceibias.n681 commonsourceibias.n631 161.3
R7480 commonsourceibias.n680 commonsourceibias.n679 161.3
R7481 commonsourceibias.n677 commonsourceibias.n632 161.3
R7482 commonsourceibias.n676 commonsourceibias.n675 161.3
R7483 commonsourceibias.n674 commonsourceibias.n633 161.3
R7484 commonsourceibias.n673 commonsourceibias.n672 161.3
R7485 commonsourceibias.n670 commonsourceibias.n634 161.3
R7486 commonsourceibias.n668 commonsourceibias.n667 161.3
R7487 commonsourceibias.n666 commonsourceibias.n635 161.3
R7488 commonsourceibias.n665 commonsourceibias.n664 161.3
R7489 commonsourceibias.n662 commonsourceibias.n636 161.3
R7490 commonsourceibias.n661 commonsourceibias.n660 161.3
R7491 commonsourceibias.n659 commonsourceibias.n637 161.3
R7492 commonsourceibias.n658 commonsourceibias.n657 161.3
R7493 commonsourceibias.n655 commonsourceibias.n638 161.3
R7494 commonsourceibias.n653 commonsourceibias.n652 161.3
R7495 commonsourceibias.n651 commonsourceibias.n639 161.3
R7496 commonsourceibias.n650 commonsourceibias.n649 161.3
R7497 commonsourceibias.n647 commonsourceibias.n640 161.3
R7498 commonsourceibias.n646 commonsourceibias.n645 161.3
R7499 commonsourceibias.n644 commonsourceibias.n641 161.3
R7500 commonsourceibias.n500 commonsourceibias.n388 161.3
R7501 commonsourceibias.n498 commonsourceibias.n497 161.3
R7502 commonsourceibias.n496 commonsourceibias.n389 161.3
R7503 commonsourceibias.n495 commonsourceibias.n494 161.3
R7504 commonsourceibias.n492 commonsourceibias.n390 161.3
R7505 commonsourceibias.n491 commonsourceibias.n490 161.3
R7506 commonsourceibias.n489 commonsourceibias.n391 161.3
R7507 commonsourceibias.n488 commonsourceibias.n487 161.3
R7508 commonsourceibias.n485 commonsourceibias.n392 161.3
R7509 commonsourceibias.n483 commonsourceibias.n482 161.3
R7510 commonsourceibias.n481 commonsourceibias.n393 161.3
R7511 commonsourceibias.n480 commonsourceibias.n479 161.3
R7512 commonsourceibias.n477 commonsourceibias.n394 161.3
R7513 commonsourceibias.n476 commonsourceibias.n475 161.3
R7514 commonsourceibias.n474 commonsourceibias.n395 161.3
R7515 commonsourceibias.n473 commonsourceibias.n472 161.3
R7516 commonsourceibias.n470 commonsourceibias.n396 161.3
R7517 commonsourceibias.n468 commonsourceibias.n467 161.3
R7518 commonsourceibias.n466 commonsourceibias.n397 161.3
R7519 commonsourceibias.n465 commonsourceibias.n464 161.3
R7520 commonsourceibias.n462 commonsourceibias.n398 161.3
R7521 commonsourceibias.n461 commonsourceibias.n460 161.3
R7522 commonsourceibias.n459 commonsourceibias.n399 161.3
R7523 commonsourceibias.n458 commonsourceibias.n457 161.3
R7524 commonsourceibias.n455 commonsourceibias.n400 161.3
R7525 commonsourceibias.n453 commonsourceibias.n452 161.3
R7526 commonsourceibias.n451 commonsourceibias.n401 161.3
R7527 commonsourceibias.n450 commonsourceibias.n449 161.3
R7528 commonsourceibias.n447 commonsourceibias.n402 161.3
R7529 commonsourceibias.n446 commonsourceibias.n445 161.3
R7530 commonsourceibias.n444 commonsourceibias.n403 161.3
R7531 commonsourceibias.n443 commonsourceibias.n442 161.3
R7532 commonsourceibias.n440 commonsourceibias.n404 161.3
R7533 commonsourceibias.n438 commonsourceibias.n437 161.3
R7534 commonsourceibias.n436 commonsourceibias.n405 161.3
R7535 commonsourceibias.n435 commonsourceibias.n434 161.3
R7536 commonsourceibias.n432 commonsourceibias.n406 161.3
R7537 commonsourceibias.n431 commonsourceibias.n430 161.3
R7538 commonsourceibias.n429 commonsourceibias.n407 161.3
R7539 commonsourceibias.n428 commonsourceibias.n427 161.3
R7540 commonsourceibias.n425 commonsourceibias.n408 161.3
R7541 commonsourceibias.n423 commonsourceibias.n422 161.3
R7542 commonsourceibias.n421 commonsourceibias.n409 161.3
R7543 commonsourceibias.n420 commonsourceibias.n419 161.3
R7544 commonsourceibias.n417 commonsourceibias.n410 161.3
R7545 commonsourceibias.n416 commonsourceibias.n415 161.3
R7546 commonsourceibias.n414 commonsourceibias.n411 161.3
R7547 commonsourceibias.n570 commonsourceibias.n569 161.3
R7548 commonsourceibias.n568 commonsourceibias.n567 161.3
R7549 commonsourceibias.n566 commonsourceibias.n516 161.3
R7550 commonsourceibias.n565 commonsourceibias.n564 161.3
R7551 commonsourceibias.n563 commonsourceibias.n562 161.3
R7552 commonsourceibias.n561 commonsourceibias.n518 161.3
R7553 commonsourceibias.n560 commonsourceibias.n559 161.3
R7554 commonsourceibias.n558 commonsourceibias.n557 161.3
R7555 commonsourceibias.n556 commonsourceibias.n520 161.3
R7556 commonsourceibias.n554 commonsourceibias.n553 161.3
R7557 commonsourceibias.n552 commonsourceibias.n521 161.3
R7558 commonsourceibias.n551 commonsourceibias.n550 161.3
R7559 commonsourceibias.n548 commonsourceibias.n522 161.3
R7560 commonsourceibias.n547 commonsourceibias.n546 161.3
R7561 commonsourceibias.n545 commonsourceibias.n523 161.3
R7562 commonsourceibias.n544 commonsourceibias.n543 161.3
R7563 commonsourceibias.n541 commonsourceibias.n524 161.3
R7564 commonsourceibias.n539 commonsourceibias.n538 161.3
R7565 commonsourceibias.n537 commonsourceibias.n525 161.3
R7566 commonsourceibias.n536 commonsourceibias.n535 161.3
R7567 commonsourceibias.n533 commonsourceibias.n526 161.3
R7568 commonsourceibias.n532 commonsourceibias.n531 161.3
R7569 commonsourceibias.n530 commonsourceibias.n527 161.3
R7570 commonsourceibias.n615 commonsourceibias.n367 161.3
R7571 commonsourceibias.n613 commonsourceibias.n612 161.3
R7572 commonsourceibias.n611 commonsourceibias.n368 161.3
R7573 commonsourceibias.n610 commonsourceibias.n609 161.3
R7574 commonsourceibias.n607 commonsourceibias.n369 161.3
R7575 commonsourceibias.n606 commonsourceibias.n605 161.3
R7576 commonsourceibias.n604 commonsourceibias.n370 161.3
R7577 commonsourceibias.n603 commonsourceibias.n602 161.3
R7578 commonsourceibias.n600 commonsourceibias.n371 161.3
R7579 commonsourceibias.n598 commonsourceibias.n597 161.3
R7580 commonsourceibias.n596 commonsourceibias.n372 161.3
R7581 commonsourceibias.n595 commonsourceibias.n594 161.3
R7582 commonsourceibias.n592 commonsourceibias.n373 161.3
R7583 commonsourceibias.n591 commonsourceibias.n590 161.3
R7584 commonsourceibias.n589 commonsourceibias.n374 161.3
R7585 commonsourceibias.n588 commonsourceibias.n587 161.3
R7586 commonsourceibias.n585 commonsourceibias.n375 161.3
R7587 commonsourceibias.n583 commonsourceibias.n582 161.3
R7588 commonsourceibias.n581 commonsourceibias.n376 161.3
R7589 commonsourceibias.n580 commonsourceibias.n579 161.3
R7590 commonsourceibias.n577 commonsourceibias.n377 161.3
R7591 commonsourceibias.n576 commonsourceibias.n575 161.3
R7592 commonsourceibias.n574 commonsourceibias.n378 161.3
R7593 commonsourceibias.n573 commonsourceibias.n572 161.3
R7594 commonsourceibias.n141 commonsourceibias.n139 81.5057
R7595 commonsourceibias.n381 commonsourceibias.n379 81.5057
R7596 commonsourceibias.n141 commonsourceibias.n140 80.9324
R7597 commonsourceibias.n143 commonsourceibias.n142 80.9324
R7598 commonsourceibias.n145 commonsourceibias.n144 80.9324
R7599 commonsourceibias.n147 commonsourceibias.n146 80.9324
R7600 commonsourceibias.n138 commonsourceibias.n137 80.9324
R7601 commonsourceibias.n136 commonsourceibias.n135 80.9324
R7602 commonsourceibias.n134 commonsourceibias.n133 80.9324
R7603 commonsourceibias.n132 commonsourceibias.n131 80.9324
R7604 commonsourceibias.n130 commonsourceibias.n129 80.9324
R7605 commonsourceibias.n504 commonsourceibias.n503 80.9324
R7606 commonsourceibias.n506 commonsourceibias.n505 80.9324
R7607 commonsourceibias.n508 commonsourceibias.n507 80.9324
R7608 commonsourceibias.n510 commonsourceibias.n509 80.9324
R7609 commonsourceibias.n512 commonsourceibias.n511 80.9324
R7610 commonsourceibias.n387 commonsourceibias.n386 80.9324
R7611 commonsourceibias.n385 commonsourceibias.n384 80.9324
R7612 commonsourceibias.n383 commonsourceibias.n382 80.9324
R7613 commonsourceibias.n381 commonsourceibias.n380 80.9324
R7614 commonsourceibias.n365 commonsourceibias.n364 80.6037
R7615 commonsourceibias.n128 commonsourceibias.n127 80.6037
R7616 commonsourceibias.n250 commonsourceibias.n249 80.6037
R7617 commonsourceibias.n732 commonsourceibias.n731 80.6037
R7618 commonsourceibias.n502 commonsourceibias.n501 80.6037
R7619 commonsourceibias.n617 commonsourceibias.n616 80.6037
R7620 commonsourceibias.n322 commonsourceibias.n321 56.5617
R7621 commonsourceibias.n336 commonsourceibias.n335 56.5617
R7622 commonsourceibias.n85 commonsourceibias.n84 56.5617
R7623 commonsourceibias.n71 commonsourceibias.n70 56.5617
R7624 commonsourceibias.n207 commonsourceibias.n206 56.5617
R7625 commonsourceibias.n193 commonsourceibias.n192 56.5617
R7626 commonsourceibias.n687 commonsourceibias.n685 56.5617
R7627 commonsourceibias.n702 commonsourceibias.n700 56.5617
R7628 commonsourceibias.n457 commonsourceibias.n455 56.5617
R7629 commonsourceibias.n472 commonsourceibias.n470 56.5617
R7630 commonsourceibias.n572 commonsourceibias.n570 56.5617
R7631 commonsourceibias.n294 commonsourceibias.n293 56.5617
R7632 commonsourceibias.n308 commonsourceibias.n307 56.5617
R7633 commonsourceibias.n350 commonsourceibias.n349 56.5617
R7634 commonsourceibias.n113 commonsourceibias.n112 56.5617
R7635 commonsourceibias.n99 commonsourceibias.n98 56.5617
R7636 commonsourceibias.n57 commonsourceibias.n56 56.5617
R7637 commonsourceibias.n235 commonsourceibias.n234 56.5617
R7638 commonsourceibias.n221 commonsourceibias.n220 56.5617
R7639 commonsourceibias.n179 commonsourceibias.n178 56.5617
R7640 commonsourceibias.n657 commonsourceibias.n655 56.5617
R7641 commonsourceibias.n672 commonsourceibias.n670 56.5617
R7642 commonsourceibias.n717 commonsourceibias.n715 56.5617
R7643 commonsourceibias.n427 commonsourceibias.n425 56.5617
R7644 commonsourceibias.n442 commonsourceibias.n440 56.5617
R7645 commonsourceibias.n487 commonsourceibias.n485 56.5617
R7646 commonsourceibias.n602 commonsourceibias.n600 56.5617
R7647 commonsourceibias.n587 commonsourceibias.n585 56.5617
R7648 commonsourceibias.n543 commonsourceibias.n541 56.5617
R7649 commonsourceibias.n557 commonsourceibias.n556 56.5617
R7650 commonsourceibias.n285 commonsourceibias.n284 51.2335
R7651 commonsourceibias.n357 commonsourceibias.n252 51.2335
R7652 commonsourceibias.n120 commonsourceibias.n15 51.2335
R7653 commonsourceibias.n48 commonsourceibias.n47 51.2335
R7654 commonsourceibias.n242 commonsourceibias.n1 51.2335
R7655 commonsourceibias.n170 commonsourceibias.n169 51.2335
R7656 commonsourceibias.n647 commonsourceibias.n646 51.2335
R7657 commonsourceibias.n724 commonsourceibias.n619 51.2335
R7658 commonsourceibias.n417 commonsourceibias.n416 51.2335
R7659 commonsourceibias.n494 commonsourceibias.n389 51.2335
R7660 commonsourceibias.n609 commonsourceibias.n368 51.2335
R7661 commonsourceibias.n533 commonsourceibias.n532 51.2335
R7662 commonsourceibias.n364 commonsourceibias.n363 50.9056
R7663 commonsourceibias.n127 commonsourceibias.n126 50.9056
R7664 commonsourceibias.n249 commonsourceibias.n248 50.9056
R7665 commonsourceibias.n731 commonsourceibias.n730 50.9056
R7666 commonsourceibias.n501 commonsourceibias.n500 50.9056
R7667 commonsourceibias.n616 commonsourceibias.n615 50.9056
R7668 commonsourceibias.n299 commonsourceibias.n298 50.2647
R7669 commonsourceibias.n343 commonsourceibias.n257 50.2647
R7670 commonsourceibias.n106 commonsourceibias.n20 50.2647
R7671 commonsourceibias.n62 commonsourceibias.n61 50.2647
R7672 commonsourceibias.n228 commonsourceibias.n6 50.2647
R7673 commonsourceibias.n184 commonsourceibias.n183 50.2647
R7674 commonsourceibias.n662 commonsourceibias.n661 50.2647
R7675 commonsourceibias.n709 commonsourceibias.n623 50.2647
R7676 commonsourceibias.n432 commonsourceibias.n431 50.2647
R7677 commonsourceibias.n479 commonsourceibias.n393 50.2647
R7678 commonsourceibias.n594 commonsourceibias.n372 50.2647
R7679 commonsourceibias.n548 commonsourceibias.n547 50.2647
R7680 commonsourceibias.n281 commonsourceibias.n280 49.9027
R7681 commonsourceibias.n44 commonsourceibias.n43 49.9027
R7682 commonsourceibias.n166 commonsourceibias.n165 49.9027
R7683 commonsourceibias.n643 commonsourceibias.n642 49.9027
R7684 commonsourceibias.n413 commonsourceibias.n412 49.9027
R7685 commonsourceibias.n529 commonsourceibias.n528 49.9027
R7686 commonsourceibias.n313 commonsourceibias.n312 49.296
R7687 commonsourceibias.n329 commonsourceibias.n262 49.296
R7688 commonsourceibias.n92 commonsourceibias.n25 49.296
R7689 commonsourceibias.n76 commonsourceibias.n75 49.296
R7690 commonsourceibias.n214 commonsourceibias.n11 49.296
R7691 commonsourceibias.n198 commonsourceibias.n197 49.296
R7692 commonsourceibias.n677 commonsourceibias.n676 49.296
R7693 commonsourceibias.n694 commonsourceibias.n627 49.296
R7694 commonsourceibias.n447 commonsourceibias.n446 49.296
R7695 commonsourceibias.n464 commonsourceibias.n397 49.296
R7696 commonsourceibias.n579 commonsourceibias.n376 49.296
R7697 commonsourceibias.n562 commonsourceibias.n561 49.296
R7698 commonsourceibias.n315 commonsourceibias.n267 48.3272
R7699 commonsourceibias.n327 commonsourceibias.n326 48.3272
R7700 commonsourceibias.n90 commonsourceibias.n89 48.3272
R7701 commonsourceibias.n78 commonsourceibias.n30 48.3272
R7702 commonsourceibias.n212 commonsourceibias.n211 48.3272
R7703 commonsourceibias.n202 commonsourceibias.n201 48.3272
R7704 commonsourceibias.n679 commonsourceibias.n631 48.3272
R7705 commonsourceibias.n692 commonsourceibias.n691 48.3272
R7706 commonsourceibias.n449 commonsourceibias.n401 48.3272
R7707 commonsourceibias.n462 commonsourceibias.n461 48.3272
R7708 commonsourceibias.n577 commonsourceibias.n576 48.3272
R7709 commonsourceibias.n566 commonsourceibias.n565 48.3272
R7710 commonsourceibias.n301 commonsourceibias.n272 47.3584
R7711 commonsourceibias.n341 commonsourceibias.n340 47.3584
R7712 commonsourceibias.n104 commonsourceibias.n103 47.3584
R7713 commonsourceibias.n64 commonsourceibias.n35 47.3584
R7714 commonsourceibias.n226 commonsourceibias.n225 47.3584
R7715 commonsourceibias.n186 commonsourceibias.n157 47.3584
R7716 commonsourceibias.n664 commonsourceibias.n635 47.3584
R7717 commonsourceibias.n707 commonsourceibias.n706 47.3584
R7718 commonsourceibias.n434 commonsourceibias.n405 47.3584
R7719 commonsourceibias.n477 commonsourceibias.n476 47.3584
R7720 commonsourceibias.n592 commonsourceibias.n591 47.3584
R7721 commonsourceibias.n550 commonsourceibias.n521 47.3584
R7722 commonsourceibias.n287 commonsourceibias.n277 46.3896
R7723 commonsourceibias.n355 commonsourceibias.n354 46.3896
R7724 commonsourceibias.n118 commonsourceibias.n117 46.3896
R7725 commonsourceibias.n50 commonsourceibias.n40 46.3896
R7726 commonsourceibias.n240 commonsourceibias.n239 46.3896
R7727 commonsourceibias.n172 commonsourceibias.n162 46.3896
R7728 commonsourceibias.n649 commonsourceibias.n639 46.3896
R7729 commonsourceibias.n722 commonsourceibias.n721 46.3896
R7730 commonsourceibias.n419 commonsourceibias.n409 46.3896
R7731 commonsourceibias.n492 commonsourceibias.n491 46.3896
R7732 commonsourceibias.n607 commonsourceibias.n606 46.3896
R7733 commonsourceibias.n535 commonsourceibias.n525 46.3896
R7734 commonsourceibias.n282 commonsourceibias.n281 44.7059
R7735 commonsourceibias.n644 commonsourceibias.n643 44.7059
R7736 commonsourceibias.n414 commonsourceibias.n413 44.7059
R7737 commonsourceibias.n530 commonsourceibias.n529 44.7059
R7738 commonsourceibias.n45 commonsourceibias.n44 44.7059
R7739 commonsourceibias.n167 commonsourceibias.n166 44.7059
R7740 commonsourceibias.n291 commonsourceibias.n277 34.7644
R7741 commonsourceibias.n354 commonsourceibias.n254 34.7644
R7742 commonsourceibias.n117 commonsourceibias.n17 34.7644
R7743 commonsourceibias.n54 commonsourceibias.n40 34.7644
R7744 commonsourceibias.n239 commonsourceibias.n3 34.7644
R7745 commonsourceibias.n176 commonsourceibias.n162 34.7644
R7746 commonsourceibias.n653 commonsourceibias.n639 34.7644
R7747 commonsourceibias.n721 commonsourceibias.n621 34.7644
R7748 commonsourceibias.n423 commonsourceibias.n409 34.7644
R7749 commonsourceibias.n491 commonsourceibias.n391 34.7644
R7750 commonsourceibias.n606 commonsourceibias.n370 34.7644
R7751 commonsourceibias.n539 commonsourceibias.n525 34.7644
R7752 commonsourceibias.n305 commonsourceibias.n272 33.7956
R7753 commonsourceibias.n340 commonsourceibias.n259 33.7956
R7754 commonsourceibias.n103 commonsourceibias.n22 33.7956
R7755 commonsourceibias.n68 commonsourceibias.n35 33.7956
R7756 commonsourceibias.n225 commonsourceibias.n8 33.7956
R7757 commonsourceibias.n190 commonsourceibias.n157 33.7956
R7758 commonsourceibias.n668 commonsourceibias.n635 33.7956
R7759 commonsourceibias.n706 commonsourceibias.n625 33.7956
R7760 commonsourceibias.n438 commonsourceibias.n405 33.7956
R7761 commonsourceibias.n476 commonsourceibias.n395 33.7956
R7762 commonsourceibias.n591 commonsourceibias.n374 33.7956
R7763 commonsourceibias.n554 commonsourceibias.n521 33.7956
R7764 commonsourceibias.n319 commonsourceibias.n267 32.8269
R7765 commonsourceibias.n326 commonsourceibias.n264 32.8269
R7766 commonsourceibias.n89 commonsourceibias.n27 32.8269
R7767 commonsourceibias.n82 commonsourceibias.n30 32.8269
R7768 commonsourceibias.n211 commonsourceibias.n13 32.8269
R7769 commonsourceibias.n203 commonsourceibias.n202 32.8269
R7770 commonsourceibias.n683 commonsourceibias.n631 32.8269
R7771 commonsourceibias.n691 commonsourceibias.n629 32.8269
R7772 commonsourceibias.n453 commonsourceibias.n401 32.8269
R7773 commonsourceibias.n461 commonsourceibias.n399 32.8269
R7774 commonsourceibias.n576 commonsourceibias.n378 32.8269
R7775 commonsourceibias.n567 commonsourceibias.n566 32.8269
R7776 commonsourceibias.n312 commonsourceibias.n269 31.8581
R7777 commonsourceibias.n333 commonsourceibias.n262 31.8581
R7778 commonsourceibias.n96 commonsourceibias.n25 31.8581
R7779 commonsourceibias.n75 commonsourceibias.n32 31.8581
R7780 commonsourceibias.n218 commonsourceibias.n11 31.8581
R7781 commonsourceibias.n197 commonsourceibias.n196 31.8581
R7782 commonsourceibias.n676 commonsourceibias.n633 31.8581
R7783 commonsourceibias.n698 commonsourceibias.n627 31.8581
R7784 commonsourceibias.n446 commonsourceibias.n403 31.8581
R7785 commonsourceibias.n468 commonsourceibias.n397 31.8581
R7786 commonsourceibias.n583 commonsourceibias.n376 31.8581
R7787 commonsourceibias.n561 commonsourceibias.n560 31.8581
R7788 commonsourceibias.n298 commonsourceibias.n274 30.8893
R7789 commonsourceibias.n347 commonsourceibias.n257 30.8893
R7790 commonsourceibias.n110 commonsourceibias.n20 30.8893
R7791 commonsourceibias.n61 commonsourceibias.n37 30.8893
R7792 commonsourceibias.n232 commonsourceibias.n6 30.8893
R7793 commonsourceibias.n183 commonsourceibias.n159 30.8893
R7794 commonsourceibias.n661 commonsourceibias.n637 30.8893
R7795 commonsourceibias.n713 commonsourceibias.n623 30.8893
R7796 commonsourceibias.n431 commonsourceibias.n407 30.8893
R7797 commonsourceibias.n483 commonsourceibias.n393 30.8893
R7798 commonsourceibias.n598 commonsourceibias.n372 30.8893
R7799 commonsourceibias.n547 commonsourceibias.n523 30.8893
R7800 commonsourceibias.n284 commonsourceibias.n279 29.9206
R7801 commonsourceibias.n361 commonsourceibias.n252 29.9206
R7802 commonsourceibias.n124 commonsourceibias.n15 29.9206
R7803 commonsourceibias.n47 commonsourceibias.n42 29.9206
R7804 commonsourceibias.n246 commonsourceibias.n1 29.9206
R7805 commonsourceibias.n169 commonsourceibias.n164 29.9206
R7806 commonsourceibias.n646 commonsourceibias.n641 29.9206
R7807 commonsourceibias.n728 commonsourceibias.n619 29.9206
R7808 commonsourceibias.n416 commonsourceibias.n411 29.9206
R7809 commonsourceibias.n498 commonsourceibias.n389 29.9206
R7810 commonsourceibias.n613 commonsourceibias.n368 29.9206
R7811 commonsourceibias.n532 commonsourceibias.n527 29.9206
R7812 commonsourceibias.n363 commonsourceibias.n362 21.8872
R7813 commonsourceibias.n126 commonsourceibias.n125 21.8872
R7814 commonsourceibias.n248 commonsourceibias.n247 21.8872
R7815 commonsourceibias.n730 commonsourceibias.n729 21.8872
R7816 commonsourceibias.n500 commonsourceibias.n499 21.8872
R7817 commonsourceibias.n615 commonsourceibias.n614 21.8872
R7818 commonsourceibias.n294 commonsourceibias.n276 21.3954
R7819 commonsourceibias.n349 commonsourceibias.n348 21.3954
R7820 commonsourceibias.n112 commonsourceibias.n111 21.3954
R7821 commonsourceibias.n57 commonsourceibias.n39 21.3954
R7822 commonsourceibias.n234 commonsourceibias.n233 21.3954
R7823 commonsourceibias.n179 commonsourceibias.n161 21.3954
R7824 commonsourceibias.n657 commonsourceibias.n656 21.3954
R7825 commonsourceibias.n715 commonsourceibias.n714 21.3954
R7826 commonsourceibias.n427 commonsourceibias.n426 21.3954
R7827 commonsourceibias.n485 commonsourceibias.n484 21.3954
R7828 commonsourceibias.n600 commonsourceibias.n599 21.3954
R7829 commonsourceibias.n543 commonsourceibias.n542 21.3954
R7830 commonsourceibias.n308 commonsourceibias.n271 20.9036
R7831 commonsourceibias.n335 commonsourceibias.n334 20.9036
R7832 commonsourceibias.n98 commonsourceibias.n97 20.9036
R7833 commonsourceibias.n71 commonsourceibias.n34 20.9036
R7834 commonsourceibias.n220 commonsourceibias.n219 20.9036
R7835 commonsourceibias.n193 commonsourceibias.n155 20.9036
R7836 commonsourceibias.n672 commonsourceibias.n671 20.9036
R7837 commonsourceibias.n700 commonsourceibias.n699 20.9036
R7838 commonsourceibias.n442 commonsourceibias.n441 20.9036
R7839 commonsourceibias.n470 commonsourceibias.n469 20.9036
R7840 commonsourceibias.n585 commonsourceibias.n584 20.9036
R7841 commonsourceibias.n557 commonsourceibias.n519 20.9036
R7842 commonsourceibias.n321 commonsourceibias.n320 20.4117
R7843 commonsourceibias.n322 commonsourceibias.n266 20.4117
R7844 commonsourceibias.n85 commonsourceibias.n29 20.4117
R7845 commonsourceibias.n84 commonsourceibias.n83 20.4117
R7846 commonsourceibias.n207 commonsourceibias.n150 20.4117
R7847 commonsourceibias.n206 commonsourceibias.n151 20.4117
R7848 commonsourceibias.n685 commonsourceibias.n684 20.4117
R7849 commonsourceibias.n687 commonsourceibias.n686 20.4117
R7850 commonsourceibias.n455 commonsourceibias.n454 20.4117
R7851 commonsourceibias.n457 commonsourceibias.n456 20.4117
R7852 commonsourceibias.n572 commonsourceibias.n571 20.4117
R7853 commonsourceibias.n570 commonsourceibias.n515 20.4117
R7854 commonsourceibias.n307 commonsourceibias.n306 19.9199
R7855 commonsourceibias.n336 commonsourceibias.n261 19.9199
R7856 commonsourceibias.n99 commonsourceibias.n24 19.9199
R7857 commonsourceibias.n70 commonsourceibias.n69 19.9199
R7858 commonsourceibias.n221 commonsourceibias.n10 19.9199
R7859 commonsourceibias.n192 commonsourceibias.n191 19.9199
R7860 commonsourceibias.n670 commonsourceibias.n669 19.9199
R7861 commonsourceibias.n702 commonsourceibias.n701 19.9199
R7862 commonsourceibias.n440 commonsourceibias.n439 19.9199
R7863 commonsourceibias.n472 commonsourceibias.n471 19.9199
R7864 commonsourceibias.n587 commonsourceibias.n586 19.9199
R7865 commonsourceibias.n556 commonsourceibias.n555 19.9199
R7866 commonsourceibias.n293 commonsourceibias.n292 19.4281
R7867 commonsourceibias.n350 commonsourceibias.n256 19.4281
R7868 commonsourceibias.n113 commonsourceibias.n19 19.4281
R7869 commonsourceibias.n56 commonsourceibias.n55 19.4281
R7870 commonsourceibias.n235 commonsourceibias.n5 19.4281
R7871 commonsourceibias.n178 commonsourceibias.n177 19.4281
R7872 commonsourceibias.n655 commonsourceibias.n654 19.4281
R7873 commonsourceibias.n717 commonsourceibias.n716 19.4281
R7874 commonsourceibias.n425 commonsourceibias.n424 19.4281
R7875 commonsourceibias.n487 commonsourceibias.n486 19.4281
R7876 commonsourceibias.n602 commonsourceibias.n601 19.4281
R7877 commonsourceibias.n541 commonsourceibias.n540 19.4281
R7878 commonsourceibias.n286 commonsourceibias.n285 13.526
R7879 commonsourceibias.n357 commonsourceibias.n356 13.526
R7880 commonsourceibias.n120 commonsourceibias.n119 13.526
R7881 commonsourceibias.n49 commonsourceibias.n48 13.526
R7882 commonsourceibias.n242 commonsourceibias.n241 13.526
R7883 commonsourceibias.n171 commonsourceibias.n170 13.526
R7884 commonsourceibias.n648 commonsourceibias.n647 13.526
R7885 commonsourceibias.n724 commonsourceibias.n723 13.526
R7886 commonsourceibias.n418 commonsourceibias.n417 13.526
R7887 commonsourceibias.n494 commonsourceibias.n493 13.526
R7888 commonsourceibias.n609 commonsourceibias.n608 13.526
R7889 commonsourceibias.n534 commonsourceibias.n533 13.526
R7890 commonsourceibias.n130 commonsourceibias.n128 13.2322
R7891 commonsourceibias.n504 commonsourceibias.n502 13.2322
R7892 commonsourceibias.n300 commonsourceibias.n299 13.0342
R7893 commonsourceibias.n343 commonsourceibias.n342 13.0342
R7894 commonsourceibias.n106 commonsourceibias.n105 13.0342
R7895 commonsourceibias.n63 commonsourceibias.n62 13.0342
R7896 commonsourceibias.n228 commonsourceibias.n227 13.0342
R7897 commonsourceibias.n185 commonsourceibias.n184 13.0342
R7898 commonsourceibias.n663 commonsourceibias.n662 13.0342
R7899 commonsourceibias.n709 commonsourceibias.n708 13.0342
R7900 commonsourceibias.n433 commonsourceibias.n432 13.0342
R7901 commonsourceibias.n479 commonsourceibias.n478 13.0342
R7902 commonsourceibias.n594 commonsourceibias.n593 13.0342
R7903 commonsourceibias.n549 commonsourceibias.n548 13.0342
R7904 commonsourceibias.n314 commonsourceibias.n313 12.5423
R7905 commonsourceibias.n329 commonsourceibias.n328 12.5423
R7906 commonsourceibias.n92 commonsourceibias.n91 12.5423
R7907 commonsourceibias.n77 commonsourceibias.n76 12.5423
R7908 commonsourceibias.n214 commonsourceibias.n213 12.5423
R7909 commonsourceibias.n198 commonsourceibias.n153 12.5423
R7910 commonsourceibias.n678 commonsourceibias.n677 12.5423
R7911 commonsourceibias.n694 commonsourceibias.n693 12.5423
R7912 commonsourceibias.n448 commonsourceibias.n447 12.5423
R7913 commonsourceibias.n464 commonsourceibias.n463 12.5423
R7914 commonsourceibias.n579 commonsourceibias.n578 12.5423
R7915 commonsourceibias.n562 commonsourceibias.n517 12.5423
R7916 commonsourceibias.n315 commonsourceibias.n314 12.0505
R7917 commonsourceibias.n328 commonsourceibias.n327 12.0505
R7918 commonsourceibias.n91 commonsourceibias.n90 12.0505
R7919 commonsourceibias.n78 commonsourceibias.n77 12.0505
R7920 commonsourceibias.n213 commonsourceibias.n212 12.0505
R7921 commonsourceibias.n201 commonsourceibias.n153 12.0505
R7922 commonsourceibias.n679 commonsourceibias.n678 12.0505
R7923 commonsourceibias.n693 commonsourceibias.n692 12.0505
R7924 commonsourceibias.n449 commonsourceibias.n448 12.0505
R7925 commonsourceibias.n463 commonsourceibias.n462 12.0505
R7926 commonsourceibias.n578 commonsourceibias.n577 12.0505
R7927 commonsourceibias.n565 commonsourceibias.n517 12.0505
R7928 commonsourceibias.n734 commonsourceibias.n366 11.9876
R7929 commonsourceibias.n301 commonsourceibias.n300 11.5587
R7930 commonsourceibias.n342 commonsourceibias.n341 11.5587
R7931 commonsourceibias.n105 commonsourceibias.n104 11.5587
R7932 commonsourceibias.n64 commonsourceibias.n63 11.5587
R7933 commonsourceibias.n227 commonsourceibias.n226 11.5587
R7934 commonsourceibias.n186 commonsourceibias.n185 11.5587
R7935 commonsourceibias.n664 commonsourceibias.n663 11.5587
R7936 commonsourceibias.n708 commonsourceibias.n707 11.5587
R7937 commonsourceibias.n434 commonsourceibias.n433 11.5587
R7938 commonsourceibias.n478 commonsourceibias.n477 11.5587
R7939 commonsourceibias.n593 commonsourceibias.n592 11.5587
R7940 commonsourceibias.n550 commonsourceibias.n549 11.5587
R7941 commonsourceibias.n287 commonsourceibias.n286 11.0668
R7942 commonsourceibias.n356 commonsourceibias.n355 11.0668
R7943 commonsourceibias.n119 commonsourceibias.n118 11.0668
R7944 commonsourceibias.n50 commonsourceibias.n49 11.0668
R7945 commonsourceibias.n241 commonsourceibias.n240 11.0668
R7946 commonsourceibias.n172 commonsourceibias.n171 11.0668
R7947 commonsourceibias.n649 commonsourceibias.n648 11.0668
R7948 commonsourceibias.n723 commonsourceibias.n722 11.0668
R7949 commonsourceibias.n419 commonsourceibias.n418 11.0668
R7950 commonsourceibias.n493 commonsourceibias.n492 11.0668
R7951 commonsourceibias.n608 commonsourceibias.n607 11.0668
R7952 commonsourceibias.n535 commonsourceibias.n534 11.0668
R7953 commonsourceibias.n734 commonsourceibias.n733 10.3347
R7954 commonsourceibias.n149 commonsourceibias.n148 9.50363
R7955 commonsourceibias.n514 commonsourceibias.n513 9.50363
R7956 commonsourceibias.n366 commonsourceibias.n250 8.75852
R7957 commonsourceibias.n733 commonsourceibias.n617 8.75852
R7958 commonsourceibias.n292 commonsourceibias.n291 5.16479
R7959 commonsourceibias.n256 commonsourceibias.n254 5.16479
R7960 commonsourceibias.n19 commonsourceibias.n17 5.16479
R7961 commonsourceibias.n55 commonsourceibias.n54 5.16479
R7962 commonsourceibias.n5 commonsourceibias.n3 5.16479
R7963 commonsourceibias.n177 commonsourceibias.n176 5.16479
R7964 commonsourceibias.n654 commonsourceibias.n653 5.16479
R7965 commonsourceibias.n716 commonsourceibias.n621 5.16479
R7966 commonsourceibias.n424 commonsourceibias.n423 5.16479
R7967 commonsourceibias.n486 commonsourceibias.n391 5.16479
R7968 commonsourceibias.n601 commonsourceibias.n370 5.16479
R7969 commonsourceibias.n540 commonsourceibias.n539 5.16479
R7970 commonsourceibias.n366 commonsourceibias.n365 5.03125
R7971 commonsourceibias.n733 commonsourceibias.n732 5.03125
R7972 commonsourceibias.n306 commonsourceibias.n305 4.67295
R7973 commonsourceibias.n261 commonsourceibias.n259 4.67295
R7974 commonsourceibias.n24 commonsourceibias.n22 4.67295
R7975 commonsourceibias.n69 commonsourceibias.n68 4.67295
R7976 commonsourceibias.n10 commonsourceibias.n8 4.67295
R7977 commonsourceibias.n191 commonsourceibias.n190 4.67295
R7978 commonsourceibias.n669 commonsourceibias.n668 4.67295
R7979 commonsourceibias.n701 commonsourceibias.n625 4.67295
R7980 commonsourceibias.n439 commonsourceibias.n438 4.67295
R7981 commonsourceibias.n471 commonsourceibias.n395 4.67295
R7982 commonsourceibias.n586 commonsourceibias.n374 4.67295
R7983 commonsourceibias.n555 commonsourceibias.n554 4.67295
R7984 commonsourceibias commonsourceibias.n734 4.20978
R7985 commonsourceibias.n320 commonsourceibias.n319 4.18111
R7986 commonsourceibias.n266 commonsourceibias.n264 4.18111
R7987 commonsourceibias.n29 commonsourceibias.n27 4.18111
R7988 commonsourceibias.n83 commonsourceibias.n82 4.18111
R7989 commonsourceibias.n150 commonsourceibias.n13 4.18111
R7990 commonsourceibias.n203 commonsourceibias.n151 4.18111
R7991 commonsourceibias.n684 commonsourceibias.n683 4.18111
R7992 commonsourceibias.n686 commonsourceibias.n629 4.18111
R7993 commonsourceibias.n454 commonsourceibias.n453 4.18111
R7994 commonsourceibias.n456 commonsourceibias.n399 4.18111
R7995 commonsourceibias.n571 commonsourceibias.n378 4.18111
R7996 commonsourceibias.n567 commonsourceibias.n515 4.18111
R7997 commonsourceibias.n271 commonsourceibias.n269 3.68928
R7998 commonsourceibias.n334 commonsourceibias.n333 3.68928
R7999 commonsourceibias.n97 commonsourceibias.n96 3.68928
R8000 commonsourceibias.n34 commonsourceibias.n32 3.68928
R8001 commonsourceibias.n219 commonsourceibias.n218 3.68928
R8002 commonsourceibias.n196 commonsourceibias.n155 3.68928
R8003 commonsourceibias.n671 commonsourceibias.n633 3.68928
R8004 commonsourceibias.n699 commonsourceibias.n698 3.68928
R8005 commonsourceibias.n441 commonsourceibias.n403 3.68928
R8006 commonsourceibias.n469 commonsourceibias.n468 3.68928
R8007 commonsourceibias.n584 commonsourceibias.n583 3.68928
R8008 commonsourceibias.n560 commonsourceibias.n519 3.68928
R8009 commonsourceibias.n276 commonsourceibias.n274 3.19744
R8010 commonsourceibias.n348 commonsourceibias.n347 3.19744
R8011 commonsourceibias.n111 commonsourceibias.n110 3.19744
R8012 commonsourceibias.n39 commonsourceibias.n37 3.19744
R8013 commonsourceibias.n233 commonsourceibias.n232 3.19744
R8014 commonsourceibias.n161 commonsourceibias.n159 3.19744
R8015 commonsourceibias.n656 commonsourceibias.n637 3.19744
R8016 commonsourceibias.n714 commonsourceibias.n713 3.19744
R8017 commonsourceibias.n426 commonsourceibias.n407 3.19744
R8018 commonsourceibias.n484 commonsourceibias.n483 3.19744
R8019 commonsourceibias.n599 commonsourceibias.n598 3.19744
R8020 commonsourceibias.n542 commonsourceibias.n523 3.19744
R8021 commonsourceibias.n139 commonsourceibias.t65 2.82907
R8022 commonsourceibias.n139 commonsourceibias.t33 2.82907
R8023 commonsourceibias.n140 commonsourceibias.t61 2.82907
R8024 commonsourceibias.n140 commonsourceibias.t53 2.82907
R8025 commonsourceibias.n142 commonsourceibias.t69 2.82907
R8026 commonsourceibias.n142 commonsourceibias.t19 2.82907
R8027 commonsourceibias.n144 commonsourceibias.t9 2.82907
R8028 commonsourceibias.n144 commonsourceibias.t29 2.82907
R8029 commonsourceibias.n146 commonsourceibias.t77 2.82907
R8030 commonsourceibias.n146 commonsourceibias.t39 2.82907
R8031 commonsourceibias.n137 commonsourceibias.t15 2.82907
R8032 commonsourceibias.n137 commonsourceibias.t55 2.82907
R8033 commonsourceibias.n135 commonsourceibias.t37 2.82907
R8034 commonsourceibias.n135 commonsourceibias.t23 2.82907
R8035 commonsourceibias.n133 commonsourceibias.t47 2.82907
R8036 commonsourceibias.n133 commonsourceibias.t17 2.82907
R8037 commonsourceibias.n131 commonsourceibias.t43 2.82907
R8038 commonsourceibias.n131 commonsourceibias.t11 2.82907
R8039 commonsourceibias.n129 commonsourceibias.t13 2.82907
R8040 commonsourceibias.n129 commonsourceibias.t67 2.82907
R8041 commonsourceibias.n503 commonsourceibias.t49 2.82907
R8042 commonsourceibias.n503 commonsourceibias.t59 2.82907
R8043 commonsourceibias.n505 commonsourceibias.t57 2.82907
R8044 commonsourceibias.n505 commonsourceibias.t31 2.82907
R8045 commonsourceibias.n507 commonsourceibias.t71 2.82907
R8046 commonsourceibias.n507 commonsourceibias.t25 2.82907
R8047 commonsourceibias.n509 commonsourceibias.t79 2.82907
R8048 commonsourceibias.n509 commonsourceibias.t51 2.82907
R8049 commonsourceibias.n511 commonsourceibias.t3 2.82907
R8050 commonsourceibias.n511 commonsourceibias.t63 2.82907
R8051 commonsourceibias.n386 commonsourceibias.t5 2.82907
R8052 commonsourceibias.n386 commonsourceibias.t75 2.82907
R8053 commonsourceibias.n384 commonsourceibias.t73 2.82907
R8054 commonsourceibias.n384 commonsourceibias.t41 2.82907
R8055 commonsourceibias.n382 commonsourceibias.t35 2.82907
R8056 commonsourceibias.n382 commonsourceibias.t27 2.82907
R8057 commonsourceibias.n380 commonsourceibias.t45 2.82907
R8058 commonsourceibias.n380 commonsourceibias.t7 2.82907
R8059 commonsourceibias.n379 commonsourceibias.t1 2.82907
R8060 commonsourceibias.n379 commonsourceibias.t21 2.82907
R8061 commonsourceibias.n280 commonsourceibias.n279 2.7056
R8062 commonsourceibias.n362 commonsourceibias.n361 2.7056
R8063 commonsourceibias.n125 commonsourceibias.n124 2.7056
R8064 commonsourceibias.n43 commonsourceibias.n42 2.7056
R8065 commonsourceibias.n247 commonsourceibias.n246 2.7056
R8066 commonsourceibias.n165 commonsourceibias.n164 2.7056
R8067 commonsourceibias.n642 commonsourceibias.n641 2.7056
R8068 commonsourceibias.n729 commonsourceibias.n728 2.7056
R8069 commonsourceibias.n412 commonsourceibias.n411 2.7056
R8070 commonsourceibias.n499 commonsourceibias.n498 2.7056
R8071 commonsourceibias.n614 commonsourceibias.n613 2.7056
R8072 commonsourceibias.n528 commonsourceibias.n527 2.7056
R8073 commonsourceibias.n132 commonsourceibias.n130 0.573776
R8074 commonsourceibias.n134 commonsourceibias.n132 0.573776
R8075 commonsourceibias.n136 commonsourceibias.n134 0.573776
R8076 commonsourceibias.n138 commonsourceibias.n136 0.573776
R8077 commonsourceibias.n147 commonsourceibias.n145 0.573776
R8078 commonsourceibias.n145 commonsourceibias.n143 0.573776
R8079 commonsourceibias.n143 commonsourceibias.n141 0.573776
R8080 commonsourceibias.n383 commonsourceibias.n381 0.573776
R8081 commonsourceibias.n385 commonsourceibias.n383 0.573776
R8082 commonsourceibias.n387 commonsourceibias.n385 0.573776
R8083 commonsourceibias.n512 commonsourceibias.n510 0.573776
R8084 commonsourceibias.n510 commonsourceibias.n508 0.573776
R8085 commonsourceibias.n508 commonsourceibias.n506 0.573776
R8086 commonsourceibias.n506 commonsourceibias.n504 0.573776
R8087 commonsourceibias.n148 commonsourceibias.n138 0.287138
R8088 commonsourceibias.n148 commonsourceibias.n147 0.287138
R8089 commonsourceibias.n513 commonsourceibias.n387 0.287138
R8090 commonsourceibias.n513 commonsourceibias.n512 0.287138
R8091 commonsourceibias.n365 commonsourceibias.n251 0.285035
R8092 commonsourceibias.n128 commonsourceibias.n14 0.285035
R8093 commonsourceibias.n250 commonsourceibias.n0 0.285035
R8094 commonsourceibias.n732 commonsourceibias.n618 0.285035
R8095 commonsourceibias.n502 commonsourceibias.n388 0.285035
R8096 commonsourceibias.n617 commonsourceibias.n367 0.285035
R8097 commonsourceibias.n360 commonsourceibias.n251 0.189894
R8098 commonsourceibias.n360 commonsourceibias.n359 0.189894
R8099 commonsourceibias.n359 commonsourceibias.n358 0.189894
R8100 commonsourceibias.n358 commonsourceibias.n253 0.189894
R8101 commonsourceibias.n353 commonsourceibias.n253 0.189894
R8102 commonsourceibias.n353 commonsourceibias.n352 0.189894
R8103 commonsourceibias.n352 commonsourceibias.n351 0.189894
R8104 commonsourceibias.n351 commonsourceibias.n255 0.189894
R8105 commonsourceibias.n346 commonsourceibias.n255 0.189894
R8106 commonsourceibias.n346 commonsourceibias.n345 0.189894
R8107 commonsourceibias.n345 commonsourceibias.n344 0.189894
R8108 commonsourceibias.n344 commonsourceibias.n258 0.189894
R8109 commonsourceibias.n339 commonsourceibias.n258 0.189894
R8110 commonsourceibias.n339 commonsourceibias.n338 0.189894
R8111 commonsourceibias.n338 commonsourceibias.n337 0.189894
R8112 commonsourceibias.n337 commonsourceibias.n260 0.189894
R8113 commonsourceibias.n332 commonsourceibias.n260 0.189894
R8114 commonsourceibias.n332 commonsourceibias.n331 0.189894
R8115 commonsourceibias.n331 commonsourceibias.n330 0.189894
R8116 commonsourceibias.n330 commonsourceibias.n263 0.189894
R8117 commonsourceibias.n325 commonsourceibias.n263 0.189894
R8118 commonsourceibias.n325 commonsourceibias.n324 0.189894
R8119 commonsourceibias.n324 commonsourceibias.n323 0.189894
R8120 commonsourceibias.n323 commonsourceibias.n265 0.189894
R8121 commonsourceibias.n318 commonsourceibias.n265 0.189894
R8122 commonsourceibias.n318 commonsourceibias.n317 0.189894
R8123 commonsourceibias.n317 commonsourceibias.n316 0.189894
R8124 commonsourceibias.n316 commonsourceibias.n268 0.189894
R8125 commonsourceibias.n311 commonsourceibias.n268 0.189894
R8126 commonsourceibias.n311 commonsourceibias.n310 0.189894
R8127 commonsourceibias.n310 commonsourceibias.n309 0.189894
R8128 commonsourceibias.n309 commonsourceibias.n270 0.189894
R8129 commonsourceibias.n304 commonsourceibias.n270 0.189894
R8130 commonsourceibias.n304 commonsourceibias.n303 0.189894
R8131 commonsourceibias.n303 commonsourceibias.n302 0.189894
R8132 commonsourceibias.n302 commonsourceibias.n273 0.189894
R8133 commonsourceibias.n297 commonsourceibias.n273 0.189894
R8134 commonsourceibias.n297 commonsourceibias.n296 0.189894
R8135 commonsourceibias.n296 commonsourceibias.n295 0.189894
R8136 commonsourceibias.n295 commonsourceibias.n275 0.189894
R8137 commonsourceibias.n290 commonsourceibias.n275 0.189894
R8138 commonsourceibias.n290 commonsourceibias.n289 0.189894
R8139 commonsourceibias.n289 commonsourceibias.n288 0.189894
R8140 commonsourceibias.n288 commonsourceibias.n278 0.189894
R8141 commonsourceibias.n283 commonsourceibias.n278 0.189894
R8142 commonsourceibias.n283 commonsourceibias.n282 0.189894
R8143 commonsourceibias.n123 commonsourceibias.n14 0.189894
R8144 commonsourceibias.n123 commonsourceibias.n122 0.189894
R8145 commonsourceibias.n122 commonsourceibias.n121 0.189894
R8146 commonsourceibias.n121 commonsourceibias.n16 0.189894
R8147 commonsourceibias.n116 commonsourceibias.n16 0.189894
R8148 commonsourceibias.n116 commonsourceibias.n115 0.189894
R8149 commonsourceibias.n115 commonsourceibias.n114 0.189894
R8150 commonsourceibias.n114 commonsourceibias.n18 0.189894
R8151 commonsourceibias.n109 commonsourceibias.n18 0.189894
R8152 commonsourceibias.n109 commonsourceibias.n108 0.189894
R8153 commonsourceibias.n108 commonsourceibias.n107 0.189894
R8154 commonsourceibias.n107 commonsourceibias.n21 0.189894
R8155 commonsourceibias.n102 commonsourceibias.n21 0.189894
R8156 commonsourceibias.n102 commonsourceibias.n101 0.189894
R8157 commonsourceibias.n101 commonsourceibias.n100 0.189894
R8158 commonsourceibias.n100 commonsourceibias.n23 0.189894
R8159 commonsourceibias.n95 commonsourceibias.n23 0.189894
R8160 commonsourceibias.n95 commonsourceibias.n94 0.189894
R8161 commonsourceibias.n94 commonsourceibias.n93 0.189894
R8162 commonsourceibias.n93 commonsourceibias.n26 0.189894
R8163 commonsourceibias.n88 commonsourceibias.n26 0.189894
R8164 commonsourceibias.n88 commonsourceibias.n87 0.189894
R8165 commonsourceibias.n87 commonsourceibias.n86 0.189894
R8166 commonsourceibias.n86 commonsourceibias.n28 0.189894
R8167 commonsourceibias.n81 commonsourceibias.n28 0.189894
R8168 commonsourceibias.n81 commonsourceibias.n80 0.189894
R8169 commonsourceibias.n80 commonsourceibias.n79 0.189894
R8170 commonsourceibias.n79 commonsourceibias.n31 0.189894
R8171 commonsourceibias.n74 commonsourceibias.n31 0.189894
R8172 commonsourceibias.n74 commonsourceibias.n73 0.189894
R8173 commonsourceibias.n73 commonsourceibias.n72 0.189894
R8174 commonsourceibias.n72 commonsourceibias.n33 0.189894
R8175 commonsourceibias.n67 commonsourceibias.n33 0.189894
R8176 commonsourceibias.n67 commonsourceibias.n66 0.189894
R8177 commonsourceibias.n66 commonsourceibias.n65 0.189894
R8178 commonsourceibias.n65 commonsourceibias.n36 0.189894
R8179 commonsourceibias.n60 commonsourceibias.n36 0.189894
R8180 commonsourceibias.n60 commonsourceibias.n59 0.189894
R8181 commonsourceibias.n59 commonsourceibias.n58 0.189894
R8182 commonsourceibias.n58 commonsourceibias.n38 0.189894
R8183 commonsourceibias.n53 commonsourceibias.n38 0.189894
R8184 commonsourceibias.n53 commonsourceibias.n52 0.189894
R8185 commonsourceibias.n52 commonsourceibias.n51 0.189894
R8186 commonsourceibias.n51 commonsourceibias.n41 0.189894
R8187 commonsourceibias.n46 commonsourceibias.n41 0.189894
R8188 commonsourceibias.n46 commonsourceibias.n45 0.189894
R8189 commonsourceibias.n205 commonsourceibias.n204 0.189894
R8190 commonsourceibias.n204 commonsourceibias.n152 0.189894
R8191 commonsourceibias.n200 commonsourceibias.n152 0.189894
R8192 commonsourceibias.n200 commonsourceibias.n199 0.189894
R8193 commonsourceibias.n199 commonsourceibias.n154 0.189894
R8194 commonsourceibias.n195 commonsourceibias.n154 0.189894
R8195 commonsourceibias.n195 commonsourceibias.n194 0.189894
R8196 commonsourceibias.n194 commonsourceibias.n156 0.189894
R8197 commonsourceibias.n189 commonsourceibias.n156 0.189894
R8198 commonsourceibias.n189 commonsourceibias.n188 0.189894
R8199 commonsourceibias.n188 commonsourceibias.n187 0.189894
R8200 commonsourceibias.n187 commonsourceibias.n158 0.189894
R8201 commonsourceibias.n182 commonsourceibias.n158 0.189894
R8202 commonsourceibias.n182 commonsourceibias.n181 0.189894
R8203 commonsourceibias.n181 commonsourceibias.n180 0.189894
R8204 commonsourceibias.n180 commonsourceibias.n160 0.189894
R8205 commonsourceibias.n175 commonsourceibias.n160 0.189894
R8206 commonsourceibias.n175 commonsourceibias.n174 0.189894
R8207 commonsourceibias.n174 commonsourceibias.n173 0.189894
R8208 commonsourceibias.n173 commonsourceibias.n163 0.189894
R8209 commonsourceibias.n168 commonsourceibias.n163 0.189894
R8210 commonsourceibias.n168 commonsourceibias.n167 0.189894
R8211 commonsourceibias.n245 commonsourceibias.n0 0.189894
R8212 commonsourceibias.n245 commonsourceibias.n244 0.189894
R8213 commonsourceibias.n244 commonsourceibias.n243 0.189894
R8214 commonsourceibias.n243 commonsourceibias.n2 0.189894
R8215 commonsourceibias.n238 commonsourceibias.n2 0.189894
R8216 commonsourceibias.n238 commonsourceibias.n237 0.189894
R8217 commonsourceibias.n237 commonsourceibias.n236 0.189894
R8218 commonsourceibias.n236 commonsourceibias.n4 0.189894
R8219 commonsourceibias.n231 commonsourceibias.n4 0.189894
R8220 commonsourceibias.n231 commonsourceibias.n230 0.189894
R8221 commonsourceibias.n230 commonsourceibias.n229 0.189894
R8222 commonsourceibias.n229 commonsourceibias.n7 0.189894
R8223 commonsourceibias.n224 commonsourceibias.n7 0.189894
R8224 commonsourceibias.n224 commonsourceibias.n223 0.189894
R8225 commonsourceibias.n223 commonsourceibias.n222 0.189894
R8226 commonsourceibias.n222 commonsourceibias.n9 0.189894
R8227 commonsourceibias.n217 commonsourceibias.n9 0.189894
R8228 commonsourceibias.n217 commonsourceibias.n216 0.189894
R8229 commonsourceibias.n216 commonsourceibias.n215 0.189894
R8230 commonsourceibias.n215 commonsourceibias.n12 0.189894
R8231 commonsourceibias.n210 commonsourceibias.n12 0.189894
R8232 commonsourceibias.n210 commonsourceibias.n209 0.189894
R8233 commonsourceibias.n209 commonsourceibias.n208 0.189894
R8234 commonsourceibias.n645 commonsourceibias.n644 0.189894
R8235 commonsourceibias.n645 commonsourceibias.n640 0.189894
R8236 commonsourceibias.n650 commonsourceibias.n640 0.189894
R8237 commonsourceibias.n651 commonsourceibias.n650 0.189894
R8238 commonsourceibias.n652 commonsourceibias.n651 0.189894
R8239 commonsourceibias.n652 commonsourceibias.n638 0.189894
R8240 commonsourceibias.n658 commonsourceibias.n638 0.189894
R8241 commonsourceibias.n659 commonsourceibias.n658 0.189894
R8242 commonsourceibias.n660 commonsourceibias.n659 0.189894
R8243 commonsourceibias.n660 commonsourceibias.n636 0.189894
R8244 commonsourceibias.n665 commonsourceibias.n636 0.189894
R8245 commonsourceibias.n666 commonsourceibias.n665 0.189894
R8246 commonsourceibias.n667 commonsourceibias.n666 0.189894
R8247 commonsourceibias.n667 commonsourceibias.n634 0.189894
R8248 commonsourceibias.n673 commonsourceibias.n634 0.189894
R8249 commonsourceibias.n674 commonsourceibias.n673 0.189894
R8250 commonsourceibias.n675 commonsourceibias.n674 0.189894
R8251 commonsourceibias.n675 commonsourceibias.n632 0.189894
R8252 commonsourceibias.n680 commonsourceibias.n632 0.189894
R8253 commonsourceibias.n681 commonsourceibias.n680 0.189894
R8254 commonsourceibias.n682 commonsourceibias.n681 0.189894
R8255 commonsourceibias.n682 commonsourceibias.n630 0.189894
R8256 commonsourceibias.n688 commonsourceibias.n630 0.189894
R8257 commonsourceibias.n689 commonsourceibias.n688 0.189894
R8258 commonsourceibias.n690 commonsourceibias.n689 0.189894
R8259 commonsourceibias.n690 commonsourceibias.n628 0.189894
R8260 commonsourceibias.n695 commonsourceibias.n628 0.189894
R8261 commonsourceibias.n696 commonsourceibias.n695 0.189894
R8262 commonsourceibias.n697 commonsourceibias.n696 0.189894
R8263 commonsourceibias.n697 commonsourceibias.n626 0.189894
R8264 commonsourceibias.n703 commonsourceibias.n626 0.189894
R8265 commonsourceibias.n704 commonsourceibias.n703 0.189894
R8266 commonsourceibias.n705 commonsourceibias.n704 0.189894
R8267 commonsourceibias.n705 commonsourceibias.n624 0.189894
R8268 commonsourceibias.n710 commonsourceibias.n624 0.189894
R8269 commonsourceibias.n711 commonsourceibias.n710 0.189894
R8270 commonsourceibias.n712 commonsourceibias.n711 0.189894
R8271 commonsourceibias.n712 commonsourceibias.n622 0.189894
R8272 commonsourceibias.n718 commonsourceibias.n622 0.189894
R8273 commonsourceibias.n719 commonsourceibias.n718 0.189894
R8274 commonsourceibias.n720 commonsourceibias.n719 0.189894
R8275 commonsourceibias.n720 commonsourceibias.n620 0.189894
R8276 commonsourceibias.n725 commonsourceibias.n620 0.189894
R8277 commonsourceibias.n726 commonsourceibias.n725 0.189894
R8278 commonsourceibias.n727 commonsourceibias.n726 0.189894
R8279 commonsourceibias.n727 commonsourceibias.n618 0.189894
R8280 commonsourceibias.n415 commonsourceibias.n414 0.189894
R8281 commonsourceibias.n415 commonsourceibias.n410 0.189894
R8282 commonsourceibias.n420 commonsourceibias.n410 0.189894
R8283 commonsourceibias.n421 commonsourceibias.n420 0.189894
R8284 commonsourceibias.n422 commonsourceibias.n421 0.189894
R8285 commonsourceibias.n422 commonsourceibias.n408 0.189894
R8286 commonsourceibias.n428 commonsourceibias.n408 0.189894
R8287 commonsourceibias.n429 commonsourceibias.n428 0.189894
R8288 commonsourceibias.n430 commonsourceibias.n429 0.189894
R8289 commonsourceibias.n430 commonsourceibias.n406 0.189894
R8290 commonsourceibias.n435 commonsourceibias.n406 0.189894
R8291 commonsourceibias.n436 commonsourceibias.n435 0.189894
R8292 commonsourceibias.n437 commonsourceibias.n436 0.189894
R8293 commonsourceibias.n437 commonsourceibias.n404 0.189894
R8294 commonsourceibias.n443 commonsourceibias.n404 0.189894
R8295 commonsourceibias.n444 commonsourceibias.n443 0.189894
R8296 commonsourceibias.n445 commonsourceibias.n444 0.189894
R8297 commonsourceibias.n445 commonsourceibias.n402 0.189894
R8298 commonsourceibias.n450 commonsourceibias.n402 0.189894
R8299 commonsourceibias.n451 commonsourceibias.n450 0.189894
R8300 commonsourceibias.n452 commonsourceibias.n451 0.189894
R8301 commonsourceibias.n452 commonsourceibias.n400 0.189894
R8302 commonsourceibias.n458 commonsourceibias.n400 0.189894
R8303 commonsourceibias.n459 commonsourceibias.n458 0.189894
R8304 commonsourceibias.n460 commonsourceibias.n459 0.189894
R8305 commonsourceibias.n460 commonsourceibias.n398 0.189894
R8306 commonsourceibias.n465 commonsourceibias.n398 0.189894
R8307 commonsourceibias.n466 commonsourceibias.n465 0.189894
R8308 commonsourceibias.n467 commonsourceibias.n466 0.189894
R8309 commonsourceibias.n467 commonsourceibias.n396 0.189894
R8310 commonsourceibias.n473 commonsourceibias.n396 0.189894
R8311 commonsourceibias.n474 commonsourceibias.n473 0.189894
R8312 commonsourceibias.n475 commonsourceibias.n474 0.189894
R8313 commonsourceibias.n475 commonsourceibias.n394 0.189894
R8314 commonsourceibias.n480 commonsourceibias.n394 0.189894
R8315 commonsourceibias.n481 commonsourceibias.n480 0.189894
R8316 commonsourceibias.n482 commonsourceibias.n481 0.189894
R8317 commonsourceibias.n482 commonsourceibias.n392 0.189894
R8318 commonsourceibias.n488 commonsourceibias.n392 0.189894
R8319 commonsourceibias.n489 commonsourceibias.n488 0.189894
R8320 commonsourceibias.n490 commonsourceibias.n489 0.189894
R8321 commonsourceibias.n490 commonsourceibias.n390 0.189894
R8322 commonsourceibias.n495 commonsourceibias.n390 0.189894
R8323 commonsourceibias.n496 commonsourceibias.n495 0.189894
R8324 commonsourceibias.n497 commonsourceibias.n496 0.189894
R8325 commonsourceibias.n497 commonsourceibias.n388 0.189894
R8326 commonsourceibias.n531 commonsourceibias.n530 0.189894
R8327 commonsourceibias.n531 commonsourceibias.n526 0.189894
R8328 commonsourceibias.n536 commonsourceibias.n526 0.189894
R8329 commonsourceibias.n537 commonsourceibias.n536 0.189894
R8330 commonsourceibias.n538 commonsourceibias.n537 0.189894
R8331 commonsourceibias.n538 commonsourceibias.n524 0.189894
R8332 commonsourceibias.n544 commonsourceibias.n524 0.189894
R8333 commonsourceibias.n545 commonsourceibias.n544 0.189894
R8334 commonsourceibias.n546 commonsourceibias.n545 0.189894
R8335 commonsourceibias.n546 commonsourceibias.n522 0.189894
R8336 commonsourceibias.n551 commonsourceibias.n522 0.189894
R8337 commonsourceibias.n552 commonsourceibias.n551 0.189894
R8338 commonsourceibias.n553 commonsourceibias.n552 0.189894
R8339 commonsourceibias.n553 commonsourceibias.n520 0.189894
R8340 commonsourceibias.n558 commonsourceibias.n520 0.189894
R8341 commonsourceibias.n559 commonsourceibias.n558 0.189894
R8342 commonsourceibias.n559 commonsourceibias.n518 0.189894
R8343 commonsourceibias.n563 commonsourceibias.n518 0.189894
R8344 commonsourceibias.n564 commonsourceibias.n563 0.189894
R8345 commonsourceibias.n564 commonsourceibias.n516 0.189894
R8346 commonsourceibias.n568 commonsourceibias.n516 0.189894
R8347 commonsourceibias.n569 commonsourceibias.n568 0.189894
R8348 commonsourceibias.n574 commonsourceibias.n573 0.189894
R8349 commonsourceibias.n575 commonsourceibias.n574 0.189894
R8350 commonsourceibias.n575 commonsourceibias.n377 0.189894
R8351 commonsourceibias.n580 commonsourceibias.n377 0.189894
R8352 commonsourceibias.n581 commonsourceibias.n580 0.189894
R8353 commonsourceibias.n582 commonsourceibias.n581 0.189894
R8354 commonsourceibias.n582 commonsourceibias.n375 0.189894
R8355 commonsourceibias.n588 commonsourceibias.n375 0.189894
R8356 commonsourceibias.n589 commonsourceibias.n588 0.189894
R8357 commonsourceibias.n590 commonsourceibias.n589 0.189894
R8358 commonsourceibias.n590 commonsourceibias.n373 0.189894
R8359 commonsourceibias.n595 commonsourceibias.n373 0.189894
R8360 commonsourceibias.n596 commonsourceibias.n595 0.189894
R8361 commonsourceibias.n597 commonsourceibias.n596 0.189894
R8362 commonsourceibias.n597 commonsourceibias.n371 0.189894
R8363 commonsourceibias.n603 commonsourceibias.n371 0.189894
R8364 commonsourceibias.n604 commonsourceibias.n603 0.189894
R8365 commonsourceibias.n605 commonsourceibias.n604 0.189894
R8366 commonsourceibias.n605 commonsourceibias.n369 0.189894
R8367 commonsourceibias.n610 commonsourceibias.n369 0.189894
R8368 commonsourceibias.n611 commonsourceibias.n610 0.189894
R8369 commonsourceibias.n612 commonsourceibias.n611 0.189894
R8370 commonsourceibias.n612 commonsourceibias.n367 0.189894
R8371 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R8372 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R8373 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R8374 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R8375 gnd.n2829 gnd.n2828 978.75
R8376 gnd.n4756 gnd.n4755 939.716
R8377 gnd.n5581 gnd.n1311 771.183
R8378 gnd.n6759 gnd.n6758 771.183
R8379 gnd.n5818 gnd.n1309 771.183
R8380 gnd.n6815 gnd.n632 771.183
R8381 gnd.n4663 gnd.n1989 766.379
R8382 gnd.n4666 gnd.n4665 766.379
R8383 gnd.n3968 gnd.n3871 766.379
R8384 gnd.n3964 gnd.n3869 766.379
R8385 gnd.n4754 gnd.n2011 756.769
R8386 gnd.n3363 gnd.n3362 756.769
R8387 gnd.n4061 gnd.n3778 756.769
R8388 gnd.n4059 gnd.n3781 756.769
R8389 gnd.n7417 gnd.n125 751.963
R8390 gnd.n7575 gnd.n7574 751.963
R8391 gnd.n6973 gnd.n517 751.963
R8392 gnd.n6621 gnd.n479 751.963
R8393 gnd.n5575 gnd.n1357 751.963
R8394 gnd.n5773 gnd.n5772 751.963
R8395 gnd.n4823 gnd.n4758 751.963
R8396 gnd.n5071 gnd.n1987 751.963
R8397 gnd.n7572 gnd.n127 732.745
R8398 gnd.n195 gnd.n123 732.745
R8399 gnd.n6976 gnd.n6975 732.745
R8400 gnd.n7048 gnd.n484 732.745
R8401 gnd.n5770 gnd.n1359 732.745
R8402 gnd.n5701 gnd.n1355 732.745
R8403 gnd.n4990 gnd.n4757 732.745
R8404 gnd.n5069 gnd.n4873 732.745
R8405 gnd.n3140 gnd.n2188 723.135
R8406 gnd.n2830 gnd.n2496 723.135
R8407 gnd.n7220 gnd.n343 723.135
R8408 gnd.n2064 gnd.n1798 723.135
R8409 gnd.n2188 gnd.n2187 585
R8410 gnd.n3142 gnd.n2188 585
R8411 gnd.n3145 gnd.n3144 585
R8412 gnd.n3144 gnd.n3143 585
R8413 gnd.n2185 gnd.n2184 585
R8414 gnd.n2184 gnd.n2183 585
R8415 gnd.n3150 gnd.n3149 585
R8416 gnd.n3151 gnd.n3150 585
R8417 gnd.n2182 gnd.n2181 585
R8418 gnd.n3152 gnd.n2182 585
R8419 gnd.n3155 gnd.n3154 585
R8420 gnd.n3154 gnd.n3153 585
R8421 gnd.n2179 gnd.n2178 585
R8422 gnd.n2178 gnd.n2177 585
R8423 gnd.n3160 gnd.n3159 585
R8424 gnd.n3161 gnd.n3160 585
R8425 gnd.n2176 gnd.n2175 585
R8426 gnd.n3162 gnd.n2176 585
R8427 gnd.n3165 gnd.n3164 585
R8428 gnd.n3164 gnd.n3163 585
R8429 gnd.n2173 gnd.n2172 585
R8430 gnd.n2172 gnd.n2171 585
R8431 gnd.n3170 gnd.n3169 585
R8432 gnd.n3171 gnd.n3170 585
R8433 gnd.n2170 gnd.n2169 585
R8434 gnd.n3172 gnd.n2170 585
R8435 gnd.n3175 gnd.n3174 585
R8436 gnd.n3174 gnd.n3173 585
R8437 gnd.n2167 gnd.n2166 585
R8438 gnd.n2166 gnd.n2165 585
R8439 gnd.n3180 gnd.n3179 585
R8440 gnd.n3181 gnd.n3180 585
R8441 gnd.n2164 gnd.n2163 585
R8442 gnd.n3182 gnd.n2164 585
R8443 gnd.n3185 gnd.n3184 585
R8444 gnd.n3184 gnd.n3183 585
R8445 gnd.n2161 gnd.n2160 585
R8446 gnd.n2160 gnd.n2159 585
R8447 gnd.n3190 gnd.n3189 585
R8448 gnd.n3191 gnd.n3190 585
R8449 gnd.n2158 gnd.n2157 585
R8450 gnd.n3192 gnd.n2158 585
R8451 gnd.n3195 gnd.n3194 585
R8452 gnd.n3194 gnd.n3193 585
R8453 gnd.n2155 gnd.n2154 585
R8454 gnd.n2154 gnd.n2153 585
R8455 gnd.n3200 gnd.n3199 585
R8456 gnd.n3201 gnd.n3200 585
R8457 gnd.n2152 gnd.n2151 585
R8458 gnd.n3202 gnd.n2152 585
R8459 gnd.n3205 gnd.n3204 585
R8460 gnd.n3204 gnd.n3203 585
R8461 gnd.n2149 gnd.n2148 585
R8462 gnd.n2148 gnd.n2147 585
R8463 gnd.n3210 gnd.n3209 585
R8464 gnd.n3211 gnd.n3210 585
R8465 gnd.n2146 gnd.n2145 585
R8466 gnd.n3212 gnd.n2146 585
R8467 gnd.n3215 gnd.n3214 585
R8468 gnd.n3214 gnd.n3213 585
R8469 gnd.n2143 gnd.n2142 585
R8470 gnd.n2142 gnd.n2141 585
R8471 gnd.n3220 gnd.n3219 585
R8472 gnd.n3221 gnd.n3220 585
R8473 gnd.n2140 gnd.n2139 585
R8474 gnd.n3222 gnd.n2140 585
R8475 gnd.n3225 gnd.n3224 585
R8476 gnd.n3224 gnd.n3223 585
R8477 gnd.n2137 gnd.n2136 585
R8478 gnd.n2136 gnd.n2135 585
R8479 gnd.n3230 gnd.n3229 585
R8480 gnd.n3231 gnd.n3230 585
R8481 gnd.n2134 gnd.n2133 585
R8482 gnd.n3232 gnd.n2134 585
R8483 gnd.n3235 gnd.n3234 585
R8484 gnd.n3234 gnd.n3233 585
R8485 gnd.n2131 gnd.n2130 585
R8486 gnd.n2130 gnd.n2129 585
R8487 gnd.n3240 gnd.n3239 585
R8488 gnd.n3241 gnd.n3240 585
R8489 gnd.n2128 gnd.n2127 585
R8490 gnd.n3242 gnd.n2128 585
R8491 gnd.n3245 gnd.n3244 585
R8492 gnd.n3244 gnd.n3243 585
R8493 gnd.n2125 gnd.n2124 585
R8494 gnd.n2124 gnd.n2123 585
R8495 gnd.n3250 gnd.n3249 585
R8496 gnd.n3251 gnd.n3250 585
R8497 gnd.n2122 gnd.n2121 585
R8498 gnd.n3252 gnd.n2122 585
R8499 gnd.n3255 gnd.n3254 585
R8500 gnd.n3254 gnd.n3253 585
R8501 gnd.n2119 gnd.n2118 585
R8502 gnd.n2118 gnd.n2117 585
R8503 gnd.n3260 gnd.n3259 585
R8504 gnd.n3261 gnd.n3260 585
R8505 gnd.n2116 gnd.n2115 585
R8506 gnd.n3262 gnd.n2116 585
R8507 gnd.n3265 gnd.n3264 585
R8508 gnd.n3264 gnd.n3263 585
R8509 gnd.n2113 gnd.n2112 585
R8510 gnd.n2112 gnd.n2111 585
R8511 gnd.n3270 gnd.n3269 585
R8512 gnd.n3271 gnd.n3270 585
R8513 gnd.n2110 gnd.n2109 585
R8514 gnd.n3272 gnd.n2110 585
R8515 gnd.n3275 gnd.n3274 585
R8516 gnd.n3274 gnd.n3273 585
R8517 gnd.n2107 gnd.n2106 585
R8518 gnd.n2106 gnd.n2105 585
R8519 gnd.n3280 gnd.n3279 585
R8520 gnd.n3281 gnd.n3280 585
R8521 gnd.n2104 gnd.n2103 585
R8522 gnd.n3282 gnd.n2104 585
R8523 gnd.n3285 gnd.n3284 585
R8524 gnd.n3284 gnd.n3283 585
R8525 gnd.n2101 gnd.n2100 585
R8526 gnd.n2100 gnd.n2099 585
R8527 gnd.n3290 gnd.n3289 585
R8528 gnd.n3291 gnd.n3290 585
R8529 gnd.n2098 gnd.n2097 585
R8530 gnd.n3292 gnd.n2098 585
R8531 gnd.n3295 gnd.n3294 585
R8532 gnd.n3294 gnd.n3293 585
R8533 gnd.n2095 gnd.n2094 585
R8534 gnd.n2094 gnd.n2093 585
R8535 gnd.n3300 gnd.n3299 585
R8536 gnd.n3301 gnd.n3300 585
R8537 gnd.n2092 gnd.n2091 585
R8538 gnd.n3302 gnd.n2092 585
R8539 gnd.n3305 gnd.n3304 585
R8540 gnd.n3304 gnd.n3303 585
R8541 gnd.n2089 gnd.n2088 585
R8542 gnd.n2088 gnd.n2087 585
R8543 gnd.n3310 gnd.n3309 585
R8544 gnd.n3311 gnd.n3310 585
R8545 gnd.n2086 gnd.n2085 585
R8546 gnd.n3312 gnd.n2086 585
R8547 gnd.n3315 gnd.n3314 585
R8548 gnd.n3314 gnd.n3313 585
R8549 gnd.n2083 gnd.n2082 585
R8550 gnd.n2082 gnd.n2081 585
R8551 gnd.n3320 gnd.n3319 585
R8552 gnd.n3321 gnd.n3320 585
R8553 gnd.n2080 gnd.n2079 585
R8554 gnd.n3322 gnd.n2080 585
R8555 gnd.n3325 gnd.n3324 585
R8556 gnd.n3324 gnd.n3323 585
R8557 gnd.n2077 gnd.n2076 585
R8558 gnd.n2076 gnd.n2075 585
R8559 gnd.n3330 gnd.n3329 585
R8560 gnd.n3331 gnd.n3330 585
R8561 gnd.n2074 gnd.n2073 585
R8562 gnd.n3332 gnd.n2074 585
R8563 gnd.n3335 gnd.n3334 585
R8564 gnd.n3334 gnd.n3333 585
R8565 gnd.n2071 gnd.n2070 585
R8566 gnd.n2070 gnd.n2069 585
R8567 gnd.n3340 gnd.n3339 585
R8568 gnd.n3341 gnd.n3340 585
R8569 gnd.n2068 gnd.n2067 585
R8570 gnd.n3342 gnd.n2068 585
R8571 gnd.n3345 gnd.n3344 585
R8572 gnd.n3344 gnd.n3343 585
R8573 gnd.n2065 gnd.n2063 585
R8574 gnd.n2063 gnd.n2062 585
R8575 gnd.n3353 gnd.n3352 585
R8576 gnd.n3354 gnd.n3353 585
R8577 gnd.n3140 gnd.n3139 585
R8578 gnd.n3141 gnd.n3140 585
R8579 gnd.n2191 gnd.n2190 585
R8580 gnd.n2190 gnd.n2189 585
R8581 gnd.n3135 gnd.n3134 585
R8582 gnd.n3134 gnd.n3133 585
R8583 gnd.n2194 gnd.n2193 585
R8584 gnd.n3132 gnd.n2194 585
R8585 gnd.n3130 gnd.n3129 585
R8586 gnd.n3131 gnd.n3130 585
R8587 gnd.n3128 gnd.n2196 585
R8588 gnd.n2196 gnd.n2195 585
R8589 gnd.n3127 gnd.n3126 585
R8590 gnd.n3126 gnd.n3125 585
R8591 gnd.n2201 gnd.n2200 585
R8592 gnd.n3124 gnd.n2201 585
R8593 gnd.n3122 gnd.n3121 585
R8594 gnd.n3123 gnd.n3122 585
R8595 gnd.n3120 gnd.n2203 585
R8596 gnd.n2203 gnd.n2202 585
R8597 gnd.n3119 gnd.n3118 585
R8598 gnd.n3118 gnd.n3117 585
R8599 gnd.n2209 gnd.n2208 585
R8600 gnd.n3116 gnd.n2209 585
R8601 gnd.n3114 gnd.n3113 585
R8602 gnd.n3115 gnd.n3114 585
R8603 gnd.n3112 gnd.n2211 585
R8604 gnd.n2211 gnd.n2210 585
R8605 gnd.n3111 gnd.n3110 585
R8606 gnd.n3110 gnd.n3109 585
R8607 gnd.n2217 gnd.n2216 585
R8608 gnd.n3108 gnd.n2217 585
R8609 gnd.n3106 gnd.n3105 585
R8610 gnd.n3107 gnd.n3106 585
R8611 gnd.n3104 gnd.n2219 585
R8612 gnd.n2219 gnd.n2218 585
R8613 gnd.n3103 gnd.n3102 585
R8614 gnd.n3102 gnd.n3101 585
R8615 gnd.n2225 gnd.n2224 585
R8616 gnd.n3100 gnd.n2225 585
R8617 gnd.n3098 gnd.n3097 585
R8618 gnd.n3099 gnd.n3098 585
R8619 gnd.n3096 gnd.n2227 585
R8620 gnd.n2227 gnd.n2226 585
R8621 gnd.n3095 gnd.n3094 585
R8622 gnd.n3094 gnd.n3093 585
R8623 gnd.n2233 gnd.n2232 585
R8624 gnd.n3092 gnd.n2233 585
R8625 gnd.n3090 gnd.n3089 585
R8626 gnd.n3091 gnd.n3090 585
R8627 gnd.n3088 gnd.n2235 585
R8628 gnd.n2235 gnd.n2234 585
R8629 gnd.n3087 gnd.n3086 585
R8630 gnd.n3086 gnd.n3085 585
R8631 gnd.n2241 gnd.n2240 585
R8632 gnd.n3084 gnd.n2241 585
R8633 gnd.n3082 gnd.n3081 585
R8634 gnd.n3083 gnd.n3082 585
R8635 gnd.n3080 gnd.n2243 585
R8636 gnd.n2243 gnd.n2242 585
R8637 gnd.n3079 gnd.n3078 585
R8638 gnd.n3078 gnd.n3077 585
R8639 gnd.n2249 gnd.n2248 585
R8640 gnd.n3076 gnd.n2249 585
R8641 gnd.n3074 gnd.n3073 585
R8642 gnd.n3075 gnd.n3074 585
R8643 gnd.n3072 gnd.n2251 585
R8644 gnd.n2251 gnd.n2250 585
R8645 gnd.n3071 gnd.n3070 585
R8646 gnd.n3070 gnd.n3069 585
R8647 gnd.n2257 gnd.n2256 585
R8648 gnd.n3068 gnd.n2257 585
R8649 gnd.n3066 gnd.n3065 585
R8650 gnd.n3067 gnd.n3066 585
R8651 gnd.n3064 gnd.n2259 585
R8652 gnd.n2259 gnd.n2258 585
R8653 gnd.n3063 gnd.n3062 585
R8654 gnd.n3062 gnd.n3061 585
R8655 gnd.n2265 gnd.n2264 585
R8656 gnd.n3060 gnd.n2265 585
R8657 gnd.n3058 gnd.n3057 585
R8658 gnd.n3059 gnd.n3058 585
R8659 gnd.n3056 gnd.n2267 585
R8660 gnd.n2267 gnd.n2266 585
R8661 gnd.n3055 gnd.n3054 585
R8662 gnd.n3054 gnd.n3053 585
R8663 gnd.n2273 gnd.n2272 585
R8664 gnd.n3052 gnd.n2273 585
R8665 gnd.n3050 gnd.n3049 585
R8666 gnd.n3051 gnd.n3050 585
R8667 gnd.n3048 gnd.n2275 585
R8668 gnd.n2275 gnd.n2274 585
R8669 gnd.n3047 gnd.n3046 585
R8670 gnd.n3046 gnd.n3045 585
R8671 gnd.n2281 gnd.n2280 585
R8672 gnd.n3044 gnd.n2281 585
R8673 gnd.n3042 gnd.n3041 585
R8674 gnd.n3043 gnd.n3042 585
R8675 gnd.n3040 gnd.n2283 585
R8676 gnd.n2283 gnd.n2282 585
R8677 gnd.n3039 gnd.n3038 585
R8678 gnd.n3038 gnd.n3037 585
R8679 gnd.n2289 gnd.n2288 585
R8680 gnd.n3036 gnd.n2289 585
R8681 gnd.n3034 gnd.n3033 585
R8682 gnd.n3035 gnd.n3034 585
R8683 gnd.n3032 gnd.n2291 585
R8684 gnd.n2291 gnd.n2290 585
R8685 gnd.n3031 gnd.n3030 585
R8686 gnd.n3030 gnd.n3029 585
R8687 gnd.n2297 gnd.n2296 585
R8688 gnd.n3028 gnd.n2297 585
R8689 gnd.n3026 gnd.n3025 585
R8690 gnd.n3027 gnd.n3026 585
R8691 gnd.n3024 gnd.n2299 585
R8692 gnd.n2299 gnd.n2298 585
R8693 gnd.n3023 gnd.n3022 585
R8694 gnd.n3022 gnd.n3021 585
R8695 gnd.n2305 gnd.n2304 585
R8696 gnd.n3020 gnd.n2305 585
R8697 gnd.n3018 gnd.n3017 585
R8698 gnd.n3019 gnd.n3018 585
R8699 gnd.n3016 gnd.n2307 585
R8700 gnd.n2307 gnd.n2306 585
R8701 gnd.n3015 gnd.n3014 585
R8702 gnd.n3014 gnd.n3013 585
R8703 gnd.n2313 gnd.n2312 585
R8704 gnd.n3012 gnd.n2313 585
R8705 gnd.n3010 gnd.n3009 585
R8706 gnd.n3011 gnd.n3010 585
R8707 gnd.n3008 gnd.n2315 585
R8708 gnd.n2315 gnd.n2314 585
R8709 gnd.n3007 gnd.n3006 585
R8710 gnd.n3006 gnd.n3005 585
R8711 gnd.n2321 gnd.n2320 585
R8712 gnd.n3004 gnd.n2321 585
R8713 gnd.n3002 gnd.n3001 585
R8714 gnd.n3003 gnd.n3002 585
R8715 gnd.n3000 gnd.n2323 585
R8716 gnd.n2323 gnd.n2322 585
R8717 gnd.n2999 gnd.n2998 585
R8718 gnd.n2998 gnd.n2997 585
R8719 gnd.n2329 gnd.n2328 585
R8720 gnd.n2996 gnd.n2329 585
R8721 gnd.n2994 gnd.n2993 585
R8722 gnd.n2995 gnd.n2994 585
R8723 gnd.n2992 gnd.n2331 585
R8724 gnd.n2331 gnd.n2330 585
R8725 gnd.n2991 gnd.n2990 585
R8726 gnd.n2990 gnd.n2989 585
R8727 gnd.n2337 gnd.n2336 585
R8728 gnd.n2988 gnd.n2337 585
R8729 gnd.n2986 gnd.n2985 585
R8730 gnd.n2987 gnd.n2986 585
R8731 gnd.n2984 gnd.n2339 585
R8732 gnd.n2339 gnd.n2338 585
R8733 gnd.n2983 gnd.n2982 585
R8734 gnd.n2982 gnd.n2981 585
R8735 gnd.n2345 gnd.n2344 585
R8736 gnd.n2980 gnd.n2345 585
R8737 gnd.n2978 gnd.n2977 585
R8738 gnd.n2979 gnd.n2978 585
R8739 gnd.n2976 gnd.n2347 585
R8740 gnd.n2347 gnd.n2346 585
R8741 gnd.n2975 gnd.n2974 585
R8742 gnd.n2974 gnd.n2973 585
R8743 gnd.n2353 gnd.n2352 585
R8744 gnd.n2972 gnd.n2353 585
R8745 gnd.n2970 gnd.n2969 585
R8746 gnd.n2971 gnd.n2970 585
R8747 gnd.n2968 gnd.n2355 585
R8748 gnd.n2355 gnd.n2354 585
R8749 gnd.n2967 gnd.n2966 585
R8750 gnd.n2966 gnd.n2965 585
R8751 gnd.n2361 gnd.n2360 585
R8752 gnd.n2964 gnd.n2361 585
R8753 gnd.n2962 gnd.n2961 585
R8754 gnd.n2963 gnd.n2962 585
R8755 gnd.n2960 gnd.n2363 585
R8756 gnd.n2363 gnd.n2362 585
R8757 gnd.n2959 gnd.n2958 585
R8758 gnd.n2958 gnd.n2957 585
R8759 gnd.n2369 gnd.n2368 585
R8760 gnd.n2956 gnd.n2369 585
R8761 gnd.n2954 gnd.n2953 585
R8762 gnd.n2955 gnd.n2954 585
R8763 gnd.n2952 gnd.n2371 585
R8764 gnd.n2371 gnd.n2370 585
R8765 gnd.n2951 gnd.n2950 585
R8766 gnd.n2950 gnd.n2949 585
R8767 gnd.n2377 gnd.n2376 585
R8768 gnd.n2948 gnd.n2377 585
R8769 gnd.n2946 gnd.n2945 585
R8770 gnd.n2947 gnd.n2946 585
R8771 gnd.n2944 gnd.n2379 585
R8772 gnd.n2379 gnd.n2378 585
R8773 gnd.n2943 gnd.n2942 585
R8774 gnd.n2942 gnd.n2941 585
R8775 gnd.n2385 gnd.n2384 585
R8776 gnd.n2940 gnd.n2385 585
R8777 gnd.n2938 gnd.n2937 585
R8778 gnd.n2939 gnd.n2938 585
R8779 gnd.n2936 gnd.n2387 585
R8780 gnd.n2387 gnd.n2386 585
R8781 gnd.n2935 gnd.n2934 585
R8782 gnd.n2934 gnd.n2933 585
R8783 gnd.n2393 gnd.n2392 585
R8784 gnd.n2932 gnd.n2393 585
R8785 gnd.n2930 gnd.n2929 585
R8786 gnd.n2931 gnd.n2930 585
R8787 gnd.n2928 gnd.n2395 585
R8788 gnd.n2395 gnd.n2394 585
R8789 gnd.n2927 gnd.n2926 585
R8790 gnd.n2926 gnd.n2925 585
R8791 gnd.n2401 gnd.n2400 585
R8792 gnd.n2924 gnd.n2401 585
R8793 gnd.n2922 gnd.n2921 585
R8794 gnd.n2923 gnd.n2922 585
R8795 gnd.n2920 gnd.n2403 585
R8796 gnd.n2403 gnd.n2402 585
R8797 gnd.n2919 gnd.n2918 585
R8798 gnd.n2918 gnd.n2917 585
R8799 gnd.n2409 gnd.n2408 585
R8800 gnd.n2916 gnd.n2409 585
R8801 gnd.n2914 gnd.n2913 585
R8802 gnd.n2915 gnd.n2914 585
R8803 gnd.n2912 gnd.n2411 585
R8804 gnd.n2411 gnd.n2410 585
R8805 gnd.n2911 gnd.n2910 585
R8806 gnd.n2910 gnd.n2909 585
R8807 gnd.n2417 gnd.n2416 585
R8808 gnd.n2908 gnd.n2417 585
R8809 gnd.n2906 gnd.n2905 585
R8810 gnd.n2907 gnd.n2906 585
R8811 gnd.n2904 gnd.n2419 585
R8812 gnd.n2419 gnd.n2418 585
R8813 gnd.n2903 gnd.n2902 585
R8814 gnd.n2902 gnd.n2901 585
R8815 gnd.n2425 gnd.n2424 585
R8816 gnd.n2900 gnd.n2425 585
R8817 gnd.n2898 gnd.n2897 585
R8818 gnd.n2899 gnd.n2898 585
R8819 gnd.n2896 gnd.n2427 585
R8820 gnd.n2427 gnd.n2426 585
R8821 gnd.n2895 gnd.n2894 585
R8822 gnd.n2894 gnd.n2893 585
R8823 gnd.n2433 gnd.n2432 585
R8824 gnd.n2892 gnd.n2433 585
R8825 gnd.n2890 gnd.n2889 585
R8826 gnd.n2891 gnd.n2890 585
R8827 gnd.n2888 gnd.n2435 585
R8828 gnd.n2435 gnd.n2434 585
R8829 gnd.n2887 gnd.n2886 585
R8830 gnd.n2886 gnd.n2885 585
R8831 gnd.n2441 gnd.n2440 585
R8832 gnd.n2884 gnd.n2441 585
R8833 gnd.n2882 gnd.n2881 585
R8834 gnd.n2883 gnd.n2882 585
R8835 gnd.n2880 gnd.n2443 585
R8836 gnd.n2443 gnd.n2442 585
R8837 gnd.n2879 gnd.n2878 585
R8838 gnd.n2878 gnd.n2877 585
R8839 gnd.n2449 gnd.n2448 585
R8840 gnd.n2876 gnd.n2449 585
R8841 gnd.n2874 gnd.n2873 585
R8842 gnd.n2875 gnd.n2874 585
R8843 gnd.n2872 gnd.n2451 585
R8844 gnd.n2451 gnd.n2450 585
R8845 gnd.n2871 gnd.n2870 585
R8846 gnd.n2870 gnd.n2869 585
R8847 gnd.n2457 gnd.n2456 585
R8848 gnd.n2868 gnd.n2457 585
R8849 gnd.n2866 gnd.n2865 585
R8850 gnd.n2867 gnd.n2866 585
R8851 gnd.n2864 gnd.n2459 585
R8852 gnd.n2459 gnd.n2458 585
R8853 gnd.n2863 gnd.n2862 585
R8854 gnd.n2862 gnd.n2861 585
R8855 gnd.n2465 gnd.n2464 585
R8856 gnd.n2860 gnd.n2465 585
R8857 gnd.n2858 gnd.n2857 585
R8858 gnd.n2859 gnd.n2858 585
R8859 gnd.n2856 gnd.n2467 585
R8860 gnd.n2467 gnd.n2466 585
R8861 gnd.n2855 gnd.n2854 585
R8862 gnd.n2854 gnd.n2853 585
R8863 gnd.n2473 gnd.n2472 585
R8864 gnd.n2852 gnd.n2473 585
R8865 gnd.n2850 gnd.n2849 585
R8866 gnd.n2851 gnd.n2850 585
R8867 gnd.n2848 gnd.n2475 585
R8868 gnd.n2475 gnd.n2474 585
R8869 gnd.n2847 gnd.n2846 585
R8870 gnd.n2846 gnd.n2845 585
R8871 gnd.n2481 gnd.n2480 585
R8872 gnd.n2844 gnd.n2481 585
R8873 gnd.n2842 gnd.n2841 585
R8874 gnd.n2843 gnd.n2842 585
R8875 gnd.n2840 gnd.n2483 585
R8876 gnd.n2483 gnd.n2482 585
R8877 gnd.n2839 gnd.n2838 585
R8878 gnd.n2838 gnd.n2837 585
R8879 gnd.n2489 gnd.n2488 585
R8880 gnd.n2836 gnd.n2489 585
R8881 gnd.n2834 gnd.n2833 585
R8882 gnd.n2835 gnd.n2834 585
R8883 gnd.n2832 gnd.n2491 585
R8884 gnd.n2491 gnd.n2490 585
R8885 gnd.n2831 gnd.n2830 585
R8886 gnd.n2830 gnd.n2829 585
R8887 gnd.n344 gnd.n342 585
R8888 gnd.n2656 gnd.n342 585
R8889 gnd.n2662 gnd.n2658 585
R8890 gnd.n2658 gnd.n2657 585
R8891 gnd.n2664 gnd.n2663 585
R8892 gnd.n2665 gnd.n2664 585
R8893 gnd.n2655 gnd.n2654 585
R8894 gnd.n2666 gnd.n2655 585
R8895 gnd.n2669 gnd.n2668 585
R8896 gnd.n2668 gnd.n2667 585
R8897 gnd.n2670 gnd.n2649 585
R8898 gnd.n2649 gnd.n2648 585
R8899 gnd.n2672 gnd.n2671 585
R8900 gnd.n2673 gnd.n2672 585
R8901 gnd.n2647 gnd.n2646 585
R8902 gnd.n2674 gnd.n2647 585
R8903 gnd.n2677 gnd.n2676 585
R8904 gnd.n2676 gnd.n2675 585
R8905 gnd.n2678 gnd.n2641 585
R8906 gnd.n2641 gnd.n2640 585
R8907 gnd.n2680 gnd.n2679 585
R8908 gnd.n2681 gnd.n2680 585
R8909 gnd.n2639 gnd.n2638 585
R8910 gnd.n2682 gnd.n2639 585
R8911 gnd.n2685 gnd.n2684 585
R8912 gnd.n2684 gnd.n2683 585
R8913 gnd.n2686 gnd.n2633 585
R8914 gnd.n2633 gnd.n2632 585
R8915 gnd.n2688 gnd.n2687 585
R8916 gnd.n2689 gnd.n2688 585
R8917 gnd.n2631 gnd.n2630 585
R8918 gnd.n2690 gnd.n2631 585
R8919 gnd.n2693 gnd.n2692 585
R8920 gnd.n2692 gnd.n2691 585
R8921 gnd.n2694 gnd.n2625 585
R8922 gnd.n2625 gnd.n2624 585
R8923 gnd.n2696 gnd.n2695 585
R8924 gnd.n2697 gnd.n2696 585
R8925 gnd.n2623 gnd.n2622 585
R8926 gnd.n2698 gnd.n2623 585
R8927 gnd.n2701 gnd.n2700 585
R8928 gnd.n2700 gnd.n2699 585
R8929 gnd.n2702 gnd.n2617 585
R8930 gnd.n2617 gnd.n2616 585
R8931 gnd.n2704 gnd.n2703 585
R8932 gnd.n2705 gnd.n2704 585
R8933 gnd.n2615 gnd.n2614 585
R8934 gnd.n2706 gnd.n2615 585
R8935 gnd.n2709 gnd.n2708 585
R8936 gnd.n2708 gnd.n2707 585
R8937 gnd.n2710 gnd.n2609 585
R8938 gnd.n2609 gnd.n2608 585
R8939 gnd.n2712 gnd.n2711 585
R8940 gnd.n2713 gnd.n2712 585
R8941 gnd.n2607 gnd.n2606 585
R8942 gnd.n2714 gnd.n2607 585
R8943 gnd.n2717 gnd.n2716 585
R8944 gnd.n2716 gnd.n2715 585
R8945 gnd.n2718 gnd.n2601 585
R8946 gnd.n2601 gnd.n2600 585
R8947 gnd.n2720 gnd.n2719 585
R8948 gnd.n2721 gnd.n2720 585
R8949 gnd.n2599 gnd.n2598 585
R8950 gnd.n2722 gnd.n2599 585
R8951 gnd.n2725 gnd.n2724 585
R8952 gnd.n2724 gnd.n2723 585
R8953 gnd.n2726 gnd.n2593 585
R8954 gnd.n2593 gnd.n2592 585
R8955 gnd.n2728 gnd.n2727 585
R8956 gnd.n2729 gnd.n2728 585
R8957 gnd.n2591 gnd.n2590 585
R8958 gnd.n2730 gnd.n2591 585
R8959 gnd.n2733 gnd.n2732 585
R8960 gnd.n2732 gnd.n2731 585
R8961 gnd.n2734 gnd.n2585 585
R8962 gnd.n2585 gnd.n2584 585
R8963 gnd.n2736 gnd.n2735 585
R8964 gnd.n2737 gnd.n2736 585
R8965 gnd.n2583 gnd.n2582 585
R8966 gnd.n2738 gnd.n2583 585
R8967 gnd.n2741 gnd.n2740 585
R8968 gnd.n2740 gnd.n2739 585
R8969 gnd.n2742 gnd.n2577 585
R8970 gnd.n2577 gnd.n2576 585
R8971 gnd.n2744 gnd.n2743 585
R8972 gnd.n2745 gnd.n2744 585
R8973 gnd.n2575 gnd.n2574 585
R8974 gnd.n2746 gnd.n2575 585
R8975 gnd.n2749 gnd.n2748 585
R8976 gnd.n2748 gnd.n2747 585
R8977 gnd.n2750 gnd.n2569 585
R8978 gnd.n2569 gnd.n2568 585
R8979 gnd.n2752 gnd.n2751 585
R8980 gnd.n2753 gnd.n2752 585
R8981 gnd.n2567 gnd.n2566 585
R8982 gnd.n2754 gnd.n2567 585
R8983 gnd.n2757 gnd.n2756 585
R8984 gnd.n2756 gnd.n2755 585
R8985 gnd.n2758 gnd.n2561 585
R8986 gnd.n2561 gnd.n2560 585
R8987 gnd.n2760 gnd.n2759 585
R8988 gnd.n2761 gnd.n2760 585
R8989 gnd.n2559 gnd.n2558 585
R8990 gnd.n2762 gnd.n2559 585
R8991 gnd.n2765 gnd.n2764 585
R8992 gnd.n2764 gnd.n2763 585
R8993 gnd.n2766 gnd.n2553 585
R8994 gnd.n2553 gnd.n2552 585
R8995 gnd.n2768 gnd.n2767 585
R8996 gnd.n2769 gnd.n2768 585
R8997 gnd.n2551 gnd.n2550 585
R8998 gnd.n2770 gnd.n2551 585
R8999 gnd.n2773 gnd.n2772 585
R9000 gnd.n2772 gnd.n2771 585
R9001 gnd.n2774 gnd.n2545 585
R9002 gnd.n2545 gnd.n2544 585
R9003 gnd.n2776 gnd.n2775 585
R9004 gnd.n2777 gnd.n2776 585
R9005 gnd.n2543 gnd.n2542 585
R9006 gnd.n2778 gnd.n2543 585
R9007 gnd.n2781 gnd.n2780 585
R9008 gnd.n2780 gnd.n2779 585
R9009 gnd.n2782 gnd.n2537 585
R9010 gnd.n2537 gnd.n2536 585
R9011 gnd.n2784 gnd.n2783 585
R9012 gnd.n2785 gnd.n2784 585
R9013 gnd.n2535 gnd.n2534 585
R9014 gnd.n2786 gnd.n2535 585
R9015 gnd.n2789 gnd.n2788 585
R9016 gnd.n2788 gnd.n2787 585
R9017 gnd.n2790 gnd.n2529 585
R9018 gnd.n2529 gnd.n2528 585
R9019 gnd.n2792 gnd.n2791 585
R9020 gnd.n2793 gnd.n2792 585
R9021 gnd.n2527 gnd.n2526 585
R9022 gnd.n2794 gnd.n2527 585
R9023 gnd.n2797 gnd.n2796 585
R9024 gnd.n2796 gnd.n2795 585
R9025 gnd.n2798 gnd.n2521 585
R9026 gnd.n2521 gnd.n2520 585
R9027 gnd.n2800 gnd.n2799 585
R9028 gnd.n2801 gnd.n2800 585
R9029 gnd.n2519 gnd.n2518 585
R9030 gnd.n2802 gnd.n2519 585
R9031 gnd.n2805 gnd.n2804 585
R9032 gnd.n2804 gnd.n2803 585
R9033 gnd.n2806 gnd.n2513 585
R9034 gnd.n2513 gnd.n2512 585
R9035 gnd.n2808 gnd.n2807 585
R9036 gnd.n2809 gnd.n2808 585
R9037 gnd.n2511 gnd.n2510 585
R9038 gnd.n2810 gnd.n2511 585
R9039 gnd.n2813 gnd.n2812 585
R9040 gnd.n2812 gnd.n2811 585
R9041 gnd.n2814 gnd.n2506 585
R9042 gnd.n2506 gnd.n2505 585
R9043 gnd.n2816 gnd.n2815 585
R9044 gnd.n2817 gnd.n2816 585
R9045 gnd.n2504 gnd.n2503 585
R9046 gnd.n2818 gnd.n2504 585
R9047 gnd.n2821 gnd.n2820 585
R9048 gnd.n2820 gnd.n2819 585
R9049 gnd.n2500 gnd.n2498 585
R9050 gnd.n2498 gnd.n2497 585
R9051 gnd.n2826 gnd.n2825 585
R9052 gnd.n2827 gnd.n2826 585
R9053 gnd.n2499 gnd.n2496 585
R9054 gnd.n2828 gnd.n2496 585
R9055 gnd.n5691 gnd.n1357 585
R9056 gnd.n5771 gnd.n1357 585
R9057 gnd.n5693 gnd.n5692 585
R9058 gnd.n5694 gnd.n5693 585
R9059 gnd.n1651 gnd.n1650 585
R9060 gnd.n5386 gnd.n1650 585
R9061 gnd.n5569 gnd.n5568 585
R9062 gnd.n5568 gnd.n5567 585
R9063 gnd.n1654 gnd.n1653 585
R9064 gnd.n5384 gnd.n1654 585
R9065 gnd.n5556 gnd.n5555 585
R9066 gnd.n5557 gnd.n5556 585
R9067 gnd.n1670 gnd.n1669 585
R9068 gnd.n5373 gnd.n1669 585
R9069 gnd.n5551 gnd.n5550 585
R9070 gnd.n5550 gnd.n5549 585
R9071 gnd.n1673 gnd.n1672 585
R9072 gnd.n5328 gnd.n1673 585
R9073 gnd.n5540 gnd.n5539 585
R9074 gnd.n5541 gnd.n5540 585
R9075 gnd.n1686 gnd.n1685 585
R9076 gnd.n5334 gnd.n1685 585
R9077 gnd.n5535 gnd.n5534 585
R9078 gnd.n5534 gnd.n5533 585
R9079 gnd.n1689 gnd.n1688 585
R9080 gnd.n5320 gnd.n1689 585
R9081 gnd.n5524 gnd.n5523 585
R9082 gnd.n5525 gnd.n5524 585
R9083 gnd.n1704 gnd.n1703 585
R9084 gnd.n5316 gnd.n1703 585
R9085 gnd.n5519 gnd.n5518 585
R9086 gnd.n5518 gnd.n5517 585
R9087 gnd.n1707 gnd.n1706 585
R9088 gnd.n5289 gnd.n1707 585
R9089 gnd.n5508 gnd.n5507 585
R9090 gnd.n5509 gnd.n5508 585
R9091 gnd.n1720 gnd.n1719 585
R9092 gnd.n5295 gnd.n1719 585
R9093 gnd.n5503 gnd.n5502 585
R9094 gnd.n5502 gnd.n5501 585
R9095 gnd.n1723 gnd.n1722 585
R9096 gnd.n5280 gnd.n1723 585
R9097 gnd.n5492 gnd.n5491 585
R9098 gnd.n5493 gnd.n5492 585
R9099 gnd.n1738 gnd.n1737 585
R9100 gnd.n5276 gnd.n1737 585
R9101 gnd.n5487 gnd.n5486 585
R9102 gnd.n5486 gnd.n5485 585
R9103 gnd.n1741 gnd.n1740 585
R9104 gnd.n5249 gnd.n1741 585
R9105 gnd.n5476 gnd.n5475 585
R9106 gnd.n5477 gnd.n5476 585
R9107 gnd.n1754 gnd.n1753 585
R9108 gnd.n5429 gnd.n1753 585
R9109 gnd.n5471 gnd.n5470 585
R9110 gnd.n5470 gnd.n5469 585
R9111 gnd.n1757 gnd.n1756 585
R9112 gnd.n5241 gnd.n1757 585
R9113 gnd.n5443 gnd.n5442 585
R9114 gnd.n5442 gnd.n5441 585
R9115 gnd.n5444 gnd.n1791 585
R9116 gnd.n5233 gnd.n1791 585
R9117 gnd.n5446 gnd.n5445 585
R9118 gnd.n5447 gnd.n5446 585
R9119 gnd.n1783 gnd.n1782 585
R9120 gnd.n1786 gnd.n1783 585
R9121 gnd.n5457 gnd.n5456 585
R9122 gnd.n5456 gnd.n5455 585
R9123 gnd.n5458 gnd.n1777 585
R9124 gnd.n1777 gnd.n1775 585
R9125 gnd.n5460 gnd.n5459 585
R9126 gnd.n5461 gnd.n5460 585
R9127 gnd.n1778 gnd.n1776 585
R9128 gnd.n5217 gnd.n1776 585
R9129 gnd.n1895 gnd.n1894 585
R9130 gnd.n1894 gnd.n1867 585
R9131 gnd.n1896 gnd.n1874 585
R9132 gnd.n5199 gnd.n1874 585
R9133 gnd.n5186 gnd.n5185 585
R9134 gnd.n5185 gnd.n5184 585
R9135 gnd.n5187 gnd.n1886 585
R9136 gnd.n1886 gnd.n1884 585
R9137 gnd.n5189 gnd.n5188 585
R9138 gnd.n5190 gnd.n5189 585
R9139 gnd.n1887 gnd.n1885 585
R9140 gnd.n5173 gnd.n1885 585
R9141 gnd.n5145 gnd.n5144 585
R9142 gnd.n5144 gnd.n1902 585
R9143 gnd.n5146 gnd.n1910 585
R9144 gnd.n5160 gnd.n1910 585
R9145 gnd.n5147 gnd.n1920 585
R9146 gnd.n1920 gnd.n1908 585
R9147 gnd.n5149 gnd.n5148 585
R9148 gnd.n5150 gnd.n5149 585
R9149 gnd.n1921 gnd.n1919 585
R9150 gnd.n1928 gnd.n1919 585
R9151 gnd.n5136 gnd.n5135 585
R9152 gnd.n5135 gnd.n5134 585
R9153 gnd.n1924 gnd.n1923 585
R9154 gnd.n1925 gnd.n1924 585
R9155 gnd.n5125 gnd.n5124 585
R9156 gnd.n5126 gnd.n5125 585
R9157 gnd.n1938 gnd.n1937 585
R9158 gnd.n1937 gnd.n1934 585
R9159 gnd.n5120 gnd.n5119 585
R9160 gnd.n5119 gnd.n5118 585
R9161 gnd.n1941 gnd.n1940 585
R9162 gnd.n1942 gnd.n1941 585
R9163 gnd.n5109 gnd.n5108 585
R9164 gnd.n5110 gnd.n5109 585
R9165 gnd.n1953 gnd.n1952 585
R9166 gnd.n1960 gnd.n1952 585
R9167 gnd.n5104 gnd.n5103 585
R9168 gnd.n5103 gnd.n5102 585
R9169 gnd.n1956 gnd.n1955 585
R9170 gnd.n1957 gnd.n1956 585
R9171 gnd.n5093 gnd.n5092 585
R9172 gnd.n5094 gnd.n5093 585
R9173 gnd.n1970 gnd.n1969 585
R9174 gnd.n1969 gnd.n1966 585
R9175 gnd.n5088 gnd.n5087 585
R9176 gnd.n5087 gnd.n5086 585
R9177 gnd.n1973 gnd.n1972 585
R9178 gnd.n1974 gnd.n1973 585
R9179 gnd.n5077 gnd.n5076 585
R9180 gnd.n5078 gnd.n5077 585
R9181 gnd.n1985 gnd.n1984 585
R9182 gnd.n4872 gnd.n1984 585
R9183 gnd.n5072 gnd.n5071 585
R9184 gnd.n5071 gnd.n5070 585
R9185 gnd.n4779 gnd.n1987 585
R9186 gnd.n4782 gnd.n4780 585
R9187 gnd.n4785 gnd.n4784 585
R9188 gnd.n4777 gnd.n4776 585
R9189 gnd.n4790 gnd.n4789 585
R9190 gnd.n4792 gnd.n4775 585
R9191 gnd.n4795 gnd.n4794 585
R9192 gnd.n4773 gnd.n4772 585
R9193 gnd.n4800 gnd.n4799 585
R9194 gnd.n4802 gnd.n4771 585
R9195 gnd.n4805 gnd.n4804 585
R9196 gnd.n4769 gnd.n4768 585
R9197 gnd.n4810 gnd.n4809 585
R9198 gnd.n4812 gnd.n4767 585
R9199 gnd.n4815 gnd.n4814 585
R9200 gnd.n4765 gnd.n4764 585
R9201 gnd.n4820 gnd.n4819 585
R9202 gnd.n4822 gnd.n4763 585
R9203 gnd.n4824 gnd.n4823 585
R9204 gnd.n4823 gnd.n4756 585
R9205 gnd.n5774 gnd.n5773 585
R9206 gnd.n5775 gnd.n1350 585
R9207 gnd.n5627 gnd.n1347 585
R9208 gnd.n5630 gnd.n5629 585
R9209 gnd.n5640 gnd.n5626 585
R9210 gnd.n5641 gnd.n5624 585
R9211 gnd.n5623 gnd.n5614 585
R9212 gnd.n5648 gnd.n5613 585
R9213 gnd.n5649 gnd.n5612 585
R9214 gnd.n5610 gnd.n5604 585
R9215 gnd.n5656 gnd.n5603 585
R9216 gnd.n5657 gnd.n5601 585
R9217 gnd.n5600 gnd.n5591 585
R9218 gnd.n5664 gnd.n5590 585
R9219 gnd.n5665 gnd.n5589 585
R9220 gnd.n5587 gnd.n5579 585
R9221 gnd.n5672 gnd.n5578 585
R9222 gnd.n5673 gnd.n5576 585
R9223 gnd.n5575 gnd.n5573 585
R9224 gnd.n5575 gnd.n1364 585
R9225 gnd.n5772 gnd.n1353 585
R9226 gnd.n5772 gnd.n5771 585
R9227 gnd.n5388 gnd.n1352 585
R9228 gnd.n5694 gnd.n1352 585
R9229 gnd.n5391 gnd.n5387 585
R9230 gnd.n5387 gnd.n5386 585
R9231 gnd.n5392 gnd.n1657 585
R9232 gnd.n5567 gnd.n1657 585
R9233 gnd.n5393 gnd.n5385 585
R9234 gnd.n5385 gnd.n5384 585
R9235 gnd.n1829 gnd.n1667 585
R9236 gnd.n5557 gnd.n1667 585
R9237 gnd.n5397 gnd.n1828 585
R9238 gnd.n5373 gnd.n1828 585
R9239 gnd.n5398 gnd.n1676 585
R9240 gnd.n5549 gnd.n1676 585
R9241 gnd.n5399 gnd.n1827 585
R9242 gnd.n5328 gnd.n1827 585
R9243 gnd.n1825 gnd.n1683 585
R9244 gnd.n5541 gnd.n1683 585
R9245 gnd.n5403 gnd.n1824 585
R9246 gnd.n5334 gnd.n1824 585
R9247 gnd.n5404 gnd.n1692 585
R9248 gnd.n5533 gnd.n1692 585
R9249 gnd.n5405 gnd.n1823 585
R9250 gnd.n5320 gnd.n1823 585
R9251 gnd.n1821 gnd.n1701 585
R9252 gnd.n5525 gnd.n1701 585
R9253 gnd.n5409 gnd.n1820 585
R9254 gnd.n5316 gnd.n1820 585
R9255 gnd.n5410 gnd.n1710 585
R9256 gnd.n5517 gnd.n1710 585
R9257 gnd.n5411 gnd.n1819 585
R9258 gnd.n5289 gnd.n1819 585
R9259 gnd.n1817 gnd.n1717 585
R9260 gnd.n5509 gnd.n1717 585
R9261 gnd.n5415 gnd.n1816 585
R9262 gnd.n5295 gnd.n1816 585
R9263 gnd.n5416 gnd.n1726 585
R9264 gnd.n5501 gnd.n1726 585
R9265 gnd.n5417 gnd.n1815 585
R9266 gnd.n5280 gnd.n1815 585
R9267 gnd.n1813 gnd.n1735 585
R9268 gnd.n5493 gnd.n1735 585
R9269 gnd.n5421 gnd.n1812 585
R9270 gnd.n5276 gnd.n1812 585
R9271 gnd.n5422 gnd.n1744 585
R9272 gnd.n5485 gnd.n1744 585
R9273 gnd.n5423 gnd.n1811 585
R9274 gnd.n5249 gnd.n1811 585
R9275 gnd.n1808 gnd.n1751 585
R9276 gnd.n5477 gnd.n1751 585
R9277 gnd.n5428 gnd.n5427 585
R9278 gnd.n5429 gnd.n5428 585
R9279 gnd.n1807 gnd.n1760 585
R9280 gnd.n5469 gnd.n1760 585
R9281 gnd.n5240 gnd.n5239 585
R9282 gnd.n5241 gnd.n5240 585
R9283 gnd.n1857 gnd.n1797 585
R9284 gnd.n5441 gnd.n1797 585
R9285 gnd.n5235 gnd.n5234 585
R9286 gnd.n5234 gnd.n5233 585
R9287 gnd.n1859 gnd.n1790 585
R9288 gnd.n5447 gnd.n1790 585
R9289 gnd.n5210 gnd.n5208 585
R9290 gnd.n5208 gnd.n1786 585
R9291 gnd.n5211 gnd.n1785 585
R9292 gnd.n5455 gnd.n1785 585
R9293 gnd.n5213 gnd.n5212 585
R9294 gnd.n5212 gnd.n1775 585
R9295 gnd.n5214 gnd.n1774 585
R9296 gnd.n5461 gnd.n1774 585
R9297 gnd.n5216 gnd.n5215 585
R9298 gnd.n5217 gnd.n5216 585
R9299 gnd.n1869 gnd.n1868 585
R9300 gnd.n1868 gnd.n1867 585
R9301 gnd.n5201 gnd.n5200 585
R9302 gnd.n5200 gnd.n5199 585
R9303 gnd.n1872 gnd.n1871 585
R9304 gnd.n5184 gnd.n1872 585
R9305 gnd.n5169 gnd.n5168 585
R9306 gnd.n5168 gnd.n1884 585
R9307 gnd.n5170 gnd.n1883 585
R9308 gnd.n5190 gnd.n1883 585
R9309 gnd.n5172 gnd.n5171 585
R9310 gnd.n5173 gnd.n5172 585
R9311 gnd.n1904 gnd.n1903 585
R9312 gnd.n1903 gnd.n1902 585
R9313 gnd.n5162 gnd.n5161 585
R9314 gnd.n5161 gnd.n5160 585
R9315 gnd.n1907 gnd.n1906 585
R9316 gnd.n1908 gnd.n1907 585
R9317 gnd.n4845 gnd.n1918 585
R9318 gnd.n5150 gnd.n1918 585
R9319 gnd.n4847 gnd.n4846 585
R9320 gnd.n4846 gnd.n1928 585
R9321 gnd.n4848 gnd.n1927 585
R9322 gnd.n5134 gnd.n1927 585
R9323 gnd.n4850 gnd.n4849 585
R9324 gnd.n4849 gnd.n1925 585
R9325 gnd.n4851 gnd.n1936 585
R9326 gnd.n5126 gnd.n1936 585
R9327 gnd.n4853 gnd.n4852 585
R9328 gnd.n4852 gnd.n1934 585
R9329 gnd.n4854 gnd.n1944 585
R9330 gnd.n5118 gnd.n1944 585
R9331 gnd.n4856 gnd.n4855 585
R9332 gnd.n4855 gnd.n1942 585
R9333 gnd.n4857 gnd.n1951 585
R9334 gnd.n5110 gnd.n1951 585
R9335 gnd.n4859 gnd.n4858 585
R9336 gnd.n4858 gnd.n1960 585
R9337 gnd.n4860 gnd.n1959 585
R9338 gnd.n5102 gnd.n1959 585
R9339 gnd.n4862 gnd.n4861 585
R9340 gnd.n4861 gnd.n1957 585
R9341 gnd.n4863 gnd.n1968 585
R9342 gnd.n5094 gnd.n1968 585
R9343 gnd.n4865 gnd.n4864 585
R9344 gnd.n4864 gnd.n1966 585
R9345 gnd.n4866 gnd.n1976 585
R9346 gnd.n5086 gnd.n1976 585
R9347 gnd.n4868 gnd.n4867 585
R9348 gnd.n4867 gnd.n1974 585
R9349 gnd.n4869 gnd.n1983 585
R9350 gnd.n5078 gnd.n1983 585
R9351 gnd.n4871 gnd.n4870 585
R9352 gnd.n4872 gnd.n4871 585
R9353 gnd.n4759 gnd.n4758 585
R9354 gnd.n5070 gnd.n4758 585
R9355 gnd.n7477 gnd.n125 585
R9356 gnd.n7573 gnd.n125 585
R9357 gnd.n7478 gnd.n7415 585
R9358 gnd.n7415 gnd.n122 585
R9359 gnd.n7479 gnd.n203 585
R9360 gnd.n7493 gnd.n203 585
R9361 gnd.n215 gnd.n213 585
R9362 gnd.n213 gnd.n202 585
R9363 gnd.n7484 gnd.n7483 585
R9364 gnd.n7485 gnd.n7484 585
R9365 gnd.n214 gnd.n212 585
R9366 gnd.n212 gnd.n209 585
R9367 gnd.n7411 gnd.n7410 585
R9368 gnd.n7410 gnd.n7409 585
R9369 gnd.n218 gnd.n217 585
R9370 gnd.n228 gnd.n218 585
R9371 gnd.n7400 gnd.n7399 585
R9372 gnd.n7401 gnd.n7400 585
R9373 gnd.n230 gnd.n229 585
R9374 gnd.n229 gnd.n225 585
R9375 gnd.n7395 gnd.n7394 585
R9376 gnd.n7394 gnd.n7393 585
R9377 gnd.n233 gnd.n232 585
R9378 gnd.n234 gnd.n233 585
R9379 gnd.n7384 gnd.n7383 585
R9380 gnd.n7385 gnd.n7384 585
R9381 gnd.n245 gnd.n244 585
R9382 gnd.n250 gnd.n244 585
R9383 gnd.n7379 gnd.n7378 585
R9384 gnd.n7378 gnd.n7377 585
R9385 gnd.n248 gnd.n247 585
R9386 gnd.n259 gnd.n248 585
R9387 gnd.n7368 gnd.n7367 585
R9388 gnd.n7369 gnd.n7368 585
R9389 gnd.n261 gnd.n260 585
R9390 gnd.n260 gnd.n256 585
R9391 gnd.n7363 gnd.n7362 585
R9392 gnd.n7362 gnd.n7361 585
R9393 gnd.n264 gnd.n263 585
R9394 gnd.n265 gnd.n264 585
R9395 gnd.n7352 gnd.n7351 585
R9396 gnd.n7353 gnd.n7352 585
R9397 gnd.n275 gnd.n274 585
R9398 gnd.n280 gnd.n274 585
R9399 gnd.n7347 gnd.n7346 585
R9400 gnd.n7346 gnd.n7345 585
R9401 gnd.n278 gnd.n277 585
R9402 gnd.n289 gnd.n278 585
R9403 gnd.n7336 gnd.n7335 585
R9404 gnd.n7337 gnd.n7336 585
R9405 gnd.n291 gnd.n290 585
R9406 gnd.n290 gnd.n286 585
R9407 gnd.n7331 gnd.n7330 585
R9408 gnd.n7330 gnd.n7329 585
R9409 gnd.n294 gnd.n293 585
R9410 gnd.n295 gnd.n294 585
R9411 gnd.n7307 gnd.n7306 585
R9412 gnd.n7306 gnd.n7305 585
R9413 gnd.n7308 gnd.n323 585
R9414 gnd.n7301 gnd.n323 585
R9415 gnd.n329 gnd.n321 585
R9416 gnd.n330 gnd.n329 585
R9417 gnd.n7312 gnd.n320 585
R9418 gnd.n7228 gnd.n320 585
R9419 gnd.n7313 gnd.n319 585
R9420 gnd.n336 gnd.n319 585
R9421 gnd.n7314 gnd.n318 585
R9422 gnd.n7222 gnd.n318 585
R9423 gnd.n315 gnd.n313 585
R9424 gnd.n7202 gnd.n313 585
R9425 gnd.n7319 gnd.n7318 585
R9426 gnd.n7320 gnd.n7319 585
R9427 gnd.n314 gnd.n312 585
R9428 gnd.n7211 gnd.n312 585
R9429 gnd.n7173 gnd.n7171 585
R9430 gnd.n7171 gnd.n349 585
R9431 gnd.n7174 gnd.n362 585
R9432 gnd.n7190 gnd.n362 585
R9433 gnd.n7175 gnd.n7170 585
R9434 gnd.n7170 gnd.n7169 585
R9435 gnd.n376 gnd.n374 585
R9436 gnd.n6930 gnd.n374 585
R9437 gnd.n7180 gnd.n7179 585
R9438 gnd.n7181 gnd.n7180 585
R9439 gnd.n375 gnd.n373 585
R9440 gnd.n7159 gnd.n373 585
R9441 gnd.n7124 gnd.n395 585
R9442 gnd.n7138 gnd.n395 585
R9443 gnd.n408 gnd.n406 585
R9444 gnd.n6938 gnd.n406 585
R9445 gnd.n7129 gnd.n7128 585
R9446 gnd.n7130 gnd.n7129 585
R9447 gnd.n407 gnd.n405 585
R9448 gnd.n6917 gnd.n405 585
R9449 gnd.n7121 gnd.n7120 585
R9450 gnd.n7120 gnd.n7119 585
R9451 gnd.n411 gnd.n410 585
R9452 gnd.n6898 gnd.n411 585
R9453 gnd.n7110 gnd.n7109 585
R9454 gnd.n7111 gnd.n7110 585
R9455 gnd.n424 gnd.n423 585
R9456 gnd.n6904 gnd.n423 585
R9457 gnd.n7105 gnd.n7104 585
R9458 gnd.n7104 gnd.n7103 585
R9459 gnd.n427 gnd.n426 585
R9460 gnd.n6890 gnd.n427 585
R9461 gnd.n7094 gnd.n7093 585
R9462 gnd.n7095 gnd.n7094 585
R9463 gnd.n442 gnd.n441 585
R9464 gnd.n6886 gnd.n441 585
R9465 gnd.n7089 gnd.n7088 585
R9466 gnd.n7088 gnd.n7087 585
R9467 gnd.n445 gnd.n444 585
R9468 gnd.n6859 gnd.n445 585
R9469 gnd.n7078 gnd.n7077 585
R9470 gnd.n7079 gnd.n7078 585
R9471 gnd.n458 gnd.n457 585
R9472 gnd.n6865 gnd.n457 585
R9473 gnd.n7073 gnd.n7072 585
R9474 gnd.n7072 gnd.n7071 585
R9475 gnd.n461 gnd.n460 585
R9476 gnd.n6850 gnd.n461 585
R9477 gnd.n7062 gnd.n7061 585
R9478 gnd.n7063 gnd.n7062 585
R9479 gnd.n476 gnd.n475 585
R9480 gnd.n6846 gnd.n475 585
R9481 gnd.n7057 gnd.n7056 585
R9482 gnd.n7056 gnd.n7055 585
R9483 gnd.n479 gnd.n478 585
R9484 gnd.n6974 gnd.n479 585
R9485 gnd.n6622 gnd.n6621 585
R9486 gnd.n6624 gnd.n6623 585
R9487 gnd.n6754 gnd.n6625 585
R9488 gnd.n6753 gnd.n6626 585
R9489 gnd.n6628 gnd.n6627 585
R9490 gnd.n6746 gnd.n6636 585
R9491 gnd.n6745 gnd.n6637 585
R9492 gnd.n6644 gnd.n6638 585
R9493 gnd.n6738 gnd.n6645 585
R9494 gnd.n6737 gnd.n6646 585
R9495 gnd.n6648 gnd.n6647 585
R9496 gnd.n6730 gnd.n6656 585
R9497 gnd.n6729 gnd.n6657 585
R9498 gnd.n6664 gnd.n6658 585
R9499 gnd.n6722 gnd.n6665 585
R9500 gnd.n6721 gnd.n6666 585
R9501 gnd.n6668 gnd.n6667 585
R9502 gnd.n6714 gnd.n6711 585
R9503 gnd.n6710 gnd.n517 585
R9504 gnd.n7046 gnd.n517 585
R9505 gnd.n7576 gnd.n7575 585
R9506 gnd.n7448 gnd.n120 585
R9507 gnd.n7450 gnd.n7449 585
R9508 gnd.n7446 gnd.n7445 585
R9509 gnd.n7454 gnd.n7444 585
R9510 gnd.n7455 gnd.n7442 585
R9511 gnd.n7456 gnd.n7441 585
R9512 gnd.n7439 gnd.n7437 585
R9513 gnd.n7460 gnd.n7436 585
R9514 gnd.n7461 gnd.n7434 585
R9515 gnd.n7462 gnd.n7433 585
R9516 gnd.n7431 gnd.n7429 585
R9517 gnd.n7466 gnd.n7428 585
R9518 gnd.n7467 gnd.n7426 585
R9519 gnd.n7468 gnd.n7425 585
R9520 gnd.n7423 gnd.n7421 585
R9521 gnd.n7472 gnd.n7420 585
R9522 gnd.n7473 gnd.n7418 585
R9523 gnd.n7474 gnd.n7417 585
R9524 gnd.n7417 gnd.n124 585
R9525 gnd.n7574 gnd.n116 585
R9526 gnd.n7574 gnd.n7573 585
R9527 gnd.n7580 gnd.n115 585
R9528 gnd.n122 gnd.n115 585
R9529 gnd.n7581 gnd.n114 585
R9530 gnd.n7493 gnd.n114 585
R9531 gnd.n7582 gnd.n113 585
R9532 gnd.n202 gnd.n113 585
R9533 gnd.n211 gnd.n111 585
R9534 gnd.n7485 gnd.n211 585
R9535 gnd.n7586 gnd.n110 585
R9536 gnd.n209 gnd.n110 585
R9537 gnd.n7587 gnd.n109 585
R9538 gnd.n7409 gnd.n109 585
R9539 gnd.n7588 gnd.n108 585
R9540 gnd.n228 gnd.n108 585
R9541 gnd.n227 gnd.n106 585
R9542 gnd.n7401 gnd.n227 585
R9543 gnd.n7592 gnd.n105 585
R9544 gnd.n225 gnd.n105 585
R9545 gnd.n7593 gnd.n104 585
R9546 gnd.n7393 gnd.n104 585
R9547 gnd.n7594 gnd.n103 585
R9548 gnd.n234 gnd.n103 585
R9549 gnd.n243 gnd.n101 585
R9550 gnd.n7385 gnd.n243 585
R9551 gnd.n7598 gnd.n100 585
R9552 gnd.n250 gnd.n100 585
R9553 gnd.n7599 gnd.n99 585
R9554 gnd.n7377 gnd.n99 585
R9555 gnd.n7600 gnd.n98 585
R9556 gnd.n259 gnd.n98 585
R9557 gnd.n258 gnd.n96 585
R9558 gnd.n7369 gnd.n258 585
R9559 gnd.n7604 gnd.n95 585
R9560 gnd.n256 gnd.n95 585
R9561 gnd.n7605 gnd.n94 585
R9562 gnd.n7361 gnd.n94 585
R9563 gnd.n7606 gnd.n93 585
R9564 gnd.n265 gnd.n93 585
R9565 gnd.n273 gnd.n91 585
R9566 gnd.n7353 gnd.n273 585
R9567 gnd.n7610 gnd.n90 585
R9568 gnd.n280 gnd.n90 585
R9569 gnd.n7611 gnd.n89 585
R9570 gnd.n7345 gnd.n89 585
R9571 gnd.n7612 gnd.n88 585
R9572 gnd.n289 gnd.n88 585
R9573 gnd.n288 gnd.n86 585
R9574 gnd.n7337 gnd.n288 585
R9575 gnd.n7616 gnd.n85 585
R9576 gnd.n286 gnd.n85 585
R9577 gnd.n7617 gnd.n84 585
R9578 gnd.n7329 gnd.n84 585
R9579 gnd.n7618 gnd.n83 585
R9580 gnd.n295 gnd.n83 585
R9581 gnd.n325 gnd.n81 585
R9582 gnd.n7305 gnd.n325 585
R9583 gnd.n7622 gnd.n80 585
R9584 gnd.n7301 gnd.n80 585
R9585 gnd.n7623 gnd.n79 585
R9586 gnd.n330 gnd.n79 585
R9587 gnd.n7624 gnd.n78 585
R9588 gnd.n7228 gnd.n78 585
R9589 gnd.n340 gnd.n76 585
R9590 gnd.n340 gnd.n336 585
R9591 gnd.n7204 gnd.n341 585
R9592 gnd.n7222 gnd.n341 585
R9593 gnd.n7205 gnd.n7203 585
R9594 gnd.n7203 gnd.n7202 585
R9595 gnd.n353 gnd.n310 585
R9596 gnd.n7320 gnd.n310 585
R9597 gnd.n7210 gnd.n7209 585
R9598 gnd.n7211 gnd.n7210 585
R9599 gnd.n352 gnd.n351 585
R9600 gnd.n351 gnd.n349 585
R9601 gnd.n382 gnd.n360 585
R9602 gnd.n7190 gnd.n360 585
R9603 gnd.n7168 gnd.n7167 585
R9604 gnd.n7169 gnd.n7168 585
R9605 gnd.n381 gnd.n380 585
R9606 gnd.n6930 gnd.n380 585
R9607 gnd.n7162 gnd.n371 585
R9608 gnd.n7181 gnd.n371 585
R9609 gnd.n7161 gnd.n7160 585
R9610 gnd.n7160 gnd.n7159 585
R9611 gnd.n385 gnd.n384 585
R9612 gnd.n7138 gnd.n385 585
R9613 gnd.n6942 gnd.n6939 585
R9614 gnd.n6939 gnd.n6938 585
R9615 gnd.n6943 gnd.n403 585
R9616 gnd.n7130 gnd.n403 585
R9617 gnd.n6944 gnd.n584 585
R9618 gnd.n6917 gnd.n584 585
R9619 gnd.n582 gnd.n414 585
R9620 gnd.n7119 gnd.n414 585
R9621 gnd.n6948 gnd.n581 585
R9622 gnd.n6898 gnd.n581 585
R9623 gnd.n6949 gnd.n421 585
R9624 gnd.n7111 gnd.n421 585
R9625 gnd.n6950 gnd.n580 585
R9626 gnd.n6904 gnd.n580 585
R9627 gnd.n578 gnd.n430 585
R9628 gnd.n7103 gnd.n430 585
R9629 gnd.n6954 gnd.n577 585
R9630 gnd.n6890 gnd.n577 585
R9631 gnd.n6955 gnd.n439 585
R9632 gnd.n7095 gnd.n439 585
R9633 gnd.n6956 gnd.n576 585
R9634 gnd.n6886 gnd.n576 585
R9635 gnd.n574 gnd.n448 585
R9636 gnd.n7087 gnd.n448 585
R9637 gnd.n6960 gnd.n573 585
R9638 gnd.n6859 gnd.n573 585
R9639 gnd.n6961 gnd.n455 585
R9640 gnd.n7079 gnd.n455 585
R9641 gnd.n6962 gnd.n572 585
R9642 gnd.n6865 gnd.n572 585
R9643 gnd.n570 gnd.n464 585
R9644 gnd.n7071 gnd.n464 585
R9645 gnd.n6966 gnd.n569 585
R9646 gnd.n6850 gnd.n569 585
R9647 gnd.n6967 gnd.n473 585
R9648 gnd.n7063 gnd.n473 585
R9649 gnd.n6968 gnd.n568 585
R9650 gnd.n6846 gnd.n568 585
R9651 gnd.n565 gnd.n482 585
R9652 gnd.n7055 gnd.n482 585
R9653 gnd.n6973 gnd.n6972 585
R9654 gnd.n6974 gnd.n6973 585
R9655 gnd.n4663 gnd.n4662 585
R9656 gnd.n4664 gnd.n4663 585
R9657 gnd.n3357 gnd.n3356 585
R9658 gnd.n3364 gnd.n3356 585
R9659 gnd.n4645 gnd.n4644 585
R9660 gnd.n4646 gnd.n4645 585
R9661 gnd.n3375 gnd.n3374 585
R9662 gnd.n3374 gnd.n3370 585
R9663 gnd.n4635 gnd.n4634 585
R9664 gnd.n4636 gnd.n4635 585
R9665 gnd.n3383 gnd.n3382 585
R9666 gnd.n3388 gnd.n3382 585
R9667 gnd.n4357 gnd.n3400 585
R9668 gnd.n3400 gnd.n3387 585
R9669 gnd.n4359 gnd.n4358 585
R9670 gnd.n4360 gnd.n4359 585
R9671 gnd.n3401 gnd.n3399 585
R9672 gnd.n3399 gnd.n3395 585
R9673 gnd.n4348 gnd.n4347 585
R9674 gnd.n4349 gnd.n4348 585
R9675 gnd.n3408 gnd.n3407 585
R9676 gnd.n3413 gnd.n3407 585
R9677 gnd.n4326 gnd.n3426 585
R9678 gnd.n3426 gnd.n3412 585
R9679 gnd.n4328 gnd.n4327 585
R9680 gnd.n4329 gnd.n4328 585
R9681 gnd.n3427 gnd.n3425 585
R9682 gnd.n3425 gnd.n3421 585
R9683 gnd.n4317 gnd.n4316 585
R9684 gnd.n4318 gnd.n4317 585
R9685 gnd.n3434 gnd.n3433 585
R9686 gnd.n3438 gnd.n3433 585
R9687 gnd.n4295 gnd.n3450 585
R9688 gnd.n3588 gnd.n3450 585
R9689 gnd.n4297 gnd.n4296 585
R9690 gnd.n4298 gnd.n4297 585
R9691 gnd.n3451 gnd.n3449 585
R9692 gnd.n3449 gnd.n3446 585
R9693 gnd.n4286 gnd.n4285 585
R9694 gnd.n4287 gnd.n4286 585
R9695 gnd.n3458 gnd.n3457 585
R9696 gnd.n3463 gnd.n3457 585
R9697 gnd.n4264 gnd.n3476 585
R9698 gnd.n3476 gnd.n3462 585
R9699 gnd.n4266 gnd.n4265 585
R9700 gnd.n4267 gnd.n4266 585
R9701 gnd.n3477 gnd.n3475 585
R9702 gnd.n3475 gnd.n3471 585
R9703 gnd.n4255 gnd.n4254 585
R9704 gnd.n4256 gnd.n4255 585
R9705 gnd.n3485 gnd.n3484 585
R9706 gnd.n3490 gnd.n3484 585
R9707 gnd.n4233 gnd.n3502 585
R9708 gnd.n3502 gnd.n3489 585
R9709 gnd.n4235 gnd.n4234 585
R9710 gnd.n4236 gnd.n4235 585
R9711 gnd.n3503 gnd.n3501 585
R9712 gnd.n3501 gnd.n3497 585
R9713 gnd.n4224 gnd.n4223 585
R9714 gnd.n4225 gnd.n4224 585
R9715 gnd.n3510 gnd.n3509 585
R9716 gnd.n3613 gnd.n3509 585
R9717 gnd.n4202 gnd.n3525 585
R9718 gnd.n3525 gnd.n3514 585
R9719 gnd.n4204 gnd.n4203 585
R9720 gnd.n4205 gnd.n4204 585
R9721 gnd.n3526 gnd.n3524 585
R9722 gnd.n4194 gnd.n3524 585
R9723 gnd.n3694 gnd.n3693 585
R9724 gnd.n3694 gnd.n3531 585
R9725 gnd.n4181 gnd.n4180 585
R9726 gnd.n4180 gnd.n4179 585
R9727 gnd.n4182 gnd.n3686 585
R9728 gnd.n4159 gnd.n3686 585
R9729 gnd.n4184 gnd.n4183 585
R9730 gnd.n4185 gnd.n4184 585
R9731 gnd.n3687 gnd.n3685 585
R9732 gnd.n4167 gnd.n3685 585
R9733 gnd.n4151 gnd.n4150 585
R9734 gnd.n4150 gnd.n3704 585
R9735 gnd.n4149 gnd.n3709 585
R9736 gnd.n4149 gnd.n4148 585
R9737 gnd.n4134 gnd.n3710 585
R9738 gnd.n3718 gnd.n3710 585
R9739 gnd.n4136 gnd.n4135 585
R9740 gnd.n4137 gnd.n4136 585
R9741 gnd.n3721 gnd.n3720 585
R9742 gnd.n3728 gnd.n3720 585
R9743 gnd.n4109 gnd.n4108 585
R9744 gnd.n4110 gnd.n4109 585
R9745 gnd.n3740 gnd.n3739 585
R9746 gnd.n3739 gnd.n3735 585
R9747 gnd.n4099 gnd.n4098 585
R9748 gnd.n4100 gnd.n4099 585
R9749 gnd.n3750 gnd.n3749 585
R9750 gnd.n3755 gnd.n3749 585
R9751 gnd.n4077 gnd.n3768 585
R9752 gnd.n3768 gnd.n3754 585
R9753 gnd.n4079 gnd.n4078 585
R9754 gnd.n4080 gnd.n4079 585
R9755 gnd.n3769 gnd.n3767 585
R9756 gnd.n3767 gnd.n3763 585
R9757 gnd.n4068 gnd.n4067 585
R9758 gnd.n4069 gnd.n4068 585
R9759 gnd.n3776 gnd.n3775 585
R9760 gnd.n3780 gnd.n3775 585
R9761 gnd.n4045 gnd.n3797 585
R9762 gnd.n3797 gnd.n3779 585
R9763 gnd.n4047 gnd.n4046 585
R9764 gnd.n4048 gnd.n4047 585
R9765 gnd.n3798 gnd.n3796 585
R9766 gnd.n3796 gnd.n3787 585
R9767 gnd.n4040 gnd.n4039 585
R9768 gnd.n4039 gnd.n4038 585
R9769 gnd.n3845 gnd.n3844 585
R9770 gnd.n3846 gnd.n3845 585
R9771 gnd.n3999 gnd.n3998 585
R9772 gnd.n4000 gnd.n3999 585
R9773 gnd.n3855 gnd.n3854 585
R9774 gnd.n3854 gnd.n3853 585
R9775 gnd.n3994 gnd.n3993 585
R9776 gnd.n3993 gnd.n3992 585
R9777 gnd.n3858 gnd.n3857 585
R9778 gnd.n3859 gnd.n3858 585
R9779 gnd.n3983 gnd.n3982 585
R9780 gnd.n3984 gnd.n3983 585
R9781 gnd.n3866 gnd.n3865 585
R9782 gnd.n3975 gnd.n3865 585
R9783 gnd.n3978 gnd.n3977 585
R9784 gnd.n3977 gnd.n3976 585
R9785 gnd.n3869 gnd.n3868 585
R9786 gnd.n3870 gnd.n3869 585
R9787 gnd.n3964 gnd.n3963 585
R9788 gnd.n3962 gnd.n3888 585
R9789 gnd.n3961 gnd.n3887 585
R9790 gnd.n3966 gnd.n3887 585
R9791 gnd.n3960 gnd.n3959 585
R9792 gnd.n3958 gnd.n3957 585
R9793 gnd.n3956 gnd.n3955 585
R9794 gnd.n3954 gnd.n3953 585
R9795 gnd.n3952 gnd.n3951 585
R9796 gnd.n3950 gnd.n3949 585
R9797 gnd.n3948 gnd.n3947 585
R9798 gnd.n3946 gnd.n3945 585
R9799 gnd.n3944 gnd.n3943 585
R9800 gnd.n3942 gnd.n3941 585
R9801 gnd.n3940 gnd.n3939 585
R9802 gnd.n3938 gnd.n3937 585
R9803 gnd.n3936 gnd.n3935 585
R9804 gnd.n3934 gnd.n3933 585
R9805 gnd.n3932 gnd.n3931 585
R9806 gnd.n3930 gnd.n3929 585
R9807 gnd.n3928 gnd.n3927 585
R9808 gnd.n3926 gnd.n3925 585
R9809 gnd.n3924 gnd.n3923 585
R9810 gnd.n3922 gnd.n3921 585
R9811 gnd.n3920 gnd.n3919 585
R9812 gnd.n3918 gnd.n3917 585
R9813 gnd.n3875 gnd.n3874 585
R9814 gnd.n3969 gnd.n3968 585
R9815 gnd.n4667 gnd.n4666 585
R9816 gnd.n4669 gnd.n4668 585
R9817 gnd.n4671 gnd.n4670 585
R9818 gnd.n4673 gnd.n4672 585
R9819 gnd.n4675 gnd.n4674 585
R9820 gnd.n4677 gnd.n4676 585
R9821 gnd.n4679 gnd.n4678 585
R9822 gnd.n4681 gnd.n4680 585
R9823 gnd.n4683 gnd.n4682 585
R9824 gnd.n4685 gnd.n4684 585
R9825 gnd.n4687 gnd.n4686 585
R9826 gnd.n4689 gnd.n4688 585
R9827 gnd.n4691 gnd.n4690 585
R9828 gnd.n4693 gnd.n4692 585
R9829 gnd.n4695 gnd.n4694 585
R9830 gnd.n4697 gnd.n4696 585
R9831 gnd.n4699 gnd.n4698 585
R9832 gnd.n4701 gnd.n4700 585
R9833 gnd.n4703 gnd.n4702 585
R9834 gnd.n4705 gnd.n4704 585
R9835 gnd.n4707 gnd.n4706 585
R9836 gnd.n4709 gnd.n4708 585
R9837 gnd.n4711 gnd.n4710 585
R9838 gnd.n4713 gnd.n4712 585
R9839 gnd.n4715 gnd.n4714 585
R9840 gnd.n4716 gnd.n2031 585
R9841 gnd.n4717 gnd.n1989 585
R9842 gnd.n4755 gnd.n1989 585
R9843 gnd.n4665 gnd.n2061 585
R9844 gnd.n4665 gnd.n4664 585
R9845 gnd.n3564 gnd.n2060 585
R9846 gnd.n3364 gnd.n2060 585
R9847 gnd.n3565 gnd.n3372 585
R9848 gnd.n4646 gnd.n3372 585
R9849 gnd.n3567 gnd.n3566 585
R9850 gnd.n3566 gnd.n3370 585
R9851 gnd.n3568 gnd.n3381 585
R9852 gnd.n4636 gnd.n3381 585
R9853 gnd.n3570 gnd.n3569 585
R9854 gnd.n3570 gnd.n3388 585
R9855 gnd.n3572 gnd.n3571 585
R9856 gnd.n3571 gnd.n3387 585
R9857 gnd.n3573 gnd.n3397 585
R9858 gnd.n4360 gnd.n3397 585
R9859 gnd.n3575 gnd.n3574 585
R9860 gnd.n3574 gnd.n3395 585
R9861 gnd.n3576 gnd.n3406 585
R9862 gnd.n4349 gnd.n3406 585
R9863 gnd.n3578 gnd.n3577 585
R9864 gnd.n3578 gnd.n3413 585
R9865 gnd.n3580 gnd.n3579 585
R9866 gnd.n3579 gnd.n3412 585
R9867 gnd.n3581 gnd.n3423 585
R9868 gnd.n4329 gnd.n3423 585
R9869 gnd.n3583 gnd.n3582 585
R9870 gnd.n3582 gnd.n3421 585
R9871 gnd.n3584 gnd.n3432 585
R9872 gnd.n4318 gnd.n3432 585
R9873 gnd.n3586 gnd.n3585 585
R9874 gnd.n3586 gnd.n3438 585
R9875 gnd.n3590 gnd.n3589 585
R9876 gnd.n3589 gnd.n3588 585
R9877 gnd.n3591 gnd.n3448 585
R9878 gnd.n4298 gnd.n3448 585
R9879 gnd.n3593 gnd.n3592 585
R9880 gnd.n3592 gnd.n3446 585
R9881 gnd.n3594 gnd.n3456 585
R9882 gnd.n4287 gnd.n3456 585
R9883 gnd.n3596 gnd.n3595 585
R9884 gnd.n3596 gnd.n3463 585
R9885 gnd.n3598 gnd.n3597 585
R9886 gnd.n3597 gnd.n3462 585
R9887 gnd.n3599 gnd.n3473 585
R9888 gnd.n4267 gnd.n3473 585
R9889 gnd.n3601 gnd.n3600 585
R9890 gnd.n3600 gnd.n3471 585
R9891 gnd.n3602 gnd.n3483 585
R9892 gnd.n4256 gnd.n3483 585
R9893 gnd.n3604 gnd.n3603 585
R9894 gnd.n3604 gnd.n3490 585
R9895 gnd.n3606 gnd.n3605 585
R9896 gnd.n3605 gnd.n3489 585
R9897 gnd.n3607 gnd.n3499 585
R9898 gnd.n4236 gnd.n3499 585
R9899 gnd.n3609 gnd.n3608 585
R9900 gnd.n3608 gnd.n3497 585
R9901 gnd.n3610 gnd.n3508 585
R9902 gnd.n4225 gnd.n3508 585
R9903 gnd.n3615 gnd.n3614 585
R9904 gnd.n3614 gnd.n3613 585
R9905 gnd.n3611 gnd.n3534 585
R9906 gnd.n3611 gnd.n3514 585
R9907 gnd.n4191 gnd.n3522 585
R9908 gnd.n4205 gnd.n3522 585
R9909 gnd.n4193 gnd.n4192 585
R9910 gnd.n4194 gnd.n4193 585
R9911 gnd.n3695 gnd.n3532 585
R9912 gnd.n3532 gnd.n3531 585
R9913 gnd.n3697 gnd.n3696 585
R9914 gnd.n4179 gnd.n3697 585
R9915 gnd.n3682 gnd.n3680 585
R9916 gnd.n4159 gnd.n3682 585
R9917 gnd.n4187 gnd.n4186 585
R9918 gnd.n4186 gnd.n4185 585
R9919 gnd.n3681 gnd.n3679 585
R9920 gnd.n4167 gnd.n3681 585
R9921 gnd.n4144 gnd.n3713 585
R9922 gnd.n3713 gnd.n3704 585
R9923 gnd.n4146 gnd.n4145 585
R9924 gnd.n4148 gnd.n4146 585
R9925 gnd.n3714 gnd.n3712 585
R9926 gnd.n3718 gnd.n3712 585
R9927 gnd.n4139 gnd.n4138 585
R9928 gnd.n4138 gnd.n4137 585
R9929 gnd.n3717 gnd.n3716 585
R9930 gnd.n3728 gnd.n3717 585
R9931 gnd.n4018 gnd.n3737 585
R9932 gnd.n4110 gnd.n3737 585
R9933 gnd.n4020 gnd.n4019 585
R9934 gnd.n4019 gnd.n3735 585
R9935 gnd.n4021 gnd.n3748 585
R9936 gnd.n4100 gnd.n3748 585
R9937 gnd.n4023 gnd.n4022 585
R9938 gnd.n4023 gnd.n3755 585
R9939 gnd.n4025 gnd.n4024 585
R9940 gnd.n4024 gnd.n3754 585
R9941 gnd.n4026 gnd.n3765 585
R9942 gnd.n4080 gnd.n3765 585
R9943 gnd.n4028 gnd.n4027 585
R9944 gnd.n4027 gnd.n3763 585
R9945 gnd.n4029 gnd.n3774 585
R9946 gnd.n4069 gnd.n3774 585
R9947 gnd.n4031 gnd.n4030 585
R9948 gnd.n4031 gnd.n3780 585
R9949 gnd.n4033 gnd.n4032 585
R9950 gnd.n4032 gnd.n3779 585
R9951 gnd.n4034 gnd.n3795 585
R9952 gnd.n4048 gnd.n3795 585
R9953 gnd.n4035 gnd.n3848 585
R9954 gnd.n3848 gnd.n3787 585
R9955 gnd.n4037 gnd.n4036 585
R9956 gnd.n4038 gnd.n4037 585
R9957 gnd.n3849 gnd.n3847 585
R9958 gnd.n3847 gnd.n3846 585
R9959 gnd.n4002 gnd.n4001 585
R9960 gnd.n4001 gnd.n4000 585
R9961 gnd.n3852 gnd.n3851 585
R9962 gnd.n3853 gnd.n3852 585
R9963 gnd.n3991 gnd.n3990 585
R9964 gnd.n3992 gnd.n3991 585
R9965 gnd.n3861 gnd.n3860 585
R9966 gnd.n3860 gnd.n3859 585
R9967 gnd.n3986 gnd.n3985 585
R9968 gnd.n3985 gnd.n3984 585
R9969 gnd.n3864 gnd.n3863 585
R9970 gnd.n3975 gnd.n3864 585
R9971 gnd.n3974 gnd.n3973 585
R9972 gnd.n3976 gnd.n3974 585
R9973 gnd.n3872 gnd.n3871 585
R9974 gnd.n3871 gnd.n3870 585
R9975 gnd.n4654 gnd.n2011 585
R9976 gnd.n2011 gnd.n1988 585
R9977 gnd.n4656 gnd.n4655 585
R9978 gnd.n4657 gnd.n4656 585
R9979 gnd.n3366 gnd.n3365 585
R9980 gnd.n3373 gnd.n3365 585
R9981 gnd.n4649 gnd.n4648 585
R9982 gnd.n4648 gnd.n4647 585
R9983 gnd.n3369 gnd.n3368 585
R9984 gnd.n4637 gnd.n3369 585
R9985 gnd.n4368 gnd.n3390 585
R9986 gnd.n3390 gnd.n3380 585
R9987 gnd.n4370 gnd.n4369 585
R9988 gnd.n4371 gnd.n4370 585
R9989 gnd.n3391 gnd.n3389 585
R9990 gnd.n3398 gnd.n3389 585
R9991 gnd.n4363 gnd.n4362 585
R9992 gnd.n4362 gnd.n4361 585
R9993 gnd.n3394 gnd.n3393 585
R9994 gnd.n4350 gnd.n3394 585
R9995 gnd.n4337 gnd.n3416 585
R9996 gnd.n3416 gnd.n3415 585
R9997 gnd.n4339 gnd.n4338 585
R9998 gnd.n4340 gnd.n4339 585
R9999 gnd.n3417 gnd.n3414 585
R10000 gnd.n3424 gnd.n3414 585
R10001 gnd.n4332 gnd.n4331 585
R10002 gnd.n4331 gnd.n4330 585
R10003 gnd.n3420 gnd.n3419 585
R10004 gnd.n4319 gnd.n3420 585
R10005 gnd.n4306 gnd.n3441 585
R10006 gnd.n3441 gnd.n3440 585
R10007 gnd.n4308 gnd.n4307 585
R10008 gnd.n4309 gnd.n4308 585
R10009 gnd.n3442 gnd.n3439 585
R10010 gnd.n3587 gnd.n3439 585
R10011 gnd.n4301 gnd.n4300 585
R10012 gnd.n4300 gnd.n4299 585
R10013 gnd.n3445 gnd.n3444 585
R10014 gnd.n4288 gnd.n3445 585
R10015 gnd.n4275 gnd.n3466 585
R10016 gnd.n3466 gnd.n3465 585
R10017 gnd.n4277 gnd.n4276 585
R10018 gnd.n4278 gnd.n4277 585
R10019 gnd.n3467 gnd.n3464 585
R10020 gnd.n3474 gnd.n3464 585
R10021 gnd.n4270 gnd.n4269 585
R10022 gnd.n4269 gnd.n4268 585
R10023 gnd.n3470 gnd.n3469 585
R10024 gnd.n4257 gnd.n3470 585
R10025 gnd.n4244 gnd.n3492 585
R10026 gnd.n3492 gnd.n3482 585
R10027 gnd.n4246 gnd.n4245 585
R10028 gnd.n4247 gnd.n4246 585
R10029 gnd.n3493 gnd.n3491 585
R10030 gnd.n3500 gnd.n3491 585
R10031 gnd.n4239 gnd.n4238 585
R10032 gnd.n4238 gnd.n4237 585
R10033 gnd.n3496 gnd.n3495 585
R10034 gnd.n4226 gnd.n3496 585
R10035 gnd.n4213 gnd.n3516 585
R10036 gnd.n3612 gnd.n3516 585
R10037 gnd.n4215 gnd.n4214 585
R10038 gnd.n4216 gnd.n4215 585
R10039 gnd.n3517 gnd.n3515 585
R10040 gnd.n3523 gnd.n3515 585
R10041 gnd.n4208 gnd.n4207 585
R10042 gnd.n4207 gnd.n4206 585
R10043 gnd.n3520 gnd.n3519 585
R10044 gnd.n4195 gnd.n3520 585
R10045 gnd.n4177 gnd.n4176 585
R10046 gnd.n4178 gnd.n4177 585
R10047 gnd.n3699 gnd.n3698 585
R10048 gnd.n4160 gnd.n3698 585
R10049 gnd.n4172 gnd.n4171 585
R10050 gnd.n4171 gnd.n3684 585
R10051 gnd.n4170 gnd.n3701 585
R10052 gnd.n4170 gnd.n3683 585
R10053 gnd.n4169 gnd.n3703 585
R10054 gnd.n4169 gnd.n4168 585
R10055 gnd.n4121 gnd.n3702 585
R10056 gnd.n4147 gnd.n3702 585
R10057 gnd.n4123 gnd.n4122 585
R10058 gnd.n4122 gnd.n3711 585
R10059 gnd.n4124 gnd.n3730 585
R10060 gnd.n3730 gnd.n3719 585
R10061 gnd.n4126 gnd.n4125 585
R10062 gnd.n4127 gnd.n4126 585
R10063 gnd.n3731 gnd.n3729 585
R10064 gnd.n3738 gnd.n3729 585
R10065 gnd.n4113 gnd.n4112 585
R10066 gnd.n4112 gnd.n4111 585
R10067 gnd.n3734 gnd.n3733 585
R10068 gnd.n4101 gnd.n3734 585
R10069 gnd.n4088 gnd.n3758 585
R10070 gnd.n3758 gnd.n3757 585
R10071 gnd.n4090 gnd.n4089 585
R10072 gnd.n4091 gnd.n4090 585
R10073 gnd.n3759 gnd.n3756 585
R10074 gnd.n3766 gnd.n3756 585
R10075 gnd.n4083 gnd.n4082 585
R10076 gnd.n4082 gnd.n4081 585
R10077 gnd.n3762 gnd.n3761 585
R10078 gnd.n4070 gnd.n3762 585
R10079 gnd.n4057 gnd.n3783 585
R10080 gnd.n3783 gnd.n3782 585
R10081 gnd.n4059 gnd.n4058 585
R10082 gnd.n4060 gnd.n4059 585
R10083 gnd.n4053 gnd.n3781 585
R10084 gnd.n4052 gnd.n4051 585
R10085 gnd.n3786 gnd.n3785 585
R10086 gnd.n4049 gnd.n3786 585
R10087 gnd.n3808 gnd.n3807 585
R10088 gnd.n3811 gnd.n3810 585
R10089 gnd.n3809 gnd.n3804 585
R10090 gnd.n3816 gnd.n3815 585
R10091 gnd.n3818 gnd.n3817 585
R10092 gnd.n3821 gnd.n3820 585
R10093 gnd.n3819 gnd.n3802 585
R10094 gnd.n3826 gnd.n3825 585
R10095 gnd.n3828 gnd.n3827 585
R10096 gnd.n3831 gnd.n3830 585
R10097 gnd.n3829 gnd.n3800 585
R10098 gnd.n3836 gnd.n3835 585
R10099 gnd.n3840 gnd.n3837 585
R10100 gnd.n3841 gnd.n3778 585
R10101 gnd.n3362 gnd.n2026 585
R10102 gnd.n4723 gnd.n4722 585
R10103 gnd.n4725 gnd.n4724 585
R10104 gnd.n4727 gnd.n4726 585
R10105 gnd.n4729 gnd.n4728 585
R10106 gnd.n4731 gnd.n4730 585
R10107 gnd.n4733 gnd.n4732 585
R10108 gnd.n4735 gnd.n4734 585
R10109 gnd.n4737 gnd.n4736 585
R10110 gnd.n4739 gnd.n4738 585
R10111 gnd.n4741 gnd.n4740 585
R10112 gnd.n4743 gnd.n4742 585
R10113 gnd.n4745 gnd.n4744 585
R10114 gnd.n4748 gnd.n4747 585
R10115 gnd.n4746 gnd.n2014 585
R10116 gnd.n4752 gnd.n2012 585
R10117 gnd.n4754 gnd.n4753 585
R10118 gnd.n4755 gnd.n4754 585
R10119 gnd.n3363 gnd.n3360 585
R10120 gnd.n3363 gnd.n1988 585
R10121 gnd.n4659 gnd.n4658 585
R10122 gnd.n4658 gnd.n4657 585
R10123 gnd.n3361 gnd.n3359 585
R10124 gnd.n3373 gnd.n3361 585
R10125 gnd.n4640 gnd.n3371 585
R10126 gnd.n4647 gnd.n3371 585
R10127 gnd.n4639 gnd.n4638 585
R10128 gnd.n4638 gnd.n4637 585
R10129 gnd.n3379 gnd.n3377 585
R10130 gnd.n3380 gnd.n3379 585
R10131 gnd.n4373 gnd.n4372 585
R10132 gnd.n4372 gnd.n4371 585
R10133 gnd.n3386 gnd.n3385 585
R10134 gnd.n3398 gnd.n3386 585
R10135 gnd.n4353 gnd.n3396 585
R10136 gnd.n4361 gnd.n3396 585
R10137 gnd.n4352 gnd.n4351 585
R10138 gnd.n4351 gnd.n4350 585
R10139 gnd.n3405 gnd.n3403 585
R10140 gnd.n3415 gnd.n3405 585
R10141 gnd.n4342 gnd.n4341 585
R10142 gnd.n4341 gnd.n4340 585
R10143 gnd.n3411 gnd.n3410 585
R10144 gnd.n3424 gnd.n3411 585
R10145 gnd.n4322 gnd.n3422 585
R10146 gnd.n4330 gnd.n3422 585
R10147 gnd.n4321 gnd.n4320 585
R10148 gnd.n4320 gnd.n4319 585
R10149 gnd.n3431 gnd.n3429 585
R10150 gnd.n3440 gnd.n3431 585
R10151 gnd.n4311 gnd.n4310 585
R10152 gnd.n4310 gnd.n4309 585
R10153 gnd.n3437 gnd.n3436 585
R10154 gnd.n3587 gnd.n3437 585
R10155 gnd.n4291 gnd.n3447 585
R10156 gnd.n4299 gnd.n3447 585
R10157 gnd.n4290 gnd.n4289 585
R10158 gnd.n4289 gnd.n4288 585
R10159 gnd.n3455 gnd.n3453 585
R10160 gnd.n3465 gnd.n3455 585
R10161 gnd.n4280 gnd.n4279 585
R10162 gnd.n4279 gnd.n4278 585
R10163 gnd.n3461 gnd.n3460 585
R10164 gnd.n3474 gnd.n3461 585
R10165 gnd.n4260 gnd.n3472 585
R10166 gnd.n4268 gnd.n3472 585
R10167 gnd.n4259 gnd.n4258 585
R10168 gnd.n4258 gnd.n4257 585
R10169 gnd.n3481 gnd.n3479 585
R10170 gnd.n3482 gnd.n3481 585
R10171 gnd.n4249 gnd.n4248 585
R10172 gnd.n4248 gnd.n4247 585
R10173 gnd.n3488 gnd.n3487 585
R10174 gnd.n3500 gnd.n3488 585
R10175 gnd.n4229 gnd.n3498 585
R10176 gnd.n4237 gnd.n3498 585
R10177 gnd.n4228 gnd.n4227 585
R10178 gnd.n4227 gnd.n4226 585
R10179 gnd.n3507 gnd.n3505 585
R10180 gnd.n3612 gnd.n3507 585
R10181 gnd.n4218 gnd.n4217 585
R10182 gnd.n4217 gnd.n4216 585
R10183 gnd.n3513 gnd.n3512 585
R10184 gnd.n3523 gnd.n3513 585
R10185 gnd.n4198 gnd.n3521 585
R10186 gnd.n4206 gnd.n3521 585
R10187 gnd.n4197 gnd.n4196 585
R10188 gnd.n4196 gnd.n4195 585
R10189 gnd.n3530 gnd.n3528 585
R10190 gnd.n4178 gnd.n3530 585
R10191 gnd.n4161 gnd.n4158 585
R10192 gnd.n4161 gnd.n4160 585
R10193 gnd.n4163 gnd.n4162 585
R10194 gnd.n4162 gnd.n3684 585
R10195 gnd.n4164 gnd.n3706 585
R10196 gnd.n3706 gnd.n3683 585
R10197 gnd.n4166 gnd.n4165 585
R10198 gnd.n4168 gnd.n4166 585
R10199 gnd.n3707 gnd.n3705 585
R10200 gnd.n4147 gnd.n3705 585
R10201 gnd.n4131 gnd.n4130 585
R10202 gnd.n4130 gnd.n3711 585
R10203 gnd.n4129 gnd.n3725 585
R10204 gnd.n4129 gnd.n3719 585
R10205 gnd.n4128 gnd.n3727 585
R10206 gnd.n4128 gnd.n4127 585
R10207 gnd.n4105 gnd.n3726 585
R10208 gnd.n3738 gnd.n3726 585
R10209 gnd.n4104 gnd.n3736 585
R10210 gnd.n4111 gnd.n3736 585
R10211 gnd.n4103 gnd.n4102 585
R10212 gnd.n4102 gnd.n4101 585
R10213 gnd.n3747 gnd.n3744 585
R10214 gnd.n3757 gnd.n3747 585
R10215 gnd.n4093 gnd.n4092 585
R10216 gnd.n4092 gnd.n4091 585
R10217 gnd.n3753 gnd.n3752 585
R10218 gnd.n3766 gnd.n3753 585
R10219 gnd.n4073 gnd.n3764 585
R10220 gnd.n4081 gnd.n3764 585
R10221 gnd.n4072 gnd.n4071 585
R10222 gnd.n4071 gnd.n4070 585
R10223 gnd.n3773 gnd.n3771 585
R10224 gnd.n3782 gnd.n3773 585
R10225 gnd.n4062 gnd.n4061 585
R10226 gnd.n4061 gnd.n4060 585
R10227 gnd.n5770 gnd.n5769 585
R10228 gnd.n5771 gnd.n5770 585
R10229 gnd.n1360 gnd.n1358 585
R10230 gnd.n5694 gnd.n1358 585
R10231 gnd.n5564 gnd.n1660 585
R10232 gnd.n5386 gnd.n1660 585
R10233 gnd.n5566 gnd.n5565 585
R10234 gnd.n5567 gnd.n5566 585
R10235 gnd.n1661 gnd.n1659 585
R10236 gnd.n5384 gnd.n1659 585
R10237 gnd.n5559 gnd.n5558 585
R10238 gnd.n5558 gnd.n5557 585
R10239 gnd.n1664 gnd.n1663 585
R10240 gnd.n5373 gnd.n1664 585
R10241 gnd.n5548 gnd.n5547 585
R10242 gnd.n5549 gnd.n5548 585
R10243 gnd.n1678 gnd.n1677 585
R10244 gnd.n5328 gnd.n1677 585
R10245 gnd.n5543 gnd.n5542 585
R10246 gnd.n5542 gnd.n5541 585
R10247 gnd.n1681 gnd.n1680 585
R10248 gnd.n5334 gnd.n1681 585
R10249 gnd.n5532 gnd.n5531 585
R10250 gnd.n5533 gnd.n5532 585
R10251 gnd.n1695 gnd.n1694 585
R10252 gnd.n5320 gnd.n1694 585
R10253 gnd.n5527 gnd.n5526 585
R10254 gnd.n5526 gnd.n5525 585
R10255 gnd.n1698 gnd.n1697 585
R10256 gnd.n5316 gnd.n1698 585
R10257 gnd.n5516 gnd.n5515 585
R10258 gnd.n5517 gnd.n5516 585
R10259 gnd.n1712 gnd.n1711 585
R10260 gnd.n5289 gnd.n1711 585
R10261 gnd.n5511 gnd.n5510 585
R10262 gnd.n5510 gnd.n5509 585
R10263 gnd.n1715 gnd.n1714 585
R10264 gnd.n5295 gnd.n1715 585
R10265 gnd.n5500 gnd.n5499 585
R10266 gnd.n5501 gnd.n5500 585
R10267 gnd.n1729 gnd.n1728 585
R10268 gnd.n5280 gnd.n1728 585
R10269 gnd.n5495 gnd.n5494 585
R10270 gnd.n5494 gnd.n5493 585
R10271 gnd.n1732 gnd.n1731 585
R10272 gnd.n5276 gnd.n1732 585
R10273 gnd.n5484 gnd.n5483 585
R10274 gnd.n5485 gnd.n5484 585
R10275 gnd.n1746 gnd.n1745 585
R10276 gnd.n5249 gnd.n1745 585
R10277 gnd.n5479 gnd.n5478 585
R10278 gnd.n5478 gnd.n5477 585
R10279 gnd.n1749 gnd.n1748 585
R10280 gnd.n5429 gnd.n1749 585
R10281 gnd.n5468 gnd.n5467 585
R10282 gnd.n5469 gnd.n5468 585
R10283 gnd.n1763 gnd.n1762 585
R10284 gnd.n5241 gnd.n1762 585
R10285 gnd.n5440 gnd.n5439 585
R10286 gnd.n5441 gnd.n5440 585
R10287 gnd.n5438 gnd.n1787 585
R10288 gnd.n5233 gnd.n1787 585
R10289 gnd.n5449 gnd.n5448 585
R10290 gnd.n5448 gnd.n5447 585
R10291 gnd.n5451 gnd.n5450 585
R10292 gnd.n5451 gnd.n1786 585
R10293 gnd.n5454 gnd.n5453 585
R10294 gnd.n5455 gnd.n5454 585
R10295 gnd.n5452 gnd.n1772 585
R10296 gnd.n1775 gnd.n1772 585
R10297 gnd.n5463 gnd.n5462 585
R10298 gnd.n5462 gnd.n5461 585
R10299 gnd.n5464 gnd.n1771 585
R10300 gnd.n5217 gnd.n1771 585
R10301 gnd.n1876 gnd.n1770 585
R10302 gnd.n1876 gnd.n1867 585
R10303 gnd.n5198 gnd.n5197 585
R10304 gnd.n5199 gnd.n5198 585
R10305 gnd.n5196 gnd.n1875 585
R10306 gnd.n5184 gnd.n1875 585
R10307 gnd.n1881 gnd.n1877 585
R10308 gnd.n1884 gnd.n1881 585
R10309 gnd.n5192 gnd.n5191 585
R10310 gnd.n5191 gnd.n5190 585
R10311 gnd.n1880 gnd.n1879 585
R10312 gnd.n5173 gnd.n1880 585
R10313 gnd.n5157 gnd.n1912 585
R10314 gnd.n1912 gnd.n1902 585
R10315 gnd.n5159 gnd.n5158 585
R10316 gnd.n5160 gnd.n5159 585
R10317 gnd.n1913 gnd.n1911 585
R10318 gnd.n1911 gnd.n1908 585
R10319 gnd.n5152 gnd.n5151 585
R10320 gnd.n5151 gnd.n5150 585
R10321 gnd.n1916 gnd.n1915 585
R10322 gnd.n1928 gnd.n1916 585
R10323 gnd.n5133 gnd.n5132 585
R10324 gnd.n5134 gnd.n5133 585
R10325 gnd.n1930 gnd.n1929 585
R10326 gnd.n1929 gnd.n1925 585
R10327 gnd.n5128 gnd.n5127 585
R10328 gnd.n5127 gnd.n5126 585
R10329 gnd.n1933 gnd.n1932 585
R10330 gnd.n1934 gnd.n1933 585
R10331 gnd.n5117 gnd.n5116 585
R10332 gnd.n5118 gnd.n5117 585
R10333 gnd.n1946 gnd.n1945 585
R10334 gnd.n1945 gnd.n1942 585
R10335 gnd.n5112 gnd.n5111 585
R10336 gnd.n5111 gnd.n5110 585
R10337 gnd.n1949 gnd.n1948 585
R10338 gnd.n1960 gnd.n1949 585
R10339 gnd.n5101 gnd.n5100 585
R10340 gnd.n5102 gnd.n5101 585
R10341 gnd.n1962 gnd.n1961 585
R10342 gnd.n1961 gnd.n1957 585
R10343 gnd.n5096 gnd.n5095 585
R10344 gnd.n5095 gnd.n5094 585
R10345 gnd.n1965 gnd.n1964 585
R10346 gnd.n1966 gnd.n1965 585
R10347 gnd.n5085 gnd.n5084 585
R10348 gnd.n5086 gnd.n5085 585
R10349 gnd.n1978 gnd.n1977 585
R10350 gnd.n1977 gnd.n1974 585
R10351 gnd.n5080 gnd.n5079 585
R10352 gnd.n5079 gnd.n5078 585
R10353 gnd.n1981 gnd.n1980 585
R10354 gnd.n4872 gnd.n1981 585
R10355 gnd.n5069 gnd.n5068 585
R10356 gnd.n5070 gnd.n5069 585
R10357 gnd.n5065 gnd.n4873 585
R10358 gnd.n5064 gnd.n5063 585
R10359 gnd.n5061 gnd.n4875 585
R10360 gnd.n5061 gnd.n4756 585
R10361 gnd.n5060 gnd.n5059 585
R10362 gnd.n5058 gnd.n5057 585
R10363 gnd.n5056 gnd.n4880 585
R10364 gnd.n5054 gnd.n5053 585
R10365 gnd.n5052 gnd.n4881 585
R10366 gnd.n5051 gnd.n5050 585
R10367 gnd.n5048 gnd.n4886 585
R10368 gnd.n5046 gnd.n5045 585
R10369 gnd.n5044 gnd.n4887 585
R10370 gnd.n5043 gnd.n5042 585
R10371 gnd.n5040 gnd.n4892 585
R10372 gnd.n5038 gnd.n5037 585
R10373 gnd.n5036 gnd.n4893 585
R10374 gnd.n5035 gnd.n5034 585
R10375 gnd.n5032 gnd.n4898 585
R10376 gnd.n5030 gnd.n5029 585
R10377 gnd.n5028 gnd.n4899 585
R10378 gnd.n5027 gnd.n5026 585
R10379 gnd.n5024 gnd.n4907 585
R10380 gnd.n5022 gnd.n5021 585
R10381 gnd.n5020 gnd.n4908 585
R10382 gnd.n5019 gnd.n5018 585
R10383 gnd.n5016 gnd.n4913 585
R10384 gnd.n5014 gnd.n5013 585
R10385 gnd.n5012 gnd.n4914 585
R10386 gnd.n5011 gnd.n5010 585
R10387 gnd.n5008 gnd.n4919 585
R10388 gnd.n5006 gnd.n5005 585
R10389 gnd.n5004 gnd.n4920 585
R10390 gnd.n5003 gnd.n5002 585
R10391 gnd.n5000 gnd.n4925 585
R10392 gnd.n4998 gnd.n4997 585
R10393 gnd.n4996 gnd.n4926 585
R10394 gnd.n4995 gnd.n4931 585
R10395 gnd.n4988 gnd.n4934 585
R10396 gnd.n4991 gnd.n4990 585
R10397 gnd.n5701 gnd.n5700 585
R10398 gnd.n5703 gnd.n1643 585
R10399 gnd.n5705 gnd.n5704 585
R10400 gnd.n5706 gnd.n1636 585
R10401 gnd.n5708 gnd.n5707 585
R10402 gnd.n5710 gnd.n1634 585
R10403 gnd.n5712 gnd.n5711 585
R10404 gnd.n5713 gnd.n1629 585
R10405 gnd.n5715 gnd.n5714 585
R10406 gnd.n5717 gnd.n1627 585
R10407 gnd.n5719 gnd.n5718 585
R10408 gnd.n5720 gnd.n1622 585
R10409 gnd.n5722 gnd.n5721 585
R10410 gnd.n5724 gnd.n1620 585
R10411 gnd.n5726 gnd.n5725 585
R10412 gnd.n5727 gnd.n1615 585
R10413 gnd.n5729 gnd.n5728 585
R10414 gnd.n5731 gnd.n1613 585
R10415 gnd.n5733 gnd.n5732 585
R10416 gnd.n5734 gnd.n1607 585
R10417 gnd.n5736 gnd.n5735 585
R10418 gnd.n5740 gnd.n1386 585
R10419 gnd.n5742 gnd.n5741 585
R10420 gnd.n5743 gnd.n1381 585
R10421 gnd.n5745 gnd.n5744 585
R10422 gnd.n5747 gnd.n1379 585
R10423 gnd.n5749 gnd.n5748 585
R10424 gnd.n5750 gnd.n1374 585
R10425 gnd.n5752 gnd.n5751 585
R10426 gnd.n5754 gnd.n1372 585
R10427 gnd.n5756 gnd.n5755 585
R10428 gnd.n5757 gnd.n1366 585
R10429 gnd.n5759 gnd.n5758 585
R10430 gnd.n5761 gnd.n1365 585
R10431 gnd.n5762 gnd.n1363 585
R10432 gnd.n5765 gnd.n5764 585
R10433 gnd.n5766 gnd.n1359 585
R10434 gnd.n1364 gnd.n1359 585
R10435 gnd.n5697 gnd.n1355 585
R10436 gnd.n5771 gnd.n1355 585
R10437 gnd.n5696 gnd.n5695 585
R10438 gnd.n5695 gnd.n5694 585
R10439 gnd.n1648 gnd.n1647 585
R10440 gnd.n5386 gnd.n1648 585
R10441 gnd.n5381 gnd.n1656 585
R10442 gnd.n5567 gnd.n1656 585
R10443 gnd.n5383 gnd.n5382 585
R10444 gnd.n5384 gnd.n5383 585
R10445 gnd.n1831 gnd.n1666 585
R10446 gnd.n5557 gnd.n1666 585
R10447 gnd.n5375 gnd.n5374 585
R10448 gnd.n5374 gnd.n5373 585
R10449 gnd.n1833 gnd.n1675 585
R10450 gnd.n5549 gnd.n1675 585
R10451 gnd.n5330 gnd.n5329 585
R10452 gnd.n5329 gnd.n5328 585
R10453 gnd.n5331 gnd.n1682 585
R10454 gnd.n5541 gnd.n1682 585
R10455 gnd.n5333 gnd.n5332 585
R10456 gnd.n5334 gnd.n5333 585
R10457 gnd.n1840 gnd.n1691 585
R10458 gnd.n5533 gnd.n1691 585
R10459 gnd.n5322 gnd.n5321 585
R10460 gnd.n5321 gnd.n5320 585
R10461 gnd.n5319 gnd.n1700 585
R10462 gnd.n5525 gnd.n1700 585
R10463 gnd.n5318 gnd.n5317 585
R10464 gnd.n5317 gnd.n5316 585
R10465 gnd.n1842 gnd.n1709 585
R10466 gnd.n5517 gnd.n1709 585
R10467 gnd.n5291 gnd.n5290 585
R10468 gnd.n5290 gnd.n5289 585
R10469 gnd.n5292 gnd.n1716 585
R10470 gnd.n5509 gnd.n1716 585
R10471 gnd.n5294 gnd.n5293 585
R10472 gnd.n5295 gnd.n5294 585
R10473 gnd.n1850 gnd.n1725 585
R10474 gnd.n5501 gnd.n1725 585
R10475 gnd.n5282 gnd.n5281 585
R10476 gnd.n5281 gnd.n5280 585
R10477 gnd.n5279 gnd.n1734 585
R10478 gnd.n5493 gnd.n1734 585
R10479 gnd.n5278 gnd.n5277 585
R10480 gnd.n5277 gnd.n5276 585
R10481 gnd.n1852 gnd.n1743 585
R10482 gnd.n5485 gnd.n1743 585
R10483 gnd.n5251 gnd.n5250 585
R10484 gnd.n5250 gnd.n5249 585
R10485 gnd.n5248 gnd.n1750 585
R10486 gnd.n5477 gnd.n1750 585
R10487 gnd.n5247 gnd.n1806 585
R10488 gnd.n5429 gnd.n1806 585
R10489 gnd.n1854 gnd.n1759 585
R10490 gnd.n5469 gnd.n1759 585
R10491 gnd.n5243 gnd.n5242 585
R10492 gnd.n5242 gnd.n5241 585
R10493 gnd.n1856 gnd.n1796 585
R10494 gnd.n5441 gnd.n1796 585
R10495 gnd.n5232 gnd.n5231 585
R10496 gnd.n5233 gnd.n5232 585
R10497 gnd.n1860 gnd.n1789 585
R10498 gnd.n5447 gnd.n1789 585
R10499 gnd.n5227 gnd.n5226 585
R10500 gnd.n5226 gnd.n1786 585
R10501 gnd.n5225 gnd.n1784 585
R10502 gnd.n5455 gnd.n1784 585
R10503 gnd.n5224 gnd.n5223 585
R10504 gnd.n5223 gnd.n1775 585
R10505 gnd.n1863 gnd.n1773 585
R10506 gnd.n5461 gnd.n1773 585
R10507 gnd.n5219 gnd.n5218 585
R10508 gnd.n5218 gnd.n5217 585
R10509 gnd.n1866 gnd.n1865 585
R10510 gnd.n1867 gnd.n1866 585
R10511 gnd.n5181 gnd.n1873 585
R10512 gnd.n5199 gnd.n1873 585
R10513 gnd.n5183 gnd.n5182 585
R10514 gnd.n5184 gnd.n5183 585
R10515 gnd.n1898 gnd.n1897 585
R10516 gnd.n1897 gnd.n1884 585
R10517 gnd.n5176 gnd.n1882 585
R10518 gnd.n5190 gnd.n1882 585
R10519 gnd.n5175 gnd.n5174 585
R10520 gnd.n5174 gnd.n5173 585
R10521 gnd.n1901 gnd.n1900 585
R10522 gnd.n1902 gnd.n1901 585
R10523 gnd.n4957 gnd.n1909 585
R10524 gnd.n5160 gnd.n1909 585
R10525 gnd.n4959 gnd.n4958 585
R10526 gnd.n4958 gnd.n1908 585
R10527 gnd.n4960 gnd.n1917 585
R10528 gnd.n5150 gnd.n1917 585
R10529 gnd.n4962 gnd.n4961 585
R10530 gnd.n4961 gnd.n1928 585
R10531 gnd.n4963 gnd.n1926 585
R10532 gnd.n5134 gnd.n1926 585
R10533 gnd.n4965 gnd.n4964 585
R10534 gnd.n4964 gnd.n1925 585
R10535 gnd.n4966 gnd.n1935 585
R10536 gnd.n5126 gnd.n1935 585
R10537 gnd.n4968 gnd.n4967 585
R10538 gnd.n4967 gnd.n1934 585
R10539 gnd.n4969 gnd.n1943 585
R10540 gnd.n5118 gnd.n1943 585
R10541 gnd.n4971 gnd.n4970 585
R10542 gnd.n4970 gnd.n1942 585
R10543 gnd.n4972 gnd.n1950 585
R10544 gnd.n5110 gnd.n1950 585
R10545 gnd.n4974 gnd.n4973 585
R10546 gnd.n4973 gnd.n1960 585
R10547 gnd.n4975 gnd.n1958 585
R10548 gnd.n5102 gnd.n1958 585
R10549 gnd.n4977 gnd.n4976 585
R10550 gnd.n4976 gnd.n1957 585
R10551 gnd.n4978 gnd.n1967 585
R10552 gnd.n5094 gnd.n1967 585
R10553 gnd.n4980 gnd.n4979 585
R10554 gnd.n4979 gnd.n1966 585
R10555 gnd.n4981 gnd.n1975 585
R10556 gnd.n5086 gnd.n1975 585
R10557 gnd.n4983 gnd.n4982 585
R10558 gnd.n4982 gnd.n1974 585
R10559 gnd.n4984 gnd.n1982 585
R10560 gnd.n5078 gnd.n1982 585
R10561 gnd.n4985 gnd.n4936 585
R10562 gnd.n4936 gnd.n4872 585
R10563 gnd.n4986 gnd.n4757 585
R10564 gnd.n5070 gnd.n4757 585
R10565 gnd.n7572 gnd.n7571 585
R10566 gnd.n7573 gnd.n7572 585
R10567 gnd.n128 gnd.n126 585
R10568 gnd.n126 gnd.n122 585
R10569 gnd.n7492 gnd.n7491 585
R10570 gnd.n7493 gnd.n7492 585
R10571 gnd.n205 gnd.n204 585
R10572 gnd.n204 gnd.n202 585
R10573 gnd.n7487 gnd.n7486 585
R10574 gnd.n7486 gnd.n7485 585
R10575 gnd.n208 gnd.n207 585
R10576 gnd.n209 gnd.n208 585
R10577 gnd.n7408 gnd.n7407 585
R10578 gnd.n7409 gnd.n7408 585
R10579 gnd.n221 gnd.n220 585
R10580 gnd.n228 gnd.n220 585
R10581 gnd.n7403 gnd.n7402 585
R10582 gnd.n7402 gnd.n7401 585
R10583 gnd.n224 gnd.n223 585
R10584 gnd.n225 gnd.n224 585
R10585 gnd.n7392 gnd.n7391 585
R10586 gnd.n7393 gnd.n7392 585
R10587 gnd.n238 gnd.n237 585
R10588 gnd.n237 gnd.n234 585
R10589 gnd.n7387 gnd.n7386 585
R10590 gnd.n7386 gnd.n7385 585
R10591 gnd.n241 gnd.n240 585
R10592 gnd.n250 gnd.n241 585
R10593 gnd.n7376 gnd.n7375 585
R10594 gnd.n7377 gnd.n7376 585
R10595 gnd.n252 gnd.n251 585
R10596 gnd.n259 gnd.n251 585
R10597 gnd.n7371 gnd.n7370 585
R10598 gnd.n7370 gnd.n7369 585
R10599 gnd.n255 gnd.n254 585
R10600 gnd.n256 gnd.n255 585
R10601 gnd.n7360 gnd.n7359 585
R10602 gnd.n7361 gnd.n7360 585
R10603 gnd.n268 gnd.n267 585
R10604 gnd.n267 gnd.n265 585
R10605 gnd.n7355 gnd.n7354 585
R10606 gnd.n7354 gnd.n7353 585
R10607 gnd.n271 gnd.n270 585
R10608 gnd.n280 gnd.n271 585
R10609 gnd.n7344 gnd.n7343 585
R10610 gnd.n7345 gnd.n7344 585
R10611 gnd.n282 gnd.n281 585
R10612 gnd.n289 gnd.n281 585
R10613 gnd.n7339 gnd.n7338 585
R10614 gnd.n7338 gnd.n7337 585
R10615 gnd.n285 gnd.n284 585
R10616 gnd.n286 gnd.n285 585
R10617 gnd.n7328 gnd.n7327 585
R10618 gnd.n7329 gnd.n7328 585
R10619 gnd.n298 gnd.n297 585
R10620 gnd.n297 gnd.n295 585
R10621 gnd.n7304 gnd.n7303 585
R10622 gnd.n7305 gnd.n7304 585
R10623 gnd.n7302 gnd.n328 585
R10624 gnd.n7302 gnd.n7301 585
R10625 gnd.n327 gnd.n326 585
R10626 gnd.n330 gnd.n326 585
R10627 gnd.n7227 gnd.n7226 585
R10628 gnd.n7228 gnd.n7227 585
R10629 gnd.n7225 gnd.n7224 585
R10630 gnd.n7224 gnd.n336 585
R10631 gnd.n7223 gnd.n338 585
R10632 gnd.n7223 gnd.n7222 585
R10633 gnd.n337 gnd.n307 585
R10634 gnd.n7202 gnd.n307 585
R10635 gnd.n7322 gnd.n7321 585
R10636 gnd.n7321 gnd.n7320 585
R10637 gnd.n7323 gnd.n306 585
R10638 gnd.n7211 gnd.n306 585
R10639 gnd.n364 gnd.n305 585
R10640 gnd.n364 gnd.n349 585
R10641 gnd.n7189 gnd.n7188 585
R10642 gnd.n7190 gnd.n7189 585
R10643 gnd.n7187 gnd.n363 585
R10644 gnd.n7169 gnd.n363 585
R10645 gnd.n369 gnd.n365 585
R10646 gnd.n6930 gnd.n369 585
R10647 gnd.n7183 gnd.n7182 585
R10648 gnd.n7182 gnd.n7181 585
R10649 gnd.n368 gnd.n367 585
R10650 gnd.n7159 gnd.n368 585
R10651 gnd.n7137 gnd.n7136 585
R10652 gnd.n7138 gnd.n7137 585
R10653 gnd.n397 gnd.n396 585
R10654 gnd.n6938 gnd.n396 585
R10655 gnd.n7132 gnd.n7131 585
R10656 gnd.n7131 gnd.n7130 585
R10657 gnd.n400 gnd.n399 585
R10658 gnd.n6917 gnd.n400 585
R10659 gnd.n7118 gnd.n7117 585
R10660 gnd.n7119 gnd.n7118 585
R10661 gnd.n416 gnd.n415 585
R10662 gnd.n6898 gnd.n415 585
R10663 gnd.n7113 gnd.n7112 585
R10664 gnd.n7112 gnd.n7111 585
R10665 gnd.n419 gnd.n418 585
R10666 gnd.n6904 gnd.n419 585
R10667 gnd.n7102 gnd.n7101 585
R10668 gnd.n7103 gnd.n7102 585
R10669 gnd.n433 gnd.n432 585
R10670 gnd.n6890 gnd.n432 585
R10671 gnd.n7097 gnd.n7096 585
R10672 gnd.n7096 gnd.n7095 585
R10673 gnd.n436 gnd.n435 585
R10674 gnd.n6886 gnd.n436 585
R10675 gnd.n7086 gnd.n7085 585
R10676 gnd.n7087 gnd.n7086 585
R10677 gnd.n450 gnd.n449 585
R10678 gnd.n6859 gnd.n449 585
R10679 gnd.n7081 gnd.n7080 585
R10680 gnd.n7080 gnd.n7079 585
R10681 gnd.n453 gnd.n452 585
R10682 gnd.n6865 gnd.n453 585
R10683 gnd.n7070 gnd.n7069 585
R10684 gnd.n7071 gnd.n7070 585
R10685 gnd.n467 gnd.n466 585
R10686 gnd.n6850 gnd.n466 585
R10687 gnd.n7065 gnd.n7064 585
R10688 gnd.n7064 gnd.n7063 585
R10689 gnd.n470 gnd.n469 585
R10690 gnd.n6846 gnd.n470 585
R10691 gnd.n7054 gnd.n7053 585
R10692 gnd.n7055 gnd.n7054 585
R10693 gnd.n485 gnd.n484 585
R10694 gnd.n6974 gnd.n484 585
R10695 gnd.n7049 gnd.n7048 585
R10696 gnd.n488 gnd.n487 585
R10697 gnd.n7045 gnd.n7044 585
R10698 gnd.n7046 gnd.n7045 585
R10699 gnd.n7043 gnd.n519 585
R10700 gnd.n7042 gnd.n7041 585
R10701 gnd.n7040 gnd.n7039 585
R10702 gnd.n7038 gnd.n7037 585
R10703 gnd.n7036 gnd.n7035 585
R10704 gnd.n7034 gnd.n7033 585
R10705 gnd.n7032 gnd.n7031 585
R10706 gnd.n7030 gnd.n7029 585
R10707 gnd.n7028 gnd.n7027 585
R10708 gnd.n7026 gnd.n7025 585
R10709 gnd.n7024 gnd.n7023 585
R10710 gnd.n7022 gnd.n7021 585
R10711 gnd.n7020 gnd.n7019 585
R10712 gnd.n7017 gnd.n7016 585
R10713 gnd.n7015 gnd.n7014 585
R10714 gnd.n7013 gnd.n7012 585
R10715 gnd.n7011 gnd.n7010 585
R10716 gnd.n7009 gnd.n7008 585
R10717 gnd.n7007 gnd.n7006 585
R10718 gnd.n7005 gnd.n7004 585
R10719 gnd.n7003 gnd.n7002 585
R10720 gnd.n7001 gnd.n7000 585
R10721 gnd.n6999 gnd.n6998 585
R10722 gnd.n6997 gnd.n6996 585
R10723 gnd.n6995 gnd.n6994 585
R10724 gnd.n6993 gnd.n6992 585
R10725 gnd.n6991 gnd.n6990 585
R10726 gnd.n6989 gnd.n6988 585
R10727 gnd.n6987 gnd.n6986 585
R10728 gnd.n6985 gnd.n6984 585
R10729 gnd.n6983 gnd.n6982 585
R10730 gnd.n6981 gnd.n557 585
R10731 gnd.n561 gnd.n558 585
R10732 gnd.n6977 gnd.n6976 585
R10733 gnd.n196 gnd.n195 585
R10734 gnd.n7501 gnd.n191 585
R10735 gnd.n7503 gnd.n7502 585
R10736 gnd.n7505 gnd.n189 585
R10737 gnd.n7507 gnd.n7506 585
R10738 gnd.n7508 gnd.n184 585
R10739 gnd.n7510 gnd.n7509 585
R10740 gnd.n7512 gnd.n182 585
R10741 gnd.n7514 gnd.n7513 585
R10742 gnd.n7515 gnd.n177 585
R10743 gnd.n7517 gnd.n7516 585
R10744 gnd.n7519 gnd.n175 585
R10745 gnd.n7521 gnd.n7520 585
R10746 gnd.n7522 gnd.n170 585
R10747 gnd.n7524 gnd.n7523 585
R10748 gnd.n7526 gnd.n168 585
R10749 gnd.n7528 gnd.n7527 585
R10750 gnd.n7529 gnd.n163 585
R10751 gnd.n7531 gnd.n7530 585
R10752 gnd.n7533 gnd.n161 585
R10753 gnd.n7535 gnd.n7534 585
R10754 gnd.n7539 gnd.n156 585
R10755 gnd.n7541 gnd.n7540 585
R10756 gnd.n7543 gnd.n154 585
R10757 gnd.n7545 gnd.n7544 585
R10758 gnd.n7546 gnd.n149 585
R10759 gnd.n7548 gnd.n7547 585
R10760 gnd.n7550 gnd.n147 585
R10761 gnd.n7552 gnd.n7551 585
R10762 gnd.n7553 gnd.n142 585
R10763 gnd.n7555 gnd.n7554 585
R10764 gnd.n7557 gnd.n140 585
R10765 gnd.n7559 gnd.n7558 585
R10766 gnd.n7560 gnd.n135 585
R10767 gnd.n7562 gnd.n7561 585
R10768 gnd.n7564 gnd.n133 585
R10769 gnd.n7566 gnd.n7565 585
R10770 gnd.n7567 gnd.n131 585
R10771 gnd.n7568 gnd.n127 585
R10772 gnd.n127 gnd.n124 585
R10773 gnd.n7497 gnd.n123 585
R10774 gnd.n7573 gnd.n123 585
R10775 gnd.n7496 gnd.n7495 585
R10776 gnd.n7495 gnd.n122 585
R10777 gnd.n7494 gnd.n200 585
R10778 gnd.n7494 gnd.n7493 585
R10779 gnd.n7261 gnd.n201 585
R10780 gnd.n202 gnd.n201 585
R10781 gnd.n7262 gnd.n210 585
R10782 gnd.n7485 gnd.n210 585
R10783 gnd.n7264 gnd.n7263 585
R10784 gnd.n7263 gnd.n209 585
R10785 gnd.n7265 gnd.n219 585
R10786 gnd.n7409 gnd.n219 585
R10787 gnd.n7267 gnd.n7266 585
R10788 gnd.n7266 gnd.n228 585
R10789 gnd.n7268 gnd.n226 585
R10790 gnd.n7401 gnd.n226 585
R10791 gnd.n7270 gnd.n7269 585
R10792 gnd.n7269 gnd.n225 585
R10793 gnd.n7271 gnd.n235 585
R10794 gnd.n7393 gnd.n235 585
R10795 gnd.n7273 gnd.n7272 585
R10796 gnd.n7272 gnd.n234 585
R10797 gnd.n7274 gnd.n242 585
R10798 gnd.n7385 gnd.n242 585
R10799 gnd.n7276 gnd.n7275 585
R10800 gnd.n7275 gnd.n250 585
R10801 gnd.n7277 gnd.n249 585
R10802 gnd.n7377 gnd.n249 585
R10803 gnd.n7279 gnd.n7278 585
R10804 gnd.n7278 gnd.n259 585
R10805 gnd.n7280 gnd.n257 585
R10806 gnd.n7369 gnd.n257 585
R10807 gnd.n7282 gnd.n7281 585
R10808 gnd.n7281 gnd.n256 585
R10809 gnd.n7283 gnd.n266 585
R10810 gnd.n7361 gnd.n266 585
R10811 gnd.n7285 gnd.n7284 585
R10812 gnd.n7284 gnd.n265 585
R10813 gnd.n7286 gnd.n272 585
R10814 gnd.n7353 gnd.n272 585
R10815 gnd.n7288 gnd.n7287 585
R10816 gnd.n7287 gnd.n280 585
R10817 gnd.n7289 gnd.n279 585
R10818 gnd.n7345 gnd.n279 585
R10819 gnd.n7291 gnd.n7290 585
R10820 gnd.n7290 gnd.n289 585
R10821 gnd.n7292 gnd.n287 585
R10822 gnd.n7337 gnd.n287 585
R10823 gnd.n7294 gnd.n7293 585
R10824 gnd.n7293 gnd.n286 585
R10825 gnd.n7295 gnd.n296 585
R10826 gnd.n7329 gnd.n296 585
R10827 gnd.n7297 gnd.n7296 585
R10828 gnd.n7296 gnd.n295 585
R10829 gnd.n7298 gnd.n324 585
R10830 gnd.n7305 gnd.n324 585
R10831 gnd.n7300 gnd.n7299 585
R10832 gnd.n7301 gnd.n7300 585
R10833 gnd.n332 gnd.n331 585
R10834 gnd.n331 gnd.n330 585
R10835 gnd.n7230 gnd.n7229 585
R10836 gnd.n7229 gnd.n7228 585
R10837 gnd.n335 gnd.n334 585
R10838 gnd.n336 gnd.n335 585
R10839 gnd.n7199 gnd.n339 585
R10840 gnd.n7222 gnd.n339 585
R10841 gnd.n7201 gnd.n7200 585
R10842 gnd.n7202 gnd.n7201 585
R10843 gnd.n355 gnd.n309 585
R10844 gnd.n7320 gnd.n309 585
R10845 gnd.n7194 gnd.n350 585
R10846 gnd.n7211 gnd.n350 585
R10847 gnd.n7193 gnd.n7192 585
R10848 gnd.n7192 gnd.n349 585
R10849 gnd.n7191 gnd.n357 585
R10850 gnd.n7191 gnd.n7190 585
R10851 gnd.n6929 gnd.n358 585
R10852 gnd.n7169 gnd.n358 585
R10853 gnd.n6932 gnd.n6931 585
R10854 gnd.n6931 gnd.n6930 585
R10855 gnd.n6933 gnd.n370 585
R10856 gnd.n7181 gnd.n370 585
R10857 gnd.n6934 gnd.n387 585
R10858 gnd.n7159 gnd.n387 585
R10859 gnd.n6935 gnd.n394 585
R10860 gnd.n7138 gnd.n394 585
R10861 gnd.n6937 gnd.n6936 585
R10862 gnd.n6938 gnd.n6937 585
R10863 gnd.n585 gnd.n402 585
R10864 gnd.n7130 gnd.n402 585
R10865 gnd.n6919 gnd.n6918 585
R10866 gnd.n6918 gnd.n6917 585
R10867 gnd.n587 gnd.n413 585
R10868 gnd.n7119 gnd.n413 585
R10869 gnd.n6900 gnd.n6899 585
R10870 gnd.n6899 gnd.n6898 585
R10871 gnd.n6901 gnd.n420 585
R10872 gnd.n7111 gnd.n420 585
R10873 gnd.n6903 gnd.n6902 585
R10874 gnd.n6904 gnd.n6903 585
R10875 gnd.n594 gnd.n429 585
R10876 gnd.n7103 gnd.n429 585
R10877 gnd.n6892 gnd.n6891 585
R10878 gnd.n6891 gnd.n6890 585
R10879 gnd.n6889 gnd.n438 585
R10880 gnd.n7095 gnd.n438 585
R10881 gnd.n6888 gnd.n6887 585
R10882 gnd.n6887 gnd.n6886 585
R10883 gnd.n596 gnd.n447 585
R10884 gnd.n7087 gnd.n447 585
R10885 gnd.n6861 gnd.n6860 585
R10886 gnd.n6860 gnd.n6859 585
R10887 gnd.n6862 gnd.n454 585
R10888 gnd.n7079 gnd.n454 585
R10889 gnd.n6864 gnd.n6863 585
R10890 gnd.n6865 gnd.n6864 585
R10891 gnd.n6841 gnd.n463 585
R10892 gnd.n7071 gnd.n463 585
R10893 gnd.n6852 gnd.n6851 585
R10894 gnd.n6851 gnd.n6850 585
R10895 gnd.n6849 gnd.n472 585
R10896 gnd.n7063 gnd.n472 585
R10897 gnd.n6848 gnd.n6847 585
R10898 gnd.n6847 gnd.n6846 585
R10899 gnd.n6843 gnd.n481 585
R10900 gnd.n7055 gnd.n481 585
R10901 gnd.n6975 gnd.n563 585
R10902 gnd.n6975 gnd.n6974 585
R10903 gnd.n675 gnd.n674 585
R10904 gnd.n675 gnd.n646 585
R10905 gnd.n6771 gnd.n6770 585
R10906 gnd.n6770 gnd.n6769 585
R10907 gnd.n6772 gnd.n672 585
R10908 gnd.n672 gnd.n655 585
R10909 gnd.n6774 gnd.n6773 585
R10910 gnd.n6775 gnd.n6774 585
R10911 gnd.n673 gnd.n671 585
R10912 gnd.n671 gnd.n670 585
R10913 gnd.n6573 gnd.n661 585
R10914 gnd.n6781 gnd.n661 585
R10915 gnd.n6575 gnd.n6574 585
R10916 gnd.n6576 gnd.n6575 585
R10917 gnd.n6572 gnd.n899 585
R10918 gnd.n899 gnd.n898 585
R10919 gnd.n6571 gnd.n6570 585
R10920 gnd.n6570 gnd.n6569 585
R10921 gnd.n901 gnd.n900 585
R10922 gnd.n901 gnd.n880 585
R10923 gnd.n6557 gnd.n908 585
R10924 gnd.n908 gnd.n879 585
R10925 gnd.n6559 gnd.n6558 585
R10926 gnd.n6560 gnd.n6559 585
R10927 gnd.n6556 gnd.n907 585
R10928 gnd.n907 gnd.n890 585
R10929 gnd.n6555 gnd.n6554 585
R10930 gnd.n6554 gnd.n888 585
R10931 gnd.n6553 gnd.n909 585
R10932 gnd.n6553 gnd.n6552 585
R10933 gnd.n6227 gnd.n910 585
R10934 gnd.n911 gnd.n910 585
R10935 gnd.n6228 gnd.n6226 585
R10936 gnd.n6226 gnd.n920 585
R10937 gnd.n6230 gnd.n6229 585
R10938 gnd.n6230 gnd.n919 585
R10939 gnd.n6231 gnd.n6225 585
R10940 gnd.n6372 gnd.n6231 585
R10941 gnd.n6376 gnd.n6375 585
R10942 gnd.n6375 gnd.n6374 585
R10943 gnd.n6377 gnd.n6223 585
R10944 gnd.n6223 gnd.n928 585
R10945 gnd.n6379 gnd.n6378 585
R10946 gnd.n6380 gnd.n6379 585
R10947 gnd.n6224 gnd.n6222 585
R10948 gnd.n6222 gnd.n939 585
R10949 gnd.n6349 gnd.n6239 585
R10950 gnd.n6239 gnd.n937 585
R10951 gnd.n6351 gnd.n6350 585
R10952 gnd.n6352 gnd.n6351 585
R10953 gnd.n6348 gnd.n6238 585
R10954 gnd.n6238 gnd.n947 585
R10955 gnd.n6347 gnd.n6346 585
R10956 gnd.n6346 gnd.n945 585
R10957 gnd.n6345 gnd.n6240 585
R10958 gnd.n6345 gnd.n6344 585
R10959 gnd.n6331 gnd.n6241 585
R10960 gnd.n6241 gnd.n955 585
R10961 gnd.n6332 gnd.n6249 585
R10962 gnd.n6249 gnd.n953 585
R10963 gnd.n6334 gnd.n6333 585
R10964 gnd.n6335 gnd.n6334 585
R10965 gnd.n6330 gnd.n6248 585
R10966 gnd.n6248 gnd.n6247 585
R10967 gnd.n6329 gnd.n6328 585
R10968 gnd.n6328 gnd.n961 585
R10969 gnd.n6327 gnd.n6250 585
R10970 gnd.n6327 gnd.n6326 585
R10971 gnd.n6312 gnd.n6251 585
R10972 gnd.n6251 gnd.n970 585
R10973 gnd.n6313 gnd.n6259 585
R10974 gnd.n6259 gnd.n968 585
R10975 gnd.n6315 gnd.n6314 585
R10976 gnd.n6316 gnd.n6315 585
R10977 gnd.n6311 gnd.n6258 585
R10978 gnd.n6258 gnd.n6256 585
R10979 gnd.n6310 gnd.n6309 585
R10980 gnd.n6309 gnd.n976 585
R10981 gnd.n6308 gnd.n6260 585
R10982 gnd.n6308 gnd.n6307 585
R10983 gnd.n6295 gnd.n6261 585
R10984 gnd.n6261 gnd.n984 585
R10985 gnd.n6297 gnd.n6296 585
R10986 gnd.n6298 gnd.n6297 585
R10987 gnd.n6294 gnd.n6268 585
R10988 gnd.n6268 gnd.n6267 585
R10989 gnd.n6293 gnd.n6292 585
R10990 gnd.n6292 gnd.n992 585
R10991 gnd.n6291 gnd.n6269 585
R10992 gnd.n6291 gnd.n990 585
R10993 gnd.n6290 gnd.n6273 585
R10994 gnd.n6290 gnd.n6289 585
R10995 gnd.n6272 gnd.n6270 585
R10996 gnd.n6270 gnd.n1000 585
R10997 gnd.n6271 gnd.n1038 585
R10998 gnd.n1038 gnd.n998 585
R10999 gnd.n6416 gnd.n1037 585
R11000 gnd.n6416 gnd.n6415 585
R11001 gnd.n6418 gnd.n6417 585
R11002 gnd.n6417 gnd.n1008 585
R11003 gnd.n6419 gnd.n1035 585
R11004 gnd.n1035 gnd.n1006 585
R11005 gnd.n6421 gnd.n6420 585
R11006 gnd.n6422 gnd.n6421 585
R11007 gnd.n1036 gnd.n1034 585
R11008 gnd.n1034 gnd.n1016 585
R11009 gnd.n1170 gnd.n1169 585
R11010 gnd.n1170 gnd.n1014 585
R11011 gnd.n1172 gnd.n1171 585
R11012 gnd.n1171 gnd.n1025 585
R11013 gnd.n1173 gnd.n1023 585
R11014 gnd.n6430 gnd.n1023 585
R11015 gnd.n1175 gnd.n1174 585
R11016 gnd.n1174 gnd.n1022 585
R11017 gnd.n1176 gnd.n1165 585
R11018 gnd.n1165 gnd.n1049 585
R11019 gnd.n1178 gnd.n1177 585
R11020 gnd.n1179 gnd.n1178 585
R11021 gnd.n1168 gnd.n1164 585
R11022 gnd.n1164 gnd.n1058 585
R11023 gnd.n1167 gnd.n1166 585
R11024 gnd.n1166 gnd.n1056 585
R11025 gnd.n1156 gnd.n1155 585
R11026 gnd.n6080 gnd.n1156 585
R11027 gnd.n6083 gnd.n6082 585
R11028 gnd.n6082 gnd.n6081 585
R11029 gnd.n6084 gnd.n1152 585
R11030 gnd.n1152 gnd.n1065 585
R11031 gnd.n6086 gnd.n6085 585
R11032 gnd.n6087 gnd.n6086 585
R11033 gnd.n1154 gnd.n1151 585
R11034 gnd.n1151 gnd.n1149 585
R11035 gnd.n1153 gnd.n1140 585
R11036 gnd.n6093 gnd.n1140 585
R11037 gnd.n6096 gnd.n1139 585
R11038 gnd.n6096 gnd.n6095 585
R11039 gnd.n6098 gnd.n6097 585
R11040 gnd.n6097 gnd.n1080 585
R11041 gnd.n6099 gnd.n1136 585
R11042 gnd.n1136 gnd.n1078 585
R11043 gnd.n6101 gnd.n6100 585
R11044 gnd.n6102 gnd.n6101 585
R11045 gnd.n1138 gnd.n1135 585
R11046 gnd.n1135 gnd.n1087 585
R11047 gnd.n1137 gnd.n1124 585
R11048 gnd.n6108 gnd.n1124 585
R11049 gnd.n6111 gnd.n1123 585
R11050 gnd.n6111 gnd.n6110 585
R11051 gnd.n6113 gnd.n6112 585
R11052 gnd.n6112 gnd.n1095 585
R11053 gnd.n6114 gnd.n1121 585
R11054 gnd.n1121 gnd.n1093 585
R11055 gnd.n6116 gnd.n6115 585
R11056 gnd.n6117 gnd.n6116 585
R11057 gnd.n1122 gnd.n1120 585
R11058 gnd.n1120 gnd.n1103 585
R11059 gnd.n5871 gnd.n5870 585
R11060 gnd.n5871 gnd.n1101 585
R11061 gnd.n5873 gnd.n5872 585
R11062 gnd.n5872 gnd.n1111 585
R11063 gnd.n5874 gnd.n1109 585
R11064 gnd.n6125 gnd.n1109 585
R11065 gnd.n5875 gnd.n5869 585
R11066 gnd.n5869 gnd.n1200 585
R11067 gnd.n5877 gnd.n5876 585
R11068 gnd.n5877 gnd.n1199 585
R11069 gnd.n5941 gnd.n5868 585
R11070 gnd.n5941 gnd.n5940 585
R11071 gnd.n5943 gnd.n5942 585
R11072 gnd.n5942 gnd.n1209 585
R11073 gnd.n5944 gnd.n5866 585
R11074 gnd.n5866 gnd.n1207 585
R11075 gnd.n5946 gnd.n5945 585
R11076 gnd.n5947 gnd.n5946 585
R11077 gnd.n5867 gnd.n5865 585
R11078 gnd.n5865 gnd.n1218 585
R11079 gnd.n5924 gnd.n5885 585
R11080 gnd.n5885 gnd.n1216 585
R11081 gnd.n5926 gnd.n5925 585
R11082 gnd.n5927 gnd.n5926 585
R11083 gnd.n5923 gnd.n5884 585
R11084 gnd.n5884 gnd.n1225 585
R11085 gnd.n5922 gnd.n5921 585
R11086 gnd.n5921 gnd.n5920 585
R11087 gnd.n5887 gnd.n5886 585
R11088 gnd.n5889 gnd.n5887 585
R11089 gnd.n5907 gnd.n5906 585
R11090 gnd.n5906 gnd.n1233 585
R11091 gnd.n5908 gnd.n5903 585
R11092 gnd.n5903 gnd.n1231 585
R11093 gnd.n5910 gnd.n5909 585
R11094 gnd.n5911 gnd.n5910 585
R11095 gnd.n5905 gnd.n5902 585
R11096 gnd.n5902 gnd.n1241 585
R11097 gnd.n5904 gnd.n1276 585
R11098 gnd.n1276 gnd.n1239 585
R11099 gnd.n5969 gnd.n1275 585
R11100 gnd.n5969 gnd.n5968 585
R11101 gnd.n5971 gnd.n5970 585
R11102 gnd.n5970 gnd.n1248 585
R11103 gnd.n5972 gnd.n1273 585
R11104 gnd.n5852 gnd.n1273 585
R11105 gnd.n5974 gnd.n5973 585
R11106 gnd.n5975 gnd.n5974 585
R11107 gnd.n1274 gnd.n1272 585
R11108 gnd.n1272 gnd.n1256 585
R11109 gnd.n1521 gnd.n1520 585
R11110 gnd.n1521 gnd.n1254 585
R11111 gnd.n1523 gnd.n1522 585
R11112 gnd.n1522 gnd.n1264 585
R11113 gnd.n1524 gnd.n1262 585
R11114 gnd.n5983 gnd.n1262 585
R11115 gnd.n1526 gnd.n1525 585
R11116 gnd.n1525 gnd.n1288 585
R11117 gnd.n1527 gnd.n1413 585
R11118 gnd.n1413 gnd.n1287 585
R11119 gnd.n1529 gnd.n1528 585
R11120 gnd.n1530 gnd.n1529 585
R11121 gnd.n1519 gnd.n1412 585
R11122 gnd.n1412 gnd.n1297 585
R11123 gnd.n1518 gnd.n1517 585
R11124 gnd.n1517 gnd.n1295 585
R11125 gnd.n1516 gnd.n1515 585
R11126 gnd.n1514 gnd.n1513 585
R11127 gnd.n1512 gnd.n1436 585
R11128 gnd.n1512 gnd.n1305 585
R11129 gnd.n1511 gnd.n1510 585
R11130 gnd.n1509 gnd.n1508 585
R11131 gnd.n1507 gnd.n1438 585
R11132 gnd.n1505 gnd.n1504 585
R11133 gnd.n1503 gnd.n1439 585
R11134 gnd.n1502 gnd.n1501 585
R11135 gnd.n1499 gnd.n1440 585
R11136 gnd.n1497 gnd.n1496 585
R11137 gnd.n1495 gnd.n1441 585
R11138 gnd.n1494 gnd.n1493 585
R11139 gnd.n1491 gnd.n1442 585
R11140 gnd.n1489 gnd.n1488 585
R11141 gnd.n1487 gnd.n1443 585
R11142 gnd.n1486 gnd.n1485 585
R11143 gnd.n1483 gnd.n1444 585
R11144 gnd.n1481 gnd.n1480 585
R11145 gnd.n1479 gnd.n1445 585
R11146 gnd.n1478 gnd.n1477 585
R11147 gnd.n1475 gnd.n1446 585
R11148 gnd.n1473 gnd.n1472 585
R11149 gnd.n1471 gnd.n1447 585
R11150 gnd.n1470 gnd.n1469 585
R11151 gnd.n1467 gnd.n1448 585
R11152 gnd.n1465 gnd.n1464 585
R11153 gnd.n1463 gnd.n1449 585
R11154 gnd.n1462 gnd.n1461 585
R11155 gnd.n1459 gnd.n1458 585
R11156 gnd.n1457 gnd.n1456 585
R11157 gnd.n1455 gnd.n1391 585
R11158 gnd.n1605 gnd.n1604 585
R11159 gnd.n1602 gnd.n1390 585
R11160 gnd.n1600 gnd.n1599 585
R11161 gnd.n1598 gnd.n1393 585
R11162 gnd.n1596 gnd.n1595 585
R11163 gnd.n1593 gnd.n1396 585
R11164 gnd.n1591 gnd.n1590 585
R11165 gnd.n1589 gnd.n1397 585
R11166 gnd.n1588 gnd.n1587 585
R11167 gnd.n1585 gnd.n1398 585
R11168 gnd.n1583 gnd.n1582 585
R11169 gnd.n1581 gnd.n1399 585
R11170 gnd.n1580 gnd.n1579 585
R11171 gnd.n1577 gnd.n1400 585
R11172 gnd.n1575 gnd.n1574 585
R11173 gnd.n1573 gnd.n1401 585
R11174 gnd.n1572 gnd.n1571 585
R11175 gnd.n1569 gnd.n1402 585
R11176 gnd.n1567 gnd.n1566 585
R11177 gnd.n1565 gnd.n1403 585
R11178 gnd.n1564 gnd.n1563 585
R11179 gnd.n1561 gnd.n1404 585
R11180 gnd.n1559 gnd.n1558 585
R11181 gnd.n1557 gnd.n1405 585
R11182 gnd.n1556 gnd.n1555 585
R11183 gnd.n1553 gnd.n1406 585
R11184 gnd.n1551 gnd.n1550 585
R11185 gnd.n1549 gnd.n1407 585
R11186 gnd.n1548 gnd.n1547 585
R11187 gnd.n1545 gnd.n1408 585
R11188 gnd.n1543 gnd.n1542 585
R11189 gnd.n1541 gnd.n1409 585
R11190 gnd.n1540 gnd.n1539 585
R11191 gnd.n866 gnd.n865 585
R11192 gnd.n863 gnd.n677 585
R11193 gnd.n862 gnd.n861 585
R11194 gnd.n860 gnd.n859 585
R11195 gnd.n858 gnd.n679 585
R11196 gnd.n856 gnd.n855 585
R11197 gnd.n854 gnd.n680 585
R11198 gnd.n853 gnd.n852 585
R11199 gnd.n850 gnd.n681 585
R11200 gnd.n848 gnd.n847 585
R11201 gnd.n846 gnd.n682 585
R11202 gnd.n845 gnd.n844 585
R11203 gnd.n842 gnd.n683 585
R11204 gnd.n840 gnd.n839 585
R11205 gnd.n838 gnd.n684 585
R11206 gnd.n837 gnd.n836 585
R11207 gnd.n834 gnd.n685 585
R11208 gnd.n832 gnd.n831 585
R11209 gnd.n830 gnd.n686 585
R11210 gnd.n829 gnd.n828 585
R11211 gnd.n826 gnd.n687 585
R11212 gnd.n824 gnd.n823 585
R11213 gnd.n822 gnd.n688 585
R11214 gnd.n821 gnd.n820 585
R11215 gnd.n818 gnd.n689 585
R11216 gnd.n816 gnd.n815 585
R11217 gnd.n814 gnd.n690 585
R11218 gnd.n813 gnd.n812 585
R11219 gnd.n810 gnd.n691 585
R11220 gnd.n808 gnd.n807 585
R11221 gnd.n803 gnd.n692 585
R11222 gnd.n802 gnd.n801 585
R11223 gnd.n799 gnd.n648 585
R11224 gnd.n796 gnd.n534 585
R11225 gnd.n795 gnd.n794 585
R11226 gnd.n793 gnd.n792 585
R11227 gnd.n791 gnd.n694 585
R11228 gnd.n789 gnd.n788 585
R11229 gnd.n784 gnd.n695 585
R11230 gnd.n783 gnd.n782 585
R11231 gnd.n780 gnd.n696 585
R11232 gnd.n778 gnd.n777 585
R11233 gnd.n776 gnd.n697 585
R11234 gnd.n775 gnd.n774 585
R11235 gnd.n772 gnd.n698 585
R11236 gnd.n770 gnd.n769 585
R11237 gnd.n768 gnd.n699 585
R11238 gnd.n767 gnd.n766 585
R11239 gnd.n764 gnd.n700 585
R11240 gnd.n762 gnd.n761 585
R11241 gnd.n760 gnd.n701 585
R11242 gnd.n759 gnd.n758 585
R11243 gnd.n756 gnd.n702 585
R11244 gnd.n754 gnd.n753 585
R11245 gnd.n752 gnd.n703 585
R11246 gnd.n751 gnd.n750 585
R11247 gnd.n748 gnd.n704 585
R11248 gnd.n746 gnd.n745 585
R11249 gnd.n744 gnd.n705 585
R11250 gnd.n743 gnd.n742 585
R11251 gnd.n740 gnd.n706 585
R11252 gnd.n738 gnd.n737 585
R11253 gnd.n736 gnd.n707 585
R11254 gnd.n735 gnd.n734 585
R11255 gnd.n732 gnd.n708 585
R11256 gnd.n730 gnd.n729 585
R11257 gnd.n867 gnd.n676 585
R11258 gnd.n676 gnd.n646 585
R11259 gnd.n869 gnd.n868 585
R11260 gnd.n6769 gnd.n869 585
R11261 gnd.n668 gnd.n667 585
R11262 gnd.n668 gnd.n655 585
R11263 gnd.n6777 gnd.n6776 585
R11264 gnd.n6776 gnd.n6775 585
R11265 gnd.n6778 gnd.n665 585
R11266 gnd.n670 gnd.n665 585
R11267 gnd.n6780 gnd.n6779 585
R11268 gnd.n6781 gnd.n6780 585
R11269 gnd.n666 gnd.n664 585
R11270 gnd.n6576 gnd.n664 585
R11271 gnd.n6565 gnd.n903 585
R11272 gnd.n903 gnd.n898 585
R11273 gnd.n6567 gnd.n6566 585
R11274 gnd.n6569 gnd.n6567 585
R11275 gnd.n6564 gnd.n902 585
R11276 gnd.n902 gnd.n880 585
R11277 gnd.n6563 gnd.n6562 585
R11278 gnd.n6562 gnd.n879 585
R11279 gnd.n6561 gnd.n904 585
R11280 gnd.n6561 gnd.n6560 585
R11281 gnd.n6361 gnd.n905 585
R11282 gnd.n905 gnd.n890 585
R11283 gnd.n6363 gnd.n6362 585
R11284 gnd.n6362 gnd.n888 585
R11285 gnd.n6364 gnd.n912 585
R11286 gnd.n6552 gnd.n912 585
R11287 gnd.n6366 gnd.n6365 585
R11288 gnd.n6366 gnd.n911 585
R11289 gnd.n6368 gnd.n6367 585
R11290 gnd.n6367 gnd.n920 585
R11291 gnd.n6369 gnd.n6233 585
R11292 gnd.n6233 gnd.n919 585
R11293 gnd.n6371 gnd.n6370 585
R11294 gnd.n6372 gnd.n6371 585
R11295 gnd.n6360 gnd.n6232 585
R11296 gnd.n6374 gnd.n6232 585
R11297 gnd.n6359 gnd.n6358 585
R11298 gnd.n6358 gnd.n928 585
R11299 gnd.n6357 gnd.n6221 585
R11300 gnd.n6380 gnd.n6221 585
R11301 gnd.n6356 gnd.n6355 585
R11302 gnd.n6355 gnd.n939 585
R11303 gnd.n6354 gnd.n6234 585
R11304 gnd.n6354 gnd.n937 585
R11305 gnd.n6353 gnd.n6236 585
R11306 gnd.n6353 gnd.n6352 585
R11307 gnd.n6340 gnd.n6235 585
R11308 gnd.n6235 gnd.n947 585
R11309 gnd.n6341 gnd.n6244 585
R11310 gnd.n6244 gnd.n945 585
R11311 gnd.n6343 gnd.n6342 585
R11312 gnd.n6344 gnd.n6343 585
R11313 gnd.n6339 gnd.n6243 585
R11314 gnd.n6243 gnd.n955 585
R11315 gnd.n6338 gnd.n6337 585
R11316 gnd.n6337 gnd.n953 585
R11317 gnd.n6336 gnd.n6245 585
R11318 gnd.n6336 gnd.n6335 585
R11319 gnd.n6321 gnd.n6246 585
R11320 gnd.n6247 gnd.n6246 585
R11321 gnd.n6322 gnd.n6253 585
R11322 gnd.n6253 gnd.n961 585
R11323 gnd.n6324 gnd.n6323 585
R11324 gnd.n6326 gnd.n6324 585
R11325 gnd.n6320 gnd.n6252 585
R11326 gnd.n6252 gnd.n970 585
R11327 gnd.n6319 gnd.n6318 585
R11328 gnd.n6318 gnd.n968 585
R11329 gnd.n6317 gnd.n6254 585
R11330 gnd.n6317 gnd.n6316 585
R11331 gnd.n6302 gnd.n6255 585
R11332 gnd.n6256 gnd.n6255 585
R11333 gnd.n6303 gnd.n6263 585
R11334 gnd.n6263 gnd.n976 585
R11335 gnd.n6305 gnd.n6304 585
R11336 gnd.n6307 gnd.n6305 585
R11337 gnd.n6301 gnd.n6262 585
R11338 gnd.n6262 gnd.n984 585
R11339 gnd.n6300 gnd.n6299 585
R11340 gnd.n6299 gnd.n6298 585
R11341 gnd.n6265 gnd.n6264 585
R11342 gnd.n6267 gnd.n6265 585
R11343 gnd.n6284 gnd.n6283 585
R11344 gnd.n6283 gnd.n992 585
R11345 gnd.n6285 gnd.n6275 585
R11346 gnd.n6275 gnd.n990 585
R11347 gnd.n6287 gnd.n6286 585
R11348 gnd.n6289 gnd.n6287 585
R11349 gnd.n6282 gnd.n6274 585
R11350 gnd.n6274 gnd.n1000 585
R11351 gnd.n6281 gnd.n6280 585
R11352 gnd.n6280 gnd.n998 585
R11353 gnd.n6279 gnd.n1039 585
R11354 gnd.n6415 gnd.n1039 585
R11355 gnd.n6278 gnd.n6277 585
R11356 gnd.n6277 gnd.n1008 585
R11357 gnd.n6276 gnd.n1031 585
R11358 gnd.n1031 gnd.n1006 585
R11359 gnd.n6423 gnd.n1032 585
R11360 gnd.n6423 gnd.n6422 585
R11361 gnd.n6424 gnd.n1030 585
R11362 gnd.n6424 gnd.n1016 585
R11363 gnd.n6426 gnd.n6425 585
R11364 gnd.n6425 gnd.n1014 585
R11365 gnd.n6427 gnd.n1028 585
R11366 gnd.n1028 gnd.n1025 585
R11367 gnd.n6429 gnd.n6428 585
R11368 gnd.n6430 gnd.n6429 585
R11369 gnd.n1029 gnd.n1027 585
R11370 gnd.n1027 gnd.n1022 585
R11371 gnd.n1162 gnd.n1161 585
R11372 gnd.n1162 gnd.n1049 585
R11373 gnd.n1180 gnd.n1160 585
R11374 gnd.n1180 gnd.n1179 585
R11375 gnd.n1182 gnd.n1181 585
R11376 gnd.n1181 gnd.n1058 585
R11377 gnd.n1183 gnd.n1158 585
R11378 gnd.n1158 gnd.n1056 585
R11379 gnd.n1185 gnd.n1184 585
R11380 gnd.n6080 gnd.n1185 585
R11381 gnd.n1159 gnd.n1157 585
R11382 gnd.n6081 gnd.n1157 585
R11383 gnd.n1148 gnd.n1147 585
R11384 gnd.n1148 gnd.n1065 585
R11385 gnd.n6089 gnd.n6088 585
R11386 gnd.n6088 gnd.n6087 585
R11387 gnd.n6090 gnd.n1143 585
R11388 gnd.n1149 gnd.n1143 585
R11389 gnd.n6092 gnd.n6091 585
R11390 gnd.n6093 gnd.n6092 585
R11391 gnd.n1146 gnd.n1141 585
R11392 gnd.n6095 gnd.n1141 585
R11393 gnd.n1145 gnd.n1144 585
R11394 gnd.n1144 gnd.n1080 585
R11395 gnd.n1133 gnd.n1132 585
R11396 gnd.n1133 gnd.n1078 585
R11397 gnd.n6104 gnd.n6103 585
R11398 gnd.n6103 gnd.n6102 585
R11399 gnd.n6105 gnd.n1127 585
R11400 gnd.n1127 gnd.n1087 585
R11401 gnd.n6107 gnd.n6106 585
R11402 gnd.n6108 gnd.n6107 585
R11403 gnd.n1131 gnd.n1125 585
R11404 gnd.n6110 gnd.n1125 585
R11405 gnd.n1130 gnd.n1129 585
R11406 gnd.n1129 gnd.n1095 585
R11407 gnd.n1128 gnd.n1117 585
R11408 gnd.n1117 gnd.n1093 585
R11409 gnd.n6118 gnd.n1118 585
R11410 gnd.n6118 gnd.n6117 585
R11411 gnd.n6119 gnd.n1116 585
R11412 gnd.n6119 gnd.n1103 585
R11413 gnd.n6121 gnd.n6120 585
R11414 gnd.n6120 gnd.n1101 585
R11415 gnd.n6122 gnd.n1114 585
R11416 gnd.n1114 gnd.n1111 585
R11417 gnd.n6124 gnd.n6123 585
R11418 gnd.n6125 gnd.n6124 585
R11419 gnd.n1115 gnd.n1113 585
R11420 gnd.n1200 gnd.n1113 585
R11421 gnd.n5936 gnd.n5879 585
R11422 gnd.n5879 gnd.n1199 585
R11423 gnd.n5938 gnd.n5937 585
R11424 gnd.n5940 gnd.n5938 585
R11425 gnd.n5935 gnd.n5878 585
R11426 gnd.n5878 gnd.n1209 585
R11427 gnd.n5934 gnd.n5933 585
R11428 gnd.n5933 gnd.n1207 585
R11429 gnd.n5932 gnd.n5864 585
R11430 gnd.n5947 gnd.n5864 585
R11431 gnd.n5931 gnd.n5930 585
R11432 gnd.n5930 gnd.n1218 585
R11433 gnd.n5929 gnd.n5880 585
R11434 gnd.n5929 gnd.n1216 585
R11435 gnd.n5928 gnd.n5882 585
R11436 gnd.n5928 gnd.n5927 585
R11437 gnd.n5917 gnd.n5881 585
R11438 gnd.n5881 gnd.n1225 585
R11439 gnd.n5919 gnd.n5918 585
R11440 gnd.n5920 gnd.n5919 585
R11441 gnd.n5916 gnd.n5890 585
R11442 gnd.n5890 gnd.n5889 585
R11443 gnd.n5915 gnd.n5914 585
R11444 gnd.n5914 gnd.n1233 585
R11445 gnd.n5913 gnd.n5891 585
R11446 gnd.n5913 gnd.n1231 585
R11447 gnd.n5912 gnd.n5900 585
R11448 gnd.n5912 gnd.n5911 585
R11449 gnd.n5899 gnd.n5892 585
R11450 gnd.n5892 gnd.n1241 585
R11451 gnd.n5898 gnd.n5897 585
R11452 gnd.n5897 gnd.n1239 585
R11453 gnd.n5896 gnd.n1277 585
R11454 gnd.n5968 gnd.n1277 585
R11455 gnd.n5895 gnd.n5894 585
R11456 gnd.n5894 gnd.n1248 585
R11457 gnd.n5893 gnd.n1270 585
R11458 gnd.n5852 gnd.n1270 585
R11459 gnd.n5976 gnd.n1271 585
R11460 gnd.n5976 gnd.n5975 585
R11461 gnd.n5977 gnd.n1269 585
R11462 gnd.n5977 gnd.n1256 585
R11463 gnd.n5979 gnd.n5978 585
R11464 gnd.n5978 gnd.n1254 585
R11465 gnd.n5980 gnd.n1267 585
R11466 gnd.n1267 gnd.n1264 585
R11467 gnd.n5982 gnd.n5981 585
R11468 gnd.n5983 gnd.n5982 585
R11469 gnd.n1268 gnd.n1266 585
R11470 gnd.n1288 gnd.n1266 585
R11471 gnd.n1533 gnd.n1532 585
R11472 gnd.n1532 gnd.n1287 585
R11473 gnd.n1534 gnd.n1531 585
R11474 gnd.n1531 gnd.n1530 585
R11475 gnd.n1536 gnd.n1535 585
R11476 gnd.n1536 gnd.n1297 585
R11477 gnd.n1537 gnd.n1410 585
R11478 gnd.n1537 gnd.n1295 585
R11479 gnd.n3351 gnd.n2064 585
R11480 gnd.n2064 gnd.n1788 585
R11481 gnd.n7220 gnd.n7219 585
R11482 gnd.n7221 gnd.n7220 585
R11483 gnd.n7216 gnd.n343 585
R11484 gnd.n343 gnd.n311 585
R11485 gnd.n7215 gnd.n7214 585
R11486 gnd.n7214 gnd.n308 585
R11487 gnd.n7213 gnd.n346 585
R11488 gnd.n7213 gnd.n7212 585
R11489 gnd.n7150 gnd.n348 585
R11490 gnd.n361 gnd.n348 585
R11491 gnd.n7152 gnd.n7151 585
R11492 gnd.n7152 gnd.n359 585
R11493 gnd.n7154 gnd.n7153 585
R11494 gnd.n7153 gnd.n379 585
R11495 gnd.n7155 gnd.n389 585
R11496 gnd.n389 gnd.n372 585
R11497 gnd.n7157 gnd.n7156 585
R11498 gnd.n7158 gnd.n7157 585
R11499 gnd.n390 gnd.n388 585
R11500 gnd.n388 gnd.n386 585
R11501 gnd.n7141 gnd.n7140 585
R11502 gnd.n7140 gnd.n7139 585
R11503 gnd.n393 gnd.n392 585
R11504 gnd.n404 gnd.n393 585
R11505 gnd.n6913 gnd.n589 585
R11506 gnd.n589 gnd.n401 585
R11507 gnd.n6915 gnd.n6914 585
R11508 gnd.n6916 gnd.n6915 585
R11509 gnd.n590 gnd.n588 585
R11510 gnd.n588 gnd.n412 585
R11511 gnd.n6908 gnd.n6907 585
R11512 gnd.n6907 gnd.n422 585
R11513 gnd.n6906 gnd.n592 585
R11514 gnd.n6906 gnd.n6905 585
R11515 gnd.n6877 gnd.n593 585
R11516 gnd.n593 gnd.n431 585
R11517 gnd.n6879 gnd.n6878 585
R11518 gnd.n6879 gnd.n428 585
R11519 gnd.n6881 gnd.n6880 585
R11520 gnd.n6880 gnd.n440 585
R11521 gnd.n6882 gnd.n599 585
R11522 gnd.n599 gnd.n437 585
R11523 gnd.n6884 gnd.n6883 585
R11524 gnd.n6885 gnd.n6884 585
R11525 gnd.n600 gnd.n598 585
R11526 gnd.n598 gnd.n446 585
R11527 gnd.n6869 gnd.n6868 585
R11528 gnd.n6868 gnd.n456 585
R11529 gnd.n6867 gnd.n602 585
R11530 gnd.n6867 gnd.n6866 585
R11531 gnd.n6840 gnd.n6839 585
R11532 gnd.n6840 gnd.n465 585
R11533 gnd.n604 gnd.n603 585
R11534 gnd.n603 gnd.n462 585
R11535 gnd.n6835 gnd.n6834 585
R11536 gnd.n6834 gnd.n474 585
R11537 gnd.n6833 gnd.n606 585
R11538 gnd.n6833 gnd.n471 585
R11539 gnd.n6832 gnd.n6831 585
R11540 gnd.n6832 gnd.n483 585
R11541 gnd.n608 gnd.n607 585
R11542 gnd.n607 gnd.n480 585
R11543 gnd.n6827 gnd.n6826 585
R11544 gnd.n6826 gnd.n564 585
R11545 gnd.n6825 gnd.n610 585
R11546 gnd.n6825 gnd.n518 585
R11547 gnd.n6824 gnd.n6823 585
R11548 gnd.n6824 gnd.n489 585
R11549 gnd.n612 gnd.n611 585
R11550 gnd.n6816 gnd.n611 585
R11551 gnd.n6819 gnd.n6818 585
R11552 gnd.n6818 gnd.n6817 585
R11553 gnd.n615 gnd.n614 585
R11554 gnd.n616 gnd.n615 585
R11555 gnd.n6805 gnd.n641 585
R11556 gnd.n641 gnd.n639 585
R11557 gnd.n6807 gnd.n6806 585
R11558 gnd.n6808 gnd.n6807 585
R11559 gnd.n642 gnd.n640 585
R11560 gnd.n6613 gnd.n640 585
R11561 gnd.n6800 gnd.n6799 585
R11562 gnd.n6799 gnd.n6798 585
R11563 gnd.n645 gnd.n644 585
R11564 gnd.n6768 gnd.n645 585
R11565 gnd.n6788 gnd.n6787 585
R11566 gnd.n6789 gnd.n6788 585
R11567 gnd.n657 gnd.n656 585
R11568 gnd.n669 gnd.n656 585
R11569 gnd.n6783 gnd.n6782 585
R11570 gnd.n6782 gnd.n6781 585
R11571 gnd.n660 gnd.n659 585
R11572 gnd.n6577 gnd.n660 585
R11573 gnd.n6597 gnd.n883 585
R11574 gnd.n6568 gnd.n883 585
R11575 gnd.n6599 gnd.n6598 585
R11576 gnd.n6600 gnd.n6599 585
R11577 gnd.n884 gnd.n882 585
R11578 gnd.n906 gnd.n882 585
R11579 gnd.n6592 gnd.n6591 585
R11580 gnd.n6591 gnd.n6590 585
R11581 gnd.n887 gnd.n886 585
R11582 gnd.n6551 gnd.n887 585
R11583 gnd.n6539 gnd.n923 585
R11584 gnd.n6523 gnd.n923 585
R11585 gnd.n6541 gnd.n6540 585
R11586 gnd.n6542 gnd.n6541 585
R11587 gnd.n924 gnd.n922 585
R11588 gnd.n6373 gnd.n922 585
R11589 gnd.n6534 gnd.n6533 585
R11590 gnd.n6533 gnd.n6532 585
R11591 gnd.n927 gnd.n926 585
R11592 gnd.n6381 gnd.n927 585
R11593 gnd.n6517 gnd.n6516 585
R11594 gnd.t4 gnd.n6517 585
R11595 gnd.n941 gnd.n940 585
R11596 gnd.n6237 gnd.n940 585
R11597 gnd.n6512 gnd.n6511 585
R11598 gnd.n6511 gnd.n6510 585
R11599 gnd.n944 gnd.n943 585
R11600 gnd.n6242 gnd.n944 585
R11601 gnd.n6501 gnd.n6500 585
R11602 gnd.n6502 gnd.n6501 585
R11603 gnd.n957 gnd.n956 585
R11604 gnd.n6335 gnd.n956 585
R11605 gnd.n6496 gnd.n6495 585
R11606 gnd.n6495 gnd.n6494 585
R11607 gnd.n960 gnd.n959 585
R11608 gnd.n6325 gnd.n960 585
R11609 gnd.n6485 gnd.n6484 585
R11610 gnd.n6486 gnd.n6485 585
R11611 gnd.n972 gnd.n971 585
R11612 gnd.n6257 gnd.n971 585
R11613 gnd.n6480 gnd.n6479 585
R11614 gnd.n6479 gnd.n6478 585
R11615 gnd.n975 gnd.n974 585
R11616 gnd.n6306 gnd.n975 585
R11617 gnd.n6469 gnd.n6468 585
R11618 gnd.n6470 gnd.n6469 585
R11619 gnd.n986 gnd.n985 585
R11620 gnd.n6266 gnd.n985 585
R11621 gnd.n6464 gnd.n6463 585
R11622 gnd.n6463 gnd.n6462 585
R11623 gnd.n989 gnd.n988 585
R11624 gnd.n6288 gnd.n989 585
R11625 gnd.n6453 gnd.n6452 585
R11626 gnd.n6454 gnd.n6453 585
R11627 gnd.n1002 gnd.n1001 585
R11628 gnd.n6414 gnd.n1001 585
R11629 gnd.n6448 gnd.n6447 585
R11630 gnd.n6447 gnd.n6446 585
R11631 gnd.n1005 gnd.n1004 585
R11632 gnd.n1033 gnd.n1005 585
R11633 gnd.n6437 gnd.n6436 585
R11634 gnd.n6438 gnd.n6437 585
R11635 gnd.n1018 gnd.n1017 585
R11636 gnd.n1044 gnd.n1017 585
R11637 gnd.n6432 gnd.n6431 585
R11638 gnd.n6431 gnd.n6430 585
R11639 gnd.n1021 gnd.n1020 585
R11640 gnd.n6192 gnd.n1021 585
R11641 gnd.n6180 gnd.n1060 585
R11642 gnd.n1163 gnd.n1060 585
R11643 gnd.n6182 gnd.n6181 585
R11644 gnd.n6183 gnd.n6182 585
R11645 gnd.n1061 gnd.n1059 585
R11646 gnd.n6079 gnd.n1059 585
R11647 gnd.n6175 gnd.n6174 585
R11648 gnd.n6174 gnd.n6173 585
R11649 gnd.n1064 gnd.n1063 585
R11650 gnd.n1150 gnd.n1064 585
R11651 gnd.n6164 gnd.n6163 585
R11652 gnd.n6165 gnd.n6164 585
R11653 gnd.n1074 gnd.n1073 585
R11654 gnd.n6094 gnd.n1073 585
R11655 gnd.n6159 gnd.n6158 585
R11656 gnd.n6158 gnd.n6157 585
R11657 gnd.n1077 gnd.n1076 585
R11658 gnd.n1134 gnd.n1077 585
R11659 gnd.n6148 gnd.n6147 585
R11660 gnd.n6149 gnd.n6148 585
R11661 gnd.n1089 gnd.n1088 585
R11662 gnd.n6109 gnd.n1088 585
R11663 gnd.n6143 gnd.n6142 585
R11664 gnd.n6142 gnd.n6141 585
R11665 gnd.n1092 gnd.n1091 585
R11666 gnd.n1119 gnd.n1092 585
R11667 gnd.n6132 gnd.n6131 585
R11668 gnd.n6133 gnd.n6132 585
R11669 gnd.n1105 gnd.n1104 585
R11670 gnd.n1194 gnd.n1104 585
R11671 gnd.n6127 gnd.n6126 585
R11672 gnd.n6126 gnd.n6125 585
R11673 gnd.n1108 gnd.n1107 585
R11674 gnd.n6049 gnd.n1108 585
R11675 gnd.n6037 gnd.n1211 585
R11676 gnd.n5939 gnd.n1211 585
R11677 gnd.n6039 gnd.n6038 585
R11678 gnd.n6040 gnd.n6039 585
R11679 gnd.n1212 gnd.n1210 585
R11680 gnd.n5948 gnd.n1210 585
R11681 gnd.n6032 gnd.n6031 585
R11682 gnd.n6031 gnd.t7 585
R11683 gnd.n1215 gnd.n1214 585
R11684 gnd.n5883 gnd.n1215 585
R11685 gnd.n6022 gnd.n6021 585
R11686 gnd.n6023 gnd.n6022 585
R11687 gnd.n1227 gnd.n1226 585
R11688 gnd.n5888 gnd.n1226 585
R11689 gnd.n6017 gnd.n6016 585
R11690 gnd.n6016 gnd.n6015 585
R11691 gnd.n1230 gnd.n1229 585
R11692 gnd.n5901 gnd.n1230 585
R11693 gnd.n6006 gnd.n6005 585
R11694 gnd.n6007 gnd.n6006 585
R11695 gnd.n1243 gnd.n1242 585
R11696 gnd.n5967 gnd.n1242 585
R11697 gnd.n6001 gnd.n6000 585
R11698 gnd.n6000 gnd.n5999 585
R11699 gnd.n1246 gnd.n1245 585
R11700 gnd.n5853 gnd.n1246 585
R11701 gnd.n5990 gnd.n5989 585
R11702 gnd.n5991 gnd.n5990 585
R11703 gnd.n1258 gnd.n1257 585
R11704 gnd.n1282 gnd.n1257 585
R11705 gnd.n5985 gnd.n5984 585
R11706 gnd.n5984 gnd.n5983 585
R11707 gnd.n1261 gnd.n1260 585
R11708 gnd.n5844 gnd.n1261 585
R11709 gnd.n5832 gnd.n1299 585
R11710 gnd.n1411 gnd.n1299 585
R11711 gnd.n5834 gnd.n5833 585
R11712 gnd.n5835 gnd.n5834 585
R11713 gnd.n1300 gnd.n1298 585
R11714 gnd.n5677 gnd.n1298 585
R11715 gnd.n5827 gnd.n5826 585
R11716 gnd.n5826 gnd.n5825 585
R11717 gnd.n1303 gnd.n1302 585
R11718 gnd.n1312 gnd.n1303 585
R11719 gnd.n5816 gnd.n5815 585
R11720 gnd.n5817 gnd.n5816 585
R11721 gnd.n1314 gnd.n1313 585
R11722 gnd.n1313 gnd.n1310 585
R11723 gnd.n5811 gnd.n5810 585
R11724 gnd.n5810 gnd.n5809 585
R11725 gnd.n1317 gnd.n1316 585
R11726 gnd.n1318 gnd.n1317 585
R11727 gnd.n5356 gnd.n5352 585
R11728 gnd.n5352 gnd.n5351 585
R11729 gnd.n5359 gnd.n5357 585
R11730 gnd.n5359 gnd.n5358 585
R11731 gnd.n5360 gnd.n5350 585
R11732 gnd.n5360 gnd.n1356 585
R11733 gnd.n5362 gnd.n5361 585
R11734 gnd.n5361 gnd.n1354 585
R11735 gnd.n5363 gnd.n5345 585
R11736 gnd.n5345 gnd.n1649 585
R11737 gnd.n5365 gnd.n5364 585
R11738 gnd.n5365 gnd.n1658 585
R11739 gnd.n5366 gnd.n5344 585
R11740 gnd.n5366 gnd.n1655 585
R11741 gnd.n5368 gnd.n5367 585
R11742 gnd.n5367 gnd.n1668 585
R11743 gnd.n5369 gnd.n1835 585
R11744 gnd.n1835 gnd.n1665 585
R11745 gnd.n5371 gnd.n5370 585
R11746 gnd.n5372 gnd.n5371 585
R11747 gnd.n1836 gnd.n1834 585
R11748 gnd.n1834 gnd.n1674 585
R11749 gnd.n5338 gnd.n5337 585
R11750 gnd.n5337 gnd.n1684 585
R11751 gnd.n5336 gnd.n1838 585
R11752 gnd.n5336 gnd.n5335 585
R11753 gnd.n5307 gnd.n1839 585
R11754 gnd.n1839 gnd.n1693 585
R11755 gnd.n5309 gnd.n5308 585
R11756 gnd.n5309 gnd.n1690 585
R11757 gnd.n5311 gnd.n5310 585
R11758 gnd.n5310 gnd.n1702 585
R11759 gnd.n5312 gnd.n1845 585
R11760 gnd.n1845 gnd.n1699 585
R11761 gnd.n5314 gnd.n5313 585
R11762 gnd.n5315 gnd.n5314 585
R11763 gnd.n1846 gnd.n1844 585
R11764 gnd.n1844 gnd.n1708 585
R11765 gnd.n5299 gnd.n5298 585
R11766 gnd.n5298 gnd.n1718 585
R11767 gnd.n5297 gnd.n1848 585
R11768 gnd.n5297 gnd.n5296 585
R11769 gnd.n5267 gnd.n1849 585
R11770 gnd.n1849 gnd.n1727 585
R11771 gnd.n5269 gnd.n5268 585
R11772 gnd.n5269 gnd.n1724 585
R11773 gnd.n5271 gnd.n5270 585
R11774 gnd.n5270 gnd.n1736 585
R11775 gnd.n5272 gnd.n5256 585
R11776 gnd.n5256 gnd.n1733 585
R11777 gnd.n5274 gnd.n5273 585
R11778 gnd.n5275 gnd.n5274 585
R11779 gnd.n5257 gnd.n5255 585
R11780 gnd.n5255 gnd.n1742 585
R11781 gnd.n5259 gnd.n1805 585
R11782 gnd.n1805 gnd.n1752 585
R11783 gnd.n5431 gnd.n1804 585
R11784 gnd.n5431 gnd.n5430 585
R11785 gnd.n5433 gnd.n5432 585
R11786 gnd.n5432 gnd.n1761 585
R11787 gnd.n5434 gnd.n1799 585
R11788 gnd.n1799 gnd.n1758 585
R11789 gnd.n5436 gnd.n5435 585
R11790 gnd.n5437 gnd.n5436 585
R11791 gnd.n1800 gnd.n1798 585
R11792 gnd.n1798 gnd.n1795 585
R11793 gnd.n6760 gnd.n6759 585
R11794 gnd.n6759 gnd.n639 585
R11795 gnd.n6761 gnd.n638 585
R11796 gnd.n6808 gnd.n638 585
R11797 gnd.n6762 gnd.n6614 585
R11798 gnd.n6614 gnd.n6613 585
R11799 gnd.n871 gnd.n647 585
R11800 gnd.n6798 gnd.n647 585
R11801 gnd.n6767 gnd.n6766 585
R11802 gnd.n6768 gnd.n6767 585
R11803 gnd.n870 gnd.n654 585
R11804 gnd.n6789 gnd.n654 585
R11805 gnd.n6609 gnd.n6608 585
R11806 gnd.n6608 gnd.n669 585
R11807 gnd.n6607 gnd.n662 585
R11808 gnd.n6781 gnd.n662 585
R11809 gnd.n6606 gnd.n874 585
R11810 gnd.n6577 gnd.n874 585
R11811 gnd.n878 gnd.n873 585
R11812 gnd.n6568 gnd.n878 585
R11813 gnd.n6602 gnd.n6601 585
R11814 gnd.n6601 gnd.n6600 585
R11815 gnd.n877 gnd.n876 585
R11816 gnd.n906 gnd.n877 585
R11817 gnd.n915 gnd.n889 585
R11818 gnd.n6590 gnd.n889 585
R11819 gnd.n6550 gnd.n6549 585
R11820 gnd.n6551 gnd.n6550 585
R11821 gnd.n914 gnd.n913 585
R11822 gnd.n6523 gnd.n913 585
R11823 gnd.n6544 gnd.n6543 585
R11824 gnd.n6543 gnd.n6542 585
R11825 gnd.n918 gnd.n917 585
R11826 gnd.n6373 gnd.n918 585
R11827 gnd.n6383 gnd.n929 585
R11828 gnd.n6532 gnd.n929 585
R11829 gnd.n6384 gnd.n6382 585
R11830 gnd.n6382 gnd.n6381 585
R11831 gnd.n6219 gnd.n938 585
R11832 gnd.t4 gnd.n938 585
R11833 gnd.n6388 gnd.n6218 585
R11834 gnd.n6237 gnd.n6218 585
R11835 gnd.n6389 gnd.n946 585
R11836 gnd.n6510 gnd.n946 585
R11837 gnd.n6390 gnd.n6217 585
R11838 gnd.n6242 gnd.n6217 585
R11839 gnd.n6215 gnd.n954 585
R11840 gnd.n6502 gnd.n954 585
R11841 gnd.n6394 gnd.n6214 585
R11842 gnd.n6335 gnd.n6214 585
R11843 gnd.n6395 gnd.n962 585
R11844 gnd.n6494 gnd.n962 585
R11845 gnd.n6396 gnd.n6213 585
R11846 gnd.n6325 gnd.n6213 585
R11847 gnd.n6211 gnd.n969 585
R11848 gnd.n6486 gnd.n969 585
R11849 gnd.n6400 gnd.n6210 585
R11850 gnd.n6257 gnd.n6210 585
R11851 gnd.n6401 gnd.n977 585
R11852 gnd.n6478 gnd.n977 585
R11853 gnd.n6402 gnd.n6209 585
R11854 gnd.n6306 gnd.n6209 585
R11855 gnd.n6207 gnd.n983 585
R11856 gnd.n6470 gnd.n983 585
R11857 gnd.n6406 gnd.n6206 585
R11858 gnd.n6266 gnd.n6206 585
R11859 gnd.n6407 gnd.n991 585
R11860 gnd.n6462 gnd.n991 585
R11861 gnd.n6408 gnd.n6205 585
R11862 gnd.n6288 gnd.n6205 585
R11863 gnd.n1041 gnd.n999 585
R11864 gnd.n6454 gnd.n999 585
R11865 gnd.n6413 gnd.n6412 585
R11866 gnd.n6414 gnd.n6413 585
R11867 gnd.n1040 gnd.n1007 585
R11868 gnd.n6446 gnd.n1007 585
R11869 gnd.n6201 gnd.n6200 585
R11870 gnd.n6200 gnd.n1033 585
R11871 gnd.n6199 gnd.n1015 585
R11872 gnd.n6438 gnd.n1015 585
R11873 gnd.n6198 gnd.n1045 585
R11874 gnd.n1045 gnd.n1044 585
R11875 gnd.n1043 gnd.n1024 585
R11876 gnd.n6430 gnd.n1024 585
R11877 gnd.n6194 gnd.n6193 585
R11878 gnd.n6193 gnd.n6192 585
R11879 gnd.n1048 gnd.n1047 585
R11880 gnd.n1163 gnd.n1048 585
R11881 gnd.n1187 gnd.n1057 585
R11882 gnd.n6183 gnd.n1057 585
R11883 gnd.n6078 gnd.n6077 585
R11884 gnd.n6079 gnd.n6078 585
R11885 gnd.n1186 gnd.n1066 585
R11886 gnd.n6173 gnd.n1066 585
R11887 gnd.n6072 gnd.n6071 585
R11888 gnd.n6071 gnd.n1150 585
R11889 gnd.n6070 gnd.n1072 585
R11890 gnd.n6165 gnd.n1072 585
R11891 gnd.n6069 gnd.n1142 585
R11892 gnd.n6094 gnd.n1142 585
R11893 gnd.n1189 gnd.n1079 585
R11894 gnd.n6157 gnd.n1079 585
R11895 gnd.n6065 gnd.n6064 585
R11896 gnd.n6064 gnd.n1134 585
R11897 gnd.n6063 gnd.n1086 585
R11898 gnd.n6149 gnd.n1086 585
R11899 gnd.n6062 gnd.n1126 585
R11900 gnd.n6109 gnd.n1126 585
R11901 gnd.n1191 gnd.n1094 585
R11902 gnd.n6141 gnd.n1094 585
R11903 gnd.n6058 gnd.n6057 585
R11904 gnd.n6057 gnd.n1119 585
R11905 gnd.n6056 gnd.n1102 585
R11906 gnd.n6133 gnd.n1102 585
R11907 gnd.n6055 gnd.n1195 585
R11908 gnd.n1195 gnd.n1194 585
R11909 gnd.n1193 gnd.n1110 585
R11910 gnd.n6125 gnd.n1110 585
R11911 gnd.n6051 gnd.n6050 585
R11912 gnd.n6050 gnd.n6049 585
R11913 gnd.n1198 gnd.n1197 585
R11914 gnd.n5939 gnd.n1198 585
R11915 gnd.n5950 gnd.n1208 585
R11916 gnd.n6040 gnd.n1208 585
R11917 gnd.n5953 gnd.n5949 585
R11918 gnd.n5949 gnd.n5948 585
R11919 gnd.n5954 gnd.n1217 585
R11920 gnd.t7 gnd.n1217 585
R11921 gnd.n5955 gnd.n5863 585
R11922 gnd.n5883 gnd.n5863 585
R11923 gnd.n5861 gnd.n1224 585
R11924 gnd.n6023 gnd.n1224 585
R11925 gnd.n5959 gnd.n5860 585
R11926 gnd.n5888 gnd.n5860 585
R11927 gnd.n5960 gnd.n1232 585
R11928 gnd.n6015 gnd.n1232 585
R11929 gnd.n5961 gnd.n5859 585
R11930 gnd.n5901 gnd.n5859 585
R11931 gnd.n1279 gnd.n1240 585
R11932 gnd.n6007 gnd.n1240 585
R11933 gnd.n5966 gnd.n5965 585
R11934 gnd.n5967 gnd.n5966 585
R11935 gnd.n1278 gnd.n1247 585
R11936 gnd.n5999 gnd.n1247 585
R11937 gnd.n5855 gnd.n5854 585
R11938 gnd.n5854 gnd.n5853 585
R11939 gnd.n5851 gnd.n1255 585
R11940 gnd.n5991 gnd.n1255 585
R11941 gnd.n5850 gnd.n1283 585
R11942 gnd.n1283 gnd.n1282 585
R11943 gnd.n1281 gnd.n1263 585
R11944 gnd.n5983 gnd.n1263 585
R11945 gnd.n5846 gnd.n5845 585
R11946 gnd.n5845 gnd.n5844 585
R11947 gnd.n1286 gnd.n1285 585
R11948 gnd.n1411 gnd.n1286 585
R11949 gnd.n5680 gnd.n1296 585
R11950 gnd.n5835 gnd.n1296 585
R11951 gnd.n5679 gnd.n5678 585
R11952 gnd.n5678 gnd.n5677 585
R11953 gnd.n5684 gnd.n1304 585
R11954 gnd.n5825 gnd.n1304 585
R11955 gnd.n5685 gnd.n5676 585
R11956 gnd.n5676 gnd.n1312 585
R11957 gnd.n5686 gnd.n1311 585
R11958 gnd.n5817 gnd.n1311 585
R11959 gnd.n5582 gnd.n5581 585
R11960 gnd.n5669 gnd.n5583 585
R11961 gnd.n5668 gnd.n5584 585
R11962 gnd.n5593 gnd.n5585 585
R11963 gnd.n5661 gnd.n5594 585
R11964 gnd.n5660 gnd.n5595 585
R11965 gnd.n5597 gnd.n5596 585
R11966 gnd.n5653 gnd.n5606 585
R11967 gnd.n5652 gnd.n5607 585
R11968 gnd.n5616 gnd.n5608 585
R11969 gnd.n5645 gnd.n5617 585
R11970 gnd.n5644 gnd.n5618 585
R11971 gnd.n5620 gnd.n5619 585
R11972 gnd.n5637 gnd.n5632 585
R11973 gnd.n5636 gnd.n5633 585
R11974 gnd.n1344 gnd.n1343 585
R11975 gnd.n5778 gnd.n1345 585
R11976 gnd.n5781 gnd.n5780 585
R11977 gnd.n5779 gnd.n1340 585
R11978 gnd.n5787 gnd.n5786 585
R11979 gnd.n5789 gnd.n5788 585
R11980 gnd.n5792 gnd.n5791 585
R11981 gnd.n5790 gnd.n1338 585
R11982 gnd.n5797 gnd.n5796 585
R11983 gnd.n5799 gnd.n5798 585
R11984 gnd.n5802 gnd.n5801 585
R11985 gnd.n1333 gnd.n1332 585
R11986 gnd.n5807 gnd.n5806 585
R11987 gnd.n1334 gnd.n1309 585
R11988 gnd.n5809 gnd.n1309 585
R11989 gnd.n6811 gnd.n632 585
R11990 gnd.n639 gnd.n632 585
R11991 gnd.n6810 gnd.n6809 585
R11992 gnd.n6809 gnd.n6808 585
R11993 gnd.n637 gnd.n636 585
R11994 gnd.n6613 gnd.n637 585
R11995 gnd.n6797 gnd.n6796 585
R11996 gnd.n6798 gnd.n6797 585
R11997 gnd.n650 gnd.n649 585
R11998 gnd.n6768 gnd.n649 585
R11999 gnd.n6791 gnd.n6790 585
R12000 gnd.n6790 gnd.n6789 585
R12001 gnd.n653 gnd.n652 585
R12002 gnd.n669 gnd.n653 585
R12003 gnd.n6579 gnd.n663 585
R12004 gnd.n6781 gnd.n663 585
R12005 gnd.n6582 gnd.n6578 585
R12006 gnd.n6578 gnd.n6577 585
R12007 gnd.n6583 gnd.n897 585
R12008 gnd.n6568 gnd.n897 585
R12009 gnd.n6584 gnd.n881 585
R12010 gnd.n6600 gnd.n881 585
R12011 gnd.n894 gnd.n892 585
R12012 gnd.n906 gnd.n892 585
R12013 gnd.n6589 gnd.n6588 585
R12014 gnd.n6590 gnd.n6589 585
R12015 gnd.n893 gnd.n891 585
R12016 gnd.n6551 gnd.n891 585
R12017 gnd.n6525 gnd.n6524 585
R12018 gnd.n6524 gnd.n6523 585
R12019 gnd.n6526 gnd.n921 585
R12020 gnd.n6542 gnd.n921 585
R12021 gnd.n933 gnd.n931 585
R12022 gnd.n6373 gnd.n931 585
R12023 gnd.n6531 gnd.n6530 585
R12024 gnd.n6532 gnd.n6531 585
R12025 gnd.n932 gnd.n930 585
R12026 gnd.n6381 gnd.n930 585
R12027 gnd.n6519 gnd.n6518 585
R12028 gnd.n6518 gnd.t4 585
R12029 gnd.n936 gnd.n935 585
R12030 gnd.n6237 gnd.n936 585
R12031 gnd.n6509 gnd.n6508 585
R12032 gnd.n6510 gnd.n6509 585
R12033 gnd.n949 gnd.n948 585
R12034 gnd.n6242 gnd.n948 585
R12035 gnd.n6504 gnd.n6503 585
R12036 gnd.n6503 gnd.n6502 585
R12037 gnd.n952 gnd.n951 585
R12038 gnd.n6335 gnd.n952 585
R12039 gnd.n6493 gnd.n6492 585
R12040 gnd.n6494 gnd.n6493 585
R12041 gnd.n964 gnd.n963 585
R12042 gnd.n6325 gnd.n963 585
R12043 gnd.n6488 gnd.n6487 585
R12044 gnd.n6487 gnd.n6486 585
R12045 gnd.n967 gnd.n966 585
R12046 gnd.n6257 gnd.n967 585
R12047 gnd.n6477 gnd.n6476 585
R12048 gnd.n6478 gnd.n6477 585
R12049 gnd.n979 gnd.n978 585
R12050 gnd.n6306 gnd.n978 585
R12051 gnd.n6472 gnd.n6471 585
R12052 gnd.n6471 gnd.n6470 585
R12053 gnd.n982 gnd.n981 585
R12054 gnd.n6266 gnd.n982 585
R12055 gnd.n6461 gnd.n6460 585
R12056 gnd.n6462 gnd.n6461 585
R12057 gnd.n994 gnd.n993 585
R12058 gnd.n6288 gnd.n993 585
R12059 gnd.n6456 gnd.n6455 585
R12060 gnd.n6455 gnd.n6454 585
R12061 gnd.n997 gnd.n996 585
R12062 gnd.n6414 gnd.n997 585
R12063 gnd.n6445 gnd.n6444 585
R12064 gnd.n6446 gnd.n6445 585
R12065 gnd.n1010 gnd.n1009 585
R12066 gnd.n1033 gnd.n1009 585
R12067 gnd.n6440 gnd.n6439 585
R12068 gnd.n6439 gnd.n6438 585
R12069 gnd.n1013 gnd.n1012 585
R12070 gnd.n1044 gnd.n1013 585
R12071 gnd.n1052 gnd.n1026 585
R12072 gnd.n6430 gnd.n1026 585
R12073 gnd.n6191 gnd.n6190 585
R12074 gnd.n6192 gnd.n6191 585
R12075 gnd.n1051 gnd.n1050 585
R12076 gnd.n1163 gnd.n1050 585
R12077 gnd.n6185 gnd.n6184 585
R12078 gnd.n6184 gnd.n6183 585
R12079 gnd.n1055 gnd.n1054 585
R12080 gnd.n6079 gnd.n1055 585
R12081 gnd.n6172 gnd.n6171 585
R12082 gnd.n6173 gnd.n6172 585
R12083 gnd.n1068 gnd.n1067 585
R12084 gnd.n1150 gnd.n1067 585
R12085 gnd.n6167 gnd.n6166 585
R12086 gnd.n6166 gnd.n6165 585
R12087 gnd.n1071 gnd.n1070 585
R12088 gnd.n6094 gnd.n1071 585
R12089 gnd.n6156 gnd.n6155 585
R12090 gnd.n6157 gnd.n6156 585
R12091 gnd.n1082 gnd.n1081 585
R12092 gnd.n1134 gnd.n1081 585
R12093 gnd.n6151 gnd.n6150 585
R12094 gnd.n6150 gnd.n6149 585
R12095 gnd.n1085 gnd.n1084 585
R12096 gnd.n6109 gnd.n1085 585
R12097 gnd.n6140 gnd.n6139 585
R12098 gnd.n6141 gnd.n6140 585
R12099 gnd.n1097 gnd.n1096 585
R12100 gnd.n1119 gnd.n1096 585
R12101 gnd.n6135 gnd.n6134 585
R12102 gnd.n6134 gnd.n6133 585
R12103 gnd.n1100 gnd.n1099 585
R12104 gnd.n1194 gnd.n1100 585
R12105 gnd.n1203 gnd.n1112 585
R12106 gnd.n6125 gnd.n1112 585
R12107 gnd.n6048 gnd.n6047 585
R12108 gnd.n6049 gnd.n6048 585
R12109 gnd.n1202 gnd.n1201 585
R12110 gnd.n5939 gnd.n1201 585
R12111 gnd.n6042 gnd.n6041 585
R12112 gnd.n6041 gnd.n6040 585
R12113 gnd.n1206 gnd.n1205 585
R12114 gnd.n5948 gnd.n1206 585
R12115 gnd.n6030 gnd.n6029 585
R12116 gnd.t7 gnd.n6030 585
R12117 gnd.n1220 gnd.n1219 585
R12118 gnd.n5883 gnd.n1219 585
R12119 gnd.n6025 gnd.n6024 585
R12120 gnd.n6024 gnd.n6023 585
R12121 gnd.n1223 gnd.n1222 585
R12122 gnd.n5888 gnd.n1223 585
R12123 gnd.n6014 gnd.n6013 585
R12124 gnd.n6015 gnd.n6014 585
R12125 gnd.n1235 gnd.n1234 585
R12126 gnd.n5901 gnd.n1234 585
R12127 gnd.n6009 gnd.n6008 585
R12128 gnd.n6008 gnd.n6007 585
R12129 gnd.n1238 gnd.n1237 585
R12130 gnd.n5967 gnd.n1238 585
R12131 gnd.n5998 gnd.n5997 585
R12132 gnd.n5999 gnd.n5998 585
R12133 gnd.n1250 gnd.n1249 585
R12134 gnd.n5853 gnd.n1249 585
R12135 gnd.n5993 gnd.n5992 585
R12136 gnd.n5992 gnd.n5991 585
R12137 gnd.n1253 gnd.n1252 585
R12138 gnd.n1282 gnd.n1253 585
R12139 gnd.n1291 gnd.n1265 585
R12140 gnd.n5983 gnd.n1265 585
R12141 gnd.n5843 gnd.n5842 585
R12142 gnd.n5844 gnd.n5843 585
R12143 gnd.n1290 gnd.n1289 585
R12144 gnd.n1411 gnd.n1289 585
R12145 gnd.n5837 gnd.n5836 585
R12146 gnd.n5836 gnd.n5835 585
R12147 gnd.n1294 gnd.n1293 585
R12148 gnd.n5677 gnd.n1294 585
R12149 gnd.n5824 gnd.n5823 585
R12150 gnd.n5825 gnd.n5824 585
R12151 gnd.n1307 gnd.n1306 585
R12152 gnd.n1312 gnd.n1306 585
R12153 gnd.n5819 gnd.n5818 585
R12154 gnd.n5818 gnd.n5817 585
R12155 gnd.n6815 gnd.n6814 585
R12156 gnd.n6817 gnd.n6815 585
R12157 gnd.n633 gnd.n631 585
R12158 gnd.n6694 gnd.n6693 585
R12159 gnd.n6695 gnd.n6692 585
R12160 gnd.n6687 gnd.n6686 585
R12161 gnd.n6699 gnd.n6685 585
R12162 gnd.n6700 gnd.n6684 585
R12163 gnd.n6701 gnd.n6683 585
R12164 gnd.n6681 gnd.n6680 585
R12165 gnd.n6705 gnd.n6679 585
R12166 gnd.n6706 gnd.n6678 585
R12167 gnd.n6707 gnd.n6677 585
R12168 gnd.n6674 gnd.n6673 585
R12169 gnd.n6717 gnd.n6672 585
R12170 gnd.n6718 gnd.n6671 585
R12171 gnd.n6670 gnd.n6662 585
R12172 gnd.n6725 gnd.n6661 585
R12173 gnd.n6726 gnd.n6660 585
R12174 gnd.n6654 gnd.n6653 585
R12175 gnd.n6733 gnd.n6652 585
R12176 gnd.n6734 gnd.n6651 585
R12177 gnd.n6650 gnd.n6642 585
R12178 gnd.n6741 gnd.n6641 585
R12179 gnd.n6742 gnd.n6640 585
R12180 gnd.n6634 gnd.n6633 585
R12181 gnd.n6749 gnd.n6632 585
R12182 gnd.n6750 gnd.n6631 585
R12183 gnd.n6630 gnd.n6616 585
R12184 gnd.n6758 gnd.n6757 585
R12185 gnd.n730 gnd.n675 506.916
R12186 gnd.n865 gnd.n676 506.916
R12187 gnd.n1539 gnd.n1537 506.916
R12188 gnd.n1517 gnd.n1516 506.916
R12189 gnd.n3142 gnd.n3141 414.56
R12190 gnd.n1394 gnd.t110 389.64
R12191 gnd.n804 gnd.t47 389.64
R12192 gnd.n1450 gnd.t57 389.64
R12193 gnd.n785 gnd.t101 389.64
R12194 gnd.n1336 gnd.t94 371.625
R12195 gnd.n118 gnd.t28 371.625
R12196 gnd.n6712 gnd.t68 371.625
R12197 gnd.n1348 gnd.t81 371.625
R12198 gnd.n537 gnd.t61 371.625
R12199 gnd.n559 gnd.t32 371.625
R12200 gnd.n197 gnd.t107 371.625
R12201 gnd.n7536 gnd.t116 371.625
R12202 gnd.n4900 gnd.t54 371.625
R12203 gnd.n4932 gnd.t24 371.625
R12204 gnd.n4761 gnd.t91 371.625
R12205 gnd.n1641 gnd.t43 371.625
R12206 gnd.n1388 gnd.t78 371.625
R12207 gnd.n6689 gnd.t74 371.625
R12208 gnd.n3838 gnd.t20 323.425
R12209 gnd.n2027 gnd.t64 323.425
R12210 gnd.n4625 gnd.n4599 289.615
R12211 gnd.n4593 gnd.n4567 289.615
R12212 gnd.n4561 gnd.n4535 289.615
R12213 gnd.n4530 gnd.n4504 289.615
R12214 gnd.n4498 gnd.n4472 289.615
R12215 gnd.n4466 gnd.n4440 289.615
R12216 gnd.n4434 gnd.n4408 289.615
R12217 gnd.n4403 gnd.n4377 289.615
R12218 gnd.n3912 gnd.t87 279.217
R12219 gnd.n2053 gnd.t36 279.217
R12220 gnd.n1420 gnd.t100 260.649
R12221 gnd.n720 gnd.t106 260.649
R12222 gnd.n1435 gnd.n1305 256.663
R12223 gnd.n1437 gnd.n1305 256.663
R12224 gnd.n1506 gnd.n1305 256.663
R12225 gnd.n1500 gnd.n1305 256.663
R12226 gnd.n1498 gnd.n1305 256.663
R12227 gnd.n1492 gnd.n1305 256.663
R12228 gnd.n1490 gnd.n1305 256.663
R12229 gnd.n1484 gnd.n1305 256.663
R12230 gnd.n1482 gnd.n1305 256.663
R12231 gnd.n1476 gnd.n1305 256.663
R12232 gnd.n1474 gnd.n1305 256.663
R12233 gnd.n1468 gnd.n1305 256.663
R12234 gnd.n1466 gnd.n1305 256.663
R12235 gnd.n1460 gnd.n1305 256.663
R12236 gnd.n1453 gnd.n1305 256.663
R12237 gnd.n1454 gnd.n1305 256.663
R12238 gnd.n1605 gnd.n1392 256.663
R12239 gnd.n1603 gnd.n1305 256.663
R12240 gnd.n1601 gnd.n1305 256.663
R12241 gnd.n1594 gnd.n1305 256.663
R12242 gnd.n1592 gnd.n1305 256.663
R12243 gnd.n1586 gnd.n1305 256.663
R12244 gnd.n1584 gnd.n1305 256.663
R12245 gnd.n1578 gnd.n1305 256.663
R12246 gnd.n1576 gnd.n1305 256.663
R12247 gnd.n1570 gnd.n1305 256.663
R12248 gnd.n1568 gnd.n1305 256.663
R12249 gnd.n1562 gnd.n1305 256.663
R12250 gnd.n1560 gnd.n1305 256.663
R12251 gnd.n1554 gnd.n1305 256.663
R12252 gnd.n1552 gnd.n1305 256.663
R12253 gnd.n1546 gnd.n1305 256.663
R12254 gnd.n1544 gnd.n1305 256.663
R12255 gnd.n1538 gnd.n1305 256.663
R12256 gnd.n864 gnd.n648 256.663
R12257 gnd.n678 gnd.n648 256.663
R12258 gnd.n857 gnd.n648 256.663
R12259 gnd.n851 gnd.n648 256.663
R12260 gnd.n849 gnd.n648 256.663
R12261 gnd.n843 gnd.n648 256.663
R12262 gnd.n841 gnd.n648 256.663
R12263 gnd.n835 gnd.n648 256.663
R12264 gnd.n833 gnd.n648 256.663
R12265 gnd.n827 gnd.n648 256.663
R12266 gnd.n825 gnd.n648 256.663
R12267 gnd.n819 gnd.n648 256.663
R12268 gnd.n817 gnd.n648 256.663
R12269 gnd.n811 gnd.n648 256.663
R12270 gnd.n809 gnd.n648 256.663
R12271 gnd.n800 gnd.n648 256.663
R12272 gnd.n798 gnd.n534 256.663
R12273 gnd.n797 gnd.n648 256.663
R12274 gnd.n693 gnd.n648 256.663
R12275 gnd.n790 gnd.n648 256.663
R12276 gnd.n781 gnd.n648 256.663
R12277 gnd.n779 gnd.n648 256.663
R12278 gnd.n773 gnd.n648 256.663
R12279 gnd.n771 gnd.n648 256.663
R12280 gnd.n765 gnd.n648 256.663
R12281 gnd.n763 gnd.n648 256.663
R12282 gnd.n757 gnd.n648 256.663
R12283 gnd.n755 gnd.n648 256.663
R12284 gnd.n749 gnd.n648 256.663
R12285 gnd.n747 gnd.n648 256.663
R12286 gnd.n741 gnd.n648 256.663
R12287 gnd.n739 gnd.n648 256.663
R12288 gnd.n733 gnd.n648 256.663
R12289 gnd.n731 gnd.n648 256.663
R12290 gnd.n4781 gnd.n4756 242.672
R12291 gnd.n4783 gnd.n4756 242.672
R12292 gnd.n4791 gnd.n4756 242.672
R12293 gnd.n4793 gnd.n4756 242.672
R12294 gnd.n4801 gnd.n4756 242.672
R12295 gnd.n4803 gnd.n4756 242.672
R12296 gnd.n4811 gnd.n4756 242.672
R12297 gnd.n4813 gnd.n4756 242.672
R12298 gnd.n4821 gnd.n4756 242.672
R12299 gnd.n1364 gnd.n1351 242.672
R12300 gnd.n5628 gnd.n1364 242.672
R12301 gnd.n5625 gnd.n1364 242.672
R12302 gnd.n5622 gnd.n1364 242.672
R12303 gnd.n5611 gnd.n1364 242.672
R12304 gnd.n5602 gnd.n1364 242.672
R12305 gnd.n5599 gnd.n1364 242.672
R12306 gnd.n5588 gnd.n1364 242.672
R12307 gnd.n5577 gnd.n1364 242.672
R12308 gnd.n7046 gnd.n508 242.672
R12309 gnd.n7046 gnd.n509 242.672
R12310 gnd.n7046 gnd.n510 242.672
R12311 gnd.n7046 gnd.n511 242.672
R12312 gnd.n7046 gnd.n512 242.672
R12313 gnd.n7046 gnd.n513 242.672
R12314 gnd.n7046 gnd.n514 242.672
R12315 gnd.n7046 gnd.n515 242.672
R12316 gnd.n7046 gnd.n516 242.672
R12317 gnd.n124 gnd.n121 242.672
R12318 gnd.n7447 gnd.n124 242.672
R12319 gnd.n7443 gnd.n124 242.672
R12320 gnd.n7440 gnd.n124 242.672
R12321 gnd.n7435 gnd.n124 242.672
R12322 gnd.n7432 gnd.n124 242.672
R12323 gnd.n7427 gnd.n124 242.672
R12324 gnd.n7424 gnd.n124 242.672
R12325 gnd.n7419 gnd.n124 242.672
R12326 gnd.n3966 gnd.n3965 242.672
R12327 gnd.n3966 gnd.n3876 242.672
R12328 gnd.n3966 gnd.n3877 242.672
R12329 gnd.n3966 gnd.n3878 242.672
R12330 gnd.n3966 gnd.n3879 242.672
R12331 gnd.n3966 gnd.n3880 242.672
R12332 gnd.n3966 gnd.n3881 242.672
R12333 gnd.n3966 gnd.n3882 242.672
R12334 gnd.n3966 gnd.n3883 242.672
R12335 gnd.n3966 gnd.n3884 242.672
R12336 gnd.n3966 gnd.n3885 242.672
R12337 gnd.n3966 gnd.n3886 242.672
R12338 gnd.n3967 gnd.n3966 242.672
R12339 gnd.n4755 gnd.n2002 242.672
R12340 gnd.n4755 gnd.n2001 242.672
R12341 gnd.n4755 gnd.n2000 242.672
R12342 gnd.n4755 gnd.n1999 242.672
R12343 gnd.n4755 gnd.n1998 242.672
R12344 gnd.n4755 gnd.n1997 242.672
R12345 gnd.n4755 gnd.n1996 242.672
R12346 gnd.n4755 gnd.n1995 242.672
R12347 gnd.n4755 gnd.n1994 242.672
R12348 gnd.n4755 gnd.n1993 242.672
R12349 gnd.n4755 gnd.n1992 242.672
R12350 gnd.n4755 gnd.n1991 242.672
R12351 gnd.n4755 gnd.n1990 242.672
R12352 gnd.n4050 gnd.n4049 242.672
R12353 gnd.n4049 gnd.n3788 242.672
R12354 gnd.n4049 gnd.n3789 242.672
R12355 gnd.n4049 gnd.n3790 242.672
R12356 gnd.n4049 gnd.n3791 242.672
R12357 gnd.n4049 gnd.n3792 242.672
R12358 gnd.n4049 gnd.n3793 242.672
R12359 gnd.n4049 gnd.n3794 242.672
R12360 gnd.n4755 gnd.n2003 242.672
R12361 gnd.n4755 gnd.n2004 242.672
R12362 gnd.n4755 gnd.n2005 242.672
R12363 gnd.n4755 gnd.n2006 242.672
R12364 gnd.n4755 gnd.n2007 242.672
R12365 gnd.n4755 gnd.n2008 242.672
R12366 gnd.n4755 gnd.n2009 242.672
R12367 gnd.n4755 gnd.n2010 242.672
R12368 gnd.n5062 gnd.n4756 242.672
R12369 gnd.n4876 gnd.n4756 242.672
R12370 gnd.n5055 gnd.n4756 242.672
R12371 gnd.n5049 gnd.n4756 242.672
R12372 gnd.n5047 gnd.n4756 242.672
R12373 gnd.n5041 gnd.n4756 242.672
R12374 gnd.n5039 gnd.n4756 242.672
R12375 gnd.n5033 gnd.n4756 242.672
R12376 gnd.n5031 gnd.n4756 242.672
R12377 gnd.n5025 gnd.n4756 242.672
R12378 gnd.n5023 gnd.n4756 242.672
R12379 gnd.n5017 gnd.n4756 242.672
R12380 gnd.n5015 gnd.n4756 242.672
R12381 gnd.n5009 gnd.n4756 242.672
R12382 gnd.n5007 gnd.n4756 242.672
R12383 gnd.n5001 gnd.n4756 242.672
R12384 gnd.n4999 gnd.n4756 242.672
R12385 gnd.n4930 gnd.n4756 242.672
R12386 gnd.n4989 gnd.n4756 242.672
R12387 gnd.n5702 gnd.n1364 242.672
R12388 gnd.n1644 gnd.n1364 242.672
R12389 gnd.n5709 gnd.n1364 242.672
R12390 gnd.n1635 gnd.n1364 242.672
R12391 gnd.n5716 gnd.n1364 242.672
R12392 gnd.n1628 gnd.n1364 242.672
R12393 gnd.n5723 gnd.n1364 242.672
R12394 gnd.n1621 gnd.n1364 242.672
R12395 gnd.n5730 gnd.n1364 242.672
R12396 gnd.n1614 gnd.n1364 242.672
R12397 gnd.n5737 gnd.n1364 242.672
R12398 gnd.n5738 gnd.n1606 242.672
R12399 gnd.n5739 gnd.n1364 242.672
R12400 gnd.n1387 gnd.n1364 242.672
R12401 gnd.n5746 gnd.n1364 242.672
R12402 gnd.n1380 gnd.n1364 242.672
R12403 gnd.n5753 gnd.n1364 242.672
R12404 gnd.n1373 gnd.n1364 242.672
R12405 gnd.n5760 gnd.n1364 242.672
R12406 gnd.n5763 gnd.n1364 242.672
R12407 gnd.n7047 gnd.n7046 242.672
R12408 gnd.n7046 gnd.n490 242.672
R12409 gnd.n7046 gnd.n491 242.672
R12410 gnd.n7046 gnd.n492 242.672
R12411 gnd.n7046 gnd.n493 242.672
R12412 gnd.n7046 gnd.n494 242.672
R12413 gnd.n7046 gnd.n495 242.672
R12414 gnd.n7046 gnd.n496 242.672
R12415 gnd.n7018 gnd.n535 242.672
R12416 gnd.n7046 gnd.n497 242.672
R12417 gnd.n7046 gnd.n498 242.672
R12418 gnd.n7046 gnd.n499 242.672
R12419 gnd.n7046 gnd.n500 242.672
R12420 gnd.n7046 gnd.n501 242.672
R12421 gnd.n7046 gnd.n502 242.672
R12422 gnd.n7046 gnd.n503 242.672
R12423 gnd.n7046 gnd.n504 242.672
R12424 gnd.n7046 gnd.n505 242.672
R12425 gnd.n7046 gnd.n506 242.672
R12426 gnd.n7046 gnd.n507 242.672
R12427 gnd.n194 gnd.n124 242.672
R12428 gnd.n7504 gnd.n124 242.672
R12429 gnd.n190 gnd.n124 242.672
R12430 gnd.n7511 gnd.n124 242.672
R12431 gnd.n183 gnd.n124 242.672
R12432 gnd.n7518 gnd.n124 242.672
R12433 gnd.n176 gnd.n124 242.672
R12434 gnd.n7525 gnd.n124 242.672
R12435 gnd.n169 gnd.n124 242.672
R12436 gnd.n7532 gnd.n124 242.672
R12437 gnd.n162 gnd.n124 242.672
R12438 gnd.n7542 gnd.n124 242.672
R12439 gnd.n155 gnd.n124 242.672
R12440 gnd.n7549 gnd.n124 242.672
R12441 gnd.n148 gnd.n124 242.672
R12442 gnd.n7556 gnd.n124 242.672
R12443 gnd.n141 gnd.n124 242.672
R12444 gnd.n7563 gnd.n124 242.672
R12445 gnd.n134 gnd.n124 242.672
R12446 gnd.n5809 gnd.n1319 242.672
R12447 gnd.n5809 gnd.n1320 242.672
R12448 gnd.n5809 gnd.n1321 242.672
R12449 gnd.n5809 gnd.n1322 242.672
R12450 gnd.n5809 gnd.n1323 242.672
R12451 gnd.n5809 gnd.n1324 242.672
R12452 gnd.n5809 gnd.n1325 242.672
R12453 gnd.n5809 gnd.n1326 242.672
R12454 gnd.n5809 gnd.n1327 242.672
R12455 gnd.n5809 gnd.n1328 242.672
R12456 gnd.n5809 gnd.n1329 242.672
R12457 gnd.n5809 gnd.n1330 242.672
R12458 gnd.n5809 gnd.n1331 242.672
R12459 gnd.n5809 gnd.n5808 242.672
R12460 gnd.n6817 gnd.n630 242.672
R12461 gnd.n6817 gnd.n629 242.672
R12462 gnd.n6817 gnd.n628 242.672
R12463 gnd.n6817 gnd.n627 242.672
R12464 gnd.n6817 gnd.n626 242.672
R12465 gnd.n6817 gnd.n625 242.672
R12466 gnd.n6817 gnd.n624 242.672
R12467 gnd.n6817 gnd.n623 242.672
R12468 gnd.n6817 gnd.n622 242.672
R12469 gnd.n6817 gnd.n621 242.672
R12470 gnd.n6817 gnd.n620 242.672
R12471 gnd.n6817 gnd.n619 242.672
R12472 gnd.n6817 gnd.n618 242.672
R12473 gnd.n6817 gnd.n617 242.672
R12474 gnd.n131 gnd.n127 240.244
R12475 gnd.n7565 gnd.n7564 240.244
R12476 gnd.n7562 gnd.n135 240.244
R12477 gnd.n7558 gnd.n7557 240.244
R12478 gnd.n7555 gnd.n142 240.244
R12479 gnd.n7551 gnd.n7550 240.244
R12480 gnd.n7548 gnd.n149 240.244
R12481 gnd.n7544 gnd.n7543 240.244
R12482 gnd.n7541 gnd.n156 240.244
R12483 gnd.n7534 gnd.n7533 240.244
R12484 gnd.n7531 gnd.n163 240.244
R12485 gnd.n7527 gnd.n7526 240.244
R12486 gnd.n7524 gnd.n170 240.244
R12487 gnd.n7520 gnd.n7519 240.244
R12488 gnd.n7517 gnd.n177 240.244
R12489 gnd.n7513 gnd.n7512 240.244
R12490 gnd.n7510 gnd.n184 240.244
R12491 gnd.n7506 gnd.n7505 240.244
R12492 gnd.n7503 gnd.n191 240.244
R12493 gnd.n6975 gnd.n481 240.244
R12494 gnd.n6847 gnd.n481 240.244
R12495 gnd.n6847 gnd.n472 240.244
R12496 gnd.n6851 gnd.n472 240.244
R12497 gnd.n6851 gnd.n463 240.244
R12498 gnd.n6864 gnd.n463 240.244
R12499 gnd.n6864 gnd.n454 240.244
R12500 gnd.n6860 gnd.n454 240.244
R12501 gnd.n6860 gnd.n447 240.244
R12502 gnd.n6887 gnd.n447 240.244
R12503 gnd.n6887 gnd.n438 240.244
R12504 gnd.n6891 gnd.n438 240.244
R12505 gnd.n6891 gnd.n429 240.244
R12506 gnd.n6903 gnd.n429 240.244
R12507 gnd.n6903 gnd.n420 240.244
R12508 gnd.n6899 gnd.n420 240.244
R12509 gnd.n6899 gnd.n413 240.244
R12510 gnd.n6918 gnd.n413 240.244
R12511 gnd.n6918 gnd.n402 240.244
R12512 gnd.n6937 gnd.n402 240.244
R12513 gnd.n6937 gnd.n394 240.244
R12514 gnd.n394 gnd.n387 240.244
R12515 gnd.n387 gnd.n370 240.244
R12516 gnd.n6931 gnd.n370 240.244
R12517 gnd.n6931 gnd.n358 240.244
R12518 gnd.n7191 gnd.n358 240.244
R12519 gnd.n7192 gnd.n7191 240.244
R12520 gnd.n7192 gnd.n350 240.244
R12521 gnd.n350 gnd.n309 240.244
R12522 gnd.n7201 gnd.n309 240.244
R12523 gnd.n7201 gnd.n339 240.244
R12524 gnd.n339 gnd.n335 240.244
R12525 gnd.n7229 gnd.n335 240.244
R12526 gnd.n7229 gnd.n331 240.244
R12527 gnd.n7300 gnd.n331 240.244
R12528 gnd.n7300 gnd.n324 240.244
R12529 gnd.n7296 gnd.n324 240.244
R12530 gnd.n7296 gnd.n296 240.244
R12531 gnd.n7293 gnd.n296 240.244
R12532 gnd.n7293 gnd.n287 240.244
R12533 gnd.n7290 gnd.n287 240.244
R12534 gnd.n7290 gnd.n279 240.244
R12535 gnd.n7287 gnd.n279 240.244
R12536 gnd.n7287 gnd.n272 240.244
R12537 gnd.n7284 gnd.n272 240.244
R12538 gnd.n7284 gnd.n266 240.244
R12539 gnd.n7281 gnd.n266 240.244
R12540 gnd.n7281 gnd.n257 240.244
R12541 gnd.n7278 gnd.n257 240.244
R12542 gnd.n7278 gnd.n249 240.244
R12543 gnd.n7275 gnd.n249 240.244
R12544 gnd.n7275 gnd.n242 240.244
R12545 gnd.n7272 gnd.n242 240.244
R12546 gnd.n7272 gnd.n235 240.244
R12547 gnd.n7269 gnd.n235 240.244
R12548 gnd.n7269 gnd.n226 240.244
R12549 gnd.n7266 gnd.n226 240.244
R12550 gnd.n7266 gnd.n219 240.244
R12551 gnd.n7263 gnd.n219 240.244
R12552 gnd.n7263 gnd.n210 240.244
R12553 gnd.n210 gnd.n201 240.244
R12554 gnd.n7494 gnd.n201 240.244
R12555 gnd.n7495 gnd.n7494 240.244
R12556 gnd.n7495 gnd.n123 240.244
R12557 gnd.n7045 gnd.n488 240.244
R12558 gnd.n7045 gnd.n519 240.244
R12559 gnd.n7041 gnd.n7040 240.244
R12560 gnd.n7037 gnd.n7036 240.244
R12561 gnd.n7033 gnd.n7032 240.244
R12562 gnd.n7029 gnd.n7028 240.244
R12563 gnd.n7025 gnd.n7024 240.244
R12564 gnd.n7021 gnd.n7020 240.244
R12565 gnd.n7016 gnd.n7015 240.244
R12566 gnd.n7012 gnd.n7011 240.244
R12567 gnd.n7008 gnd.n7007 240.244
R12568 gnd.n7004 gnd.n7003 240.244
R12569 gnd.n7000 gnd.n6999 240.244
R12570 gnd.n6996 gnd.n6995 240.244
R12571 gnd.n6992 gnd.n6991 240.244
R12572 gnd.n6988 gnd.n6987 240.244
R12573 gnd.n6984 gnd.n6983 240.244
R12574 gnd.n558 gnd.n557 240.244
R12575 gnd.n7054 gnd.n484 240.244
R12576 gnd.n7054 gnd.n470 240.244
R12577 gnd.n7064 gnd.n470 240.244
R12578 gnd.n7064 gnd.n466 240.244
R12579 gnd.n7070 gnd.n466 240.244
R12580 gnd.n7070 gnd.n453 240.244
R12581 gnd.n7080 gnd.n453 240.244
R12582 gnd.n7080 gnd.n449 240.244
R12583 gnd.n7086 gnd.n449 240.244
R12584 gnd.n7086 gnd.n436 240.244
R12585 gnd.n7096 gnd.n436 240.244
R12586 gnd.n7096 gnd.n432 240.244
R12587 gnd.n7102 gnd.n432 240.244
R12588 gnd.n7102 gnd.n419 240.244
R12589 gnd.n7112 gnd.n419 240.244
R12590 gnd.n7112 gnd.n415 240.244
R12591 gnd.n7118 gnd.n415 240.244
R12592 gnd.n7118 gnd.n400 240.244
R12593 gnd.n7131 gnd.n400 240.244
R12594 gnd.n7131 gnd.n396 240.244
R12595 gnd.n7137 gnd.n396 240.244
R12596 gnd.n7137 gnd.n368 240.244
R12597 gnd.n7182 gnd.n368 240.244
R12598 gnd.n7182 gnd.n369 240.244
R12599 gnd.n369 gnd.n363 240.244
R12600 gnd.n7189 gnd.n363 240.244
R12601 gnd.n7189 gnd.n364 240.244
R12602 gnd.n364 gnd.n306 240.244
R12603 gnd.n7321 gnd.n306 240.244
R12604 gnd.n7321 gnd.n307 240.244
R12605 gnd.n7223 gnd.n307 240.244
R12606 gnd.n7224 gnd.n7223 240.244
R12607 gnd.n7227 gnd.n7224 240.244
R12608 gnd.n7227 gnd.n326 240.244
R12609 gnd.n7302 gnd.n326 240.244
R12610 gnd.n7304 gnd.n7302 240.244
R12611 gnd.n7304 gnd.n297 240.244
R12612 gnd.n7328 gnd.n297 240.244
R12613 gnd.n7328 gnd.n285 240.244
R12614 gnd.n7338 gnd.n285 240.244
R12615 gnd.n7338 gnd.n281 240.244
R12616 gnd.n7344 gnd.n281 240.244
R12617 gnd.n7344 gnd.n271 240.244
R12618 gnd.n7354 gnd.n271 240.244
R12619 gnd.n7354 gnd.n267 240.244
R12620 gnd.n7360 gnd.n267 240.244
R12621 gnd.n7360 gnd.n255 240.244
R12622 gnd.n7370 gnd.n255 240.244
R12623 gnd.n7370 gnd.n251 240.244
R12624 gnd.n7376 gnd.n251 240.244
R12625 gnd.n7376 gnd.n241 240.244
R12626 gnd.n7386 gnd.n241 240.244
R12627 gnd.n7386 gnd.n237 240.244
R12628 gnd.n7392 gnd.n237 240.244
R12629 gnd.n7392 gnd.n224 240.244
R12630 gnd.n7402 gnd.n224 240.244
R12631 gnd.n7402 gnd.n220 240.244
R12632 gnd.n7408 gnd.n220 240.244
R12633 gnd.n7408 gnd.n208 240.244
R12634 gnd.n7486 gnd.n208 240.244
R12635 gnd.n7486 gnd.n204 240.244
R12636 gnd.n7492 gnd.n204 240.244
R12637 gnd.n7492 gnd.n126 240.244
R12638 gnd.n7572 gnd.n126 240.244
R12639 gnd.n5764 gnd.n1359 240.244
R12640 gnd.n5762 gnd.n5761 240.244
R12641 gnd.n5759 gnd.n1366 240.244
R12642 gnd.n5755 gnd.n5754 240.244
R12643 gnd.n5752 gnd.n1374 240.244
R12644 gnd.n5748 gnd.n5747 240.244
R12645 gnd.n5745 gnd.n1381 240.244
R12646 gnd.n5741 gnd.n5740 240.244
R12647 gnd.n5736 gnd.n1607 240.244
R12648 gnd.n5732 gnd.n5731 240.244
R12649 gnd.n5729 gnd.n1615 240.244
R12650 gnd.n5725 gnd.n5724 240.244
R12651 gnd.n5722 gnd.n1622 240.244
R12652 gnd.n5718 gnd.n5717 240.244
R12653 gnd.n5715 gnd.n1629 240.244
R12654 gnd.n5711 gnd.n5710 240.244
R12655 gnd.n5708 gnd.n1636 240.244
R12656 gnd.n5704 gnd.n5703 240.244
R12657 gnd.n4936 gnd.n4757 240.244
R12658 gnd.n4936 gnd.n1982 240.244
R12659 gnd.n4982 gnd.n1982 240.244
R12660 gnd.n4982 gnd.n1975 240.244
R12661 gnd.n4979 gnd.n1975 240.244
R12662 gnd.n4979 gnd.n1967 240.244
R12663 gnd.n4976 gnd.n1967 240.244
R12664 gnd.n4976 gnd.n1958 240.244
R12665 gnd.n4973 gnd.n1958 240.244
R12666 gnd.n4973 gnd.n1950 240.244
R12667 gnd.n4970 gnd.n1950 240.244
R12668 gnd.n4970 gnd.n1943 240.244
R12669 gnd.n4967 gnd.n1943 240.244
R12670 gnd.n4967 gnd.n1935 240.244
R12671 gnd.n4964 gnd.n1935 240.244
R12672 gnd.n4964 gnd.n1926 240.244
R12673 gnd.n4961 gnd.n1926 240.244
R12674 gnd.n4961 gnd.n1917 240.244
R12675 gnd.n4958 gnd.n1917 240.244
R12676 gnd.n4958 gnd.n1909 240.244
R12677 gnd.n1909 gnd.n1901 240.244
R12678 gnd.n5174 gnd.n1901 240.244
R12679 gnd.n5174 gnd.n1882 240.244
R12680 gnd.n1897 gnd.n1882 240.244
R12681 gnd.n5183 gnd.n1897 240.244
R12682 gnd.n5183 gnd.n1873 240.244
R12683 gnd.n1873 gnd.n1866 240.244
R12684 gnd.n5218 gnd.n1866 240.244
R12685 gnd.n5218 gnd.n1773 240.244
R12686 gnd.n5223 gnd.n1773 240.244
R12687 gnd.n5223 gnd.n1784 240.244
R12688 gnd.n5226 gnd.n1784 240.244
R12689 gnd.n5226 gnd.n1789 240.244
R12690 gnd.n5232 gnd.n1789 240.244
R12691 gnd.n5232 gnd.n1796 240.244
R12692 gnd.n5242 gnd.n1796 240.244
R12693 gnd.n5242 gnd.n1759 240.244
R12694 gnd.n1806 gnd.n1759 240.244
R12695 gnd.n1806 gnd.n1750 240.244
R12696 gnd.n5250 gnd.n1750 240.244
R12697 gnd.n5250 gnd.n1743 240.244
R12698 gnd.n5277 gnd.n1743 240.244
R12699 gnd.n5277 gnd.n1734 240.244
R12700 gnd.n5281 gnd.n1734 240.244
R12701 gnd.n5281 gnd.n1725 240.244
R12702 gnd.n5294 gnd.n1725 240.244
R12703 gnd.n5294 gnd.n1716 240.244
R12704 gnd.n5290 gnd.n1716 240.244
R12705 gnd.n5290 gnd.n1709 240.244
R12706 gnd.n5317 gnd.n1709 240.244
R12707 gnd.n5317 gnd.n1700 240.244
R12708 gnd.n5321 gnd.n1700 240.244
R12709 gnd.n5321 gnd.n1691 240.244
R12710 gnd.n5333 gnd.n1691 240.244
R12711 gnd.n5333 gnd.n1682 240.244
R12712 gnd.n5329 gnd.n1682 240.244
R12713 gnd.n5329 gnd.n1675 240.244
R12714 gnd.n5374 gnd.n1675 240.244
R12715 gnd.n5374 gnd.n1666 240.244
R12716 gnd.n5383 gnd.n1666 240.244
R12717 gnd.n5383 gnd.n1656 240.244
R12718 gnd.n1656 gnd.n1648 240.244
R12719 gnd.n5695 gnd.n1648 240.244
R12720 gnd.n5695 gnd.n1355 240.244
R12721 gnd.n5063 gnd.n5061 240.244
R12722 gnd.n5061 gnd.n5060 240.244
R12723 gnd.n5057 gnd.n5056 240.244
R12724 gnd.n5054 gnd.n4881 240.244
R12725 gnd.n5050 gnd.n5048 240.244
R12726 gnd.n5046 gnd.n4887 240.244
R12727 gnd.n5042 gnd.n5040 240.244
R12728 gnd.n5038 gnd.n4893 240.244
R12729 gnd.n5034 gnd.n5032 240.244
R12730 gnd.n5030 gnd.n4899 240.244
R12731 gnd.n5026 gnd.n5024 240.244
R12732 gnd.n5022 gnd.n4908 240.244
R12733 gnd.n5018 gnd.n5016 240.244
R12734 gnd.n5014 gnd.n4914 240.244
R12735 gnd.n5010 gnd.n5008 240.244
R12736 gnd.n5006 gnd.n4920 240.244
R12737 gnd.n5002 gnd.n5000 240.244
R12738 gnd.n4998 gnd.n4926 240.244
R12739 gnd.n4988 gnd.n4931 240.244
R12740 gnd.n5069 gnd.n1981 240.244
R12741 gnd.n5079 gnd.n1981 240.244
R12742 gnd.n5079 gnd.n1977 240.244
R12743 gnd.n5085 gnd.n1977 240.244
R12744 gnd.n5085 gnd.n1965 240.244
R12745 gnd.n5095 gnd.n1965 240.244
R12746 gnd.n5095 gnd.n1961 240.244
R12747 gnd.n5101 gnd.n1961 240.244
R12748 gnd.n5101 gnd.n1949 240.244
R12749 gnd.n5111 gnd.n1949 240.244
R12750 gnd.n5111 gnd.n1945 240.244
R12751 gnd.n5117 gnd.n1945 240.244
R12752 gnd.n5117 gnd.n1933 240.244
R12753 gnd.n5127 gnd.n1933 240.244
R12754 gnd.n5127 gnd.n1929 240.244
R12755 gnd.n5133 gnd.n1929 240.244
R12756 gnd.n5133 gnd.n1916 240.244
R12757 gnd.n5151 gnd.n1916 240.244
R12758 gnd.n5151 gnd.n1911 240.244
R12759 gnd.n5159 gnd.n1911 240.244
R12760 gnd.n5159 gnd.n1912 240.244
R12761 gnd.n1912 gnd.n1880 240.244
R12762 gnd.n5191 gnd.n1880 240.244
R12763 gnd.n5191 gnd.n1881 240.244
R12764 gnd.n1881 gnd.n1875 240.244
R12765 gnd.n5198 gnd.n1875 240.244
R12766 gnd.n5198 gnd.n1876 240.244
R12767 gnd.n1876 gnd.n1771 240.244
R12768 gnd.n5462 gnd.n1771 240.244
R12769 gnd.n5462 gnd.n1772 240.244
R12770 gnd.n5454 gnd.n1772 240.244
R12771 gnd.n5454 gnd.n5451 240.244
R12772 gnd.n5451 gnd.n5448 240.244
R12773 gnd.n5448 gnd.n1787 240.244
R12774 gnd.n5440 gnd.n1787 240.244
R12775 gnd.n5440 gnd.n1762 240.244
R12776 gnd.n5468 gnd.n1762 240.244
R12777 gnd.n5468 gnd.n1749 240.244
R12778 gnd.n5478 gnd.n1749 240.244
R12779 gnd.n5478 gnd.n1745 240.244
R12780 gnd.n5484 gnd.n1745 240.244
R12781 gnd.n5484 gnd.n1732 240.244
R12782 gnd.n5494 gnd.n1732 240.244
R12783 gnd.n5494 gnd.n1728 240.244
R12784 gnd.n5500 gnd.n1728 240.244
R12785 gnd.n5500 gnd.n1715 240.244
R12786 gnd.n5510 gnd.n1715 240.244
R12787 gnd.n5510 gnd.n1711 240.244
R12788 gnd.n5516 gnd.n1711 240.244
R12789 gnd.n5516 gnd.n1698 240.244
R12790 gnd.n5526 gnd.n1698 240.244
R12791 gnd.n5526 gnd.n1694 240.244
R12792 gnd.n5532 gnd.n1694 240.244
R12793 gnd.n5532 gnd.n1681 240.244
R12794 gnd.n5542 gnd.n1681 240.244
R12795 gnd.n5542 gnd.n1677 240.244
R12796 gnd.n5548 gnd.n1677 240.244
R12797 gnd.n5548 gnd.n1664 240.244
R12798 gnd.n5558 gnd.n1664 240.244
R12799 gnd.n5558 gnd.n1659 240.244
R12800 gnd.n5566 gnd.n1659 240.244
R12801 gnd.n5566 gnd.n1660 240.244
R12802 gnd.n1660 gnd.n1358 240.244
R12803 gnd.n5770 gnd.n1358 240.244
R12804 gnd.n4754 gnd.n2012 240.244
R12805 gnd.n4747 gnd.n4746 240.244
R12806 gnd.n4744 gnd.n4743 240.244
R12807 gnd.n4740 gnd.n4739 240.244
R12808 gnd.n4736 gnd.n4735 240.244
R12809 gnd.n4732 gnd.n4731 240.244
R12810 gnd.n4728 gnd.n4727 240.244
R12811 gnd.n4724 gnd.n4723 240.244
R12812 gnd.n4061 gnd.n3773 240.244
R12813 gnd.n4071 gnd.n3773 240.244
R12814 gnd.n4071 gnd.n3764 240.244
R12815 gnd.n3764 gnd.n3753 240.244
R12816 gnd.n4092 gnd.n3753 240.244
R12817 gnd.n4092 gnd.n3747 240.244
R12818 gnd.n4102 gnd.n3747 240.244
R12819 gnd.n4102 gnd.n3736 240.244
R12820 gnd.n3736 gnd.n3726 240.244
R12821 gnd.n4128 gnd.n3726 240.244
R12822 gnd.n4129 gnd.n4128 240.244
R12823 gnd.n4130 gnd.n4129 240.244
R12824 gnd.n4130 gnd.n3705 240.244
R12825 gnd.n4166 gnd.n3705 240.244
R12826 gnd.n4166 gnd.n3706 240.244
R12827 gnd.n4162 gnd.n3706 240.244
R12828 gnd.n4162 gnd.n4161 240.244
R12829 gnd.n4161 gnd.n3530 240.244
R12830 gnd.n4196 gnd.n3530 240.244
R12831 gnd.n4196 gnd.n3521 240.244
R12832 gnd.n3521 gnd.n3513 240.244
R12833 gnd.n4217 gnd.n3513 240.244
R12834 gnd.n4217 gnd.n3507 240.244
R12835 gnd.n4227 gnd.n3507 240.244
R12836 gnd.n4227 gnd.n3498 240.244
R12837 gnd.n3498 gnd.n3488 240.244
R12838 gnd.n4248 gnd.n3488 240.244
R12839 gnd.n4248 gnd.n3481 240.244
R12840 gnd.n4258 gnd.n3481 240.244
R12841 gnd.n4258 gnd.n3472 240.244
R12842 gnd.n3472 gnd.n3461 240.244
R12843 gnd.n4279 gnd.n3461 240.244
R12844 gnd.n4279 gnd.n3455 240.244
R12845 gnd.n4289 gnd.n3455 240.244
R12846 gnd.n4289 gnd.n3447 240.244
R12847 gnd.n3447 gnd.n3437 240.244
R12848 gnd.n4310 gnd.n3437 240.244
R12849 gnd.n4310 gnd.n3431 240.244
R12850 gnd.n4320 gnd.n3431 240.244
R12851 gnd.n4320 gnd.n3422 240.244
R12852 gnd.n3422 gnd.n3411 240.244
R12853 gnd.n4341 gnd.n3411 240.244
R12854 gnd.n4341 gnd.n3405 240.244
R12855 gnd.n4351 gnd.n3405 240.244
R12856 gnd.n4351 gnd.n3396 240.244
R12857 gnd.n3396 gnd.n3386 240.244
R12858 gnd.n4372 gnd.n3386 240.244
R12859 gnd.n4372 gnd.n3379 240.244
R12860 gnd.n4638 gnd.n3379 240.244
R12861 gnd.n4638 gnd.n3371 240.244
R12862 gnd.n3371 gnd.n3361 240.244
R12863 gnd.n4658 gnd.n3361 240.244
R12864 gnd.n4658 gnd.n3363 240.244
R12865 gnd.n4051 gnd.n3786 240.244
R12866 gnd.n3807 gnd.n3786 240.244
R12867 gnd.n3810 gnd.n3809 240.244
R12868 gnd.n3817 gnd.n3816 240.244
R12869 gnd.n3820 gnd.n3819 240.244
R12870 gnd.n3827 gnd.n3826 240.244
R12871 gnd.n3830 gnd.n3829 240.244
R12872 gnd.n3837 gnd.n3836 240.244
R12873 gnd.n4059 gnd.n3783 240.244
R12874 gnd.n3783 gnd.n3762 240.244
R12875 gnd.n4082 gnd.n3762 240.244
R12876 gnd.n4082 gnd.n3756 240.244
R12877 gnd.n4090 gnd.n3756 240.244
R12878 gnd.n4090 gnd.n3758 240.244
R12879 gnd.n3758 gnd.n3734 240.244
R12880 gnd.n4112 gnd.n3734 240.244
R12881 gnd.n4112 gnd.n3729 240.244
R12882 gnd.n4126 gnd.n3729 240.244
R12883 gnd.n4126 gnd.n3730 240.244
R12884 gnd.n4122 gnd.n3730 240.244
R12885 gnd.n4122 gnd.n3702 240.244
R12886 gnd.n4169 gnd.n3702 240.244
R12887 gnd.n4170 gnd.n4169 240.244
R12888 gnd.n4171 gnd.n4170 240.244
R12889 gnd.n4171 gnd.n3698 240.244
R12890 gnd.n4177 gnd.n3698 240.244
R12891 gnd.n4177 gnd.n3520 240.244
R12892 gnd.n4207 gnd.n3520 240.244
R12893 gnd.n4207 gnd.n3515 240.244
R12894 gnd.n4215 gnd.n3515 240.244
R12895 gnd.n4215 gnd.n3516 240.244
R12896 gnd.n3516 gnd.n3496 240.244
R12897 gnd.n4238 gnd.n3496 240.244
R12898 gnd.n4238 gnd.n3491 240.244
R12899 gnd.n4246 gnd.n3491 240.244
R12900 gnd.n4246 gnd.n3492 240.244
R12901 gnd.n3492 gnd.n3470 240.244
R12902 gnd.n4269 gnd.n3470 240.244
R12903 gnd.n4269 gnd.n3464 240.244
R12904 gnd.n4277 gnd.n3464 240.244
R12905 gnd.n4277 gnd.n3466 240.244
R12906 gnd.n3466 gnd.n3445 240.244
R12907 gnd.n4300 gnd.n3445 240.244
R12908 gnd.n4300 gnd.n3439 240.244
R12909 gnd.n4308 gnd.n3439 240.244
R12910 gnd.n4308 gnd.n3441 240.244
R12911 gnd.n3441 gnd.n3420 240.244
R12912 gnd.n4331 gnd.n3420 240.244
R12913 gnd.n4331 gnd.n3414 240.244
R12914 gnd.n4339 gnd.n3414 240.244
R12915 gnd.n4339 gnd.n3416 240.244
R12916 gnd.n3416 gnd.n3394 240.244
R12917 gnd.n4362 gnd.n3394 240.244
R12918 gnd.n4362 gnd.n3389 240.244
R12919 gnd.n4370 gnd.n3389 240.244
R12920 gnd.n4370 gnd.n3390 240.244
R12921 gnd.n3390 gnd.n3369 240.244
R12922 gnd.n4648 gnd.n3369 240.244
R12923 gnd.n4648 gnd.n3365 240.244
R12924 gnd.n4656 gnd.n3365 240.244
R12925 gnd.n4656 gnd.n2011 240.244
R12926 gnd.n2031 gnd.n1989 240.244
R12927 gnd.n4714 gnd.n4713 240.244
R12928 gnd.n4710 gnd.n4709 240.244
R12929 gnd.n4706 gnd.n4705 240.244
R12930 gnd.n4702 gnd.n4701 240.244
R12931 gnd.n4698 gnd.n4697 240.244
R12932 gnd.n4694 gnd.n4693 240.244
R12933 gnd.n4690 gnd.n4689 240.244
R12934 gnd.n4686 gnd.n4685 240.244
R12935 gnd.n4682 gnd.n4681 240.244
R12936 gnd.n4678 gnd.n4677 240.244
R12937 gnd.n4674 gnd.n4673 240.244
R12938 gnd.n4670 gnd.n4669 240.244
R12939 gnd.n3974 gnd.n3871 240.244
R12940 gnd.n3974 gnd.n3864 240.244
R12941 gnd.n3985 gnd.n3864 240.244
R12942 gnd.n3985 gnd.n3860 240.244
R12943 gnd.n3991 gnd.n3860 240.244
R12944 gnd.n3991 gnd.n3852 240.244
R12945 gnd.n4001 gnd.n3852 240.244
R12946 gnd.n4001 gnd.n3847 240.244
R12947 gnd.n4037 gnd.n3847 240.244
R12948 gnd.n4037 gnd.n3848 240.244
R12949 gnd.n3848 gnd.n3795 240.244
R12950 gnd.n4032 gnd.n3795 240.244
R12951 gnd.n4032 gnd.n4031 240.244
R12952 gnd.n4031 gnd.n3774 240.244
R12953 gnd.n4027 gnd.n3774 240.244
R12954 gnd.n4027 gnd.n3765 240.244
R12955 gnd.n4024 gnd.n3765 240.244
R12956 gnd.n4024 gnd.n4023 240.244
R12957 gnd.n4023 gnd.n3748 240.244
R12958 gnd.n4019 gnd.n3748 240.244
R12959 gnd.n4019 gnd.n3737 240.244
R12960 gnd.n3737 gnd.n3717 240.244
R12961 gnd.n4138 gnd.n3717 240.244
R12962 gnd.n4138 gnd.n3712 240.244
R12963 gnd.n4146 gnd.n3712 240.244
R12964 gnd.n4146 gnd.n3713 240.244
R12965 gnd.n3713 gnd.n3681 240.244
R12966 gnd.n4186 gnd.n3681 240.244
R12967 gnd.n4186 gnd.n3682 240.244
R12968 gnd.n3697 gnd.n3682 240.244
R12969 gnd.n3697 gnd.n3532 240.244
R12970 gnd.n4193 gnd.n3532 240.244
R12971 gnd.n4193 gnd.n3522 240.244
R12972 gnd.n3611 gnd.n3522 240.244
R12973 gnd.n3614 gnd.n3611 240.244
R12974 gnd.n3614 gnd.n3508 240.244
R12975 gnd.n3608 gnd.n3508 240.244
R12976 gnd.n3608 gnd.n3499 240.244
R12977 gnd.n3605 gnd.n3499 240.244
R12978 gnd.n3605 gnd.n3604 240.244
R12979 gnd.n3604 gnd.n3483 240.244
R12980 gnd.n3600 gnd.n3483 240.244
R12981 gnd.n3600 gnd.n3473 240.244
R12982 gnd.n3597 gnd.n3473 240.244
R12983 gnd.n3597 gnd.n3596 240.244
R12984 gnd.n3596 gnd.n3456 240.244
R12985 gnd.n3592 gnd.n3456 240.244
R12986 gnd.n3592 gnd.n3448 240.244
R12987 gnd.n3589 gnd.n3448 240.244
R12988 gnd.n3589 gnd.n3586 240.244
R12989 gnd.n3586 gnd.n3432 240.244
R12990 gnd.n3582 gnd.n3432 240.244
R12991 gnd.n3582 gnd.n3423 240.244
R12992 gnd.n3579 gnd.n3423 240.244
R12993 gnd.n3579 gnd.n3578 240.244
R12994 gnd.n3578 gnd.n3406 240.244
R12995 gnd.n3574 gnd.n3406 240.244
R12996 gnd.n3574 gnd.n3397 240.244
R12997 gnd.n3571 gnd.n3397 240.244
R12998 gnd.n3571 gnd.n3570 240.244
R12999 gnd.n3570 gnd.n3381 240.244
R13000 gnd.n3566 gnd.n3381 240.244
R13001 gnd.n3566 gnd.n3372 240.244
R13002 gnd.n3372 gnd.n2060 240.244
R13003 gnd.n4665 gnd.n2060 240.244
R13004 gnd.n3888 gnd.n3887 240.244
R13005 gnd.n3959 gnd.n3887 240.244
R13006 gnd.n3957 gnd.n3956 240.244
R13007 gnd.n3953 gnd.n3952 240.244
R13008 gnd.n3949 gnd.n3948 240.244
R13009 gnd.n3945 gnd.n3944 240.244
R13010 gnd.n3941 gnd.n3940 240.244
R13011 gnd.n3937 gnd.n3936 240.244
R13012 gnd.n3933 gnd.n3932 240.244
R13013 gnd.n3929 gnd.n3928 240.244
R13014 gnd.n3925 gnd.n3924 240.244
R13015 gnd.n3921 gnd.n3920 240.244
R13016 gnd.n3917 gnd.n3875 240.244
R13017 gnd.n3977 gnd.n3869 240.244
R13018 gnd.n3977 gnd.n3865 240.244
R13019 gnd.n3983 gnd.n3865 240.244
R13020 gnd.n3983 gnd.n3858 240.244
R13021 gnd.n3993 gnd.n3858 240.244
R13022 gnd.n3993 gnd.n3854 240.244
R13023 gnd.n3999 gnd.n3854 240.244
R13024 gnd.n3999 gnd.n3845 240.244
R13025 gnd.n4039 gnd.n3845 240.244
R13026 gnd.n4039 gnd.n3796 240.244
R13027 gnd.n4047 gnd.n3796 240.244
R13028 gnd.n4047 gnd.n3797 240.244
R13029 gnd.n3797 gnd.n3775 240.244
R13030 gnd.n4068 gnd.n3775 240.244
R13031 gnd.n4068 gnd.n3767 240.244
R13032 gnd.n4079 gnd.n3767 240.244
R13033 gnd.n4079 gnd.n3768 240.244
R13034 gnd.n3768 gnd.n3749 240.244
R13035 gnd.n4099 gnd.n3749 240.244
R13036 gnd.n4099 gnd.n3739 240.244
R13037 gnd.n4109 gnd.n3739 240.244
R13038 gnd.n4109 gnd.n3720 240.244
R13039 gnd.n4136 gnd.n3720 240.244
R13040 gnd.n4136 gnd.n3710 240.244
R13041 gnd.n4149 gnd.n3710 240.244
R13042 gnd.n4150 gnd.n4149 240.244
R13043 gnd.n4150 gnd.n3685 240.244
R13044 gnd.n4184 gnd.n3685 240.244
R13045 gnd.n4184 gnd.n3686 240.244
R13046 gnd.n4180 gnd.n3686 240.244
R13047 gnd.n4180 gnd.n3694 240.244
R13048 gnd.n3694 gnd.n3524 240.244
R13049 gnd.n4204 gnd.n3524 240.244
R13050 gnd.n4204 gnd.n3525 240.244
R13051 gnd.n3525 gnd.n3509 240.244
R13052 gnd.n4224 gnd.n3509 240.244
R13053 gnd.n4224 gnd.n3501 240.244
R13054 gnd.n4235 gnd.n3501 240.244
R13055 gnd.n4235 gnd.n3502 240.244
R13056 gnd.n3502 gnd.n3484 240.244
R13057 gnd.n4255 gnd.n3484 240.244
R13058 gnd.n4255 gnd.n3475 240.244
R13059 gnd.n4266 gnd.n3475 240.244
R13060 gnd.n4266 gnd.n3476 240.244
R13061 gnd.n3476 gnd.n3457 240.244
R13062 gnd.n4286 gnd.n3457 240.244
R13063 gnd.n4286 gnd.n3449 240.244
R13064 gnd.n4297 gnd.n3449 240.244
R13065 gnd.n4297 gnd.n3450 240.244
R13066 gnd.n3450 gnd.n3433 240.244
R13067 gnd.n4317 gnd.n3433 240.244
R13068 gnd.n4317 gnd.n3425 240.244
R13069 gnd.n4328 gnd.n3425 240.244
R13070 gnd.n4328 gnd.n3426 240.244
R13071 gnd.n3426 gnd.n3407 240.244
R13072 gnd.n4348 gnd.n3407 240.244
R13073 gnd.n4348 gnd.n3399 240.244
R13074 gnd.n4359 gnd.n3399 240.244
R13075 gnd.n4359 gnd.n3400 240.244
R13076 gnd.n3400 gnd.n3382 240.244
R13077 gnd.n4635 gnd.n3382 240.244
R13078 gnd.n4635 gnd.n3374 240.244
R13079 gnd.n4645 gnd.n3374 240.244
R13080 gnd.n4645 gnd.n3356 240.244
R13081 gnd.n4663 gnd.n3356 240.244
R13082 gnd.n7418 gnd.n7417 240.244
R13083 gnd.n7423 gnd.n7420 240.244
R13084 gnd.n7426 gnd.n7425 240.244
R13085 gnd.n7431 gnd.n7428 240.244
R13086 gnd.n7434 gnd.n7433 240.244
R13087 gnd.n7439 gnd.n7436 240.244
R13088 gnd.n7442 gnd.n7441 240.244
R13089 gnd.n7446 gnd.n7444 240.244
R13090 gnd.n7449 gnd.n7448 240.244
R13091 gnd.n6973 gnd.n482 240.244
R13092 gnd.n568 gnd.n482 240.244
R13093 gnd.n568 gnd.n473 240.244
R13094 gnd.n569 gnd.n473 240.244
R13095 gnd.n569 gnd.n464 240.244
R13096 gnd.n572 gnd.n464 240.244
R13097 gnd.n572 gnd.n455 240.244
R13098 gnd.n573 gnd.n455 240.244
R13099 gnd.n573 gnd.n448 240.244
R13100 gnd.n576 gnd.n448 240.244
R13101 gnd.n576 gnd.n439 240.244
R13102 gnd.n577 gnd.n439 240.244
R13103 gnd.n577 gnd.n430 240.244
R13104 gnd.n580 gnd.n430 240.244
R13105 gnd.n580 gnd.n421 240.244
R13106 gnd.n581 gnd.n421 240.244
R13107 gnd.n581 gnd.n414 240.244
R13108 gnd.n584 gnd.n414 240.244
R13109 gnd.n584 gnd.n403 240.244
R13110 gnd.n6939 gnd.n403 240.244
R13111 gnd.n6939 gnd.n385 240.244
R13112 gnd.n7160 gnd.n385 240.244
R13113 gnd.n7160 gnd.n371 240.244
R13114 gnd.n380 gnd.n371 240.244
R13115 gnd.n7168 gnd.n380 240.244
R13116 gnd.n7168 gnd.n360 240.244
R13117 gnd.n360 gnd.n351 240.244
R13118 gnd.n7210 gnd.n351 240.244
R13119 gnd.n7210 gnd.n310 240.244
R13120 gnd.n7203 gnd.n310 240.244
R13121 gnd.n7203 gnd.n341 240.244
R13122 gnd.n341 gnd.n340 240.244
R13123 gnd.n340 gnd.n78 240.244
R13124 gnd.n79 gnd.n78 240.244
R13125 gnd.n80 gnd.n79 240.244
R13126 gnd.n325 gnd.n80 240.244
R13127 gnd.n325 gnd.n83 240.244
R13128 gnd.n84 gnd.n83 240.244
R13129 gnd.n85 gnd.n84 240.244
R13130 gnd.n288 gnd.n85 240.244
R13131 gnd.n288 gnd.n88 240.244
R13132 gnd.n89 gnd.n88 240.244
R13133 gnd.n90 gnd.n89 240.244
R13134 gnd.n273 gnd.n90 240.244
R13135 gnd.n273 gnd.n93 240.244
R13136 gnd.n94 gnd.n93 240.244
R13137 gnd.n95 gnd.n94 240.244
R13138 gnd.n258 gnd.n95 240.244
R13139 gnd.n258 gnd.n98 240.244
R13140 gnd.n99 gnd.n98 240.244
R13141 gnd.n100 gnd.n99 240.244
R13142 gnd.n243 gnd.n100 240.244
R13143 gnd.n243 gnd.n103 240.244
R13144 gnd.n104 gnd.n103 240.244
R13145 gnd.n105 gnd.n104 240.244
R13146 gnd.n227 gnd.n105 240.244
R13147 gnd.n227 gnd.n108 240.244
R13148 gnd.n109 gnd.n108 240.244
R13149 gnd.n110 gnd.n109 240.244
R13150 gnd.n211 gnd.n110 240.244
R13151 gnd.n211 gnd.n113 240.244
R13152 gnd.n114 gnd.n113 240.244
R13153 gnd.n115 gnd.n114 240.244
R13154 gnd.n7574 gnd.n115 240.244
R13155 gnd.n6625 gnd.n6624 240.244
R13156 gnd.n6627 gnd.n6626 240.244
R13157 gnd.n6637 gnd.n6636 240.244
R13158 gnd.n6645 gnd.n6644 240.244
R13159 gnd.n6647 gnd.n6646 240.244
R13160 gnd.n6657 gnd.n6656 240.244
R13161 gnd.n6665 gnd.n6664 240.244
R13162 gnd.n6667 gnd.n6666 240.244
R13163 gnd.n6711 gnd.n517 240.244
R13164 gnd.n7056 gnd.n479 240.244
R13165 gnd.n7056 gnd.n475 240.244
R13166 gnd.n7062 gnd.n475 240.244
R13167 gnd.n7062 gnd.n461 240.244
R13168 gnd.n7072 gnd.n461 240.244
R13169 gnd.n7072 gnd.n457 240.244
R13170 gnd.n7078 gnd.n457 240.244
R13171 gnd.n7078 gnd.n445 240.244
R13172 gnd.n7088 gnd.n445 240.244
R13173 gnd.n7088 gnd.n441 240.244
R13174 gnd.n7094 gnd.n441 240.244
R13175 gnd.n7094 gnd.n427 240.244
R13176 gnd.n7104 gnd.n427 240.244
R13177 gnd.n7104 gnd.n423 240.244
R13178 gnd.n7110 gnd.n423 240.244
R13179 gnd.n7110 gnd.n411 240.244
R13180 gnd.n7120 gnd.n411 240.244
R13181 gnd.n7120 gnd.n405 240.244
R13182 gnd.n7129 gnd.n405 240.244
R13183 gnd.n7129 gnd.n406 240.244
R13184 gnd.n406 gnd.n395 240.244
R13185 gnd.n395 gnd.n373 240.244
R13186 gnd.n7180 gnd.n373 240.244
R13187 gnd.n7180 gnd.n374 240.244
R13188 gnd.n7170 gnd.n374 240.244
R13189 gnd.n7170 gnd.n362 240.244
R13190 gnd.n7171 gnd.n362 240.244
R13191 gnd.n7171 gnd.n312 240.244
R13192 gnd.n7319 gnd.n312 240.244
R13193 gnd.n7319 gnd.n313 240.244
R13194 gnd.n318 gnd.n313 240.244
R13195 gnd.n319 gnd.n318 240.244
R13196 gnd.n320 gnd.n319 240.244
R13197 gnd.n329 gnd.n320 240.244
R13198 gnd.n329 gnd.n323 240.244
R13199 gnd.n7306 gnd.n323 240.244
R13200 gnd.n7306 gnd.n294 240.244
R13201 gnd.n7330 gnd.n294 240.244
R13202 gnd.n7330 gnd.n290 240.244
R13203 gnd.n7336 gnd.n290 240.244
R13204 gnd.n7336 gnd.n278 240.244
R13205 gnd.n7346 gnd.n278 240.244
R13206 gnd.n7346 gnd.n274 240.244
R13207 gnd.n7352 gnd.n274 240.244
R13208 gnd.n7352 gnd.n264 240.244
R13209 gnd.n7362 gnd.n264 240.244
R13210 gnd.n7362 gnd.n260 240.244
R13211 gnd.n7368 gnd.n260 240.244
R13212 gnd.n7368 gnd.n248 240.244
R13213 gnd.n7378 gnd.n248 240.244
R13214 gnd.n7378 gnd.n244 240.244
R13215 gnd.n7384 gnd.n244 240.244
R13216 gnd.n7384 gnd.n233 240.244
R13217 gnd.n7394 gnd.n233 240.244
R13218 gnd.n7394 gnd.n229 240.244
R13219 gnd.n7400 gnd.n229 240.244
R13220 gnd.n7400 gnd.n218 240.244
R13221 gnd.n7410 gnd.n218 240.244
R13222 gnd.n7410 gnd.n212 240.244
R13223 gnd.n7484 gnd.n212 240.244
R13224 gnd.n7484 gnd.n213 240.244
R13225 gnd.n213 gnd.n203 240.244
R13226 gnd.n7415 gnd.n203 240.244
R13227 gnd.n7415 gnd.n125 240.244
R13228 gnd.n5576 gnd.n5575 240.244
R13229 gnd.n5587 gnd.n5578 240.244
R13230 gnd.n5590 gnd.n5589 240.244
R13231 gnd.n5601 gnd.n5600 240.244
R13232 gnd.n5610 gnd.n5603 240.244
R13233 gnd.n5613 gnd.n5612 240.244
R13234 gnd.n5624 gnd.n5623 240.244
R13235 gnd.n5629 gnd.n5626 240.244
R13236 gnd.n5627 gnd.n1350 240.244
R13237 gnd.n4871 gnd.n4758 240.244
R13238 gnd.n4871 gnd.n1983 240.244
R13239 gnd.n4867 gnd.n1983 240.244
R13240 gnd.n4867 gnd.n1976 240.244
R13241 gnd.n4864 gnd.n1976 240.244
R13242 gnd.n4864 gnd.n1968 240.244
R13243 gnd.n4861 gnd.n1968 240.244
R13244 gnd.n4861 gnd.n1959 240.244
R13245 gnd.n4858 gnd.n1959 240.244
R13246 gnd.n4858 gnd.n1951 240.244
R13247 gnd.n4855 gnd.n1951 240.244
R13248 gnd.n4855 gnd.n1944 240.244
R13249 gnd.n4852 gnd.n1944 240.244
R13250 gnd.n4852 gnd.n1936 240.244
R13251 gnd.n4849 gnd.n1936 240.244
R13252 gnd.n4849 gnd.n1927 240.244
R13253 gnd.n4846 gnd.n1927 240.244
R13254 gnd.n4846 gnd.n1918 240.244
R13255 gnd.n1918 gnd.n1907 240.244
R13256 gnd.n5161 gnd.n1907 240.244
R13257 gnd.n5161 gnd.n1903 240.244
R13258 gnd.n5172 gnd.n1903 240.244
R13259 gnd.n5172 gnd.n1883 240.244
R13260 gnd.n5168 gnd.n1883 240.244
R13261 gnd.n5168 gnd.n1872 240.244
R13262 gnd.n5200 gnd.n1872 240.244
R13263 gnd.n5200 gnd.n1868 240.244
R13264 gnd.n5216 gnd.n1868 240.244
R13265 gnd.n5216 gnd.n1774 240.244
R13266 gnd.n5212 gnd.n1774 240.244
R13267 gnd.n5212 gnd.n1785 240.244
R13268 gnd.n5208 gnd.n1785 240.244
R13269 gnd.n5208 gnd.n1790 240.244
R13270 gnd.n5234 gnd.n1790 240.244
R13271 gnd.n5234 gnd.n1797 240.244
R13272 gnd.n5240 gnd.n1797 240.244
R13273 gnd.n5240 gnd.n1760 240.244
R13274 gnd.n5428 gnd.n1760 240.244
R13275 gnd.n5428 gnd.n1751 240.244
R13276 gnd.n1811 gnd.n1751 240.244
R13277 gnd.n1811 gnd.n1744 240.244
R13278 gnd.n1812 gnd.n1744 240.244
R13279 gnd.n1812 gnd.n1735 240.244
R13280 gnd.n1815 gnd.n1735 240.244
R13281 gnd.n1815 gnd.n1726 240.244
R13282 gnd.n1816 gnd.n1726 240.244
R13283 gnd.n1816 gnd.n1717 240.244
R13284 gnd.n1819 gnd.n1717 240.244
R13285 gnd.n1819 gnd.n1710 240.244
R13286 gnd.n1820 gnd.n1710 240.244
R13287 gnd.n1820 gnd.n1701 240.244
R13288 gnd.n1823 gnd.n1701 240.244
R13289 gnd.n1823 gnd.n1692 240.244
R13290 gnd.n1824 gnd.n1692 240.244
R13291 gnd.n1824 gnd.n1683 240.244
R13292 gnd.n1827 gnd.n1683 240.244
R13293 gnd.n1827 gnd.n1676 240.244
R13294 gnd.n1828 gnd.n1676 240.244
R13295 gnd.n1828 gnd.n1667 240.244
R13296 gnd.n5385 gnd.n1667 240.244
R13297 gnd.n5385 gnd.n1657 240.244
R13298 gnd.n5387 gnd.n1657 240.244
R13299 gnd.n5387 gnd.n1352 240.244
R13300 gnd.n5772 gnd.n1352 240.244
R13301 gnd.n4784 gnd.n4782 240.244
R13302 gnd.n4790 gnd.n4776 240.244
R13303 gnd.n4794 gnd.n4792 240.244
R13304 gnd.n4800 gnd.n4772 240.244
R13305 gnd.n4804 gnd.n4802 240.244
R13306 gnd.n4810 gnd.n4768 240.244
R13307 gnd.n4814 gnd.n4812 240.244
R13308 gnd.n4820 gnd.n4764 240.244
R13309 gnd.n4823 gnd.n4822 240.244
R13310 gnd.n5071 gnd.n1984 240.244
R13311 gnd.n5077 gnd.n1984 240.244
R13312 gnd.n5077 gnd.n1973 240.244
R13313 gnd.n5087 gnd.n1973 240.244
R13314 gnd.n5087 gnd.n1969 240.244
R13315 gnd.n5093 gnd.n1969 240.244
R13316 gnd.n5093 gnd.n1956 240.244
R13317 gnd.n5103 gnd.n1956 240.244
R13318 gnd.n5103 gnd.n1952 240.244
R13319 gnd.n5109 gnd.n1952 240.244
R13320 gnd.n5109 gnd.n1941 240.244
R13321 gnd.n5119 gnd.n1941 240.244
R13322 gnd.n5119 gnd.n1937 240.244
R13323 gnd.n5125 gnd.n1937 240.244
R13324 gnd.n5125 gnd.n1924 240.244
R13325 gnd.n5135 gnd.n1924 240.244
R13326 gnd.n5135 gnd.n1919 240.244
R13327 gnd.n5149 gnd.n1919 240.244
R13328 gnd.n5149 gnd.n1920 240.244
R13329 gnd.n1920 gnd.n1910 240.244
R13330 gnd.n5144 gnd.n1910 240.244
R13331 gnd.n5144 gnd.n1885 240.244
R13332 gnd.n5189 gnd.n1885 240.244
R13333 gnd.n5189 gnd.n1886 240.244
R13334 gnd.n5185 gnd.n1886 240.244
R13335 gnd.n5185 gnd.n1874 240.244
R13336 gnd.n1894 gnd.n1874 240.244
R13337 gnd.n1894 gnd.n1776 240.244
R13338 gnd.n5460 gnd.n1776 240.244
R13339 gnd.n5460 gnd.n1777 240.244
R13340 gnd.n5456 gnd.n1777 240.244
R13341 gnd.n5456 gnd.n1783 240.244
R13342 gnd.n5446 gnd.n1783 240.244
R13343 gnd.n5446 gnd.n1791 240.244
R13344 gnd.n5442 gnd.n1791 240.244
R13345 gnd.n5442 gnd.n1757 240.244
R13346 gnd.n5470 gnd.n1757 240.244
R13347 gnd.n5470 gnd.n1753 240.244
R13348 gnd.n5476 gnd.n1753 240.244
R13349 gnd.n5476 gnd.n1741 240.244
R13350 gnd.n5486 gnd.n1741 240.244
R13351 gnd.n5486 gnd.n1737 240.244
R13352 gnd.n5492 gnd.n1737 240.244
R13353 gnd.n5492 gnd.n1723 240.244
R13354 gnd.n5502 gnd.n1723 240.244
R13355 gnd.n5502 gnd.n1719 240.244
R13356 gnd.n5508 gnd.n1719 240.244
R13357 gnd.n5508 gnd.n1707 240.244
R13358 gnd.n5518 gnd.n1707 240.244
R13359 gnd.n5518 gnd.n1703 240.244
R13360 gnd.n5524 gnd.n1703 240.244
R13361 gnd.n5524 gnd.n1689 240.244
R13362 gnd.n5534 gnd.n1689 240.244
R13363 gnd.n5534 gnd.n1685 240.244
R13364 gnd.n5540 gnd.n1685 240.244
R13365 gnd.n5540 gnd.n1673 240.244
R13366 gnd.n5550 gnd.n1673 240.244
R13367 gnd.n5550 gnd.n1669 240.244
R13368 gnd.n5556 gnd.n1669 240.244
R13369 gnd.n5556 gnd.n1654 240.244
R13370 gnd.n5568 gnd.n1654 240.244
R13371 gnd.n5568 gnd.n1650 240.244
R13372 gnd.n5693 gnd.n1650 240.244
R13373 gnd.n5693 gnd.n1357 240.244
R13374 gnd.n3140 gnd.n2190 240.244
R13375 gnd.n3134 gnd.n2190 240.244
R13376 gnd.n3134 gnd.n2194 240.244
R13377 gnd.n3130 gnd.n2194 240.244
R13378 gnd.n3130 gnd.n2196 240.244
R13379 gnd.n3126 gnd.n2196 240.244
R13380 gnd.n3126 gnd.n2201 240.244
R13381 gnd.n3122 gnd.n2201 240.244
R13382 gnd.n3122 gnd.n2203 240.244
R13383 gnd.n3118 gnd.n2203 240.244
R13384 gnd.n3118 gnd.n2209 240.244
R13385 gnd.n3114 gnd.n2209 240.244
R13386 gnd.n3114 gnd.n2211 240.244
R13387 gnd.n3110 gnd.n2211 240.244
R13388 gnd.n3110 gnd.n2217 240.244
R13389 gnd.n3106 gnd.n2217 240.244
R13390 gnd.n3106 gnd.n2219 240.244
R13391 gnd.n3102 gnd.n2219 240.244
R13392 gnd.n3102 gnd.n2225 240.244
R13393 gnd.n3098 gnd.n2225 240.244
R13394 gnd.n3098 gnd.n2227 240.244
R13395 gnd.n3094 gnd.n2227 240.244
R13396 gnd.n3094 gnd.n2233 240.244
R13397 gnd.n3090 gnd.n2233 240.244
R13398 gnd.n3090 gnd.n2235 240.244
R13399 gnd.n3086 gnd.n2235 240.244
R13400 gnd.n3086 gnd.n2241 240.244
R13401 gnd.n3082 gnd.n2241 240.244
R13402 gnd.n3082 gnd.n2243 240.244
R13403 gnd.n3078 gnd.n2243 240.244
R13404 gnd.n3078 gnd.n2249 240.244
R13405 gnd.n3074 gnd.n2249 240.244
R13406 gnd.n3074 gnd.n2251 240.244
R13407 gnd.n3070 gnd.n2251 240.244
R13408 gnd.n3070 gnd.n2257 240.244
R13409 gnd.n3066 gnd.n2257 240.244
R13410 gnd.n3066 gnd.n2259 240.244
R13411 gnd.n3062 gnd.n2259 240.244
R13412 gnd.n3062 gnd.n2265 240.244
R13413 gnd.n3058 gnd.n2265 240.244
R13414 gnd.n3058 gnd.n2267 240.244
R13415 gnd.n3054 gnd.n2267 240.244
R13416 gnd.n3054 gnd.n2273 240.244
R13417 gnd.n3050 gnd.n2273 240.244
R13418 gnd.n3050 gnd.n2275 240.244
R13419 gnd.n3046 gnd.n2275 240.244
R13420 gnd.n3046 gnd.n2281 240.244
R13421 gnd.n3042 gnd.n2281 240.244
R13422 gnd.n3042 gnd.n2283 240.244
R13423 gnd.n3038 gnd.n2283 240.244
R13424 gnd.n3038 gnd.n2289 240.244
R13425 gnd.n3034 gnd.n2289 240.244
R13426 gnd.n3034 gnd.n2291 240.244
R13427 gnd.n3030 gnd.n2291 240.244
R13428 gnd.n3030 gnd.n2297 240.244
R13429 gnd.n3026 gnd.n2297 240.244
R13430 gnd.n3026 gnd.n2299 240.244
R13431 gnd.n3022 gnd.n2299 240.244
R13432 gnd.n3022 gnd.n2305 240.244
R13433 gnd.n3018 gnd.n2305 240.244
R13434 gnd.n3018 gnd.n2307 240.244
R13435 gnd.n3014 gnd.n2307 240.244
R13436 gnd.n3014 gnd.n2313 240.244
R13437 gnd.n3010 gnd.n2313 240.244
R13438 gnd.n3010 gnd.n2315 240.244
R13439 gnd.n3006 gnd.n2315 240.244
R13440 gnd.n3006 gnd.n2321 240.244
R13441 gnd.n3002 gnd.n2321 240.244
R13442 gnd.n3002 gnd.n2323 240.244
R13443 gnd.n2998 gnd.n2323 240.244
R13444 gnd.n2998 gnd.n2329 240.244
R13445 gnd.n2994 gnd.n2329 240.244
R13446 gnd.n2994 gnd.n2331 240.244
R13447 gnd.n2990 gnd.n2331 240.244
R13448 gnd.n2990 gnd.n2337 240.244
R13449 gnd.n2986 gnd.n2337 240.244
R13450 gnd.n2986 gnd.n2339 240.244
R13451 gnd.n2982 gnd.n2339 240.244
R13452 gnd.n2982 gnd.n2345 240.244
R13453 gnd.n2978 gnd.n2345 240.244
R13454 gnd.n2978 gnd.n2347 240.244
R13455 gnd.n2974 gnd.n2347 240.244
R13456 gnd.n2974 gnd.n2353 240.244
R13457 gnd.n2970 gnd.n2353 240.244
R13458 gnd.n2970 gnd.n2355 240.244
R13459 gnd.n2966 gnd.n2355 240.244
R13460 gnd.n2966 gnd.n2361 240.244
R13461 gnd.n2962 gnd.n2361 240.244
R13462 gnd.n2962 gnd.n2363 240.244
R13463 gnd.n2958 gnd.n2363 240.244
R13464 gnd.n2958 gnd.n2369 240.244
R13465 gnd.n2954 gnd.n2369 240.244
R13466 gnd.n2954 gnd.n2371 240.244
R13467 gnd.n2950 gnd.n2371 240.244
R13468 gnd.n2950 gnd.n2377 240.244
R13469 gnd.n2946 gnd.n2377 240.244
R13470 gnd.n2946 gnd.n2379 240.244
R13471 gnd.n2942 gnd.n2379 240.244
R13472 gnd.n2942 gnd.n2385 240.244
R13473 gnd.n2938 gnd.n2385 240.244
R13474 gnd.n2938 gnd.n2387 240.244
R13475 gnd.n2934 gnd.n2387 240.244
R13476 gnd.n2934 gnd.n2393 240.244
R13477 gnd.n2930 gnd.n2393 240.244
R13478 gnd.n2930 gnd.n2395 240.244
R13479 gnd.n2926 gnd.n2395 240.244
R13480 gnd.n2926 gnd.n2401 240.244
R13481 gnd.n2922 gnd.n2401 240.244
R13482 gnd.n2922 gnd.n2403 240.244
R13483 gnd.n2918 gnd.n2403 240.244
R13484 gnd.n2918 gnd.n2409 240.244
R13485 gnd.n2914 gnd.n2409 240.244
R13486 gnd.n2914 gnd.n2411 240.244
R13487 gnd.n2910 gnd.n2411 240.244
R13488 gnd.n2910 gnd.n2417 240.244
R13489 gnd.n2906 gnd.n2417 240.244
R13490 gnd.n2906 gnd.n2419 240.244
R13491 gnd.n2902 gnd.n2419 240.244
R13492 gnd.n2902 gnd.n2425 240.244
R13493 gnd.n2898 gnd.n2425 240.244
R13494 gnd.n2898 gnd.n2427 240.244
R13495 gnd.n2894 gnd.n2427 240.244
R13496 gnd.n2894 gnd.n2433 240.244
R13497 gnd.n2890 gnd.n2433 240.244
R13498 gnd.n2890 gnd.n2435 240.244
R13499 gnd.n2886 gnd.n2435 240.244
R13500 gnd.n2886 gnd.n2441 240.244
R13501 gnd.n2882 gnd.n2441 240.244
R13502 gnd.n2882 gnd.n2443 240.244
R13503 gnd.n2878 gnd.n2443 240.244
R13504 gnd.n2878 gnd.n2449 240.244
R13505 gnd.n2874 gnd.n2449 240.244
R13506 gnd.n2874 gnd.n2451 240.244
R13507 gnd.n2870 gnd.n2451 240.244
R13508 gnd.n2870 gnd.n2457 240.244
R13509 gnd.n2866 gnd.n2457 240.244
R13510 gnd.n2866 gnd.n2459 240.244
R13511 gnd.n2862 gnd.n2459 240.244
R13512 gnd.n2862 gnd.n2465 240.244
R13513 gnd.n2858 gnd.n2465 240.244
R13514 gnd.n2858 gnd.n2467 240.244
R13515 gnd.n2854 gnd.n2467 240.244
R13516 gnd.n2854 gnd.n2473 240.244
R13517 gnd.n2850 gnd.n2473 240.244
R13518 gnd.n2850 gnd.n2475 240.244
R13519 gnd.n2846 gnd.n2475 240.244
R13520 gnd.n2846 gnd.n2481 240.244
R13521 gnd.n2842 gnd.n2481 240.244
R13522 gnd.n2842 gnd.n2483 240.244
R13523 gnd.n2838 gnd.n2483 240.244
R13524 gnd.n2838 gnd.n2489 240.244
R13525 gnd.n2834 gnd.n2489 240.244
R13526 gnd.n2834 gnd.n2491 240.244
R13527 gnd.n2830 gnd.n2491 240.244
R13528 gnd.n2826 gnd.n2496 240.244
R13529 gnd.n2826 gnd.n2498 240.244
R13530 gnd.n2820 gnd.n2498 240.244
R13531 gnd.n2820 gnd.n2504 240.244
R13532 gnd.n2816 gnd.n2504 240.244
R13533 gnd.n2816 gnd.n2506 240.244
R13534 gnd.n2812 gnd.n2506 240.244
R13535 gnd.n2812 gnd.n2511 240.244
R13536 gnd.n2808 gnd.n2511 240.244
R13537 gnd.n2808 gnd.n2513 240.244
R13538 gnd.n2804 gnd.n2513 240.244
R13539 gnd.n2804 gnd.n2519 240.244
R13540 gnd.n2800 gnd.n2519 240.244
R13541 gnd.n2800 gnd.n2521 240.244
R13542 gnd.n2796 gnd.n2521 240.244
R13543 gnd.n2796 gnd.n2527 240.244
R13544 gnd.n2792 gnd.n2527 240.244
R13545 gnd.n2792 gnd.n2529 240.244
R13546 gnd.n2788 gnd.n2529 240.244
R13547 gnd.n2788 gnd.n2535 240.244
R13548 gnd.n2784 gnd.n2535 240.244
R13549 gnd.n2784 gnd.n2537 240.244
R13550 gnd.n2780 gnd.n2537 240.244
R13551 gnd.n2780 gnd.n2543 240.244
R13552 gnd.n2776 gnd.n2543 240.244
R13553 gnd.n2776 gnd.n2545 240.244
R13554 gnd.n2772 gnd.n2545 240.244
R13555 gnd.n2772 gnd.n2551 240.244
R13556 gnd.n2768 gnd.n2551 240.244
R13557 gnd.n2768 gnd.n2553 240.244
R13558 gnd.n2764 gnd.n2553 240.244
R13559 gnd.n2764 gnd.n2559 240.244
R13560 gnd.n2760 gnd.n2559 240.244
R13561 gnd.n2760 gnd.n2561 240.244
R13562 gnd.n2756 gnd.n2561 240.244
R13563 gnd.n2756 gnd.n2567 240.244
R13564 gnd.n2752 gnd.n2567 240.244
R13565 gnd.n2752 gnd.n2569 240.244
R13566 gnd.n2748 gnd.n2569 240.244
R13567 gnd.n2748 gnd.n2575 240.244
R13568 gnd.n2744 gnd.n2575 240.244
R13569 gnd.n2744 gnd.n2577 240.244
R13570 gnd.n2740 gnd.n2577 240.244
R13571 gnd.n2740 gnd.n2583 240.244
R13572 gnd.n2736 gnd.n2583 240.244
R13573 gnd.n2736 gnd.n2585 240.244
R13574 gnd.n2732 gnd.n2585 240.244
R13575 gnd.n2732 gnd.n2591 240.244
R13576 gnd.n2728 gnd.n2591 240.244
R13577 gnd.n2728 gnd.n2593 240.244
R13578 gnd.n2724 gnd.n2593 240.244
R13579 gnd.n2724 gnd.n2599 240.244
R13580 gnd.n2720 gnd.n2599 240.244
R13581 gnd.n2720 gnd.n2601 240.244
R13582 gnd.n2716 gnd.n2601 240.244
R13583 gnd.n2716 gnd.n2607 240.244
R13584 gnd.n2712 gnd.n2607 240.244
R13585 gnd.n2712 gnd.n2609 240.244
R13586 gnd.n2708 gnd.n2609 240.244
R13587 gnd.n2708 gnd.n2615 240.244
R13588 gnd.n2704 gnd.n2615 240.244
R13589 gnd.n2704 gnd.n2617 240.244
R13590 gnd.n2700 gnd.n2617 240.244
R13591 gnd.n2700 gnd.n2623 240.244
R13592 gnd.n2696 gnd.n2623 240.244
R13593 gnd.n2696 gnd.n2625 240.244
R13594 gnd.n2692 gnd.n2625 240.244
R13595 gnd.n2692 gnd.n2631 240.244
R13596 gnd.n2688 gnd.n2631 240.244
R13597 gnd.n2688 gnd.n2633 240.244
R13598 gnd.n2684 gnd.n2633 240.244
R13599 gnd.n2684 gnd.n2639 240.244
R13600 gnd.n2680 gnd.n2639 240.244
R13601 gnd.n2680 gnd.n2641 240.244
R13602 gnd.n2676 gnd.n2641 240.244
R13603 gnd.n2676 gnd.n2647 240.244
R13604 gnd.n2672 gnd.n2647 240.244
R13605 gnd.n2672 gnd.n2649 240.244
R13606 gnd.n2668 gnd.n2649 240.244
R13607 gnd.n2668 gnd.n2655 240.244
R13608 gnd.n2664 gnd.n2655 240.244
R13609 gnd.n2664 gnd.n2658 240.244
R13610 gnd.n2658 gnd.n342 240.244
R13611 gnd.n7220 gnd.n342 240.244
R13612 gnd.n5436 gnd.n1798 240.244
R13613 gnd.n5436 gnd.n1799 240.244
R13614 gnd.n5432 gnd.n1799 240.244
R13615 gnd.n5432 gnd.n5431 240.244
R13616 gnd.n5431 gnd.n1805 240.244
R13617 gnd.n5255 gnd.n1805 240.244
R13618 gnd.n5274 gnd.n5255 240.244
R13619 gnd.n5274 gnd.n5256 240.244
R13620 gnd.n5270 gnd.n5256 240.244
R13621 gnd.n5270 gnd.n5269 240.244
R13622 gnd.n5269 gnd.n1849 240.244
R13623 gnd.n5297 gnd.n1849 240.244
R13624 gnd.n5298 gnd.n5297 240.244
R13625 gnd.n5298 gnd.n1844 240.244
R13626 gnd.n5314 gnd.n1844 240.244
R13627 gnd.n5314 gnd.n1845 240.244
R13628 gnd.n5310 gnd.n1845 240.244
R13629 gnd.n5310 gnd.n5309 240.244
R13630 gnd.n5309 gnd.n1839 240.244
R13631 gnd.n5336 gnd.n1839 240.244
R13632 gnd.n5337 gnd.n5336 240.244
R13633 gnd.n5337 gnd.n1834 240.244
R13634 gnd.n5371 gnd.n1834 240.244
R13635 gnd.n5371 gnd.n1835 240.244
R13636 gnd.n5367 gnd.n1835 240.244
R13637 gnd.n5367 gnd.n5366 240.244
R13638 gnd.n5366 gnd.n5365 240.244
R13639 gnd.n5365 gnd.n5345 240.244
R13640 gnd.n5361 gnd.n5345 240.244
R13641 gnd.n5361 gnd.n5360 240.244
R13642 gnd.n5360 gnd.n5359 240.244
R13643 gnd.n5359 gnd.n5352 240.244
R13644 gnd.n5352 gnd.n1317 240.244
R13645 gnd.n5810 gnd.n1317 240.244
R13646 gnd.n5810 gnd.n1313 240.244
R13647 gnd.n5816 gnd.n1313 240.244
R13648 gnd.n5816 gnd.n1303 240.244
R13649 gnd.n5826 gnd.n1303 240.244
R13650 gnd.n5826 gnd.n1298 240.244
R13651 gnd.n5834 gnd.n1298 240.244
R13652 gnd.n5834 gnd.n1299 240.244
R13653 gnd.n1299 gnd.n1261 240.244
R13654 gnd.n5984 gnd.n1261 240.244
R13655 gnd.n5984 gnd.n1257 240.244
R13656 gnd.n5990 gnd.n1257 240.244
R13657 gnd.n5990 gnd.n1246 240.244
R13658 gnd.n6000 gnd.n1246 240.244
R13659 gnd.n6000 gnd.n1242 240.244
R13660 gnd.n6006 gnd.n1242 240.244
R13661 gnd.n6006 gnd.n1230 240.244
R13662 gnd.n6016 gnd.n1230 240.244
R13663 gnd.n6016 gnd.n1226 240.244
R13664 gnd.n6022 gnd.n1226 240.244
R13665 gnd.n6022 gnd.n1215 240.244
R13666 gnd.n6031 gnd.n1215 240.244
R13667 gnd.n6031 gnd.n1210 240.244
R13668 gnd.n6039 gnd.n1210 240.244
R13669 gnd.n6039 gnd.n1211 240.244
R13670 gnd.n1211 gnd.n1108 240.244
R13671 gnd.n6126 gnd.n1108 240.244
R13672 gnd.n6126 gnd.n1104 240.244
R13673 gnd.n6132 gnd.n1104 240.244
R13674 gnd.n6132 gnd.n1092 240.244
R13675 gnd.n6142 gnd.n1092 240.244
R13676 gnd.n6142 gnd.n1088 240.244
R13677 gnd.n6148 gnd.n1088 240.244
R13678 gnd.n6148 gnd.n1077 240.244
R13679 gnd.n6158 gnd.n1077 240.244
R13680 gnd.n6158 gnd.n1073 240.244
R13681 gnd.n6164 gnd.n1073 240.244
R13682 gnd.n6164 gnd.n1064 240.244
R13683 gnd.n6174 gnd.n1064 240.244
R13684 gnd.n6174 gnd.n1059 240.244
R13685 gnd.n6182 gnd.n1059 240.244
R13686 gnd.n6182 gnd.n1060 240.244
R13687 gnd.n1060 gnd.n1021 240.244
R13688 gnd.n6431 gnd.n1021 240.244
R13689 gnd.n6431 gnd.n1017 240.244
R13690 gnd.n6437 gnd.n1017 240.244
R13691 gnd.n6437 gnd.n1005 240.244
R13692 gnd.n6447 gnd.n1005 240.244
R13693 gnd.n6447 gnd.n1001 240.244
R13694 gnd.n6453 gnd.n1001 240.244
R13695 gnd.n6453 gnd.n989 240.244
R13696 gnd.n6463 gnd.n989 240.244
R13697 gnd.n6463 gnd.n985 240.244
R13698 gnd.n6469 gnd.n985 240.244
R13699 gnd.n6469 gnd.n975 240.244
R13700 gnd.n6479 gnd.n975 240.244
R13701 gnd.n6479 gnd.n971 240.244
R13702 gnd.n6485 gnd.n971 240.244
R13703 gnd.n6485 gnd.n960 240.244
R13704 gnd.n6495 gnd.n960 240.244
R13705 gnd.n6495 gnd.n956 240.244
R13706 gnd.n6501 gnd.n956 240.244
R13707 gnd.n6501 gnd.n944 240.244
R13708 gnd.n6511 gnd.n944 240.244
R13709 gnd.n6511 gnd.n940 240.244
R13710 gnd.n6517 gnd.n940 240.244
R13711 gnd.n6517 gnd.n927 240.244
R13712 gnd.n6533 gnd.n927 240.244
R13713 gnd.n6533 gnd.n922 240.244
R13714 gnd.n6541 gnd.n922 240.244
R13715 gnd.n6541 gnd.n923 240.244
R13716 gnd.n923 gnd.n887 240.244
R13717 gnd.n6591 gnd.n887 240.244
R13718 gnd.n6591 gnd.n882 240.244
R13719 gnd.n6599 gnd.n882 240.244
R13720 gnd.n6599 gnd.n883 240.244
R13721 gnd.n883 gnd.n660 240.244
R13722 gnd.n6782 gnd.n660 240.244
R13723 gnd.n6782 gnd.n656 240.244
R13724 gnd.n6788 gnd.n656 240.244
R13725 gnd.n6788 gnd.n645 240.244
R13726 gnd.n6799 gnd.n645 240.244
R13727 gnd.n6799 gnd.n640 240.244
R13728 gnd.n6807 gnd.n640 240.244
R13729 gnd.n6807 gnd.n641 240.244
R13730 gnd.n641 gnd.n615 240.244
R13731 gnd.n6818 gnd.n615 240.244
R13732 gnd.n6818 gnd.n611 240.244
R13733 gnd.n6824 gnd.n611 240.244
R13734 gnd.n6825 gnd.n6824 240.244
R13735 gnd.n6826 gnd.n6825 240.244
R13736 gnd.n6826 gnd.n607 240.244
R13737 gnd.n6832 gnd.n607 240.244
R13738 gnd.n6833 gnd.n6832 240.244
R13739 gnd.n6834 gnd.n6833 240.244
R13740 gnd.n6834 gnd.n603 240.244
R13741 gnd.n6840 gnd.n603 240.244
R13742 gnd.n6867 gnd.n6840 240.244
R13743 gnd.n6868 gnd.n6867 240.244
R13744 gnd.n6868 gnd.n598 240.244
R13745 gnd.n6884 gnd.n598 240.244
R13746 gnd.n6884 gnd.n599 240.244
R13747 gnd.n6880 gnd.n599 240.244
R13748 gnd.n6880 gnd.n6879 240.244
R13749 gnd.n6879 gnd.n593 240.244
R13750 gnd.n6906 gnd.n593 240.244
R13751 gnd.n6907 gnd.n6906 240.244
R13752 gnd.n6907 gnd.n588 240.244
R13753 gnd.n6915 gnd.n588 240.244
R13754 gnd.n6915 gnd.n589 240.244
R13755 gnd.n589 gnd.n393 240.244
R13756 gnd.n7140 gnd.n393 240.244
R13757 gnd.n7140 gnd.n388 240.244
R13758 gnd.n7157 gnd.n388 240.244
R13759 gnd.n7157 gnd.n389 240.244
R13760 gnd.n7153 gnd.n389 240.244
R13761 gnd.n7153 gnd.n7152 240.244
R13762 gnd.n7152 gnd.n348 240.244
R13763 gnd.n7213 gnd.n348 240.244
R13764 gnd.n7214 gnd.n7213 240.244
R13765 gnd.n7214 gnd.n343 240.244
R13766 gnd.n3144 gnd.n2188 240.244
R13767 gnd.n3144 gnd.n2184 240.244
R13768 gnd.n3150 gnd.n2184 240.244
R13769 gnd.n3150 gnd.n2182 240.244
R13770 gnd.n3154 gnd.n2182 240.244
R13771 gnd.n3154 gnd.n2178 240.244
R13772 gnd.n3160 gnd.n2178 240.244
R13773 gnd.n3160 gnd.n2176 240.244
R13774 gnd.n3164 gnd.n2176 240.244
R13775 gnd.n3164 gnd.n2172 240.244
R13776 gnd.n3170 gnd.n2172 240.244
R13777 gnd.n3170 gnd.n2170 240.244
R13778 gnd.n3174 gnd.n2170 240.244
R13779 gnd.n3174 gnd.n2166 240.244
R13780 gnd.n3180 gnd.n2166 240.244
R13781 gnd.n3180 gnd.n2164 240.244
R13782 gnd.n3184 gnd.n2164 240.244
R13783 gnd.n3184 gnd.n2160 240.244
R13784 gnd.n3190 gnd.n2160 240.244
R13785 gnd.n3190 gnd.n2158 240.244
R13786 gnd.n3194 gnd.n2158 240.244
R13787 gnd.n3194 gnd.n2154 240.244
R13788 gnd.n3200 gnd.n2154 240.244
R13789 gnd.n3200 gnd.n2152 240.244
R13790 gnd.n3204 gnd.n2152 240.244
R13791 gnd.n3204 gnd.n2148 240.244
R13792 gnd.n3210 gnd.n2148 240.244
R13793 gnd.n3210 gnd.n2146 240.244
R13794 gnd.n3214 gnd.n2146 240.244
R13795 gnd.n3214 gnd.n2142 240.244
R13796 gnd.n3220 gnd.n2142 240.244
R13797 gnd.n3220 gnd.n2140 240.244
R13798 gnd.n3224 gnd.n2140 240.244
R13799 gnd.n3224 gnd.n2136 240.244
R13800 gnd.n3230 gnd.n2136 240.244
R13801 gnd.n3230 gnd.n2134 240.244
R13802 gnd.n3234 gnd.n2134 240.244
R13803 gnd.n3234 gnd.n2130 240.244
R13804 gnd.n3240 gnd.n2130 240.244
R13805 gnd.n3240 gnd.n2128 240.244
R13806 gnd.n3244 gnd.n2128 240.244
R13807 gnd.n3244 gnd.n2124 240.244
R13808 gnd.n3250 gnd.n2124 240.244
R13809 gnd.n3250 gnd.n2122 240.244
R13810 gnd.n3254 gnd.n2122 240.244
R13811 gnd.n3254 gnd.n2118 240.244
R13812 gnd.n3260 gnd.n2118 240.244
R13813 gnd.n3260 gnd.n2116 240.244
R13814 gnd.n3264 gnd.n2116 240.244
R13815 gnd.n3264 gnd.n2112 240.244
R13816 gnd.n3270 gnd.n2112 240.244
R13817 gnd.n3270 gnd.n2110 240.244
R13818 gnd.n3274 gnd.n2110 240.244
R13819 gnd.n3274 gnd.n2106 240.244
R13820 gnd.n3280 gnd.n2106 240.244
R13821 gnd.n3280 gnd.n2104 240.244
R13822 gnd.n3284 gnd.n2104 240.244
R13823 gnd.n3284 gnd.n2100 240.244
R13824 gnd.n3290 gnd.n2100 240.244
R13825 gnd.n3290 gnd.n2098 240.244
R13826 gnd.n3294 gnd.n2098 240.244
R13827 gnd.n3294 gnd.n2094 240.244
R13828 gnd.n3300 gnd.n2094 240.244
R13829 gnd.n3300 gnd.n2092 240.244
R13830 gnd.n3304 gnd.n2092 240.244
R13831 gnd.n3304 gnd.n2088 240.244
R13832 gnd.n3310 gnd.n2088 240.244
R13833 gnd.n3310 gnd.n2086 240.244
R13834 gnd.n3314 gnd.n2086 240.244
R13835 gnd.n3314 gnd.n2082 240.244
R13836 gnd.n3320 gnd.n2082 240.244
R13837 gnd.n3320 gnd.n2080 240.244
R13838 gnd.n3324 gnd.n2080 240.244
R13839 gnd.n3324 gnd.n2076 240.244
R13840 gnd.n3330 gnd.n2076 240.244
R13841 gnd.n3330 gnd.n2074 240.244
R13842 gnd.n3334 gnd.n2074 240.244
R13843 gnd.n3334 gnd.n2070 240.244
R13844 gnd.n3340 gnd.n2070 240.244
R13845 gnd.n3340 gnd.n2068 240.244
R13846 gnd.n3344 gnd.n2068 240.244
R13847 gnd.n3344 gnd.n2063 240.244
R13848 gnd.n3353 gnd.n2063 240.244
R13849 gnd.n3353 gnd.n2064 240.244
R13850 gnd.n5676 gnd.n1311 240.244
R13851 gnd.n5676 gnd.n1304 240.244
R13852 gnd.n5678 gnd.n1304 240.244
R13853 gnd.n5678 gnd.n1296 240.244
R13854 gnd.n1296 gnd.n1286 240.244
R13855 gnd.n5845 gnd.n1286 240.244
R13856 gnd.n5845 gnd.n1263 240.244
R13857 gnd.n1283 gnd.n1263 240.244
R13858 gnd.n1283 gnd.n1255 240.244
R13859 gnd.n5854 gnd.n1255 240.244
R13860 gnd.n5854 gnd.n1247 240.244
R13861 gnd.n5966 gnd.n1247 240.244
R13862 gnd.n5966 gnd.n1240 240.244
R13863 gnd.n5859 gnd.n1240 240.244
R13864 gnd.n5859 gnd.n1232 240.244
R13865 gnd.n5860 gnd.n1232 240.244
R13866 gnd.n5860 gnd.n1224 240.244
R13867 gnd.n5863 gnd.n1224 240.244
R13868 gnd.n5863 gnd.n1217 240.244
R13869 gnd.n5949 gnd.n1217 240.244
R13870 gnd.n5949 gnd.n1208 240.244
R13871 gnd.n1208 gnd.n1198 240.244
R13872 gnd.n6050 gnd.n1198 240.244
R13873 gnd.n6050 gnd.n1110 240.244
R13874 gnd.n1195 gnd.n1110 240.244
R13875 gnd.n1195 gnd.n1102 240.244
R13876 gnd.n6057 gnd.n1102 240.244
R13877 gnd.n6057 gnd.n1094 240.244
R13878 gnd.n1126 gnd.n1094 240.244
R13879 gnd.n1126 gnd.n1086 240.244
R13880 gnd.n6064 gnd.n1086 240.244
R13881 gnd.n6064 gnd.n1079 240.244
R13882 gnd.n1142 gnd.n1079 240.244
R13883 gnd.n1142 gnd.n1072 240.244
R13884 gnd.n6071 gnd.n1072 240.244
R13885 gnd.n6071 gnd.n1066 240.244
R13886 gnd.n6078 gnd.n1066 240.244
R13887 gnd.n6078 gnd.n1057 240.244
R13888 gnd.n1057 gnd.n1048 240.244
R13889 gnd.n6193 gnd.n1048 240.244
R13890 gnd.n6193 gnd.n1024 240.244
R13891 gnd.n1045 gnd.n1024 240.244
R13892 gnd.n1045 gnd.n1015 240.244
R13893 gnd.n6200 gnd.n1015 240.244
R13894 gnd.n6200 gnd.n1007 240.244
R13895 gnd.n6413 gnd.n1007 240.244
R13896 gnd.n6413 gnd.n999 240.244
R13897 gnd.n6205 gnd.n999 240.244
R13898 gnd.n6205 gnd.n991 240.244
R13899 gnd.n6206 gnd.n991 240.244
R13900 gnd.n6206 gnd.n983 240.244
R13901 gnd.n6209 gnd.n983 240.244
R13902 gnd.n6209 gnd.n977 240.244
R13903 gnd.n6210 gnd.n977 240.244
R13904 gnd.n6210 gnd.n969 240.244
R13905 gnd.n6213 gnd.n969 240.244
R13906 gnd.n6213 gnd.n962 240.244
R13907 gnd.n6214 gnd.n962 240.244
R13908 gnd.n6214 gnd.n954 240.244
R13909 gnd.n6217 gnd.n954 240.244
R13910 gnd.n6217 gnd.n946 240.244
R13911 gnd.n6218 gnd.n946 240.244
R13912 gnd.n6218 gnd.n938 240.244
R13913 gnd.n6382 gnd.n938 240.244
R13914 gnd.n6382 gnd.n929 240.244
R13915 gnd.n929 gnd.n918 240.244
R13916 gnd.n6543 gnd.n918 240.244
R13917 gnd.n6543 gnd.n913 240.244
R13918 gnd.n6550 gnd.n913 240.244
R13919 gnd.n6550 gnd.n889 240.244
R13920 gnd.n889 gnd.n877 240.244
R13921 gnd.n6601 gnd.n877 240.244
R13922 gnd.n6601 gnd.n878 240.244
R13923 gnd.n878 gnd.n874 240.244
R13924 gnd.n874 gnd.n662 240.244
R13925 gnd.n6608 gnd.n662 240.244
R13926 gnd.n6608 gnd.n654 240.244
R13927 gnd.n6767 gnd.n654 240.244
R13928 gnd.n6767 gnd.n647 240.244
R13929 gnd.n6614 gnd.n647 240.244
R13930 gnd.n6614 gnd.n638 240.244
R13931 gnd.n6759 gnd.n638 240.244
R13932 gnd.n5584 gnd.n5583 240.244
R13933 gnd.n5594 gnd.n5593 240.244
R13934 gnd.n5596 gnd.n5595 240.244
R13935 gnd.n5607 gnd.n5606 240.244
R13936 gnd.n5617 gnd.n5616 240.244
R13937 gnd.n5619 gnd.n5618 240.244
R13938 gnd.n5633 gnd.n5632 240.244
R13939 gnd.n1345 gnd.n1344 240.244
R13940 gnd.n5780 gnd.n5779 240.244
R13941 gnd.n5788 gnd.n5787 240.244
R13942 gnd.n5791 gnd.n5790 240.244
R13943 gnd.n5798 gnd.n5797 240.244
R13944 gnd.n5801 gnd.n1332 240.244
R13945 gnd.n5807 gnd.n1309 240.244
R13946 gnd.n5818 gnd.n1306 240.244
R13947 gnd.n5824 gnd.n1306 240.244
R13948 gnd.n5824 gnd.n1294 240.244
R13949 gnd.n5836 gnd.n1294 240.244
R13950 gnd.n5836 gnd.n1289 240.244
R13951 gnd.n5843 gnd.n1289 240.244
R13952 gnd.n5843 gnd.n1265 240.244
R13953 gnd.n1265 gnd.n1253 240.244
R13954 gnd.n5992 gnd.n1253 240.244
R13955 gnd.n5992 gnd.n1249 240.244
R13956 gnd.n5998 gnd.n1249 240.244
R13957 gnd.n5998 gnd.n1238 240.244
R13958 gnd.n6008 gnd.n1238 240.244
R13959 gnd.n6008 gnd.n1234 240.244
R13960 gnd.n6014 gnd.n1234 240.244
R13961 gnd.n6014 gnd.n1223 240.244
R13962 gnd.n6024 gnd.n1223 240.244
R13963 gnd.n6024 gnd.n1219 240.244
R13964 gnd.n6030 gnd.n1219 240.244
R13965 gnd.n6030 gnd.n1206 240.244
R13966 gnd.n6041 gnd.n1206 240.244
R13967 gnd.n6041 gnd.n1201 240.244
R13968 gnd.n6048 gnd.n1201 240.244
R13969 gnd.n6048 gnd.n1112 240.244
R13970 gnd.n1112 gnd.n1100 240.244
R13971 gnd.n6134 gnd.n1100 240.244
R13972 gnd.n6134 gnd.n1096 240.244
R13973 gnd.n6140 gnd.n1096 240.244
R13974 gnd.n6140 gnd.n1085 240.244
R13975 gnd.n6150 gnd.n1085 240.244
R13976 gnd.n6150 gnd.n1081 240.244
R13977 gnd.n6156 gnd.n1081 240.244
R13978 gnd.n6156 gnd.n1071 240.244
R13979 gnd.n6166 gnd.n1071 240.244
R13980 gnd.n6166 gnd.n1067 240.244
R13981 gnd.n6172 gnd.n1067 240.244
R13982 gnd.n6172 gnd.n1055 240.244
R13983 gnd.n6184 gnd.n1055 240.244
R13984 gnd.n6184 gnd.n1050 240.244
R13985 gnd.n6191 gnd.n1050 240.244
R13986 gnd.n6191 gnd.n1026 240.244
R13987 gnd.n1026 gnd.n1013 240.244
R13988 gnd.n6439 gnd.n1013 240.244
R13989 gnd.n6439 gnd.n1009 240.244
R13990 gnd.n6445 gnd.n1009 240.244
R13991 gnd.n6445 gnd.n997 240.244
R13992 gnd.n6455 gnd.n997 240.244
R13993 gnd.n6455 gnd.n993 240.244
R13994 gnd.n6461 gnd.n993 240.244
R13995 gnd.n6461 gnd.n982 240.244
R13996 gnd.n6471 gnd.n982 240.244
R13997 gnd.n6471 gnd.n978 240.244
R13998 gnd.n6477 gnd.n978 240.244
R13999 gnd.n6477 gnd.n967 240.244
R14000 gnd.n6487 gnd.n967 240.244
R14001 gnd.n6487 gnd.n963 240.244
R14002 gnd.n6493 gnd.n963 240.244
R14003 gnd.n6493 gnd.n952 240.244
R14004 gnd.n6503 gnd.n952 240.244
R14005 gnd.n6503 gnd.n948 240.244
R14006 gnd.n6509 gnd.n948 240.244
R14007 gnd.n6509 gnd.n936 240.244
R14008 gnd.n6518 gnd.n936 240.244
R14009 gnd.n6518 gnd.n930 240.244
R14010 gnd.n6531 gnd.n930 240.244
R14011 gnd.n6531 gnd.n931 240.244
R14012 gnd.n931 gnd.n921 240.244
R14013 gnd.n6524 gnd.n921 240.244
R14014 gnd.n6524 gnd.n891 240.244
R14015 gnd.n6589 gnd.n891 240.244
R14016 gnd.n6589 gnd.n892 240.244
R14017 gnd.n892 gnd.n881 240.244
R14018 gnd.n897 gnd.n881 240.244
R14019 gnd.n6578 gnd.n897 240.244
R14020 gnd.n6578 gnd.n663 240.244
R14021 gnd.n663 gnd.n653 240.244
R14022 gnd.n6790 gnd.n653 240.244
R14023 gnd.n6790 gnd.n649 240.244
R14024 gnd.n6797 gnd.n649 240.244
R14025 gnd.n6797 gnd.n637 240.244
R14026 gnd.n6809 gnd.n637 240.244
R14027 gnd.n6809 gnd.n632 240.244
R14028 gnd.n6631 gnd.n6630 240.244
R14029 gnd.n6633 gnd.n6632 240.244
R14030 gnd.n6641 gnd.n6640 240.244
R14031 gnd.n6651 gnd.n6650 240.244
R14032 gnd.n6653 gnd.n6652 240.244
R14033 gnd.n6661 gnd.n6660 240.244
R14034 gnd.n6671 gnd.n6670 240.244
R14035 gnd.n6673 gnd.n6672 240.244
R14036 gnd.n6678 gnd.n6677 240.244
R14037 gnd.n6680 gnd.n6679 240.244
R14038 gnd.n6684 gnd.n6683 240.244
R14039 gnd.n6686 gnd.n6685 240.244
R14040 gnd.n6693 gnd.n6692 240.244
R14041 gnd.n6815 gnd.n631 240.244
R14042 gnd.n1420 gnd.n1419 240.132
R14043 gnd.n720 gnd.n719 240.132
R14044 gnd.n3141 gnd.n2189 225.874
R14045 gnd.n3133 gnd.n2189 225.874
R14046 gnd.n3133 gnd.n3132 225.874
R14047 gnd.n3132 gnd.n3131 225.874
R14048 gnd.n3131 gnd.n2195 225.874
R14049 gnd.n3125 gnd.n2195 225.874
R14050 gnd.n3125 gnd.n3124 225.874
R14051 gnd.n3124 gnd.n3123 225.874
R14052 gnd.n3123 gnd.n2202 225.874
R14053 gnd.n3117 gnd.n2202 225.874
R14054 gnd.n3117 gnd.n3116 225.874
R14055 gnd.n3116 gnd.n3115 225.874
R14056 gnd.n3115 gnd.n2210 225.874
R14057 gnd.n3109 gnd.n2210 225.874
R14058 gnd.n3109 gnd.n3108 225.874
R14059 gnd.n3108 gnd.n3107 225.874
R14060 gnd.n3107 gnd.n2218 225.874
R14061 gnd.n3101 gnd.n2218 225.874
R14062 gnd.n3101 gnd.n3100 225.874
R14063 gnd.n3100 gnd.n3099 225.874
R14064 gnd.n3099 gnd.n2226 225.874
R14065 gnd.n3093 gnd.n2226 225.874
R14066 gnd.n3093 gnd.n3092 225.874
R14067 gnd.n3092 gnd.n3091 225.874
R14068 gnd.n3091 gnd.n2234 225.874
R14069 gnd.n3085 gnd.n2234 225.874
R14070 gnd.n3085 gnd.n3084 225.874
R14071 gnd.n3084 gnd.n3083 225.874
R14072 gnd.n3083 gnd.n2242 225.874
R14073 gnd.n3077 gnd.n2242 225.874
R14074 gnd.n3077 gnd.n3076 225.874
R14075 gnd.n3076 gnd.n3075 225.874
R14076 gnd.n3075 gnd.n2250 225.874
R14077 gnd.n3069 gnd.n2250 225.874
R14078 gnd.n3069 gnd.n3068 225.874
R14079 gnd.n3068 gnd.n3067 225.874
R14080 gnd.n3067 gnd.n2258 225.874
R14081 gnd.n3061 gnd.n2258 225.874
R14082 gnd.n3061 gnd.n3060 225.874
R14083 gnd.n3060 gnd.n3059 225.874
R14084 gnd.n3059 gnd.n2266 225.874
R14085 gnd.n3053 gnd.n2266 225.874
R14086 gnd.n3053 gnd.n3052 225.874
R14087 gnd.n3052 gnd.n3051 225.874
R14088 gnd.n3051 gnd.n2274 225.874
R14089 gnd.n3045 gnd.n2274 225.874
R14090 gnd.n3045 gnd.n3044 225.874
R14091 gnd.n3044 gnd.n3043 225.874
R14092 gnd.n3043 gnd.n2282 225.874
R14093 gnd.n3037 gnd.n2282 225.874
R14094 gnd.n3037 gnd.n3036 225.874
R14095 gnd.n3036 gnd.n3035 225.874
R14096 gnd.n3035 gnd.n2290 225.874
R14097 gnd.n3029 gnd.n2290 225.874
R14098 gnd.n3029 gnd.n3028 225.874
R14099 gnd.n3028 gnd.n3027 225.874
R14100 gnd.n3027 gnd.n2298 225.874
R14101 gnd.n3021 gnd.n2298 225.874
R14102 gnd.n3021 gnd.n3020 225.874
R14103 gnd.n3020 gnd.n3019 225.874
R14104 gnd.n3019 gnd.n2306 225.874
R14105 gnd.n3013 gnd.n2306 225.874
R14106 gnd.n3013 gnd.n3012 225.874
R14107 gnd.n3012 gnd.n3011 225.874
R14108 gnd.n3011 gnd.n2314 225.874
R14109 gnd.n3005 gnd.n2314 225.874
R14110 gnd.n3005 gnd.n3004 225.874
R14111 gnd.n3004 gnd.n3003 225.874
R14112 gnd.n3003 gnd.n2322 225.874
R14113 gnd.n2997 gnd.n2322 225.874
R14114 gnd.n2997 gnd.n2996 225.874
R14115 gnd.n2996 gnd.n2995 225.874
R14116 gnd.n2995 gnd.n2330 225.874
R14117 gnd.n2989 gnd.n2330 225.874
R14118 gnd.n2989 gnd.n2988 225.874
R14119 gnd.n2988 gnd.n2987 225.874
R14120 gnd.n2987 gnd.n2338 225.874
R14121 gnd.n2981 gnd.n2338 225.874
R14122 gnd.n2981 gnd.n2980 225.874
R14123 gnd.n2980 gnd.n2979 225.874
R14124 gnd.n2979 gnd.n2346 225.874
R14125 gnd.n2973 gnd.n2346 225.874
R14126 gnd.n2973 gnd.n2972 225.874
R14127 gnd.n2972 gnd.n2971 225.874
R14128 gnd.n2971 gnd.n2354 225.874
R14129 gnd.n2965 gnd.n2354 225.874
R14130 gnd.n2965 gnd.n2964 225.874
R14131 gnd.n2964 gnd.n2963 225.874
R14132 gnd.n2963 gnd.n2362 225.874
R14133 gnd.n2957 gnd.n2362 225.874
R14134 gnd.n2957 gnd.n2956 225.874
R14135 gnd.n2956 gnd.n2955 225.874
R14136 gnd.n2955 gnd.n2370 225.874
R14137 gnd.n2949 gnd.n2370 225.874
R14138 gnd.n2949 gnd.n2948 225.874
R14139 gnd.n2948 gnd.n2947 225.874
R14140 gnd.n2947 gnd.n2378 225.874
R14141 gnd.n2941 gnd.n2378 225.874
R14142 gnd.n2941 gnd.n2940 225.874
R14143 gnd.n2940 gnd.n2939 225.874
R14144 gnd.n2939 gnd.n2386 225.874
R14145 gnd.n2933 gnd.n2386 225.874
R14146 gnd.n2933 gnd.n2932 225.874
R14147 gnd.n2932 gnd.n2931 225.874
R14148 gnd.n2931 gnd.n2394 225.874
R14149 gnd.n2925 gnd.n2394 225.874
R14150 gnd.n2925 gnd.n2924 225.874
R14151 gnd.n2924 gnd.n2923 225.874
R14152 gnd.n2923 gnd.n2402 225.874
R14153 gnd.n2917 gnd.n2402 225.874
R14154 gnd.n2917 gnd.n2916 225.874
R14155 gnd.n2916 gnd.n2915 225.874
R14156 gnd.n2915 gnd.n2410 225.874
R14157 gnd.n2909 gnd.n2410 225.874
R14158 gnd.n2909 gnd.n2908 225.874
R14159 gnd.n2908 gnd.n2907 225.874
R14160 gnd.n2907 gnd.n2418 225.874
R14161 gnd.n2901 gnd.n2418 225.874
R14162 gnd.n2901 gnd.n2900 225.874
R14163 gnd.n2900 gnd.n2899 225.874
R14164 gnd.n2899 gnd.n2426 225.874
R14165 gnd.n2893 gnd.n2426 225.874
R14166 gnd.n2893 gnd.n2892 225.874
R14167 gnd.n2892 gnd.n2891 225.874
R14168 gnd.n2891 gnd.n2434 225.874
R14169 gnd.n2885 gnd.n2434 225.874
R14170 gnd.n2885 gnd.n2884 225.874
R14171 gnd.n2884 gnd.n2883 225.874
R14172 gnd.n2883 gnd.n2442 225.874
R14173 gnd.n2877 gnd.n2442 225.874
R14174 gnd.n2877 gnd.n2876 225.874
R14175 gnd.n2876 gnd.n2875 225.874
R14176 gnd.n2875 gnd.n2450 225.874
R14177 gnd.n2869 gnd.n2450 225.874
R14178 gnd.n2869 gnd.n2868 225.874
R14179 gnd.n2868 gnd.n2867 225.874
R14180 gnd.n2867 gnd.n2458 225.874
R14181 gnd.n2861 gnd.n2458 225.874
R14182 gnd.n2861 gnd.n2860 225.874
R14183 gnd.n2860 gnd.n2859 225.874
R14184 gnd.n2859 gnd.n2466 225.874
R14185 gnd.n2853 gnd.n2466 225.874
R14186 gnd.n2853 gnd.n2852 225.874
R14187 gnd.n2852 gnd.n2851 225.874
R14188 gnd.n2851 gnd.n2474 225.874
R14189 gnd.n2845 gnd.n2474 225.874
R14190 gnd.n2845 gnd.n2844 225.874
R14191 gnd.n2844 gnd.n2843 225.874
R14192 gnd.n2843 gnd.n2482 225.874
R14193 gnd.n2837 gnd.n2482 225.874
R14194 gnd.n2837 gnd.n2836 225.874
R14195 gnd.n2836 gnd.n2835 225.874
R14196 gnd.n2835 gnd.n2490 225.874
R14197 gnd.n2829 gnd.n2490 225.874
R14198 gnd.n3912 gnd.t90 224.174
R14199 gnd.n2053 gnd.t38 224.174
R14200 gnd.n535 gnd.n496 199.319
R14201 gnd.n535 gnd.n497 199.319
R14202 gnd.n5739 gnd.n5738 199.319
R14203 gnd.n5738 gnd.n5737 199.319
R14204 gnd.n1421 gnd.n1418 186.49
R14205 gnd.n721 gnd.n718 186.49
R14206 gnd.n4626 gnd.n4625 185
R14207 gnd.n4624 gnd.n4623 185
R14208 gnd.n4603 gnd.n4602 185
R14209 gnd.n4618 gnd.n4617 185
R14210 gnd.n4616 gnd.n4615 185
R14211 gnd.n4607 gnd.n4606 185
R14212 gnd.n4610 gnd.n4609 185
R14213 gnd.n4594 gnd.n4593 185
R14214 gnd.n4592 gnd.n4591 185
R14215 gnd.n4571 gnd.n4570 185
R14216 gnd.n4586 gnd.n4585 185
R14217 gnd.n4584 gnd.n4583 185
R14218 gnd.n4575 gnd.n4574 185
R14219 gnd.n4578 gnd.n4577 185
R14220 gnd.n4562 gnd.n4561 185
R14221 gnd.n4560 gnd.n4559 185
R14222 gnd.n4539 gnd.n4538 185
R14223 gnd.n4554 gnd.n4553 185
R14224 gnd.n4552 gnd.n4551 185
R14225 gnd.n4543 gnd.n4542 185
R14226 gnd.n4546 gnd.n4545 185
R14227 gnd.n4531 gnd.n4530 185
R14228 gnd.n4529 gnd.n4528 185
R14229 gnd.n4508 gnd.n4507 185
R14230 gnd.n4523 gnd.n4522 185
R14231 gnd.n4521 gnd.n4520 185
R14232 gnd.n4512 gnd.n4511 185
R14233 gnd.n4515 gnd.n4514 185
R14234 gnd.n4499 gnd.n4498 185
R14235 gnd.n4497 gnd.n4496 185
R14236 gnd.n4476 gnd.n4475 185
R14237 gnd.n4491 gnd.n4490 185
R14238 gnd.n4489 gnd.n4488 185
R14239 gnd.n4480 gnd.n4479 185
R14240 gnd.n4483 gnd.n4482 185
R14241 gnd.n4467 gnd.n4466 185
R14242 gnd.n4465 gnd.n4464 185
R14243 gnd.n4444 gnd.n4443 185
R14244 gnd.n4459 gnd.n4458 185
R14245 gnd.n4457 gnd.n4456 185
R14246 gnd.n4448 gnd.n4447 185
R14247 gnd.n4451 gnd.n4450 185
R14248 gnd.n4435 gnd.n4434 185
R14249 gnd.n4433 gnd.n4432 185
R14250 gnd.n4412 gnd.n4411 185
R14251 gnd.n4427 gnd.n4426 185
R14252 gnd.n4425 gnd.n4424 185
R14253 gnd.n4416 gnd.n4415 185
R14254 gnd.n4419 gnd.n4418 185
R14255 gnd.n4404 gnd.n4403 185
R14256 gnd.n4402 gnd.n4401 185
R14257 gnd.n4381 gnd.n4380 185
R14258 gnd.n4396 gnd.n4395 185
R14259 gnd.n4394 gnd.n4393 185
R14260 gnd.n4385 gnd.n4384 185
R14261 gnd.n4388 gnd.n4387 185
R14262 gnd.n3913 gnd.t89 178.987
R14263 gnd.n2054 gnd.t39 178.987
R14264 gnd.n1 gnd.t176 170.774
R14265 gnd.n7 gnd.t3 170.103
R14266 gnd.n6 gnd.t171 170.103
R14267 gnd.n5 gnd.t122 170.103
R14268 gnd.n4 gnd.t185 170.103
R14269 gnd.n3 gnd.t6 170.103
R14270 gnd.n2 gnd.t162 170.103
R14271 gnd.n1 gnd.t191 170.103
R14272 gnd.n734 gnd.n732 163.367
R14273 gnd.n738 gnd.n707 163.367
R14274 gnd.n742 gnd.n740 163.367
R14275 gnd.n746 gnd.n705 163.367
R14276 gnd.n750 gnd.n748 163.367
R14277 gnd.n754 gnd.n703 163.367
R14278 gnd.n758 gnd.n756 163.367
R14279 gnd.n762 gnd.n701 163.367
R14280 gnd.n766 gnd.n764 163.367
R14281 gnd.n770 gnd.n699 163.367
R14282 gnd.n774 gnd.n772 163.367
R14283 gnd.n778 gnd.n697 163.367
R14284 gnd.n782 gnd.n780 163.367
R14285 gnd.n789 gnd.n695 163.367
R14286 gnd.n792 gnd.n791 163.367
R14287 gnd.n796 gnd.n795 163.367
R14288 gnd.n801 gnd.n799 163.367
R14289 gnd.n808 gnd.n692 163.367
R14290 gnd.n812 gnd.n810 163.367
R14291 gnd.n816 gnd.n690 163.367
R14292 gnd.n820 gnd.n818 163.367
R14293 gnd.n824 gnd.n688 163.367
R14294 gnd.n828 gnd.n826 163.367
R14295 gnd.n832 gnd.n686 163.367
R14296 gnd.n836 gnd.n834 163.367
R14297 gnd.n840 gnd.n684 163.367
R14298 gnd.n844 gnd.n842 163.367
R14299 gnd.n848 gnd.n682 163.367
R14300 gnd.n852 gnd.n850 163.367
R14301 gnd.n856 gnd.n680 163.367
R14302 gnd.n859 gnd.n858 163.367
R14303 gnd.n863 gnd.n862 163.367
R14304 gnd.n1537 gnd.n1536 163.367
R14305 gnd.n1536 gnd.n1531 163.367
R14306 gnd.n1532 gnd.n1531 163.367
R14307 gnd.n1532 gnd.n1266 163.367
R14308 gnd.n5982 gnd.n1266 163.367
R14309 gnd.n5982 gnd.n1267 163.367
R14310 gnd.n5978 gnd.n1267 163.367
R14311 gnd.n5978 gnd.n5977 163.367
R14312 gnd.n5977 gnd.n5976 163.367
R14313 gnd.n5976 gnd.n1270 163.367
R14314 gnd.n5894 gnd.n1270 163.367
R14315 gnd.n5894 gnd.n1277 163.367
R14316 gnd.n5897 gnd.n1277 163.367
R14317 gnd.n5897 gnd.n5892 163.367
R14318 gnd.n5912 gnd.n5892 163.367
R14319 gnd.n5913 gnd.n5912 163.367
R14320 gnd.n5914 gnd.n5913 163.367
R14321 gnd.n5914 gnd.n5890 163.367
R14322 gnd.n5919 gnd.n5890 163.367
R14323 gnd.n5919 gnd.n5881 163.367
R14324 gnd.n5928 gnd.n5881 163.367
R14325 gnd.n5929 gnd.n5928 163.367
R14326 gnd.n5930 gnd.n5929 163.367
R14327 gnd.n5930 gnd.n5864 163.367
R14328 gnd.n5933 gnd.n5864 163.367
R14329 gnd.n5933 gnd.n5878 163.367
R14330 gnd.n5938 gnd.n5878 163.367
R14331 gnd.n5938 gnd.n5879 163.367
R14332 gnd.n5879 gnd.n1113 163.367
R14333 gnd.n6124 gnd.n1113 163.367
R14334 gnd.n6124 gnd.n1114 163.367
R14335 gnd.n6120 gnd.n1114 163.367
R14336 gnd.n6120 gnd.n6119 163.367
R14337 gnd.n6119 gnd.n6118 163.367
R14338 gnd.n6118 gnd.n1117 163.367
R14339 gnd.n1129 gnd.n1117 163.367
R14340 gnd.n1129 gnd.n1125 163.367
R14341 gnd.n6107 gnd.n1125 163.367
R14342 gnd.n6107 gnd.n1127 163.367
R14343 gnd.n6103 gnd.n1127 163.367
R14344 gnd.n6103 gnd.n1133 163.367
R14345 gnd.n1144 gnd.n1133 163.367
R14346 gnd.n1144 gnd.n1141 163.367
R14347 gnd.n6092 gnd.n1141 163.367
R14348 gnd.n6092 gnd.n1143 163.367
R14349 gnd.n6088 gnd.n1143 163.367
R14350 gnd.n6088 gnd.n1148 163.367
R14351 gnd.n1157 gnd.n1148 163.367
R14352 gnd.n1185 gnd.n1157 163.367
R14353 gnd.n1185 gnd.n1158 163.367
R14354 gnd.n1181 gnd.n1158 163.367
R14355 gnd.n1181 gnd.n1180 163.367
R14356 gnd.n1180 gnd.n1162 163.367
R14357 gnd.n1162 gnd.n1027 163.367
R14358 gnd.n6429 gnd.n1027 163.367
R14359 gnd.n6429 gnd.n1028 163.367
R14360 gnd.n6425 gnd.n1028 163.367
R14361 gnd.n6425 gnd.n6424 163.367
R14362 gnd.n6424 gnd.n6423 163.367
R14363 gnd.n6423 gnd.n1031 163.367
R14364 gnd.n6277 gnd.n1031 163.367
R14365 gnd.n6277 gnd.n1039 163.367
R14366 gnd.n6280 gnd.n1039 163.367
R14367 gnd.n6280 gnd.n6274 163.367
R14368 gnd.n6287 gnd.n6274 163.367
R14369 gnd.n6287 gnd.n6275 163.367
R14370 gnd.n6283 gnd.n6275 163.367
R14371 gnd.n6283 gnd.n6265 163.367
R14372 gnd.n6299 gnd.n6265 163.367
R14373 gnd.n6299 gnd.n6262 163.367
R14374 gnd.n6305 gnd.n6262 163.367
R14375 gnd.n6305 gnd.n6263 163.367
R14376 gnd.n6263 gnd.n6255 163.367
R14377 gnd.n6317 gnd.n6255 163.367
R14378 gnd.n6318 gnd.n6317 163.367
R14379 gnd.n6318 gnd.n6252 163.367
R14380 gnd.n6324 gnd.n6252 163.367
R14381 gnd.n6324 gnd.n6253 163.367
R14382 gnd.n6253 gnd.n6246 163.367
R14383 gnd.n6336 gnd.n6246 163.367
R14384 gnd.n6337 gnd.n6336 163.367
R14385 gnd.n6337 gnd.n6243 163.367
R14386 gnd.n6343 gnd.n6243 163.367
R14387 gnd.n6343 gnd.n6244 163.367
R14388 gnd.n6244 gnd.n6235 163.367
R14389 gnd.n6353 gnd.n6235 163.367
R14390 gnd.n6354 gnd.n6353 163.367
R14391 gnd.n6355 gnd.n6354 163.367
R14392 gnd.n6355 gnd.n6221 163.367
R14393 gnd.n6358 gnd.n6221 163.367
R14394 gnd.n6358 gnd.n6232 163.367
R14395 gnd.n6371 gnd.n6232 163.367
R14396 gnd.n6371 gnd.n6233 163.367
R14397 gnd.n6367 gnd.n6233 163.367
R14398 gnd.n6367 gnd.n6366 163.367
R14399 gnd.n6366 gnd.n912 163.367
R14400 gnd.n6362 gnd.n912 163.367
R14401 gnd.n6362 gnd.n905 163.367
R14402 gnd.n6561 gnd.n905 163.367
R14403 gnd.n6562 gnd.n6561 163.367
R14404 gnd.n6562 gnd.n902 163.367
R14405 gnd.n6567 gnd.n902 163.367
R14406 gnd.n6567 gnd.n903 163.367
R14407 gnd.n903 gnd.n664 163.367
R14408 gnd.n6780 gnd.n664 163.367
R14409 gnd.n6780 gnd.n665 163.367
R14410 gnd.n6776 gnd.n665 163.367
R14411 gnd.n6776 gnd.n668 163.367
R14412 gnd.n869 gnd.n668 163.367
R14413 gnd.n869 gnd.n676 163.367
R14414 gnd.n1513 gnd.n1512 163.367
R14415 gnd.n1512 gnd.n1511 163.367
R14416 gnd.n1508 gnd.n1507 163.367
R14417 gnd.n1505 gnd.n1439 163.367
R14418 gnd.n1501 gnd.n1499 163.367
R14419 gnd.n1497 gnd.n1441 163.367
R14420 gnd.n1493 gnd.n1491 163.367
R14421 gnd.n1489 gnd.n1443 163.367
R14422 gnd.n1485 gnd.n1483 163.367
R14423 gnd.n1481 gnd.n1445 163.367
R14424 gnd.n1477 gnd.n1475 163.367
R14425 gnd.n1473 gnd.n1447 163.367
R14426 gnd.n1469 gnd.n1467 163.367
R14427 gnd.n1465 gnd.n1449 163.367
R14428 gnd.n1461 gnd.n1459 163.367
R14429 gnd.n1456 gnd.n1455 163.367
R14430 gnd.n1604 gnd.n1602 163.367
R14431 gnd.n1600 gnd.n1393 163.367
R14432 gnd.n1595 gnd.n1593 163.367
R14433 gnd.n1591 gnd.n1397 163.367
R14434 gnd.n1587 gnd.n1585 163.367
R14435 gnd.n1583 gnd.n1399 163.367
R14436 gnd.n1579 gnd.n1577 163.367
R14437 gnd.n1575 gnd.n1401 163.367
R14438 gnd.n1571 gnd.n1569 163.367
R14439 gnd.n1567 gnd.n1403 163.367
R14440 gnd.n1563 gnd.n1561 163.367
R14441 gnd.n1559 gnd.n1405 163.367
R14442 gnd.n1555 gnd.n1553 163.367
R14443 gnd.n1551 gnd.n1407 163.367
R14444 gnd.n1547 gnd.n1545 163.367
R14445 gnd.n1543 gnd.n1409 163.367
R14446 gnd.n1517 gnd.n1412 163.367
R14447 gnd.n1529 gnd.n1412 163.367
R14448 gnd.n1529 gnd.n1413 163.367
R14449 gnd.n1525 gnd.n1413 163.367
R14450 gnd.n1525 gnd.n1262 163.367
R14451 gnd.n1522 gnd.n1262 163.367
R14452 gnd.n1522 gnd.n1521 163.367
R14453 gnd.n1521 gnd.n1272 163.367
R14454 gnd.n5974 gnd.n1272 163.367
R14455 gnd.n5974 gnd.n1273 163.367
R14456 gnd.n5970 gnd.n1273 163.367
R14457 gnd.n5970 gnd.n5969 163.367
R14458 gnd.n5969 gnd.n1276 163.367
R14459 gnd.n5902 gnd.n1276 163.367
R14460 gnd.n5910 gnd.n5902 163.367
R14461 gnd.n5910 gnd.n5903 163.367
R14462 gnd.n5906 gnd.n5903 163.367
R14463 gnd.n5906 gnd.n5887 163.367
R14464 gnd.n5921 gnd.n5887 163.367
R14465 gnd.n5921 gnd.n5884 163.367
R14466 gnd.n5926 gnd.n5884 163.367
R14467 gnd.n5926 gnd.n5885 163.367
R14468 gnd.n5885 gnd.n5865 163.367
R14469 gnd.n5946 gnd.n5865 163.367
R14470 gnd.n5946 gnd.n5866 163.367
R14471 gnd.n5942 gnd.n5866 163.367
R14472 gnd.n5942 gnd.n5941 163.367
R14473 gnd.n5941 gnd.n5877 163.367
R14474 gnd.n5877 gnd.n5869 163.367
R14475 gnd.n5869 gnd.n1109 163.367
R14476 gnd.n5872 gnd.n1109 163.367
R14477 gnd.n5872 gnd.n5871 163.367
R14478 gnd.n5871 gnd.n1120 163.367
R14479 gnd.n6116 gnd.n1120 163.367
R14480 gnd.n6116 gnd.n1121 163.367
R14481 gnd.n6112 gnd.n1121 163.367
R14482 gnd.n6112 gnd.n6111 163.367
R14483 gnd.n6111 gnd.n1124 163.367
R14484 gnd.n1135 gnd.n1124 163.367
R14485 gnd.n6101 gnd.n1135 163.367
R14486 gnd.n6101 gnd.n1136 163.367
R14487 gnd.n6097 gnd.n1136 163.367
R14488 gnd.n6097 gnd.n6096 163.367
R14489 gnd.n6096 gnd.n1140 163.367
R14490 gnd.n1151 gnd.n1140 163.367
R14491 gnd.n6086 gnd.n1151 163.367
R14492 gnd.n6086 gnd.n1152 163.367
R14493 gnd.n6082 gnd.n1152 163.367
R14494 gnd.n6082 gnd.n1156 163.367
R14495 gnd.n1166 gnd.n1156 163.367
R14496 gnd.n1166 gnd.n1164 163.367
R14497 gnd.n1178 gnd.n1164 163.367
R14498 gnd.n1178 gnd.n1165 163.367
R14499 gnd.n1174 gnd.n1165 163.367
R14500 gnd.n1174 gnd.n1023 163.367
R14501 gnd.n1171 gnd.n1023 163.367
R14502 gnd.n1171 gnd.n1170 163.367
R14503 gnd.n1170 gnd.n1034 163.367
R14504 gnd.n6421 gnd.n1034 163.367
R14505 gnd.n6421 gnd.n1035 163.367
R14506 gnd.n6417 gnd.n1035 163.367
R14507 gnd.n6417 gnd.n6416 163.367
R14508 gnd.n6416 gnd.n1038 163.367
R14509 gnd.n6270 gnd.n1038 163.367
R14510 gnd.n6290 gnd.n6270 163.367
R14511 gnd.n6291 gnd.n6290 163.367
R14512 gnd.n6292 gnd.n6291 163.367
R14513 gnd.n6292 gnd.n6268 163.367
R14514 gnd.n6297 gnd.n6268 163.367
R14515 gnd.n6297 gnd.n6261 163.367
R14516 gnd.n6308 gnd.n6261 163.367
R14517 gnd.n6309 gnd.n6308 163.367
R14518 gnd.n6309 gnd.n6258 163.367
R14519 gnd.n6315 gnd.n6258 163.367
R14520 gnd.n6315 gnd.n6259 163.367
R14521 gnd.n6259 gnd.n6251 163.367
R14522 gnd.n6327 gnd.n6251 163.367
R14523 gnd.n6328 gnd.n6327 163.367
R14524 gnd.n6328 gnd.n6248 163.367
R14525 gnd.n6334 gnd.n6248 163.367
R14526 gnd.n6334 gnd.n6249 163.367
R14527 gnd.n6249 gnd.n6241 163.367
R14528 gnd.n6345 gnd.n6241 163.367
R14529 gnd.n6346 gnd.n6345 163.367
R14530 gnd.n6346 gnd.n6238 163.367
R14531 gnd.n6351 gnd.n6238 163.367
R14532 gnd.n6351 gnd.n6239 163.367
R14533 gnd.n6239 gnd.n6222 163.367
R14534 gnd.n6379 gnd.n6222 163.367
R14535 gnd.n6379 gnd.n6223 163.367
R14536 gnd.n6375 gnd.n6223 163.367
R14537 gnd.n6375 gnd.n6231 163.367
R14538 gnd.n6231 gnd.n6230 163.367
R14539 gnd.n6230 gnd.n6226 163.367
R14540 gnd.n6226 gnd.n910 163.367
R14541 gnd.n6553 gnd.n910 163.367
R14542 gnd.n6554 gnd.n6553 163.367
R14543 gnd.n6554 gnd.n907 163.367
R14544 gnd.n6559 gnd.n907 163.367
R14545 gnd.n6559 gnd.n908 163.367
R14546 gnd.n908 gnd.n901 163.367
R14547 gnd.n6570 gnd.n901 163.367
R14548 gnd.n6570 gnd.n899 163.367
R14549 gnd.n6575 gnd.n899 163.367
R14550 gnd.n6575 gnd.n661 163.367
R14551 gnd.n671 gnd.n661 163.367
R14552 gnd.n6774 gnd.n671 163.367
R14553 gnd.n6774 gnd.n672 163.367
R14554 gnd.n6770 gnd.n672 163.367
R14555 gnd.n6770 gnd.n675 163.367
R14556 gnd.n727 gnd.n726 156.462
R14557 gnd.n4566 gnd.n4534 153.042
R14558 gnd.n4630 gnd.n4629 152.079
R14559 gnd.n4598 gnd.n4597 152.079
R14560 gnd.n4566 gnd.n4565 152.079
R14561 gnd.n1426 gnd.n1425 152
R14562 gnd.n1427 gnd.n1416 152
R14563 gnd.n1429 gnd.n1428 152
R14564 gnd.n1431 gnd.n1414 152
R14565 gnd.n1433 gnd.n1432 152
R14566 gnd.n725 gnd.n709 152
R14567 gnd.n717 gnd.n710 152
R14568 gnd.n716 gnd.n715 152
R14569 gnd.n714 gnd.n711 152
R14570 gnd.n712 gnd.t104 150.546
R14571 gnd.t129 gnd.n4608 147.661
R14572 gnd.t135 gnd.n4576 147.661
R14573 gnd.t189 gnd.n4544 147.661
R14574 gnd.t132 gnd.n4513 147.661
R14575 gnd.t160 gnd.n4481 147.661
R14576 gnd.t353 gnd.n4449 147.661
R14577 gnd.t10 gnd.n4417 147.661
R14578 gnd.t158 gnd.n4386 147.661
R14579 gnd.n798 gnd.n797 143.351
R14580 gnd.n1454 gnd.n1392 143.351
R14581 gnd.n1603 gnd.n1392 143.351
R14582 gnd.n1423 gnd.t14 130.484
R14583 gnd.n1432 gnd.t98 126.766
R14584 gnd.n1430 gnd.t17 126.766
R14585 gnd.n1416 gnd.t51 126.766
R14586 gnd.n1424 gnd.t113 126.766
R14587 gnd.n713 gnd.t84 126.766
R14588 gnd.n715 gnd.t11 126.766
R14589 gnd.n724 gnd.t71 126.766
R14590 gnd.n726 gnd.t40 126.766
R14591 gnd.n4625 gnd.n4624 104.615
R14592 gnd.n4624 gnd.n4602 104.615
R14593 gnd.n4617 gnd.n4602 104.615
R14594 gnd.n4617 gnd.n4616 104.615
R14595 gnd.n4616 gnd.n4606 104.615
R14596 gnd.n4609 gnd.n4606 104.615
R14597 gnd.n4593 gnd.n4592 104.615
R14598 gnd.n4592 gnd.n4570 104.615
R14599 gnd.n4585 gnd.n4570 104.615
R14600 gnd.n4585 gnd.n4584 104.615
R14601 gnd.n4584 gnd.n4574 104.615
R14602 gnd.n4577 gnd.n4574 104.615
R14603 gnd.n4561 gnd.n4560 104.615
R14604 gnd.n4560 gnd.n4538 104.615
R14605 gnd.n4553 gnd.n4538 104.615
R14606 gnd.n4553 gnd.n4552 104.615
R14607 gnd.n4552 gnd.n4542 104.615
R14608 gnd.n4545 gnd.n4542 104.615
R14609 gnd.n4530 gnd.n4529 104.615
R14610 gnd.n4529 gnd.n4507 104.615
R14611 gnd.n4522 gnd.n4507 104.615
R14612 gnd.n4522 gnd.n4521 104.615
R14613 gnd.n4521 gnd.n4511 104.615
R14614 gnd.n4514 gnd.n4511 104.615
R14615 gnd.n4498 gnd.n4497 104.615
R14616 gnd.n4497 gnd.n4475 104.615
R14617 gnd.n4490 gnd.n4475 104.615
R14618 gnd.n4490 gnd.n4489 104.615
R14619 gnd.n4489 gnd.n4479 104.615
R14620 gnd.n4482 gnd.n4479 104.615
R14621 gnd.n4466 gnd.n4465 104.615
R14622 gnd.n4465 gnd.n4443 104.615
R14623 gnd.n4458 gnd.n4443 104.615
R14624 gnd.n4458 gnd.n4457 104.615
R14625 gnd.n4457 gnd.n4447 104.615
R14626 gnd.n4450 gnd.n4447 104.615
R14627 gnd.n4434 gnd.n4433 104.615
R14628 gnd.n4433 gnd.n4411 104.615
R14629 gnd.n4426 gnd.n4411 104.615
R14630 gnd.n4426 gnd.n4425 104.615
R14631 gnd.n4425 gnd.n4415 104.615
R14632 gnd.n4418 gnd.n4415 104.615
R14633 gnd.n4403 gnd.n4402 104.615
R14634 gnd.n4402 gnd.n4380 104.615
R14635 gnd.n4395 gnd.n4380 104.615
R14636 gnd.n4395 gnd.n4394 104.615
R14637 gnd.n4394 gnd.n4384 104.615
R14638 gnd.n4387 gnd.n4384 104.615
R14639 gnd.n3838 gnd.t23 100.632
R14640 gnd.n2027 gnd.t66 100.632
R14641 gnd.n7565 gnd.n134 99.6594
R14642 gnd.n7563 gnd.n7562 99.6594
R14643 gnd.n7558 gnd.n141 99.6594
R14644 gnd.n7556 gnd.n7555 99.6594
R14645 gnd.n7551 gnd.n148 99.6594
R14646 gnd.n7549 gnd.n7548 99.6594
R14647 gnd.n7544 gnd.n155 99.6594
R14648 gnd.n7542 gnd.n7541 99.6594
R14649 gnd.n7534 gnd.n162 99.6594
R14650 gnd.n7532 gnd.n7531 99.6594
R14651 gnd.n7527 gnd.n169 99.6594
R14652 gnd.n7525 gnd.n7524 99.6594
R14653 gnd.n7520 gnd.n176 99.6594
R14654 gnd.n7518 gnd.n7517 99.6594
R14655 gnd.n7513 gnd.n183 99.6594
R14656 gnd.n7511 gnd.n7510 99.6594
R14657 gnd.n7506 gnd.n190 99.6594
R14658 gnd.n7504 gnd.n7503 99.6594
R14659 gnd.n195 gnd.n194 99.6594
R14660 gnd.n7048 gnd.n7047 99.6594
R14661 gnd.n519 gnd.n490 99.6594
R14662 gnd.n7040 gnd.n491 99.6594
R14663 gnd.n7036 gnd.n492 99.6594
R14664 gnd.n7032 gnd.n493 99.6594
R14665 gnd.n7028 gnd.n494 99.6594
R14666 gnd.n7024 gnd.n495 99.6594
R14667 gnd.n7020 gnd.n496 99.6594
R14668 gnd.n7015 gnd.n498 99.6594
R14669 gnd.n7011 gnd.n499 99.6594
R14670 gnd.n7007 gnd.n500 99.6594
R14671 gnd.n7003 gnd.n501 99.6594
R14672 gnd.n6999 gnd.n502 99.6594
R14673 gnd.n6995 gnd.n503 99.6594
R14674 gnd.n6991 gnd.n504 99.6594
R14675 gnd.n6987 gnd.n505 99.6594
R14676 gnd.n6983 gnd.n506 99.6594
R14677 gnd.n558 gnd.n507 99.6594
R14678 gnd.n5763 gnd.n5762 99.6594
R14679 gnd.n5760 gnd.n5759 99.6594
R14680 gnd.n5755 gnd.n1373 99.6594
R14681 gnd.n5753 gnd.n5752 99.6594
R14682 gnd.n5748 gnd.n1380 99.6594
R14683 gnd.n5746 gnd.n5745 99.6594
R14684 gnd.n5741 gnd.n1387 99.6594
R14685 gnd.n5737 gnd.n5736 99.6594
R14686 gnd.n5732 gnd.n1614 99.6594
R14687 gnd.n5730 gnd.n5729 99.6594
R14688 gnd.n5725 gnd.n1621 99.6594
R14689 gnd.n5723 gnd.n5722 99.6594
R14690 gnd.n5718 gnd.n1628 99.6594
R14691 gnd.n5716 gnd.n5715 99.6594
R14692 gnd.n5711 gnd.n1635 99.6594
R14693 gnd.n5709 gnd.n5708 99.6594
R14694 gnd.n5704 gnd.n1644 99.6594
R14695 gnd.n5702 gnd.n5701 99.6594
R14696 gnd.n5062 gnd.n4873 99.6594
R14697 gnd.n5060 gnd.n4876 99.6594
R14698 gnd.n5056 gnd.n5055 99.6594
R14699 gnd.n5049 gnd.n4881 99.6594
R14700 gnd.n5048 gnd.n5047 99.6594
R14701 gnd.n5041 gnd.n4887 99.6594
R14702 gnd.n5040 gnd.n5039 99.6594
R14703 gnd.n5033 gnd.n4893 99.6594
R14704 gnd.n5032 gnd.n5031 99.6594
R14705 gnd.n5025 gnd.n4899 99.6594
R14706 gnd.n5024 gnd.n5023 99.6594
R14707 gnd.n5017 gnd.n4908 99.6594
R14708 gnd.n5016 gnd.n5015 99.6594
R14709 gnd.n5009 gnd.n4914 99.6594
R14710 gnd.n5008 gnd.n5007 99.6594
R14711 gnd.n5001 gnd.n4920 99.6594
R14712 gnd.n5000 gnd.n4999 99.6594
R14713 gnd.n4930 gnd.n4926 99.6594
R14714 gnd.n4989 gnd.n4988 99.6594
R14715 gnd.n4746 gnd.n2010 99.6594
R14716 gnd.n4744 gnd.n2009 99.6594
R14717 gnd.n4740 gnd.n2008 99.6594
R14718 gnd.n4736 gnd.n2007 99.6594
R14719 gnd.n4732 gnd.n2006 99.6594
R14720 gnd.n4728 gnd.n2005 99.6594
R14721 gnd.n4724 gnd.n2004 99.6594
R14722 gnd.n3362 gnd.n2003 99.6594
R14723 gnd.n4050 gnd.n3781 99.6594
R14724 gnd.n3807 gnd.n3788 99.6594
R14725 gnd.n3809 gnd.n3789 99.6594
R14726 gnd.n3817 gnd.n3790 99.6594
R14727 gnd.n3819 gnd.n3791 99.6594
R14728 gnd.n3827 gnd.n3792 99.6594
R14729 gnd.n3829 gnd.n3793 99.6594
R14730 gnd.n3837 gnd.n3794 99.6594
R14731 gnd.n4714 gnd.n1990 99.6594
R14732 gnd.n4710 gnd.n1991 99.6594
R14733 gnd.n4706 gnd.n1992 99.6594
R14734 gnd.n4702 gnd.n1993 99.6594
R14735 gnd.n4698 gnd.n1994 99.6594
R14736 gnd.n4694 gnd.n1995 99.6594
R14737 gnd.n4690 gnd.n1996 99.6594
R14738 gnd.n4686 gnd.n1997 99.6594
R14739 gnd.n4682 gnd.n1998 99.6594
R14740 gnd.n4678 gnd.n1999 99.6594
R14741 gnd.n4674 gnd.n2000 99.6594
R14742 gnd.n4670 gnd.n2001 99.6594
R14743 gnd.n4666 gnd.n2002 99.6594
R14744 gnd.n3965 gnd.n3964 99.6594
R14745 gnd.n3959 gnd.n3876 99.6594
R14746 gnd.n3956 gnd.n3877 99.6594
R14747 gnd.n3952 gnd.n3878 99.6594
R14748 gnd.n3948 gnd.n3879 99.6594
R14749 gnd.n3944 gnd.n3880 99.6594
R14750 gnd.n3940 gnd.n3881 99.6594
R14751 gnd.n3936 gnd.n3882 99.6594
R14752 gnd.n3932 gnd.n3883 99.6594
R14753 gnd.n3928 gnd.n3884 99.6594
R14754 gnd.n3924 gnd.n3885 99.6594
R14755 gnd.n3920 gnd.n3886 99.6594
R14756 gnd.n3967 gnd.n3875 99.6594
R14757 gnd.n7420 gnd.n7419 99.6594
R14758 gnd.n7425 gnd.n7424 99.6594
R14759 gnd.n7428 gnd.n7427 99.6594
R14760 gnd.n7433 gnd.n7432 99.6594
R14761 gnd.n7436 gnd.n7435 99.6594
R14762 gnd.n7441 gnd.n7440 99.6594
R14763 gnd.n7444 gnd.n7443 99.6594
R14764 gnd.n7449 gnd.n7447 99.6594
R14765 gnd.n7575 gnd.n121 99.6594
R14766 gnd.n6621 gnd.n508 99.6594
R14767 gnd.n6625 gnd.n509 99.6594
R14768 gnd.n6627 gnd.n510 99.6594
R14769 gnd.n6637 gnd.n511 99.6594
R14770 gnd.n6645 gnd.n512 99.6594
R14771 gnd.n6647 gnd.n513 99.6594
R14772 gnd.n6657 gnd.n514 99.6594
R14773 gnd.n6665 gnd.n515 99.6594
R14774 gnd.n6667 gnd.n516 99.6594
R14775 gnd.n5578 gnd.n5577 99.6594
R14776 gnd.n5589 gnd.n5588 99.6594
R14777 gnd.n5600 gnd.n5599 99.6594
R14778 gnd.n5603 gnd.n5602 99.6594
R14779 gnd.n5612 gnd.n5611 99.6594
R14780 gnd.n5623 gnd.n5622 99.6594
R14781 gnd.n5626 gnd.n5625 99.6594
R14782 gnd.n5628 gnd.n5627 99.6594
R14783 gnd.n5773 gnd.n1351 99.6594
R14784 gnd.n4781 gnd.n1987 99.6594
R14785 gnd.n4784 gnd.n4783 99.6594
R14786 gnd.n4791 gnd.n4790 99.6594
R14787 gnd.n4794 gnd.n4793 99.6594
R14788 gnd.n4801 gnd.n4800 99.6594
R14789 gnd.n4804 gnd.n4803 99.6594
R14790 gnd.n4811 gnd.n4810 99.6594
R14791 gnd.n4814 gnd.n4813 99.6594
R14792 gnd.n4821 gnd.n4820 99.6594
R14793 gnd.n4782 gnd.n4781 99.6594
R14794 gnd.n4783 gnd.n4776 99.6594
R14795 gnd.n4792 gnd.n4791 99.6594
R14796 gnd.n4793 gnd.n4772 99.6594
R14797 gnd.n4802 gnd.n4801 99.6594
R14798 gnd.n4803 gnd.n4768 99.6594
R14799 gnd.n4812 gnd.n4811 99.6594
R14800 gnd.n4813 gnd.n4764 99.6594
R14801 gnd.n4822 gnd.n4821 99.6594
R14802 gnd.n1351 gnd.n1350 99.6594
R14803 gnd.n5629 gnd.n5628 99.6594
R14804 gnd.n5625 gnd.n5624 99.6594
R14805 gnd.n5622 gnd.n5613 99.6594
R14806 gnd.n5611 gnd.n5610 99.6594
R14807 gnd.n5602 gnd.n5601 99.6594
R14808 gnd.n5599 gnd.n5590 99.6594
R14809 gnd.n5588 gnd.n5587 99.6594
R14810 gnd.n5577 gnd.n5576 99.6594
R14811 gnd.n6624 gnd.n508 99.6594
R14812 gnd.n6626 gnd.n509 99.6594
R14813 gnd.n6636 gnd.n510 99.6594
R14814 gnd.n6644 gnd.n511 99.6594
R14815 gnd.n6646 gnd.n512 99.6594
R14816 gnd.n6656 gnd.n513 99.6594
R14817 gnd.n6664 gnd.n514 99.6594
R14818 gnd.n6666 gnd.n515 99.6594
R14819 gnd.n6711 gnd.n516 99.6594
R14820 gnd.n7448 gnd.n121 99.6594
R14821 gnd.n7447 gnd.n7446 99.6594
R14822 gnd.n7443 gnd.n7442 99.6594
R14823 gnd.n7440 gnd.n7439 99.6594
R14824 gnd.n7435 gnd.n7434 99.6594
R14825 gnd.n7432 gnd.n7431 99.6594
R14826 gnd.n7427 gnd.n7426 99.6594
R14827 gnd.n7424 gnd.n7423 99.6594
R14828 gnd.n7419 gnd.n7418 99.6594
R14829 gnd.n3965 gnd.n3888 99.6594
R14830 gnd.n3957 gnd.n3876 99.6594
R14831 gnd.n3953 gnd.n3877 99.6594
R14832 gnd.n3949 gnd.n3878 99.6594
R14833 gnd.n3945 gnd.n3879 99.6594
R14834 gnd.n3941 gnd.n3880 99.6594
R14835 gnd.n3937 gnd.n3881 99.6594
R14836 gnd.n3933 gnd.n3882 99.6594
R14837 gnd.n3929 gnd.n3883 99.6594
R14838 gnd.n3925 gnd.n3884 99.6594
R14839 gnd.n3921 gnd.n3885 99.6594
R14840 gnd.n3917 gnd.n3886 99.6594
R14841 gnd.n3968 gnd.n3967 99.6594
R14842 gnd.n4669 gnd.n2002 99.6594
R14843 gnd.n4673 gnd.n2001 99.6594
R14844 gnd.n4677 gnd.n2000 99.6594
R14845 gnd.n4681 gnd.n1999 99.6594
R14846 gnd.n4685 gnd.n1998 99.6594
R14847 gnd.n4689 gnd.n1997 99.6594
R14848 gnd.n4693 gnd.n1996 99.6594
R14849 gnd.n4697 gnd.n1995 99.6594
R14850 gnd.n4701 gnd.n1994 99.6594
R14851 gnd.n4705 gnd.n1993 99.6594
R14852 gnd.n4709 gnd.n1992 99.6594
R14853 gnd.n4713 gnd.n1991 99.6594
R14854 gnd.n2031 gnd.n1990 99.6594
R14855 gnd.n4051 gnd.n4050 99.6594
R14856 gnd.n3810 gnd.n3788 99.6594
R14857 gnd.n3816 gnd.n3789 99.6594
R14858 gnd.n3820 gnd.n3790 99.6594
R14859 gnd.n3826 gnd.n3791 99.6594
R14860 gnd.n3830 gnd.n3792 99.6594
R14861 gnd.n3836 gnd.n3793 99.6594
R14862 gnd.n3794 gnd.n3778 99.6594
R14863 gnd.n4723 gnd.n2003 99.6594
R14864 gnd.n4727 gnd.n2004 99.6594
R14865 gnd.n4731 gnd.n2005 99.6594
R14866 gnd.n4735 gnd.n2006 99.6594
R14867 gnd.n4739 gnd.n2007 99.6594
R14868 gnd.n4743 gnd.n2008 99.6594
R14869 gnd.n4747 gnd.n2009 99.6594
R14870 gnd.n2012 gnd.n2010 99.6594
R14871 gnd.n5063 gnd.n5062 99.6594
R14872 gnd.n5057 gnd.n4876 99.6594
R14873 gnd.n5055 gnd.n5054 99.6594
R14874 gnd.n5050 gnd.n5049 99.6594
R14875 gnd.n5047 gnd.n5046 99.6594
R14876 gnd.n5042 gnd.n5041 99.6594
R14877 gnd.n5039 gnd.n5038 99.6594
R14878 gnd.n5034 gnd.n5033 99.6594
R14879 gnd.n5031 gnd.n5030 99.6594
R14880 gnd.n5026 gnd.n5025 99.6594
R14881 gnd.n5023 gnd.n5022 99.6594
R14882 gnd.n5018 gnd.n5017 99.6594
R14883 gnd.n5015 gnd.n5014 99.6594
R14884 gnd.n5010 gnd.n5009 99.6594
R14885 gnd.n5007 gnd.n5006 99.6594
R14886 gnd.n5002 gnd.n5001 99.6594
R14887 gnd.n4999 gnd.n4998 99.6594
R14888 gnd.n4931 gnd.n4930 99.6594
R14889 gnd.n4990 gnd.n4989 99.6594
R14890 gnd.n5703 gnd.n5702 99.6594
R14891 gnd.n1644 gnd.n1636 99.6594
R14892 gnd.n5710 gnd.n5709 99.6594
R14893 gnd.n1635 gnd.n1629 99.6594
R14894 gnd.n5717 gnd.n5716 99.6594
R14895 gnd.n1628 gnd.n1622 99.6594
R14896 gnd.n5724 gnd.n5723 99.6594
R14897 gnd.n1621 gnd.n1615 99.6594
R14898 gnd.n5731 gnd.n5730 99.6594
R14899 gnd.n1614 gnd.n1607 99.6594
R14900 gnd.n5740 gnd.n5739 99.6594
R14901 gnd.n1387 gnd.n1381 99.6594
R14902 gnd.n5747 gnd.n5746 99.6594
R14903 gnd.n1380 gnd.n1374 99.6594
R14904 gnd.n5754 gnd.n5753 99.6594
R14905 gnd.n1373 gnd.n1366 99.6594
R14906 gnd.n5761 gnd.n5760 99.6594
R14907 gnd.n5764 gnd.n5763 99.6594
R14908 gnd.n7047 gnd.n488 99.6594
R14909 gnd.n7041 gnd.n490 99.6594
R14910 gnd.n7037 gnd.n491 99.6594
R14911 gnd.n7033 gnd.n492 99.6594
R14912 gnd.n7029 gnd.n493 99.6594
R14913 gnd.n7025 gnd.n494 99.6594
R14914 gnd.n7021 gnd.n495 99.6594
R14915 gnd.n7016 gnd.n497 99.6594
R14916 gnd.n7012 gnd.n498 99.6594
R14917 gnd.n7008 gnd.n499 99.6594
R14918 gnd.n7004 gnd.n500 99.6594
R14919 gnd.n7000 gnd.n501 99.6594
R14920 gnd.n6996 gnd.n502 99.6594
R14921 gnd.n6992 gnd.n503 99.6594
R14922 gnd.n6988 gnd.n504 99.6594
R14923 gnd.n6984 gnd.n505 99.6594
R14924 gnd.n557 gnd.n506 99.6594
R14925 gnd.n6976 gnd.n507 99.6594
R14926 gnd.n194 gnd.n191 99.6594
R14927 gnd.n7505 gnd.n7504 99.6594
R14928 gnd.n190 gnd.n184 99.6594
R14929 gnd.n7512 gnd.n7511 99.6594
R14930 gnd.n183 gnd.n177 99.6594
R14931 gnd.n7519 gnd.n7518 99.6594
R14932 gnd.n176 gnd.n170 99.6594
R14933 gnd.n7526 gnd.n7525 99.6594
R14934 gnd.n169 gnd.n163 99.6594
R14935 gnd.n7533 gnd.n7532 99.6594
R14936 gnd.n162 gnd.n156 99.6594
R14937 gnd.n7543 gnd.n7542 99.6594
R14938 gnd.n155 gnd.n149 99.6594
R14939 gnd.n7550 gnd.n7549 99.6594
R14940 gnd.n148 gnd.n142 99.6594
R14941 gnd.n7557 gnd.n7556 99.6594
R14942 gnd.n141 gnd.n135 99.6594
R14943 gnd.n7564 gnd.n7563 99.6594
R14944 gnd.n134 gnd.n131 99.6594
R14945 gnd.n5581 gnd.n1319 99.6594
R14946 gnd.n5584 gnd.n1320 99.6594
R14947 gnd.n5594 gnd.n1321 99.6594
R14948 gnd.n5596 gnd.n1322 99.6594
R14949 gnd.n5607 gnd.n1323 99.6594
R14950 gnd.n5617 gnd.n1324 99.6594
R14951 gnd.n5619 gnd.n1325 99.6594
R14952 gnd.n5633 gnd.n1326 99.6594
R14953 gnd.n1345 gnd.n1327 99.6594
R14954 gnd.n5779 gnd.n1328 99.6594
R14955 gnd.n5788 gnd.n1329 99.6594
R14956 gnd.n5790 gnd.n1330 99.6594
R14957 gnd.n5798 gnd.n1331 99.6594
R14958 gnd.n5808 gnd.n1332 99.6594
R14959 gnd.n5583 gnd.n1319 99.6594
R14960 gnd.n5593 gnd.n1320 99.6594
R14961 gnd.n5595 gnd.n1321 99.6594
R14962 gnd.n5606 gnd.n1322 99.6594
R14963 gnd.n5616 gnd.n1323 99.6594
R14964 gnd.n5618 gnd.n1324 99.6594
R14965 gnd.n5632 gnd.n1325 99.6594
R14966 gnd.n1344 gnd.n1326 99.6594
R14967 gnd.n5780 gnd.n1327 99.6594
R14968 gnd.n5787 gnd.n1328 99.6594
R14969 gnd.n5791 gnd.n1329 99.6594
R14970 gnd.n5797 gnd.n1330 99.6594
R14971 gnd.n5801 gnd.n1331 99.6594
R14972 gnd.n5808 gnd.n5807 99.6594
R14973 gnd.n6758 gnd.n617 99.6594
R14974 gnd.n6631 gnd.n618 99.6594
R14975 gnd.n6633 gnd.n619 99.6594
R14976 gnd.n6641 gnd.n620 99.6594
R14977 gnd.n6651 gnd.n621 99.6594
R14978 gnd.n6653 gnd.n622 99.6594
R14979 gnd.n6661 gnd.n623 99.6594
R14980 gnd.n6671 gnd.n624 99.6594
R14981 gnd.n6673 gnd.n625 99.6594
R14982 gnd.n6678 gnd.n626 99.6594
R14983 gnd.n6680 gnd.n627 99.6594
R14984 gnd.n6684 gnd.n628 99.6594
R14985 gnd.n6686 gnd.n629 99.6594
R14986 gnd.n6693 gnd.n630 99.6594
R14987 gnd.n631 gnd.n630 99.6594
R14988 gnd.n6692 gnd.n629 99.6594
R14989 gnd.n6685 gnd.n628 99.6594
R14990 gnd.n6683 gnd.n627 99.6594
R14991 gnd.n6679 gnd.n626 99.6594
R14992 gnd.n6677 gnd.n625 99.6594
R14993 gnd.n6672 gnd.n624 99.6594
R14994 gnd.n6670 gnd.n623 99.6594
R14995 gnd.n6660 gnd.n622 99.6594
R14996 gnd.n6652 gnd.n621 99.6594
R14997 gnd.n6650 gnd.n620 99.6594
R14998 gnd.n6640 gnd.n619 99.6594
R14999 gnd.n6632 gnd.n618 99.6594
R15000 gnd.n6630 gnd.n617 99.6594
R15001 gnd.n1336 gnd.t97 98.63
R15002 gnd.n118 gnd.t30 98.63
R15003 gnd.n6712 gnd.t70 98.63
R15004 gnd.n1348 gnd.t82 98.63
R15005 gnd.n537 gnd.t63 98.63
R15006 gnd.n559 gnd.t35 98.63
R15007 gnd.n197 gnd.t108 98.63
R15008 gnd.n7536 gnd.t117 98.63
R15009 gnd.n4900 gnd.t56 98.63
R15010 gnd.n4932 gnd.t27 98.63
R15011 gnd.n4761 gnd.t93 98.63
R15012 gnd.n1641 gnd.t45 98.63
R15013 gnd.n1388 gnd.t79 98.63
R15014 gnd.n6689 gnd.t76 98.63
R15015 gnd.n1394 gnd.t112 96.6984
R15016 gnd.n804 gnd.t49 96.6984
R15017 gnd.n1450 gnd.t60 96.6906
R15018 gnd.n785 gnd.t102 96.6906
R15019 gnd.n2828 gnd.n2827 89.3769
R15020 gnd.n2827 gnd.n2497 89.3769
R15021 gnd.n2819 gnd.n2497 89.3769
R15022 gnd.n2819 gnd.n2818 89.3769
R15023 gnd.n2818 gnd.n2817 89.3769
R15024 gnd.n2817 gnd.n2505 89.3769
R15025 gnd.n2811 gnd.n2505 89.3769
R15026 gnd.n2811 gnd.n2810 89.3769
R15027 gnd.n2810 gnd.n2809 89.3769
R15028 gnd.n2809 gnd.n2512 89.3769
R15029 gnd.n2803 gnd.n2512 89.3769
R15030 gnd.n2803 gnd.n2802 89.3769
R15031 gnd.n2802 gnd.n2801 89.3769
R15032 gnd.n2801 gnd.n2520 89.3769
R15033 gnd.n2795 gnd.n2520 89.3769
R15034 gnd.n2795 gnd.n2794 89.3769
R15035 gnd.n2794 gnd.n2793 89.3769
R15036 gnd.n2793 gnd.n2528 89.3769
R15037 gnd.n2787 gnd.n2528 89.3769
R15038 gnd.n2787 gnd.n2786 89.3769
R15039 gnd.n2786 gnd.n2785 89.3769
R15040 gnd.n2785 gnd.n2536 89.3769
R15041 gnd.n2779 gnd.n2536 89.3769
R15042 gnd.n2779 gnd.n2778 89.3769
R15043 gnd.n2778 gnd.n2777 89.3769
R15044 gnd.n2777 gnd.n2544 89.3769
R15045 gnd.n2771 gnd.n2544 89.3769
R15046 gnd.n2771 gnd.n2770 89.3769
R15047 gnd.n2770 gnd.n2769 89.3769
R15048 gnd.n2769 gnd.n2552 89.3769
R15049 gnd.n2763 gnd.n2552 89.3769
R15050 gnd.n2763 gnd.n2762 89.3769
R15051 gnd.n2762 gnd.n2761 89.3769
R15052 gnd.n2761 gnd.n2560 89.3769
R15053 gnd.n2755 gnd.n2560 89.3769
R15054 gnd.n2755 gnd.n2754 89.3769
R15055 gnd.n2754 gnd.n2753 89.3769
R15056 gnd.n2753 gnd.n2568 89.3769
R15057 gnd.n2747 gnd.n2568 89.3769
R15058 gnd.n2747 gnd.n2746 89.3769
R15059 gnd.n2746 gnd.n2745 89.3769
R15060 gnd.n2745 gnd.n2576 89.3769
R15061 gnd.n2739 gnd.n2576 89.3769
R15062 gnd.n2739 gnd.n2738 89.3769
R15063 gnd.n2738 gnd.n2737 89.3769
R15064 gnd.n2737 gnd.n2584 89.3769
R15065 gnd.n2731 gnd.n2584 89.3769
R15066 gnd.n2731 gnd.n2730 89.3769
R15067 gnd.n2730 gnd.n2729 89.3769
R15068 gnd.n2729 gnd.n2592 89.3769
R15069 gnd.n2723 gnd.n2592 89.3769
R15070 gnd.n2723 gnd.n2722 89.3769
R15071 gnd.n2722 gnd.n2721 89.3769
R15072 gnd.n2721 gnd.n2600 89.3769
R15073 gnd.n2715 gnd.n2600 89.3769
R15074 gnd.n2715 gnd.n2714 89.3769
R15075 gnd.n2714 gnd.n2713 89.3769
R15076 gnd.n2713 gnd.n2608 89.3769
R15077 gnd.n2707 gnd.n2608 89.3769
R15078 gnd.n2707 gnd.n2706 89.3769
R15079 gnd.n2706 gnd.n2705 89.3769
R15080 gnd.n2705 gnd.n2616 89.3769
R15081 gnd.n2699 gnd.n2616 89.3769
R15082 gnd.n2699 gnd.n2698 89.3769
R15083 gnd.n2698 gnd.n2697 89.3769
R15084 gnd.n2697 gnd.n2624 89.3769
R15085 gnd.n2691 gnd.n2624 89.3769
R15086 gnd.n2691 gnd.n2690 89.3769
R15087 gnd.n2690 gnd.n2689 89.3769
R15088 gnd.n2689 gnd.n2632 89.3769
R15089 gnd.n2683 gnd.n2632 89.3769
R15090 gnd.n2683 gnd.n2682 89.3769
R15091 gnd.n2682 gnd.n2681 89.3769
R15092 gnd.n2681 gnd.n2640 89.3769
R15093 gnd.n2675 gnd.n2640 89.3769
R15094 gnd.n2675 gnd.n2674 89.3769
R15095 gnd.n2674 gnd.n2673 89.3769
R15096 gnd.n2673 gnd.n2648 89.3769
R15097 gnd.n2667 gnd.n2648 89.3769
R15098 gnd.n2667 gnd.n2666 89.3769
R15099 gnd.n2666 gnd.n2665 89.3769
R15100 gnd.n2665 gnd.n2657 89.3769
R15101 gnd.n2657 gnd.n2656 89.3769
R15102 gnd.n1423 gnd.n1422 81.8399
R15103 gnd.n3839 gnd.t22 74.8376
R15104 gnd.n2028 gnd.t67 74.8376
R15105 gnd.n1395 gnd.t111 72.8438
R15106 gnd.n805 gnd.t50 72.8438
R15107 gnd.n1424 gnd.n1417 72.8411
R15108 gnd.n1430 gnd.n1415 72.8411
R15109 gnd.n724 gnd.n723 72.8411
R15110 gnd.n1337 gnd.t96 72.836
R15111 gnd.n1451 gnd.t59 72.836
R15112 gnd.n786 gnd.t103 72.836
R15113 gnd.n119 gnd.t31 72.836
R15114 gnd.n6713 gnd.t69 72.836
R15115 gnd.n1349 gnd.t83 72.836
R15116 gnd.n538 gnd.t62 72.836
R15117 gnd.n560 gnd.t34 72.836
R15118 gnd.n198 gnd.t109 72.836
R15119 gnd.n7537 gnd.t118 72.836
R15120 gnd.n4901 gnd.t55 72.836
R15121 gnd.n4933 gnd.t26 72.836
R15122 gnd.n4762 gnd.t92 72.836
R15123 gnd.n1642 gnd.t46 72.836
R15124 gnd.n1389 gnd.t80 72.836
R15125 gnd.n6690 gnd.t77 72.836
R15126 gnd.n732 gnd.n731 71.676
R15127 gnd.n733 gnd.n707 71.676
R15128 gnd.n740 gnd.n739 71.676
R15129 gnd.n741 gnd.n705 71.676
R15130 gnd.n748 gnd.n747 71.676
R15131 gnd.n749 gnd.n703 71.676
R15132 gnd.n756 gnd.n755 71.676
R15133 gnd.n757 gnd.n701 71.676
R15134 gnd.n764 gnd.n763 71.676
R15135 gnd.n765 gnd.n699 71.676
R15136 gnd.n772 gnd.n771 71.676
R15137 gnd.n773 gnd.n697 71.676
R15138 gnd.n780 gnd.n779 71.676
R15139 gnd.n781 gnd.n695 71.676
R15140 gnd.n791 gnd.n790 71.676
R15141 gnd.n795 gnd.n693 71.676
R15142 gnd.n799 gnd.n798 71.676
R15143 gnd.n800 gnd.n692 71.676
R15144 gnd.n810 gnd.n809 71.676
R15145 gnd.n811 gnd.n690 71.676
R15146 gnd.n818 gnd.n817 71.676
R15147 gnd.n819 gnd.n688 71.676
R15148 gnd.n826 gnd.n825 71.676
R15149 gnd.n827 gnd.n686 71.676
R15150 gnd.n834 gnd.n833 71.676
R15151 gnd.n835 gnd.n684 71.676
R15152 gnd.n842 gnd.n841 71.676
R15153 gnd.n843 gnd.n682 71.676
R15154 gnd.n850 gnd.n849 71.676
R15155 gnd.n851 gnd.n680 71.676
R15156 gnd.n858 gnd.n857 71.676
R15157 gnd.n862 gnd.n678 71.676
R15158 gnd.n865 gnd.n864 71.676
R15159 gnd.n1516 gnd.n1435 71.676
R15160 gnd.n1511 gnd.n1437 71.676
R15161 gnd.n1507 gnd.n1506 71.676
R15162 gnd.n1500 gnd.n1439 71.676
R15163 gnd.n1499 gnd.n1498 71.676
R15164 gnd.n1492 gnd.n1441 71.676
R15165 gnd.n1491 gnd.n1490 71.676
R15166 gnd.n1484 gnd.n1443 71.676
R15167 gnd.n1483 gnd.n1482 71.676
R15168 gnd.n1476 gnd.n1445 71.676
R15169 gnd.n1475 gnd.n1474 71.676
R15170 gnd.n1468 gnd.n1447 71.676
R15171 gnd.n1467 gnd.n1466 71.676
R15172 gnd.n1460 gnd.n1449 71.676
R15173 gnd.n1459 gnd.n1453 71.676
R15174 gnd.n1455 gnd.n1454 71.676
R15175 gnd.n1602 gnd.n1601 71.676
R15176 gnd.n1594 gnd.n1393 71.676
R15177 gnd.n1593 gnd.n1592 71.676
R15178 gnd.n1586 gnd.n1397 71.676
R15179 gnd.n1585 gnd.n1584 71.676
R15180 gnd.n1578 gnd.n1399 71.676
R15181 gnd.n1577 gnd.n1576 71.676
R15182 gnd.n1570 gnd.n1401 71.676
R15183 gnd.n1569 gnd.n1568 71.676
R15184 gnd.n1562 gnd.n1403 71.676
R15185 gnd.n1561 gnd.n1560 71.676
R15186 gnd.n1554 gnd.n1405 71.676
R15187 gnd.n1553 gnd.n1552 71.676
R15188 gnd.n1546 gnd.n1407 71.676
R15189 gnd.n1545 gnd.n1544 71.676
R15190 gnd.n1538 gnd.n1409 71.676
R15191 gnd.n1513 gnd.n1435 71.676
R15192 gnd.n1508 gnd.n1437 71.676
R15193 gnd.n1506 gnd.n1505 71.676
R15194 gnd.n1501 gnd.n1500 71.676
R15195 gnd.n1498 gnd.n1497 71.676
R15196 gnd.n1493 gnd.n1492 71.676
R15197 gnd.n1490 gnd.n1489 71.676
R15198 gnd.n1485 gnd.n1484 71.676
R15199 gnd.n1482 gnd.n1481 71.676
R15200 gnd.n1477 gnd.n1476 71.676
R15201 gnd.n1474 gnd.n1473 71.676
R15202 gnd.n1469 gnd.n1468 71.676
R15203 gnd.n1466 gnd.n1465 71.676
R15204 gnd.n1461 gnd.n1460 71.676
R15205 gnd.n1456 gnd.n1453 71.676
R15206 gnd.n1604 gnd.n1603 71.676
R15207 gnd.n1601 gnd.n1600 71.676
R15208 gnd.n1595 gnd.n1594 71.676
R15209 gnd.n1592 gnd.n1591 71.676
R15210 gnd.n1587 gnd.n1586 71.676
R15211 gnd.n1584 gnd.n1583 71.676
R15212 gnd.n1579 gnd.n1578 71.676
R15213 gnd.n1576 gnd.n1575 71.676
R15214 gnd.n1571 gnd.n1570 71.676
R15215 gnd.n1568 gnd.n1567 71.676
R15216 gnd.n1563 gnd.n1562 71.676
R15217 gnd.n1560 gnd.n1559 71.676
R15218 gnd.n1555 gnd.n1554 71.676
R15219 gnd.n1552 gnd.n1551 71.676
R15220 gnd.n1547 gnd.n1546 71.676
R15221 gnd.n1544 gnd.n1543 71.676
R15222 gnd.n1539 gnd.n1538 71.676
R15223 gnd.n864 gnd.n863 71.676
R15224 gnd.n859 gnd.n678 71.676
R15225 gnd.n857 gnd.n856 71.676
R15226 gnd.n852 gnd.n851 71.676
R15227 gnd.n849 gnd.n848 71.676
R15228 gnd.n844 gnd.n843 71.676
R15229 gnd.n841 gnd.n840 71.676
R15230 gnd.n836 gnd.n835 71.676
R15231 gnd.n833 gnd.n832 71.676
R15232 gnd.n828 gnd.n827 71.676
R15233 gnd.n825 gnd.n824 71.676
R15234 gnd.n820 gnd.n819 71.676
R15235 gnd.n817 gnd.n816 71.676
R15236 gnd.n812 gnd.n811 71.676
R15237 gnd.n809 gnd.n808 71.676
R15238 gnd.n801 gnd.n800 71.676
R15239 gnd.n797 gnd.n796 71.676
R15240 gnd.n792 gnd.n693 71.676
R15241 gnd.n790 gnd.n789 71.676
R15242 gnd.n782 gnd.n781 71.676
R15243 gnd.n779 gnd.n778 71.676
R15244 gnd.n774 gnd.n773 71.676
R15245 gnd.n771 gnd.n770 71.676
R15246 gnd.n766 gnd.n765 71.676
R15247 gnd.n763 gnd.n762 71.676
R15248 gnd.n758 gnd.n757 71.676
R15249 gnd.n755 gnd.n754 71.676
R15250 gnd.n750 gnd.n749 71.676
R15251 gnd.n747 gnd.n746 71.676
R15252 gnd.n742 gnd.n741 71.676
R15253 gnd.n739 gnd.n738 71.676
R15254 gnd.n734 gnd.n733 71.676
R15255 gnd.n731 gnd.n730 71.676
R15256 gnd.n8 gnd.t153 69.1507
R15257 gnd.n14 gnd.t155 68.4792
R15258 gnd.n13 gnd.t178 68.4792
R15259 gnd.n12 gnd.t168 68.4792
R15260 gnd.n11 gnd.t126 68.4792
R15261 gnd.n10 gnd.t164 68.4792
R15262 gnd.n9 gnd.t355 68.4792
R15263 gnd.n8 gnd.t124 68.4792
R15264 gnd.n3966 gnd.n3870 64.369
R15265 gnd.n1597 gnd.n1395 59.5399
R15266 gnd.n806 gnd.n805 59.5399
R15267 gnd.n1452 gnd.n1451 59.5399
R15268 gnd.n787 gnd.n786 59.5399
R15269 gnd.n1434 gnd.n1433 59.1804
R15270 gnd.n4755 gnd.n1988 57.3586
R15271 gnd.n3657 gnd.t195 56.607
R15272 gnd.n56 gnd.t325 56.607
R15273 gnd.n3618 gnd.t279 56.407
R15274 gnd.n3637 gnd.t253 56.407
R15275 gnd.n17 gnd.t317 56.407
R15276 gnd.n36 gnd.t287 56.407
R15277 gnd.n3674 gnd.t263 55.8337
R15278 gnd.n3635 gnd.t302 55.8337
R15279 gnd.n3654 gnd.t276 55.8337
R15280 gnd.n73 gnd.t334 55.8337
R15281 gnd.n34 gnd.t318 55.8337
R15282 gnd.n53 gnd.t289 55.8337
R15283 gnd.n1421 gnd.n1420 54.358
R15284 gnd.n721 gnd.n720 54.358
R15285 gnd.n2656 gnd.n236 53.6263
R15286 gnd.n3657 gnd.n3656 53.0052
R15287 gnd.n3659 gnd.n3658 53.0052
R15288 gnd.n3661 gnd.n3660 53.0052
R15289 gnd.n3663 gnd.n3662 53.0052
R15290 gnd.n3665 gnd.n3664 53.0052
R15291 gnd.n3667 gnd.n3666 53.0052
R15292 gnd.n3669 gnd.n3668 53.0052
R15293 gnd.n3671 gnd.n3670 53.0052
R15294 gnd.n3673 gnd.n3672 53.0052
R15295 gnd.n3618 gnd.n3617 53.0052
R15296 gnd.n3620 gnd.n3619 53.0052
R15297 gnd.n3622 gnd.n3621 53.0052
R15298 gnd.n3624 gnd.n3623 53.0052
R15299 gnd.n3626 gnd.n3625 53.0052
R15300 gnd.n3628 gnd.n3627 53.0052
R15301 gnd.n3630 gnd.n3629 53.0052
R15302 gnd.n3632 gnd.n3631 53.0052
R15303 gnd.n3634 gnd.n3633 53.0052
R15304 gnd.n3637 gnd.n3636 53.0052
R15305 gnd.n3639 gnd.n3638 53.0052
R15306 gnd.n3641 gnd.n3640 53.0052
R15307 gnd.n3643 gnd.n3642 53.0052
R15308 gnd.n3645 gnd.n3644 53.0052
R15309 gnd.n3647 gnd.n3646 53.0052
R15310 gnd.n3649 gnd.n3648 53.0052
R15311 gnd.n3651 gnd.n3650 53.0052
R15312 gnd.n3653 gnd.n3652 53.0052
R15313 gnd.n72 gnd.n71 53.0052
R15314 gnd.n70 gnd.n69 53.0052
R15315 gnd.n68 gnd.n67 53.0052
R15316 gnd.n66 gnd.n65 53.0052
R15317 gnd.n64 gnd.n63 53.0052
R15318 gnd.n62 gnd.n61 53.0052
R15319 gnd.n60 gnd.n59 53.0052
R15320 gnd.n58 gnd.n57 53.0052
R15321 gnd.n56 gnd.n55 53.0052
R15322 gnd.n33 gnd.n32 53.0052
R15323 gnd.n31 gnd.n30 53.0052
R15324 gnd.n29 gnd.n28 53.0052
R15325 gnd.n27 gnd.n26 53.0052
R15326 gnd.n25 gnd.n24 53.0052
R15327 gnd.n23 gnd.n22 53.0052
R15328 gnd.n21 gnd.n20 53.0052
R15329 gnd.n19 gnd.n18 53.0052
R15330 gnd.n17 gnd.n16 53.0052
R15331 gnd.n52 gnd.n51 53.0052
R15332 gnd.n50 gnd.n49 53.0052
R15333 gnd.n48 gnd.n47 53.0052
R15334 gnd.n46 gnd.n45 53.0052
R15335 gnd.n44 gnd.n43 53.0052
R15336 gnd.n42 gnd.n41 53.0052
R15337 gnd.n40 gnd.n39 53.0052
R15338 gnd.n38 gnd.n37 53.0052
R15339 gnd.n36 gnd.n35 53.0052
R15340 gnd.n712 gnd.n711 52.4801
R15341 gnd.n4609 gnd.t129 52.3082
R15342 gnd.n4577 gnd.t135 52.3082
R15343 gnd.n4545 gnd.t189 52.3082
R15344 gnd.n4514 gnd.t132 52.3082
R15345 gnd.n4482 gnd.t160 52.3082
R15346 gnd.n4450 gnd.t353 52.3082
R15347 gnd.n4418 gnd.t10 52.3082
R15348 gnd.n4387 gnd.t158 52.3082
R15349 gnd.n5070 gnd.n4756 51.6227
R15350 gnd.n7573 gnd.n124 51.6227
R15351 gnd.n4439 gnd.n4407 51.4173
R15352 gnd.n4503 gnd.n4502 50.455
R15353 gnd.n4471 gnd.n4470 50.455
R15354 gnd.n4439 gnd.n4438 50.455
R15355 gnd.n7018 gnd.n534 45.6325
R15356 gnd.n1606 gnd.n1605 45.6325
R15357 gnd.n3913 gnd.n3912 45.1884
R15358 gnd.n2054 gnd.n2053 45.1884
R15359 gnd.n728 gnd.n727 44.3322
R15360 gnd.n1424 gnd.n1423 44.3189
R15361 gnd.n5800 gnd.n1337 42.2793
R15362 gnd.n3914 gnd.n3913 42.2793
R15363 gnd.n2055 gnd.n2054 42.2793
R15364 gnd.n3840 gnd.n3839 42.2793
R15365 gnd.n4722 gnd.n2028 42.2793
R15366 gnd.n120 gnd.n119 42.2793
R15367 gnd.n6714 gnd.n6713 42.2793
R15368 gnd.n5775 gnd.n1349 42.2793
R15369 gnd.n561 gnd.n560 42.2793
R15370 gnd.n7501 gnd.n198 42.2793
R15371 gnd.n7538 gnd.n7537 42.2793
R15372 gnd.n4902 gnd.n4901 42.2793
R15373 gnd.n4934 gnd.n4933 42.2793
R15374 gnd.n4763 gnd.n4762 42.2793
R15375 gnd.n1643 gnd.n1642 42.2793
R15376 gnd.n6691 gnd.n6690 42.2793
R15377 gnd.n1422 gnd.n1421 41.6274
R15378 gnd.n722 gnd.n721 41.6274
R15379 gnd.n1431 gnd.n1430 40.8975
R15380 gnd.n725 gnd.n724 40.8975
R15381 gnd.n7018 gnd.n538 36.9518
R15382 gnd.n1606 gnd.n1389 36.9518
R15383 gnd.n1430 gnd.n1429 35.055
R15384 gnd.n1425 gnd.n1424 35.055
R15385 gnd.n714 gnd.n713 35.055
R15386 gnd.n724 gnd.n710 35.055
R15387 gnd.n867 gnd.n866 32.9371
R15388 gnd.n1540 gnd.n1410 32.9371
R15389 gnd.n3143 gnd.n3142 32.6173
R15390 gnd.n3143 gnd.n2183 32.6173
R15391 gnd.n3151 gnd.n2183 32.6173
R15392 gnd.n3152 gnd.n3151 32.6173
R15393 gnd.n3153 gnd.n3152 32.6173
R15394 gnd.n3153 gnd.n2177 32.6173
R15395 gnd.n3161 gnd.n2177 32.6173
R15396 gnd.n3162 gnd.n3161 32.6173
R15397 gnd.n3163 gnd.n3162 32.6173
R15398 gnd.n3163 gnd.n2171 32.6173
R15399 gnd.n3171 gnd.n2171 32.6173
R15400 gnd.n3172 gnd.n3171 32.6173
R15401 gnd.n3173 gnd.n3172 32.6173
R15402 gnd.n3173 gnd.n2165 32.6173
R15403 gnd.n3181 gnd.n2165 32.6173
R15404 gnd.n3182 gnd.n3181 32.6173
R15405 gnd.n3183 gnd.n3182 32.6173
R15406 gnd.n3183 gnd.n2159 32.6173
R15407 gnd.n3191 gnd.n2159 32.6173
R15408 gnd.n3192 gnd.n3191 32.6173
R15409 gnd.n3193 gnd.n3192 32.6173
R15410 gnd.n3193 gnd.n2153 32.6173
R15411 gnd.n3201 gnd.n2153 32.6173
R15412 gnd.n3202 gnd.n3201 32.6173
R15413 gnd.n3203 gnd.n3202 32.6173
R15414 gnd.n3203 gnd.n2147 32.6173
R15415 gnd.n3211 gnd.n2147 32.6173
R15416 gnd.n3212 gnd.n3211 32.6173
R15417 gnd.n3213 gnd.n3212 32.6173
R15418 gnd.n3213 gnd.n2141 32.6173
R15419 gnd.n3221 gnd.n2141 32.6173
R15420 gnd.n3222 gnd.n3221 32.6173
R15421 gnd.n3223 gnd.n3222 32.6173
R15422 gnd.n3223 gnd.n2135 32.6173
R15423 gnd.n3231 gnd.n2135 32.6173
R15424 gnd.n3232 gnd.n3231 32.6173
R15425 gnd.n3233 gnd.n3232 32.6173
R15426 gnd.n3233 gnd.n2129 32.6173
R15427 gnd.n3241 gnd.n2129 32.6173
R15428 gnd.n3242 gnd.n3241 32.6173
R15429 gnd.n3243 gnd.n3242 32.6173
R15430 gnd.n3243 gnd.n2123 32.6173
R15431 gnd.n3251 gnd.n2123 32.6173
R15432 gnd.n3252 gnd.n3251 32.6173
R15433 gnd.n3253 gnd.n3252 32.6173
R15434 gnd.n3253 gnd.n2117 32.6173
R15435 gnd.n3261 gnd.n2117 32.6173
R15436 gnd.n3262 gnd.n3261 32.6173
R15437 gnd.n3263 gnd.n3262 32.6173
R15438 gnd.n3263 gnd.n2111 32.6173
R15439 gnd.n3271 gnd.n2111 32.6173
R15440 gnd.n3272 gnd.n3271 32.6173
R15441 gnd.n3273 gnd.n3272 32.6173
R15442 gnd.n3273 gnd.n2105 32.6173
R15443 gnd.n3281 gnd.n2105 32.6173
R15444 gnd.n3282 gnd.n3281 32.6173
R15445 gnd.n3283 gnd.n3282 32.6173
R15446 gnd.n3283 gnd.n2099 32.6173
R15447 gnd.n3291 gnd.n2099 32.6173
R15448 gnd.n3292 gnd.n3291 32.6173
R15449 gnd.n3293 gnd.n3292 32.6173
R15450 gnd.n3293 gnd.n2093 32.6173
R15451 gnd.n3301 gnd.n2093 32.6173
R15452 gnd.n3302 gnd.n3301 32.6173
R15453 gnd.n3303 gnd.n3302 32.6173
R15454 gnd.n3303 gnd.n2087 32.6173
R15455 gnd.n3311 gnd.n2087 32.6173
R15456 gnd.n3312 gnd.n3311 32.6173
R15457 gnd.n3313 gnd.n3312 32.6173
R15458 gnd.n3313 gnd.n2081 32.6173
R15459 gnd.n3321 gnd.n2081 32.6173
R15460 gnd.n3322 gnd.n3321 32.6173
R15461 gnd.n3323 gnd.n3322 32.6173
R15462 gnd.n3323 gnd.n2075 32.6173
R15463 gnd.n3331 gnd.n2075 32.6173
R15464 gnd.n3332 gnd.n3331 32.6173
R15465 gnd.n3333 gnd.n3332 32.6173
R15466 gnd.n3333 gnd.n2069 32.6173
R15467 gnd.n3341 gnd.n2069 32.6173
R15468 gnd.n3342 gnd.n3341 32.6173
R15469 gnd.n3343 gnd.n3342 32.6173
R15470 gnd.n3343 gnd.n2062 32.6173
R15471 gnd.n3354 gnd.n2062 32.6173
R15472 gnd.n3976 gnd.n3870 31.8661
R15473 gnd.n3976 gnd.n3975 31.8661
R15474 gnd.n3984 gnd.n3859 31.8661
R15475 gnd.n3992 gnd.n3859 31.8661
R15476 gnd.n3992 gnd.n3853 31.8661
R15477 gnd.n4000 gnd.n3853 31.8661
R15478 gnd.n4000 gnd.n3846 31.8661
R15479 gnd.n4038 gnd.n3846 31.8661
R15480 gnd.n4048 gnd.n3779 31.8661
R15481 gnd.n5070 gnd.n4872 31.8661
R15482 gnd.n5078 gnd.n1974 31.8661
R15483 gnd.n5086 gnd.n1974 31.8661
R15484 gnd.n5086 gnd.n1966 31.8661
R15485 gnd.n5094 gnd.n1966 31.8661
R15486 gnd.n5102 gnd.n1957 31.8661
R15487 gnd.n5102 gnd.n1960 31.8661
R15488 gnd.n5110 gnd.n1942 31.8661
R15489 gnd.n5118 gnd.n1942 31.8661
R15490 gnd.n5126 gnd.n1934 31.8661
R15491 gnd.n5134 gnd.n1925 31.8661
R15492 gnd.n5134 gnd.n1928 31.8661
R15493 gnd.n5150 gnd.n1908 31.8661
R15494 gnd.n5160 gnd.n1908 31.8661
R15495 gnd.n5173 gnd.n1902 31.8661
R15496 gnd.n5190 gnd.n1884 31.8661
R15497 gnd.n5184 gnd.n1884 31.8661
R15498 gnd.n5199 gnd.n1867 31.8661
R15499 gnd.n5217 gnd.n1867 31.8661
R15500 gnd.n5461 gnd.n1775 31.8661
R15501 gnd.n5455 gnd.n1786 31.8661
R15502 gnd.n5358 gnd.n1356 31.8661
R15503 gnd.n5351 gnd.n1318 31.8661
R15504 gnd.n5809 gnd.n1318 31.8661
R15505 gnd.n5809 gnd.n1310 31.8661
R15506 gnd.n5817 gnd.n1310 31.8661
R15507 gnd.n5817 gnd.n1312 31.8661
R15508 gnd.n6808 gnd.n639 31.8661
R15509 gnd.n639 gnd.n616 31.8661
R15510 gnd.n6817 gnd.n616 31.8661
R15511 gnd.n6817 gnd.n6816 31.8661
R15512 gnd.n6816 gnd.n489 31.8661
R15513 gnd.n564 gnd.n518 31.8661
R15514 gnd.n7228 gnd.n336 31.8661
R15515 gnd.n7301 gnd.n330 31.8661
R15516 gnd.n7305 gnd.n295 31.8661
R15517 gnd.n7329 gnd.n295 31.8661
R15518 gnd.n7337 gnd.n286 31.8661
R15519 gnd.n7337 gnd.n289 31.8661
R15520 gnd.n7345 gnd.n280 31.8661
R15521 gnd.n7353 gnd.n265 31.8661
R15522 gnd.n7361 gnd.n265 31.8661
R15523 gnd.n7369 gnd.n256 31.8661
R15524 gnd.n7369 gnd.n259 31.8661
R15525 gnd.n7377 gnd.n250 31.8661
R15526 gnd.n7385 gnd.n234 31.8661
R15527 gnd.n7393 gnd.n234 31.8661
R15528 gnd.n7401 gnd.n225 31.8661
R15529 gnd.n7401 gnd.n228 31.8661
R15530 gnd.n7409 gnd.n209 31.8661
R15531 gnd.n7485 gnd.n209 31.8661
R15532 gnd.n7485 gnd.n202 31.8661
R15533 gnd.n7493 gnd.n202 31.8661
R15534 gnd.n7573 gnd.n122 31.8661
R15535 gnd.n5461 gnd.t247 31.5474
R15536 gnd.n7301 gnd.t314 31.5474
R15537 gnd.t282 gnd.n1902 30.9101
R15538 gnd.n280 gnd.t239 30.9101
R15539 gnd.t227 gnd.n1934 30.2728
R15540 gnd.n250 gnd.t213 30.2728
R15541 gnd.n4872 gnd.t25 28.3609
R15542 gnd.t29 gnd.n122 28.3609
R15543 gnd.n5351 gnd.n1364 27.4049
R15544 gnd.n7046 gnd.n489 27.4049
R15545 gnd.n1337 gnd.n1336 25.7944
R15546 gnd.n3839 gnd.n3838 25.7944
R15547 gnd.n2028 gnd.n2027 25.7944
R15548 gnd.n119 gnd.n118 25.7944
R15549 gnd.n6713 gnd.n6712 25.7944
R15550 gnd.n1349 gnd.n1348 25.7944
R15551 gnd.n538 gnd.n537 25.7944
R15552 gnd.n560 gnd.n559 25.7944
R15553 gnd.n198 gnd.n197 25.7944
R15554 gnd.n7537 gnd.n7536 25.7944
R15555 gnd.n4901 gnd.n4900 25.7944
R15556 gnd.n4933 gnd.n4932 25.7944
R15557 gnd.n4762 gnd.n4761 25.7944
R15558 gnd.n1642 gnd.n1641 25.7944
R15559 gnd.n1389 gnd.n1388 25.7944
R15560 gnd.n6690 gnd.n6689 25.7944
R15561 gnd.n4060 gnd.n3780 24.8557
R15562 gnd.n4070 gnd.n3763 24.8557
R15563 gnd.n3766 gnd.n3754 24.8557
R15564 gnd.n4091 gnd.n3755 24.8557
R15565 gnd.n4101 gnd.n3735 24.8557
R15566 gnd.n4111 gnd.n4110 24.8557
R15567 gnd.n3719 gnd.n3718 24.8557
R15568 gnd.n4148 gnd.n3711 24.8557
R15569 gnd.n4147 gnd.n3704 24.8557
R15570 gnd.n4185 gnd.n3683 24.8557
R15571 gnd.n4159 gnd.n3684 24.8557
R15572 gnd.n4178 gnd.n3531 24.8557
R15573 gnd.n4195 gnd.n4194 24.8557
R15574 gnd.n4206 gnd.n4205 24.8557
R15575 gnd.n3523 gnd.n3514 24.8557
R15576 gnd.n4226 gnd.n3497 24.8557
R15577 gnd.n3500 gnd.n3489 24.8557
R15578 gnd.n4247 gnd.n3490 24.8557
R15579 gnd.n4256 gnd.n3482 24.8557
R15580 gnd.n4257 gnd.n3471 24.8557
R15581 gnd.n3474 gnd.n3462 24.8557
R15582 gnd.n4278 gnd.n3463 24.8557
R15583 gnd.n4288 gnd.n3446 24.8557
R15584 gnd.n4299 gnd.n4298 24.8557
R15585 gnd.n3588 gnd.n3587 24.8557
R15586 gnd.n4309 gnd.n3438 24.8557
R15587 gnd.n4319 gnd.n3421 24.8557
R15588 gnd.n4330 gnd.n4329 24.8557
R15589 gnd.n4340 gnd.n3413 24.8557
R15590 gnd.n4350 gnd.n3395 24.8557
R15591 gnd.n4361 gnd.n4360 24.8557
R15592 gnd.n4371 gnd.n3388 24.8557
R15593 gnd.n4636 gnd.n3380 24.8557
R15594 gnd.n4637 gnd.n3370 24.8557
R15595 gnd.n1395 gnd.n1394 23.855
R15596 gnd.n805 gnd.n804 23.855
R15597 gnd.n1451 gnd.n1450 23.855
R15598 gnd.n786 gnd.n785 23.855
R15599 gnd.n4081 gnd.t157 23.2624
R15600 gnd.n5094 gnd.t262 23.2624
R15601 gnd.n5677 gnd.n1305 23.2624
R15602 gnd.n6798 gnd.n648 23.2624
R15603 gnd.n7409 gnd.t288 23.2624
R15604 gnd.n3782 gnd.t21 22.6251
R15605 gnd.n5126 gnd.t231 22.6251
R15606 gnd.n7377 gnd.t196 22.6251
R15607 gnd.n5173 gnd.t204 21.9878
R15608 gnd.n7345 gnd.t255 21.9878
R15609 gnd.n5983 gnd.n1264 21.6691
R15610 gnd.n5975 gnd.n1256 21.6691
R15611 gnd.n5911 gnd.n1241 21.6691
R15612 gnd.n5927 gnd.n1225 21.6691
R15613 gnd.n5947 gnd.n1218 21.6691
R15614 gnd.n6125 gnd.n1111 21.6691
R15615 gnd.n6110 gnd.n1095 21.6691
R15616 gnd.n6102 gnd.n1087 21.6691
R15617 gnd.n6095 gnd.n1080 21.6691
R15618 gnd.n6087 gnd.n1149 21.6691
R15619 gnd.n6081 gnd.n6080 21.6691
R15620 gnd.n6430 gnd.n1022 21.6691
R15621 gnd.n6430 gnd.n1025 21.6691
R15622 gnd.n6415 gnd.n1008 21.6691
R15623 gnd.n6289 gnd.n1000 21.6691
R15624 gnd.n6267 gnd.n992 21.6691
R15625 gnd.n6307 gnd.n984 21.6691
R15626 gnd.n6316 gnd.n6256 21.6691
R15627 gnd.n6335 gnd.n6247 21.6691
R15628 gnd.n6352 gnd.n937 21.6691
R15629 gnd.n6380 gnd.n928 21.6691
R15630 gnd.n6552 gnd.n911 21.6691
R15631 gnd.n6569 gnd.n880 21.6691
R15632 gnd.n6769 gnd.n655 21.6691
R15633 gnd.t131 gnd.n3787 21.3504
R15634 gnd.t206 gnd.n1775 21.3504
R15635 gnd.n1788 gnd.n1786 21.3504
R15636 gnd.n5233 gnd.t229 21.3504
R15637 gnd.n7202 gnd.t218 21.3504
R15638 gnd.n7221 gnd.n336 21.3504
R15639 gnd.t305 gnd.n330 21.3504
R15640 gnd.n1518 gnd.n1434 20.7615
R15641 gnd.n728 gnd.n674 20.7615
R15642 gnd.t140 gnd.n3412 20.7131
R15643 gnd.n5199 gnd.t245 20.7131
R15644 gnd.n7329 gnd.t258 20.7131
R15645 gnd.t18 gnd.n1297 20.3945
R15646 gnd.n1411 gnd.n1287 20.3945
R15647 gnd.n5991 gnd.n1254 20.3945
R15648 gnd.n5939 gnd.n1199 20.3945
R15649 gnd.n6133 gnd.n1101 20.3945
R15650 gnd.n1163 gnd.n1049 20.3945
R15651 gnd.n6438 gnd.n1014 20.3945
R15652 gnd.n6325 gnd.n961 20.3945
R15653 gnd.n6242 gnd.n955 20.3945
R15654 gnd.n4287 gnd.t142 20.0758
R15655 gnd.n5150 gnd.t265 20.0758
R15656 gnd.t154 gnd.t48 20.0758
R15657 gnd.n7361 gnd.t296 20.0758
R15658 gnd.n1418 gnd.t115 19.8005
R15659 gnd.n1418 gnd.t16 19.8005
R15660 gnd.n1419 gnd.t19 19.8005
R15661 gnd.n1419 gnd.t53 19.8005
R15662 gnd.n718 gnd.t73 19.8005
R15663 gnd.n718 gnd.t42 19.8005
R15664 gnd.n719 gnd.t86 19.8005
R15665 gnd.n719 gnd.t13 19.8005
R15666 gnd.n3355 gnd.n3354 19.5706
R15667 gnd.n1415 gnd.n1414 19.5087
R15668 gnd.n1428 gnd.n1415 19.5087
R15669 gnd.n1426 gnd.n1417 19.5087
R15670 gnd.n723 gnd.n717 19.5087
R15671 gnd.t144 gnd.n4236 19.4385
R15672 gnd.n5110 gnd.t208 19.4385
R15673 gnd.n5819 gnd.n1307 19.3944
R15674 gnd.n5823 gnd.n1307 19.3944
R15675 gnd.n5823 gnd.n1293 19.3944
R15676 gnd.n5837 gnd.n1293 19.3944
R15677 gnd.n5837 gnd.n1290 19.3944
R15678 gnd.n5842 gnd.n1290 19.3944
R15679 gnd.n5842 gnd.n1291 19.3944
R15680 gnd.n1291 gnd.n1252 19.3944
R15681 gnd.n5993 gnd.n1252 19.3944
R15682 gnd.n5993 gnd.n1250 19.3944
R15683 gnd.n5997 gnd.n1250 19.3944
R15684 gnd.n5997 gnd.n1237 19.3944
R15685 gnd.n6009 gnd.n1237 19.3944
R15686 gnd.n6009 gnd.n1235 19.3944
R15687 gnd.n6013 gnd.n1235 19.3944
R15688 gnd.n6013 gnd.n1222 19.3944
R15689 gnd.n6025 gnd.n1222 19.3944
R15690 gnd.n6025 gnd.n1220 19.3944
R15691 gnd.n6029 gnd.n1220 19.3944
R15692 gnd.n6029 gnd.n1205 19.3944
R15693 gnd.n6042 gnd.n1205 19.3944
R15694 gnd.n6042 gnd.n1202 19.3944
R15695 gnd.n6047 gnd.n1202 19.3944
R15696 gnd.n6047 gnd.n1203 19.3944
R15697 gnd.n1203 gnd.n1099 19.3944
R15698 gnd.n6135 gnd.n1099 19.3944
R15699 gnd.n6135 gnd.n1097 19.3944
R15700 gnd.n6139 gnd.n1097 19.3944
R15701 gnd.n6139 gnd.n1084 19.3944
R15702 gnd.n6151 gnd.n1084 19.3944
R15703 gnd.n6151 gnd.n1082 19.3944
R15704 gnd.n6155 gnd.n1082 19.3944
R15705 gnd.n6155 gnd.n1070 19.3944
R15706 gnd.n6167 gnd.n1070 19.3944
R15707 gnd.n6167 gnd.n1068 19.3944
R15708 gnd.n6171 gnd.n1068 19.3944
R15709 gnd.n6171 gnd.n1054 19.3944
R15710 gnd.n6185 gnd.n1054 19.3944
R15711 gnd.n6185 gnd.n1051 19.3944
R15712 gnd.n6190 gnd.n1051 19.3944
R15713 gnd.n6190 gnd.n1052 19.3944
R15714 gnd.n1052 gnd.n1012 19.3944
R15715 gnd.n6440 gnd.n1012 19.3944
R15716 gnd.n6440 gnd.n1010 19.3944
R15717 gnd.n6444 gnd.n1010 19.3944
R15718 gnd.n6444 gnd.n996 19.3944
R15719 gnd.n6456 gnd.n996 19.3944
R15720 gnd.n6456 gnd.n994 19.3944
R15721 gnd.n6460 gnd.n994 19.3944
R15722 gnd.n6460 gnd.n981 19.3944
R15723 gnd.n6472 gnd.n981 19.3944
R15724 gnd.n6472 gnd.n979 19.3944
R15725 gnd.n6476 gnd.n979 19.3944
R15726 gnd.n6476 gnd.n966 19.3944
R15727 gnd.n6488 gnd.n966 19.3944
R15728 gnd.n6488 gnd.n964 19.3944
R15729 gnd.n6492 gnd.n964 19.3944
R15730 gnd.n6492 gnd.n951 19.3944
R15731 gnd.n6504 gnd.n951 19.3944
R15732 gnd.n6504 gnd.n949 19.3944
R15733 gnd.n6508 gnd.n949 19.3944
R15734 gnd.n6508 gnd.n935 19.3944
R15735 gnd.n6519 gnd.n935 19.3944
R15736 gnd.n6519 gnd.n932 19.3944
R15737 gnd.n6530 gnd.n932 19.3944
R15738 gnd.n6530 gnd.n933 19.3944
R15739 gnd.n6526 gnd.n933 19.3944
R15740 gnd.n6526 gnd.n6525 19.3944
R15741 gnd.n6525 gnd.n893 19.3944
R15742 gnd.n6588 gnd.n893 19.3944
R15743 gnd.n6588 gnd.n894 19.3944
R15744 gnd.n6584 gnd.n894 19.3944
R15745 gnd.n6584 gnd.n6583 19.3944
R15746 gnd.n6583 gnd.n6582 19.3944
R15747 gnd.n6582 gnd.n6579 19.3944
R15748 gnd.n6579 gnd.n652 19.3944
R15749 gnd.n6791 gnd.n652 19.3944
R15750 gnd.n6791 gnd.n650 19.3944
R15751 gnd.n6796 gnd.n650 19.3944
R15752 gnd.n6796 gnd.n636 19.3944
R15753 gnd.n6810 gnd.n636 19.3944
R15754 gnd.n6811 gnd.n6810 19.3944
R15755 gnd.n5802 gnd.n1333 19.3944
R15756 gnd.n5806 gnd.n1333 19.3944
R15757 gnd.n5806 gnd.n1334 19.3944
R15758 gnd.n5669 gnd.n5582 19.3944
R15759 gnd.n5669 gnd.n5668 19.3944
R15760 gnd.n5668 gnd.n5585 19.3944
R15761 gnd.n5661 gnd.n5585 19.3944
R15762 gnd.n5661 gnd.n5660 19.3944
R15763 gnd.n5660 gnd.n5597 19.3944
R15764 gnd.n5653 gnd.n5597 19.3944
R15765 gnd.n5653 gnd.n5652 19.3944
R15766 gnd.n5652 gnd.n5608 19.3944
R15767 gnd.n5645 gnd.n5608 19.3944
R15768 gnd.n5645 gnd.n5644 19.3944
R15769 gnd.n5644 gnd.n5620 19.3944
R15770 gnd.n5637 gnd.n5620 19.3944
R15771 gnd.n5637 gnd.n5636 19.3944
R15772 gnd.n5636 gnd.n1343 19.3944
R15773 gnd.n5778 gnd.n1343 19.3944
R15774 gnd.n5781 gnd.n5778 19.3944
R15775 gnd.n5781 gnd.n1340 19.3944
R15776 gnd.n5786 gnd.n1340 19.3944
R15777 gnd.n5789 gnd.n5786 19.3944
R15778 gnd.n5792 gnd.n5789 19.3944
R15779 gnd.n5792 gnd.n1338 19.3944
R15780 gnd.n5796 gnd.n1338 19.3944
R15781 gnd.n5799 gnd.n5796 19.3944
R15782 gnd.n3963 gnd.n3962 19.3944
R15783 gnd.n3962 gnd.n3961 19.3944
R15784 gnd.n3961 gnd.n3960 19.3944
R15785 gnd.n3960 gnd.n3958 19.3944
R15786 gnd.n3958 gnd.n3955 19.3944
R15787 gnd.n3955 gnd.n3954 19.3944
R15788 gnd.n3954 gnd.n3951 19.3944
R15789 gnd.n3951 gnd.n3950 19.3944
R15790 gnd.n3950 gnd.n3947 19.3944
R15791 gnd.n3947 gnd.n3946 19.3944
R15792 gnd.n3946 gnd.n3943 19.3944
R15793 gnd.n3943 gnd.n3942 19.3944
R15794 gnd.n3942 gnd.n3939 19.3944
R15795 gnd.n3939 gnd.n3938 19.3944
R15796 gnd.n3938 gnd.n3935 19.3944
R15797 gnd.n3935 gnd.n3934 19.3944
R15798 gnd.n3934 gnd.n3931 19.3944
R15799 gnd.n3931 gnd.n3930 19.3944
R15800 gnd.n3930 gnd.n3927 19.3944
R15801 gnd.n3927 gnd.n3926 19.3944
R15802 gnd.n3926 gnd.n3923 19.3944
R15803 gnd.n3923 gnd.n3922 19.3944
R15804 gnd.n3919 gnd.n3918 19.3944
R15805 gnd.n3918 gnd.n3874 19.3944
R15806 gnd.n3969 gnd.n3874 19.3944
R15807 gnd.n4672 gnd.n4671 19.3944
R15808 gnd.n4671 gnd.n4668 19.3944
R15809 gnd.n4668 gnd.n4667 19.3944
R15810 gnd.n4717 gnd.n4716 19.3944
R15811 gnd.n4716 gnd.n4715 19.3944
R15812 gnd.n4715 gnd.n4712 19.3944
R15813 gnd.n4712 gnd.n4711 19.3944
R15814 gnd.n4711 gnd.n4708 19.3944
R15815 gnd.n4708 gnd.n4707 19.3944
R15816 gnd.n4707 gnd.n4704 19.3944
R15817 gnd.n4704 gnd.n4703 19.3944
R15818 gnd.n4703 gnd.n4700 19.3944
R15819 gnd.n4700 gnd.n4699 19.3944
R15820 gnd.n4699 gnd.n4696 19.3944
R15821 gnd.n4696 gnd.n4695 19.3944
R15822 gnd.n4695 gnd.n4692 19.3944
R15823 gnd.n4692 gnd.n4691 19.3944
R15824 gnd.n4691 gnd.n4688 19.3944
R15825 gnd.n4688 gnd.n4687 19.3944
R15826 gnd.n4687 gnd.n4684 19.3944
R15827 gnd.n4684 gnd.n4683 19.3944
R15828 gnd.n4683 gnd.n4680 19.3944
R15829 gnd.n4680 gnd.n4679 19.3944
R15830 gnd.n4679 gnd.n4676 19.3944
R15831 gnd.n4676 gnd.n4675 19.3944
R15832 gnd.n4062 gnd.n3771 19.3944
R15833 gnd.n4072 gnd.n3771 19.3944
R15834 gnd.n4073 gnd.n4072 19.3944
R15835 gnd.n4073 gnd.n3752 19.3944
R15836 gnd.n4093 gnd.n3752 19.3944
R15837 gnd.n4093 gnd.n3744 19.3944
R15838 gnd.n4103 gnd.n3744 19.3944
R15839 gnd.n4104 gnd.n4103 19.3944
R15840 gnd.n4105 gnd.n4104 19.3944
R15841 gnd.n4105 gnd.n3727 19.3944
R15842 gnd.n3727 gnd.n3725 19.3944
R15843 gnd.n4131 gnd.n3725 19.3944
R15844 gnd.n4131 gnd.n3707 19.3944
R15845 gnd.n4165 gnd.n3707 19.3944
R15846 gnd.n4165 gnd.n4164 19.3944
R15847 gnd.n4164 gnd.n4163 19.3944
R15848 gnd.n4163 gnd.n4158 19.3944
R15849 gnd.n4158 gnd.n3528 19.3944
R15850 gnd.n4197 gnd.n3528 19.3944
R15851 gnd.n4198 gnd.n4197 19.3944
R15852 gnd.n4198 gnd.n3512 19.3944
R15853 gnd.n4218 gnd.n3512 19.3944
R15854 gnd.n4218 gnd.n3505 19.3944
R15855 gnd.n4228 gnd.n3505 19.3944
R15856 gnd.n4229 gnd.n4228 19.3944
R15857 gnd.n4229 gnd.n3487 19.3944
R15858 gnd.n4249 gnd.n3487 19.3944
R15859 gnd.n4249 gnd.n3479 19.3944
R15860 gnd.n4259 gnd.n3479 19.3944
R15861 gnd.n4260 gnd.n4259 19.3944
R15862 gnd.n4260 gnd.n3460 19.3944
R15863 gnd.n4280 gnd.n3460 19.3944
R15864 gnd.n4280 gnd.n3453 19.3944
R15865 gnd.n4290 gnd.n3453 19.3944
R15866 gnd.n4291 gnd.n4290 19.3944
R15867 gnd.n4291 gnd.n3436 19.3944
R15868 gnd.n4311 gnd.n3436 19.3944
R15869 gnd.n4311 gnd.n3429 19.3944
R15870 gnd.n4321 gnd.n3429 19.3944
R15871 gnd.n4322 gnd.n4321 19.3944
R15872 gnd.n4322 gnd.n3410 19.3944
R15873 gnd.n4342 gnd.n3410 19.3944
R15874 gnd.n4342 gnd.n3403 19.3944
R15875 gnd.n4352 gnd.n3403 19.3944
R15876 gnd.n4353 gnd.n4352 19.3944
R15877 gnd.n4353 gnd.n3385 19.3944
R15878 gnd.n4373 gnd.n3385 19.3944
R15879 gnd.n4373 gnd.n3377 19.3944
R15880 gnd.n4639 gnd.n3377 19.3944
R15881 gnd.n4640 gnd.n4639 19.3944
R15882 gnd.n4640 gnd.n3359 19.3944
R15883 gnd.n4659 gnd.n3359 19.3944
R15884 gnd.n4659 gnd.n3360 19.3944
R15885 gnd.n4053 gnd.n4052 19.3944
R15886 gnd.n4052 gnd.n3785 19.3944
R15887 gnd.n3808 gnd.n3785 19.3944
R15888 gnd.n3811 gnd.n3808 19.3944
R15889 gnd.n3811 gnd.n3804 19.3944
R15890 gnd.n3815 gnd.n3804 19.3944
R15891 gnd.n3818 gnd.n3815 19.3944
R15892 gnd.n3821 gnd.n3818 19.3944
R15893 gnd.n3821 gnd.n3802 19.3944
R15894 gnd.n3825 gnd.n3802 19.3944
R15895 gnd.n3828 gnd.n3825 19.3944
R15896 gnd.n3831 gnd.n3828 19.3944
R15897 gnd.n3831 gnd.n3800 19.3944
R15898 gnd.n3835 gnd.n3800 19.3944
R15899 gnd.n4058 gnd.n4057 19.3944
R15900 gnd.n4057 gnd.n3761 19.3944
R15901 gnd.n4083 gnd.n3761 19.3944
R15902 gnd.n4083 gnd.n3759 19.3944
R15903 gnd.n4089 gnd.n3759 19.3944
R15904 gnd.n4089 gnd.n4088 19.3944
R15905 gnd.n4088 gnd.n3733 19.3944
R15906 gnd.n4113 gnd.n3733 19.3944
R15907 gnd.n4113 gnd.n3731 19.3944
R15908 gnd.n4125 gnd.n3731 19.3944
R15909 gnd.n4125 gnd.n4124 19.3944
R15910 gnd.n4124 gnd.n4123 19.3944
R15911 gnd.n4123 gnd.n4121 19.3944
R15912 gnd.n4121 gnd.n3703 19.3944
R15913 gnd.n3703 gnd.n3701 19.3944
R15914 gnd.n4172 gnd.n3701 19.3944
R15915 gnd.n4172 gnd.n3699 19.3944
R15916 gnd.n4176 gnd.n3699 19.3944
R15917 gnd.n4176 gnd.n3519 19.3944
R15918 gnd.n4208 gnd.n3519 19.3944
R15919 gnd.n4208 gnd.n3517 19.3944
R15920 gnd.n4214 gnd.n3517 19.3944
R15921 gnd.n4214 gnd.n4213 19.3944
R15922 gnd.n4213 gnd.n3495 19.3944
R15923 gnd.n4239 gnd.n3495 19.3944
R15924 gnd.n4239 gnd.n3493 19.3944
R15925 gnd.n4245 gnd.n3493 19.3944
R15926 gnd.n4245 gnd.n4244 19.3944
R15927 gnd.n4244 gnd.n3469 19.3944
R15928 gnd.n4270 gnd.n3469 19.3944
R15929 gnd.n4270 gnd.n3467 19.3944
R15930 gnd.n4276 gnd.n3467 19.3944
R15931 gnd.n4276 gnd.n4275 19.3944
R15932 gnd.n4275 gnd.n3444 19.3944
R15933 gnd.n4301 gnd.n3444 19.3944
R15934 gnd.n4301 gnd.n3442 19.3944
R15935 gnd.n4307 gnd.n3442 19.3944
R15936 gnd.n4307 gnd.n4306 19.3944
R15937 gnd.n4306 gnd.n3419 19.3944
R15938 gnd.n4332 gnd.n3419 19.3944
R15939 gnd.n4332 gnd.n3417 19.3944
R15940 gnd.n4338 gnd.n3417 19.3944
R15941 gnd.n4338 gnd.n4337 19.3944
R15942 gnd.n4337 gnd.n3393 19.3944
R15943 gnd.n4363 gnd.n3393 19.3944
R15944 gnd.n4363 gnd.n3391 19.3944
R15945 gnd.n4369 gnd.n3391 19.3944
R15946 gnd.n4369 gnd.n4368 19.3944
R15947 gnd.n4368 gnd.n3368 19.3944
R15948 gnd.n4649 gnd.n3368 19.3944
R15949 gnd.n4649 gnd.n3366 19.3944
R15950 gnd.n4655 gnd.n3366 19.3944
R15951 gnd.n4655 gnd.n4654 19.3944
R15952 gnd.n4753 gnd.n4752 19.3944
R15953 gnd.n4752 gnd.n2014 19.3944
R15954 gnd.n4748 gnd.n2014 19.3944
R15955 gnd.n4748 gnd.n4745 19.3944
R15956 gnd.n4745 gnd.n4742 19.3944
R15957 gnd.n4742 gnd.n4741 19.3944
R15958 gnd.n4741 gnd.n4738 19.3944
R15959 gnd.n4738 gnd.n4737 19.3944
R15960 gnd.n4737 gnd.n4734 19.3944
R15961 gnd.n4734 gnd.n4733 19.3944
R15962 gnd.n4733 gnd.n4730 19.3944
R15963 gnd.n4730 gnd.n4729 19.3944
R15964 gnd.n4729 gnd.n4726 19.3944
R15965 gnd.n4726 gnd.n4725 19.3944
R15966 gnd.n3973 gnd.n3872 19.3944
R15967 gnd.n3973 gnd.n3863 19.3944
R15968 gnd.n3986 gnd.n3863 19.3944
R15969 gnd.n3986 gnd.n3861 19.3944
R15970 gnd.n3990 gnd.n3861 19.3944
R15971 gnd.n3990 gnd.n3851 19.3944
R15972 gnd.n4002 gnd.n3851 19.3944
R15973 gnd.n4002 gnd.n3849 19.3944
R15974 gnd.n4036 gnd.n3849 19.3944
R15975 gnd.n4036 gnd.n4035 19.3944
R15976 gnd.n4035 gnd.n4034 19.3944
R15977 gnd.n4034 gnd.n4033 19.3944
R15978 gnd.n4033 gnd.n4030 19.3944
R15979 gnd.n4030 gnd.n4029 19.3944
R15980 gnd.n4029 gnd.n4028 19.3944
R15981 gnd.n4028 gnd.n4026 19.3944
R15982 gnd.n4026 gnd.n4025 19.3944
R15983 gnd.n4025 gnd.n4022 19.3944
R15984 gnd.n4022 gnd.n4021 19.3944
R15985 gnd.n4021 gnd.n4020 19.3944
R15986 gnd.n4020 gnd.n4018 19.3944
R15987 gnd.n4018 gnd.n3716 19.3944
R15988 gnd.n4139 gnd.n3716 19.3944
R15989 gnd.n4139 gnd.n3714 19.3944
R15990 gnd.n4145 gnd.n3714 19.3944
R15991 gnd.n4145 gnd.n4144 19.3944
R15992 gnd.n4144 gnd.n3679 19.3944
R15993 gnd.n4187 gnd.n3679 19.3944
R15994 gnd.n4187 gnd.n3680 19.3944
R15995 gnd.n3696 gnd.n3695 19.3944
R15996 gnd.n4192 gnd.n4191 19.3944
R15997 gnd.n3615 gnd.n3534 19.3944
R15998 gnd.n3610 gnd.n3609 19.3944
R15999 gnd.n3609 gnd.n3607 19.3944
R16000 gnd.n3607 gnd.n3606 19.3944
R16001 gnd.n3606 gnd.n3603 19.3944
R16002 gnd.n3603 gnd.n3602 19.3944
R16003 gnd.n3602 gnd.n3601 19.3944
R16004 gnd.n3601 gnd.n3599 19.3944
R16005 gnd.n3599 gnd.n3598 19.3944
R16006 gnd.n3598 gnd.n3595 19.3944
R16007 gnd.n3595 gnd.n3594 19.3944
R16008 gnd.n3594 gnd.n3593 19.3944
R16009 gnd.n3593 gnd.n3591 19.3944
R16010 gnd.n3591 gnd.n3590 19.3944
R16011 gnd.n3590 gnd.n3585 19.3944
R16012 gnd.n3585 gnd.n3584 19.3944
R16013 gnd.n3584 gnd.n3583 19.3944
R16014 gnd.n3583 gnd.n3581 19.3944
R16015 gnd.n3581 gnd.n3580 19.3944
R16016 gnd.n3580 gnd.n3577 19.3944
R16017 gnd.n3577 gnd.n3576 19.3944
R16018 gnd.n3576 gnd.n3575 19.3944
R16019 gnd.n3575 gnd.n3573 19.3944
R16020 gnd.n3573 gnd.n3572 19.3944
R16021 gnd.n3572 gnd.n3569 19.3944
R16022 gnd.n3569 gnd.n3568 19.3944
R16023 gnd.n3568 gnd.n3567 19.3944
R16024 gnd.n3567 gnd.n3565 19.3944
R16025 gnd.n3565 gnd.n3564 19.3944
R16026 gnd.n3564 gnd.n2061 19.3944
R16027 gnd.n3978 gnd.n3868 19.3944
R16028 gnd.n3978 gnd.n3866 19.3944
R16029 gnd.n3982 gnd.n3866 19.3944
R16030 gnd.n3982 gnd.n3857 19.3944
R16031 gnd.n3994 gnd.n3857 19.3944
R16032 gnd.n3994 gnd.n3855 19.3944
R16033 gnd.n3998 gnd.n3855 19.3944
R16034 gnd.n3998 gnd.n3844 19.3944
R16035 gnd.n4040 gnd.n3844 19.3944
R16036 gnd.n4040 gnd.n3798 19.3944
R16037 gnd.n4046 gnd.n3798 19.3944
R16038 gnd.n4046 gnd.n4045 19.3944
R16039 gnd.n4045 gnd.n3776 19.3944
R16040 gnd.n4067 gnd.n3776 19.3944
R16041 gnd.n4067 gnd.n3769 19.3944
R16042 gnd.n4078 gnd.n3769 19.3944
R16043 gnd.n4078 gnd.n4077 19.3944
R16044 gnd.n4077 gnd.n3750 19.3944
R16045 gnd.n4098 gnd.n3750 19.3944
R16046 gnd.n4098 gnd.n3740 19.3944
R16047 gnd.n4108 gnd.n3740 19.3944
R16048 gnd.n4108 gnd.n3721 19.3944
R16049 gnd.n4135 gnd.n3721 19.3944
R16050 gnd.n4135 gnd.n4134 19.3944
R16051 gnd.n4134 gnd.n3709 19.3944
R16052 gnd.n4151 gnd.n3709 19.3944
R16053 gnd.n4151 gnd.n3687 19.3944
R16054 gnd.n4183 gnd.n3687 19.3944
R16055 gnd.n4183 gnd.n4182 19.3944
R16056 gnd.n4182 gnd.n4181 19.3944
R16057 gnd.n4181 gnd.n3693 19.3944
R16058 gnd.n3693 gnd.n3526 19.3944
R16059 gnd.n4203 gnd.n3526 19.3944
R16060 gnd.n4203 gnd.n4202 19.3944
R16061 gnd.n4202 gnd.n3510 19.3944
R16062 gnd.n4223 gnd.n3510 19.3944
R16063 gnd.n4223 gnd.n3503 19.3944
R16064 gnd.n4234 gnd.n3503 19.3944
R16065 gnd.n4234 gnd.n4233 19.3944
R16066 gnd.n4233 gnd.n3485 19.3944
R16067 gnd.n4254 gnd.n3485 19.3944
R16068 gnd.n4254 gnd.n3477 19.3944
R16069 gnd.n4265 gnd.n3477 19.3944
R16070 gnd.n4265 gnd.n4264 19.3944
R16071 gnd.n4264 gnd.n3458 19.3944
R16072 gnd.n4285 gnd.n3458 19.3944
R16073 gnd.n4285 gnd.n3451 19.3944
R16074 gnd.n4296 gnd.n3451 19.3944
R16075 gnd.n4296 gnd.n4295 19.3944
R16076 gnd.n4295 gnd.n3434 19.3944
R16077 gnd.n4316 gnd.n3434 19.3944
R16078 gnd.n4316 gnd.n3427 19.3944
R16079 gnd.n4327 gnd.n3427 19.3944
R16080 gnd.n4327 gnd.n4326 19.3944
R16081 gnd.n4326 gnd.n3408 19.3944
R16082 gnd.n4347 gnd.n3408 19.3944
R16083 gnd.n4347 gnd.n3401 19.3944
R16084 gnd.n4358 gnd.n3401 19.3944
R16085 gnd.n4358 gnd.n4357 19.3944
R16086 gnd.n4357 gnd.n3383 19.3944
R16087 gnd.n4634 gnd.n3383 19.3944
R16088 gnd.n4634 gnd.n3375 19.3944
R16089 gnd.n4644 gnd.n3375 19.3944
R16090 gnd.n4644 gnd.n3357 19.3944
R16091 gnd.n4662 gnd.n3357 19.3944
R16092 gnd.n6972 gnd.n565 19.3944
R16093 gnd.n6968 gnd.n565 19.3944
R16094 gnd.n6968 gnd.n6967 19.3944
R16095 gnd.n6967 gnd.n6966 19.3944
R16096 gnd.n6966 gnd.n570 19.3944
R16097 gnd.n6962 gnd.n570 19.3944
R16098 gnd.n6962 gnd.n6961 19.3944
R16099 gnd.n6961 gnd.n6960 19.3944
R16100 gnd.n6960 gnd.n574 19.3944
R16101 gnd.n6956 gnd.n574 19.3944
R16102 gnd.n6956 gnd.n6955 19.3944
R16103 gnd.n6955 gnd.n6954 19.3944
R16104 gnd.n6954 gnd.n578 19.3944
R16105 gnd.n6950 gnd.n578 19.3944
R16106 gnd.n6950 gnd.n6949 19.3944
R16107 gnd.n6949 gnd.n6948 19.3944
R16108 gnd.n6948 gnd.n582 19.3944
R16109 gnd.n6944 gnd.n582 19.3944
R16110 gnd.n6944 gnd.n6943 19.3944
R16111 gnd.n6943 gnd.n6942 19.3944
R16112 gnd.n6942 gnd.n384 19.3944
R16113 gnd.n7161 gnd.n384 19.3944
R16114 gnd.n7162 gnd.n7161 19.3944
R16115 gnd.n7162 gnd.n381 19.3944
R16116 gnd.n7167 gnd.n381 19.3944
R16117 gnd.n7167 gnd.n382 19.3944
R16118 gnd.n382 gnd.n352 19.3944
R16119 gnd.n7209 gnd.n352 19.3944
R16120 gnd.n7209 gnd.n353 19.3944
R16121 gnd.n7205 gnd.n353 19.3944
R16122 gnd.n7205 gnd.n7204 19.3944
R16123 gnd.n7204 gnd.n76 19.3944
R16124 gnd.n7624 gnd.n76 19.3944
R16125 gnd.n7624 gnd.n7623 19.3944
R16126 gnd.n7623 gnd.n7622 19.3944
R16127 gnd.n7622 gnd.n81 19.3944
R16128 gnd.n7618 gnd.n81 19.3944
R16129 gnd.n7618 gnd.n7617 19.3944
R16130 gnd.n7617 gnd.n7616 19.3944
R16131 gnd.n7616 gnd.n86 19.3944
R16132 gnd.n7612 gnd.n86 19.3944
R16133 gnd.n7612 gnd.n7611 19.3944
R16134 gnd.n7611 gnd.n7610 19.3944
R16135 gnd.n7610 gnd.n91 19.3944
R16136 gnd.n7606 gnd.n91 19.3944
R16137 gnd.n7606 gnd.n7605 19.3944
R16138 gnd.n7605 gnd.n7604 19.3944
R16139 gnd.n7604 gnd.n96 19.3944
R16140 gnd.n7600 gnd.n96 19.3944
R16141 gnd.n7600 gnd.n7599 19.3944
R16142 gnd.n7599 gnd.n7598 19.3944
R16143 gnd.n7598 gnd.n101 19.3944
R16144 gnd.n7594 gnd.n101 19.3944
R16145 gnd.n7594 gnd.n7593 19.3944
R16146 gnd.n7593 gnd.n7592 19.3944
R16147 gnd.n7592 gnd.n106 19.3944
R16148 gnd.n7588 gnd.n106 19.3944
R16149 gnd.n7588 gnd.n7587 19.3944
R16150 gnd.n7587 gnd.n7586 19.3944
R16151 gnd.n7586 gnd.n111 19.3944
R16152 gnd.n7582 gnd.n111 19.3944
R16153 gnd.n7582 gnd.n7581 19.3944
R16154 gnd.n7581 gnd.n7580 19.3944
R16155 gnd.n7580 gnd.n116 19.3944
R16156 gnd.n7474 gnd.n7473 19.3944
R16157 gnd.n7473 gnd.n7472 19.3944
R16158 gnd.n7472 gnd.n7421 19.3944
R16159 gnd.n7468 gnd.n7421 19.3944
R16160 gnd.n7468 gnd.n7467 19.3944
R16161 gnd.n7467 gnd.n7466 19.3944
R16162 gnd.n7466 gnd.n7429 19.3944
R16163 gnd.n7462 gnd.n7429 19.3944
R16164 gnd.n7462 gnd.n7461 19.3944
R16165 gnd.n7461 gnd.n7460 19.3944
R16166 gnd.n7460 gnd.n7437 19.3944
R16167 gnd.n7456 gnd.n7437 19.3944
R16168 gnd.n7456 gnd.n7455 19.3944
R16169 gnd.n7455 gnd.n7454 19.3944
R16170 gnd.n7454 gnd.n7445 19.3944
R16171 gnd.n7450 gnd.n7445 19.3944
R16172 gnd.n6623 gnd.n6622 19.3944
R16173 gnd.n6754 gnd.n6623 19.3944
R16174 gnd.n6754 gnd.n6753 19.3944
R16175 gnd.n6753 gnd.n6628 19.3944
R16176 gnd.n6746 gnd.n6628 19.3944
R16177 gnd.n6746 gnd.n6745 19.3944
R16178 gnd.n6745 gnd.n6638 19.3944
R16179 gnd.n6738 gnd.n6638 19.3944
R16180 gnd.n6738 gnd.n6737 19.3944
R16181 gnd.n6737 gnd.n6648 19.3944
R16182 gnd.n6730 gnd.n6648 19.3944
R16183 gnd.n6730 gnd.n6729 19.3944
R16184 gnd.n6729 gnd.n6658 19.3944
R16185 gnd.n6722 gnd.n6658 19.3944
R16186 gnd.n6722 gnd.n6721 19.3944
R16187 gnd.n6721 gnd.n6668 19.3944
R16188 gnd.n7057 gnd.n478 19.3944
R16189 gnd.n7057 gnd.n476 19.3944
R16190 gnd.n7061 gnd.n476 19.3944
R16191 gnd.n7061 gnd.n460 19.3944
R16192 gnd.n7073 gnd.n460 19.3944
R16193 gnd.n7073 gnd.n458 19.3944
R16194 gnd.n7077 gnd.n458 19.3944
R16195 gnd.n7077 gnd.n444 19.3944
R16196 gnd.n7089 gnd.n444 19.3944
R16197 gnd.n7089 gnd.n442 19.3944
R16198 gnd.n7093 gnd.n442 19.3944
R16199 gnd.n7093 gnd.n426 19.3944
R16200 gnd.n7105 gnd.n426 19.3944
R16201 gnd.n7105 gnd.n424 19.3944
R16202 gnd.n7109 gnd.n424 19.3944
R16203 gnd.n7109 gnd.n410 19.3944
R16204 gnd.n7121 gnd.n410 19.3944
R16205 gnd.n7121 gnd.n407 19.3944
R16206 gnd.n7128 gnd.n407 19.3944
R16207 gnd.n7128 gnd.n408 19.3944
R16208 gnd.n7124 gnd.n408 19.3944
R16209 gnd.n7124 gnd.n375 19.3944
R16210 gnd.n7179 gnd.n375 19.3944
R16211 gnd.n7179 gnd.n376 19.3944
R16212 gnd.n7175 gnd.n376 19.3944
R16213 gnd.n7175 gnd.n7174 19.3944
R16214 gnd.n7174 gnd.n7173 19.3944
R16215 gnd.n7173 gnd.n314 19.3944
R16216 gnd.n7318 gnd.n314 19.3944
R16217 gnd.n7318 gnd.n315 19.3944
R16218 gnd.n7314 gnd.n315 19.3944
R16219 gnd.n7314 gnd.n7313 19.3944
R16220 gnd.n7313 gnd.n7312 19.3944
R16221 gnd.n7312 gnd.n321 19.3944
R16222 gnd.n7308 gnd.n321 19.3944
R16223 gnd.n7308 gnd.n7307 19.3944
R16224 gnd.n7307 gnd.n293 19.3944
R16225 gnd.n7331 gnd.n293 19.3944
R16226 gnd.n7331 gnd.n291 19.3944
R16227 gnd.n7335 gnd.n291 19.3944
R16228 gnd.n7335 gnd.n277 19.3944
R16229 gnd.n7347 gnd.n277 19.3944
R16230 gnd.n7347 gnd.n275 19.3944
R16231 gnd.n7351 gnd.n275 19.3944
R16232 gnd.n7351 gnd.n263 19.3944
R16233 gnd.n7363 gnd.n263 19.3944
R16234 gnd.n7363 gnd.n261 19.3944
R16235 gnd.n7367 gnd.n261 19.3944
R16236 gnd.n7367 gnd.n247 19.3944
R16237 gnd.n7379 gnd.n247 19.3944
R16238 gnd.n7379 gnd.n245 19.3944
R16239 gnd.n7383 gnd.n245 19.3944
R16240 gnd.n7383 gnd.n232 19.3944
R16241 gnd.n7395 gnd.n232 19.3944
R16242 gnd.n7395 gnd.n230 19.3944
R16243 gnd.n7399 gnd.n230 19.3944
R16244 gnd.n7399 gnd.n217 19.3944
R16245 gnd.n7411 gnd.n217 19.3944
R16246 gnd.n7411 gnd.n214 19.3944
R16247 gnd.n7483 gnd.n214 19.3944
R16248 gnd.n7483 gnd.n215 19.3944
R16249 gnd.n7479 gnd.n215 19.3944
R16250 gnd.n7479 gnd.n7478 19.3944
R16251 gnd.n7478 gnd.n7477 19.3944
R16252 gnd.n5673 gnd.n5573 19.3944
R16253 gnd.n5673 gnd.n5672 19.3944
R16254 gnd.n5672 gnd.n5579 19.3944
R16255 gnd.n5665 gnd.n5579 19.3944
R16256 gnd.n5665 gnd.n5664 19.3944
R16257 gnd.n5664 gnd.n5591 19.3944
R16258 gnd.n5657 gnd.n5591 19.3944
R16259 gnd.n5657 gnd.n5656 19.3944
R16260 gnd.n5656 gnd.n5604 19.3944
R16261 gnd.n5649 gnd.n5604 19.3944
R16262 gnd.n5649 gnd.n5648 19.3944
R16263 gnd.n5648 gnd.n5614 19.3944
R16264 gnd.n5641 gnd.n5614 19.3944
R16265 gnd.n5641 gnd.n5640 19.3944
R16266 gnd.n5640 gnd.n5630 19.3944
R16267 gnd.n5630 gnd.n1347 19.3944
R16268 gnd.n5435 gnd.n1800 19.3944
R16269 gnd.n5435 gnd.n5434 19.3944
R16270 gnd.n5434 gnd.n5433 19.3944
R16271 gnd.n5433 gnd.n1804 19.3944
R16272 gnd.n5259 gnd.n1804 19.3944
R16273 gnd.n5259 gnd.n5257 19.3944
R16274 gnd.n5273 gnd.n5257 19.3944
R16275 gnd.n5273 gnd.n5272 19.3944
R16276 gnd.n5272 gnd.n5271 19.3944
R16277 gnd.n5271 gnd.n5268 19.3944
R16278 gnd.n5268 gnd.n5267 19.3944
R16279 gnd.n5267 gnd.n1848 19.3944
R16280 gnd.n5299 gnd.n1848 19.3944
R16281 gnd.n5299 gnd.n1846 19.3944
R16282 gnd.n5313 gnd.n1846 19.3944
R16283 gnd.n5313 gnd.n5312 19.3944
R16284 gnd.n5312 gnd.n5311 19.3944
R16285 gnd.n5311 gnd.n5308 19.3944
R16286 gnd.n5308 gnd.n5307 19.3944
R16287 gnd.n5307 gnd.n1838 19.3944
R16288 gnd.n5338 gnd.n1838 19.3944
R16289 gnd.n5338 gnd.n1836 19.3944
R16290 gnd.n5370 gnd.n1836 19.3944
R16291 gnd.n5370 gnd.n5369 19.3944
R16292 gnd.n5369 gnd.n5368 19.3944
R16293 gnd.n5368 gnd.n5344 19.3944
R16294 gnd.n5364 gnd.n5344 19.3944
R16295 gnd.n5364 gnd.n5363 19.3944
R16296 gnd.n5363 gnd.n5362 19.3944
R16297 gnd.n5362 gnd.n5350 19.3944
R16298 gnd.n5357 gnd.n5350 19.3944
R16299 gnd.n5357 gnd.n5356 19.3944
R16300 gnd.n5356 gnd.n1316 19.3944
R16301 gnd.n5811 gnd.n1316 19.3944
R16302 gnd.n5811 gnd.n1314 19.3944
R16303 gnd.n5815 gnd.n1314 19.3944
R16304 gnd.n5815 gnd.n1302 19.3944
R16305 gnd.n5827 gnd.n1302 19.3944
R16306 gnd.n5827 gnd.n1300 19.3944
R16307 gnd.n5833 gnd.n1300 19.3944
R16308 gnd.n5833 gnd.n5832 19.3944
R16309 gnd.n5832 gnd.n1260 19.3944
R16310 gnd.n5985 gnd.n1260 19.3944
R16311 gnd.n5985 gnd.n1258 19.3944
R16312 gnd.n5989 gnd.n1258 19.3944
R16313 gnd.n5989 gnd.n1245 19.3944
R16314 gnd.n6001 gnd.n1245 19.3944
R16315 gnd.n6001 gnd.n1243 19.3944
R16316 gnd.n6005 gnd.n1243 19.3944
R16317 gnd.n6005 gnd.n1229 19.3944
R16318 gnd.n6017 gnd.n1229 19.3944
R16319 gnd.n6017 gnd.n1227 19.3944
R16320 gnd.n6021 gnd.n1227 19.3944
R16321 gnd.n6021 gnd.n1214 19.3944
R16322 gnd.n6032 gnd.n1214 19.3944
R16323 gnd.n6032 gnd.n1212 19.3944
R16324 gnd.n6038 gnd.n1212 19.3944
R16325 gnd.n6038 gnd.n6037 19.3944
R16326 gnd.n6037 gnd.n1107 19.3944
R16327 gnd.n6127 gnd.n1107 19.3944
R16328 gnd.n6127 gnd.n1105 19.3944
R16329 gnd.n6131 gnd.n1105 19.3944
R16330 gnd.n6131 gnd.n1091 19.3944
R16331 gnd.n6143 gnd.n1091 19.3944
R16332 gnd.n6143 gnd.n1089 19.3944
R16333 gnd.n6147 gnd.n1089 19.3944
R16334 gnd.n6147 gnd.n1076 19.3944
R16335 gnd.n6159 gnd.n1076 19.3944
R16336 gnd.n6159 gnd.n1074 19.3944
R16337 gnd.n6163 gnd.n1074 19.3944
R16338 gnd.n6163 gnd.n1063 19.3944
R16339 gnd.n6175 gnd.n1063 19.3944
R16340 gnd.n6175 gnd.n1061 19.3944
R16341 gnd.n6181 gnd.n1061 19.3944
R16342 gnd.n6181 gnd.n6180 19.3944
R16343 gnd.n6180 gnd.n1020 19.3944
R16344 gnd.n6432 gnd.n1020 19.3944
R16345 gnd.n6432 gnd.n1018 19.3944
R16346 gnd.n6436 gnd.n1018 19.3944
R16347 gnd.n6436 gnd.n1004 19.3944
R16348 gnd.n6448 gnd.n1004 19.3944
R16349 gnd.n6448 gnd.n1002 19.3944
R16350 gnd.n6452 gnd.n1002 19.3944
R16351 gnd.n6452 gnd.n988 19.3944
R16352 gnd.n6464 gnd.n988 19.3944
R16353 gnd.n6464 gnd.n986 19.3944
R16354 gnd.n6468 gnd.n986 19.3944
R16355 gnd.n6468 gnd.n974 19.3944
R16356 gnd.n6480 gnd.n974 19.3944
R16357 gnd.n6480 gnd.n972 19.3944
R16358 gnd.n6484 gnd.n972 19.3944
R16359 gnd.n6484 gnd.n959 19.3944
R16360 gnd.n6496 gnd.n959 19.3944
R16361 gnd.n6496 gnd.n957 19.3944
R16362 gnd.n6500 gnd.n957 19.3944
R16363 gnd.n6500 gnd.n943 19.3944
R16364 gnd.n6512 gnd.n943 19.3944
R16365 gnd.n6512 gnd.n941 19.3944
R16366 gnd.n6516 gnd.n941 19.3944
R16367 gnd.n6516 gnd.n926 19.3944
R16368 gnd.n6534 gnd.n926 19.3944
R16369 gnd.n6534 gnd.n924 19.3944
R16370 gnd.n6540 gnd.n924 19.3944
R16371 gnd.n6540 gnd.n6539 19.3944
R16372 gnd.n6539 gnd.n886 19.3944
R16373 gnd.n6592 gnd.n886 19.3944
R16374 gnd.n6592 gnd.n884 19.3944
R16375 gnd.n6598 gnd.n884 19.3944
R16376 gnd.n6598 gnd.n6597 19.3944
R16377 gnd.n6597 gnd.n659 19.3944
R16378 gnd.n6783 gnd.n659 19.3944
R16379 gnd.n6783 gnd.n657 19.3944
R16380 gnd.n6787 gnd.n657 19.3944
R16381 gnd.n6787 gnd.n644 19.3944
R16382 gnd.n6800 gnd.n644 19.3944
R16383 gnd.n6800 gnd.n642 19.3944
R16384 gnd.n6806 gnd.n642 19.3944
R16385 gnd.n6806 gnd.n6805 19.3944
R16386 gnd.n6805 gnd.n614 19.3944
R16387 gnd.n6819 gnd.n614 19.3944
R16388 gnd.n6819 gnd.n612 19.3944
R16389 gnd.n6823 gnd.n612 19.3944
R16390 gnd.n6823 gnd.n610 19.3944
R16391 gnd.n6827 gnd.n610 19.3944
R16392 gnd.n6827 gnd.n608 19.3944
R16393 gnd.n6831 gnd.n608 19.3944
R16394 gnd.n6831 gnd.n606 19.3944
R16395 gnd.n6835 gnd.n606 19.3944
R16396 gnd.n6835 gnd.n604 19.3944
R16397 gnd.n6839 gnd.n604 19.3944
R16398 gnd.n6839 gnd.n602 19.3944
R16399 gnd.n6869 gnd.n602 19.3944
R16400 gnd.n6869 gnd.n600 19.3944
R16401 gnd.n6883 gnd.n600 19.3944
R16402 gnd.n6883 gnd.n6882 19.3944
R16403 gnd.n6882 gnd.n6881 19.3944
R16404 gnd.n6881 gnd.n6878 19.3944
R16405 gnd.n6878 gnd.n6877 19.3944
R16406 gnd.n6877 gnd.n592 19.3944
R16407 gnd.n6908 gnd.n592 19.3944
R16408 gnd.n6908 gnd.n590 19.3944
R16409 gnd.n6914 gnd.n590 19.3944
R16410 gnd.n6914 gnd.n6913 19.3944
R16411 gnd.n6913 gnd.n392 19.3944
R16412 gnd.n7141 gnd.n392 19.3944
R16413 gnd.n7141 gnd.n390 19.3944
R16414 gnd.n7156 gnd.n390 19.3944
R16415 gnd.n7156 gnd.n7155 19.3944
R16416 gnd.n7155 gnd.n7154 19.3944
R16417 gnd.n7154 gnd.n7151 19.3944
R16418 gnd.n7151 gnd.n7150 19.3944
R16419 gnd.n7150 gnd.n346 19.3944
R16420 gnd.n7215 gnd.n346 19.3944
R16421 gnd.n7216 gnd.n7215 19.3944
R16422 gnd.n2825 gnd.n2499 19.3944
R16423 gnd.n2825 gnd.n2500 19.3944
R16424 gnd.n2821 gnd.n2500 19.3944
R16425 gnd.n2821 gnd.n2503 19.3944
R16426 gnd.n2815 gnd.n2503 19.3944
R16427 gnd.n2815 gnd.n2814 19.3944
R16428 gnd.n2814 gnd.n2813 19.3944
R16429 gnd.n2813 gnd.n2510 19.3944
R16430 gnd.n2807 gnd.n2510 19.3944
R16431 gnd.n2807 gnd.n2806 19.3944
R16432 gnd.n2806 gnd.n2805 19.3944
R16433 gnd.n2805 gnd.n2518 19.3944
R16434 gnd.n2799 gnd.n2518 19.3944
R16435 gnd.n2799 gnd.n2798 19.3944
R16436 gnd.n2798 gnd.n2797 19.3944
R16437 gnd.n2797 gnd.n2526 19.3944
R16438 gnd.n2791 gnd.n2526 19.3944
R16439 gnd.n2791 gnd.n2790 19.3944
R16440 gnd.n2790 gnd.n2789 19.3944
R16441 gnd.n2789 gnd.n2534 19.3944
R16442 gnd.n2783 gnd.n2534 19.3944
R16443 gnd.n2783 gnd.n2782 19.3944
R16444 gnd.n2782 gnd.n2781 19.3944
R16445 gnd.n2781 gnd.n2542 19.3944
R16446 gnd.n2775 gnd.n2542 19.3944
R16447 gnd.n2775 gnd.n2774 19.3944
R16448 gnd.n2774 gnd.n2773 19.3944
R16449 gnd.n2773 gnd.n2550 19.3944
R16450 gnd.n2767 gnd.n2550 19.3944
R16451 gnd.n2767 gnd.n2766 19.3944
R16452 gnd.n2766 gnd.n2765 19.3944
R16453 gnd.n2765 gnd.n2558 19.3944
R16454 gnd.n2759 gnd.n2558 19.3944
R16455 gnd.n2759 gnd.n2758 19.3944
R16456 gnd.n2758 gnd.n2757 19.3944
R16457 gnd.n2757 gnd.n2566 19.3944
R16458 gnd.n2751 gnd.n2566 19.3944
R16459 gnd.n2751 gnd.n2750 19.3944
R16460 gnd.n2750 gnd.n2749 19.3944
R16461 gnd.n2749 gnd.n2574 19.3944
R16462 gnd.n2743 gnd.n2574 19.3944
R16463 gnd.n2743 gnd.n2742 19.3944
R16464 gnd.n2742 gnd.n2741 19.3944
R16465 gnd.n2741 gnd.n2582 19.3944
R16466 gnd.n2735 gnd.n2582 19.3944
R16467 gnd.n2735 gnd.n2734 19.3944
R16468 gnd.n2734 gnd.n2733 19.3944
R16469 gnd.n2733 gnd.n2590 19.3944
R16470 gnd.n2727 gnd.n2590 19.3944
R16471 gnd.n2727 gnd.n2726 19.3944
R16472 gnd.n2726 gnd.n2725 19.3944
R16473 gnd.n2725 gnd.n2598 19.3944
R16474 gnd.n2719 gnd.n2598 19.3944
R16475 gnd.n2719 gnd.n2718 19.3944
R16476 gnd.n2718 gnd.n2717 19.3944
R16477 gnd.n2717 gnd.n2606 19.3944
R16478 gnd.n2711 gnd.n2606 19.3944
R16479 gnd.n2711 gnd.n2710 19.3944
R16480 gnd.n2710 gnd.n2709 19.3944
R16481 gnd.n2709 gnd.n2614 19.3944
R16482 gnd.n2703 gnd.n2614 19.3944
R16483 gnd.n2703 gnd.n2702 19.3944
R16484 gnd.n2702 gnd.n2701 19.3944
R16485 gnd.n2701 gnd.n2622 19.3944
R16486 gnd.n2695 gnd.n2622 19.3944
R16487 gnd.n2695 gnd.n2694 19.3944
R16488 gnd.n2694 gnd.n2693 19.3944
R16489 gnd.n2693 gnd.n2630 19.3944
R16490 gnd.n2687 gnd.n2630 19.3944
R16491 gnd.n2687 gnd.n2686 19.3944
R16492 gnd.n2686 gnd.n2685 19.3944
R16493 gnd.n2685 gnd.n2638 19.3944
R16494 gnd.n2679 gnd.n2638 19.3944
R16495 gnd.n2679 gnd.n2678 19.3944
R16496 gnd.n2678 gnd.n2677 19.3944
R16497 gnd.n2677 gnd.n2646 19.3944
R16498 gnd.n2671 gnd.n2646 19.3944
R16499 gnd.n2671 gnd.n2670 19.3944
R16500 gnd.n2670 gnd.n2669 19.3944
R16501 gnd.n2669 gnd.n2654 19.3944
R16502 gnd.n2663 gnd.n2654 19.3944
R16503 gnd.n2663 gnd.n2662 19.3944
R16504 gnd.n2662 gnd.n344 19.3944
R16505 gnd.n7219 gnd.n344 19.3944
R16506 gnd.n3139 gnd.n2191 19.3944
R16507 gnd.n3135 gnd.n2191 19.3944
R16508 gnd.n3135 gnd.n2193 19.3944
R16509 gnd.n3129 gnd.n2193 19.3944
R16510 gnd.n3129 gnd.n3128 19.3944
R16511 gnd.n3128 gnd.n3127 19.3944
R16512 gnd.n3127 gnd.n2200 19.3944
R16513 gnd.n3121 gnd.n2200 19.3944
R16514 gnd.n3121 gnd.n3120 19.3944
R16515 gnd.n3120 gnd.n3119 19.3944
R16516 gnd.n3119 gnd.n2208 19.3944
R16517 gnd.n3113 gnd.n2208 19.3944
R16518 gnd.n3113 gnd.n3112 19.3944
R16519 gnd.n3112 gnd.n3111 19.3944
R16520 gnd.n3111 gnd.n2216 19.3944
R16521 gnd.n3105 gnd.n2216 19.3944
R16522 gnd.n3105 gnd.n3104 19.3944
R16523 gnd.n3104 gnd.n3103 19.3944
R16524 gnd.n3103 gnd.n2224 19.3944
R16525 gnd.n3097 gnd.n2224 19.3944
R16526 gnd.n3097 gnd.n3096 19.3944
R16527 gnd.n3096 gnd.n3095 19.3944
R16528 gnd.n3095 gnd.n2232 19.3944
R16529 gnd.n3089 gnd.n2232 19.3944
R16530 gnd.n3089 gnd.n3088 19.3944
R16531 gnd.n3088 gnd.n3087 19.3944
R16532 gnd.n3087 gnd.n2240 19.3944
R16533 gnd.n3081 gnd.n2240 19.3944
R16534 gnd.n3081 gnd.n3080 19.3944
R16535 gnd.n3080 gnd.n3079 19.3944
R16536 gnd.n3079 gnd.n2248 19.3944
R16537 gnd.n3073 gnd.n2248 19.3944
R16538 gnd.n3073 gnd.n3072 19.3944
R16539 gnd.n3072 gnd.n3071 19.3944
R16540 gnd.n3071 gnd.n2256 19.3944
R16541 gnd.n3065 gnd.n2256 19.3944
R16542 gnd.n3065 gnd.n3064 19.3944
R16543 gnd.n3064 gnd.n3063 19.3944
R16544 gnd.n3063 gnd.n2264 19.3944
R16545 gnd.n3057 gnd.n2264 19.3944
R16546 gnd.n3057 gnd.n3056 19.3944
R16547 gnd.n3056 gnd.n3055 19.3944
R16548 gnd.n3055 gnd.n2272 19.3944
R16549 gnd.n3049 gnd.n2272 19.3944
R16550 gnd.n3049 gnd.n3048 19.3944
R16551 gnd.n3048 gnd.n3047 19.3944
R16552 gnd.n3047 gnd.n2280 19.3944
R16553 gnd.n3041 gnd.n2280 19.3944
R16554 gnd.n3041 gnd.n3040 19.3944
R16555 gnd.n3040 gnd.n3039 19.3944
R16556 gnd.n3039 gnd.n2288 19.3944
R16557 gnd.n3033 gnd.n2288 19.3944
R16558 gnd.n3033 gnd.n3032 19.3944
R16559 gnd.n3032 gnd.n3031 19.3944
R16560 gnd.n3031 gnd.n2296 19.3944
R16561 gnd.n3025 gnd.n2296 19.3944
R16562 gnd.n3025 gnd.n3024 19.3944
R16563 gnd.n3024 gnd.n3023 19.3944
R16564 gnd.n3023 gnd.n2304 19.3944
R16565 gnd.n3017 gnd.n2304 19.3944
R16566 gnd.n3017 gnd.n3016 19.3944
R16567 gnd.n3016 gnd.n3015 19.3944
R16568 gnd.n3015 gnd.n2312 19.3944
R16569 gnd.n3009 gnd.n2312 19.3944
R16570 gnd.n3009 gnd.n3008 19.3944
R16571 gnd.n3008 gnd.n3007 19.3944
R16572 gnd.n3007 gnd.n2320 19.3944
R16573 gnd.n3001 gnd.n2320 19.3944
R16574 gnd.n3001 gnd.n3000 19.3944
R16575 gnd.n3000 gnd.n2999 19.3944
R16576 gnd.n2999 gnd.n2328 19.3944
R16577 gnd.n2993 gnd.n2328 19.3944
R16578 gnd.n2993 gnd.n2992 19.3944
R16579 gnd.n2992 gnd.n2991 19.3944
R16580 gnd.n2991 gnd.n2336 19.3944
R16581 gnd.n2985 gnd.n2336 19.3944
R16582 gnd.n2985 gnd.n2984 19.3944
R16583 gnd.n2984 gnd.n2983 19.3944
R16584 gnd.n2983 gnd.n2344 19.3944
R16585 gnd.n2977 gnd.n2344 19.3944
R16586 gnd.n2977 gnd.n2976 19.3944
R16587 gnd.n2976 gnd.n2975 19.3944
R16588 gnd.n2975 gnd.n2352 19.3944
R16589 gnd.n2969 gnd.n2352 19.3944
R16590 gnd.n2969 gnd.n2968 19.3944
R16591 gnd.n2968 gnd.n2967 19.3944
R16592 gnd.n2967 gnd.n2360 19.3944
R16593 gnd.n2961 gnd.n2360 19.3944
R16594 gnd.n2961 gnd.n2960 19.3944
R16595 gnd.n2960 gnd.n2959 19.3944
R16596 gnd.n2959 gnd.n2368 19.3944
R16597 gnd.n2953 gnd.n2368 19.3944
R16598 gnd.n2953 gnd.n2952 19.3944
R16599 gnd.n2952 gnd.n2951 19.3944
R16600 gnd.n2951 gnd.n2376 19.3944
R16601 gnd.n2945 gnd.n2376 19.3944
R16602 gnd.n2945 gnd.n2944 19.3944
R16603 gnd.n2944 gnd.n2943 19.3944
R16604 gnd.n2943 gnd.n2384 19.3944
R16605 gnd.n2937 gnd.n2384 19.3944
R16606 gnd.n2937 gnd.n2936 19.3944
R16607 gnd.n2936 gnd.n2935 19.3944
R16608 gnd.n2935 gnd.n2392 19.3944
R16609 gnd.n2929 gnd.n2392 19.3944
R16610 gnd.n2929 gnd.n2928 19.3944
R16611 gnd.n2928 gnd.n2927 19.3944
R16612 gnd.n2927 gnd.n2400 19.3944
R16613 gnd.n2921 gnd.n2400 19.3944
R16614 gnd.n2921 gnd.n2920 19.3944
R16615 gnd.n2920 gnd.n2919 19.3944
R16616 gnd.n2919 gnd.n2408 19.3944
R16617 gnd.n2913 gnd.n2408 19.3944
R16618 gnd.n2913 gnd.n2912 19.3944
R16619 gnd.n2912 gnd.n2911 19.3944
R16620 gnd.n2911 gnd.n2416 19.3944
R16621 gnd.n2905 gnd.n2416 19.3944
R16622 gnd.n2905 gnd.n2904 19.3944
R16623 gnd.n2904 gnd.n2903 19.3944
R16624 gnd.n2903 gnd.n2424 19.3944
R16625 gnd.n2897 gnd.n2424 19.3944
R16626 gnd.n2897 gnd.n2896 19.3944
R16627 gnd.n2896 gnd.n2895 19.3944
R16628 gnd.n2895 gnd.n2432 19.3944
R16629 gnd.n2889 gnd.n2432 19.3944
R16630 gnd.n2889 gnd.n2888 19.3944
R16631 gnd.n2888 gnd.n2887 19.3944
R16632 gnd.n2887 gnd.n2440 19.3944
R16633 gnd.n2881 gnd.n2440 19.3944
R16634 gnd.n2881 gnd.n2880 19.3944
R16635 gnd.n2880 gnd.n2879 19.3944
R16636 gnd.n2879 gnd.n2448 19.3944
R16637 gnd.n2873 gnd.n2448 19.3944
R16638 gnd.n2873 gnd.n2872 19.3944
R16639 gnd.n2872 gnd.n2871 19.3944
R16640 gnd.n2871 gnd.n2456 19.3944
R16641 gnd.n2865 gnd.n2456 19.3944
R16642 gnd.n2865 gnd.n2864 19.3944
R16643 gnd.n2864 gnd.n2863 19.3944
R16644 gnd.n2863 gnd.n2464 19.3944
R16645 gnd.n2857 gnd.n2464 19.3944
R16646 gnd.n2857 gnd.n2856 19.3944
R16647 gnd.n2856 gnd.n2855 19.3944
R16648 gnd.n2855 gnd.n2472 19.3944
R16649 gnd.n2849 gnd.n2472 19.3944
R16650 gnd.n2849 gnd.n2848 19.3944
R16651 gnd.n2848 gnd.n2847 19.3944
R16652 gnd.n2847 gnd.n2480 19.3944
R16653 gnd.n2841 gnd.n2480 19.3944
R16654 gnd.n2841 gnd.n2840 19.3944
R16655 gnd.n2840 gnd.n2839 19.3944
R16656 gnd.n2839 gnd.n2488 19.3944
R16657 gnd.n2833 gnd.n2488 19.3944
R16658 gnd.n2833 gnd.n2832 19.3944
R16659 gnd.n2832 gnd.n2831 19.3944
R16660 gnd.n7049 gnd.n487 19.3944
R16661 gnd.n7044 gnd.n487 19.3944
R16662 gnd.n7044 gnd.n7043 19.3944
R16663 gnd.n7043 gnd.n7042 19.3944
R16664 gnd.n7042 gnd.n7039 19.3944
R16665 gnd.n7039 gnd.n7038 19.3944
R16666 gnd.n7038 gnd.n7035 19.3944
R16667 gnd.n7035 gnd.n7034 19.3944
R16668 gnd.n7034 gnd.n7031 19.3944
R16669 gnd.n7031 gnd.n7030 19.3944
R16670 gnd.n7030 gnd.n7027 19.3944
R16671 gnd.n7027 gnd.n7026 19.3944
R16672 gnd.n7026 gnd.n7023 19.3944
R16673 gnd.n7023 gnd.n7022 19.3944
R16674 gnd.n7022 gnd.n7019 19.3944
R16675 gnd.n7017 gnd.n7014 19.3944
R16676 gnd.n7014 gnd.n7013 19.3944
R16677 gnd.n7013 gnd.n7010 19.3944
R16678 gnd.n7010 gnd.n7009 19.3944
R16679 gnd.n7009 gnd.n7006 19.3944
R16680 gnd.n7006 gnd.n7005 19.3944
R16681 gnd.n7005 gnd.n7002 19.3944
R16682 gnd.n7002 gnd.n7001 19.3944
R16683 gnd.n7001 gnd.n6998 19.3944
R16684 gnd.n6998 gnd.n6997 19.3944
R16685 gnd.n6997 gnd.n6994 19.3944
R16686 gnd.n6994 gnd.n6993 19.3944
R16687 gnd.n6993 gnd.n6990 19.3944
R16688 gnd.n6990 gnd.n6989 19.3944
R16689 gnd.n6989 gnd.n6986 19.3944
R16690 gnd.n6986 gnd.n6985 19.3944
R16691 gnd.n6985 gnd.n6982 19.3944
R16692 gnd.n6982 gnd.n6981 19.3944
R16693 gnd.n6843 gnd.n563 19.3944
R16694 gnd.n6848 gnd.n6843 19.3944
R16695 gnd.n6849 gnd.n6848 19.3944
R16696 gnd.n6852 gnd.n6849 19.3944
R16697 gnd.n6852 gnd.n6841 19.3944
R16698 gnd.n6863 gnd.n6841 19.3944
R16699 gnd.n6863 gnd.n6862 19.3944
R16700 gnd.n6862 gnd.n6861 19.3944
R16701 gnd.n6861 gnd.n596 19.3944
R16702 gnd.n6888 gnd.n596 19.3944
R16703 gnd.n6889 gnd.n6888 19.3944
R16704 gnd.n6892 gnd.n6889 19.3944
R16705 gnd.n6892 gnd.n594 19.3944
R16706 gnd.n6902 gnd.n594 19.3944
R16707 gnd.n6902 gnd.n6901 19.3944
R16708 gnd.n6901 gnd.n6900 19.3944
R16709 gnd.n6900 gnd.n587 19.3944
R16710 gnd.n6919 gnd.n587 19.3944
R16711 gnd.n6919 gnd.n585 19.3944
R16712 gnd.n6936 gnd.n585 19.3944
R16713 gnd.n6936 gnd.n6935 19.3944
R16714 gnd.n6935 gnd.n6934 19.3944
R16715 gnd.n6934 gnd.n6933 19.3944
R16716 gnd.n6933 gnd.n6932 19.3944
R16717 gnd.n6932 gnd.n6929 19.3944
R16718 gnd.n6929 gnd.n357 19.3944
R16719 gnd.n7193 gnd.n357 19.3944
R16720 gnd.n7194 gnd.n7193 19.3944
R16721 gnd.n7194 gnd.n355 19.3944
R16722 gnd.n7200 gnd.n355 19.3944
R16723 gnd.n7200 gnd.n7199 19.3944
R16724 gnd.n7199 gnd.n334 19.3944
R16725 gnd.n7230 gnd.n334 19.3944
R16726 gnd.n7230 gnd.n332 19.3944
R16727 gnd.n7299 gnd.n332 19.3944
R16728 gnd.n7299 gnd.n7298 19.3944
R16729 gnd.n7298 gnd.n7297 19.3944
R16730 gnd.n7297 gnd.n7295 19.3944
R16731 gnd.n7295 gnd.n7294 19.3944
R16732 gnd.n7294 gnd.n7292 19.3944
R16733 gnd.n7292 gnd.n7291 19.3944
R16734 gnd.n7291 gnd.n7289 19.3944
R16735 gnd.n7289 gnd.n7288 19.3944
R16736 gnd.n7288 gnd.n7286 19.3944
R16737 gnd.n7286 gnd.n7285 19.3944
R16738 gnd.n7285 gnd.n7283 19.3944
R16739 gnd.n7283 gnd.n7282 19.3944
R16740 gnd.n7282 gnd.n7280 19.3944
R16741 gnd.n7280 gnd.n7279 19.3944
R16742 gnd.n7279 gnd.n7277 19.3944
R16743 gnd.n7277 gnd.n7276 19.3944
R16744 gnd.n7276 gnd.n7274 19.3944
R16745 gnd.n7274 gnd.n7273 19.3944
R16746 gnd.n7273 gnd.n7271 19.3944
R16747 gnd.n7271 gnd.n7270 19.3944
R16748 gnd.n7270 gnd.n7268 19.3944
R16749 gnd.n7268 gnd.n7267 19.3944
R16750 gnd.n7267 gnd.n7265 19.3944
R16751 gnd.n7265 gnd.n7264 19.3944
R16752 gnd.n7264 gnd.n7262 19.3944
R16753 gnd.n7262 gnd.n7261 19.3944
R16754 gnd.n7261 gnd.n200 19.3944
R16755 gnd.n7496 gnd.n200 19.3944
R16756 gnd.n7497 gnd.n7496 19.3944
R16757 gnd.n7535 gnd.n161 19.3944
R16758 gnd.n7530 gnd.n161 19.3944
R16759 gnd.n7530 gnd.n7529 19.3944
R16760 gnd.n7529 gnd.n7528 19.3944
R16761 gnd.n7528 gnd.n168 19.3944
R16762 gnd.n7523 gnd.n168 19.3944
R16763 gnd.n7523 gnd.n7522 19.3944
R16764 gnd.n7522 gnd.n7521 19.3944
R16765 gnd.n7521 gnd.n175 19.3944
R16766 gnd.n7516 gnd.n175 19.3944
R16767 gnd.n7516 gnd.n7515 19.3944
R16768 gnd.n7515 gnd.n7514 19.3944
R16769 gnd.n7514 gnd.n182 19.3944
R16770 gnd.n7509 gnd.n182 19.3944
R16771 gnd.n7509 gnd.n7508 19.3944
R16772 gnd.n7508 gnd.n7507 19.3944
R16773 gnd.n7507 gnd.n189 19.3944
R16774 gnd.n7502 gnd.n189 19.3944
R16775 gnd.n7568 gnd.n7567 19.3944
R16776 gnd.n7567 gnd.n7566 19.3944
R16777 gnd.n7566 gnd.n133 19.3944
R16778 gnd.n7561 gnd.n133 19.3944
R16779 gnd.n7561 gnd.n7560 19.3944
R16780 gnd.n7560 gnd.n7559 19.3944
R16781 gnd.n7559 gnd.n140 19.3944
R16782 gnd.n7554 gnd.n140 19.3944
R16783 gnd.n7554 gnd.n7553 19.3944
R16784 gnd.n7553 gnd.n7552 19.3944
R16785 gnd.n7552 gnd.n147 19.3944
R16786 gnd.n7547 gnd.n147 19.3944
R16787 gnd.n7547 gnd.n7546 19.3944
R16788 gnd.n7546 gnd.n7545 19.3944
R16789 gnd.n7545 gnd.n154 19.3944
R16790 gnd.n7540 gnd.n154 19.3944
R16791 gnd.n7540 gnd.n7539 19.3944
R16792 gnd.n7053 gnd.n485 19.3944
R16793 gnd.n7053 gnd.n469 19.3944
R16794 gnd.n7065 gnd.n469 19.3944
R16795 gnd.n7065 gnd.n467 19.3944
R16796 gnd.n7069 gnd.n467 19.3944
R16797 gnd.n7069 gnd.n452 19.3944
R16798 gnd.n7081 gnd.n452 19.3944
R16799 gnd.n7081 gnd.n450 19.3944
R16800 gnd.n7085 gnd.n450 19.3944
R16801 gnd.n7085 gnd.n435 19.3944
R16802 gnd.n7097 gnd.n435 19.3944
R16803 gnd.n7097 gnd.n433 19.3944
R16804 gnd.n7101 gnd.n433 19.3944
R16805 gnd.n7101 gnd.n418 19.3944
R16806 gnd.n7113 gnd.n418 19.3944
R16807 gnd.n7113 gnd.n416 19.3944
R16808 gnd.n7117 gnd.n416 19.3944
R16809 gnd.n7117 gnd.n399 19.3944
R16810 gnd.n7132 gnd.n399 19.3944
R16811 gnd.n7132 gnd.n397 19.3944
R16812 gnd.n7136 gnd.n397 19.3944
R16813 gnd.n7136 gnd.n367 19.3944
R16814 gnd.n7183 gnd.n367 19.3944
R16815 gnd.n7183 gnd.n365 19.3944
R16816 gnd.n7187 gnd.n365 19.3944
R16817 gnd.n7188 gnd.n7187 19.3944
R16818 gnd.n7188 gnd.n305 19.3944
R16819 gnd.n7323 gnd.n7322 19.3944
R16820 gnd.n338 gnd.n337 19.3944
R16821 gnd.n7226 gnd.n7225 19.3944
R16822 gnd.n328 gnd.n327 19.3944
R16823 gnd.n7303 gnd.n298 19.3944
R16824 gnd.n7327 gnd.n298 19.3944
R16825 gnd.n7327 gnd.n284 19.3944
R16826 gnd.n7339 gnd.n284 19.3944
R16827 gnd.n7339 gnd.n282 19.3944
R16828 gnd.n7343 gnd.n282 19.3944
R16829 gnd.n7343 gnd.n270 19.3944
R16830 gnd.n7355 gnd.n270 19.3944
R16831 gnd.n7355 gnd.n268 19.3944
R16832 gnd.n7359 gnd.n268 19.3944
R16833 gnd.n7359 gnd.n254 19.3944
R16834 gnd.n7371 gnd.n254 19.3944
R16835 gnd.n7371 gnd.n252 19.3944
R16836 gnd.n7375 gnd.n252 19.3944
R16837 gnd.n7375 gnd.n240 19.3944
R16838 gnd.n7387 gnd.n240 19.3944
R16839 gnd.n7387 gnd.n238 19.3944
R16840 gnd.n7391 gnd.n238 19.3944
R16841 gnd.n7391 gnd.n223 19.3944
R16842 gnd.n7403 gnd.n223 19.3944
R16843 gnd.n7403 gnd.n221 19.3944
R16844 gnd.n7407 gnd.n221 19.3944
R16845 gnd.n7407 gnd.n207 19.3944
R16846 gnd.n7487 gnd.n207 19.3944
R16847 gnd.n7487 gnd.n205 19.3944
R16848 gnd.n7491 gnd.n205 19.3944
R16849 gnd.n7491 gnd.n128 19.3944
R16850 gnd.n7571 gnd.n128 19.3944
R16851 gnd.n5065 gnd.n5064 19.3944
R16852 gnd.n5064 gnd.n4875 19.3944
R16853 gnd.n5059 gnd.n4875 19.3944
R16854 gnd.n5059 gnd.n5058 19.3944
R16855 gnd.n5058 gnd.n4880 19.3944
R16856 gnd.n5053 gnd.n4880 19.3944
R16857 gnd.n5053 gnd.n5052 19.3944
R16858 gnd.n5052 gnd.n5051 19.3944
R16859 gnd.n5051 gnd.n4886 19.3944
R16860 gnd.n5045 gnd.n4886 19.3944
R16861 gnd.n5045 gnd.n5044 19.3944
R16862 gnd.n5044 gnd.n5043 19.3944
R16863 gnd.n5043 gnd.n4892 19.3944
R16864 gnd.n5037 gnd.n4892 19.3944
R16865 gnd.n5037 gnd.n5036 19.3944
R16866 gnd.n5036 gnd.n5035 19.3944
R16867 gnd.n5035 gnd.n4898 19.3944
R16868 gnd.n5029 gnd.n5028 19.3944
R16869 gnd.n5028 gnd.n5027 19.3944
R16870 gnd.n5027 gnd.n4907 19.3944
R16871 gnd.n5021 gnd.n4907 19.3944
R16872 gnd.n5021 gnd.n5020 19.3944
R16873 gnd.n5020 gnd.n5019 19.3944
R16874 gnd.n5019 gnd.n4913 19.3944
R16875 gnd.n5013 gnd.n4913 19.3944
R16876 gnd.n5013 gnd.n5012 19.3944
R16877 gnd.n5012 gnd.n5011 19.3944
R16878 gnd.n5011 gnd.n4919 19.3944
R16879 gnd.n5005 gnd.n4919 19.3944
R16880 gnd.n5005 gnd.n5004 19.3944
R16881 gnd.n5004 gnd.n5003 19.3944
R16882 gnd.n5003 gnd.n4925 19.3944
R16883 gnd.n4997 gnd.n4925 19.3944
R16884 gnd.n4997 gnd.n4996 19.3944
R16885 gnd.n4996 gnd.n4995 19.3944
R16886 gnd.n5072 gnd.n1985 19.3944
R16887 gnd.n5076 gnd.n1985 19.3944
R16888 gnd.n5076 gnd.n1972 19.3944
R16889 gnd.n5088 gnd.n1972 19.3944
R16890 gnd.n5088 gnd.n1970 19.3944
R16891 gnd.n5092 gnd.n1970 19.3944
R16892 gnd.n5092 gnd.n1955 19.3944
R16893 gnd.n5104 gnd.n1955 19.3944
R16894 gnd.n5104 gnd.n1953 19.3944
R16895 gnd.n5108 gnd.n1953 19.3944
R16896 gnd.n5108 gnd.n1940 19.3944
R16897 gnd.n5120 gnd.n1940 19.3944
R16898 gnd.n5120 gnd.n1938 19.3944
R16899 gnd.n5124 gnd.n1938 19.3944
R16900 gnd.n5124 gnd.n1923 19.3944
R16901 gnd.n5136 gnd.n1923 19.3944
R16902 gnd.n5136 gnd.n1921 19.3944
R16903 gnd.n5148 gnd.n1921 19.3944
R16904 gnd.n5148 gnd.n5147 19.3944
R16905 gnd.n5147 gnd.n5146 19.3944
R16906 gnd.n5146 gnd.n5145 19.3944
R16907 gnd.n5145 gnd.n1887 19.3944
R16908 gnd.n5188 gnd.n1887 19.3944
R16909 gnd.n5188 gnd.n5187 19.3944
R16910 gnd.n5187 gnd.n5186 19.3944
R16911 gnd.n5186 gnd.n1896 19.3944
R16912 gnd.n1896 gnd.n1895 19.3944
R16913 gnd.n1895 gnd.n1778 19.3944
R16914 gnd.n5459 gnd.n1778 19.3944
R16915 gnd.n5459 gnd.n5458 19.3944
R16916 gnd.n5458 gnd.n5457 19.3944
R16917 gnd.n5457 gnd.n1782 19.3944
R16918 gnd.n5445 gnd.n1782 19.3944
R16919 gnd.n5445 gnd.n5444 19.3944
R16920 gnd.n5444 gnd.n5443 19.3944
R16921 gnd.n5443 gnd.n1756 19.3944
R16922 gnd.n5471 gnd.n1756 19.3944
R16923 gnd.n5471 gnd.n1754 19.3944
R16924 gnd.n5475 gnd.n1754 19.3944
R16925 gnd.n5475 gnd.n1740 19.3944
R16926 gnd.n5487 gnd.n1740 19.3944
R16927 gnd.n5487 gnd.n1738 19.3944
R16928 gnd.n5491 gnd.n1738 19.3944
R16929 gnd.n5491 gnd.n1722 19.3944
R16930 gnd.n5503 gnd.n1722 19.3944
R16931 gnd.n5503 gnd.n1720 19.3944
R16932 gnd.n5507 gnd.n1720 19.3944
R16933 gnd.n5507 gnd.n1706 19.3944
R16934 gnd.n5519 gnd.n1706 19.3944
R16935 gnd.n5519 gnd.n1704 19.3944
R16936 gnd.n5523 gnd.n1704 19.3944
R16937 gnd.n5523 gnd.n1688 19.3944
R16938 gnd.n5535 gnd.n1688 19.3944
R16939 gnd.n5535 gnd.n1686 19.3944
R16940 gnd.n5539 gnd.n1686 19.3944
R16941 gnd.n5539 gnd.n1672 19.3944
R16942 gnd.n5551 gnd.n1672 19.3944
R16943 gnd.n5551 gnd.n1670 19.3944
R16944 gnd.n5555 gnd.n1670 19.3944
R16945 gnd.n5555 gnd.n1653 19.3944
R16946 gnd.n5569 gnd.n1653 19.3944
R16947 gnd.n5569 gnd.n1651 19.3944
R16948 gnd.n5692 gnd.n1651 19.3944
R16949 gnd.n5692 gnd.n5691 19.3944
R16950 gnd.n4780 gnd.n4779 19.3944
R16951 gnd.n4785 gnd.n4780 19.3944
R16952 gnd.n4785 gnd.n4777 19.3944
R16953 gnd.n4789 gnd.n4777 19.3944
R16954 gnd.n4789 gnd.n4775 19.3944
R16955 gnd.n4795 gnd.n4775 19.3944
R16956 gnd.n4795 gnd.n4773 19.3944
R16957 gnd.n4799 gnd.n4773 19.3944
R16958 gnd.n4799 gnd.n4771 19.3944
R16959 gnd.n4805 gnd.n4771 19.3944
R16960 gnd.n4805 gnd.n4769 19.3944
R16961 gnd.n4809 gnd.n4769 19.3944
R16962 gnd.n4809 gnd.n4767 19.3944
R16963 gnd.n4815 gnd.n4767 19.3944
R16964 gnd.n4815 gnd.n4765 19.3944
R16965 gnd.n4819 gnd.n4765 19.3944
R16966 gnd.n4870 gnd.n4759 19.3944
R16967 gnd.n4870 gnd.n4869 19.3944
R16968 gnd.n4869 gnd.n4868 19.3944
R16969 gnd.n4868 gnd.n4866 19.3944
R16970 gnd.n4866 gnd.n4865 19.3944
R16971 gnd.n4865 gnd.n4863 19.3944
R16972 gnd.n4863 gnd.n4862 19.3944
R16973 gnd.n4862 gnd.n4860 19.3944
R16974 gnd.n4860 gnd.n4859 19.3944
R16975 gnd.n4859 gnd.n4857 19.3944
R16976 gnd.n4857 gnd.n4856 19.3944
R16977 gnd.n4856 gnd.n4854 19.3944
R16978 gnd.n4854 gnd.n4853 19.3944
R16979 gnd.n4853 gnd.n4851 19.3944
R16980 gnd.n4851 gnd.n4850 19.3944
R16981 gnd.n4850 gnd.n4848 19.3944
R16982 gnd.n4848 gnd.n4847 19.3944
R16983 gnd.n4847 gnd.n4845 19.3944
R16984 gnd.n4845 gnd.n1906 19.3944
R16985 gnd.n5162 gnd.n1906 19.3944
R16986 gnd.n5162 gnd.n1904 19.3944
R16987 gnd.n5171 gnd.n1904 19.3944
R16988 gnd.n5171 gnd.n5170 19.3944
R16989 gnd.n5170 gnd.n5169 19.3944
R16990 gnd.n5169 gnd.n1871 19.3944
R16991 gnd.n5201 gnd.n1871 19.3944
R16992 gnd.n5201 gnd.n1869 19.3944
R16993 gnd.n5215 gnd.n1869 19.3944
R16994 gnd.n5215 gnd.n5214 19.3944
R16995 gnd.n5214 gnd.n5213 19.3944
R16996 gnd.n5213 gnd.n5211 19.3944
R16997 gnd.n5211 gnd.n5210 19.3944
R16998 gnd.n5210 gnd.n1859 19.3944
R16999 gnd.n5235 gnd.n1859 19.3944
R17000 gnd.n5235 gnd.n1857 19.3944
R17001 gnd.n5239 gnd.n1857 19.3944
R17002 gnd.n5239 gnd.n1807 19.3944
R17003 gnd.n5427 gnd.n1807 19.3944
R17004 gnd.n5427 gnd.n1808 19.3944
R17005 gnd.n5423 gnd.n1808 19.3944
R17006 gnd.n5423 gnd.n5422 19.3944
R17007 gnd.n5422 gnd.n5421 19.3944
R17008 gnd.n5421 gnd.n1813 19.3944
R17009 gnd.n5417 gnd.n1813 19.3944
R17010 gnd.n5417 gnd.n5416 19.3944
R17011 gnd.n5416 gnd.n5415 19.3944
R17012 gnd.n5415 gnd.n1817 19.3944
R17013 gnd.n5411 gnd.n1817 19.3944
R17014 gnd.n5411 gnd.n5410 19.3944
R17015 gnd.n5410 gnd.n5409 19.3944
R17016 gnd.n5409 gnd.n1821 19.3944
R17017 gnd.n5405 gnd.n1821 19.3944
R17018 gnd.n5405 gnd.n5404 19.3944
R17019 gnd.n5404 gnd.n5403 19.3944
R17020 gnd.n5403 gnd.n1825 19.3944
R17021 gnd.n5399 gnd.n1825 19.3944
R17022 gnd.n5399 gnd.n5398 19.3944
R17023 gnd.n5398 gnd.n5397 19.3944
R17024 gnd.n5397 gnd.n1829 19.3944
R17025 gnd.n5393 gnd.n1829 19.3944
R17026 gnd.n5393 gnd.n5392 19.3944
R17027 gnd.n5392 gnd.n5391 19.3944
R17028 gnd.n5391 gnd.n5388 19.3944
R17029 gnd.n5388 gnd.n1353 19.3944
R17030 gnd.n4986 gnd.n4985 19.3944
R17031 gnd.n4985 gnd.n4984 19.3944
R17032 gnd.n4984 gnd.n4983 19.3944
R17033 gnd.n4983 gnd.n4981 19.3944
R17034 gnd.n4981 gnd.n4980 19.3944
R17035 gnd.n4980 gnd.n4978 19.3944
R17036 gnd.n4978 gnd.n4977 19.3944
R17037 gnd.n4977 gnd.n4975 19.3944
R17038 gnd.n4975 gnd.n4974 19.3944
R17039 gnd.n4974 gnd.n4972 19.3944
R17040 gnd.n4972 gnd.n4971 19.3944
R17041 gnd.n4971 gnd.n4969 19.3944
R17042 gnd.n4969 gnd.n4968 19.3944
R17043 gnd.n4968 gnd.n4966 19.3944
R17044 gnd.n4966 gnd.n4965 19.3944
R17045 gnd.n4965 gnd.n4963 19.3944
R17046 gnd.n4963 gnd.n4962 19.3944
R17047 gnd.n4962 gnd.n4960 19.3944
R17048 gnd.n4960 gnd.n4959 19.3944
R17049 gnd.n4959 gnd.n4957 19.3944
R17050 gnd.n4957 gnd.n1900 19.3944
R17051 gnd.n5175 gnd.n1900 19.3944
R17052 gnd.n5176 gnd.n5175 19.3944
R17053 gnd.n5176 gnd.n1898 19.3944
R17054 gnd.n5182 gnd.n1898 19.3944
R17055 gnd.n5182 gnd.n5181 19.3944
R17056 gnd.n5181 gnd.n1865 19.3944
R17057 gnd.n5219 gnd.n1865 19.3944
R17058 gnd.n5219 gnd.n1863 19.3944
R17059 gnd.n5224 gnd.n1863 19.3944
R17060 gnd.n5225 gnd.n5224 19.3944
R17061 gnd.n5227 gnd.n5225 19.3944
R17062 gnd.n5227 gnd.n1860 19.3944
R17063 gnd.n5231 gnd.n1860 19.3944
R17064 gnd.n5231 gnd.n1856 19.3944
R17065 gnd.n5243 gnd.n1856 19.3944
R17066 gnd.n5243 gnd.n1854 19.3944
R17067 gnd.n5247 gnd.n1854 19.3944
R17068 gnd.n5248 gnd.n5247 19.3944
R17069 gnd.n5251 gnd.n5248 19.3944
R17070 gnd.n5251 gnd.n1852 19.3944
R17071 gnd.n5278 gnd.n1852 19.3944
R17072 gnd.n5279 gnd.n5278 19.3944
R17073 gnd.n5282 gnd.n5279 19.3944
R17074 gnd.n5282 gnd.n1850 19.3944
R17075 gnd.n5293 gnd.n1850 19.3944
R17076 gnd.n5293 gnd.n5292 19.3944
R17077 gnd.n5292 gnd.n5291 19.3944
R17078 gnd.n5291 gnd.n1842 19.3944
R17079 gnd.n5318 gnd.n1842 19.3944
R17080 gnd.n5319 gnd.n5318 19.3944
R17081 gnd.n5322 gnd.n5319 19.3944
R17082 gnd.n5322 gnd.n1840 19.3944
R17083 gnd.n5332 gnd.n1840 19.3944
R17084 gnd.n5332 gnd.n5331 19.3944
R17085 gnd.n5331 gnd.n5330 19.3944
R17086 gnd.n5330 gnd.n1833 19.3944
R17087 gnd.n5375 gnd.n1833 19.3944
R17088 gnd.n5375 gnd.n1831 19.3944
R17089 gnd.n5382 gnd.n1831 19.3944
R17090 gnd.n5382 gnd.n5381 19.3944
R17091 gnd.n5381 gnd.n1647 19.3944
R17092 gnd.n5696 gnd.n1647 19.3944
R17093 gnd.n5697 gnd.n5696 19.3944
R17094 gnd.n5735 gnd.n5734 19.3944
R17095 gnd.n5734 gnd.n5733 19.3944
R17096 gnd.n5733 gnd.n1613 19.3944
R17097 gnd.n5728 gnd.n1613 19.3944
R17098 gnd.n5728 gnd.n5727 19.3944
R17099 gnd.n5727 gnd.n5726 19.3944
R17100 gnd.n5726 gnd.n1620 19.3944
R17101 gnd.n5721 gnd.n1620 19.3944
R17102 gnd.n5721 gnd.n5720 19.3944
R17103 gnd.n5720 gnd.n5719 19.3944
R17104 gnd.n5719 gnd.n1627 19.3944
R17105 gnd.n5714 gnd.n1627 19.3944
R17106 gnd.n5714 gnd.n5713 19.3944
R17107 gnd.n5713 gnd.n5712 19.3944
R17108 gnd.n5712 gnd.n1634 19.3944
R17109 gnd.n5707 gnd.n1634 19.3944
R17110 gnd.n5707 gnd.n5706 19.3944
R17111 gnd.n5706 gnd.n5705 19.3944
R17112 gnd.n5766 gnd.n5765 19.3944
R17113 gnd.n5765 gnd.n1363 19.3944
R17114 gnd.n1365 gnd.n1363 19.3944
R17115 gnd.n5758 gnd.n1365 19.3944
R17116 gnd.n5758 gnd.n5757 19.3944
R17117 gnd.n5757 gnd.n5756 19.3944
R17118 gnd.n5756 gnd.n1372 19.3944
R17119 gnd.n5751 gnd.n1372 19.3944
R17120 gnd.n5751 gnd.n5750 19.3944
R17121 gnd.n5750 gnd.n5749 19.3944
R17122 gnd.n5749 gnd.n1379 19.3944
R17123 gnd.n5744 gnd.n1379 19.3944
R17124 gnd.n5744 gnd.n5743 19.3944
R17125 gnd.n5743 gnd.n5742 19.3944
R17126 gnd.n5742 gnd.n1386 19.3944
R17127 gnd.n5068 gnd.n1980 19.3944
R17128 gnd.n5080 gnd.n1980 19.3944
R17129 gnd.n5080 gnd.n1978 19.3944
R17130 gnd.n5084 gnd.n1978 19.3944
R17131 gnd.n5084 gnd.n1964 19.3944
R17132 gnd.n5096 gnd.n1964 19.3944
R17133 gnd.n5096 gnd.n1962 19.3944
R17134 gnd.n5100 gnd.n1962 19.3944
R17135 gnd.n5100 gnd.n1948 19.3944
R17136 gnd.n5112 gnd.n1948 19.3944
R17137 gnd.n5112 gnd.n1946 19.3944
R17138 gnd.n5116 gnd.n1946 19.3944
R17139 gnd.n5116 gnd.n1932 19.3944
R17140 gnd.n5128 gnd.n1932 19.3944
R17141 gnd.n5128 gnd.n1930 19.3944
R17142 gnd.n5132 gnd.n1930 19.3944
R17143 gnd.n5132 gnd.n1915 19.3944
R17144 gnd.n5152 gnd.n1915 19.3944
R17145 gnd.n5152 gnd.n1913 19.3944
R17146 gnd.n5158 gnd.n1913 19.3944
R17147 gnd.n5158 gnd.n5157 19.3944
R17148 gnd.n5157 gnd.n1879 19.3944
R17149 gnd.n5192 gnd.n1879 19.3944
R17150 gnd.n5192 gnd.n1877 19.3944
R17151 gnd.n5196 gnd.n1877 19.3944
R17152 gnd.n5197 gnd.n5196 19.3944
R17153 gnd.n5197 gnd.n1770 19.3944
R17154 gnd.n5464 gnd.n5463 19.3944
R17155 gnd.n5453 gnd.n5452 19.3944
R17156 gnd.n5450 gnd.n5449 19.3944
R17157 gnd.n5439 gnd.n5438 19.3944
R17158 gnd.n5467 gnd.n1763 19.3944
R17159 gnd.n5467 gnd.n1748 19.3944
R17160 gnd.n5479 gnd.n1748 19.3944
R17161 gnd.n5479 gnd.n1746 19.3944
R17162 gnd.n5483 gnd.n1746 19.3944
R17163 gnd.n5483 gnd.n1731 19.3944
R17164 gnd.n5495 gnd.n1731 19.3944
R17165 gnd.n5495 gnd.n1729 19.3944
R17166 gnd.n5499 gnd.n1729 19.3944
R17167 gnd.n5499 gnd.n1714 19.3944
R17168 gnd.n5511 gnd.n1714 19.3944
R17169 gnd.n5511 gnd.n1712 19.3944
R17170 gnd.n5515 gnd.n1712 19.3944
R17171 gnd.n5515 gnd.n1697 19.3944
R17172 gnd.n5527 gnd.n1697 19.3944
R17173 gnd.n5527 gnd.n1695 19.3944
R17174 gnd.n5531 gnd.n1695 19.3944
R17175 gnd.n5531 gnd.n1680 19.3944
R17176 gnd.n5543 gnd.n1680 19.3944
R17177 gnd.n5543 gnd.n1678 19.3944
R17178 gnd.n5547 gnd.n1678 19.3944
R17179 gnd.n5547 gnd.n1663 19.3944
R17180 gnd.n5559 gnd.n1663 19.3944
R17181 gnd.n5559 gnd.n1661 19.3944
R17182 gnd.n5565 gnd.n1661 19.3944
R17183 gnd.n5565 gnd.n5564 19.3944
R17184 gnd.n5564 gnd.n1360 19.3944
R17185 gnd.n5769 gnd.n1360 19.3944
R17186 gnd.n3145 gnd.n2187 19.3944
R17187 gnd.n3145 gnd.n2185 19.3944
R17188 gnd.n3149 gnd.n2185 19.3944
R17189 gnd.n3149 gnd.n2181 19.3944
R17190 gnd.n3155 gnd.n2181 19.3944
R17191 gnd.n3155 gnd.n2179 19.3944
R17192 gnd.n3159 gnd.n2179 19.3944
R17193 gnd.n3159 gnd.n2175 19.3944
R17194 gnd.n3165 gnd.n2175 19.3944
R17195 gnd.n3165 gnd.n2173 19.3944
R17196 gnd.n3169 gnd.n2173 19.3944
R17197 gnd.n3169 gnd.n2169 19.3944
R17198 gnd.n3175 gnd.n2169 19.3944
R17199 gnd.n3175 gnd.n2167 19.3944
R17200 gnd.n3179 gnd.n2167 19.3944
R17201 gnd.n3179 gnd.n2163 19.3944
R17202 gnd.n3185 gnd.n2163 19.3944
R17203 gnd.n3185 gnd.n2161 19.3944
R17204 gnd.n3189 gnd.n2161 19.3944
R17205 gnd.n3189 gnd.n2157 19.3944
R17206 gnd.n3195 gnd.n2157 19.3944
R17207 gnd.n3195 gnd.n2155 19.3944
R17208 gnd.n3199 gnd.n2155 19.3944
R17209 gnd.n3199 gnd.n2151 19.3944
R17210 gnd.n3205 gnd.n2151 19.3944
R17211 gnd.n3205 gnd.n2149 19.3944
R17212 gnd.n3209 gnd.n2149 19.3944
R17213 gnd.n3209 gnd.n2145 19.3944
R17214 gnd.n3215 gnd.n2145 19.3944
R17215 gnd.n3215 gnd.n2143 19.3944
R17216 gnd.n3219 gnd.n2143 19.3944
R17217 gnd.n3219 gnd.n2139 19.3944
R17218 gnd.n3225 gnd.n2139 19.3944
R17219 gnd.n3225 gnd.n2137 19.3944
R17220 gnd.n3229 gnd.n2137 19.3944
R17221 gnd.n3229 gnd.n2133 19.3944
R17222 gnd.n3235 gnd.n2133 19.3944
R17223 gnd.n3235 gnd.n2131 19.3944
R17224 gnd.n3239 gnd.n2131 19.3944
R17225 gnd.n3239 gnd.n2127 19.3944
R17226 gnd.n3245 gnd.n2127 19.3944
R17227 gnd.n3245 gnd.n2125 19.3944
R17228 gnd.n3249 gnd.n2125 19.3944
R17229 gnd.n3249 gnd.n2121 19.3944
R17230 gnd.n3255 gnd.n2121 19.3944
R17231 gnd.n3255 gnd.n2119 19.3944
R17232 gnd.n3259 gnd.n2119 19.3944
R17233 gnd.n3259 gnd.n2115 19.3944
R17234 gnd.n3265 gnd.n2115 19.3944
R17235 gnd.n3265 gnd.n2113 19.3944
R17236 gnd.n3269 gnd.n2113 19.3944
R17237 gnd.n3269 gnd.n2109 19.3944
R17238 gnd.n3275 gnd.n2109 19.3944
R17239 gnd.n3275 gnd.n2107 19.3944
R17240 gnd.n3279 gnd.n2107 19.3944
R17241 gnd.n3279 gnd.n2103 19.3944
R17242 gnd.n3285 gnd.n2103 19.3944
R17243 gnd.n3285 gnd.n2101 19.3944
R17244 gnd.n3289 gnd.n2101 19.3944
R17245 gnd.n3289 gnd.n2097 19.3944
R17246 gnd.n3295 gnd.n2097 19.3944
R17247 gnd.n3295 gnd.n2095 19.3944
R17248 gnd.n3299 gnd.n2095 19.3944
R17249 gnd.n3299 gnd.n2091 19.3944
R17250 gnd.n3305 gnd.n2091 19.3944
R17251 gnd.n3305 gnd.n2089 19.3944
R17252 gnd.n3309 gnd.n2089 19.3944
R17253 gnd.n3309 gnd.n2085 19.3944
R17254 gnd.n3315 gnd.n2085 19.3944
R17255 gnd.n3315 gnd.n2083 19.3944
R17256 gnd.n3319 gnd.n2083 19.3944
R17257 gnd.n3319 gnd.n2079 19.3944
R17258 gnd.n3325 gnd.n2079 19.3944
R17259 gnd.n3325 gnd.n2077 19.3944
R17260 gnd.n3329 gnd.n2077 19.3944
R17261 gnd.n3329 gnd.n2073 19.3944
R17262 gnd.n3335 gnd.n2073 19.3944
R17263 gnd.n3335 gnd.n2071 19.3944
R17264 gnd.n3339 gnd.n2071 19.3944
R17265 gnd.n3339 gnd.n2067 19.3944
R17266 gnd.n3345 gnd.n2067 19.3944
R17267 gnd.n3345 gnd.n2065 19.3944
R17268 gnd.n3352 gnd.n2065 19.3944
R17269 gnd.n3352 gnd.n3351 19.3944
R17270 gnd.n5686 gnd.n5685 19.3944
R17271 gnd.n5685 gnd.n5684 19.3944
R17272 gnd.n5684 gnd.n5679 19.3944
R17273 gnd.n5680 gnd.n5679 19.3944
R17274 gnd.n5680 gnd.n1285 19.3944
R17275 gnd.n5846 gnd.n1285 19.3944
R17276 gnd.n5846 gnd.n1281 19.3944
R17277 gnd.n5850 gnd.n1281 19.3944
R17278 gnd.n5851 gnd.n5850 19.3944
R17279 gnd.n5855 gnd.n5851 19.3944
R17280 gnd.n5855 gnd.n1278 19.3944
R17281 gnd.n5965 gnd.n1278 19.3944
R17282 gnd.n5965 gnd.n1279 19.3944
R17283 gnd.n5961 gnd.n1279 19.3944
R17284 gnd.n5961 gnd.n5960 19.3944
R17285 gnd.n5960 gnd.n5959 19.3944
R17286 gnd.n5959 gnd.n5861 19.3944
R17287 gnd.n5955 gnd.n5861 19.3944
R17288 gnd.n5955 gnd.n5954 19.3944
R17289 gnd.n5954 gnd.n5953 19.3944
R17290 gnd.n5953 gnd.n5950 19.3944
R17291 gnd.n5950 gnd.n1197 19.3944
R17292 gnd.n6051 gnd.n1197 19.3944
R17293 gnd.n6051 gnd.n1193 19.3944
R17294 gnd.n6055 gnd.n1193 19.3944
R17295 gnd.n6056 gnd.n6055 19.3944
R17296 gnd.n6058 gnd.n6056 19.3944
R17297 gnd.n6058 gnd.n1191 19.3944
R17298 gnd.n6062 gnd.n1191 19.3944
R17299 gnd.n6063 gnd.n6062 19.3944
R17300 gnd.n6065 gnd.n6063 19.3944
R17301 gnd.n6065 gnd.n1189 19.3944
R17302 gnd.n6069 gnd.n1189 19.3944
R17303 gnd.n6070 gnd.n6069 19.3944
R17304 gnd.n6072 gnd.n6070 19.3944
R17305 gnd.n6072 gnd.n1186 19.3944
R17306 gnd.n6077 gnd.n1186 19.3944
R17307 gnd.n6077 gnd.n1187 19.3944
R17308 gnd.n1187 gnd.n1047 19.3944
R17309 gnd.n6194 gnd.n1047 19.3944
R17310 gnd.n6194 gnd.n1043 19.3944
R17311 gnd.n6198 gnd.n1043 19.3944
R17312 gnd.n6199 gnd.n6198 19.3944
R17313 gnd.n6201 gnd.n6199 19.3944
R17314 gnd.n6201 gnd.n1040 19.3944
R17315 gnd.n6412 gnd.n1040 19.3944
R17316 gnd.n6412 gnd.n1041 19.3944
R17317 gnd.n6408 gnd.n1041 19.3944
R17318 gnd.n6408 gnd.n6407 19.3944
R17319 gnd.n6407 gnd.n6406 19.3944
R17320 gnd.n6406 gnd.n6207 19.3944
R17321 gnd.n6402 gnd.n6207 19.3944
R17322 gnd.n6402 gnd.n6401 19.3944
R17323 gnd.n6401 gnd.n6400 19.3944
R17324 gnd.n6400 gnd.n6211 19.3944
R17325 gnd.n6396 gnd.n6211 19.3944
R17326 gnd.n6396 gnd.n6395 19.3944
R17327 gnd.n6395 gnd.n6394 19.3944
R17328 gnd.n6394 gnd.n6215 19.3944
R17329 gnd.n6390 gnd.n6215 19.3944
R17330 gnd.n6390 gnd.n6389 19.3944
R17331 gnd.n6389 gnd.n6388 19.3944
R17332 gnd.n6388 gnd.n6219 19.3944
R17333 gnd.n6384 gnd.n6219 19.3944
R17334 gnd.n6384 gnd.n6383 19.3944
R17335 gnd.n6383 gnd.n917 19.3944
R17336 gnd.n6544 gnd.n917 19.3944
R17337 gnd.n6544 gnd.n914 19.3944
R17338 gnd.n6549 gnd.n914 19.3944
R17339 gnd.n6549 gnd.n915 19.3944
R17340 gnd.n915 gnd.n876 19.3944
R17341 gnd.n6602 gnd.n876 19.3944
R17342 gnd.n6602 gnd.n873 19.3944
R17343 gnd.n6606 gnd.n873 19.3944
R17344 gnd.n6607 gnd.n6606 19.3944
R17345 gnd.n6609 gnd.n6607 19.3944
R17346 gnd.n6609 gnd.n870 19.3944
R17347 gnd.n6766 gnd.n870 19.3944
R17348 gnd.n6766 gnd.n871 19.3944
R17349 gnd.n6762 gnd.n871 19.3944
R17350 gnd.n6762 gnd.n6761 19.3944
R17351 gnd.n6761 gnd.n6760 19.3944
R17352 gnd.n6695 gnd.n6694 19.3944
R17353 gnd.n6694 gnd.n633 19.3944
R17354 gnd.n6814 gnd.n633 19.3944
R17355 gnd.n6757 gnd.n6616 19.3944
R17356 gnd.n6750 gnd.n6616 19.3944
R17357 gnd.n6750 gnd.n6749 19.3944
R17358 gnd.n6749 gnd.n6634 19.3944
R17359 gnd.n6742 gnd.n6634 19.3944
R17360 gnd.n6742 gnd.n6741 19.3944
R17361 gnd.n6741 gnd.n6642 19.3944
R17362 gnd.n6734 gnd.n6642 19.3944
R17363 gnd.n6734 gnd.n6733 19.3944
R17364 gnd.n6733 gnd.n6654 19.3944
R17365 gnd.n6726 gnd.n6654 19.3944
R17366 gnd.n6726 gnd.n6725 19.3944
R17367 gnd.n6725 gnd.n6662 19.3944
R17368 gnd.n6718 gnd.n6662 19.3944
R17369 gnd.n6718 gnd.n6717 19.3944
R17370 gnd.n6717 gnd.n6674 19.3944
R17371 gnd.n6707 gnd.n6674 19.3944
R17372 gnd.n6707 gnd.n6706 19.3944
R17373 gnd.n6706 gnd.n6705 19.3944
R17374 gnd.n6705 gnd.n6681 19.3944
R17375 gnd.n6701 gnd.n6681 19.3944
R17376 gnd.n6701 gnd.n6700 19.3944
R17377 gnd.n6700 gnd.n6699 19.3944
R17378 gnd.n6699 gnd.n6687 19.3944
R17379 gnd.n1200 gnd.t156 19.1199
R17380 gnd.n6141 gnd.n1093 19.1199
R17381 gnd.n6079 gnd.n1056 19.1199
R17382 gnd.n6446 gnd.n1006 19.1199
R17383 gnd.n6257 gnd.n968 19.1199
R17384 gnd.t130 gnd.n953 19.1199
R17385 gnd.n6798 gnd.n646 19.1199
R17386 gnd.n4179 gnd.t149 18.8012
R17387 gnd.n3612 gnd.t134 18.8012
R17388 gnd.n4049 gnd.n4048 18.4825
R17389 gnd.n6576 gnd.t85 18.4825
R17390 gnd.n7019 gnd.n7018 18.4247
R17391 gnd.n1606 gnd.n1386 18.4247
R17392 gnd.n7450 gnd.n120 18.2308
R17393 gnd.n6714 gnd.n6668 18.2308
R17394 gnd.n5775 gnd.n1347 18.2308
R17395 gnd.n4819 gnd.n4763 18.2308
R17396 gnd.t139 gnd.n3728 18.1639
R17397 gnd.n5852 gnd.t152 18.1639
R17398 gnd.t2 gnd.n879 18.1639
R17399 gnd.n6007 gnd.n1239 17.8452
R17400 gnd.n5883 gnd.n1216 17.8452
R17401 gnd.n1150 gnd.n1065 17.8452
R17402 gnd.n6454 gnd.n998 17.8452
R17403 gnd.n6381 gnd.n939 17.8452
R17404 gnd.n6551 gnd.n888 17.8452
R17405 gnd.n3757 gnd.t147 17.5266
R17406 gnd.n6149 gnd.t354 17.5266
R17407 gnd.n6306 gnd.t121 17.5266
R17408 gnd.n4657 gnd.n3355 17.2079
R17409 gnd.t120 gnd.n1248 17.2079
R17410 gnd.n6560 gnd.t169 17.2079
R17411 gnd.n7393 gnd.n236 17.2079
R17412 gnd.n4168 gnd.t143 16.8893
R17413 gnd.n5441 gnd.n1795 16.5706
R17414 gnd.n5469 gnd.n1758 16.5706
R17415 gnd.n5429 gnd.n1761 16.5706
R17416 gnd.n5249 gnd.n1752 16.5706
R17417 gnd.n5485 gnd.n1742 16.5706
R17418 gnd.n5276 gnd.n5275 16.5706
R17419 gnd.n5493 gnd.n1733 16.5706
R17420 gnd.n5501 gnd.n1724 16.5706
R17421 gnd.n5295 gnd.n1727 16.5706
R17422 gnd.n5289 gnd.n1718 16.5706
R17423 gnd.n5517 gnd.n1708 16.5706
R17424 gnd.n5316 gnd.n5315 16.5706
R17425 gnd.n5525 gnd.n1699 16.5706
R17426 gnd.n5533 gnd.n1690 16.5706
R17427 gnd.n5334 gnd.n1693 16.5706
R17428 gnd.n5328 gnd.n1684 16.5706
R17429 gnd.n5549 gnd.n1674 16.5706
R17430 gnd.n5373 gnd.n5372 16.5706
R17431 gnd.n5557 gnd.n1665 16.5706
R17432 gnd.n5384 gnd.n1668 16.5706
R17433 gnd.n5567 gnd.n1655 16.5706
R17434 gnd.n5386 gnd.n1658 16.5706
R17435 gnd.n5694 gnd.n1649 16.5706
R17436 gnd.n5771 gnd.n1354 16.5706
R17437 gnd.n6015 gnd.n1231 16.5706
R17438 gnd.n5920 gnd.n5888 16.5706
R17439 gnd.n6157 gnd.n1078 16.5706
R17440 gnd.n6094 gnd.n6093 16.5706
R17441 gnd.n6462 gnd.n990 16.5706
R17442 gnd.n6298 gnd.n6266 16.5706
R17443 gnd.n6374 gnd.n6373 16.5706
R17444 gnd.n6542 gnd.n920 16.5706
R17445 gnd.n6974 gnd.n480 16.5706
R17446 gnd.n7055 gnd.n483 16.5706
R17447 gnd.n6846 gnd.n471 16.5706
R17448 gnd.n7063 gnd.n474 16.5706
R17449 gnd.n6850 gnd.n462 16.5706
R17450 gnd.n7071 gnd.n465 16.5706
R17451 gnd.n6866 gnd.n6865 16.5706
R17452 gnd.n7079 gnd.n456 16.5706
R17453 gnd.n6859 gnd.n446 16.5706
R17454 gnd.n6886 gnd.n437 16.5706
R17455 gnd.n7095 gnd.n440 16.5706
R17456 gnd.n7103 gnd.n431 16.5706
R17457 gnd.n6905 gnd.n6904 16.5706
R17458 gnd.n7111 gnd.n422 16.5706
R17459 gnd.n6898 gnd.n412 16.5706
R17460 gnd.n6917 gnd.n401 16.5706
R17461 gnd.n7130 gnd.n404 16.5706
R17462 gnd.n7138 gnd.n386 16.5706
R17463 gnd.n7159 gnd.n7158 16.5706
R17464 gnd.n7181 gnd.n372 16.5706
R17465 gnd.n6930 gnd.n379 16.5706
R17466 gnd.n7190 gnd.n361 16.5706
R17467 gnd.n7212 gnd.n349 16.5706
R17468 gnd.n7320 gnd.n311 16.5706
R17469 gnd.n3984 gnd.t88 16.2519
R17470 gnd.n4216 gnd.t141 16.2519
R17471 gnd.n5437 gnd.t198 16.2519
R17472 gnd.n1312 gnd.t95 16.2519
R17473 gnd.n6808 gnd.t75 16.2519
R17474 gnd.t298 gnd.n308 16.2519
R17475 gnd.n5940 gnd.t0 15.9333
R17476 gnd.n6344 gnd.t127 15.9333
R17477 gnd.n4610 gnd.n4608 15.6674
R17478 gnd.n4578 gnd.n4576 15.6674
R17479 gnd.n4546 gnd.n4544 15.6674
R17480 gnd.n4515 gnd.n4513 15.6674
R17481 gnd.n4483 gnd.n4481 15.6674
R17482 gnd.n4451 gnd.n4449 15.6674
R17483 gnd.n4419 gnd.n4417 15.6674
R17484 gnd.n4388 gnd.n4386 15.6674
R17485 gnd.n3975 gnd.t88 15.6146
R17486 gnd.t37 gnd.n4646 15.6146
R17487 gnd.t65 gnd.n3364 15.6146
R17488 gnd.t200 gnd.n1736 15.6146
R17489 gnd.n5825 gnd.t95 15.6146
R17490 gnd.n6613 gnd.t75 15.6146
R17491 gnd.n7139 gnd.t243 15.6146
R17492 gnd.n5233 gnd.n1795 15.296
R17493 gnd.n5441 gnd.n5437 15.296
R17494 gnd.n5241 gnd.n1758 15.296
R17495 gnd.n5469 gnd.n1761 15.296
R17496 gnd.n5430 gnd.n5429 15.296
R17497 gnd.n5477 gnd.n1752 15.296
R17498 gnd.n5249 gnd.n1742 15.296
R17499 gnd.n5276 gnd.n1733 15.296
R17500 gnd.n5493 gnd.n1736 15.296
R17501 gnd.n5280 gnd.n1724 15.296
R17502 gnd.n5501 gnd.n1727 15.296
R17503 gnd.n5296 gnd.n5295 15.296
R17504 gnd.n5509 gnd.n1718 15.296
R17505 gnd.n5289 gnd.n1708 15.296
R17506 gnd.n5316 gnd.n1699 15.296
R17507 gnd.n5525 gnd.n1702 15.296
R17508 gnd.n5320 gnd.n1690 15.296
R17509 gnd.n5533 gnd.n1693 15.296
R17510 gnd.n5335 gnd.n5334 15.296
R17511 gnd.n5541 gnd.n1684 15.296
R17512 gnd.n5328 gnd.n1674 15.296
R17513 gnd.n5373 gnd.n1665 15.296
R17514 gnd.n5557 gnd.n1668 15.296
R17515 gnd.n5384 gnd.n1655 15.296
R17516 gnd.n5567 gnd.n1658 15.296
R17517 gnd.n5694 gnd.n1354 15.296
R17518 gnd.n5771 gnd.n1356 15.296
R17519 gnd.n6974 gnd.n564 15.296
R17520 gnd.n7055 gnd.n480 15.296
R17521 gnd.n7063 gnd.n471 15.296
R17522 gnd.n6850 gnd.n474 15.296
R17523 gnd.n7071 gnd.n462 15.296
R17524 gnd.n6865 gnd.n465 15.296
R17525 gnd.n6859 gnd.n456 15.296
R17526 gnd.n7087 gnd.n446 15.296
R17527 gnd.n6886 gnd.n6885 15.296
R17528 gnd.n7095 gnd.n437 15.296
R17529 gnd.n6890 gnd.n440 15.296
R17530 gnd.n7103 gnd.n428 15.296
R17531 gnd.n6904 gnd.n431 15.296
R17532 gnd.n6898 gnd.n422 15.296
R17533 gnd.n7119 gnd.n412 15.296
R17534 gnd.n6917 gnd.n6916 15.296
R17535 gnd.n7130 gnd.n401 15.296
R17536 gnd.n6938 gnd.n404 15.296
R17537 gnd.n7139 gnd.n7138 15.296
R17538 gnd.n7159 gnd.n386 15.296
R17539 gnd.n6930 gnd.n372 15.296
R17540 gnd.n7169 gnd.n379 15.296
R17541 gnd.n7190 gnd.n359 15.296
R17542 gnd.n361 gnd.n349 15.296
R17543 gnd.n7212 gnd.n7211 15.296
R17544 gnd.n7320 gnd.n308 15.296
R17545 gnd.n7202 gnd.n311 15.296
R17546 gnd.n713 gnd.n712 15.0827
R17547 gnd.n1422 gnd.n1417 15.0481
R17548 gnd.n723 gnd.n722 15.0481
R17549 gnd.n3440 gnd.t148 14.9773
R17550 gnd.t216 gnd.n1702 14.9773
R17551 gnd.t308 gnd.n428 14.9773
R17552 gnd.n6023 gnd.t166 14.6587
R17553 gnd.n6532 gnd.t179 14.6587
R17554 gnd.n3415 gnd.t159 14.34
R17555 gnd.n3398 gnd.t146 14.34
R17556 gnd.n5967 gnd.n1239 14.0214
R17557 gnd.t7 gnd.n1216 14.0214
R17558 gnd.n6109 gnd.n6108 14.0214
R17559 gnd.n6173 gnd.n1065 14.0214
R17560 gnd.n6414 gnd.n998 14.0214
R17561 gnd.n6478 gnd.n976 14.0214
R17562 gnd.t4 gnd.n939 14.0214
R17563 gnd.n6590 gnd.n888 14.0214
R17564 gnd.n6789 gnd.t12 14.0214
R17565 gnd.n4137 gnd.t188 13.7027
R17566 gnd.t190 gnd.n1233 13.7027
R17567 gnd.t177 gnd.n919 13.7027
R17568 gnd.n3841 gnd.n3840 13.5763
R17569 gnd.n4722 gnd.n2026 13.5763
R17570 gnd.n6981 gnd.n561 13.5763
R17571 gnd.n7502 gnd.n7501 13.5763
R17572 gnd.n4995 gnd.n4934 13.5763
R17573 gnd.n5705 gnd.n1643 13.5763
R17574 gnd.n4049 gnd.n3787 13.384
R17575 gnd.n1433 gnd.n1414 13.1884
R17576 gnd.n1428 gnd.n1427 13.1884
R17577 gnd.n1427 gnd.n1426 13.1884
R17578 gnd.n716 gnd.n711 13.1884
R17579 gnd.n717 gnd.n716 13.1884
R17580 gnd.n1429 gnd.n1416 13.146
R17581 gnd.n1425 gnd.n1416 13.146
R17582 gnd.n715 gnd.n714 13.146
R17583 gnd.n715 gnd.n710 13.146
R17584 gnd.n4611 gnd.n4607 12.8005
R17585 gnd.n4579 gnd.n4575 12.8005
R17586 gnd.n4547 gnd.n4543 12.8005
R17587 gnd.n4516 gnd.n4512 12.8005
R17588 gnd.n4484 gnd.n4480 12.8005
R17589 gnd.n4452 gnd.n4448 12.8005
R17590 gnd.n4420 gnd.n4416 12.8005
R17591 gnd.n4389 gnd.n4385 12.8005
R17592 gnd.n5835 gnd.n1295 12.7467
R17593 gnd.t52 gnd.t58 12.7467
R17594 gnd.n5853 gnd.n5852 12.7467
R17595 gnd.t187 gnd.n1231 12.7467
R17596 gnd.n6040 gnd.n1207 12.7467
R17597 gnd.n1119 gnd.n1093 12.7467
R17598 gnd.n6183 gnd.n1056 12.7467
R17599 gnd.t180 gnd.n1058 12.7467
R17600 gnd.n6422 gnd.t173 12.7467
R17601 gnd.n1033 gnd.n1006 12.7467
R17602 gnd.n6486 gnd.n968 12.7467
R17603 gnd.n6510 gnd.n947 12.7467
R17604 gnd.t172 gnd.n920 12.7467
R17605 gnd.n6600 gnd.n879 12.7467
R17606 gnd.t105 gnd.n898 12.7467
R17607 gnd.n1960 gnd.t208 12.4281
R17608 gnd.n5541 gnd.t220 12.4281
R17609 gnd.t123 gnd.n1207 12.4281
R17610 gnd.t170 gnd.n947 12.4281
R17611 gnd.n7087 gnd.t235 12.4281
R17612 gnd.t222 gnd.n225 12.4281
R17613 gnd.n3840 gnd.n3835 12.4126
R17614 gnd.n4725 gnd.n4722 12.4126
R17615 gnd.n6977 gnd.n561 12.4126
R17616 gnd.n7501 gnd.n196 12.4126
R17617 gnd.n4991 gnd.n4934 12.4126
R17618 gnd.n5700 gnd.n1643 12.4126
R17619 gnd.n1515 gnd.n1434 12.1761
R17620 gnd.n729 gnd.n728 12.1761
R17621 gnd.n4615 gnd.n4614 12.0247
R17622 gnd.n4583 gnd.n4582 12.0247
R17623 gnd.n4551 gnd.n4550 12.0247
R17624 gnd.n4520 gnd.n4519 12.0247
R17625 gnd.n4488 gnd.n4487 12.0247
R17626 gnd.n4456 gnd.n4455 12.0247
R17627 gnd.n4424 gnd.n4423 12.0247
R17628 gnd.n4393 gnd.n4392 12.0247
R17629 gnd.n1928 gnd.t265 11.7908
R17630 gnd.n5509 gnd.t237 11.7908
R17631 gnd.t44 gnd.n1649 11.7908
R17632 gnd.t33 gnd.n483 11.7908
R17633 gnd.n7119 gnd.t271 11.7908
R17634 gnd.t296 gnd.n256 11.7908
R17635 gnd.n5844 gnd.n1287 11.4721
R17636 gnd.n6049 gnd.n1199 11.4721
R17637 gnd.n1194 gnd.n1101 11.4721
R17638 gnd.n6192 gnd.n1049 11.4721
R17639 gnd.n1044 gnd.n1014 11.4721
R17640 gnd.n6494 gnd.n961 11.4721
R17641 gnd.n6502 gnd.n955 11.4721
R17642 gnd.n6577 gnd.n898 11.4721
R17643 gnd.n6775 gnd.n669 11.4721
R17644 gnd.n4618 gnd.n4605 11.249
R17645 gnd.n4586 gnd.n4573 11.249
R17646 gnd.n4554 gnd.n4541 11.249
R17647 gnd.n4523 gnd.n4510 11.249
R17648 gnd.n4491 gnd.n4478 11.249
R17649 gnd.n4459 gnd.n4446 11.249
R17650 gnd.n4427 gnd.n4414 11.249
R17651 gnd.n4396 gnd.n4383 11.249
R17652 gnd.n4127 gnd.t188 11.1535
R17653 gnd.n5184 gnd.t245 11.1535
R17654 gnd.n5477 gnd.t251 11.1535
R17655 gnd.n7169 gnd.t291 11.1535
R17656 gnd.t258 gnd.n286 11.1535
R17657 gnd.t99 gnd.n1295 10.8348
R17658 gnd.t182 gnd.n1103 10.8348
R17659 gnd.n6117 gnd.t182 10.8348
R17660 gnd.t1 gnd.n970 10.8348
R17661 gnd.n6326 gnd.t1 10.8348
R17662 gnd.n803 gnd.n802 10.6151
R17663 gnd.n807 gnd.n803 10.6151
R17664 gnd.n813 gnd.n691 10.6151
R17665 gnd.n814 gnd.n813 10.6151
R17666 gnd.n815 gnd.n814 10.6151
R17667 gnd.n815 gnd.n689 10.6151
R17668 gnd.n821 gnd.n689 10.6151
R17669 gnd.n822 gnd.n821 10.6151
R17670 gnd.n823 gnd.n822 10.6151
R17671 gnd.n823 gnd.n687 10.6151
R17672 gnd.n829 gnd.n687 10.6151
R17673 gnd.n830 gnd.n829 10.6151
R17674 gnd.n831 gnd.n830 10.6151
R17675 gnd.n831 gnd.n685 10.6151
R17676 gnd.n837 gnd.n685 10.6151
R17677 gnd.n838 gnd.n837 10.6151
R17678 gnd.n839 gnd.n838 10.6151
R17679 gnd.n839 gnd.n683 10.6151
R17680 gnd.n845 gnd.n683 10.6151
R17681 gnd.n846 gnd.n845 10.6151
R17682 gnd.n847 gnd.n846 10.6151
R17683 gnd.n847 gnd.n681 10.6151
R17684 gnd.n853 gnd.n681 10.6151
R17685 gnd.n854 gnd.n853 10.6151
R17686 gnd.n855 gnd.n854 10.6151
R17687 gnd.n855 gnd.n679 10.6151
R17688 gnd.n860 gnd.n679 10.6151
R17689 gnd.n861 gnd.n860 10.6151
R17690 gnd.n861 gnd.n677 10.6151
R17691 gnd.n866 gnd.n677 10.6151
R17692 gnd.n1535 gnd.n1410 10.6151
R17693 gnd.n1535 gnd.n1534 10.6151
R17694 gnd.n1534 gnd.n1533 10.6151
R17695 gnd.n1533 gnd.n1268 10.6151
R17696 gnd.n5981 gnd.n1268 10.6151
R17697 gnd.n5981 gnd.n5980 10.6151
R17698 gnd.n5980 gnd.n5979 10.6151
R17699 gnd.n5979 gnd.n1269 10.6151
R17700 gnd.n1271 gnd.n1269 10.6151
R17701 gnd.n5893 gnd.n1271 10.6151
R17702 gnd.n5895 gnd.n5893 10.6151
R17703 gnd.n5896 gnd.n5895 10.6151
R17704 gnd.n5898 gnd.n5896 10.6151
R17705 gnd.n5899 gnd.n5898 10.6151
R17706 gnd.n5900 gnd.n5899 10.6151
R17707 gnd.n5900 gnd.n5891 10.6151
R17708 gnd.n5915 gnd.n5891 10.6151
R17709 gnd.n5916 gnd.n5915 10.6151
R17710 gnd.n5918 gnd.n5916 10.6151
R17711 gnd.n5918 gnd.n5917 10.6151
R17712 gnd.n5917 gnd.n5882 10.6151
R17713 gnd.n5882 gnd.n5880 10.6151
R17714 gnd.n5931 gnd.n5880 10.6151
R17715 gnd.n5932 gnd.n5931 10.6151
R17716 gnd.n5934 gnd.n5932 10.6151
R17717 gnd.n5935 gnd.n5934 10.6151
R17718 gnd.n5937 gnd.n5935 10.6151
R17719 gnd.n5937 gnd.n5936 10.6151
R17720 gnd.n5936 gnd.n1115 10.6151
R17721 gnd.n6123 gnd.n1115 10.6151
R17722 gnd.n6123 gnd.n6122 10.6151
R17723 gnd.n6122 gnd.n6121 10.6151
R17724 gnd.n6121 gnd.n1116 10.6151
R17725 gnd.n1118 gnd.n1116 10.6151
R17726 gnd.n1128 gnd.n1118 10.6151
R17727 gnd.n1130 gnd.n1128 10.6151
R17728 gnd.n1131 gnd.n1130 10.6151
R17729 gnd.n6106 gnd.n1131 10.6151
R17730 gnd.n6106 gnd.n6105 10.6151
R17731 gnd.n6105 gnd.n6104 10.6151
R17732 gnd.n6104 gnd.n1132 10.6151
R17733 gnd.n1145 gnd.n1132 10.6151
R17734 gnd.n1146 gnd.n1145 10.6151
R17735 gnd.n6091 gnd.n1146 10.6151
R17736 gnd.n6091 gnd.n6090 10.6151
R17737 gnd.n6090 gnd.n6089 10.6151
R17738 gnd.n6089 gnd.n1147 10.6151
R17739 gnd.n1159 gnd.n1147 10.6151
R17740 gnd.n1184 gnd.n1159 10.6151
R17741 gnd.n1184 gnd.n1183 10.6151
R17742 gnd.n1183 gnd.n1182 10.6151
R17743 gnd.n1182 gnd.n1160 10.6151
R17744 gnd.n1161 gnd.n1160 10.6151
R17745 gnd.n1161 gnd.n1029 10.6151
R17746 gnd.n6428 gnd.n1029 10.6151
R17747 gnd.n6428 gnd.n6427 10.6151
R17748 gnd.n6427 gnd.n6426 10.6151
R17749 gnd.n6426 gnd.n1030 10.6151
R17750 gnd.n1032 gnd.n1030 10.6151
R17751 gnd.n6276 gnd.n1032 10.6151
R17752 gnd.n6278 gnd.n6276 10.6151
R17753 gnd.n6279 gnd.n6278 10.6151
R17754 gnd.n6281 gnd.n6279 10.6151
R17755 gnd.n6282 gnd.n6281 10.6151
R17756 gnd.n6286 gnd.n6282 10.6151
R17757 gnd.n6286 gnd.n6285 10.6151
R17758 gnd.n6285 gnd.n6284 10.6151
R17759 gnd.n6284 gnd.n6264 10.6151
R17760 gnd.n6300 gnd.n6264 10.6151
R17761 gnd.n6301 gnd.n6300 10.6151
R17762 gnd.n6304 gnd.n6301 10.6151
R17763 gnd.n6304 gnd.n6303 10.6151
R17764 gnd.n6303 gnd.n6302 10.6151
R17765 gnd.n6302 gnd.n6254 10.6151
R17766 gnd.n6319 gnd.n6254 10.6151
R17767 gnd.n6320 gnd.n6319 10.6151
R17768 gnd.n6323 gnd.n6320 10.6151
R17769 gnd.n6323 gnd.n6322 10.6151
R17770 gnd.n6322 gnd.n6321 10.6151
R17771 gnd.n6321 gnd.n6245 10.6151
R17772 gnd.n6338 gnd.n6245 10.6151
R17773 gnd.n6339 gnd.n6338 10.6151
R17774 gnd.n6342 gnd.n6339 10.6151
R17775 gnd.n6342 gnd.n6341 10.6151
R17776 gnd.n6341 gnd.n6340 10.6151
R17777 gnd.n6340 gnd.n6236 10.6151
R17778 gnd.n6236 gnd.n6234 10.6151
R17779 gnd.n6356 gnd.n6234 10.6151
R17780 gnd.n6357 gnd.n6356 10.6151
R17781 gnd.n6359 gnd.n6357 10.6151
R17782 gnd.n6360 gnd.n6359 10.6151
R17783 gnd.n6370 gnd.n6360 10.6151
R17784 gnd.n6370 gnd.n6369 10.6151
R17785 gnd.n6369 gnd.n6368 10.6151
R17786 gnd.n6368 gnd.n6365 10.6151
R17787 gnd.n6365 gnd.n6364 10.6151
R17788 gnd.n6364 gnd.n6363 10.6151
R17789 gnd.n6363 gnd.n6361 10.6151
R17790 gnd.n6361 gnd.n904 10.6151
R17791 gnd.n6563 gnd.n904 10.6151
R17792 gnd.n6564 gnd.n6563 10.6151
R17793 gnd.n6566 gnd.n6564 10.6151
R17794 gnd.n6566 gnd.n6565 10.6151
R17795 gnd.n6565 gnd.n666 10.6151
R17796 gnd.n6779 gnd.n666 10.6151
R17797 gnd.n6779 gnd.n6778 10.6151
R17798 gnd.n6778 gnd.n6777 10.6151
R17799 gnd.n6777 gnd.n667 10.6151
R17800 gnd.n868 gnd.n667 10.6151
R17801 gnd.n868 gnd.n867 10.6151
R17802 gnd.n1599 gnd.n1390 10.6151
R17803 gnd.n1599 gnd.n1598 10.6151
R17804 gnd.n1596 gnd.n1396 10.6151
R17805 gnd.n1590 gnd.n1396 10.6151
R17806 gnd.n1590 gnd.n1589 10.6151
R17807 gnd.n1589 gnd.n1588 10.6151
R17808 gnd.n1588 gnd.n1398 10.6151
R17809 gnd.n1582 gnd.n1398 10.6151
R17810 gnd.n1582 gnd.n1581 10.6151
R17811 gnd.n1581 gnd.n1580 10.6151
R17812 gnd.n1580 gnd.n1400 10.6151
R17813 gnd.n1574 gnd.n1400 10.6151
R17814 gnd.n1574 gnd.n1573 10.6151
R17815 gnd.n1573 gnd.n1572 10.6151
R17816 gnd.n1572 gnd.n1402 10.6151
R17817 gnd.n1566 gnd.n1402 10.6151
R17818 gnd.n1566 gnd.n1565 10.6151
R17819 gnd.n1565 gnd.n1564 10.6151
R17820 gnd.n1564 gnd.n1404 10.6151
R17821 gnd.n1558 gnd.n1404 10.6151
R17822 gnd.n1558 gnd.n1557 10.6151
R17823 gnd.n1557 gnd.n1556 10.6151
R17824 gnd.n1556 gnd.n1406 10.6151
R17825 gnd.n1550 gnd.n1406 10.6151
R17826 gnd.n1550 gnd.n1549 10.6151
R17827 gnd.n1549 gnd.n1548 10.6151
R17828 gnd.n1548 gnd.n1408 10.6151
R17829 gnd.n1542 gnd.n1408 10.6151
R17830 gnd.n1542 gnd.n1541 10.6151
R17831 gnd.n1541 gnd.n1540 10.6151
R17832 gnd.n1515 gnd.n1514 10.6151
R17833 gnd.n1514 gnd.n1436 10.6151
R17834 gnd.n1510 gnd.n1436 10.6151
R17835 gnd.n1510 gnd.n1509 10.6151
R17836 gnd.n1509 gnd.n1438 10.6151
R17837 gnd.n1504 gnd.n1438 10.6151
R17838 gnd.n1504 gnd.n1503 10.6151
R17839 gnd.n1503 gnd.n1502 10.6151
R17840 gnd.n1502 gnd.n1440 10.6151
R17841 gnd.n1496 gnd.n1440 10.6151
R17842 gnd.n1496 gnd.n1495 10.6151
R17843 gnd.n1495 gnd.n1494 10.6151
R17844 gnd.n1494 gnd.n1442 10.6151
R17845 gnd.n1488 gnd.n1442 10.6151
R17846 gnd.n1488 gnd.n1487 10.6151
R17847 gnd.n1487 gnd.n1486 10.6151
R17848 gnd.n1486 gnd.n1444 10.6151
R17849 gnd.n1480 gnd.n1444 10.6151
R17850 gnd.n1480 gnd.n1479 10.6151
R17851 gnd.n1479 gnd.n1478 10.6151
R17852 gnd.n1478 gnd.n1446 10.6151
R17853 gnd.n1472 gnd.n1446 10.6151
R17854 gnd.n1472 gnd.n1471 10.6151
R17855 gnd.n1471 gnd.n1470 10.6151
R17856 gnd.n1470 gnd.n1448 10.6151
R17857 gnd.n1464 gnd.n1448 10.6151
R17858 gnd.n1464 gnd.n1463 10.6151
R17859 gnd.n1463 gnd.n1462 10.6151
R17860 gnd.n1458 gnd.n1457 10.6151
R17861 gnd.n1457 gnd.n1391 10.6151
R17862 gnd.n729 gnd.n708 10.6151
R17863 gnd.n735 gnd.n708 10.6151
R17864 gnd.n736 gnd.n735 10.6151
R17865 gnd.n737 gnd.n736 10.6151
R17866 gnd.n737 gnd.n706 10.6151
R17867 gnd.n743 gnd.n706 10.6151
R17868 gnd.n744 gnd.n743 10.6151
R17869 gnd.n745 gnd.n744 10.6151
R17870 gnd.n745 gnd.n704 10.6151
R17871 gnd.n751 gnd.n704 10.6151
R17872 gnd.n752 gnd.n751 10.6151
R17873 gnd.n753 gnd.n752 10.6151
R17874 gnd.n753 gnd.n702 10.6151
R17875 gnd.n759 gnd.n702 10.6151
R17876 gnd.n760 gnd.n759 10.6151
R17877 gnd.n761 gnd.n760 10.6151
R17878 gnd.n761 gnd.n700 10.6151
R17879 gnd.n767 gnd.n700 10.6151
R17880 gnd.n768 gnd.n767 10.6151
R17881 gnd.n769 gnd.n768 10.6151
R17882 gnd.n769 gnd.n698 10.6151
R17883 gnd.n775 gnd.n698 10.6151
R17884 gnd.n776 gnd.n775 10.6151
R17885 gnd.n777 gnd.n776 10.6151
R17886 gnd.n777 gnd.n696 10.6151
R17887 gnd.n783 gnd.n696 10.6151
R17888 gnd.n784 gnd.n783 10.6151
R17889 gnd.n788 gnd.n784 10.6151
R17890 gnd.n793 gnd.n694 10.6151
R17891 gnd.n794 gnd.n793 10.6151
R17892 gnd.n1519 gnd.n1518 10.6151
R17893 gnd.n1528 gnd.n1519 10.6151
R17894 gnd.n1528 gnd.n1527 10.6151
R17895 gnd.n1527 gnd.n1526 10.6151
R17896 gnd.n1526 gnd.n1524 10.6151
R17897 gnd.n1524 gnd.n1523 10.6151
R17898 gnd.n1523 gnd.n1520 10.6151
R17899 gnd.n1520 gnd.n1274 10.6151
R17900 gnd.n5973 gnd.n1274 10.6151
R17901 gnd.n5973 gnd.n5972 10.6151
R17902 gnd.n5972 gnd.n5971 10.6151
R17903 gnd.n5971 gnd.n1275 10.6151
R17904 gnd.n5904 gnd.n1275 10.6151
R17905 gnd.n5905 gnd.n5904 10.6151
R17906 gnd.n5909 gnd.n5905 10.6151
R17907 gnd.n5909 gnd.n5908 10.6151
R17908 gnd.n5908 gnd.n5907 10.6151
R17909 gnd.n5907 gnd.n5886 10.6151
R17910 gnd.n5922 gnd.n5886 10.6151
R17911 gnd.n5923 gnd.n5922 10.6151
R17912 gnd.n5925 gnd.n5923 10.6151
R17913 gnd.n5925 gnd.n5924 10.6151
R17914 gnd.n5924 gnd.n5867 10.6151
R17915 gnd.n5945 gnd.n5867 10.6151
R17916 gnd.n5945 gnd.n5944 10.6151
R17917 gnd.n5944 gnd.n5943 10.6151
R17918 gnd.n5943 gnd.n5868 10.6151
R17919 gnd.n5876 gnd.n5868 10.6151
R17920 gnd.n5876 gnd.n5875 10.6151
R17921 gnd.n5875 gnd.n5874 10.6151
R17922 gnd.n5874 gnd.n5873 10.6151
R17923 gnd.n5873 gnd.n5870 10.6151
R17924 gnd.n5870 gnd.n1122 10.6151
R17925 gnd.n6115 gnd.n1122 10.6151
R17926 gnd.n6115 gnd.n6114 10.6151
R17927 gnd.n6114 gnd.n6113 10.6151
R17928 gnd.n6113 gnd.n1123 10.6151
R17929 gnd.n1137 gnd.n1123 10.6151
R17930 gnd.n1138 gnd.n1137 10.6151
R17931 gnd.n6100 gnd.n1138 10.6151
R17932 gnd.n6100 gnd.n6099 10.6151
R17933 gnd.n6099 gnd.n6098 10.6151
R17934 gnd.n6098 gnd.n1139 10.6151
R17935 gnd.n1153 gnd.n1139 10.6151
R17936 gnd.n1154 gnd.n1153 10.6151
R17937 gnd.n6085 gnd.n1154 10.6151
R17938 gnd.n6085 gnd.n6084 10.6151
R17939 gnd.n6084 gnd.n6083 10.6151
R17940 gnd.n6083 gnd.n1155 10.6151
R17941 gnd.n1167 gnd.n1155 10.6151
R17942 gnd.n1168 gnd.n1167 10.6151
R17943 gnd.n1177 gnd.n1168 10.6151
R17944 gnd.n1177 gnd.n1176 10.6151
R17945 gnd.n1176 gnd.n1175 10.6151
R17946 gnd.n1175 gnd.n1173 10.6151
R17947 gnd.n1173 gnd.n1172 10.6151
R17948 gnd.n1172 gnd.n1169 10.6151
R17949 gnd.n1169 gnd.n1036 10.6151
R17950 gnd.n6420 gnd.n1036 10.6151
R17951 gnd.n6420 gnd.n6419 10.6151
R17952 gnd.n6419 gnd.n6418 10.6151
R17953 gnd.n6418 gnd.n1037 10.6151
R17954 gnd.n6271 gnd.n1037 10.6151
R17955 gnd.n6272 gnd.n6271 10.6151
R17956 gnd.n6273 gnd.n6272 10.6151
R17957 gnd.n6273 gnd.n6269 10.6151
R17958 gnd.n6293 gnd.n6269 10.6151
R17959 gnd.n6294 gnd.n6293 10.6151
R17960 gnd.n6296 gnd.n6294 10.6151
R17961 gnd.n6296 gnd.n6295 10.6151
R17962 gnd.n6295 gnd.n6260 10.6151
R17963 gnd.n6310 gnd.n6260 10.6151
R17964 gnd.n6311 gnd.n6310 10.6151
R17965 gnd.n6314 gnd.n6311 10.6151
R17966 gnd.n6314 gnd.n6313 10.6151
R17967 gnd.n6313 gnd.n6312 10.6151
R17968 gnd.n6312 gnd.n6250 10.6151
R17969 gnd.n6329 gnd.n6250 10.6151
R17970 gnd.n6330 gnd.n6329 10.6151
R17971 gnd.n6333 gnd.n6330 10.6151
R17972 gnd.n6333 gnd.n6332 10.6151
R17973 gnd.n6332 gnd.n6331 10.6151
R17974 gnd.n6331 gnd.n6240 10.6151
R17975 gnd.n6347 gnd.n6240 10.6151
R17976 gnd.n6348 gnd.n6347 10.6151
R17977 gnd.n6350 gnd.n6348 10.6151
R17978 gnd.n6350 gnd.n6349 10.6151
R17979 gnd.n6349 gnd.n6224 10.6151
R17980 gnd.n6378 gnd.n6224 10.6151
R17981 gnd.n6378 gnd.n6377 10.6151
R17982 gnd.n6377 gnd.n6376 10.6151
R17983 gnd.n6376 gnd.n6225 10.6151
R17984 gnd.n6229 gnd.n6225 10.6151
R17985 gnd.n6229 gnd.n6228 10.6151
R17986 gnd.n6228 gnd.n6227 10.6151
R17987 gnd.n6227 gnd.n909 10.6151
R17988 gnd.n6555 gnd.n909 10.6151
R17989 gnd.n6556 gnd.n6555 10.6151
R17990 gnd.n6558 gnd.n6556 10.6151
R17991 gnd.n6558 gnd.n6557 10.6151
R17992 gnd.n6557 gnd.n900 10.6151
R17993 gnd.n6571 gnd.n900 10.6151
R17994 gnd.n6572 gnd.n6571 10.6151
R17995 gnd.n6574 gnd.n6572 10.6151
R17996 gnd.n6574 gnd.n6573 10.6151
R17997 gnd.n6573 gnd.n673 10.6151
R17998 gnd.n6773 gnd.n673 10.6151
R17999 gnd.n6773 gnd.n6772 10.6151
R18000 gnd.n6772 gnd.n6771 10.6151
R18001 gnd.n6771 gnd.n674 10.6151
R18002 gnd.n4038 gnd.t131 10.5161
R18003 gnd.n4349 gnd.t159 10.5161
R18004 gnd.t146 gnd.n3387 10.5161
R18005 gnd.n5455 gnd.t206 10.5161
R18006 gnd.n5447 gnd.n1788 10.5161
R18007 gnd.n5447 gnd.t229 10.5161
R18008 gnd.n7222 gnd.t218 10.5161
R18009 gnd.n7222 gnd.n7221 10.5161
R18010 gnd.n7228 gnd.t305 10.5161
R18011 gnd.n4619 gnd.n4603 10.4732
R18012 gnd.n4587 gnd.n4571 10.4732
R18013 gnd.n4555 gnd.n4539 10.4732
R18014 gnd.n4524 gnd.n4508 10.4732
R18015 gnd.n4492 gnd.n4476 10.4732
R18016 gnd.n4460 gnd.n4444 10.4732
R18017 gnd.n4428 gnd.n4412 10.4732
R18018 gnd.n4397 gnd.n4381 10.4732
R18019 gnd.n5844 gnd.n1288 10.1975
R18020 gnd.n1282 gnd.n1264 10.1975
R18021 gnd.n6049 gnd.n1200 10.1975
R18022 gnd.n6192 gnd.n1022 10.1975
R18023 gnd.n1044 gnd.n1025 10.1975
R18024 gnd.n6502 gnd.n953 10.1975
R18025 gnd.n6577 gnd.n6576 10.1975
R18026 gnd.n670 gnd.n669 10.1975
R18027 gnd.n4318 gnd.t148 9.87883
R18028 gnd.n5190 gnd.t204 9.87883
R18029 gnd.n5485 gnd.t210 9.87883
R18030 gnd.n7181 gnd.t225 9.87883
R18031 gnd.n289 gnd.t255 9.87883
R18032 gnd.n7627 gnd.n74 9.81789
R18033 gnd.n4623 gnd.n4622 9.69747
R18034 gnd.n4591 gnd.n4590 9.69747
R18035 gnd.n4559 gnd.n4558 9.69747
R18036 gnd.n4528 gnd.n4527 9.69747
R18037 gnd.n4496 gnd.n4495 9.69747
R18038 gnd.n4464 gnd.n4463 9.69747
R18039 gnd.n4432 gnd.n4431 9.69747
R18040 gnd.n4401 gnd.n4400 9.69747
R18041 gnd.n1134 gnd.t183 9.56018
R18042 gnd.n6470 gnd.t181 9.56018
R18043 gnd.n5689 gnd.n5573 9.45599
R18044 gnd.n6622 gnd.n6620 9.45599
R18045 gnd.n4629 gnd.n4628 9.45567
R18046 gnd.n4597 gnd.n4596 9.45567
R18047 gnd.n4565 gnd.n4564 9.45567
R18048 gnd.n4534 gnd.n4533 9.45567
R18049 gnd.n4502 gnd.n4501 9.45567
R18050 gnd.n4470 gnd.n4469 9.45567
R18051 gnd.n4438 gnd.n4437 9.45567
R18052 gnd.n4407 gnd.n4406 9.45567
R18053 gnd.n3676 gnd.n3675 9.39724
R18054 gnd.n4628 gnd.n4627 9.3005
R18055 gnd.n4601 gnd.n4600 9.3005
R18056 gnd.n4622 gnd.n4621 9.3005
R18057 gnd.n4620 gnd.n4619 9.3005
R18058 gnd.n4605 gnd.n4604 9.3005
R18059 gnd.n4614 gnd.n4613 9.3005
R18060 gnd.n4612 gnd.n4611 9.3005
R18061 gnd.n4596 gnd.n4595 9.3005
R18062 gnd.n4569 gnd.n4568 9.3005
R18063 gnd.n4590 gnd.n4589 9.3005
R18064 gnd.n4588 gnd.n4587 9.3005
R18065 gnd.n4573 gnd.n4572 9.3005
R18066 gnd.n4582 gnd.n4581 9.3005
R18067 gnd.n4580 gnd.n4579 9.3005
R18068 gnd.n4564 gnd.n4563 9.3005
R18069 gnd.n4537 gnd.n4536 9.3005
R18070 gnd.n4558 gnd.n4557 9.3005
R18071 gnd.n4556 gnd.n4555 9.3005
R18072 gnd.n4541 gnd.n4540 9.3005
R18073 gnd.n4550 gnd.n4549 9.3005
R18074 gnd.n4548 gnd.n4547 9.3005
R18075 gnd.n4533 gnd.n4532 9.3005
R18076 gnd.n4506 gnd.n4505 9.3005
R18077 gnd.n4527 gnd.n4526 9.3005
R18078 gnd.n4525 gnd.n4524 9.3005
R18079 gnd.n4510 gnd.n4509 9.3005
R18080 gnd.n4519 gnd.n4518 9.3005
R18081 gnd.n4517 gnd.n4516 9.3005
R18082 gnd.n4501 gnd.n4500 9.3005
R18083 gnd.n4474 gnd.n4473 9.3005
R18084 gnd.n4495 gnd.n4494 9.3005
R18085 gnd.n4493 gnd.n4492 9.3005
R18086 gnd.n4478 gnd.n4477 9.3005
R18087 gnd.n4487 gnd.n4486 9.3005
R18088 gnd.n4485 gnd.n4484 9.3005
R18089 gnd.n4469 gnd.n4468 9.3005
R18090 gnd.n4442 gnd.n4441 9.3005
R18091 gnd.n4463 gnd.n4462 9.3005
R18092 gnd.n4461 gnd.n4460 9.3005
R18093 gnd.n4446 gnd.n4445 9.3005
R18094 gnd.n4455 gnd.n4454 9.3005
R18095 gnd.n4453 gnd.n4452 9.3005
R18096 gnd.n4437 gnd.n4436 9.3005
R18097 gnd.n4410 gnd.n4409 9.3005
R18098 gnd.n4431 gnd.n4430 9.3005
R18099 gnd.n4429 gnd.n4428 9.3005
R18100 gnd.n4414 gnd.n4413 9.3005
R18101 gnd.n4423 gnd.n4422 9.3005
R18102 gnd.n4421 gnd.n4420 9.3005
R18103 gnd.n4406 gnd.n4405 9.3005
R18104 gnd.n4379 gnd.n4378 9.3005
R18105 gnd.n4400 gnd.n4399 9.3005
R18106 gnd.n4398 gnd.n4397 9.3005
R18107 gnd.n4383 gnd.n4382 9.3005
R18108 gnd.n4392 gnd.n4391 9.3005
R18109 gnd.n4390 gnd.n4389 9.3005
R18110 gnd.n4752 gnd.n4751 9.3005
R18111 gnd.n4750 gnd.n2014 9.3005
R18112 gnd.n4749 gnd.n4748 9.3005
R18113 gnd.n4745 gnd.n2015 9.3005
R18114 gnd.n4742 gnd.n2016 9.3005
R18115 gnd.n4741 gnd.n2017 9.3005
R18116 gnd.n4738 gnd.n2018 9.3005
R18117 gnd.n4737 gnd.n2019 9.3005
R18118 gnd.n4734 gnd.n2020 9.3005
R18119 gnd.n4733 gnd.n2021 9.3005
R18120 gnd.n4730 gnd.n2022 9.3005
R18121 gnd.n4729 gnd.n2023 9.3005
R18122 gnd.n4726 gnd.n2024 9.3005
R18123 gnd.n4725 gnd.n2025 9.3005
R18124 gnd.n4722 gnd.n4721 9.3005
R18125 gnd.n4720 gnd.n2026 9.3005
R18126 gnd.n4753 gnd.n2013 9.3005
R18127 gnd.n4057 gnd.n4056 9.3005
R18128 gnd.n3761 gnd.n3760 9.3005
R18129 gnd.n4084 gnd.n4083 9.3005
R18130 gnd.n4085 gnd.n3759 9.3005
R18131 gnd.n4089 gnd.n4086 9.3005
R18132 gnd.n4088 gnd.n4087 9.3005
R18133 gnd.n3733 gnd.n3732 9.3005
R18134 gnd.n4114 gnd.n4113 9.3005
R18135 gnd.n4115 gnd.n3731 9.3005
R18136 gnd.n4125 gnd.n4116 9.3005
R18137 gnd.n4124 gnd.n4117 9.3005
R18138 gnd.n4123 gnd.n4118 9.3005
R18139 gnd.n4121 gnd.n4120 9.3005
R18140 gnd.n4119 gnd.n3703 9.3005
R18141 gnd.n3701 gnd.n3700 9.3005
R18142 gnd.n4173 gnd.n4172 9.3005
R18143 gnd.n4174 gnd.n3699 9.3005
R18144 gnd.n4176 gnd.n4175 9.3005
R18145 gnd.n3519 gnd.n3518 9.3005
R18146 gnd.n4209 gnd.n4208 9.3005
R18147 gnd.n4210 gnd.n3517 9.3005
R18148 gnd.n4214 gnd.n4211 9.3005
R18149 gnd.n4213 gnd.n4212 9.3005
R18150 gnd.n3495 gnd.n3494 9.3005
R18151 gnd.n4240 gnd.n4239 9.3005
R18152 gnd.n4241 gnd.n3493 9.3005
R18153 gnd.n4245 gnd.n4242 9.3005
R18154 gnd.n4244 gnd.n4243 9.3005
R18155 gnd.n3469 gnd.n3468 9.3005
R18156 gnd.n4271 gnd.n4270 9.3005
R18157 gnd.n4272 gnd.n3467 9.3005
R18158 gnd.n4276 gnd.n4273 9.3005
R18159 gnd.n4275 gnd.n4274 9.3005
R18160 gnd.n3444 gnd.n3443 9.3005
R18161 gnd.n4302 gnd.n4301 9.3005
R18162 gnd.n4303 gnd.n3442 9.3005
R18163 gnd.n4307 gnd.n4304 9.3005
R18164 gnd.n4306 gnd.n4305 9.3005
R18165 gnd.n3419 gnd.n3418 9.3005
R18166 gnd.n4333 gnd.n4332 9.3005
R18167 gnd.n4334 gnd.n3417 9.3005
R18168 gnd.n4338 gnd.n4335 9.3005
R18169 gnd.n4337 gnd.n4336 9.3005
R18170 gnd.n3393 gnd.n3392 9.3005
R18171 gnd.n4364 gnd.n4363 9.3005
R18172 gnd.n4365 gnd.n3391 9.3005
R18173 gnd.n4369 gnd.n4366 9.3005
R18174 gnd.n4368 gnd.n4367 9.3005
R18175 gnd.n3368 gnd.n3367 9.3005
R18176 gnd.n4650 gnd.n4649 9.3005
R18177 gnd.n4651 gnd.n3366 9.3005
R18178 gnd.n4655 gnd.n4652 9.3005
R18179 gnd.n4654 gnd.n4653 9.3005
R18180 gnd.n4058 gnd.n4055 9.3005
R18181 gnd.n3840 gnd.n3799 9.3005
R18182 gnd.n3835 gnd.n3834 9.3005
R18183 gnd.n3833 gnd.n3800 9.3005
R18184 gnd.n3832 gnd.n3831 9.3005
R18185 gnd.n3828 gnd.n3801 9.3005
R18186 gnd.n3825 gnd.n3824 9.3005
R18187 gnd.n3823 gnd.n3802 9.3005
R18188 gnd.n3822 gnd.n3821 9.3005
R18189 gnd.n3818 gnd.n3803 9.3005
R18190 gnd.n3815 gnd.n3814 9.3005
R18191 gnd.n3813 gnd.n3804 9.3005
R18192 gnd.n3812 gnd.n3811 9.3005
R18193 gnd.n3808 gnd.n3806 9.3005
R18194 gnd.n3805 gnd.n3785 9.3005
R18195 gnd.n4052 gnd.n3784 9.3005
R18196 gnd.n4054 gnd.n4053 9.3005
R18197 gnd.n3842 gnd.n3841 9.3005
R18198 gnd.n4065 gnd.n3771 9.3005
R18199 gnd.n4072 gnd.n3772 9.3005
R18200 gnd.n4074 gnd.n4073 9.3005
R18201 gnd.n4075 gnd.n3752 9.3005
R18202 gnd.n4094 gnd.n4093 9.3005
R18203 gnd.n4096 gnd.n3744 9.3005
R18204 gnd.n4103 gnd.n3746 9.3005
R18205 gnd.n4104 gnd.n3741 9.3005
R18206 gnd.n4106 gnd.n4105 9.3005
R18207 gnd.n3742 gnd.n3727 9.3005
R18208 gnd.n3725 gnd.n3723 9.3005
R18209 gnd.n4132 gnd.n4131 9.3005
R18210 gnd.n3708 gnd.n3707 9.3005
R18211 gnd.n4165 gnd.n4153 9.3005
R18212 gnd.n4164 gnd.n4155 9.3005
R18213 gnd.n4163 gnd.n4156 9.3005
R18214 gnd.n4158 gnd.n4157 9.3005
R18215 gnd.n3691 gnd.n3528 9.3005
R18216 gnd.n4197 gnd.n3529 9.3005
R18217 gnd.n4199 gnd.n4198 9.3005
R18218 gnd.n4200 gnd.n3512 9.3005
R18219 gnd.n4219 gnd.n4218 9.3005
R18220 gnd.n4221 gnd.n3505 9.3005
R18221 gnd.n4228 gnd.n3506 9.3005
R18222 gnd.n4230 gnd.n4229 9.3005
R18223 gnd.n4231 gnd.n3487 9.3005
R18224 gnd.n4250 gnd.n4249 9.3005
R18225 gnd.n4252 gnd.n3479 9.3005
R18226 gnd.n4259 gnd.n3480 9.3005
R18227 gnd.n4261 gnd.n4260 9.3005
R18228 gnd.n4262 gnd.n3460 9.3005
R18229 gnd.n4281 gnd.n4280 9.3005
R18230 gnd.n4283 gnd.n3453 9.3005
R18231 gnd.n4290 gnd.n3454 9.3005
R18232 gnd.n4292 gnd.n4291 9.3005
R18233 gnd.n4293 gnd.n3436 9.3005
R18234 gnd.n4312 gnd.n4311 9.3005
R18235 gnd.n4314 gnd.n3429 9.3005
R18236 gnd.n4321 gnd.n3430 9.3005
R18237 gnd.n4323 gnd.n4322 9.3005
R18238 gnd.n4324 gnd.n3410 9.3005
R18239 gnd.n4343 gnd.n4342 9.3005
R18240 gnd.n4345 gnd.n3403 9.3005
R18241 gnd.n4352 gnd.n3404 9.3005
R18242 gnd.n4354 gnd.n4353 9.3005
R18243 gnd.n4355 gnd.n3385 9.3005
R18244 gnd.n4374 gnd.n4373 9.3005
R18245 gnd.n4376 gnd.n3377 9.3005
R18246 gnd.n4639 gnd.n3378 9.3005
R18247 gnd.n4641 gnd.n4640 9.3005
R18248 gnd.n4642 gnd.n3359 9.3005
R18249 gnd.n4660 gnd.n4659 9.3005
R18250 gnd.n3360 gnd.n2029 9.3005
R18251 gnd.n4063 gnd.n4062 9.3005
R18252 gnd.n4716 gnd.n2030 9.3005
R18253 gnd.n4715 gnd.n2032 9.3005
R18254 gnd.n4712 gnd.n2033 9.3005
R18255 gnd.n4711 gnd.n2034 9.3005
R18256 gnd.n4708 gnd.n2035 9.3005
R18257 gnd.n4707 gnd.n2036 9.3005
R18258 gnd.n4704 gnd.n2037 9.3005
R18259 gnd.n4703 gnd.n2038 9.3005
R18260 gnd.n4700 gnd.n2039 9.3005
R18261 gnd.n4699 gnd.n2040 9.3005
R18262 gnd.n4696 gnd.n2041 9.3005
R18263 gnd.n4695 gnd.n2042 9.3005
R18264 gnd.n4692 gnd.n2043 9.3005
R18265 gnd.n4691 gnd.n2044 9.3005
R18266 gnd.n4688 gnd.n2045 9.3005
R18267 gnd.n4687 gnd.n2046 9.3005
R18268 gnd.n4684 gnd.n2047 9.3005
R18269 gnd.n4683 gnd.n2048 9.3005
R18270 gnd.n4680 gnd.n2049 9.3005
R18271 gnd.n4679 gnd.n2050 9.3005
R18272 gnd.n4676 gnd.n2051 9.3005
R18273 gnd.n4675 gnd.n2052 9.3005
R18274 gnd.n4672 gnd.n2056 9.3005
R18275 gnd.n4671 gnd.n2057 9.3005
R18276 gnd.n4668 gnd.n2058 9.3005
R18277 gnd.n4667 gnd.n2059 9.3005
R18278 gnd.n4718 gnd.n4717 9.3005
R18279 gnd.n3609 gnd.n3535 9.3005
R18280 gnd.n3607 gnd.n3536 9.3005
R18281 gnd.n3606 gnd.n3537 9.3005
R18282 gnd.n3603 gnd.n3538 9.3005
R18283 gnd.n3602 gnd.n3539 9.3005
R18284 gnd.n3601 gnd.n3540 9.3005
R18285 gnd.n3599 gnd.n3541 9.3005
R18286 gnd.n3598 gnd.n3542 9.3005
R18287 gnd.n3595 gnd.n3543 9.3005
R18288 gnd.n3594 gnd.n3544 9.3005
R18289 gnd.n3593 gnd.n3545 9.3005
R18290 gnd.n3591 gnd.n3546 9.3005
R18291 gnd.n3590 gnd.n3547 9.3005
R18292 gnd.n3585 gnd.n3548 9.3005
R18293 gnd.n3584 gnd.n3549 9.3005
R18294 gnd.n3583 gnd.n3550 9.3005
R18295 gnd.n3581 gnd.n3551 9.3005
R18296 gnd.n3580 gnd.n3552 9.3005
R18297 gnd.n3577 gnd.n3553 9.3005
R18298 gnd.n3576 gnd.n3554 9.3005
R18299 gnd.n3575 gnd.n3555 9.3005
R18300 gnd.n3573 gnd.n3556 9.3005
R18301 gnd.n3572 gnd.n3557 9.3005
R18302 gnd.n3569 gnd.n3558 9.3005
R18303 gnd.n3568 gnd.n3559 9.3005
R18304 gnd.n3567 gnd.n3560 9.3005
R18305 gnd.n3565 gnd.n3561 9.3005
R18306 gnd.n3564 gnd.n3563 9.3005
R18307 gnd.n3562 gnd.n2061 9.3005
R18308 gnd.n3973 gnd.n3972 9.3005
R18309 gnd.n3863 gnd.n3862 9.3005
R18310 gnd.n3987 gnd.n3986 9.3005
R18311 gnd.n3988 gnd.n3861 9.3005
R18312 gnd.n3990 gnd.n3989 9.3005
R18313 gnd.n3851 gnd.n3850 9.3005
R18314 gnd.n4003 gnd.n4002 9.3005
R18315 gnd.n4004 gnd.n3849 9.3005
R18316 gnd.n4036 gnd.n4005 9.3005
R18317 gnd.n4035 gnd.n4006 9.3005
R18318 gnd.n4034 gnd.n4007 9.3005
R18319 gnd.n4033 gnd.n4008 9.3005
R18320 gnd.n4030 gnd.n4009 9.3005
R18321 gnd.n4029 gnd.n4010 9.3005
R18322 gnd.n4028 gnd.n4011 9.3005
R18323 gnd.n4026 gnd.n4012 9.3005
R18324 gnd.n4025 gnd.n4013 9.3005
R18325 gnd.n4022 gnd.n4014 9.3005
R18326 gnd.n4021 gnd.n4015 9.3005
R18327 gnd.n4020 gnd.n4016 9.3005
R18328 gnd.n4018 gnd.n4017 9.3005
R18329 gnd.n3716 gnd.n3715 9.3005
R18330 gnd.n4140 gnd.n4139 9.3005
R18331 gnd.n4141 gnd.n3714 9.3005
R18332 gnd.n4145 gnd.n4142 9.3005
R18333 gnd.n4144 gnd.n4143 9.3005
R18334 gnd.n3679 gnd.n3678 9.3005
R18335 gnd.n4188 gnd.n4187 9.3005
R18336 gnd.n3971 gnd.n3872 9.3005
R18337 gnd.n3874 gnd.n3873 9.3005
R18338 gnd.n3918 gnd.n3916 9.3005
R18339 gnd.n3919 gnd.n3915 9.3005
R18340 gnd.n3922 gnd.n3911 9.3005
R18341 gnd.n3923 gnd.n3910 9.3005
R18342 gnd.n3926 gnd.n3909 9.3005
R18343 gnd.n3927 gnd.n3908 9.3005
R18344 gnd.n3930 gnd.n3907 9.3005
R18345 gnd.n3931 gnd.n3906 9.3005
R18346 gnd.n3934 gnd.n3905 9.3005
R18347 gnd.n3935 gnd.n3904 9.3005
R18348 gnd.n3938 gnd.n3903 9.3005
R18349 gnd.n3939 gnd.n3902 9.3005
R18350 gnd.n3942 gnd.n3901 9.3005
R18351 gnd.n3943 gnd.n3900 9.3005
R18352 gnd.n3946 gnd.n3899 9.3005
R18353 gnd.n3947 gnd.n3898 9.3005
R18354 gnd.n3950 gnd.n3897 9.3005
R18355 gnd.n3951 gnd.n3896 9.3005
R18356 gnd.n3954 gnd.n3895 9.3005
R18357 gnd.n3955 gnd.n3894 9.3005
R18358 gnd.n3958 gnd.n3893 9.3005
R18359 gnd.n3960 gnd.n3892 9.3005
R18360 gnd.n3961 gnd.n3891 9.3005
R18361 gnd.n3962 gnd.n3890 9.3005
R18362 gnd.n3963 gnd.n3889 9.3005
R18363 gnd.n3970 gnd.n3969 9.3005
R18364 gnd.n3979 gnd.n3978 9.3005
R18365 gnd.n3980 gnd.n3866 9.3005
R18366 gnd.n3982 gnd.n3981 9.3005
R18367 gnd.n3857 gnd.n3856 9.3005
R18368 gnd.n3995 gnd.n3994 9.3005
R18369 gnd.n3996 gnd.n3855 9.3005
R18370 gnd.n3998 gnd.n3997 9.3005
R18371 gnd.n3844 gnd.n3843 9.3005
R18372 gnd.n4041 gnd.n4040 9.3005
R18373 gnd.n4042 gnd.n3798 9.3005
R18374 gnd.n4046 gnd.n4044 9.3005
R18375 gnd.n4045 gnd.n3777 9.3005
R18376 gnd.n4064 gnd.n3776 9.3005
R18377 gnd.n4067 gnd.n4066 9.3005
R18378 gnd.n3770 gnd.n3769 9.3005
R18379 gnd.n4078 gnd.n4076 9.3005
R18380 gnd.n4077 gnd.n3751 9.3005
R18381 gnd.n4095 gnd.n3750 9.3005
R18382 gnd.n4098 gnd.n4097 9.3005
R18383 gnd.n3745 gnd.n3740 9.3005
R18384 gnd.n4108 gnd.n4107 9.3005
R18385 gnd.n3743 gnd.n3721 9.3005
R18386 gnd.n4135 gnd.n3722 9.3005
R18387 gnd.n4134 gnd.n4133 9.3005
R18388 gnd.n3724 gnd.n3709 9.3005
R18389 gnd.n4152 gnd.n4151 9.3005
R18390 gnd.n4154 gnd.n3687 9.3005
R18391 gnd.n4183 gnd.n3688 9.3005
R18392 gnd.n4182 gnd.n3689 9.3005
R18393 gnd.n4181 gnd.n3690 9.3005
R18394 gnd.n3693 gnd.n3692 9.3005
R18395 gnd.n3527 gnd.n3526 9.3005
R18396 gnd.n4203 gnd.n4201 9.3005
R18397 gnd.n4202 gnd.n3511 9.3005
R18398 gnd.n4220 gnd.n3510 9.3005
R18399 gnd.n4223 gnd.n4222 9.3005
R18400 gnd.n3504 gnd.n3503 9.3005
R18401 gnd.n4234 gnd.n4232 9.3005
R18402 gnd.n4233 gnd.n3486 9.3005
R18403 gnd.n4251 gnd.n3485 9.3005
R18404 gnd.n4254 gnd.n4253 9.3005
R18405 gnd.n3478 gnd.n3477 9.3005
R18406 gnd.n4265 gnd.n4263 9.3005
R18407 gnd.n4264 gnd.n3459 9.3005
R18408 gnd.n4282 gnd.n3458 9.3005
R18409 gnd.n4285 gnd.n4284 9.3005
R18410 gnd.n3452 gnd.n3451 9.3005
R18411 gnd.n4296 gnd.n4294 9.3005
R18412 gnd.n4295 gnd.n3435 9.3005
R18413 gnd.n4313 gnd.n3434 9.3005
R18414 gnd.n4316 gnd.n4315 9.3005
R18415 gnd.n3428 gnd.n3427 9.3005
R18416 gnd.n4327 gnd.n4325 9.3005
R18417 gnd.n4326 gnd.n3409 9.3005
R18418 gnd.n4344 gnd.n3408 9.3005
R18419 gnd.n4347 gnd.n4346 9.3005
R18420 gnd.n3402 gnd.n3401 9.3005
R18421 gnd.n4358 gnd.n4356 9.3005
R18422 gnd.n4357 gnd.n3384 9.3005
R18423 gnd.n4375 gnd.n3383 9.3005
R18424 gnd.n4634 gnd.n4633 9.3005
R18425 gnd.n3376 gnd.n3375 9.3005
R18426 gnd.n4644 gnd.n4643 9.3005
R18427 gnd.n3358 gnd.n3357 9.3005
R18428 gnd.n4662 gnd.n4661 9.3005
R18429 gnd.n3868 gnd.n3867 9.3005
R18430 gnd.n3139 gnd.n3138 9.3005
R18431 gnd.n3137 gnd.n2191 9.3005
R18432 gnd.n3136 gnd.n3135 9.3005
R18433 gnd.n2193 gnd.n2192 9.3005
R18434 gnd.n3129 gnd.n2197 9.3005
R18435 gnd.n3128 gnd.n2198 9.3005
R18436 gnd.n3127 gnd.n2199 9.3005
R18437 gnd.n2204 gnd.n2200 9.3005
R18438 gnd.n3121 gnd.n2205 9.3005
R18439 gnd.n3120 gnd.n2206 9.3005
R18440 gnd.n3119 gnd.n2207 9.3005
R18441 gnd.n2212 gnd.n2208 9.3005
R18442 gnd.n3113 gnd.n2213 9.3005
R18443 gnd.n3112 gnd.n2214 9.3005
R18444 gnd.n3111 gnd.n2215 9.3005
R18445 gnd.n2220 gnd.n2216 9.3005
R18446 gnd.n3105 gnd.n2221 9.3005
R18447 gnd.n3104 gnd.n2222 9.3005
R18448 gnd.n3103 gnd.n2223 9.3005
R18449 gnd.n2228 gnd.n2224 9.3005
R18450 gnd.n3097 gnd.n2229 9.3005
R18451 gnd.n3096 gnd.n2230 9.3005
R18452 gnd.n3095 gnd.n2231 9.3005
R18453 gnd.n2236 gnd.n2232 9.3005
R18454 gnd.n3089 gnd.n2237 9.3005
R18455 gnd.n3088 gnd.n2238 9.3005
R18456 gnd.n3087 gnd.n2239 9.3005
R18457 gnd.n2244 gnd.n2240 9.3005
R18458 gnd.n3081 gnd.n2245 9.3005
R18459 gnd.n3080 gnd.n2246 9.3005
R18460 gnd.n3079 gnd.n2247 9.3005
R18461 gnd.n2252 gnd.n2248 9.3005
R18462 gnd.n3073 gnd.n2253 9.3005
R18463 gnd.n3072 gnd.n2254 9.3005
R18464 gnd.n3071 gnd.n2255 9.3005
R18465 gnd.n2260 gnd.n2256 9.3005
R18466 gnd.n3065 gnd.n2261 9.3005
R18467 gnd.n3064 gnd.n2262 9.3005
R18468 gnd.n3063 gnd.n2263 9.3005
R18469 gnd.n2268 gnd.n2264 9.3005
R18470 gnd.n3057 gnd.n2269 9.3005
R18471 gnd.n3056 gnd.n2270 9.3005
R18472 gnd.n3055 gnd.n2271 9.3005
R18473 gnd.n2276 gnd.n2272 9.3005
R18474 gnd.n3049 gnd.n2277 9.3005
R18475 gnd.n3048 gnd.n2278 9.3005
R18476 gnd.n3047 gnd.n2279 9.3005
R18477 gnd.n2284 gnd.n2280 9.3005
R18478 gnd.n3041 gnd.n2285 9.3005
R18479 gnd.n3040 gnd.n2286 9.3005
R18480 gnd.n3039 gnd.n2287 9.3005
R18481 gnd.n2292 gnd.n2288 9.3005
R18482 gnd.n3033 gnd.n2293 9.3005
R18483 gnd.n3032 gnd.n2294 9.3005
R18484 gnd.n3031 gnd.n2295 9.3005
R18485 gnd.n2300 gnd.n2296 9.3005
R18486 gnd.n3025 gnd.n2301 9.3005
R18487 gnd.n3024 gnd.n2302 9.3005
R18488 gnd.n3023 gnd.n2303 9.3005
R18489 gnd.n2308 gnd.n2304 9.3005
R18490 gnd.n3017 gnd.n2309 9.3005
R18491 gnd.n3016 gnd.n2310 9.3005
R18492 gnd.n3015 gnd.n2311 9.3005
R18493 gnd.n2316 gnd.n2312 9.3005
R18494 gnd.n3009 gnd.n2317 9.3005
R18495 gnd.n3008 gnd.n2318 9.3005
R18496 gnd.n3007 gnd.n2319 9.3005
R18497 gnd.n2324 gnd.n2320 9.3005
R18498 gnd.n3001 gnd.n2325 9.3005
R18499 gnd.n3000 gnd.n2326 9.3005
R18500 gnd.n2999 gnd.n2327 9.3005
R18501 gnd.n2332 gnd.n2328 9.3005
R18502 gnd.n2993 gnd.n2333 9.3005
R18503 gnd.n2992 gnd.n2334 9.3005
R18504 gnd.n2991 gnd.n2335 9.3005
R18505 gnd.n2340 gnd.n2336 9.3005
R18506 gnd.n2985 gnd.n2341 9.3005
R18507 gnd.n2984 gnd.n2342 9.3005
R18508 gnd.n2983 gnd.n2343 9.3005
R18509 gnd.n2348 gnd.n2344 9.3005
R18510 gnd.n2977 gnd.n2349 9.3005
R18511 gnd.n2976 gnd.n2350 9.3005
R18512 gnd.n2975 gnd.n2351 9.3005
R18513 gnd.n2356 gnd.n2352 9.3005
R18514 gnd.n2969 gnd.n2357 9.3005
R18515 gnd.n2968 gnd.n2358 9.3005
R18516 gnd.n2967 gnd.n2359 9.3005
R18517 gnd.n2364 gnd.n2360 9.3005
R18518 gnd.n2961 gnd.n2365 9.3005
R18519 gnd.n2960 gnd.n2366 9.3005
R18520 gnd.n2959 gnd.n2367 9.3005
R18521 gnd.n2372 gnd.n2368 9.3005
R18522 gnd.n2953 gnd.n2373 9.3005
R18523 gnd.n2952 gnd.n2374 9.3005
R18524 gnd.n2951 gnd.n2375 9.3005
R18525 gnd.n2380 gnd.n2376 9.3005
R18526 gnd.n2945 gnd.n2381 9.3005
R18527 gnd.n2944 gnd.n2382 9.3005
R18528 gnd.n2943 gnd.n2383 9.3005
R18529 gnd.n2388 gnd.n2384 9.3005
R18530 gnd.n2937 gnd.n2389 9.3005
R18531 gnd.n2936 gnd.n2390 9.3005
R18532 gnd.n2935 gnd.n2391 9.3005
R18533 gnd.n2396 gnd.n2392 9.3005
R18534 gnd.n2929 gnd.n2397 9.3005
R18535 gnd.n2928 gnd.n2398 9.3005
R18536 gnd.n2927 gnd.n2399 9.3005
R18537 gnd.n2404 gnd.n2400 9.3005
R18538 gnd.n2921 gnd.n2405 9.3005
R18539 gnd.n2920 gnd.n2406 9.3005
R18540 gnd.n2919 gnd.n2407 9.3005
R18541 gnd.n2412 gnd.n2408 9.3005
R18542 gnd.n2913 gnd.n2413 9.3005
R18543 gnd.n2912 gnd.n2414 9.3005
R18544 gnd.n2911 gnd.n2415 9.3005
R18545 gnd.n2420 gnd.n2416 9.3005
R18546 gnd.n2905 gnd.n2421 9.3005
R18547 gnd.n2904 gnd.n2422 9.3005
R18548 gnd.n2903 gnd.n2423 9.3005
R18549 gnd.n2428 gnd.n2424 9.3005
R18550 gnd.n2897 gnd.n2429 9.3005
R18551 gnd.n2896 gnd.n2430 9.3005
R18552 gnd.n2895 gnd.n2431 9.3005
R18553 gnd.n2436 gnd.n2432 9.3005
R18554 gnd.n2889 gnd.n2437 9.3005
R18555 gnd.n2888 gnd.n2438 9.3005
R18556 gnd.n2887 gnd.n2439 9.3005
R18557 gnd.n2444 gnd.n2440 9.3005
R18558 gnd.n2881 gnd.n2445 9.3005
R18559 gnd.n2880 gnd.n2446 9.3005
R18560 gnd.n2879 gnd.n2447 9.3005
R18561 gnd.n2452 gnd.n2448 9.3005
R18562 gnd.n2873 gnd.n2453 9.3005
R18563 gnd.n2872 gnd.n2454 9.3005
R18564 gnd.n2871 gnd.n2455 9.3005
R18565 gnd.n2460 gnd.n2456 9.3005
R18566 gnd.n2865 gnd.n2461 9.3005
R18567 gnd.n2864 gnd.n2462 9.3005
R18568 gnd.n2863 gnd.n2463 9.3005
R18569 gnd.n2468 gnd.n2464 9.3005
R18570 gnd.n2857 gnd.n2469 9.3005
R18571 gnd.n2856 gnd.n2470 9.3005
R18572 gnd.n2855 gnd.n2471 9.3005
R18573 gnd.n2476 gnd.n2472 9.3005
R18574 gnd.n2849 gnd.n2477 9.3005
R18575 gnd.n2848 gnd.n2478 9.3005
R18576 gnd.n2847 gnd.n2479 9.3005
R18577 gnd.n2484 gnd.n2480 9.3005
R18578 gnd.n2841 gnd.n2485 9.3005
R18579 gnd.n2840 gnd.n2486 9.3005
R18580 gnd.n2839 gnd.n2487 9.3005
R18581 gnd.n2492 gnd.n2488 9.3005
R18582 gnd.n2833 gnd.n2493 9.3005
R18583 gnd.n2832 gnd.n2494 9.3005
R18584 gnd.n2831 gnd.n2495 9.3005
R18585 gnd.n2825 gnd.n2824 9.3005
R18586 gnd.n2823 gnd.n2500 9.3005
R18587 gnd.n2822 gnd.n2821 9.3005
R18588 gnd.n2503 gnd.n2502 9.3005
R18589 gnd.n2815 gnd.n2507 9.3005
R18590 gnd.n2814 gnd.n2508 9.3005
R18591 gnd.n2813 gnd.n2509 9.3005
R18592 gnd.n2514 gnd.n2510 9.3005
R18593 gnd.n2807 gnd.n2515 9.3005
R18594 gnd.n2806 gnd.n2516 9.3005
R18595 gnd.n2805 gnd.n2517 9.3005
R18596 gnd.n2522 gnd.n2518 9.3005
R18597 gnd.n2799 gnd.n2523 9.3005
R18598 gnd.n2798 gnd.n2524 9.3005
R18599 gnd.n2797 gnd.n2525 9.3005
R18600 gnd.n2530 gnd.n2526 9.3005
R18601 gnd.n2791 gnd.n2531 9.3005
R18602 gnd.n2790 gnd.n2532 9.3005
R18603 gnd.n2789 gnd.n2533 9.3005
R18604 gnd.n2538 gnd.n2534 9.3005
R18605 gnd.n2783 gnd.n2539 9.3005
R18606 gnd.n2782 gnd.n2540 9.3005
R18607 gnd.n2781 gnd.n2541 9.3005
R18608 gnd.n2546 gnd.n2542 9.3005
R18609 gnd.n2775 gnd.n2547 9.3005
R18610 gnd.n2774 gnd.n2548 9.3005
R18611 gnd.n2773 gnd.n2549 9.3005
R18612 gnd.n2554 gnd.n2550 9.3005
R18613 gnd.n2767 gnd.n2555 9.3005
R18614 gnd.n2766 gnd.n2556 9.3005
R18615 gnd.n2765 gnd.n2557 9.3005
R18616 gnd.n2562 gnd.n2558 9.3005
R18617 gnd.n2759 gnd.n2563 9.3005
R18618 gnd.n2758 gnd.n2564 9.3005
R18619 gnd.n2757 gnd.n2565 9.3005
R18620 gnd.n2570 gnd.n2566 9.3005
R18621 gnd.n2751 gnd.n2571 9.3005
R18622 gnd.n2750 gnd.n2572 9.3005
R18623 gnd.n2749 gnd.n2573 9.3005
R18624 gnd.n2578 gnd.n2574 9.3005
R18625 gnd.n2743 gnd.n2579 9.3005
R18626 gnd.n2742 gnd.n2580 9.3005
R18627 gnd.n2741 gnd.n2581 9.3005
R18628 gnd.n2586 gnd.n2582 9.3005
R18629 gnd.n2735 gnd.n2587 9.3005
R18630 gnd.n2734 gnd.n2588 9.3005
R18631 gnd.n2733 gnd.n2589 9.3005
R18632 gnd.n2594 gnd.n2590 9.3005
R18633 gnd.n2727 gnd.n2595 9.3005
R18634 gnd.n2726 gnd.n2596 9.3005
R18635 gnd.n2725 gnd.n2597 9.3005
R18636 gnd.n2602 gnd.n2598 9.3005
R18637 gnd.n2719 gnd.n2603 9.3005
R18638 gnd.n2718 gnd.n2604 9.3005
R18639 gnd.n2717 gnd.n2605 9.3005
R18640 gnd.n2610 gnd.n2606 9.3005
R18641 gnd.n2711 gnd.n2611 9.3005
R18642 gnd.n2710 gnd.n2612 9.3005
R18643 gnd.n2709 gnd.n2613 9.3005
R18644 gnd.n2618 gnd.n2614 9.3005
R18645 gnd.n2703 gnd.n2619 9.3005
R18646 gnd.n2702 gnd.n2620 9.3005
R18647 gnd.n2701 gnd.n2621 9.3005
R18648 gnd.n2626 gnd.n2622 9.3005
R18649 gnd.n2695 gnd.n2627 9.3005
R18650 gnd.n2694 gnd.n2628 9.3005
R18651 gnd.n2693 gnd.n2629 9.3005
R18652 gnd.n2634 gnd.n2630 9.3005
R18653 gnd.n2687 gnd.n2635 9.3005
R18654 gnd.n2686 gnd.n2636 9.3005
R18655 gnd.n2685 gnd.n2637 9.3005
R18656 gnd.n2642 gnd.n2638 9.3005
R18657 gnd.n2679 gnd.n2643 9.3005
R18658 gnd.n2678 gnd.n2644 9.3005
R18659 gnd.n2677 gnd.n2645 9.3005
R18660 gnd.n2650 gnd.n2646 9.3005
R18661 gnd.n2671 gnd.n2651 9.3005
R18662 gnd.n2670 gnd.n2652 9.3005
R18663 gnd.n2669 gnd.n2653 9.3005
R18664 gnd.n2659 gnd.n2654 9.3005
R18665 gnd.n2663 gnd.n2660 9.3005
R18666 gnd.n2662 gnd.n2661 9.3005
R18667 gnd.n345 gnd.n344 9.3005
R18668 gnd.n7219 gnd.n7218 9.3005
R18669 gnd.n2501 gnd.n2499 9.3005
R18670 gnd.n7567 gnd.n130 9.3005
R18671 gnd.n7566 gnd.n132 9.3005
R18672 gnd.n136 gnd.n133 9.3005
R18673 gnd.n7561 gnd.n137 9.3005
R18674 gnd.n7560 gnd.n138 9.3005
R18675 gnd.n7559 gnd.n139 9.3005
R18676 gnd.n143 gnd.n140 9.3005
R18677 gnd.n7554 gnd.n144 9.3005
R18678 gnd.n7553 gnd.n145 9.3005
R18679 gnd.n7552 gnd.n146 9.3005
R18680 gnd.n150 gnd.n147 9.3005
R18681 gnd.n7547 gnd.n151 9.3005
R18682 gnd.n7546 gnd.n152 9.3005
R18683 gnd.n7545 gnd.n153 9.3005
R18684 gnd.n157 gnd.n154 9.3005
R18685 gnd.n7540 gnd.n158 9.3005
R18686 gnd.n7539 gnd.n159 9.3005
R18687 gnd.n7535 gnd.n160 9.3005
R18688 gnd.n164 gnd.n161 9.3005
R18689 gnd.n7530 gnd.n165 9.3005
R18690 gnd.n7529 gnd.n166 9.3005
R18691 gnd.n7528 gnd.n167 9.3005
R18692 gnd.n171 gnd.n168 9.3005
R18693 gnd.n7523 gnd.n172 9.3005
R18694 gnd.n7522 gnd.n173 9.3005
R18695 gnd.n7521 gnd.n174 9.3005
R18696 gnd.n178 gnd.n175 9.3005
R18697 gnd.n7516 gnd.n179 9.3005
R18698 gnd.n7515 gnd.n180 9.3005
R18699 gnd.n7514 gnd.n181 9.3005
R18700 gnd.n185 gnd.n182 9.3005
R18701 gnd.n7509 gnd.n186 9.3005
R18702 gnd.n7508 gnd.n187 9.3005
R18703 gnd.n7507 gnd.n188 9.3005
R18704 gnd.n192 gnd.n189 9.3005
R18705 gnd.n7502 gnd.n193 9.3005
R18706 gnd.n7501 gnd.n7500 9.3005
R18707 gnd.n7499 gnd.n196 9.3005
R18708 gnd.n7569 gnd.n7568 9.3005
R18709 gnd.n6844 gnd.n6843 9.3005
R18710 gnd.n6848 gnd.n6845 9.3005
R18711 gnd.n6849 gnd.n6842 9.3005
R18712 gnd.n6853 gnd.n6852 9.3005
R18713 gnd.n6854 gnd.n6841 9.3005
R18714 gnd.n6863 gnd.n6855 9.3005
R18715 gnd.n6862 gnd.n6856 9.3005
R18716 gnd.n6861 gnd.n6858 9.3005
R18717 gnd.n6857 gnd.n596 9.3005
R18718 gnd.n6888 gnd.n597 9.3005
R18719 gnd.n6889 gnd.n595 9.3005
R18720 gnd.n6893 gnd.n6892 9.3005
R18721 gnd.n6894 gnd.n594 9.3005
R18722 gnd.n6902 gnd.n6895 9.3005
R18723 gnd.n6901 gnd.n6896 9.3005
R18724 gnd.n6900 gnd.n6897 9.3005
R18725 gnd.n587 gnd.n586 9.3005
R18726 gnd.n6920 gnd.n6919 9.3005
R18727 gnd.n6921 gnd.n585 9.3005
R18728 gnd.n6936 gnd.n6922 9.3005
R18729 gnd.n6935 gnd.n6923 9.3005
R18730 gnd.n6934 gnd.n6924 9.3005
R18731 gnd.n6933 gnd.n6925 9.3005
R18732 gnd.n6932 gnd.n6926 9.3005
R18733 gnd.n6929 gnd.n6928 9.3005
R18734 gnd.n6927 gnd.n357 9.3005
R18735 gnd.n7193 gnd.n356 9.3005
R18736 gnd.n7195 gnd.n7194 9.3005
R18737 gnd.n7196 gnd.n355 9.3005
R18738 gnd.n7200 gnd.n7197 9.3005
R18739 gnd.n7199 gnd.n7198 9.3005
R18740 gnd.n334 gnd.n333 9.3005
R18741 gnd.n7231 gnd.n7230 9.3005
R18742 gnd.n7232 gnd.n332 9.3005
R18743 gnd.n7299 gnd.n7233 9.3005
R18744 gnd.n7298 gnd.n7234 9.3005
R18745 gnd.n7297 gnd.n7235 9.3005
R18746 gnd.n7295 gnd.n7236 9.3005
R18747 gnd.n7294 gnd.n7237 9.3005
R18748 gnd.n7292 gnd.n7238 9.3005
R18749 gnd.n7291 gnd.n7239 9.3005
R18750 gnd.n7289 gnd.n7240 9.3005
R18751 gnd.n7288 gnd.n7241 9.3005
R18752 gnd.n7286 gnd.n7242 9.3005
R18753 gnd.n7285 gnd.n7243 9.3005
R18754 gnd.n7283 gnd.n7244 9.3005
R18755 gnd.n7282 gnd.n7245 9.3005
R18756 gnd.n7280 gnd.n7246 9.3005
R18757 gnd.n7279 gnd.n7247 9.3005
R18758 gnd.n7277 gnd.n7248 9.3005
R18759 gnd.n7276 gnd.n7249 9.3005
R18760 gnd.n7274 gnd.n7250 9.3005
R18761 gnd.n7273 gnd.n7251 9.3005
R18762 gnd.n7271 gnd.n7252 9.3005
R18763 gnd.n7270 gnd.n7253 9.3005
R18764 gnd.n7268 gnd.n7254 9.3005
R18765 gnd.n7267 gnd.n7255 9.3005
R18766 gnd.n7265 gnd.n7256 9.3005
R18767 gnd.n7264 gnd.n7257 9.3005
R18768 gnd.n7262 gnd.n7258 9.3005
R18769 gnd.n7261 gnd.n7260 9.3005
R18770 gnd.n7259 gnd.n200 9.3005
R18771 gnd.n7496 gnd.n199 9.3005
R18772 gnd.n7498 gnd.n7497 9.3005
R18773 gnd.n563 gnd.n562 9.3005
R18774 gnd.n6981 gnd.n6980 9.3005
R18775 gnd.n6982 gnd.n556 9.3005
R18776 gnd.n6985 gnd.n555 9.3005
R18777 gnd.n6986 gnd.n554 9.3005
R18778 gnd.n6989 gnd.n553 9.3005
R18779 gnd.n6990 gnd.n552 9.3005
R18780 gnd.n6993 gnd.n551 9.3005
R18781 gnd.n6994 gnd.n550 9.3005
R18782 gnd.n6997 gnd.n549 9.3005
R18783 gnd.n6998 gnd.n548 9.3005
R18784 gnd.n7001 gnd.n547 9.3005
R18785 gnd.n7002 gnd.n546 9.3005
R18786 gnd.n7005 gnd.n545 9.3005
R18787 gnd.n7006 gnd.n544 9.3005
R18788 gnd.n7009 gnd.n543 9.3005
R18789 gnd.n7010 gnd.n542 9.3005
R18790 gnd.n7013 gnd.n541 9.3005
R18791 gnd.n7014 gnd.n540 9.3005
R18792 gnd.n7017 gnd.n539 9.3005
R18793 gnd.n7019 gnd.n533 9.3005
R18794 gnd.n7022 gnd.n532 9.3005
R18795 gnd.n7023 gnd.n531 9.3005
R18796 gnd.n7026 gnd.n530 9.3005
R18797 gnd.n7027 gnd.n529 9.3005
R18798 gnd.n7030 gnd.n528 9.3005
R18799 gnd.n7031 gnd.n527 9.3005
R18800 gnd.n7034 gnd.n526 9.3005
R18801 gnd.n7035 gnd.n525 9.3005
R18802 gnd.n7038 gnd.n524 9.3005
R18803 gnd.n7039 gnd.n523 9.3005
R18804 gnd.n7042 gnd.n522 9.3005
R18805 gnd.n7043 gnd.n521 9.3005
R18806 gnd.n7044 gnd.n520 9.3005
R18807 gnd.n487 gnd.n486 9.3005
R18808 gnd.n7050 gnd.n7049 9.3005
R18809 gnd.n6979 gnd.n561 9.3005
R18810 gnd.n6978 gnd.n6977 9.3005
R18811 gnd.n7053 gnd.n7052 9.3005
R18812 gnd.n469 gnd.n468 9.3005
R18813 gnd.n7066 gnd.n7065 9.3005
R18814 gnd.n7067 gnd.n467 9.3005
R18815 gnd.n7069 gnd.n7068 9.3005
R18816 gnd.n452 gnd.n451 9.3005
R18817 gnd.n7082 gnd.n7081 9.3005
R18818 gnd.n7083 gnd.n450 9.3005
R18819 gnd.n7085 gnd.n7084 9.3005
R18820 gnd.n435 gnd.n434 9.3005
R18821 gnd.n7098 gnd.n7097 9.3005
R18822 gnd.n7099 gnd.n433 9.3005
R18823 gnd.n7101 gnd.n7100 9.3005
R18824 gnd.n418 gnd.n417 9.3005
R18825 gnd.n7114 gnd.n7113 9.3005
R18826 gnd.n7115 gnd.n416 9.3005
R18827 gnd.n7117 gnd.n7116 9.3005
R18828 gnd.n399 gnd.n398 9.3005
R18829 gnd.n7133 gnd.n7132 9.3005
R18830 gnd.n7134 gnd.n397 9.3005
R18831 gnd.n7136 gnd.n7135 9.3005
R18832 gnd.n367 gnd.n366 9.3005
R18833 gnd.n7184 gnd.n7183 9.3005
R18834 gnd.n7185 gnd.n365 9.3005
R18835 gnd.n7187 gnd.n7186 9.3005
R18836 gnd.n7188 gnd.n299 9.3005
R18837 gnd.n7327 gnd.n7326 9.3005
R18838 gnd.n284 gnd.n283 9.3005
R18839 gnd.n7340 gnd.n7339 9.3005
R18840 gnd.n7341 gnd.n282 9.3005
R18841 gnd.n7343 gnd.n7342 9.3005
R18842 gnd.n270 gnd.n269 9.3005
R18843 gnd.n7356 gnd.n7355 9.3005
R18844 gnd.n7357 gnd.n268 9.3005
R18845 gnd.n7359 gnd.n7358 9.3005
R18846 gnd.n254 gnd.n253 9.3005
R18847 gnd.n7372 gnd.n7371 9.3005
R18848 gnd.n7373 gnd.n252 9.3005
R18849 gnd.n7375 gnd.n7374 9.3005
R18850 gnd.n240 gnd.n239 9.3005
R18851 gnd.n7388 gnd.n7387 9.3005
R18852 gnd.n7389 gnd.n238 9.3005
R18853 gnd.n7391 gnd.n7390 9.3005
R18854 gnd.n223 gnd.n222 9.3005
R18855 gnd.n7404 gnd.n7403 9.3005
R18856 gnd.n7405 gnd.n221 9.3005
R18857 gnd.n7407 gnd.n7406 9.3005
R18858 gnd.n207 gnd.n206 9.3005
R18859 gnd.n7488 gnd.n7487 9.3005
R18860 gnd.n7489 gnd.n205 9.3005
R18861 gnd.n7491 gnd.n7490 9.3005
R18862 gnd.n129 gnd.n128 9.3005
R18863 gnd.n7571 gnd.n7570 9.3005
R18864 gnd.n7051 gnd.n485 9.3005
R18865 gnd.n7325 gnd.n298 9.3005
R18866 gnd.n7148 gnd.n346 9.3005
R18867 gnd.n7215 gnd.n347 9.3005
R18868 gnd.n7217 gnd.n7216 9.3005
R18869 gnd.n5433 gnd.n1803 9.3005
R18870 gnd.n5258 gnd.n1804 9.3005
R18871 gnd.n5260 gnd.n5259 9.3005
R18872 gnd.n5261 gnd.n5257 9.3005
R18873 gnd.n5273 gnd.n5262 9.3005
R18874 gnd.n5272 gnd.n5263 9.3005
R18875 gnd.n5271 gnd.n5264 9.3005
R18876 gnd.n5268 gnd.n5265 9.3005
R18877 gnd.n5267 gnd.n5266 9.3005
R18878 gnd.n1848 gnd.n1847 9.3005
R18879 gnd.n5300 gnd.n5299 9.3005
R18880 gnd.n5301 gnd.n1846 9.3005
R18881 gnd.n5313 gnd.n5302 9.3005
R18882 gnd.n5312 gnd.n5303 9.3005
R18883 gnd.n5311 gnd.n5304 9.3005
R18884 gnd.n5308 gnd.n5305 9.3005
R18885 gnd.n5307 gnd.n5306 9.3005
R18886 gnd.n1838 gnd.n1837 9.3005
R18887 gnd.n5339 gnd.n5338 9.3005
R18888 gnd.n5340 gnd.n1836 9.3005
R18889 gnd.n5370 gnd.n5341 9.3005
R18890 gnd.n5369 gnd.n5342 9.3005
R18891 gnd.n5368 gnd.n5343 9.3005
R18892 gnd.n5346 gnd.n5344 9.3005
R18893 gnd.n5364 gnd.n5347 9.3005
R18894 gnd.n5363 gnd.n5348 9.3005
R18895 gnd.n5362 gnd.n5349 9.3005
R18896 gnd.n5353 gnd.n5350 9.3005
R18897 gnd.n5357 gnd.n5354 9.3005
R18898 gnd.n5356 gnd.n5355 9.3005
R18899 gnd.n1316 gnd.n1315 9.3005
R18900 gnd.n5812 gnd.n5811 9.3005
R18901 gnd.n5813 gnd.n1314 9.3005
R18902 gnd.n5815 gnd.n5814 9.3005
R18903 gnd.n1302 gnd.n1301 9.3005
R18904 gnd.n5828 gnd.n5827 9.3005
R18905 gnd.n5829 gnd.n1300 9.3005
R18906 gnd.n5833 gnd.n5830 9.3005
R18907 gnd.n5832 gnd.n5831 9.3005
R18908 gnd.n1260 gnd.n1259 9.3005
R18909 gnd.n5986 gnd.n5985 9.3005
R18910 gnd.n5987 gnd.n1258 9.3005
R18911 gnd.n5989 gnd.n5988 9.3005
R18912 gnd.n1245 gnd.n1244 9.3005
R18913 gnd.n6002 gnd.n6001 9.3005
R18914 gnd.n6003 gnd.n1243 9.3005
R18915 gnd.n6005 gnd.n6004 9.3005
R18916 gnd.n1229 gnd.n1228 9.3005
R18917 gnd.n6018 gnd.n6017 9.3005
R18918 gnd.n6019 gnd.n1227 9.3005
R18919 gnd.n6021 gnd.n6020 9.3005
R18920 gnd.n1214 gnd.n1213 9.3005
R18921 gnd.n6033 gnd.n6032 9.3005
R18922 gnd.n6034 gnd.n1212 9.3005
R18923 gnd.n6038 gnd.n6035 9.3005
R18924 gnd.n6037 gnd.n6036 9.3005
R18925 gnd.n1107 gnd.n1106 9.3005
R18926 gnd.n6128 gnd.n6127 9.3005
R18927 gnd.n6129 gnd.n1105 9.3005
R18928 gnd.n6131 gnd.n6130 9.3005
R18929 gnd.n1091 gnd.n1090 9.3005
R18930 gnd.n6144 gnd.n6143 9.3005
R18931 gnd.n6145 gnd.n1089 9.3005
R18932 gnd.n6147 gnd.n6146 9.3005
R18933 gnd.n1076 gnd.n1075 9.3005
R18934 gnd.n6160 gnd.n6159 9.3005
R18935 gnd.n6161 gnd.n1074 9.3005
R18936 gnd.n6163 gnd.n6162 9.3005
R18937 gnd.n1063 gnd.n1062 9.3005
R18938 gnd.n6176 gnd.n6175 9.3005
R18939 gnd.n6177 gnd.n1061 9.3005
R18940 gnd.n6181 gnd.n6178 9.3005
R18941 gnd.n6180 gnd.n6179 9.3005
R18942 gnd.n1020 gnd.n1019 9.3005
R18943 gnd.n6433 gnd.n6432 9.3005
R18944 gnd.n6434 gnd.n1018 9.3005
R18945 gnd.n6436 gnd.n6435 9.3005
R18946 gnd.n1004 gnd.n1003 9.3005
R18947 gnd.n6449 gnd.n6448 9.3005
R18948 gnd.n6450 gnd.n1002 9.3005
R18949 gnd.n6452 gnd.n6451 9.3005
R18950 gnd.n988 gnd.n987 9.3005
R18951 gnd.n6465 gnd.n6464 9.3005
R18952 gnd.n6466 gnd.n986 9.3005
R18953 gnd.n6468 gnd.n6467 9.3005
R18954 gnd.n974 gnd.n973 9.3005
R18955 gnd.n6481 gnd.n6480 9.3005
R18956 gnd.n6482 gnd.n972 9.3005
R18957 gnd.n6484 gnd.n6483 9.3005
R18958 gnd.n959 gnd.n958 9.3005
R18959 gnd.n6497 gnd.n6496 9.3005
R18960 gnd.n6498 gnd.n957 9.3005
R18961 gnd.n6500 gnd.n6499 9.3005
R18962 gnd.n943 gnd.n942 9.3005
R18963 gnd.n6513 gnd.n6512 9.3005
R18964 gnd.n6514 gnd.n941 9.3005
R18965 gnd.n6516 gnd.n6515 9.3005
R18966 gnd.n926 gnd.n925 9.3005
R18967 gnd.n6535 gnd.n6534 9.3005
R18968 gnd.n6536 gnd.n924 9.3005
R18969 gnd.n6540 gnd.n6537 9.3005
R18970 gnd.n6539 gnd.n6538 9.3005
R18971 gnd.n886 gnd.n885 9.3005
R18972 gnd.n6593 gnd.n6592 9.3005
R18973 gnd.n6594 gnd.n884 9.3005
R18974 gnd.n6598 gnd.n6595 9.3005
R18975 gnd.n6597 gnd.n6596 9.3005
R18976 gnd.n659 gnd.n658 9.3005
R18977 gnd.n6784 gnd.n6783 9.3005
R18978 gnd.n6785 gnd.n657 9.3005
R18979 gnd.n6787 gnd.n6786 9.3005
R18980 gnd.n644 gnd.n643 9.3005
R18981 gnd.n6801 gnd.n6800 9.3005
R18982 gnd.n6802 gnd.n642 9.3005
R18983 gnd.n6806 gnd.n6803 9.3005
R18984 gnd.n6805 gnd.n6804 9.3005
R18985 gnd.n614 gnd.n613 9.3005
R18986 gnd.n6820 gnd.n6819 9.3005
R18987 gnd.n6821 gnd.n612 9.3005
R18988 gnd.n6823 gnd.n6822 9.3005
R18989 gnd.n610 gnd.n609 9.3005
R18990 gnd.n6828 gnd.n6827 9.3005
R18991 gnd.n6829 gnd.n608 9.3005
R18992 gnd.n6831 gnd.n6830 9.3005
R18993 gnd.n606 gnd.n605 9.3005
R18994 gnd.n6836 gnd.n6835 9.3005
R18995 gnd.n6837 gnd.n604 9.3005
R18996 gnd.n6839 gnd.n6838 9.3005
R18997 gnd.n602 gnd.n601 9.3005
R18998 gnd.n6870 gnd.n6869 9.3005
R18999 gnd.n6871 gnd.n600 9.3005
R19000 gnd.n6883 gnd.n6872 9.3005
R19001 gnd.n6882 gnd.n6873 9.3005
R19002 gnd.n6881 gnd.n6874 9.3005
R19003 gnd.n6878 gnd.n6875 9.3005
R19004 gnd.n6877 gnd.n6876 9.3005
R19005 gnd.n592 gnd.n591 9.3005
R19006 gnd.n6909 gnd.n6908 9.3005
R19007 gnd.n6910 gnd.n590 9.3005
R19008 gnd.n6914 gnd.n6911 9.3005
R19009 gnd.n6913 gnd.n6912 9.3005
R19010 gnd.n392 gnd.n391 9.3005
R19011 gnd.n7142 gnd.n7141 9.3005
R19012 gnd.n7143 gnd.n390 9.3005
R19013 gnd.n7156 gnd.n7144 9.3005
R19014 gnd.n7155 gnd.n7145 9.3005
R19015 gnd.n7154 gnd.n7146 9.3005
R19016 gnd.n7151 gnd.n7147 9.3005
R19017 gnd.n7150 gnd.n7149 9.3005
R19018 gnd.n5210 gnd.n5209 9.3005
R19019 gnd.n4870 gnd.n4827 9.3005
R19020 gnd.n4869 gnd.n4828 9.3005
R19021 gnd.n4868 gnd.n4829 9.3005
R19022 gnd.n4866 gnd.n4830 9.3005
R19023 gnd.n4865 gnd.n4831 9.3005
R19024 gnd.n4863 gnd.n4832 9.3005
R19025 gnd.n4862 gnd.n4833 9.3005
R19026 gnd.n4860 gnd.n4834 9.3005
R19027 gnd.n4859 gnd.n4835 9.3005
R19028 gnd.n4857 gnd.n4836 9.3005
R19029 gnd.n4856 gnd.n4837 9.3005
R19030 gnd.n4854 gnd.n4838 9.3005
R19031 gnd.n4853 gnd.n4839 9.3005
R19032 gnd.n4851 gnd.n4840 9.3005
R19033 gnd.n4850 gnd.n4841 9.3005
R19034 gnd.n4848 gnd.n4842 9.3005
R19035 gnd.n4847 gnd.n4843 9.3005
R19036 gnd.n4845 gnd.n4844 9.3005
R19037 gnd.n1906 gnd.n1905 9.3005
R19038 gnd.n5163 gnd.n5162 9.3005
R19039 gnd.n5164 gnd.n1904 9.3005
R19040 gnd.n5171 gnd.n5165 9.3005
R19041 gnd.n5170 gnd.n5166 9.3005
R19042 gnd.n5169 gnd.n5167 9.3005
R19043 gnd.n1871 gnd.n1870 9.3005
R19044 gnd.n5202 gnd.n5201 9.3005
R19045 gnd.n5203 gnd.n1869 9.3005
R19046 gnd.n5215 gnd.n5204 9.3005
R19047 gnd.n5214 gnd.n5205 9.3005
R19048 gnd.n5213 gnd.n5206 9.3005
R19049 gnd.n5211 gnd.n5207 9.3005
R19050 gnd.n4826 gnd.n4759 9.3005
R19051 gnd.n4819 gnd.n4818 9.3005
R19052 gnd.n4817 gnd.n4765 9.3005
R19053 gnd.n4816 gnd.n4815 9.3005
R19054 gnd.n4767 gnd.n4766 9.3005
R19055 gnd.n4809 gnd.n4808 9.3005
R19056 gnd.n4807 gnd.n4769 9.3005
R19057 gnd.n4806 gnd.n4805 9.3005
R19058 gnd.n4771 gnd.n4770 9.3005
R19059 gnd.n4799 gnd.n4798 9.3005
R19060 gnd.n4797 gnd.n4773 9.3005
R19061 gnd.n4796 gnd.n4795 9.3005
R19062 gnd.n4775 gnd.n4774 9.3005
R19063 gnd.n4789 gnd.n4788 9.3005
R19064 gnd.n4787 gnd.n4777 9.3005
R19065 gnd.n4786 gnd.n4785 9.3005
R19066 gnd.n4780 gnd.n4778 9.3005
R19067 gnd.n4779 gnd.n1986 9.3005
R19068 gnd.n4763 gnd.n4760 9.3005
R19069 gnd.n4825 gnd.n4824 9.3005
R19070 gnd.n5074 gnd.n1985 9.3005
R19071 gnd.n5076 gnd.n5075 9.3005
R19072 gnd.n1972 gnd.n1971 9.3005
R19073 gnd.n5089 gnd.n5088 9.3005
R19074 gnd.n5090 gnd.n1970 9.3005
R19075 gnd.n5092 gnd.n5091 9.3005
R19076 gnd.n1955 gnd.n1954 9.3005
R19077 gnd.n5105 gnd.n5104 9.3005
R19078 gnd.n5106 gnd.n1953 9.3005
R19079 gnd.n5108 gnd.n5107 9.3005
R19080 gnd.n1940 gnd.n1939 9.3005
R19081 gnd.n5121 gnd.n5120 9.3005
R19082 gnd.n5122 gnd.n1938 9.3005
R19083 gnd.n5124 gnd.n5123 9.3005
R19084 gnd.n1923 gnd.n1922 9.3005
R19085 gnd.n5137 gnd.n5136 9.3005
R19086 gnd.n5138 gnd.n1921 9.3005
R19087 gnd.n5148 gnd.n5139 9.3005
R19088 gnd.n5147 gnd.n5140 9.3005
R19089 gnd.n5146 gnd.n5141 9.3005
R19090 gnd.n5145 gnd.n5143 9.3005
R19091 gnd.n5142 gnd.n1887 9.3005
R19092 gnd.n5188 gnd.n1888 9.3005
R19093 gnd.n5187 gnd.n1889 9.3005
R19094 gnd.n5186 gnd.n1890 9.3005
R19095 gnd.n1896 gnd.n1891 9.3005
R19096 gnd.n1895 gnd.n1893 9.3005
R19097 gnd.n1892 gnd.n1778 9.3005
R19098 gnd.n5459 gnd.n1779 9.3005
R19099 gnd.n5458 gnd.n1780 9.3005
R19100 gnd.n5457 gnd.n1781 9.3005
R19101 gnd.n1861 gnd.n1782 9.3005
R19102 gnd.n5445 gnd.n1792 9.3005
R19103 gnd.n5444 gnd.n1793 9.3005
R19104 gnd.n5443 gnd.n1794 9.3005
R19105 gnd.n1756 gnd.n1755 9.3005
R19106 gnd.n5472 gnd.n5471 9.3005
R19107 gnd.n5473 gnd.n1754 9.3005
R19108 gnd.n5475 gnd.n5474 9.3005
R19109 gnd.n1740 gnd.n1739 9.3005
R19110 gnd.n5488 gnd.n5487 9.3005
R19111 gnd.n5489 gnd.n1738 9.3005
R19112 gnd.n5491 gnd.n5490 9.3005
R19113 gnd.n1722 gnd.n1721 9.3005
R19114 gnd.n5504 gnd.n5503 9.3005
R19115 gnd.n5505 gnd.n1720 9.3005
R19116 gnd.n5507 gnd.n5506 9.3005
R19117 gnd.n1706 gnd.n1705 9.3005
R19118 gnd.n5520 gnd.n5519 9.3005
R19119 gnd.n5521 gnd.n1704 9.3005
R19120 gnd.n5523 gnd.n5522 9.3005
R19121 gnd.n1688 gnd.n1687 9.3005
R19122 gnd.n5536 gnd.n5535 9.3005
R19123 gnd.n5537 gnd.n1686 9.3005
R19124 gnd.n5539 gnd.n5538 9.3005
R19125 gnd.n1672 gnd.n1671 9.3005
R19126 gnd.n5552 gnd.n5551 9.3005
R19127 gnd.n5553 gnd.n1670 9.3005
R19128 gnd.n5555 gnd.n5554 9.3005
R19129 gnd.n1653 gnd.n1652 9.3005
R19130 gnd.n5570 gnd.n5569 9.3005
R19131 gnd.n5571 gnd.n1651 9.3005
R19132 gnd.n5692 gnd.n5572 9.3005
R19133 gnd.n5691 gnd.n5690 9.3005
R19134 gnd.n5073 gnd.n5072 9.3005
R19135 gnd.n1608 gnd.n1386 9.3005
R19136 gnd.n5742 gnd.n1385 9.3005
R19137 gnd.n5743 gnd.n1384 9.3005
R19138 gnd.n5744 gnd.n1383 9.3005
R19139 gnd.n1382 gnd.n1379 9.3005
R19140 gnd.n5749 gnd.n1378 9.3005
R19141 gnd.n5750 gnd.n1377 9.3005
R19142 gnd.n5751 gnd.n1376 9.3005
R19143 gnd.n1375 gnd.n1372 9.3005
R19144 gnd.n5756 gnd.n1371 9.3005
R19145 gnd.n5757 gnd.n1370 9.3005
R19146 gnd.n5758 gnd.n1369 9.3005
R19147 gnd.n1368 gnd.n1365 9.3005
R19148 gnd.n1367 gnd.n1363 9.3005
R19149 gnd.n5765 gnd.n1362 9.3005
R19150 gnd.n5767 gnd.n5766 9.3005
R19151 gnd.n5734 gnd.n1611 9.3005
R19152 gnd.n5733 gnd.n1612 9.3005
R19153 gnd.n1616 gnd.n1613 9.3005
R19154 gnd.n5728 gnd.n1617 9.3005
R19155 gnd.n5727 gnd.n1618 9.3005
R19156 gnd.n5726 gnd.n1619 9.3005
R19157 gnd.n1623 gnd.n1620 9.3005
R19158 gnd.n5721 gnd.n1624 9.3005
R19159 gnd.n5720 gnd.n1625 9.3005
R19160 gnd.n5719 gnd.n1626 9.3005
R19161 gnd.n1630 gnd.n1627 9.3005
R19162 gnd.n5714 gnd.n1631 9.3005
R19163 gnd.n5713 gnd.n1632 9.3005
R19164 gnd.n5712 gnd.n1633 9.3005
R19165 gnd.n1637 gnd.n1634 9.3005
R19166 gnd.n5707 gnd.n1638 9.3005
R19167 gnd.n5706 gnd.n1639 9.3005
R19168 gnd.n5705 gnd.n1640 9.3005
R19169 gnd.n1645 gnd.n1643 9.3005
R19170 gnd.n5700 gnd.n5699 9.3005
R19171 gnd.n5735 gnd.n1610 9.3005
R19172 gnd.n4985 gnd.n4935 9.3005
R19173 gnd.n4984 gnd.n4937 9.3005
R19174 gnd.n4983 gnd.n4938 9.3005
R19175 gnd.n4981 gnd.n4939 9.3005
R19176 gnd.n4980 gnd.n4940 9.3005
R19177 gnd.n4978 gnd.n4941 9.3005
R19178 gnd.n4977 gnd.n4942 9.3005
R19179 gnd.n4975 gnd.n4943 9.3005
R19180 gnd.n4974 gnd.n4944 9.3005
R19181 gnd.n4972 gnd.n4945 9.3005
R19182 gnd.n4971 gnd.n4946 9.3005
R19183 gnd.n4969 gnd.n4947 9.3005
R19184 gnd.n4968 gnd.n4948 9.3005
R19185 gnd.n4966 gnd.n4949 9.3005
R19186 gnd.n4965 gnd.n4950 9.3005
R19187 gnd.n4963 gnd.n4951 9.3005
R19188 gnd.n4962 gnd.n4952 9.3005
R19189 gnd.n4960 gnd.n4953 9.3005
R19190 gnd.n4959 gnd.n4954 9.3005
R19191 gnd.n4957 gnd.n4956 9.3005
R19192 gnd.n4955 gnd.n1900 9.3005
R19193 gnd.n5175 gnd.n1899 9.3005
R19194 gnd.n5177 gnd.n5176 9.3005
R19195 gnd.n5178 gnd.n1898 9.3005
R19196 gnd.n5182 gnd.n5179 9.3005
R19197 gnd.n5181 gnd.n5180 9.3005
R19198 gnd.n1865 gnd.n1864 9.3005
R19199 gnd.n5220 gnd.n5219 9.3005
R19200 gnd.n5221 gnd.n1863 9.3005
R19201 gnd.n5224 gnd.n5222 9.3005
R19202 gnd.n5225 gnd.n1862 9.3005
R19203 gnd.n5228 gnd.n5227 9.3005
R19204 gnd.n5229 gnd.n1860 9.3005
R19205 gnd.n5231 gnd.n5230 9.3005
R19206 gnd.n1856 gnd.n1855 9.3005
R19207 gnd.n5244 gnd.n5243 9.3005
R19208 gnd.n5245 gnd.n1854 9.3005
R19209 gnd.n5247 gnd.n5246 9.3005
R19210 gnd.n5248 gnd.n1853 9.3005
R19211 gnd.n5252 gnd.n5251 9.3005
R19212 gnd.n5253 gnd.n1852 9.3005
R19213 gnd.n5278 gnd.n5254 9.3005
R19214 gnd.n5279 gnd.n1851 9.3005
R19215 gnd.n5283 gnd.n5282 9.3005
R19216 gnd.n5284 gnd.n1850 9.3005
R19217 gnd.n5293 gnd.n5285 9.3005
R19218 gnd.n5292 gnd.n5286 9.3005
R19219 gnd.n5291 gnd.n5288 9.3005
R19220 gnd.n5287 gnd.n1842 9.3005
R19221 gnd.n5318 gnd.n1843 9.3005
R19222 gnd.n5319 gnd.n1841 9.3005
R19223 gnd.n5323 gnd.n5322 9.3005
R19224 gnd.n5324 gnd.n1840 9.3005
R19225 gnd.n5332 gnd.n5325 9.3005
R19226 gnd.n5331 gnd.n5326 9.3005
R19227 gnd.n5330 gnd.n5327 9.3005
R19228 gnd.n1833 gnd.n1832 9.3005
R19229 gnd.n5376 gnd.n5375 9.3005
R19230 gnd.n5377 gnd.n1831 9.3005
R19231 gnd.n5382 gnd.n5378 9.3005
R19232 gnd.n5381 gnd.n5380 9.3005
R19233 gnd.n5379 gnd.n1647 9.3005
R19234 gnd.n5696 gnd.n1646 9.3005
R19235 gnd.n5698 gnd.n5697 9.3005
R19236 gnd.n4987 gnd.n4986 9.3005
R19237 gnd.n4995 gnd.n4994 9.3005
R19238 gnd.n4996 gnd.n4929 9.3005
R19239 gnd.n4997 gnd.n4928 9.3005
R19240 gnd.n4927 gnd.n4925 9.3005
R19241 gnd.n5003 gnd.n4924 9.3005
R19242 gnd.n5004 gnd.n4923 9.3005
R19243 gnd.n5005 gnd.n4922 9.3005
R19244 gnd.n4921 gnd.n4919 9.3005
R19245 gnd.n5011 gnd.n4918 9.3005
R19246 gnd.n5012 gnd.n4917 9.3005
R19247 gnd.n5013 gnd.n4916 9.3005
R19248 gnd.n4915 gnd.n4913 9.3005
R19249 gnd.n5019 gnd.n4912 9.3005
R19250 gnd.n5020 gnd.n4911 9.3005
R19251 gnd.n5021 gnd.n4910 9.3005
R19252 gnd.n4909 gnd.n4907 9.3005
R19253 gnd.n5027 gnd.n4906 9.3005
R19254 gnd.n5028 gnd.n4905 9.3005
R19255 gnd.n5029 gnd.n4904 9.3005
R19256 gnd.n4903 gnd.n4898 9.3005
R19257 gnd.n5035 gnd.n4897 9.3005
R19258 gnd.n5036 gnd.n4896 9.3005
R19259 gnd.n5037 gnd.n4895 9.3005
R19260 gnd.n4894 gnd.n4892 9.3005
R19261 gnd.n5043 gnd.n4891 9.3005
R19262 gnd.n5044 gnd.n4890 9.3005
R19263 gnd.n5045 gnd.n4889 9.3005
R19264 gnd.n4888 gnd.n4886 9.3005
R19265 gnd.n5051 gnd.n4885 9.3005
R19266 gnd.n5052 gnd.n4884 9.3005
R19267 gnd.n5053 gnd.n4883 9.3005
R19268 gnd.n4882 gnd.n4880 9.3005
R19269 gnd.n5058 gnd.n4879 9.3005
R19270 gnd.n5059 gnd.n4878 9.3005
R19271 gnd.n4877 gnd.n4875 9.3005
R19272 gnd.n5064 gnd.n4874 9.3005
R19273 gnd.n5066 gnd.n5065 9.3005
R19274 gnd.n4993 gnd.n4934 9.3005
R19275 gnd.n4992 gnd.n4991 9.3005
R19276 gnd.n1980 gnd.n1979 9.3005
R19277 gnd.n5081 gnd.n5080 9.3005
R19278 gnd.n5082 gnd.n1978 9.3005
R19279 gnd.n5084 gnd.n5083 9.3005
R19280 gnd.n1964 gnd.n1963 9.3005
R19281 gnd.n5097 gnd.n5096 9.3005
R19282 gnd.n5098 gnd.n1962 9.3005
R19283 gnd.n5100 gnd.n5099 9.3005
R19284 gnd.n1948 gnd.n1947 9.3005
R19285 gnd.n5113 gnd.n5112 9.3005
R19286 gnd.n5114 gnd.n1946 9.3005
R19287 gnd.n5116 gnd.n5115 9.3005
R19288 gnd.n1932 gnd.n1931 9.3005
R19289 gnd.n5129 gnd.n5128 9.3005
R19290 gnd.n5130 gnd.n1930 9.3005
R19291 gnd.n5132 gnd.n5131 9.3005
R19292 gnd.n1915 gnd.n1914 9.3005
R19293 gnd.n5153 gnd.n5152 9.3005
R19294 gnd.n5154 gnd.n1913 9.3005
R19295 gnd.n5158 gnd.n5155 9.3005
R19296 gnd.n5157 gnd.n5156 9.3005
R19297 gnd.n1879 gnd.n1878 9.3005
R19298 gnd.n5193 gnd.n5192 9.3005
R19299 gnd.n5194 gnd.n1877 9.3005
R19300 gnd.n5196 gnd.n5195 9.3005
R19301 gnd.n5197 gnd.n1764 9.3005
R19302 gnd.n1748 gnd.n1747 9.3005
R19303 gnd.n5480 gnd.n5479 9.3005
R19304 gnd.n5481 gnd.n1746 9.3005
R19305 gnd.n5483 gnd.n5482 9.3005
R19306 gnd.n1731 gnd.n1730 9.3005
R19307 gnd.n5496 gnd.n5495 9.3005
R19308 gnd.n5497 gnd.n1729 9.3005
R19309 gnd.n5499 gnd.n5498 9.3005
R19310 gnd.n1714 gnd.n1713 9.3005
R19311 gnd.n5512 gnd.n5511 9.3005
R19312 gnd.n5513 gnd.n1712 9.3005
R19313 gnd.n5515 gnd.n5514 9.3005
R19314 gnd.n1697 gnd.n1696 9.3005
R19315 gnd.n5528 gnd.n5527 9.3005
R19316 gnd.n5529 gnd.n1695 9.3005
R19317 gnd.n5531 gnd.n5530 9.3005
R19318 gnd.n1680 gnd.n1679 9.3005
R19319 gnd.n5544 gnd.n5543 9.3005
R19320 gnd.n5545 gnd.n1678 9.3005
R19321 gnd.n5547 gnd.n5546 9.3005
R19322 gnd.n1663 gnd.n1662 9.3005
R19323 gnd.n5560 gnd.n5559 9.3005
R19324 gnd.n5561 gnd.n1661 9.3005
R19325 gnd.n5565 gnd.n5562 9.3005
R19326 gnd.n5564 gnd.n5563 9.3005
R19327 gnd.n1361 gnd.n1360 9.3005
R19328 gnd.n5769 gnd.n5768 9.3005
R19329 gnd.n5068 gnd.n5067 9.3005
R19330 gnd.n5467 gnd.n5466 9.3005
R19331 gnd.n5435 gnd.n1801 9.3005
R19332 gnd.n5434 gnd.n1802 9.3005
R19333 gnd.n3349 gnd.n1800 9.3005
R19334 gnd.n3352 gnd.n3348 9.3005
R19335 gnd.n3347 gnd.n2065 9.3005
R19336 gnd.n3346 gnd.n3345 9.3005
R19337 gnd.n2067 gnd.n2066 9.3005
R19338 gnd.n3339 gnd.n3338 9.3005
R19339 gnd.n3337 gnd.n2071 9.3005
R19340 gnd.n3336 gnd.n3335 9.3005
R19341 gnd.n2073 gnd.n2072 9.3005
R19342 gnd.n3329 gnd.n3328 9.3005
R19343 gnd.n3327 gnd.n2077 9.3005
R19344 gnd.n3326 gnd.n3325 9.3005
R19345 gnd.n2079 gnd.n2078 9.3005
R19346 gnd.n3319 gnd.n3318 9.3005
R19347 gnd.n3317 gnd.n2083 9.3005
R19348 gnd.n3316 gnd.n3315 9.3005
R19349 gnd.n2085 gnd.n2084 9.3005
R19350 gnd.n3309 gnd.n3308 9.3005
R19351 gnd.n3307 gnd.n2089 9.3005
R19352 gnd.n3306 gnd.n3305 9.3005
R19353 gnd.n2091 gnd.n2090 9.3005
R19354 gnd.n3299 gnd.n3298 9.3005
R19355 gnd.n3297 gnd.n2095 9.3005
R19356 gnd.n3296 gnd.n3295 9.3005
R19357 gnd.n2097 gnd.n2096 9.3005
R19358 gnd.n3289 gnd.n3288 9.3005
R19359 gnd.n3287 gnd.n2101 9.3005
R19360 gnd.n3286 gnd.n3285 9.3005
R19361 gnd.n2103 gnd.n2102 9.3005
R19362 gnd.n3279 gnd.n3278 9.3005
R19363 gnd.n3277 gnd.n2107 9.3005
R19364 gnd.n3276 gnd.n3275 9.3005
R19365 gnd.n2109 gnd.n2108 9.3005
R19366 gnd.n3269 gnd.n3268 9.3005
R19367 gnd.n3267 gnd.n2113 9.3005
R19368 gnd.n3266 gnd.n3265 9.3005
R19369 gnd.n2115 gnd.n2114 9.3005
R19370 gnd.n3259 gnd.n3258 9.3005
R19371 gnd.n3257 gnd.n2119 9.3005
R19372 gnd.n3256 gnd.n3255 9.3005
R19373 gnd.n2121 gnd.n2120 9.3005
R19374 gnd.n3249 gnd.n3248 9.3005
R19375 gnd.n3247 gnd.n2125 9.3005
R19376 gnd.n3246 gnd.n3245 9.3005
R19377 gnd.n2127 gnd.n2126 9.3005
R19378 gnd.n3239 gnd.n3238 9.3005
R19379 gnd.n3237 gnd.n2131 9.3005
R19380 gnd.n3236 gnd.n3235 9.3005
R19381 gnd.n2133 gnd.n2132 9.3005
R19382 gnd.n3229 gnd.n3228 9.3005
R19383 gnd.n3227 gnd.n2137 9.3005
R19384 gnd.n3226 gnd.n3225 9.3005
R19385 gnd.n2139 gnd.n2138 9.3005
R19386 gnd.n3219 gnd.n3218 9.3005
R19387 gnd.n3217 gnd.n2143 9.3005
R19388 gnd.n3216 gnd.n3215 9.3005
R19389 gnd.n2145 gnd.n2144 9.3005
R19390 gnd.n3209 gnd.n3208 9.3005
R19391 gnd.n3207 gnd.n2149 9.3005
R19392 gnd.n3206 gnd.n3205 9.3005
R19393 gnd.n2151 gnd.n2150 9.3005
R19394 gnd.n3199 gnd.n3198 9.3005
R19395 gnd.n3197 gnd.n2155 9.3005
R19396 gnd.n3196 gnd.n3195 9.3005
R19397 gnd.n2157 gnd.n2156 9.3005
R19398 gnd.n3189 gnd.n3188 9.3005
R19399 gnd.n3187 gnd.n2161 9.3005
R19400 gnd.n3186 gnd.n3185 9.3005
R19401 gnd.n2163 gnd.n2162 9.3005
R19402 gnd.n3179 gnd.n3178 9.3005
R19403 gnd.n3177 gnd.n2167 9.3005
R19404 gnd.n3176 gnd.n3175 9.3005
R19405 gnd.n2169 gnd.n2168 9.3005
R19406 gnd.n3169 gnd.n3168 9.3005
R19407 gnd.n3167 gnd.n2173 9.3005
R19408 gnd.n3166 gnd.n3165 9.3005
R19409 gnd.n2175 gnd.n2174 9.3005
R19410 gnd.n3159 gnd.n3158 9.3005
R19411 gnd.n3157 gnd.n2179 9.3005
R19412 gnd.n3156 gnd.n3155 9.3005
R19413 gnd.n2181 gnd.n2180 9.3005
R19414 gnd.n3149 gnd.n3148 9.3005
R19415 gnd.n3147 gnd.n2185 9.3005
R19416 gnd.n3146 gnd.n3145 9.3005
R19417 gnd.n2187 gnd.n2186 9.3005
R19418 gnd.n3351 gnd.n3350 9.3005
R19419 gnd.n6618 gnd.n6616 9.3005
R19420 gnd.n6751 gnd.n6750 9.3005
R19421 gnd.n6749 gnd.n6748 9.3005
R19422 gnd.n6635 gnd.n6634 9.3005
R19423 gnd.n6743 gnd.n6742 9.3005
R19424 gnd.n6741 gnd.n6740 9.3005
R19425 gnd.n6643 gnd.n6642 9.3005
R19426 gnd.n6735 gnd.n6734 9.3005
R19427 gnd.n6733 gnd.n6732 9.3005
R19428 gnd.n6655 gnd.n6654 9.3005
R19429 gnd.n6727 gnd.n6726 9.3005
R19430 gnd.n6725 gnd.n6724 9.3005
R19431 gnd.n6663 gnd.n6662 9.3005
R19432 gnd.n6719 gnd.n6718 9.3005
R19433 gnd.n6717 gnd.n6716 9.3005
R19434 gnd.n6675 gnd.n6674 9.3005
R19435 gnd.n6708 gnd.n6707 9.3005
R19436 gnd.n6706 gnd.n6676 9.3005
R19437 gnd.n6757 gnd.n6756 9.3005
R19438 gnd.n6669 gnd.n6668 9.3005
R19439 gnd.n6721 gnd.n6720 9.3005
R19440 gnd.n6723 gnd.n6722 9.3005
R19441 gnd.n6659 gnd.n6658 9.3005
R19442 gnd.n6729 gnd.n6728 9.3005
R19443 gnd.n6731 gnd.n6730 9.3005
R19444 gnd.n6649 gnd.n6648 9.3005
R19445 gnd.n6737 gnd.n6736 9.3005
R19446 gnd.n6739 gnd.n6738 9.3005
R19447 gnd.n6639 gnd.n6638 9.3005
R19448 gnd.n6745 gnd.n6744 9.3005
R19449 gnd.n6747 gnd.n6746 9.3005
R19450 gnd.n6629 gnd.n6628 9.3005
R19451 gnd.n6753 gnd.n6752 9.3005
R19452 gnd.n6755 gnd.n6754 9.3005
R19453 gnd.n6623 gnd.n6617 9.3005
R19454 gnd.n6715 gnd.n6714 9.3005
R19455 gnd.n6710 gnd.n6709 9.3005
R19456 gnd.n6705 gnd.n6704 9.3005
R19457 gnd.n6703 gnd.n6681 9.3005
R19458 gnd.n6702 gnd.n6701 9.3005
R19459 gnd.n6700 gnd.n6682 9.3005
R19460 gnd.n6699 gnd.n6698 9.3005
R19461 gnd.n6697 gnd.n6687 9.3005
R19462 gnd.n6696 gnd.n6695 9.3005
R19463 gnd.n6694 gnd.n6688 9.3005
R19464 gnd.n634 gnd.n633 9.3005
R19465 gnd.n6814 gnd.n6813 9.3005
R19466 gnd.n5821 gnd.n1307 9.3005
R19467 gnd.n5823 gnd.n5822 9.3005
R19468 gnd.n1293 gnd.n1292 9.3005
R19469 gnd.n5838 gnd.n5837 9.3005
R19470 gnd.n5839 gnd.n1290 9.3005
R19471 gnd.n5842 gnd.n5841 9.3005
R19472 gnd.n5840 gnd.n1291 9.3005
R19473 gnd.n1252 gnd.n1251 9.3005
R19474 gnd.n5994 gnd.n5993 9.3005
R19475 gnd.n5995 gnd.n1250 9.3005
R19476 gnd.n5997 gnd.n5996 9.3005
R19477 gnd.n1237 gnd.n1236 9.3005
R19478 gnd.n6010 gnd.n6009 9.3005
R19479 gnd.n6011 gnd.n1235 9.3005
R19480 gnd.n6013 gnd.n6012 9.3005
R19481 gnd.n1222 gnd.n1221 9.3005
R19482 gnd.n6026 gnd.n6025 9.3005
R19483 gnd.n6027 gnd.n1220 9.3005
R19484 gnd.n6029 gnd.n6028 9.3005
R19485 gnd.n1205 gnd.n1204 9.3005
R19486 gnd.n6043 gnd.n6042 9.3005
R19487 gnd.n6044 gnd.n1202 9.3005
R19488 gnd.n6047 gnd.n6046 9.3005
R19489 gnd.n6045 gnd.n1203 9.3005
R19490 gnd.n1099 gnd.n1098 9.3005
R19491 gnd.n6136 gnd.n6135 9.3005
R19492 gnd.n6137 gnd.n1097 9.3005
R19493 gnd.n6139 gnd.n6138 9.3005
R19494 gnd.n1084 gnd.n1083 9.3005
R19495 gnd.n6152 gnd.n6151 9.3005
R19496 gnd.n6153 gnd.n1082 9.3005
R19497 gnd.n6155 gnd.n6154 9.3005
R19498 gnd.n1070 gnd.n1069 9.3005
R19499 gnd.n6168 gnd.n6167 9.3005
R19500 gnd.n6169 gnd.n1068 9.3005
R19501 gnd.n6171 gnd.n6170 9.3005
R19502 gnd.n1054 gnd.n1053 9.3005
R19503 gnd.n6186 gnd.n6185 9.3005
R19504 gnd.n6187 gnd.n1051 9.3005
R19505 gnd.n6190 gnd.n6189 9.3005
R19506 gnd.n6188 gnd.n1052 9.3005
R19507 gnd.n1012 gnd.n1011 9.3005
R19508 gnd.n6441 gnd.n6440 9.3005
R19509 gnd.n6442 gnd.n1010 9.3005
R19510 gnd.n6444 gnd.n6443 9.3005
R19511 gnd.n996 gnd.n995 9.3005
R19512 gnd.n6457 gnd.n6456 9.3005
R19513 gnd.n6458 gnd.n994 9.3005
R19514 gnd.n6460 gnd.n6459 9.3005
R19515 gnd.n981 gnd.n980 9.3005
R19516 gnd.n6473 gnd.n6472 9.3005
R19517 gnd.n6474 gnd.n979 9.3005
R19518 gnd.n6476 gnd.n6475 9.3005
R19519 gnd.n966 gnd.n965 9.3005
R19520 gnd.n6489 gnd.n6488 9.3005
R19521 gnd.n6490 gnd.n964 9.3005
R19522 gnd.n6492 gnd.n6491 9.3005
R19523 gnd.n951 gnd.n950 9.3005
R19524 gnd.n6505 gnd.n6504 9.3005
R19525 gnd.n6506 gnd.n949 9.3005
R19526 gnd.n6508 gnd.n6507 9.3005
R19527 gnd.n935 gnd.n934 9.3005
R19528 gnd.n6520 gnd.n6519 9.3005
R19529 gnd.n6521 gnd.n932 9.3005
R19530 gnd.n6530 gnd.n6529 9.3005
R19531 gnd.n6528 gnd.n933 9.3005
R19532 gnd.n6527 gnd.n6526 9.3005
R19533 gnd.n6525 gnd.n6522 9.3005
R19534 gnd.n895 gnd.n893 9.3005
R19535 gnd.n6588 gnd.n6587 9.3005
R19536 gnd.n6586 gnd.n894 9.3005
R19537 gnd.n6585 gnd.n6584 9.3005
R19538 gnd.n6583 gnd.n896 9.3005
R19539 gnd.n6582 gnd.n6581 9.3005
R19540 gnd.n6580 gnd.n6579 9.3005
R19541 gnd.n652 gnd.n651 9.3005
R19542 gnd.n6792 gnd.n6791 9.3005
R19543 gnd.n6793 gnd.n650 9.3005
R19544 gnd.n6796 gnd.n6795 9.3005
R19545 gnd.n6794 gnd.n636 9.3005
R19546 gnd.n6810 gnd.n635 9.3005
R19547 gnd.n6812 gnd.n6811 9.3005
R19548 gnd.n5820 gnd.n5819 9.3005
R19549 gnd.n5806 gnd.n5805 9.3005
R19550 gnd.n5804 gnd.n1333 9.3005
R19551 gnd.n5803 gnd.n5802 9.3005
R19552 gnd.n5799 gnd.n1335 9.3005
R19553 gnd.n5796 gnd.n5795 9.3005
R19554 gnd.n5794 gnd.n1338 9.3005
R19555 gnd.n5793 gnd.n5792 9.3005
R19556 gnd.n5789 gnd.n1339 9.3005
R19557 gnd.n5786 gnd.n5785 9.3005
R19558 gnd.n1334 gnd.n1308 9.3005
R19559 gnd.n1859 gnd.n1858 9.3005
R19560 gnd.n5236 gnd.n5235 9.3005
R19561 gnd.n5237 gnd.n1857 9.3005
R19562 gnd.n5239 gnd.n5238 9.3005
R19563 gnd.n1809 gnd.n1807 9.3005
R19564 gnd.n5427 gnd.n5426 9.3005
R19565 gnd.n5425 gnd.n1808 9.3005
R19566 gnd.n5424 gnd.n5423 9.3005
R19567 gnd.n5422 gnd.n1810 9.3005
R19568 gnd.n5421 gnd.n5420 9.3005
R19569 gnd.n5419 gnd.n1813 9.3005
R19570 gnd.n5418 gnd.n5417 9.3005
R19571 gnd.n5416 gnd.n1814 9.3005
R19572 gnd.n5415 gnd.n5414 9.3005
R19573 gnd.n5413 gnd.n1817 9.3005
R19574 gnd.n5412 gnd.n5411 9.3005
R19575 gnd.n5410 gnd.n1818 9.3005
R19576 gnd.n5409 gnd.n5408 9.3005
R19577 gnd.n5407 gnd.n1821 9.3005
R19578 gnd.n5406 gnd.n5405 9.3005
R19579 gnd.n5404 gnd.n1822 9.3005
R19580 gnd.n5403 gnd.n5402 9.3005
R19581 gnd.n5401 gnd.n1825 9.3005
R19582 gnd.n5400 gnd.n5399 9.3005
R19583 gnd.n5398 gnd.n1826 9.3005
R19584 gnd.n5397 gnd.n5396 9.3005
R19585 gnd.n5395 gnd.n1829 9.3005
R19586 gnd.n5394 gnd.n5393 9.3005
R19587 gnd.n5392 gnd.n1830 9.3005
R19588 gnd.n5391 gnd.n5390 9.3005
R19589 gnd.n5389 gnd.n5388 9.3005
R19590 gnd.n1353 gnd.n1341 9.3005
R19591 gnd.n5783 gnd.n1340 9.3005
R19592 gnd.n5782 gnd.n5781 9.3005
R19593 gnd.n5778 gnd.n5777 9.3005
R19594 gnd.n1346 gnd.n1343 9.3005
R19595 gnd.n5636 gnd.n5635 9.3005
R19596 gnd.n5638 gnd.n5637 9.3005
R19597 gnd.n5621 gnd.n5620 9.3005
R19598 gnd.n5644 gnd.n5643 9.3005
R19599 gnd.n5646 gnd.n5645 9.3005
R19600 gnd.n5609 gnd.n5608 9.3005
R19601 gnd.n5652 gnd.n5651 9.3005
R19602 gnd.n5654 gnd.n5653 9.3005
R19603 gnd.n5598 gnd.n5597 9.3005
R19604 gnd.n5660 gnd.n5659 9.3005
R19605 gnd.n5662 gnd.n5661 9.3005
R19606 gnd.n5586 gnd.n5585 9.3005
R19607 gnd.n5668 gnd.n5667 9.3005
R19608 gnd.n5670 gnd.n5669 9.3005
R19609 gnd.n5582 gnd.n5574 9.3005
R19610 gnd.n5674 gnd.n5673 9.3005
R19611 gnd.n5672 gnd.n5671 9.3005
R19612 gnd.n5580 gnd.n5579 9.3005
R19613 gnd.n5666 gnd.n5665 9.3005
R19614 gnd.n5664 gnd.n5663 9.3005
R19615 gnd.n5592 gnd.n5591 9.3005
R19616 gnd.n5658 gnd.n5657 9.3005
R19617 gnd.n5656 gnd.n5655 9.3005
R19618 gnd.n5605 gnd.n5604 9.3005
R19619 gnd.n5650 gnd.n5649 9.3005
R19620 gnd.n5648 gnd.n5647 9.3005
R19621 gnd.n5615 gnd.n5614 9.3005
R19622 gnd.n5642 gnd.n5641 9.3005
R19623 gnd.n5640 gnd.n5639 9.3005
R19624 gnd.n5631 gnd.n5630 9.3005
R19625 gnd.n5634 gnd.n1347 9.3005
R19626 gnd.n5776 gnd.n5775 9.3005
R19627 gnd.n5774 gnd.n1342 9.3005
R19628 gnd.n5685 gnd.n5675 9.3005
R19629 gnd.n5684 gnd.n5683 9.3005
R19630 gnd.n5682 gnd.n5679 9.3005
R19631 gnd.n5681 gnd.n5680 9.3005
R19632 gnd.n1285 gnd.n1284 9.3005
R19633 gnd.n5847 gnd.n5846 9.3005
R19634 gnd.n5848 gnd.n1281 9.3005
R19635 gnd.n5850 gnd.n5849 9.3005
R19636 gnd.n5851 gnd.n1280 9.3005
R19637 gnd.n5856 gnd.n5855 9.3005
R19638 gnd.n5857 gnd.n1278 9.3005
R19639 gnd.n5965 gnd.n5964 9.3005
R19640 gnd.n5963 gnd.n1279 9.3005
R19641 gnd.n5962 gnd.n5961 9.3005
R19642 gnd.n5960 gnd.n5858 9.3005
R19643 gnd.n5959 gnd.n5958 9.3005
R19644 gnd.n5957 gnd.n5861 9.3005
R19645 gnd.n5956 gnd.n5955 9.3005
R19646 gnd.n5954 gnd.n5862 9.3005
R19647 gnd.n5953 gnd.n5952 9.3005
R19648 gnd.n5951 gnd.n5950 9.3005
R19649 gnd.n1197 gnd.n1196 9.3005
R19650 gnd.n6052 gnd.n6051 9.3005
R19651 gnd.n6053 gnd.n1193 9.3005
R19652 gnd.n6055 gnd.n6054 9.3005
R19653 gnd.n6056 gnd.n1192 9.3005
R19654 gnd.n6059 gnd.n6058 9.3005
R19655 gnd.n6060 gnd.n1191 9.3005
R19656 gnd.n6062 gnd.n6061 9.3005
R19657 gnd.n6063 gnd.n1190 9.3005
R19658 gnd.n6066 gnd.n6065 9.3005
R19659 gnd.n6067 gnd.n1189 9.3005
R19660 gnd.n6069 gnd.n6068 9.3005
R19661 gnd.n6070 gnd.n1188 9.3005
R19662 gnd.n6073 gnd.n6072 9.3005
R19663 gnd.n6074 gnd.n1186 9.3005
R19664 gnd.n6077 gnd.n6076 9.3005
R19665 gnd.n6075 gnd.n1187 9.3005
R19666 gnd.n1047 gnd.n1046 9.3005
R19667 gnd.n6195 gnd.n6194 9.3005
R19668 gnd.n6196 gnd.n1043 9.3005
R19669 gnd.n6198 gnd.n6197 9.3005
R19670 gnd.n6199 gnd.n1042 9.3005
R19671 gnd.n6202 gnd.n6201 9.3005
R19672 gnd.n6203 gnd.n1040 9.3005
R19673 gnd.n6412 gnd.n6411 9.3005
R19674 gnd.n6410 gnd.n1041 9.3005
R19675 gnd.n6409 gnd.n6408 9.3005
R19676 gnd.n6407 gnd.n6204 9.3005
R19677 gnd.n6406 gnd.n6405 9.3005
R19678 gnd.n6404 gnd.n6207 9.3005
R19679 gnd.n6403 gnd.n6402 9.3005
R19680 gnd.n6401 gnd.n6208 9.3005
R19681 gnd.n6400 gnd.n6399 9.3005
R19682 gnd.n6398 gnd.n6211 9.3005
R19683 gnd.n6397 gnd.n6396 9.3005
R19684 gnd.n6395 gnd.n6212 9.3005
R19685 gnd.n6394 gnd.n6393 9.3005
R19686 gnd.n6392 gnd.n6215 9.3005
R19687 gnd.n6391 gnd.n6390 9.3005
R19688 gnd.n6389 gnd.n6216 9.3005
R19689 gnd.n6388 gnd.n6387 9.3005
R19690 gnd.n6386 gnd.n6219 9.3005
R19691 gnd.n6385 gnd.n6384 9.3005
R19692 gnd.n6383 gnd.n6220 9.3005
R19693 gnd.n917 gnd.n916 9.3005
R19694 gnd.n6545 gnd.n6544 9.3005
R19695 gnd.n6546 gnd.n914 9.3005
R19696 gnd.n6549 gnd.n6548 9.3005
R19697 gnd.n6547 gnd.n915 9.3005
R19698 gnd.n876 gnd.n875 9.3005
R19699 gnd.n6603 gnd.n6602 9.3005
R19700 gnd.n6604 gnd.n873 9.3005
R19701 gnd.n6606 gnd.n6605 9.3005
R19702 gnd.n6607 gnd.n872 9.3005
R19703 gnd.n6610 gnd.n6609 9.3005
R19704 gnd.n6611 gnd.n870 9.3005
R19705 gnd.n6766 gnd.n6765 9.3005
R19706 gnd.n6764 gnd.n871 9.3005
R19707 gnd.n6763 gnd.n6762 9.3005
R19708 gnd.n6761 gnd.n6612 9.3005
R19709 gnd.n6760 gnd.n6615 9.3005
R19710 gnd.n5687 gnd.n5686 9.3005
R19711 gnd.n7058 gnd.n7057 9.3005
R19712 gnd.n7059 gnd.n476 9.3005
R19713 gnd.n7061 gnd.n7060 9.3005
R19714 gnd.n460 gnd.n459 9.3005
R19715 gnd.n7074 gnd.n7073 9.3005
R19716 gnd.n7075 gnd.n458 9.3005
R19717 gnd.n7077 gnd.n7076 9.3005
R19718 gnd.n444 gnd.n443 9.3005
R19719 gnd.n7090 gnd.n7089 9.3005
R19720 gnd.n7091 gnd.n442 9.3005
R19721 gnd.n7093 gnd.n7092 9.3005
R19722 gnd.n426 gnd.n425 9.3005
R19723 gnd.n7106 gnd.n7105 9.3005
R19724 gnd.n7107 gnd.n424 9.3005
R19725 gnd.n7109 gnd.n7108 9.3005
R19726 gnd.n410 gnd.n409 9.3005
R19727 gnd.n7122 gnd.n7121 9.3005
R19728 gnd.n7123 gnd.n407 9.3005
R19729 gnd.n7128 gnd.n7127 9.3005
R19730 gnd.n7126 gnd.n408 9.3005
R19731 gnd.n7125 gnd.n7124 9.3005
R19732 gnd.n377 gnd.n375 9.3005
R19733 gnd.n7179 gnd.n7178 9.3005
R19734 gnd.n7177 gnd.n376 9.3005
R19735 gnd.n7176 gnd.n7175 9.3005
R19736 gnd.n7174 gnd.n378 9.3005
R19737 gnd.n7173 gnd.n7172 9.3005
R19738 gnd.n316 gnd.n314 9.3005
R19739 gnd.n7318 gnd.n7317 9.3005
R19740 gnd.n7316 gnd.n315 9.3005
R19741 gnd.n7315 gnd.n7314 9.3005
R19742 gnd.n7313 gnd.n317 9.3005
R19743 gnd.n7312 gnd.n7311 9.3005
R19744 gnd.n7310 gnd.n321 9.3005
R19745 gnd.n7309 gnd.n7308 9.3005
R19746 gnd.n7307 gnd.n322 9.3005
R19747 gnd.n293 gnd.n292 9.3005
R19748 gnd.n7332 gnd.n7331 9.3005
R19749 gnd.n7333 gnd.n291 9.3005
R19750 gnd.n7335 gnd.n7334 9.3005
R19751 gnd.n277 gnd.n276 9.3005
R19752 gnd.n7348 gnd.n7347 9.3005
R19753 gnd.n7349 gnd.n275 9.3005
R19754 gnd.n7351 gnd.n7350 9.3005
R19755 gnd.n263 gnd.n262 9.3005
R19756 gnd.n7364 gnd.n7363 9.3005
R19757 gnd.n7365 gnd.n261 9.3005
R19758 gnd.n7367 gnd.n7366 9.3005
R19759 gnd.n247 gnd.n246 9.3005
R19760 gnd.n7380 gnd.n7379 9.3005
R19761 gnd.n7381 gnd.n245 9.3005
R19762 gnd.n7383 gnd.n7382 9.3005
R19763 gnd.n232 gnd.n231 9.3005
R19764 gnd.n7396 gnd.n7395 9.3005
R19765 gnd.n7397 gnd.n230 9.3005
R19766 gnd.n7399 gnd.n7398 9.3005
R19767 gnd.n217 gnd.n216 9.3005
R19768 gnd.n7412 gnd.n7411 9.3005
R19769 gnd.n7413 gnd.n214 9.3005
R19770 gnd.n7483 gnd.n7482 9.3005
R19771 gnd.n7481 gnd.n215 9.3005
R19772 gnd.n7480 gnd.n7479 9.3005
R19773 gnd.n7478 gnd.n7414 9.3005
R19774 gnd.n7477 gnd.n7476 9.3005
R19775 gnd.n478 gnd.n477 9.3005
R19776 gnd.n7473 gnd.n7416 9.3005
R19777 gnd.n7472 gnd.n7471 9.3005
R19778 gnd.n7470 gnd.n7421 9.3005
R19779 gnd.n7469 gnd.n7468 9.3005
R19780 gnd.n7467 gnd.n7422 9.3005
R19781 gnd.n7466 gnd.n7465 9.3005
R19782 gnd.n7464 gnd.n7429 9.3005
R19783 gnd.n7463 gnd.n7462 9.3005
R19784 gnd.n7461 gnd.n7430 9.3005
R19785 gnd.n7460 gnd.n7459 9.3005
R19786 gnd.n7458 gnd.n7437 9.3005
R19787 gnd.n7457 gnd.n7456 9.3005
R19788 gnd.n7455 gnd.n7438 9.3005
R19789 gnd.n7454 gnd.n7453 9.3005
R19790 gnd.n7452 gnd.n7445 9.3005
R19791 gnd.n7451 gnd.n7450 9.3005
R19792 gnd.n120 gnd.n117 9.3005
R19793 gnd.n7577 gnd.n7576 9.3005
R19794 gnd.n7475 gnd.n7474 9.3005
R19795 gnd.n6970 gnd.n565 9.3005
R19796 gnd.n6969 gnd.n6968 9.3005
R19797 gnd.n6967 gnd.n567 9.3005
R19798 gnd.n6966 gnd.n6965 9.3005
R19799 gnd.n6964 gnd.n570 9.3005
R19800 gnd.n6963 gnd.n6962 9.3005
R19801 gnd.n6961 gnd.n571 9.3005
R19802 gnd.n6960 gnd.n6959 9.3005
R19803 gnd.n6958 gnd.n574 9.3005
R19804 gnd.n6957 gnd.n6956 9.3005
R19805 gnd.n6955 gnd.n575 9.3005
R19806 gnd.n6954 gnd.n6953 9.3005
R19807 gnd.n6952 gnd.n578 9.3005
R19808 gnd.n6951 gnd.n6950 9.3005
R19809 gnd.n6949 gnd.n579 9.3005
R19810 gnd.n6948 gnd.n6947 9.3005
R19811 gnd.n6946 gnd.n582 9.3005
R19812 gnd.n6945 gnd.n6944 9.3005
R19813 gnd.n6943 gnd.n583 9.3005
R19814 gnd.n6942 gnd.n6941 9.3005
R19815 gnd.n6940 gnd.n384 9.3005
R19816 gnd.n7161 gnd.n383 9.3005
R19817 gnd.n7163 gnd.n7162 9.3005
R19818 gnd.n7164 gnd.n381 9.3005
R19819 gnd.n7167 gnd.n7166 9.3005
R19820 gnd.n7165 gnd.n382 9.3005
R19821 gnd.n354 gnd.n352 9.3005
R19822 gnd.n7209 gnd.n7208 9.3005
R19823 gnd.n7207 gnd.n353 9.3005
R19824 gnd.n7206 gnd.n7205 9.3005
R19825 gnd.n7204 gnd.n75 9.3005
R19826 gnd.n7626 gnd.n76 9.3005
R19827 gnd.n7625 gnd.n7624 9.3005
R19828 gnd.n7623 gnd.n77 9.3005
R19829 gnd.n7622 gnd.n7621 9.3005
R19830 gnd.n7620 gnd.n81 9.3005
R19831 gnd.n7619 gnd.n7618 9.3005
R19832 gnd.n7617 gnd.n82 9.3005
R19833 gnd.n7616 gnd.n7615 9.3005
R19834 gnd.n7614 gnd.n86 9.3005
R19835 gnd.n7613 gnd.n7612 9.3005
R19836 gnd.n7611 gnd.n87 9.3005
R19837 gnd.n7610 gnd.n7609 9.3005
R19838 gnd.n7608 gnd.n91 9.3005
R19839 gnd.n7607 gnd.n7606 9.3005
R19840 gnd.n7605 gnd.n92 9.3005
R19841 gnd.n7604 gnd.n7603 9.3005
R19842 gnd.n7602 gnd.n96 9.3005
R19843 gnd.n7601 gnd.n7600 9.3005
R19844 gnd.n7599 gnd.n97 9.3005
R19845 gnd.n7598 gnd.n7597 9.3005
R19846 gnd.n7596 gnd.n101 9.3005
R19847 gnd.n7595 gnd.n7594 9.3005
R19848 gnd.n7593 gnd.n102 9.3005
R19849 gnd.n7592 gnd.n7591 9.3005
R19850 gnd.n7590 gnd.n106 9.3005
R19851 gnd.n7589 gnd.n7588 9.3005
R19852 gnd.n7587 gnd.n107 9.3005
R19853 gnd.n7586 gnd.n7585 9.3005
R19854 gnd.n7584 gnd.n111 9.3005
R19855 gnd.n7583 gnd.n7582 9.3005
R19856 gnd.n7581 gnd.n112 9.3005
R19857 gnd.n7580 gnd.n7579 9.3005
R19858 gnd.n7578 gnd.n116 9.3005
R19859 gnd.n6972 gnd.n6971 9.3005
R19860 gnd.t150 gnd.n4267 9.24152
R19861 gnd.n4647 gnd.t37 9.24152
R19862 gnd.n3373 gnd.t65 9.24152
R19863 gnd.t231 gnd.n1925 9.24152
R19864 gnd.n5517 gnd.t192 9.24152
R19865 gnd.n7111 gnd.t202 9.24152
R19866 gnd.n259 gnd.t196 9.24152
R19867 gnd.t352 gnd.t150 8.92286
R19868 gnd.n5835 gnd.n1297 8.92286
R19869 gnd.n6040 gnd.n1209 8.92286
R19870 gnd.n6117 gnd.n1119 8.92286
R19871 gnd.n6183 gnd.n1058 8.92286
R19872 gnd.n6422 gnd.n1033 8.92286
R19873 gnd.n6486 gnd.n970 8.92286
R19874 gnd.n6510 gnd.n945 8.92286
R19875 gnd.n6600 gnd.n880 8.92286
R19876 gnd.n6769 gnd.n6768 8.92286
R19877 gnd.n4626 gnd.n4601 8.92171
R19878 gnd.n4594 gnd.n4569 8.92171
R19879 gnd.n4562 gnd.n4537 8.92171
R19880 gnd.n4531 gnd.n4506 8.92171
R19881 gnd.n4499 gnd.n4474 8.92171
R19882 gnd.n4467 gnd.n4442 8.92171
R19883 gnd.n4435 gnd.n4410 8.92171
R19884 gnd.n4404 gnd.n4379 8.92171
R19885 gnd.n727 gnd.n709 8.72777
R19886 gnd.n3613 gnd.t141 8.60421
R19887 gnd.t262 gnd.n1957 8.60421
R19888 gnd.n5549 gnd.t194 8.60421
R19889 gnd.n5825 gnd.n1305 8.60421
R19890 gnd.n1179 gnd.t163 8.60421
R19891 gnd.t184 gnd.n1016 8.60421
R19892 gnd.n7079 gnd.t286 8.60421
R19893 gnd.n228 gnd.t288 8.60421
R19894 gnd.n3655 gnd.n3635 8.43467
R19895 gnd.n54 gnd.n34 8.43467
R19896 gnd.n5209 gnd.n0 8.41456
R19897 gnd.n7627 gnd.n7626 8.41456
R19898 gnd.n5677 gnd.t99 8.28555
R19899 gnd.n4627 gnd.n4599 8.14595
R19900 gnd.n4595 gnd.n4567 8.14595
R19901 gnd.n4563 gnd.n4535 8.14595
R19902 gnd.n4532 gnd.n4504 8.14595
R19903 gnd.n4500 gnd.n4472 8.14595
R19904 gnd.n4468 gnd.n4440 8.14595
R19905 gnd.n4436 gnd.n4408 8.14595
R19906 gnd.n4405 gnd.n4377 8.14595
R19907 gnd.n4632 gnd.n4631 7.97301
R19908 gnd.t143 gnd.n4167 7.9669
R19909 gnd.n5889 gnd.t190 7.9669
R19910 gnd.n6372 gnd.t177 7.9669
R19911 gnd.n7576 gnd.n120 7.75808
R19912 gnd.n6714 gnd.n6710 7.75808
R19913 gnd.n5775 gnd.n5774 7.75808
R19914 gnd.n4824 gnd.n4763 7.75808
R19915 gnd.n4664 gnd.n3355 7.64824
R19916 gnd.n1282 gnd.t114 7.64824
R19917 gnd.n5968 gnd.n5967 7.64824
R19918 gnd.t7 gnd.n1218 7.64824
R19919 gnd.n6093 gnd.t133 7.64824
R19920 gnd.n6165 gnd.t133 7.64824
R19921 gnd.n6288 gnd.t165 7.64824
R19922 gnd.t165 gnd.n990 7.64824
R19923 gnd.t4 gnd.n937 7.64824
R19924 gnd.n6590 gnd.n890 7.64824
R19925 gnd.n6568 gnd.t105 7.64824
R19926 gnd.n4100 gnd.t147 7.32958
R19927 gnd.t175 gnd.t52 7.32958
R19928 gnd.n1432 gnd.n1431 7.30353
R19929 gnd.n726 gnd.n725 7.30353
R19930 gnd.n4060 gnd.n3779 7.01093
R19931 gnd.n3782 gnd.n3780 7.01093
R19932 gnd.n4070 gnd.n4069 7.01093
R19933 gnd.n4081 gnd.n3763 7.01093
R19934 gnd.n4080 gnd.n3766 7.01093
R19935 gnd.n4091 gnd.n3754 7.01093
R19936 gnd.n3757 gnd.n3755 7.01093
R19937 gnd.n4101 gnd.n4100 7.01093
R19938 gnd.n4111 gnd.n3735 7.01093
R19939 gnd.n4110 gnd.n3738 7.01093
R19940 gnd.n4127 gnd.n3728 7.01093
R19941 gnd.n4137 gnd.n3719 7.01093
R19942 gnd.n4148 gnd.n4147 7.01093
R19943 gnd.n4168 gnd.n3704 7.01093
R19944 gnd.n4167 gnd.n3683 7.01093
R19945 gnd.n4185 gnd.n3684 7.01093
R19946 gnd.n4179 gnd.n4178 7.01093
R19947 gnd.n4195 gnd.n3531 7.01093
R19948 gnd.n4205 gnd.n3523 7.01093
R19949 gnd.n4216 gnd.n3514 7.01093
R19950 gnd.n3613 gnd.n3612 7.01093
R19951 gnd.n4226 gnd.n4225 7.01093
R19952 gnd.n4237 gnd.n3497 7.01093
R19953 gnd.n4236 gnd.n3500 7.01093
R19954 gnd.n4247 gnd.n3489 7.01093
R19955 gnd.n4257 gnd.n4256 7.01093
R19956 gnd.n4268 gnd.n3471 7.01093
R19957 gnd.n4267 gnd.n3474 7.01093
R19958 gnd.n4278 gnd.n3462 7.01093
R19959 gnd.n3465 gnd.n3463 7.01093
R19960 gnd.n4288 gnd.n4287 7.01093
R19961 gnd.n4299 gnd.n3446 7.01093
R19962 gnd.n3440 gnd.n3438 7.01093
R19963 gnd.n4319 gnd.n4318 7.01093
R19964 gnd.n4330 gnd.n3421 7.01093
R19965 gnd.n4329 gnd.n3424 7.01093
R19966 gnd.n4340 gnd.n3412 7.01093
R19967 gnd.n3415 gnd.n3413 7.01093
R19968 gnd.n4361 gnd.n3395 7.01093
R19969 gnd.n4360 gnd.n3398 7.01093
R19970 gnd.n4371 gnd.n3387 7.01093
R19971 gnd.n3388 gnd.n3380 7.01093
R19972 gnd.n4637 gnd.n4636 7.01093
R19973 gnd.n4647 gnd.n3370 7.01093
R19974 gnd.n4646 gnd.n3373 7.01093
R19975 gnd.n4657 gnd.n3364 7.01093
R19976 gnd.n4664 gnd.n1988 7.01093
R19977 gnd.n6173 gnd.t8 7.01093
R19978 gnd.t186 gnd.n6414 7.01093
R19979 gnd.n6768 gnd.t72 7.01093
R19980 gnd.n3738 gnd.t139 6.69227
R19981 gnd.n4268 gnd.t352 6.69227
R19982 gnd.n4350 gnd.t138 6.69227
R19983 gnd.n5372 gnd.t194 6.69227
R19984 gnd.n5948 gnd.t123 6.69227
R19985 gnd.n6237 gnd.t170 6.69227
R19986 gnd.n6866 gnd.t286 6.69227
R19987 gnd.n807 gnd.n806 6.5566
R19988 gnd.n1598 gnd.n1597 6.5566
R19989 gnd.n1458 gnd.n1452 6.5566
R19990 gnd.n787 gnd.n694 6.5566
R19991 gnd.n5911 gnd.n5901 6.37362
R19992 gnd.n6023 gnd.n1225 6.37362
R19993 gnd.n6102 gnd.n1134 6.37362
R19994 gnd.n6470 gnd.n984 6.37362
R19995 gnd.n6532 gnd.n928 6.37362
R19996 gnd.n6523 gnd.n911 6.37362
R19997 gnd.n6775 gnd.t12 6.37362
R19998 gnd.n5802 gnd.n5800 6.20656
R19999 gnd.n7538 gnd.n7535 6.20656
R20000 gnd.n5029 gnd.n4902 6.20656
R20001 gnd.n6695 gnd.n6691 6.20656
R20002 gnd.t9 gnd.n4159 6.05496
R20003 gnd.n4160 gnd.t149 6.05496
R20004 gnd.n4225 gnd.t134 6.05496
R20005 gnd.n3587 gnd.t145 6.05496
R20006 gnd.n5315 gnd.t192 6.05496
R20007 gnd.n6905 gnd.t202 6.05496
R20008 gnd.n4629 gnd.n4599 5.81868
R20009 gnd.n4597 gnd.n4567 5.81868
R20010 gnd.n4565 gnd.n4535 5.81868
R20011 gnd.n4534 gnd.n4504 5.81868
R20012 gnd.n4502 gnd.n4472 5.81868
R20013 gnd.n4470 gnd.n4440 5.81868
R20014 gnd.n4438 gnd.n4408 5.81868
R20015 gnd.n4407 gnd.n4377 5.81868
R20016 gnd.n5975 gnd.t15 5.73631
R20017 gnd.t0 gnd.n1209 5.73631
R20018 gnd.t183 gnd.n1078 5.73631
R20019 gnd.n6298 gnd.t181 5.73631
R20020 gnd.t127 gnd.n945 5.73631
R20021 gnd.t72 gnd.n646 5.73631
R20022 gnd.n802 gnd.n534 5.62001
R20023 gnd.n1605 gnd.n1390 5.62001
R20024 gnd.n1605 gnd.n1391 5.62001
R20025 gnd.n794 gnd.n534 5.62001
R20026 gnd.n3919 gnd.n3914 5.4308
R20027 gnd.n4672 gnd.n2055 5.4308
R20028 gnd.n4237 gnd.t144 5.41765
R20029 gnd.t151 gnd.n3482 5.41765
R20030 gnd.n4309 gnd.t128 5.41765
R20031 gnd.n5430 gnd.t251 5.41765
R20032 gnd.n5275 gnd.t210 5.41765
R20033 gnd.n1194 gnd.t161 5.41765
R20034 gnd.n6494 gnd.t167 5.41765
R20035 gnd.n7158 gnd.t225 5.41765
R20036 gnd.t291 gnd.n359 5.41765
R20037 gnd.n6015 gnd.n1233 5.09899
R20038 gnd.n5889 gnd.n5888 5.09899
R20039 gnd.t119 gnd.n6109 5.09899
R20040 gnd.n6157 gnd.n1080 5.09899
R20041 gnd.n6095 gnd.n6094 5.09899
R20042 gnd.n6462 gnd.n992 5.09899
R20043 gnd.n6267 gnd.n6266 5.09899
R20044 gnd.n6478 gnd.t174 5.09899
R20045 gnd.n6373 gnd.n6372 5.09899
R20046 gnd.n6542 gnd.n919 5.09899
R20047 gnd.n4627 gnd.n4626 5.04292
R20048 gnd.n4595 gnd.n4594 5.04292
R20049 gnd.n4563 gnd.n4562 5.04292
R20050 gnd.n4532 gnd.n4531 5.04292
R20051 gnd.n4500 gnd.n4499 5.04292
R20052 gnd.n4468 gnd.n4467 5.04292
R20053 gnd.n4436 gnd.n4435 5.04292
R20054 gnd.n4405 gnd.n4404 5.04292
R20055 gnd.n3675 gnd.n3674 4.82753
R20056 gnd.n74 gnd.n73 4.82753
R20057 gnd.n4206 gnd.t136 4.78034
R20058 gnd.n3465 gnd.t142 4.78034
R20059 gnd.n5296 gnd.t237 4.78034
R20060 gnd.t161 gnd.n1111 4.78034
R20061 gnd.n6247 gnd.t167 4.78034
R20062 gnd.t41 gnd.n648 4.78034
R20063 gnd.n6916 gnd.t271 4.78034
R20064 gnd.n3680 gnd.n3677 4.74817
R20065 gnd.n4192 gnd.n3533 4.74817
R20066 gnd.n4190 gnd.n3534 4.74817
R20067 gnd.n3616 gnd.n3610 4.74817
R20068 gnd.n3696 gnd.n3677 4.74817
R20069 gnd.n3695 gnd.n3533 4.74817
R20070 gnd.n4191 gnd.n4190 4.74817
R20071 gnd.n3616 gnd.n3615 4.74817
R20072 gnd.n7324 gnd.n7323 4.74817
R20073 gnd.n337 gnd.n304 4.74817
R20074 gnd.n7225 gnd.n303 4.74817
R20075 gnd.n327 gnd.n302 4.74817
R20076 gnd.n7303 gnd.n301 4.74817
R20077 gnd.n7324 gnd.n305 4.74817
R20078 gnd.n7322 gnd.n304 4.74817
R20079 gnd.n338 gnd.n303 4.74817
R20080 gnd.n7226 gnd.n302 4.74817
R20081 gnd.n328 gnd.n301 4.74817
R20082 gnd.n5465 gnd.n5464 4.74817
R20083 gnd.n5452 gnd.n1769 4.74817
R20084 gnd.n5450 gnd.n1768 4.74817
R20085 gnd.n5438 gnd.n1767 4.74817
R20086 gnd.n1766 gnd.n1763 4.74817
R20087 gnd.n5465 gnd.n1770 4.74817
R20088 gnd.n5463 gnd.n1769 4.74817
R20089 gnd.n5453 gnd.n1768 4.74817
R20090 gnd.n5449 gnd.n1767 4.74817
R20091 gnd.n5439 gnd.n1766 4.74817
R20092 gnd.n3655 gnd.n3654 4.7074
R20093 gnd.n54 gnd.n53 4.7074
R20094 gnd.n3675 gnd.n3655 4.65959
R20095 gnd.n74 gnd.n54 4.65959
R20096 gnd.n7018 gnd.n536 4.6132
R20097 gnd.n1609 gnd.n1606 4.6132
R20098 gnd.n5358 gnd.n1364 4.46168
R20099 gnd.n5968 gnd.t120 4.46168
R20100 gnd.t169 gnd.n890 4.46168
R20101 gnd.n7046 gnd.n518 4.46168
R20102 gnd.n722 gnd.n709 4.46111
R20103 gnd.n4612 gnd.n4608 4.38594
R20104 gnd.n4580 gnd.n4576 4.38594
R20105 gnd.n4548 gnd.n4544 4.38594
R20106 gnd.n4517 gnd.n4513 4.38594
R20107 gnd.n4485 gnd.n4481 4.38594
R20108 gnd.n4453 gnd.n4449 4.38594
R20109 gnd.n4421 gnd.n4417 4.38594
R20110 gnd.n4390 gnd.n4386 4.38594
R20111 gnd.n4623 gnd.n4601 4.26717
R20112 gnd.n4591 gnd.n4569 4.26717
R20113 gnd.n4559 gnd.n4537 4.26717
R20114 gnd.n4528 gnd.n4506 4.26717
R20115 gnd.n4496 gnd.n4474 4.26717
R20116 gnd.n4464 gnd.n4442 4.26717
R20117 gnd.n4432 gnd.n4410 4.26717
R20118 gnd.n4401 gnd.n4379 4.26717
R20119 gnd.t137 gnd.n3711 4.14303
R20120 gnd.n3424 gnd.t140 4.14303
R20121 gnd.n5335 gnd.t220 4.14303
R20122 gnd.n1149 gnd.t5 4.14303
R20123 gnd.n6289 gnd.t125 4.14303
R20124 gnd.n6885 gnd.t235 4.14303
R20125 gnd.n4631 gnd.n4630 4.08274
R20126 gnd.n806 gnd.n691 4.05904
R20127 gnd.n1597 gnd.n1596 4.05904
R20128 gnd.n1462 gnd.n1452 4.05904
R20129 gnd.n788 gnd.n787 4.05904
R20130 gnd.n15 gnd.n7 3.99943
R20131 gnd.t114 gnd.n1254 3.82437
R20132 gnd.n6007 gnd.n1241 3.82437
R20133 gnd.n5927 gnd.n5883 3.82437
R20134 gnd.n6149 gnd.n1087 3.82437
R20135 gnd.n6087 gnd.n1150 3.82437
R20136 gnd.n6454 gnd.n1000 3.82437
R20137 gnd.n6307 gnd.n6306 3.82437
R20138 gnd.n6381 gnd.n6380 3.82437
R20139 gnd.n6552 gnd.n6551 3.82437
R20140 gnd.n6613 gnd.t41 3.82437
R20141 gnd.n4631 gnd.n4503 3.70378
R20142 gnd.n4189 gnd.n3676 3.65935
R20143 gnd.n15 gnd.n14 3.60163
R20144 gnd.n5078 gnd.t25 3.50571
R20145 gnd.n5386 gnd.t44 3.50571
R20146 gnd.n6846 gnd.t33 3.50571
R20147 gnd.n7493 gnd.t29 3.50571
R20148 gnd.n4622 gnd.n4603 3.49141
R20149 gnd.n4590 gnd.n4571 3.49141
R20150 gnd.n4558 gnd.n4539 3.49141
R20151 gnd.n4527 gnd.n4508 3.49141
R20152 gnd.n4495 gnd.n4476 3.49141
R20153 gnd.n4463 gnd.n4444 3.49141
R20154 gnd.n4431 gnd.n4412 3.49141
R20155 gnd.n4400 gnd.n4381 3.49141
R20156 gnd.n5853 gnd.t15 3.18706
R20157 gnd.n6781 gnd.t85 3.18706
R20158 gnd.n3718 gnd.t137 2.8684
R20159 gnd.n3656 gnd.t331 2.82907
R20160 gnd.n3656 gnd.t277 2.82907
R20161 gnd.n3658 gnd.t316 2.82907
R20162 gnd.n3658 gnd.t193 2.82907
R20163 gnd.n3660 gnd.t224 2.82907
R20164 gnd.n3660 gnd.t201 2.82907
R20165 gnd.n3662 gnd.t199 2.82907
R20166 gnd.n3662 gnd.t344 2.82907
R20167 gnd.n3664 gnd.t207 2.82907
R20168 gnd.n3664 gnd.t268 2.82907
R20169 gnd.n3666 gnd.t303 2.82907
R20170 gnd.n3666 gnd.t248 2.82907
R20171 gnd.n3668 gnd.t283 2.82907
R20172 gnd.n3668 gnd.t205 2.82907
R20173 gnd.n3670 gnd.t254 2.82907
R20174 gnd.n3670 gnd.t336 2.82907
R20175 gnd.n3672 gnd.t311 2.82907
R20176 gnd.n3672 gnd.t310 2.82907
R20177 gnd.n3617 gnd.t217 2.82907
R20178 gnd.n3617 gnd.t250 2.82907
R20179 gnd.n3619 gnd.t267 2.82907
R20180 gnd.n3619 gnd.t332 2.82907
R20181 gnd.n3621 gnd.t242 2.82907
R20182 gnd.n3621 gnd.t234 2.82907
R20183 gnd.n3623 gnd.t290 2.82907
R20184 gnd.n3623 gnd.t278 2.82907
R20185 gnd.n3625 gnd.t337 2.82907
R20186 gnd.n3625 gnd.t257 2.82907
R20187 gnd.n3627 gnd.t273 2.82907
R20188 gnd.n3627 gnd.t304 2.82907
R20189 gnd.n3629 gnd.t320 2.82907
R20190 gnd.n3629 gnd.t241 2.82907
R20191 gnd.n3631 gnd.t249 2.82907
R20192 gnd.n3631 gnd.t285 2.82907
R20193 gnd.n3633 gnd.t209 2.82907
R20194 gnd.n3633 gnd.t228 2.82907
R20195 gnd.n3636 gnd.t343 2.82907
R20196 gnd.n3636 gnd.t221 2.82907
R20197 gnd.n3638 gnd.t238 2.82907
R20198 gnd.n3638 gnd.t307 2.82907
R20199 gnd.n3640 gnd.t211 2.82907
R20200 gnd.n3640 gnd.t350 2.82907
R20201 gnd.n3642 gnd.t260 2.82907
R20202 gnd.n3642 gnd.t252 2.82907
R20203 gnd.n3644 gnd.t321 2.82907
R20204 gnd.n3644 gnd.t230 2.82907
R20205 gnd.n3646 gnd.t246 2.82907
R20206 gnd.n3646 gnd.t275 2.82907
R20207 gnd.n3648 gnd.t293 2.82907
R20208 gnd.n3648 gnd.t212 2.82907
R20209 gnd.n3650 gnd.t232 2.82907
R20210 gnd.n3650 gnd.t266 2.82907
R20211 gnd.n3652 gnd.t340 2.82907
R20212 gnd.n3652 gnd.t348 2.82907
R20213 gnd.n71 gnd.t215 2.82907
R20214 gnd.n71 gnd.t233 2.82907
R20215 gnd.n69 gnd.t297 2.82907
R20216 gnd.n69 gnd.t197 2.82907
R20217 gnd.n67 gnd.t330 2.82907
R20218 gnd.n67 gnd.t240 2.82907
R20219 gnd.n65 gnd.t351 2.82907
R20220 gnd.n65 gnd.t259 2.82907
R20221 gnd.n63 gnd.t219 2.82907
R20222 gnd.n63 gnd.t342 2.82907
R20223 gnd.n61 gnd.t312 2.82907
R20224 gnd.n61 gnd.t326 2.82907
R20225 gnd.n59 gnd.t328 2.82907
R20226 gnd.n59 gnd.t349 2.82907
R20227 gnd.n57 gnd.t322 2.82907
R20228 gnd.n57 gnd.t272 2.82907
R20229 gnd.n55 gnd.t236 2.82907
R20230 gnd.n55 gnd.t309 2.82907
R20231 gnd.n32 gnd.t214 2.82907
R20232 gnd.n32 gnd.t223 2.82907
R20233 gnd.n30 gnd.t327 2.82907
R20234 gnd.n30 gnd.t295 2.82907
R20235 gnd.n28 gnd.t280 2.82907
R20236 gnd.n28 gnd.t345 2.82907
R20237 gnd.n26 gnd.t335 2.82907
R20238 gnd.n26 gnd.t313 2.82907
R20239 gnd.n24 gnd.t294 2.82907
R20240 gnd.n24 gnd.t324 2.82907
R20241 gnd.n22 gnd.t319 2.82907
R20242 gnd.n22 gnd.t329 2.82907
R20243 gnd.n20 gnd.t270 2.82907
R20244 gnd.n20 gnd.t226 2.82907
R20245 gnd.n18 gnd.t203 2.82907
R20246 gnd.n18 gnd.t301 2.82907
R20247 gnd.n16 gnd.t284 2.82907
R20248 gnd.n16 gnd.t338 2.82907
R20249 gnd.n51 gnd.t341 2.82907
R20250 gnd.n51 gnd.t347 2.82907
R20251 gnd.n49 gnd.t300 2.82907
R20252 gnd.n49 gnd.t269 2.82907
R20253 gnd.n47 gnd.t256 2.82907
R20254 gnd.n47 gnd.t323 2.82907
R20255 gnd.n45 gnd.t315 2.82907
R20256 gnd.n45 gnd.t281 2.82907
R20257 gnd.n43 gnd.t261 2.82907
R20258 gnd.n43 gnd.t306 2.82907
R20259 gnd.n41 gnd.t292 2.82907
R20260 gnd.n41 gnd.t299 2.82907
R20261 gnd.n39 gnd.t244 2.82907
R20262 gnd.n39 gnd.t346 2.82907
R20263 gnd.n37 gnd.t339 2.82907
R20264 gnd.n37 gnd.t274 2.82907
R20265 gnd.n35 gnd.t264 2.82907
R20266 gnd.n35 gnd.t333 2.82907
R20267 gnd.n4619 gnd.n4618 2.71565
R20268 gnd.n4587 gnd.n4586 2.71565
R20269 gnd.n4555 gnd.n4554 2.71565
R20270 gnd.n4524 gnd.n4523 2.71565
R20271 gnd.n4492 gnd.n4491 2.71565
R20272 gnd.n4460 gnd.n4459 2.71565
R20273 gnd.n4428 gnd.n4427 2.71565
R20274 gnd.n4397 gnd.n4396 2.71565
R20275 gnd.n5999 gnd.n1248 2.54975
R20276 gnd.n5901 gnd.t187 2.54975
R20277 gnd.n5948 gnd.n5947 2.54975
R20278 gnd.n6125 gnd.t156 2.54975
R20279 gnd.n6141 gnd.n1095 2.54975
R20280 gnd.n6110 gnd.t119 2.54975
R20281 gnd.n6080 gnd.n6079 2.54975
R20282 gnd.n6446 gnd.n1008 2.54975
R20283 gnd.n6256 gnd.t174 2.54975
R20284 gnd.n6316 gnd.n6257 2.54975
R20285 gnd.n6335 gnd.t130 2.54975
R20286 gnd.n6352 gnd.n6237 2.54975
R20287 gnd.n6523 gnd.t172 2.54975
R20288 gnd.n6560 gnd.n906 2.54975
R20289 gnd.n4189 gnd.n3677 2.27742
R20290 gnd.n4189 gnd.n3533 2.27742
R20291 gnd.n4190 gnd.n4189 2.27742
R20292 gnd.n4189 gnd.n3616 2.27742
R20293 gnd.n7325 gnd.n7324 2.27742
R20294 gnd.n7325 gnd.n304 2.27742
R20295 gnd.n7325 gnd.n303 2.27742
R20296 gnd.n7325 gnd.n302 2.27742
R20297 gnd.n7325 gnd.n301 2.27742
R20298 gnd.n5466 gnd.n5465 2.27742
R20299 gnd.n5466 gnd.n1769 2.27742
R20300 gnd.n5466 gnd.n1768 2.27742
R20301 gnd.n5466 gnd.n1767 2.27742
R20302 gnd.n5466 gnd.n1766 2.27742
R20303 gnd.n4069 gnd.t21 2.23109
R20304 gnd.n4194 gnd.t136 2.23109
R20305 gnd.n6165 gnd.t5 2.23109
R20306 gnd.t125 gnd.n6288 2.23109
R20307 gnd.n236 gnd.t222 2.23109
R20308 gnd.n4615 gnd.n4605 1.93989
R20309 gnd.n4583 gnd.n4573 1.93989
R20310 gnd.n4551 gnd.n4541 1.93989
R20311 gnd.n4520 gnd.n4510 1.93989
R20312 gnd.n4488 gnd.n4478 1.93989
R20313 gnd.n4456 gnd.n4446 1.93989
R20314 gnd.n4424 gnd.n4414 1.93989
R20315 gnd.n4393 gnd.n4383 1.93989
R20316 gnd.t157 gnd.n4080 1.59378
R20317 gnd.n3490 gnd.t151 1.59378
R20318 gnd.n3588 gnd.t128 1.59378
R20319 gnd.n5118 gnd.t227 1.59378
R20320 gnd.n5320 gnd.t216 1.59378
R20321 gnd.n6890 gnd.t308 1.59378
R20322 gnd.n7385 gnd.t213 1.59378
R20323 gnd.n1530 gnd.t18 1.27512
R20324 gnd.n1530 gnd.n1411 1.27512
R20325 gnd.n5991 gnd.n1256 1.27512
R20326 gnd.n5940 gnd.n5939 1.27512
R20327 gnd.n6133 gnd.n1103 1.27512
R20328 gnd.n1179 gnd.n1163 1.27512
R20329 gnd.n6438 gnd.n1016 1.27512
R20330 gnd.n6326 gnd.n6325 1.27512
R20331 gnd.n6344 gnd.n6242 1.27512
R20332 gnd.n6569 gnd.n6568 1.27512
R20333 gnd.n6789 gnd.n655 1.27512
R20334 gnd.n3922 gnd.n3914 1.16414
R20335 gnd.n4675 gnd.n2055 1.16414
R20336 gnd.n4614 gnd.n4607 1.16414
R20337 gnd.n4582 gnd.n4575 1.16414
R20338 gnd.n4550 gnd.n4543 1.16414
R20339 gnd.n4519 gnd.n4512 1.16414
R20340 gnd.n4487 gnd.n4480 1.16414
R20341 gnd.n4455 gnd.n4448 1.16414
R20342 gnd.n4423 gnd.n4416 1.16414
R20343 gnd.n4392 gnd.n4385 1.16414
R20344 gnd.n7018 gnd.n7017 0.970197
R20345 gnd.n5735 gnd.n1606 0.970197
R20346 gnd.n4598 gnd.n4566 0.962709
R20347 gnd.n4630 gnd.n4598 0.962709
R20348 gnd.n4471 gnd.n4439 0.962709
R20349 gnd.n4503 gnd.n4471 0.962709
R20350 gnd.n4160 gnd.t9 0.956468
R20351 gnd.n4298 gnd.t145 0.956468
R20352 gnd.n5160 gnd.t282 0.956468
R20353 gnd.n5280 gnd.t200 0.956468
R20354 gnd.n1288 gnd.t175 0.956468
R20355 gnd.n5999 gnd.t152 0.956468
R20356 gnd.n906 gnd.t2 0.956468
R20357 gnd.n670 gnd.t154 0.956468
R20358 gnd.n6938 gnd.t243 0.956468
R20359 gnd.n7353 gnd.t239 0.956468
R20360 gnd.n3667 gnd.n3665 0.773756
R20361 gnd.n66 gnd.n64 0.773756
R20362 gnd.n3674 gnd.n3673 0.773756
R20363 gnd.n3673 gnd.n3671 0.773756
R20364 gnd.n3671 gnd.n3669 0.773756
R20365 gnd.n3669 gnd.n3667 0.773756
R20366 gnd.n3665 gnd.n3663 0.773756
R20367 gnd.n3663 gnd.n3661 0.773756
R20368 gnd.n3661 gnd.n3659 0.773756
R20369 gnd.n3659 gnd.n3657 0.773756
R20370 gnd.n58 gnd.n56 0.773756
R20371 gnd.n60 gnd.n58 0.773756
R20372 gnd.n62 gnd.n60 0.773756
R20373 gnd.n64 gnd.n62 0.773756
R20374 gnd.n68 gnd.n66 0.773756
R20375 gnd.n70 gnd.n68 0.773756
R20376 gnd.n72 gnd.n70 0.773756
R20377 gnd.n73 gnd.n72 0.773756
R20378 gnd.n2 gnd.n1 0.672012
R20379 gnd.n3 gnd.n2 0.672012
R20380 gnd.n4 gnd.n3 0.672012
R20381 gnd.n5 gnd.n4 0.672012
R20382 gnd.n6 gnd.n5 0.672012
R20383 gnd.n7 gnd.n6 0.672012
R20384 gnd.n9 gnd.n8 0.672012
R20385 gnd.n10 gnd.n9 0.672012
R20386 gnd.n11 gnd.n10 0.672012
R20387 gnd.n12 gnd.n11 0.672012
R20388 gnd.n13 gnd.n12 0.672012
R20389 gnd.n14 gnd.n13 0.672012
R20390 gnd.n5983 gnd.t58 0.637812
R20391 gnd.n5920 gnd.t166 0.637812
R20392 gnd.n6081 gnd.t8 0.637812
R20393 gnd.n6415 gnd.t186 0.637812
R20394 gnd.n6374 gnd.t179 0.637812
R20395 gnd.n6781 gnd.t48 0.637812
R20396 gnd.n7628 gnd.n7627 0.63688
R20397 gnd gnd.n0 0.634843
R20398 gnd.n3635 gnd.n3634 0.573776
R20399 gnd.n3634 gnd.n3632 0.573776
R20400 gnd.n3632 gnd.n3630 0.573776
R20401 gnd.n3630 gnd.n3628 0.573776
R20402 gnd.n3628 gnd.n3626 0.573776
R20403 gnd.n3626 gnd.n3624 0.573776
R20404 gnd.n3624 gnd.n3622 0.573776
R20405 gnd.n3622 gnd.n3620 0.573776
R20406 gnd.n3620 gnd.n3618 0.573776
R20407 gnd.n3654 gnd.n3653 0.573776
R20408 gnd.n3653 gnd.n3651 0.573776
R20409 gnd.n3651 gnd.n3649 0.573776
R20410 gnd.n3649 gnd.n3647 0.573776
R20411 gnd.n3647 gnd.n3645 0.573776
R20412 gnd.n3645 gnd.n3643 0.573776
R20413 gnd.n3643 gnd.n3641 0.573776
R20414 gnd.n3641 gnd.n3639 0.573776
R20415 gnd.n3639 gnd.n3637 0.573776
R20416 gnd.n19 gnd.n17 0.573776
R20417 gnd.n21 gnd.n19 0.573776
R20418 gnd.n23 gnd.n21 0.573776
R20419 gnd.n25 gnd.n23 0.573776
R20420 gnd.n27 gnd.n25 0.573776
R20421 gnd.n29 gnd.n27 0.573776
R20422 gnd.n31 gnd.n29 0.573776
R20423 gnd.n33 gnd.n31 0.573776
R20424 gnd.n34 gnd.n33 0.573776
R20425 gnd.n38 gnd.n36 0.573776
R20426 gnd.n40 gnd.n38 0.573776
R20427 gnd.n42 gnd.n40 0.573776
R20428 gnd.n44 gnd.n42 0.573776
R20429 gnd.n46 gnd.n44 0.573776
R20430 gnd.n48 gnd.n46 0.573776
R20431 gnd.n50 gnd.n48 0.573776
R20432 gnd.n52 gnd.n50 0.573776
R20433 gnd.n53 gnd.n52 0.573776
R20434 gnd.n7325 gnd.n300 0.5435
R20435 gnd.n5466 gnd.n1765 0.5435
R20436 gnd.n5688 gnd.n5687 0.523366
R20437 gnd.n6619 gnd.n6615 0.523366
R20438 gnd.n6813 gnd.n6812 0.489829
R20439 gnd.n5820 gnd.n1308 0.489829
R20440 gnd.n3562 gnd.n2059 0.486781
R20441 gnd.n3971 gnd.n3970 0.48678
R20442 gnd.n4653 gnd.n2013 0.480683
R20443 gnd.n4055 gnd.n4054 0.480683
R20444 gnd.n4826 gnd.n4825 0.477634
R20445 gnd.n5073 gnd.n1986 0.477634
R20446 gnd.n7476 gnd.n7475 0.477634
R20447 gnd.n7578 gnd.n7577 0.477634
R20448 gnd.n7570 gnd.n7569 0.465439
R20449 gnd.n7499 gnd.n7498 0.465439
R20450 gnd.n6978 gnd.n562 0.465439
R20451 gnd.n7051 gnd.n7050 0.465439
R20452 gnd.n5768 gnd.n5767 0.465439
R20453 gnd.n5699 gnd.n5698 0.465439
R20454 gnd.n4992 gnd.n4987 0.465439
R20455 gnd.n5067 gnd.n5066 0.465439
R20456 gnd.n3138 gnd.n2186 0.459342
R20457 gnd.n2501 gnd.n2495 0.459342
R20458 gnd.n7218 gnd.n7217 0.459342
R20459 gnd.n3350 gnd.n3349 0.459342
R20460 gnd.n5800 gnd.n5799 0.388379
R20461 gnd.n4611 gnd.n4610 0.388379
R20462 gnd.n4579 gnd.n4578 0.388379
R20463 gnd.n4547 gnd.n4546 0.388379
R20464 gnd.n4516 gnd.n4515 0.388379
R20465 gnd.n4484 gnd.n4483 0.388379
R20466 gnd.n4452 gnd.n4451 0.388379
R20467 gnd.n4420 gnd.n4419 0.388379
R20468 gnd.n4389 gnd.n4388 0.388379
R20469 gnd.n7539 gnd.n7538 0.388379
R20470 gnd.n4902 gnd.n4898 0.388379
R20471 gnd.n6691 gnd.n6687 0.388379
R20472 gnd.n5690 gnd.n5689 0.377553
R20473 gnd.n6620 gnd.n477 0.377553
R20474 gnd.n7628 gnd.n15 0.374463
R20475 gnd.t138 gnd.n4349 0.319156
R20476 gnd.n5217 gnd.t247 0.319156
R20477 gnd.n5241 gnd.t198 0.319156
R20478 gnd.n6108 gnd.t354 0.319156
R20479 gnd.t163 gnd.t180 0.319156
R20480 gnd.t173 gnd.t184 0.319156
R20481 gnd.t121 gnd.n976 0.319156
R20482 gnd.n7211 gnd.t298 0.319156
R20483 gnd.n7305 gnd.t314 0.319156
R20484 gnd.n3889 gnd.n3867 0.311721
R20485 gnd gnd.n7628 0.295112
R20486 gnd.n4720 gnd.n4719 0.268793
R20487 gnd.n5784 gnd.n1341 0.247451
R20488 gnd.n6971 gnd.n566 0.247451
R20489 gnd.n4719 gnd.n4718 0.241354
R20490 gnd.n536 gnd.n533 0.229039
R20491 gnd.n539 gnd.n536 0.229039
R20492 gnd.n1609 gnd.n1608 0.229039
R20493 gnd.n1610 gnd.n1609 0.229039
R20494 gnd.n3676 gnd.n0 0.210825
R20495 gnd.n4043 gnd.n3842 0.206293
R20496 gnd.n4628 gnd.n4600 0.155672
R20497 gnd.n4621 gnd.n4600 0.155672
R20498 gnd.n4621 gnd.n4620 0.155672
R20499 gnd.n4620 gnd.n4604 0.155672
R20500 gnd.n4613 gnd.n4604 0.155672
R20501 gnd.n4613 gnd.n4612 0.155672
R20502 gnd.n4596 gnd.n4568 0.155672
R20503 gnd.n4589 gnd.n4568 0.155672
R20504 gnd.n4589 gnd.n4588 0.155672
R20505 gnd.n4588 gnd.n4572 0.155672
R20506 gnd.n4581 gnd.n4572 0.155672
R20507 gnd.n4581 gnd.n4580 0.155672
R20508 gnd.n4564 gnd.n4536 0.155672
R20509 gnd.n4557 gnd.n4536 0.155672
R20510 gnd.n4557 gnd.n4556 0.155672
R20511 gnd.n4556 gnd.n4540 0.155672
R20512 gnd.n4549 gnd.n4540 0.155672
R20513 gnd.n4549 gnd.n4548 0.155672
R20514 gnd.n4533 gnd.n4505 0.155672
R20515 gnd.n4526 gnd.n4505 0.155672
R20516 gnd.n4526 gnd.n4525 0.155672
R20517 gnd.n4525 gnd.n4509 0.155672
R20518 gnd.n4518 gnd.n4509 0.155672
R20519 gnd.n4518 gnd.n4517 0.155672
R20520 gnd.n4501 gnd.n4473 0.155672
R20521 gnd.n4494 gnd.n4473 0.155672
R20522 gnd.n4494 gnd.n4493 0.155672
R20523 gnd.n4493 gnd.n4477 0.155672
R20524 gnd.n4486 gnd.n4477 0.155672
R20525 gnd.n4486 gnd.n4485 0.155672
R20526 gnd.n4469 gnd.n4441 0.155672
R20527 gnd.n4462 gnd.n4441 0.155672
R20528 gnd.n4462 gnd.n4461 0.155672
R20529 gnd.n4461 gnd.n4445 0.155672
R20530 gnd.n4454 gnd.n4445 0.155672
R20531 gnd.n4454 gnd.n4453 0.155672
R20532 gnd.n4437 gnd.n4409 0.155672
R20533 gnd.n4430 gnd.n4409 0.155672
R20534 gnd.n4430 gnd.n4429 0.155672
R20535 gnd.n4429 gnd.n4413 0.155672
R20536 gnd.n4422 gnd.n4413 0.155672
R20537 gnd.n4422 gnd.n4421 0.155672
R20538 gnd.n4406 gnd.n4378 0.155672
R20539 gnd.n4399 gnd.n4378 0.155672
R20540 gnd.n4399 gnd.n4398 0.155672
R20541 gnd.n4398 gnd.n4382 0.155672
R20542 gnd.n4391 gnd.n4382 0.155672
R20543 gnd.n4391 gnd.n4390 0.155672
R20544 gnd.n4751 gnd.n2013 0.152939
R20545 gnd.n4751 gnd.n4750 0.152939
R20546 gnd.n4750 gnd.n4749 0.152939
R20547 gnd.n4749 gnd.n2015 0.152939
R20548 gnd.n2016 gnd.n2015 0.152939
R20549 gnd.n2017 gnd.n2016 0.152939
R20550 gnd.n2018 gnd.n2017 0.152939
R20551 gnd.n2019 gnd.n2018 0.152939
R20552 gnd.n2020 gnd.n2019 0.152939
R20553 gnd.n2021 gnd.n2020 0.152939
R20554 gnd.n2022 gnd.n2021 0.152939
R20555 gnd.n2023 gnd.n2022 0.152939
R20556 gnd.n2024 gnd.n2023 0.152939
R20557 gnd.n2025 gnd.n2024 0.152939
R20558 gnd.n4721 gnd.n2025 0.152939
R20559 gnd.n4721 gnd.n4720 0.152939
R20560 gnd.n4056 gnd.n4055 0.152939
R20561 gnd.n4056 gnd.n3760 0.152939
R20562 gnd.n4084 gnd.n3760 0.152939
R20563 gnd.n4085 gnd.n4084 0.152939
R20564 gnd.n4086 gnd.n4085 0.152939
R20565 gnd.n4087 gnd.n4086 0.152939
R20566 gnd.n4087 gnd.n3732 0.152939
R20567 gnd.n4114 gnd.n3732 0.152939
R20568 gnd.n4115 gnd.n4114 0.152939
R20569 gnd.n4116 gnd.n4115 0.152939
R20570 gnd.n4117 gnd.n4116 0.152939
R20571 gnd.n4118 gnd.n4117 0.152939
R20572 gnd.n4120 gnd.n4118 0.152939
R20573 gnd.n4120 gnd.n4119 0.152939
R20574 gnd.n4119 gnd.n3700 0.152939
R20575 gnd.n4173 gnd.n3700 0.152939
R20576 gnd.n4174 gnd.n4173 0.152939
R20577 gnd.n4175 gnd.n4174 0.152939
R20578 gnd.n4175 gnd.n3518 0.152939
R20579 gnd.n4209 gnd.n3518 0.152939
R20580 gnd.n4210 gnd.n4209 0.152939
R20581 gnd.n4211 gnd.n4210 0.152939
R20582 gnd.n4212 gnd.n4211 0.152939
R20583 gnd.n4212 gnd.n3494 0.152939
R20584 gnd.n4240 gnd.n3494 0.152939
R20585 gnd.n4241 gnd.n4240 0.152939
R20586 gnd.n4242 gnd.n4241 0.152939
R20587 gnd.n4243 gnd.n4242 0.152939
R20588 gnd.n4243 gnd.n3468 0.152939
R20589 gnd.n4271 gnd.n3468 0.152939
R20590 gnd.n4272 gnd.n4271 0.152939
R20591 gnd.n4273 gnd.n4272 0.152939
R20592 gnd.n4274 gnd.n4273 0.152939
R20593 gnd.n4274 gnd.n3443 0.152939
R20594 gnd.n4302 gnd.n3443 0.152939
R20595 gnd.n4303 gnd.n4302 0.152939
R20596 gnd.n4304 gnd.n4303 0.152939
R20597 gnd.n4305 gnd.n4304 0.152939
R20598 gnd.n4305 gnd.n3418 0.152939
R20599 gnd.n4333 gnd.n3418 0.152939
R20600 gnd.n4334 gnd.n4333 0.152939
R20601 gnd.n4335 gnd.n4334 0.152939
R20602 gnd.n4336 gnd.n4335 0.152939
R20603 gnd.n4336 gnd.n3392 0.152939
R20604 gnd.n4364 gnd.n3392 0.152939
R20605 gnd.n4365 gnd.n4364 0.152939
R20606 gnd.n4366 gnd.n4365 0.152939
R20607 gnd.n4367 gnd.n4366 0.152939
R20608 gnd.n4367 gnd.n3367 0.152939
R20609 gnd.n4650 gnd.n3367 0.152939
R20610 gnd.n4651 gnd.n4650 0.152939
R20611 gnd.n4652 gnd.n4651 0.152939
R20612 gnd.n4653 gnd.n4652 0.152939
R20613 gnd.n4054 gnd.n3784 0.152939
R20614 gnd.n3805 gnd.n3784 0.152939
R20615 gnd.n3806 gnd.n3805 0.152939
R20616 gnd.n3812 gnd.n3806 0.152939
R20617 gnd.n3813 gnd.n3812 0.152939
R20618 gnd.n3814 gnd.n3813 0.152939
R20619 gnd.n3814 gnd.n3803 0.152939
R20620 gnd.n3822 gnd.n3803 0.152939
R20621 gnd.n3823 gnd.n3822 0.152939
R20622 gnd.n3824 gnd.n3823 0.152939
R20623 gnd.n3824 gnd.n3801 0.152939
R20624 gnd.n3832 gnd.n3801 0.152939
R20625 gnd.n3833 gnd.n3832 0.152939
R20626 gnd.n3834 gnd.n3833 0.152939
R20627 gnd.n3834 gnd.n3799 0.152939
R20628 gnd.n3842 gnd.n3799 0.152939
R20629 gnd.n4718 gnd.n2030 0.152939
R20630 gnd.n2032 gnd.n2030 0.152939
R20631 gnd.n2033 gnd.n2032 0.152939
R20632 gnd.n2034 gnd.n2033 0.152939
R20633 gnd.n2035 gnd.n2034 0.152939
R20634 gnd.n2036 gnd.n2035 0.152939
R20635 gnd.n2037 gnd.n2036 0.152939
R20636 gnd.n2038 gnd.n2037 0.152939
R20637 gnd.n2039 gnd.n2038 0.152939
R20638 gnd.n2040 gnd.n2039 0.152939
R20639 gnd.n2041 gnd.n2040 0.152939
R20640 gnd.n2042 gnd.n2041 0.152939
R20641 gnd.n2043 gnd.n2042 0.152939
R20642 gnd.n2044 gnd.n2043 0.152939
R20643 gnd.n2045 gnd.n2044 0.152939
R20644 gnd.n2046 gnd.n2045 0.152939
R20645 gnd.n2047 gnd.n2046 0.152939
R20646 gnd.n2048 gnd.n2047 0.152939
R20647 gnd.n2049 gnd.n2048 0.152939
R20648 gnd.n2050 gnd.n2049 0.152939
R20649 gnd.n2051 gnd.n2050 0.152939
R20650 gnd.n2052 gnd.n2051 0.152939
R20651 gnd.n2056 gnd.n2052 0.152939
R20652 gnd.n2057 gnd.n2056 0.152939
R20653 gnd.n2058 gnd.n2057 0.152939
R20654 gnd.n2059 gnd.n2058 0.152939
R20655 gnd.n3536 gnd.n3535 0.152939
R20656 gnd.n3537 gnd.n3536 0.152939
R20657 gnd.n3538 gnd.n3537 0.152939
R20658 gnd.n3539 gnd.n3538 0.152939
R20659 gnd.n3540 gnd.n3539 0.152939
R20660 gnd.n3541 gnd.n3540 0.152939
R20661 gnd.n3542 gnd.n3541 0.152939
R20662 gnd.n3543 gnd.n3542 0.152939
R20663 gnd.n3544 gnd.n3543 0.152939
R20664 gnd.n3545 gnd.n3544 0.152939
R20665 gnd.n3546 gnd.n3545 0.152939
R20666 gnd.n3547 gnd.n3546 0.152939
R20667 gnd.n3548 gnd.n3547 0.152939
R20668 gnd.n3549 gnd.n3548 0.152939
R20669 gnd.n3550 gnd.n3549 0.152939
R20670 gnd.n3551 gnd.n3550 0.152939
R20671 gnd.n3552 gnd.n3551 0.152939
R20672 gnd.n3553 gnd.n3552 0.152939
R20673 gnd.n3554 gnd.n3553 0.152939
R20674 gnd.n3555 gnd.n3554 0.152939
R20675 gnd.n3556 gnd.n3555 0.152939
R20676 gnd.n3557 gnd.n3556 0.152939
R20677 gnd.n3558 gnd.n3557 0.152939
R20678 gnd.n3559 gnd.n3558 0.152939
R20679 gnd.n3560 gnd.n3559 0.152939
R20680 gnd.n3561 gnd.n3560 0.152939
R20681 gnd.n3563 gnd.n3561 0.152939
R20682 gnd.n3563 gnd.n3562 0.152939
R20683 gnd.n3972 gnd.n3971 0.152939
R20684 gnd.n3972 gnd.n3862 0.152939
R20685 gnd.n3987 gnd.n3862 0.152939
R20686 gnd.n3988 gnd.n3987 0.152939
R20687 gnd.n3989 gnd.n3988 0.152939
R20688 gnd.n3989 gnd.n3850 0.152939
R20689 gnd.n4003 gnd.n3850 0.152939
R20690 gnd.n4004 gnd.n4003 0.152939
R20691 gnd.n4005 gnd.n4004 0.152939
R20692 gnd.n4006 gnd.n4005 0.152939
R20693 gnd.n4007 gnd.n4006 0.152939
R20694 gnd.n4008 gnd.n4007 0.152939
R20695 gnd.n4009 gnd.n4008 0.152939
R20696 gnd.n4010 gnd.n4009 0.152939
R20697 gnd.n4011 gnd.n4010 0.152939
R20698 gnd.n4012 gnd.n4011 0.152939
R20699 gnd.n4013 gnd.n4012 0.152939
R20700 gnd.n4014 gnd.n4013 0.152939
R20701 gnd.n4015 gnd.n4014 0.152939
R20702 gnd.n4016 gnd.n4015 0.152939
R20703 gnd.n4017 gnd.n4016 0.152939
R20704 gnd.n4017 gnd.n3715 0.152939
R20705 gnd.n4140 gnd.n3715 0.152939
R20706 gnd.n4141 gnd.n4140 0.152939
R20707 gnd.n4142 gnd.n4141 0.152939
R20708 gnd.n4143 gnd.n4142 0.152939
R20709 gnd.n4143 gnd.n3678 0.152939
R20710 gnd.n4188 gnd.n3678 0.152939
R20711 gnd.n3890 gnd.n3889 0.152939
R20712 gnd.n3891 gnd.n3890 0.152939
R20713 gnd.n3892 gnd.n3891 0.152939
R20714 gnd.n3893 gnd.n3892 0.152939
R20715 gnd.n3894 gnd.n3893 0.152939
R20716 gnd.n3895 gnd.n3894 0.152939
R20717 gnd.n3896 gnd.n3895 0.152939
R20718 gnd.n3897 gnd.n3896 0.152939
R20719 gnd.n3898 gnd.n3897 0.152939
R20720 gnd.n3899 gnd.n3898 0.152939
R20721 gnd.n3900 gnd.n3899 0.152939
R20722 gnd.n3901 gnd.n3900 0.152939
R20723 gnd.n3902 gnd.n3901 0.152939
R20724 gnd.n3903 gnd.n3902 0.152939
R20725 gnd.n3904 gnd.n3903 0.152939
R20726 gnd.n3905 gnd.n3904 0.152939
R20727 gnd.n3906 gnd.n3905 0.152939
R20728 gnd.n3907 gnd.n3906 0.152939
R20729 gnd.n3908 gnd.n3907 0.152939
R20730 gnd.n3909 gnd.n3908 0.152939
R20731 gnd.n3910 gnd.n3909 0.152939
R20732 gnd.n3911 gnd.n3910 0.152939
R20733 gnd.n3915 gnd.n3911 0.152939
R20734 gnd.n3916 gnd.n3915 0.152939
R20735 gnd.n3916 gnd.n3873 0.152939
R20736 gnd.n3970 gnd.n3873 0.152939
R20737 gnd.n3138 gnd.n3137 0.152939
R20738 gnd.n3137 gnd.n3136 0.152939
R20739 gnd.n3136 gnd.n2192 0.152939
R20740 gnd.n2197 gnd.n2192 0.152939
R20741 gnd.n2198 gnd.n2197 0.152939
R20742 gnd.n2199 gnd.n2198 0.152939
R20743 gnd.n2204 gnd.n2199 0.152939
R20744 gnd.n2205 gnd.n2204 0.152939
R20745 gnd.n2206 gnd.n2205 0.152939
R20746 gnd.n2207 gnd.n2206 0.152939
R20747 gnd.n2212 gnd.n2207 0.152939
R20748 gnd.n2213 gnd.n2212 0.152939
R20749 gnd.n2214 gnd.n2213 0.152939
R20750 gnd.n2215 gnd.n2214 0.152939
R20751 gnd.n2220 gnd.n2215 0.152939
R20752 gnd.n2221 gnd.n2220 0.152939
R20753 gnd.n2222 gnd.n2221 0.152939
R20754 gnd.n2223 gnd.n2222 0.152939
R20755 gnd.n2228 gnd.n2223 0.152939
R20756 gnd.n2229 gnd.n2228 0.152939
R20757 gnd.n2230 gnd.n2229 0.152939
R20758 gnd.n2231 gnd.n2230 0.152939
R20759 gnd.n2236 gnd.n2231 0.152939
R20760 gnd.n2237 gnd.n2236 0.152939
R20761 gnd.n2238 gnd.n2237 0.152939
R20762 gnd.n2239 gnd.n2238 0.152939
R20763 gnd.n2244 gnd.n2239 0.152939
R20764 gnd.n2245 gnd.n2244 0.152939
R20765 gnd.n2246 gnd.n2245 0.152939
R20766 gnd.n2247 gnd.n2246 0.152939
R20767 gnd.n2252 gnd.n2247 0.152939
R20768 gnd.n2253 gnd.n2252 0.152939
R20769 gnd.n2254 gnd.n2253 0.152939
R20770 gnd.n2255 gnd.n2254 0.152939
R20771 gnd.n2260 gnd.n2255 0.152939
R20772 gnd.n2261 gnd.n2260 0.152939
R20773 gnd.n2262 gnd.n2261 0.152939
R20774 gnd.n2263 gnd.n2262 0.152939
R20775 gnd.n2268 gnd.n2263 0.152939
R20776 gnd.n2269 gnd.n2268 0.152939
R20777 gnd.n2270 gnd.n2269 0.152939
R20778 gnd.n2271 gnd.n2270 0.152939
R20779 gnd.n2276 gnd.n2271 0.152939
R20780 gnd.n2277 gnd.n2276 0.152939
R20781 gnd.n2278 gnd.n2277 0.152939
R20782 gnd.n2279 gnd.n2278 0.152939
R20783 gnd.n2284 gnd.n2279 0.152939
R20784 gnd.n2285 gnd.n2284 0.152939
R20785 gnd.n2286 gnd.n2285 0.152939
R20786 gnd.n2287 gnd.n2286 0.152939
R20787 gnd.n2292 gnd.n2287 0.152939
R20788 gnd.n2293 gnd.n2292 0.152939
R20789 gnd.n2294 gnd.n2293 0.152939
R20790 gnd.n2295 gnd.n2294 0.152939
R20791 gnd.n2300 gnd.n2295 0.152939
R20792 gnd.n2301 gnd.n2300 0.152939
R20793 gnd.n2302 gnd.n2301 0.152939
R20794 gnd.n2303 gnd.n2302 0.152939
R20795 gnd.n2308 gnd.n2303 0.152939
R20796 gnd.n2309 gnd.n2308 0.152939
R20797 gnd.n2310 gnd.n2309 0.152939
R20798 gnd.n2311 gnd.n2310 0.152939
R20799 gnd.n2316 gnd.n2311 0.152939
R20800 gnd.n2317 gnd.n2316 0.152939
R20801 gnd.n2318 gnd.n2317 0.152939
R20802 gnd.n2319 gnd.n2318 0.152939
R20803 gnd.n2324 gnd.n2319 0.152939
R20804 gnd.n2325 gnd.n2324 0.152939
R20805 gnd.n2326 gnd.n2325 0.152939
R20806 gnd.n2327 gnd.n2326 0.152939
R20807 gnd.n2332 gnd.n2327 0.152939
R20808 gnd.n2333 gnd.n2332 0.152939
R20809 gnd.n2334 gnd.n2333 0.152939
R20810 gnd.n2335 gnd.n2334 0.152939
R20811 gnd.n2340 gnd.n2335 0.152939
R20812 gnd.n2341 gnd.n2340 0.152939
R20813 gnd.n2342 gnd.n2341 0.152939
R20814 gnd.n2343 gnd.n2342 0.152939
R20815 gnd.n2348 gnd.n2343 0.152939
R20816 gnd.n2349 gnd.n2348 0.152939
R20817 gnd.n2350 gnd.n2349 0.152939
R20818 gnd.n2351 gnd.n2350 0.152939
R20819 gnd.n2356 gnd.n2351 0.152939
R20820 gnd.n2357 gnd.n2356 0.152939
R20821 gnd.n2358 gnd.n2357 0.152939
R20822 gnd.n2359 gnd.n2358 0.152939
R20823 gnd.n2364 gnd.n2359 0.152939
R20824 gnd.n2365 gnd.n2364 0.152939
R20825 gnd.n2366 gnd.n2365 0.152939
R20826 gnd.n2367 gnd.n2366 0.152939
R20827 gnd.n2372 gnd.n2367 0.152939
R20828 gnd.n2373 gnd.n2372 0.152939
R20829 gnd.n2374 gnd.n2373 0.152939
R20830 gnd.n2375 gnd.n2374 0.152939
R20831 gnd.n2380 gnd.n2375 0.152939
R20832 gnd.n2381 gnd.n2380 0.152939
R20833 gnd.n2382 gnd.n2381 0.152939
R20834 gnd.n2383 gnd.n2382 0.152939
R20835 gnd.n2388 gnd.n2383 0.152939
R20836 gnd.n2389 gnd.n2388 0.152939
R20837 gnd.n2390 gnd.n2389 0.152939
R20838 gnd.n2391 gnd.n2390 0.152939
R20839 gnd.n2396 gnd.n2391 0.152939
R20840 gnd.n2397 gnd.n2396 0.152939
R20841 gnd.n2398 gnd.n2397 0.152939
R20842 gnd.n2399 gnd.n2398 0.152939
R20843 gnd.n2404 gnd.n2399 0.152939
R20844 gnd.n2405 gnd.n2404 0.152939
R20845 gnd.n2406 gnd.n2405 0.152939
R20846 gnd.n2407 gnd.n2406 0.152939
R20847 gnd.n2412 gnd.n2407 0.152939
R20848 gnd.n2413 gnd.n2412 0.152939
R20849 gnd.n2414 gnd.n2413 0.152939
R20850 gnd.n2415 gnd.n2414 0.152939
R20851 gnd.n2420 gnd.n2415 0.152939
R20852 gnd.n2421 gnd.n2420 0.152939
R20853 gnd.n2422 gnd.n2421 0.152939
R20854 gnd.n2423 gnd.n2422 0.152939
R20855 gnd.n2428 gnd.n2423 0.152939
R20856 gnd.n2429 gnd.n2428 0.152939
R20857 gnd.n2430 gnd.n2429 0.152939
R20858 gnd.n2431 gnd.n2430 0.152939
R20859 gnd.n2436 gnd.n2431 0.152939
R20860 gnd.n2437 gnd.n2436 0.152939
R20861 gnd.n2438 gnd.n2437 0.152939
R20862 gnd.n2439 gnd.n2438 0.152939
R20863 gnd.n2444 gnd.n2439 0.152939
R20864 gnd.n2445 gnd.n2444 0.152939
R20865 gnd.n2446 gnd.n2445 0.152939
R20866 gnd.n2447 gnd.n2446 0.152939
R20867 gnd.n2452 gnd.n2447 0.152939
R20868 gnd.n2453 gnd.n2452 0.152939
R20869 gnd.n2454 gnd.n2453 0.152939
R20870 gnd.n2455 gnd.n2454 0.152939
R20871 gnd.n2460 gnd.n2455 0.152939
R20872 gnd.n2461 gnd.n2460 0.152939
R20873 gnd.n2462 gnd.n2461 0.152939
R20874 gnd.n2463 gnd.n2462 0.152939
R20875 gnd.n2468 gnd.n2463 0.152939
R20876 gnd.n2469 gnd.n2468 0.152939
R20877 gnd.n2470 gnd.n2469 0.152939
R20878 gnd.n2471 gnd.n2470 0.152939
R20879 gnd.n2476 gnd.n2471 0.152939
R20880 gnd.n2477 gnd.n2476 0.152939
R20881 gnd.n2478 gnd.n2477 0.152939
R20882 gnd.n2479 gnd.n2478 0.152939
R20883 gnd.n2484 gnd.n2479 0.152939
R20884 gnd.n2485 gnd.n2484 0.152939
R20885 gnd.n2486 gnd.n2485 0.152939
R20886 gnd.n2487 gnd.n2486 0.152939
R20887 gnd.n2492 gnd.n2487 0.152939
R20888 gnd.n2493 gnd.n2492 0.152939
R20889 gnd.n2494 gnd.n2493 0.152939
R20890 gnd.n2495 gnd.n2494 0.152939
R20891 gnd.n2824 gnd.n2501 0.152939
R20892 gnd.n2824 gnd.n2823 0.152939
R20893 gnd.n2823 gnd.n2822 0.152939
R20894 gnd.n2822 gnd.n2502 0.152939
R20895 gnd.n2507 gnd.n2502 0.152939
R20896 gnd.n2508 gnd.n2507 0.152939
R20897 gnd.n2509 gnd.n2508 0.152939
R20898 gnd.n2514 gnd.n2509 0.152939
R20899 gnd.n2515 gnd.n2514 0.152939
R20900 gnd.n2516 gnd.n2515 0.152939
R20901 gnd.n2517 gnd.n2516 0.152939
R20902 gnd.n2522 gnd.n2517 0.152939
R20903 gnd.n2523 gnd.n2522 0.152939
R20904 gnd.n2524 gnd.n2523 0.152939
R20905 gnd.n2525 gnd.n2524 0.152939
R20906 gnd.n2530 gnd.n2525 0.152939
R20907 gnd.n2531 gnd.n2530 0.152939
R20908 gnd.n2532 gnd.n2531 0.152939
R20909 gnd.n2533 gnd.n2532 0.152939
R20910 gnd.n2538 gnd.n2533 0.152939
R20911 gnd.n2539 gnd.n2538 0.152939
R20912 gnd.n2540 gnd.n2539 0.152939
R20913 gnd.n2541 gnd.n2540 0.152939
R20914 gnd.n2546 gnd.n2541 0.152939
R20915 gnd.n2547 gnd.n2546 0.152939
R20916 gnd.n2548 gnd.n2547 0.152939
R20917 gnd.n2549 gnd.n2548 0.152939
R20918 gnd.n2554 gnd.n2549 0.152939
R20919 gnd.n2555 gnd.n2554 0.152939
R20920 gnd.n2556 gnd.n2555 0.152939
R20921 gnd.n2557 gnd.n2556 0.152939
R20922 gnd.n2562 gnd.n2557 0.152939
R20923 gnd.n2563 gnd.n2562 0.152939
R20924 gnd.n2564 gnd.n2563 0.152939
R20925 gnd.n2565 gnd.n2564 0.152939
R20926 gnd.n2570 gnd.n2565 0.152939
R20927 gnd.n2571 gnd.n2570 0.152939
R20928 gnd.n2572 gnd.n2571 0.152939
R20929 gnd.n2573 gnd.n2572 0.152939
R20930 gnd.n2578 gnd.n2573 0.152939
R20931 gnd.n2579 gnd.n2578 0.152939
R20932 gnd.n2580 gnd.n2579 0.152939
R20933 gnd.n2581 gnd.n2580 0.152939
R20934 gnd.n2586 gnd.n2581 0.152939
R20935 gnd.n2587 gnd.n2586 0.152939
R20936 gnd.n2588 gnd.n2587 0.152939
R20937 gnd.n2589 gnd.n2588 0.152939
R20938 gnd.n2594 gnd.n2589 0.152939
R20939 gnd.n2595 gnd.n2594 0.152939
R20940 gnd.n2596 gnd.n2595 0.152939
R20941 gnd.n2597 gnd.n2596 0.152939
R20942 gnd.n2602 gnd.n2597 0.152939
R20943 gnd.n2603 gnd.n2602 0.152939
R20944 gnd.n2604 gnd.n2603 0.152939
R20945 gnd.n2605 gnd.n2604 0.152939
R20946 gnd.n2610 gnd.n2605 0.152939
R20947 gnd.n2611 gnd.n2610 0.152939
R20948 gnd.n2612 gnd.n2611 0.152939
R20949 gnd.n2613 gnd.n2612 0.152939
R20950 gnd.n2618 gnd.n2613 0.152939
R20951 gnd.n2619 gnd.n2618 0.152939
R20952 gnd.n2620 gnd.n2619 0.152939
R20953 gnd.n2621 gnd.n2620 0.152939
R20954 gnd.n2626 gnd.n2621 0.152939
R20955 gnd.n2627 gnd.n2626 0.152939
R20956 gnd.n2628 gnd.n2627 0.152939
R20957 gnd.n2629 gnd.n2628 0.152939
R20958 gnd.n2634 gnd.n2629 0.152939
R20959 gnd.n2635 gnd.n2634 0.152939
R20960 gnd.n2636 gnd.n2635 0.152939
R20961 gnd.n2637 gnd.n2636 0.152939
R20962 gnd.n2642 gnd.n2637 0.152939
R20963 gnd.n2643 gnd.n2642 0.152939
R20964 gnd.n2644 gnd.n2643 0.152939
R20965 gnd.n2645 gnd.n2644 0.152939
R20966 gnd.n2650 gnd.n2645 0.152939
R20967 gnd.n2651 gnd.n2650 0.152939
R20968 gnd.n2652 gnd.n2651 0.152939
R20969 gnd.n2653 gnd.n2652 0.152939
R20970 gnd.n2659 gnd.n2653 0.152939
R20971 gnd.n2660 gnd.n2659 0.152939
R20972 gnd.n2661 gnd.n2660 0.152939
R20973 gnd.n2661 gnd.n345 0.152939
R20974 gnd.n7218 gnd.n345 0.152939
R20975 gnd.n7326 gnd.n7325 0.152939
R20976 gnd.n7326 gnd.n283 0.152939
R20977 gnd.n7340 gnd.n283 0.152939
R20978 gnd.n7341 gnd.n7340 0.152939
R20979 gnd.n7342 gnd.n7341 0.152939
R20980 gnd.n7342 gnd.n269 0.152939
R20981 gnd.n7356 gnd.n269 0.152939
R20982 gnd.n7357 gnd.n7356 0.152939
R20983 gnd.n7358 gnd.n7357 0.152939
R20984 gnd.n7358 gnd.n253 0.152939
R20985 gnd.n7372 gnd.n253 0.152939
R20986 gnd.n7373 gnd.n7372 0.152939
R20987 gnd.n7374 gnd.n7373 0.152939
R20988 gnd.n7374 gnd.n239 0.152939
R20989 gnd.n7388 gnd.n239 0.152939
R20990 gnd.n7389 gnd.n7388 0.152939
R20991 gnd.n7390 gnd.n7389 0.152939
R20992 gnd.n7390 gnd.n222 0.152939
R20993 gnd.n7404 gnd.n222 0.152939
R20994 gnd.n7405 gnd.n7404 0.152939
R20995 gnd.n7406 gnd.n7405 0.152939
R20996 gnd.n7406 gnd.n206 0.152939
R20997 gnd.n7488 gnd.n206 0.152939
R20998 gnd.n7489 gnd.n7488 0.152939
R20999 gnd.n7490 gnd.n7489 0.152939
R21000 gnd.n7490 gnd.n129 0.152939
R21001 gnd.n7570 gnd.n129 0.152939
R21002 gnd.n7569 gnd.n130 0.152939
R21003 gnd.n132 gnd.n130 0.152939
R21004 gnd.n136 gnd.n132 0.152939
R21005 gnd.n137 gnd.n136 0.152939
R21006 gnd.n138 gnd.n137 0.152939
R21007 gnd.n139 gnd.n138 0.152939
R21008 gnd.n143 gnd.n139 0.152939
R21009 gnd.n144 gnd.n143 0.152939
R21010 gnd.n145 gnd.n144 0.152939
R21011 gnd.n146 gnd.n145 0.152939
R21012 gnd.n150 gnd.n146 0.152939
R21013 gnd.n151 gnd.n150 0.152939
R21014 gnd.n152 gnd.n151 0.152939
R21015 gnd.n153 gnd.n152 0.152939
R21016 gnd.n157 gnd.n153 0.152939
R21017 gnd.n158 gnd.n157 0.152939
R21018 gnd.n159 gnd.n158 0.152939
R21019 gnd.n160 gnd.n159 0.152939
R21020 gnd.n164 gnd.n160 0.152939
R21021 gnd.n165 gnd.n164 0.152939
R21022 gnd.n166 gnd.n165 0.152939
R21023 gnd.n167 gnd.n166 0.152939
R21024 gnd.n171 gnd.n167 0.152939
R21025 gnd.n172 gnd.n171 0.152939
R21026 gnd.n173 gnd.n172 0.152939
R21027 gnd.n174 gnd.n173 0.152939
R21028 gnd.n178 gnd.n174 0.152939
R21029 gnd.n179 gnd.n178 0.152939
R21030 gnd.n180 gnd.n179 0.152939
R21031 gnd.n181 gnd.n180 0.152939
R21032 gnd.n185 gnd.n181 0.152939
R21033 gnd.n186 gnd.n185 0.152939
R21034 gnd.n187 gnd.n186 0.152939
R21035 gnd.n188 gnd.n187 0.152939
R21036 gnd.n192 gnd.n188 0.152939
R21037 gnd.n193 gnd.n192 0.152939
R21038 gnd.n7500 gnd.n193 0.152939
R21039 gnd.n7500 gnd.n7499 0.152939
R21040 gnd.n6844 gnd.n562 0.152939
R21041 gnd.n6845 gnd.n6844 0.152939
R21042 gnd.n6845 gnd.n6842 0.152939
R21043 gnd.n6853 gnd.n6842 0.152939
R21044 gnd.n6854 gnd.n6853 0.152939
R21045 gnd.n6855 gnd.n6854 0.152939
R21046 gnd.n6856 gnd.n6855 0.152939
R21047 gnd.n6858 gnd.n6856 0.152939
R21048 gnd.n6858 gnd.n6857 0.152939
R21049 gnd.n6857 gnd.n597 0.152939
R21050 gnd.n597 gnd.n595 0.152939
R21051 gnd.n6893 gnd.n595 0.152939
R21052 gnd.n6894 gnd.n6893 0.152939
R21053 gnd.n6895 gnd.n6894 0.152939
R21054 gnd.n6896 gnd.n6895 0.152939
R21055 gnd.n6897 gnd.n6896 0.152939
R21056 gnd.n6897 gnd.n586 0.152939
R21057 gnd.n6920 gnd.n586 0.152939
R21058 gnd.n6921 gnd.n6920 0.152939
R21059 gnd.n6922 gnd.n6921 0.152939
R21060 gnd.n6923 gnd.n6922 0.152939
R21061 gnd.n6924 gnd.n6923 0.152939
R21062 gnd.n6925 gnd.n6924 0.152939
R21063 gnd.n6926 gnd.n6925 0.152939
R21064 gnd.n6928 gnd.n6926 0.152939
R21065 gnd.n6928 gnd.n6927 0.152939
R21066 gnd.n6927 gnd.n356 0.152939
R21067 gnd.n7195 gnd.n356 0.152939
R21068 gnd.n7196 gnd.n7195 0.152939
R21069 gnd.n7197 gnd.n7196 0.152939
R21070 gnd.n7198 gnd.n7197 0.152939
R21071 gnd.n7198 gnd.n333 0.152939
R21072 gnd.n7231 gnd.n333 0.152939
R21073 gnd.n7232 gnd.n7231 0.152939
R21074 gnd.n7233 gnd.n7232 0.152939
R21075 gnd.n7234 gnd.n7233 0.152939
R21076 gnd.n7235 gnd.n7234 0.152939
R21077 gnd.n7236 gnd.n7235 0.152939
R21078 gnd.n7237 gnd.n7236 0.152939
R21079 gnd.n7238 gnd.n7237 0.152939
R21080 gnd.n7239 gnd.n7238 0.152939
R21081 gnd.n7240 gnd.n7239 0.152939
R21082 gnd.n7241 gnd.n7240 0.152939
R21083 gnd.n7242 gnd.n7241 0.152939
R21084 gnd.n7243 gnd.n7242 0.152939
R21085 gnd.n7244 gnd.n7243 0.152939
R21086 gnd.n7245 gnd.n7244 0.152939
R21087 gnd.n7246 gnd.n7245 0.152939
R21088 gnd.n7247 gnd.n7246 0.152939
R21089 gnd.n7248 gnd.n7247 0.152939
R21090 gnd.n7249 gnd.n7248 0.152939
R21091 gnd.n7250 gnd.n7249 0.152939
R21092 gnd.n7251 gnd.n7250 0.152939
R21093 gnd.n7252 gnd.n7251 0.152939
R21094 gnd.n7253 gnd.n7252 0.152939
R21095 gnd.n7254 gnd.n7253 0.152939
R21096 gnd.n7255 gnd.n7254 0.152939
R21097 gnd.n7256 gnd.n7255 0.152939
R21098 gnd.n7257 gnd.n7256 0.152939
R21099 gnd.n7258 gnd.n7257 0.152939
R21100 gnd.n7260 gnd.n7258 0.152939
R21101 gnd.n7260 gnd.n7259 0.152939
R21102 gnd.n7259 gnd.n199 0.152939
R21103 gnd.n7498 gnd.n199 0.152939
R21104 gnd.n7050 gnd.n486 0.152939
R21105 gnd.n520 gnd.n486 0.152939
R21106 gnd.n521 gnd.n520 0.152939
R21107 gnd.n522 gnd.n521 0.152939
R21108 gnd.n523 gnd.n522 0.152939
R21109 gnd.n524 gnd.n523 0.152939
R21110 gnd.n525 gnd.n524 0.152939
R21111 gnd.n526 gnd.n525 0.152939
R21112 gnd.n527 gnd.n526 0.152939
R21113 gnd.n528 gnd.n527 0.152939
R21114 gnd.n529 gnd.n528 0.152939
R21115 gnd.n530 gnd.n529 0.152939
R21116 gnd.n531 gnd.n530 0.152939
R21117 gnd.n532 gnd.n531 0.152939
R21118 gnd.n533 gnd.n532 0.152939
R21119 gnd.n540 gnd.n539 0.152939
R21120 gnd.n541 gnd.n540 0.152939
R21121 gnd.n542 gnd.n541 0.152939
R21122 gnd.n543 gnd.n542 0.152939
R21123 gnd.n544 gnd.n543 0.152939
R21124 gnd.n545 gnd.n544 0.152939
R21125 gnd.n546 gnd.n545 0.152939
R21126 gnd.n547 gnd.n546 0.152939
R21127 gnd.n548 gnd.n547 0.152939
R21128 gnd.n549 gnd.n548 0.152939
R21129 gnd.n550 gnd.n549 0.152939
R21130 gnd.n551 gnd.n550 0.152939
R21131 gnd.n552 gnd.n551 0.152939
R21132 gnd.n553 gnd.n552 0.152939
R21133 gnd.n554 gnd.n553 0.152939
R21134 gnd.n555 gnd.n554 0.152939
R21135 gnd.n556 gnd.n555 0.152939
R21136 gnd.n6980 gnd.n556 0.152939
R21137 gnd.n6980 gnd.n6979 0.152939
R21138 gnd.n6979 gnd.n6978 0.152939
R21139 gnd.n7052 gnd.n7051 0.152939
R21140 gnd.n7052 gnd.n468 0.152939
R21141 gnd.n7066 gnd.n468 0.152939
R21142 gnd.n7067 gnd.n7066 0.152939
R21143 gnd.n7068 gnd.n7067 0.152939
R21144 gnd.n7068 gnd.n451 0.152939
R21145 gnd.n7082 gnd.n451 0.152939
R21146 gnd.n7083 gnd.n7082 0.152939
R21147 gnd.n7084 gnd.n7083 0.152939
R21148 gnd.n7084 gnd.n434 0.152939
R21149 gnd.n7098 gnd.n434 0.152939
R21150 gnd.n7099 gnd.n7098 0.152939
R21151 gnd.n7100 gnd.n7099 0.152939
R21152 gnd.n7100 gnd.n417 0.152939
R21153 gnd.n7114 gnd.n417 0.152939
R21154 gnd.n7115 gnd.n7114 0.152939
R21155 gnd.n7116 gnd.n7115 0.152939
R21156 gnd.n7116 gnd.n398 0.152939
R21157 gnd.n7133 gnd.n398 0.152939
R21158 gnd.n7134 gnd.n7133 0.152939
R21159 gnd.n7135 gnd.n7134 0.152939
R21160 gnd.n7135 gnd.n366 0.152939
R21161 gnd.n7184 gnd.n366 0.152939
R21162 gnd.n7185 gnd.n7184 0.152939
R21163 gnd.n7186 gnd.n7185 0.152939
R21164 gnd.n7186 gnd.n299 0.152939
R21165 gnd.n7325 gnd.n299 0.152939
R21166 gnd.n7149 gnd.n7148 0.152939
R21167 gnd.n7148 gnd.n347 0.152939
R21168 gnd.n1803 gnd.n1802 0.152939
R21169 gnd.n5258 gnd.n1803 0.152939
R21170 gnd.n5260 gnd.n5258 0.152939
R21171 gnd.n5261 gnd.n5260 0.152939
R21172 gnd.n5262 gnd.n5261 0.152939
R21173 gnd.n5263 gnd.n5262 0.152939
R21174 gnd.n5264 gnd.n5263 0.152939
R21175 gnd.n5265 gnd.n5264 0.152939
R21176 gnd.n5266 gnd.n5265 0.152939
R21177 gnd.n5266 gnd.n1847 0.152939
R21178 gnd.n5300 gnd.n1847 0.152939
R21179 gnd.n5301 gnd.n5300 0.152939
R21180 gnd.n5302 gnd.n5301 0.152939
R21181 gnd.n5303 gnd.n5302 0.152939
R21182 gnd.n5304 gnd.n5303 0.152939
R21183 gnd.n5305 gnd.n5304 0.152939
R21184 gnd.n5306 gnd.n5305 0.152939
R21185 gnd.n5306 gnd.n1837 0.152939
R21186 gnd.n5339 gnd.n1837 0.152939
R21187 gnd.n5340 gnd.n5339 0.152939
R21188 gnd.n5341 gnd.n5340 0.152939
R21189 gnd.n5342 gnd.n5341 0.152939
R21190 gnd.n5343 gnd.n5342 0.152939
R21191 gnd.n5346 gnd.n5343 0.152939
R21192 gnd.n5347 gnd.n5346 0.152939
R21193 gnd.n5348 gnd.n5347 0.152939
R21194 gnd.n5349 gnd.n5348 0.152939
R21195 gnd.n5353 gnd.n5349 0.152939
R21196 gnd.n5354 gnd.n5353 0.152939
R21197 gnd.n5355 gnd.n5354 0.152939
R21198 gnd.n5355 gnd.n1315 0.152939
R21199 gnd.n5812 gnd.n1315 0.152939
R21200 gnd.n5813 gnd.n5812 0.152939
R21201 gnd.n5814 gnd.n5813 0.152939
R21202 gnd.n5814 gnd.n1301 0.152939
R21203 gnd.n5828 gnd.n1301 0.152939
R21204 gnd.n5829 gnd.n5828 0.152939
R21205 gnd.n5830 gnd.n5829 0.152939
R21206 gnd.n5831 gnd.n5830 0.152939
R21207 gnd.n5831 gnd.n1259 0.152939
R21208 gnd.n5986 gnd.n1259 0.152939
R21209 gnd.n5987 gnd.n5986 0.152939
R21210 gnd.n5988 gnd.n5987 0.152939
R21211 gnd.n5988 gnd.n1244 0.152939
R21212 gnd.n6002 gnd.n1244 0.152939
R21213 gnd.n6003 gnd.n6002 0.152939
R21214 gnd.n6004 gnd.n6003 0.152939
R21215 gnd.n6004 gnd.n1228 0.152939
R21216 gnd.n6018 gnd.n1228 0.152939
R21217 gnd.n6019 gnd.n6018 0.152939
R21218 gnd.n6020 gnd.n6019 0.152939
R21219 gnd.n6020 gnd.n1213 0.152939
R21220 gnd.n6033 gnd.n1213 0.152939
R21221 gnd.n6034 gnd.n6033 0.152939
R21222 gnd.n6035 gnd.n6034 0.152939
R21223 gnd.n6036 gnd.n6035 0.152939
R21224 gnd.n6036 gnd.n1106 0.152939
R21225 gnd.n6128 gnd.n1106 0.152939
R21226 gnd.n6129 gnd.n6128 0.152939
R21227 gnd.n6130 gnd.n6129 0.152939
R21228 gnd.n6130 gnd.n1090 0.152939
R21229 gnd.n6144 gnd.n1090 0.152939
R21230 gnd.n6145 gnd.n6144 0.152939
R21231 gnd.n6146 gnd.n6145 0.152939
R21232 gnd.n6146 gnd.n1075 0.152939
R21233 gnd.n6160 gnd.n1075 0.152939
R21234 gnd.n6161 gnd.n6160 0.152939
R21235 gnd.n6162 gnd.n6161 0.152939
R21236 gnd.n6162 gnd.n1062 0.152939
R21237 gnd.n6176 gnd.n1062 0.152939
R21238 gnd.n6177 gnd.n6176 0.152939
R21239 gnd.n6178 gnd.n6177 0.152939
R21240 gnd.n6179 gnd.n6178 0.152939
R21241 gnd.n6179 gnd.n1019 0.152939
R21242 gnd.n6433 gnd.n1019 0.152939
R21243 gnd.n6434 gnd.n6433 0.152939
R21244 gnd.n6435 gnd.n6434 0.152939
R21245 gnd.n6435 gnd.n1003 0.152939
R21246 gnd.n6449 gnd.n1003 0.152939
R21247 gnd.n6450 gnd.n6449 0.152939
R21248 gnd.n6451 gnd.n6450 0.152939
R21249 gnd.n6451 gnd.n987 0.152939
R21250 gnd.n6465 gnd.n987 0.152939
R21251 gnd.n6466 gnd.n6465 0.152939
R21252 gnd.n6467 gnd.n6466 0.152939
R21253 gnd.n6467 gnd.n973 0.152939
R21254 gnd.n6481 gnd.n973 0.152939
R21255 gnd.n6482 gnd.n6481 0.152939
R21256 gnd.n6483 gnd.n6482 0.152939
R21257 gnd.n6483 gnd.n958 0.152939
R21258 gnd.n6497 gnd.n958 0.152939
R21259 gnd.n6498 gnd.n6497 0.152939
R21260 gnd.n6499 gnd.n6498 0.152939
R21261 gnd.n6499 gnd.n942 0.152939
R21262 gnd.n6513 gnd.n942 0.152939
R21263 gnd.n6514 gnd.n6513 0.152939
R21264 gnd.n6515 gnd.n6514 0.152939
R21265 gnd.n6515 gnd.n925 0.152939
R21266 gnd.n6535 gnd.n925 0.152939
R21267 gnd.n6536 gnd.n6535 0.152939
R21268 gnd.n6537 gnd.n6536 0.152939
R21269 gnd.n6538 gnd.n6537 0.152939
R21270 gnd.n6538 gnd.n885 0.152939
R21271 gnd.n6593 gnd.n885 0.152939
R21272 gnd.n6594 gnd.n6593 0.152939
R21273 gnd.n6595 gnd.n6594 0.152939
R21274 gnd.n6596 gnd.n6595 0.152939
R21275 gnd.n6596 gnd.n658 0.152939
R21276 gnd.n6784 gnd.n658 0.152939
R21277 gnd.n6785 gnd.n6784 0.152939
R21278 gnd.n6786 gnd.n6785 0.152939
R21279 gnd.n6786 gnd.n643 0.152939
R21280 gnd.n6801 gnd.n643 0.152939
R21281 gnd.n6802 gnd.n6801 0.152939
R21282 gnd.n6803 gnd.n6802 0.152939
R21283 gnd.n6804 gnd.n6803 0.152939
R21284 gnd.n6804 gnd.n613 0.152939
R21285 gnd.n6820 gnd.n613 0.152939
R21286 gnd.n6821 gnd.n6820 0.152939
R21287 gnd.n6822 gnd.n6821 0.152939
R21288 gnd.n6822 gnd.n609 0.152939
R21289 gnd.n6828 gnd.n609 0.152939
R21290 gnd.n6829 gnd.n6828 0.152939
R21291 gnd.n6830 gnd.n6829 0.152939
R21292 gnd.n6830 gnd.n605 0.152939
R21293 gnd.n6836 gnd.n605 0.152939
R21294 gnd.n6837 gnd.n6836 0.152939
R21295 gnd.n6838 gnd.n6837 0.152939
R21296 gnd.n6838 gnd.n601 0.152939
R21297 gnd.n6870 gnd.n601 0.152939
R21298 gnd.n6871 gnd.n6870 0.152939
R21299 gnd.n6872 gnd.n6871 0.152939
R21300 gnd.n6873 gnd.n6872 0.152939
R21301 gnd.n6874 gnd.n6873 0.152939
R21302 gnd.n6875 gnd.n6874 0.152939
R21303 gnd.n6876 gnd.n6875 0.152939
R21304 gnd.n6876 gnd.n591 0.152939
R21305 gnd.n6909 gnd.n591 0.152939
R21306 gnd.n6910 gnd.n6909 0.152939
R21307 gnd.n6911 gnd.n6910 0.152939
R21308 gnd.n6912 gnd.n6911 0.152939
R21309 gnd.n6912 gnd.n391 0.152939
R21310 gnd.n7142 gnd.n391 0.152939
R21311 gnd.n7143 gnd.n7142 0.152939
R21312 gnd.n7144 gnd.n7143 0.152939
R21313 gnd.n7145 gnd.n7144 0.152939
R21314 gnd.n7146 gnd.n7145 0.152939
R21315 gnd.n7147 gnd.n7146 0.152939
R21316 gnd.n7149 gnd.n7147 0.152939
R21317 gnd.n4827 gnd.n4826 0.152939
R21318 gnd.n4828 gnd.n4827 0.152939
R21319 gnd.n4829 gnd.n4828 0.152939
R21320 gnd.n4830 gnd.n4829 0.152939
R21321 gnd.n4831 gnd.n4830 0.152939
R21322 gnd.n4832 gnd.n4831 0.152939
R21323 gnd.n4833 gnd.n4832 0.152939
R21324 gnd.n4834 gnd.n4833 0.152939
R21325 gnd.n4835 gnd.n4834 0.152939
R21326 gnd.n4836 gnd.n4835 0.152939
R21327 gnd.n4837 gnd.n4836 0.152939
R21328 gnd.n4838 gnd.n4837 0.152939
R21329 gnd.n4839 gnd.n4838 0.152939
R21330 gnd.n4840 gnd.n4839 0.152939
R21331 gnd.n4841 gnd.n4840 0.152939
R21332 gnd.n4842 gnd.n4841 0.152939
R21333 gnd.n4843 gnd.n4842 0.152939
R21334 gnd.n4844 gnd.n4843 0.152939
R21335 gnd.n4844 gnd.n1905 0.152939
R21336 gnd.n5163 gnd.n1905 0.152939
R21337 gnd.n5164 gnd.n5163 0.152939
R21338 gnd.n5165 gnd.n5164 0.152939
R21339 gnd.n5166 gnd.n5165 0.152939
R21340 gnd.n5167 gnd.n5166 0.152939
R21341 gnd.n5167 gnd.n1870 0.152939
R21342 gnd.n5202 gnd.n1870 0.152939
R21343 gnd.n5203 gnd.n5202 0.152939
R21344 gnd.n5204 gnd.n5203 0.152939
R21345 gnd.n5205 gnd.n5204 0.152939
R21346 gnd.n5206 gnd.n5205 0.152939
R21347 gnd.n5207 gnd.n5206 0.152939
R21348 gnd.n4778 gnd.n1986 0.152939
R21349 gnd.n4786 gnd.n4778 0.152939
R21350 gnd.n4787 gnd.n4786 0.152939
R21351 gnd.n4788 gnd.n4787 0.152939
R21352 gnd.n4788 gnd.n4774 0.152939
R21353 gnd.n4796 gnd.n4774 0.152939
R21354 gnd.n4797 gnd.n4796 0.152939
R21355 gnd.n4798 gnd.n4797 0.152939
R21356 gnd.n4798 gnd.n4770 0.152939
R21357 gnd.n4806 gnd.n4770 0.152939
R21358 gnd.n4807 gnd.n4806 0.152939
R21359 gnd.n4808 gnd.n4807 0.152939
R21360 gnd.n4808 gnd.n4766 0.152939
R21361 gnd.n4816 gnd.n4766 0.152939
R21362 gnd.n4817 gnd.n4816 0.152939
R21363 gnd.n4818 gnd.n4817 0.152939
R21364 gnd.n4818 gnd.n4760 0.152939
R21365 gnd.n4825 gnd.n4760 0.152939
R21366 gnd.n5074 gnd.n5073 0.152939
R21367 gnd.n5075 gnd.n5074 0.152939
R21368 gnd.n5075 gnd.n1971 0.152939
R21369 gnd.n5089 gnd.n1971 0.152939
R21370 gnd.n5090 gnd.n5089 0.152939
R21371 gnd.n5091 gnd.n5090 0.152939
R21372 gnd.n5091 gnd.n1954 0.152939
R21373 gnd.n5105 gnd.n1954 0.152939
R21374 gnd.n5106 gnd.n5105 0.152939
R21375 gnd.n5107 gnd.n5106 0.152939
R21376 gnd.n5107 gnd.n1939 0.152939
R21377 gnd.n5121 gnd.n1939 0.152939
R21378 gnd.n5122 gnd.n5121 0.152939
R21379 gnd.n5123 gnd.n5122 0.152939
R21380 gnd.n5123 gnd.n1922 0.152939
R21381 gnd.n5137 gnd.n1922 0.152939
R21382 gnd.n5138 gnd.n5137 0.152939
R21383 gnd.n5139 gnd.n5138 0.152939
R21384 gnd.n5140 gnd.n5139 0.152939
R21385 gnd.n5141 gnd.n5140 0.152939
R21386 gnd.n5143 gnd.n5141 0.152939
R21387 gnd.n5143 gnd.n5142 0.152939
R21388 gnd.n5142 gnd.n1888 0.152939
R21389 gnd.n1889 gnd.n1888 0.152939
R21390 gnd.n1890 gnd.n1889 0.152939
R21391 gnd.n1891 gnd.n1890 0.152939
R21392 gnd.n1893 gnd.n1891 0.152939
R21393 gnd.n1893 gnd.n1892 0.152939
R21394 gnd.n1892 gnd.n1779 0.152939
R21395 gnd.n1780 gnd.n1779 0.152939
R21396 gnd.n1781 gnd.n1780 0.152939
R21397 gnd.n1861 gnd.n1781 0.152939
R21398 gnd.n1861 gnd.n1792 0.152939
R21399 gnd.n1793 gnd.n1792 0.152939
R21400 gnd.n1794 gnd.n1793 0.152939
R21401 gnd.n1794 gnd.n1755 0.152939
R21402 gnd.n5472 gnd.n1755 0.152939
R21403 gnd.n5473 gnd.n5472 0.152939
R21404 gnd.n5474 gnd.n5473 0.152939
R21405 gnd.n5474 gnd.n1739 0.152939
R21406 gnd.n5488 gnd.n1739 0.152939
R21407 gnd.n5489 gnd.n5488 0.152939
R21408 gnd.n5490 gnd.n5489 0.152939
R21409 gnd.n5490 gnd.n1721 0.152939
R21410 gnd.n5504 gnd.n1721 0.152939
R21411 gnd.n5505 gnd.n5504 0.152939
R21412 gnd.n5506 gnd.n5505 0.152939
R21413 gnd.n5506 gnd.n1705 0.152939
R21414 gnd.n5520 gnd.n1705 0.152939
R21415 gnd.n5521 gnd.n5520 0.152939
R21416 gnd.n5522 gnd.n5521 0.152939
R21417 gnd.n5522 gnd.n1687 0.152939
R21418 gnd.n5536 gnd.n1687 0.152939
R21419 gnd.n5537 gnd.n5536 0.152939
R21420 gnd.n5538 gnd.n5537 0.152939
R21421 gnd.n5538 gnd.n1671 0.152939
R21422 gnd.n5552 gnd.n1671 0.152939
R21423 gnd.n5553 gnd.n5552 0.152939
R21424 gnd.n5554 gnd.n5553 0.152939
R21425 gnd.n5554 gnd.n1652 0.152939
R21426 gnd.n5570 gnd.n1652 0.152939
R21427 gnd.n5571 gnd.n5570 0.152939
R21428 gnd.n5572 gnd.n5571 0.152939
R21429 gnd.n5690 gnd.n5572 0.152939
R21430 gnd.n5466 gnd.n1747 0.152939
R21431 gnd.n5480 gnd.n1747 0.152939
R21432 gnd.n5481 gnd.n5480 0.152939
R21433 gnd.n5482 gnd.n5481 0.152939
R21434 gnd.n5482 gnd.n1730 0.152939
R21435 gnd.n5496 gnd.n1730 0.152939
R21436 gnd.n5497 gnd.n5496 0.152939
R21437 gnd.n5498 gnd.n5497 0.152939
R21438 gnd.n5498 gnd.n1713 0.152939
R21439 gnd.n5512 gnd.n1713 0.152939
R21440 gnd.n5513 gnd.n5512 0.152939
R21441 gnd.n5514 gnd.n5513 0.152939
R21442 gnd.n5514 gnd.n1696 0.152939
R21443 gnd.n5528 gnd.n1696 0.152939
R21444 gnd.n5529 gnd.n5528 0.152939
R21445 gnd.n5530 gnd.n5529 0.152939
R21446 gnd.n5530 gnd.n1679 0.152939
R21447 gnd.n5544 gnd.n1679 0.152939
R21448 gnd.n5545 gnd.n5544 0.152939
R21449 gnd.n5546 gnd.n5545 0.152939
R21450 gnd.n5546 gnd.n1662 0.152939
R21451 gnd.n5560 gnd.n1662 0.152939
R21452 gnd.n5561 gnd.n5560 0.152939
R21453 gnd.n5562 gnd.n5561 0.152939
R21454 gnd.n5563 gnd.n5562 0.152939
R21455 gnd.n5563 gnd.n1361 0.152939
R21456 gnd.n5768 gnd.n1361 0.152939
R21457 gnd.n5767 gnd.n1362 0.152939
R21458 gnd.n1367 gnd.n1362 0.152939
R21459 gnd.n1368 gnd.n1367 0.152939
R21460 gnd.n1369 gnd.n1368 0.152939
R21461 gnd.n1370 gnd.n1369 0.152939
R21462 gnd.n1371 gnd.n1370 0.152939
R21463 gnd.n1375 gnd.n1371 0.152939
R21464 gnd.n1376 gnd.n1375 0.152939
R21465 gnd.n1377 gnd.n1376 0.152939
R21466 gnd.n1378 gnd.n1377 0.152939
R21467 gnd.n1382 gnd.n1378 0.152939
R21468 gnd.n1383 gnd.n1382 0.152939
R21469 gnd.n1384 gnd.n1383 0.152939
R21470 gnd.n1385 gnd.n1384 0.152939
R21471 gnd.n1608 gnd.n1385 0.152939
R21472 gnd.n1611 gnd.n1610 0.152939
R21473 gnd.n1612 gnd.n1611 0.152939
R21474 gnd.n1616 gnd.n1612 0.152939
R21475 gnd.n1617 gnd.n1616 0.152939
R21476 gnd.n1618 gnd.n1617 0.152939
R21477 gnd.n1619 gnd.n1618 0.152939
R21478 gnd.n1623 gnd.n1619 0.152939
R21479 gnd.n1624 gnd.n1623 0.152939
R21480 gnd.n1625 gnd.n1624 0.152939
R21481 gnd.n1626 gnd.n1625 0.152939
R21482 gnd.n1630 gnd.n1626 0.152939
R21483 gnd.n1631 gnd.n1630 0.152939
R21484 gnd.n1632 gnd.n1631 0.152939
R21485 gnd.n1633 gnd.n1632 0.152939
R21486 gnd.n1637 gnd.n1633 0.152939
R21487 gnd.n1638 gnd.n1637 0.152939
R21488 gnd.n1639 gnd.n1638 0.152939
R21489 gnd.n1640 gnd.n1639 0.152939
R21490 gnd.n1645 gnd.n1640 0.152939
R21491 gnd.n5699 gnd.n1645 0.152939
R21492 gnd.n4987 gnd.n4935 0.152939
R21493 gnd.n4937 gnd.n4935 0.152939
R21494 gnd.n4938 gnd.n4937 0.152939
R21495 gnd.n4939 gnd.n4938 0.152939
R21496 gnd.n4940 gnd.n4939 0.152939
R21497 gnd.n4941 gnd.n4940 0.152939
R21498 gnd.n4942 gnd.n4941 0.152939
R21499 gnd.n4943 gnd.n4942 0.152939
R21500 gnd.n4944 gnd.n4943 0.152939
R21501 gnd.n4945 gnd.n4944 0.152939
R21502 gnd.n4946 gnd.n4945 0.152939
R21503 gnd.n4947 gnd.n4946 0.152939
R21504 gnd.n4948 gnd.n4947 0.152939
R21505 gnd.n4949 gnd.n4948 0.152939
R21506 gnd.n4950 gnd.n4949 0.152939
R21507 gnd.n4951 gnd.n4950 0.152939
R21508 gnd.n4952 gnd.n4951 0.152939
R21509 gnd.n4953 gnd.n4952 0.152939
R21510 gnd.n4954 gnd.n4953 0.152939
R21511 gnd.n4956 gnd.n4954 0.152939
R21512 gnd.n4956 gnd.n4955 0.152939
R21513 gnd.n4955 gnd.n1899 0.152939
R21514 gnd.n5177 gnd.n1899 0.152939
R21515 gnd.n5178 gnd.n5177 0.152939
R21516 gnd.n5179 gnd.n5178 0.152939
R21517 gnd.n5180 gnd.n5179 0.152939
R21518 gnd.n5180 gnd.n1864 0.152939
R21519 gnd.n5220 gnd.n1864 0.152939
R21520 gnd.n5221 gnd.n5220 0.152939
R21521 gnd.n5222 gnd.n5221 0.152939
R21522 gnd.n5222 gnd.n1862 0.152939
R21523 gnd.n5228 gnd.n1862 0.152939
R21524 gnd.n5229 gnd.n5228 0.152939
R21525 gnd.n5230 gnd.n5229 0.152939
R21526 gnd.n5230 gnd.n1855 0.152939
R21527 gnd.n5244 gnd.n1855 0.152939
R21528 gnd.n5245 gnd.n5244 0.152939
R21529 gnd.n5246 gnd.n5245 0.152939
R21530 gnd.n5246 gnd.n1853 0.152939
R21531 gnd.n5252 gnd.n1853 0.152939
R21532 gnd.n5253 gnd.n5252 0.152939
R21533 gnd.n5254 gnd.n5253 0.152939
R21534 gnd.n5254 gnd.n1851 0.152939
R21535 gnd.n5283 gnd.n1851 0.152939
R21536 gnd.n5284 gnd.n5283 0.152939
R21537 gnd.n5285 gnd.n5284 0.152939
R21538 gnd.n5286 gnd.n5285 0.152939
R21539 gnd.n5288 gnd.n5286 0.152939
R21540 gnd.n5288 gnd.n5287 0.152939
R21541 gnd.n5287 gnd.n1843 0.152939
R21542 gnd.n1843 gnd.n1841 0.152939
R21543 gnd.n5323 gnd.n1841 0.152939
R21544 gnd.n5324 gnd.n5323 0.152939
R21545 gnd.n5325 gnd.n5324 0.152939
R21546 gnd.n5326 gnd.n5325 0.152939
R21547 gnd.n5327 gnd.n5326 0.152939
R21548 gnd.n5327 gnd.n1832 0.152939
R21549 gnd.n5376 gnd.n1832 0.152939
R21550 gnd.n5377 gnd.n5376 0.152939
R21551 gnd.n5378 gnd.n5377 0.152939
R21552 gnd.n5380 gnd.n5378 0.152939
R21553 gnd.n5380 gnd.n5379 0.152939
R21554 gnd.n5379 gnd.n1646 0.152939
R21555 gnd.n5698 gnd.n1646 0.152939
R21556 gnd.n5066 gnd.n4874 0.152939
R21557 gnd.n4877 gnd.n4874 0.152939
R21558 gnd.n4878 gnd.n4877 0.152939
R21559 gnd.n4879 gnd.n4878 0.152939
R21560 gnd.n4882 gnd.n4879 0.152939
R21561 gnd.n4883 gnd.n4882 0.152939
R21562 gnd.n4884 gnd.n4883 0.152939
R21563 gnd.n4885 gnd.n4884 0.152939
R21564 gnd.n4888 gnd.n4885 0.152939
R21565 gnd.n4889 gnd.n4888 0.152939
R21566 gnd.n4890 gnd.n4889 0.152939
R21567 gnd.n4891 gnd.n4890 0.152939
R21568 gnd.n4894 gnd.n4891 0.152939
R21569 gnd.n4895 gnd.n4894 0.152939
R21570 gnd.n4896 gnd.n4895 0.152939
R21571 gnd.n4897 gnd.n4896 0.152939
R21572 gnd.n4903 gnd.n4897 0.152939
R21573 gnd.n4904 gnd.n4903 0.152939
R21574 gnd.n4905 gnd.n4904 0.152939
R21575 gnd.n4906 gnd.n4905 0.152939
R21576 gnd.n4909 gnd.n4906 0.152939
R21577 gnd.n4910 gnd.n4909 0.152939
R21578 gnd.n4911 gnd.n4910 0.152939
R21579 gnd.n4912 gnd.n4911 0.152939
R21580 gnd.n4915 gnd.n4912 0.152939
R21581 gnd.n4916 gnd.n4915 0.152939
R21582 gnd.n4917 gnd.n4916 0.152939
R21583 gnd.n4918 gnd.n4917 0.152939
R21584 gnd.n4921 gnd.n4918 0.152939
R21585 gnd.n4922 gnd.n4921 0.152939
R21586 gnd.n4923 gnd.n4922 0.152939
R21587 gnd.n4924 gnd.n4923 0.152939
R21588 gnd.n4927 gnd.n4924 0.152939
R21589 gnd.n4928 gnd.n4927 0.152939
R21590 gnd.n4929 gnd.n4928 0.152939
R21591 gnd.n4994 gnd.n4929 0.152939
R21592 gnd.n4994 gnd.n4993 0.152939
R21593 gnd.n4993 gnd.n4992 0.152939
R21594 gnd.n5067 gnd.n1979 0.152939
R21595 gnd.n5081 gnd.n1979 0.152939
R21596 gnd.n5082 gnd.n5081 0.152939
R21597 gnd.n5083 gnd.n5082 0.152939
R21598 gnd.n5083 gnd.n1963 0.152939
R21599 gnd.n5097 gnd.n1963 0.152939
R21600 gnd.n5098 gnd.n5097 0.152939
R21601 gnd.n5099 gnd.n5098 0.152939
R21602 gnd.n5099 gnd.n1947 0.152939
R21603 gnd.n5113 gnd.n1947 0.152939
R21604 gnd.n5114 gnd.n5113 0.152939
R21605 gnd.n5115 gnd.n5114 0.152939
R21606 gnd.n5115 gnd.n1931 0.152939
R21607 gnd.n5129 gnd.n1931 0.152939
R21608 gnd.n5130 gnd.n5129 0.152939
R21609 gnd.n5131 gnd.n5130 0.152939
R21610 gnd.n5131 gnd.n1914 0.152939
R21611 gnd.n5153 gnd.n1914 0.152939
R21612 gnd.n5154 gnd.n5153 0.152939
R21613 gnd.n5155 gnd.n5154 0.152939
R21614 gnd.n5156 gnd.n5155 0.152939
R21615 gnd.n5156 gnd.n1878 0.152939
R21616 gnd.n5193 gnd.n1878 0.152939
R21617 gnd.n5194 gnd.n5193 0.152939
R21618 gnd.n5195 gnd.n5194 0.152939
R21619 gnd.n5195 gnd.n1764 0.152939
R21620 gnd.n5466 gnd.n1764 0.152939
R21621 gnd.n1802 gnd.n1801 0.152939
R21622 gnd.n3146 gnd.n2186 0.152939
R21623 gnd.n3147 gnd.n3146 0.152939
R21624 gnd.n3148 gnd.n3147 0.152939
R21625 gnd.n3148 gnd.n2180 0.152939
R21626 gnd.n3156 gnd.n2180 0.152939
R21627 gnd.n3157 gnd.n3156 0.152939
R21628 gnd.n3158 gnd.n3157 0.152939
R21629 gnd.n3158 gnd.n2174 0.152939
R21630 gnd.n3166 gnd.n2174 0.152939
R21631 gnd.n3167 gnd.n3166 0.152939
R21632 gnd.n3168 gnd.n3167 0.152939
R21633 gnd.n3168 gnd.n2168 0.152939
R21634 gnd.n3176 gnd.n2168 0.152939
R21635 gnd.n3177 gnd.n3176 0.152939
R21636 gnd.n3178 gnd.n3177 0.152939
R21637 gnd.n3178 gnd.n2162 0.152939
R21638 gnd.n3186 gnd.n2162 0.152939
R21639 gnd.n3187 gnd.n3186 0.152939
R21640 gnd.n3188 gnd.n3187 0.152939
R21641 gnd.n3188 gnd.n2156 0.152939
R21642 gnd.n3196 gnd.n2156 0.152939
R21643 gnd.n3197 gnd.n3196 0.152939
R21644 gnd.n3198 gnd.n3197 0.152939
R21645 gnd.n3198 gnd.n2150 0.152939
R21646 gnd.n3206 gnd.n2150 0.152939
R21647 gnd.n3207 gnd.n3206 0.152939
R21648 gnd.n3208 gnd.n3207 0.152939
R21649 gnd.n3208 gnd.n2144 0.152939
R21650 gnd.n3216 gnd.n2144 0.152939
R21651 gnd.n3217 gnd.n3216 0.152939
R21652 gnd.n3218 gnd.n3217 0.152939
R21653 gnd.n3218 gnd.n2138 0.152939
R21654 gnd.n3226 gnd.n2138 0.152939
R21655 gnd.n3227 gnd.n3226 0.152939
R21656 gnd.n3228 gnd.n3227 0.152939
R21657 gnd.n3228 gnd.n2132 0.152939
R21658 gnd.n3236 gnd.n2132 0.152939
R21659 gnd.n3237 gnd.n3236 0.152939
R21660 gnd.n3238 gnd.n3237 0.152939
R21661 gnd.n3238 gnd.n2126 0.152939
R21662 gnd.n3246 gnd.n2126 0.152939
R21663 gnd.n3247 gnd.n3246 0.152939
R21664 gnd.n3248 gnd.n3247 0.152939
R21665 gnd.n3248 gnd.n2120 0.152939
R21666 gnd.n3256 gnd.n2120 0.152939
R21667 gnd.n3257 gnd.n3256 0.152939
R21668 gnd.n3258 gnd.n3257 0.152939
R21669 gnd.n3258 gnd.n2114 0.152939
R21670 gnd.n3266 gnd.n2114 0.152939
R21671 gnd.n3267 gnd.n3266 0.152939
R21672 gnd.n3268 gnd.n3267 0.152939
R21673 gnd.n3268 gnd.n2108 0.152939
R21674 gnd.n3276 gnd.n2108 0.152939
R21675 gnd.n3277 gnd.n3276 0.152939
R21676 gnd.n3278 gnd.n3277 0.152939
R21677 gnd.n3278 gnd.n2102 0.152939
R21678 gnd.n3286 gnd.n2102 0.152939
R21679 gnd.n3287 gnd.n3286 0.152939
R21680 gnd.n3288 gnd.n3287 0.152939
R21681 gnd.n3288 gnd.n2096 0.152939
R21682 gnd.n3296 gnd.n2096 0.152939
R21683 gnd.n3297 gnd.n3296 0.152939
R21684 gnd.n3298 gnd.n3297 0.152939
R21685 gnd.n3298 gnd.n2090 0.152939
R21686 gnd.n3306 gnd.n2090 0.152939
R21687 gnd.n3307 gnd.n3306 0.152939
R21688 gnd.n3308 gnd.n3307 0.152939
R21689 gnd.n3308 gnd.n2084 0.152939
R21690 gnd.n3316 gnd.n2084 0.152939
R21691 gnd.n3317 gnd.n3316 0.152939
R21692 gnd.n3318 gnd.n3317 0.152939
R21693 gnd.n3318 gnd.n2078 0.152939
R21694 gnd.n3326 gnd.n2078 0.152939
R21695 gnd.n3327 gnd.n3326 0.152939
R21696 gnd.n3328 gnd.n3327 0.152939
R21697 gnd.n3328 gnd.n2072 0.152939
R21698 gnd.n3336 gnd.n2072 0.152939
R21699 gnd.n3337 gnd.n3336 0.152939
R21700 gnd.n3338 gnd.n3337 0.152939
R21701 gnd.n3338 gnd.n2066 0.152939
R21702 gnd.n3346 gnd.n2066 0.152939
R21703 gnd.n3347 gnd.n3346 0.152939
R21704 gnd.n3348 gnd.n3347 0.152939
R21705 gnd.n3350 gnd.n3348 0.152939
R21706 gnd.n6704 gnd.n6703 0.152939
R21707 gnd.n6703 gnd.n6702 0.152939
R21708 gnd.n6702 gnd.n6682 0.152939
R21709 gnd.n6698 gnd.n6682 0.152939
R21710 gnd.n6698 gnd.n6697 0.152939
R21711 gnd.n6697 gnd.n6696 0.152939
R21712 gnd.n6696 gnd.n6688 0.152939
R21713 gnd.n6688 gnd.n634 0.152939
R21714 gnd.n6813 gnd.n634 0.152939
R21715 gnd.n5821 gnd.n5820 0.152939
R21716 gnd.n5822 gnd.n5821 0.152939
R21717 gnd.n5822 gnd.n1292 0.152939
R21718 gnd.n5838 gnd.n1292 0.152939
R21719 gnd.n5839 gnd.n5838 0.152939
R21720 gnd.n5841 gnd.n5839 0.152939
R21721 gnd.n5841 gnd.n5840 0.152939
R21722 gnd.n5840 gnd.n1251 0.152939
R21723 gnd.n5994 gnd.n1251 0.152939
R21724 gnd.n5995 gnd.n5994 0.152939
R21725 gnd.n5996 gnd.n5995 0.152939
R21726 gnd.n5996 gnd.n1236 0.152939
R21727 gnd.n6010 gnd.n1236 0.152939
R21728 gnd.n6011 gnd.n6010 0.152939
R21729 gnd.n6012 gnd.n6011 0.152939
R21730 gnd.n6012 gnd.n1221 0.152939
R21731 gnd.n6026 gnd.n1221 0.152939
R21732 gnd.n6027 gnd.n6026 0.152939
R21733 gnd.n6028 gnd.n6027 0.152939
R21734 gnd.n6028 gnd.n1204 0.152939
R21735 gnd.n6043 gnd.n1204 0.152939
R21736 gnd.n6044 gnd.n6043 0.152939
R21737 gnd.n6046 gnd.n6044 0.152939
R21738 gnd.n6046 gnd.n6045 0.152939
R21739 gnd.n6045 gnd.n1098 0.152939
R21740 gnd.n6136 gnd.n1098 0.152939
R21741 gnd.n6137 gnd.n6136 0.152939
R21742 gnd.n6138 gnd.n6137 0.152939
R21743 gnd.n6138 gnd.n1083 0.152939
R21744 gnd.n6152 gnd.n1083 0.152939
R21745 gnd.n6153 gnd.n6152 0.152939
R21746 gnd.n6154 gnd.n6153 0.152939
R21747 gnd.n6154 gnd.n1069 0.152939
R21748 gnd.n6168 gnd.n1069 0.152939
R21749 gnd.n6169 gnd.n6168 0.152939
R21750 gnd.n6170 gnd.n6169 0.152939
R21751 gnd.n6170 gnd.n1053 0.152939
R21752 gnd.n6186 gnd.n1053 0.152939
R21753 gnd.n6187 gnd.n6186 0.152939
R21754 gnd.n6189 gnd.n6187 0.152939
R21755 gnd.n6189 gnd.n6188 0.152939
R21756 gnd.n6188 gnd.n1011 0.152939
R21757 gnd.n6441 gnd.n1011 0.152939
R21758 gnd.n6442 gnd.n6441 0.152939
R21759 gnd.n6443 gnd.n6442 0.152939
R21760 gnd.n6443 gnd.n995 0.152939
R21761 gnd.n6457 gnd.n995 0.152939
R21762 gnd.n6458 gnd.n6457 0.152939
R21763 gnd.n6459 gnd.n6458 0.152939
R21764 gnd.n6459 gnd.n980 0.152939
R21765 gnd.n6473 gnd.n980 0.152939
R21766 gnd.n6474 gnd.n6473 0.152939
R21767 gnd.n6475 gnd.n6474 0.152939
R21768 gnd.n6475 gnd.n965 0.152939
R21769 gnd.n6489 gnd.n965 0.152939
R21770 gnd.n6490 gnd.n6489 0.152939
R21771 gnd.n6491 gnd.n6490 0.152939
R21772 gnd.n6491 gnd.n950 0.152939
R21773 gnd.n6505 gnd.n950 0.152939
R21774 gnd.n6506 gnd.n6505 0.152939
R21775 gnd.n6507 gnd.n6506 0.152939
R21776 gnd.n6507 gnd.n934 0.152939
R21777 gnd.n6520 gnd.n934 0.152939
R21778 gnd.n6521 gnd.n6520 0.152939
R21779 gnd.n6529 gnd.n6521 0.152939
R21780 gnd.n6529 gnd.n6528 0.152939
R21781 gnd.n6528 gnd.n6527 0.152939
R21782 gnd.n6527 gnd.n6522 0.152939
R21783 gnd.n6522 gnd.n895 0.152939
R21784 gnd.n6587 gnd.n895 0.152939
R21785 gnd.n6587 gnd.n6586 0.152939
R21786 gnd.n6586 gnd.n6585 0.152939
R21787 gnd.n6585 gnd.n896 0.152939
R21788 gnd.n6581 gnd.n896 0.152939
R21789 gnd.n6581 gnd.n6580 0.152939
R21790 gnd.n6580 gnd.n651 0.152939
R21791 gnd.n6792 gnd.n651 0.152939
R21792 gnd.n6793 gnd.n6792 0.152939
R21793 gnd.n6795 gnd.n6793 0.152939
R21794 gnd.n6795 gnd.n6794 0.152939
R21795 gnd.n6794 gnd.n635 0.152939
R21796 gnd.n6812 gnd.n635 0.152939
R21797 gnd.n5785 gnd.n1339 0.152939
R21798 gnd.n5793 gnd.n1339 0.152939
R21799 gnd.n5794 gnd.n5793 0.152939
R21800 gnd.n5795 gnd.n5794 0.152939
R21801 gnd.n5795 gnd.n1335 0.152939
R21802 gnd.n5803 gnd.n1335 0.152939
R21803 gnd.n5804 gnd.n5803 0.152939
R21804 gnd.n5805 gnd.n5804 0.152939
R21805 gnd.n5805 gnd.n1308 0.152939
R21806 gnd.n5236 gnd.n1858 0.152939
R21807 gnd.n5237 gnd.n5236 0.152939
R21808 gnd.n5238 gnd.n5237 0.152939
R21809 gnd.n5238 gnd.n1809 0.152939
R21810 gnd.n5426 gnd.n1809 0.152939
R21811 gnd.n5426 gnd.n5425 0.152939
R21812 gnd.n5425 gnd.n5424 0.152939
R21813 gnd.n5424 gnd.n1810 0.152939
R21814 gnd.n5420 gnd.n1810 0.152939
R21815 gnd.n5420 gnd.n5419 0.152939
R21816 gnd.n5419 gnd.n5418 0.152939
R21817 gnd.n5418 gnd.n1814 0.152939
R21818 gnd.n5414 gnd.n1814 0.152939
R21819 gnd.n5414 gnd.n5413 0.152939
R21820 gnd.n5413 gnd.n5412 0.152939
R21821 gnd.n5412 gnd.n1818 0.152939
R21822 gnd.n5408 gnd.n1818 0.152939
R21823 gnd.n5408 gnd.n5407 0.152939
R21824 gnd.n5407 gnd.n5406 0.152939
R21825 gnd.n5406 gnd.n1822 0.152939
R21826 gnd.n5402 gnd.n1822 0.152939
R21827 gnd.n5402 gnd.n5401 0.152939
R21828 gnd.n5401 gnd.n5400 0.152939
R21829 gnd.n5400 gnd.n1826 0.152939
R21830 gnd.n5396 gnd.n1826 0.152939
R21831 gnd.n5396 gnd.n5395 0.152939
R21832 gnd.n5395 gnd.n5394 0.152939
R21833 gnd.n5394 gnd.n1830 0.152939
R21834 gnd.n5390 gnd.n1830 0.152939
R21835 gnd.n5390 gnd.n5389 0.152939
R21836 gnd.n5389 gnd.n1341 0.152939
R21837 gnd.n5687 gnd.n5675 0.152939
R21838 gnd.n5683 gnd.n5675 0.152939
R21839 gnd.n5683 gnd.n5682 0.152939
R21840 gnd.n5682 gnd.n5681 0.152939
R21841 gnd.n5681 gnd.n1284 0.152939
R21842 gnd.n5847 gnd.n1284 0.152939
R21843 gnd.n5848 gnd.n5847 0.152939
R21844 gnd.n5849 gnd.n5848 0.152939
R21845 gnd.n5849 gnd.n1280 0.152939
R21846 gnd.n5856 gnd.n1280 0.152939
R21847 gnd.n5857 gnd.n5856 0.152939
R21848 gnd.n5964 gnd.n5857 0.152939
R21849 gnd.n5964 gnd.n5963 0.152939
R21850 gnd.n5963 gnd.n5962 0.152939
R21851 gnd.n5962 gnd.n5858 0.152939
R21852 gnd.n5958 gnd.n5858 0.152939
R21853 gnd.n5958 gnd.n5957 0.152939
R21854 gnd.n5957 gnd.n5956 0.152939
R21855 gnd.n5956 gnd.n5862 0.152939
R21856 gnd.n5952 gnd.n5862 0.152939
R21857 gnd.n5952 gnd.n5951 0.152939
R21858 gnd.n5951 gnd.n1196 0.152939
R21859 gnd.n6052 gnd.n1196 0.152939
R21860 gnd.n6053 gnd.n6052 0.152939
R21861 gnd.n6054 gnd.n6053 0.152939
R21862 gnd.n6054 gnd.n1192 0.152939
R21863 gnd.n6059 gnd.n1192 0.152939
R21864 gnd.n6060 gnd.n6059 0.152939
R21865 gnd.n6061 gnd.n6060 0.152939
R21866 gnd.n6061 gnd.n1190 0.152939
R21867 gnd.n6066 gnd.n1190 0.152939
R21868 gnd.n6067 gnd.n6066 0.152939
R21869 gnd.n6068 gnd.n6067 0.152939
R21870 gnd.n6068 gnd.n1188 0.152939
R21871 gnd.n6073 gnd.n1188 0.152939
R21872 gnd.n6074 gnd.n6073 0.152939
R21873 gnd.n6076 gnd.n6074 0.152939
R21874 gnd.n6076 gnd.n6075 0.152939
R21875 gnd.n6075 gnd.n1046 0.152939
R21876 gnd.n6195 gnd.n1046 0.152939
R21877 gnd.n6196 gnd.n6195 0.152939
R21878 gnd.n6197 gnd.n6196 0.152939
R21879 gnd.n6197 gnd.n1042 0.152939
R21880 gnd.n6202 gnd.n1042 0.152939
R21881 gnd.n6203 gnd.n6202 0.152939
R21882 gnd.n6411 gnd.n6203 0.152939
R21883 gnd.n6411 gnd.n6410 0.152939
R21884 gnd.n6410 gnd.n6409 0.152939
R21885 gnd.n6409 gnd.n6204 0.152939
R21886 gnd.n6405 gnd.n6204 0.152939
R21887 gnd.n6405 gnd.n6404 0.152939
R21888 gnd.n6404 gnd.n6403 0.152939
R21889 gnd.n6403 gnd.n6208 0.152939
R21890 gnd.n6399 gnd.n6208 0.152939
R21891 gnd.n6399 gnd.n6398 0.152939
R21892 gnd.n6398 gnd.n6397 0.152939
R21893 gnd.n6397 gnd.n6212 0.152939
R21894 gnd.n6393 gnd.n6212 0.152939
R21895 gnd.n6393 gnd.n6392 0.152939
R21896 gnd.n6392 gnd.n6391 0.152939
R21897 gnd.n6391 gnd.n6216 0.152939
R21898 gnd.n6387 gnd.n6216 0.152939
R21899 gnd.n6387 gnd.n6386 0.152939
R21900 gnd.n6386 gnd.n6385 0.152939
R21901 gnd.n6385 gnd.n6220 0.152939
R21902 gnd.n6220 gnd.n916 0.152939
R21903 gnd.n6545 gnd.n916 0.152939
R21904 gnd.n6546 gnd.n6545 0.152939
R21905 gnd.n6548 gnd.n6546 0.152939
R21906 gnd.n6548 gnd.n6547 0.152939
R21907 gnd.n6547 gnd.n875 0.152939
R21908 gnd.n6603 gnd.n875 0.152939
R21909 gnd.n6604 gnd.n6603 0.152939
R21910 gnd.n6605 gnd.n6604 0.152939
R21911 gnd.n6605 gnd.n872 0.152939
R21912 gnd.n6610 gnd.n872 0.152939
R21913 gnd.n6611 gnd.n6610 0.152939
R21914 gnd.n6765 gnd.n6611 0.152939
R21915 gnd.n6765 gnd.n6764 0.152939
R21916 gnd.n6764 gnd.n6763 0.152939
R21917 gnd.n6763 gnd.n6612 0.152939
R21918 gnd.n6615 gnd.n6612 0.152939
R21919 gnd.n7058 gnd.n477 0.152939
R21920 gnd.n7059 gnd.n7058 0.152939
R21921 gnd.n7060 gnd.n7059 0.152939
R21922 gnd.n7060 gnd.n459 0.152939
R21923 gnd.n7074 gnd.n459 0.152939
R21924 gnd.n7075 gnd.n7074 0.152939
R21925 gnd.n7076 gnd.n7075 0.152939
R21926 gnd.n7076 gnd.n443 0.152939
R21927 gnd.n7090 gnd.n443 0.152939
R21928 gnd.n7091 gnd.n7090 0.152939
R21929 gnd.n7092 gnd.n7091 0.152939
R21930 gnd.n7092 gnd.n425 0.152939
R21931 gnd.n7106 gnd.n425 0.152939
R21932 gnd.n7107 gnd.n7106 0.152939
R21933 gnd.n7108 gnd.n7107 0.152939
R21934 gnd.n7108 gnd.n409 0.152939
R21935 gnd.n7122 gnd.n409 0.152939
R21936 gnd.n7123 gnd.n7122 0.152939
R21937 gnd.n7127 gnd.n7123 0.152939
R21938 gnd.n7127 gnd.n7126 0.152939
R21939 gnd.n7126 gnd.n7125 0.152939
R21940 gnd.n7125 gnd.n377 0.152939
R21941 gnd.n7178 gnd.n377 0.152939
R21942 gnd.n7178 gnd.n7177 0.152939
R21943 gnd.n7177 gnd.n7176 0.152939
R21944 gnd.n7176 gnd.n378 0.152939
R21945 gnd.n7172 gnd.n378 0.152939
R21946 gnd.n7172 gnd.n316 0.152939
R21947 gnd.n7317 gnd.n316 0.152939
R21948 gnd.n7317 gnd.n7316 0.152939
R21949 gnd.n7316 gnd.n7315 0.152939
R21950 gnd.n7315 gnd.n317 0.152939
R21951 gnd.n7311 gnd.n317 0.152939
R21952 gnd.n7311 gnd.n7310 0.152939
R21953 gnd.n7310 gnd.n7309 0.152939
R21954 gnd.n7309 gnd.n322 0.152939
R21955 gnd.n322 gnd.n292 0.152939
R21956 gnd.n7332 gnd.n292 0.152939
R21957 gnd.n7333 gnd.n7332 0.152939
R21958 gnd.n7334 gnd.n7333 0.152939
R21959 gnd.n7334 gnd.n276 0.152939
R21960 gnd.n7348 gnd.n276 0.152939
R21961 gnd.n7349 gnd.n7348 0.152939
R21962 gnd.n7350 gnd.n7349 0.152939
R21963 gnd.n7350 gnd.n262 0.152939
R21964 gnd.n7364 gnd.n262 0.152939
R21965 gnd.n7365 gnd.n7364 0.152939
R21966 gnd.n7366 gnd.n7365 0.152939
R21967 gnd.n7366 gnd.n246 0.152939
R21968 gnd.n7380 gnd.n246 0.152939
R21969 gnd.n7381 gnd.n7380 0.152939
R21970 gnd.n7382 gnd.n7381 0.152939
R21971 gnd.n7382 gnd.n231 0.152939
R21972 gnd.n7396 gnd.n231 0.152939
R21973 gnd.n7397 gnd.n7396 0.152939
R21974 gnd.n7398 gnd.n7397 0.152939
R21975 gnd.n7398 gnd.n216 0.152939
R21976 gnd.n7412 gnd.n216 0.152939
R21977 gnd.n7413 gnd.n7412 0.152939
R21978 gnd.n7482 gnd.n7413 0.152939
R21979 gnd.n7482 gnd.n7481 0.152939
R21980 gnd.n7481 gnd.n7480 0.152939
R21981 gnd.n7480 gnd.n7414 0.152939
R21982 gnd.n7476 gnd.n7414 0.152939
R21983 gnd.n7475 gnd.n7416 0.152939
R21984 gnd.n7471 gnd.n7416 0.152939
R21985 gnd.n7471 gnd.n7470 0.152939
R21986 gnd.n7470 gnd.n7469 0.152939
R21987 gnd.n7469 gnd.n7422 0.152939
R21988 gnd.n7465 gnd.n7422 0.152939
R21989 gnd.n7465 gnd.n7464 0.152939
R21990 gnd.n7464 gnd.n7463 0.152939
R21991 gnd.n7463 gnd.n7430 0.152939
R21992 gnd.n7459 gnd.n7430 0.152939
R21993 gnd.n7459 gnd.n7458 0.152939
R21994 gnd.n7458 gnd.n7457 0.152939
R21995 gnd.n7457 gnd.n7438 0.152939
R21996 gnd.n7453 gnd.n7438 0.152939
R21997 gnd.n7453 gnd.n7452 0.152939
R21998 gnd.n7452 gnd.n7451 0.152939
R21999 gnd.n7451 gnd.n117 0.152939
R22000 gnd.n7577 gnd.n117 0.152939
R22001 gnd.n6971 gnd.n6970 0.152939
R22002 gnd.n6970 gnd.n6969 0.152939
R22003 gnd.n6969 gnd.n567 0.152939
R22004 gnd.n6965 gnd.n567 0.152939
R22005 gnd.n6965 gnd.n6964 0.152939
R22006 gnd.n6964 gnd.n6963 0.152939
R22007 gnd.n6963 gnd.n571 0.152939
R22008 gnd.n6959 gnd.n571 0.152939
R22009 gnd.n6959 gnd.n6958 0.152939
R22010 gnd.n6958 gnd.n6957 0.152939
R22011 gnd.n6957 gnd.n575 0.152939
R22012 gnd.n6953 gnd.n575 0.152939
R22013 gnd.n6953 gnd.n6952 0.152939
R22014 gnd.n6952 gnd.n6951 0.152939
R22015 gnd.n6951 gnd.n579 0.152939
R22016 gnd.n6947 gnd.n579 0.152939
R22017 gnd.n6947 gnd.n6946 0.152939
R22018 gnd.n6946 gnd.n6945 0.152939
R22019 gnd.n6945 gnd.n583 0.152939
R22020 gnd.n6941 gnd.n583 0.152939
R22021 gnd.n6941 gnd.n6940 0.152939
R22022 gnd.n6940 gnd.n383 0.152939
R22023 gnd.n7163 gnd.n383 0.152939
R22024 gnd.n7164 gnd.n7163 0.152939
R22025 gnd.n7166 gnd.n7164 0.152939
R22026 gnd.n7166 gnd.n7165 0.152939
R22027 gnd.n7165 gnd.n354 0.152939
R22028 gnd.n7208 gnd.n354 0.152939
R22029 gnd.n7208 gnd.n7207 0.152939
R22030 gnd.n7207 gnd.n7206 0.152939
R22031 gnd.n7206 gnd.n75 0.152939
R22032 gnd.n7626 gnd.n75 0.152939
R22033 gnd.n7626 gnd.n7625 0.152939
R22034 gnd.n7625 gnd.n77 0.152939
R22035 gnd.n7621 gnd.n77 0.152939
R22036 gnd.n7621 gnd.n7620 0.152939
R22037 gnd.n7620 gnd.n7619 0.152939
R22038 gnd.n7619 gnd.n82 0.152939
R22039 gnd.n7615 gnd.n82 0.152939
R22040 gnd.n7615 gnd.n7614 0.152939
R22041 gnd.n7614 gnd.n7613 0.152939
R22042 gnd.n7613 gnd.n87 0.152939
R22043 gnd.n7609 gnd.n87 0.152939
R22044 gnd.n7609 gnd.n7608 0.152939
R22045 gnd.n7608 gnd.n7607 0.152939
R22046 gnd.n7607 gnd.n92 0.152939
R22047 gnd.n7603 gnd.n92 0.152939
R22048 gnd.n7603 gnd.n7602 0.152939
R22049 gnd.n7602 gnd.n7601 0.152939
R22050 gnd.n7601 gnd.n97 0.152939
R22051 gnd.n7597 gnd.n97 0.152939
R22052 gnd.n7597 gnd.n7596 0.152939
R22053 gnd.n7596 gnd.n7595 0.152939
R22054 gnd.n7595 gnd.n102 0.152939
R22055 gnd.n7591 gnd.n102 0.152939
R22056 gnd.n7591 gnd.n7590 0.152939
R22057 gnd.n7590 gnd.n7589 0.152939
R22058 gnd.n7589 gnd.n107 0.152939
R22059 gnd.n7585 gnd.n107 0.152939
R22060 gnd.n7585 gnd.n7584 0.152939
R22061 gnd.n7584 gnd.n7583 0.152939
R22062 gnd.n7583 gnd.n112 0.152939
R22063 gnd.n7579 gnd.n112 0.152939
R22064 gnd.n7579 gnd.n7578 0.152939
R22065 gnd.n6704 gnd.n566 0.151415
R22066 gnd.n5785 gnd.n5784 0.151415
R22067 gnd.n5209 gnd.n5207 0.145814
R22068 gnd.n5209 gnd.n1858 0.145814
R22069 gnd.n347 gnd.n300 0.130073
R22070 gnd.n1801 gnd.n1765 0.130073
R22071 gnd.n4189 gnd.n3535 0.0767195
R22072 gnd.n4189 gnd.n4188 0.0767195
R22073 gnd.n5689 gnd.n5688 0.063
R22074 gnd.n6620 gnd.n6619 0.063
R22075 gnd.n4719 gnd.n2029 0.0477147
R22076 gnd.n3979 gnd.n3867 0.0442063
R22077 gnd.n3980 gnd.n3979 0.0442063
R22078 gnd.n3981 gnd.n3980 0.0442063
R22079 gnd.n3981 gnd.n3856 0.0442063
R22080 gnd.n3995 gnd.n3856 0.0442063
R22081 gnd.n3996 gnd.n3995 0.0442063
R22082 gnd.n3997 gnd.n3996 0.0442063
R22083 gnd.n3997 gnd.n3843 0.0442063
R22084 gnd.n4041 gnd.n3843 0.0442063
R22085 gnd.n4042 gnd.n4041 0.0442063
R22086 gnd.n4044 gnd.n3777 0.0344674
R22087 gnd.n6708 gnd.n6676 0.0344674
R22088 gnd.n5783 gnd.n5782 0.0344674
R22089 gnd.n4064 gnd.n4063 0.0269946
R22090 gnd.n4066 gnd.n4065 0.0269946
R22091 gnd.n3772 gnd.n3770 0.0269946
R22092 gnd.n4076 gnd.n4074 0.0269946
R22093 gnd.n4075 gnd.n3751 0.0269946
R22094 gnd.n4095 gnd.n4094 0.0269946
R22095 gnd.n4097 gnd.n4096 0.0269946
R22096 gnd.n3746 gnd.n3745 0.0269946
R22097 gnd.n4107 gnd.n3741 0.0269946
R22098 gnd.n4106 gnd.n3743 0.0269946
R22099 gnd.n3742 gnd.n3722 0.0269946
R22100 gnd.n4133 gnd.n3723 0.0269946
R22101 gnd.n4132 gnd.n3724 0.0269946
R22102 gnd.n4152 gnd.n3708 0.0269946
R22103 gnd.n4154 gnd.n4153 0.0269946
R22104 gnd.n4155 gnd.n3688 0.0269946
R22105 gnd.n4156 gnd.n3689 0.0269946
R22106 gnd.n4157 gnd.n3690 0.0269946
R22107 gnd.n3692 gnd.n3691 0.0269946
R22108 gnd.n3529 gnd.n3527 0.0269946
R22109 gnd.n4201 gnd.n4199 0.0269946
R22110 gnd.n4200 gnd.n3511 0.0269946
R22111 gnd.n4220 gnd.n4219 0.0269946
R22112 gnd.n4222 gnd.n4221 0.0269946
R22113 gnd.n3506 gnd.n3504 0.0269946
R22114 gnd.n4232 gnd.n4230 0.0269946
R22115 gnd.n4231 gnd.n3486 0.0269946
R22116 gnd.n4251 gnd.n4250 0.0269946
R22117 gnd.n4253 gnd.n4252 0.0269946
R22118 gnd.n3480 gnd.n3478 0.0269946
R22119 gnd.n4263 gnd.n4261 0.0269946
R22120 gnd.n4262 gnd.n3459 0.0269946
R22121 gnd.n4282 gnd.n4281 0.0269946
R22122 gnd.n4284 gnd.n4283 0.0269946
R22123 gnd.n3454 gnd.n3452 0.0269946
R22124 gnd.n4294 gnd.n4292 0.0269946
R22125 gnd.n4293 gnd.n3435 0.0269946
R22126 gnd.n4313 gnd.n4312 0.0269946
R22127 gnd.n4315 gnd.n4314 0.0269946
R22128 gnd.n3430 gnd.n3428 0.0269946
R22129 gnd.n4325 gnd.n4323 0.0269946
R22130 gnd.n4324 gnd.n3409 0.0269946
R22131 gnd.n4344 gnd.n4343 0.0269946
R22132 gnd.n4346 gnd.n4345 0.0269946
R22133 gnd.n3404 gnd.n3402 0.0269946
R22134 gnd.n4356 gnd.n4354 0.0269946
R22135 gnd.n4355 gnd.n3384 0.0269946
R22136 gnd.n4375 gnd.n4374 0.0269946
R22137 gnd.n3378 gnd.n3376 0.0269946
R22138 gnd.n4643 gnd.n4641 0.0269946
R22139 gnd.n4642 gnd.n3358 0.0269946
R22140 gnd.n4661 gnd.n4660 0.0269946
R22141 gnd.n6619 gnd.n6617 0.0246168
R22142 gnd.n5688 gnd.n5674 0.0246168
R22143 gnd.n7217 gnd.n300 0.0233659
R22144 gnd.n3349 gnd.n1765 0.0233659
R22145 gnd.n4044 gnd.n4043 0.0202011
R22146 gnd.n6756 gnd.n6617 0.0174837
R22147 gnd.n6756 gnd.n6755 0.0174837
R22148 gnd.n6755 gnd.n6618 0.0174837
R22149 gnd.n6752 gnd.n6618 0.0174837
R22150 gnd.n6752 gnd.n6751 0.0174837
R22151 gnd.n6751 gnd.n6629 0.0174837
R22152 gnd.n6748 gnd.n6629 0.0174837
R22153 gnd.n6748 gnd.n6747 0.0174837
R22154 gnd.n6747 gnd.n6635 0.0174837
R22155 gnd.n6744 gnd.n6635 0.0174837
R22156 gnd.n6744 gnd.n6743 0.0174837
R22157 gnd.n6743 gnd.n6639 0.0174837
R22158 gnd.n6740 gnd.n6639 0.0174837
R22159 gnd.n6740 gnd.n6739 0.0174837
R22160 gnd.n6739 gnd.n6643 0.0174837
R22161 gnd.n6736 gnd.n6643 0.0174837
R22162 gnd.n6736 gnd.n6735 0.0174837
R22163 gnd.n6735 gnd.n6649 0.0174837
R22164 gnd.n6732 gnd.n6649 0.0174837
R22165 gnd.n6732 gnd.n6731 0.0174837
R22166 gnd.n6731 gnd.n6655 0.0174837
R22167 gnd.n6728 gnd.n6655 0.0174837
R22168 gnd.n6728 gnd.n6727 0.0174837
R22169 gnd.n6727 gnd.n6659 0.0174837
R22170 gnd.n6724 gnd.n6659 0.0174837
R22171 gnd.n6724 gnd.n6723 0.0174837
R22172 gnd.n6723 gnd.n6663 0.0174837
R22173 gnd.n6720 gnd.n6663 0.0174837
R22174 gnd.n6720 gnd.n6719 0.0174837
R22175 gnd.n6719 gnd.n6669 0.0174837
R22176 gnd.n6716 gnd.n6669 0.0174837
R22177 gnd.n6716 gnd.n6715 0.0174837
R22178 gnd.n6715 gnd.n6675 0.0174837
R22179 gnd.n6709 gnd.n6675 0.0174837
R22180 gnd.n6709 gnd.n6708 0.0174837
R22181 gnd.n5674 gnd.n5574 0.0174837
R22182 gnd.n5671 gnd.n5574 0.0174837
R22183 gnd.n5671 gnd.n5670 0.0174837
R22184 gnd.n5670 gnd.n5580 0.0174837
R22185 gnd.n5667 gnd.n5580 0.0174837
R22186 gnd.n5667 gnd.n5666 0.0174837
R22187 gnd.n5666 gnd.n5586 0.0174837
R22188 gnd.n5663 gnd.n5586 0.0174837
R22189 gnd.n5663 gnd.n5662 0.0174837
R22190 gnd.n5662 gnd.n5592 0.0174837
R22191 gnd.n5659 gnd.n5592 0.0174837
R22192 gnd.n5659 gnd.n5658 0.0174837
R22193 gnd.n5658 gnd.n5598 0.0174837
R22194 gnd.n5655 gnd.n5598 0.0174837
R22195 gnd.n5655 gnd.n5654 0.0174837
R22196 gnd.n5654 gnd.n5605 0.0174837
R22197 gnd.n5651 gnd.n5605 0.0174837
R22198 gnd.n5651 gnd.n5650 0.0174837
R22199 gnd.n5650 gnd.n5609 0.0174837
R22200 gnd.n5647 gnd.n5609 0.0174837
R22201 gnd.n5647 gnd.n5646 0.0174837
R22202 gnd.n5646 gnd.n5615 0.0174837
R22203 gnd.n5643 gnd.n5615 0.0174837
R22204 gnd.n5643 gnd.n5642 0.0174837
R22205 gnd.n5642 gnd.n5621 0.0174837
R22206 gnd.n5639 gnd.n5621 0.0174837
R22207 gnd.n5639 gnd.n5638 0.0174837
R22208 gnd.n5638 gnd.n5631 0.0174837
R22209 gnd.n5635 gnd.n5631 0.0174837
R22210 gnd.n5635 gnd.n5634 0.0174837
R22211 gnd.n5634 gnd.n1346 0.0174837
R22212 gnd.n5776 gnd.n1346 0.0174837
R22213 gnd.n5777 gnd.n5776 0.0174837
R22214 gnd.n5777 gnd.n1342 0.0174837
R22215 gnd.n5782 gnd.n1342 0.0174837
R22216 gnd.n4043 gnd.n4042 0.0148637
R22217 gnd.n4632 gnd.n4376 0.0144266
R22218 gnd.n4633 gnd.n4632 0.0130679
R22219 gnd.n4063 gnd.n3777 0.00797283
R22220 gnd.n4065 gnd.n4064 0.00797283
R22221 gnd.n4066 gnd.n3772 0.00797283
R22222 gnd.n4074 gnd.n3770 0.00797283
R22223 gnd.n4076 gnd.n4075 0.00797283
R22224 gnd.n4094 gnd.n3751 0.00797283
R22225 gnd.n4096 gnd.n4095 0.00797283
R22226 gnd.n4097 gnd.n3746 0.00797283
R22227 gnd.n3745 gnd.n3741 0.00797283
R22228 gnd.n4107 gnd.n4106 0.00797283
R22229 gnd.n3743 gnd.n3742 0.00797283
R22230 gnd.n3723 gnd.n3722 0.00797283
R22231 gnd.n4133 gnd.n4132 0.00797283
R22232 gnd.n3724 gnd.n3708 0.00797283
R22233 gnd.n4153 gnd.n4152 0.00797283
R22234 gnd.n4155 gnd.n4154 0.00797283
R22235 gnd.n4156 gnd.n3688 0.00797283
R22236 gnd.n4157 gnd.n3689 0.00797283
R22237 gnd.n3691 gnd.n3690 0.00797283
R22238 gnd.n3692 gnd.n3529 0.00797283
R22239 gnd.n4199 gnd.n3527 0.00797283
R22240 gnd.n4201 gnd.n4200 0.00797283
R22241 gnd.n4219 gnd.n3511 0.00797283
R22242 gnd.n4221 gnd.n4220 0.00797283
R22243 gnd.n4222 gnd.n3506 0.00797283
R22244 gnd.n4230 gnd.n3504 0.00797283
R22245 gnd.n4232 gnd.n4231 0.00797283
R22246 gnd.n4250 gnd.n3486 0.00797283
R22247 gnd.n4252 gnd.n4251 0.00797283
R22248 gnd.n4253 gnd.n3480 0.00797283
R22249 gnd.n4261 gnd.n3478 0.00797283
R22250 gnd.n4263 gnd.n4262 0.00797283
R22251 gnd.n4281 gnd.n3459 0.00797283
R22252 gnd.n4283 gnd.n4282 0.00797283
R22253 gnd.n4284 gnd.n3454 0.00797283
R22254 gnd.n4292 gnd.n3452 0.00797283
R22255 gnd.n4294 gnd.n4293 0.00797283
R22256 gnd.n4312 gnd.n3435 0.00797283
R22257 gnd.n4314 gnd.n4313 0.00797283
R22258 gnd.n4315 gnd.n3430 0.00797283
R22259 gnd.n4323 gnd.n3428 0.00797283
R22260 gnd.n4325 gnd.n4324 0.00797283
R22261 gnd.n4343 gnd.n3409 0.00797283
R22262 gnd.n4345 gnd.n4344 0.00797283
R22263 gnd.n4346 gnd.n3404 0.00797283
R22264 gnd.n4354 gnd.n3402 0.00797283
R22265 gnd.n4356 gnd.n4355 0.00797283
R22266 gnd.n4374 gnd.n3384 0.00797283
R22267 gnd.n4376 gnd.n4375 0.00797283
R22268 gnd.n4633 gnd.n3378 0.00797283
R22269 gnd.n4641 gnd.n3376 0.00797283
R22270 gnd.n4643 gnd.n4642 0.00797283
R22271 gnd.n4660 gnd.n3358 0.00797283
R22272 gnd.n4661 gnd.n2029 0.00797283
R22273 gnd.n333 gnd.n317 0.00433921
R22274 gnd.n5228 gnd.n1861 0.00433921
R22275 gnd.n6676 gnd.n566 0.000839674
R22276 gnd.n5784 gnd.n5783 0.000839674
R22277 plus.n76 plus.t11 250.337
R22278 plus.n15 plus.t14 250.337
R22279 plus.n124 plus.t1 243.97
R22280 plus.n120 plus.t24 231.093
R22281 plus.n59 plus.t20 231.093
R22282 plus.n124 plus.n123 223.454
R22283 plus.n126 plus.n125 223.454
R22284 plus.n77 plus.t5 187.445
R22285 plus.n74 plus.t22 187.445
R22286 plus.n72 plus.t21 187.445
R22287 plus.n89 plus.t16 187.445
R22288 plus.n95 plus.t17 187.445
R22289 plus.n68 plus.t13 187.445
R22290 plus.n66 plus.t15 187.445
R22291 plus.n107 plus.t10 187.445
R22292 plus.n113 plus.t26 187.445
R22293 plus.n62 plus.t28 187.445
R22294 plus.n1 plus.t23 187.445
R22295 plus.n52 plus.t6 187.445
R22296 plus.n46 plus.t12 187.445
R22297 plus.n5 plus.t8 187.445
R22298 plus.n7 plus.t7 187.445
R22299 plus.n34 plus.t19 187.445
R22300 plus.n28 plus.t18 187.445
R22301 plus.n11 plus.t27 187.445
R22302 plus.n13 plus.t25 187.445
R22303 plus.n16 plus.t9 187.445
R22304 plus.n121 plus.n120 161.3
R22305 plus.n119 plus.n61 161.3
R22306 plus.n118 plus.n117 161.3
R22307 plus.n116 plus.n115 161.3
R22308 plus.n114 plus.n63 161.3
R22309 plus.n112 plus.n111 161.3
R22310 plus.n110 plus.n64 161.3
R22311 plus.n109 plus.n108 161.3
R22312 plus.n106 plus.n65 161.3
R22313 plus.n105 plus.n104 161.3
R22314 plus.n103 plus.n102 161.3
R22315 plus.n101 plus.n67 161.3
R22316 plus.n100 plus.n99 161.3
R22317 plus.n98 plus.n97 161.3
R22318 plus.n96 plus.n69 161.3
R22319 plus.n94 plus.n93 161.3
R22320 plus.n92 plus.n70 161.3
R22321 plus.n91 plus.n90 161.3
R22322 plus.n88 plus.n71 161.3
R22323 plus.n87 plus.n86 161.3
R22324 plus.n85 plus.n84 161.3
R22325 plus.n83 plus.n73 161.3
R22326 plus.n82 plus.n81 161.3
R22327 plus.n80 plus.n79 161.3
R22328 plus.n78 plus.n75 161.3
R22329 plus.n17 plus.n14 161.3
R22330 plus.n19 plus.n18 161.3
R22331 plus.n21 plus.n20 161.3
R22332 plus.n22 plus.n12 161.3
R22333 plus.n24 plus.n23 161.3
R22334 plus.n26 plus.n25 161.3
R22335 plus.n27 plus.n10 161.3
R22336 plus.n30 plus.n29 161.3
R22337 plus.n31 plus.n9 161.3
R22338 plus.n33 plus.n32 161.3
R22339 plus.n35 plus.n8 161.3
R22340 plus.n37 plus.n36 161.3
R22341 plus.n39 plus.n38 161.3
R22342 plus.n40 plus.n6 161.3
R22343 plus.n42 plus.n41 161.3
R22344 plus.n44 plus.n43 161.3
R22345 plus.n45 plus.n4 161.3
R22346 plus.n48 plus.n47 161.3
R22347 plus.n49 plus.n3 161.3
R22348 plus.n51 plus.n50 161.3
R22349 plus.n53 plus.n2 161.3
R22350 plus.n55 plus.n54 161.3
R22351 plus.n57 plus.n56 161.3
R22352 plus.n58 plus.n0 161.3
R22353 plus.n60 plus.n59 161.3
R22354 plus.n88 plus.n87 56.5617
R22355 plus.n97 plus.n96 56.5617
R22356 plus.n106 plus.n105 56.5617
R22357 plus.n45 plus.n44 56.5617
R22358 plus.n36 plus.n35 56.5617
R22359 plus.n27 plus.n26 56.5617
R22360 plus.n79 plus.n78 56.5617
R22361 plus.n115 plus.n114 56.5617
R22362 plus.n54 plus.n53 56.5617
R22363 plus.n18 plus.n17 56.5617
R22364 plus.n119 plus.n118 50.2647
R22365 plus.n58 plus.n57 50.2647
R22366 plus.n84 plus.n83 46.3896
R22367 plus.n108 plus.n64 46.3896
R22368 plus.n47 plus.n3 46.3896
R22369 plus.n23 plus.n22 46.3896
R22370 plus.n76 plus.n75 43.1929
R22371 plus.n15 plus.n14 43.1929
R22372 plus.n94 plus.n70 42.5146
R22373 plus.n101 plus.n100 42.5146
R22374 plus.n40 plus.n39 42.5146
R22375 plus.n33 plus.n9 42.5146
R22376 plus.n77 plus.n76 40.6041
R22377 plus.n16 plus.n15 40.6041
R22378 plus.n90 plus.n70 38.6395
R22379 plus.n102 plus.n101 38.6395
R22380 plus.n41 plus.n40 38.6395
R22381 plus.n29 plus.n9 38.6395
R22382 plus.n122 plus.n121 35.2031
R22383 plus.n83 plus.n82 34.7644
R22384 plus.n112 plus.n64 34.7644
R22385 plus.n51 plus.n3 34.7644
R22386 plus.n22 plus.n21 34.7644
R22387 plus.n79 plus.n74 21.8872
R22388 plus.n114 plus.n113 21.8872
R22389 plus.n53 plus.n52 21.8872
R22390 plus.n18 plus.n13 21.8872
R22391 plus.n89 plus.n88 19.9199
R22392 plus.n105 plus.n66 19.9199
R22393 plus.n44 plus.n5 19.9199
R22394 plus.n28 plus.n27 19.9199
R22395 plus.n123 plus.t2 19.8005
R22396 plus.n123 plus.t4 19.8005
R22397 plus.n125 plus.t3 19.8005
R22398 plus.n125 plus.t0 19.8005
R22399 plus.n96 plus.n95 17.9525
R22400 plus.n97 plus.n68 17.9525
R22401 plus.n36 plus.n7 17.9525
R22402 plus.n35 plus.n34 17.9525
R22403 plus.n87 plus.n72 15.9852
R22404 plus.n107 plus.n106 15.9852
R22405 plus.n46 plus.n45 15.9852
R22406 plus.n26 plus.n11 15.9852
R22407 plus plus.n127 15.0684
R22408 plus.n78 plus.n77 14.0178
R22409 plus.n115 plus.n62 14.0178
R22410 plus.n54 plus.n1 14.0178
R22411 plus.n17 plus.n16 14.0178
R22412 plus.n122 plus.n60 11.9342
R22413 plus.n118 plus.n62 10.575
R22414 plus.n57 plus.n1 10.575
R22415 plus.n120 plus.n119 9.49444
R22416 plus.n59 plus.n58 9.49444
R22417 plus.n84 plus.n72 8.60764
R22418 plus.n108 plus.n107 8.60764
R22419 plus.n47 plus.n46 8.60764
R22420 plus.n23 plus.n11 8.60764
R22421 plus.n95 plus.n94 6.6403
R22422 plus.n100 plus.n68 6.6403
R22423 plus.n39 plus.n7 6.6403
R22424 plus.n34 plus.n33 6.6403
R22425 plus.n127 plus.n126 5.40567
R22426 plus.n90 plus.n89 4.67295
R22427 plus.n102 plus.n66 4.67295
R22428 plus.n41 plus.n5 4.67295
R22429 plus.n29 plus.n28 4.67295
R22430 plus.n82 plus.n74 2.7056
R22431 plus.n113 plus.n112 2.7056
R22432 plus.n52 plus.n51 2.7056
R22433 plus.n21 plus.n13 2.7056
R22434 plus.n127 plus.n122 1.188
R22435 plus.n126 plus.n124 0.716017
R22436 plus.n80 plus.n75 0.189894
R22437 plus.n81 plus.n80 0.189894
R22438 plus.n81 plus.n73 0.189894
R22439 plus.n85 plus.n73 0.189894
R22440 plus.n86 plus.n85 0.189894
R22441 plus.n86 plus.n71 0.189894
R22442 plus.n91 plus.n71 0.189894
R22443 plus.n92 plus.n91 0.189894
R22444 plus.n93 plus.n92 0.189894
R22445 plus.n93 plus.n69 0.189894
R22446 plus.n98 plus.n69 0.189894
R22447 plus.n99 plus.n98 0.189894
R22448 plus.n99 plus.n67 0.189894
R22449 plus.n103 plus.n67 0.189894
R22450 plus.n104 plus.n103 0.189894
R22451 plus.n104 plus.n65 0.189894
R22452 plus.n109 plus.n65 0.189894
R22453 plus.n110 plus.n109 0.189894
R22454 plus.n111 plus.n110 0.189894
R22455 plus.n111 plus.n63 0.189894
R22456 plus.n116 plus.n63 0.189894
R22457 plus.n117 plus.n116 0.189894
R22458 plus.n117 plus.n61 0.189894
R22459 plus.n121 plus.n61 0.189894
R22460 plus.n60 plus.n0 0.189894
R22461 plus.n56 plus.n0 0.189894
R22462 plus.n56 plus.n55 0.189894
R22463 plus.n55 plus.n2 0.189894
R22464 plus.n50 plus.n2 0.189894
R22465 plus.n50 plus.n49 0.189894
R22466 plus.n49 plus.n48 0.189894
R22467 plus.n48 plus.n4 0.189894
R22468 plus.n43 plus.n4 0.189894
R22469 plus.n43 plus.n42 0.189894
R22470 plus.n42 plus.n6 0.189894
R22471 plus.n38 plus.n6 0.189894
R22472 plus.n38 plus.n37 0.189894
R22473 plus.n37 plus.n8 0.189894
R22474 plus.n32 plus.n8 0.189894
R22475 plus.n32 plus.n31 0.189894
R22476 plus.n31 plus.n30 0.189894
R22477 plus.n30 plus.n10 0.189894
R22478 plus.n25 plus.n10 0.189894
R22479 plus.n25 plus.n24 0.189894
R22480 plus.n24 plus.n12 0.189894
R22481 plus.n20 plus.n12 0.189894
R22482 plus.n20 plus.n19 0.189894
R22483 plus.n19 plus.n14 0.189894
R22484 a_n3106_n452.n1 a_n3106_n452.t2 214.321
R22485 a_n3106_n452.n14 a_n3106_n452.t37 214.321
R22486 a_n3106_n452.n15 a_n3106_n452.t30 214.321
R22487 a_n3106_n452.n16 a_n3106_n452.t45 214.321
R22488 a_n3106_n452.n17 a_n3106_n452.t3 214.321
R22489 a_n3106_n452.n18 a_n3106_n452.t35 214.321
R22490 a_n3106_n452.n19 a_n3106_n452.t53 214.321
R22491 a_n3106_n452.n20 a_n3106_n452.t38 214.321
R22492 a_n3106_n452.n0 a_n3106_n452.t23 55.8337
R22493 a_n3106_n452.n2 a_n3106_n452.t55 55.8337
R22494 a_n3106_n452.n13 a_n3106_n452.t39 55.8337
R22495 a_n3106_n452.n47 a_n3106_n452.t10 55.8335
R22496 a_n3106_n452.n45 a_n3106_n452.t46 55.8335
R22497 a_n3106_n452.n34 a_n3106_n452.t44 55.8335
R22498 a_n3106_n452.n33 a_n3106_n452.t20 55.8335
R22499 a_n3106_n452.n22 a_n3106_n452.t14 55.8335
R22500 a_n3106_n452.n49 a_n3106_n452.n48 53.0052
R22501 a_n3106_n452.n51 a_n3106_n452.n50 53.0052
R22502 a_n3106_n452.n53 a_n3106_n452.n52 53.0052
R22503 a_n3106_n452.n55 a_n3106_n452.n54 53.0052
R22504 a_n3106_n452.n4 a_n3106_n452.n3 53.0052
R22505 a_n3106_n452.n6 a_n3106_n452.n5 53.0052
R22506 a_n3106_n452.n8 a_n3106_n452.n7 53.0052
R22507 a_n3106_n452.n10 a_n3106_n452.n9 53.0052
R22508 a_n3106_n452.n12 a_n3106_n452.n11 53.0052
R22509 a_n3106_n452.n44 a_n3106_n452.n43 53.0051
R22510 a_n3106_n452.n42 a_n3106_n452.n41 53.0051
R22511 a_n3106_n452.n40 a_n3106_n452.n39 53.0051
R22512 a_n3106_n452.n38 a_n3106_n452.n37 53.0051
R22513 a_n3106_n452.n36 a_n3106_n452.n35 53.0051
R22514 a_n3106_n452.n32 a_n3106_n452.n31 53.0051
R22515 a_n3106_n452.n30 a_n3106_n452.n29 53.0051
R22516 a_n3106_n452.n28 a_n3106_n452.n27 53.0051
R22517 a_n3106_n452.n26 a_n3106_n452.n25 53.0051
R22518 a_n3106_n452.n24 a_n3106_n452.n23 53.0051
R22519 a_n3106_n452.n57 a_n3106_n452.n56 53.0051
R22520 a_n3106_n452.n21 a_n3106_n452.n13 12.2417
R22521 a_n3106_n452.n47 a_n3106_n452.n46 12.2417
R22522 a_n3106_n452.n22 a_n3106_n452.n21 5.16214
R22523 a_n3106_n452.n46 a_n3106_n452.n45 5.16214
R22524 a_n3106_n452.n48 a_n3106_n452.t8 2.82907
R22525 a_n3106_n452.n48 a_n3106_n452.t6 2.82907
R22526 a_n3106_n452.n50 a_n3106_n452.t19 2.82907
R22527 a_n3106_n452.n50 a_n3106_n452.t24 2.82907
R22528 a_n3106_n452.n52 a_n3106_n452.t17 2.82907
R22529 a_n3106_n452.n52 a_n3106_n452.t21 2.82907
R22530 a_n3106_n452.n54 a_n3106_n452.t13 2.82907
R22531 a_n3106_n452.n54 a_n3106_n452.t18 2.82907
R22532 a_n3106_n452.n3 a_n3106_n452.t48 2.82907
R22533 a_n3106_n452.n3 a_n3106_n452.t5 2.82907
R22534 a_n3106_n452.n5 a_n3106_n452.t40 2.82907
R22535 a_n3106_n452.n5 a_n3106_n452.t47 2.82907
R22536 a_n3106_n452.n7 a_n3106_n452.t34 2.82907
R22537 a_n3106_n452.n7 a_n3106_n452.t43 2.82907
R22538 a_n3106_n452.n9 a_n3106_n452.t4 2.82907
R22539 a_n3106_n452.n9 a_n3106_n452.t0 2.82907
R22540 a_n3106_n452.n11 a_n3106_n452.t51 2.82907
R22541 a_n3106_n452.n11 a_n3106_n452.t36 2.82907
R22542 a_n3106_n452.n43 a_n3106_n452.t52 2.82907
R22543 a_n3106_n452.n43 a_n3106_n452.t50 2.82907
R22544 a_n3106_n452.n41 a_n3106_n452.t32 2.82907
R22545 a_n3106_n452.n41 a_n3106_n452.t33 2.82907
R22546 a_n3106_n452.n39 a_n3106_n452.t1 2.82907
R22547 a_n3106_n452.n39 a_n3106_n452.t31 2.82907
R22548 a_n3106_n452.n37 a_n3106_n452.t41 2.82907
R22549 a_n3106_n452.n37 a_n3106_n452.t54 2.82907
R22550 a_n3106_n452.n35 a_n3106_n452.t49 2.82907
R22551 a_n3106_n452.n35 a_n3106_n452.t42 2.82907
R22552 a_n3106_n452.n31 a_n3106_n452.t9 2.82907
R22553 a_n3106_n452.n31 a_n3106_n452.t25 2.82907
R22554 a_n3106_n452.n29 a_n3106_n452.t16 2.82907
R22555 a_n3106_n452.n29 a_n3106_n452.t7 2.82907
R22556 a_n3106_n452.n27 a_n3106_n452.t27 2.82907
R22557 a_n3106_n452.n27 a_n3106_n452.t15 2.82907
R22558 a_n3106_n452.n25 a_n3106_n452.t22 2.82907
R22559 a_n3106_n452.n25 a_n3106_n452.t26 2.82907
R22560 a_n3106_n452.n23 a_n3106_n452.t11 2.82907
R22561 a_n3106_n452.n23 a_n3106_n452.t28 2.82907
R22562 a_n3106_n452.t29 a_n3106_n452.n57 2.82907
R22563 a_n3106_n452.n57 a_n3106_n452.t12 2.82907
R22564 a_n3106_n452.n46 a_n3106_n452.n1 2.54197
R22565 a_n3106_n452.n21 a_n3106_n452.n20 2.0129
R22566 a_n3106_n452.n20 a_n3106_n452.n19 0.672012
R22567 a_n3106_n452.n19 a_n3106_n452.n18 0.672012
R22568 a_n3106_n452.n18 a_n3106_n452.n17 0.672012
R22569 a_n3106_n452.n17 a_n3106_n452.n16 0.672012
R22570 a_n3106_n452.n16 a_n3106_n452.n15 0.672012
R22571 a_n3106_n452.n15 a_n3106_n452.n14 0.672012
R22572 a_n3106_n452.n14 a_n3106_n452.n1 0.672012
R22573 a_n3106_n452.n24 a_n3106_n452.n22 0.530672
R22574 a_n3106_n452.n26 a_n3106_n452.n24 0.530672
R22575 a_n3106_n452.n28 a_n3106_n452.n26 0.530672
R22576 a_n3106_n452.n30 a_n3106_n452.n28 0.530672
R22577 a_n3106_n452.n32 a_n3106_n452.n30 0.530672
R22578 a_n3106_n452.n33 a_n3106_n452.n32 0.530672
R22579 a_n3106_n452.n36 a_n3106_n452.n34 0.530672
R22580 a_n3106_n452.n38 a_n3106_n452.n36 0.530672
R22581 a_n3106_n452.n40 a_n3106_n452.n38 0.530672
R22582 a_n3106_n452.n42 a_n3106_n452.n40 0.530672
R22583 a_n3106_n452.n44 a_n3106_n452.n42 0.530672
R22584 a_n3106_n452.n45 a_n3106_n452.n44 0.530672
R22585 a_n3106_n452.n13 a_n3106_n452.n12 0.530672
R22586 a_n3106_n452.n12 a_n3106_n452.n10 0.530672
R22587 a_n3106_n452.n10 a_n3106_n452.n8 0.530672
R22588 a_n3106_n452.n8 a_n3106_n452.n6 0.530672
R22589 a_n3106_n452.n6 a_n3106_n452.n4 0.530672
R22590 a_n3106_n452.n4 a_n3106_n452.n2 0.530672
R22591 a_n3106_n452.n56 a_n3106_n452.n0 0.530672
R22592 a_n3106_n452.n56 a_n3106_n452.n55 0.530672
R22593 a_n3106_n452.n55 a_n3106_n452.n53 0.530672
R22594 a_n3106_n452.n53 a_n3106_n452.n51 0.530672
R22595 a_n3106_n452.n51 a_n3106_n452.n49 0.530672
R22596 a_n3106_n452.n49 a_n3106_n452.n47 0.530672
R22597 a_n3106_n452.n34 a_n3106_n452.n33 0.235414
R22598 a_n3106_n452.n2 a_n3106_n452.n0 0.235414
R22599 outputibias.n27 outputibias.n1 289.615
R22600 outputibias.n58 outputibias.n32 289.615
R22601 outputibias.n90 outputibias.n64 289.615
R22602 outputibias.n122 outputibias.n96 289.615
R22603 outputibias.n28 outputibias.n27 185
R22604 outputibias.n26 outputibias.n25 185
R22605 outputibias.n5 outputibias.n4 185
R22606 outputibias.n20 outputibias.n19 185
R22607 outputibias.n18 outputibias.n17 185
R22608 outputibias.n9 outputibias.n8 185
R22609 outputibias.n12 outputibias.n11 185
R22610 outputibias.n59 outputibias.n58 185
R22611 outputibias.n57 outputibias.n56 185
R22612 outputibias.n36 outputibias.n35 185
R22613 outputibias.n51 outputibias.n50 185
R22614 outputibias.n49 outputibias.n48 185
R22615 outputibias.n40 outputibias.n39 185
R22616 outputibias.n43 outputibias.n42 185
R22617 outputibias.n91 outputibias.n90 185
R22618 outputibias.n89 outputibias.n88 185
R22619 outputibias.n68 outputibias.n67 185
R22620 outputibias.n83 outputibias.n82 185
R22621 outputibias.n81 outputibias.n80 185
R22622 outputibias.n72 outputibias.n71 185
R22623 outputibias.n75 outputibias.n74 185
R22624 outputibias.n123 outputibias.n122 185
R22625 outputibias.n121 outputibias.n120 185
R22626 outputibias.n100 outputibias.n99 185
R22627 outputibias.n115 outputibias.n114 185
R22628 outputibias.n113 outputibias.n112 185
R22629 outputibias.n104 outputibias.n103 185
R22630 outputibias.n107 outputibias.n106 185
R22631 outputibias.n0 outputibias.t9 178.945
R22632 outputibias.n133 outputibias.t10 177.018
R22633 outputibias.n132 outputibias.t11 177.018
R22634 outputibias.n0 outputibias.t8 177.018
R22635 outputibias.t7 outputibias.n10 147.661
R22636 outputibias.t1 outputibias.n41 147.661
R22637 outputibias.t3 outputibias.n73 147.661
R22638 outputibias.t5 outputibias.n105 147.661
R22639 outputibias.n128 outputibias.t6 132.363
R22640 outputibias.n128 outputibias.t0 130.436
R22641 outputibias.n129 outputibias.t2 130.436
R22642 outputibias.n130 outputibias.t4 130.436
R22643 outputibias.n27 outputibias.n26 104.615
R22644 outputibias.n26 outputibias.n4 104.615
R22645 outputibias.n19 outputibias.n4 104.615
R22646 outputibias.n19 outputibias.n18 104.615
R22647 outputibias.n18 outputibias.n8 104.615
R22648 outputibias.n11 outputibias.n8 104.615
R22649 outputibias.n58 outputibias.n57 104.615
R22650 outputibias.n57 outputibias.n35 104.615
R22651 outputibias.n50 outputibias.n35 104.615
R22652 outputibias.n50 outputibias.n49 104.615
R22653 outputibias.n49 outputibias.n39 104.615
R22654 outputibias.n42 outputibias.n39 104.615
R22655 outputibias.n90 outputibias.n89 104.615
R22656 outputibias.n89 outputibias.n67 104.615
R22657 outputibias.n82 outputibias.n67 104.615
R22658 outputibias.n82 outputibias.n81 104.615
R22659 outputibias.n81 outputibias.n71 104.615
R22660 outputibias.n74 outputibias.n71 104.615
R22661 outputibias.n122 outputibias.n121 104.615
R22662 outputibias.n121 outputibias.n99 104.615
R22663 outputibias.n114 outputibias.n99 104.615
R22664 outputibias.n114 outputibias.n113 104.615
R22665 outputibias.n113 outputibias.n103 104.615
R22666 outputibias.n106 outputibias.n103 104.615
R22667 outputibias.n63 outputibias.n31 95.6354
R22668 outputibias.n63 outputibias.n62 94.6732
R22669 outputibias.n95 outputibias.n94 94.6732
R22670 outputibias.n127 outputibias.n126 94.6732
R22671 outputibias.n11 outputibias.t7 52.3082
R22672 outputibias.n42 outputibias.t1 52.3082
R22673 outputibias.n74 outputibias.t3 52.3082
R22674 outputibias.n106 outputibias.t5 52.3082
R22675 outputibias.n12 outputibias.n10 15.6674
R22676 outputibias.n43 outputibias.n41 15.6674
R22677 outputibias.n75 outputibias.n73 15.6674
R22678 outputibias.n107 outputibias.n105 15.6674
R22679 outputibias.n13 outputibias.n9 12.8005
R22680 outputibias.n44 outputibias.n40 12.8005
R22681 outputibias.n76 outputibias.n72 12.8005
R22682 outputibias.n108 outputibias.n104 12.8005
R22683 outputibias.n17 outputibias.n16 12.0247
R22684 outputibias.n48 outputibias.n47 12.0247
R22685 outputibias.n80 outputibias.n79 12.0247
R22686 outputibias.n112 outputibias.n111 12.0247
R22687 outputibias.n20 outputibias.n7 11.249
R22688 outputibias.n51 outputibias.n38 11.249
R22689 outputibias.n83 outputibias.n70 11.249
R22690 outputibias.n115 outputibias.n102 11.249
R22691 outputibias.n21 outputibias.n5 10.4732
R22692 outputibias.n52 outputibias.n36 10.4732
R22693 outputibias.n84 outputibias.n68 10.4732
R22694 outputibias.n116 outputibias.n100 10.4732
R22695 outputibias.n25 outputibias.n24 9.69747
R22696 outputibias.n56 outputibias.n55 9.69747
R22697 outputibias.n88 outputibias.n87 9.69747
R22698 outputibias.n120 outputibias.n119 9.69747
R22699 outputibias.n31 outputibias.n30 9.45567
R22700 outputibias.n62 outputibias.n61 9.45567
R22701 outputibias.n94 outputibias.n93 9.45567
R22702 outputibias.n126 outputibias.n125 9.45567
R22703 outputibias.n30 outputibias.n29 9.3005
R22704 outputibias.n3 outputibias.n2 9.3005
R22705 outputibias.n24 outputibias.n23 9.3005
R22706 outputibias.n22 outputibias.n21 9.3005
R22707 outputibias.n7 outputibias.n6 9.3005
R22708 outputibias.n16 outputibias.n15 9.3005
R22709 outputibias.n14 outputibias.n13 9.3005
R22710 outputibias.n61 outputibias.n60 9.3005
R22711 outputibias.n34 outputibias.n33 9.3005
R22712 outputibias.n55 outputibias.n54 9.3005
R22713 outputibias.n53 outputibias.n52 9.3005
R22714 outputibias.n38 outputibias.n37 9.3005
R22715 outputibias.n47 outputibias.n46 9.3005
R22716 outputibias.n45 outputibias.n44 9.3005
R22717 outputibias.n93 outputibias.n92 9.3005
R22718 outputibias.n66 outputibias.n65 9.3005
R22719 outputibias.n87 outputibias.n86 9.3005
R22720 outputibias.n85 outputibias.n84 9.3005
R22721 outputibias.n70 outputibias.n69 9.3005
R22722 outputibias.n79 outputibias.n78 9.3005
R22723 outputibias.n77 outputibias.n76 9.3005
R22724 outputibias.n125 outputibias.n124 9.3005
R22725 outputibias.n98 outputibias.n97 9.3005
R22726 outputibias.n119 outputibias.n118 9.3005
R22727 outputibias.n117 outputibias.n116 9.3005
R22728 outputibias.n102 outputibias.n101 9.3005
R22729 outputibias.n111 outputibias.n110 9.3005
R22730 outputibias.n109 outputibias.n108 9.3005
R22731 outputibias.n28 outputibias.n3 8.92171
R22732 outputibias.n59 outputibias.n34 8.92171
R22733 outputibias.n91 outputibias.n66 8.92171
R22734 outputibias.n123 outputibias.n98 8.92171
R22735 outputibias.n29 outputibias.n1 8.14595
R22736 outputibias.n60 outputibias.n32 8.14595
R22737 outputibias.n92 outputibias.n64 8.14595
R22738 outputibias.n124 outputibias.n96 8.14595
R22739 outputibias.n31 outputibias.n1 5.81868
R22740 outputibias.n62 outputibias.n32 5.81868
R22741 outputibias.n94 outputibias.n64 5.81868
R22742 outputibias.n126 outputibias.n96 5.81868
R22743 outputibias.n131 outputibias.n130 5.20947
R22744 outputibias.n29 outputibias.n28 5.04292
R22745 outputibias.n60 outputibias.n59 5.04292
R22746 outputibias.n92 outputibias.n91 5.04292
R22747 outputibias.n124 outputibias.n123 5.04292
R22748 outputibias.n131 outputibias.n127 4.42209
R22749 outputibias.n14 outputibias.n10 4.38594
R22750 outputibias.n45 outputibias.n41 4.38594
R22751 outputibias.n77 outputibias.n73 4.38594
R22752 outputibias.n109 outputibias.n105 4.38594
R22753 outputibias.n132 outputibias.n131 4.28454
R22754 outputibias.n25 outputibias.n3 4.26717
R22755 outputibias.n56 outputibias.n34 4.26717
R22756 outputibias.n88 outputibias.n66 4.26717
R22757 outputibias.n120 outputibias.n98 4.26717
R22758 outputibias.n24 outputibias.n5 3.49141
R22759 outputibias.n55 outputibias.n36 3.49141
R22760 outputibias.n87 outputibias.n68 3.49141
R22761 outputibias.n119 outputibias.n100 3.49141
R22762 outputibias.n21 outputibias.n20 2.71565
R22763 outputibias.n52 outputibias.n51 2.71565
R22764 outputibias.n84 outputibias.n83 2.71565
R22765 outputibias.n116 outputibias.n115 2.71565
R22766 outputibias.n17 outputibias.n7 1.93989
R22767 outputibias.n48 outputibias.n38 1.93989
R22768 outputibias.n80 outputibias.n70 1.93989
R22769 outputibias.n112 outputibias.n102 1.93989
R22770 outputibias.n130 outputibias.n129 1.9266
R22771 outputibias.n129 outputibias.n128 1.9266
R22772 outputibias.n133 outputibias.n132 1.92658
R22773 outputibias.n134 outputibias.n133 1.29913
R22774 outputibias.n16 outputibias.n9 1.16414
R22775 outputibias.n47 outputibias.n40 1.16414
R22776 outputibias.n79 outputibias.n72 1.16414
R22777 outputibias.n111 outputibias.n104 1.16414
R22778 outputibias.n127 outputibias.n95 0.962709
R22779 outputibias.n95 outputibias.n63 0.962709
R22780 outputibias.n13 outputibias.n12 0.388379
R22781 outputibias.n44 outputibias.n43 0.388379
R22782 outputibias.n76 outputibias.n75 0.388379
R22783 outputibias.n108 outputibias.n107 0.388379
R22784 outputibias.n134 outputibias.n0 0.337251
R22785 outputibias outputibias.n134 0.302375
R22786 outputibias.n30 outputibias.n2 0.155672
R22787 outputibias.n23 outputibias.n2 0.155672
R22788 outputibias.n23 outputibias.n22 0.155672
R22789 outputibias.n22 outputibias.n6 0.155672
R22790 outputibias.n15 outputibias.n6 0.155672
R22791 outputibias.n15 outputibias.n14 0.155672
R22792 outputibias.n61 outputibias.n33 0.155672
R22793 outputibias.n54 outputibias.n33 0.155672
R22794 outputibias.n54 outputibias.n53 0.155672
R22795 outputibias.n53 outputibias.n37 0.155672
R22796 outputibias.n46 outputibias.n37 0.155672
R22797 outputibias.n46 outputibias.n45 0.155672
R22798 outputibias.n93 outputibias.n65 0.155672
R22799 outputibias.n86 outputibias.n65 0.155672
R22800 outputibias.n86 outputibias.n85 0.155672
R22801 outputibias.n85 outputibias.n69 0.155672
R22802 outputibias.n78 outputibias.n69 0.155672
R22803 outputibias.n78 outputibias.n77 0.155672
R22804 outputibias.n125 outputibias.n97 0.155672
R22805 outputibias.n118 outputibias.n97 0.155672
R22806 outputibias.n118 outputibias.n117 0.155672
R22807 outputibias.n117 outputibias.n101 0.155672
R22808 outputibias.n110 outputibias.n101 0.155672
R22809 outputibias.n110 outputibias.n109 0.155672
R22810 a_n2650_8322.n25 a_n2650_8322.t29 74.6477
R22811 a_n2650_8322.n11 a_n2650_8322.t9 74.6477
R22812 a_n2650_8322.n1 a_n2650_8322.t31 74.6474
R22813 a_n2650_8322.n18 a_n2650_8322.t14 74.2899
R22814 a_n2650_8322.n8 a_n2650_8322.t28 74.2899
R22815 a_n2650_8322.n12 a_n2650_8322.t7 74.2899
R22816 a_n2650_8322.n13 a_n2650_8322.t10 74.2899
R22817 a_n2650_8322.n16 a_n2650_8322.t11 74.2899
R22818 a_n2650_8322.n24 a_n2650_8322.n23 70.6783
R22819 a_n2650_8322.n22 a_n2650_8322.n21 70.6783
R22820 a_n2650_8322.n20 a_n2650_8322.n19 70.6783
R22821 a_n2650_8322.n1 a_n2650_8322.n0 70.6783
R22822 a_n2650_8322.n3 a_n2650_8322.n2 70.6783
R22823 a_n2650_8322.n5 a_n2650_8322.n4 70.6783
R22824 a_n2650_8322.n7 a_n2650_8322.n6 70.6783
R22825 a_n2650_8322.n11 a_n2650_8322.n10 70.6783
R22826 a_n2650_8322.n15 a_n2650_8322.n14 70.6783
R22827 a_n2650_8322.n26 a_n2650_8322.n25 70.6782
R22828 a_n2650_8322.n18 a_n2650_8322.n17 24.1867
R22829 a_n2650_8322.n9 a_n2650_8322.t5 9.92253
R22830 a_n2650_8322.n17 a_n2650_8322.n16 7.67184
R22831 a_n2650_8322.n9 a_n2650_8322.n8 6.55222
R22832 a_n2650_8322.n17 a_n2650_8322.n9 5.3452
R22833 a_n2650_8322.n23 a_n2650_8322.t16 3.61217
R22834 a_n2650_8322.n23 a_n2650_8322.t15 3.61217
R22835 a_n2650_8322.n21 a_n2650_8322.t27 3.61217
R22836 a_n2650_8322.n21 a_n2650_8322.t21 3.61217
R22837 a_n2650_8322.n19 a_n2650_8322.t25 3.61217
R22838 a_n2650_8322.n19 a_n2650_8322.t23 3.61217
R22839 a_n2650_8322.n0 a_n2650_8322.t26 3.61217
R22840 a_n2650_8322.n0 a_n2650_8322.t22 3.61217
R22841 a_n2650_8322.n2 a_n2650_8322.t20 3.61217
R22842 a_n2650_8322.n2 a_n2650_8322.t33 3.61217
R22843 a_n2650_8322.n4 a_n2650_8322.t30 3.61217
R22844 a_n2650_8322.n4 a_n2650_8322.t19 3.61217
R22845 a_n2650_8322.n6 a_n2650_8322.t17 3.61217
R22846 a_n2650_8322.n6 a_n2650_8322.t18 3.61217
R22847 a_n2650_8322.n10 a_n2650_8322.t12 3.61217
R22848 a_n2650_8322.n10 a_n2650_8322.t13 3.61217
R22849 a_n2650_8322.n14 a_n2650_8322.t8 3.61217
R22850 a_n2650_8322.n14 a_n2650_8322.t6 3.61217
R22851 a_n2650_8322.t32 a_n2650_8322.n26 3.61217
R22852 a_n2650_8322.n26 a_n2650_8322.t24 3.61217
R22853 a_n2650_8322.n8 a_n2650_8322.n7 0.358259
R22854 a_n2650_8322.n7 a_n2650_8322.n5 0.358259
R22855 a_n2650_8322.n5 a_n2650_8322.n3 0.358259
R22856 a_n2650_8322.n3 a_n2650_8322.n1 0.358259
R22857 a_n2650_8322.n16 a_n2650_8322.n15 0.358259
R22858 a_n2650_8322.n15 a_n2650_8322.n13 0.358259
R22859 a_n2650_8322.n12 a_n2650_8322.n11 0.358259
R22860 a_n2650_8322.n20 a_n2650_8322.n18 0.358259
R22861 a_n2650_8322.n22 a_n2650_8322.n20 0.358259
R22862 a_n2650_8322.n24 a_n2650_8322.n22 0.358259
R22863 a_n2650_8322.n25 a_n2650_8322.n24 0.358259
R22864 a_n2650_8322.n13 a_n2650_8322.n12 0.101793
R22865 a_n2650_8322.t4 a_n2650_8322.t2 0.0788333
R22866 a_n2650_8322.t0 a_n2650_8322.t1 0.0788333
R22867 a_n2650_8322.t5 a_n2650_8322.t3 0.0788333
R22868 a_n2650_8322.t0 a_n2650_8322.t4 0.0318333
R22869 a_n2650_8322.t5 a_n2650_8322.t1 0.0318333
R22870 a_n2650_8322.t2 a_n2650_8322.t1 0.0318333
R22871 a_n2650_8322.t3 a_n2650_8322.t0 0.0318333
R22872 output.n41 output.n15 289.615
R22873 output.n72 output.n46 289.615
R22874 output.n104 output.n78 289.615
R22875 output.n136 output.n110 289.615
R22876 output.n77 output.n45 197.26
R22877 output.n77 output.n76 196.298
R22878 output.n109 output.n108 196.298
R22879 output.n141 output.n140 196.298
R22880 output.n42 output.n41 185
R22881 output.n40 output.n39 185
R22882 output.n19 output.n18 185
R22883 output.n34 output.n33 185
R22884 output.n32 output.n31 185
R22885 output.n23 output.n22 185
R22886 output.n26 output.n25 185
R22887 output.n73 output.n72 185
R22888 output.n71 output.n70 185
R22889 output.n50 output.n49 185
R22890 output.n65 output.n64 185
R22891 output.n63 output.n62 185
R22892 output.n54 output.n53 185
R22893 output.n57 output.n56 185
R22894 output.n105 output.n104 185
R22895 output.n103 output.n102 185
R22896 output.n82 output.n81 185
R22897 output.n97 output.n96 185
R22898 output.n95 output.n94 185
R22899 output.n86 output.n85 185
R22900 output.n89 output.n88 185
R22901 output.n137 output.n136 185
R22902 output.n135 output.n134 185
R22903 output.n114 output.n113 185
R22904 output.n129 output.n128 185
R22905 output.n127 output.n126 185
R22906 output.n118 output.n117 185
R22907 output.n121 output.n120 185
R22908 output.t2 output.n24 147.661
R22909 output.t3 output.n55 147.661
R22910 output.t1 output.n87 147.661
R22911 output.t0 output.n119 147.661
R22912 output.n41 output.n40 104.615
R22913 output.n40 output.n18 104.615
R22914 output.n33 output.n18 104.615
R22915 output.n33 output.n32 104.615
R22916 output.n32 output.n22 104.615
R22917 output.n25 output.n22 104.615
R22918 output.n72 output.n71 104.615
R22919 output.n71 output.n49 104.615
R22920 output.n64 output.n49 104.615
R22921 output.n64 output.n63 104.615
R22922 output.n63 output.n53 104.615
R22923 output.n56 output.n53 104.615
R22924 output.n104 output.n103 104.615
R22925 output.n103 output.n81 104.615
R22926 output.n96 output.n81 104.615
R22927 output.n96 output.n95 104.615
R22928 output.n95 output.n85 104.615
R22929 output.n88 output.n85 104.615
R22930 output.n136 output.n135 104.615
R22931 output.n135 output.n113 104.615
R22932 output.n128 output.n113 104.615
R22933 output.n128 output.n127 104.615
R22934 output.n127 output.n117 104.615
R22935 output.n120 output.n117 104.615
R22936 output.n1 output.t14 77.056
R22937 output.n14 output.t15 76.6694
R22938 output.n1 output.n0 72.7095
R22939 output.n3 output.n2 72.7095
R22940 output.n5 output.n4 72.7095
R22941 output.n7 output.n6 72.7095
R22942 output.n9 output.n8 72.7095
R22943 output.n11 output.n10 72.7095
R22944 output.n13 output.n12 72.7095
R22945 output.n25 output.t2 52.3082
R22946 output.n56 output.t3 52.3082
R22947 output.n88 output.t1 52.3082
R22948 output.n120 output.t0 52.3082
R22949 output.n26 output.n24 15.6674
R22950 output.n57 output.n55 15.6674
R22951 output.n89 output.n87 15.6674
R22952 output.n121 output.n119 15.6674
R22953 output.n27 output.n23 12.8005
R22954 output.n58 output.n54 12.8005
R22955 output.n90 output.n86 12.8005
R22956 output.n122 output.n118 12.8005
R22957 output.n31 output.n30 12.0247
R22958 output.n62 output.n61 12.0247
R22959 output.n94 output.n93 12.0247
R22960 output.n126 output.n125 12.0247
R22961 output.n34 output.n21 11.249
R22962 output.n65 output.n52 11.249
R22963 output.n97 output.n84 11.249
R22964 output.n129 output.n116 11.249
R22965 output.n35 output.n19 10.4732
R22966 output.n66 output.n50 10.4732
R22967 output.n98 output.n82 10.4732
R22968 output.n130 output.n114 10.4732
R22969 output.n39 output.n38 9.69747
R22970 output.n70 output.n69 9.69747
R22971 output.n102 output.n101 9.69747
R22972 output.n134 output.n133 9.69747
R22973 output.n45 output.n44 9.45567
R22974 output.n76 output.n75 9.45567
R22975 output.n108 output.n107 9.45567
R22976 output.n140 output.n139 9.45567
R22977 output.n44 output.n43 9.3005
R22978 output.n17 output.n16 9.3005
R22979 output.n38 output.n37 9.3005
R22980 output.n36 output.n35 9.3005
R22981 output.n21 output.n20 9.3005
R22982 output.n30 output.n29 9.3005
R22983 output.n28 output.n27 9.3005
R22984 output.n75 output.n74 9.3005
R22985 output.n48 output.n47 9.3005
R22986 output.n69 output.n68 9.3005
R22987 output.n67 output.n66 9.3005
R22988 output.n52 output.n51 9.3005
R22989 output.n61 output.n60 9.3005
R22990 output.n59 output.n58 9.3005
R22991 output.n107 output.n106 9.3005
R22992 output.n80 output.n79 9.3005
R22993 output.n101 output.n100 9.3005
R22994 output.n99 output.n98 9.3005
R22995 output.n84 output.n83 9.3005
R22996 output.n93 output.n92 9.3005
R22997 output.n91 output.n90 9.3005
R22998 output.n139 output.n138 9.3005
R22999 output.n112 output.n111 9.3005
R23000 output.n133 output.n132 9.3005
R23001 output.n131 output.n130 9.3005
R23002 output.n116 output.n115 9.3005
R23003 output.n125 output.n124 9.3005
R23004 output.n123 output.n122 9.3005
R23005 output.n42 output.n17 8.92171
R23006 output.n73 output.n48 8.92171
R23007 output.n105 output.n80 8.92171
R23008 output.n137 output.n112 8.92171
R23009 output output.n141 8.15037
R23010 output.n43 output.n15 8.14595
R23011 output.n74 output.n46 8.14595
R23012 output.n106 output.n78 8.14595
R23013 output.n138 output.n110 8.14595
R23014 output.n45 output.n15 5.81868
R23015 output.n76 output.n46 5.81868
R23016 output.n108 output.n78 5.81868
R23017 output.n140 output.n110 5.81868
R23018 output.n43 output.n42 5.04292
R23019 output.n74 output.n73 5.04292
R23020 output.n106 output.n105 5.04292
R23021 output.n138 output.n137 5.04292
R23022 output.n28 output.n24 4.38594
R23023 output.n59 output.n55 4.38594
R23024 output.n91 output.n87 4.38594
R23025 output.n123 output.n119 4.38594
R23026 output.n39 output.n17 4.26717
R23027 output.n70 output.n48 4.26717
R23028 output.n102 output.n80 4.26717
R23029 output.n134 output.n112 4.26717
R23030 output.n0 output.t8 3.9605
R23031 output.n0 output.t6 3.9605
R23032 output.n2 output.t13 3.9605
R23033 output.n2 output.t16 3.9605
R23034 output.n4 output.t18 3.9605
R23035 output.n4 output.t10 3.9605
R23036 output.n6 output.t12 3.9605
R23037 output.n6 output.t19 3.9605
R23038 output.n8 output.t4 3.9605
R23039 output.n8 output.t9 3.9605
R23040 output.n10 output.t11 3.9605
R23041 output.n10 output.t17 3.9605
R23042 output.n12 output.t7 3.9605
R23043 output.n12 output.t5 3.9605
R23044 output.n38 output.n19 3.49141
R23045 output.n69 output.n50 3.49141
R23046 output.n101 output.n82 3.49141
R23047 output.n133 output.n114 3.49141
R23048 output.n35 output.n34 2.71565
R23049 output.n66 output.n65 2.71565
R23050 output.n98 output.n97 2.71565
R23051 output.n130 output.n129 2.71565
R23052 output.n31 output.n21 1.93989
R23053 output.n62 output.n52 1.93989
R23054 output.n94 output.n84 1.93989
R23055 output.n126 output.n116 1.93989
R23056 output.n30 output.n23 1.16414
R23057 output.n61 output.n54 1.16414
R23058 output.n93 output.n86 1.16414
R23059 output.n125 output.n118 1.16414
R23060 output.n141 output.n109 0.962709
R23061 output.n109 output.n77 0.962709
R23062 output.n27 output.n26 0.388379
R23063 output.n58 output.n57 0.388379
R23064 output.n90 output.n89 0.388379
R23065 output.n122 output.n121 0.388379
R23066 output.n14 output.n13 0.387128
R23067 output.n13 output.n11 0.387128
R23068 output.n11 output.n9 0.387128
R23069 output.n9 output.n7 0.387128
R23070 output.n7 output.n5 0.387128
R23071 output.n5 output.n3 0.387128
R23072 output.n3 output.n1 0.387128
R23073 output.n44 output.n16 0.155672
R23074 output.n37 output.n16 0.155672
R23075 output.n37 output.n36 0.155672
R23076 output.n36 output.n20 0.155672
R23077 output.n29 output.n20 0.155672
R23078 output.n29 output.n28 0.155672
R23079 output.n75 output.n47 0.155672
R23080 output.n68 output.n47 0.155672
R23081 output.n68 output.n67 0.155672
R23082 output.n67 output.n51 0.155672
R23083 output.n60 output.n51 0.155672
R23084 output.n60 output.n59 0.155672
R23085 output.n107 output.n79 0.155672
R23086 output.n100 output.n79 0.155672
R23087 output.n100 output.n99 0.155672
R23088 output.n99 output.n83 0.155672
R23089 output.n92 output.n83 0.155672
R23090 output.n92 output.n91 0.155672
R23091 output.n139 output.n111 0.155672
R23092 output.n132 output.n111 0.155672
R23093 output.n132 output.n131 0.155672
R23094 output.n131 output.n115 0.155672
R23095 output.n124 output.n115 0.155672
R23096 output.n124 output.n123 0.155672
R23097 output output.n14 0.126227
R23098 minus.n76 minus.t28 250.337
R23099 minus.n15 minus.t20 250.337
R23100 minus.n126 minus.t1 243.255
R23101 minus.n120 minus.t8 231.093
R23102 minus.n59 minus.t10 231.093
R23103 minus.n125 minus.n123 224.169
R23104 minus.n125 minus.n124 223.454
R23105 minus.n62 minus.t12 187.445
R23106 minus.n113 minus.t18 187.445
R23107 minus.n107 minus.t25 187.445
R23108 minus.n66 minus.t22 187.445
R23109 minus.n68 minus.t19 187.445
R23110 minus.n95 minus.t7 187.445
R23111 minus.n89 minus.t6 187.445
R23112 minus.n72 minus.t16 187.445
R23113 minus.n74 minus.t15 187.445
R23114 minus.n77 minus.t23 187.445
R23115 minus.n16 minus.t14 187.445
R23116 minus.n13 minus.t9 187.445
R23117 minus.n11 minus.t5 187.445
R23118 minus.n28 minus.t26 187.445
R23119 minus.n34 minus.t27 187.445
R23120 minus.n7 minus.t21 187.445
R23121 minus.n5 minus.t24 187.445
R23122 minus.n46 minus.t17 187.445
R23123 minus.n52 minus.t11 187.445
R23124 minus.n1 minus.t13 187.445
R23125 minus.n78 minus.n75 161.3
R23126 minus.n80 minus.n79 161.3
R23127 minus.n82 minus.n81 161.3
R23128 minus.n83 minus.n73 161.3
R23129 minus.n85 minus.n84 161.3
R23130 minus.n87 minus.n86 161.3
R23131 minus.n88 minus.n71 161.3
R23132 minus.n91 minus.n90 161.3
R23133 minus.n92 minus.n70 161.3
R23134 minus.n94 minus.n93 161.3
R23135 minus.n96 minus.n69 161.3
R23136 minus.n98 minus.n97 161.3
R23137 minus.n100 minus.n99 161.3
R23138 minus.n101 minus.n67 161.3
R23139 minus.n103 minus.n102 161.3
R23140 minus.n105 minus.n104 161.3
R23141 minus.n106 minus.n65 161.3
R23142 minus.n109 minus.n108 161.3
R23143 minus.n110 minus.n64 161.3
R23144 minus.n112 minus.n111 161.3
R23145 minus.n114 minus.n63 161.3
R23146 minus.n116 minus.n115 161.3
R23147 minus.n118 minus.n117 161.3
R23148 minus.n119 minus.n61 161.3
R23149 minus.n121 minus.n120 161.3
R23150 minus.n60 minus.n59 161.3
R23151 minus.n58 minus.n0 161.3
R23152 minus.n57 minus.n56 161.3
R23153 minus.n55 minus.n54 161.3
R23154 minus.n53 minus.n2 161.3
R23155 minus.n51 minus.n50 161.3
R23156 minus.n49 minus.n3 161.3
R23157 minus.n48 minus.n47 161.3
R23158 minus.n45 minus.n4 161.3
R23159 minus.n44 minus.n43 161.3
R23160 minus.n42 minus.n41 161.3
R23161 minus.n40 minus.n6 161.3
R23162 minus.n39 minus.n38 161.3
R23163 minus.n37 minus.n36 161.3
R23164 minus.n35 minus.n8 161.3
R23165 minus.n33 minus.n32 161.3
R23166 minus.n31 minus.n9 161.3
R23167 minus.n30 minus.n29 161.3
R23168 minus.n27 minus.n10 161.3
R23169 minus.n26 minus.n25 161.3
R23170 minus.n24 minus.n23 161.3
R23171 minus.n22 minus.n12 161.3
R23172 minus.n21 minus.n20 161.3
R23173 minus.n19 minus.n18 161.3
R23174 minus.n17 minus.n14 161.3
R23175 minus.n106 minus.n105 56.5617
R23176 minus.n97 minus.n96 56.5617
R23177 minus.n88 minus.n87 56.5617
R23178 minus.n27 minus.n26 56.5617
R23179 minus.n36 minus.n35 56.5617
R23180 minus.n45 minus.n44 56.5617
R23181 minus.n115 minus.n114 56.5617
R23182 minus.n79 minus.n78 56.5617
R23183 minus.n18 minus.n17 56.5617
R23184 minus.n54 minus.n53 56.5617
R23185 minus.n119 minus.n118 50.2647
R23186 minus.n58 minus.n57 50.2647
R23187 minus.n108 minus.n64 46.3896
R23188 minus.n84 minus.n83 46.3896
R23189 minus.n23 minus.n22 46.3896
R23190 minus.n47 minus.n3 46.3896
R23191 minus.n76 minus.n75 43.1929
R23192 minus.n15 minus.n14 43.1929
R23193 minus.n101 minus.n100 42.5146
R23194 minus.n94 minus.n70 42.5146
R23195 minus.n33 minus.n9 42.5146
R23196 minus.n40 minus.n39 42.5146
R23197 minus.n77 minus.n76 40.6041
R23198 minus.n16 minus.n15 40.6041
R23199 minus.n102 minus.n101 38.6395
R23200 minus.n90 minus.n70 38.6395
R23201 minus.n29 minus.n9 38.6395
R23202 minus.n41 minus.n40 38.6395
R23203 minus.n122 minus.n121 35.4191
R23204 minus.n112 minus.n64 34.7644
R23205 minus.n83 minus.n82 34.7644
R23206 minus.n22 minus.n21 34.7644
R23207 minus.n51 minus.n3 34.7644
R23208 minus.n114 minus.n113 21.8872
R23209 minus.n79 minus.n74 21.8872
R23210 minus.n18 minus.n13 21.8872
R23211 minus.n53 minus.n52 21.8872
R23212 minus.n105 minus.n66 19.9199
R23213 minus.n89 minus.n88 19.9199
R23214 minus.n28 minus.n27 19.9199
R23215 minus.n44 minus.n5 19.9199
R23216 minus.n124 minus.t0 19.8005
R23217 minus.n124 minus.t2 19.8005
R23218 minus.n123 minus.t4 19.8005
R23219 minus.n123 minus.t3 19.8005
R23220 minus.n97 minus.n68 17.9525
R23221 minus.n96 minus.n95 17.9525
R23222 minus.n35 minus.n34 17.9525
R23223 minus.n36 minus.n7 17.9525
R23224 minus.n107 minus.n106 15.9852
R23225 minus.n87 minus.n72 15.9852
R23226 minus.n26 minus.n11 15.9852
R23227 minus.n46 minus.n45 15.9852
R23228 minus.n115 minus.n62 14.0178
R23229 minus.n78 minus.n77 14.0178
R23230 minus.n17 minus.n16 14.0178
R23231 minus.n54 minus.n1 14.0178
R23232 minus.n122 minus.n60 12.1501
R23233 minus minus.n127 11.5812
R23234 minus.n118 minus.n62 10.575
R23235 minus.n57 minus.n1 10.575
R23236 minus.n120 minus.n119 9.49444
R23237 minus.n59 minus.n58 9.49444
R23238 minus.n108 minus.n107 8.60764
R23239 minus.n84 minus.n72 8.60764
R23240 minus.n23 minus.n11 8.60764
R23241 minus.n47 minus.n46 8.60764
R23242 minus.n100 minus.n68 6.6403
R23243 minus.n95 minus.n94 6.6403
R23244 minus.n34 minus.n33 6.6403
R23245 minus.n39 minus.n7 6.6403
R23246 minus.n127 minus.n126 4.80222
R23247 minus.n102 minus.n66 4.67295
R23248 minus.n90 minus.n89 4.67295
R23249 minus.n29 minus.n28 4.67295
R23250 minus.n41 minus.n5 4.67295
R23251 minus.n113 minus.n112 2.7056
R23252 minus.n82 minus.n74 2.7056
R23253 minus.n21 minus.n13 2.7056
R23254 minus.n52 minus.n51 2.7056
R23255 minus.n127 minus.n122 0.972091
R23256 minus.n126 minus.n125 0.716017
R23257 minus.n121 minus.n61 0.189894
R23258 minus.n117 minus.n61 0.189894
R23259 minus.n117 minus.n116 0.189894
R23260 minus.n116 minus.n63 0.189894
R23261 minus.n111 minus.n63 0.189894
R23262 minus.n111 minus.n110 0.189894
R23263 minus.n110 minus.n109 0.189894
R23264 minus.n109 minus.n65 0.189894
R23265 minus.n104 minus.n65 0.189894
R23266 minus.n104 minus.n103 0.189894
R23267 minus.n103 minus.n67 0.189894
R23268 minus.n99 minus.n67 0.189894
R23269 minus.n99 minus.n98 0.189894
R23270 minus.n98 minus.n69 0.189894
R23271 minus.n93 minus.n69 0.189894
R23272 minus.n93 minus.n92 0.189894
R23273 minus.n92 minus.n91 0.189894
R23274 minus.n91 minus.n71 0.189894
R23275 minus.n86 minus.n71 0.189894
R23276 minus.n86 minus.n85 0.189894
R23277 minus.n85 minus.n73 0.189894
R23278 minus.n81 minus.n73 0.189894
R23279 minus.n81 minus.n80 0.189894
R23280 minus.n80 minus.n75 0.189894
R23281 minus.n19 minus.n14 0.189894
R23282 minus.n20 minus.n19 0.189894
R23283 minus.n20 minus.n12 0.189894
R23284 minus.n24 minus.n12 0.189894
R23285 minus.n25 minus.n24 0.189894
R23286 minus.n25 minus.n10 0.189894
R23287 minus.n30 minus.n10 0.189894
R23288 minus.n31 minus.n30 0.189894
R23289 minus.n32 minus.n31 0.189894
R23290 minus.n32 minus.n8 0.189894
R23291 minus.n37 minus.n8 0.189894
R23292 minus.n38 minus.n37 0.189894
R23293 minus.n38 minus.n6 0.189894
R23294 minus.n42 minus.n6 0.189894
R23295 minus.n43 minus.n42 0.189894
R23296 minus.n43 minus.n4 0.189894
R23297 minus.n48 minus.n4 0.189894
R23298 minus.n49 minus.n48 0.189894
R23299 minus.n50 minus.n49 0.189894
R23300 minus.n50 minus.n2 0.189894
R23301 minus.n55 minus.n2 0.189894
R23302 minus.n56 minus.n55 0.189894
R23303 minus.n56 minus.n0 0.189894
R23304 minus.n60 minus.n0 0.189894
R23305 diffpairibias.n0 diffpairibias.t18 436.822
R23306 diffpairibias.n21 diffpairibias.t19 435.479
R23307 diffpairibias.n20 diffpairibias.t16 435.479
R23308 diffpairibias.n19 diffpairibias.t17 435.479
R23309 diffpairibias.n18 diffpairibias.t21 435.479
R23310 diffpairibias.n0 diffpairibias.t22 435.479
R23311 diffpairibias.n1 diffpairibias.t20 435.479
R23312 diffpairibias.n2 diffpairibias.t23 435.479
R23313 diffpairibias.n10 diffpairibias.t0 377.536
R23314 diffpairibias.n10 diffpairibias.t8 376.193
R23315 diffpairibias.n11 diffpairibias.t10 376.193
R23316 diffpairibias.n12 diffpairibias.t6 376.193
R23317 diffpairibias.n13 diffpairibias.t2 376.193
R23318 diffpairibias.n14 diffpairibias.t12 376.193
R23319 diffpairibias.n15 diffpairibias.t4 376.193
R23320 diffpairibias.n16 diffpairibias.t14 376.193
R23321 diffpairibias.n3 diffpairibias.t1 113.368
R23322 diffpairibias.n3 diffpairibias.t9 112.698
R23323 diffpairibias.n4 diffpairibias.t11 112.698
R23324 diffpairibias.n5 diffpairibias.t7 112.698
R23325 diffpairibias.n6 diffpairibias.t3 112.698
R23326 diffpairibias.n7 diffpairibias.t13 112.698
R23327 diffpairibias.n8 diffpairibias.t5 112.698
R23328 diffpairibias.n9 diffpairibias.t15 112.698
R23329 diffpairibias.n17 diffpairibias.n16 4.77242
R23330 diffpairibias.n17 diffpairibias.n9 4.30807
R23331 diffpairibias.n18 diffpairibias.n17 4.13945
R23332 diffpairibias.n16 diffpairibias.n15 1.34352
R23333 diffpairibias.n15 diffpairibias.n14 1.34352
R23334 diffpairibias.n14 diffpairibias.n13 1.34352
R23335 diffpairibias.n13 diffpairibias.n12 1.34352
R23336 diffpairibias.n12 diffpairibias.n11 1.34352
R23337 diffpairibias.n11 diffpairibias.n10 1.34352
R23338 diffpairibias.n2 diffpairibias.n1 1.34352
R23339 diffpairibias.n1 diffpairibias.n0 1.34352
R23340 diffpairibias.n19 diffpairibias.n18 1.34352
R23341 diffpairibias.n20 diffpairibias.n19 1.34352
R23342 diffpairibias.n21 diffpairibias.n20 1.34352
R23343 diffpairibias.n22 diffpairibias.n21 0.862419
R23344 diffpairibias diffpairibias.n22 0.684875
R23345 diffpairibias.n9 diffpairibias.n8 0.672012
R23346 diffpairibias.n8 diffpairibias.n7 0.672012
R23347 diffpairibias.n7 diffpairibias.n6 0.672012
R23348 diffpairibias.n6 diffpairibias.n5 0.672012
R23349 diffpairibias.n5 diffpairibias.n4 0.672012
R23350 diffpairibias.n4 diffpairibias.n3 0.672012
R23351 diffpairibias.n22 diffpairibias.n2 0.190907
C0 minus diffpairibias 5.39e-19
C1 commonsourceibias output 0.006808f
C2 CSoutput minus 2.80108f
C3 vdd plus 0.079456f
C4 commonsourceibias outputibias 0.003832f
C5 plus diffpairibias 4.4e-19
C6 vdd commonsourceibias 0.004218f
C7 CSoutput plus 0.9147f
C8 commonsourceibias diffpairibias 0.052851f
C9 CSoutput commonsourceibias 44.9728f
C10 minus plus 10.4342f
C11 minus commonsourceibias 0.515369f
C12 plus commonsourceibias 0.498793f
C13 output outputibias 2.34152f
C14 vdd output 7.23429f
C15 CSoutput output 6.13571f
C16 CSoutput outputibias 0.032386f
C17 vdd CSoutput 68.27061f
C18 diffpairibias gnd 48.95304f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.180656p
C22 plus gnd 39.3442f
C23 minus gnd 31.211967f
C24 CSoutput gnd 0.114563p
C25 vdd gnd 0.415267p
C26 diffpairibias.t18 gnd 0.087401f
C27 diffpairibias.t22 gnd 0.087239f
C28 diffpairibias.n0 gnd 0.102784f
C29 diffpairibias.t20 gnd 0.087239f
C30 diffpairibias.n1 gnd 0.050171f
C31 diffpairibias.t23 gnd 0.087239f
C32 diffpairibias.n2 gnd 0.039841f
C33 diffpairibias.t1 gnd 0.083757f
C34 diffpairibias.t9 gnd 0.083392f
C35 diffpairibias.n3 gnd 0.131682f
C36 diffpairibias.t11 gnd 0.083392f
C37 diffpairibias.n4 gnd 0.07027f
C38 diffpairibias.t7 gnd 0.083392f
C39 diffpairibias.n5 gnd 0.07027f
C40 diffpairibias.t3 gnd 0.083392f
C41 diffpairibias.n6 gnd 0.07027f
C42 diffpairibias.t13 gnd 0.083392f
C43 diffpairibias.n7 gnd 0.07027f
C44 diffpairibias.t5 gnd 0.083392f
C45 diffpairibias.n8 gnd 0.07027f
C46 diffpairibias.t15 gnd 0.083392f
C47 diffpairibias.n9 gnd 0.099771f
C48 diffpairibias.t0 gnd 0.08427f
C49 diffpairibias.t8 gnd 0.084123f
C50 diffpairibias.n10 gnd 0.091784f
C51 diffpairibias.t10 gnd 0.084123f
C52 diffpairibias.n11 gnd 0.050681f
C53 diffpairibias.t6 gnd 0.084123f
C54 diffpairibias.n12 gnd 0.050681f
C55 diffpairibias.t2 gnd 0.084123f
C56 diffpairibias.n13 gnd 0.050681f
C57 diffpairibias.t12 gnd 0.084123f
C58 diffpairibias.n14 gnd 0.050681f
C59 diffpairibias.t4 gnd 0.084123f
C60 diffpairibias.n15 gnd 0.050681f
C61 diffpairibias.t14 gnd 0.084123f
C62 diffpairibias.n16 gnd 0.059977f
C63 diffpairibias.n17 gnd 0.226448f
C64 diffpairibias.t21 gnd 0.087239f
C65 diffpairibias.n18 gnd 0.050181f
C66 diffpairibias.t17 gnd 0.087239f
C67 diffpairibias.n19 gnd 0.050171f
C68 diffpairibias.t16 gnd 0.087239f
C69 diffpairibias.n20 gnd 0.050171f
C70 diffpairibias.t19 gnd 0.087239f
C71 diffpairibias.n21 gnd 0.045859f
C72 diffpairibias.n22 gnd 0.046268f
C73 minus.n0 gnd 0.030662f
C74 minus.t13 gnd 0.515581f
C75 minus.n1 gnd 0.208524f
C76 minus.n2 gnd 0.030662f
C77 minus.t11 gnd 0.515581f
C78 minus.n3 gnd 0.026202f
C79 minus.n4 gnd 0.030662f
C80 minus.t17 gnd 0.515581f
C81 minus.t24 gnd 0.515581f
C82 minus.n5 gnd 0.208524f
C83 minus.n6 gnd 0.030662f
C84 minus.t21 gnd 0.515581f
C85 minus.n7 gnd 0.208524f
C86 minus.n8 gnd 0.030662f
C87 minus.t27 gnd 0.515581f
C88 minus.n9 gnd 0.024922f
C89 minus.n10 gnd 0.030662f
C90 minus.t26 gnd 0.515581f
C91 minus.t5 gnd 0.515581f
C92 minus.n11 gnd 0.208524f
C93 minus.n12 gnd 0.030662f
C94 minus.t9 gnd 0.515581f
C95 minus.n13 gnd 0.208524f
C96 minus.n14 gnd 0.130127f
C97 minus.t14 gnd 0.515581f
C98 minus.t20 gnd 0.576771f
C99 minus.n15 gnd 0.243785f
C100 minus.n16 gnd 0.238799f
C101 minus.n17 gnd 0.039289f
C102 minus.n18 gnd 0.034698f
C103 minus.n19 gnd 0.030662f
C104 minus.n20 gnd 0.030662f
C105 minus.n21 gnd 0.036642f
C106 minus.n22 gnd 0.026202f
C107 minus.n23 gnd 0.039934f
C108 minus.n24 gnd 0.030662f
C109 minus.n25 gnd 0.030662f
C110 minus.n26 gnd 0.038141f
C111 minus.n27 gnd 0.035846f
C112 minus.n28 gnd 0.208524f
C113 minus.n29 gnd 0.038409f
C114 minus.n30 gnd 0.030662f
C115 minus.n31 gnd 0.030662f
C116 minus.n32 gnd 0.030662f
C117 minus.n33 gnd 0.039446f
C118 minus.n34 gnd 0.208524f
C119 minus.n35 gnd 0.036993f
C120 minus.n36 gnd 0.036993f
C121 minus.n37 gnd 0.030662f
C122 minus.n38 gnd 0.030662f
C123 minus.n39 gnd 0.039446f
C124 minus.n40 gnd 0.024922f
C125 minus.n41 gnd 0.038409f
C126 minus.n42 gnd 0.030662f
C127 minus.n43 gnd 0.030662f
C128 minus.n44 gnd 0.035846f
C129 minus.n45 gnd 0.038141f
C130 minus.n46 gnd 0.208524f
C131 minus.n47 gnd 0.039934f
C132 minus.n48 gnd 0.030662f
C133 minus.n49 gnd 0.030662f
C134 minus.n50 gnd 0.030662f
C135 minus.n51 gnd 0.036642f
C136 minus.n52 gnd 0.208524f
C137 minus.n53 gnd 0.034698f
C138 minus.n54 gnd 0.039289f
C139 minus.n55 gnd 0.030662f
C140 minus.n56 gnd 0.030662f
C141 minus.n57 gnd 0.04f
C142 minus.n58 gnd 0.011144f
C143 minus.t10 gnd 0.557601f
C144 minus.n59 gnd 0.241436f
C145 minus.n60 gnd 0.359197f
C146 minus.n61 gnd 0.030662f
C147 minus.t8 gnd 0.557601f
C148 minus.t12 gnd 0.515581f
C149 minus.n62 gnd 0.208524f
C150 minus.n63 gnd 0.030662f
C151 minus.t18 gnd 0.515581f
C152 minus.n64 gnd 0.026202f
C153 minus.n65 gnd 0.030662f
C154 minus.t25 gnd 0.515581f
C155 minus.t22 gnd 0.515581f
C156 minus.n66 gnd 0.208524f
C157 minus.n67 gnd 0.030662f
C158 minus.t19 gnd 0.515581f
C159 minus.n68 gnd 0.208524f
C160 minus.n69 gnd 0.030662f
C161 minus.t7 gnd 0.515581f
C162 minus.n70 gnd 0.024922f
C163 minus.n71 gnd 0.030662f
C164 minus.t6 gnd 0.515581f
C165 minus.t16 gnd 0.515581f
C166 minus.n72 gnd 0.208524f
C167 minus.n73 gnd 0.030662f
C168 minus.t15 gnd 0.515581f
C169 minus.n74 gnd 0.208524f
C170 minus.n75 gnd 0.130127f
C171 minus.t23 gnd 0.515581f
C172 minus.t28 gnd 0.576771f
C173 minus.n76 gnd 0.243785f
C174 minus.n77 gnd 0.238799f
C175 minus.n78 gnd 0.039289f
C176 minus.n79 gnd 0.034698f
C177 minus.n80 gnd 0.030662f
C178 minus.n81 gnd 0.030662f
C179 minus.n82 gnd 0.036642f
C180 minus.n83 gnd 0.026202f
C181 minus.n84 gnd 0.039934f
C182 minus.n85 gnd 0.030662f
C183 minus.n86 gnd 0.030662f
C184 minus.n87 gnd 0.038141f
C185 minus.n88 gnd 0.035846f
C186 minus.n89 gnd 0.208524f
C187 minus.n90 gnd 0.038409f
C188 minus.n91 gnd 0.030662f
C189 minus.n92 gnd 0.030662f
C190 minus.n93 gnd 0.030662f
C191 minus.n94 gnd 0.039446f
C192 minus.n95 gnd 0.208524f
C193 minus.n96 gnd 0.036993f
C194 minus.n97 gnd 0.036993f
C195 minus.n98 gnd 0.030662f
C196 minus.n99 gnd 0.030662f
C197 minus.n100 gnd 0.039446f
C198 minus.n101 gnd 0.024922f
C199 minus.n102 gnd 0.038409f
C200 minus.n103 gnd 0.030662f
C201 minus.n104 gnd 0.030662f
C202 minus.n105 gnd 0.035846f
C203 minus.n106 gnd 0.038141f
C204 minus.n107 gnd 0.208524f
C205 minus.n108 gnd 0.039934f
C206 minus.n109 gnd 0.030662f
C207 minus.n110 gnd 0.030662f
C208 minus.n111 gnd 0.030662f
C209 minus.n112 gnd 0.036642f
C210 minus.n113 gnd 0.208524f
C211 minus.n114 gnd 0.034698f
C212 minus.n115 gnd 0.039289f
C213 minus.n116 gnd 0.030662f
C214 minus.n117 gnd 0.030662f
C215 minus.n118 gnd 0.04f
C216 minus.n119 gnd 0.011144f
C217 minus.n120 gnd 0.241436f
C218 minus.n121 gnd 1.11855f
C219 minus.n122 gnd 1.64306f
C220 minus.t4 gnd 0.009452f
C221 minus.t3 gnd 0.009452f
C222 minus.n123 gnd 0.031081f
C223 minus.t0 gnd 0.009452f
C224 minus.t2 gnd 0.009452f
C225 minus.n124 gnd 0.030655f
C226 minus.n125 gnd 0.26163f
C227 minus.t1 gnd 0.05261f
C228 minus.n126 gnd 0.142769f
C229 minus.n127 gnd 1.95331f
C230 output.t14 gnd 0.464308f
C231 output.t8 gnd 0.044422f
C232 output.t6 gnd 0.044422f
C233 output.n0 gnd 0.364624f
C234 output.n1 gnd 0.614102f
C235 output.t13 gnd 0.044422f
C236 output.t16 gnd 0.044422f
C237 output.n2 gnd 0.364624f
C238 output.n3 gnd 0.350265f
C239 output.t18 gnd 0.044422f
C240 output.t10 gnd 0.044422f
C241 output.n4 gnd 0.364624f
C242 output.n5 gnd 0.350265f
C243 output.t12 gnd 0.044422f
C244 output.t19 gnd 0.044422f
C245 output.n6 gnd 0.364624f
C246 output.n7 gnd 0.350265f
C247 output.t4 gnd 0.044422f
C248 output.t9 gnd 0.044422f
C249 output.n8 gnd 0.364624f
C250 output.n9 gnd 0.350265f
C251 output.t11 gnd 0.044422f
C252 output.t17 gnd 0.044422f
C253 output.n10 gnd 0.364624f
C254 output.n11 gnd 0.350265f
C255 output.t7 gnd 0.044422f
C256 output.t5 gnd 0.044422f
C257 output.n12 gnd 0.364624f
C258 output.n13 gnd 0.350265f
C259 output.t15 gnd 0.462979f
C260 output.n14 gnd 0.28994f
C261 output.n15 gnd 0.015803f
C262 output.n16 gnd 0.011243f
C263 output.n17 gnd 0.006041f
C264 output.n18 gnd 0.01428f
C265 output.n19 gnd 0.006397f
C266 output.n20 gnd 0.011243f
C267 output.n21 gnd 0.006041f
C268 output.n22 gnd 0.01428f
C269 output.n23 gnd 0.006397f
C270 output.n24 gnd 0.048111f
C271 output.t2 gnd 0.023274f
C272 output.n25 gnd 0.01071f
C273 output.n26 gnd 0.008435f
C274 output.n27 gnd 0.006041f
C275 output.n28 gnd 0.267512f
C276 output.n29 gnd 0.011243f
C277 output.n30 gnd 0.006041f
C278 output.n31 gnd 0.006397f
C279 output.n32 gnd 0.01428f
C280 output.n33 gnd 0.01428f
C281 output.n34 gnd 0.006397f
C282 output.n35 gnd 0.006041f
C283 output.n36 gnd 0.011243f
C284 output.n37 gnd 0.011243f
C285 output.n38 gnd 0.006041f
C286 output.n39 gnd 0.006397f
C287 output.n40 gnd 0.01428f
C288 output.n41 gnd 0.030913f
C289 output.n42 gnd 0.006397f
C290 output.n43 gnd 0.006041f
C291 output.n44 gnd 0.025987f
C292 output.n45 gnd 0.097665f
C293 output.n46 gnd 0.015803f
C294 output.n47 gnd 0.011243f
C295 output.n48 gnd 0.006041f
C296 output.n49 gnd 0.01428f
C297 output.n50 gnd 0.006397f
C298 output.n51 gnd 0.011243f
C299 output.n52 gnd 0.006041f
C300 output.n53 gnd 0.01428f
C301 output.n54 gnd 0.006397f
C302 output.n55 gnd 0.048111f
C303 output.t3 gnd 0.023274f
C304 output.n56 gnd 0.01071f
C305 output.n57 gnd 0.008435f
C306 output.n58 gnd 0.006041f
C307 output.n59 gnd 0.267512f
C308 output.n60 gnd 0.011243f
C309 output.n61 gnd 0.006041f
C310 output.n62 gnd 0.006397f
C311 output.n63 gnd 0.01428f
C312 output.n64 gnd 0.01428f
C313 output.n65 gnd 0.006397f
C314 output.n66 gnd 0.006041f
C315 output.n67 gnd 0.011243f
C316 output.n68 gnd 0.011243f
C317 output.n69 gnd 0.006041f
C318 output.n70 gnd 0.006397f
C319 output.n71 gnd 0.01428f
C320 output.n72 gnd 0.030913f
C321 output.n73 gnd 0.006397f
C322 output.n74 gnd 0.006041f
C323 output.n75 gnd 0.025987f
C324 output.n76 gnd 0.09306f
C325 output.n77 gnd 1.65264f
C326 output.n78 gnd 0.015803f
C327 output.n79 gnd 0.011243f
C328 output.n80 gnd 0.006041f
C329 output.n81 gnd 0.01428f
C330 output.n82 gnd 0.006397f
C331 output.n83 gnd 0.011243f
C332 output.n84 gnd 0.006041f
C333 output.n85 gnd 0.01428f
C334 output.n86 gnd 0.006397f
C335 output.n87 gnd 0.048111f
C336 output.t1 gnd 0.023274f
C337 output.n88 gnd 0.01071f
C338 output.n89 gnd 0.008435f
C339 output.n90 gnd 0.006041f
C340 output.n91 gnd 0.267512f
C341 output.n92 gnd 0.011243f
C342 output.n93 gnd 0.006041f
C343 output.n94 gnd 0.006397f
C344 output.n95 gnd 0.01428f
C345 output.n96 gnd 0.01428f
C346 output.n97 gnd 0.006397f
C347 output.n98 gnd 0.006041f
C348 output.n99 gnd 0.011243f
C349 output.n100 gnd 0.011243f
C350 output.n101 gnd 0.006041f
C351 output.n102 gnd 0.006397f
C352 output.n103 gnd 0.01428f
C353 output.n104 gnd 0.030913f
C354 output.n105 gnd 0.006397f
C355 output.n106 gnd 0.006041f
C356 output.n107 gnd 0.025987f
C357 output.n108 gnd 0.09306f
C358 output.n109 gnd 0.713089f
C359 output.n110 gnd 0.015803f
C360 output.n111 gnd 0.011243f
C361 output.n112 gnd 0.006041f
C362 output.n113 gnd 0.01428f
C363 output.n114 gnd 0.006397f
C364 output.n115 gnd 0.011243f
C365 output.n116 gnd 0.006041f
C366 output.n117 gnd 0.01428f
C367 output.n118 gnd 0.006397f
C368 output.n119 gnd 0.048111f
C369 output.t0 gnd 0.023274f
C370 output.n120 gnd 0.01071f
C371 output.n121 gnd 0.008435f
C372 output.n122 gnd 0.006041f
C373 output.n123 gnd 0.267512f
C374 output.n124 gnd 0.011243f
C375 output.n125 gnd 0.006041f
C376 output.n126 gnd 0.006397f
C377 output.n127 gnd 0.01428f
C378 output.n128 gnd 0.01428f
C379 output.n129 gnd 0.006397f
C380 output.n130 gnd 0.006041f
C381 output.n131 gnd 0.011243f
C382 output.n132 gnd 0.011243f
C383 output.n133 gnd 0.006041f
C384 output.n134 gnd 0.006397f
C385 output.n135 gnd 0.01428f
C386 output.n136 gnd 0.030913f
C387 output.n137 gnd 0.006397f
C388 output.n138 gnd 0.006041f
C389 output.n139 gnd 0.025987f
C390 output.n140 gnd 0.09306f
C391 output.n141 gnd 1.67353f
C392 a_n2650_8322.t24 gnd 0.09797f
C393 a_n2650_8322.t1 gnd 20.3248f
C394 a_n2650_8322.t2 gnd 20.1823f
C395 a_n2650_8322.t4 gnd 20.1823f
C396 a_n2650_8322.t0 gnd 20.3248f
C397 a_n2650_8322.t3 gnd 20.1823f
C398 a_n2650_8322.t5 gnd 29.385302f
C399 a_n2650_8322.t31 gnd 0.917342f
C400 a_n2650_8322.t26 gnd 0.09797f
C401 a_n2650_8322.t22 gnd 0.09797f
C402 a_n2650_8322.n0 gnd 0.690103f
C403 a_n2650_8322.n1 gnd 0.77109f
C404 a_n2650_8322.t20 gnd 0.09797f
C405 a_n2650_8322.t33 gnd 0.09797f
C406 a_n2650_8322.n2 gnd 0.690103f
C407 a_n2650_8322.n3 gnd 0.39178f
C408 a_n2650_8322.t30 gnd 0.09797f
C409 a_n2650_8322.t19 gnd 0.09797f
C410 a_n2650_8322.n4 gnd 0.690103f
C411 a_n2650_8322.n5 gnd 0.39178f
C412 a_n2650_8322.t17 gnd 0.09797f
C413 a_n2650_8322.t18 gnd 0.09797f
C414 a_n2650_8322.n6 gnd 0.690103f
C415 a_n2650_8322.n7 gnd 0.39178f
C416 a_n2650_8322.t28 gnd 0.915517f
C417 a_n2650_8322.n8 gnd 0.995819f
C418 a_n2650_8322.n9 gnd 3.63884f
C419 a_n2650_8322.t9 gnd 0.917344f
C420 a_n2650_8322.t12 gnd 0.09797f
C421 a_n2650_8322.t13 gnd 0.09797f
C422 a_n2650_8322.n10 gnd 0.690103f
C423 a_n2650_8322.n11 gnd 0.771088f
C424 a_n2650_8322.t7 gnd 0.915517f
C425 a_n2650_8322.n12 gnd 0.388022f
C426 a_n2650_8322.t10 gnd 0.915517f
C427 a_n2650_8322.n13 gnd 0.388022f
C428 a_n2650_8322.t8 gnd 0.09797f
C429 a_n2650_8322.t6 gnd 0.09797f
C430 a_n2650_8322.n14 gnd 0.690103f
C431 a_n2650_8322.n15 gnd 0.39178f
C432 a_n2650_8322.t11 gnd 0.915517f
C433 a_n2650_8322.n16 gnd 1.27304f
C434 a_n2650_8322.n17 gnd 2.08003f
C435 a_n2650_8322.t14 gnd 0.915517f
C436 a_n2650_8322.n18 gnd 1.70845f
C437 a_n2650_8322.t25 gnd 0.09797f
C438 a_n2650_8322.t23 gnd 0.09797f
C439 a_n2650_8322.n19 gnd 0.690103f
C440 a_n2650_8322.n20 gnd 0.39178f
C441 a_n2650_8322.t27 gnd 0.09797f
C442 a_n2650_8322.t21 gnd 0.09797f
C443 a_n2650_8322.n21 gnd 0.690103f
C444 a_n2650_8322.n22 gnd 0.39178f
C445 a_n2650_8322.t16 gnd 0.09797f
C446 a_n2650_8322.t15 gnd 0.09797f
C447 a_n2650_8322.n23 gnd 0.690103f
C448 a_n2650_8322.n24 gnd 0.39178f
C449 a_n2650_8322.t29 gnd 0.917344f
C450 a_n2650_8322.n25 gnd 0.771086f
C451 a_n2650_8322.n26 gnd 0.690105f
C452 a_n2650_8322.t32 gnd 0.09797f
C453 outputibias.t8 gnd 0.11477f
C454 outputibias.t9 gnd 0.115567f
C455 outputibias.n0 gnd 0.130108f
C456 outputibias.n1 gnd 0.001372f
C457 outputibias.n2 gnd 9.76e-19
C458 outputibias.n3 gnd 5.24e-19
C459 outputibias.n4 gnd 0.001239f
C460 outputibias.n5 gnd 5.55e-19
C461 outputibias.n6 gnd 9.76e-19
C462 outputibias.n7 gnd 5.24e-19
C463 outputibias.n8 gnd 0.001239f
C464 outputibias.n9 gnd 5.55e-19
C465 outputibias.n10 gnd 0.004176f
C466 outputibias.t7 gnd 0.00202f
C467 outputibias.n11 gnd 9.3e-19
C468 outputibias.n12 gnd 7.32e-19
C469 outputibias.n13 gnd 5.24e-19
C470 outputibias.n14 gnd 0.02322f
C471 outputibias.n15 gnd 9.76e-19
C472 outputibias.n16 gnd 5.24e-19
C473 outputibias.n17 gnd 5.55e-19
C474 outputibias.n18 gnd 0.001239f
C475 outputibias.n19 gnd 0.001239f
C476 outputibias.n20 gnd 5.55e-19
C477 outputibias.n21 gnd 5.24e-19
C478 outputibias.n22 gnd 9.76e-19
C479 outputibias.n23 gnd 9.76e-19
C480 outputibias.n24 gnd 5.24e-19
C481 outputibias.n25 gnd 5.55e-19
C482 outputibias.n26 gnd 0.001239f
C483 outputibias.n27 gnd 0.002683f
C484 outputibias.n28 gnd 5.55e-19
C485 outputibias.n29 gnd 5.24e-19
C486 outputibias.n30 gnd 0.002256f
C487 outputibias.n31 gnd 0.005781f
C488 outputibias.n32 gnd 0.001372f
C489 outputibias.n33 gnd 9.76e-19
C490 outputibias.n34 gnd 5.24e-19
C491 outputibias.n35 gnd 0.001239f
C492 outputibias.n36 gnd 5.55e-19
C493 outputibias.n37 gnd 9.76e-19
C494 outputibias.n38 gnd 5.24e-19
C495 outputibias.n39 gnd 0.001239f
C496 outputibias.n40 gnd 5.55e-19
C497 outputibias.n41 gnd 0.004176f
C498 outputibias.t1 gnd 0.00202f
C499 outputibias.n42 gnd 9.3e-19
C500 outputibias.n43 gnd 7.32e-19
C501 outputibias.n44 gnd 5.24e-19
C502 outputibias.n45 gnd 0.02322f
C503 outputibias.n46 gnd 9.76e-19
C504 outputibias.n47 gnd 5.24e-19
C505 outputibias.n48 gnd 5.55e-19
C506 outputibias.n49 gnd 0.001239f
C507 outputibias.n50 gnd 0.001239f
C508 outputibias.n51 gnd 5.55e-19
C509 outputibias.n52 gnd 5.24e-19
C510 outputibias.n53 gnd 9.76e-19
C511 outputibias.n54 gnd 9.76e-19
C512 outputibias.n55 gnd 5.24e-19
C513 outputibias.n56 gnd 5.55e-19
C514 outputibias.n57 gnd 0.001239f
C515 outputibias.n58 gnd 0.002683f
C516 outputibias.n59 gnd 5.55e-19
C517 outputibias.n60 gnd 5.24e-19
C518 outputibias.n61 gnd 0.002256f
C519 outputibias.n62 gnd 0.005197f
C520 outputibias.n63 gnd 0.121892f
C521 outputibias.n64 gnd 0.001372f
C522 outputibias.n65 gnd 9.76e-19
C523 outputibias.n66 gnd 5.24e-19
C524 outputibias.n67 gnd 0.001239f
C525 outputibias.n68 gnd 5.55e-19
C526 outputibias.n69 gnd 9.76e-19
C527 outputibias.n70 gnd 5.24e-19
C528 outputibias.n71 gnd 0.001239f
C529 outputibias.n72 gnd 5.55e-19
C530 outputibias.n73 gnd 0.004176f
C531 outputibias.t3 gnd 0.00202f
C532 outputibias.n74 gnd 9.3e-19
C533 outputibias.n75 gnd 7.32e-19
C534 outputibias.n76 gnd 5.24e-19
C535 outputibias.n77 gnd 0.02322f
C536 outputibias.n78 gnd 9.76e-19
C537 outputibias.n79 gnd 5.24e-19
C538 outputibias.n80 gnd 5.55e-19
C539 outputibias.n81 gnd 0.001239f
C540 outputibias.n82 gnd 0.001239f
C541 outputibias.n83 gnd 5.55e-19
C542 outputibias.n84 gnd 5.24e-19
C543 outputibias.n85 gnd 9.76e-19
C544 outputibias.n86 gnd 9.76e-19
C545 outputibias.n87 gnd 5.24e-19
C546 outputibias.n88 gnd 5.55e-19
C547 outputibias.n89 gnd 0.001239f
C548 outputibias.n90 gnd 0.002683f
C549 outputibias.n91 gnd 5.55e-19
C550 outputibias.n92 gnd 5.24e-19
C551 outputibias.n93 gnd 0.002256f
C552 outputibias.n94 gnd 0.005197f
C553 outputibias.n95 gnd 0.064513f
C554 outputibias.n96 gnd 0.001372f
C555 outputibias.n97 gnd 9.76e-19
C556 outputibias.n98 gnd 5.24e-19
C557 outputibias.n99 gnd 0.001239f
C558 outputibias.n100 gnd 5.55e-19
C559 outputibias.n101 gnd 9.76e-19
C560 outputibias.n102 gnd 5.24e-19
C561 outputibias.n103 gnd 0.001239f
C562 outputibias.n104 gnd 5.55e-19
C563 outputibias.n105 gnd 0.004176f
C564 outputibias.t5 gnd 0.00202f
C565 outputibias.n106 gnd 9.3e-19
C566 outputibias.n107 gnd 7.32e-19
C567 outputibias.n108 gnd 5.24e-19
C568 outputibias.n109 gnd 0.02322f
C569 outputibias.n110 gnd 9.76e-19
C570 outputibias.n111 gnd 5.24e-19
C571 outputibias.n112 gnd 5.55e-19
C572 outputibias.n113 gnd 0.001239f
C573 outputibias.n114 gnd 0.001239f
C574 outputibias.n115 gnd 5.55e-19
C575 outputibias.n116 gnd 5.24e-19
C576 outputibias.n117 gnd 9.76e-19
C577 outputibias.n118 gnd 9.76e-19
C578 outputibias.n119 gnd 5.24e-19
C579 outputibias.n120 gnd 5.55e-19
C580 outputibias.n121 gnd 0.001239f
C581 outputibias.n122 gnd 0.002683f
C582 outputibias.n123 gnd 5.55e-19
C583 outputibias.n124 gnd 5.24e-19
C584 outputibias.n125 gnd 0.002256f
C585 outputibias.n126 gnd 0.005197f
C586 outputibias.n127 gnd 0.084814f
C587 outputibias.t4 gnd 0.108319f
C588 outputibias.t2 gnd 0.108319f
C589 outputibias.t0 gnd 0.108319f
C590 outputibias.t6 gnd 0.109238f
C591 outputibias.n128 gnd 0.134674f
C592 outputibias.n129 gnd 0.07244f
C593 outputibias.n130 gnd 0.079818f
C594 outputibias.n131 gnd 0.164901f
C595 outputibias.t11 gnd 0.11477f
C596 outputibias.n132 gnd 0.067481f
C597 outputibias.t10 gnd 0.11477f
C598 outputibias.n133 gnd 0.065115f
C599 outputibias.n134 gnd 0.029159f
C600 a_n3106_n452.t12 gnd 0.10001f
C601 a_n3106_n452.t23 gnd 1.03942f
C602 a_n3106_n452.n0 gnd 0.392946f
C603 a_n3106_n452.t2 gnd 1.29145f
C604 a_n3106_n452.n1 gnd 1.22854f
C605 a_n3106_n452.t55 gnd 1.03942f
C606 a_n3106_n452.n2 gnd 0.392946f
C607 a_n3106_n452.t48 gnd 0.10001f
C608 a_n3106_n452.t5 gnd 0.10001f
C609 a_n3106_n452.n3 gnd 0.816794f
C610 a_n3106_n452.n4 gnd 0.411618f
C611 a_n3106_n452.t40 gnd 0.10001f
C612 a_n3106_n452.t47 gnd 0.10001f
C613 a_n3106_n452.n5 gnd 0.816794f
C614 a_n3106_n452.n6 gnd 0.411618f
C615 a_n3106_n452.t34 gnd 0.10001f
C616 a_n3106_n452.t43 gnd 0.10001f
C617 a_n3106_n452.n7 gnd 0.816794f
C618 a_n3106_n452.n8 gnd 0.411618f
C619 a_n3106_n452.t4 gnd 0.10001f
C620 a_n3106_n452.t0 gnd 0.10001f
C621 a_n3106_n452.n9 gnd 0.816794f
C622 a_n3106_n452.n10 gnd 0.411618f
C623 a_n3106_n452.t51 gnd 0.10001f
C624 a_n3106_n452.t36 gnd 0.10001f
C625 a_n3106_n452.n11 gnd 0.816794f
C626 a_n3106_n452.n12 gnd 0.411618f
C627 a_n3106_n452.t39 gnd 1.03942f
C628 a_n3106_n452.n13 gnd 0.972974f
C629 a_n3106_n452.t37 gnd 1.29145f
C630 a_n3106_n452.n14 gnd 0.909591f
C631 a_n3106_n452.t30 gnd 1.29145f
C632 a_n3106_n452.n15 gnd 0.909591f
C633 a_n3106_n452.t45 gnd 1.29145f
C634 a_n3106_n452.n16 gnd 0.909591f
C635 a_n3106_n452.t3 gnd 1.29145f
C636 a_n3106_n452.n17 gnd 0.909591f
C637 a_n3106_n452.t35 gnd 1.29145f
C638 a_n3106_n452.n18 gnd 0.909591f
C639 a_n3106_n452.t53 gnd 1.29145f
C640 a_n3106_n452.n19 gnd 0.909591f
C641 a_n3106_n452.t38 gnd 1.29145f
C642 a_n3106_n452.n20 gnd 0.789472f
C643 a_n3106_n452.n21 gnd 0.948419f
C644 a_n3106_n452.t14 gnd 1.03941f
C645 a_n3106_n452.n22 gnd 0.645631f
C646 a_n3106_n452.t11 gnd 0.10001f
C647 a_n3106_n452.t28 gnd 0.10001f
C648 a_n3106_n452.n23 gnd 0.816793f
C649 a_n3106_n452.n24 gnd 0.41162f
C650 a_n3106_n452.t22 gnd 0.10001f
C651 a_n3106_n452.t26 gnd 0.10001f
C652 a_n3106_n452.n25 gnd 0.816793f
C653 a_n3106_n452.n26 gnd 0.41162f
C654 a_n3106_n452.t27 gnd 0.10001f
C655 a_n3106_n452.t15 gnd 0.10001f
C656 a_n3106_n452.n27 gnd 0.816793f
C657 a_n3106_n452.n28 gnd 0.41162f
C658 a_n3106_n452.t16 gnd 0.10001f
C659 a_n3106_n452.t7 gnd 0.10001f
C660 a_n3106_n452.n29 gnd 0.816793f
C661 a_n3106_n452.n30 gnd 0.41162f
C662 a_n3106_n452.t9 gnd 0.10001f
C663 a_n3106_n452.t25 gnd 0.10001f
C664 a_n3106_n452.n31 gnd 0.816793f
C665 a_n3106_n452.n32 gnd 0.41162f
C666 a_n3106_n452.t20 gnd 1.03941f
C667 a_n3106_n452.n33 gnd 0.39295f
C668 a_n3106_n452.t44 gnd 1.03941f
C669 a_n3106_n452.n34 gnd 0.39295f
C670 a_n3106_n452.t49 gnd 0.10001f
C671 a_n3106_n452.t42 gnd 0.10001f
C672 a_n3106_n452.n35 gnd 0.816793f
C673 a_n3106_n452.n36 gnd 0.41162f
C674 a_n3106_n452.t41 gnd 0.10001f
C675 a_n3106_n452.t54 gnd 0.10001f
C676 a_n3106_n452.n37 gnd 0.816793f
C677 a_n3106_n452.n38 gnd 0.41162f
C678 a_n3106_n452.t1 gnd 0.10001f
C679 a_n3106_n452.t31 gnd 0.10001f
C680 a_n3106_n452.n39 gnd 0.816793f
C681 a_n3106_n452.n40 gnd 0.41162f
C682 a_n3106_n452.t32 gnd 0.10001f
C683 a_n3106_n452.t33 gnd 0.10001f
C684 a_n3106_n452.n41 gnd 0.816793f
C685 a_n3106_n452.n42 gnd 0.41162f
C686 a_n3106_n452.t52 gnd 0.10001f
C687 a_n3106_n452.t50 gnd 0.10001f
C688 a_n3106_n452.n43 gnd 0.816793f
C689 a_n3106_n452.n44 gnd 0.41162f
C690 a_n3106_n452.t46 gnd 1.03941f
C691 a_n3106_n452.n45 gnd 0.645631f
C692 a_n3106_n452.n46 gnd 1.05146f
C693 a_n3106_n452.t10 gnd 1.03941f
C694 a_n3106_n452.n47 gnd 0.972978f
C695 a_n3106_n452.t8 gnd 0.10001f
C696 a_n3106_n452.t6 gnd 0.10001f
C697 a_n3106_n452.n48 gnd 0.816794f
C698 a_n3106_n452.n49 gnd 0.411618f
C699 a_n3106_n452.t19 gnd 0.10001f
C700 a_n3106_n452.t24 gnd 0.10001f
C701 a_n3106_n452.n50 gnd 0.816794f
C702 a_n3106_n452.n51 gnd 0.411618f
C703 a_n3106_n452.t17 gnd 0.10001f
C704 a_n3106_n452.t21 gnd 0.10001f
C705 a_n3106_n452.n52 gnd 0.816794f
C706 a_n3106_n452.n53 gnd 0.411618f
C707 a_n3106_n452.t13 gnd 0.10001f
C708 a_n3106_n452.t18 gnd 0.10001f
C709 a_n3106_n452.n54 gnd 0.816794f
C710 a_n3106_n452.n55 gnd 0.411618f
C711 a_n3106_n452.n56 gnd 0.411617f
C712 a_n3106_n452.n57 gnd 0.816796f
C713 a_n3106_n452.t29 gnd 0.10001f
C714 plus.n0 gnd 0.022838f
C715 plus.t20 gnd 0.415311f
C716 plus.t23 gnd 0.384014f
C717 plus.n1 gnd 0.155312f
C718 plus.n2 gnd 0.022838f
C719 plus.t6 gnd 0.384014f
C720 plus.n3 gnd 0.019515f
C721 plus.n4 gnd 0.022838f
C722 plus.t12 gnd 0.384014f
C723 plus.t8 gnd 0.384014f
C724 plus.n5 gnd 0.155312f
C725 plus.n6 gnd 0.022838f
C726 plus.t7 gnd 0.384014f
C727 plus.n7 gnd 0.155312f
C728 plus.n8 gnd 0.022838f
C729 plus.t19 gnd 0.384014f
C730 plus.n9 gnd 0.018562f
C731 plus.n10 gnd 0.022838f
C732 plus.t18 gnd 0.384014f
C733 plus.t27 gnd 0.384014f
C734 plus.n11 gnd 0.155312f
C735 plus.n12 gnd 0.022838f
C736 plus.t25 gnd 0.384014f
C737 plus.n13 gnd 0.155312f
C738 plus.n14 gnd 0.096921f
C739 plus.t9 gnd 0.384014f
C740 plus.t14 gnd 0.429589f
C741 plus.n15 gnd 0.181575f
C742 plus.n16 gnd 0.177861f
C743 plus.n17 gnd 0.029263f
C744 plus.n18 gnd 0.025844f
C745 plus.n19 gnd 0.022838f
C746 plus.n20 gnd 0.022838f
C747 plus.n21 gnd 0.027291f
C748 plus.n22 gnd 0.019515f
C749 plus.n23 gnd 0.029743f
C750 plus.n24 gnd 0.022838f
C751 plus.n25 gnd 0.022838f
C752 plus.n26 gnd 0.028408f
C753 plus.n27 gnd 0.026698f
C754 plus.n28 gnd 0.155312f
C755 plus.n29 gnd 0.028608f
C756 plus.n30 gnd 0.022838f
C757 plus.n31 gnd 0.022838f
C758 plus.n32 gnd 0.022838f
C759 plus.n33 gnd 0.02938f
C760 plus.n34 gnd 0.155312f
C761 plus.n35 gnd 0.027553f
C762 plus.n36 gnd 0.027553f
C763 plus.n37 gnd 0.022838f
C764 plus.n38 gnd 0.022838f
C765 plus.n39 gnd 0.02938f
C766 plus.n40 gnd 0.018562f
C767 plus.n41 gnd 0.028608f
C768 plus.n42 gnd 0.022838f
C769 plus.n43 gnd 0.022838f
C770 plus.n44 gnd 0.026698f
C771 plus.n45 gnd 0.028408f
C772 plus.n46 gnd 0.155312f
C773 plus.n47 gnd 0.029743f
C774 plus.n48 gnd 0.022838f
C775 plus.n49 gnd 0.022838f
C776 plus.n50 gnd 0.022838f
C777 plus.n51 gnd 0.027291f
C778 plus.n52 gnd 0.155312f
C779 plus.n53 gnd 0.025844f
C780 plus.n54 gnd 0.029263f
C781 plus.n55 gnd 0.022838f
C782 plus.n56 gnd 0.022838f
C783 plus.n57 gnd 0.029793f
C784 plus.n58 gnd 0.0083f
C785 plus.n59 gnd 0.179825f
C786 plus.n60 gnd 0.261661f
C787 plus.n61 gnd 0.022838f
C788 plus.t28 gnd 0.384014f
C789 plus.n62 gnd 0.155312f
C790 plus.n63 gnd 0.022838f
C791 plus.t26 gnd 0.384014f
C792 plus.n64 gnd 0.019515f
C793 plus.n65 gnd 0.022838f
C794 plus.t10 gnd 0.384014f
C795 plus.t15 gnd 0.384014f
C796 plus.n66 gnd 0.155312f
C797 plus.n67 gnd 0.022838f
C798 plus.t13 gnd 0.384014f
C799 plus.n68 gnd 0.155312f
C800 plus.n69 gnd 0.022838f
C801 plus.t17 gnd 0.384014f
C802 plus.n70 gnd 0.018562f
C803 plus.n71 gnd 0.022838f
C804 plus.t16 gnd 0.384014f
C805 plus.t21 gnd 0.384014f
C806 plus.n72 gnd 0.155312f
C807 plus.n73 gnd 0.022838f
C808 plus.t22 gnd 0.384014f
C809 plus.n74 gnd 0.155312f
C810 plus.n75 gnd 0.096921f
C811 plus.t5 gnd 0.384014f
C812 plus.t11 gnd 0.429589f
C813 plus.n76 gnd 0.181575f
C814 plus.n77 gnd 0.177861f
C815 plus.n78 gnd 0.029263f
C816 plus.n79 gnd 0.025844f
C817 plus.n80 gnd 0.022838f
C818 plus.n81 gnd 0.022838f
C819 plus.n82 gnd 0.027291f
C820 plus.n83 gnd 0.019515f
C821 plus.n84 gnd 0.029743f
C822 plus.n85 gnd 0.022838f
C823 plus.n86 gnd 0.022838f
C824 plus.n87 gnd 0.028408f
C825 plus.n88 gnd 0.026698f
C826 plus.n89 gnd 0.155312f
C827 plus.n90 gnd 0.028608f
C828 plus.n91 gnd 0.022838f
C829 plus.n92 gnd 0.022838f
C830 plus.n93 gnd 0.022838f
C831 plus.n94 gnd 0.02938f
C832 plus.n95 gnd 0.155312f
C833 plus.n96 gnd 0.027553f
C834 plus.n97 gnd 0.027553f
C835 plus.n98 gnd 0.022838f
C836 plus.n99 gnd 0.022838f
C837 plus.n100 gnd 0.02938f
C838 plus.n101 gnd 0.018562f
C839 plus.n102 gnd 0.028608f
C840 plus.n103 gnd 0.022838f
C841 plus.n104 gnd 0.022838f
C842 plus.n105 gnd 0.026698f
C843 plus.n106 gnd 0.028408f
C844 plus.n107 gnd 0.155312f
C845 plus.n108 gnd 0.029743f
C846 plus.n109 gnd 0.022838f
C847 plus.n110 gnd 0.022838f
C848 plus.n111 gnd 0.022838f
C849 plus.n112 gnd 0.027291f
C850 plus.n113 gnd 0.155312f
C851 plus.n114 gnd 0.025844f
C852 plus.n115 gnd 0.029263f
C853 plus.n116 gnd 0.022838f
C854 plus.n117 gnd 0.022838f
C855 plus.n118 gnd 0.029793f
C856 plus.n119 gnd 0.0083f
C857 plus.t24 gnd 0.415311f
C858 plus.n120 gnd 0.179825f
C859 plus.n121 gnd 0.823978f
C860 plus.n122 gnd 1.21471f
C861 plus.t1 gnd 0.039425f
C862 plus.t2 gnd 0.00704f
C863 plus.t4 gnd 0.00704f
C864 plus.n123 gnd 0.022833f
C865 plus.n124 gnd 0.177252f
C866 plus.t3 gnd 0.00704f
C867 plus.t0 gnd 0.00704f
C868 plus.n125 gnd 0.022833f
C869 plus.n126 gnd 0.133049f
C870 plus.n127 gnd 3.03081f
C871 commonsourceibias.n0 gnd 0.010705f
C872 commonsourceibias.t118 gnd 0.162096f
C873 commonsourceibias.t135 gnd 0.149881f
C874 commonsourceibias.n1 gnd 0.007808f
C875 commonsourceibias.n2 gnd 0.008022f
C876 commonsourceibias.t92 gnd 0.149881f
C877 commonsourceibias.n3 gnd 0.010321f
C878 commonsourceibias.n4 gnd 0.008022f
C879 commonsourceibias.t90 gnd 0.149881f
C880 commonsourceibias.n5 gnd 0.059802f
C881 commonsourceibias.t127 gnd 0.149881f
C882 commonsourceibias.n6 gnd 0.007564f
C883 commonsourceibias.n7 gnd 0.008022f
C884 commonsourceibias.t143 gnd 0.149881f
C885 commonsourceibias.n8 gnd 0.010168f
C886 commonsourceibias.n9 gnd 0.008022f
C887 commonsourceibias.t84 gnd 0.149881f
C888 commonsourceibias.n10 gnd 0.059802f
C889 commonsourceibias.t115 gnd 0.149881f
C890 commonsourceibias.n11 gnd 0.007348f
C891 commonsourceibias.n12 gnd 0.008022f
C892 commonsourceibias.t111 gnd 0.149881f
C893 commonsourceibias.n13 gnd 0.009997f
C894 commonsourceibias.n14 gnd 0.010705f
C895 commonsourceibias.t12 gnd 0.162096f
C896 commonsourceibias.t66 gnd 0.149881f
C897 commonsourceibias.n15 gnd 0.007808f
C898 commonsourceibias.n16 gnd 0.008022f
C899 commonsourceibias.t42 gnd 0.149881f
C900 commonsourceibias.n17 gnd 0.010321f
C901 commonsourceibias.n18 gnd 0.008022f
C902 commonsourceibias.t10 gnd 0.149881f
C903 commonsourceibias.n19 gnd 0.059802f
C904 commonsourceibias.t46 gnd 0.149881f
C905 commonsourceibias.n20 gnd 0.007564f
C906 commonsourceibias.n21 gnd 0.008022f
C907 commonsourceibias.t16 gnd 0.149881f
C908 commonsourceibias.n22 gnd 0.010168f
C909 commonsourceibias.n23 gnd 0.008022f
C910 commonsourceibias.t36 gnd 0.149881f
C911 commonsourceibias.n24 gnd 0.059802f
C912 commonsourceibias.t22 gnd 0.149881f
C913 commonsourceibias.n25 gnd 0.007348f
C914 commonsourceibias.n26 gnd 0.008022f
C915 commonsourceibias.t14 gnd 0.149881f
C916 commonsourceibias.n27 gnd 0.009997f
C917 commonsourceibias.n28 gnd 0.008022f
C918 commonsourceibias.t54 gnd 0.149881f
C919 commonsourceibias.n29 gnd 0.059802f
C920 commonsourceibias.t76 gnd 0.149881f
C921 commonsourceibias.n30 gnd 0.007159f
C922 commonsourceibias.n31 gnd 0.008022f
C923 commonsourceibias.t38 gnd 0.149881f
C924 commonsourceibias.n32 gnd 0.009806f
C925 commonsourceibias.n33 gnd 0.008022f
C926 commonsourceibias.t8 gnd 0.149881f
C927 commonsourceibias.n34 gnd 0.059802f
C928 commonsourceibias.t28 gnd 0.149881f
C929 commonsourceibias.n35 gnd 0.006995f
C930 commonsourceibias.n36 gnd 0.008022f
C931 commonsourceibias.t68 gnd 0.149881f
C932 commonsourceibias.n37 gnd 0.009595f
C933 commonsourceibias.n38 gnd 0.008022f
C934 commonsourceibias.t18 gnd 0.149881f
C935 commonsourceibias.n39 gnd 0.059802f
C936 commonsourceibias.t60 gnd 0.149881f
C937 commonsourceibias.n40 gnd 0.006855f
C938 commonsourceibias.n41 gnd 0.008022f
C939 commonsourceibias.t52 gnd 0.149881f
C940 commonsourceibias.n42 gnd 0.00936f
C941 commonsourceibias.t32 gnd 0.16664f
C942 commonsourceibias.t64 gnd 0.149881f
C943 commonsourceibias.n43 gnd 0.065328f
C944 commonsourceibias.n44 gnd 0.07169f
C945 commonsourceibias.n45 gnd 0.033265f
C946 commonsourceibias.n46 gnd 0.008022f
C947 commonsourceibias.n47 gnd 0.007808f
C948 commonsourceibias.n48 gnd 0.01119f
C949 commonsourceibias.n49 gnd 0.059802f
C950 commonsourceibias.n50 gnd 0.011182f
C951 commonsourceibias.n51 gnd 0.008022f
C952 commonsourceibias.n52 gnd 0.008022f
C953 commonsourceibias.n53 gnd 0.008022f
C954 commonsourceibias.n54 gnd 0.010321f
C955 commonsourceibias.n55 gnd 0.059802f
C956 commonsourceibias.n56 gnd 0.010563f
C957 commonsourceibias.n57 gnd 0.010263f
C958 commonsourceibias.n58 gnd 0.008022f
C959 commonsourceibias.n59 gnd 0.008022f
C960 commonsourceibias.n60 gnd 0.008022f
C961 commonsourceibias.n61 gnd 0.007564f
C962 commonsourceibias.n62 gnd 0.0112f
C963 commonsourceibias.n63 gnd 0.059802f
C964 commonsourceibias.n64 gnd 0.011196f
C965 commonsourceibias.n65 gnd 0.008022f
C966 commonsourceibias.n66 gnd 0.008022f
C967 commonsourceibias.n67 gnd 0.008022f
C968 commonsourceibias.n68 gnd 0.010168f
C969 commonsourceibias.n69 gnd 0.059802f
C970 commonsourceibias.n70 gnd 0.010488f
C971 commonsourceibias.n71 gnd 0.010338f
C972 commonsourceibias.n72 gnd 0.008022f
C973 commonsourceibias.n73 gnd 0.008022f
C974 commonsourceibias.n74 gnd 0.008022f
C975 commonsourceibias.n75 gnd 0.007348f
C976 commonsourceibias.n76 gnd 0.011204f
C977 commonsourceibias.n77 gnd 0.059802f
C978 commonsourceibias.n78 gnd 0.011203f
C979 commonsourceibias.n79 gnd 0.008022f
C980 commonsourceibias.n80 gnd 0.008022f
C981 commonsourceibias.n81 gnd 0.008022f
C982 commonsourceibias.n82 gnd 0.009997f
C983 commonsourceibias.n83 gnd 0.059802f
C984 commonsourceibias.n84 gnd 0.010413f
C985 commonsourceibias.n85 gnd 0.010413f
C986 commonsourceibias.n86 gnd 0.008022f
C987 commonsourceibias.n87 gnd 0.008022f
C988 commonsourceibias.n88 gnd 0.008022f
C989 commonsourceibias.n89 gnd 0.007159f
C990 commonsourceibias.n90 gnd 0.011203f
C991 commonsourceibias.n91 gnd 0.059802f
C992 commonsourceibias.n92 gnd 0.011204f
C993 commonsourceibias.n93 gnd 0.008022f
C994 commonsourceibias.n94 gnd 0.008022f
C995 commonsourceibias.n95 gnd 0.008022f
C996 commonsourceibias.n96 gnd 0.009806f
C997 commonsourceibias.n97 gnd 0.059802f
C998 commonsourceibias.n98 gnd 0.010338f
C999 commonsourceibias.n99 gnd 0.010488f
C1000 commonsourceibias.n100 gnd 0.008022f
C1001 commonsourceibias.n101 gnd 0.008022f
C1002 commonsourceibias.n102 gnd 0.008022f
C1003 commonsourceibias.n103 gnd 0.006995f
C1004 commonsourceibias.n104 gnd 0.011196f
C1005 commonsourceibias.n105 gnd 0.059802f
C1006 commonsourceibias.n106 gnd 0.0112f
C1007 commonsourceibias.n107 gnd 0.008022f
C1008 commonsourceibias.n108 gnd 0.008022f
C1009 commonsourceibias.n109 gnd 0.008022f
C1010 commonsourceibias.n110 gnd 0.009595f
C1011 commonsourceibias.n111 gnd 0.059802f
C1012 commonsourceibias.n112 gnd 0.010263f
C1013 commonsourceibias.n113 gnd 0.010563f
C1014 commonsourceibias.n114 gnd 0.008022f
C1015 commonsourceibias.n115 gnd 0.008022f
C1016 commonsourceibias.n116 gnd 0.008022f
C1017 commonsourceibias.n117 gnd 0.006855f
C1018 commonsourceibias.n118 gnd 0.011182f
C1019 commonsourceibias.n119 gnd 0.059802f
C1020 commonsourceibias.n120 gnd 0.01119f
C1021 commonsourceibias.n121 gnd 0.008022f
C1022 commonsourceibias.n122 gnd 0.008022f
C1023 commonsourceibias.n123 gnd 0.008022f
C1024 commonsourceibias.n124 gnd 0.00936f
C1025 commonsourceibias.n125 gnd 0.059802f
C1026 commonsourceibias.n126 gnd 0.009843f
C1027 commonsourceibias.n127 gnd 0.071758f
C1028 commonsourceibias.n128 gnd 0.079928f
C1029 commonsourceibias.t13 gnd 0.017311f
C1030 commonsourceibias.t67 gnd 0.017311f
C1031 commonsourceibias.n129 gnd 0.152968f
C1032 commonsourceibias.n130 gnd 0.132319f
C1033 commonsourceibias.t43 gnd 0.017311f
C1034 commonsourceibias.t11 gnd 0.017311f
C1035 commonsourceibias.n131 gnd 0.152968f
C1036 commonsourceibias.n132 gnd 0.070264f
C1037 commonsourceibias.t47 gnd 0.017311f
C1038 commonsourceibias.t17 gnd 0.017311f
C1039 commonsourceibias.n133 gnd 0.152968f
C1040 commonsourceibias.n134 gnd 0.070264f
C1041 commonsourceibias.t37 gnd 0.017311f
C1042 commonsourceibias.t23 gnd 0.017311f
C1043 commonsourceibias.n135 gnd 0.152968f
C1044 commonsourceibias.n136 gnd 0.070264f
C1045 commonsourceibias.t15 gnd 0.017311f
C1046 commonsourceibias.t55 gnd 0.017311f
C1047 commonsourceibias.n137 gnd 0.152968f
C1048 commonsourceibias.n138 gnd 0.058702f
C1049 commonsourceibias.t65 gnd 0.017311f
C1050 commonsourceibias.t33 gnd 0.017311f
C1051 commonsourceibias.n139 gnd 0.15348f
C1052 commonsourceibias.t61 gnd 0.017311f
C1053 commonsourceibias.t53 gnd 0.017311f
C1054 commonsourceibias.n140 gnd 0.152968f
C1055 commonsourceibias.n141 gnd 0.142538f
C1056 commonsourceibias.t69 gnd 0.017311f
C1057 commonsourceibias.t19 gnd 0.017311f
C1058 commonsourceibias.n142 gnd 0.152968f
C1059 commonsourceibias.n143 gnd 0.070264f
C1060 commonsourceibias.t9 gnd 0.017311f
C1061 commonsourceibias.t29 gnd 0.017311f
C1062 commonsourceibias.n144 gnd 0.152968f
C1063 commonsourceibias.n145 gnd 0.070264f
C1064 commonsourceibias.t77 gnd 0.017311f
C1065 commonsourceibias.t39 gnd 0.017311f
C1066 commonsourceibias.n146 gnd 0.152968f
C1067 commonsourceibias.n147 gnd 0.058702f
C1068 commonsourceibias.n148 gnd 0.071082f
C1069 commonsourceibias.n149 gnd 0.05192f
C1070 commonsourceibias.t131 gnd 0.149881f
C1071 commonsourceibias.n150 gnd 0.059802f
C1072 commonsourceibias.t106 gnd 0.149881f
C1073 commonsourceibias.n151 gnd 0.059802f
C1074 commonsourceibias.n152 gnd 0.008022f
C1075 commonsourceibias.t103 gnd 0.149881f
C1076 commonsourceibias.n153 gnd 0.059802f
C1077 commonsourceibias.n154 gnd 0.008022f
C1078 commonsourceibias.t121 gnd 0.149881f
C1079 commonsourceibias.n155 gnd 0.059802f
C1080 commonsourceibias.n156 gnd 0.008022f
C1081 commonsourceibias.t138 gnd 0.149881f
C1082 commonsourceibias.n157 gnd 0.006995f
C1083 commonsourceibias.n158 gnd 0.008022f
C1084 commonsourceibias.t95 gnd 0.149881f
C1085 commonsourceibias.n159 gnd 0.009595f
C1086 commonsourceibias.n160 gnd 0.008022f
C1087 commonsourceibias.t110 gnd 0.149881f
C1088 commonsourceibias.n161 gnd 0.059802f
C1089 commonsourceibias.t130 gnd 0.149881f
C1090 commonsourceibias.n162 gnd 0.006855f
C1091 commonsourceibias.n163 gnd 0.008022f
C1092 commonsourceibias.t87 gnd 0.149881f
C1093 commonsourceibias.n164 gnd 0.00936f
C1094 commonsourceibias.t117 gnd 0.16664f
C1095 commonsourceibias.t83 gnd 0.149881f
C1096 commonsourceibias.n165 gnd 0.065328f
C1097 commonsourceibias.n166 gnd 0.07169f
C1098 commonsourceibias.n167 gnd 0.033265f
C1099 commonsourceibias.n168 gnd 0.008022f
C1100 commonsourceibias.n169 gnd 0.007808f
C1101 commonsourceibias.n170 gnd 0.01119f
C1102 commonsourceibias.n171 gnd 0.059802f
C1103 commonsourceibias.n172 gnd 0.011182f
C1104 commonsourceibias.n173 gnd 0.008022f
C1105 commonsourceibias.n174 gnd 0.008022f
C1106 commonsourceibias.n175 gnd 0.008022f
C1107 commonsourceibias.n176 gnd 0.010321f
C1108 commonsourceibias.n177 gnd 0.059802f
C1109 commonsourceibias.n178 gnd 0.010563f
C1110 commonsourceibias.n179 gnd 0.010263f
C1111 commonsourceibias.n180 gnd 0.008022f
C1112 commonsourceibias.n181 gnd 0.008022f
C1113 commonsourceibias.n182 gnd 0.008022f
C1114 commonsourceibias.n183 gnd 0.007564f
C1115 commonsourceibias.n184 gnd 0.0112f
C1116 commonsourceibias.n185 gnd 0.059802f
C1117 commonsourceibias.n186 gnd 0.011196f
C1118 commonsourceibias.n187 gnd 0.008022f
C1119 commonsourceibias.n188 gnd 0.008022f
C1120 commonsourceibias.n189 gnd 0.008022f
C1121 commonsourceibias.n190 gnd 0.010168f
C1122 commonsourceibias.n191 gnd 0.059802f
C1123 commonsourceibias.n192 gnd 0.010488f
C1124 commonsourceibias.n193 gnd 0.010338f
C1125 commonsourceibias.n194 gnd 0.008022f
C1126 commonsourceibias.n195 gnd 0.008022f
C1127 commonsourceibias.n196 gnd 0.009806f
C1128 commonsourceibias.n197 gnd 0.007348f
C1129 commonsourceibias.n198 gnd 0.011204f
C1130 commonsourceibias.n199 gnd 0.008022f
C1131 commonsourceibias.n200 gnd 0.008022f
C1132 commonsourceibias.n201 gnd 0.011203f
C1133 commonsourceibias.n202 gnd 0.007159f
C1134 commonsourceibias.n203 gnd 0.009997f
C1135 commonsourceibias.n204 gnd 0.008022f
C1136 commonsourceibias.n205 gnd 0.007008f
C1137 commonsourceibias.n206 gnd 0.010413f
C1138 commonsourceibias.n207 gnd 0.010413f
C1139 commonsourceibias.n208 gnd 0.007008f
C1140 commonsourceibias.n209 gnd 0.008022f
C1141 commonsourceibias.n210 gnd 0.008022f
C1142 commonsourceibias.n211 gnd 0.007159f
C1143 commonsourceibias.n212 gnd 0.011203f
C1144 commonsourceibias.n213 gnd 0.059802f
C1145 commonsourceibias.n214 gnd 0.011204f
C1146 commonsourceibias.n215 gnd 0.008022f
C1147 commonsourceibias.n216 gnd 0.008022f
C1148 commonsourceibias.n217 gnd 0.008022f
C1149 commonsourceibias.n218 gnd 0.009806f
C1150 commonsourceibias.n219 gnd 0.059802f
C1151 commonsourceibias.n220 gnd 0.010338f
C1152 commonsourceibias.n221 gnd 0.010488f
C1153 commonsourceibias.n222 gnd 0.008022f
C1154 commonsourceibias.n223 gnd 0.008022f
C1155 commonsourceibias.n224 gnd 0.008022f
C1156 commonsourceibias.n225 gnd 0.006995f
C1157 commonsourceibias.n226 gnd 0.011196f
C1158 commonsourceibias.n227 gnd 0.059802f
C1159 commonsourceibias.n228 gnd 0.0112f
C1160 commonsourceibias.n229 gnd 0.008022f
C1161 commonsourceibias.n230 gnd 0.008022f
C1162 commonsourceibias.n231 gnd 0.008022f
C1163 commonsourceibias.n232 gnd 0.009595f
C1164 commonsourceibias.n233 gnd 0.059802f
C1165 commonsourceibias.n234 gnd 0.010263f
C1166 commonsourceibias.n235 gnd 0.010563f
C1167 commonsourceibias.n236 gnd 0.008022f
C1168 commonsourceibias.n237 gnd 0.008022f
C1169 commonsourceibias.n238 gnd 0.008022f
C1170 commonsourceibias.n239 gnd 0.006855f
C1171 commonsourceibias.n240 gnd 0.011182f
C1172 commonsourceibias.n241 gnd 0.059802f
C1173 commonsourceibias.n242 gnd 0.01119f
C1174 commonsourceibias.n243 gnd 0.008022f
C1175 commonsourceibias.n244 gnd 0.008022f
C1176 commonsourceibias.n245 gnd 0.008022f
C1177 commonsourceibias.n246 gnd 0.00936f
C1178 commonsourceibias.n247 gnd 0.059802f
C1179 commonsourceibias.n248 gnd 0.009843f
C1180 commonsourceibias.n249 gnd 0.071758f
C1181 commonsourceibias.n250 gnd 0.046883f
C1182 commonsourceibias.n251 gnd 0.010705f
C1183 commonsourceibias.t120 gnd 0.149881f
C1184 commonsourceibias.n252 gnd 0.007808f
C1185 commonsourceibias.n253 gnd 0.008022f
C1186 commonsourceibias.t81 gnd 0.149881f
C1187 commonsourceibias.n254 gnd 0.010321f
C1188 commonsourceibias.n255 gnd 0.008022f
C1189 commonsourceibias.t159 gnd 0.149881f
C1190 commonsourceibias.n256 gnd 0.059802f
C1191 commonsourceibias.t109 gnd 0.149881f
C1192 commonsourceibias.n257 gnd 0.007564f
C1193 commonsourceibias.n258 gnd 0.008022f
C1194 commonsourceibias.t129 gnd 0.149881f
C1195 commonsourceibias.n259 gnd 0.010168f
C1196 commonsourceibias.n260 gnd 0.008022f
C1197 commonsourceibias.t151 gnd 0.149881f
C1198 commonsourceibias.n261 gnd 0.059802f
C1199 commonsourceibias.t100 gnd 0.149881f
C1200 commonsourceibias.n262 gnd 0.007348f
C1201 commonsourceibias.n263 gnd 0.008022f
C1202 commonsourceibias.t96 gnd 0.149881f
C1203 commonsourceibias.n264 gnd 0.009997f
C1204 commonsourceibias.n265 gnd 0.008022f
C1205 commonsourceibias.t113 gnd 0.149881f
C1206 commonsourceibias.n266 gnd 0.059802f
C1207 commonsourceibias.t94 gnd 0.149881f
C1208 commonsourceibias.n267 gnd 0.007159f
C1209 commonsourceibias.n268 gnd 0.008022f
C1210 commonsourceibias.t91 gnd 0.149881f
C1211 commonsourceibias.n269 gnd 0.009806f
C1212 commonsourceibias.n270 gnd 0.008022f
C1213 commonsourceibias.t104 gnd 0.149881f
C1214 commonsourceibias.n271 gnd 0.059802f
C1215 commonsourceibias.t122 gnd 0.149881f
C1216 commonsourceibias.n272 gnd 0.006995f
C1217 commonsourceibias.n273 gnd 0.008022f
C1218 commonsourceibias.t85 gnd 0.149881f
C1219 commonsourceibias.n274 gnd 0.009595f
C1220 commonsourceibias.n275 gnd 0.008022f
C1221 commonsourceibias.t97 gnd 0.149881f
C1222 commonsourceibias.n276 gnd 0.059802f
C1223 commonsourceibias.t112 gnd 0.149881f
C1224 commonsourceibias.n277 gnd 0.006855f
C1225 commonsourceibias.n278 gnd 0.008022f
C1226 commonsourceibias.t155 gnd 0.149881f
C1227 commonsourceibias.n279 gnd 0.00936f
C1228 commonsourceibias.t101 gnd 0.16664f
C1229 commonsourceibias.t152 gnd 0.149881f
C1230 commonsourceibias.n280 gnd 0.065328f
C1231 commonsourceibias.n281 gnd 0.07169f
C1232 commonsourceibias.n282 gnd 0.033265f
C1233 commonsourceibias.n283 gnd 0.008022f
C1234 commonsourceibias.n284 gnd 0.007808f
C1235 commonsourceibias.n285 gnd 0.01119f
C1236 commonsourceibias.n286 gnd 0.059802f
C1237 commonsourceibias.n287 gnd 0.011182f
C1238 commonsourceibias.n288 gnd 0.008022f
C1239 commonsourceibias.n289 gnd 0.008022f
C1240 commonsourceibias.n290 gnd 0.008022f
C1241 commonsourceibias.n291 gnd 0.010321f
C1242 commonsourceibias.n292 gnd 0.059802f
C1243 commonsourceibias.n293 gnd 0.010563f
C1244 commonsourceibias.n294 gnd 0.010263f
C1245 commonsourceibias.n295 gnd 0.008022f
C1246 commonsourceibias.n296 gnd 0.008022f
C1247 commonsourceibias.n297 gnd 0.008022f
C1248 commonsourceibias.n298 gnd 0.007564f
C1249 commonsourceibias.n299 gnd 0.0112f
C1250 commonsourceibias.n300 gnd 0.059802f
C1251 commonsourceibias.n301 gnd 0.011196f
C1252 commonsourceibias.n302 gnd 0.008022f
C1253 commonsourceibias.n303 gnd 0.008022f
C1254 commonsourceibias.n304 gnd 0.008022f
C1255 commonsourceibias.n305 gnd 0.010168f
C1256 commonsourceibias.n306 gnd 0.059802f
C1257 commonsourceibias.n307 gnd 0.010488f
C1258 commonsourceibias.n308 gnd 0.010338f
C1259 commonsourceibias.n309 gnd 0.008022f
C1260 commonsourceibias.n310 gnd 0.008022f
C1261 commonsourceibias.n311 gnd 0.008022f
C1262 commonsourceibias.n312 gnd 0.007348f
C1263 commonsourceibias.n313 gnd 0.011204f
C1264 commonsourceibias.n314 gnd 0.059802f
C1265 commonsourceibias.n315 gnd 0.011203f
C1266 commonsourceibias.n316 gnd 0.008022f
C1267 commonsourceibias.n317 gnd 0.008022f
C1268 commonsourceibias.n318 gnd 0.008022f
C1269 commonsourceibias.n319 gnd 0.009997f
C1270 commonsourceibias.n320 gnd 0.059802f
C1271 commonsourceibias.n321 gnd 0.010413f
C1272 commonsourceibias.n322 gnd 0.010413f
C1273 commonsourceibias.n323 gnd 0.008022f
C1274 commonsourceibias.n324 gnd 0.008022f
C1275 commonsourceibias.n325 gnd 0.008022f
C1276 commonsourceibias.n326 gnd 0.007159f
C1277 commonsourceibias.n327 gnd 0.011203f
C1278 commonsourceibias.n328 gnd 0.059802f
C1279 commonsourceibias.n329 gnd 0.011204f
C1280 commonsourceibias.n330 gnd 0.008022f
C1281 commonsourceibias.n331 gnd 0.008022f
C1282 commonsourceibias.n332 gnd 0.008022f
C1283 commonsourceibias.n333 gnd 0.009806f
C1284 commonsourceibias.n334 gnd 0.059802f
C1285 commonsourceibias.n335 gnd 0.010338f
C1286 commonsourceibias.n336 gnd 0.010488f
C1287 commonsourceibias.n337 gnd 0.008022f
C1288 commonsourceibias.n338 gnd 0.008022f
C1289 commonsourceibias.n339 gnd 0.008022f
C1290 commonsourceibias.n340 gnd 0.006995f
C1291 commonsourceibias.n341 gnd 0.011196f
C1292 commonsourceibias.n342 gnd 0.059802f
C1293 commonsourceibias.n343 gnd 0.0112f
C1294 commonsourceibias.n344 gnd 0.008022f
C1295 commonsourceibias.n345 gnd 0.008022f
C1296 commonsourceibias.n346 gnd 0.008022f
C1297 commonsourceibias.n347 gnd 0.009595f
C1298 commonsourceibias.n348 gnd 0.059802f
C1299 commonsourceibias.n349 gnd 0.010263f
C1300 commonsourceibias.n350 gnd 0.010563f
C1301 commonsourceibias.n351 gnd 0.008022f
C1302 commonsourceibias.n352 gnd 0.008022f
C1303 commonsourceibias.n353 gnd 0.008022f
C1304 commonsourceibias.n354 gnd 0.006855f
C1305 commonsourceibias.n355 gnd 0.011182f
C1306 commonsourceibias.n356 gnd 0.059802f
C1307 commonsourceibias.n357 gnd 0.01119f
C1308 commonsourceibias.n358 gnd 0.008022f
C1309 commonsourceibias.n359 gnd 0.008022f
C1310 commonsourceibias.n360 gnd 0.008022f
C1311 commonsourceibias.n361 gnd 0.00936f
C1312 commonsourceibias.n362 gnd 0.059802f
C1313 commonsourceibias.n363 gnd 0.009843f
C1314 commonsourceibias.t102 gnd 0.162096f
C1315 commonsourceibias.n364 gnd 0.071758f
C1316 commonsourceibias.n365 gnd 0.024957f
C1317 commonsourceibias.n366 gnd 0.404135f
C1318 commonsourceibias.n367 gnd 0.010705f
C1319 commonsourceibias.t139 gnd 0.162096f
C1320 commonsourceibias.t153 gnd 0.149881f
C1321 commonsourceibias.n368 gnd 0.007808f
C1322 commonsourceibias.n369 gnd 0.008022f
C1323 commonsourceibias.t86 gnd 0.149881f
C1324 commonsourceibias.n370 gnd 0.010321f
C1325 commonsourceibias.n371 gnd 0.008022f
C1326 commonsourceibias.t146 gnd 0.149881f
C1327 commonsourceibias.n372 gnd 0.007564f
C1328 commonsourceibias.n373 gnd 0.008022f
C1329 commonsourceibias.t80 gnd 0.149881f
C1330 commonsourceibias.n374 gnd 0.010168f
C1331 commonsourceibias.n375 gnd 0.008022f
C1332 commonsourceibias.t140 gnd 0.149881f
C1333 commonsourceibias.n376 gnd 0.007348f
C1334 commonsourceibias.n377 gnd 0.008022f
C1335 commonsourceibias.t133 gnd 0.149881f
C1336 commonsourceibias.n378 gnd 0.009997f
C1337 commonsourceibias.t1 gnd 0.017311f
C1338 commonsourceibias.t21 gnd 0.017311f
C1339 commonsourceibias.n379 gnd 0.15348f
C1340 commonsourceibias.t45 gnd 0.017311f
C1341 commonsourceibias.t7 gnd 0.017311f
C1342 commonsourceibias.n380 gnd 0.152968f
C1343 commonsourceibias.n381 gnd 0.142538f
C1344 commonsourceibias.t35 gnd 0.017311f
C1345 commonsourceibias.t27 gnd 0.017311f
C1346 commonsourceibias.n382 gnd 0.152968f
C1347 commonsourceibias.n383 gnd 0.070264f
C1348 commonsourceibias.t73 gnd 0.017311f
C1349 commonsourceibias.t41 gnd 0.017311f
C1350 commonsourceibias.n384 gnd 0.152968f
C1351 commonsourceibias.n385 gnd 0.070264f
C1352 commonsourceibias.t5 gnd 0.017311f
C1353 commonsourceibias.t75 gnd 0.017311f
C1354 commonsourceibias.n386 gnd 0.152968f
C1355 commonsourceibias.n387 gnd 0.058702f
C1356 commonsourceibias.n388 gnd 0.010705f
C1357 commonsourceibias.t48 gnd 0.149881f
C1358 commonsourceibias.n389 gnd 0.007808f
C1359 commonsourceibias.n390 gnd 0.008022f
C1360 commonsourceibias.t30 gnd 0.149881f
C1361 commonsourceibias.n391 gnd 0.010321f
C1362 commonsourceibias.n392 gnd 0.008022f
C1363 commonsourceibias.t24 gnd 0.149881f
C1364 commonsourceibias.n393 gnd 0.007564f
C1365 commonsourceibias.n394 gnd 0.008022f
C1366 commonsourceibias.t70 gnd 0.149881f
C1367 commonsourceibias.n395 gnd 0.010168f
C1368 commonsourceibias.n396 gnd 0.008022f
C1369 commonsourceibias.t78 gnd 0.149881f
C1370 commonsourceibias.n397 gnd 0.007348f
C1371 commonsourceibias.n398 gnd 0.008022f
C1372 commonsourceibias.t62 gnd 0.149881f
C1373 commonsourceibias.n399 gnd 0.009997f
C1374 commonsourceibias.n400 gnd 0.008022f
C1375 commonsourceibias.t74 gnd 0.149881f
C1376 commonsourceibias.n401 gnd 0.007159f
C1377 commonsourceibias.n402 gnd 0.008022f
C1378 commonsourceibias.t4 gnd 0.149881f
C1379 commonsourceibias.n403 gnd 0.009806f
C1380 commonsourceibias.n404 gnd 0.008022f
C1381 commonsourceibias.t72 gnd 0.149881f
C1382 commonsourceibias.n405 gnd 0.006995f
C1383 commonsourceibias.n406 gnd 0.008022f
C1384 commonsourceibias.t26 gnd 0.149881f
C1385 commonsourceibias.n407 gnd 0.009595f
C1386 commonsourceibias.n408 gnd 0.008022f
C1387 commonsourceibias.t6 gnd 0.149881f
C1388 commonsourceibias.n409 gnd 0.006855f
C1389 commonsourceibias.n410 gnd 0.008022f
C1390 commonsourceibias.t44 gnd 0.149881f
C1391 commonsourceibias.n411 gnd 0.00936f
C1392 commonsourceibias.t0 gnd 0.16664f
C1393 commonsourceibias.t20 gnd 0.149881f
C1394 commonsourceibias.n412 gnd 0.065328f
C1395 commonsourceibias.n413 gnd 0.07169f
C1396 commonsourceibias.n414 gnd 0.033265f
C1397 commonsourceibias.n415 gnd 0.008022f
C1398 commonsourceibias.n416 gnd 0.007808f
C1399 commonsourceibias.n417 gnd 0.01119f
C1400 commonsourceibias.n418 gnd 0.059802f
C1401 commonsourceibias.n419 gnd 0.011182f
C1402 commonsourceibias.n420 gnd 0.008022f
C1403 commonsourceibias.n421 gnd 0.008022f
C1404 commonsourceibias.n422 gnd 0.008022f
C1405 commonsourceibias.n423 gnd 0.010321f
C1406 commonsourceibias.n424 gnd 0.059802f
C1407 commonsourceibias.n425 gnd 0.010563f
C1408 commonsourceibias.t34 gnd 0.149881f
C1409 commonsourceibias.n426 gnd 0.059802f
C1410 commonsourceibias.n427 gnd 0.010263f
C1411 commonsourceibias.n428 gnd 0.008022f
C1412 commonsourceibias.n429 gnd 0.008022f
C1413 commonsourceibias.n430 gnd 0.008022f
C1414 commonsourceibias.n431 gnd 0.007564f
C1415 commonsourceibias.n432 gnd 0.0112f
C1416 commonsourceibias.n433 gnd 0.059802f
C1417 commonsourceibias.n434 gnd 0.011196f
C1418 commonsourceibias.n435 gnd 0.008022f
C1419 commonsourceibias.n436 gnd 0.008022f
C1420 commonsourceibias.n437 gnd 0.008022f
C1421 commonsourceibias.n438 gnd 0.010168f
C1422 commonsourceibias.n439 gnd 0.059802f
C1423 commonsourceibias.n440 gnd 0.010488f
C1424 commonsourceibias.t40 gnd 0.149881f
C1425 commonsourceibias.n441 gnd 0.059802f
C1426 commonsourceibias.n442 gnd 0.010338f
C1427 commonsourceibias.n443 gnd 0.008022f
C1428 commonsourceibias.n444 gnd 0.008022f
C1429 commonsourceibias.n445 gnd 0.008022f
C1430 commonsourceibias.n446 gnd 0.007348f
C1431 commonsourceibias.n447 gnd 0.011204f
C1432 commonsourceibias.n448 gnd 0.059802f
C1433 commonsourceibias.n449 gnd 0.011203f
C1434 commonsourceibias.n450 gnd 0.008022f
C1435 commonsourceibias.n451 gnd 0.008022f
C1436 commonsourceibias.n452 gnd 0.008022f
C1437 commonsourceibias.n453 gnd 0.009997f
C1438 commonsourceibias.n454 gnd 0.059802f
C1439 commonsourceibias.n455 gnd 0.010413f
C1440 commonsourceibias.t2 gnd 0.149881f
C1441 commonsourceibias.n456 gnd 0.059802f
C1442 commonsourceibias.n457 gnd 0.010413f
C1443 commonsourceibias.n458 gnd 0.008022f
C1444 commonsourceibias.n459 gnd 0.008022f
C1445 commonsourceibias.n460 gnd 0.008022f
C1446 commonsourceibias.n461 gnd 0.007159f
C1447 commonsourceibias.n462 gnd 0.011203f
C1448 commonsourceibias.n463 gnd 0.059802f
C1449 commonsourceibias.n464 gnd 0.011204f
C1450 commonsourceibias.n465 gnd 0.008022f
C1451 commonsourceibias.n466 gnd 0.008022f
C1452 commonsourceibias.n467 gnd 0.008022f
C1453 commonsourceibias.n468 gnd 0.009806f
C1454 commonsourceibias.n469 gnd 0.059802f
C1455 commonsourceibias.n470 gnd 0.010338f
C1456 commonsourceibias.t50 gnd 0.149881f
C1457 commonsourceibias.n471 gnd 0.059802f
C1458 commonsourceibias.n472 gnd 0.010488f
C1459 commonsourceibias.n473 gnd 0.008022f
C1460 commonsourceibias.n474 gnd 0.008022f
C1461 commonsourceibias.n475 gnd 0.008022f
C1462 commonsourceibias.n476 gnd 0.006995f
C1463 commonsourceibias.n477 gnd 0.011196f
C1464 commonsourceibias.n478 gnd 0.059802f
C1465 commonsourceibias.n479 gnd 0.0112f
C1466 commonsourceibias.n480 gnd 0.008022f
C1467 commonsourceibias.n481 gnd 0.008022f
C1468 commonsourceibias.n482 gnd 0.008022f
C1469 commonsourceibias.n483 gnd 0.009595f
C1470 commonsourceibias.n484 gnd 0.059802f
C1471 commonsourceibias.n485 gnd 0.010263f
C1472 commonsourceibias.t56 gnd 0.149881f
C1473 commonsourceibias.n486 gnd 0.059802f
C1474 commonsourceibias.n487 gnd 0.010563f
C1475 commonsourceibias.n488 gnd 0.008022f
C1476 commonsourceibias.n489 gnd 0.008022f
C1477 commonsourceibias.n490 gnd 0.008022f
C1478 commonsourceibias.n491 gnd 0.006855f
C1479 commonsourceibias.n492 gnd 0.011182f
C1480 commonsourceibias.n493 gnd 0.059802f
C1481 commonsourceibias.n494 gnd 0.01119f
C1482 commonsourceibias.n495 gnd 0.008022f
C1483 commonsourceibias.n496 gnd 0.008022f
C1484 commonsourceibias.n497 gnd 0.008022f
C1485 commonsourceibias.n498 gnd 0.00936f
C1486 commonsourceibias.n499 gnd 0.059802f
C1487 commonsourceibias.n500 gnd 0.009843f
C1488 commonsourceibias.t58 gnd 0.162096f
C1489 commonsourceibias.n501 gnd 0.071758f
C1490 commonsourceibias.n502 gnd 0.079928f
C1491 commonsourceibias.t49 gnd 0.017311f
C1492 commonsourceibias.t59 gnd 0.017311f
C1493 commonsourceibias.n503 gnd 0.152968f
C1494 commonsourceibias.n504 gnd 0.132319f
C1495 commonsourceibias.t57 gnd 0.017311f
C1496 commonsourceibias.t31 gnd 0.017311f
C1497 commonsourceibias.n505 gnd 0.152968f
C1498 commonsourceibias.n506 gnd 0.070264f
C1499 commonsourceibias.t71 gnd 0.017311f
C1500 commonsourceibias.t25 gnd 0.017311f
C1501 commonsourceibias.n507 gnd 0.152968f
C1502 commonsourceibias.n508 gnd 0.070264f
C1503 commonsourceibias.t79 gnd 0.017311f
C1504 commonsourceibias.t51 gnd 0.017311f
C1505 commonsourceibias.n509 gnd 0.152968f
C1506 commonsourceibias.n510 gnd 0.070264f
C1507 commonsourceibias.t3 gnd 0.017311f
C1508 commonsourceibias.t63 gnd 0.017311f
C1509 commonsourceibias.n511 gnd 0.152968f
C1510 commonsourceibias.n512 gnd 0.058702f
C1511 commonsourceibias.n513 gnd 0.071082f
C1512 commonsourceibias.n514 gnd 0.05192f
C1513 commonsourceibias.t98 gnd 0.149881f
C1514 commonsourceibias.n515 gnd 0.059802f
C1515 commonsourceibias.n516 gnd 0.008022f
C1516 commonsourceibias.t126 gnd 0.149881f
C1517 commonsourceibias.n517 gnd 0.059802f
C1518 commonsourceibias.n518 gnd 0.008022f
C1519 commonsourceibias.t142 gnd 0.149881f
C1520 commonsourceibias.n519 gnd 0.059802f
C1521 commonsourceibias.n520 gnd 0.008022f
C1522 commonsourceibias.t156 gnd 0.149881f
C1523 commonsourceibias.n521 gnd 0.006995f
C1524 commonsourceibias.n522 gnd 0.008022f
C1525 commonsourceibias.t114 gnd 0.149881f
C1526 commonsourceibias.n523 gnd 0.009595f
C1527 commonsourceibias.n524 gnd 0.008022f
C1528 commonsourceibias.t148 gnd 0.149881f
C1529 commonsourceibias.n525 gnd 0.006855f
C1530 commonsourceibias.n526 gnd 0.008022f
C1531 commonsourceibias.t82 gnd 0.149881f
C1532 commonsourceibias.n527 gnd 0.00936f
C1533 commonsourceibias.t125 gnd 0.16664f
C1534 commonsourceibias.t89 gnd 0.149881f
C1535 commonsourceibias.n528 gnd 0.065328f
C1536 commonsourceibias.n529 gnd 0.07169f
C1537 commonsourceibias.n530 gnd 0.033265f
C1538 commonsourceibias.n531 gnd 0.008022f
C1539 commonsourceibias.n532 gnd 0.007808f
C1540 commonsourceibias.n533 gnd 0.01119f
C1541 commonsourceibias.n534 gnd 0.059802f
C1542 commonsourceibias.n535 gnd 0.011182f
C1543 commonsourceibias.n536 gnd 0.008022f
C1544 commonsourceibias.n537 gnd 0.008022f
C1545 commonsourceibias.n538 gnd 0.008022f
C1546 commonsourceibias.n539 gnd 0.010321f
C1547 commonsourceibias.n540 gnd 0.059802f
C1548 commonsourceibias.n541 gnd 0.010563f
C1549 commonsourceibias.t134 gnd 0.149881f
C1550 commonsourceibias.n542 gnd 0.059802f
C1551 commonsourceibias.n543 gnd 0.010263f
C1552 commonsourceibias.n544 gnd 0.008022f
C1553 commonsourceibias.n545 gnd 0.008022f
C1554 commonsourceibias.n546 gnd 0.008022f
C1555 commonsourceibias.n547 gnd 0.007564f
C1556 commonsourceibias.n548 gnd 0.0112f
C1557 commonsourceibias.n549 gnd 0.059802f
C1558 commonsourceibias.n550 gnd 0.011196f
C1559 commonsourceibias.n551 gnd 0.008022f
C1560 commonsourceibias.n552 gnd 0.008022f
C1561 commonsourceibias.n553 gnd 0.008022f
C1562 commonsourceibias.n554 gnd 0.010168f
C1563 commonsourceibias.n555 gnd 0.059802f
C1564 commonsourceibias.n556 gnd 0.010488f
C1565 commonsourceibias.n557 gnd 0.010338f
C1566 commonsourceibias.n558 gnd 0.008022f
C1567 commonsourceibias.n559 gnd 0.008022f
C1568 commonsourceibias.n560 gnd 0.009806f
C1569 commonsourceibias.n561 gnd 0.007348f
C1570 commonsourceibias.n562 gnd 0.011204f
C1571 commonsourceibias.n563 gnd 0.008022f
C1572 commonsourceibias.n564 gnd 0.008022f
C1573 commonsourceibias.n565 gnd 0.011203f
C1574 commonsourceibias.n566 gnd 0.007159f
C1575 commonsourceibias.n567 gnd 0.009997f
C1576 commonsourceibias.n568 gnd 0.008022f
C1577 commonsourceibias.n569 gnd 0.007008f
C1578 commonsourceibias.n570 gnd 0.010413f
C1579 commonsourceibias.t149 gnd 0.149881f
C1580 commonsourceibias.n571 gnd 0.059802f
C1581 commonsourceibias.n572 gnd 0.010413f
C1582 commonsourceibias.n573 gnd 0.007008f
C1583 commonsourceibias.n574 gnd 0.008022f
C1584 commonsourceibias.n575 gnd 0.008022f
C1585 commonsourceibias.n576 gnd 0.007159f
C1586 commonsourceibias.n577 gnd 0.011203f
C1587 commonsourceibias.n578 gnd 0.059802f
C1588 commonsourceibias.n579 gnd 0.011204f
C1589 commonsourceibias.n580 gnd 0.008022f
C1590 commonsourceibias.n581 gnd 0.008022f
C1591 commonsourceibias.n582 gnd 0.008022f
C1592 commonsourceibias.n583 gnd 0.009806f
C1593 commonsourceibias.n584 gnd 0.059802f
C1594 commonsourceibias.n585 gnd 0.010338f
C1595 commonsourceibias.t157 gnd 0.149881f
C1596 commonsourceibias.n586 gnd 0.059802f
C1597 commonsourceibias.n587 gnd 0.010488f
C1598 commonsourceibias.n588 gnd 0.008022f
C1599 commonsourceibias.n589 gnd 0.008022f
C1600 commonsourceibias.n590 gnd 0.008022f
C1601 commonsourceibias.n591 gnd 0.006995f
C1602 commonsourceibias.n592 gnd 0.011196f
C1603 commonsourceibias.n593 gnd 0.059802f
C1604 commonsourceibias.n594 gnd 0.0112f
C1605 commonsourceibias.n595 gnd 0.008022f
C1606 commonsourceibias.n596 gnd 0.008022f
C1607 commonsourceibias.n597 gnd 0.008022f
C1608 commonsourceibias.n598 gnd 0.009595f
C1609 commonsourceibias.n599 gnd 0.059802f
C1610 commonsourceibias.n600 gnd 0.010263f
C1611 commonsourceibias.t105 gnd 0.149881f
C1612 commonsourceibias.n601 gnd 0.059802f
C1613 commonsourceibias.n602 gnd 0.010563f
C1614 commonsourceibias.n603 gnd 0.008022f
C1615 commonsourceibias.n604 gnd 0.008022f
C1616 commonsourceibias.n605 gnd 0.008022f
C1617 commonsourceibias.n606 gnd 0.006855f
C1618 commonsourceibias.n607 gnd 0.011182f
C1619 commonsourceibias.n608 gnd 0.059802f
C1620 commonsourceibias.n609 gnd 0.01119f
C1621 commonsourceibias.n610 gnd 0.008022f
C1622 commonsourceibias.n611 gnd 0.008022f
C1623 commonsourceibias.n612 gnd 0.008022f
C1624 commonsourceibias.n613 gnd 0.00936f
C1625 commonsourceibias.n614 gnd 0.059802f
C1626 commonsourceibias.n615 gnd 0.009843f
C1627 commonsourceibias.n616 gnd 0.071758f
C1628 commonsourceibias.n617 gnd 0.046883f
C1629 commonsourceibias.n618 gnd 0.010705f
C1630 commonsourceibias.t141 gnd 0.149881f
C1631 commonsourceibias.n619 gnd 0.007808f
C1632 commonsourceibias.n620 gnd 0.008022f
C1633 commonsourceibias.t154 gnd 0.149881f
C1634 commonsourceibias.n621 gnd 0.010321f
C1635 commonsourceibias.n622 gnd 0.008022f
C1636 commonsourceibias.t132 gnd 0.149881f
C1637 commonsourceibias.n623 gnd 0.007564f
C1638 commonsourceibias.n624 gnd 0.008022f
C1639 commonsourceibias.t147 gnd 0.149881f
C1640 commonsourceibias.n625 gnd 0.010168f
C1641 commonsourceibias.n626 gnd 0.008022f
C1642 commonsourceibias.t124 gnd 0.149881f
C1643 commonsourceibias.n627 gnd 0.007348f
C1644 commonsourceibias.n628 gnd 0.008022f
C1645 commonsourceibias.t116 gnd 0.149881f
C1646 commonsourceibias.n629 gnd 0.009997f
C1647 commonsourceibias.n630 gnd 0.008022f
C1648 commonsourceibias.t88 gnd 0.149881f
C1649 commonsourceibias.n631 gnd 0.007159f
C1650 commonsourceibias.n632 gnd 0.008022f
C1651 commonsourceibias.t107 gnd 0.149881f
C1652 commonsourceibias.n633 gnd 0.009806f
C1653 commonsourceibias.n634 gnd 0.008022f
C1654 commonsourceibias.t145 gnd 0.149881f
C1655 commonsourceibias.n635 gnd 0.006995f
C1656 commonsourceibias.n636 gnd 0.008022f
C1657 commonsourceibias.t99 gnd 0.149881f
C1658 commonsourceibias.n637 gnd 0.009595f
C1659 commonsourceibias.n638 gnd 0.008022f
C1660 commonsourceibias.t137 gnd 0.149881f
C1661 commonsourceibias.n639 gnd 0.006855f
C1662 commonsourceibias.n640 gnd 0.008022f
C1663 commonsourceibias.t150 gnd 0.149881f
C1664 commonsourceibias.n641 gnd 0.00936f
C1665 commonsourceibias.t108 gnd 0.16664f
C1666 commonsourceibias.t158 gnd 0.149881f
C1667 commonsourceibias.n642 gnd 0.065328f
C1668 commonsourceibias.n643 gnd 0.07169f
C1669 commonsourceibias.n644 gnd 0.033265f
C1670 commonsourceibias.n645 gnd 0.008022f
C1671 commonsourceibias.n646 gnd 0.007808f
C1672 commonsourceibias.n647 gnd 0.01119f
C1673 commonsourceibias.n648 gnd 0.059802f
C1674 commonsourceibias.n649 gnd 0.011182f
C1675 commonsourceibias.n650 gnd 0.008022f
C1676 commonsourceibias.n651 gnd 0.008022f
C1677 commonsourceibias.n652 gnd 0.008022f
C1678 commonsourceibias.n653 gnd 0.010321f
C1679 commonsourceibias.n654 gnd 0.059802f
C1680 commonsourceibias.n655 gnd 0.010563f
C1681 commonsourceibias.t119 gnd 0.149881f
C1682 commonsourceibias.n656 gnd 0.059802f
C1683 commonsourceibias.n657 gnd 0.010263f
C1684 commonsourceibias.n658 gnd 0.008022f
C1685 commonsourceibias.n659 gnd 0.008022f
C1686 commonsourceibias.n660 gnd 0.008022f
C1687 commonsourceibias.n661 gnd 0.007564f
C1688 commonsourceibias.n662 gnd 0.0112f
C1689 commonsourceibias.n663 gnd 0.059802f
C1690 commonsourceibias.n664 gnd 0.011196f
C1691 commonsourceibias.n665 gnd 0.008022f
C1692 commonsourceibias.n666 gnd 0.008022f
C1693 commonsourceibias.n667 gnd 0.008022f
C1694 commonsourceibias.n668 gnd 0.010168f
C1695 commonsourceibias.n669 gnd 0.059802f
C1696 commonsourceibias.n670 gnd 0.010488f
C1697 commonsourceibias.t128 gnd 0.149881f
C1698 commonsourceibias.n671 gnd 0.059802f
C1699 commonsourceibias.n672 gnd 0.010338f
C1700 commonsourceibias.n673 gnd 0.008022f
C1701 commonsourceibias.n674 gnd 0.008022f
C1702 commonsourceibias.n675 gnd 0.008022f
C1703 commonsourceibias.n676 gnd 0.007348f
C1704 commonsourceibias.n677 gnd 0.011204f
C1705 commonsourceibias.n678 gnd 0.059802f
C1706 commonsourceibias.n679 gnd 0.011203f
C1707 commonsourceibias.n680 gnd 0.008022f
C1708 commonsourceibias.n681 gnd 0.008022f
C1709 commonsourceibias.n682 gnd 0.008022f
C1710 commonsourceibias.n683 gnd 0.009997f
C1711 commonsourceibias.n684 gnd 0.059802f
C1712 commonsourceibias.n685 gnd 0.010413f
C1713 commonsourceibias.t136 gnd 0.149881f
C1714 commonsourceibias.n686 gnd 0.059802f
C1715 commonsourceibias.n687 gnd 0.010413f
C1716 commonsourceibias.n688 gnd 0.008022f
C1717 commonsourceibias.n689 gnd 0.008022f
C1718 commonsourceibias.n690 gnd 0.008022f
C1719 commonsourceibias.n691 gnd 0.007159f
C1720 commonsourceibias.n692 gnd 0.011203f
C1721 commonsourceibias.n693 gnd 0.059802f
C1722 commonsourceibias.n694 gnd 0.011204f
C1723 commonsourceibias.n695 gnd 0.008022f
C1724 commonsourceibias.n696 gnd 0.008022f
C1725 commonsourceibias.n697 gnd 0.008022f
C1726 commonsourceibias.n698 gnd 0.009806f
C1727 commonsourceibias.n699 gnd 0.059802f
C1728 commonsourceibias.n700 gnd 0.010338f
C1729 commonsourceibias.t144 gnd 0.149881f
C1730 commonsourceibias.n701 gnd 0.059802f
C1731 commonsourceibias.n702 gnd 0.010488f
C1732 commonsourceibias.n703 gnd 0.008022f
C1733 commonsourceibias.n704 gnd 0.008022f
C1734 commonsourceibias.n705 gnd 0.008022f
C1735 commonsourceibias.n706 gnd 0.006995f
C1736 commonsourceibias.n707 gnd 0.011196f
C1737 commonsourceibias.n708 gnd 0.059802f
C1738 commonsourceibias.n709 gnd 0.0112f
C1739 commonsourceibias.n710 gnd 0.008022f
C1740 commonsourceibias.n711 gnd 0.008022f
C1741 commonsourceibias.n712 gnd 0.008022f
C1742 commonsourceibias.n713 gnd 0.009595f
C1743 commonsourceibias.n714 gnd 0.059802f
C1744 commonsourceibias.n715 gnd 0.010263f
C1745 commonsourceibias.t93 gnd 0.149881f
C1746 commonsourceibias.n716 gnd 0.059802f
C1747 commonsourceibias.n717 gnd 0.010563f
C1748 commonsourceibias.n718 gnd 0.008022f
C1749 commonsourceibias.n719 gnd 0.008022f
C1750 commonsourceibias.n720 gnd 0.008022f
C1751 commonsourceibias.n721 gnd 0.006855f
C1752 commonsourceibias.n722 gnd 0.011182f
C1753 commonsourceibias.n723 gnd 0.059802f
C1754 commonsourceibias.n724 gnd 0.01119f
C1755 commonsourceibias.n725 gnd 0.008022f
C1756 commonsourceibias.n726 gnd 0.008022f
C1757 commonsourceibias.n727 gnd 0.008022f
C1758 commonsourceibias.n728 gnd 0.00936f
C1759 commonsourceibias.n729 gnd 0.059802f
C1760 commonsourceibias.n730 gnd 0.009843f
C1761 commonsourceibias.t123 gnd 0.162096f
C1762 commonsourceibias.n731 gnd 0.071758f
C1763 commonsourceibias.n732 gnd 0.024957f
C1764 commonsourceibias.n733 gnd 0.221543f
C1765 commonsourceibias.n734 gnd 4.49224f
C1766 CSoutput.n0 gnd 0.03683f
C1767 CSoutput.t146 gnd 0.243625f
C1768 CSoutput.n1 gnd 0.110009f
C1769 CSoutput.n2 gnd 0.03683f
C1770 CSoutput.t144 gnd 0.243625f
C1771 CSoutput.n3 gnd 0.029191f
C1772 CSoutput.n4 gnd 0.03683f
C1773 CSoutput.t137 gnd 0.243625f
C1774 CSoutput.n5 gnd 0.025172f
C1775 CSoutput.n6 gnd 0.03683f
C1776 CSoutput.t141 gnd 0.243625f
C1777 CSoutput.t130 gnd 0.243625f
C1778 CSoutput.n7 gnd 0.10881f
C1779 CSoutput.n8 gnd 0.03683f
C1780 CSoutput.t129 gnd 0.243625f
C1781 CSoutput.n9 gnd 0.024f
C1782 CSoutput.n10 gnd 0.03683f
C1783 CSoutput.t138 gnd 0.243625f
C1784 CSoutput.t143 gnd 0.243625f
C1785 CSoutput.n11 gnd 0.10881f
C1786 CSoutput.n12 gnd 0.03683f
C1787 CSoutput.t149 gnd 0.243625f
C1788 CSoutput.n13 gnd 0.025172f
C1789 CSoutput.n14 gnd 0.03683f
C1790 CSoutput.t131 gnd 0.243625f
C1791 CSoutput.t140 gnd 0.243625f
C1792 CSoutput.n15 gnd 0.10881f
C1793 CSoutput.n16 gnd 0.03683f
C1794 CSoutput.t147 gnd 0.243625f
C1795 CSoutput.n17 gnd 0.026885f
C1796 CSoutput.t134 gnd 0.291138f
C1797 CSoutput.t145 gnd 0.243625f
C1798 CSoutput.n18 gnd 0.138908f
C1799 CSoutput.n19 gnd 0.134789f
C1800 CSoutput.n20 gnd 0.156371f
C1801 CSoutput.n21 gnd 0.03683f
C1802 CSoutput.n22 gnd 0.030739f
C1803 CSoutput.n23 gnd 0.10881f
C1804 CSoutput.n24 gnd 0.029631f
C1805 CSoutput.n25 gnd 0.029191f
C1806 CSoutput.n26 gnd 0.03683f
C1807 CSoutput.n27 gnd 0.03683f
C1808 CSoutput.n28 gnd 0.030503f
C1809 CSoutput.n29 gnd 0.025898f
C1810 CSoutput.n30 gnd 0.111232f
C1811 CSoutput.n31 gnd 0.026254f
C1812 CSoutput.n32 gnd 0.03683f
C1813 CSoutput.n33 gnd 0.03683f
C1814 CSoutput.n34 gnd 0.03683f
C1815 CSoutput.n35 gnd 0.030178f
C1816 CSoutput.n36 gnd 0.10881f
C1817 CSoutput.n37 gnd 0.028861f
C1818 CSoutput.n38 gnd 0.029962f
C1819 CSoutput.n39 gnd 0.03683f
C1820 CSoutput.n40 gnd 0.03683f
C1821 CSoutput.n41 gnd 0.030733f
C1822 CSoutput.n42 gnd 0.02809f
C1823 CSoutput.n43 gnd 0.10881f
C1824 CSoutput.n44 gnd 0.028802f
C1825 CSoutput.n45 gnd 0.03683f
C1826 CSoutput.n46 gnd 0.03683f
C1827 CSoutput.n47 gnd 0.03683f
C1828 CSoutput.n48 gnd 0.028802f
C1829 CSoutput.n49 gnd 0.10881f
C1830 CSoutput.n50 gnd 0.02809f
C1831 CSoutput.n51 gnd 0.030733f
C1832 CSoutput.n52 gnd 0.03683f
C1833 CSoutput.n53 gnd 0.03683f
C1834 CSoutput.n54 gnd 0.029962f
C1835 CSoutput.n55 gnd 0.028861f
C1836 CSoutput.n56 gnd 0.10881f
C1837 CSoutput.n57 gnd 0.030178f
C1838 CSoutput.n58 gnd 0.03683f
C1839 CSoutput.n59 gnd 0.03683f
C1840 CSoutput.n60 gnd 0.03683f
C1841 CSoutput.n61 gnd 0.026254f
C1842 CSoutput.n62 gnd 0.111232f
C1843 CSoutput.n63 gnd 0.025898f
C1844 CSoutput.t133 gnd 0.243625f
C1845 CSoutput.n64 gnd 0.10881f
C1846 CSoutput.n65 gnd 0.030503f
C1847 CSoutput.n66 gnd 0.03683f
C1848 CSoutput.n67 gnd 0.03683f
C1849 CSoutput.n68 gnd 0.03683f
C1850 CSoutput.n69 gnd 0.029631f
C1851 CSoutput.n70 gnd 0.10881f
C1852 CSoutput.n71 gnd 0.030739f
C1853 CSoutput.n72 gnd 0.026885f
C1854 CSoutput.n73 gnd 0.03683f
C1855 CSoutput.n74 gnd 0.03683f
C1856 CSoutput.n75 gnd 0.027881f
C1857 CSoutput.n76 gnd 0.016559f
C1858 CSoutput.t136 gnd 0.27373f
C1859 CSoutput.n77 gnd 0.135978f
C1860 CSoutput.n78 gnd 0.581838f
C1861 CSoutput.t26 gnd 0.045941f
C1862 CSoutput.t51 gnd 0.045941f
C1863 CSoutput.n79 gnd 0.355688f
C1864 CSoutput.t28 gnd 0.045941f
C1865 CSoutput.t41 gnd 0.045941f
C1866 CSoutput.n80 gnd 0.355054f
C1867 CSoutput.n81 gnd 0.360379f
C1868 CSoutput.t70 gnd 0.045941f
C1869 CSoutput.t47 gnd 0.045941f
C1870 CSoutput.n82 gnd 0.355054f
C1871 CSoutput.n83 gnd 0.17758f
C1872 CSoutput.t30 gnd 0.045941f
C1873 CSoutput.t61 gnd 0.045941f
C1874 CSoutput.n84 gnd 0.355054f
C1875 CSoutput.n85 gnd 0.32564f
C1876 CSoutput.t35 gnd 0.045941f
C1877 CSoutput.t66 gnd 0.045941f
C1878 CSoutput.n86 gnd 0.355688f
C1879 CSoutput.t55 gnd 0.045941f
C1880 CSoutput.t54 gnd 0.045941f
C1881 CSoutput.n87 gnd 0.355054f
C1882 CSoutput.n88 gnd 0.360379f
C1883 CSoutput.t50 gnd 0.045941f
C1884 CSoutput.t33 gnd 0.045941f
C1885 CSoutput.n89 gnd 0.355054f
C1886 CSoutput.n90 gnd 0.17758f
C1887 CSoutput.t25 gnd 0.045941f
C1888 CSoutput.t49 gnd 0.045941f
C1889 CSoutput.n91 gnd 0.355054f
C1890 CSoutput.n92 gnd 0.264816f
C1891 CSoutput.n93 gnd 0.333931f
C1892 CSoutput.t43 gnd 0.045941f
C1893 CSoutput.t71 gnd 0.045941f
C1894 CSoutput.n94 gnd 0.355688f
C1895 CSoutput.t57 gnd 0.045941f
C1896 CSoutput.t58 gnd 0.045941f
C1897 CSoutput.n95 gnd 0.355054f
C1898 CSoutput.n96 gnd 0.360379f
C1899 CSoutput.t52 gnd 0.045941f
C1900 CSoutput.t42 gnd 0.045941f
C1901 CSoutput.n97 gnd 0.355054f
C1902 CSoutput.n98 gnd 0.17758f
C1903 CSoutput.t32 gnd 0.045941f
C1904 CSoutput.t53 gnd 0.045941f
C1905 CSoutput.n99 gnd 0.355054f
C1906 CSoutput.n100 gnd 0.264816f
C1907 CSoutput.n101 gnd 0.37325f
C1908 CSoutput.n102 gnd 7.31535f
C1909 CSoutput.n104 gnd 0.651523f
C1910 CSoutput.n105 gnd 0.488642f
C1911 CSoutput.n106 gnd 0.651523f
C1912 CSoutput.n107 gnd 0.651523f
C1913 CSoutput.n108 gnd 1.7541f
C1914 CSoutput.n109 gnd 0.651523f
C1915 CSoutput.n110 gnd 0.651523f
C1916 CSoutput.t139 gnd 0.814404f
C1917 CSoutput.n111 gnd 0.651523f
C1918 CSoutput.n112 gnd 0.651523f
C1919 CSoutput.n116 gnd 0.651523f
C1920 CSoutput.n120 gnd 0.651523f
C1921 CSoutput.n121 gnd 0.651523f
C1922 CSoutput.n123 gnd 0.651523f
C1923 CSoutput.n128 gnd 0.651523f
C1924 CSoutput.n130 gnd 0.651523f
C1925 CSoutput.n131 gnd 0.651523f
C1926 CSoutput.n133 gnd 0.651523f
C1927 CSoutput.n134 gnd 0.651523f
C1928 CSoutput.n136 gnd 0.651523f
C1929 CSoutput.t132 gnd 10.8869f
C1930 CSoutput.n138 gnd 0.651523f
C1931 CSoutput.n139 gnd 0.488642f
C1932 CSoutput.n140 gnd 0.651523f
C1933 CSoutput.n141 gnd 0.651523f
C1934 CSoutput.n142 gnd 1.7541f
C1935 CSoutput.n143 gnd 0.651523f
C1936 CSoutput.n144 gnd 0.651523f
C1937 CSoutput.t148 gnd 0.814404f
C1938 CSoutput.n145 gnd 0.651523f
C1939 CSoutput.n146 gnd 0.651523f
C1940 CSoutput.n150 gnd 0.651523f
C1941 CSoutput.n154 gnd 0.651523f
C1942 CSoutput.n155 gnd 0.651523f
C1943 CSoutput.n157 gnd 0.651523f
C1944 CSoutput.n162 gnd 0.651523f
C1945 CSoutput.n164 gnd 0.651523f
C1946 CSoutput.n165 gnd 0.651523f
C1947 CSoutput.n167 gnd 0.651523f
C1948 CSoutput.n168 gnd 0.651523f
C1949 CSoutput.n170 gnd 0.651523f
C1950 CSoutput.n171 gnd 0.488642f
C1951 CSoutput.n173 gnd 0.651523f
C1952 CSoutput.n174 gnd 0.488642f
C1953 CSoutput.n175 gnd 0.651523f
C1954 CSoutput.n176 gnd 0.651523f
C1955 CSoutput.n177 gnd 1.7541f
C1956 CSoutput.n178 gnd 0.651523f
C1957 CSoutput.n179 gnd 0.651523f
C1958 CSoutput.t142 gnd 0.814404f
C1959 CSoutput.n180 gnd 0.651523f
C1960 CSoutput.n181 gnd 1.7541f
C1961 CSoutput.n183 gnd 0.651523f
C1962 CSoutput.n184 gnd 0.651523f
C1963 CSoutput.n186 gnd 0.651523f
C1964 CSoutput.n187 gnd 0.651523f
C1965 CSoutput.t128 gnd 10.7095f
C1966 CSoutput.t135 gnd 10.8869f
C1967 CSoutput.n193 gnd 2.04392f
C1968 CSoutput.n194 gnd 8.3262f
C1969 CSoutput.n195 gnd 8.6746f
C1970 CSoutput.n200 gnd 2.21412f
C1971 CSoutput.n206 gnd 0.651523f
C1972 CSoutput.n208 gnd 0.651523f
C1973 CSoutput.n210 gnd 0.651523f
C1974 CSoutput.n212 gnd 0.651523f
C1975 CSoutput.n214 gnd 0.651523f
C1976 CSoutput.n220 gnd 0.651523f
C1977 CSoutput.n227 gnd 1.19529f
C1978 CSoutput.n228 gnd 1.19529f
C1979 CSoutput.n229 gnd 0.651523f
C1980 CSoutput.n230 gnd 0.651523f
C1981 CSoutput.n232 gnd 0.488642f
C1982 CSoutput.n233 gnd 0.418478f
C1983 CSoutput.n235 gnd 0.488642f
C1984 CSoutput.n236 gnd 0.418478f
C1985 CSoutput.n237 gnd 0.488642f
C1986 CSoutput.n239 gnd 0.651523f
C1987 CSoutput.n241 gnd 1.7541f
C1988 CSoutput.n242 gnd 2.04392f
C1989 CSoutput.n243 gnd 7.657959f
C1990 CSoutput.n245 gnd 0.488642f
C1991 CSoutput.n246 gnd 1.25731f
C1992 CSoutput.n247 gnd 0.488642f
C1993 CSoutput.n249 gnd 0.651523f
C1994 CSoutput.n251 gnd 1.7541f
C1995 CSoutput.n252 gnd 3.82071f
C1996 CSoutput.t59 gnd 0.045941f
C1997 CSoutput.t24 gnd 0.045941f
C1998 CSoutput.n253 gnd 0.355688f
C1999 CSoutput.t40 gnd 0.045941f
C2000 CSoutput.t29 gnd 0.045941f
C2001 CSoutput.n254 gnd 0.355054f
C2002 CSoutput.n255 gnd 0.360379f
C2003 CSoutput.t48 gnd 0.045941f
C2004 CSoutput.t37 gnd 0.045941f
C2005 CSoutput.n256 gnd 0.355054f
C2006 CSoutput.n257 gnd 0.17758f
C2007 CSoutput.t62 gnd 0.045941f
C2008 CSoutput.t31 gnd 0.045941f
C2009 CSoutput.n258 gnd 0.355054f
C2010 CSoutput.n259 gnd 0.32564f
C2011 CSoutput.t39 gnd 0.045941f
C2012 CSoutput.t65 gnd 0.045941f
C2013 CSoutput.n260 gnd 0.355688f
C2014 CSoutput.t36 gnd 0.045941f
C2015 CSoutput.t38 gnd 0.045941f
C2016 CSoutput.n261 gnd 0.355054f
C2017 CSoutput.n262 gnd 0.360379f
C2018 CSoutput.t63 gnd 0.045941f
C2019 CSoutput.t64 gnd 0.045941f
C2020 CSoutput.n263 gnd 0.355054f
C2021 CSoutput.n264 gnd 0.17758f
C2022 CSoutput.t27 gnd 0.045941f
C2023 CSoutput.t56 gnd 0.045941f
C2024 CSoutput.n265 gnd 0.355054f
C2025 CSoutput.n266 gnd 0.264816f
C2026 CSoutput.n267 gnd 0.333931f
C2027 CSoutput.t46 gnd 0.045941f
C2028 CSoutput.t69 gnd 0.045941f
C2029 CSoutput.n268 gnd 0.355688f
C2030 CSoutput.t44 gnd 0.045941f
C2031 CSoutput.t45 gnd 0.045941f
C2032 CSoutput.n269 gnd 0.355054f
C2033 CSoutput.n270 gnd 0.360379f
C2034 CSoutput.t67 gnd 0.045941f
C2035 CSoutput.t68 gnd 0.045941f
C2036 CSoutput.n271 gnd 0.355054f
C2037 CSoutput.n272 gnd 0.17758f
C2038 CSoutput.t34 gnd 0.045941f
C2039 CSoutput.t60 gnd 0.045941f
C2040 CSoutput.n273 gnd 0.355053f
C2041 CSoutput.n274 gnd 0.264817f
C2042 CSoutput.n275 gnd 0.37325f
C2043 CSoutput.n276 gnd 10.2443f
C2044 CSoutput.t99 gnd 0.040198f
C2045 CSoutput.t117 gnd 0.040198f
C2046 CSoutput.n277 gnd 0.356393f
C2047 CSoutput.t16 gnd 0.040198f
C2048 CSoutput.t84 gnd 0.040198f
C2049 CSoutput.n278 gnd 0.355205f
C2050 CSoutput.n279 gnd 0.330984f
C2051 CSoutput.t75 gnd 0.040198f
C2052 CSoutput.t9 gnd 0.040198f
C2053 CSoutput.n280 gnd 0.355205f
C2054 CSoutput.n281 gnd 0.16316f
C2055 CSoutput.t72 gnd 0.040198f
C2056 CSoutput.t98 gnd 0.040198f
C2057 CSoutput.n282 gnd 0.355205f
C2058 CSoutput.n283 gnd 0.16316f
C2059 CSoutput.t97 gnd 0.040198f
C2060 CSoutput.t18 gnd 0.040198f
C2061 CSoutput.n284 gnd 0.355205f
C2062 CSoutput.n285 gnd 0.16316f
C2063 CSoutput.t120 gnd 0.040198f
C2064 CSoutput.t85 gnd 0.040198f
C2065 CSoutput.n286 gnd 0.355205f
C2066 CSoutput.n287 gnd 0.16316f
C2067 CSoutput.t93 gnd 0.040198f
C2068 CSoutput.t103 gnd 0.040198f
C2069 CSoutput.n288 gnd 0.355205f
C2070 CSoutput.n289 gnd 0.16316f
C2071 CSoutput.t110 gnd 0.040198f
C2072 CSoutput.t114 gnd 0.040198f
C2073 CSoutput.n290 gnd 0.355205f
C2074 CSoutput.n291 gnd 0.16316f
C2075 CSoutput.t82 gnd 0.040198f
C2076 CSoutput.t4 gnd 0.040198f
C2077 CSoutput.n292 gnd 0.355205f
C2078 CSoutput.n293 gnd 0.16316f
C2079 CSoutput.t109 gnd 0.040198f
C2080 CSoutput.t7 gnd 0.040198f
C2081 CSoutput.n294 gnd 0.355205f
C2082 CSoutput.n295 gnd 0.3009f
C2083 CSoutput.t96 gnd 0.040198f
C2084 CSoutput.t88 gnd 0.040198f
C2085 CSoutput.n296 gnd 0.356393f
C2086 CSoutput.t15 gnd 0.040198f
C2087 CSoutput.t13 gnd 0.040198f
C2088 CSoutput.n297 gnd 0.355205f
C2089 CSoutput.n298 gnd 0.330984f
C2090 CSoutput.t124 gnd 0.040198f
C2091 CSoutput.t116 gnd 0.040198f
C2092 CSoutput.n299 gnd 0.355205f
C2093 CSoutput.n300 gnd 0.16316f
C2094 CSoutput.t10 gnd 0.040198f
C2095 CSoutput.t81 gnd 0.040198f
C2096 CSoutput.n301 gnd 0.355205f
C2097 CSoutput.n302 gnd 0.16316f
C2098 CSoutput.t77 gnd 0.040198f
C2099 CSoutput.t125 gnd 0.040198f
C2100 CSoutput.n303 gnd 0.355205f
C2101 CSoutput.n304 gnd 0.16316f
C2102 CSoutput.t108 gnd 0.040198f
C2103 CSoutput.t92 gnd 0.040198f
C2104 CSoutput.n305 gnd 0.355205f
C2105 CSoutput.n306 gnd 0.16316f
C2106 CSoutput.t78 gnd 0.040198f
C2107 CSoutput.t17 gnd 0.040198f
C2108 CSoutput.n307 gnd 0.355205f
C2109 CSoutput.n308 gnd 0.16316f
C2110 CSoutput.t94 gnd 0.040198f
C2111 CSoutput.t73 gnd 0.040198f
C2112 CSoutput.n309 gnd 0.355205f
C2113 CSoutput.n310 gnd 0.16316f
C2114 CSoutput.t87 gnd 0.040198f
C2115 CSoutput.t22 gnd 0.040198f
C2116 CSoutput.n311 gnd 0.355205f
C2117 CSoutput.n312 gnd 0.16316f
C2118 CSoutput.t2 gnd 0.040198f
C2119 CSoutput.t6 gnd 0.040198f
C2120 CSoutput.n313 gnd 0.355205f
C2121 CSoutput.n314 gnd 0.247711f
C2122 CSoutput.n315 gnd 0.460267f
C2123 CSoutput.n316 gnd 10.924f
C2124 CSoutput.t20 gnd 0.040198f
C2125 CSoutput.t102 gnd 0.040198f
C2126 CSoutput.n317 gnd 0.356393f
C2127 CSoutput.t74 gnd 0.040198f
C2128 CSoutput.t0 gnd 0.040198f
C2129 CSoutput.n318 gnd 0.355205f
C2130 CSoutput.n319 gnd 0.330984f
C2131 CSoutput.t91 gnd 0.040198f
C2132 CSoutput.t118 gnd 0.040198f
C2133 CSoutput.n320 gnd 0.355205f
C2134 CSoutput.n321 gnd 0.16316f
C2135 CSoutput.t104 gnd 0.040198f
C2136 CSoutput.t3 gnd 0.040198f
C2137 CSoutput.n322 gnd 0.355205f
C2138 CSoutput.n323 gnd 0.16316f
C2139 CSoutput.t19 gnd 0.040198f
C2140 CSoutput.t89 gnd 0.040198f
C2141 CSoutput.n324 gnd 0.355205f
C2142 CSoutput.n325 gnd 0.16316f
C2143 CSoutput.t76 gnd 0.040198f
C2144 CSoutput.t119 gnd 0.040198f
C2145 CSoutput.n326 gnd 0.355205f
C2146 CSoutput.n327 gnd 0.16316f
C2147 CSoutput.t123 gnd 0.040198f
C2148 CSoutput.t14 gnd 0.040198f
C2149 CSoutput.n328 gnd 0.355205f
C2150 CSoutput.n329 gnd 0.16316f
C2151 CSoutput.t126 gnd 0.040198f
C2152 CSoutput.t115 gnd 0.040198f
C2153 CSoutput.n330 gnd 0.355205f
C2154 CSoutput.n331 gnd 0.16316f
C2155 CSoutput.t107 gnd 0.040198f
C2156 CSoutput.t83 gnd 0.040198f
C2157 CSoutput.n332 gnd 0.355205f
C2158 CSoutput.n333 gnd 0.16316f
C2159 CSoutput.t79 gnd 0.040198f
C2160 CSoutput.t105 gnd 0.040198f
C2161 CSoutput.n334 gnd 0.355205f
C2162 CSoutput.n335 gnd 0.3009f
C2163 CSoutput.t90 gnd 0.040198f
C2164 CSoutput.t8 gnd 0.040198f
C2165 CSoutput.n336 gnd 0.356393f
C2166 CSoutput.t5 gnd 0.040198f
C2167 CSoutput.t21 gnd 0.040198f
C2168 CSoutput.n337 gnd 0.355205f
C2169 CSoutput.n338 gnd 0.330984f
C2170 CSoutput.t23 gnd 0.040198f
C2171 CSoutput.t100 gnd 0.040198f
C2172 CSoutput.n339 gnd 0.355205f
C2173 CSoutput.n340 gnd 0.16316f
C2174 CSoutput.t111 gnd 0.040198f
C2175 CSoutput.t80 gnd 0.040198f
C2176 CSoutput.n341 gnd 0.355205f
C2177 CSoutput.n342 gnd 0.16316f
C2178 CSoutput.t127 gnd 0.040198f
C2179 CSoutput.t1 gnd 0.040198f
C2180 CSoutput.n343 gnd 0.355205f
C2181 CSoutput.n344 gnd 0.16316f
C2182 CSoutput.t113 gnd 0.040198f
C2183 CSoutput.t95 gnd 0.040198f
C2184 CSoutput.n345 gnd 0.355205f
C2185 CSoutput.n346 gnd 0.16316f
C2186 CSoutput.t122 gnd 0.040198f
C2187 CSoutput.t121 gnd 0.040198f
C2188 CSoutput.n347 gnd 0.355205f
C2189 CSoutput.n348 gnd 0.16316f
C2190 CSoutput.t106 gnd 0.040198f
C2191 CSoutput.t112 gnd 0.040198f
C2192 CSoutput.n349 gnd 0.355205f
C2193 CSoutput.n350 gnd 0.16316f
C2194 CSoutput.t11 gnd 0.040198f
C2195 CSoutput.t101 gnd 0.040198f
C2196 CSoutput.n351 gnd 0.355205f
C2197 CSoutput.n352 gnd 0.16316f
C2198 CSoutput.t86 gnd 0.040198f
C2199 CSoutput.t12 gnd 0.040198f
C2200 CSoutput.n353 gnd 0.355205f
C2201 CSoutput.n354 gnd 0.247711f
C2202 CSoutput.n355 gnd 0.460267f
C2203 CSoutput.n356 gnd 6.47139f
C2204 CSoutput.n357 gnd 11.981299f
C2205 a_n6972_8799.n0 gnd 4.28018f
C2206 a_n6972_8799.n1 gnd 2.09493f
C2207 a_n6972_8799.n2 gnd 3.51776f
C2208 a_n6972_8799.n3 gnd 0.877192f
C2209 a_n6972_8799.n4 gnd 0.207515f
C2210 a_n6972_8799.n5 gnd 0.28608f
C2211 a_n6972_8799.n6 gnd 0.217052f
C2212 a_n6972_8799.n7 gnd 0.207515f
C2213 a_n6972_8799.n8 gnd 0.28608f
C2214 a_n6972_8799.n9 gnd 0.217052f
C2215 a_n6972_8799.n10 gnd 0.207515f
C2216 a_n6972_8799.n11 gnd 0.450837f
C2217 a_n6972_8799.n12 gnd 0.217052f
C2218 a_n6972_8799.n13 gnd 0.207515f
C2219 a_n6972_8799.n14 gnd 0.32081f
C2220 a_n6972_8799.n15 gnd 0.182323f
C2221 a_n6972_8799.n16 gnd 0.207515f
C2222 a_n6972_8799.n17 gnd 0.32081f
C2223 a_n6972_8799.n18 gnd 0.182323f
C2224 a_n6972_8799.n19 gnd 0.207515f
C2225 a_n6972_8799.n20 gnd 0.32081f
C2226 a_n6972_8799.n21 gnd 0.34708f
C2227 a_n6972_8799.n22 gnd 1.52091f
C2228 a_n6972_8799.n23 gnd 2.71756f
C2229 a_n6972_8799.n24 gnd 3.99645f
C2230 a_n6972_8799.n25 gnd 1.52091f
C2231 a_n6972_8799.n26 gnd 0.249828f
C2232 a_n6972_8799.n27 gnd 0.004664f
C2233 a_n6972_8799.n28 gnd 0.010087f
C2234 a_n6972_8799.n29 gnd 0.010087f
C2235 a_n6972_8799.n30 gnd 0.004664f
C2236 a_n6972_8799.n31 gnd 0.249828f
C2237 a_n6972_8799.n32 gnd 0.004664f
C2238 a_n6972_8799.n33 gnd 0.010087f
C2239 a_n6972_8799.n34 gnd 0.010087f
C2240 a_n6972_8799.n35 gnd 0.004664f
C2241 a_n6972_8799.n36 gnd 0.249828f
C2242 a_n6972_8799.n37 gnd 0.004664f
C2243 a_n6972_8799.n38 gnd 0.010087f
C2244 a_n6972_8799.n39 gnd 0.010087f
C2245 a_n6972_8799.n40 gnd 0.004664f
C2246 a_n6972_8799.n41 gnd 0.004664f
C2247 a_n6972_8799.n42 gnd 0.010087f
C2248 a_n6972_8799.n43 gnd 0.010087f
C2249 a_n6972_8799.n44 gnd 0.004664f
C2250 a_n6972_8799.n45 gnd 0.249828f
C2251 a_n6972_8799.n46 gnd 0.004664f
C2252 a_n6972_8799.n47 gnd 0.010087f
C2253 a_n6972_8799.n48 gnd 0.010087f
C2254 a_n6972_8799.n49 gnd 0.004664f
C2255 a_n6972_8799.n50 gnd 0.249828f
C2256 a_n6972_8799.n51 gnd 0.004664f
C2257 a_n6972_8799.n52 gnd 0.010087f
C2258 a_n6972_8799.n53 gnd 0.010087f
C2259 a_n6972_8799.n54 gnd 0.004664f
C2260 a_n6972_8799.n55 gnd 0.249828f
C2261 a_n6972_8799.t36 gnd 0.143935f
C2262 a_n6972_8799.t33 gnd 0.143935f
C2263 a_n6972_8799.t30 gnd 0.143935f
C2264 a_n6972_8799.n56 gnd 1.13523f
C2265 a_n6972_8799.t18 gnd 0.143935f
C2266 a_n6972_8799.t20 gnd 0.143935f
C2267 a_n6972_8799.n57 gnd 1.13336f
C2268 a_n6972_8799.t32 gnd 0.143935f
C2269 a_n6972_8799.t24 gnd 0.143935f
C2270 a_n6972_8799.n58 gnd 1.13336f
C2271 a_n6972_8799.t19 gnd 0.143935f
C2272 a_n6972_8799.t27 gnd 0.143935f
C2273 a_n6972_8799.n59 gnd 1.13336f
C2274 a_n6972_8799.t31 gnd 0.143935f
C2275 a_n6972_8799.t21 gnd 0.143935f
C2276 a_n6972_8799.n60 gnd 1.13336f
C2277 a_n6972_8799.t11 gnd 0.111949f
C2278 a_n6972_8799.t43 gnd 0.111949f
C2279 a_n6972_8799.n61 gnd 0.992138f
C2280 a_n6972_8799.t8 gnd 0.111949f
C2281 a_n6972_8799.t37 gnd 0.111949f
C2282 a_n6972_8799.n62 gnd 0.989221f
C2283 a_n6972_8799.t12 gnd 0.111949f
C2284 a_n6972_8799.t1 gnd 0.111949f
C2285 a_n6972_8799.n63 gnd 0.989221f
C2286 a_n6972_8799.t3 gnd 0.111949f
C2287 a_n6972_8799.t40 gnd 0.111949f
C2288 a_n6972_8799.n64 gnd 0.992137f
C2289 a_n6972_8799.t41 gnd 0.111949f
C2290 a_n6972_8799.t42 gnd 0.111949f
C2291 a_n6972_8799.n65 gnd 0.98922f
C2292 a_n6972_8799.t7 gnd 0.111949f
C2293 a_n6972_8799.t39 gnd 0.111949f
C2294 a_n6972_8799.n66 gnd 0.98922f
C2295 a_n6972_8799.t4 gnd 0.111949f
C2296 a_n6972_8799.t14 gnd 0.111949f
C2297 a_n6972_8799.n67 gnd 0.992137f
C2298 a_n6972_8799.t15 gnd 0.111949f
C2299 a_n6972_8799.t6 gnd 0.111949f
C2300 a_n6972_8799.n68 gnd 0.98922f
C2301 a_n6972_8799.t16 gnd 0.111949f
C2302 a_n6972_8799.t2 gnd 0.111949f
C2303 a_n6972_8799.n69 gnd 0.98922f
C2304 a_n6972_8799.t10 gnd 0.111949f
C2305 a_n6972_8799.t9 gnd 0.111949f
C2306 a_n6972_8799.n70 gnd 0.989221f
C2307 a_n6972_8799.t0 gnd 0.111949f
C2308 a_n6972_8799.t13 gnd 0.111949f
C2309 a_n6972_8799.n71 gnd 0.989221f
C2310 a_n6972_8799.t38 gnd 0.111949f
C2311 a_n6972_8799.t5 gnd 0.111949f
C2312 a_n6972_8799.n72 gnd 0.989221f
C2313 a_n6972_8799.t57 gnd 0.596819f
C2314 a_n6972_8799.n73 gnd 0.268236f
C2315 a_n6972_8799.t73 gnd 0.596819f
C2316 a_n6972_8799.t62 gnd 0.596819f
C2317 a_n6972_8799.t83 gnd 0.608115f
C2318 a_n6972_8799.n74 gnd 0.250196f
C2319 a_n6972_8799.n75 gnd 0.270621f
C2320 a_n6972_8799.t63 gnd 0.596819f
C2321 a_n6972_8799.n76 gnd 0.268236f
C2322 a_n6972_8799.n77 gnd 0.263832f
C2323 a_n6972_8799.t58 gnd 0.596819f
C2324 a_n6972_8799.n78 gnd 0.263832f
C2325 a_n6972_8799.t72 gnd 0.596819f
C2326 a_n6972_8799.n79 gnd 0.270621f
C2327 a_n6972_8799.t44 gnd 0.608105f
C2328 a_n6972_8799.t61 gnd 0.596819f
C2329 a_n6972_8799.n80 gnd 0.268236f
C2330 a_n6972_8799.t82 gnd 0.596819f
C2331 a_n6972_8799.t66 gnd 0.596819f
C2332 a_n6972_8799.t90 gnd 0.608115f
C2333 a_n6972_8799.n81 gnd 0.250196f
C2334 a_n6972_8799.n82 gnd 0.270621f
C2335 a_n6972_8799.t65 gnd 0.596819f
C2336 a_n6972_8799.n83 gnd 0.268236f
C2337 a_n6972_8799.n84 gnd 0.263832f
C2338 a_n6972_8799.t60 gnd 0.596819f
C2339 a_n6972_8799.n85 gnd 0.263832f
C2340 a_n6972_8799.t80 gnd 0.596819f
C2341 a_n6972_8799.n86 gnd 0.270621f
C2342 a_n6972_8799.t49 gnd 0.608105f
C2343 a_n6972_8799.n87 gnd 0.897596f
C2344 a_n6972_8799.t74 gnd 0.596819f
C2345 a_n6972_8799.n88 gnd 0.268236f
C2346 a_n6972_8799.t68 gnd 0.596819f
C2347 a_n6972_8799.t54 gnd 0.596819f
C2348 a_n6972_8799.t85 gnd 0.608115f
C2349 a_n6972_8799.n89 gnd 0.250196f
C2350 a_n6972_8799.n90 gnd 0.270621f
C2351 a_n6972_8799.t45 gnd 0.596819f
C2352 a_n6972_8799.n91 gnd 0.268236f
C2353 a_n6972_8799.n92 gnd 0.263832f
C2354 a_n6972_8799.t87 gnd 0.596819f
C2355 a_n6972_8799.n93 gnd 0.263832f
C2356 a_n6972_8799.t89 gnd 0.596819f
C2357 a_n6972_8799.n94 gnd 0.270621f
C2358 a_n6972_8799.t64 gnd 0.608105f
C2359 a_n6972_8799.n95 gnd 1.80286f
C2360 a_n6972_8799.t69 gnd 0.608105f
C2361 a_n6972_8799.t46 gnd 0.596819f
C2362 a_n6972_8799.t71 gnd 0.596819f
C2363 a_n6972_8799.n96 gnd 0.268236f
C2364 a_n6972_8799.t70 gnd 0.596819f
C2365 a_n6972_8799.t48 gnd 0.596819f
C2366 a_n6972_8799.t47 gnd 0.596819f
C2367 a_n6972_8799.n97 gnd 0.268236f
C2368 a_n6972_8799.t55 gnd 0.608115f
C2369 a_n6972_8799.n98 gnd 0.250196f
C2370 a_n6972_8799.t81 gnd 0.596819f
C2371 a_n6972_8799.n99 gnd 0.270621f
C2372 a_n6972_8799.n100 gnd 0.263832f
C2373 a_n6972_8799.n101 gnd 0.263832f
C2374 a_n6972_8799.n102 gnd 0.270621f
C2375 a_n6972_8799.t76 gnd 0.608105f
C2376 a_n6972_8799.t50 gnd 0.596819f
C2377 a_n6972_8799.t79 gnd 0.596819f
C2378 a_n6972_8799.n103 gnd 0.268236f
C2379 a_n6972_8799.t77 gnd 0.596819f
C2380 a_n6972_8799.t52 gnd 0.596819f
C2381 a_n6972_8799.t51 gnd 0.596819f
C2382 a_n6972_8799.n104 gnd 0.268236f
C2383 a_n6972_8799.t59 gnd 0.608115f
C2384 a_n6972_8799.n105 gnd 0.250196f
C2385 a_n6972_8799.t88 gnd 0.596819f
C2386 a_n6972_8799.n106 gnd 0.270621f
C2387 a_n6972_8799.n107 gnd 0.263832f
C2388 a_n6972_8799.n108 gnd 0.263832f
C2389 a_n6972_8799.n109 gnd 0.270621f
C2390 a_n6972_8799.n110 gnd 0.897596f
C2391 a_n6972_8799.t56 gnd 0.608105f
C2392 a_n6972_8799.t91 gnd 0.596819f
C2393 a_n6972_8799.t75 gnd 0.596819f
C2394 a_n6972_8799.n111 gnd 0.268236f
C2395 a_n6972_8799.t86 gnd 0.596819f
C2396 a_n6972_8799.t67 gnd 0.596819f
C2397 a_n6972_8799.t78 gnd 0.596819f
C2398 a_n6972_8799.n112 gnd 0.268236f
C2399 a_n6972_8799.t84 gnd 0.608115f
C2400 a_n6972_8799.n113 gnd 0.250196f
C2401 a_n6972_8799.t53 gnd 0.596819f
C2402 a_n6972_8799.n114 gnd 0.270621f
C2403 a_n6972_8799.n115 gnd 0.263832f
C2404 a_n6972_8799.n116 gnd 0.263832f
C2405 a_n6972_8799.n117 gnd 0.270621f
C2406 a_n6972_8799.n118 gnd 1.24031f
C2407 a_n6972_8799.n119 gnd 15.629401f
C2408 a_n6972_8799.n120 gnd 4.36785f
C2409 a_n6972_8799.n121 gnd 6.97062f
C2410 a_n6972_8799.t25 gnd 0.143935f
C2411 a_n6972_8799.t35 gnd 0.143935f
C2412 a_n6972_8799.n122 gnd 1.13336f
C2413 a_n6972_8799.t28 gnd 0.143935f
C2414 a_n6972_8799.t22 gnd 0.143935f
C2415 a_n6972_8799.n123 gnd 1.13336f
C2416 a_n6972_8799.t23 gnd 0.143935f
C2417 a_n6972_8799.t26 gnd 0.143935f
C2418 a_n6972_8799.n124 gnd 1.13336f
C2419 a_n6972_8799.t29 gnd 0.143935f
C2420 a_n6972_8799.t34 gnd 0.143935f
C2421 a_n6972_8799.n125 gnd 1.13336f
C2422 a_n6972_8799.n126 gnd 1.13524f
C2423 a_n6972_8799.t17 gnd 0.143935f
C2424 vdd.t190 gnd 0.030489f
C2425 vdd.t171 gnd 0.030489f
C2426 vdd.n0 gnd 0.24047f
C2427 vdd.t152 gnd 0.030489f
C2428 vdd.t185 gnd 0.030489f
C2429 vdd.n1 gnd 0.240073f
C2430 vdd.n2 gnd 0.221393f
C2431 vdd.t168 gnd 0.030489f
C2432 vdd.t194 gnd 0.030489f
C2433 vdd.n3 gnd 0.240073f
C2434 vdd.n4 gnd 0.111967f
C2435 vdd.t192 gnd 0.030489f
C2436 vdd.t173 gnd 0.030489f
C2437 vdd.n5 gnd 0.240073f
C2438 vdd.n6 gnd 0.10506f
C2439 vdd.t200 gnd 0.030489f
C2440 vdd.t166 gnd 0.030489f
C2441 vdd.n7 gnd 0.24047f
C2442 vdd.t176 gnd 0.030489f
C2443 vdd.t196 gnd 0.030489f
C2444 vdd.n8 gnd 0.240073f
C2445 vdd.n9 gnd 0.221393f
C2446 vdd.t182 gnd 0.030489f
C2447 vdd.t155 gnd 0.030489f
C2448 vdd.n10 gnd 0.240073f
C2449 vdd.n11 gnd 0.111967f
C2450 vdd.t163 gnd 0.030489f
C2451 vdd.t180 gnd 0.030489f
C2452 vdd.n12 gnd 0.240073f
C2453 vdd.n13 gnd 0.10506f
C2454 vdd.n14 gnd 0.074276f
C2455 vdd.t111 gnd 0.016938f
C2456 vdd.t132 gnd 0.016938f
C2457 vdd.n15 gnd 0.155909f
C2458 vdd.t26 gnd 0.016938f
C2459 vdd.t109 gnd 0.016938f
C2460 vdd.n16 gnd 0.155453f
C2461 vdd.n17 gnd 0.270537f
C2462 vdd.t136 gnd 0.016938f
C2463 vdd.t133 gnd 0.016938f
C2464 vdd.n18 gnd 0.155453f
C2465 vdd.n19 gnd 0.111925f
C2466 vdd.t27 gnd 0.016938f
C2467 vdd.t110 gnd 0.016938f
C2468 vdd.n20 gnd 0.155909f
C2469 vdd.t4 gnd 0.016938f
C2470 vdd.t105 gnd 0.016938f
C2471 vdd.n21 gnd 0.155453f
C2472 vdd.n22 gnd 0.270537f
C2473 vdd.t115 gnd 0.016938f
C2474 vdd.t5 gnd 0.016938f
C2475 vdd.n23 gnd 0.155453f
C2476 vdd.n24 gnd 0.111925f
C2477 vdd.t137 gnd 0.016938f
C2478 vdd.t104 gnd 0.016938f
C2479 vdd.n25 gnd 0.155453f
C2480 vdd.t113 gnd 0.016938f
C2481 vdd.t114 gnd 0.016938f
C2482 vdd.n26 gnd 0.155453f
C2483 vdd.n27 gnd 18.0956f
C2484 vdd.n28 gnd 6.85786f
C2485 vdd.n29 gnd 0.00462f
C2486 vdd.n30 gnd 0.004287f
C2487 vdd.n31 gnd 0.002371f
C2488 vdd.n32 gnd 0.005445f
C2489 vdd.n33 gnd 0.002304f
C2490 vdd.n34 gnd 0.002439f
C2491 vdd.n35 gnd 0.004287f
C2492 vdd.n36 gnd 0.002304f
C2493 vdd.n37 gnd 0.005445f
C2494 vdd.n38 gnd 0.002439f
C2495 vdd.n39 gnd 0.004287f
C2496 vdd.n40 gnd 0.002304f
C2497 vdd.n41 gnd 0.004084f
C2498 vdd.n42 gnd 0.004096f
C2499 vdd.t108 gnd 0.011698f
C2500 vdd.n43 gnd 0.026027f
C2501 vdd.n44 gnd 0.135453f
C2502 vdd.n45 gnd 0.002304f
C2503 vdd.n46 gnd 0.002439f
C2504 vdd.n47 gnd 0.005445f
C2505 vdd.n48 gnd 0.005445f
C2506 vdd.n49 gnd 0.002439f
C2507 vdd.n50 gnd 0.002304f
C2508 vdd.n51 gnd 0.004287f
C2509 vdd.n52 gnd 0.004287f
C2510 vdd.n53 gnd 0.002304f
C2511 vdd.n54 gnd 0.002439f
C2512 vdd.n55 gnd 0.005445f
C2513 vdd.n56 gnd 0.005445f
C2514 vdd.n57 gnd 0.002439f
C2515 vdd.n58 gnd 0.002304f
C2516 vdd.n59 gnd 0.004287f
C2517 vdd.n60 gnd 0.004287f
C2518 vdd.n61 gnd 0.002304f
C2519 vdd.n62 gnd 0.002439f
C2520 vdd.n63 gnd 0.005445f
C2521 vdd.n64 gnd 0.005445f
C2522 vdd.n65 gnd 0.012873f
C2523 vdd.n66 gnd 0.002371f
C2524 vdd.n67 gnd 0.002304f
C2525 vdd.n68 gnd 0.01108f
C2526 vdd.n69 gnd 0.007736f
C2527 vdd.t142 gnd 0.027101f
C2528 vdd.t25 gnd 0.027101f
C2529 vdd.n70 gnd 0.186258f
C2530 vdd.n71 gnd 0.146463f
C2531 vdd.t145 gnd 0.027101f
C2532 vdd.t135 gnd 0.027101f
C2533 vdd.n72 gnd 0.186258f
C2534 vdd.n73 gnd 0.118195f
C2535 vdd.t20 gnd 0.027101f
C2536 vdd.t125 gnd 0.027101f
C2537 vdd.n74 gnd 0.186258f
C2538 vdd.n75 gnd 0.118195f
C2539 vdd.n76 gnd 0.00462f
C2540 vdd.n77 gnd 0.004287f
C2541 vdd.n78 gnd 0.002371f
C2542 vdd.n79 gnd 0.005445f
C2543 vdd.n80 gnd 0.002304f
C2544 vdd.n81 gnd 0.002439f
C2545 vdd.n82 gnd 0.004287f
C2546 vdd.n83 gnd 0.002304f
C2547 vdd.n84 gnd 0.005445f
C2548 vdd.n85 gnd 0.002439f
C2549 vdd.n86 gnd 0.004287f
C2550 vdd.n87 gnd 0.002304f
C2551 vdd.n88 gnd 0.004084f
C2552 vdd.n89 gnd 0.004096f
C2553 vdd.t23 gnd 0.011698f
C2554 vdd.n90 gnd 0.026027f
C2555 vdd.n91 gnd 0.135453f
C2556 vdd.n92 gnd 0.002304f
C2557 vdd.n93 gnd 0.002439f
C2558 vdd.n94 gnd 0.005445f
C2559 vdd.n95 gnd 0.005445f
C2560 vdd.n96 gnd 0.002439f
C2561 vdd.n97 gnd 0.002304f
C2562 vdd.n98 gnd 0.004287f
C2563 vdd.n99 gnd 0.004287f
C2564 vdd.n100 gnd 0.002304f
C2565 vdd.n101 gnd 0.002439f
C2566 vdd.n102 gnd 0.005445f
C2567 vdd.n103 gnd 0.005445f
C2568 vdd.n104 gnd 0.002439f
C2569 vdd.n105 gnd 0.002304f
C2570 vdd.n106 gnd 0.004287f
C2571 vdd.n107 gnd 0.004287f
C2572 vdd.n108 gnd 0.002304f
C2573 vdd.n109 gnd 0.002439f
C2574 vdd.n110 gnd 0.005445f
C2575 vdd.n111 gnd 0.005445f
C2576 vdd.n112 gnd 0.012873f
C2577 vdd.n113 gnd 0.002371f
C2578 vdd.n114 gnd 0.002304f
C2579 vdd.n115 gnd 0.01108f
C2580 vdd.n116 gnd 0.007493f
C2581 vdd.n117 gnd 0.087938f
C2582 vdd.n118 gnd 0.00462f
C2583 vdd.n119 gnd 0.004287f
C2584 vdd.n120 gnd 0.002371f
C2585 vdd.n121 gnd 0.005445f
C2586 vdd.n122 gnd 0.002304f
C2587 vdd.n123 gnd 0.002439f
C2588 vdd.n124 gnd 0.004287f
C2589 vdd.n125 gnd 0.002304f
C2590 vdd.n126 gnd 0.005445f
C2591 vdd.n127 gnd 0.002439f
C2592 vdd.n128 gnd 0.004287f
C2593 vdd.n129 gnd 0.002304f
C2594 vdd.n130 gnd 0.004084f
C2595 vdd.n131 gnd 0.004096f
C2596 vdd.t14 gnd 0.011698f
C2597 vdd.n132 gnd 0.026027f
C2598 vdd.n133 gnd 0.135453f
C2599 vdd.n134 gnd 0.002304f
C2600 vdd.n135 gnd 0.002439f
C2601 vdd.n136 gnd 0.005445f
C2602 vdd.n137 gnd 0.005445f
C2603 vdd.n138 gnd 0.002439f
C2604 vdd.n139 gnd 0.002304f
C2605 vdd.n140 gnd 0.004287f
C2606 vdd.n141 gnd 0.004287f
C2607 vdd.n142 gnd 0.002304f
C2608 vdd.n143 gnd 0.002439f
C2609 vdd.n144 gnd 0.005445f
C2610 vdd.n145 gnd 0.005445f
C2611 vdd.n146 gnd 0.002439f
C2612 vdd.n147 gnd 0.002304f
C2613 vdd.n148 gnd 0.004287f
C2614 vdd.n149 gnd 0.004287f
C2615 vdd.n150 gnd 0.002304f
C2616 vdd.n151 gnd 0.002439f
C2617 vdd.n152 gnd 0.005445f
C2618 vdd.n153 gnd 0.005445f
C2619 vdd.n154 gnd 0.012873f
C2620 vdd.n155 gnd 0.002371f
C2621 vdd.n156 gnd 0.002304f
C2622 vdd.n157 gnd 0.01108f
C2623 vdd.n158 gnd 0.007736f
C2624 vdd.t141 gnd 0.027101f
C2625 vdd.t129 gnd 0.027101f
C2626 vdd.n159 gnd 0.186258f
C2627 vdd.n160 gnd 0.146463f
C2628 vdd.t19 gnd 0.027101f
C2629 vdd.t206 gnd 0.027101f
C2630 vdd.n161 gnd 0.186258f
C2631 vdd.n162 gnd 0.118195f
C2632 vdd.t11 gnd 0.027101f
C2633 vdd.t143 gnd 0.027101f
C2634 vdd.n163 gnd 0.186258f
C2635 vdd.n164 gnd 0.118195f
C2636 vdd.n165 gnd 0.00462f
C2637 vdd.n166 gnd 0.004287f
C2638 vdd.n167 gnd 0.002371f
C2639 vdd.n168 gnd 0.005445f
C2640 vdd.n169 gnd 0.002304f
C2641 vdd.n170 gnd 0.002439f
C2642 vdd.n171 gnd 0.004287f
C2643 vdd.n172 gnd 0.002304f
C2644 vdd.n173 gnd 0.005445f
C2645 vdd.n174 gnd 0.002439f
C2646 vdd.n175 gnd 0.004287f
C2647 vdd.n176 gnd 0.002304f
C2648 vdd.n177 gnd 0.004084f
C2649 vdd.n178 gnd 0.004096f
C2650 vdd.t146 gnd 0.011698f
C2651 vdd.n179 gnd 0.026027f
C2652 vdd.n180 gnd 0.135453f
C2653 vdd.n181 gnd 0.002304f
C2654 vdd.n182 gnd 0.002439f
C2655 vdd.n183 gnd 0.005445f
C2656 vdd.n184 gnd 0.005445f
C2657 vdd.n185 gnd 0.002439f
C2658 vdd.n186 gnd 0.002304f
C2659 vdd.n187 gnd 0.004287f
C2660 vdd.n188 gnd 0.004287f
C2661 vdd.n189 gnd 0.002304f
C2662 vdd.n190 gnd 0.002439f
C2663 vdd.n191 gnd 0.005445f
C2664 vdd.n192 gnd 0.005445f
C2665 vdd.n193 gnd 0.002439f
C2666 vdd.n194 gnd 0.002304f
C2667 vdd.n195 gnd 0.004287f
C2668 vdd.n196 gnd 0.004287f
C2669 vdd.n197 gnd 0.002304f
C2670 vdd.n198 gnd 0.002439f
C2671 vdd.n199 gnd 0.005445f
C2672 vdd.n200 gnd 0.005445f
C2673 vdd.n201 gnd 0.012873f
C2674 vdd.n202 gnd 0.002371f
C2675 vdd.n203 gnd 0.002304f
C2676 vdd.n204 gnd 0.01108f
C2677 vdd.n205 gnd 0.007493f
C2678 vdd.n206 gnd 0.052314f
C2679 vdd.n207 gnd 0.188501f
C2680 vdd.n208 gnd 0.00462f
C2681 vdd.n209 gnd 0.004287f
C2682 vdd.n210 gnd 0.002371f
C2683 vdd.n211 gnd 0.005445f
C2684 vdd.n212 gnd 0.002304f
C2685 vdd.n213 gnd 0.002439f
C2686 vdd.n214 gnd 0.004287f
C2687 vdd.n215 gnd 0.002304f
C2688 vdd.n216 gnd 0.005445f
C2689 vdd.n217 gnd 0.002439f
C2690 vdd.n218 gnd 0.004287f
C2691 vdd.n219 gnd 0.002304f
C2692 vdd.n220 gnd 0.004084f
C2693 vdd.n221 gnd 0.004096f
C2694 vdd.t3 gnd 0.011698f
C2695 vdd.n222 gnd 0.026027f
C2696 vdd.n223 gnd 0.135453f
C2697 vdd.n224 gnd 0.002304f
C2698 vdd.n225 gnd 0.002439f
C2699 vdd.n226 gnd 0.005445f
C2700 vdd.n227 gnd 0.005445f
C2701 vdd.n228 gnd 0.002439f
C2702 vdd.n229 gnd 0.002304f
C2703 vdd.n230 gnd 0.004287f
C2704 vdd.n231 gnd 0.004287f
C2705 vdd.n232 gnd 0.002304f
C2706 vdd.n233 gnd 0.002439f
C2707 vdd.n234 gnd 0.005445f
C2708 vdd.n235 gnd 0.005445f
C2709 vdd.n236 gnd 0.002439f
C2710 vdd.n237 gnd 0.002304f
C2711 vdd.n238 gnd 0.004287f
C2712 vdd.n239 gnd 0.004287f
C2713 vdd.n240 gnd 0.002304f
C2714 vdd.n241 gnd 0.002439f
C2715 vdd.n242 gnd 0.005445f
C2716 vdd.n243 gnd 0.005445f
C2717 vdd.n244 gnd 0.012873f
C2718 vdd.n245 gnd 0.002371f
C2719 vdd.n246 gnd 0.002304f
C2720 vdd.n247 gnd 0.01108f
C2721 vdd.n248 gnd 0.007736f
C2722 vdd.t140 gnd 0.027101f
C2723 vdd.t116 gnd 0.027101f
C2724 vdd.n249 gnd 0.186258f
C2725 vdd.n250 gnd 0.146463f
C2726 vdd.t128 gnd 0.027101f
C2727 vdd.t118 gnd 0.027101f
C2728 vdd.n251 gnd 0.186258f
C2729 vdd.n252 gnd 0.118195f
C2730 vdd.t148 gnd 0.027101f
C2731 vdd.t207 gnd 0.027101f
C2732 vdd.n253 gnd 0.186258f
C2733 vdd.n254 gnd 0.118195f
C2734 vdd.n255 gnd 0.00462f
C2735 vdd.n256 gnd 0.004287f
C2736 vdd.n257 gnd 0.002371f
C2737 vdd.n258 gnd 0.005445f
C2738 vdd.n259 gnd 0.002304f
C2739 vdd.n260 gnd 0.002439f
C2740 vdd.n261 gnd 0.004287f
C2741 vdd.n262 gnd 0.002304f
C2742 vdd.n263 gnd 0.005445f
C2743 vdd.n264 gnd 0.002439f
C2744 vdd.n265 gnd 0.004287f
C2745 vdd.n266 gnd 0.002304f
C2746 vdd.n267 gnd 0.004084f
C2747 vdd.n268 gnd 0.004096f
C2748 vdd.t9 gnd 0.011698f
C2749 vdd.n269 gnd 0.026027f
C2750 vdd.n270 gnd 0.135453f
C2751 vdd.n271 gnd 0.002304f
C2752 vdd.n272 gnd 0.002439f
C2753 vdd.n273 gnd 0.005445f
C2754 vdd.n274 gnd 0.005445f
C2755 vdd.n275 gnd 0.002439f
C2756 vdd.n276 gnd 0.002304f
C2757 vdd.n277 gnd 0.004287f
C2758 vdd.n278 gnd 0.004287f
C2759 vdd.n279 gnd 0.002304f
C2760 vdd.n280 gnd 0.002439f
C2761 vdd.n281 gnd 0.005445f
C2762 vdd.n282 gnd 0.005445f
C2763 vdd.n283 gnd 0.002439f
C2764 vdd.n284 gnd 0.002304f
C2765 vdd.n285 gnd 0.004287f
C2766 vdd.n286 gnd 0.004287f
C2767 vdd.n287 gnd 0.002304f
C2768 vdd.n288 gnd 0.002439f
C2769 vdd.n289 gnd 0.005445f
C2770 vdd.n290 gnd 0.005445f
C2771 vdd.n291 gnd 0.012873f
C2772 vdd.n292 gnd 0.002371f
C2773 vdd.n293 gnd 0.002304f
C2774 vdd.n294 gnd 0.01108f
C2775 vdd.n295 gnd 0.007493f
C2776 vdd.n296 gnd 0.052314f
C2777 vdd.n297 gnd 0.204031f
C2778 vdd.n298 gnd 0.00647f
C2779 vdd.n299 gnd 0.008418f
C2780 vdd.n300 gnd 0.006775f
C2781 vdd.n301 gnd 0.006775f
C2782 vdd.n302 gnd 0.008418f
C2783 vdd.n303 gnd 0.008418f
C2784 vdd.n304 gnd 0.615084f
C2785 vdd.n305 gnd 0.008418f
C2786 vdd.n306 gnd 0.008418f
C2787 vdd.n307 gnd 0.008418f
C2788 vdd.n308 gnd 0.666699f
C2789 vdd.n309 gnd 0.008418f
C2790 vdd.n310 gnd 0.008418f
C2791 vdd.n311 gnd 0.008418f
C2792 vdd.n312 gnd 0.008418f
C2793 vdd.n313 gnd 0.006775f
C2794 vdd.n314 gnd 0.008418f
C2795 vdd.t124 gnd 0.430129f
C2796 vdd.n315 gnd 0.008418f
C2797 vdd.n316 gnd 0.008418f
C2798 vdd.n317 gnd 0.008418f
C2799 vdd.n318 gnd 0.860257f
C2800 vdd.n319 gnd 0.008418f
C2801 vdd.n320 gnd 0.008418f
C2802 vdd.n321 gnd 0.008418f
C2803 vdd.n322 gnd 0.008418f
C2804 vdd.n323 gnd 0.008418f
C2805 vdd.n324 gnd 0.006775f
C2806 vdd.n325 gnd 0.008418f
C2807 vdd.n326 gnd 0.008418f
C2808 vdd.n327 gnd 0.008418f
C2809 vdd.n328 gnd 0.020514f
C2810 vdd.n329 gnd 2.05602f
C2811 vdd.n330 gnd 0.020985f
C2812 vdd.n331 gnd 0.008418f
C2813 vdd.n332 gnd 0.008418f
C2814 vdd.n334 gnd 0.008418f
C2815 vdd.n335 gnd 0.008418f
C2816 vdd.n336 gnd 0.006775f
C2817 vdd.n337 gnd 0.006775f
C2818 vdd.n338 gnd 0.008418f
C2819 vdd.n339 gnd 0.008418f
C2820 vdd.n340 gnd 0.008418f
C2821 vdd.n341 gnd 0.008418f
C2822 vdd.n342 gnd 0.008418f
C2823 vdd.n343 gnd 0.008418f
C2824 vdd.n344 gnd 0.006775f
C2825 vdd.n346 gnd 0.008418f
C2826 vdd.n347 gnd 0.008418f
C2827 vdd.n348 gnd 0.008418f
C2828 vdd.n349 gnd 0.008418f
C2829 vdd.n350 gnd 0.008418f
C2830 vdd.n351 gnd 0.006775f
C2831 vdd.n353 gnd 0.008418f
C2832 vdd.n354 gnd 0.008418f
C2833 vdd.n355 gnd 0.008418f
C2834 vdd.n356 gnd 0.008418f
C2835 vdd.n357 gnd 0.008418f
C2836 vdd.n358 gnd 0.006775f
C2837 vdd.n360 gnd 0.008418f
C2838 vdd.n361 gnd 0.008418f
C2839 vdd.n362 gnd 0.008418f
C2840 vdd.n363 gnd 0.008418f
C2841 vdd.n364 gnd 0.005657f
C2842 vdd.t103 gnd 0.103561f
C2843 vdd.t102 gnd 0.110678f
C2844 vdd.t101 gnd 0.135249f
C2845 vdd.n365 gnd 0.17337f
C2846 vdd.n366 gnd 0.14634f
C2847 vdd.n368 gnd 0.008418f
C2848 vdd.n369 gnd 0.008418f
C2849 vdd.n370 gnd 0.006775f
C2850 vdd.n371 gnd 0.008418f
C2851 vdd.n373 gnd 0.008418f
C2852 vdd.n374 gnd 0.008418f
C2853 vdd.n375 gnd 0.008418f
C2854 vdd.n376 gnd 0.008418f
C2855 vdd.n377 gnd 0.006775f
C2856 vdd.n379 gnd 0.008418f
C2857 vdd.n380 gnd 0.008418f
C2858 vdd.n381 gnd 0.008418f
C2859 vdd.n382 gnd 0.008418f
C2860 vdd.n383 gnd 0.008418f
C2861 vdd.n384 gnd 0.006775f
C2862 vdd.n386 gnd 0.008418f
C2863 vdd.n387 gnd 0.008418f
C2864 vdd.n388 gnd 0.008418f
C2865 vdd.n389 gnd 0.008418f
C2866 vdd.n390 gnd 0.008418f
C2867 vdd.n391 gnd 0.006775f
C2868 vdd.n393 gnd 0.008418f
C2869 vdd.n394 gnd 0.008418f
C2870 vdd.n395 gnd 0.008418f
C2871 vdd.n396 gnd 0.008418f
C2872 vdd.n397 gnd 0.008418f
C2873 vdd.n398 gnd 0.006775f
C2874 vdd.n400 gnd 0.008418f
C2875 vdd.n401 gnd 0.008418f
C2876 vdd.n402 gnd 0.008418f
C2877 vdd.n403 gnd 0.008418f
C2878 vdd.n404 gnd 0.006708f
C2879 vdd.t100 gnd 0.103561f
C2880 vdd.t99 gnd 0.110678f
C2881 vdd.t98 gnd 0.135249f
C2882 vdd.n405 gnd 0.17337f
C2883 vdd.n406 gnd 0.14634f
C2884 vdd.n408 gnd 0.008418f
C2885 vdd.n409 gnd 0.008418f
C2886 vdd.n410 gnd 0.006775f
C2887 vdd.n411 gnd 0.008418f
C2888 vdd.n413 gnd 0.008418f
C2889 vdd.n414 gnd 0.008418f
C2890 vdd.n415 gnd 0.008418f
C2891 vdd.n416 gnd 0.008418f
C2892 vdd.n417 gnd 0.006775f
C2893 vdd.n419 gnd 0.008418f
C2894 vdd.n420 gnd 0.008418f
C2895 vdd.n421 gnd 0.008418f
C2896 vdd.n422 gnd 0.008418f
C2897 vdd.n423 gnd 0.008418f
C2898 vdd.n424 gnd 0.006775f
C2899 vdd.n426 gnd 0.008418f
C2900 vdd.n427 gnd 0.008418f
C2901 vdd.n428 gnd 0.008418f
C2902 vdd.n429 gnd 0.008418f
C2903 vdd.n430 gnd 0.008418f
C2904 vdd.n431 gnd 0.006775f
C2905 vdd.n433 gnd 0.008418f
C2906 vdd.n434 gnd 0.008418f
C2907 vdd.n435 gnd 0.008418f
C2908 vdd.n436 gnd 0.008418f
C2909 vdd.n437 gnd 0.008418f
C2910 vdd.n438 gnd 0.006775f
C2911 vdd.n440 gnd 0.008418f
C2912 vdd.n441 gnd 0.008418f
C2913 vdd.n442 gnd 0.008418f
C2914 vdd.n443 gnd 0.008418f
C2915 vdd.n444 gnd 0.008418f
C2916 vdd.n445 gnd 0.008418f
C2917 vdd.n446 gnd 0.006775f
C2918 vdd.n447 gnd 0.008418f
C2919 vdd.n448 gnd 0.008418f
C2920 vdd.n449 gnd 0.006775f
C2921 vdd.n450 gnd 0.008418f
C2922 vdd.n451 gnd 0.006775f
C2923 vdd.n452 gnd 0.008418f
C2924 vdd.n453 gnd 0.006775f
C2925 vdd.n454 gnd 0.008418f
C2926 vdd.n455 gnd 0.008418f
C2927 vdd.n456 gnd 0.46884f
C2928 vdd.t18 gnd 0.430129f
C2929 vdd.n457 gnd 0.008418f
C2930 vdd.n458 gnd 0.006775f
C2931 vdd.n459 gnd 0.008418f
C2932 vdd.n460 gnd 0.006775f
C2933 vdd.n461 gnd 0.008418f
C2934 vdd.t139 gnd 0.430129f
C2935 vdd.n462 gnd 0.008418f
C2936 vdd.n463 gnd 0.006775f
C2937 vdd.n464 gnd 0.008418f
C2938 vdd.n465 gnd 0.006775f
C2939 vdd.n466 gnd 0.008418f
C2940 vdd.t2 gnd 0.430129f
C2941 vdd.n467 gnd 0.537661f
C2942 vdd.n468 gnd 0.008418f
C2943 vdd.n469 gnd 0.006775f
C2944 vdd.n470 gnd 0.008418f
C2945 vdd.n471 gnd 0.006775f
C2946 vdd.n472 gnd 0.008418f
C2947 vdd.n473 gnd 0.860257f
C2948 vdd.n474 gnd 0.008418f
C2949 vdd.n475 gnd 0.006775f
C2950 vdd.n476 gnd 0.020514f
C2951 vdd.n477 gnd 0.005623f
C2952 vdd.n478 gnd 0.020514f
C2953 vdd.t37 gnd 0.430129f
C2954 vdd.n479 gnd 0.020514f
C2955 vdd.n480 gnd 0.005623f
C2956 vdd.n481 gnd 0.007239f
C2957 vdd.n482 gnd 0.006775f
C2958 vdd.n483 gnd 0.008418f
C2959 vdd.n484 gnd 8.74882f
C2960 vdd.n515 gnd 0.020985f
C2961 vdd.n516 gnd 1.18285f
C2962 vdd.n517 gnd 0.008418f
C2963 vdd.n518 gnd 0.006775f
C2964 vdd.n519 gnd 0.005387f
C2965 vdd.n520 gnd 0.026869f
C2966 vdd.n521 gnd 0.006775f
C2967 vdd.n522 gnd 0.008418f
C2968 vdd.n523 gnd 0.008418f
C2969 vdd.n524 gnd 0.008418f
C2970 vdd.n525 gnd 0.008418f
C2971 vdd.n526 gnd 0.008418f
C2972 vdd.n527 gnd 0.008418f
C2973 vdd.n528 gnd 0.008418f
C2974 vdd.n529 gnd 0.008418f
C2975 vdd.n530 gnd 0.008418f
C2976 vdd.n531 gnd 0.008418f
C2977 vdd.n532 gnd 0.008418f
C2978 vdd.n533 gnd 0.008418f
C2979 vdd.n534 gnd 0.008418f
C2980 vdd.n535 gnd 0.008418f
C2981 vdd.n536 gnd 0.005657f
C2982 vdd.n537 gnd 0.008418f
C2983 vdd.n538 gnd 0.008418f
C2984 vdd.n539 gnd 0.008418f
C2985 vdd.n540 gnd 0.008418f
C2986 vdd.n541 gnd 0.008418f
C2987 vdd.n542 gnd 0.008418f
C2988 vdd.n543 gnd 0.008418f
C2989 vdd.n544 gnd 0.008418f
C2990 vdd.n545 gnd 0.008418f
C2991 vdd.n546 gnd 0.008418f
C2992 vdd.n547 gnd 0.008418f
C2993 vdd.n548 gnd 0.008418f
C2994 vdd.n549 gnd 0.008418f
C2995 vdd.n550 gnd 0.008418f
C2996 vdd.n551 gnd 0.008418f
C2997 vdd.n552 gnd 0.008418f
C2998 vdd.n553 gnd 0.008418f
C2999 vdd.n554 gnd 0.008418f
C3000 vdd.n555 gnd 0.008418f
C3001 vdd.n556 gnd 0.006708f
C3002 vdd.t38 gnd 0.103561f
C3003 vdd.t39 gnd 0.110678f
C3004 vdd.t36 gnd 0.135249f
C3005 vdd.n557 gnd 0.17337f
C3006 vdd.n558 gnd 0.145662f
C3007 vdd.n559 gnd 0.008418f
C3008 vdd.n560 gnd 0.008418f
C3009 vdd.n561 gnd 0.008418f
C3010 vdd.n562 gnd 0.008418f
C3011 vdd.n563 gnd 0.008418f
C3012 vdd.n564 gnd 0.008418f
C3013 vdd.n565 gnd 0.008418f
C3014 vdd.n566 gnd 0.008418f
C3015 vdd.n567 gnd 0.008418f
C3016 vdd.n568 gnd 0.008418f
C3017 vdd.n569 gnd 0.008418f
C3018 vdd.n570 gnd 0.008418f
C3019 vdd.n571 gnd 0.008418f
C3020 vdd.n572 gnd 0.005387f
C3021 vdd.n575 gnd 0.005724f
C3022 vdd.n576 gnd 0.005724f
C3023 vdd.n577 gnd 0.005724f
C3024 vdd.n578 gnd 0.005724f
C3025 vdd.n579 gnd 0.005724f
C3026 vdd.n580 gnd 0.005724f
C3027 vdd.n582 gnd 0.005724f
C3028 vdd.n583 gnd 0.005724f
C3029 vdd.n585 gnd 0.005724f
C3030 vdd.n586 gnd 0.004167f
C3031 vdd.n588 gnd 0.005724f
C3032 vdd.t43 gnd 0.23131f
C3033 vdd.t42 gnd 0.236774f
C3034 vdd.t40 gnd 0.151008f
C3035 vdd.n589 gnd 0.081612f
C3036 vdd.n590 gnd 0.046293f
C3037 vdd.n591 gnd 0.008181f
C3038 vdd.n592 gnd 0.013123f
C3039 vdd.n594 gnd 0.005724f
C3040 vdd.n595 gnd 0.584975f
C3041 vdd.n596 gnd 0.012397f
C3042 vdd.n597 gnd 0.012397f
C3043 vdd.n598 gnd 0.005724f
C3044 vdd.n599 gnd 0.013193f
C3045 vdd.n600 gnd 0.005724f
C3046 vdd.n601 gnd 0.005724f
C3047 vdd.n602 gnd 0.005724f
C3048 vdd.n603 gnd 0.005724f
C3049 vdd.n604 gnd 0.005724f
C3050 vdd.n606 gnd 0.005724f
C3051 vdd.n607 gnd 0.005724f
C3052 vdd.n609 gnd 0.005724f
C3053 vdd.n610 gnd 0.005724f
C3054 vdd.n612 gnd 0.005724f
C3055 vdd.n613 gnd 0.005724f
C3056 vdd.n615 gnd 0.005724f
C3057 vdd.n616 gnd 0.005724f
C3058 vdd.n618 gnd 0.005724f
C3059 vdd.n619 gnd 0.005724f
C3060 vdd.n621 gnd 0.005724f
C3061 vdd.t70 gnd 0.23131f
C3062 vdd.t69 gnd 0.236774f
C3063 vdd.t68 gnd 0.151008f
C3064 vdd.n622 gnd 0.081612f
C3065 vdd.n623 gnd 0.046293f
C3066 vdd.n624 gnd 0.005724f
C3067 vdd.n626 gnd 0.005724f
C3068 vdd.n627 gnd 0.005724f
C3069 vdd.t41 gnd 0.292487f
C3070 vdd.n628 gnd 0.005724f
C3071 vdd.n629 gnd 0.005724f
C3072 vdd.n630 gnd 0.005724f
C3073 vdd.n631 gnd 0.005724f
C3074 vdd.n632 gnd 0.005724f
C3075 vdd.n633 gnd 0.584975f
C3076 vdd.n634 gnd 0.005724f
C3077 vdd.n635 gnd 0.005724f
C3078 vdd.n636 gnd 0.477443f
C3079 vdd.n637 gnd 0.005724f
C3080 vdd.n638 gnd 0.005724f
C3081 vdd.n639 gnd 0.005724f
C3082 vdd.n640 gnd 0.005724f
C3083 vdd.n641 gnd 0.584975f
C3084 vdd.n642 gnd 0.005724f
C3085 vdd.n643 gnd 0.005724f
C3086 vdd.n644 gnd 0.005724f
C3087 vdd.n645 gnd 0.005724f
C3088 vdd.n646 gnd 0.005724f
C3089 vdd.t177 gnd 0.292487f
C3090 vdd.n647 gnd 0.005724f
C3091 vdd.n648 gnd 0.005724f
C3092 vdd.n649 gnd 0.005724f
C3093 vdd.n650 gnd 0.005724f
C3094 vdd.n651 gnd 0.005724f
C3095 vdd.t183 gnd 0.292487f
C3096 vdd.n652 gnd 0.005724f
C3097 vdd.n653 gnd 0.005724f
C3098 vdd.n654 gnd 0.580674f
C3099 vdd.n655 gnd 0.005724f
C3100 vdd.n656 gnd 0.005724f
C3101 vdd.n657 gnd 0.005724f
C3102 vdd.t186 gnd 0.292487f
C3103 vdd.n658 gnd 0.005724f
C3104 vdd.n659 gnd 0.005724f
C3105 vdd.n660 gnd 0.451635f
C3106 vdd.n661 gnd 0.005724f
C3107 vdd.n662 gnd 0.005724f
C3108 vdd.n663 gnd 0.005724f
C3109 vdd.n664 gnd 0.391417f
C3110 vdd.n665 gnd 0.005724f
C3111 vdd.n666 gnd 0.005724f
C3112 vdd.n667 gnd 0.322596f
C3113 vdd.n668 gnd 0.005724f
C3114 vdd.n669 gnd 0.005724f
C3115 vdd.n670 gnd 0.005724f
C3116 vdd.n671 gnd 0.481744f
C3117 vdd.n672 gnd 0.005724f
C3118 vdd.n673 gnd 0.005724f
C3119 vdd.t156 gnd 0.292487f
C3120 vdd.n674 gnd 0.005724f
C3121 vdd.t56 gnd 0.236774f
C3122 vdd.t54 gnd 0.151008f
C3123 vdd.t57 gnd 0.236774f
C3124 vdd.n675 gnd 0.133077f
C3125 vdd.n676 gnd 0.005724f
C3126 vdd.n677 gnd 0.005724f
C3127 vdd.n678 gnd 0.584975f
C3128 vdd.n679 gnd 0.005724f
C3129 vdd.n680 gnd 0.005724f
C3130 vdd.t55 gnd 0.227968f
C3131 vdd.t158 gnd 0.103231f
C3132 vdd.n681 gnd 0.005724f
C3133 vdd.n682 gnd 0.005724f
C3134 vdd.n683 gnd 0.005724f
C3135 vdd.t169 gnd 0.292487f
C3136 vdd.n684 gnd 0.005724f
C3137 vdd.n685 gnd 0.005724f
C3138 vdd.n686 gnd 0.005724f
C3139 vdd.n687 gnd 0.005724f
C3140 vdd.n688 gnd 0.005724f
C3141 vdd.t187 gnd 0.292487f
C3142 vdd.n689 gnd 0.005724f
C3143 vdd.n690 gnd 0.005724f
C3144 vdd.n691 gnd 0.520456f
C3145 vdd.n692 gnd 0.005724f
C3146 vdd.n693 gnd 0.005724f
C3147 vdd.n694 gnd 0.005724f
C3148 vdd.n695 gnd 0.322596f
C3149 vdd.n696 gnd 0.005724f
C3150 vdd.n697 gnd 0.005724f
C3151 vdd.t165 gnd 0.292487f
C3152 vdd.n698 gnd 0.005724f
C3153 vdd.n699 gnd 0.005724f
C3154 vdd.n700 gnd 0.005724f
C3155 vdd.n701 gnd 0.451635f
C3156 vdd.n702 gnd 0.005724f
C3157 vdd.n703 gnd 0.005724f
C3158 vdd.t149 gnd 0.215064f
C3159 vdd.t199 gnd 0.262378f
C3160 vdd.n704 gnd 0.005724f
C3161 vdd.n705 gnd 0.005724f
C3162 vdd.n706 gnd 0.005724f
C3163 vdd.t195 gnd 0.292487f
C3164 vdd.n707 gnd 0.005724f
C3165 vdd.n708 gnd 0.005724f
C3166 vdd.t188 gnd 0.292487f
C3167 vdd.n709 gnd 0.005724f
C3168 vdd.n710 gnd 0.005724f
C3169 vdd.n711 gnd 0.005724f
C3170 vdd.t175 gnd 0.292487f
C3171 vdd.n712 gnd 0.005724f
C3172 vdd.n713 gnd 0.005724f
C3173 vdd.t153 gnd 0.292487f
C3174 vdd.n714 gnd 0.005724f
C3175 vdd.n715 gnd 0.005724f
C3176 vdd.n716 gnd 0.005724f
C3177 vdd.n717 gnd 0.584975f
C3178 vdd.n718 gnd 0.005724f
C3179 vdd.n719 gnd 0.005724f
C3180 vdd.n720 gnd 0.404321f
C3181 vdd.n721 gnd 0.005724f
C3182 vdd.n722 gnd 0.005724f
C3183 vdd.n723 gnd 0.005724f
C3184 vdd.t154 gnd 0.292487f
C3185 vdd.n724 gnd 0.005724f
C3186 vdd.n725 gnd 0.005724f
C3187 vdd.n726 gnd 0.005724f
C3188 vdd.n727 gnd 0.005724f
C3189 vdd.n728 gnd 0.005724f
C3190 vdd.t181 gnd 0.292487f
C3191 vdd.n729 gnd 0.005724f
C3192 vdd.n730 gnd 0.005724f
C3193 vdd.t79 gnd 0.292487f
C3194 vdd.n731 gnd 0.005724f
C3195 vdd.n732 gnd 0.013193f
C3196 vdd.n733 gnd 0.013193f
C3197 vdd.t179 gnd 0.516154f
C3198 vdd.n734 gnd 0.012397f
C3199 vdd.n735 gnd 0.012397f
C3200 vdd.n736 gnd 0.326898f
C3201 vdd.n737 gnd 0.013193f
C3202 vdd.n738 gnd 0.005724f
C3203 vdd.n739 gnd 0.005724f
C3204 vdd.t191 gnd 0.516154f
C3205 vdd.n757 gnd 0.013193f
C3206 vdd.n775 gnd 0.012397f
C3207 vdd.n776 gnd 0.005724f
C3208 vdd.n777 gnd 0.012397f
C3209 vdd.t94 gnd 0.23131f
C3210 vdd.t93 gnd 0.236774f
C3211 vdd.t92 gnd 0.151008f
C3212 vdd.n778 gnd 0.081612f
C3213 vdd.n779 gnd 0.046293f
C3214 vdd.n780 gnd 0.013123f
C3215 vdd.n781 gnd 0.005724f
C3216 vdd.n782 gnd 0.326898f
C3217 vdd.n783 gnd 0.012397f
C3218 vdd.n784 gnd 0.005724f
C3219 vdd.n785 gnd 0.013193f
C3220 vdd.n786 gnd 0.005724f
C3221 vdd.t77 gnd 0.23131f
C3222 vdd.t76 gnd 0.236774f
C3223 vdd.t74 gnd 0.151008f
C3224 vdd.n787 gnd 0.081612f
C3225 vdd.n788 gnd 0.046293f
C3226 vdd.n789 gnd 0.008181f
C3227 vdd.n790 gnd 0.005724f
C3228 vdd.n791 gnd 0.005724f
C3229 vdd.t75 gnd 0.292487f
C3230 vdd.n792 gnd 0.005724f
C3231 vdd.t193 gnd 0.292487f
C3232 vdd.n793 gnd 0.005724f
C3233 vdd.n794 gnd 0.005724f
C3234 vdd.n795 gnd 0.005724f
C3235 vdd.n796 gnd 0.005724f
C3236 vdd.n797 gnd 0.005724f
C3237 vdd.n798 gnd 0.584975f
C3238 vdd.n799 gnd 0.005724f
C3239 vdd.n800 gnd 0.005724f
C3240 vdd.t167 gnd 0.292487f
C3241 vdd.n801 gnd 0.005724f
C3242 vdd.n802 gnd 0.005724f
C3243 vdd.n803 gnd 0.005724f
C3244 vdd.n804 gnd 0.005724f
C3245 vdd.n805 gnd 0.404321f
C3246 vdd.n806 gnd 0.005724f
C3247 vdd.n807 gnd 0.005724f
C3248 vdd.n808 gnd 0.005724f
C3249 vdd.n809 gnd 0.005724f
C3250 vdd.n810 gnd 0.005724f
C3251 vdd.t150 gnd 0.292487f
C3252 vdd.n811 gnd 0.005724f
C3253 vdd.n812 gnd 0.005724f
C3254 vdd.t184 gnd 0.292487f
C3255 vdd.n813 gnd 0.005724f
C3256 vdd.n814 gnd 0.005724f
C3257 vdd.n815 gnd 0.005724f
C3258 vdd.t174 gnd 0.292487f
C3259 vdd.n816 gnd 0.005724f
C3260 vdd.n817 gnd 0.005724f
C3261 vdd.t151 gnd 0.292487f
C3262 vdd.n818 gnd 0.005724f
C3263 vdd.n819 gnd 0.005724f
C3264 vdd.n820 gnd 0.005724f
C3265 vdd.t170 gnd 0.262378f
C3266 vdd.n821 gnd 0.005724f
C3267 vdd.n822 gnd 0.005724f
C3268 vdd.n823 gnd 0.451635f
C3269 vdd.n824 gnd 0.005724f
C3270 vdd.n825 gnd 0.005724f
C3271 vdd.n826 gnd 0.005724f
C3272 vdd.t189 gnd 0.292487f
C3273 vdd.n827 gnd 0.005724f
C3274 vdd.n828 gnd 0.005724f
C3275 vdd.t159 gnd 0.215064f
C3276 vdd.n829 gnd 0.322596f
C3277 vdd.n830 gnd 0.005724f
C3278 vdd.n831 gnd 0.005724f
C3279 vdd.n832 gnd 0.005724f
C3280 vdd.n833 gnd 0.520456f
C3281 vdd.n834 gnd 0.005724f
C3282 vdd.n835 gnd 0.005724f
C3283 vdd.t197 gnd 0.292487f
C3284 vdd.n836 gnd 0.005724f
C3285 vdd.n837 gnd 0.005724f
C3286 vdd.n838 gnd 0.005724f
C3287 vdd.n839 gnd 0.584975f
C3288 vdd.n840 gnd 0.005724f
C3289 vdd.n841 gnd 0.005724f
C3290 vdd.t164 gnd 0.292487f
C3291 vdd.n842 gnd 0.005724f
C3292 vdd.n843 gnd 0.005724f
C3293 vdd.n844 gnd 0.005724f
C3294 vdd.t157 gnd 0.103231f
C3295 vdd.n845 gnd 0.005724f
C3296 vdd.n846 gnd 0.005724f
C3297 vdd.n847 gnd 0.005724f
C3298 vdd.t87 gnd 0.236774f
C3299 vdd.t85 gnd 0.151008f
C3300 vdd.t88 gnd 0.236774f
C3301 vdd.n848 gnd 0.133077f
C3302 vdd.n849 gnd 0.005724f
C3303 vdd.n850 gnd 0.005724f
C3304 vdd.t178 gnd 0.292487f
C3305 vdd.n851 gnd 0.005724f
C3306 vdd.n852 gnd 0.005724f
C3307 vdd.t86 gnd 0.227968f
C3308 vdd.n853 gnd 0.481744f
C3309 vdd.n854 gnd 0.005724f
C3310 vdd.n855 gnd 0.005724f
C3311 vdd.n856 gnd 0.005724f
C3312 vdd.n857 gnd 0.322596f
C3313 vdd.n858 gnd 0.005724f
C3314 vdd.n859 gnd 0.005724f
C3315 vdd.n860 gnd 0.391417f
C3316 vdd.n861 gnd 0.005724f
C3317 vdd.n862 gnd 0.005724f
C3318 vdd.n863 gnd 0.005724f
C3319 vdd.n864 gnd 0.451635f
C3320 vdd.n865 gnd 0.005724f
C3321 vdd.n866 gnd 0.005724f
C3322 vdd.t161 gnd 0.292487f
C3323 vdd.n867 gnd 0.005724f
C3324 vdd.n868 gnd 0.005724f
C3325 vdd.n869 gnd 0.005724f
C3326 vdd.n870 gnd 0.580674f
C3327 vdd.n871 gnd 0.005724f
C3328 vdd.n872 gnd 0.005724f
C3329 vdd.t160 gnd 0.292487f
C3330 vdd.n873 gnd 0.005724f
C3331 vdd.n874 gnd 0.005724f
C3332 vdd.n875 gnd 0.005724f
C3333 vdd.n876 gnd 0.584975f
C3334 vdd.n877 gnd 0.005724f
C3335 vdd.n878 gnd 0.005724f
C3336 vdd.t198 gnd 0.292487f
C3337 vdd.n879 gnd 0.005724f
C3338 vdd.n880 gnd 0.005724f
C3339 vdd.n881 gnd 0.005724f
C3340 vdd.n882 gnd 0.584975f
C3341 vdd.n883 gnd 0.005724f
C3342 vdd.n884 gnd 0.005724f
C3343 vdd.n885 gnd 0.005724f
C3344 vdd.n886 gnd 0.005724f
C3345 vdd.n887 gnd 0.005724f
C3346 vdd.n888 gnd 0.477443f
C3347 vdd.n889 gnd 0.005724f
C3348 vdd.n890 gnd 0.005724f
C3349 vdd.n891 gnd 0.005724f
C3350 vdd.n892 gnd 0.005724f
C3351 vdd.n893 gnd 0.005724f
C3352 vdd.n894 gnd 0.584975f
C3353 vdd.n895 gnd 0.005724f
C3354 vdd.n896 gnd 0.005724f
C3355 vdd.t45 gnd 0.292487f
C3356 vdd.n897 gnd 0.005724f
C3357 vdd.n898 gnd 0.013193f
C3358 vdd.n899 gnd 0.013193f
C3359 vdd.n900 gnd 8.74882f
C3360 vdd.n901 gnd 0.012397f
C3361 vdd.n902 gnd 0.012397f
C3362 vdd.n903 gnd 0.013193f
C3363 vdd.n904 gnd 0.005724f
C3364 vdd.n906 gnd 0.005724f
C3365 vdd.n907 gnd 0.005724f
C3366 vdd.n908 gnd 0.005724f
C3367 vdd.n909 gnd 0.005724f
C3368 vdd.n910 gnd 0.005724f
C3369 vdd.n911 gnd 0.005724f
C3370 vdd.n912 gnd 0.030118f
C3371 vdd.n913 gnd 0.005724f
C3372 vdd.n914 gnd 0.005724f
C3373 vdd.n915 gnd 0.005724f
C3374 vdd.n916 gnd 0.005724f
C3375 vdd.n917 gnd 0.005724f
C3376 vdd.n918 gnd 0.005724f
C3377 vdd.n919 gnd 0.005724f
C3378 vdd.t96 gnd 0.23131f
C3379 vdd.t97 gnd 0.236774f
C3380 vdd.t95 gnd 0.151008f
C3381 vdd.n920 gnd 0.081612f
C3382 vdd.n921 gnd 0.046293f
C3383 vdd.n922 gnd 0.005724f
C3384 vdd.n923 gnd 0.005724f
C3385 vdd.n924 gnd 0.005724f
C3386 vdd.n925 gnd 0.005724f
C3387 vdd.t46 gnd 0.23131f
C3388 vdd.t47 gnd 0.236774f
C3389 vdd.t44 gnd 0.151008f
C3390 vdd.n926 gnd 0.081612f
C3391 vdd.n927 gnd 0.046293f
C3392 vdd.n928 gnd 0.005724f
C3393 vdd.n929 gnd 0.005724f
C3394 vdd.n930 gnd 0.005724f
C3395 vdd.n931 gnd 0.005724f
C3396 vdd.n932 gnd 0.005724f
C3397 vdd.n933 gnd 0.005724f
C3398 vdd.n934 gnd 0.005387f
C3399 vdd.n937 gnd 0.020985f
C3400 vdd.n938 gnd 0.006775f
C3401 vdd.n939 gnd 0.008418f
C3402 vdd.n941 gnd 0.008418f
C3403 vdd.n942 gnd 0.005623f
C3404 vdd.t62 gnd 0.430129f
C3405 vdd.n943 gnd 9.09292f
C3406 vdd.n944 gnd 0.008418f
C3407 vdd.n945 gnd 0.020985f
C3408 vdd.n946 gnd 0.006775f
C3409 vdd.n947 gnd 0.008418f
C3410 vdd.n948 gnd 0.006775f
C3411 vdd.n949 gnd 0.008418f
C3412 vdd.n950 gnd 0.860257f
C3413 vdd.n951 gnd 0.008418f
C3414 vdd.n952 gnd 0.006775f
C3415 vdd.n953 gnd 0.006775f
C3416 vdd.n954 gnd 0.008418f
C3417 vdd.n955 gnd 0.006775f
C3418 vdd.n956 gnd 0.008418f
C3419 vdd.t15 gnd 0.430129f
C3420 vdd.n957 gnd 0.008418f
C3421 vdd.n958 gnd 0.006775f
C3422 vdd.n959 gnd 0.008418f
C3423 vdd.n960 gnd 0.006775f
C3424 vdd.n961 gnd 0.008418f
C3425 vdd.t21 gnd 0.430129f
C3426 vdd.n962 gnd 0.008418f
C3427 vdd.n963 gnd 0.006775f
C3428 vdd.n964 gnd 0.008418f
C3429 vdd.n965 gnd 0.006775f
C3430 vdd.n966 gnd 0.008418f
C3431 vdd.n967 gnd 0.675302f
C3432 vdd.n968 gnd 0.714014f
C3433 vdd.t0 gnd 0.430129f
C3434 vdd.n969 gnd 0.008418f
C3435 vdd.n970 gnd 0.006775f
C3436 vdd.n971 gnd 0.00462f
C3437 vdd.n972 gnd 0.004287f
C3438 vdd.n973 gnd 0.002371f
C3439 vdd.n974 gnd 0.005445f
C3440 vdd.n975 gnd 0.002304f
C3441 vdd.n976 gnd 0.002439f
C3442 vdd.n977 gnd 0.004287f
C3443 vdd.n978 gnd 0.002304f
C3444 vdd.n979 gnd 0.005445f
C3445 vdd.n980 gnd 0.002439f
C3446 vdd.n981 gnd 0.004287f
C3447 vdd.n982 gnd 0.002304f
C3448 vdd.n983 gnd 0.004084f
C3449 vdd.n984 gnd 0.004096f
C3450 vdd.t203 gnd 0.011698f
C3451 vdd.n985 gnd 0.026027f
C3452 vdd.n986 gnd 0.135453f
C3453 vdd.n987 gnd 0.002304f
C3454 vdd.n988 gnd 0.002439f
C3455 vdd.n989 gnd 0.005445f
C3456 vdd.n990 gnd 0.005445f
C3457 vdd.n991 gnd 0.002439f
C3458 vdd.n992 gnd 0.002304f
C3459 vdd.n993 gnd 0.004287f
C3460 vdd.n994 gnd 0.004287f
C3461 vdd.n995 gnd 0.002304f
C3462 vdd.n996 gnd 0.002439f
C3463 vdd.n997 gnd 0.005445f
C3464 vdd.n998 gnd 0.005445f
C3465 vdd.n999 gnd 0.002439f
C3466 vdd.n1000 gnd 0.002304f
C3467 vdd.n1001 gnd 0.004287f
C3468 vdd.n1002 gnd 0.004287f
C3469 vdd.n1003 gnd 0.002304f
C3470 vdd.n1004 gnd 0.002439f
C3471 vdd.n1005 gnd 0.005445f
C3472 vdd.n1006 gnd 0.005445f
C3473 vdd.n1007 gnd 0.012873f
C3474 vdd.n1008 gnd 0.002371f
C3475 vdd.n1009 gnd 0.002304f
C3476 vdd.n1010 gnd 0.01108f
C3477 vdd.n1011 gnd 0.007736f
C3478 vdd.t134 gnd 0.027101f
C3479 vdd.t204 gnd 0.027101f
C3480 vdd.n1012 gnd 0.186258f
C3481 vdd.n1013 gnd 0.146463f
C3482 vdd.t123 gnd 0.027101f
C3483 vdd.t119 gnd 0.027101f
C3484 vdd.n1014 gnd 0.186258f
C3485 vdd.n1015 gnd 0.118195f
C3486 vdd.t131 gnd 0.027101f
C3487 vdd.t130 gnd 0.027101f
C3488 vdd.n1016 gnd 0.186258f
C3489 vdd.n1017 gnd 0.118195f
C3490 vdd.n1018 gnd 0.00462f
C3491 vdd.n1019 gnd 0.004287f
C3492 vdd.n1020 gnd 0.002371f
C3493 vdd.n1021 gnd 0.005445f
C3494 vdd.n1022 gnd 0.002304f
C3495 vdd.n1023 gnd 0.002439f
C3496 vdd.n1024 gnd 0.004287f
C3497 vdd.n1025 gnd 0.002304f
C3498 vdd.n1026 gnd 0.005445f
C3499 vdd.n1027 gnd 0.002439f
C3500 vdd.n1028 gnd 0.004287f
C3501 vdd.n1029 gnd 0.002304f
C3502 vdd.n1030 gnd 0.004084f
C3503 vdd.n1031 gnd 0.004096f
C3504 vdd.t144 gnd 0.011698f
C3505 vdd.n1032 gnd 0.026027f
C3506 vdd.n1033 gnd 0.135453f
C3507 vdd.n1034 gnd 0.002304f
C3508 vdd.n1035 gnd 0.002439f
C3509 vdd.n1036 gnd 0.005445f
C3510 vdd.n1037 gnd 0.005445f
C3511 vdd.n1038 gnd 0.002439f
C3512 vdd.n1039 gnd 0.002304f
C3513 vdd.n1040 gnd 0.004287f
C3514 vdd.n1041 gnd 0.004287f
C3515 vdd.n1042 gnd 0.002304f
C3516 vdd.n1043 gnd 0.002439f
C3517 vdd.n1044 gnd 0.005445f
C3518 vdd.n1045 gnd 0.005445f
C3519 vdd.n1046 gnd 0.002439f
C3520 vdd.n1047 gnd 0.002304f
C3521 vdd.n1048 gnd 0.004287f
C3522 vdd.n1049 gnd 0.004287f
C3523 vdd.n1050 gnd 0.002304f
C3524 vdd.n1051 gnd 0.002439f
C3525 vdd.n1052 gnd 0.005445f
C3526 vdd.n1053 gnd 0.005445f
C3527 vdd.n1054 gnd 0.012873f
C3528 vdd.n1055 gnd 0.002371f
C3529 vdd.n1056 gnd 0.002304f
C3530 vdd.n1057 gnd 0.01108f
C3531 vdd.n1058 gnd 0.007493f
C3532 vdd.n1059 gnd 0.087938f
C3533 vdd.n1060 gnd 0.00462f
C3534 vdd.n1061 gnd 0.004287f
C3535 vdd.n1062 gnd 0.002371f
C3536 vdd.n1063 gnd 0.005445f
C3537 vdd.n1064 gnd 0.002304f
C3538 vdd.n1065 gnd 0.002439f
C3539 vdd.n1066 gnd 0.004287f
C3540 vdd.n1067 gnd 0.002304f
C3541 vdd.n1068 gnd 0.005445f
C3542 vdd.n1069 gnd 0.002439f
C3543 vdd.n1070 gnd 0.004287f
C3544 vdd.n1071 gnd 0.002304f
C3545 vdd.n1072 gnd 0.004084f
C3546 vdd.n1073 gnd 0.004096f
C3547 vdd.t112 gnd 0.011698f
C3548 vdd.n1074 gnd 0.026027f
C3549 vdd.n1075 gnd 0.135453f
C3550 vdd.n1076 gnd 0.002304f
C3551 vdd.n1077 gnd 0.002439f
C3552 vdd.n1078 gnd 0.005445f
C3553 vdd.n1079 gnd 0.005445f
C3554 vdd.n1080 gnd 0.002439f
C3555 vdd.n1081 gnd 0.002304f
C3556 vdd.n1082 gnd 0.004287f
C3557 vdd.n1083 gnd 0.004287f
C3558 vdd.n1084 gnd 0.002304f
C3559 vdd.n1085 gnd 0.002439f
C3560 vdd.n1086 gnd 0.005445f
C3561 vdd.n1087 gnd 0.005445f
C3562 vdd.n1088 gnd 0.002439f
C3563 vdd.n1089 gnd 0.002304f
C3564 vdd.n1090 gnd 0.004287f
C3565 vdd.n1091 gnd 0.004287f
C3566 vdd.n1092 gnd 0.002304f
C3567 vdd.n1093 gnd 0.002439f
C3568 vdd.n1094 gnd 0.005445f
C3569 vdd.n1095 gnd 0.005445f
C3570 vdd.n1096 gnd 0.012873f
C3571 vdd.n1097 gnd 0.002371f
C3572 vdd.n1098 gnd 0.002304f
C3573 vdd.n1099 gnd 0.01108f
C3574 vdd.n1100 gnd 0.007736f
C3575 vdd.t1 gnd 0.027101f
C3576 vdd.t120 gnd 0.027101f
C3577 vdd.n1101 gnd 0.186258f
C3578 vdd.n1102 gnd 0.146463f
C3579 vdd.t107 gnd 0.027101f
C3580 vdd.t7 gnd 0.027101f
C3581 vdd.n1103 gnd 0.186258f
C3582 vdd.n1104 gnd 0.118195f
C3583 vdd.t205 gnd 0.027101f
C3584 vdd.t147 gnd 0.027101f
C3585 vdd.n1105 gnd 0.186258f
C3586 vdd.n1106 gnd 0.118195f
C3587 vdd.n1107 gnd 0.00462f
C3588 vdd.n1108 gnd 0.004287f
C3589 vdd.n1109 gnd 0.002371f
C3590 vdd.n1110 gnd 0.005445f
C3591 vdd.n1111 gnd 0.002304f
C3592 vdd.n1112 gnd 0.002439f
C3593 vdd.n1113 gnd 0.004287f
C3594 vdd.n1114 gnd 0.002304f
C3595 vdd.n1115 gnd 0.005445f
C3596 vdd.n1116 gnd 0.002439f
C3597 vdd.n1117 gnd 0.004287f
C3598 vdd.n1118 gnd 0.002304f
C3599 vdd.n1119 gnd 0.004084f
C3600 vdd.n1120 gnd 0.004096f
C3601 vdd.t201 gnd 0.011698f
C3602 vdd.n1121 gnd 0.026027f
C3603 vdd.n1122 gnd 0.135453f
C3604 vdd.n1123 gnd 0.002304f
C3605 vdd.n1124 gnd 0.002439f
C3606 vdd.n1125 gnd 0.005445f
C3607 vdd.n1126 gnd 0.005445f
C3608 vdd.n1127 gnd 0.002439f
C3609 vdd.n1128 gnd 0.002304f
C3610 vdd.n1129 gnd 0.004287f
C3611 vdd.n1130 gnd 0.004287f
C3612 vdd.n1131 gnd 0.002304f
C3613 vdd.n1132 gnd 0.002439f
C3614 vdd.n1133 gnd 0.005445f
C3615 vdd.n1134 gnd 0.005445f
C3616 vdd.n1135 gnd 0.002439f
C3617 vdd.n1136 gnd 0.002304f
C3618 vdd.n1137 gnd 0.004287f
C3619 vdd.n1138 gnd 0.004287f
C3620 vdd.n1139 gnd 0.002304f
C3621 vdd.n1140 gnd 0.002439f
C3622 vdd.n1141 gnd 0.005445f
C3623 vdd.n1142 gnd 0.005445f
C3624 vdd.n1143 gnd 0.012873f
C3625 vdd.n1144 gnd 0.002371f
C3626 vdd.n1145 gnd 0.002304f
C3627 vdd.n1146 gnd 0.01108f
C3628 vdd.n1147 gnd 0.007493f
C3629 vdd.n1148 gnd 0.052314f
C3630 vdd.n1149 gnd 0.188501f
C3631 vdd.n1150 gnd 0.00462f
C3632 vdd.n1151 gnd 0.004287f
C3633 vdd.n1152 gnd 0.002371f
C3634 vdd.n1153 gnd 0.005445f
C3635 vdd.n1154 gnd 0.002304f
C3636 vdd.n1155 gnd 0.002439f
C3637 vdd.n1156 gnd 0.004287f
C3638 vdd.n1157 gnd 0.002304f
C3639 vdd.n1158 gnd 0.005445f
C3640 vdd.n1159 gnd 0.002439f
C3641 vdd.n1160 gnd 0.004287f
C3642 vdd.n1161 gnd 0.002304f
C3643 vdd.n1162 gnd 0.004084f
C3644 vdd.n1163 gnd 0.004096f
C3645 vdd.t16 gnd 0.011698f
C3646 vdd.n1164 gnd 0.026027f
C3647 vdd.n1165 gnd 0.135453f
C3648 vdd.n1166 gnd 0.002304f
C3649 vdd.n1167 gnd 0.002439f
C3650 vdd.n1168 gnd 0.005445f
C3651 vdd.n1169 gnd 0.005445f
C3652 vdd.n1170 gnd 0.002439f
C3653 vdd.n1171 gnd 0.002304f
C3654 vdd.n1172 gnd 0.004287f
C3655 vdd.n1173 gnd 0.004287f
C3656 vdd.n1174 gnd 0.002304f
C3657 vdd.n1175 gnd 0.002439f
C3658 vdd.n1176 gnd 0.005445f
C3659 vdd.n1177 gnd 0.005445f
C3660 vdd.n1178 gnd 0.002439f
C3661 vdd.n1179 gnd 0.002304f
C3662 vdd.n1180 gnd 0.004287f
C3663 vdd.n1181 gnd 0.004287f
C3664 vdd.n1182 gnd 0.002304f
C3665 vdd.n1183 gnd 0.002439f
C3666 vdd.n1184 gnd 0.005445f
C3667 vdd.n1185 gnd 0.005445f
C3668 vdd.n1186 gnd 0.012873f
C3669 vdd.n1187 gnd 0.002371f
C3670 vdd.n1188 gnd 0.002304f
C3671 vdd.n1189 gnd 0.01108f
C3672 vdd.n1190 gnd 0.007736f
C3673 vdd.t17 gnd 0.027101f
C3674 vdd.t22 gnd 0.027101f
C3675 vdd.n1191 gnd 0.186258f
C3676 vdd.n1192 gnd 0.146463f
C3677 vdd.t138 gnd 0.027101f
C3678 vdd.t202 gnd 0.027101f
C3679 vdd.n1193 gnd 0.186258f
C3680 vdd.n1194 gnd 0.118195f
C3681 vdd.t127 gnd 0.027101f
C3682 vdd.t13 gnd 0.027101f
C3683 vdd.n1195 gnd 0.186258f
C3684 vdd.n1196 gnd 0.118195f
C3685 vdd.n1197 gnd 0.00462f
C3686 vdd.n1198 gnd 0.004287f
C3687 vdd.n1199 gnd 0.002371f
C3688 vdd.n1200 gnd 0.005445f
C3689 vdd.n1201 gnd 0.002304f
C3690 vdd.n1202 gnd 0.002439f
C3691 vdd.n1203 gnd 0.004287f
C3692 vdd.n1204 gnd 0.002304f
C3693 vdd.n1205 gnd 0.005445f
C3694 vdd.n1206 gnd 0.002439f
C3695 vdd.n1207 gnd 0.004287f
C3696 vdd.n1208 gnd 0.002304f
C3697 vdd.n1209 gnd 0.004084f
C3698 vdd.n1210 gnd 0.004096f
C3699 vdd.t122 gnd 0.011698f
C3700 vdd.n1211 gnd 0.026027f
C3701 vdd.n1212 gnd 0.135453f
C3702 vdd.n1213 gnd 0.002304f
C3703 vdd.n1214 gnd 0.002439f
C3704 vdd.n1215 gnd 0.005445f
C3705 vdd.n1216 gnd 0.005445f
C3706 vdd.n1217 gnd 0.002439f
C3707 vdd.n1218 gnd 0.002304f
C3708 vdd.n1219 gnd 0.004287f
C3709 vdd.n1220 gnd 0.004287f
C3710 vdd.n1221 gnd 0.002304f
C3711 vdd.n1222 gnd 0.002439f
C3712 vdd.n1223 gnd 0.005445f
C3713 vdd.n1224 gnd 0.005445f
C3714 vdd.n1225 gnd 0.002439f
C3715 vdd.n1226 gnd 0.002304f
C3716 vdd.n1227 gnd 0.004287f
C3717 vdd.n1228 gnd 0.004287f
C3718 vdd.n1229 gnd 0.002304f
C3719 vdd.n1230 gnd 0.002439f
C3720 vdd.n1231 gnd 0.005445f
C3721 vdd.n1232 gnd 0.005445f
C3722 vdd.n1233 gnd 0.012873f
C3723 vdd.n1234 gnd 0.002371f
C3724 vdd.n1235 gnd 0.002304f
C3725 vdd.n1236 gnd 0.01108f
C3726 vdd.n1237 gnd 0.007493f
C3727 vdd.n1238 gnd 0.052314f
C3728 vdd.n1239 gnd 0.204031f
C3729 vdd.n1240 gnd 1.9179f
C3730 vdd.n1241 gnd 0.496513f
C3731 vdd.n1242 gnd 0.006775f
C3732 vdd.n1243 gnd 0.008418f
C3733 vdd.n1244 gnd 0.529058f
C3734 vdd.n1245 gnd 0.008418f
C3735 vdd.n1246 gnd 0.006775f
C3736 vdd.n1247 gnd 0.008418f
C3737 vdd.n1248 gnd 0.006775f
C3738 vdd.n1249 gnd 0.008418f
C3739 vdd.t12 gnd 0.430129f
C3740 vdd.t106 gnd 0.430129f
C3741 vdd.n1250 gnd 0.008418f
C3742 vdd.n1251 gnd 0.006775f
C3743 vdd.n1252 gnd 0.008418f
C3744 vdd.n1253 gnd 0.006775f
C3745 vdd.n1254 gnd 0.008418f
C3746 vdd.t126 gnd 0.430129f
C3747 vdd.n1255 gnd 0.008418f
C3748 vdd.n1256 gnd 0.006775f
C3749 vdd.n1257 gnd 0.008418f
C3750 vdd.n1258 gnd 0.006775f
C3751 vdd.n1259 gnd 0.008418f
C3752 vdd.t121 gnd 0.430129f
C3753 vdd.n1260 gnd 0.623687f
C3754 vdd.n1261 gnd 0.008418f
C3755 vdd.n1262 gnd 0.006775f
C3756 vdd.n1263 gnd 0.008418f
C3757 vdd.n1264 gnd 0.006775f
C3758 vdd.n1265 gnd 0.008418f
C3759 vdd.n1266 gnd 0.860257f
C3760 vdd.n1267 gnd 0.008418f
C3761 vdd.n1268 gnd 0.006775f
C3762 vdd.n1269 gnd 0.020514f
C3763 vdd.n1270 gnd 0.005623f
C3764 vdd.n1271 gnd 0.020514f
C3765 vdd.t33 gnd 0.430129f
C3766 vdd.n1272 gnd 0.020514f
C3767 vdd.n1273 gnd 0.005623f
C3768 vdd.n1274 gnd 0.008418f
C3769 vdd.n1275 gnd 0.006775f
C3770 vdd.n1276 gnd 0.008418f
C3771 vdd.n1307 gnd 0.020985f
C3772 vdd.n1308 gnd 1.26888f
C3773 vdd.n1309 gnd 0.008418f
C3774 vdd.n1310 gnd 0.006775f
C3775 vdd.n1311 gnd 0.008418f
C3776 vdd.n1312 gnd 0.008418f
C3777 vdd.n1313 gnd 0.008418f
C3778 vdd.n1314 gnd 0.008418f
C3779 vdd.n1315 gnd 0.008418f
C3780 vdd.n1316 gnd 0.006775f
C3781 vdd.n1317 gnd 0.008418f
C3782 vdd.n1318 gnd 0.008418f
C3783 vdd.n1319 gnd 0.008418f
C3784 vdd.n1320 gnd 0.008418f
C3785 vdd.n1321 gnd 0.008418f
C3786 vdd.n1322 gnd 0.006775f
C3787 vdd.n1323 gnd 0.008418f
C3788 vdd.n1324 gnd 0.008418f
C3789 vdd.n1325 gnd 0.008418f
C3790 vdd.n1326 gnd 0.008418f
C3791 vdd.n1327 gnd 0.008418f
C3792 vdd.n1328 gnd 0.006775f
C3793 vdd.n1329 gnd 0.008418f
C3794 vdd.n1330 gnd 0.008418f
C3795 vdd.n1331 gnd 0.008418f
C3796 vdd.n1332 gnd 0.008418f
C3797 vdd.n1333 gnd 0.008418f
C3798 vdd.t66 gnd 0.103561f
C3799 vdd.t67 gnd 0.110678f
C3800 vdd.t65 gnd 0.135249f
C3801 vdd.n1334 gnd 0.17337f
C3802 vdd.n1335 gnd 0.14634f
C3803 vdd.n1336 gnd 0.014499f
C3804 vdd.n1337 gnd 0.008418f
C3805 vdd.n1338 gnd 0.008418f
C3806 vdd.n1339 gnd 0.008418f
C3807 vdd.n1340 gnd 0.008418f
C3808 vdd.n1341 gnd 0.008418f
C3809 vdd.n1342 gnd 0.006775f
C3810 vdd.n1343 gnd 0.008418f
C3811 vdd.n1344 gnd 0.008418f
C3812 vdd.n1345 gnd 0.008418f
C3813 vdd.n1346 gnd 0.008418f
C3814 vdd.n1347 gnd 0.008418f
C3815 vdd.n1348 gnd 0.006775f
C3816 vdd.n1349 gnd 0.008418f
C3817 vdd.n1350 gnd 0.008418f
C3818 vdd.n1351 gnd 0.008418f
C3819 vdd.n1352 gnd 0.008418f
C3820 vdd.n1353 gnd 0.008418f
C3821 vdd.n1354 gnd 0.006775f
C3822 vdd.n1355 gnd 0.008418f
C3823 vdd.n1356 gnd 0.008418f
C3824 vdd.n1357 gnd 0.008418f
C3825 vdd.n1358 gnd 0.008418f
C3826 vdd.n1359 gnd 0.008418f
C3827 vdd.n1360 gnd 0.006775f
C3828 vdd.n1361 gnd 0.008418f
C3829 vdd.n1362 gnd 0.008418f
C3830 vdd.n1363 gnd 0.008418f
C3831 vdd.n1364 gnd 0.008418f
C3832 vdd.n1365 gnd 0.008418f
C3833 vdd.n1366 gnd 0.006775f
C3834 vdd.n1367 gnd 0.008418f
C3835 vdd.n1368 gnd 0.008418f
C3836 vdd.n1369 gnd 0.008418f
C3837 vdd.n1370 gnd 0.008418f
C3838 vdd.n1371 gnd 0.006775f
C3839 vdd.n1372 gnd 0.008418f
C3840 vdd.n1373 gnd 0.008418f
C3841 vdd.n1374 gnd 0.008418f
C3842 vdd.n1375 gnd 0.008418f
C3843 vdd.n1376 gnd 0.008418f
C3844 vdd.n1377 gnd 0.006775f
C3845 vdd.n1378 gnd 0.008418f
C3846 vdd.n1379 gnd 0.008418f
C3847 vdd.n1380 gnd 0.008418f
C3848 vdd.n1381 gnd 0.008418f
C3849 vdd.n1382 gnd 0.008418f
C3850 vdd.n1383 gnd 0.006775f
C3851 vdd.n1384 gnd 0.008418f
C3852 vdd.n1385 gnd 0.008418f
C3853 vdd.n1386 gnd 0.008418f
C3854 vdd.n1387 gnd 0.008418f
C3855 vdd.n1388 gnd 0.008418f
C3856 vdd.n1389 gnd 0.006775f
C3857 vdd.n1390 gnd 0.008418f
C3858 vdd.n1391 gnd 0.008418f
C3859 vdd.n1392 gnd 0.008418f
C3860 vdd.n1393 gnd 0.008418f
C3861 vdd.n1394 gnd 0.008418f
C3862 vdd.n1395 gnd 0.006775f
C3863 vdd.n1396 gnd 0.008418f
C3864 vdd.n1397 gnd 0.008418f
C3865 vdd.n1398 gnd 0.008418f
C3866 vdd.n1399 gnd 0.008418f
C3867 vdd.t34 gnd 0.103561f
C3868 vdd.t35 gnd 0.110678f
C3869 vdd.t32 gnd 0.135249f
C3870 vdd.n1400 gnd 0.17337f
C3871 vdd.n1401 gnd 0.14634f
C3872 vdd.n1402 gnd 0.011111f
C3873 vdd.n1403 gnd 0.003218f
C3874 vdd.n1404 gnd 0.020985f
C3875 vdd.n1405 gnd 0.008418f
C3876 vdd.n1406 gnd 0.003557f
C3877 vdd.n1407 gnd 0.006775f
C3878 vdd.n1408 gnd 0.006775f
C3879 vdd.n1409 gnd 0.008418f
C3880 vdd.n1410 gnd 0.008418f
C3881 vdd.n1411 gnd 0.008418f
C3882 vdd.n1412 gnd 0.006775f
C3883 vdd.n1413 gnd 0.006775f
C3884 vdd.n1414 gnd 0.006775f
C3885 vdd.n1415 gnd 0.008418f
C3886 vdd.n1416 gnd 0.008418f
C3887 vdd.n1417 gnd 0.008418f
C3888 vdd.n1418 gnd 0.006775f
C3889 vdd.n1419 gnd 0.006775f
C3890 vdd.n1420 gnd 0.006775f
C3891 vdd.n1421 gnd 0.008418f
C3892 vdd.n1422 gnd 0.008418f
C3893 vdd.n1423 gnd 0.008418f
C3894 vdd.n1424 gnd 0.006775f
C3895 vdd.n1425 gnd 0.006775f
C3896 vdd.n1426 gnd 0.006775f
C3897 vdd.n1427 gnd 0.008418f
C3898 vdd.n1428 gnd 0.008418f
C3899 vdd.n1429 gnd 0.008418f
C3900 vdd.n1430 gnd 0.006775f
C3901 vdd.n1431 gnd 0.006775f
C3902 vdd.n1432 gnd 0.006775f
C3903 vdd.n1433 gnd 0.008418f
C3904 vdd.n1434 gnd 0.008418f
C3905 vdd.n1435 gnd 0.008418f
C3906 vdd.n1436 gnd 0.006708f
C3907 vdd.n1437 gnd 0.008418f
C3908 vdd.t49 gnd 0.103561f
C3909 vdd.t50 gnd 0.110678f
C3910 vdd.t48 gnd 0.135249f
C3911 vdd.n1438 gnd 0.17337f
C3912 vdd.n1439 gnd 0.14634f
C3913 vdd.n1440 gnd 0.014499f
C3914 vdd.n1441 gnd 0.004607f
C3915 vdd.n1442 gnd 0.008418f
C3916 vdd.n1443 gnd 0.008418f
C3917 vdd.n1444 gnd 0.008418f
C3918 vdd.n1445 gnd 0.006775f
C3919 vdd.n1446 gnd 0.006775f
C3920 vdd.n1447 gnd 0.006775f
C3921 vdd.n1448 gnd 0.008418f
C3922 vdd.n1449 gnd 0.008418f
C3923 vdd.n1450 gnd 0.008418f
C3924 vdd.n1451 gnd 0.006775f
C3925 vdd.n1452 gnd 0.006775f
C3926 vdd.n1453 gnd 0.006775f
C3927 vdd.n1454 gnd 0.008418f
C3928 vdd.n1455 gnd 0.008418f
C3929 vdd.n1456 gnd 0.008418f
C3930 vdd.n1457 gnd 0.006775f
C3931 vdd.n1458 gnd 0.006775f
C3932 vdd.n1459 gnd 0.006775f
C3933 vdd.n1460 gnd 0.008418f
C3934 vdd.n1461 gnd 0.008418f
C3935 vdd.n1462 gnd 0.008418f
C3936 vdd.n1463 gnd 0.006775f
C3937 vdd.n1464 gnd 0.006775f
C3938 vdd.n1465 gnd 0.006775f
C3939 vdd.n1466 gnd 0.008418f
C3940 vdd.n1467 gnd 0.008418f
C3941 vdd.n1468 gnd 0.008418f
C3942 vdd.n1469 gnd 0.006775f
C3943 vdd.n1470 gnd 0.006775f
C3944 vdd.n1471 gnd 0.005657f
C3945 vdd.n1472 gnd 0.008418f
C3946 vdd.n1473 gnd 0.008418f
C3947 vdd.n1474 gnd 0.008418f
C3948 vdd.n1475 gnd 0.005657f
C3949 vdd.n1476 gnd 0.006775f
C3950 vdd.n1477 gnd 0.006775f
C3951 vdd.n1478 gnd 0.008418f
C3952 vdd.n1479 gnd 0.008418f
C3953 vdd.n1480 gnd 0.008418f
C3954 vdd.n1481 gnd 0.006775f
C3955 vdd.n1482 gnd 0.006775f
C3956 vdd.n1483 gnd 0.006775f
C3957 vdd.n1484 gnd 0.008418f
C3958 vdd.n1485 gnd 0.008418f
C3959 vdd.n1486 gnd 0.008418f
C3960 vdd.n1487 gnd 0.006775f
C3961 vdd.n1488 gnd 0.006775f
C3962 vdd.n1489 gnd 0.006775f
C3963 vdd.n1490 gnd 0.008418f
C3964 vdd.n1491 gnd 0.008418f
C3965 vdd.n1492 gnd 0.008418f
C3966 vdd.n1493 gnd 0.006775f
C3967 vdd.n1494 gnd 0.006775f
C3968 vdd.n1495 gnd 0.006775f
C3969 vdd.n1496 gnd 0.008418f
C3970 vdd.n1497 gnd 0.008418f
C3971 vdd.n1498 gnd 0.008418f
C3972 vdd.n1499 gnd 0.006775f
C3973 vdd.n1500 gnd 0.008418f
C3974 vdd.n1501 gnd 2.05602f
C3975 vdd.n1503 gnd 0.020985f
C3976 vdd.n1504 gnd 0.005623f
C3977 vdd.n1505 gnd 0.020985f
C3978 vdd.n1506 gnd 0.020514f
C3979 vdd.n1507 gnd 0.008418f
C3980 vdd.n1508 gnd 0.006775f
C3981 vdd.n1509 gnd 0.008418f
C3982 vdd.n1510 gnd 0.451635f
C3983 vdd.n1511 gnd 0.008418f
C3984 vdd.n1512 gnd 0.006775f
C3985 vdd.n1513 gnd 0.008418f
C3986 vdd.n1514 gnd 0.008418f
C3987 vdd.n1515 gnd 0.008418f
C3988 vdd.n1516 gnd 0.006775f
C3989 vdd.n1517 gnd 0.008418f
C3990 vdd.n1518 gnd 0.76993f
C3991 vdd.n1519 gnd 0.860257f
C3992 vdd.n1520 gnd 0.008418f
C3993 vdd.n1521 gnd 0.006775f
C3994 vdd.n1522 gnd 0.008418f
C3995 vdd.n1523 gnd 0.008418f
C3996 vdd.n1524 gnd 0.008418f
C3997 vdd.n1525 gnd 0.006775f
C3998 vdd.n1526 gnd 0.008418f
C3999 vdd.n1527 gnd 0.520456f
C4000 vdd.n1528 gnd 0.008418f
C4001 vdd.n1529 gnd 0.006775f
C4002 vdd.n1530 gnd 0.008418f
C4003 vdd.n1531 gnd 0.008418f
C4004 vdd.n1532 gnd 0.008418f
C4005 vdd.n1533 gnd 0.006775f
C4006 vdd.n1534 gnd 0.008418f
C4007 vdd.n1535 gnd 0.477443f
C4008 vdd.n1536 gnd 0.666699f
C4009 vdd.n1537 gnd 0.008418f
C4010 vdd.n1538 gnd 0.006775f
C4011 vdd.n1539 gnd 0.008418f
C4012 vdd.n1540 gnd 0.008418f
C4013 vdd.n1541 gnd 0.00647f
C4014 vdd.n1542 gnd 0.008418f
C4015 vdd.n1543 gnd 0.006775f
C4016 vdd.n1544 gnd 0.008418f
C4017 vdd.n1545 gnd 0.714014f
C4018 vdd.n1546 gnd 0.008418f
C4019 vdd.n1547 gnd 0.006775f
C4020 vdd.n1548 gnd 0.008418f
C4021 vdd.n1549 gnd 0.008418f
C4022 vdd.n1550 gnd 0.008418f
C4023 vdd.n1551 gnd 0.006775f
C4024 vdd.n1552 gnd 0.008418f
C4025 vdd.t6 gnd 0.430129f
C4026 vdd.n1553 gnd 0.615084f
C4027 vdd.n1554 gnd 0.008418f
C4028 vdd.n1555 gnd 0.006775f
C4029 vdd.n1556 gnd 0.00647f
C4030 vdd.n1557 gnd 0.008418f
C4031 vdd.n1558 gnd 0.008418f
C4032 vdd.n1559 gnd 0.006775f
C4033 vdd.n1560 gnd 0.008418f
C4034 vdd.n1561 gnd 0.46884f
C4035 vdd.n1562 gnd 0.008418f
C4036 vdd.n1563 gnd 0.006775f
C4037 vdd.n1564 gnd 0.008418f
C4038 vdd.n1565 gnd 0.008418f
C4039 vdd.n1566 gnd 0.008418f
C4040 vdd.n1567 gnd 0.006775f
C4041 vdd.n1568 gnd 0.008418f
C4042 vdd.n1569 gnd 0.606481f
C4043 vdd.n1570 gnd 0.537661f
C4044 vdd.n1571 gnd 0.008418f
C4045 vdd.n1572 gnd 0.006775f
C4046 vdd.n1573 gnd 0.008418f
C4047 vdd.n1574 gnd 0.008418f
C4048 vdd.n1575 gnd 0.008418f
C4049 vdd.n1576 gnd 0.006775f
C4050 vdd.n1577 gnd 0.008418f
C4051 vdd.n1578 gnd 0.683905f
C4052 vdd.n1579 gnd 0.008418f
C4053 vdd.n1580 gnd 0.006775f
C4054 vdd.n1581 gnd 0.008418f
C4055 vdd.n1582 gnd 0.008418f
C4056 vdd.n1583 gnd 0.020514f
C4057 vdd.n1584 gnd 0.008418f
C4058 vdd.n1585 gnd 0.008418f
C4059 vdd.n1586 gnd 0.006775f
C4060 vdd.n1587 gnd 0.008418f
C4061 vdd.n1588 gnd 0.537661f
C4062 vdd.n1589 gnd 0.860257f
C4063 vdd.n1590 gnd 0.008418f
C4064 vdd.n1591 gnd 0.006775f
C4065 vdd.n1592 gnd 0.008418f
C4066 vdd.n1593 gnd 0.008418f
C4067 vdd.n1594 gnd 0.007239f
C4068 vdd.n1595 gnd 0.006775f
C4069 vdd.n1597 gnd 0.008418f
C4070 vdd.n1599 gnd 0.006775f
C4071 vdd.n1600 gnd 0.008418f
C4072 vdd.n1601 gnd 0.006775f
C4073 vdd.n1603 gnd 0.008418f
C4074 vdd.n1604 gnd 0.006775f
C4075 vdd.n1605 gnd 0.008418f
C4076 vdd.n1606 gnd 0.008418f
C4077 vdd.n1607 gnd 0.008418f
C4078 vdd.n1608 gnd 0.008418f
C4079 vdd.n1609 gnd 0.008418f
C4080 vdd.n1610 gnd 0.006775f
C4081 vdd.n1612 gnd 0.008418f
C4082 vdd.n1613 gnd 0.008418f
C4083 vdd.n1614 gnd 0.008418f
C4084 vdd.n1615 gnd 0.008418f
C4085 vdd.n1616 gnd 0.008418f
C4086 vdd.n1617 gnd 0.006775f
C4087 vdd.n1619 gnd 0.008418f
C4088 vdd.n1620 gnd 0.008418f
C4089 vdd.n1621 gnd 0.008418f
C4090 vdd.n1622 gnd 0.008418f
C4091 vdd.n1623 gnd 0.005657f
C4092 vdd.t84 gnd 0.103561f
C4093 vdd.t83 gnd 0.110678f
C4094 vdd.t82 gnd 0.135249f
C4095 vdd.n1624 gnd 0.17337f
C4096 vdd.n1625 gnd 0.145662f
C4097 vdd.n1627 gnd 0.008418f
C4098 vdd.n1628 gnd 0.008418f
C4099 vdd.n1629 gnd 0.006775f
C4100 vdd.n1630 gnd 0.008418f
C4101 vdd.n1632 gnd 0.008418f
C4102 vdd.n1633 gnd 0.008418f
C4103 vdd.n1634 gnd 0.008418f
C4104 vdd.n1635 gnd 0.008418f
C4105 vdd.n1636 gnd 0.006775f
C4106 vdd.n1638 gnd 0.008418f
C4107 vdd.n1639 gnd 0.008418f
C4108 vdd.n1640 gnd 0.008418f
C4109 vdd.n1641 gnd 0.008418f
C4110 vdd.n1642 gnd 0.008418f
C4111 vdd.n1643 gnd 0.006775f
C4112 vdd.n1645 gnd 0.008418f
C4113 vdd.n1646 gnd 0.008418f
C4114 vdd.n1647 gnd 0.008418f
C4115 vdd.n1648 gnd 0.008418f
C4116 vdd.n1649 gnd 0.008418f
C4117 vdd.n1650 gnd 0.006775f
C4118 vdd.n1652 gnd 0.008418f
C4119 vdd.n1653 gnd 0.008418f
C4120 vdd.n1654 gnd 0.008418f
C4121 vdd.n1655 gnd 0.008418f
C4122 vdd.n1656 gnd 0.008418f
C4123 vdd.n1657 gnd 0.006775f
C4124 vdd.n1659 gnd 0.008418f
C4125 vdd.n1660 gnd 0.008418f
C4126 vdd.n1661 gnd 0.008418f
C4127 vdd.n1662 gnd 0.008418f
C4128 vdd.n1663 gnd 0.006708f
C4129 vdd.t73 gnd 0.103561f
C4130 vdd.t72 gnd 0.110678f
C4131 vdd.t71 gnd 0.135249f
C4132 vdd.n1664 gnd 0.17337f
C4133 vdd.n1665 gnd 0.145662f
C4134 vdd.n1667 gnd 0.008418f
C4135 vdd.n1668 gnd 0.008418f
C4136 vdd.n1669 gnd 0.006775f
C4137 vdd.n1670 gnd 0.008418f
C4138 vdd.n1672 gnd 0.008418f
C4139 vdd.n1673 gnd 0.008418f
C4140 vdd.n1674 gnd 0.008418f
C4141 vdd.n1675 gnd 0.008418f
C4142 vdd.n1676 gnd 0.006775f
C4143 vdd.n1678 gnd 0.008418f
C4144 vdd.n1679 gnd 0.008418f
C4145 vdd.n1680 gnd 0.008418f
C4146 vdd.n1681 gnd 0.008418f
C4147 vdd.n1682 gnd 0.008418f
C4148 vdd.n1683 gnd 0.006775f
C4149 vdd.n1685 gnd 0.008418f
C4150 vdd.n1686 gnd 0.008418f
C4151 vdd.n1687 gnd 0.008418f
C4152 vdd.n1688 gnd 0.008418f
C4153 vdd.n1689 gnd 0.008418f
C4154 vdd.n1690 gnd 0.008418f
C4155 vdd.n1691 gnd 0.006775f
C4156 vdd.n1693 gnd 0.008418f
C4157 vdd.n1695 gnd 0.008418f
C4158 vdd.n1696 gnd 0.006775f
C4159 vdd.n1697 gnd 0.006775f
C4160 vdd.n1698 gnd 0.008418f
C4161 vdd.n1700 gnd 0.008418f
C4162 vdd.n1701 gnd 0.006775f
C4163 vdd.n1702 gnd 0.006775f
C4164 vdd.n1703 gnd 0.008418f
C4165 vdd.n1705 gnd 0.008418f
C4166 vdd.n1706 gnd 0.008418f
C4167 vdd.n1707 gnd 0.006775f
C4168 vdd.n1708 gnd 0.006775f
C4169 vdd.n1709 gnd 0.006775f
C4170 vdd.n1710 gnd 0.008418f
C4171 vdd.n1712 gnd 0.008418f
C4172 vdd.n1713 gnd 0.008418f
C4173 vdd.n1714 gnd 0.006775f
C4174 vdd.n1715 gnd 0.006775f
C4175 vdd.n1716 gnd 0.006775f
C4176 vdd.n1717 gnd 0.008418f
C4177 vdd.n1719 gnd 0.008418f
C4178 vdd.n1720 gnd 0.008418f
C4179 vdd.n1721 gnd 0.006775f
C4180 vdd.n1722 gnd 0.006775f
C4181 vdd.n1723 gnd 0.006775f
C4182 vdd.n1724 gnd 0.008418f
C4183 vdd.n1726 gnd 0.008418f
C4184 vdd.n1727 gnd 0.008418f
C4185 vdd.n1728 gnd 0.006775f
C4186 vdd.n1729 gnd 0.008418f
C4187 vdd.n1730 gnd 0.008418f
C4188 vdd.n1731 gnd 0.008418f
C4189 vdd.n1732 gnd 0.013822f
C4190 vdd.n1733 gnd 0.004607f
C4191 vdd.n1734 gnd 0.006775f
C4192 vdd.n1735 gnd 0.008418f
C4193 vdd.n1737 gnd 0.008418f
C4194 vdd.n1738 gnd 0.008418f
C4195 vdd.n1739 gnd 0.006775f
C4196 vdd.n1740 gnd 0.006775f
C4197 vdd.n1741 gnd 0.006775f
C4198 vdd.n1742 gnd 0.008418f
C4199 vdd.n1744 gnd 0.008418f
C4200 vdd.n1745 gnd 0.008418f
C4201 vdd.n1746 gnd 0.006775f
C4202 vdd.n1747 gnd 0.006775f
C4203 vdd.n1748 gnd 0.006775f
C4204 vdd.n1749 gnd 0.008418f
C4205 vdd.n1751 gnd 0.008418f
C4206 vdd.n1752 gnd 0.008418f
C4207 vdd.n1753 gnd 0.006775f
C4208 vdd.n1754 gnd 0.006775f
C4209 vdd.n1755 gnd 0.006775f
C4210 vdd.n1756 gnd 0.008418f
C4211 vdd.n1758 gnd 0.008418f
C4212 vdd.n1759 gnd 0.008418f
C4213 vdd.n1760 gnd 0.006775f
C4214 vdd.n1761 gnd 0.006775f
C4215 vdd.n1762 gnd 0.006775f
C4216 vdd.n1763 gnd 0.008418f
C4217 vdd.n1765 gnd 0.008418f
C4218 vdd.n1766 gnd 0.008418f
C4219 vdd.n1767 gnd 0.006775f
C4220 vdd.n1768 gnd 0.008418f
C4221 vdd.n1769 gnd 0.008418f
C4222 vdd.n1770 gnd 0.008418f
C4223 vdd.n1771 gnd 0.013822f
C4224 vdd.n1772 gnd 0.005657f
C4225 vdd.n1773 gnd 0.006775f
C4226 vdd.n1774 gnd 0.008418f
C4227 vdd.n1776 gnd 0.008418f
C4228 vdd.n1777 gnd 0.008418f
C4229 vdd.n1778 gnd 0.006775f
C4230 vdd.n1779 gnd 0.006775f
C4231 vdd.n1780 gnd 0.006775f
C4232 vdd.n1781 gnd 0.008418f
C4233 vdd.n1783 gnd 0.008418f
C4234 vdd.n1784 gnd 0.008418f
C4235 vdd.n1785 gnd 0.006775f
C4236 vdd.n1786 gnd 0.006775f
C4237 vdd.n1787 gnd 0.006775f
C4238 vdd.n1788 gnd 0.008418f
C4239 vdd.n1790 gnd 0.008418f
C4240 vdd.n1791 gnd 0.008418f
C4241 vdd.n1793 gnd 0.008418f
C4242 vdd.n1794 gnd 0.006775f
C4243 vdd.n1795 gnd 0.005387f
C4244 vdd.n1796 gnd 0.76575f
C4245 vdd.n1798 gnd 0.006775f
C4246 vdd.n1799 gnd 0.006775f
C4247 vdd.n1800 gnd 0.008418f
C4248 vdd.n1802 gnd 0.008418f
C4249 vdd.n1803 gnd 0.008418f
C4250 vdd.n1804 gnd 0.006775f
C4251 vdd.n1805 gnd 0.005623f
C4252 vdd.n1806 gnd 0.020985f
C4253 vdd.n1807 gnd 0.020514f
C4254 vdd.n1808 gnd 0.005623f
C4255 vdd.n1809 gnd 0.020514f
C4256 vdd.n1810 gnd 1.18285f
C4257 vdd.n1811 gnd 0.020514f
C4258 vdd.n1812 gnd 0.020985f
C4259 vdd.n1813 gnd 0.003218f
C4260 vdd.t64 gnd 0.103561f
C4261 vdd.t63 gnd 0.110678f
C4262 vdd.t61 gnd 0.135249f
C4263 vdd.n1814 gnd 0.17337f
C4264 vdd.n1815 gnd 0.145662f
C4265 vdd.n1816 gnd 0.010434f
C4266 vdd.n1817 gnd 0.003557f
C4267 vdd.n1818 gnd 0.007239f
C4268 vdd.n1819 gnd 0.76575f
C4269 vdd.n1820 gnd 0.030118f
C4270 vdd.n1821 gnd 0.005724f
C4271 vdd.n1822 gnd 0.005724f
C4272 vdd.n1823 gnd 0.005724f
C4273 vdd.n1824 gnd 0.005724f
C4274 vdd.n1825 gnd 0.005724f
C4275 vdd.n1826 gnd 0.005724f
C4276 vdd.n1827 gnd 0.005724f
C4277 vdd.n1828 gnd 0.005724f
C4278 vdd.n1830 gnd 0.005724f
C4279 vdd.n1832 gnd 0.005724f
C4280 vdd.n1833 gnd 0.005724f
C4281 vdd.n1834 gnd 0.005724f
C4282 vdd.n1835 gnd 0.005724f
C4283 vdd.n1836 gnd 0.005724f
C4284 vdd.n1838 gnd 0.005724f
C4285 vdd.n1840 gnd 0.005724f
C4286 vdd.n1841 gnd 0.005724f
C4287 vdd.n1842 gnd 0.005724f
C4288 vdd.n1843 gnd 0.005724f
C4289 vdd.n1844 gnd 0.005724f
C4290 vdd.n1846 gnd 0.005724f
C4291 vdd.n1848 gnd 0.005724f
C4292 vdd.n1849 gnd 0.005724f
C4293 vdd.n1850 gnd 0.005724f
C4294 vdd.n1851 gnd 0.005724f
C4295 vdd.n1852 gnd 0.005724f
C4296 vdd.n1854 gnd 0.005724f
C4297 vdd.n1856 gnd 0.005724f
C4298 vdd.n1857 gnd 0.005724f
C4299 vdd.n1858 gnd 0.005724f
C4300 vdd.n1859 gnd 0.005724f
C4301 vdd.n1860 gnd 0.005724f
C4302 vdd.n1862 gnd 0.005724f
C4303 vdd.n1864 gnd 0.005724f
C4304 vdd.n1865 gnd 0.005724f
C4305 vdd.n1866 gnd 0.005724f
C4306 vdd.n1867 gnd 0.005724f
C4307 vdd.n1868 gnd 0.005724f
C4308 vdd.n1870 gnd 0.005724f
C4309 vdd.n1872 gnd 0.005724f
C4310 vdd.n1873 gnd 0.005724f
C4311 vdd.n1874 gnd 0.005724f
C4312 vdd.n1875 gnd 0.005724f
C4313 vdd.n1876 gnd 0.005724f
C4314 vdd.n1878 gnd 0.005724f
C4315 vdd.n1880 gnd 0.005724f
C4316 vdd.n1881 gnd 0.005724f
C4317 vdd.n1882 gnd 0.005724f
C4318 vdd.n1883 gnd 0.005724f
C4319 vdd.n1884 gnd 0.005724f
C4320 vdd.n1886 gnd 0.005724f
C4321 vdd.n1888 gnd 0.005724f
C4322 vdd.n1889 gnd 0.005724f
C4323 vdd.n1890 gnd 0.004167f
C4324 vdd.n1891 gnd 0.008181f
C4325 vdd.n1892 gnd 0.004419f
C4326 vdd.n1893 gnd 0.005724f
C4327 vdd.n1895 gnd 0.005724f
C4328 vdd.n1896 gnd 0.013193f
C4329 vdd.n1897 gnd 0.013193f
C4330 vdd.n1898 gnd 0.012397f
C4331 vdd.n1899 gnd 0.005724f
C4332 vdd.n1900 gnd 0.005724f
C4333 vdd.n1901 gnd 0.005724f
C4334 vdd.n1902 gnd 0.005724f
C4335 vdd.n1903 gnd 0.005724f
C4336 vdd.n1904 gnd 0.005724f
C4337 vdd.n1905 gnd 0.005724f
C4338 vdd.n1906 gnd 0.005724f
C4339 vdd.n1907 gnd 0.005724f
C4340 vdd.n1908 gnd 0.005724f
C4341 vdd.n1909 gnd 0.005724f
C4342 vdd.n1910 gnd 0.005724f
C4343 vdd.n1911 gnd 0.005724f
C4344 vdd.n1912 gnd 0.005724f
C4345 vdd.n1913 gnd 0.005724f
C4346 vdd.n1914 gnd 0.005724f
C4347 vdd.n1915 gnd 0.005724f
C4348 vdd.n1916 gnd 0.005724f
C4349 vdd.n1917 gnd 0.005724f
C4350 vdd.n1918 gnd 0.005724f
C4351 vdd.n1919 gnd 0.005724f
C4352 vdd.n1920 gnd 0.005724f
C4353 vdd.n1921 gnd 0.005724f
C4354 vdd.n1922 gnd 0.005724f
C4355 vdd.n1923 gnd 0.005724f
C4356 vdd.n1924 gnd 0.005724f
C4357 vdd.n1925 gnd 0.005724f
C4358 vdd.n1926 gnd 0.005724f
C4359 vdd.n1927 gnd 0.005724f
C4360 vdd.n1928 gnd 0.005724f
C4361 vdd.n1929 gnd 0.005724f
C4362 vdd.n1930 gnd 0.005724f
C4363 vdd.n1931 gnd 0.005724f
C4364 vdd.n1932 gnd 0.005724f
C4365 vdd.n1933 gnd 0.005724f
C4366 vdd.n1934 gnd 0.005724f
C4367 vdd.n1935 gnd 0.005724f
C4368 vdd.n1936 gnd 0.005724f
C4369 vdd.n1937 gnd 0.005724f
C4370 vdd.n1938 gnd 0.005724f
C4371 vdd.n1939 gnd 0.005724f
C4372 vdd.n1940 gnd 0.005724f
C4373 vdd.n1941 gnd 0.005724f
C4374 vdd.n1942 gnd 0.005724f
C4375 vdd.n1943 gnd 0.005724f
C4376 vdd.n1944 gnd 0.005724f
C4377 vdd.n1945 gnd 0.005724f
C4378 vdd.n1946 gnd 0.005724f
C4379 vdd.n1947 gnd 0.005724f
C4380 vdd.n1948 gnd 0.348404f
C4381 vdd.n1949 gnd 0.005724f
C4382 vdd.n1950 gnd 0.005724f
C4383 vdd.n1951 gnd 0.005724f
C4384 vdd.n1952 gnd 0.005724f
C4385 vdd.n1953 gnd 0.005724f
C4386 vdd.n1954 gnd 0.005724f
C4387 vdd.n1955 gnd 0.005724f
C4388 vdd.n1956 gnd 0.005724f
C4389 vdd.n1957 gnd 0.005724f
C4390 vdd.n1958 gnd 0.005724f
C4391 vdd.n1959 gnd 0.005724f
C4392 vdd.n1960 gnd 0.529058f
C4393 vdd.n1961 gnd 0.005724f
C4394 vdd.n1962 gnd 0.005724f
C4395 vdd.n1963 gnd 0.005724f
C4396 vdd.n1964 gnd 0.005724f
C4397 vdd.n1965 gnd 0.005724f
C4398 vdd.n1966 gnd 0.005724f
C4399 vdd.n1967 gnd 0.005724f
C4400 vdd.n1968 gnd 0.005724f
C4401 vdd.n1969 gnd 0.005724f
C4402 vdd.n1970 gnd 0.005724f
C4403 vdd.n1971 gnd 0.005724f
C4404 vdd.n1972 gnd 0.184955f
C4405 vdd.n1973 gnd 0.005724f
C4406 vdd.n1974 gnd 0.005724f
C4407 vdd.n1975 gnd 0.005724f
C4408 vdd.n1976 gnd 0.005724f
C4409 vdd.n1977 gnd 0.005724f
C4410 vdd.n1978 gnd 0.005724f
C4411 vdd.n1979 gnd 0.005724f
C4412 vdd.n1980 gnd 0.005724f
C4413 vdd.n1981 gnd 0.005724f
C4414 vdd.n1982 gnd 0.005724f
C4415 vdd.n1983 gnd 0.005724f
C4416 vdd.n1984 gnd 0.005724f
C4417 vdd.n1985 gnd 0.005724f
C4418 vdd.n1986 gnd 0.005724f
C4419 vdd.n1987 gnd 0.005724f
C4420 vdd.n1988 gnd 0.005724f
C4421 vdd.n1989 gnd 0.005724f
C4422 vdd.n1990 gnd 0.005724f
C4423 vdd.n1991 gnd 0.005724f
C4424 vdd.n1992 gnd 0.005724f
C4425 vdd.n1993 gnd 0.005724f
C4426 vdd.n1994 gnd 0.005724f
C4427 vdd.n1995 gnd 0.005724f
C4428 vdd.n1996 gnd 0.005724f
C4429 vdd.n1997 gnd 0.005724f
C4430 vdd.n1998 gnd 0.005724f
C4431 vdd.n1999 gnd 0.005724f
C4432 vdd.n2000 gnd 0.005724f
C4433 vdd.n2001 gnd 0.005724f
C4434 vdd.n2002 gnd 0.005724f
C4435 vdd.n2003 gnd 0.005724f
C4436 vdd.n2004 gnd 0.005724f
C4437 vdd.n2005 gnd 0.005724f
C4438 vdd.n2006 gnd 0.005724f
C4439 vdd.n2007 gnd 0.005724f
C4440 vdd.n2008 gnd 0.012397f
C4441 vdd.n2009 gnd 0.013193f
C4442 vdd.n2010 gnd 0.013193f
C4443 vdd.n2012 gnd 0.005724f
C4444 vdd.n2014 gnd 0.005724f
C4445 vdd.n2015 gnd 0.004419f
C4446 vdd.n2016 gnd 0.008181f
C4447 vdd.n2017 gnd 0.004167f
C4448 vdd.n2018 gnd 0.005724f
C4449 vdd.n2019 gnd 0.005724f
C4450 vdd.n2021 gnd 0.005724f
C4451 vdd.n2023 gnd 0.005724f
C4452 vdd.n2024 gnd 0.005724f
C4453 vdd.n2025 gnd 0.005724f
C4454 vdd.n2026 gnd 0.005724f
C4455 vdd.n2027 gnd 0.005724f
C4456 vdd.n2029 gnd 0.005724f
C4457 vdd.n2031 gnd 0.005724f
C4458 vdd.n2032 gnd 0.005724f
C4459 vdd.n2033 gnd 0.005724f
C4460 vdd.n2034 gnd 0.005724f
C4461 vdd.n2035 gnd 0.005724f
C4462 vdd.n2037 gnd 0.005724f
C4463 vdd.n2039 gnd 0.005724f
C4464 vdd.n2040 gnd 0.005724f
C4465 vdd.n2041 gnd 0.005724f
C4466 vdd.n2042 gnd 0.005724f
C4467 vdd.n2043 gnd 0.005724f
C4468 vdd.n2045 gnd 0.005724f
C4469 vdd.n2047 gnd 0.005724f
C4470 vdd.n2048 gnd 0.005724f
C4471 vdd.n2049 gnd 0.005724f
C4472 vdd.n2050 gnd 0.005724f
C4473 vdd.n2051 gnd 0.005724f
C4474 vdd.n2053 gnd 0.005724f
C4475 vdd.n2055 gnd 0.005724f
C4476 vdd.n2056 gnd 0.005724f
C4477 vdd.n2057 gnd 0.005724f
C4478 vdd.n2058 gnd 0.005724f
C4479 vdd.n2059 gnd 0.005724f
C4480 vdd.n2061 gnd 0.005724f
C4481 vdd.n2063 gnd 0.005724f
C4482 vdd.n2064 gnd 0.005724f
C4483 vdd.n2065 gnd 0.005724f
C4484 vdd.n2066 gnd 0.005724f
C4485 vdd.n2067 gnd 0.005724f
C4486 vdd.n2069 gnd 0.005724f
C4487 vdd.n2070 gnd 0.005724f
C4488 vdd.n2071 gnd 0.005724f
C4489 vdd.n2072 gnd 0.005724f
C4490 vdd.n2073 gnd 0.005724f
C4491 vdd.n2074 gnd 0.005724f
C4492 vdd.n2076 gnd 0.005724f
C4493 vdd.n2077 gnd 0.005724f
C4494 vdd.n2078 gnd 0.013193f
C4495 vdd.n2079 gnd 0.012397f
C4496 vdd.n2080 gnd 0.012397f
C4497 vdd.n2081 gnd 0.808642f
C4498 vdd.n2082 gnd 0.012397f
C4499 vdd.n2083 gnd 0.012397f
C4500 vdd.n2084 gnd 0.005724f
C4501 vdd.n2085 gnd 0.005724f
C4502 vdd.n2086 gnd 0.005724f
C4503 vdd.n2087 gnd 0.40002f
C4504 vdd.n2088 gnd 0.005724f
C4505 vdd.n2089 gnd 0.005724f
C4506 vdd.n2090 gnd 0.005724f
C4507 vdd.n2091 gnd 0.005724f
C4508 vdd.n2092 gnd 0.005724f
C4509 vdd.n2093 gnd 0.584975f
C4510 vdd.n2094 gnd 0.005724f
C4511 vdd.n2095 gnd 0.005724f
C4512 vdd.n2096 gnd 0.005724f
C4513 vdd.n2097 gnd 0.005724f
C4514 vdd.n2098 gnd 0.005724f
C4515 vdd.n2099 gnd 0.584975f
C4516 vdd.n2100 gnd 0.005724f
C4517 vdd.n2101 gnd 0.005724f
C4518 vdd.n2102 gnd 0.005724f
C4519 vdd.n2103 gnd 0.005724f
C4520 vdd.n2104 gnd 0.005724f
C4521 vdd.n2105 gnd 0.296789f
C4522 vdd.n2106 gnd 0.005724f
C4523 vdd.n2107 gnd 0.005724f
C4524 vdd.n2108 gnd 0.005724f
C4525 vdd.n2109 gnd 0.005724f
C4526 vdd.n2110 gnd 0.005724f
C4527 vdd.n2111 gnd 0.425827f
C4528 vdd.n2112 gnd 0.005724f
C4529 vdd.n2113 gnd 0.005724f
C4530 vdd.n2114 gnd 0.005724f
C4531 vdd.n2115 gnd 0.005724f
C4532 vdd.n2116 gnd 0.005724f
C4533 vdd.n2117 gnd 0.554866f
C4534 vdd.n2118 gnd 0.005724f
C4535 vdd.n2119 gnd 0.005724f
C4536 vdd.n2120 gnd 0.005724f
C4537 vdd.n2121 gnd 0.005724f
C4538 vdd.n2122 gnd 0.005724f
C4539 vdd.n2123 gnd 0.584975f
C4540 vdd.n2124 gnd 0.005724f
C4541 vdd.n2125 gnd 0.005724f
C4542 vdd.n2126 gnd 0.005724f
C4543 vdd.n2127 gnd 0.005724f
C4544 vdd.n2128 gnd 0.005724f
C4545 vdd.n2129 gnd 0.486045f
C4546 vdd.n2130 gnd 0.005724f
C4547 vdd.n2131 gnd 0.005724f
C4548 vdd.n2132 gnd 0.004714f
C4549 vdd.n2133 gnd 0.016582f
C4550 vdd.n2134 gnd 0.003872f
C4551 vdd.n2135 gnd 0.005724f
C4552 vdd.n2136 gnd 0.357007f
C4553 vdd.n2137 gnd 0.005724f
C4554 vdd.n2138 gnd 0.005724f
C4555 vdd.n2139 gnd 0.005724f
C4556 vdd.n2140 gnd 0.005724f
C4557 vdd.n2141 gnd 0.005724f
C4558 vdd.n2142 gnd 0.357007f
C4559 vdd.n2143 gnd 0.005724f
C4560 vdd.n2144 gnd 0.005724f
C4561 vdd.n2145 gnd 0.005724f
C4562 vdd.n2146 gnd 0.005724f
C4563 vdd.n2147 gnd 0.005724f
C4564 vdd.n2148 gnd 0.486045f
C4565 vdd.n2149 gnd 0.005724f
C4566 vdd.n2150 gnd 0.005724f
C4567 vdd.n2151 gnd 0.005724f
C4568 vdd.n2152 gnd 0.005724f
C4569 vdd.n2153 gnd 0.005724f
C4570 vdd.n2154 gnd 0.498949f
C4571 vdd.n2155 gnd 0.005724f
C4572 vdd.n2156 gnd 0.005724f
C4573 vdd.n2157 gnd 0.005724f
C4574 vdd.n2158 gnd 0.005724f
C4575 vdd.n2159 gnd 0.005724f
C4576 vdd.n2160 gnd 0.369911f
C4577 vdd.n2161 gnd 0.005724f
C4578 vdd.n2162 gnd 0.005724f
C4579 vdd.n2163 gnd 0.005724f
C4580 vdd.n2164 gnd 0.005724f
C4581 vdd.n2165 gnd 0.005724f
C4582 vdd.n2166 gnd 0.184955f
C4583 vdd.n2167 gnd 0.005724f
C4584 vdd.n2168 gnd 0.005724f
C4585 vdd.n2169 gnd 0.005724f
C4586 vdd.n2170 gnd 0.005724f
C4587 vdd.n2171 gnd 0.005724f
C4588 vdd.n2172 gnd 0.184955f
C4589 vdd.n2173 gnd 0.005724f
C4590 vdd.n2174 gnd 0.005724f
C4591 vdd.n2175 gnd 0.005724f
C4592 vdd.n2176 gnd 0.005724f
C4593 vdd.n2177 gnd 0.005724f
C4594 vdd.n2178 gnd 0.584975f
C4595 vdd.n2179 gnd 0.005724f
C4596 vdd.n2180 gnd 0.005724f
C4597 vdd.n2181 gnd 0.005724f
C4598 vdd.n2182 gnd 0.005724f
C4599 vdd.n2183 gnd 0.005724f
C4600 vdd.n2184 gnd 0.005724f
C4601 vdd.n2185 gnd 0.005724f
C4602 vdd.n2186 gnd 0.421526f
C4603 vdd.n2187 gnd 0.005724f
C4604 vdd.n2188 gnd 0.005724f
C4605 vdd.n2189 gnd 0.005724f
C4606 vdd.n2190 gnd 0.005724f
C4607 vdd.n2191 gnd 0.005724f
C4608 vdd.n2192 gnd 0.005724f
C4609 vdd.n2193 gnd 0.365609f
C4610 vdd.n2194 gnd 0.005724f
C4611 vdd.n2195 gnd 0.005724f
C4612 vdd.n2196 gnd 0.005724f
C4613 vdd.n2197 gnd 0.013123f
C4614 vdd.n2198 gnd 0.012468f
C4615 vdd.n2199 gnd 0.005724f
C4616 vdd.n2200 gnd 0.005724f
C4617 vdd.n2201 gnd 0.004419f
C4618 vdd.n2202 gnd 0.005724f
C4619 vdd.n2203 gnd 0.005724f
C4620 vdd.n2204 gnd 0.004167f
C4621 vdd.n2205 gnd 0.005724f
C4622 vdd.n2206 gnd 0.005724f
C4623 vdd.n2207 gnd 0.005724f
C4624 vdd.n2208 gnd 0.005724f
C4625 vdd.n2209 gnd 0.005724f
C4626 vdd.n2210 gnd 0.005724f
C4627 vdd.n2211 gnd 0.005724f
C4628 vdd.n2212 gnd 0.005724f
C4629 vdd.n2213 gnd 0.005724f
C4630 vdd.n2214 gnd 0.005724f
C4631 vdd.n2215 gnd 0.005724f
C4632 vdd.n2216 gnd 0.005724f
C4633 vdd.n2217 gnd 0.005724f
C4634 vdd.n2218 gnd 0.005724f
C4635 vdd.n2219 gnd 0.005724f
C4636 vdd.n2220 gnd 0.005724f
C4637 vdd.n2221 gnd 0.005724f
C4638 vdd.n2222 gnd 0.005724f
C4639 vdd.n2223 gnd 0.005724f
C4640 vdd.n2224 gnd 0.005724f
C4641 vdd.n2225 gnd 0.005724f
C4642 vdd.n2226 gnd 0.005724f
C4643 vdd.n2227 gnd 0.005724f
C4644 vdd.n2228 gnd 0.005724f
C4645 vdd.n2229 gnd 0.005724f
C4646 vdd.n2230 gnd 0.005724f
C4647 vdd.n2231 gnd 0.005724f
C4648 vdd.n2232 gnd 0.005724f
C4649 vdd.n2233 gnd 0.005724f
C4650 vdd.n2234 gnd 0.005724f
C4651 vdd.n2235 gnd 0.005724f
C4652 vdd.n2236 gnd 0.005724f
C4653 vdd.n2237 gnd 0.005724f
C4654 vdd.n2238 gnd 0.005724f
C4655 vdd.n2239 gnd 0.005724f
C4656 vdd.n2240 gnd 0.005724f
C4657 vdd.n2241 gnd 0.005724f
C4658 vdd.n2242 gnd 0.005724f
C4659 vdd.n2243 gnd 0.005724f
C4660 vdd.n2244 gnd 0.005724f
C4661 vdd.n2245 gnd 0.005724f
C4662 vdd.n2246 gnd 0.005724f
C4663 vdd.n2247 gnd 0.005724f
C4664 vdd.n2248 gnd 0.005724f
C4665 vdd.n2249 gnd 0.005724f
C4666 vdd.n2250 gnd 0.005724f
C4667 vdd.n2251 gnd 0.005724f
C4668 vdd.n2252 gnd 0.005724f
C4669 vdd.n2253 gnd 0.005724f
C4670 vdd.n2254 gnd 0.005724f
C4671 vdd.n2255 gnd 0.005724f
C4672 vdd.n2256 gnd 0.005724f
C4673 vdd.n2257 gnd 0.005724f
C4674 vdd.n2258 gnd 0.005724f
C4675 vdd.n2259 gnd 0.005724f
C4676 vdd.n2260 gnd 0.005724f
C4677 vdd.n2261 gnd 0.005724f
C4678 vdd.n2262 gnd 0.005724f
C4679 vdd.n2263 gnd 0.005724f
C4680 vdd.n2264 gnd 0.005724f
C4681 vdd.n2265 gnd 0.013193f
C4682 vdd.n2266 gnd 0.012397f
C4683 vdd.n2267 gnd 0.012397f
C4684 vdd.n2268 gnd 0.679603f
C4685 vdd.n2269 gnd 0.012397f
C4686 vdd.n2270 gnd 0.013193f
C4687 vdd.n2271 gnd 0.012468f
C4688 vdd.n2272 gnd 0.005724f
C4689 vdd.n2273 gnd 0.005724f
C4690 vdd.n2274 gnd 0.005724f
C4691 vdd.n2275 gnd 0.004419f
C4692 vdd.n2276 gnd 0.008181f
C4693 vdd.n2277 gnd 0.004167f
C4694 vdd.n2278 gnd 0.005724f
C4695 vdd.n2279 gnd 0.005724f
C4696 vdd.n2280 gnd 0.005724f
C4697 vdd.n2281 gnd 0.005724f
C4698 vdd.n2282 gnd 0.005724f
C4699 vdd.n2283 gnd 0.005724f
C4700 vdd.n2284 gnd 0.005724f
C4701 vdd.n2285 gnd 0.005724f
C4702 vdd.n2286 gnd 0.005724f
C4703 vdd.n2287 gnd 0.005724f
C4704 vdd.n2288 gnd 0.005724f
C4705 vdd.n2289 gnd 0.005724f
C4706 vdd.n2290 gnd 0.005724f
C4707 vdd.n2291 gnd 0.005724f
C4708 vdd.n2292 gnd 0.005724f
C4709 vdd.n2293 gnd 0.005724f
C4710 vdd.n2294 gnd 0.005724f
C4711 vdd.n2295 gnd 0.005724f
C4712 vdd.n2296 gnd 0.005724f
C4713 vdd.n2297 gnd 0.005724f
C4714 vdd.n2298 gnd 0.005724f
C4715 vdd.n2299 gnd 0.005724f
C4716 vdd.n2300 gnd 0.005724f
C4717 vdd.n2301 gnd 0.005724f
C4718 vdd.n2302 gnd 0.005724f
C4719 vdd.n2303 gnd 0.005724f
C4720 vdd.n2304 gnd 0.005724f
C4721 vdd.n2305 gnd 0.005724f
C4722 vdd.n2306 gnd 0.005724f
C4723 vdd.n2307 gnd 0.005724f
C4724 vdd.n2308 gnd 0.005724f
C4725 vdd.n2309 gnd 0.005724f
C4726 vdd.n2310 gnd 0.005724f
C4727 vdd.n2311 gnd 0.005724f
C4728 vdd.n2312 gnd 0.005724f
C4729 vdd.n2313 gnd 0.005724f
C4730 vdd.n2314 gnd 0.005724f
C4731 vdd.n2315 gnd 0.005724f
C4732 vdd.n2316 gnd 0.005724f
C4733 vdd.n2317 gnd 0.005724f
C4734 vdd.n2318 gnd 0.005724f
C4735 vdd.n2319 gnd 0.005724f
C4736 vdd.n2320 gnd 0.005724f
C4737 vdd.n2321 gnd 0.005724f
C4738 vdd.n2322 gnd 0.005724f
C4739 vdd.n2323 gnd 0.005724f
C4740 vdd.n2324 gnd 0.005724f
C4741 vdd.n2325 gnd 0.005724f
C4742 vdd.n2326 gnd 0.005724f
C4743 vdd.n2327 gnd 0.005724f
C4744 vdd.n2328 gnd 0.005724f
C4745 vdd.n2329 gnd 0.005724f
C4746 vdd.n2330 gnd 0.005724f
C4747 vdd.n2331 gnd 0.005724f
C4748 vdd.n2332 gnd 0.005724f
C4749 vdd.n2333 gnd 0.005724f
C4750 vdd.n2334 gnd 0.005724f
C4751 vdd.n2335 gnd 0.005724f
C4752 vdd.n2336 gnd 0.005724f
C4753 vdd.n2337 gnd 0.005724f
C4754 vdd.n2338 gnd 0.013193f
C4755 vdd.n2339 gnd 0.013193f
C4756 vdd.n2340 gnd 0.714014f
C4757 vdd.t172 gnd 2.53776f
C4758 vdd.t162 gnd 2.53776f
C4759 vdd.n2374 gnd 0.005724f
C4760 vdd.t90 gnd 0.23131f
C4761 vdd.t91 gnd 0.236774f
C4762 vdd.t89 gnd 0.151008f
C4763 vdd.n2375 gnd 0.081612f
C4764 vdd.n2376 gnd 0.046293f
C4765 vdd.n2377 gnd 0.008181f
C4766 vdd.n2378 gnd 0.005724f
C4767 vdd.n2379 gnd 0.005724f
C4768 vdd.n2380 gnd 0.005724f
C4769 vdd.n2381 gnd 0.005724f
C4770 vdd.n2382 gnd 0.005724f
C4771 vdd.n2383 gnd 0.005724f
C4772 vdd.n2384 gnd 0.005724f
C4773 vdd.n2385 gnd 0.005724f
C4774 vdd.n2386 gnd 0.005724f
C4775 vdd.n2387 gnd 0.005724f
C4776 vdd.n2388 gnd 0.005724f
C4777 vdd.n2389 gnd 0.005724f
C4778 vdd.n2390 gnd 0.005724f
C4779 vdd.n2391 gnd 0.005724f
C4780 vdd.n2392 gnd 0.005724f
C4781 vdd.n2393 gnd 0.005724f
C4782 vdd.n2394 gnd 0.005724f
C4783 vdd.n2395 gnd 0.005724f
C4784 vdd.n2396 gnd 0.005724f
C4785 vdd.n2397 gnd 0.005724f
C4786 vdd.n2398 gnd 0.005724f
C4787 vdd.n2399 gnd 0.005724f
C4788 vdd.n2400 gnd 0.005724f
C4789 vdd.n2401 gnd 0.005724f
C4790 vdd.n2402 gnd 0.005724f
C4791 vdd.n2403 gnd 0.005724f
C4792 vdd.n2404 gnd 0.005724f
C4793 vdd.n2405 gnd 0.005724f
C4794 vdd.n2406 gnd 0.005724f
C4795 vdd.n2407 gnd 0.005724f
C4796 vdd.n2408 gnd 0.005724f
C4797 vdd.n2409 gnd 0.005724f
C4798 vdd.n2410 gnd 0.005724f
C4799 vdd.n2411 gnd 0.005724f
C4800 vdd.n2412 gnd 0.005724f
C4801 vdd.n2413 gnd 0.005724f
C4802 vdd.n2414 gnd 0.005724f
C4803 vdd.n2415 gnd 0.005724f
C4804 vdd.n2416 gnd 0.005724f
C4805 vdd.n2417 gnd 0.005724f
C4806 vdd.n2418 gnd 0.005724f
C4807 vdd.n2419 gnd 0.005724f
C4808 vdd.n2420 gnd 0.005724f
C4809 vdd.n2421 gnd 0.005724f
C4810 vdd.n2422 gnd 0.005724f
C4811 vdd.n2423 gnd 0.005724f
C4812 vdd.n2424 gnd 0.005724f
C4813 vdd.n2425 gnd 0.005724f
C4814 vdd.n2426 gnd 0.005724f
C4815 vdd.n2427 gnd 0.005724f
C4816 vdd.n2428 gnd 0.005724f
C4817 vdd.n2429 gnd 0.005724f
C4818 vdd.n2430 gnd 0.005724f
C4819 vdd.n2431 gnd 0.005724f
C4820 vdd.n2432 gnd 0.005724f
C4821 vdd.n2433 gnd 0.005724f
C4822 vdd.n2434 gnd 0.005724f
C4823 vdd.n2435 gnd 0.005724f
C4824 vdd.n2436 gnd 0.005724f
C4825 vdd.n2437 gnd 0.005724f
C4826 vdd.n2438 gnd 0.004167f
C4827 vdd.n2439 gnd 0.005724f
C4828 vdd.n2440 gnd 0.005724f
C4829 vdd.n2441 gnd 0.004419f
C4830 vdd.n2442 gnd 0.005724f
C4831 vdd.n2443 gnd 0.005724f
C4832 vdd.t80 gnd 0.23131f
C4833 vdd.t81 gnd 0.236774f
C4834 vdd.t78 gnd 0.151008f
C4835 vdd.n2444 gnd 0.081612f
C4836 vdd.n2445 gnd 0.046293f
C4837 vdd.n2446 gnd 0.005724f
C4838 vdd.n2447 gnd 0.005724f
C4839 vdd.n2448 gnd 0.005724f
C4840 vdd.n2449 gnd 0.005724f
C4841 vdd.n2450 gnd 0.005724f
C4842 vdd.n2451 gnd 0.005724f
C4843 vdd.n2452 gnd 0.005724f
C4844 vdd.n2453 gnd 0.005724f
C4845 vdd.n2454 gnd 0.005724f
C4846 vdd.n2455 gnd 0.005724f
C4847 vdd.n2456 gnd 0.005724f
C4848 vdd.n2457 gnd 0.005724f
C4849 vdd.n2458 gnd 0.005724f
C4850 vdd.n2459 gnd 0.005724f
C4851 vdd.n2460 gnd 0.005724f
C4852 vdd.n2461 gnd 0.005724f
C4853 vdd.n2462 gnd 0.005724f
C4854 vdd.n2463 gnd 0.005724f
C4855 vdd.n2464 gnd 0.005724f
C4856 vdd.n2465 gnd 0.005724f
C4857 vdd.n2466 gnd 0.005724f
C4858 vdd.n2467 gnd 0.005724f
C4859 vdd.n2468 gnd 0.005724f
C4860 vdd.n2469 gnd 0.005724f
C4861 vdd.n2470 gnd 0.005724f
C4862 vdd.n2471 gnd 0.005724f
C4863 vdd.n2472 gnd 0.005724f
C4864 vdd.n2473 gnd 0.005724f
C4865 vdd.n2474 gnd 0.005724f
C4866 vdd.n2475 gnd 0.005724f
C4867 vdd.n2476 gnd 0.005724f
C4868 vdd.n2477 gnd 0.005724f
C4869 vdd.n2478 gnd 0.005724f
C4870 vdd.n2479 gnd 0.005724f
C4871 vdd.n2480 gnd 0.005724f
C4872 vdd.n2481 gnd 0.005724f
C4873 vdd.n2482 gnd 0.005724f
C4874 vdd.n2483 gnd 0.005724f
C4875 vdd.n2484 gnd 0.005724f
C4876 vdd.n2485 gnd 0.005724f
C4877 vdd.n2486 gnd 0.005724f
C4878 vdd.n2487 gnd 0.005724f
C4879 vdd.n2488 gnd 0.005724f
C4880 vdd.n2489 gnd 0.005724f
C4881 vdd.n2490 gnd 0.005724f
C4882 vdd.n2491 gnd 0.005724f
C4883 vdd.n2492 gnd 0.005724f
C4884 vdd.n2493 gnd 0.005724f
C4885 vdd.n2494 gnd 0.005724f
C4886 vdd.n2495 gnd 0.005724f
C4887 vdd.n2496 gnd 0.005724f
C4888 vdd.n2497 gnd 0.005724f
C4889 vdd.n2498 gnd 0.005724f
C4890 vdd.n2499 gnd 0.005724f
C4891 vdd.n2500 gnd 0.005724f
C4892 vdd.n2501 gnd 0.005724f
C4893 vdd.n2502 gnd 0.005724f
C4894 vdd.n2503 gnd 0.004167f
C4895 vdd.n2504 gnd 0.008181f
C4896 vdd.n2505 gnd 0.004419f
C4897 vdd.n2506 gnd 0.005724f
C4898 vdd.n2507 gnd 0.005724f
C4899 vdd.n2508 gnd 0.005724f
C4900 vdd.n2509 gnd 0.013193f
C4901 vdd.n2510 gnd 0.013193f
C4902 vdd.n2511 gnd 0.012397f
C4903 vdd.n2512 gnd 0.005724f
C4904 vdd.n2513 gnd 0.005724f
C4905 vdd.n2514 gnd 0.005724f
C4906 vdd.n2515 gnd 0.005724f
C4907 vdd.n2516 gnd 0.005724f
C4908 vdd.n2517 gnd 0.005724f
C4909 vdd.n2518 gnd 0.005724f
C4910 vdd.n2519 gnd 0.005724f
C4911 vdd.n2520 gnd 0.005724f
C4912 vdd.n2521 gnd 0.005724f
C4913 vdd.n2522 gnd 0.005724f
C4914 vdd.n2523 gnd 0.005724f
C4915 vdd.n2524 gnd 0.005724f
C4916 vdd.n2525 gnd 0.005724f
C4917 vdd.n2526 gnd 0.005724f
C4918 vdd.n2527 gnd 0.005724f
C4919 vdd.n2528 gnd 0.005724f
C4920 vdd.n2529 gnd 0.005724f
C4921 vdd.n2530 gnd 0.005724f
C4922 vdd.n2531 gnd 0.005724f
C4923 vdd.n2532 gnd 0.005724f
C4924 vdd.n2533 gnd 0.005724f
C4925 vdd.n2534 gnd 0.005724f
C4926 vdd.n2535 gnd 0.005724f
C4927 vdd.n2536 gnd 0.005724f
C4928 vdd.n2537 gnd 0.005724f
C4929 vdd.n2538 gnd 0.005724f
C4930 vdd.n2539 gnd 0.005724f
C4931 vdd.n2540 gnd 0.005724f
C4932 vdd.n2541 gnd 0.005724f
C4933 vdd.n2542 gnd 0.005724f
C4934 vdd.n2543 gnd 0.005724f
C4935 vdd.n2544 gnd 0.005724f
C4936 vdd.n2545 gnd 0.005724f
C4937 vdd.n2546 gnd 0.005724f
C4938 vdd.n2547 gnd 0.005724f
C4939 vdd.n2548 gnd 0.005724f
C4940 vdd.n2549 gnd 0.005724f
C4941 vdd.n2550 gnd 0.005724f
C4942 vdd.n2551 gnd 0.005724f
C4943 vdd.n2552 gnd 0.005724f
C4944 vdd.n2553 gnd 0.005724f
C4945 vdd.n2554 gnd 0.005724f
C4946 vdd.n2555 gnd 0.005724f
C4947 vdd.n2556 gnd 0.005724f
C4948 vdd.n2557 gnd 0.005724f
C4949 vdd.n2558 gnd 0.005724f
C4950 vdd.n2559 gnd 0.005724f
C4951 vdd.n2560 gnd 0.005724f
C4952 vdd.n2561 gnd 0.005724f
C4953 vdd.n2562 gnd 0.005724f
C4954 vdd.n2563 gnd 0.005724f
C4955 vdd.n2564 gnd 0.005724f
C4956 vdd.n2565 gnd 0.005724f
C4957 vdd.n2566 gnd 0.005724f
C4958 vdd.n2567 gnd 0.005724f
C4959 vdd.n2568 gnd 0.005724f
C4960 vdd.n2569 gnd 0.005724f
C4961 vdd.n2570 gnd 0.005724f
C4962 vdd.n2571 gnd 0.005724f
C4963 vdd.n2572 gnd 0.005724f
C4964 vdd.n2573 gnd 0.005724f
C4965 vdd.n2574 gnd 0.005724f
C4966 vdd.n2575 gnd 0.005724f
C4967 vdd.n2576 gnd 0.005724f
C4968 vdd.n2577 gnd 0.005724f
C4969 vdd.n2578 gnd 0.005724f
C4970 vdd.n2579 gnd 0.005724f
C4971 vdd.n2580 gnd 0.005724f
C4972 vdd.n2581 gnd 0.005724f
C4973 vdd.n2582 gnd 0.005724f
C4974 vdd.n2583 gnd 0.005724f
C4975 vdd.n2584 gnd 0.005724f
C4976 vdd.n2585 gnd 0.005724f
C4977 vdd.n2586 gnd 0.005724f
C4978 vdd.n2587 gnd 0.005724f
C4979 vdd.n2588 gnd 0.005724f
C4980 vdd.n2589 gnd 0.005724f
C4981 vdd.n2590 gnd 0.005724f
C4982 vdd.n2591 gnd 0.184955f
C4983 vdd.n2592 gnd 0.005724f
C4984 vdd.n2593 gnd 0.005724f
C4985 vdd.n2594 gnd 0.005724f
C4986 vdd.n2595 gnd 0.005724f
C4987 vdd.n2596 gnd 0.005724f
C4988 vdd.n2597 gnd 0.005724f
C4989 vdd.n2598 gnd 0.005724f
C4990 vdd.n2599 gnd 0.005724f
C4991 vdd.n2600 gnd 0.005724f
C4992 vdd.n2601 gnd 0.005724f
C4993 vdd.n2602 gnd 0.005724f
C4994 vdd.n2603 gnd 0.529058f
C4995 vdd.n2604 gnd 0.005724f
C4996 vdd.n2605 gnd 0.005724f
C4997 vdd.n2606 gnd 0.005724f
C4998 vdd.n2607 gnd 0.005724f
C4999 vdd.n2608 gnd 0.005724f
C5000 vdd.n2609 gnd 0.005724f
C5001 vdd.n2610 gnd 0.005724f
C5002 vdd.n2611 gnd 0.005724f
C5003 vdd.n2612 gnd 0.005724f
C5004 vdd.n2613 gnd 0.005724f
C5005 vdd.n2614 gnd 0.005724f
C5006 vdd.n2615 gnd 0.348404f
C5007 vdd.n2616 gnd 0.005724f
C5008 vdd.n2617 gnd 0.005724f
C5009 vdd.n2618 gnd 0.005724f
C5010 vdd.n2619 gnd 0.005724f
C5011 vdd.n2620 gnd 0.005724f
C5012 vdd.n2621 gnd 0.012397f
C5013 vdd.n2622 gnd 0.013193f
C5014 vdd.n2623 gnd 0.013193f
C5015 vdd.n2624 gnd 0.714014f
C5016 vdd.n2626 gnd 0.005724f
C5017 vdd.n2627 gnd 0.005724f
C5018 vdd.n2628 gnd 0.013193f
C5019 vdd.n2629 gnd 0.012397f
C5020 vdd.n2630 gnd 0.012397f
C5021 vdd.n2631 gnd 0.679603f
C5022 vdd.n2632 gnd 0.012397f
C5023 vdd.n2633 gnd 0.012397f
C5024 vdd.n2634 gnd 0.005724f
C5025 vdd.n2635 gnd 0.005724f
C5026 vdd.n2636 gnd 0.005724f
C5027 vdd.n2637 gnd 0.365609f
C5028 vdd.n2638 gnd 0.005724f
C5029 vdd.n2639 gnd 0.005724f
C5030 vdd.n2640 gnd 0.005724f
C5031 vdd.n2641 gnd 0.005724f
C5032 vdd.n2642 gnd 0.005724f
C5033 vdd.n2643 gnd 0.421526f
C5034 vdd.n2644 gnd 0.005724f
C5035 vdd.n2645 gnd 0.005724f
C5036 vdd.n2646 gnd 0.005724f
C5037 vdd.n2647 gnd 0.005724f
C5038 vdd.n2648 gnd 0.005724f
C5039 vdd.n2649 gnd 0.584975f
C5040 vdd.n2650 gnd 0.005724f
C5041 vdd.n2651 gnd 0.005724f
C5042 vdd.n2652 gnd 0.005724f
C5043 vdd.n2653 gnd 0.005724f
C5044 vdd.n2654 gnd 0.005724f
C5045 vdd.n2655 gnd 0.184955f
C5046 vdd.n2656 gnd 0.005724f
C5047 vdd.n2657 gnd 0.005724f
C5048 vdd.n2658 gnd 0.005724f
C5049 vdd.n2659 gnd 0.005724f
C5050 vdd.n2660 gnd 0.005724f
C5051 vdd.n2661 gnd 0.184955f
C5052 vdd.n2662 gnd 0.005724f
C5053 vdd.n2663 gnd 0.005724f
C5054 vdd.n2664 gnd 0.005724f
C5055 vdd.n2665 gnd 0.005724f
C5056 vdd.n2666 gnd 0.005724f
C5057 vdd.n2667 gnd 0.369911f
C5058 vdd.n2668 gnd 0.005724f
C5059 vdd.n2669 gnd 0.005724f
C5060 vdd.n2670 gnd 0.005724f
C5061 vdd.n2671 gnd 0.005724f
C5062 vdd.n2672 gnd 0.005724f
C5063 vdd.n2673 gnd 0.498949f
C5064 vdd.n2674 gnd 0.005724f
C5065 vdd.n2675 gnd 0.005724f
C5066 vdd.n2676 gnd 0.005724f
C5067 vdd.n2677 gnd 0.005724f
C5068 vdd.n2678 gnd 0.005724f
C5069 vdd.n2679 gnd 0.486045f
C5070 vdd.n2680 gnd 0.005724f
C5071 vdd.n2681 gnd 0.005724f
C5072 vdd.n2682 gnd 0.005724f
C5073 vdd.n2683 gnd 0.005724f
C5074 vdd.n2684 gnd 0.005724f
C5075 vdd.n2685 gnd 0.357007f
C5076 vdd.n2686 gnd 0.005724f
C5077 vdd.n2687 gnd 0.005724f
C5078 vdd.n2688 gnd 0.005724f
C5079 vdd.n2689 gnd 0.005724f
C5080 vdd.n2690 gnd 0.005724f
C5081 vdd.n2691 gnd 0.357007f
C5082 vdd.n2692 gnd 0.005724f
C5083 vdd.n2693 gnd 0.003872f
C5084 vdd.n2694 gnd 0.016582f
C5085 vdd.n2695 gnd 0.004714f
C5086 vdd.n2696 gnd 0.005724f
C5087 vdd.n2697 gnd 0.005724f
C5088 vdd.n2698 gnd 0.486045f
C5089 vdd.n2699 gnd 0.005724f
C5090 vdd.n2700 gnd 0.005724f
C5091 vdd.n2701 gnd 0.005724f
C5092 vdd.n2702 gnd 0.005724f
C5093 vdd.n2703 gnd 0.005724f
C5094 vdd.n2704 gnd 0.584975f
C5095 vdd.n2705 gnd 0.005724f
C5096 vdd.n2706 gnd 0.005724f
C5097 vdd.n2707 gnd 0.005724f
C5098 vdd.n2708 gnd 0.005724f
C5099 vdd.n2709 gnd 0.005724f
C5100 vdd.n2710 gnd 0.554866f
C5101 vdd.n2711 gnd 0.005724f
C5102 vdd.n2712 gnd 0.005724f
C5103 vdd.n2713 gnd 0.005724f
C5104 vdd.n2714 gnd 0.005724f
C5105 vdd.n2715 gnd 0.005724f
C5106 vdd.n2716 gnd 0.425827f
C5107 vdd.n2717 gnd 0.005724f
C5108 vdd.n2718 gnd 0.005724f
C5109 vdd.n2719 gnd 0.005724f
C5110 vdd.n2720 gnd 0.005724f
C5111 vdd.n2721 gnd 0.005724f
C5112 vdd.n2722 gnd 0.296789f
C5113 vdd.n2723 gnd 0.005724f
C5114 vdd.n2724 gnd 0.005724f
C5115 vdd.n2725 gnd 0.005724f
C5116 vdd.n2726 gnd 0.005724f
C5117 vdd.n2727 gnd 0.005724f
C5118 vdd.n2728 gnd 0.584975f
C5119 vdd.n2729 gnd 0.005724f
C5120 vdd.n2730 gnd 0.005724f
C5121 vdd.n2731 gnd 0.005724f
C5122 vdd.n2732 gnd 0.005724f
C5123 vdd.n2733 gnd 0.005724f
C5124 vdd.n2734 gnd 0.005724f
C5125 vdd.n2736 gnd 0.005724f
C5126 vdd.n2737 gnd 0.005724f
C5127 vdd.n2739 gnd 0.005724f
C5128 vdd.n2740 gnd 0.005724f
C5129 vdd.n2743 gnd 0.005724f
C5130 vdd.n2744 gnd 0.005724f
C5131 vdd.n2745 gnd 0.005724f
C5132 vdd.n2746 gnd 0.005724f
C5133 vdd.n2748 gnd 0.005724f
C5134 vdd.n2749 gnd 0.005724f
C5135 vdd.n2750 gnd 0.005724f
C5136 vdd.n2751 gnd 0.005724f
C5137 vdd.n2752 gnd 0.005724f
C5138 vdd.n2753 gnd 0.005724f
C5139 vdd.n2755 gnd 0.005724f
C5140 vdd.n2756 gnd 0.005724f
C5141 vdd.n2757 gnd 0.005724f
C5142 vdd.n2758 gnd 0.005724f
C5143 vdd.n2759 gnd 0.005724f
C5144 vdd.n2760 gnd 0.005724f
C5145 vdd.n2762 gnd 0.005724f
C5146 vdd.n2763 gnd 0.005724f
C5147 vdd.n2764 gnd 0.005724f
C5148 vdd.n2765 gnd 0.005724f
C5149 vdd.n2766 gnd 0.005724f
C5150 vdd.n2767 gnd 0.005724f
C5151 vdd.n2769 gnd 0.005724f
C5152 vdd.n2770 gnd 0.013193f
C5153 vdd.n2771 gnd 0.013193f
C5154 vdd.n2772 gnd 0.012397f
C5155 vdd.n2773 gnd 0.005724f
C5156 vdd.n2774 gnd 0.005724f
C5157 vdd.n2775 gnd 0.005724f
C5158 vdd.n2776 gnd 0.005724f
C5159 vdd.n2777 gnd 0.005724f
C5160 vdd.n2778 gnd 0.005724f
C5161 vdd.n2779 gnd 0.584975f
C5162 vdd.n2780 gnd 0.005724f
C5163 vdd.n2781 gnd 0.005724f
C5164 vdd.n2782 gnd 0.005724f
C5165 vdd.n2783 gnd 0.005724f
C5166 vdd.n2784 gnd 0.005724f
C5167 vdd.n2785 gnd 0.40002f
C5168 vdd.n2786 gnd 0.005724f
C5169 vdd.n2787 gnd 0.005724f
C5170 vdd.n2788 gnd 0.005724f
C5171 vdd.n2789 gnd 0.013123f
C5172 vdd.n2790 gnd 0.012468f
C5173 vdd.n2791 gnd 0.013193f
C5174 vdd.n2793 gnd 0.005724f
C5175 vdd.n2794 gnd 0.005724f
C5176 vdd.n2795 gnd 0.004419f
C5177 vdd.n2796 gnd 0.008181f
C5178 vdd.n2797 gnd 0.004167f
C5179 vdd.n2798 gnd 0.005724f
C5180 vdd.n2799 gnd 0.005724f
C5181 vdd.n2801 gnd 0.005724f
C5182 vdd.n2802 gnd 0.005724f
C5183 vdd.n2803 gnd 0.005724f
C5184 vdd.n2804 gnd 0.005724f
C5185 vdd.n2805 gnd 0.005724f
C5186 vdd.n2806 gnd 0.005724f
C5187 vdd.n2808 gnd 0.005724f
C5188 vdd.n2809 gnd 0.005724f
C5189 vdd.n2810 gnd 0.005724f
C5190 vdd.n2811 gnd 0.005724f
C5191 vdd.n2812 gnd 0.005724f
C5192 vdd.n2813 gnd 0.005724f
C5193 vdd.n2815 gnd 0.005724f
C5194 vdd.n2816 gnd 0.005724f
C5195 vdd.n2817 gnd 0.005724f
C5196 vdd.n2818 gnd 0.005724f
C5197 vdd.n2819 gnd 0.005724f
C5198 vdd.n2820 gnd 0.005724f
C5199 vdd.n2822 gnd 0.005724f
C5200 vdd.n2823 gnd 0.005724f
C5201 vdd.n2824 gnd 0.005724f
C5202 vdd.n2826 gnd 0.005724f
C5203 vdd.n2827 gnd 0.005724f
C5204 vdd.n2828 gnd 0.005724f
C5205 vdd.n2829 gnd 0.005724f
C5206 vdd.n2830 gnd 0.005724f
C5207 vdd.n2831 gnd 0.005724f
C5208 vdd.n2833 gnd 0.005724f
C5209 vdd.n2834 gnd 0.005724f
C5210 vdd.n2835 gnd 0.005724f
C5211 vdd.n2836 gnd 0.005724f
C5212 vdd.n2837 gnd 0.005724f
C5213 vdd.n2838 gnd 0.005724f
C5214 vdd.n2840 gnd 0.005724f
C5215 vdd.n2841 gnd 0.005724f
C5216 vdd.n2842 gnd 0.005724f
C5217 vdd.n2843 gnd 0.005724f
C5218 vdd.n2844 gnd 0.005724f
C5219 vdd.n2845 gnd 0.005724f
C5220 vdd.n2847 gnd 0.005724f
C5221 vdd.n2848 gnd 0.005724f
C5222 vdd.n2850 gnd 0.005724f
C5223 vdd.n2851 gnd 0.005724f
C5224 vdd.n2852 gnd 0.013193f
C5225 vdd.n2853 gnd 0.012397f
C5226 vdd.n2854 gnd 0.012397f
C5227 vdd.n2855 gnd 0.808642f
C5228 vdd.n2856 gnd 0.012397f
C5229 vdd.n2857 gnd 0.013193f
C5230 vdd.n2858 gnd 0.012468f
C5231 vdd.n2859 gnd 0.005724f
C5232 vdd.n2860 gnd 0.004419f
C5233 vdd.n2861 gnd 0.005724f
C5234 vdd.n2863 gnd 0.005724f
C5235 vdd.n2864 gnd 0.005724f
C5236 vdd.n2865 gnd 0.005724f
C5237 vdd.n2866 gnd 0.005724f
C5238 vdd.n2867 gnd 0.005724f
C5239 vdd.n2868 gnd 0.005724f
C5240 vdd.n2870 gnd 0.005724f
C5241 vdd.n2871 gnd 0.005724f
C5242 vdd.n2872 gnd 0.005724f
C5243 vdd.n2873 gnd 0.005724f
C5244 vdd.n2874 gnd 0.005724f
C5245 vdd.n2875 gnd 0.005724f
C5246 vdd.n2877 gnd 0.005724f
C5247 vdd.n2878 gnd 0.005724f
C5248 vdd.n2879 gnd 0.005724f
C5249 vdd.n2880 gnd 0.005724f
C5250 vdd.n2881 gnd 0.005724f
C5251 vdd.n2882 gnd 0.005724f
C5252 vdd.n2884 gnd 0.005724f
C5253 vdd.n2885 gnd 0.005724f
C5254 vdd.n2887 gnd 0.005724f
C5255 vdd.n2888 gnd 0.026869f
C5256 vdd.n2889 gnd 0.768998f
C5257 vdd.n2890 gnd 0.007239f
C5258 vdd.n2891 gnd 0.020985f
C5259 vdd.n2892 gnd 0.003218f
C5260 vdd.t59 gnd 0.103561f
C5261 vdd.t60 gnd 0.110678f
C5262 vdd.t58 gnd 0.135249f
C5263 vdd.n2893 gnd 0.17337f
C5264 vdd.n2894 gnd 0.145662f
C5265 vdd.n2895 gnd 0.010434f
C5266 vdd.n2896 gnd 0.008418f
C5267 vdd.n2897 gnd 0.003557f
C5268 vdd.n2898 gnd 0.006775f
C5269 vdd.n2899 gnd 0.008418f
C5270 vdd.n2900 gnd 0.008418f
C5271 vdd.n2901 gnd 0.006775f
C5272 vdd.n2902 gnd 0.006775f
C5273 vdd.n2903 gnd 0.008418f
C5274 vdd.n2904 gnd 0.008418f
C5275 vdd.n2905 gnd 0.006775f
C5276 vdd.n2906 gnd 0.006775f
C5277 vdd.n2907 gnd 0.008418f
C5278 vdd.n2908 gnd 0.008418f
C5279 vdd.n2909 gnd 0.006775f
C5280 vdd.n2910 gnd 0.006775f
C5281 vdd.n2911 gnd 0.008418f
C5282 vdd.n2912 gnd 0.008418f
C5283 vdd.n2913 gnd 0.006775f
C5284 vdd.n2914 gnd 0.006775f
C5285 vdd.n2915 gnd 0.008418f
C5286 vdd.n2916 gnd 0.008418f
C5287 vdd.n2917 gnd 0.006775f
C5288 vdd.n2918 gnd 0.006775f
C5289 vdd.n2919 gnd 0.008418f
C5290 vdd.n2920 gnd 0.008418f
C5291 vdd.n2921 gnd 0.006775f
C5292 vdd.n2922 gnd 0.006775f
C5293 vdd.n2923 gnd 0.008418f
C5294 vdd.n2924 gnd 0.008418f
C5295 vdd.n2925 gnd 0.006775f
C5296 vdd.n2926 gnd 0.006775f
C5297 vdd.n2927 gnd 0.008418f
C5298 vdd.n2928 gnd 0.008418f
C5299 vdd.n2929 gnd 0.006775f
C5300 vdd.n2930 gnd 0.006775f
C5301 vdd.n2931 gnd 0.008418f
C5302 vdd.n2932 gnd 0.008418f
C5303 vdd.n2933 gnd 0.006775f
C5304 vdd.n2934 gnd 0.008418f
C5305 vdd.n2935 gnd 0.008418f
C5306 vdd.n2936 gnd 0.006775f
C5307 vdd.n2937 gnd 0.008418f
C5308 vdd.n2938 gnd 0.008418f
C5309 vdd.n2939 gnd 0.008418f
C5310 vdd.n2940 gnd 0.013822f
C5311 vdd.n2941 gnd 0.008418f
C5312 vdd.n2942 gnd 0.008418f
C5313 vdd.n2943 gnd 0.004607f
C5314 vdd.n2944 gnd 0.006775f
C5315 vdd.n2945 gnd 0.008418f
C5316 vdd.n2946 gnd 0.008418f
C5317 vdd.n2947 gnd 0.006775f
C5318 vdd.n2948 gnd 0.006775f
C5319 vdd.n2949 gnd 0.008418f
C5320 vdd.n2950 gnd 0.008418f
C5321 vdd.n2951 gnd 0.006775f
C5322 vdd.n2952 gnd 0.006775f
C5323 vdd.n2953 gnd 0.008418f
C5324 vdd.n2954 gnd 0.008418f
C5325 vdd.n2955 gnd 0.006775f
C5326 vdd.n2956 gnd 0.006775f
C5327 vdd.n2957 gnd 0.008418f
C5328 vdd.n2958 gnd 0.008418f
C5329 vdd.n2959 gnd 0.006775f
C5330 vdd.n2960 gnd 0.006775f
C5331 vdd.n2961 gnd 0.008418f
C5332 vdd.n2962 gnd 0.008418f
C5333 vdd.n2963 gnd 0.006775f
C5334 vdd.n2964 gnd 0.006775f
C5335 vdd.n2965 gnd 0.008418f
C5336 vdd.n2966 gnd 0.008418f
C5337 vdd.n2967 gnd 0.006775f
C5338 vdd.n2968 gnd 0.006775f
C5339 vdd.n2969 gnd 0.008418f
C5340 vdd.n2970 gnd 0.008418f
C5341 vdd.n2971 gnd 0.006775f
C5342 vdd.n2972 gnd 0.006775f
C5343 vdd.n2973 gnd 0.008418f
C5344 vdd.n2974 gnd 0.008418f
C5345 vdd.n2975 gnd 0.006775f
C5346 vdd.n2976 gnd 0.006775f
C5347 vdd.n2977 gnd 0.008418f
C5348 vdd.n2978 gnd 0.008418f
C5349 vdd.n2979 gnd 0.006775f
C5350 vdd.n2980 gnd 0.008418f
C5351 vdd.n2981 gnd 0.008418f
C5352 vdd.n2982 gnd 0.006775f
C5353 vdd.n2983 gnd 0.008418f
C5354 vdd.n2984 gnd 0.008418f
C5355 vdd.n2985 gnd 0.008418f
C5356 vdd.t52 gnd 0.103561f
C5357 vdd.t53 gnd 0.110678f
C5358 vdd.t51 gnd 0.135249f
C5359 vdd.n2986 gnd 0.17337f
C5360 vdd.n2987 gnd 0.145662f
C5361 vdd.n2988 gnd 0.013822f
C5362 vdd.n2989 gnd 0.008418f
C5363 vdd.n2990 gnd 0.008418f
C5364 vdd.n2991 gnd 0.005657f
C5365 vdd.n2992 gnd 0.006775f
C5366 vdd.n2993 gnd 0.008418f
C5367 vdd.n2994 gnd 0.008418f
C5368 vdd.n2995 gnd 0.006775f
C5369 vdd.n2996 gnd 0.006775f
C5370 vdd.n2997 gnd 0.008418f
C5371 vdd.n2998 gnd 0.008418f
C5372 vdd.n2999 gnd 0.006775f
C5373 vdd.n3000 gnd 0.006775f
C5374 vdd.n3001 gnd 0.008418f
C5375 vdd.n3002 gnd 0.008418f
C5376 vdd.n3003 gnd 0.006775f
C5377 vdd.n3004 gnd 0.006775f
C5378 vdd.n3005 gnd 0.008418f
C5379 vdd.n3006 gnd 0.008418f
C5380 vdd.n3007 gnd 0.006775f
C5381 vdd.n3008 gnd 0.006775f
C5382 vdd.n3009 gnd 0.008418f
C5383 vdd.n3010 gnd 0.008418f
C5384 vdd.n3011 gnd 0.006775f
C5385 vdd.n3012 gnd 0.006775f
C5386 vdd.n3013 gnd 0.008418f
C5387 vdd.n3014 gnd 0.008418f
C5388 vdd.n3015 gnd 0.006775f
C5389 vdd.n3016 gnd 0.006775f
C5390 vdd.n3018 gnd 0.768998f
C5391 vdd.n3020 gnd 0.006775f
C5392 vdd.n3021 gnd 0.008418f
C5393 vdd.n3022 gnd 9.09292f
C5394 vdd.n3024 gnd 0.020985f
C5395 vdd.n3025 gnd 0.005623f
C5396 vdd.n3026 gnd 0.020985f
C5397 vdd.n3027 gnd 0.020514f
C5398 vdd.n3028 gnd 0.008418f
C5399 vdd.n3029 gnd 0.006775f
C5400 vdd.n3030 gnd 0.008418f
C5401 vdd.n3031 gnd 0.537661f
C5402 vdd.n3032 gnd 0.008418f
C5403 vdd.n3033 gnd 0.006775f
C5404 vdd.n3034 gnd 0.008418f
C5405 vdd.n3035 gnd 0.008418f
C5406 vdd.n3036 gnd 0.008418f
C5407 vdd.n3037 gnd 0.006775f
C5408 vdd.n3038 gnd 0.008418f
C5409 vdd.n3039 gnd 0.683905f
C5410 vdd.n3040 gnd 0.860257f
C5411 vdd.n3041 gnd 0.008418f
C5412 vdd.n3042 gnd 0.006775f
C5413 vdd.n3043 gnd 0.008418f
C5414 vdd.n3044 gnd 0.008418f
C5415 vdd.n3045 gnd 0.008418f
C5416 vdd.n3046 gnd 0.006775f
C5417 vdd.n3047 gnd 0.008418f
C5418 vdd.n3048 gnd 0.606481f
C5419 vdd.n3049 gnd 0.008418f
C5420 vdd.n3050 gnd 0.006775f
C5421 vdd.n3051 gnd 0.008418f
C5422 vdd.n3052 gnd 0.008418f
C5423 vdd.n3053 gnd 0.008418f
C5424 vdd.n3054 gnd 0.006775f
C5425 vdd.n3055 gnd 0.008418f
C5426 vdd.t24 gnd 0.430129f
C5427 vdd.n3056 gnd 0.714014f
C5428 vdd.n3057 gnd 0.008418f
C5429 vdd.n3058 gnd 0.006775f
C5430 vdd.n3059 gnd 0.008418f
C5431 vdd.n3060 gnd 0.008418f
C5432 vdd.n3061 gnd 0.008418f
C5433 vdd.n3062 gnd 0.006775f
C5434 vdd.n3063 gnd 0.008418f
C5435 vdd.n3064 gnd 0.675302f
C5436 vdd.n3065 gnd 0.008418f
C5437 vdd.n3066 gnd 0.006775f
C5438 vdd.n3067 gnd 0.008418f
C5439 vdd.n3068 gnd 0.008418f
C5440 vdd.n3069 gnd 0.008418f
C5441 vdd.n3070 gnd 0.006775f
C5442 vdd.n3071 gnd 0.006775f
C5443 vdd.n3072 gnd 0.006775f
C5444 vdd.n3073 gnd 0.008418f
C5445 vdd.n3074 gnd 0.008418f
C5446 vdd.n3075 gnd 0.008418f
C5447 vdd.n3076 gnd 0.006775f
C5448 vdd.n3077 gnd 0.006775f
C5449 vdd.n3078 gnd 0.006775f
C5450 vdd.n3079 gnd 0.008418f
C5451 vdd.n3080 gnd 0.008418f
C5452 vdd.n3081 gnd 0.008418f
C5453 vdd.n3082 gnd 0.006775f
C5454 vdd.n3083 gnd 0.006775f
C5455 vdd.n3084 gnd 0.005623f
C5456 vdd.n3085 gnd 0.020514f
C5457 vdd.n3086 gnd 0.020985f
C5458 vdd.n3088 gnd 0.020985f
C5459 vdd.n3089 gnd 0.003218f
C5460 vdd.t31 gnd 0.103561f
C5461 vdd.t30 gnd 0.110678f
C5462 vdd.t28 gnd 0.135249f
C5463 vdd.n3090 gnd 0.17337f
C5464 vdd.n3091 gnd 0.14634f
C5465 vdd.n3092 gnd 0.011111f
C5466 vdd.n3093 gnd 0.003557f
C5467 vdd.n3094 gnd 0.006775f
C5468 vdd.n3095 gnd 0.008418f
C5469 vdd.n3097 gnd 0.008418f
C5470 vdd.n3098 gnd 0.008418f
C5471 vdd.n3099 gnd 0.006775f
C5472 vdd.n3100 gnd 0.006775f
C5473 vdd.n3101 gnd 0.006775f
C5474 vdd.n3102 gnd 0.008418f
C5475 vdd.n3104 gnd 0.008418f
C5476 vdd.n3105 gnd 0.008418f
C5477 vdd.n3106 gnd 0.006775f
C5478 vdd.n3107 gnd 0.006775f
C5479 vdd.n3108 gnd 0.006775f
C5480 vdd.n3109 gnd 0.008418f
C5481 vdd.n3111 gnd 0.008418f
C5482 vdd.n3112 gnd 0.008418f
C5483 vdd.n3113 gnd 0.006775f
C5484 vdd.n3114 gnd 0.006775f
C5485 vdd.n3115 gnd 0.006775f
C5486 vdd.n3116 gnd 0.008418f
C5487 vdd.n3118 gnd 0.008418f
C5488 vdd.n3119 gnd 0.008418f
C5489 vdd.n3120 gnd 0.006775f
C5490 vdd.n3121 gnd 0.006775f
C5491 vdd.n3122 gnd 0.006775f
C5492 vdd.n3123 gnd 0.008418f
C5493 vdd.n3125 gnd 0.008418f
C5494 vdd.n3126 gnd 0.008418f
C5495 vdd.n3127 gnd 0.006775f
C5496 vdd.n3128 gnd 0.008418f
C5497 vdd.n3129 gnd 0.008418f
C5498 vdd.n3130 gnd 0.008418f
C5499 vdd.n3131 gnd 0.014499f
C5500 vdd.n3132 gnd 0.004607f
C5501 vdd.n3133 gnd 0.006775f
C5502 vdd.n3134 gnd 0.008418f
C5503 vdd.n3136 gnd 0.008418f
C5504 vdd.n3137 gnd 0.008418f
C5505 vdd.n3138 gnd 0.006775f
C5506 vdd.n3139 gnd 0.006775f
C5507 vdd.n3140 gnd 0.006775f
C5508 vdd.n3141 gnd 0.008418f
C5509 vdd.n3143 gnd 0.008418f
C5510 vdd.n3144 gnd 0.008418f
C5511 vdd.n3145 gnd 0.006775f
C5512 vdd.n3146 gnd 0.006775f
C5513 vdd.n3147 gnd 0.006775f
C5514 vdd.n3148 gnd 0.008418f
C5515 vdd.n3150 gnd 0.008418f
C5516 vdd.n3151 gnd 0.008418f
C5517 vdd.n3152 gnd 0.006775f
C5518 vdd.n3153 gnd 0.006775f
C5519 vdd.n3154 gnd 0.006775f
C5520 vdd.n3155 gnd 0.008418f
C5521 vdd.n3157 gnd 0.008418f
C5522 vdd.n3158 gnd 0.008418f
C5523 vdd.n3159 gnd 0.006775f
C5524 vdd.n3160 gnd 0.006775f
C5525 vdd.n3161 gnd 0.006775f
C5526 vdd.n3162 gnd 0.008418f
C5527 vdd.n3164 gnd 0.008418f
C5528 vdd.n3165 gnd 0.008418f
C5529 vdd.n3166 gnd 0.006775f
C5530 vdd.n3167 gnd 0.008418f
C5531 vdd.n3168 gnd 0.008418f
C5532 vdd.n3169 gnd 0.008418f
C5533 vdd.n3170 gnd 0.014499f
C5534 vdd.n3171 gnd 0.005657f
C5535 vdd.n3172 gnd 0.006775f
C5536 vdd.n3173 gnd 0.008418f
C5537 vdd.n3175 gnd 0.008418f
C5538 vdd.n3176 gnd 0.008418f
C5539 vdd.n3177 gnd 0.006775f
C5540 vdd.n3178 gnd 0.006775f
C5541 vdd.n3179 gnd 0.006775f
C5542 vdd.n3180 gnd 0.008418f
C5543 vdd.n3182 gnd 0.008418f
C5544 vdd.n3183 gnd 0.008418f
C5545 vdd.n3184 gnd 0.006775f
C5546 vdd.n3185 gnd 0.006775f
C5547 vdd.n3186 gnd 0.006775f
C5548 vdd.n3187 gnd 0.008418f
C5549 vdd.n3189 gnd 0.008418f
C5550 vdd.n3190 gnd 0.008418f
C5551 vdd.n3191 gnd 0.006775f
C5552 vdd.n3192 gnd 0.006775f
C5553 vdd.n3193 gnd 0.006775f
C5554 vdd.n3194 gnd 0.008418f
C5555 vdd.n3196 gnd 0.008418f
C5556 vdd.n3197 gnd 0.008418f
C5557 vdd.n3199 gnd 0.008418f
C5558 vdd.n3200 gnd 0.006775f
C5559 vdd.n3201 gnd 0.006775f
C5560 vdd.n3202 gnd 0.005623f
C5561 vdd.n3203 gnd 0.020985f
C5562 vdd.n3204 gnd 0.020514f
C5563 vdd.n3205 gnd 0.005623f
C5564 vdd.n3206 gnd 0.020514f
C5565 vdd.n3207 gnd 1.26888f
C5566 vdd.t29 gnd 0.430129f
C5567 vdd.n3208 gnd 0.451635f
C5568 vdd.n3209 gnd 0.860257f
C5569 vdd.n3210 gnd 0.008418f
C5570 vdd.n3211 gnd 0.006775f
C5571 vdd.n3212 gnd 0.006775f
C5572 vdd.n3213 gnd 0.006775f
C5573 vdd.n3214 gnd 0.008418f
C5574 vdd.n3215 gnd 0.76993f
C5575 vdd.t8 gnd 0.430129f
C5576 vdd.n3216 gnd 0.520456f
C5577 vdd.n3217 gnd 0.623687f
C5578 vdd.n3218 gnd 0.008418f
C5579 vdd.n3219 gnd 0.006775f
C5580 vdd.n3220 gnd 0.006775f
C5581 vdd.n3221 gnd 0.006775f
C5582 vdd.n3222 gnd 0.008418f
C5583 vdd.n3223 gnd 0.477443f
C5584 vdd.t10 gnd 0.430129f
C5585 vdd.n3224 gnd 0.714014f
C5586 vdd.t117 gnd 0.430129f
C5587 vdd.n3225 gnd 0.529058f
C5588 vdd.n3226 gnd 0.008418f
C5589 vdd.n3227 gnd 0.006775f
C5590 vdd.n3228 gnd 0.00647f
C5591 vdd.n3229 gnd 0.496513f
C5592 vdd.n3230 gnd 1.90852f
C5593 a_n2472_13878.t18 gnd 0.187389f
C5594 a_n2472_13878.t20 gnd 0.187389f
C5595 a_n2472_13878.t12 gnd 0.187389f
C5596 a_n2472_13878.n0 gnd 1.47709f
C5597 a_n2472_13878.t17 gnd 0.187389f
C5598 a_n2472_13878.t11 gnd 0.187389f
C5599 a_n2472_13878.n1 gnd 1.47552f
C5600 a_n2472_13878.n2 gnd 2.06176f
C5601 a_n2472_13878.t7 gnd 0.187389f
C5602 a_n2472_13878.t9 gnd 0.187389f
C5603 a_n2472_13878.n3 gnd 1.47552f
C5604 a_n2472_13878.n4 gnd 1.00568f
C5605 a_n2472_13878.t19 gnd 0.187389f
C5606 a_n2472_13878.t8 gnd 0.187389f
C5607 a_n2472_13878.n5 gnd 1.47552f
C5608 a_n2472_13878.n6 gnd 1.00568f
C5609 a_n2472_13878.t16 gnd 0.187389f
C5610 a_n2472_13878.t6 gnd 0.187389f
C5611 a_n2472_13878.n7 gnd 1.47552f
C5612 a_n2472_13878.n8 gnd 4.40118f
C5613 a_n2472_13878.t1 gnd 1.75461f
C5614 a_n2472_13878.t25 gnd 0.187389f
C5615 a_n2472_13878.t26 gnd 0.187389f
C5616 a_n2472_13878.n9 gnd 1.31997f
C5617 a_n2472_13878.n10 gnd 1.47487f
C5618 a_n2472_13878.t27 gnd 1.75112f
C5619 a_n2472_13878.n11 gnd 0.742173f
C5620 a_n2472_13878.t2 gnd 1.75112f
C5621 a_n2472_13878.n12 gnd 0.742173f
C5622 a_n2472_13878.t0 gnd 0.187389f
C5623 a_n2472_13878.t3 gnd 0.187389f
C5624 a_n2472_13878.n13 gnd 1.31997f
C5625 a_n2472_13878.n14 gnd 0.749361f
C5626 a_n2472_13878.t4 gnd 1.75112f
C5627 a_n2472_13878.n15 gnd 2.43496f
C5628 a_n2472_13878.n16 gnd 3.22551f
C5629 a_n2472_13878.t21 gnd 0.187389f
C5630 a_n2472_13878.t10 gnd 0.187389f
C5631 a_n2472_13878.n17 gnd 1.47552f
C5632 a_n2472_13878.n18 gnd 2.21835f
C5633 a_n2472_13878.t13 gnd 0.187389f
C5634 a_n2472_13878.t14 gnd 0.187389f
C5635 a_n2472_13878.n19 gnd 1.47552f
C5636 a_n2472_13878.n20 gnd 0.653766f
C5637 a_n2472_13878.t22 gnd 0.187389f
C5638 a_n2472_13878.t23 gnd 0.187389f
C5639 a_n2472_13878.n21 gnd 1.47552f
C5640 a_n2472_13878.n22 gnd 0.653766f
C5641 a_n2472_13878.t5 gnd 0.187389f
C5642 a_n2472_13878.t15 gnd 0.187389f
C5643 a_n2472_13878.n23 gnd 1.47552f
C5644 a_n2472_13878.n24 gnd 1.32631f
C5645 a_n2472_13878.n25 gnd 1.47797f
C5646 a_n2472_13878.t24 gnd 0.187389f
C5647 a_n2848_n452.n0 gnd 4.32595f
C5648 a_n2848_n452.n1 gnd 3.093f
C5649 a_n2848_n452.n2 gnd 3.95526f
C5650 a_n2848_n452.n3 gnd 0.896217f
C5651 a_n2848_n452.n4 gnd 0.896219f
C5652 a_n2848_n452.n5 gnd 0.212016f
C5653 a_n2848_n452.n6 gnd 0.918052f
C5654 a_n2848_n452.n7 gnd 0.212016f
C5655 a_n2848_n452.n8 gnd 0.493974f
C5656 a_n2848_n452.n9 gnd 0.44097f
C5657 a_n2848_n452.n10 gnd 2.93735f
C5658 a_n2848_n452.n11 gnd 0.212016f
C5659 a_n2848_n452.n12 gnd 0.788457f
C5660 a_n2848_n452.n13 gnd 0.788376f
C5661 a_n2848_n452.n14 gnd 0.201168f
C5662 a_n2848_n452.n15 gnd 0.148164f
C5663 a_n2848_n452.n16 gnd 0.232867f
C5664 a_n2848_n452.n17 gnd 0.179863f
C5665 a_n2848_n452.n18 gnd 0.201168f
C5666 a_n2848_n452.n19 gnd 0.148164f
C5667 a_n2848_n452.n20 gnd 0.84138f
C5668 a_n2848_n452.n21 gnd 0.212016f
C5669 a_n2848_n452.n22 gnd 0.684161f
C5670 a_n2848_n452.n23 gnd 0.212016f
C5671 a_n2848_n452.n24 gnd 0.493974f
C5672 a_n2848_n452.n25 gnd 0.212016f
C5673 a_n2848_n452.n26 gnd 0.546979f
C5674 a_n2848_n452.n27 gnd 0.212016f
C5675 a_n2848_n452.n28 gnd 0.87769f
C5676 a_n2848_n452.n29 gnd 1.7455f
C5677 a_n2848_n452.n30 gnd 1.17615f
C5678 a_n2848_n452.n31 gnd 1.15743f
C5679 a_n2848_n452.n32 gnd 1.17615f
C5680 a_n2848_n452.n33 gnd 2.19723f
C5681 a_n2848_n452.n34 gnd 0.008507f
C5682 a_n2848_n452.n35 gnd 4.1e-19
C5683 a_n2848_n452.n37 gnd 0.008209f
C5684 a_n2848_n452.n38 gnd 0.011936f
C5685 a_n2848_n452.n39 gnd 0.007897f
C5686 a_n2848_n452.n40 gnd 0.280073f
C5687 a_n2848_n452.n41 gnd 0.008507f
C5688 a_n2848_n452.n42 gnd 4.1e-19
C5689 a_n2848_n452.n44 gnd 0.008209f
C5690 a_n2848_n452.n45 gnd 0.011936f
C5691 a_n2848_n452.n46 gnd 0.007897f
C5692 a_n2848_n452.n47 gnd 0.280073f
C5693 a_n2848_n452.n48 gnd 0.008209f
C5694 a_n2848_n452.n49 gnd 0.280073f
C5695 a_n2848_n452.n50 gnd 0.008209f
C5696 a_n2848_n452.n51 gnd 0.280073f
C5697 a_n2848_n452.n52 gnd 0.008209f
C5698 a_n2848_n452.n53 gnd 0.280073f
C5699 a_n2848_n452.n54 gnd 0.008209f
C5700 a_n2848_n452.n55 gnd 1.54395f
C5701 a_n2848_n452.n56 gnd 0.280073f
C5702 a_n2848_n452.n57 gnd 0.008507f
C5703 a_n2848_n452.n58 gnd 4.1e-19
C5704 a_n2848_n452.n60 gnd 0.007897f
C5705 a_n2848_n452.n61 gnd 0.280073f
C5706 a_n2848_n452.n62 gnd 0.008507f
C5707 a_n2848_n452.n63 gnd 4.1e-19
C5708 a_n2848_n452.n65 gnd 0.008209f
C5709 a_n2848_n452.n66 gnd 0.011936f
C5710 a_n2848_n452.n67 gnd 0.007897f
C5711 a_n2848_n452.n68 gnd 0.280073f
C5712 a_n2848_n452.n69 gnd 0.296926f
C5713 a_n2848_n452.t25 gnd 1.37696f
C5714 a_n2848_n452.t53 gnd 0.147057f
C5715 a_n2848_n452.t45 gnd 0.147057f
C5716 a_n2848_n452.n71 gnd 1.03587f
C5717 a_n2848_n452.t57 gnd 0.147057f
C5718 a_n2848_n452.t37 gnd 0.147057f
C5719 a_n2848_n452.n72 gnd 1.03587f
C5720 a_n2848_n452.t59 gnd 0.147057f
C5721 a_n2848_n452.t51 gnd 0.147057f
C5722 a_n2848_n452.n73 gnd 1.03587f
C5723 a_n2848_n452.t49 gnd 0.147057f
C5724 a_n2848_n452.t27 gnd 0.147057f
C5725 a_n2848_n452.n74 gnd 1.03587f
C5726 a_n2848_n452.t48 gnd 0.684036f
C5727 a_n2848_n452.n75 gnd 0.297182f
C5728 a_n2848_n452.t58 gnd 0.684036f
C5729 a_n2848_n452.t44 gnd 0.684036f
C5730 a_n2848_n452.n76 gnd 0.30061f
C5731 a_n2848_n452.t24 gnd 0.684036f
C5732 a_n2848_n452.t75 gnd 0.684036f
C5733 a_n2848_n452.n77 gnd 0.297182f
C5734 a_n2848_n452.t90 gnd 0.684036f
C5735 a_n2848_n452.t93 gnd 0.684036f
C5736 a_n2848_n452.n78 gnd 0.30061f
C5737 a_n2848_n452.t70 gnd 0.684036f
C5738 a_n2848_n452.t28 gnd 0.684036f
C5739 a_n2848_n452.t30 gnd 0.684036f
C5740 a_n2848_n452.t40 gnd 0.684036f
C5741 a_n2848_n452.n79 gnd 0.30061f
C5742 a_n2848_n452.t46 gnd 0.684036f
C5743 a_n2848_n452.t38 gnd 0.684036f
C5744 a_n2848_n452.t32 gnd 0.684036f
C5745 a_n2848_n452.t34 gnd 0.684036f
C5746 a_n2848_n452.t98 gnd 0.684036f
C5747 a_n2848_n452.t77 gnd 0.684036f
C5748 a_n2848_n452.t82 gnd 0.684036f
C5749 a_n2848_n452.n80 gnd 0.30061f
C5750 a_n2848_n452.t71 gnd 0.684036f
C5751 a_n2848_n452.t87 gnd 0.684036f
C5752 a_n2848_n452.t95 gnd 0.684036f
C5753 a_n2848_n452.n81 gnd 0.296926f
C5754 a_n2848_n452.t96 gnd 0.684036f
C5755 a_n2848_n452.t66 gnd 0.684036f
C5756 a_n2848_n452.t79 gnd 0.684036f
C5757 a_n2848_n452.n82 gnd 0.300731f
C5758 a_n2848_n452.t69 gnd 0.695498f
C5759 a_n2848_n452.n83 gnd 0.297182f
C5760 a_n2848_n452.n84 gnd 0.291698f
C5761 a_n2848_n452.n85 gnd 0.300746f
C5762 a_n2848_n452.n86 gnd 0.303315f
C5763 a_n2848_n452.n87 gnd 0.2966f
C5764 a_n2848_n452.n88 gnd 0.291534f
C5765 a_n2848_n452.t42 gnd 0.695498f
C5766 a_n2848_n452.t60 gnd 0.684036f
C5767 a_n2848_n452.n89 gnd 0.300731f
C5768 a_n2848_n452.n90 gnd 0.29709f
C5769 a_n2848_n452.n91 gnd 0.012028f
C5770 a_n2848_n452.t54 gnd 0.684036f
C5771 a_n2848_n452.n92 gnd 0.291698f
C5772 a_n2848_n452.t14 gnd 0.114377f
C5773 a_n2848_n452.t18 gnd 0.114377f
C5774 a_n2848_n452.n93 gnd 1.01366f
C5775 a_n2848_n452.t12 gnd 0.114377f
C5776 a_n2848_n452.t11 gnd 0.114377f
C5777 a_n2848_n452.n94 gnd 1.01068f
C5778 a_n2848_n452.t62 gnd 0.114377f
C5779 a_n2848_n452.t1 gnd 0.114377f
C5780 a_n2848_n452.n95 gnd 1.01068f
C5781 a_n2848_n452.t19 gnd 0.114377f
C5782 a_n2848_n452.t15 gnd 0.114377f
C5783 a_n2848_n452.n96 gnd 1.01366f
C5784 a_n2848_n452.t6 gnd 0.114377f
C5785 a_n2848_n452.t21 gnd 0.114377f
C5786 a_n2848_n452.n97 gnd 1.01068f
C5787 a_n2848_n452.t4 gnd 0.114377f
C5788 a_n2848_n452.t5 gnd 0.114377f
C5789 a_n2848_n452.n98 gnd 1.01068f
C5790 a_n2848_n452.t9 gnd 0.114377f
C5791 a_n2848_n452.t20 gnd 0.114377f
C5792 a_n2848_n452.n99 gnd 1.01068f
C5793 a_n2848_n452.t8 gnd 0.114377f
C5794 a_n2848_n452.t2 gnd 0.114377f
C5795 a_n2848_n452.n100 gnd 1.01068f
C5796 a_n2848_n452.t0 gnd 0.114377f
C5797 a_n2848_n452.t7 gnd 0.114377f
C5798 a_n2848_n452.n101 gnd 1.01068f
C5799 a_n2848_n452.t3 gnd 0.114377f
C5800 a_n2848_n452.t63 gnd 0.114377f
C5801 a_n2848_n452.n102 gnd 1.01366f
C5802 a_n2848_n452.t16 gnd 0.114377f
C5803 a_n2848_n452.t17 gnd 0.114377f
C5804 a_n2848_n452.n103 gnd 1.01068f
C5805 a_n2848_n452.t13 gnd 0.114377f
C5806 a_n2848_n452.t10 gnd 0.114377f
C5807 a_n2848_n452.n104 gnd 1.01068f
C5808 a_n2848_n452.n105 gnd 0.012028f
C5809 a_n2848_n452.n106 gnd 0.296926f
C5810 a_n2848_n452.n107 gnd 0.303315f
C5811 a_n2848_n452.n108 gnd 0.2966f
C5812 a_n2848_n452.n109 gnd 0.291534f
C5813 a_n2848_n452.t43 gnd 1.37696f
C5814 a_n2848_n452.t35 gnd 0.147057f
C5815 a_n2848_n452.t61 gnd 0.147057f
C5816 a_n2848_n452.n110 gnd 1.03587f
C5817 a_n2848_n452.t33 gnd 0.147057f
C5818 a_n2848_n452.t55 gnd 0.147057f
C5819 a_n2848_n452.n111 gnd 1.03587f
C5820 a_n2848_n452.t47 gnd 0.147057f
C5821 a_n2848_n452.t39 gnd 0.147057f
C5822 a_n2848_n452.n112 gnd 1.03587f
C5823 a_n2848_n452.t31 gnd 0.147057f
C5824 a_n2848_n452.t41 gnd 0.147057f
C5825 a_n2848_n452.n113 gnd 1.03587f
C5826 a_n2848_n452.t29 gnd 1.37422f
C5827 a_n2848_n452.n114 gnd 1.41993f
C5828 a_n2848_n452.n115 gnd 0.924414f
C5829 a_n2848_n452.t76 gnd 0.684036f
C5830 a_n2848_n452.t86 gnd 0.684036f
C5831 a_n2848_n452.t99 gnd 0.684036f
C5832 a_n2848_n452.n116 gnd 0.300746f
C5833 a_n2848_n452.t88 gnd 0.684036f
C5834 a_n2848_n452.t73 gnd 0.684036f
C5835 a_n2848_n452.t72 gnd 0.684036f
C5836 a_n2848_n452.n117 gnd 0.300746f
C5837 a_n2848_n452.t92 gnd 0.684036f
C5838 a_n2848_n452.t81 gnd 0.684036f
C5839 a_n2848_n452.t80 gnd 0.684036f
C5840 a_n2848_n452.n118 gnd 0.300746f
C5841 a_n2848_n452.t84 gnd 0.684036f
C5842 a_n2848_n452.t74 gnd 0.684036f
C5843 a_n2848_n452.t64 gnd 0.684036f
C5844 a_n2848_n452.n119 gnd 0.300746f
C5845 a_n2848_n452.t89 gnd 0.695498f
C5846 a_n2848_n452.n120 gnd 0.296926f
C5847 a_n2848_n452.n121 gnd 0.291534f
C5848 a_n2848_n452.t97 gnd 0.695498f
C5849 a_n2848_n452.n122 gnd 0.296926f
C5850 a_n2848_n452.n123 gnd 0.291534f
C5851 a_n2848_n452.t83 gnd 0.695498f
C5852 a_n2848_n452.n124 gnd 0.296926f
C5853 a_n2848_n452.n125 gnd 0.291534f
C5854 a_n2848_n452.t78 gnd 0.695498f
C5855 a_n2848_n452.n126 gnd 0.296926f
C5856 a_n2848_n452.n127 gnd 0.291534f
C5857 a_n2848_n452.n128 gnd 1.21807f
C5858 a_n2848_n452.n129 gnd 0.291534f
C5859 a_n2848_n452.t94 gnd 0.684036f
C5860 a_n2848_n452.n130 gnd 0.2966f
C5861 a_n2848_n452.t68 gnd 0.684036f
C5862 a_n2848_n452.n131 gnd 0.303315f
C5863 a_n2848_n452.t91 gnd 0.684036f
C5864 a_n2848_n452.n132 gnd 0.300746f
C5865 a_n2848_n452.n133 gnd 0.296926f
C5866 a_n2848_n452.t65 gnd 0.684036f
C5867 a_n2848_n452.n134 gnd 0.291698f
C5868 a_n2848_n452.t85 gnd 0.684036f
C5869 a_n2848_n452.n135 gnd 0.300731f
C5870 a_n2848_n452.t67 gnd 0.695498f
C5871 a_n2848_n452.n136 gnd 0.291534f
C5872 a_n2848_n452.t52 gnd 0.684036f
C5873 a_n2848_n452.n137 gnd 0.2966f
C5874 a_n2848_n452.t56 gnd 0.684036f
C5875 a_n2848_n452.n138 gnd 0.303315f
C5876 a_n2848_n452.t36 gnd 0.684036f
C5877 a_n2848_n452.n139 gnd 0.300746f
C5878 a_n2848_n452.n140 gnd 0.296926f
C5879 a_n2848_n452.t50 gnd 0.684036f
C5880 a_n2848_n452.n141 gnd 0.291698f
C5881 a_n2848_n452.t26 gnd 0.684036f
C5882 a_n2848_n452.n142 gnd 0.300731f
C5883 a_n2848_n452.t22 gnd 0.695498f
C5884 a_n2848_n452.n143 gnd 1.25017f
C5885 a_n2848_n452.t23 gnd 1.37422f
.ends

