* NGSPICE file created from opamp.ext - technology: sky130A

.subckt opamp output vdd plus minus commonsourceibias outputibias diffpairibias gnd CSoutput
Cload output gnd 0.0p
X0 a_n1986_8322.t20 a_n2848_n452.t48 vdd.t275 vdd.t274 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X1 gnd.t306 gnd.t303 gnd.t305 gnd.t304 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X2 a_n1808_13878.t19 a_n2848_n452.t37 a_n2848_n452.t38 vdd.t271 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X3 outputibias.t7 outputibias.t6 gnd.t180 gnd.t179 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X4 a_n7636_8799.t35 plus.t5 a_n3827_n3924.t42 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X5 vdd.t83 a_n7636_8799.t36 CSoutput.t125 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X6 a_n3827_n3924.t23 diffpairibias.t20 gnd.t312 gnd.t311 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X7 gnd.t353 commonsourceibias.t80 CSoutput.t196 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X8 gnd.t302 gnd.t300 gnd.t301 gnd.t279 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X9 a_n3827_n3924.t41 plus.t6 a_n7636_8799.t34 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X10 commonsourceibias.t79 commonsourceibias.t78 gnd.t152 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X11 commonsourceibias.t77 commonsourceibias.t76 gnd.t328 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X12 a_n2848_n452.t34 a_n2848_n452.t33 a_n1808_13878.t18 vdd.t255 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X13 vdd.t219 vdd.t217 vdd.t218 vdd.t195 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X14 CSoutput.t124 a_n7636_8799.t37 vdd.t84 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X15 gnd.t299 gnd.t297 gnd.t298 gnd.t279 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X16 a_n1808_13878.t17 a_n2848_n452.t25 a_n2848_n452.t26 vdd.t261 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X17 a_n1808_13878.t7 a_n2848_n452.t49 vdd.t273 vdd.t272 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X18 vdd.t79 a_n7636_8799.t38 CSoutput.t123 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X19 CSoutput.t122 a_n7636_8799.t39 vdd.t81 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X20 gnd.t296 gnd.t294 gnd.t295 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X21 CSoutput.t197 commonsourceibias.t81 gnd.t354 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X22 gnd.t10 commonsourceibias.t74 commonsourceibias.t75 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X23 CSoutput.t121 a_n7636_8799.t40 vdd.t89 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X24 CSoutput.t4 commonsourceibias.t82 gnd.t37 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X25 gnd.t293 gnd.t291 gnd.t292 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X26 vdd.t216 vdd.t214 vdd.t215 vdd.t167 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X27 commonsourceibias.t73 commonsourceibias.t72 gnd.t47 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X28 a_n2848_n452.t6 minus.t5 a_n3827_n3924.t8 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X29 a_n1986_8322.t8 a_n2848_n452.t50 a_n7636_8799.t11 vdd.t270 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X30 a_n7636_8799.t33 plus.t7 a_n3827_n3924.t54 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X31 CSoutput.t5 commonsourceibias.t83 gnd.t39 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X32 a_n2848_n452.t45 minus.t6 a_n3827_n3924.t29 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X33 plus.t4 gnd.t288 gnd.t290 gnd.t289 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X34 CSoutput.t120 a_n7636_8799.t41 vdd.t90 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X35 output.t15 CSoutput.t200 vdd.t9 gnd.t44 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X36 vdd.t294 a_n7636_8799.t42 CSoutput.t119 vdd.t224 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X37 commonsourceibias.t71 commonsourceibias.t70 gnd.t189 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X38 vdd.t295 a_n7636_8799.t43 CSoutput.t118 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X39 vdd.t292 a_n7636_8799.t44 CSoutput.t117 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X40 CSoutput.t116 a_n7636_8799.t45 vdd.t293 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X41 a_n3827_n3924.t53 plus.t8 a_n7636_8799.t32 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X42 a_n7636_8799.t10 a_n2848_n452.t51 a_n1986_8322.t7 vdd.t271 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X43 vdd.t290 a_n7636_8799.t46 CSoutput.t115 vdd.t227 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X44 a_n3827_n3924.t16 diffpairibias.t21 gnd.t130 gnd.t129 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X45 CSoutput.t176 commonsourceibias.t84 gnd.t176 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X46 CSoutput.t114 a_n7636_8799.t47 vdd.t291 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X47 a_n3827_n3924.t30 minus.t7 a_n2848_n452.t46 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X48 gnd.t177 commonsourceibias.t85 CSoutput.t177 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X49 gnd.t287 gnd.t285 gnd.t286 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X50 gnd.t23 commonsourceibias.t68 commonsourceibias.t69 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X51 commonsourceibias.t67 commonsourceibias.t66 gnd.t190 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X52 vdd.t213 vdd.t211 vdd.t212 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X53 CSoutput.t113 a_n7636_8799.t48 vdd.t288 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X54 CSoutput.t112 a_n7636_8799.t49 vdd.t289 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X55 gnd.t118 commonsourceibias.t86 CSoutput.t150 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X56 vdd.t10 CSoutput.t201 output.t14 gnd.t45 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X57 gnd.t120 commonsourceibias.t87 CSoutput.t151 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X58 gnd.t284 gnd.t282 gnd.t283 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X59 gnd.t148 commonsourceibias.t88 CSoutput.t166 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X60 CSoutput.t111 a_n7636_8799.t50 vdd.t230 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X61 a_n3827_n3924.t52 plus.t9 a_n7636_8799.t31 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X62 gnd.t329 commonsourceibias.t64 commonsourceibias.t65 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X63 diffpairibias.t19 diffpairibias.t18 gnd.t195 gnd.t194 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X64 a_n3827_n3924.t51 plus.t10 a_n7636_8799.t30 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X65 a_n1808_13878.t16 a_n2848_n452.t43 a_n2848_n452.t44 vdd.t237 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X66 commonsourceibias.t63 commonsourceibias.t62 gnd.t121 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X67 vdd.t231 a_n7636_8799.t51 CSoutput.t110 vdd.t227 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X68 vdd.t210 vdd.t208 vdd.t209 vdd.t167 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X69 a_n3827_n3924.t10 minus.t8 a_n2848_n452.t7 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X70 output.t13 CSoutput.t202 vdd.t11 gnd.t46 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0.825 ps=5.33 w=5 l=1
X71 CSoutput.t109 a_n7636_8799.t52 vdd.t284 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X72 a_n2848_n452.t32 a_n2848_n452.t31 a_n1808_13878.t15 vdd.t247 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X73 CSoutput.t108 a_n7636_8799.t53 vdd.t285 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X74 vdd.t207 vdd.t205 vdd.t206 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X75 commonsourceibias.t61 commonsourceibias.t60 gnd.t178 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X76 vdd.t225 a_n7636_8799.t54 CSoutput.t107 vdd.t224 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X77 gnd.t281 gnd.t278 gnd.t280 gnd.t279 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X78 diffpairibias.t17 diffpairibias.t16 gnd.t3 gnd.t2 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X79 gnd.t41 commonsourceibias.t58 commonsourceibias.t59 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X80 CSoutput.t167 commonsourceibias.t89 gnd.t150 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X81 CSoutput.t106 a_n7636_8799.t55 vdd.t226 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X82 vdd.t286 a_n7636_8799.t56 CSoutput.t105 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X83 vdd.t287 a_n7636_8799.t57 CSoutput.t104 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X84 CSoutput.t182 commonsourceibias.t90 gnd.t185 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X85 vdd.t228 a_n7636_8799.t58 CSoutput.t103 vdd.t227 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X86 vdd.t229 a_n7636_8799.t59 CSoutput.t102 vdd.t72 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X87 CSoutput.t101 a_n7636_8799.t60 vdd.t282 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X88 CSoutput.t100 a_n7636_8799.t61 vdd.t283 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X89 a_n3827_n3924.t7 minus.t9 a_n2848_n452.t5 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X90 gnd.t355 commonsourceibias.t56 commonsourceibias.t57 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X91 CSoutput.t183 commonsourceibias.t91 gnd.t187 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X92 a_n3827_n3924.t46 plus.t11 a_n7636_8799.t29 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X93 CSoutput.t180 commonsourceibias.t92 gnd.t183 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X94 output.t12 CSoutput.t203 vdd.t141 gnd.t334 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X95 vdd.t142 CSoutput.t204 output.t11 gnd.t335 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=1.95 ps=10.78 w=5 l=1
X96 a_n7636_8799.t28 plus.t12 a_n3827_n3924.t45 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X97 CSoutput.t181 commonsourceibias.t93 gnd.t184 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X98 vdd.t222 a_n7636_8799.t62 CSoutput.t99 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X99 CSoutput.t164 commonsourceibias.t94 gnd.t145 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X100 CSoutput.t98 a_n7636_8799.t63 vdd.t223 vdd.t99 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X101 a_n3827_n3924.t13 diffpairibias.t22 gnd.t85 gnd.t84 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X102 CSoutput.t97 a_n7636_8799.t64 vdd.t102 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X103 CSoutput.t96 a_n7636_8799.t65 vdd.t104 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X104 CSoutput.t95 a_n7636_8799.t66 vdd.t100 vdd.t99 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X105 a_n3827_n3924.t48 plus.t13 a_n7636_8799.t27 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X106 vdd.t101 a_n7636_8799.t67 CSoutput.t94 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X107 gnd.t76 commonsourceibias.t54 commonsourceibias.t55 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X108 gnd.t12 commonsourceibias.t52 commonsourceibias.t53 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X109 gnd.t48 commonsourceibias.t50 commonsourceibias.t51 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X110 vdd.t97 a_n7636_8799.t68 CSoutput.t93 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X111 output.t19 outputibias.t8 gnd.t126 gnd.t125 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X112 a_n2848_n452.t22 a_n2848_n452.t21 a_n1808_13878.t14 vdd.t270 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X113 CSoutput.t205 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X114 vdd.t98 a_n7636_8799.t69 CSoutput.t92 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X115 vdd.t220 a_n7636_8799.t70 CSoutput.t91 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X116 a_n7636_8799.t9 a_n2848_n452.t52 a_n1986_8322.t12 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X117 a_n2848_n452.t24 a_n2848_n452.t23 a_n1808_13878.t13 vdd.t232 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X118 gnd.t277 gnd.t274 gnd.t276 gnd.t275 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X119 a_n2848_n452.t18 minus.t10 a_n3827_n3924.t25 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X120 vdd.t221 a_n7636_8799.t71 CSoutput.t90 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X121 diffpairibias.t15 diffpairibias.t14 gnd.t308 gnd.t307 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X122 output.t18 outputibias.t9 gnd.t25 gnd.t24 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X123 gnd.t146 commonsourceibias.t95 CSoutput.t165 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X124 vdd.t127 a_n7636_8799.t72 CSoutput.t89 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X125 gnd.t143 commonsourceibias.t96 CSoutput.t162 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X126 gnd.t144 commonsourceibias.t97 CSoutput.t163 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X127 gnd.t141 commonsourceibias.t98 CSoutput.t160 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X128 CSoutput.t88 a_n7636_8799.t73 vdd.t128 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X129 gnd.t142 commonsourceibias.t99 CSoutput.t161 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X130 gnd.t140 commonsourceibias.t100 CSoutput.t159 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X131 gnd.t273 gnd.t271 gnd.t272 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X132 vdd.t204 vdd.t202 vdd.t203 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X133 vdd.t94 a_n7636_8799.t74 CSoutput.t87 vdd.t72 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X134 a_n3827_n3924.t55 diffpairibias.t23 gnd.t357 gnd.t356 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X135 vdd.t143 CSoutput.t206 output.t10 gnd.t336 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X136 CSoutput.t86 a_n7636_8799.t75 vdd.t96 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X137 vdd.t201 vdd.t198 vdd.t200 vdd.t199 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X138 gnd.t270 gnd.t268 gnd.t269 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X139 CSoutput.t193 commonsourceibias.t101 gnd.t347 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X140 gnd.t267 gnd.t265 minus.t4 gnd.t266 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X141 gnd.t348 commonsourceibias.t48 commonsourceibias.t49 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X142 vdd.t197 vdd.t194 vdd.t196 vdd.t195 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X143 vdd.t193 vdd.t191 vdd.t192 vdd.t184 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X144 vdd.t269 a_n2848_n452.t53 a_n1986_8322.t19 vdd.t268 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X145 gnd.t346 commonsourceibias.t102 CSoutput.t192 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X146 a_n1986_8322.t18 a_n2848_n452.t54 vdd.t267 vdd.t266 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X147 CSoutput.t85 a_n7636_8799.t76 vdd.t106 vdd.t99 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X148 CSoutput.t84 a_n7636_8799.t77 vdd.t107 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X149 vdd.t58 a_n7636_8799.t78 CSoutput.t83 vdd.t57 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X150 gnd.t324 commonsourceibias.t46 commonsourceibias.t47 gnd.t119 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X151 gnd.t264 gnd.t262 plus.t3 gnd.t263 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X152 vdd.t265 a_n2848_n452.t55 a_n1808_13878.t6 vdd.t264 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X153 a_n7636_8799.t26 plus.t14 a_n3827_n3924.t47 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X154 a_n2848_n452.t12 minus.t11 a_n3827_n3924.t17 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X155 vdd.t190 vdd.t187 vdd.t189 vdd.t188 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X156 a_n7636_8799.t25 plus.t15 a_n3827_n3924.t50 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X157 diffpairibias.t13 diffpairibias.t12 gnd.t133 gnd.t132 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X158 CSoutput.t207 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X159 a_n2848_n452.t8 minus.t12 a_n3827_n3924.t11 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X160 CSoutput.t191 commonsourceibias.t103 gnd.t345 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X161 vdd.t186 vdd.t183 vdd.t185 vdd.t184 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X162 vdd.t60 a_n7636_8799.t79 CSoutput.t82 vdd.t59 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X163 CSoutput.t187 commonsourceibias.t104 gnd.t341 gnd.t186 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X164 commonsourceibias.t45 commonsourceibias.t44 gnd.t191 gnd.t149 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X165 CSoutput.t190 commonsourceibias.t105 gnd.t344 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X166 vdd.t182 vdd.t179 vdd.t181 vdd.t180 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X167 a_n7636_8799.t8 a_n2848_n452.t56 a_n1986_8322.t11 vdd.t239 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X168 gnd.t343 commonsourceibias.t106 CSoutput.t189 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X169 CSoutput.t170 commonsourceibias.t107 gnd.t169 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X170 a_n1986_8322.t17 a_n2848_n452.t57 vdd.t263 vdd.t262 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X171 CSoutput.t81 a_n7636_8799.t80 vdd.t124 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X172 vdd.t126 a_n7636_8799.t81 CSoutput.t80 vdd.t125 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X173 vdd.t132 a_n7636_8799.t82 CSoutput.t79 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X174 a_n2848_n452.t36 a_n2848_n452.t35 a_n1808_13878.t12 vdd.t250 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X175 a_n3827_n3924.t26 minus.t13 a_n2848_n452.t19 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X176 CSoutput.t188 commonsourceibias.t108 gnd.t342 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X177 a_n7636_8799.t7 a_n2848_n452.t58 a_n1986_8322.t2 vdd.t261 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X178 CSoutput.t78 a_n7636_8799.t83 vdd.t133 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X179 gnd.t75 commonsourceibias.t109 CSoutput.t138 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X180 gnd.t91 commonsourceibias.t42 commonsourceibias.t43 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X181 a_n1808_13878.t11 a_n2848_n452.t29 a_n2848_n452.t30 vdd.t260 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X182 gnd.t68 commonsourceibias.t110 CSoutput.t134 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X183 a_n2848_n452.t3 minus.t14 a_n3827_n3924.t4 gnd.t29 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X184 a_n3827_n3924.t49 plus.t16 a_n7636_8799.t24 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X185 commonsourceibias.t41 commonsourceibias.t40 gnd.t325 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X186 gnd.t193 commonsourceibias.t38 commonsourceibias.t39 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X187 vdd.t259 a_n2848_n452.t59 a_n1986_8322.t16 vdd.t258 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X188 CSoutput.t77 a_n7636_8799.t84 vdd.t27 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X189 vdd.t29 a_n7636_8799.t85 CSoutput.t76 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X190 gnd.t92 commonsourceibias.t36 commonsourceibias.t37 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X191 a_n3827_n3924.t56 diffpairibias.t24 gnd.t359 gnd.t358 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X192 commonsourceibias.t35 commonsourceibias.t34 gnd.t326 gnd.t38 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X193 a_n3827_n3924.t18 diffpairibias.t25 gnd.t159 gnd.t158 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X194 gnd.t74 commonsourceibias.t111 CSoutput.t137 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X195 a_n7636_8799.t23 plus.t17 a_n3827_n3924.t34 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X196 CSoutput.t75 a_n7636_8799.t86 vdd.t21 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X197 gnd.t66 commonsourceibias.t112 CSoutput.t133 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X198 vdd.t23 a_n7636_8799.t87 CSoutput.t74 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X199 gnd.t73 commonsourceibias.t113 CSoutput.t136 gnd.t40 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X200 gnd.t64 commonsourceibias.t114 CSoutput.t132 gnd.t22 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X201 vdd.t130 a_n7636_8799.t88 CSoutput.t73 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X202 a_n7636_8799.t22 plus.t18 a_n3827_n3924.t33 gnd.t77 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X203 gnd.t170 commonsourceibias.t115 CSoutput.t171 gnd.t9 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X204 CSoutput.t208 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X205 CSoutput.t173 commonsourceibias.t116 gnd.t172 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X206 vdd.t131 a_n7636_8799.t89 CSoutput.t72 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X207 vdd.t122 a_n7636_8799.t90 CSoutput.t71 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X208 commonsourceibias.t33 commonsourceibias.t32 gnd.t93 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X209 vdd.t139 CSoutput.t209 output.t9 gnd.t333 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X210 CSoutput.t168 commonsourceibias.t117 gnd.t165 gnd.t151 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X211 minus.t3 gnd.t259 gnd.t261 gnd.t260 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X212 CSoutput.t210 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X213 gnd.t323 commonsourceibias.t118 CSoutput.t186 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X214 CSoutput.t185 commonsourceibias.t119 gnd.t322 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X215 gnd.t258 gnd.t256 gnd.t257 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X216 diffpairibias.t11 diffpairibias.t10 gnd.t1 gnd.t0 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X217 a_n2848_n452.t13 minus.t15 a_n3827_n3924.t19 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X218 gnd.t321 commonsourceibias.t120 CSoutput.t184 gnd.t192 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X219 output.t17 outputibias.t10 gnd.t95 gnd.t94 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X220 gnd.t69 commonsourceibias.t30 commonsourceibias.t31 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X221 CSoutput.t70 a_n7636_8799.t91 vdd.t123 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X222 gnd.t314 commonsourceibias.t28 commonsourceibias.t29 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X223 a_n3827_n3924.t36 plus.t19 a_n7636_8799.t21 gnd.t161 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X224 CSoutput.t69 a_n7636_8799.t92 vdd.t77 vdd.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X225 CSoutput.t68 a_n7636_8799.t93 vdd.t78 vdd.t70 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X226 commonsourceibias.t27 commonsourceibias.t26 gnd.t108 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X227 CSoutput.t195 commonsourceibias.t121 gnd.t352 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X228 a_n1808_13878.t5 a_n2848_n452.t60 vdd.t236 vdd.t235 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X229 diffpairibias.t9 diffpairibias.t8 gnd.t59 gnd.t58 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X230 vdd.t178 vdd.t176 vdd.t177 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X231 vdd.t257 a_n2848_n452.t61 a_n1808_13878.t4 vdd.t256 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X232 vdd.t175 vdd.t173 vdd.t174 vdd.t160 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X233 CSoutput.t67 a_n7636_8799.t94 vdd.t120 vdd.t26 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X234 gnd.t153 commonsourceibias.t24 commonsourceibias.t25 gnd.t117 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X235 CSoutput.t199 commonsourceibias.t122 gnd.t361 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X236 vdd.t121 a_n7636_8799.t95 CSoutput.t66 vdd.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X237 a_n3827_n3924.t22 minus.t16 a_n2848_n452.t16 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X238 vdd.t172 vdd.t170 vdd.t171 vdd.t160 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X239 diffpairibias.t7 diffpairibias.t6 gnd.t310 gnd.t309 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X240 gnd.t175 commonsourceibias.t123 CSoutput.t175 gnd.t174 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=1
X241 CSoutput.t65 a_n7636_8799.t96 vdd.t45 vdd.t20 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X242 a_n3827_n3924.t2 minus.t17 a_n2848_n452.t2 gnd.t6 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X243 vdd.t46 a_n7636_8799.t97 CSoutput.t64 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X244 vdd.t55 a_n7636_8799.t98 CSoutput.t63 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X245 CSoutput.t169 commonsourceibias.t124 gnd.t168 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X246 a_n3827_n3924.t35 plus.t20 a_n7636_8799.t20 gnd.t62 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X247 CSoutput.t158 commonsourceibias.t125 gnd.t139 gnd.t107 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X248 gnd.t255 gnd.t252 gnd.t254 gnd.t253 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=0 ps=0 w=6 l=2
X249 gnd.t57 commonsourceibias.t126 CSoutput.t130 gnd.t56 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X250 a_n3827_n3924.t27 minus.t18 a_n2848_n452.t20 gnd.t197 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X251 CSoutput.t62 a_n7636_8799.t99 vdd.t56 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X252 a_n1986_8322.t1 a_n2848_n452.t62 a_n7636_8799.t6 vdd.t255 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X253 gnd.t251 gnd.t248 gnd.t250 gnd.t249 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X254 gnd.t138 commonsourceibias.t127 CSoutput.t157 gnd.t67 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X255 vdd.t280 a_n7636_8799.t100 CSoutput.t61 vdd.t224 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X256 CSoutput.t60 a_n7636_8799.t101 vdd.t281 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X257 vdd.t0 CSoutput.t211 output.t8 gnd.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X258 CSoutput.t149 commonsourceibias.t128 gnd.t106 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X259 vdd.t73 a_n7636_8799.t102 CSoutput.t59 vdd.t72 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X260 vdd.t254 a_n2848_n452.t63 a_n1986_8322.t15 vdd.t253 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X261 commonsourceibias.t23 commonsourceibias.t22 gnd.t110 gnd.t109 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X262 vdd.t75 a_n7636_8799.t103 CSoutput.t58 vdd.t74 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X263 CSoutput.t2 commonsourceibias.t129 gnd.t21 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X264 vdd.t34 a_n7636_8799.t104 CSoutput.t57 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X265 gnd.t247 gnd.t244 gnd.t246 gnd.t245 sky130_fd_pr__nfet_01v8_lvt ad=1.95 pd=10.78 as=0 ps=0 w=5 l=1
X266 gnd.t243 gnd.t241 gnd.t242 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X267 a_n1808_13878.t3 a_n2848_n452.t64 vdd.t252 vdd.t251 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X268 a_n3827_n3924.t28 diffpairibias.t26 gnd.t350 gnd.t349 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X269 minus.t2 gnd.t238 gnd.t240 gnd.t239 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X270 a_n7636_8799.t19 plus.t21 a_n3827_n3924.t38 gnd.t28 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X271 gnd.t55 commonsourceibias.t130 CSoutput.t129 gnd.t54 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X272 vdd.t91 a_n7636_8799.t105 CSoutput.t56 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X273 a_n2848_n452.t47 minus.t19 a_n3827_n3924.t57 gnd.t196 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X274 CSoutput.t55 a_n7636_8799.t106 vdd.t92 vdd.t70 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X275 CSoutput.t54 a_n7636_8799.t107 vdd.t135 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X276 a_n3827_n3924.t24 minus.t20 a_n2848_n452.t17 gnd.t313 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=1.155 ps=7.33 w=7 l=0.9
X277 vdd.t169 vdd.t166 vdd.t168 vdd.t167 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X278 gnd.t104 commonsourceibias.t131 CSoutput.t148 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X279 vdd.t165 vdd.t163 vdd.t164 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X280 CSoutput.t3 commonsourceibias.t132 gnd.t35 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X281 a_n1986_8322.t10 a_n2848_n452.t65 a_n7636_8799.t5 vdd.t250 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X282 vdd.t162 vdd.t159 vdd.t161 vdd.t160 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X283 vdd.t249 a_n2848_n452.t66 a_n1986_8322.t14 vdd.t248 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X284 CSoutput.t53 a_n7636_8799.t108 vdd.t71 vdd.t70 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X285 vdd.t119 a_n7636_8799.t109 CSoutput.t52 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X286 CSoutput.t51 a_n7636_8799.t110 vdd.t278 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X287 CSoutput.t135 commonsourceibias.t133 gnd.t72 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X288 a_n3827_n3924.t0 minus.t21 a_n2848_n452.t0 gnd.t4 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X289 vdd.t13 a_n7636_8799.t111 CSoutput.t50 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X290 vdd.t110 a_n7636_8799.t112 CSoutput.t49 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X291 gnd.t53 commonsourceibias.t134 CSoutput.t128 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X292 a_n3827_n3924.t15 minus.t22 a_n2848_n452.t11 gnd.t116 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X293 gnd.t19 commonsourceibias.t135 CSoutput.t1 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X294 CSoutput.t140 commonsourceibias.t136 gnd.t82 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X295 diffpairibias.t5 diffpairibias.t4 gnd.t340 gnd.t339 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X296 output.t7 CSoutput.t212 vdd.t1 gnd.t14 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X297 vdd.t158 vdd.t155 vdd.t157 vdd.t156 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=0 ps=0 w=9 l=0.5
X298 commonsourceibias.t21 commonsourceibias.t20 gnd.t154 gnd.t81 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X299 gnd.t8 commonsourceibias.t137 CSoutput.t0 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X300 CSoutput.t194 commonsourceibias.t138 gnd.t351 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X301 gnd.t315 commonsourceibias.t18 commonsourceibias.t19 gnd.t65 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X302 vdd.t53 a_n7636_8799.t113 CSoutput.t48 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X303 CSoutput.t47 a_n7636_8799.t114 vdd.t118 vdd.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X304 a_n3827_n3924.t9 diffpairibias.t27 gnd.t61 gnd.t60 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X305 CSoutput.t46 a_n7636_8799.t115 vdd.t69 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X306 a_n1808_13878.t10 a_n2848_n452.t27 a_n2848_n452.t28 vdd.t242 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X307 CSoutput.t198 commonsourceibias.t139 gnd.t360 gnd.t188 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X308 a_n1986_8322.t9 a_n2848_n452.t67 a_n7636_8799.t4 vdd.t247 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X309 CSoutput.t213 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X310 gnd.t237 gnd.t234 gnd.t236 gnd.t235 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X311 CSoutput.t174 commonsourceibias.t140 gnd.t173 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X312 a_n3827_n3924.t12 minus.t23 a_n2848_n452.t9 gnd.t83 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X313 CSoutput.t45 a_n7636_8799.t116 vdd.t44 vdd.t43 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X314 CSoutput.t44 a_n7636_8799.t117 vdd.t42 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X315 vdd.t12 a_n7636_8799.t118 CSoutput.t43 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X316 gnd.t316 commonsourceibias.t16 commonsourceibias.t17 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X317 output.t16 outputibias.t11 gnd.t163 gnd.t162 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X318 CSoutput.t156 commonsourceibias.t141 gnd.t137 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X319 vdd.t17 a_n7636_8799.t119 CSoutput.t42 vdd.t16 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X320 a_n1986_8322.t13 a_n2848_n452.t68 vdd.t246 vdd.t245 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X321 gnd.t136 commonsourceibias.t142 CSoutput.t155 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X322 CSoutput.t41 a_n7636_8799.t120 vdd.t4 vdd.t3 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X323 gnd.t233 gnd.t230 gnd.t232 gnd.t231 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=0.9
X324 output.t6 CSoutput.t214 vdd.t2 gnd.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X325 gnd.t229 gnd.t227 plus.t2 gnd.t228 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X326 CSoutput.t147 commonsourceibias.t143 gnd.t103 gnd.t102 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X327 commonsourceibias.t15 commonsourceibias.t14 gnd.t112 gnd.t111 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=1
X328 vdd.t244 a_n2848_n452.t69 a_n1808_13878.t2 vdd.t243 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X329 commonsourceibias.t13 commonsourceibias.t12 gnd.t71 gnd.t70 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X330 CSoutput.t40 a_n7636_8799.t121 vdd.t25 vdd.t24 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X331 CSoutput.t152 commonsourceibias.t144 gnd.t128 gnd.t105 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X332 gnd.t317 commonsourceibias.t10 commonsourceibias.t11 gnd.t18 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X333 CSoutput.t39 a_n7636_8799.t122 vdd.t277 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X334 gnd.t101 commonsourceibias.t145 CSoutput.t146 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X335 CSoutput.t154 commonsourceibias.t146 gnd.t135 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X336 vdd.t8 a_n7636_8799.t123 CSoutput.t38 vdd.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X337 output.t5 CSoutput.t215 vdd.t47 gnd.t122 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X338 vdd.t109 a_n7636_8799.t124 CSoutput.t37 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X339 vdd.t48 CSoutput.t216 output.t4 gnd.t123 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X340 vdd.t154 vdd.t151 vdd.t153 vdd.t152 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X341 gnd.t226 gnd.t223 gnd.t225 gnd.t224 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X342 a_n3827_n3924.t37 plus.t22 a_n7636_8799.t18 gnd.t33 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X343 a_n1986_8322.t4 a_n2848_n452.t70 a_n7636_8799.t3 vdd.t238 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X344 vdd.t150 vdd.t148 vdd.t149 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X345 commonsourceibias.t9 commonsourceibias.t8 gnd.t114 gnd.t113 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X346 a_n2848_n452.t15 minus.t24 a_n3827_n3924.t21 gnd.t96 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X347 CSoutput.t36 a_n7636_8799.t125 vdd.t51 vdd.t50 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X348 a_n7636_8799.t2 a_n2848_n452.t71 a_n1986_8322.t3 vdd.t242 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X349 a_n7636_8799.t17 plus.t23 a_n3827_n3924.t44 gnd.t78 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X350 gnd.t222 gnd.t220 minus.t1 gnd.t221 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X351 vdd.t19 a_n7636_8799.t126 CSoutput.t35 vdd.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X352 a_n1808_13878.t1 a_n2848_n452.t72 vdd.t241 vdd.t240 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X353 a_n2848_n452.t14 minus.t25 a_n3827_n3924.t20 gnd.t160 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X354 vdd.t140 a_n7636_8799.t127 CSoutput.t34 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X355 gnd.t155 commonsourceibias.t6 commonsourceibias.t7 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X356 CSoutput.t33 a_n7636_8799.t128 vdd.t33 vdd.t32 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X357 commonsourceibias.t5 commonsourceibias.t4 gnd.t318 gnd.t20 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X358 gnd.t99 commonsourceibias.t147 CSoutput.t145 gnd.t11 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X359 CSoutput.t153 commonsourceibias.t148 gnd.t134 gnd.t34 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X360 CSoutput.t217 a_n1986_8322.t0 sky130_fd_pr__cap_mim_m3_1 l=12 w=12
X361 gnd.t98 commonsourceibias.t149 CSoutput.t144 gnd.t97 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X362 vdd.t112 a_n7636_8799.t129 CSoutput.t32 vdd.t54 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X363 CSoutput.t31 a_n7636_8799.t130 vdd.t111 vdd.t41 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X364 CSoutput.t30 a_n7636_8799.t131 vdd.t129 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X365 CSoutput.t29 a_n7636_8799.t132 vdd.t31 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X366 CSoutput.t28 a_n7636_8799.t133 vdd.t276 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X367 a_n3827_n3924.t6 minus.t26 a_n2848_n452.t4 gnd.t32 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X368 a_n1808_13878.t9 a_n2848_n452.t41 a_n2848_n452.t42 vdd.t239 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=1.485 ps=9.33 w=9 l=0.5
X369 a_n3827_n3924.t3 diffpairibias.t28 gnd.t27 gnd.t26 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X370 gnd.t63 commonsourceibias.t150 CSoutput.t131 gnd.t52 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X371 vdd.t279 a_n7636_8799.t134 CSoutput.t27 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X372 output.t3 CSoutput.t218 vdd.t49 gnd.t124 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X373 gnd.t219 gnd.t216 gnd.t218 gnd.t217 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X374 a_n7636_8799.t16 plus.t24 a_n3827_n3924.t43 gnd.t127 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X375 gnd.t51 commonsourceibias.t151 CSoutput.t127 gnd.t7 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X376 CSoutput.t26 a_n7636_8799.t135 vdd.t108 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X377 gnd.t215 gnd.t212 gnd.t214 gnd.t213 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X378 CSoutput.t143 commonsourceibias.t152 gnd.t90 gnd.t36 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X379 CSoutput.t139 commonsourceibias.t153 gnd.t80 gnd.t79 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X380 commonsourceibias.t3 commonsourceibias.t2 gnd.t157 gnd.t156 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X381 vdd.t68 a_n7636_8799.t136 CSoutput.t25 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X382 outputibias.t5 outputibias.t4 gnd.t320 gnd.t319 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X383 vdd.t66 a_n7636_8799.t137 CSoutput.t24 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X384 diffpairibias.t3 diffpairibias.t2 gnd.t338 gnd.t337 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X385 output.t2 CSoutput.t219 vdd.t136 gnd.t330 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X386 CSoutput.t23 a_n7636_8799.t138 vdd.t40 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X387 a_n2848_n452.t40 a_n2848_n452.t39 a_n1808_13878.t8 vdd.t238 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X388 a_n2848_n452.t10 minus.t27 a_n3827_n3924.t14 gnd.t115 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X389 vdd.t93 a_n7636_8799.t139 CSoutput.t22 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X390 a_n7636_8799.t1 a_n2848_n452.t73 a_n1986_8322.t6 vdd.t237 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X391 gnd.t211 gnd.t209 plus.t1 gnd.t210 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X392 CSoutput.t21 a_n7636_8799.t140 vdd.t105 vdd.t95 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X393 vdd.t117 a_n7636_8799.t141 CSoutput.t20 vdd.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X394 outputibias.t3 outputibias.t2 gnd.t17 gnd.t16 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X395 diffpairibias.t1 diffpairibias.t0 gnd.t363 gnd.t362 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X396 vdd.t116 a_n7636_8799.t142 CSoutput.t19 vdd.t115 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X397 vdd.t147 vdd.t144 vdd.t146 vdd.t145 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.5
X398 CSoutput.t18 a_n7636_8799.t143 vdd.t65 vdd.t64 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X399 CSoutput.t126 commonsourceibias.t154 gnd.t50 gnd.t49 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X400 outputibias.t1 outputibias.t0 gnd.t167 gnd.t166 sky130_fd_pr__nfet_01v8 ad=2.34 pd=12.78 as=2.34 ps=12.78 w=6 l=2
X401 vdd.t38 a_n7636_8799.t144 CSoutput.t17 vdd.t37 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X402 gnd.t89 commonsourceibias.t155 CSoutput.t142 gnd.t88 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X403 plus.t0 gnd.t206 gnd.t208 gnd.t207 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X404 CSoutput.t179 commonsourceibias.t156 gnd.t182 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X405 gnd.t87 commonsourceibias.t157 CSoutput.t141 gnd.t86 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X406 a_n7636_8799.t15 plus.t25 a_n3827_n3924.t32 gnd.t164 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X407 gnd.t205 gnd.t202 gnd.t204 gnd.t203 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=0 ps=0 w=7 l=1
X408 gnd.t201 gnd.t199 minus.t0 gnd.t200 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X409 vdd.t137 CSoutput.t220 output.t1 gnd.t331 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X410 a_n2848_n452.t1 minus.t28 a_n3827_n3924.t1 gnd.t5 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=2.73 ps=14.78 w=7 l=0.9
X411 vdd.t234 a_n2848_n452.t74 a_n1808_13878.t0 vdd.t233 sky130_fd_pr__pfet_01v8_lvt ad=1.485 pd=9.33 as=3.51 ps=18.78 w=9 l=0.5
X412 gnd.t181 commonsourceibias.t158 CSoutput.t178 gnd.t100 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X413 a_n7636_8799.t14 plus.t26 a_n3827_n3924.t31 gnd.t131 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X414 CSoutput.t16 a_n7636_8799.t145 vdd.t36 vdd.t30 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X415 CSoutput.t15 a_n7636_8799.t146 vdd.t6 vdd.t5 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X416 vdd.t86 a_n7636_8799.t147 CSoutput.t14 vdd.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X417 vdd.t88 a_n7636_8799.t148 CSoutput.t13 vdd.t87 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X418 CSoutput.t12 a_n7636_8799.t149 vdd.t15 vdd.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X419 gnd.t171 commonsourceibias.t159 CSoutput.t172 gnd.t147 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X420 vdd.t138 CSoutput.t221 output.t0 gnd.t332 sky130_fd_pr__nfet_01v8_lvt ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=1
X421 CSoutput.t11 a_n7636_8799.t150 vdd.t134 vdd.t80 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X422 a_n1986_8322.t5 a_n2848_n452.t75 a_n7636_8799.t0 vdd.t232 sky130_fd_pr__pfet_01v8_lvt ad=3.51 pd=18.78 as=1.485 ps=9.33 w=9 l=0.5
X423 commonsourceibias.t1 commonsourceibias.t0 gnd.t43 gnd.t42 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=1
X424 a_n3827_n3924.t40 plus.t27 a_n7636_8799.t13 gnd.t198 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
X425 vdd.t63 a_n7636_8799.t151 CSoutput.t10 vdd.t52 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X426 vdd.t114 a_n7636_8799.t152 CSoutput.t9 vdd.t67 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X427 a_n3827_n3924.t5 diffpairibias.t29 gnd.t31 gnd.t30 sky130_fd_pr__nfet_01v8 ad=2.73 pd=14.78 as=2.73 ps=14.78 w=7 l=1
X428 CSoutput.t8 a_n7636_8799.t153 vdd.t62 vdd.t61 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=3.12 ps=16.78 w=8 l=0.5
X429 vdd.t35 a_n7636_8799.t154 CSoutput.t7 vdd.t22 sky130_fd_pr__pfet_01v8_lvt ad=3.12 pd=16.78 as=1.32 ps=8.33 w=8 l=0.5
X430 CSoutput.t6 a_n7636_8799.t155 vdd.t113 vdd.t39 sky130_fd_pr__pfet_01v8_lvt ad=1.32 pd=8.33 as=1.32 ps=8.33 w=8 l=0.5
X431 a_n3827_n3924.t39 plus.t28 a_n7636_8799.t12 gnd.t327 sky130_fd_pr__nfet_01v8 ad=1.155 pd=7.33 as=1.155 ps=7.33 w=7 l=0.9
R0 a_n2848_n452.n5 a_n2848_n452.t75 539.01
R1 a_n2848_n452.n97 a_n2848_n452.t58 512.366
R2 a_n2848_n452.n96 a_n2848_n452.t62 512.366
R3 a_n2848_n452.n70 a_n2848_n452.t52 512.366
R4 a_n2848_n452.n95 a_n2848_n452.t67 512.366
R5 a_n2848_n452.n1 a_n2848_n452.t39 533.058
R6 a_n2848_n452.n101 a_n2848_n452.t27 512.366
R7 a_n2848_n452.n100 a_n2848_n452.t21 512.366
R8 a_n2848_n452.n69 a_n2848_n452.t41 512.366
R9 a_n2848_n452.n98 a_n2848_n452.t35 512.366
R10 a_n2848_n452.n19 a_n2848_n452.t23 539.01
R11 a_n2848_n452.n78 a_n2848_n452.t25 512.366
R12 a_n2848_n452.n79 a_n2848_n452.t33 512.366
R13 a_n2848_n452.n73 a_n2848_n452.t29 512.366
R14 a_n2848_n452.n80 a_n2848_n452.t31 512.366
R15 a_n2848_n452.n23 a_n2848_n452.t70 539.01
R16 a_n2848_n452.n75 a_n2848_n452.t71 512.366
R17 a_n2848_n452.n76 a_n2848_n452.t50 512.366
R18 a_n2848_n452.n74 a_n2848_n452.t56 512.366
R19 a_n2848_n452.n77 a_n2848_n452.t65 512.366
R20 a_n2848_n452.n92 a_n2848_n452.t64 512.366
R21 a_n2848_n452.n82 a_n2848_n452.t55 512.366
R22 a_n2848_n452.n93 a_n2848_n452.t49 512.366
R23 a_n2848_n452.n90 a_n2848_n452.t72 512.366
R24 a_n2848_n452.n83 a_n2848_n452.t61 512.366
R25 a_n2848_n452.n91 a_n2848_n452.t60 512.366
R26 a_n2848_n452.n88 a_n2848_n452.t68 512.366
R27 a_n2848_n452.n84 a_n2848_n452.t53 512.366
R28 a_n2848_n452.n89 a_n2848_n452.t54 512.366
R29 a_n2848_n452.n86 a_n2848_n452.t57 512.366
R30 a_n2848_n452.n85 a_n2848_n452.t66 512.366
R31 a_n2848_n452.n87 a_n2848_n452.t48 512.366
R32 a_n2848_n452.n50 a_n2848_n452.n3 70.3058
R33 a_n2848_n452.n47 a_n2848_n452.n6 70.3058
R34 a_n2848_n452.n16 a_n2848_n452.n37 70.3058
R35 a_n2848_n452.n20 a_n2848_n452.n34 70.3058
R36 a_n2848_n452.n33 a_n2848_n452.n21 70.1674
R37 a_n2848_n452.n33 a_n2848_n452.n74 20.9683
R38 a_n2848_n452.n21 a_n2848_n452.n32 75.0448
R39 a_n2848_n452.n76 a_n2848_n452.n32 11.2134
R40 a_n2848_n452.n22 a_n2848_n452.n23 44.8194
R41 a_n2848_n452.n36 a_n2848_n452.n17 70.1674
R42 a_n2848_n452.n36 a_n2848_n452.n73 20.9683
R43 a_n2848_n452.n17 a_n2848_n452.n35 75.0448
R44 a_n2848_n452.n79 a_n2848_n452.n35 11.2134
R45 a_n2848_n452.n18 a_n2848_n452.n19 44.8194
R46 a_n2848_n452.n7 a_n2848_n452.n45 70.1674
R47 a_n2848_n452.n9 a_n2848_n452.n43 70.1674
R48 a_n2848_n452.n11 a_n2848_n452.n41 70.1674
R49 a_n2848_n452.n14 a_n2848_n452.n39 70.1674
R50 a_n2848_n452.n87 a_n2848_n452.n39 20.9683
R51 a_n2848_n452.n38 a_n2848_n452.n15 75.0448
R52 a_n2848_n452.n38 a_n2848_n452.n85 11.2134
R53 a_n2848_n452.n15 a_n2848_n452.n86 161.3
R54 a_n2848_n452.n89 a_n2848_n452.n41 20.9683
R55 a_n2848_n452.n40 a_n2848_n452.n12 75.0448
R56 a_n2848_n452.n40 a_n2848_n452.n84 11.2134
R57 a_n2848_n452.n12 a_n2848_n452.n88 161.3
R58 a_n2848_n452.n91 a_n2848_n452.n43 20.9683
R59 a_n2848_n452.n42 a_n2848_n452.n10 75.0448
R60 a_n2848_n452.n42 a_n2848_n452.n83 11.2134
R61 a_n2848_n452.n10 a_n2848_n452.n90 161.3
R62 a_n2848_n452.n93 a_n2848_n452.n45 20.9683
R63 a_n2848_n452.n44 a_n2848_n452.n8 75.0448
R64 a_n2848_n452.n44 a_n2848_n452.n82 11.2134
R65 a_n2848_n452.n8 a_n2848_n452.n92 161.3
R66 a_n2848_n452.n6 a_n2848_n452.n46 70.1674
R67 a_n2848_n452.n46 a_n2848_n452.n69 20.9683
R68 a_n2848_n452.n99 a_n2848_n452.n0 161.3
R69 a_n2848_n452.n4 a_n2848_n452.n49 70.1674
R70 a_n2848_n452.n49 a_n2848_n452.n70 20.9683
R71 a_n2848_n452.n48 a_n2848_n452.n4 75.0448
R72 a_n2848_n452.n96 a_n2848_n452.n48 11.2134
R73 a_n2848_n452.n2 a_n2848_n452.n5 44.8194
R74 a_n2848_n452.n100 a_n2848_n452.n51 20.9683
R75 a_n2848_n452.n51 a_n2848_n452.n0 70.1674
R76 a_n2848_n452.n0 a_n2848_n452.n1 70.3058
R77 a_n2848_n452.n67 a_n2848_n452.n65 81.4626
R78 a_n2848_n452.n58 a_n2848_n452.n56 81.4626
R79 a_n2848_n452.n54 a_n2848_n452.n52 81.4626
R80 a_n2848_n452.n67 a_n2848_n452.n66 80.9324
R81 a_n2848_n452.n31 a_n2848_n452.n68 80.9324
R82 a_n2848_n452.n30 a_n2848_n452.n64 80.9324
R83 a_n2848_n452.n63 a_n2848_n452.n62 80.9324
R84 a_n2848_n452.n61 a_n2848_n452.n60 80.9324
R85 a_n2848_n452.n58 a_n2848_n452.n57 80.9324
R86 a_n2848_n452.n29 a_n2848_n452.n59 80.9324
R87 a_n2848_n452.n28 a_n2848_n452.n55 80.9324
R88 a_n2848_n452.n54 a_n2848_n452.n53 80.9324
R89 a_n2848_n452.n27 a_n2848_n452.t38 74.6477
R90 a_n2848_n452.n24 a_n2848_n452.t24 74.6477
R91 a_n2848_n452.n26 a_n2848_n452.t40 74.2899
R92 a_n2848_n452.n25 a_n2848_n452.t44 74.2897
R93 a_n2848_n452.n27 a_n2848_n452.n103 70.6783
R94 a_n2848_n452.n25 a_n2848_n452.n72 70.6783
R95 a_n2848_n452.n24 a_n2848_n452.n71 70.6783
R96 a_n2848_n452.n104 a_n2848_n452.n27 70.6782
R97 a_n2848_n452.n97 a_n2848_n452.n96 48.2005
R98 a_n2848_n452.n95 a_n2848_n452.n49 20.9683
R99 a_n2848_n452.n101 a_n2848_n452.n51 20.9683
R100 a_n2848_n452.n98 a_n2848_n452.n46 20.9683
R101 a_n2848_n452.n79 a_n2848_n452.n78 48.2005
R102 a_n2848_n452.n80 a_n2848_n452.n36 20.9683
R103 a_n2848_n452.n76 a_n2848_n452.n75 48.2005
R104 a_n2848_n452.n77 a_n2848_n452.n33 20.9683
R105 a_n2848_n452.n92 a_n2848_n452.n82 48.2005
R106 a_n2848_n452.t69 a_n2848_n452.n45 533.335
R107 a_n2848_n452.n90 a_n2848_n452.n83 48.2005
R108 a_n2848_n452.t74 a_n2848_n452.n43 533.335
R109 a_n2848_n452.n88 a_n2848_n452.n84 48.2005
R110 a_n2848_n452.t63 a_n2848_n452.n41 533.335
R111 a_n2848_n452.n86 a_n2848_n452.n85 48.2005
R112 a_n2848_n452.t59 a_n2848_n452.n39 533.335
R113 a_n2848_n452.n50 a_n2848_n452.t73 533.058
R114 a_n2848_n452.n47 a_n2848_n452.t37 533.058
R115 a_n2848_n452.t43 a_n2848_n452.n37 533.058
R116 a_n2848_n452.t51 a_n2848_n452.n34 533.058
R117 a_n2848_n452.n61 a_n2848_n452.n29 33.585
R118 a_n2848_n452.n48 a_n2848_n452.n70 35.3134
R119 a_n2848_n452.n100 a_n2848_n452.n99 24.1005
R120 a_n2848_n452.n99 a_n2848_n452.n69 24.1005
R121 a_n2848_n452.n73 a_n2848_n452.n35 35.3134
R122 a_n2848_n452.n74 a_n2848_n452.n32 35.3134
R123 a_n2848_n452.n93 a_n2848_n452.n44 35.3134
R124 a_n2848_n452.n91 a_n2848_n452.n42 35.3134
R125 a_n2848_n452.n89 a_n2848_n452.n40 35.3134
R126 a_n2848_n452.n87 a_n2848_n452.n38 35.3134
R127 a_n2848_n452.n0 a_n2848_n452.n31 23.891
R128 a_n2848_n452.n22 a_n2848_n452.n13 12.046
R129 a_n2848_n452.n3 a_n2848_n452.n94 11.8414
R130 a_n2848_n452.n102 a_n2848_n452.n0 10.5365
R131 a_n2848_n452.n81 a_n2848_n452.n25 9.50122
R132 a_n2848_n452.n15 a_n2848_n452.n13 7.47588
R133 a_n2848_n452.n94 a_n2848_n452.n7 7.47588
R134 a_n2848_n452.n81 a_n2848_n452.n16 6.70126
R135 a_n2848_n452.n26 a_n2848_n452.n102 5.65783
R136 a_n2848_n452.n94 a_n2848_n452.n81 5.3452
R137 a_n2848_n452.n18 a_n2848_n452.n20 3.95126
R138 a_n2848_n452.n6 a_n2848_n452.n2 3.95126
R139 a_n2848_n452.n103 a_n2848_n452.t42 3.61217
R140 a_n2848_n452.n103 a_n2848_n452.t36 3.61217
R141 a_n2848_n452.n72 a_n2848_n452.t30 3.61217
R142 a_n2848_n452.n72 a_n2848_n452.t32 3.61217
R143 a_n2848_n452.n71 a_n2848_n452.t26 3.61217
R144 a_n2848_n452.n71 a_n2848_n452.t34 3.61217
R145 a_n2848_n452.n104 a_n2848_n452.t28 3.61217
R146 a_n2848_n452.t22 a_n2848_n452.n104 3.61217
R147 a_n2848_n452.n65 a_n2848_n452.t9 2.82907
R148 a_n2848_n452.n65 a_n2848_n452.t1 2.82907
R149 a_n2848_n452.n66 a_n2848_n452.t16 2.82907
R150 a_n2848_n452.n66 a_n2848_n452.t13 2.82907
R151 a_n2848_n452.n68 a_n2848_n452.t46 2.82907
R152 a_n2848_n452.n68 a_n2848_n452.t45 2.82907
R153 a_n2848_n452.n64 a_n2848_n452.t11 2.82907
R154 a_n2848_n452.n64 a_n2848_n452.t47 2.82907
R155 a_n2848_n452.n62 a_n2848_n452.t20 2.82907
R156 a_n2848_n452.n62 a_n2848_n452.t14 2.82907
R157 a_n2848_n452.n60 a_n2848_n452.t7 2.82907
R158 a_n2848_n452.n60 a_n2848_n452.t8 2.82907
R159 a_n2848_n452.n56 a_n2848_n452.t19 2.82907
R160 a_n2848_n452.n56 a_n2848_n452.t18 2.82907
R161 a_n2848_n452.n57 a_n2848_n452.t2 2.82907
R162 a_n2848_n452.n57 a_n2848_n452.t12 2.82907
R163 a_n2848_n452.n59 a_n2848_n452.t0 2.82907
R164 a_n2848_n452.n59 a_n2848_n452.t15 2.82907
R165 a_n2848_n452.n55 a_n2848_n452.t4 2.82907
R166 a_n2848_n452.n55 a_n2848_n452.t10 2.82907
R167 a_n2848_n452.n53 a_n2848_n452.t5 2.82907
R168 a_n2848_n452.n53 a_n2848_n452.t6 2.82907
R169 a_n2848_n452.n52 a_n2848_n452.t17 2.82907
R170 a_n2848_n452.n52 a_n2848_n452.t3 2.82907
R171 a_n2848_n452.n102 a_n2848_n452.n13 1.30542
R172 a_n2848_n452.n10 a_n2848_n452.n11 1.04595
R173 a_n2848_n452.n5 a_n2848_n452.n97 13.657
R174 a_n2848_n452.n95 a_n2848_n452.n50 21.4216
R175 a_n2848_n452.n1 a_n2848_n452.n101 21.4216
R176 a_n2848_n452.n98 a_n2848_n452.n47 21.4216
R177 a_n2848_n452.n78 a_n2848_n452.n19 13.657
R178 a_n2848_n452.n37 a_n2848_n452.n80 21.4216
R179 a_n2848_n452.n75 a_n2848_n452.n23 13.657
R180 a_n2848_n452.n34 a_n2848_n452.n77 21.4216
R181 a_n2848_n452.n0 a_n2848_n452.n6 1.47777
R182 a_n2848_n452.n22 a_n2848_n452.n21 0.758076
R183 a_n2848_n452.n21 a_n2848_n452.n20 0.758076
R184 a_n2848_n452.n18 a_n2848_n452.n17 0.758076
R185 a_n2848_n452.n17 a_n2848_n452.n16 0.758076
R186 a_n2848_n452.n15 a_n2848_n452.n14 0.758076
R187 a_n2848_n452.n12 a_n2848_n452.n11 0.758076
R188 a_n2848_n452.n10 a_n2848_n452.n9 0.758076
R189 a_n2848_n452.n8 a_n2848_n452.n7 0.758076
R190 a_n2848_n452.n4 a_n2848_n452.n2 0.758076
R191 a_n2848_n452.n4 a_n2848_n452.n3 0.758076
R192 a_n2848_n452.n27 a_n2848_n452.n26 0.716017
R193 a_n2848_n452.n25 a_n2848_n452.n24 0.716017
R194 a_n2848_n452.n12 a_n2848_n452.n14 0.67853
R195 a_n2848_n452.n8 a_n2848_n452.n9 0.67853
R196 a_n2848_n452.n28 a_n2848_n452.n54 0.530672
R197 a_n2848_n452.n29 a_n2848_n452.n58 0.530672
R198 a_n2848_n452.n63 a_n2848_n452.n61 0.530672
R199 a_n2848_n452.n30 a_n2848_n452.n63 0.530672
R200 a_n2848_n452.n31 a_n2848_n452.n67 0.530672
R201 a_n2848_n452.n31 a_n2848_n452.n30 0.530672
R202 a_n2848_n452.n29 a_n2848_n452.n28 0.530672
R203 vdd.n327 vdd.n291 756.745
R204 vdd.n268 vdd.n232 756.745
R205 vdd.n225 vdd.n189 756.745
R206 vdd.n166 vdd.n130 756.745
R207 vdd.n124 vdd.n88 756.745
R208 vdd.n65 vdd.n29 756.745
R209 vdd.n1746 vdd.n1710 756.745
R210 vdd.n1805 vdd.n1769 756.745
R211 vdd.n1644 vdd.n1608 756.745
R212 vdd.n1703 vdd.n1667 756.745
R213 vdd.n1543 vdd.n1507 756.745
R214 vdd.n1602 vdd.n1566 756.745
R215 vdd.n2177 vdd.t194 640.208
R216 vdd.n965 vdd.t179 640.208
R217 vdd.n2151 vdd.t217 640.208
R218 vdd.n957 vdd.t205 640.208
R219 vdd.n2922 vdd.t155 640.208
R220 vdd.n2642 vdd.t202 640.208
R221 vdd.n832 vdd.t183 640.208
R222 vdd.n2639 vdd.t187 640.208
R223 vdd.n799 vdd.t191 640.208
R224 vdd.n1027 vdd.t198 640.208
R225 vdd.n1317 vdd.t170 592.009
R226 vdd.n1355 vdd.t159 592.009
R227 vdd.n1251 vdd.t173 592.009
R228 vdd.n2333 vdd.t151 592.009
R229 vdd.n1970 vdd.t163 592.009
R230 vdd.n1930 vdd.t176 592.009
R231 vdd.n426 vdd.t166 592.009
R232 vdd.n440 vdd.t208 592.009
R233 vdd.n452 vdd.t214 592.009
R234 vdd.n768 vdd.t144 592.009
R235 vdd.n3184 vdd.t148 592.009
R236 vdd.n688 vdd.t211 592.009
R237 vdd.n328 vdd.n327 585
R238 vdd.n326 vdd.n293 585
R239 vdd.n325 vdd.n324 585
R240 vdd.n296 vdd.n294 585
R241 vdd.n319 vdd.n318 585
R242 vdd.n317 vdd.n316 585
R243 vdd.n300 vdd.n299 585
R244 vdd.n311 vdd.n310 585
R245 vdd.n309 vdd.n308 585
R246 vdd.n304 vdd.n303 585
R247 vdd.n269 vdd.n268 585
R248 vdd.n267 vdd.n234 585
R249 vdd.n266 vdd.n265 585
R250 vdd.n237 vdd.n235 585
R251 vdd.n260 vdd.n259 585
R252 vdd.n258 vdd.n257 585
R253 vdd.n241 vdd.n240 585
R254 vdd.n252 vdd.n251 585
R255 vdd.n250 vdd.n249 585
R256 vdd.n245 vdd.n244 585
R257 vdd.n226 vdd.n225 585
R258 vdd.n224 vdd.n191 585
R259 vdd.n223 vdd.n222 585
R260 vdd.n194 vdd.n192 585
R261 vdd.n217 vdd.n216 585
R262 vdd.n215 vdd.n214 585
R263 vdd.n198 vdd.n197 585
R264 vdd.n209 vdd.n208 585
R265 vdd.n207 vdd.n206 585
R266 vdd.n202 vdd.n201 585
R267 vdd.n167 vdd.n166 585
R268 vdd.n165 vdd.n132 585
R269 vdd.n164 vdd.n163 585
R270 vdd.n135 vdd.n133 585
R271 vdd.n158 vdd.n157 585
R272 vdd.n156 vdd.n155 585
R273 vdd.n139 vdd.n138 585
R274 vdd.n150 vdd.n149 585
R275 vdd.n148 vdd.n147 585
R276 vdd.n143 vdd.n142 585
R277 vdd.n125 vdd.n124 585
R278 vdd.n123 vdd.n90 585
R279 vdd.n122 vdd.n121 585
R280 vdd.n93 vdd.n91 585
R281 vdd.n116 vdd.n115 585
R282 vdd.n114 vdd.n113 585
R283 vdd.n97 vdd.n96 585
R284 vdd.n108 vdd.n107 585
R285 vdd.n106 vdd.n105 585
R286 vdd.n101 vdd.n100 585
R287 vdd.n66 vdd.n65 585
R288 vdd.n64 vdd.n31 585
R289 vdd.n63 vdd.n62 585
R290 vdd.n34 vdd.n32 585
R291 vdd.n57 vdd.n56 585
R292 vdd.n55 vdd.n54 585
R293 vdd.n38 vdd.n37 585
R294 vdd.n49 vdd.n48 585
R295 vdd.n47 vdd.n46 585
R296 vdd.n42 vdd.n41 585
R297 vdd.n1747 vdd.n1746 585
R298 vdd.n1745 vdd.n1712 585
R299 vdd.n1744 vdd.n1743 585
R300 vdd.n1715 vdd.n1713 585
R301 vdd.n1738 vdd.n1737 585
R302 vdd.n1736 vdd.n1735 585
R303 vdd.n1719 vdd.n1718 585
R304 vdd.n1730 vdd.n1729 585
R305 vdd.n1728 vdd.n1727 585
R306 vdd.n1723 vdd.n1722 585
R307 vdd.n1806 vdd.n1805 585
R308 vdd.n1804 vdd.n1771 585
R309 vdd.n1803 vdd.n1802 585
R310 vdd.n1774 vdd.n1772 585
R311 vdd.n1797 vdd.n1796 585
R312 vdd.n1795 vdd.n1794 585
R313 vdd.n1778 vdd.n1777 585
R314 vdd.n1789 vdd.n1788 585
R315 vdd.n1787 vdd.n1786 585
R316 vdd.n1782 vdd.n1781 585
R317 vdd.n1645 vdd.n1644 585
R318 vdd.n1643 vdd.n1610 585
R319 vdd.n1642 vdd.n1641 585
R320 vdd.n1613 vdd.n1611 585
R321 vdd.n1636 vdd.n1635 585
R322 vdd.n1634 vdd.n1633 585
R323 vdd.n1617 vdd.n1616 585
R324 vdd.n1628 vdd.n1627 585
R325 vdd.n1626 vdd.n1625 585
R326 vdd.n1621 vdd.n1620 585
R327 vdd.n1704 vdd.n1703 585
R328 vdd.n1702 vdd.n1669 585
R329 vdd.n1701 vdd.n1700 585
R330 vdd.n1672 vdd.n1670 585
R331 vdd.n1695 vdd.n1694 585
R332 vdd.n1693 vdd.n1692 585
R333 vdd.n1676 vdd.n1675 585
R334 vdd.n1687 vdd.n1686 585
R335 vdd.n1685 vdd.n1684 585
R336 vdd.n1680 vdd.n1679 585
R337 vdd.n1544 vdd.n1543 585
R338 vdd.n1542 vdd.n1509 585
R339 vdd.n1541 vdd.n1540 585
R340 vdd.n1512 vdd.n1510 585
R341 vdd.n1535 vdd.n1534 585
R342 vdd.n1533 vdd.n1532 585
R343 vdd.n1516 vdd.n1515 585
R344 vdd.n1527 vdd.n1526 585
R345 vdd.n1525 vdd.n1524 585
R346 vdd.n1520 vdd.n1519 585
R347 vdd.n1603 vdd.n1602 585
R348 vdd.n1601 vdd.n1568 585
R349 vdd.n1600 vdd.n1599 585
R350 vdd.n1571 vdd.n1569 585
R351 vdd.n1594 vdd.n1593 585
R352 vdd.n1592 vdd.n1591 585
R353 vdd.n1575 vdd.n1574 585
R354 vdd.n1586 vdd.n1585 585
R355 vdd.n1584 vdd.n1583 585
R356 vdd.n1579 vdd.n1578 585
R357 vdd.n3356 vdd.n392 509.269
R358 vdd.n3352 vdd.n393 509.269
R359 vdd.n3224 vdd.n685 509.269
R360 vdd.n3221 vdd.n684 509.269
R361 vdd.n2328 vdd.n1075 509.269
R362 vdd.n2331 vdd.n2330 509.269
R363 vdd.n1224 vdd.n1188 509.269
R364 vdd.n1420 vdd.n1189 509.269
R365 vdd.n305 vdd.t104 329.043
R366 vdd.n246 vdd.t23 329.043
R367 vdd.n203 vdd.t107 329.043
R368 vdd.n144 vdd.t46 329.043
R369 vdd.n102 vdd.t118 329.043
R370 vdd.n43 vdd.t35 329.043
R371 vdd.n1724 vdd.t291 329.043
R372 vdd.n1783 vdd.t66 329.043
R373 vdd.n1622 vdd.t282 329.043
R374 vdd.n1681 vdd.t63 329.043
R375 vdd.n1521 vdd.t62 329.043
R376 vdd.n1580 vdd.t53 329.043
R377 vdd.n1317 vdd.t172 319.788
R378 vdd.n1355 vdd.t162 319.788
R379 vdd.n1251 vdd.t175 319.788
R380 vdd.n2333 vdd.t153 319.788
R381 vdd.n1970 vdd.t164 319.788
R382 vdd.n1930 vdd.t177 319.788
R383 vdd.n426 vdd.t168 319.788
R384 vdd.n440 vdd.t209 319.788
R385 vdd.n452 vdd.t215 319.788
R386 vdd.n768 vdd.t147 319.788
R387 vdd.n3184 vdd.t150 319.788
R388 vdd.n688 vdd.t213 319.788
R389 vdd.n1318 vdd.t171 303.69
R390 vdd.n1356 vdd.t161 303.69
R391 vdd.n1252 vdd.t174 303.69
R392 vdd.n2334 vdd.t154 303.69
R393 vdd.n1971 vdd.t165 303.69
R394 vdd.n1931 vdd.t178 303.69
R395 vdd.n427 vdd.t169 303.69
R396 vdd.n441 vdd.t210 303.69
R397 vdd.n453 vdd.t216 303.69
R398 vdd.n769 vdd.t146 303.69
R399 vdd.n3185 vdd.t149 303.69
R400 vdd.n689 vdd.t212 303.69
R401 vdd.n2865 vdd.n913 297.074
R402 vdd.n3058 vdd.n809 297.074
R403 vdd.n2995 vdd.n806 297.074
R404 vdd.n2788 vdd.n914 297.074
R405 vdd.n2603 vdd.n954 297.074
R406 vdd.n2534 vdd.n2533 297.074
R407 vdd.n2280 vdd.n1050 297.074
R408 vdd.n2376 vdd.n1048 297.074
R409 vdd.n2974 vdd.n807 297.074
R410 vdd.n3061 vdd.n3060 297.074
R411 vdd.n2637 vdd.n915 297.074
R412 vdd.n2863 vdd.n916 297.074
R413 vdd.n2531 vdd.n963 297.074
R414 vdd.n961 vdd.n936 297.074
R415 vdd.n2217 vdd.n1051 297.074
R416 vdd.n2374 vdd.n1052 297.074
R417 vdd.n2976 vdd.n807 185
R418 vdd.n3059 vdd.n807 185
R419 vdd.n2978 vdd.n2977 185
R420 vdd.n2977 vdd.n805 185
R421 vdd.n2979 vdd.n839 185
R422 vdd.n2989 vdd.n839 185
R423 vdd.n2980 vdd.n848 185
R424 vdd.n848 vdd.n846 185
R425 vdd.n2982 vdd.n2981 185
R426 vdd.n2983 vdd.n2982 185
R427 vdd.n2935 vdd.n847 185
R428 vdd.n847 vdd.n843 185
R429 vdd.n2934 vdd.n2933 185
R430 vdd.n2933 vdd.n2932 185
R431 vdd.n850 vdd.n849 185
R432 vdd.n851 vdd.n850 185
R433 vdd.n2925 vdd.n2924 185
R434 vdd.n2926 vdd.n2925 185
R435 vdd.n2921 vdd.n860 185
R436 vdd.n860 vdd.n857 185
R437 vdd.n2920 vdd.n2919 185
R438 vdd.n2919 vdd.n2918 185
R439 vdd.n862 vdd.n861 185
R440 vdd.n870 vdd.n862 185
R441 vdd.n2911 vdd.n2910 185
R442 vdd.n2912 vdd.n2911 185
R443 vdd.n2909 vdd.n871 185
R444 vdd.n2760 vdd.n871 185
R445 vdd.n2908 vdd.n2907 185
R446 vdd.n2907 vdd.n2906 185
R447 vdd.n873 vdd.n872 185
R448 vdd.n874 vdd.n873 185
R449 vdd.n2899 vdd.n2898 185
R450 vdd.n2900 vdd.n2899 185
R451 vdd.n2897 vdd.n883 185
R452 vdd.n883 vdd.n880 185
R453 vdd.n2896 vdd.n2895 185
R454 vdd.n2895 vdd.n2894 185
R455 vdd.n885 vdd.n884 185
R456 vdd.n893 vdd.n885 185
R457 vdd.n2887 vdd.n2886 185
R458 vdd.n2888 vdd.n2887 185
R459 vdd.n2885 vdd.n894 185
R460 vdd.n900 vdd.n894 185
R461 vdd.n2884 vdd.n2883 185
R462 vdd.n2883 vdd.n2882 185
R463 vdd.n896 vdd.n895 185
R464 vdd.n897 vdd.n896 185
R465 vdd.n2875 vdd.n2874 185
R466 vdd.n2876 vdd.n2875 185
R467 vdd.n2873 vdd.n906 185
R468 vdd.n2781 vdd.n906 185
R469 vdd.n2872 vdd.n2871 185
R470 vdd.n2871 vdd.n2870 185
R471 vdd.n908 vdd.n907 185
R472 vdd.t235 vdd.n908 185
R473 vdd.n2863 vdd.n2862 185
R474 vdd.n2864 vdd.n2863 185
R475 vdd.n2861 vdd.n916 185
R476 vdd.n2860 vdd.n2859 185
R477 vdd.n918 vdd.n917 185
R478 vdd.n2646 vdd.n2645 185
R479 vdd.n2648 vdd.n2647 185
R480 vdd.n2650 vdd.n2649 185
R481 vdd.n2652 vdd.n2651 185
R482 vdd.n2654 vdd.n2653 185
R483 vdd.n2656 vdd.n2655 185
R484 vdd.n2658 vdd.n2657 185
R485 vdd.n2660 vdd.n2659 185
R486 vdd.n2662 vdd.n2661 185
R487 vdd.n2664 vdd.n2663 185
R488 vdd.n2666 vdd.n2665 185
R489 vdd.n2668 vdd.n2667 185
R490 vdd.n2670 vdd.n2669 185
R491 vdd.n2672 vdd.n2671 185
R492 vdd.n2674 vdd.n2673 185
R493 vdd.n2676 vdd.n2675 185
R494 vdd.n2678 vdd.n2677 185
R495 vdd.n2680 vdd.n2679 185
R496 vdd.n2682 vdd.n2681 185
R497 vdd.n2684 vdd.n2683 185
R498 vdd.n2686 vdd.n2685 185
R499 vdd.n2688 vdd.n2687 185
R500 vdd.n2690 vdd.n2689 185
R501 vdd.n2692 vdd.n2691 185
R502 vdd.n2694 vdd.n2693 185
R503 vdd.n2696 vdd.n2695 185
R504 vdd.n2698 vdd.n2697 185
R505 vdd.n2700 vdd.n2699 185
R506 vdd.n2702 vdd.n2701 185
R507 vdd.n2704 vdd.n2703 185
R508 vdd.n2706 vdd.n2705 185
R509 vdd.n2707 vdd.n2637 185
R510 vdd.n2857 vdd.n2637 185
R511 vdd.n3062 vdd.n3061 185
R512 vdd.n3063 vdd.n798 185
R513 vdd.n3065 vdd.n3064 185
R514 vdd.n3067 vdd.n796 185
R515 vdd.n3069 vdd.n3068 185
R516 vdd.n3070 vdd.n795 185
R517 vdd.n3072 vdd.n3071 185
R518 vdd.n3074 vdd.n793 185
R519 vdd.n3076 vdd.n3075 185
R520 vdd.n3077 vdd.n792 185
R521 vdd.n3079 vdd.n3078 185
R522 vdd.n3081 vdd.n790 185
R523 vdd.n3083 vdd.n3082 185
R524 vdd.n3084 vdd.n789 185
R525 vdd.n3086 vdd.n3085 185
R526 vdd.n3088 vdd.n788 185
R527 vdd.n3089 vdd.n786 185
R528 vdd.n3092 vdd.n3091 185
R529 vdd.n787 vdd.n785 185
R530 vdd.n2948 vdd.n2947 185
R531 vdd.n2950 vdd.n2949 185
R532 vdd.n2952 vdd.n2944 185
R533 vdd.n2954 vdd.n2953 185
R534 vdd.n2955 vdd.n2943 185
R535 vdd.n2957 vdd.n2956 185
R536 vdd.n2959 vdd.n2941 185
R537 vdd.n2961 vdd.n2960 185
R538 vdd.n2962 vdd.n2940 185
R539 vdd.n2964 vdd.n2963 185
R540 vdd.n2966 vdd.n2938 185
R541 vdd.n2968 vdd.n2967 185
R542 vdd.n2969 vdd.n2937 185
R543 vdd.n2971 vdd.n2970 185
R544 vdd.n2973 vdd.n2936 185
R545 vdd.n2975 vdd.n2974 185
R546 vdd.n2974 vdd.n692 185
R547 vdd.n3060 vdd.n802 185
R548 vdd.n3060 vdd.n3059 185
R549 vdd.n2712 vdd.n804 185
R550 vdd.n805 vdd.n804 185
R551 vdd.n2713 vdd.n838 185
R552 vdd.n2989 vdd.n838 185
R553 vdd.n2715 vdd.n2714 185
R554 vdd.n2714 vdd.n846 185
R555 vdd.n2716 vdd.n845 185
R556 vdd.n2983 vdd.n845 185
R557 vdd.n2718 vdd.n2717 185
R558 vdd.n2717 vdd.n843 185
R559 vdd.n2719 vdd.n853 185
R560 vdd.n2932 vdd.n853 185
R561 vdd.n2721 vdd.n2720 185
R562 vdd.n2720 vdd.n851 185
R563 vdd.n2722 vdd.n859 185
R564 vdd.n2926 vdd.n859 185
R565 vdd.n2724 vdd.n2723 185
R566 vdd.n2723 vdd.n857 185
R567 vdd.n2725 vdd.n864 185
R568 vdd.n2918 vdd.n864 185
R569 vdd.n2727 vdd.n2726 185
R570 vdd.n2726 vdd.n870 185
R571 vdd.n2728 vdd.n869 185
R572 vdd.n2912 vdd.n869 185
R573 vdd.n2762 vdd.n2761 185
R574 vdd.n2761 vdd.n2760 185
R575 vdd.n2763 vdd.n876 185
R576 vdd.n2906 vdd.n876 185
R577 vdd.n2765 vdd.n2764 185
R578 vdd.n2764 vdd.n874 185
R579 vdd.n2766 vdd.n882 185
R580 vdd.n2900 vdd.n882 185
R581 vdd.n2768 vdd.n2767 185
R582 vdd.n2767 vdd.n880 185
R583 vdd.n2769 vdd.n887 185
R584 vdd.n2894 vdd.n887 185
R585 vdd.n2771 vdd.n2770 185
R586 vdd.n2770 vdd.n893 185
R587 vdd.n2772 vdd.n892 185
R588 vdd.n2888 vdd.n892 185
R589 vdd.n2774 vdd.n2773 185
R590 vdd.n2773 vdd.n900 185
R591 vdd.n2775 vdd.n899 185
R592 vdd.n2882 vdd.n899 185
R593 vdd.n2777 vdd.n2776 185
R594 vdd.n2776 vdd.n897 185
R595 vdd.n2778 vdd.n905 185
R596 vdd.n2876 vdd.n905 185
R597 vdd.n2780 vdd.n2779 185
R598 vdd.n2781 vdd.n2780 185
R599 vdd.n2711 vdd.n910 185
R600 vdd.n2870 vdd.n910 185
R601 vdd.n2710 vdd.n2709 185
R602 vdd.n2709 vdd.t235 185
R603 vdd.n2708 vdd.n915 185
R604 vdd.n2864 vdd.n915 185
R605 vdd.n2328 vdd.n2327 185
R606 vdd.n2329 vdd.n2328 185
R607 vdd.n1076 vdd.n1074 185
R608 vdd.n1894 vdd.n1074 185
R609 vdd.n1897 vdd.n1896 185
R610 vdd.n1896 vdd.n1895 185
R611 vdd.n1079 vdd.n1078 185
R612 vdd.n1080 vdd.n1079 185
R613 vdd.n1883 vdd.n1882 185
R614 vdd.n1884 vdd.n1883 185
R615 vdd.n1088 vdd.n1087 185
R616 vdd.n1875 vdd.n1087 185
R617 vdd.n1878 vdd.n1877 185
R618 vdd.n1877 vdd.n1876 185
R619 vdd.n1091 vdd.n1090 185
R620 vdd.n1098 vdd.n1091 185
R621 vdd.n1866 vdd.n1865 185
R622 vdd.n1867 vdd.n1866 185
R623 vdd.n1100 vdd.n1099 185
R624 vdd.n1099 vdd.n1097 185
R625 vdd.n1861 vdd.n1860 185
R626 vdd.n1860 vdd.n1859 185
R627 vdd.n1103 vdd.n1102 185
R628 vdd.n1104 vdd.n1103 185
R629 vdd.n1850 vdd.n1849 185
R630 vdd.n1851 vdd.n1850 185
R631 vdd.n1111 vdd.n1110 185
R632 vdd.n1842 vdd.n1110 185
R633 vdd.n1845 vdd.n1844 185
R634 vdd.n1844 vdd.n1843 185
R635 vdd.n1114 vdd.n1113 185
R636 vdd.n1120 vdd.n1114 185
R637 vdd.n1833 vdd.n1832 185
R638 vdd.n1834 vdd.n1833 185
R639 vdd.n1122 vdd.n1121 185
R640 vdd.n1825 vdd.n1121 185
R641 vdd.n1828 vdd.n1827 185
R642 vdd.n1827 vdd.n1826 185
R643 vdd.n1125 vdd.n1124 185
R644 vdd.n1126 vdd.n1125 185
R645 vdd.n1816 vdd.n1815 185
R646 vdd.n1817 vdd.n1816 185
R647 vdd.n1134 vdd.n1133 185
R648 vdd.n1133 vdd.n1132 185
R649 vdd.n1504 vdd.n1503 185
R650 vdd.n1503 vdd.n1502 185
R651 vdd.n1137 vdd.n1136 185
R652 vdd.n1143 vdd.n1137 185
R653 vdd.n1493 vdd.n1492 185
R654 vdd.n1494 vdd.n1493 185
R655 vdd.n1145 vdd.n1144 185
R656 vdd.n1485 vdd.n1144 185
R657 vdd.n1488 vdd.n1487 185
R658 vdd.n1487 vdd.n1486 185
R659 vdd.n1148 vdd.n1147 185
R660 vdd.n1155 vdd.n1148 185
R661 vdd.n1476 vdd.n1475 185
R662 vdd.n1477 vdd.n1476 185
R663 vdd.n1157 vdd.n1156 185
R664 vdd.n1156 vdd.n1154 185
R665 vdd.n1471 vdd.n1470 185
R666 vdd.n1470 vdd.n1469 185
R667 vdd.n1160 vdd.n1159 185
R668 vdd.n1161 vdd.n1160 185
R669 vdd.n1460 vdd.n1459 185
R670 vdd.n1461 vdd.n1460 185
R671 vdd.n1168 vdd.n1167 185
R672 vdd.n1452 vdd.n1167 185
R673 vdd.n1455 vdd.n1454 185
R674 vdd.n1454 vdd.n1453 185
R675 vdd.n1171 vdd.n1170 185
R676 vdd.n1177 vdd.n1171 185
R677 vdd.n1443 vdd.n1442 185
R678 vdd.n1444 vdd.n1443 185
R679 vdd.n1179 vdd.n1178 185
R680 vdd.n1435 vdd.n1178 185
R681 vdd.n1438 vdd.n1437 185
R682 vdd.n1437 vdd.n1436 185
R683 vdd.n1182 vdd.n1181 185
R684 vdd.n1183 vdd.n1182 185
R685 vdd.n1426 vdd.n1425 185
R686 vdd.n1427 vdd.n1426 185
R687 vdd.n1190 vdd.n1189 185
R688 vdd.n1225 vdd.n1189 185
R689 vdd.n1421 vdd.n1420 185
R690 vdd.n1193 vdd.n1192 185
R691 vdd.n1417 vdd.n1416 185
R692 vdd.n1418 vdd.n1417 185
R693 vdd.n1227 vdd.n1226 185
R694 vdd.n1412 vdd.n1229 185
R695 vdd.n1411 vdd.n1230 185
R696 vdd.n1410 vdd.n1231 185
R697 vdd.n1233 vdd.n1232 185
R698 vdd.n1406 vdd.n1235 185
R699 vdd.n1405 vdd.n1236 185
R700 vdd.n1404 vdd.n1237 185
R701 vdd.n1239 vdd.n1238 185
R702 vdd.n1400 vdd.n1241 185
R703 vdd.n1399 vdd.n1242 185
R704 vdd.n1398 vdd.n1243 185
R705 vdd.n1245 vdd.n1244 185
R706 vdd.n1394 vdd.n1247 185
R707 vdd.n1393 vdd.n1248 185
R708 vdd.n1392 vdd.n1249 185
R709 vdd.n1253 vdd.n1250 185
R710 vdd.n1388 vdd.n1255 185
R711 vdd.n1387 vdd.n1256 185
R712 vdd.n1386 vdd.n1257 185
R713 vdd.n1259 vdd.n1258 185
R714 vdd.n1382 vdd.n1261 185
R715 vdd.n1381 vdd.n1262 185
R716 vdd.n1380 vdd.n1263 185
R717 vdd.n1265 vdd.n1264 185
R718 vdd.n1376 vdd.n1267 185
R719 vdd.n1375 vdd.n1268 185
R720 vdd.n1374 vdd.n1269 185
R721 vdd.n1271 vdd.n1270 185
R722 vdd.n1370 vdd.n1273 185
R723 vdd.n1369 vdd.n1274 185
R724 vdd.n1368 vdd.n1275 185
R725 vdd.n1277 vdd.n1276 185
R726 vdd.n1364 vdd.n1279 185
R727 vdd.n1363 vdd.n1280 185
R728 vdd.n1362 vdd.n1281 185
R729 vdd.n1283 vdd.n1282 185
R730 vdd.n1358 vdd.n1285 185
R731 vdd.n1357 vdd.n1354 185
R732 vdd.n1353 vdd.n1286 185
R733 vdd.n1288 vdd.n1287 185
R734 vdd.n1349 vdd.n1290 185
R735 vdd.n1348 vdd.n1291 185
R736 vdd.n1347 vdd.n1292 185
R737 vdd.n1294 vdd.n1293 185
R738 vdd.n1343 vdd.n1296 185
R739 vdd.n1342 vdd.n1297 185
R740 vdd.n1341 vdd.n1298 185
R741 vdd.n1300 vdd.n1299 185
R742 vdd.n1337 vdd.n1302 185
R743 vdd.n1336 vdd.n1303 185
R744 vdd.n1335 vdd.n1304 185
R745 vdd.n1306 vdd.n1305 185
R746 vdd.n1331 vdd.n1308 185
R747 vdd.n1330 vdd.n1309 185
R748 vdd.n1329 vdd.n1310 185
R749 vdd.n1312 vdd.n1311 185
R750 vdd.n1325 vdd.n1314 185
R751 vdd.n1324 vdd.n1315 185
R752 vdd.n1323 vdd.n1316 185
R753 vdd.n1320 vdd.n1224 185
R754 vdd.n1418 vdd.n1224 185
R755 vdd.n2332 vdd.n2331 185
R756 vdd.n2336 vdd.n1069 185
R757 vdd.n1999 vdd.n1068 185
R758 vdd.n2002 vdd.n2001 185
R759 vdd.n2004 vdd.n2003 185
R760 vdd.n2007 vdd.n2006 185
R761 vdd.n2009 vdd.n2008 185
R762 vdd.n2011 vdd.n1997 185
R763 vdd.n2013 vdd.n2012 185
R764 vdd.n2014 vdd.n1991 185
R765 vdd.n2016 vdd.n2015 185
R766 vdd.n2018 vdd.n1989 185
R767 vdd.n2020 vdd.n2019 185
R768 vdd.n2021 vdd.n1984 185
R769 vdd.n2023 vdd.n2022 185
R770 vdd.n2025 vdd.n1982 185
R771 vdd.n2027 vdd.n2026 185
R772 vdd.n2028 vdd.n1978 185
R773 vdd.n2030 vdd.n2029 185
R774 vdd.n2032 vdd.n1975 185
R775 vdd.n2034 vdd.n2033 185
R776 vdd.n1976 vdd.n1969 185
R777 vdd.n2038 vdd.n1973 185
R778 vdd.n2039 vdd.n1965 185
R779 vdd.n2041 vdd.n2040 185
R780 vdd.n2043 vdd.n1963 185
R781 vdd.n2045 vdd.n2044 185
R782 vdd.n2046 vdd.n1958 185
R783 vdd.n2048 vdd.n2047 185
R784 vdd.n2050 vdd.n1956 185
R785 vdd.n2052 vdd.n2051 185
R786 vdd.n2053 vdd.n1951 185
R787 vdd.n2055 vdd.n2054 185
R788 vdd.n2057 vdd.n1949 185
R789 vdd.n2059 vdd.n2058 185
R790 vdd.n2060 vdd.n1944 185
R791 vdd.n2062 vdd.n2061 185
R792 vdd.n2064 vdd.n1942 185
R793 vdd.n2066 vdd.n2065 185
R794 vdd.n2067 vdd.n1938 185
R795 vdd.n2069 vdd.n2068 185
R796 vdd.n2071 vdd.n1935 185
R797 vdd.n2073 vdd.n2072 185
R798 vdd.n1936 vdd.n1929 185
R799 vdd.n2077 vdd.n1933 185
R800 vdd.n2078 vdd.n1925 185
R801 vdd.n2080 vdd.n2079 185
R802 vdd.n2082 vdd.n1923 185
R803 vdd.n2084 vdd.n2083 185
R804 vdd.n2085 vdd.n1918 185
R805 vdd.n2087 vdd.n2086 185
R806 vdd.n2089 vdd.n1916 185
R807 vdd.n2091 vdd.n2090 185
R808 vdd.n2092 vdd.n1911 185
R809 vdd.n2094 vdd.n2093 185
R810 vdd.n2096 vdd.n1910 185
R811 vdd.n2097 vdd.n1907 185
R812 vdd.n2100 vdd.n2099 185
R813 vdd.n1909 vdd.n1905 185
R814 vdd.n2317 vdd.n1903 185
R815 vdd.n2319 vdd.n2318 185
R816 vdd.n2321 vdd.n1901 185
R817 vdd.n2323 vdd.n2322 185
R818 vdd.n2324 vdd.n1075 185
R819 vdd.n2330 vdd.n1072 185
R820 vdd.n2330 vdd.n2329 185
R821 vdd.n1083 vdd.n1071 185
R822 vdd.n1894 vdd.n1071 185
R823 vdd.n1893 vdd.n1892 185
R824 vdd.n1895 vdd.n1893 185
R825 vdd.n1082 vdd.n1081 185
R826 vdd.n1081 vdd.n1080 185
R827 vdd.n1886 vdd.n1885 185
R828 vdd.n1885 vdd.n1884 185
R829 vdd.n1086 vdd.n1085 185
R830 vdd.n1875 vdd.n1086 185
R831 vdd.n1874 vdd.n1873 185
R832 vdd.n1876 vdd.n1874 185
R833 vdd.n1093 vdd.n1092 185
R834 vdd.n1098 vdd.n1092 185
R835 vdd.n1869 vdd.n1868 185
R836 vdd.n1868 vdd.n1867 185
R837 vdd.n1096 vdd.n1095 185
R838 vdd.n1097 vdd.n1096 185
R839 vdd.n1858 vdd.n1857 185
R840 vdd.n1859 vdd.n1858 185
R841 vdd.n1106 vdd.n1105 185
R842 vdd.n1105 vdd.n1104 185
R843 vdd.n1853 vdd.n1852 185
R844 vdd.n1852 vdd.n1851 185
R845 vdd.n1109 vdd.n1108 185
R846 vdd.n1842 vdd.n1109 185
R847 vdd.n1841 vdd.n1840 185
R848 vdd.n1843 vdd.n1841 185
R849 vdd.n1116 vdd.n1115 185
R850 vdd.n1120 vdd.n1115 185
R851 vdd.n1836 vdd.n1835 185
R852 vdd.n1835 vdd.n1834 185
R853 vdd.n1119 vdd.n1118 185
R854 vdd.n1825 vdd.n1119 185
R855 vdd.n1824 vdd.n1823 185
R856 vdd.n1826 vdd.n1824 185
R857 vdd.n1128 vdd.n1127 185
R858 vdd.n1127 vdd.n1126 185
R859 vdd.n1819 vdd.n1818 185
R860 vdd.n1818 vdd.n1817 185
R861 vdd.n1131 vdd.n1130 185
R862 vdd.n1132 vdd.n1131 185
R863 vdd.n1501 vdd.n1500 185
R864 vdd.n1502 vdd.n1501 185
R865 vdd.n1139 vdd.n1138 185
R866 vdd.n1143 vdd.n1138 185
R867 vdd.n1496 vdd.n1495 185
R868 vdd.n1495 vdd.n1494 185
R869 vdd.n1142 vdd.n1141 185
R870 vdd.n1485 vdd.n1142 185
R871 vdd.n1484 vdd.n1483 185
R872 vdd.n1486 vdd.n1484 185
R873 vdd.n1150 vdd.n1149 185
R874 vdd.n1155 vdd.n1149 185
R875 vdd.n1479 vdd.n1478 185
R876 vdd.n1478 vdd.n1477 185
R877 vdd.n1153 vdd.n1152 185
R878 vdd.n1154 vdd.n1153 185
R879 vdd.n1468 vdd.n1467 185
R880 vdd.n1469 vdd.n1468 185
R881 vdd.n1163 vdd.n1162 185
R882 vdd.n1162 vdd.n1161 185
R883 vdd.n1463 vdd.n1462 185
R884 vdd.n1462 vdd.n1461 185
R885 vdd.n1166 vdd.n1165 185
R886 vdd.n1452 vdd.n1166 185
R887 vdd.n1451 vdd.n1450 185
R888 vdd.n1453 vdd.n1451 185
R889 vdd.n1173 vdd.n1172 185
R890 vdd.n1177 vdd.n1172 185
R891 vdd.n1446 vdd.n1445 185
R892 vdd.n1445 vdd.n1444 185
R893 vdd.n1176 vdd.n1175 185
R894 vdd.n1435 vdd.n1176 185
R895 vdd.n1434 vdd.n1433 185
R896 vdd.n1436 vdd.n1434 185
R897 vdd.n1185 vdd.n1184 185
R898 vdd.n1184 vdd.n1183 185
R899 vdd.n1429 vdd.n1428 185
R900 vdd.n1428 vdd.n1427 185
R901 vdd.n1188 vdd.n1187 185
R902 vdd.n1225 vdd.n1188 185
R903 vdd.n956 vdd.n954 185
R904 vdd.n2532 vdd.n954 185
R905 vdd.n2454 vdd.n973 185
R906 vdd.n973 vdd.t268 185
R907 vdd.n2456 vdd.n2455 185
R908 vdd.n2457 vdd.n2456 185
R909 vdd.n2453 vdd.n972 185
R910 vdd.n2156 vdd.n972 185
R911 vdd.n2452 vdd.n2451 185
R912 vdd.n2451 vdd.n2450 185
R913 vdd.n975 vdd.n974 185
R914 vdd.n976 vdd.n975 185
R915 vdd.n2441 vdd.n2440 185
R916 vdd.n2442 vdd.n2441 185
R917 vdd.n2439 vdd.n986 185
R918 vdd.n986 vdd.n983 185
R919 vdd.n2438 vdd.n2437 185
R920 vdd.n2437 vdd.n2436 185
R921 vdd.n988 vdd.n987 185
R922 vdd.n989 vdd.n988 185
R923 vdd.n2429 vdd.n2428 185
R924 vdd.n2430 vdd.n2429 185
R925 vdd.n2427 vdd.n997 185
R926 vdd.n1002 vdd.n997 185
R927 vdd.n2426 vdd.n2425 185
R928 vdd.n2425 vdd.n2424 185
R929 vdd.n999 vdd.n998 185
R930 vdd.n1008 vdd.n999 185
R931 vdd.n2417 vdd.n2416 185
R932 vdd.n2418 vdd.n2417 185
R933 vdd.n2415 vdd.n1009 185
R934 vdd.n2257 vdd.n1009 185
R935 vdd.n2414 vdd.n2413 185
R936 vdd.n2413 vdd.n2412 185
R937 vdd.n1011 vdd.n1010 185
R938 vdd.n1012 vdd.n1011 185
R939 vdd.n2405 vdd.n2404 185
R940 vdd.n2406 vdd.n2405 185
R941 vdd.n2403 vdd.n1021 185
R942 vdd.n1021 vdd.n1018 185
R943 vdd.n2402 vdd.n2401 185
R944 vdd.n2401 vdd.n2400 185
R945 vdd.n1023 vdd.n1022 185
R946 vdd.n1033 vdd.n1023 185
R947 vdd.n2392 vdd.n2391 185
R948 vdd.n2393 vdd.n2392 185
R949 vdd.n2390 vdd.n1034 185
R950 vdd.n1034 vdd.n1030 185
R951 vdd.n2389 vdd.n2388 185
R952 vdd.n2388 vdd.n2387 185
R953 vdd.n1036 vdd.n1035 185
R954 vdd.n1037 vdd.n1036 185
R955 vdd.n2380 vdd.n2379 185
R956 vdd.n2381 vdd.n2380 185
R957 vdd.n2378 vdd.n1046 185
R958 vdd.n1046 vdd.n1043 185
R959 vdd.n2377 vdd.n2376 185
R960 vdd.n2376 vdd.n2375 185
R961 vdd.n1048 vdd.n1047 185
R962 vdd.n2112 vdd.n2111 185
R963 vdd.n2113 vdd.n2109 185
R964 vdd.n2109 vdd.n1049 185
R965 vdd.n2115 vdd.n2114 185
R966 vdd.n2117 vdd.n2108 185
R967 vdd.n2120 vdd.n2119 185
R968 vdd.n2121 vdd.n2107 185
R969 vdd.n2123 vdd.n2122 185
R970 vdd.n2125 vdd.n2106 185
R971 vdd.n2128 vdd.n2127 185
R972 vdd.n2129 vdd.n2105 185
R973 vdd.n2131 vdd.n2130 185
R974 vdd.n2133 vdd.n2104 185
R975 vdd.n2136 vdd.n2135 185
R976 vdd.n2137 vdd.n2103 185
R977 vdd.n2139 vdd.n2138 185
R978 vdd.n2141 vdd.n2102 185
R979 vdd.n2314 vdd.n2142 185
R980 vdd.n2313 vdd.n2312 185
R981 vdd.n2310 vdd.n2143 185
R982 vdd.n2308 vdd.n2307 185
R983 vdd.n2306 vdd.n2144 185
R984 vdd.n2305 vdd.n2304 185
R985 vdd.n2302 vdd.n2145 185
R986 vdd.n2300 vdd.n2299 185
R987 vdd.n2298 vdd.n2146 185
R988 vdd.n2297 vdd.n2296 185
R989 vdd.n2294 vdd.n2147 185
R990 vdd.n2292 vdd.n2291 185
R991 vdd.n2290 vdd.n2148 185
R992 vdd.n2289 vdd.n2288 185
R993 vdd.n2286 vdd.n2149 185
R994 vdd.n2284 vdd.n2283 185
R995 vdd.n2282 vdd.n2150 185
R996 vdd.n2281 vdd.n2280 185
R997 vdd.n2535 vdd.n2534 185
R998 vdd.n2537 vdd.n2536 185
R999 vdd.n2539 vdd.n2538 185
R1000 vdd.n2542 vdd.n2541 185
R1001 vdd.n2544 vdd.n2543 185
R1002 vdd.n2546 vdd.n2545 185
R1003 vdd.n2548 vdd.n2547 185
R1004 vdd.n2550 vdd.n2549 185
R1005 vdd.n2552 vdd.n2551 185
R1006 vdd.n2554 vdd.n2553 185
R1007 vdd.n2556 vdd.n2555 185
R1008 vdd.n2558 vdd.n2557 185
R1009 vdd.n2560 vdd.n2559 185
R1010 vdd.n2562 vdd.n2561 185
R1011 vdd.n2564 vdd.n2563 185
R1012 vdd.n2566 vdd.n2565 185
R1013 vdd.n2568 vdd.n2567 185
R1014 vdd.n2570 vdd.n2569 185
R1015 vdd.n2572 vdd.n2571 185
R1016 vdd.n2574 vdd.n2573 185
R1017 vdd.n2576 vdd.n2575 185
R1018 vdd.n2578 vdd.n2577 185
R1019 vdd.n2580 vdd.n2579 185
R1020 vdd.n2582 vdd.n2581 185
R1021 vdd.n2584 vdd.n2583 185
R1022 vdd.n2586 vdd.n2585 185
R1023 vdd.n2588 vdd.n2587 185
R1024 vdd.n2590 vdd.n2589 185
R1025 vdd.n2592 vdd.n2591 185
R1026 vdd.n2594 vdd.n2593 185
R1027 vdd.n2596 vdd.n2595 185
R1028 vdd.n2598 vdd.n2597 185
R1029 vdd.n2600 vdd.n2599 185
R1030 vdd.n2601 vdd.n955 185
R1031 vdd.n2603 vdd.n2602 185
R1032 vdd.n2604 vdd.n2603 185
R1033 vdd.n2533 vdd.n959 185
R1034 vdd.n2533 vdd.n2532 185
R1035 vdd.n2154 vdd.n960 185
R1036 vdd.t268 vdd.n960 185
R1037 vdd.n2155 vdd.n970 185
R1038 vdd.n2457 vdd.n970 185
R1039 vdd.n2158 vdd.n2157 185
R1040 vdd.n2157 vdd.n2156 185
R1041 vdd.n2159 vdd.n977 185
R1042 vdd.n2450 vdd.n977 185
R1043 vdd.n2161 vdd.n2160 185
R1044 vdd.n2160 vdd.n976 185
R1045 vdd.n2162 vdd.n984 185
R1046 vdd.n2442 vdd.n984 185
R1047 vdd.n2164 vdd.n2163 185
R1048 vdd.n2163 vdd.n983 185
R1049 vdd.n2165 vdd.n990 185
R1050 vdd.n2436 vdd.n990 185
R1051 vdd.n2167 vdd.n2166 185
R1052 vdd.n2166 vdd.n989 185
R1053 vdd.n2168 vdd.n995 185
R1054 vdd.n2430 vdd.n995 185
R1055 vdd.n2170 vdd.n2169 185
R1056 vdd.n2169 vdd.n1002 185
R1057 vdd.n2171 vdd.n1000 185
R1058 vdd.n2424 vdd.n1000 185
R1059 vdd.n2173 vdd.n2172 185
R1060 vdd.n2172 vdd.n1008 185
R1061 vdd.n2174 vdd.n1006 185
R1062 vdd.n2418 vdd.n1006 185
R1063 vdd.n2259 vdd.n2258 185
R1064 vdd.n2258 vdd.n2257 185
R1065 vdd.n2260 vdd.n1013 185
R1066 vdd.n2412 vdd.n1013 185
R1067 vdd.n2262 vdd.n2261 185
R1068 vdd.n2261 vdd.n1012 185
R1069 vdd.n2263 vdd.n1019 185
R1070 vdd.n2406 vdd.n1019 185
R1071 vdd.n2265 vdd.n2264 185
R1072 vdd.n2264 vdd.n1018 185
R1073 vdd.n2266 vdd.n1024 185
R1074 vdd.n2400 vdd.n1024 185
R1075 vdd.n2268 vdd.n2267 185
R1076 vdd.n2267 vdd.n1033 185
R1077 vdd.n2269 vdd.n1031 185
R1078 vdd.n2393 vdd.n1031 185
R1079 vdd.n2271 vdd.n2270 185
R1080 vdd.n2270 vdd.n1030 185
R1081 vdd.n2272 vdd.n1038 185
R1082 vdd.n2387 vdd.n1038 185
R1083 vdd.n2274 vdd.n2273 185
R1084 vdd.n2273 vdd.n1037 185
R1085 vdd.n2275 vdd.n1044 185
R1086 vdd.n2381 vdd.n1044 185
R1087 vdd.n2277 vdd.n2276 185
R1088 vdd.n2276 vdd.n1043 185
R1089 vdd.n2278 vdd.n1050 185
R1090 vdd.n2375 vdd.n1050 185
R1091 vdd.n3357 vdd.n3356 185
R1092 vdd.n3356 vdd.n3355 185
R1093 vdd.n3358 vdd.n387 185
R1094 vdd.n387 vdd.n386 185
R1095 vdd.n3360 vdd.n3359 185
R1096 vdd.n3361 vdd.n3360 185
R1097 vdd.n382 vdd.n381 185
R1098 vdd.n3362 vdd.n382 185
R1099 vdd.n3365 vdd.n3364 185
R1100 vdd.n3364 vdd.n3363 185
R1101 vdd.n3366 vdd.n376 185
R1102 vdd.n376 vdd.n375 185
R1103 vdd.n3368 vdd.n3367 185
R1104 vdd.n3369 vdd.n3368 185
R1105 vdd.n371 vdd.n370 185
R1106 vdd.n3370 vdd.n371 185
R1107 vdd.n3373 vdd.n3372 185
R1108 vdd.n3372 vdd.n3371 185
R1109 vdd.n3374 vdd.n365 185
R1110 vdd.n3331 vdd.n365 185
R1111 vdd.n3376 vdd.n3375 185
R1112 vdd.n3377 vdd.n3376 185
R1113 vdd.n360 vdd.n359 185
R1114 vdd.n3378 vdd.n360 185
R1115 vdd.n3381 vdd.n3380 185
R1116 vdd.n3380 vdd.n3379 185
R1117 vdd.n3382 vdd.n354 185
R1118 vdd.n361 vdd.n354 185
R1119 vdd.n3384 vdd.n3383 185
R1120 vdd.n3385 vdd.n3384 185
R1121 vdd.n350 vdd.n349 185
R1122 vdd.n3386 vdd.n350 185
R1123 vdd.n3389 vdd.n3388 185
R1124 vdd.n3388 vdd.n3387 185
R1125 vdd.n3390 vdd.n345 185
R1126 vdd.n345 vdd.n344 185
R1127 vdd.n3392 vdd.n3391 185
R1128 vdd.n3393 vdd.n3392 185
R1129 vdd.n339 vdd.n337 185
R1130 vdd.n3394 vdd.n339 185
R1131 vdd.n3397 vdd.n3396 185
R1132 vdd.n3396 vdd.n3395 185
R1133 vdd.n338 vdd.n336 185
R1134 vdd.n340 vdd.n338 185
R1135 vdd.n3307 vdd.n3306 185
R1136 vdd.n3308 vdd.n3307 185
R1137 vdd.n635 vdd.n634 185
R1138 vdd.n634 vdd.n633 185
R1139 vdd.n3302 vdd.n3301 185
R1140 vdd.n3301 vdd.n3300 185
R1141 vdd.n638 vdd.n637 185
R1142 vdd.n644 vdd.n638 185
R1143 vdd.n3288 vdd.n3287 185
R1144 vdd.n3289 vdd.n3288 185
R1145 vdd.n646 vdd.n645 185
R1146 vdd.n3280 vdd.n645 185
R1147 vdd.n3283 vdd.n3282 185
R1148 vdd.n3282 vdd.n3281 185
R1149 vdd.n649 vdd.n648 185
R1150 vdd.n656 vdd.n649 185
R1151 vdd.n3271 vdd.n3270 185
R1152 vdd.n3272 vdd.n3271 185
R1153 vdd.n658 vdd.n657 185
R1154 vdd.n657 vdd.n655 185
R1155 vdd.n3266 vdd.n3265 185
R1156 vdd.n3265 vdd.n3264 185
R1157 vdd.n661 vdd.n660 185
R1158 vdd.n662 vdd.n661 185
R1159 vdd.n3255 vdd.n3254 185
R1160 vdd.n3256 vdd.n3255 185
R1161 vdd.n669 vdd.n668 185
R1162 vdd.n3247 vdd.n668 185
R1163 vdd.n3250 vdd.n3249 185
R1164 vdd.n3249 vdd.n3248 185
R1165 vdd.n672 vdd.n671 185
R1166 vdd.n679 vdd.n672 185
R1167 vdd.n3238 vdd.n3237 185
R1168 vdd.n3239 vdd.n3238 185
R1169 vdd.n681 vdd.n680 185
R1170 vdd.n680 vdd.n678 185
R1171 vdd.n3233 vdd.n3232 185
R1172 vdd.n3232 vdd.n3231 185
R1173 vdd.n684 vdd.n683 185
R1174 vdd.n723 vdd.n684 185
R1175 vdd.n3221 vdd.n3220 185
R1176 vdd.n3219 vdd.n725 185
R1177 vdd.n3218 vdd.n724 185
R1178 vdd.n3223 vdd.n724 185
R1179 vdd.n729 vdd.n728 185
R1180 vdd.n733 vdd.n732 185
R1181 vdd.n3214 vdd.n734 185
R1182 vdd.n3213 vdd.n3212 185
R1183 vdd.n3211 vdd.n3210 185
R1184 vdd.n3209 vdd.n3208 185
R1185 vdd.n3207 vdd.n3206 185
R1186 vdd.n3205 vdd.n3204 185
R1187 vdd.n3203 vdd.n3202 185
R1188 vdd.n3201 vdd.n3200 185
R1189 vdd.n3199 vdd.n3198 185
R1190 vdd.n3197 vdd.n3196 185
R1191 vdd.n3195 vdd.n3194 185
R1192 vdd.n3193 vdd.n3192 185
R1193 vdd.n3191 vdd.n3190 185
R1194 vdd.n3189 vdd.n3188 185
R1195 vdd.n3187 vdd.n3186 185
R1196 vdd.n3178 vdd.n747 185
R1197 vdd.n3180 vdd.n3179 185
R1198 vdd.n3177 vdd.n3176 185
R1199 vdd.n3175 vdd.n3174 185
R1200 vdd.n3173 vdd.n3172 185
R1201 vdd.n3171 vdd.n3170 185
R1202 vdd.n3169 vdd.n3168 185
R1203 vdd.n3167 vdd.n3166 185
R1204 vdd.n3165 vdd.n3164 185
R1205 vdd.n3163 vdd.n3162 185
R1206 vdd.n3161 vdd.n3160 185
R1207 vdd.n3159 vdd.n3158 185
R1208 vdd.n3157 vdd.n3156 185
R1209 vdd.n3155 vdd.n3154 185
R1210 vdd.n3153 vdd.n3152 185
R1211 vdd.n3151 vdd.n3150 185
R1212 vdd.n3149 vdd.n3148 185
R1213 vdd.n3147 vdd.n3146 185
R1214 vdd.n3145 vdd.n3144 185
R1215 vdd.n3143 vdd.n3142 185
R1216 vdd.n3141 vdd.n3140 185
R1217 vdd.n3139 vdd.n3138 185
R1218 vdd.n3132 vdd.n767 185
R1219 vdd.n3134 vdd.n3133 185
R1220 vdd.n3131 vdd.n3130 185
R1221 vdd.n3129 vdd.n3128 185
R1222 vdd.n3127 vdd.n3126 185
R1223 vdd.n3125 vdd.n3124 185
R1224 vdd.n3123 vdd.n3122 185
R1225 vdd.n3121 vdd.n3120 185
R1226 vdd.n3119 vdd.n3118 185
R1227 vdd.n3117 vdd.n3116 185
R1228 vdd.n3115 vdd.n3114 185
R1229 vdd.n3113 vdd.n3112 185
R1230 vdd.n3111 vdd.n3110 185
R1231 vdd.n3109 vdd.n3108 185
R1232 vdd.n3107 vdd.n3106 185
R1233 vdd.n3105 vdd.n3104 185
R1234 vdd.n3103 vdd.n3102 185
R1235 vdd.n3101 vdd.n3100 185
R1236 vdd.n3099 vdd.n3098 185
R1237 vdd.n3097 vdd.n3096 185
R1238 vdd.n3095 vdd.n691 185
R1239 vdd.n3225 vdd.n3224 185
R1240 vdd.n3224 vdd.n3223 185
R1241 vdd.n3352 vdd.n3351 185
R1242 vdd.n618 vdd.n425 185
R1243 vdd.n617 vdd.n616 185
R1244 vdd.n615 vdd.n614 185
R1245 vdd.n613 vdd.n430 185
R1246 vdd.n609 vdd.n608 185
R1247 vdd.n607 vdd.n606 185
R1248 vdd.n605 vdd.n604 185
R1249 vdd.n603 vdd.n432 185
R1250 vdd.n599 vdd.n598 185
R1251 vdd.n597 vdd.n596 185
R1252 vdd.n595 vdd.n594 185
R1253 vdd.n593 vdd.n434 185
R1254 vdd.n589 vdd.n588 185
R1255 vdd.n587 vdd.n586 185
R1256 vdd.n585 vdd.n584 185
R1257 vdd.n583 vdd.n436 185
R1258 vdd.n579 vdd.n578 185
R1259 vdd.n577 vdd.n576 185
R1260 vdd.n575 vdd.n574 185
R1261 vdd.n573 vdd.n438 185
R1262 vdd.n569 vdd.n568 185
R1263 vdd.n567 vdd.n566 185
R1264 vdd.n565 vdd.n564 185
R1265 vdd.n563 vdd.n442 185
R1266 vdd.n559 vdd.n558 185
R1267 vdd.n557 vdd.n556 185
R1268 vdd.n555 vdd.n554 185
R1269 vdd.n553 vdd.n444 185
R1270 vdd.n549 vdd.n548 185
R1271 vdd.n547 vdd.n546 185
R1272 vdd.n545 vdd.n544 185
R1273 vdd.n543 vdd.n446 185
R1274 vdd.n539 vdd.n538 185
R1275 vdd.n537 vdd.n536 185
R1276 vdd.n535 vdd.n534 185
R1277 vdd.n533 vdd.n448 185
R1278 vdd.n529 vdd.n528 185
R1279 vdd.n527 vdd.n526 185
R1280 vdd.n525 vdd.n524 185
R1281 vdd.n523 vdd.n450 185
R1282 vdd.n519 vdd.n518 185
R1283 vdd.n517 vdd.n516 185
R1284 vdd.n515 vdd.n514 185
R1285 vdd.n513 vdd.n454 185
R1286 vdd.n509 vdd.n508 185
R1287 vdd.n507 vdd.n506 185
R1288 vdd.n505 vdd.n504 185
R1289 vdd.n503 vdd.n456 185
R1290 vdd.n499 vdd.n498 185
R1291 vdd.n497 vdd.n496 185
R1292 vdd.n495 vdd.n494 185
R1293 vdd.n493 vdd.n458 185
R1294 vdd.n489 vdd.n488 185
R1295 vdd.n487 vdd.n486 185
R1296 vdd.n485 vdd.n484 185
R1297 vdd.n483 vdd.n460 185
R1298 vdd.n479 vdd.n478 185
R1299 vdd.n477 vdd.n476 185
R1300 vdd.n475 vdd.n474 185
R1301 vdd.n473 vdd.n462 185
R1302 vdd.n469 vdd.n468 185
R1303 vdd.n467 vdd.n466 185
R1304 vdd.n465 vdd.n392 185
R1305 vdd.n3348 vdd.n393 185
R1306 vdd.n3355 vdd.n393 185
R1307 vdd.n3347 vdd.n3346 185
R1308 vdd.n3346 vdd.n386 185
R1309 vdd.n3345 vdd.n385 185
R1310 vdd.n3361 vdd.n385 185
R1311 vdd.n621 vdd.n384 185
R1312 vdd.n3362 vdd.n384 185
R1313 vdd.n3341 vdd.n383 185
R1314 vdd.n3363 vdd.n383 185
R1315 vdd.n3340 vdd.n3339 185
R1316 vdd.n3339 vdd.n375 185
R1317 vdd.n3338 vdd.n374 185
R1318 vdd.n3369 vdd.n374 185
R1319 vdd.n623 vdd.n373 185
R1320 vdd.n3370 vdd.n373 185
R1321 vdd.n3334 vdd.n372 185
R1322 vdd.n3371 vdd.n372 185
R1323 vdd.n3333 vdd.n3332 185
R1324 vdd.n3332 vdd.n3331 185
R1325 vdd.n3330 vdd.n364 185
R1326 vdd.n3377 vdd.n364 185
R1327 vdd.n625 vdd.n363 185
R1328 vdd.n3378 vdd.n363 185
R1329 vdd.n3326 vdd.n362 185
R1330 vdd.n3379 vdd.n362 185
R1331 vdd.n3325 vdd.n3324 185
R1332 vdd.n3324 vdd.n361 185
R1333 vdd.n3323 vdd.n353 185
R1334 vdd.n3385 vdd.n353 185
R1335 vdd.n627 vdd.n352 185
R1336 vdd.n3386 vdd.n352 185
R1337 vdd.n3319 vdd.n351 185
R1338 vdd.n3387 vdd.n351 185
R1339 vdd.n3318 vdd.n3317 185
R1340 vdd.n3317 vdd.n344 185
R1341 vdd.n3316 vdd.n343 185
R1342 vdd.n3393 vdd.n343 185
R1343 vdd.n629 vdd.n342 185
R1344 vdd.n3394 vdd.n342 185
R1345 vdd.n3312 vdd.n341 185
R1346 vdd.n3395 vdd.n341 185
R1347 vdd.n3311 vdd.n3310 185
R1348 vdd.n3310 vdd.n340 185
R1349 vdd.n3309 vdd.n631 185
R1350 vdd.n3309 vdd.n3308 185
R1351 vdd.n3297 vdd.n632 185
R1352 vdd.n633 vdd.n632 185
R1353 vdd.n3299 vdd.n3298 185
R1354 vdd.n3300 vdd.n3299 185
R1355 vdd.n640 vdd.n639 185
R1356 vdd.n644 vdd.n639 185
R1357 vdd.n3291 vdd.n3290 185
R1358 vdd.n3290 vdd.n3289 185
R1359 vdd.n643 vdd.n642 185
R1360 vdd.n3280 vdd.n643 185
R1361 vdd.n3279 vdd.n3278 185
R1362 vdd.n3281 vdd.n3279 185
R1363 vdd.n651 vdd.n650 185
R1364 vdd.n656 vdd.n650 185
R1365 vdd.n3274 vdd.n3273 185
R1366 vdd.n3273 vdd.n3272 185
R1367 vdd.n654 vdd.n653 185
R1368 vdd.n655 vdd.n654 185
R1369 vdd.n3263 vdd.n3262 185
R1370 vdd.n3264 vdd.n3263 185
R1371 vdd.n664 vdd.n663 185
R1372 vdd.n663 vdd.n662 185
R1373 vdd.n3258 vdd.n3257 185
R1374 vdd.n3257 vdd.n3256 185
R1375 vdd.n667 vdd.n666 185
R1376 vdd.n3247 vdd.n667 185
R1377 vdd.n3246 vdd.n3245 185
R1378 vdd.n3248 vdd.n3246 185
R1379 vdd.n674 vdd.n673 185
R1380 vdd.n679 vdd.n673 185
R1381 vdd.n3241 vdd.n3240 185
R1382 vdd.n3240 vdd.n3239 185
R1383 vdd.n677 vdd.n676 185
R1384 vdd.n678 vdd.n677 185
R1385 vdd.n3230 vdd.n3229 185
R1386 vdd.n3231 vdd.n3230 185
R1387 vdd.n686 vdd.n685 185
R1388 vdd.n723 vdd.n685 185
R1389 vdd.n913 vdd.n912 185
R1390 vdd.n2855 vdd.n2854 185
R1391 vdd.n2853 vdd.n2638 185
R1392 vdd.n2857 vdd.n2638 185
R1393 vdd.n2852 vdd.n2851 185
R1394 vdd.n2850 vdd.n2849 185
R1395 vdd.n2848 vdd.n2847 185
R1396 vdd.n2846 vdd.n2845 185
R1397 vdd.n2844 vdd.n2843 185
R1398 vdd.n2842 vdd.n2841 185
R1399 vdd.n2840 vdd.n2839 185
R1400 vdd.n2838 vdd.n2837 185
R1401 vdd.n2836 vdd.n2835 185
R1402 vdd.n2834 vdd.n2833 185
R1403 vdd.n2832 vdd.n2831 185
R1404 vdd.n2830 vdd.n2829 185
R1405 vdd.n2828 vdd.n2827 185
R1406 vdd.n2826 vdd.n2825 185
R1407 vdd.n2824 vdd.n2823 185
R1408 vdd.n2822 vdd.n2821 185
R1409 vdd.n2820 vdd.n2819 185
R1410 vdd.n2818 vdd.n2817 185
R1411 vdd.n2816 vdd.n2815 185
R1412 vdd.n2814 vdd.n2813 185
R1413 vdd.n2812 vdd.n2811 185
R1414 vdd.n2810 vdd.n2809 185
R1415 vdd.n2808 vdd.n2807 185
R1416 vdd.n2806 vdd.n2805 185
R1417 vdd.n2804 vdd.n2803 185
R1418 vdd.n2802 vdd.n2801 185
R1419 vdd.n2800 vdd.n2799 185
R1420 vdd.n2798 vdd.n2797 185
R1421 vdd.n2796 vdd.n2795 185
R1422 vdd.n2793 vdd.n2792 185
R1423 vdd.n2791 vdd.n2790 185
R1424 vdd.n2789 vdd.n2788 185
R1425 vdd.n2995 vdd.n2994 185
R1426 vdd.n2997 vdd.n834 185
R1427 vdd.n2999 vdd.n2998 185
R1428 vdd.n3001 vdd.n831 185
R1429 vdd.n3003 vdd.n3002 185
R1430 vdd.n3005 vdd.n829 185
R1431 vdd.n3007 vdd.n3006 185
R1432 vdd.n3008 vdd.n828 185
R1433 vdd.n3010 vdd.n3009 185
R1434 vdd.n3012 vdd.n826 185
R1435 vdd.n3014 vdd.n3013 185
R1436 vdd.n3015 vdd.n825 185
R1437 vdd.n3017 vdd.n3016 185
R1438 vdd.n3019 vdd.n823 185
R1439 vdd.n3021 vdd.n3020 185
R1440 vdd.n3022 vdd.n822 185
R1441 vdd.n3024 vdd.n3023 185
R1442 vdd.n3026 vdd.n731 185
R1443 vdd.n3028 vdd.n3027 185
R1444 vdd.n3030 vdd.n820 185
R1445 vdd.n3032 vdd.n3031 185
R1446 vdd.n3033 vdd.n819 185
R1447 vdd.n3035 vdd.n3034 185
R1448 vdd.n3037 vdd.n817 185
R1449 vdd.n3039 vdd.n3038 185
R1450 vdd.n3040 vdd.n816 185
R1451 vdd.n3042 vdd.n3041 185
R1452 vdd.n3044 vdd.n814 185
R1453 vdd.n3046 vdd.n3045 185
R1454 vdd.n3047 vdd.n813 185
R1455 vdd.n3049 vdd.n3048 185
R1456 vdd.n3051 vdd.n812 185
R1457 vdd.n3052 vdd.n811 185
R1458 vdd.n3055 vdd.n3054 185
R1459 vdd.n3056 vdd.n809 185
R1460 vdd.n809 vdd.n692 185
R1461 vdd.n2993 vdd.n806 185
R1462 vdd.n3059 vdd.n806 185
R1463 vdd.n2992 vdd.n2991 185
R1464 vdd.n2991 vdd.n805 185
R1465 vdd.n2990 vdd.n836 185
R1466 vdd.n2990 vdd.n2989 185
R1467 vdd.n2744 vdd.n837 185
R1468 vdd.n846 vdd.n837 185
R1469 vdd.n2745 vdd.n844 185
R1470 vdd.n2983 vdd.n844 185
R1471 vdd.n2747 vdd.n2746 185
R1472 vdd.n2746 vdd.n843 185
R1473 vdd.n2748 vdd.n852 185
R1474 vdd.n2932 vdd.n852 185
R1475 vdd.n2750 vdd.n2749 185
R1476 vdd.n2749 vdd.n851 185
R1477 vdd.n2751 vdd.n858 185
R1478 vdd.n2926 vdd.n858 185
R1479 vdd.n2753 vdd.n2752 185
R1480 vdd.n2752 vdd.n857 185
R1481 vdd.n2754 vdd.n863 185
R1482 vdd.n2918 vdd.n863 185
R1483 vdd.n2756 vdd.n2755 185
R1484 vdd.n2755 vdd.n870 185
R1485 vdd.n2757 vdd.n868 185
R1486 vdd.n2912 vdd.n868 185
R1487 vdd.n2759 vdd.n2758 185
R1488 vdd.n2760 vdd.n2759 185
R1489 vdd.n2743 vdd.n875 185
R1490 vdd.n2906 vdd.n875 185
R1491 vdd.n2742 vdd.n2741 185
R1492 vdd.n2741 vdd.n874 185
R1493 vdd.n2740 vdd.n881 185
R1494 vdd.n2900 vdd.n881 185
R1495 vdd.n2739 vdd.n2738 185
R1496 vdd.n2738 vdd.n880 185
R1497 vdd.n2737 vdd.n886 185
R1498 vdd.n2894 vdd.n886 185
R1499 vdd.n2736 vdd.n2735 185
R1500 vdd.n2735 vdd.n893 185
R1501 vdd.n2734 vdd.n891 185
R1502 vdd.n2888 vdd.n891 185
R1503 vdd.n2733 vdd.n2732 185
R1504 vdd.n2732 vdd.n900 185
R1505 vdd.n2731 vdd.n898 185
R1506 vdd.n2882 vdd.n898 185
R1507 vdd.n2730 vdd.n2729 185
R1508 vdd.n2729 vdd.n897 185
R1509 vdd.n2641 vdd.n904 185
R1510 vdd.n2876 vdd.n904 185
R1511 vdd.n2783 vdd.n2782 185
R1512 vdd.n2782 vdd.n2781 185
R1513 vdd.n2784 vdd.n909 185
R1514 vdd.n2870 vdd.n909 185
R1515 vdd.n2786 vdd.n2785 185
R1516 vdd.n2785 vdd.t235 185
R1517 vdd.n2787 vdd.n914 185
R1518 vdd.n2864 vdd.n914 185
R1519 vdd.n2866 vdd.n2865 185
R1520 vdd.n2865 vdd.n2864 185
R1521 vdd.n2867 vdd.n911 185
R1522 vdd.n911 vdd.t235 185
R1523 vdd.n2869 vdd.n2868 185
R1524 vdd.n2870 vdd.n2869 185
R1525 vdd.n903 vdd.n902 185
R1526 vdd.n2781 vdd.n903 185
R1527 vdd.n2878 vdd.n2877 185
R1528 vdd.n2877 vdd.n2876 185
R1529 vdd.n2879 vdd.n901 185
R1530 vdd.n901 vdd.n897 185
R1531 vdd.n2881 vdd.n2880 185
R1532 vdd.n2882 vdd.n2881 185
R1533 vdd.n890 vdd.n889 185
R1534 vdd.n900 vdd.n890 185
R1535 vdd.n2890 vdd.n2889 185
R1536 vdd.n2889 vdd.n2888 185
R1537 vdd.n2891 vdd.n888 185
R1538 vdd.n893 vdd.n888 185
R1539 vdd.n2893 vdd.n2892 185
R1540 vdd.n2894 vdd.n2893 185
R1541 vdd.n879 vdd.n878 185
R1542 vdd.n880 vdd.n879 185
R1543 vdd.n2902 vdd.n2901 185
R1544 vdd.n2901 vdd.n2900 185
R1545 vdd.n2903 vdd.n877 185
R1546 vdd.n877 vdd.n874 185
R1547 vdd.n2905 vdd.n2904 185
R1548 vdd.n2906 vdd.n2905 185
R1549 vdd.n867 vdd.n866 185
R1550 vdd.n2760 vdd.n867 185
R1551 vdd.n2914 vdd.n2913 185
R1552 vdd.n2913 vdd.n2912 185
R1553 vdd.n2915 vdd.n865 185
R1554 vdd.n870 vdd.n865 185
R1555 vdd.n2917 vdd.n2916 185
R1556 vdd.n2918 vdd.n2917 185
R1557 vdd.n856 vdd.n855 185
R1558 vdd.n857 vdd.n856 185
R1559 vdd.n2928 vdd.n2927 185
R1560 vdd.n2927 vdd.n2926 185
R1561 vdd.n2929 vdd.n854 185
R1562 vdd.n854 vdd.n851 185
R1563 vdd.n2931 vdd.n2930 185
R1564 vdd.n2932 vdd.n2931 185
R1565 vdd.n842 vdd.n841 185
R1566 vdd.n843 vdd.n842 185
R1567 vdd.n2985 vdd.n2984 185
R1568 vdd.n2984 vdd.n2983 185
R1569 vdd.n2986 vdd.n840 185
R1570 vdd.n846 vdd.n840 185
R1571 vdd.n2988 vdd.n2987 185
R1572 vdd.n2989 vdd.n2988 185
R1573 vdd.n810 vdd.n808 185
R1574 vdd.n808 vdd.n805 185
R1575 vdd.n3058 vdd.n3057 185
R1576 vdd.n3059 vdd.n3058 185
R1577 vdd.n2531 vdd.n2530 185
R1578 vdd.n2532 vdd.n2531 185
R1579 vdd.n964 vdd.n962 185
R1580 vdd.n962 vdd.t268 185
R1581 vdd.n2446 vdd.n971 185
R1582 vdd.n2457 vdd.n971 185
R1583 vdd.n2447 vdd.n980 185
R1584 vdd.n2156 vdd.n980 185
R1585 vdd.n2449 vdd.n2448 185
R1586 vdd.n2450 vdd.n2449 185
R1587 vdd.n2445 vdd.n979 185
R1588 vdd.n979 vdd.n976 185
R1589 vdd.n2444 vdd.n2443 185
R1590 vdd.n2443 vdd.n2442 185
R1591 vdd.n982 vdd.n981 185
R1592 vdd.n983 vdd.n982 185
R1593 vdd.n2435 vdd.n2434 185
R1594 vdd.n2436 vdd.n2435 185
R1595 vdd.n2433 vdd.n992 185
R1596 vdd.n992 vdd.n989 185
R1597 vdd.n2432 vdd.n2431 185
R1598 vdd.n2431 vdd.n2430 185
R1599 vdd.n994 vdd.n993 185
R1600 vdd.n1002 vdd.n994 185
R1601 vdd.n2423 vdd.n2422 185
R1602 vdd.n2424 vdd.n2423 185
R1603 vdd.n2421 vdd.n1003 185
R1604 vdd.n1008 vdd.n1003 185
R1605 vdd.n2420 vdd.n2419 185
R1606 vdd.n2419 vdd.n2418 185
R1607 vdd.n1005 vdd.n1004 185
R1608 vdd.n2257 vdd.n1005 185
R1609 vdd.n2411 vdd.n2410 185
R1610 vdd.n2412 vdd.n2411 185
R1611 vdd.n2409 vdd.n1015 185
R1612 vdd.n1015 vdd.n1012 185
R1613 vdd.n2408 vdd.n2407 185
R1614 vdd.n2407 vdd.n2406 185
R1615 vdd.n1017 vdd.n1016 185
R1616 vdd.n1018 vdd.n1017 185
R1617 vdd.n2399 vdd.n2398 185
R1618 vdd.n2400 vdd.n2399 185
R1619 vdd.n2396 vdd.n1026 185
R1620 vdd.n1033 vdd.n1026 185
R1621 vdd.n2395 vdd.n2394 185
R1622 vdd.n2394 vdd.n2393 185
R1623 vdd.n1029 vdd.n1028 185
R1624 vdd.n1030 vdd.n1029 185
R1625 vdd.n2386 vdd.n2385 185
R1626 vdd.n2387 vdd.n2386 185
R1627 vdd.n2384 vdd.n1040 185
R1628 vdd.n1040 vdd.n1037 185
R1629 vdd.n2383 vdd.n2382 185
R1630 vdd.n2382 vdd.n2381 185
R1631 vdd.n1042 vdd.n1041 185
R1632 vdd.n1043 vdd.n1042 185
R1633 vdd.n2374 vdd.n2373 185
R1634 vdd.n2375 vdd.n2374 185
R1635 vdd.n2462 vdd.n936 185
R1636 vdd.n2604 vdd.n936 185
R1637 vdd.n2464 vdd.n2463 185
R1638 vdd.n2466 vdd.n2465 185
R1639 vdd.n2468 vdd.n2467 185
R1640 vdd.n2470 vdd.n2469 185
R1641 vdd.n2472 vdd.n2471 185
R1642 vdd.n2474 vdd.n2473 185
R1643 vdd.n2476 vdd.n2475 185
R1644 vdd.n2478 vdd.n2477 185
R1645 vdd.n2480 vdd.n2479 185
R1646 vdd.n2482 vdd.n2481 185
R1647 vdd.n2484 vdd.n2483 185
R1648 vdd.n2486 vdd.n2485 185
R1649 vdd.n2488 vdd.n2487 185
R1650 vdd.n2490 vdd.n2489 185
R1651 vdd.n2492 vdd.n2491 185
R1652 vdd.n2494 vdd.n2493 185
R1653 vdd.n2496 vdd.n2495 185
R1654 vdd.n2498 vdd.n2497 185
R1655 vdd.n2500 vdd.n2499 185
R1656 vdd.n2502 vdd.n2501 185
R1657 vdd.n2504 vdd.n2503 185
R1658 vdd.n2506 vdd.n2505 185
R1659 vdd.n2508 vdd.n2507 185
R1660 vdd.n2510 vdd.n2509 185
R1661 vdd.n2512 vdd.n2511 185
R1662 vdd.n2514 vdd.n2513 185
R1663 vdd.n2516 vdd.n2515 185
R1664 vdd.n2518 vdd.n2517 185
R1665 vdd.n2520 vdd.n2519 185
R1666 vdd.n2522 vdd.n2521 185
R1667 vdd.n2524 vdd.n2523 185
R1668 vdd.n2526 vdd.n2525 185
R1669 vdd.n2528 vdd.n2527 185
R1670 vdd.n2529 vdd.n963 185
R1671 vdd.n2461 vdd.n961 185
R1672 vdd.n2532 vdd.n961 185
R1673 vdd.n2460 vdd.n2459 185
R1674 vdd.n2459 vdd.t268 185
R1675 vdd.n2458 vdd.n968 185
R1676 vdd.n2458 vdd.n2457 185
R1677 vdd.n2238 vdd.n969 185
R1678 vdd.n2156 vdd.n969 185
R1679 vdd.n2239 vdd.n978 185
R1680 vdd.n2450 vdd.n978 185
R1681 vdd.n2241 vdd.n2240 185
R1682 vdd.n2240 vdd.n976 185
R1683 vdd.n2242 vdd.n985 185
R1684 vdd.n2442 vdd.n985 185
R1685 vdd.n2244 vdd.n2243 185
R1686 vdd.n2243 vdd.n983 185
R1687 vdd.n2245 vdd.n991 185
R1688 vdd.n2436 vdd.n991 185
R1689 vdd.n2247 vdd.n2246 185
R1690 vdd.n2246 vdd.n989 185
R1691 vdd.n2248 vdd.n996 185
R1692 vdd.n2430 vdd.n996 185
R1693 vdd.n2250 vdd.n2249 185
R1694 vdd.n2249 vdd.n1002 185
R1695 vdd.n2251 vdd.n1001 185
R1696 vdd.n2424 vdd.n1001 185
R1697 vdd.n2253 vdd.n2252 185
R1698 vdd.n2252 vdd.n1008 185
R1699 vdd.n2254 vdd.n1007 185
R1700 vdd.n2418 vdd.n1007 185
R1701 vdd.n2256 vdd.n2255 185
R1702 vdd.n2257 vdd.n2256 185
R1703 vdd.n2237 vdd.n1014 185
R1704 vdd.n2412 vdd.n1014 185
R1705 vdd.n2236 vdd.n2235 185
R1706 vdd.n2235 vdd.n1012 185
R1707 vdd.n2234 vdd.n1020 185
R1708 vdd.n2406 vdd.n1020 185
R1709 vdd.n2233 vdd.n2232 185
R1710 vdd.n2232 vdd.n1018 185
R1711 vdd.n2231 vdd.n1025 185
R1712 vdd.n2400 vdd.n1025 185
R1713 vdd.n2230 vdd.n2229 185
R1714 vdd.n2229 vdd.n1033 185
R1715 vdd.n2228 vdd.n1032 185
R1716 vdd.n2393 vdd.n1032 185
R1717 vdd.n2227 vdd.n2226 185
R1718 vdd.n2226 vdd.n1030 185
R1719 vdd.n2225 vdd.n1039 185
R1720 vdd.n2387 vdd.n1039 185
R1721 vdd.n2224 vdd.n2223 185
R1722 vdd.n2223 vdd.n1037 185
R1723 vdd.n2222 vdd.n1045 185
R1724 vdd.n2381 vdd.n1045 185
R1725 vdd.n2221 vdd.n2220 185
R1726 vdd.n2220 vdd.n1043 185
R1727 vdd.n2219 vdd.n1051 185
R1728 vdd.n2375 vdd.n1051 185
R1729 vdd.n2372 vdd.n1052 185
R1730 vdd.n2371 vdd.n2370 185
R1731 vdd.n2368 vdd.n1053 185
R1732 vdd.n2366 vdd.n2365 185
R1733 vdd.n2364 vdd.n1054 185
R1734 vdd.n2363 vdd.n2362 185
R1735 vdd.n2360 vdd.n1055 185
R1736 vdd.n2358 vdd.n2357 185
R1737 vdd.n2356 vdd.n1056 185
R1738 vdd.n2355 vdd.n2354 185
R1739 vdd.n2352 vdd.n1057 185
R1740 vdd.n2350 vdd.n2349 185
R1741 vdd.n2348 vdd.n1058 185
R1742 vdd.n2347 vdd.n2346 185
R1743 vdd.n2344 vdd.n1059 185
R1744 vdd.n2342 vdd.n2341 185
R1745 vdd.n2340 vdd.n1060 185
R1746 vdd.n2339 vdd.n1062 185
R1747 vdd.n2184 vdd.n1063 185
R1748 vdd.n2187 vdd.n2186 185
R1749 vdd.n2189 vdd.n2188 185
R1750 vdd.n2191 vdd.n2183 185
R1751 vdd.n2194 vdd.n2193 185
R1752 vdd.n2195 vdd.n2182 185
R1753 vdd.n2197 vdd.n2196 185
R1754 vdd.n2199 vdd.n2181 185
R1755 vdd.n2202 vdd.n2201 185
R1756 vdd.n2203 vdd.n2180 185
R1757 vdd.n2205 vdd.n2204 185
R1758 vdd.n2207 vdd.n2179 185
R1759 vdd.n2210 vdd.n2209 185
R1760 vdd.n2211 vdd.n2176 185
R1761 vdd.n2214 vdd.n2213 185
R1762 vdd.n2216 vdd.n2175 185
R1763 vdd.n2218 vdd.n2217 185
R1764 vdd.n2217 vdd.n1049 185
R1765 vdd.n327 vdd.n326 171.744
R1766 vdd.n326 vdd.n325 171.744
R1767 vdd.n325 vdd.n294 171.744
R1768 vdd.n318 vdd.n294 171.744
R1769 vdd.n318 vdd.n317 171.744
R1770 vdd.n317 vdd.n299 171.744
R1771 vdd.n310 vdd.n299 171.744
R1772 vdd.n310 vdd.n309 171.744
R1773 vdd.n309 vdd.n303 171.744
R1774 vdd.n268 vdd.n267 171.744
R1775 vdd.n267 vdd.n266 171.744
R1776 vdd.n266 vdd.n235 171.744
R1777 vdd.n259 vdd.n235 171.744
R1778 vdd.n259 vdd.n258 171.744
R1779 vdd.n258 vdd.n240 171.744
R1780 vdd.n251 vdd.n240 171.744
R1781 vdd.n251 vdd.n250 171.744
R1782 vdd.n250 vdd.n244 171.744
R1783 vdd.n225 vdd.n224 171.744
R1784 vdd.n224 vdd.n223 171.744
R1785 vdd.n223 vdd.n192 171.744
R1786 vdd.n216 vdd.n192 171.744
R1787 vdd.n216 vdd.n215 171.744
R1788 vdd.n215 vdd.n197 171.744
R1789 vdd.n208 vdd.n197 171.744
R1790 vdd.n208 vdd.n207 171.744
R1791 vdd.n207 vdd.n201 171.744
R1792 vdd.n166 vdd.n165 171.744
R1793 vdd.n165 vdd.n164 171.744
R1794 vdd.n164 vdd.n133 171.744
R1795 vdd.n157 vdd.n133 171.744
R1796 vdd.n157 vdd.n156 171.744
R1797 vdd.n156 vdd.n138 171.744
R1798 vdd.n149 vdd.n138 171.744
R1799 vdd.n149 vdd.n148 171.744
R1800 vdd.n148 vdd.n142 171.744
R1801 vdd.n124 vdd.n123 171.744
R1802 vdd.n123 vdd.n122 171.744
R1803 vdd.n122 vdd.n91 171.744
R1804 vdd.n115 vdd.n91 171.744
R1805 vdd.n115 vdd.n114 171.744
R1806 vdd.n114 vdd.n96 171.744
R1807 vdd.n107 vdd.n96 171.744
R1808 vdd.n107 vdd.n106 171.744
R1809 vdd.n106 vdd.n100 171.744
R1810 vdd.n65 vdd.n64 171.744
R1811 vdd.n64 vdd.n63 171.744
R1812 vdd.n63 vdd.n32 171.744
R1813 vdd.n56 vdd.n32 171.744
R1814 vdd.n56 vdd.n55 171.744
R1815 vdd.n55 vdd.n37 171.744
R1816 vdd.n48 vdd.n37 171.744
R1817 vdd.n48 vdd.n47 171.744
R1818 vdd.n47 vdd.n41 171.744
R1819 vdd.n1746 vdd.n1745 171.744
R1820 vdd.n1745 vdd.n1744 171.744
R1821 vdd.n1744 vdd.n1713 171.744
R1822 vdd.n1737 vdd.n1713 171.744
R1823 vdd.n1737 vdd.n1736 171.744
R1824 vdd.n1736 vdd.n1718 171.744
R1825 vdd.n1729 vdd.n1718 171.744
R1826 vdd.n1729 vdd.n1728 171.744
R1827 vdd.n1728 vdd.n1722 171.744
R1828 vdd.n1805 vdd.n1804 171.744
R1829 vdd.n1804 vdd.n1803 171.744
R1830 vdd.n1803 vdd.n1772 171.744
R1831 vdd.n1796 vdd.n1772 171.744
R1832 vdd.n1796 vdd.n1795 171.744
R1833 vdd.n1795 vdd.n1777 171.744
R1834 vdd.n1788 vdd.n1777 171.744
R1835 vdd.n1788 vdd.n1787 171.744
R1836 vdd.n1787 vdd.n1781 171.744
R1837 vdd.n1644 vdd.n1643 171.744
R1838 vdd.n1643 vdd.n1642 171.744
R1839 vdd.n1642 vdd.n1611 171.744
R1840 vdd.n1635 vdd.n1611 171.744
R1841 vdd.n1635 vdd.n1634 171.744
R1842 vdd.n1634 vdd.n1616 171.744
R1843 vdd.n1627 vdd.n1616 171.744
R1844 vdd.n1627 vdd.n1626 171.744
R1845 vdd.n1626 vdd.n1620 171.744
R1846 vdd.n1703 vdd.n1702 171.744
R1847 vdd.n1702 vdd.n1701 171.744
R1848 vdd.n1701 vdd.n1670 171.744
R1849 vdd.n1694 vdd.n1670 171.744
R1850 vdd.n1694 vdd.n1693 171.744
R1851 vdd.n1693 vdd.n1675 171.744
R1852 vdd.n1686 vdd.n1675 171.744
R1853 vdd.n1686 vdd.n1685 171.744
R1854 vdd.n1685 vdd.n1679 171.744
R1855 vdd.n1543 vdd.n1542 171.744
R1856 vdd.n1542 vdd.n1541 171.744
R1857 vdd.n1541 vdd.n1510 171.744
R1858 vdd.n1534 vdd.n1510 171.744
R1859 vdd.n1534 vdd.n1533 171.744
R1860 vdd.n1533 vdd.n1515 171.744
R1861 vdd.n1526 vdd.n1515 171.744
R1862 vdd.n1526 vdd.n1525 171.744
R1863 vdd.n1525 vdd.n1519 171.744
R1864 vdd.n1602 vdd.n1601 171.744
R1865 vdd.n1601 vdd.n1600 171.744
R1866 vdd.n1600 vdd.n1569 171.744
R1867 vdd.n1593 vdd.n1569 171.744
R1868 vdd.n1593 vdd.n1592 171.744
R1869 vdd.n1592 vdd.n1574 171.744
R1870 vdd.n1585 vdd.n1574 171.744
R1871 vdd.n1585 vdd.n1584 171.744
R1872 vdd.n1584 vdd.n1578 171.744
R1873 vdd.n468 vdd.n467 146.341
R1874 vdd.n474 vdd.n473 146.341
R1875 vdd.n478 vdd.n477 146.341
R1876 vdd.n484 vdd.n483 146.341
R1877 vdd.n488 vdd.n487 146.341
R1878 vdd.n494 vdd.n493 146.341
R1879 vdd.n498 vdd.n497 146.341
R1880 vdd.n504 vdd.n503 146.341
R1881 vdd.n508 vdd.n507 146.341
R1882 vdd.n514 vdd.n513 146.341
R1883 vdd.n518 vdd.n517 146.341
R1884 vdd.n524 vdd.n523 146.341
R1885 vdd.n528 vdd.n527 146.341
R1886 vdd.n534 vdd.n533 146.341
R1887 vdd.n538 vdd.n537 146.341
R1888 vdd.n544 vdd.n543 146.341
R1889 vdd.n548 vdd.n547 146.341
R1890 vdd.n554 vdd.n553 146.341
R1891 vdd.n558 vdd.n557 146.341
R1892 vdd.n564 vdd.n563 146.341
R1893 vdd.n568 vdd.n567 146.341
R1894 vdd.n574 vdd.n573 146.341
R1895 vdd.n578 vdd.n577 146.341
R1896 vdd.n584 vdd.n583 146.341
R1897 vdd.n588 vdd.n587 146.341
R1898 vdd.n594 vdd.n593 146.341
R1899 vdd.n598 vdd.n597 146.341
R1900 vdd.n604 vdd.n603 146.341
R1901 vdd.n608 vdd.n607 146.341
R1902 vdd.n614 vdd.n613 146.341
R1903 vdd.n616 vdd.n425 146.341
R1904 vdd.n3230 vdd.n685 146.341
R1905 vdd.n3230 vdd.n677 146.341
R1906 vdd.n3240 vdd.n677 146.341
R1907 vdd.n3240 vdd.n673 146.341
R1908 vdd.n3246 vdd.n673 146.341
R1909 vdd.n3246 vdd.n667 146.341
R1910 vdd.n3257 vdd.n667 146.341
R1911 vdd.n3257 vdd.n663 146.341
R1912 vdd.n3263 vdd.n663 146.341
R1913 vdd.n3263 vdd.n654 146.341
R1914 vdd.n3273 vdd.n654 146.341
R1915 vdd.n3273 vdd.n650 146.341
R1916 vdd.n3279 vdd.n650 146.341
R1917 vdd.n3279 vdd.n643 146.341
R1918 vdd.n3290 vdd.n643 146.341
R1919 vdd.n3290 vdd.n639 146.341
R1920 vdd.n3299 vdd.n639 146.341
R1921 vdd.n3299 vdd.n632 146.341
R1922 vdd.n3309 vdd.n632 146.341
R1923 vdd.n3310 vdd.n3309 146.341
R1924 vdd.n3310 vdd.n341 146.341
R1925 vdd.n342 vdd.n341 146.341
R1926 vdd.n343 vdd.n342 146.341
R1927 vdd.n3317 vdd.n343 146.341
R1928 vdd.n3317 vdd.n351 146.341
R1929 vdd.n352 vdd.n351 146.341
R1930 vdd.n353 vdd.n352 146.341
R1931 vdd.n3324 vdd.n353 146.341
R1932 vdd.n3324 vdd.n362 146.341
R1933 vdd.n363 vdd.n362 146.341
R1934 vdd.n364 vdd.n363 146.341
R1935 vdd.n3332 vdd.n364 146.341
R1936 vdd.n3332 vdd.n372 146.341
R1937 vdd.n373 vdd.n372 146.341
R1938 vdd.n374 vdd.n373 146.341
R1939 vdd.n3339 vdd.n374 146.341
R1940 vdd.n3339 vdd.n383 146.341
R1941 vdd.n384 vdd.n383 146.341
R1942 vdd.n385 vdd.n384 146.341
R1943 vdd.n3346 vdd.n385 146.341
R1944 vdd.n3346 vdd.n393 146.341
R1945 vdd.n725 vdd.n724 146.341
R1946 vdd.n728 vdd.n724 146.341
R1947 vdd.n734 vdd.n733 146.341
R1948 vdd.n3212 vdd.n3211 146.341
R1949 vdd.n3208 vdd.n3207 146.341
R1950 vdd.n3204 vdd.n3203 146.341
R1951 vdd.n3200 vdd.n3199 146.341
R1952 vdd.n3196 vdd.n3195 146.341
R1953 vdd.n3192 vdd.n3191 146.341
R1954 vdd.n3188 vdd.n3187 146.341
R1955 vdd.n3179 vdd.n3178 146.341
R1956 vdd.n3176 vdd.n3175 146.341
R1957 vdd.n3172 vdd.n3171 146.341
R1958 vdd.n3168 vdd.n3167 146.341
R1959 vdd.n3164 vdd.n3163 146.341
R1960 vdd.n3160 vdd.n3159 146.341
R1961 vdd.n3156 vdd.n3155 146.341
R1962 vdd.n3152 vdd.n3151 146.341
R1963 vdd.n3148 vdd.n3147 146.341
R1964 vdd.n3144 vdd.n3143 146.341
R1965 vdd.n3140 vdd.n3139 146.341
R1966 vdd.n3133 vdd.n3132 146.341
R1967 vdd.n3130 vdd.n3129 146.341
R1968 vdd.n3126 vdd.n3125 146.341
R1969 vdd.n3122 vdd.n3121 146.341
R1970 vdd.n3118 vdd.n3117 146.341
R1971 vdd.n3114 vdd.n3113 146.341
R1972 vdd.n3110 vdd.n3109 146.341
R1973 vdd.n3106 vdd.n3105 146.341
R1974 vdd.n3102 vdd.n3101 146.341
R1975 vdd.n3098 vdd.n3097 146.341
R1976 vdd.n3224 vdd.n691 146.341
R1977 vdd.n3232 vdd.n684 146.341
R1978 vdd.n3232 vdd.n680 146.341
R1979 vdd.n3238 vdd.n680 146.341
R1980 vdd.n3238 vdd.n672 146.341
R1981 vdd.n3249 vdd.n672 146.341
R1982 vdd.n3249 vdd.n668 146.341
R1983 vdd.n3255 vdd.n668 146.341
R1984 vdd.n3255 vdd.n661 146.341
R1985 vdd.n3265 vdd.n661 146.341
R1986 vdd.n3265 vdd.n657 146.341
R1987 vdd.n3271 vdd.n657 146.341
R1988 vdd.n3271 vdd.n649 146.341
R1989 vdd.n3282 vdd.n649 146.341
R1990 vdd.n3282 vdd.n645 146.341
R1991 vdd.n3288 vdd.n645 146.341
R1992 vdd.n3288 vdd.n638 146.341
R1993 vdd.n3301 vdd.n638 146.341
R1994 vdd.n3301 vdd.n634 146.341
R1995 vdd.n3307 vdd.n634 146.341
R1996 vdd.n3307 vdd.n338 146.341
R1997 vdd.n3396 vdd.n338 146.341
R1998 vdd.n3396 vdd.n339 146.341
R1999 vdd.n3392 vdd.n339 146.341
R2000 vdd.n3392 vdd.n345 146.341
R2001 vdd.n3388 vdd.n345 146.341
R2002 vdd.n3388 vdd.n350 146.341
R2003 vdd.n3384 vdd.n350 146.341
R2004 vdd.n3384 vdd.n354 146.341
R2005 vdd.n3380 vdd.n354 146.341
R2006 vdd.n3380 vdd.n360 146.341
R2007 vdd.n3376 vdd.n360 146.341
R2008 vdd.n3376 vdd.n365 146.341
R2009 vdd.n3372 vdd.n365 146.341
R2010 vdd.n3372 vdd.n371 146.341
R2011 vdd.n3368 vdd.n371 146.341
R2012 vdd.n3368 vdd.n376 146.341
R2013 vdd.n3364 vdd.n376 146.341
R2014 vdd.n3364 vdd.n382 146.341
R2015 vdd.n3360 vdd.n382 146.341
R2016 vdd.n3360 vdd.n387 146.341
R2017 vdd.n3356 vdd.n387 146.341
R2018 vdd.n2322 vdd.n2321 146.341
R2019 vdd.n2319 vdd.n1903 146.341
R2020 vdd.n2099 vdd.n1909 146.341
R2021 vdd.n2097 vdd.n2096 146.341
R2022 vdd.n2094 vdd.n1911 146.341
R2023 vdd.n2090 vdd.n2089 146.341
R2024 vdd.n2087 vdd.n1918 146.341
R2025 vdd.n2083 vdd.n2082 146.341
R2026 vdd.n2080 vdd.n1925 146.341
R2027 vdd.n1936 vdd.n1933 146.341
R2028 vdd.n2072 vdd.n2071 146.341
R2029 vdd.n2069 vdd.n1938 146.341
R2030 vdd.n2065 vdd.n2064 146.341
R2031 vdd.n2062 vdd.n1944 146.341
R2032 vdd.n2058 vdd.n2057 146.341
R2033 vdd.n2055 vdd.n1951 146.341
R2034 vdd.n2051 vdd.n2050 146.341
R2035 vdd.n2048 vdd.n1958 146.341
R2036 vdd.n2044 vdd.n2043 146.341
R2037 vdd.n2041 vdd.n1965 146.341
R2038 vdd.n1976 vdd.n1973 146.341
R2039 vdd.n2033 vdd.n2032 146.341
R2040 vdd.n2030 vdd.n1978 146.341
R2041 vdd.n2026 vdd.n2025 146.341
R2042 vdd.n2023 vdd.n1984 146.341
R2043 vdd.n2019 vdd.n2018 146.341
R2044 vdd.n2016 vdd.n1991 146.341
R2045 vdd.n2012 vdd.n2011 146.341
R2046 vdd.n2009 vdd.n2006 146.341
R2047 vdd.n2004 vdd.n2001 146.341
R2048 vdd.n1999 vdd.n1069 146.341
R2049 vdd.n1428 vdd.n1188 146.341
R2050 vdd.n1428 vdd.n1184 146.341
R2051 vdd.n1434 vdd.n1184 146.341
R2052 vdd.n1434 vdd.n1176 146.341
R2053 vdd.n1445 vdd.n1176 146.341
R2054 vdd.n1445 vdd.n1172 146.341
R2055 vdd.n1451 vdd.n1172 146.341
R2056 vdd.n1451 vdd.n1166 146.341
R2057 vdd.n1462 vdd.n1166 146.341
R2058 vdd.n1462 vdd.n1162 146.341
R2059 vdd.n1468 vdd.n1162 146.341
R2060 vdd.n1468 vdd.n1153 146.341
R2061 vdd.n1478 vdd.n1153 146.341
R2062 vdd.n1478 vdd.n1149 146.341
R2063 vdd.n1484 vdd.n1149 146.341
R2064 vdd.n1484 vdd.n1142 146.341
R2065 vdd.n1495 vdd.n1142 146.341
R2066 vdd.n1495 vdd.n1138 146.341
R2067 vdd.n1501 vdd.n1138 146.341
R2068 vdd.n1501 vdd.n1131 146.341
R2069 vdd.n1818 vdd.n1131 146.341
R2070 vdd.n1818 vdd.n1127 146.341
R2071 vdd.n1824 vdd.n1127 146.341
R2072 vdd.n1824 vdd.n1119 146.341
R2073 vdd.n1835 vdd.n1119 146.341
R2074 vdd.n1835 vdd.n1115 146.341
R2075 vdd.n1841 vdd.n1115 146.341
R2076 vdd.n1841 vdd.n1109 146.341
R2077 vdd.n1852 vdd.n1109 146.341
R2078 vdd.n1852 vdd.n1105 146.341
R2079 vdd.n1858 vdd.n1105 146.341
R2080 vdd.n1858 vdd.n1096 146.341
R2081 vdd.n1868 vdd.n1096 146.341
R2082 vdd.n1868 vdd.n1092 146.341
R2083 vdd.n1874 vdd.n1092 146.341
R2084 vdd.n1874 vdd.n1086 146.341
R2085 vdd.n1885 vdd.n1086 146.341
R2086 vdd.n1885 vdd.n1081 146.341
R2087 vdd.n1893 vdd.n1081 146.341
R2088 vdd.n1893 vdd.n1071 146.341
R2089 vdd.n2330 vdd.n1071 146.341
R2090 vdd.n1417 vdd.n1193 146.341
R2091 vdd.n1417 vdd.n1226 146.341
R2092 vdd.n1230 vdd.n1229 146.341
R2093 vdd.n1232 vdd.n1231 146.341
R2094 vdd.n1236 vdd.n1235 146.341
R2095 vdd.n1238 vdd.n1237 146.341
R2096 vdd.n1242 vdd.n1241 146.341
R2097 vdd.n1244 vdd.n1243 146.341
R2098 vdd.n1248 vdd.n1247 146.341
R2099 vdd.n1250 vdd.n1249 146.341
R2100 vdd.n1256 vdd.n1255 146.341
R2101 vdd.n1258 vdd.n1257 146.341
R2102 vdd.n1262 vdd.n1261 146.341
R2103 vdd.n1264 vdd.n1263 146.341
R2104 vdd.n1268 vdd.n1267 146.341
R2105 vdd.n1270 vdd.n1269 146.341
R2106 vdd.n1274 vdd.n1273 146.341
R2107 vdd.n1276 vdd.n1275 146.341
R2108 vdd.n1280 vdd.n1279 146.341
R2109 vdd.n1282 vdd.n1281 146.341
R2110 vdd.n1354 vdd.n1285 146.341
R2111 vdd.n1287 vdd.n1286 146.341
R2112 vdd.n1291 vdd.n1290 146.341
R2113 vdd.n1293 vdd.n1292 146.341
R2114 vdd.n1297 vdd.n1296 146.341
R2115 vdd.n1299 vdd.n1298 146.341
R2116 vdd.n1303 vdd.n1302 146.341
R2117 vdd.n1305 vdd.n1304 146.341
R2118 vdd.n1309 vdd.n1308 146.341
R2119 vdd.n1311 vdd.n1310 146.341
R2120 vdd.n1315 vdd.n1314 146.341
R2121 vdd.n1316 vdd.n1224 146.341
R2122 vdd.n1426 vdd.n1189 146.341
R2123 vdd.n1426 vdd.n1182 146.341
R2124 vdd.n1437 vdd.n1182 146.341
R2125 vdd.n1437 vdd.n1178 146.341
R2126 vdd.n1443 vdd.n1178 146.341
R2127 vdd.n1443 vdd.n1171 146.341
R2128 vdd.n1454 vdd.n1171 146.341
R2129 vdd.n1454 vdd.n1167 146.341
R2130 vdd.n1460 vdd.n1167 146.341
R2131 vdd.n1460 vdd.n1160 146.341
R2132 vdd.n1470 vdd.n1160 146.341
R2133 vdd.n1470 vdd.n1156 146.341
R2134 vdd.n1476 vdd.n1156 146.341
R2135 vdd.n1476 vdd.n1148 146.341
R2136 vdd.n1487 vdd.n1148 146.341
R2137 vdd.n1487 vdd.n1144 146.341
R2138 vdd.n1493 vdd.n1144 146.341
R2139 vdd.n1493 vdd.n1137 146.341
R2140 vdd.n1503 vdd.n1137 146.341
R2141 vdd.n1503 vdd.n1133 146.341
R2142 vdd.n1816 vdd.n1133 146.341
R2143 vdd.n1816 vdd.n1125 146.341
R2144 vdd.n1827 vdd.n1125 146.341
R2145 vdd.n1827 vdd.n1121 146.341
R2146 vdd.n1833 vdd.n1121 146.341
R2147 vdd.n1833 vdd.n1114 146.341
R2148 vdd.n1844 vdd.n1114 146.341
R2149 vdd.n1844 vdd.n1110 146.341
R2150 vdd.n1850 vdd.n1110 146.341
R2151 vdd.n1850 vdd.n1103 146.341
R2152 vdd.n1860 vdd.n1103 146.341
R2153 vdd.n1860 vdd.n1099 146.341
R2154 vdd.n1866 vdd.n1099 146.341
R2155 vdd.n1866 vdd.n1091 146.341
R2156 vdd.n1877 vdd.n1091 146.341
R2157 vdd.n1877 vdd.n1087 146.341
R2158 vdd.n1883 vdd.n1087 146.341
R2159 vdd.n1883 vdd.n1079 146.341
R2160 vdd.n1896 vdd.n1079 146.341
R2161 vdd.n1896 vdd.n1074 146.341
R2162 vdd.n2328 vdd.n1074 146.341
R2163 vdd.n1073 vdd.n1049 141.707
R2164 vdd.n3223 vdd.n692 141.707
R2165 vdd.n2177 vdd.t197 127.284
R2166 vdd.n965 vdd.t181 127.284
R2167 vdd.n2151 vdd.t219 127.284
R2168 vdd.n957 vdd.t206 127.284
R2169 vdd.n2922 vdd.t157 127.284
R2170 vdd.n2922 vdd.t158 127.284
R2171 vdd.n2642 vdd.t204 127.284
R2172 vdd.n832 vdd.t185 127.284
R2173 vdd.n2639 vdd.t190 127.284
R2174 vdd.n799 vdd.t192 127.284
R2175 vdd.n1027 vdd.t200 127.284
R2176 vdd.n1027 vdd.t201 127.284
R2177 vdd.n22 vdd.n20 117.314
R2178 vdd.n17 vdd.n15 117.314
R2179 vdd.n27 vdd.n26 116.927
R2180 vdd.n24 vdd.n23 116.927
R2181 vdd.n22 vdd.n21 116.927
R2182 vdd.n17 vdd.n16 116.927
R2183 vdd.n19 vdd.n18 116.927
R2184 vdd.n27 vdd.n25 116.927
R2185 vdd.n2178 vdd.t196 111.188
R2186 vdd.n966 vdd.t182 111.188
R2187 vdd.n2152 vdd.t218 111.188
R2188 vdd.n958 vdd.t207 111.188
R2189 vdd.n2643 vdd.t203 111.188
R2190 vdd.n833 vdd.t186 111.188
R2191 vdd.n2640 vdd.t189 111.188
R2192 vdd.n800 vdd.t193 111.188
R2193 vdd.n2865 vdd.n911 99.5127
R2194 vdd.n2869 vdd.n911 99.5127
R2195 vdd.n2869 vdd.n903 99.5127
R2196 vdd.n2877 vdd.n903 99.5127
R2197 vdd.n2877 vdd.n901 99.5127
R2198 vdd.n2881 vdd.n901 99.5127
R2199 vdd.n2881 vdd.n890 99.5127
R2200 vdd.n2889 vdd.n890 99.5127
R2201 vdd.n2889 vdd.n888 99.5127
R2202 vdd.n2893 vdd.n888 99.5127
R2203 vdd.n2893 vdd.n879 99.5127
R2204 vdd.n2901 vdd.n879 99.5127
R2205 vdd.n2901 vdd.n877 99.5127
R2206 vdd.n2905 vdd.n877 99.5127
R2207 vdd.n2905 vdd.n867 99.5127
R2208 vdd.n2913 vdd.n867 99.5127
R2209 vdd.n2913 vdd.n865 99.5127
R2210 vdd.n2917 vdd.n865 99.5127
R2211 vdd.n2917 vdd.n856 99.5127
R2212 vdd.n2927 vdd.n856 99.5127
R2213 vdd.n2927 vdd.n854 99.5127
R2214 vdd.n2931 vdd.n854 99.5127
R2215 vdd.n2931 vdd.n842 99.5127
R2216 vdd.n2984 vdd.n842 99.5127
R2217 vdd.n2984 vdd.n840 99.5127
R2218 vdd.n2988 vdd.n840 99.5127
R2219 vdd.n2988 vdd.n808 99.5127
R2220 vdd.n3058 vdd.n808 99.5127
R2221 vdd.n3054 vdd.n809 99.5127
R2222 vdd.n3052 vdd.n3051 99.5127
R2223 vdd.n3049 vdd.n813 99.5127
R2224 vdd.n3045 vdd.n3044 99.5127
R2225 vdd.n3042 vdd.n816 99.5127
R2226 vdd.n3038 vdd.n3037 99.5127
R2227 vdd.n3035 vdd.n819 99.5127
R2228 vdd.n3031 vdd.n3030 99.5127
R2229 vdd.n3028 vdd.n3026 99.5127
R2230 vdd.n3024 vdd.n822 99.5127
R2231 vdd.n3020 vdd.n3019 99.5127
R2232 vdd.n3017 vdd.n825 99.5127
R2233 vdd.n3013 vdd.n3012 99.5127
R2234 vdd.n3010 vdd.n828 99.5127
R2235 vdd.n3006 vdd.n3005 99.5127
R2236 vdd.n3003 vdd.n831 99.5127
R2237 vdd.n2998 vdd.n2997 99.5127
R2238 vdd.n2785 vdd.n914 99.5127
R2239 vdd.n2785 vdd.n909 99.5127
R2240 vdd.n2782 vdd.n909 99.5127
R2241 vdd.n2782 vdd.n904 99.5127
R2242 vdd.n2729 vdd.n904 99.5127
R2243 vdd.n2729 vdd.n898 99.5127
R2244 vdd.n2732 vdd.n898 99.5127
R2245 vdd.n2732 vdd.n891 99.5127
R2246 vdd.n2735 vdd.n891 99.5127
R2247 vdd.n2735 vdd.n886 99.5127
R2248 vdd.n2738 vdd.n886 99.5127
R2249 vdd.n2738 vdd.n881 99.5127
R2250 vdd.n2741 vdd.n881 99.5127
R2251 vdd.n2741 vdd.n875 99.5127
R2252 vdd.n2759 vdd.n875 99.5127
R2253 vdd.n2759 vdd.n868 99.5127
R2254 vdd.n2755 vdd.n868 99.5127
R2255 vdd.n2755 vdd.n863 99.5127
R2256 vdd.n2752 vdd.n863 99.5127
R2257 vdd.n2752 vdd.n858 99.5127
R2258 vdd.n2749 vdd.n858 99.5127
R2259 vdd.n2749 vdd.n852 99.5127
R2260 vdd.n2746 vdd.n852 99.5127
R2261 vdd.n2746 vdd.n844 99.5127
R2262 vdd.n844 vdd.n837 99.5127
R2263 vdd.n2990 vdd.n837 99.5127
R2264 vdd.n2991 vdd.n2990 99.5127
R2265 vdd.n2991 vdd.n806 99.5127
R2266 vdd.n2855 vdd.n2638 99.5127
R2267 vdd.n2851 vdd.n2638 99.5127
R2268 vdd.n2849 vdd.n2848 99.5127
R2269 vdd.n2845 vdd.n2844 99.5127
R2270 vdd.n2841 vdd.n2840 99.5127
R2271 vdd.n2837 vdd.n2836 99.5127
R2272 vdd.n2833 vdd.n2832 99.5127
R2273 vdd.n2829 vdd.n2828 99.5127
R2274 vdd.n2825 vdd.n2824 99.5127
R2275 vdd.n2821 vdd.n2820 99.5127
R2276 vdd.n2817 vdd.n2816 99.5127
R2277 vdd.n2813 vdd.n2812 99.5127
R2278 vdd.n2809 vdd.n2808 99.5127
R2279 vdd.n2805 vdd.n2804 99.5127
R2280 vdd.n2801 vdd.n2800 99.5127
R2281 vdd.n2797 vdd.n2796 99.5127
R2282 vdd.n2792 vdd.n2791 99.5127
R2283 vdd.n2603 vdd.n955 99.5127
R2284 vdd.n2599 vdd.n2598 99.5127
R2285 vdd.n2595 vdd.n2594 99.5127
R2286 vdd.n2591 vdd.n2590 99.5127
R2287 vdd.n2587 vdd.n2586 99.5127
R2288 vdd.n2583 vdd.n2582 99.5127
R2289 vdd.n2579 vdd.n2578 99.5127
R2290 vdd.n2575 vdd.n2574 99.5127
R2291 vdd.n2571 vdd.n2570 99.5127
R2292 vdd.n2567 vdd.n2566 99.5127
R2293 vdd.n2563 vdd.n2562 99.5127
R2294 vdd.n2559 vdd.n2558 99.5127
R2295 vdd.n2555 vdd.n2554 99.5127
R2296 vdd.n2551 vdd.n2550 99.5127
R2297 vdd.n2547 vdd.n2546 99.5127
R2298 vdd.n2543 vdd.n2542 99.5127
R2299 vdd.n2538 vdd.n2537 99.5127
R2300 vdd.n2276 vdd.n1050 99.5127
R2301 vdd.n2276 vdd.n1044 99.5127
R2302 vdd.n2273 vdd.n1044 99.5127
R2303 vdd.n2273 vdd.n1038 99.5127
R2304 vdd.n2270 vdd.n1038 99.5127
R2305 vdd.n2270 vdd.n1031 99.5127
R2306 vdd.n2267 vdd.n1031 99.5127
R2307 vdd.n2267 vdd.n1024 99.5127
R2308 vdd.n2264 vdd.n1024 99.5127
R2309 vdd.n2264 vdd.n1019 99.5127
R2310 vdd.n2261 vdd.n1019 99.5127
R2311 vdd.n2261 vdd.n1013 99.5127
R2312 vdd.n2258 vdd.n1013 99.5127
R2313 vdd.n2258 vdd.n1006 99.5127
R2314 vdd.n2172 vdd.n1006 99.5127
R2315 vdd.n2172 vdd.n1000 99.5127
R2316 vdd.n2169 vdd.n1000 99.5127
R2317 vdd.n2169 vdd.n995 99.5127
R2318 vdd.n2166 vdd.n995 99.5127
R2319 vdd.n2166 vdd.n990 99.5127
R2320 vdd.n2163 vdd.n990 99.5127
R2321 vdd.n2163 vdd.n984 99.5127
R2322 vdd.n2160 vdd.n984 99.5127
R2323 vdd.n2160 vdd.n977 99.5127
R2324 vdd.n2157 vdd.n977 99.5127
R2325 vdd.n2157 vdd.n970 99.5127
R2326 vdd.n970 vdd.n960 99.5127
R2327 vdd.n2533 vdd.n960 99.5127
R2328 vdd.n2111 vdd.n2109 99.5127
R2329 vdd.n2115 vdd.n2109 99.5127
R2330 vdd.n2119 vdd.n2117 99.5127
R2331 vdd.n2123 vdd.n2107 99.5127
R2332 vdd.n2127 vdd.n2125 99.5127
R2333 vdd.n2131 vdd.n2105 99.5127
R2334 vdd.n2135 vdd.n2133 99.5127
R2335 vdd.n2139 vdd.n2103 99.5127
R2336 vdd.n2142 vdd.n2141 99.5127
R2337 vdd.n2312 vdd.n2310 99.5127
R2338 vdd.n2308 vdd.n2144 99.5127
R2339 vdd.n2304 vdd.n2302 99.5127
R2340 vdd.n2300 vdd.n2146 99.5127
R2341 vdd.n2296 vdd.n2294 99.5127
R2342 vdd.n2292 vdd.n2148 99.5127
R2343 vdd.n2288 vdd.n2286 99.5127
R2344 vdd.n2284 vdd.n2150 99.5127
R2345 vdd.n2376 vdd.n1046 99.5127
R2346 vdd.n2380 vdd.n1046 99.5127
R2347 vdd.n2380 vdd.n1036 99.5127
R2348 vdd.n2388 vdd.n1036 99.5127
R2349 vdd.n2388 vdd.n1034 99.5127
R2350 vdd.n2392 vdd.n1034 99.5127
R2351 vdd.n2392 vdd.n1023 99.5127
R2352 vdd.n2401 vdd.n1023 99.5127
R2353 vdd.n2401 vdd.n1021 99.5127
R2354 vdd.n2405 vdd.n1021 99.5127
R2355 vdd.n2405 vdd.n1011 99.5127
R2356 vdd.n2413 vdd.n1011 99.5127
R2357 vdd.n2413 vdd.n1009 99.5127
R2358 vdd.n2417 vdd.n1009 99.5127
R2359 vdd.n2417 vdd.n999 99.5127
R2360 vdd.n2425 vdd.n999 99.5127
R2361 vdd.n2425 vdd.n997 99.5127
R2362 vdd.n2429 vdd.n997 99.5127
R2363 vdd.n2429 vdd.n988 99.5127
R2364 vdd.n2437 vdd.n988 99.5127
R2365 vdd.n2437 vdd.n986 99.5127
R2366 vdd.n2441 vdd.n986 99.5127
R2367 vdd.n2441 vdd.n975 99.5127
R2368 vdd.n2451 vdd.n975 99.5127
R2369 vdd.n2451 vdd.n972 99.5127
R2370 vdd.n2456 vdd.n972 99.5127
R2371 vdd.n2456 vdd.n973 99.5127
R2372 vdd.n973 vdd.n954 99.5127
R2373 vdd.n2974 vdd.n2973 99.5127
R2374 vdd.n2971 vdd.n2937 99.5127
R2375 vdd.n2967 vdd.n2966 99.5127
R2376 vdd.n2964 vdd.n2940 99.5127
R2377 vdd.n2960 vdd.n2959 99.5127
R2378 vdd.n2957 vdd.n2943 99.5127
R2379 vdd.n2953 vdd.n2952 99.5127
R2380 vdd.n2950 vdd.n2947 99.5127
R2381 vdd.n3091 vdd.n787 99.5127
R2382 vdd.n3089 vdd.n3088 99.5127
R2383 vdd.n3086 vdd.n789 99.5127
R2384 vdd.n3082 vdd.n3081 99.5127
R2385 vdd.n3079 vdd.n792 99.5127
R2386 vdd.n3075 vdd.n3074 99.5127
R2387 vdd.n3072 vdd.n795 99.5127
R2388 vdd.n3068 vdd.n3067 99.5127
R2389 vdd.n3065 vdd.n798 99.5127
R2390 vdd.n2709 vdd.n915 99.5127
R2391 vdd.n2709 vdd.n910 99.5127
R2392 vdd.n2780 vdd.n910 99.5127
R2393 vdd.n2780 vdd.n905 99.5127
R2394 vdd.n2776 vdd.n905 99.5127
R2395 vdd.n2776 vdd.n899 99.5127
R2396 vdd.n2773 vdd.n899 99.5127
R2397 vdd.n2773 vdd.n892 99.5127
R2398 vdd.n2770 vdd.n892 99.5127
R2399 vdd.n2770 vdd.n887 99.5127
R2400 vdd.n2767 vdd.n887 99.5127
R2401 vdd.n2767 vdd.n882 99.5127
R2402 vdd.n2764 vdd.n882 99.5127
R2403 vdd.n2764 vdd.n876 99.5127
R2404 vdd.n2761 vdd.n876 99.5127
R2405 vdd.n2761 vdd.n869 99.5127
R2406 vdd.n2726 vdd.n869 99.5127
R2407 vdd.n2726 vdd.n864 99.5127
R2408 vdd.n2723 vdd.n864 99.5127
R2409 vdd.n2723 vdd.n859 99.5127
R2410 vdd.n2720 vdd.n859 99.5127
R2411 vdd.n2720 vdd.n853 99.5127
R2412 vdd.n2717 vdd.n853 99.5127
R2413 vdd.n2717 vdd.n845 99.5127
R2414 vdd.n2714 vdd.n845 99.5127
R2415 vdd.n2714 vdd.n838 99.5127
R2416 vdd.n838 vdd.n804 99.5127
R2417 vdd.n3060 vdd.n804 99.5127
R2418 vdd.n2859 vdd.n918 99.5127
R2419 vdd.n2647 vdd.n2646 99.5127
R2420 vdd.n2651 vdd.n2650 99.5127
R2421 vdd.n2655 vdd.n2654 99.5127
R2422 vdd.n2659 vdd.n2658 99.5127
R2423 vdd.n2663 vdd.n2662 99.5127
R2424 vdd.n2667 vdd.n2666 99.5127
R2425 vdd.n2671 vdd.n2670 99.5127
R2426 vdd.n2675 vdd.n2674 99.5127
R2427 vdd.n2679 vdd.n2678 99.5127
R2428 vdd.n2683 vdd.n2682 99.5127
R2429 vdd.n2687 vdd.n2686 99.5127
R2430 vdd.n2691 vdd.n2690 99.5127
R2431 vdd.n2695 vdd.n2694 99.5127
R2432 vdd.n2699 vdd.n2698 99.5127
R2433 vdd.n2703 vdd.n2702 99.5127
R2434 vdd.n2705 vdd.n2637 99.5127
R2435 vdd.n2863 vdd.n908 99.5127
R2436 vdd.n2871 vdd.n908 99.5127
R2437 vdd.n2871 vdd.n906 99.5127
R2438 vdd.n2875 vdd.n906 99.5127
R2439 vdd.n2875 vdd.n896 99.5127
R2440 vdd.n2883 vdd.n896 99.5127
R2441 vdd.n2883 vdd.n894 99.5127
R2442 vdd.n2887 vdd.n894 99.5127
R2443 vdd.n2887 vdd.n885 99.5127
R2444 vdd.n2895 vdd.n885 99.5127
R2445 vdd.n2895 vdd.n883 99.5127
R2446 vdd.n2899 vdd.n883 99.5127
R2447 vdd.n2899 vdd.n873 99.5127
R2448 vdd.n2907 vdd.n873 99.5127
R2449 vdd.n2907 vdd.n871 99.5127
R2450 vdd.n2911 vdd.n871 99.5127
R2451 vdd.n2911 vdd.n862 99.5127
R2452 vdd.n2919 vdd.n862 99.5127
R2453 vdd.n2919 vdd.n860 99.5127
R2454 vdd.n2925 vdd.n860 99.5127
R2455 vdd.n2925 vdd.n850 99.5127
R2456 vdd.n2933 vdd.n850 99.5127
R2457 vdd.n2933 vdd.n847 99.5127
R2458 vdd.n2982 vdd.n847 99.5127
R2459 vdd.n2982 vdd.n848 99.5127
R2460 vdd.n848 vdd.n839 99.5127
R2461 vdd.n2977 vdd.n839 99.5127
R2462 vdd.n2977 vdd.n807 99.5127
R2463 vdd.n2527 vdd.n2526 99.5127
R2464 vdd.n2523 vdd.n2522 99.5127
R2465 vdd.n2519 vdd.n2518 99.5127
R2466 vdd.n2515 vdd.n2514 99.5127
R2467 vdd.n2511 vdd.n2510 99.5127
R2468 vdd.n2507 vdd.n2506 99.5127
R2469 vdd.n2503 vdd.n2502 99.5127
R2470 vdd.n2499 vdd.n2498 99.5127
R2471 vdd.n2495 vdd.n2494 99.5127
R2472 vdd.n2491 vdd.n2490 99.5127
R2473 vdd.n2487 vdd.n2486 99.5127
R2474 vdd.n2483 vdd.n2482 99.5127
R2475 vdd.n2479 vdd.n2478 99.5127
R2476 vdd.n2475 vdd.n2474 99.5127
R2477 vdd.n2471 vdd.n2470 99.5127
R2478 vdd.n2467 vdd.n2466 99.5127
R2479 vdd.n2463 vdd.n936 99.5127
R2480 vdd.n2220 vdd.n1051 99.5127
R2481 vdd.n2220 vdd.n1045 99.5127
R2482 vdd.n2223 vdd.n1045 99.5127
R2483 vdd.n2223 vdd.n1039 99.5127
R2484 vdd.n2226 vdd.n1039 99.5127
R2485 vdd.n2226 vdd.n1032 99.5127
R2486 vdd.n2229 vdd.n1032 99.5127
R2487 vdd.n2229 vdd.n1025 99.5127
R2488 vdd.n2232 vdd.n1025 99.5127
R2489 vdd.n2232 vdd.n1020 99.5127
R2490 vdd.n2235 vdd.n1020 99.5127
R2491 vdd.n2235 vdd.n1014 99.5127
R2492 vdd.n2256 vdd.n1014 99.5127
R2493 vdd.n2256 vdd.n1007 99.5127
R2494 vdd.n2252 vdd.n1007 99.5127
R2495 vdd.n2252 vdd.n1001 99.5127
R2496 vdd.n2249 vdd.n1001 99.5127
R2497 vdd.n2249 vdd.n996 99.5127
R2498 vdd.n2246 vdd.n996 99.5127
R2499 vdd.n2246 vdd.n991 99.5127
R2500 vdd.n2243 vdd.n991 99.5127
R2501 vdd.n2243 vdd.n985 99.5127
R2502 vdd.n2240 vdd.n985 99.5127
R2503 vdd.n2240 vdd.n978 99.5127
R2504 vdd.n978 vdd.n969 99.5127
R2505 vdd.n2458 vdd.n969 99.5127
R2506 vdd.n2459 vdd.n2458 99.5127
R2507 vdd.n2459 vdd.n961 99.5127
R2508 vdd.n2370 vdd.n2368 99.5127
R2509 vdd.n2366 vdd.n1054 99.5127
R2510 vdd.n2362 vdd.n2360 99.5127
R2511 vdd.n2358 vdd.n1056 99.5127
R2512 vdd.n2354 vdd.n2352 99.5127
R2513 vdd.n2350 vdd.n1058 99.5127
R2514 vdd.n2346 vdd.n2344 99.5127
R2515 vdd.n2342 vdd.n1060 99.5127
R2516 vdd.n2184 vdd.n1062 99.5127
R2517 vdd.n2189 vdd.n2186 99.5127
R2518 vdd.n2193 vdd.n2191 99.5127
R2519 vdd.n2197 vdd.n2182 99.5127
R2520 vdd.n2201 vdd.n2199 99.5127
R2521 vdd.n2205 vdd.n2180 99.5127
R2522 vdd.n2209 vdd.n2207 99.5127
R2523 vdd.n2214 vdd.n2176 99.5127
R2524 vdd.n2217 vdd.n2216 99.5127
R2525 vdd.n2374 vdd.n1042 99.5127
R2526 vdd.n2382 vdd.n1042 99.5127
R2527 vdd.n2382 vdd.n1040 99.5127
R2528 vdd.n2386 vdd.n1040 99.5127
R2529 vdd.n2386 vdd.n1029 99.5127
R2530 vdd.n2394 vdd.n1029 99.5127
R2531 vdd.n2394 vdd.n1026 99.5127
R2532 vdd.n2399 vdd.n1026 99.5127
R2533 vdd.n2399 vdd.n1017 99.5127
R2534 vdd.n2407 vdd.n1017 99.5127
R2535 vdd.n2407 vdd.n1015 99.5127
R2536 vdd.n2411 vdd.n1015 99.5127
R2537 vdd.n2411 vdd.n1005 99.5127
R2538 vdd.n2419 vdd.n1005 99.5127
R2539 vdd.n2419 vdd.n1003 99.5127
R2540 vdd.n2423 vdd.n1003 99.5127
R2541 vdd.n2423 vdd.n994 99.5127
R2542 vdd.n2431 vdd.n994 99.5127
R2543 vdd.n2431 vdd.n992 99.5127
R2544 vdd.n2435 vdd.n992 99.5127
R2545 vdd.n2435 vdd.n982 99.5127
R2546 vdd.n2443 vdd.n982 99.5127
R2547 vdd.n2443 vdd.n979 99.5127
R2548 vdd.n2449 vdd.n979 99.5127
R2549 vdd.n2449 vdd.n980 99.5127
R2550 vdd.n980 vdd.n971 99.5127
R2551 vdd.n971 vdd.n962 99.5127
R2552 vdd.n2531 vdd.n962 99.5127
R2553 vdd.n9 vdd.n7 98.9633
R2554 vdd.n2 vdd.n0 98.9633
R2555 vdd.n9 vdd.n8 98.6055
R2556 vdd.n11 vdd.n10 98.6055
R2557 vdd.n13 vdd.n12 98.6055
R2558 vdd.n6 vdd.n5 98.6055
R2559 vdd.n4 vdd.n3 98.6055
R2560 vdd.n2 vdd.n1 98.6055
R2561 vdd.t104 vdd.n303 85.8723
R2562 vdd.t23 vdd.n244 85.8723
R2563 vdd.t107 vdd.n201 85.8723
R2564 vdd.t46 vdd.n142 85.8723
R2565 vdd.t118 vdd.n100 85.8723
R2566 vdd.t35 vdd.n41 85.8723
R2567 vdd.t291 vdd.n1722 85.8723
R2568 vdd.t66 vdd.n1781 85.8723
R2569 vdd.t282 vdd.n1620 85.8723
R2570 vdd.t63 vdd.n1679 85.8723
R2571 vdd.t62 vdd.n1519 85.8723
R2572 vdd.t53 vdd.n1578 85.8723
R2573 vdd.n2923 vdd.n2922 78.546
R2574 vdd.n2397 vdd.n1027 78.546
R2575 vdd.n290 vdd.n289 75.1835
R2576 vdd.n288 vdd.n287 75.1835
R2577 vdd.n286 vdd.n285 75.1835
R2578 vdd.n284 vdd.n283 75.1835
R2579 vdd.n282 vdd.n281 75.1835
R2580 vdd.n280 vdd.n279 75.1835
R2581 vdd.n278 vdd.n277 75.1835
R2582 vdd.n276 vdd.n275 75.1835
R2583 vdd.n274 vdd.n273 75.1835
R2584 vdd.n188 vdd.n187 75.1835
R2585 vdd.n186 vdd.n185 75.1835
R2586 vdd.n184 vdd.n183 75.1835
R2587 vdd.n182 vdd.n181 75.1835
R2588 vdd.n180 vdd.n179 75.1835
R2589 vdd.n178 vdd.n177 75.1835
R2590 vdd.n176 vdd.n175 75.1835
R2591 vdd.n174 vdd.n173 75.1835
R2592 vdd.n172 vdd.n171 75.1835
R2593 vdd.n87 vdd.n86 75.1835
R2594 vdd.n85 vdd.n84 75.1835
R2595 vdd.n83 vdd.n82 75.1835
R2596 vdd.n81 vdd.n80 75.1835
R2597 vdd.n79 vdd.n78 75.1835
R2598 vdd.n77 vdd.n76 75.1835
R2599 vdd.n75 vdd.n74 75.1835
R2600 vdd.n73 vdd.n72 75.1835
R2601 vdd.n71 vdd.n70 75.1835
R2602 vdd.n1752 vdd.n1751 75.1835
R2603 vdd.n1754 vdd.n1753 75.1835
R2604 vdd.n1756 vdd.n1755 75.1835
R2605 vdd.n1758 vdd.n1757 75.1835
R2606 vdd.n1760 vdd.n1759 75.1835
R2607 vdd.n1762 vdd.n1761 75.1835
R2608 vdd.n1764 vdd.n1763 75.1835
R2609 vdd.n1766 vdd.n1765 75.1835
R2610 vdd.n1768 vdd.n1767 75.1835
R2611 vdd.n1650 vdd.n1649 75.1835
R2612 vdd.n1652 vdd.n1651 75.1835
R2613 vdd.n1654 vdd.n1653 75.1835
R2614 vdd.n1656 vdd.n1655 75.1835
R2615 vdd.n1658 vdd.n1657 75.1835
R2616 vdd.n1660 vdd.n1659 75.1835
R2617 vdd.n1662 vdd.n1661 75.1835
R2618 vdd.n1664 vdd.n1663 75.1835
R2619 vdd.n1666 vdd.n1665 75.1835
R2620 vdd.n1549 vdd.n1548 75.1835
R2621 vdd.n1551 vdd.n1550 75.1835
R2622 vdd.n1553 vdd.n1552 75.1835
R2623 vdd.n1555 vdd.n1554 75.1835
R2624 vdd.n1557 vdd.n1556 75.1835
R2625 vdd.n1559 vdd.n1558 75.1835
R2626 vdd.n1561 vdd.n1560 75.1835
R2627 vdd.n1563 vdd.n1562 75.1835
R2628 vdd.n1565 vdd.n1564 75.1835
R2629 vdd.n2858 vdd.n2857 72.8958
R2630 vdd.n2857 vdd.n2621 72.8958
R2631 vdd.n2857 vdd.n2622 72.8958
R2632 vdd.n2857 vdd.n2623 72.8958
R2633 vdd.n2857 vdd.n2624 72.8958
R2634 vdd.n2857 vdd.n2625 72.8958
R2635 vdd.n2857 vdd.n2626 72.8958
R2636 vdd.n2857 vdd.n2627 72.8958
R2637 vdd.n2857 vdd.n2628 72.8958
R2638 vdd.n2857 vdd.n2629 72.8958
R2639 vdd.n2857 vdd.n2630 72.8958
R2640 vdd.n2857 vdd.n2631 72.8958
R2641 vdd.n2857 vdd.n2632 72.8958
R2642 vdd.n2857 vdd.n2633 72.8958
R2643 vdd.n2857 vdd.n2634 72.8958
R2644 vdd.n2857 vdd.n2635 72.8958
R2645 vdd.n2857 vdd.n2636 72.8958
R2646 vdd.n803 vdd.n692 72.8958
R2647 vdd.n3066 vdd.n692 72.8958
R2648 vdd.n797 vdd.n692 72.8958
R2649 vdd.n3073 vdd.n692 72.8958
R2650 vdd.n794 vdd.n692 72.8958
R2651 vdd.n3080 vdd.n692 72.8958
R2652 vdd.n791 vdd.n692 72.8958
R2653 vdd.n3087 vdd.n692 72.8958
R2654 vdd.n3090 vdd.n692 72.8958
R2655 vdd.n2946 vdd.n692 72.8958
R2656 vdd.n2951 vdd.n692 72.8958
R2657 vdd.n2945 vdd.n692 72.8958
R2658 vdd.n2958 vdd.n692 72.8958
R2659 vdd.n2942 vdd.n692 72.8958
R2660 vdd.n2965 vdd.n692 72.8958
R2661 vdd.n2939 vdd.n692 72.8958
R2662 vdd.n2972 vdd.n692 72.8958
R2663 vdd.n2110 vdd.n1049 72.8958
R2664 vdd.n2116 vdd.n1049 72.8958
R2665 vdd.n2118 vdd.n1049 72.8958
R2666 vdd.n2124 vdd.n1049 72.8958
R2667 vdd.n2126 vdd.n1049 72.8958
R2668 vdd.n2132 vdd.n1049 72.8958
R2669 vdd.n2134 vdd.n1049 72.8958
R2670 vdd.n2140 vdd.n1049 72.8958
R2671 vdd.n2311 vdd.n1049 72.8958
R2672 vdd.n2309 vdd.n1049 72.8958
R2673 vdd.n2303 vdd.n1049 72.8958
R2674 vdd.n2301 vdd.n1049 72.8958
R2675 vdd.n2295 vdd.n1049 72.8958
R2676 vdd.n2293 vdd.n1049 72.8958
R2677 vdd.n2287 vdd.n1049 72.8958
R2678 vdd.n2285 vdd.n1049 72.8958
R2679 vdd.n2279 vdd.n1049 72.8958
R2680 vdd.n2604 vdd.n937 72.8958
R2681 vdd.n2604 vdd.n938 72.8958
R2682 vdd.n2604 vdd.n939 72.8958
R2683 vdd.n2604 vdd.n940 72.8958
R2684 vdd.n2604 vdd.n941 72.8958
R2685 vdd.n2604 vdd.n942 72.8958
R2686 vdd.n2604 vdd.n943 72.8958
R2687 vdd.n2604 vdd.n944 72.8958
R2688 vdd.n2604 vdd.n945 72.8958
R2689 vdd.n2604 vdd.n946 72.8958
R2690 vdd.n2604 vdd.n947 72.8958
R2691 vdd.n2604 vdd.n948 72.8958
R2692 vdd.n2604 vdd.n949 72.8958
R2693 vdd.n2604 vdd.n950 72.8958
R2694 vdd.n2604 vdd.n951 72.8958
R2695 vdd.n2604 vdd.n952 72.8958
R2696 vdd.n2604 vdd.n953 72.8958
R2697 vdd.n2857 vdd.n2856 72.8958
R2698 vdd.n2857 vdd.n2605 72.8958
R2699 vdd.n2857 vdd.n2606 72.8958
R2700 vdd.n2857 vdd.n2607 72.8958
R2701 vdd.n2857 vdd.n2608 72.8958
R2702 vdd.n2857 vdd.n2609 72.8958
R2703 vdd.n2857 vdd.n2610 72.8958
R2704 vdd.n2857 vdd.n2611 72.8958
R2705 vdd.n2857 vdd.n2612 72.8958
R2706 vdd.n2857 vdd.n2613 72.8958
R2707 vdd.n2857 vdd.n2614 72.8958
R2708 vdd.n2857 vdd.n2615 72.8958
R2709 vdd.n2857 vdd.n2616 72.8958
R2710 vdd.n2857 vdd.n2617 72.8958
R2711 vdd.n2857 vdd.n2618 72.8958
R2712 vdd.n2857 vdd.n2619 72.8958
R2713 vdd.n2857 vdd.n2620 72.8958
R2714 vdd.n2996 vdd.n692 72.8958
R2715 vdd.n835 vdd.n692 72.8958
R2716 vdd.n3004 vdd.n692 72.8958
R2717 vdd.n830 vdd.n692 72.8958
R2718 vdd.n3011 vdd.n692 72.8958
R2719 vdd.n827 vdd.n692 72.8958
R2720 vdd.n3018 vdd.n692 72.8958
R2721 vdd.n824 vdd.n692 72.8958
R2722 vdd.n3025 vdd.n692 72.8958
R2723 vdd.n3029 vdd.n692 72.8958
R2724 vdd.n821 vdd.n692 72.8958
R2725 vdd.n3036 vdd.n692 72.8958
R2726 vdd.n818 vdd.n692 72.8958
R2727 vdd.n3043 vdd.n692 72.8958
R2728 vdd.n815 vdd.n692 72.8958
R2729 vdd.n3050 vdd.n692 72.8958
R2730 vdd.n3053 vdd.n692 72.8958
R2731 vdd.n2604 vdd.n935 72.8958
R2732 vdd.n2604 vdd.n934 72.8958
R2733 vdd.n2604 vdd.n933 72.8958
R2734 vdd.n2604 vdd.n932 72.8958
R2735 vdd.n2604 vdd.n931 72.8958
R2736 vdd.n2604 vdd.n930 72.8958
R2737 vdd.n2604 vdd.n929 72.8958
R2738 vdd.n2604 vdd.n928 72.8958
R2739 vdd.n2604 vdd.n927 72.8958
R2740 vdd.n2604 vdd.n926 72.8958
R2741 vdd.n2604 vdd.n925 72.8958
R2742 vdd.n2604 vdd.n924 72.8958
R2743 vdd.n2604 vdd.n923 72.8958
R2744 vdd.n2604 vdd.n922 72.8958
R2745 vdd.n2604 vdd.n921 72.8958
R2746 vdd.n2604 vdd.n920 72.8958
R2747 vdd.n2604 vdd.n919 72.8958
R2748 vdd.n2369 vdd.n1049 72.8958
R2749 vdd.n2367 vdd.n1049 72.8958
R2750 vdd.n2361 vdd.n1049 72.8958
R2751 vdd.n2359 vdd.n1049 72.8958
R2752 vdd.n2353 vdd.n1049 72.8958
R2753 vdd.n2351 vdd.n1049 72.8958
R2754 vdd.n2345 vdd.n1049 72.8958
R2755 vdd.n2343 vdd.n1049 72.8958
R2756 vdd.n1061 vdd.n1049 72.8958
R2757 vdd.n2185 vdd.n1049 72.8958
R2758 vdd.n2190 vdd.n1049 72.8958
R2759 vdd.n2192 vdd.n1049 72.8958
R2760 vdd.n2198 vdd.n1049 72.8958
R2761 vdd.n2200 vdd.n1049 72.8958
R2762 vdd.n2206 vdd.n1049 72.8958
R2763 vdd.n2208 vdd.n1049 72.8958
R2764 vdd.n2215 vdd.n1049 72.8958
R2765 vdd.n1419 vdd.n1418 66.2847
R2766 vdd.n1418 vdd.n1194 66.2847
R2767 vdd.n1418 vdd.n1195 66.2847
R2768 vdd.n1418 vdd.n1196 66.2847
R2769 vdd.n1418 vdd.n1197 66.2847
R2770 vdd.n1418 vdd.n1198 66.2847
R2771 vdd.n1418 vdd.n1199 66.2847
R2772 vdd.n1418 vdd.n1200 66.2847
R2773 vdd.n1418 vdd.n1201 66.2847
R2774 vdd.n1418 vdd.n1202 66.2847
R2775 vdd.n1418 vdd.n1203 66.2847
R2776 vdd.n1418 vdd.n1204 66.2847
R2777 vdd.n1418 vdd.n1205 66.2847
R2778 vdd.n1418 vdd.n1206 66.2847
R2779 vdd.n1418 vdd.n1207 66.2847
R2780 vdd.n1418 vdd.n1208 66.2847
R2781 vdd.n1418 vdd.n1209 66.2847
R2782 vdd.n1418 vdd.n1210 66.2847
R2783 vdd.n1418 vdd.n1211 66.2847
R2784 vdd.n1418 vdd.n1212 66.2847
R2785 vdd.n1418 vdd.n1213 66.2847
R2786 vdd.n1418 vdd.n1214 66.2847
R2787 vdd.n1418 vdd.n1215 66.2847
R2788 vdd.n1418 vdd.n1216 66.2847
R2789 vdd.n1418 vdd.n1217 66.2847
R2790 vdd.n1418 vdd.n1218 66.2847
R2791 vdd.n1418 vdd.n1219 66.2847
R2792 vdd.n1418 vdd.n1220 66.2847
R2793 vdd.n1418 vdd.n1221 66.2847
R2794 vdd.n1418 vdd.n1222 66.2847
R2795 vdd.n1418 vdd.n1223 66.2847
R2796 vdd.n1073 vdd.n1070 66.2847
R2797 vdd.n2000 vdd.n1073 66.2847
R2798 vdd.n2005 vdd.n1073 66.2847
R2799 vdd.n2010 vdd.n1073 66.2847
R2800 vdd.n1998 vdd.n1073 66.2847
R2801 vdd.n2017 vdd.n1073 66.2847
R2802 vdd.n1990 vdd.n1073 66.2847
R2803 vdd.n2024 vdd.n1073 66.2847
R2804 vdd.n1983 vdd.n1073 66.2847
R2805 vdd.n2031 vdd.n1073 66.2847
R2806 vdd.n1977 vdd.n1073 66.2847
R2807 vdd.n1972 vdd.n1073 66.2847
R2808 vdd.n2042 vdd.n1073 66.2847
R2809 vdd.n1964 vdd.n1073 66.2847
R2810 vdd.n2049 vdd.n1073 66.2847
R2811 vdd.n1957 vdd.n1073 66.2847
R2812 vdd.n2056 vdd.n1073 66.2847
R2813 vdd.n1950 vdd.n1073 66.2847
R2814 vdd.n2063 vdd.n1073 66.2847
R2815 vdd.n1943 vdd.n1073 66.2847
R2816 vdd.n2070 vdd.n1073 66.2847
R2817 vdd.n1937 vdd.n1073 66.2847
R2818 vdd.n1932 vdd.n1073 66.2847
R2819 vdd.n2081 vdd.n1073 66.2847
R2820 vdd.n1924 vdd.n1073 66.2847
R2821 vdd.n2088 vdd.n1073 66.2847
R2822 vdd.n1917 vdd.n1073 66.2847
R2823 vdd.n2095 vdd.n1073 66.2847
R2824 vdd.n2098 vdd.n1073 66.2847
R2825 vdd.n1908 vdd.n1073 66.2847
R2826 vdd.n2320 vdd.n1073 66.2847
R2827 vdd.n1902 vdd.n1073 66.2847
R2828 vdd.n3223 vdd.n3222 66.2847
R2829 vdd.n3223 vdd.n693 66.2847
R2830 vdd.n3223 vdd.n694 66.2847
R2831 vdd.n3223 vdd.n695 66.2847
R2832 vdd.n3223 vdd.n696 66.2847
R2833 vdd.n3223 vdd.n697 66.2847
R2834 vdd.n3223 vdd.n698 66.2847
R2835 vdd.n3223 vdd.n699 66.2847
R2836 vdd.n3223 vdd.n700 66.2847
R2837 vdd.n3223 vdd.n701 66.2847
R2838 vdd.n3223 vdd.n702 66.2847
R2839 vdd.n3223 vdd.n703 66.2847
R2840 vdd.n3223 vdd.n704 66.2847
R2841 vdd.n3223 vdd.n705 66.2847
R2842 vdd.n3223 vdd.n706 66.2847
R2843 vdd.n3223 vdd.n707 66.2847
R2844 vdd.n3223 vdd.n708 66.2847
R2845 vdd.n3223 vdd.n709 66.2847
R2846 vdd.n3223 vdd.n710 66.2847
R2847 vdd.n3223 vdd.n711 66.2847
R2848 vdd.n3223 vdd.n712 66.2847
R2849 vdd.n3223 vdd.n713 66.2847
R2850 vdd.n3223 vdd.n714 66.2847
R2851 vdd.n3223 vdd.n715 66.2847
R2852 vdd.n3223 vdd.n716 66.2847
R2853 vdd.n3223 vdd.n717 66.2847
R2854 vdd.n3223 vdd.n718 66.2847
R2855 vdd.n3223 vdd.n719 66.2847
R2856 vdd.n3223 vdd.n720 66.2847
R2857 vdd.n3223 vdd.n721 66.2847
R2858 vdd.n3223 vdd.n722 66.2847
R2859 vdd.n3354 vdd.n3353 66.2847
R2860 vdd.n3354 vdd.n424 66.2847
R2861 vdd.n3354 vdd.n423 66.2847
R2862 vdd.n3354 vdd.n422 66.2847
R2863 vdd.n3354 vdd.n421 66.2847
R2864 vdd.n3354 vdd.n420 66.2847
R2865 vdd.n3354 vdd.n419 66.2847
R2866 vdd.n3354 vdd.n418 66.2847
R2867 vdd.n3354 vdd.n417 66.2847
R2868 vdd.n3354 vdd.n416 66.2847
R2869 vdd.n3354 vdd.n415 66.2847
R2870 vdd.n3354 vdd.n414 66.2847
R2871 vdd.n3354 vdd.n413 66.2847
R2872 vdd.n3354 vdd.n412 66.2847
R2873 vdd.n3354 vdd.n411 66.2847
R2874 vdd.n3354 vdd.n410 66.2847
R2875 vdd.n3354 vdd.n409 66.2847
R2876 vdd.n3354 vdd.n408 66.2847
R2877 vdd.n3354 vdd.n407 66.2847
R2878 vdd.n3354 vdd.n406 66.2847
R2879 vdd.n3354 vdd.n405 66.2847
R2880 vdd.n3354 vdd.n404 66.2847
R2881 vdd.n3354 vdd.n403 66.2847
R2882 vdd.n3354 vdd.n402 66.2847
R2883 vdd.n3354 vdd.n401 66.2847
R2884 vdd.n3354 vdd.n400 66.2847
R2885 vdd.n3354 vdd.n399 66.2847
R2886 vdd.n3354 vdd.n398 66.2847
R2887 vdd.n3354 vdd.n397 66.2847
R2888 vdd.n3354 vdd.n396 66.2847
R2889 vdd.n3354 vdd.n395 66.2847
R2890 vdd.n3354 vdd.n394 66.2847
R2891 vdd.n467 vdd.n394 52.4337
R2892 vdd.n473 vdd.n395 52.4337
R2893 vdd.n477 vdd.n396 52.4337
R2894 vdd.n483 vdd.n397 52.4337
R2895 vdd.n487 vdd.n398 52.4337
R2896 vdd.n493 vdd.n399 52.4337
R2897 vdd.n497 vdd.n400 52.4337
R2898 vdd.n503 vdd.n401 52.4337
R2899 vdd.n507 vdd.n402 52.4337
R2900 vdd.n513 vdd.n403 52.4337
R2901 vdd.n517 vdd.n404 52.4337
R2902 vdd.n523 vdd.n405 52.4337
R2903 vdd.n527 vdd.n406 52.4337
R2904 vdd.n533 vdd.n407 52.4337
R2905 vdd.n537 vdd.n408 52.4337
R2906 vdd.n543 vdd.n409 52.4337
R2907 vdd.n547 vdd.n410 52.4337
R2908 vdd.n553 vdd.n411 52.4337
R2909 vdd.n557 vdd.n412 52.4337
R2910 vdd.n563 vdd.n413 52.4337
R2911 vdd.n567 vdd.n414 52.4337
R2912 vdd.n573 vdd.n415 52.4337
R2913 vdd.n577 vdd.n416 52.4337
R2914 vdd.n583 vdd.n417 52.4337
R2915 vdd.n587 vdd.n418 52.4337
R2916 vdd.n593 vdd.n419 52.4337
R2917 vdd.n597 vdd.n420 52.4337
R2918 vdd.n603 vdd.n421 52.4337
R2919 vdd.n607 vdd.n422 52.4337
R2920 vdd.n613 vdd.n423 52.4337
R2921 vdd.n616 vdd.n424 52.4337
R2922 vdd.n3353 vdd.n3352 52.4337
R2923 vdd.n3222 vdd.n3221 52.4337
R2924 vdd.n728 vdd.n693 52.4337
R2925 vdd.n734 vdd.n694 52.4337
R2926 vdd.n3211 vdd.n695 52.4337
R2927 vdd.n3207 vdd.n696 52.4337
R2928 vdd.n3203 vdd.n697 52.4337
R2929 vdd.n3199 vdd.n698 52.4337
R2930 vdd.n3195 vdd.n699 52.4337
R2931 vdd.n3191 vdd.n700 52.4337
R2932 vdd.n3187 vdd.n701 52.4337
R2933 vdd.n3179 vdd.n702 52.4337
R2934 vdd.n3175 vdd.n703 52.4337
R2935 vdd.n3171 vdd.n704 52.4337
R2936 vdd.n3167 vdd.n705 52.4337
R2937 vdd.n3163 vdd.n706 52.4337
R2938 vdd.n3159 vdd.n707 52.4337
R2939 vdd.n3155 vdd.n708 52.4337
R2940 vdd.n3151 vdd.n709 52.4337
R2941 vdd.n3147 vdd.n710 52.4337
R2942 vdd.n3143 vdd.n711 52.4337
R2943 vdd.n3139 vdd.n712 52.4337
R2944 vdd.n3133 vdd.n713 52.4337
R2945 vdd.n3129 vdd.n714 52.4337
R2946 vdd.n3125 vdd.n715 52.4337
R2947 vdd.n3121 vdd.n716 52.4337
R2948 vdd.n3117 vdd.n717 52.4337
R2949 vdd.n3113 vdd.n718 52.4337
R2950 vdd.n3109 vdd.n719 52.4337
R2951 vdd.n3105 vdd.n720 52.4337
R2952 vdd.n3101 vdd.n721 52.4337
R2953 vdd.n3097 vdd.n722 52.4337
R2954 vdd.n2322 vdd.n1902 52.4337
R2955 vdd.n2320 vdd.n2319 52.4337
R2956 vdd.n1909 vdd.n1908 52.4337
R2957 vdd.n2098 vdd.n2097 52.4337
R2958 vdd.n2095 vdd.n2094 52.4337
R2959 vdd.n2090 vdd.n1917 52.4337
R2960 vdd.n2088 vdd.n2087 52.4337
R2961 vdd.n2083 vdd.n1924 52.4337
R2962 vdd.n2081 vdd.n2080 52.4337
R2963 vdd.n1933 vdd.n1932 52.4337
R2964 vdd.n2072 vdd.n1937 52.4337
R2965 vdd.n2070 vdd.n2069 52.4337
R2966 vdd.n2065 vdd.n1943 52.4337
R2967 vdd.n2063 vdd.n2062 52.4337
R2968 vdd.n2058 vdd.n1950 52.4337
R2969 vdd.n2056 vdd.n2055 52.4337
R2970 vdd.n2051 vdd.n1957 52.4337
R2971 vdd.n2049 vdd.n2048 52.4337
R2972 vdd.n2044 vdd.n1964 52.4337
R2973 vdd.n2042 vdd.n2041 52.4337
R2974 vdd.n1973 vdd.n1972 52.4337
R2975 vdd.n2033 vdd.n1977 52.4337
R2976 vdd.n2031 vdd.n2030 52.4337
R2977 vdd.n2026 vdd.n1983 52.4337
R2978 vdd.n2024 vdd.n2023 52.4337
R2979 vdd.n2019 vdd.n1990 52.4337
R2980 vdd.n2017 vdd.n2016 52.4337
R2981 vdd.n2012 vdd.n1998 52.4337
R2982 vdd.n2010 vdd.n2009 52.4337
R2983 vdd.n2005 vdd.n2004 52.4337
R2984 vdd.n2000 vdd.n1999 52.4337
R2985 vdd.n2331 vdd.n1070 52.4337
R2986 vdd.n1420 vdd.n1419 52.4337
R2987 vdd.n1226 vdd.n1194 52.4337
R2988 vdd.n1230 vdd.n1195 52.4337
R2989 vdd.n1232 vdd.n1196 52.4337
R2990 vdd.n1236 vdd.n1197 52.4337
R2991 vdd.n1238 vdd.n1198 52.4337
R2992 vdd.n1242 vdd.n1199 52.4337
R2993 vdd.n1244 vdd.n1200 52.4337
R2994 vdd.n1248 vdd.n1201 52.4337
R2995 vdd.n1250 vdd.n1202 52.4337
R2996 vdd.n1256 vdd.n1203 52.4337
R2997 vdd.n1258 vdd.n1204 52.4337
R2998 vdd.n1262 vdd.n1205 52.4337
R2999 vdd.n1264 vdd.n1206 52.4337
R3000 vdd.n1268 vdd.n1207 52.4337
R3001 vdd.n1270 vdd.n1208 52.4337
R3002 vdd.n1274 vdd.n1209 52.4337
R3003 vdd.n1276 vdd.n1210 52.4337
R3004 vdd.n1280 vdd.n1211 52.4337
R3005 vdd.n1282 vdd.n1212 52.4337
R3006 vdd.n1354 vdd.n1213 52.4337
R3007 vdd.n1287 vdd.n1214 52.4337
R3008 vdd.n1291 vdd.n1215 52.4337
R3009 vdd.n1293 vdd.n1216 52.4337
R3010 vdd.n1297 vdd.n1217 52.4337
R3011 vdd.n1299 vdd.n1218 52.4337
R3012 vdd.n1303 vdd.n1219 52.4337
R3013 vdd.n1305 vdd.n1220 52.4337
R3014 vdd.n1309 vdd.n1221 52.4337
R3015 vdd.n1311 vdd.n1222 52.4337
R3016 vdd.n1315 vdd.n1223 52.4337
R3017 vdd.n1419 vdd.n1193 52.4337
R3018 vdd.n1229 vdd.n1194 52.4337
R3019 vdd.n1231 vdd.n1195 52.4337
R3020 vdd.n1235 vdd.n1196 52.4337
R3021 vdd.n1237 vdd.n1197 52.4337
R3022 vdd.n1241 vdd.n1198 52.4337
R3023 vdd.n1243 vdd.n1199 52.4337
R3024 vdd.n1247 vdd.n1200 52.4337
R3025 vdd.n1249 vdd.n1201 52.4337
R3026 vdd.n1255 vdd.n1202 52.4337
R3027 vdd.n1257 vdd.n1203 52.4337
R3028 vdd.n1261 vdd.n1204 52.4337
R3029 vdd.n1263 vdd.n1205 52.4337
R3030 vdd.n1267 vdd.n1206 52.4337
R3031 vdd.n1269 vdd.n1207 52.4337
R3032 vdd.n1273 vdd.n1208 52.4337
R3033 vdd.n1275 vdd.n1209 52.4337
R3034 vdd.n1279 vdd.n1210 52.4337
R3035 vdd.n1281 vdd.n1211 52.4337
R3036 vdd.n1285 vdd.n1212 52.4337
R3037 vdd.n1286 vdd.n1213 52.4337
R3038 vdd.n1290 vdd.n1214 52.4337
R3039 vdd.n1292 vdd.n1215 52.4337
R3040 vdd.n1296 vdd.n1216 52.4337
R3041 vdd.n1298 vdd.n1217 52.4337
R3042 vdd.n1302 vdd.n1218 52.4337
R3043 vdd.n1304 vdd.n1219 52.4337
R3044 vdd.n1308 vdd.n1220 52.4337
R3045 vdd.n1310 vdd.n1221 52.4337
R3046 vdd.n1314 vdd.n1222 52.4337
R3047 vdd.n1316 vdd.n1223 52.4337
R3048 vdd.n1070 vdd.n1069 52.4337
R3049 vdd.n2001 vdd.n2000 52.4337
R3050 vdd.n2006 vdd.n2005 52.4337
R3051 vdd.n2011 vdd.n2010 52.4337
R3052 vdd.n1998 vdd.n1991 52.4337
R3053 vdd.n2018 vdd.n2017 52.4337
R3054 vdd.n1990 vdd.n1984 52.4337
R3055 vdd.n2025 vdd.n2024 52.4337
R3056 vdd.n1983 vdd.n1978 52.4337
R3057 vdd.n2032 vdd.n2031 52.4337
R3058 vdd.n1977 vdd.n1976 52.4337
R3059 vdd.n1972 vdd.n1965 52.4337
R3060 vdd.n2043 vdd.n2042 52.4337
R3061 vdd.n1964 vdd.n1958 52.4337
R3062 vdd.n2050 vdd.n2049 52.4337
R3063 vdd.n1957 vdd.n1951 52.4337
R3064 vdd.n2057 vdd.n2056 52.4337
R3065 vdd.n1950 vdd.n1944 52.4337
R3066 vdd.n2064 vdd.n2063 52.4337
R3067 vdd.n1943 vdd.n1938 52.4337
R3068 vdd.n2071 vdd.n2070 52.4337
R3069 vdd.n1937 vdd.n1936 52.4337
R3070 vdd.n1932 vdd.n1925 52.4337
R3071 vdd.n2082 vdd.n2081 52.4337
R3072 vdd.n1924 vdd.n1918 52.4337
R3073 vdd.n2089 vdd.n2088 52.4337
R3074 vdd.n1917 vdd.n1911 52.4337
R3075 vdd.n2096 vdd.n2095 52.4337
R3076 vdd.n2099 vdd.n2098 52.4337
R3077 vdd.n1908 vdd.n1903 52.4337
R3078 vdd.n2321 vdd.n2320 52.4337
R3079 vdd.n1902 vdd.n1075 52.4337
R3080 vdd.n3222 vdd.n725 52.4337
R3081 vdd.n733 vdd.n693 52.4337
R3082 vdd.n3212 vdd.n694 52.4337
R3083 vdd.n3208 vdd.n695 52.4337
R3084 vdd.n3204 vdd.n696 52.4337
R3085 vdd.n3200 vdd.n697 52.4337
R3086 vdd.n3196 vdd.n698 52.4337
R3087 vdd.n3192 vdd.n699 52.4337
R3088 vdd.n3188 vdd.n700 52.4337
R3089 vdd.n3178 vdd.n701 52.4337
R3090 vdd.n3176 vdd.n702 52.4337
R3091 vdd.n3172 vdd.n703 52.4337
R3092 vdd.n3168 vdd.n704 52.4337
R3093 vdd.n3164 vdd.n705 52.4337
R3094 vdd.n3160 vdd.n706 52.4337
R3095 vdd.n3156 vdd.n707 52.4337
R3096 vdd.n3152 vdd.n708 52.4337
R3097 vdd.n3148 vdd.n709 52.4337
R3098 vdd.n3144 vdd.n710 52.4337
R3099 vdd.n3140 vdd.n711 52.4337
R3100 vdd.n3132 vdd.n712 52.4337
R3101 vdd.n3130 vdd.n713 52.4337
R3102 vdd.n3126 vdd.n714 52.4337
R3103 vdd.n3122 vdd.n715 52.4337
R3104 vdd.n3118 vdd.n716 52.4337
R3105 vdd.n3114 vdd.n717 52.4337
R3106 vdd.n3110 vdd.n718 52.4337
R3107 vdd.n3106 vdd.n719 52.4337
R3108 vdd.n3102 vdd.n720 52.4337
R3109 vdd.n3098 vdd.n721 52.4337
R3110 vdd.n722 vdd.n691 52.4337
R3111 vdd.n3353 vdd.n425 52.4337
R3112 vdd.n614 vdd.n424 52.4337
R3113 vdd.n608 vdd.n423 52.4337
R3114 vdd.n604 vdd.n422 52.4337
R3115 vdd.n598 vdd.n421 52.4337
R3116 vdd.n594 vdd.n420 52.4337
R3117 vdd.n588 vdd.n419 52.4337
R3118 vdd.n584 vdd.n418 52.4337
R3119 vdd.n578 vdd.n417 52.4337
R3120 vdd.n574 vdd.n416 52.4337
R3121 vdd.n568 vdd.n415 52.4337
R3122 vdd.n564 vdd.n414 52.4337
R3123 vdd.n558 vdd.n413 52.4337
R3124 vdd.n554 vdd.n412 52.4337
R3125 vdd.n548 vdd.n411 52.4337
R3126 vdd.n544 vdd.n410 52.4337
R3127 vdd.n538 vdd.n409 52.4337
R3128 vdd.n534 vdd.n408 52.4337
R3129 vdd.n528 vdd.n407 52.4337
R3130 vdd.n524 vdd.n406 52.4337
R3131 vdd.n518 vdd.n405 52.4337
R3132 vdd.n514 vdd.n404 52.4337
R3133 vdd.n508 vdd.n403 52.4337
R3134 vdd.n504 vdd.n402 52.4337
R3135 vdd.n498 vdd.n401 52.4337
R3136 vdd.n494 vdd.n400 52.4337
R3137 vdd.n488 vdd.n399 52.4337
R3138 vdd.n484 vdd.n398 52.4337
R3139 vdd.n478 vdd.n397 52.4337
R3140 vdd.n474 vdd.n396 52.4337
R3141 vdd.n468 vdd.n395 52.4337
R3142 vdd.n394 vdd.n392 52.4337
R3143 vdd.t240 vdd.t253 51.4683
R3144 vdd.n274 vdd.n272 42.0461
R3145 vdd.n172 vdd.n170 42.0461
R3146 vdd.n71 vdd.n69 42.0461
R3147 vdd.n1752 vdd.n1750 42.0461
R3148 vdd.n1650 vdd.n1648 42.0461
R3149 vdd.n1549 vdd.n1547 42.0461
R3150 vdd.n332 vdd.n331 41.6884
R3151 vdd.n230 vdd.n229 41.6884
R3152 vdd.n129 vdd.n128 41.6884
R3153 vdd.n1810 vdd.n1809 41.6884
R3154 vdd.n1708 vdd.n1707 41.6884
R3155 vdd.n1607 vdd.n1606 41.6884
R3156 vdd.n1319 vdd.n1318 41.1157
R3157 vdd.n1357 vdd.n1356 41.1157
R3158 vdd.n1253 vdd.n1252 41.1157
R3159 vdd.n428 vdd.n427 41.1157
R3160 vdd.n566 vdd.n441 41.1157
R3161 vdd.n454 vdd.n453 41.1157
R3162 vdd.n3053 vdd.n3052 39.2114
R3163 vdd.n3050 vdd.n3049 39.2114
R3164 vdd.n3045 vdd.n815 39.2114
R3165 vdd.n3043 vdd.n3042 39.2114
R3166 vdd.n3038 vdd.n818 39.2114
R3167 vdd.n3036 vdd.n3035 39.2114
R3168 vdd.n3031 vdd.n821 39.2114
R3169 vdd.n3029 vdd.n3028 39.2114
R3170 vdd.n3025 vdd.n3024 39.2114
R3171 vdd.n3020 vdd.n824 39.2114
R3172 vdd.n3018 vdd.n3017 39.2114
R3173 vdd.n3013 vdd.n827 39.2114
R3174 vdd.n3011 vdd.n3010 39.2114
R3175 vdd.n3006 vdd.n830 39.2114
R3176 vdd.n3004 vdd.n3003 39.2114
R3177 vdd.n2998 vdd.n835 39.2114
R3178 vdd.n2996 vdd.n2995 39.2114
R3179 vdd.n2856 vdd.n913 39.2114
R3180 vdd.n2851 vdd.n2605 39.2114
R3181 vdd.n2848 vdd.n2606 39.2114
R3182 vdd.n2844 vdd.n2607 39.2114
R3183 vdd.n2840 vdd.n2608 39.2114
R3184 vdd.n2836 vdd.n2609 39.2114
R3185 vdd.n2832 vdd.n2610 39.2114
R3186 vdd.n2828 vdd.n2611 39.2114
R3187 vdd.n2824 vdd.n2612 39.2114
R3188 vdd.n2820 vdd.n2613 39.2114
R3189 vdd.n2816 vdd.n2614 39.2114
R3190 vdd.n2812 vdd.n2615 39.2114
R3191 vdd.n2808 vdd.n2616 39.2114
R3192 vdd.n2804 vdd.n2617 39.2114
R3193 vdd.n2800 vdd.n2618 39.2114
R3194 vdd.n2796 vdd.n2619 39.2114
R3195 vdd.n2791 vdd.n2620 39.2114
R3196 vdd.n2599 vdd.n953 39.2114
R3197 vdd.n2595 vdd.n952 39.2114
R3198 vdd.n2591 vdd.n951 39.2114
R3199 vdd.n2587 vdd.n950 39.2114
R3200 vdd.n2583 vdd.n949 39.2114
R3201 vdd.n2579 vdd.n948 39.2114
R3202 vdd.n2575 vdd.n947 39.2114
R3203 vdd.n2571 vdd.n946 39.2114
R3204 vdd.n2567 vdd.n945 39.2114
R3205 vdd.n2563 vdd.n944 39.2114
R3206 vdd.n2559 vdd.n943 39.2114
R3207 vdd.n2555 vdd.n942 39.2114
R3208 vdd.n2551 vdd.n941 39.2114
R3209 vdd.n2547 vdd.n940 39.2114
R3210 vdd.n2543 vdd.n939 39.2114
R3211 vdd.n2538 vdd.n938 39.2114
R3212 vdd.n2534 vdd.n937 39.2114
R3213 vdd.n2110 vdd.n1048 39.2114
R3214 vdd.n2116 vdd.n2115 39.2114
R3215 vdd.n2119 vdd.n2118 39.2114
R3216 vdd.n2124 vdd.n2123 39.2114
R3217 vdd.n2127 vdd.n2126 39.2114
R3218 vdd.n2132 vdd.n2131 39.2114
R3219 vdd.n2135 vdd.n2134 39.2114
R3220 vdd.n2140 vdd.n2139 39.2114
R3221 vdd.n2311 vdd.n2142 39.2114
R3222 vdd.n2310 vdd.n2309 39.2114
R3223 vdd.n2303 vdd.n2144 39.2114
R3224 vdd.n2302 vdd.n2301 39.2114
R3225 vdd.n2295 vdd.n2146 39.2114
R3226 vdd.n2294 vdd.n2293 39.2114
R3227 vdd.n2287 vdd.n2148 39.2114
R3228 vdd.n2286 vdd.n2285 39.2114
R3229 vdd.n2279 vdd.n2150 39.2114
R3230 vdd.n2972 vdd.n2971 39.2114
R3231 vdd.n2967 vdd.n2939 39.2114
R3232 vdd.n2965 vdd.n2964 39.2114
R3233 vdd.n2960 vdd.n2942 39.2114
R3234 vdd.n2958 vdd.n2957 39.2114
R3235 vdd.n2953 vdd.n2945 39.2114
R3236 vdd.n2951 vdd.n2950 39.2114
R3237 vdd.n2946 vdd.n787 39.2114
R3238 vdd.n3090 vdd.n3089 39.2114
R3239 vdd.n3087 vdd.n3086 39.2114
R3240 vdd.n3082 vdd.n791 39.2114
R3241 vdd.n3080 vdd.n3079 39.2114
R3242 vdd.n3075 vdd.n794 39.2114
R3243 vdd.n3073 vdd.n3072 39.2114
R3244 vdd.n3068 vdd.n797 39.2114
R3245 vdd.n3066 vdd.n3065 39.2114
R3246 vdd.n3061 vdd.n803 39.2114
R3247 vdd.n2858 vdd.n916 39.2114
R3248 vdd.n2621 vdd.n918 39.2114
R3249 vdd.n2647 vdd.n2622 39.2114
R3250 vdd.n2651 vdd.n2623 39.2114
R3251 vdd.n2655 vdd.n2624 39.2114
R3252 vdd.n2659 vdd.n2625 39.2114
R3253 vdd.n2663 vdd.n2626 39.2114
R3254 vdd.n2667 vdd.n2627 39.2114
R3255 vdd.n2671 vdd.n2628 39.2114
R3256 vdd.n2675 vdd.n2629 39.2114
R3257 vdd.n2679 vdd.n2630 39.2114
R3258 vdd.n2683 vdd.n2631 39.2114
R3259 vdd.n2687 vdd.n2632 39.2114
R3260 vdd.n2691 vdd.n2633 39.2114
R3261 vdd.n2695 vdd.n2634 39.2114
R3262 vdd.n2699 vdd.n2635 39.2114
R3263 vdd.n2703 vdd.n2636 39.2114
R3264 vdd.n2859 vdd.n2858 39.2114
R3265 vdd.n2646 vdd.n2621 39.2114
R3266 vdd.n2650 vdd.n2622 39.2114
R3267 vdd.n2654 vdd.n2623 39.2114
R3268 vdd.n2658 vdd.n2624 39.2114
R3269 vdd.n2662 vdd.n2625 39.2114
R3270 vdd.n2666 vdd.n2626 39.2114
R3271 vdd.n2670 vdd.n2627 39.2114
R3272 vdd.n2674 vdd.n2628 39.2114
R3273 vdd.n2678 vdd.n2629 39.2114
R3274 vdd.n2682 vdd.n2630 39.2114
R3275 vdd.n2686 vdd.n2631 39.2114
R3276 vdd.n2690 vdd.n2632 39.2114
R3277 vdd.n2694 vdd.n2633 39.2114
R3278 vdd.n2698 vdd.n2634 39.2114
R3279 vdd.n2702 vdd.n2635 39.2114
R3280 vdd.n2705 vdd.n2636 39.2114
R3281 vdd.n803 vdd.n798 39.2114
R3282 vdd.n3067 vdd.n3066 39.2114
R3283 vdd.n797 vdd.n795 39.2114
R3284 vdd.n3074 vdd.n3073 39.2114
R3285 vdd.n794 vdd.n792 39.2114
R3286 vdd.n3081 vdd.n3080 39.2114
R3287 vdd.n791 vdd.n789 39.2114
R3288 vdd.n3088 vdd.n3087 39.2114
R3289 vdd.n3091 vdd.n3090 39.2114
R3290 vdd.n2947 vdd.n2946 39.2114
R3291 vdd.n2952 vdd.n2951 39.2114
R3292 vdd.n2945 vdd.n2943 39.2114
R3293 vdd.n2959 vdd.n2958 39.2114
R3294 vdd.n2942 vdd.n2940 39.2114
R3295 vdd.n2966 vdd.n2965 39.2114
R3296 vdd.n2939 vdd.n2937 39.2114
R3297 vdd.n2973 vdd.n2972 39.2114
R3298 vdd.n2111 vdd.n2110 39.2114
R3299 vdd.n2117 vdd.n2116 39.2114
R3300 vdd.n2118 vdd.n2107 39.2114
R3301 vdd.n2125 vdd.n2124 39.2114
R3302 vdd.n2126 vdd.n2105 39.2114
R3303 vdd.n2133 vdd.n2132 39.2114
R3304 vdd.n2134 vdd.n2103 39.2114
R3305 vdd.n2141 vdd.n2140 39.2114
R3306 vdd.n2312 vdd.n2311 39.2114
R3307 vdd.n2309 vdd.n2308 39.2114
R3308 vdd.n2304 vdd.n2303 39.2114
R3309 vdd.n2301 vdd.n2300 39.2114
R3310 vdd.n2296 vdd.n2295 39.2114
R3311 vdd.n2293 vdd.n2292 39.2114
R3312 vdd.n2288 vdd.n2287 39.2114
R3313 vdd.n2285 vdd.n2284 39.2114
R3314 vdd.n2280 vdd.n2279 39.2114
R3315 vdd.n2537 vdd.n937 39.2114
R3316 vdd.n2542 vdd.n938 39.2114
R3317 vdd.n2546 vdd.n939 39.2114
R3318 vdd.n2550 vdd.n940 39.2114
R3319 vdd.n2554 vdd.n941 39.2114
R3320 vdd.n2558 vdd.n942 39.2114
R3321 vdd.n2562 vdd.n943 39.2114
R3322 vdd.n2566 vdd.n944 39.2114
R3323 vdd.n2570 vdd.n945 39.2114
R3324 vdd.n2574 vdd.n946 39.2114
R3325 vdd.n2578 vdd.n947 39.2114
R3326 vdd.n2582 vdd.n948 39.2114
R3327 vdd.n2586 vdd.n949 39.2114
R3328 vdd.n2590 vdd.n950 39.2114
R3329 vdd.n2594 vdd.n951 39.2114
R3330 vdd.n2598 vdd.n952 39.2114
R3331 vdd.n955 vdd.n953 39.2114
R3332 vdd.n2856 vdd.n2855 39.2114
R3333 vdd.n2849 vdd.n2605 39.2114
R3334 vdd.n2845 vdd.n2606 39.2114
R3335 vdd.n2841 vdd.n2607 39.2114
R3336 vdd.n2837 vdd.n2608 39.2114
R3337 vdd.n2833 vdd.n2609 39.2114
R3338 vdd.n2829 vdd.n2610 39.2114
R3339 vdd.n2825 vdd.n2611 39.2114
R3340 vdd.n2821 vdd.n2612 39.2114
R3341 vdd.n2817 vdd.n2613 39.2114
R3342 vdd.n2813 vdd.n2614 39.2114
R3343 vdd.n2809 vdd.n2615 39.2114
R3344 vdd.n2805 vdd.n2616 39.2114
R3345 vdd.n2801 vdd.n2617 39.2114
R3346 vdd.n2797 vdd.n2618 39.2114
R3347 vdd.n2792 vdd.n2619 39.2114
R3348 vdd.n2788 vdd.n2620 39.2114
R3349 vdd.n2997 vdd.n2996 39.2114
R3350 vdd.n835 vdd.n831 39.2114
R3351 vdd.n3005 vdd.n3004 39.2114
R3352 vdd.n830 vdd.n828 39.2114
R3353 vdd.n3012 vdd.n3011 39.2114
R3354 vdd.n827 vdd.n825 39.2114
R3355 vdd.n3019 vdd.n3018 39.2114
R3356 vdd.n824 vdd.n822 39.2114
R3357 vdd.n3026 vdd.n3025 39.2114
R3358 vdd.n3030 vdd.n3029 39.2114
R3359 vdd.n821 vdd.n819 39.2114
R3360 vdd.n3037 vdd.n3036 39.2114
R3361 vdd.n818 vdd.n816 39.2114
R3362 vdd.n3044 vdd.n3043 39.2114
R3363 vdd.n815 vdd.n813 39.2114
R3364 vdd.n3051 vdd.n3050 39.2114
R3365 vdd.n3054 vdd.n3053 39.2114
R3366 vdd.n963 vdd.n919 39.2114
R3367 vdd.n2526 vdd.n920 39.2114
R3368 vdd.n2522 vdd.n921 39.2114
R3369 vdd.n2518 vdd.n922 39.2114
R3370 vdd.n2514 vdd.n923 39.2114
R3371 vdd.n2510 vdd.n924 39.2114
R3372 vdd.n2506 vdd.n925 39.2114
R3373 vdd.n2502 vdd.n926 39.2114
R3374 vdd.n2498 vdd.n927 39.2114
R3375 vdd.n2494 vdd.n928 39.2114
R3376 vdd.n2490 vdd.n929 39.2114
R3377 vdd.n2486 vdd.n930 39.2114
R3378 vdd.n2482 vdd.n931 39.2114
R3379 vdd.n2478 vdd.n932 39.2114
R3380 vdd.n2474 vdd.n933 39.2114
R3381 vdd.n2470 vdd.n934 39.2114
R3382 vdd.n2466 vdd.n935 39.2114
R3383 vdd.n2369 vdd.n1052 39.2114
R3384 vdd.n2368 vdd.n2367 39.2114
R3385 vdd.n2361 vdd.n1054 39.2114
R3386 vdd.n2360 vdd.n2359 39.2114
R3387 vdd.n2353 vdd.n1056 39.2114
R3388 vdd.n2352 vdd.n2351 39.2114
R3389 vdd.n2345 vdd.n1058 39.2114
R3390 vdd.n2344 vdd.n2343 39.2114
R3391 vdd.n1061 vdd.n1060 39.2114
R3392 vdd.n2185 vdd.n2184 39.2114
R3393 vdd.n2190 vdd.n2189 39.2114
R3394 vdd.n2193 vdd.n2192 39.2114
R3395 vdd.n2198 vdd.n2197 39.2114
R3396 vdd.n2201 vdd.n2200 39.2114
R3397 vdd.n2206 vdd.n2205 39.2114
R3398 vdd.n2209 vdd.n2208 39.2114
R3399 vdd.n2215 vdd.n2214 39.2114
R3400 vdd.n2463 vdd.n935 39.2114
R3401 vdd.n2467 vdd.n934 39.2114
R3402 vdd.n2471 vdd.n933 39.2114
R3403 vdd.n2475 vdd.n932 39.2114
R3404 vdd.n2479 vdd.n931 39.2114
R3405 vdd.n2483 vdd.n930 39.2114
R3406 vdd.n2487 vdd.n929 39.2114
R3407 vdd.n2491 vdd.n928 39.2114
R3408 vdd.n2495 vdd.n927 39.2114
R3409 vdd.n2499 vdd.n926 39.2114
R3410 vdd.n2503 vdd.n925 39.2114
R3411 vdd.n2507 vdd.n924 39.2114
R3412 vdd.n2511 vdd.n923 39.2114
R3413 vdd.n2515 vdd.n922 39.2114
R3414 vdd.n2519 vdd.n921 39.2114
R3415 vdd.n2523 vdd.n920 39.2114
R3416 vdd.n2527 vdd.n919 39.2114
R3417 vdd.n2370 vdd.n2369 39.2114
R3418 vdd.n2367 vdd.n2366 39.2114
R3419 vdd.n2362 vdd.n2361 39.2114
R3420 vdd.n2359 vdd.n2358 39.2114
R3421 vdd.n2354 vdd.n2353 39.2114
R3422 vdd.n2351 vdd.n2350 39.2114
R3423 vdd.n2346 vdd.n2345 39.2114
R3424 vdd.n2343 vdd.n2342 39.2114
R3425 vdd.n1062 vdd.n1061 39.2114
R3426 vdd.n2186 vdd.n2185 39.2114
R3427 vdd.n2191 vdd.n2190 39.2114
R3428 vdd.n2192 vdd.n2182 39.2114
R3429 vdd.n2199 vdd.n2198 39.2114
R3430 vdd.n2200 vdd.n2180 39.2114
R3431 vdd.n2207 vdd.n2206 39.2114
R3432 vdd.n2208 vdd.n2176 39.2114
R3433 vdd.n2216 vdd.n2215 39.2114
R3434 vdd.n2335 vdd.n2334 37.2369
R3435 vdd.n2038 vdd.n1971 37.2369
R3436 vdd.n2077 vdd.n1931 37.2369
R3437 vdd.n3138 vdd.n769 37.2369
R3438 vdd.n3186 vdd.n3185 37.2369
R3439 vdd.n690 vdd.n689 37.2369
R3440 vdd.n2377 vdd.n1047 31.6883
R3441 vdd.n2602 vdd.n956 31.6883
R3442 vdd.n2535 vdd.n959 31.6883
R3443 vdd.n2281 vdd.n2278 31.6883
R3444 vdd.n2789 vdd.n2787 31.6883
R3445 vdd.n2994 vdd.n2993 31.6883
R3446 vdd.n2866 vdd.n912 31.6883
R3447 vdd.n3057 vdd.n3056 31.6883
R3448 vdd.n2976 vdd.n2975 31.6883
R3449 vdd.n3062 vdd.n802 31.6883
R3450 vdd.n2708 vdd.n2707 31.6883
R3451 vdd.n2862 vdd.n2861 31.6883
R3452 vdd.n2373 vdd.n2372 31.6883
R3453 vdd.n2530 vdd.n2529 31.6883
R3454 vdd.n2462 vdd.n2461 31.6883
R3455 vdd.n2219 vdd.n2218 31.6883
R3456 vdd.n2212 vdd.n2178 30.449
R3457 vdd.n967 vdd.n966 30.449
R3458 vdd.n2153 vdd.n2152 30.449
R3459 vdd.n2540 vdd.n958 30.449
R3460 vdd.n2644 vdd.n2643 30.449
R3461 vdd.n3000 vdd.n833 30.449
R3462 vdd.n2794 vdd.n2640 30.449
R3463 vdd.n801 vdd.n800 30.449
R3464 vdd.n1418 vdd.n1225 22.2201
R3465 vdd.n2329 vdd.n1073 22.2201
R3466 vdd.n3223 vdd.n723 22.2201
R3467 vdd.n3355 vdd.n3354 22.2201
R3468 vdd.n1429 vdd.n1187 19.3944
R3469 vdd.n1429 vdd.n1185 19.3944
R3470 vdd.n1433 vdd.n1185 19.3944
R3471 vdd.n1433 vdd.n1175 19.3944
R3472 vdd.n1446 vdd.n1175 19.3944
R3473 vdd.n1446 vdd.n1173 19.3944
R3474 vdd.n1450 vdd.n1173 19.3944
R3475 vdd.n1450 vdd.n1165 19.3944
R3476 vdd.n1463 vdd.n1165 19.3944
R3477 vdd.n1463 vdd.n1163 19.3944
R3478 vdd.n1467 vdd.n1163 19.3944
R3479 vdd.n1467 vdd.n1152 19.3944
R3480 vdd.n1479 vdd.n1152 19.3944
R3481 vdd.n1479 vdd.n1150 19.3944
R3482 vdd.n1483 vdd.n1150 19.3944
R3483 vdd.n1483 vdd.n1141 19.3944
R3484 vdd.n1496 vdd.n1141 19.3944
R3485 vdd.n1496 vdd.n1139 19.3944
R3486 vdd.n1500 vdd.n1139 19.3944
R3487 vdd.n1500 vdd.n1130 19.3944
R3488 vdd.n1819 vdd.n1130 19.3944
R3489 vdd.n1819 vdd.n1128 19.3944
R3490 vdd.n1823 vdd.n1128 19.3944
R3491 vdd.n1823 vdd.n1118 19.3944
R3492 vdd.n1836 vdd.n1118 19.3944
R3493 vdd.n1836 vdd.n1116 19.3944
R3494 vdd.n1840 vdd.n1116 19.3944
R3495 vdd.n1840 vdd.n1108 19.3944
R3496 vdd.n1853 vdd.n1108 19.3944
R3497 vdd.n1853 vdd.n1106 19.3944
R3498 vdd.n1857 vdd.n1106 19.3944
R3499 vdd.n1857 vdd.n1095 19.3944
R3500 vdd.n1869 vdd.n1095 19.3944
R3501 vdd.n1869 vdd.n1093 19.3944
R3502 vdd.n1873 vdd.n1093 19.3944
R3503 vdd.n1873 vdd.n1085 19.3944
R3504 vdd.n1886 vdd.n1085 19.3944
R3505 vdd.n1886 vdd.n1082 19.3944
R3506 vdd.n1892 vdd.n1082 19.3944
R3507 vdd.n1892 vdd.n1083 19.3944
R3508 vdd.n1083 vdd.n1072 19.3944
R3509 vdd.n1353 vdd.n1288 19.3944
R3510 vdd.n1349 vdd.n1288 19.3944
R3511 vdd.n1349 vdd.n1348 19.3944
R3512 vdd.n1348 vdd.n1347 19.3944
R3513 vdd.n1347 vdd.n1294 19.3944
R3514 vdd.n1343 vdd.n1294 19.3944
R3515 vdd.n1343 vdd.n1342 19.3944
R3516 vdd.n1342 vdd.n1341 19.3944
R3517 vdd.n1341 vdd.n1300 19.3944
R3518 vdd.n1337 vdd.n1300 19.3944
R3519 vdd.n1337 vdd.n1336 19.3944
R3520 vdd.n1336 vdd.n1335 19.3944
R3521 vdd.n1335 vdd.n1306 19.3944
R3522 vdd.n1331 vdd.n1306 19.3944
R3523 vdd.n1331 vdd.n1330 19.3944
R3524 vdd.n1330 vdd.n1329 19.3944
R3525 vdd.n1329 vdd.n1312 19.3944
R3526 vdd.n1325 vdd.n1312 19.3944
R3527 vdd.n1325 vdd.n1324 19.3944
R3528 vdd.n1324 vdd.n1323 19.3944
R3529 vdd.n1388 vdd.n1387 19.3944
R3530 vdd.n1387 vdd.n1386 19.3944
R3531 vdd.n1386 vdd.n1259 19.3944
R3532 vdd.n1382 vdd.n1259 19.3944
R3533 vdd.n1382 vdd.n1381 19.3944
R3534 vdd.n1381 vdd.n1380 19.3944
R3535 vdd.n1380 vdd.n1265 19.3944
R3536 vdd.n1376 vdd.n1265 19.3944
R3537 vdd.n1376 vdd.n1375 19.3944
R3538 vdd.n1375 vdd.n1374 19.3944
R3539 vdd.n1374 vdd.n1271 19.3944
R3540 vdd.n1370 vdd.n1271 19.3944
R3541 vdd.n1370 vdd.n1369 19.3944
R3542 vdd.n1369 vdd.n1368 19.3944
R3543 vdd.n1368 vdd.n1277 19.3944
R3544 vdd.n1364 vdd.n1277 19.3944
R3545 vdd.n1364 vdd.n1363 19.3944
R3546 vdd.n1363 vdd.n1362 19.3944
R3547 vdd.n1362 vdd.n1283 19.3944
R3548 vdd.n1358 vdd.n1283 19.3944
R3549 vdd.n1421 vdd.n1192 19.3944
R3550 vdd.n1416 vdd.n1192 19.3944
R3551 vdd.n1416 vdd.n1227 19.3944
R3552 vdd.n1412 vdd.n1227 19.3944
R3553 vdd.n1412 vdd.n1411 19.3944
R3554 vdd.n1411 vdd.n1410 19.3944
R3555 vdd.n1410 vdd.n1233 19.3944
R3556 vdd.n1406 vdd.n1233 19.3944
R3557 vdd.n1406 vdd.n1405 19.3944
R3558 vdd.n1405 vdd.n1404 19.3944
R3559 vdd.n1404 vdd.n1239 19.3944
R3560 vdd.n1400 vdd.n1239 19.3944
R3561 vdd.n1400 vdd.n1399 19.3944
R3562 vdd.n1399 vdd.n1398 19.3944
R3563 vdd.n1398 vdd.n1245 19.3944
R3564 vdd.n1394 vdd.n1245 19.3944
R3565 vdd.n1394 vdd.n1393 19.3944
R3566 vdd.n1393 vdd.n1392 19.3944
R3567 vdd.n2034 vdd.n1969 19.3944
R3568 vdd.n2034 vdd.n1975 19.3944
R3569 vdd.n2029 vdd.n1975 19.3944
R3570 vdd.n2029 vdd.n2028 19.3944
R3571 vdd.n2028 vdd.n2027 19.3944
R3572 vdd.n2027 vdd.n1982 19.3944
R3573 vdd.n2022 vdd.n1982 19.3944
R3574 vdd.n2022 vdd.n2021 19.3944
R3575 vdd.n2021 vdd.n2020 19.3944
R3576 vdd.n2020 vdd.n1989 19.3944
R3577 vdd.n2015 vdd.n1989 19.3944
R3578 vdd.n2015 vdd.n2014 19.3944
R3579 vdd.n2014 vdd.n2013 19.3944
R3580 vdd.n2013 vdd.n1997 19.3944
R3581 vdd.n2008 vdd.n1997 19.3944
R3582 vdd.n2008 vdd.n2007 19.3944
R3583 vdd.n2003 vdd.n2002 19.3944
R3584 vdd.n2336 vdd.n1068 19.3944
R3585 vdd.n2073 vdd.n1929 19.3944
R3586 vdd.n2073 vdd.n1935 19.3944
R3587 vdd.n2068 vdd.n1935 19.3944
R3588 vdd.n2068 vdd.n2067 19.3944
R3589 vdd.n2067 vdd.n2066 19.3944
R3590 vdd.n2066 vdd.n1942 19.3944
R3591 vdd.n2061 vdd.n1942 19.3944
R3592 vdd.n2061 vdd.n2060 19.3944
R3593 vdd.n2060 vdd.n2059 19.3944
R3594 vdd.n2059 vdd.n1949 19.3944
R3595 vdd.n2054 vdd.n1949 19.3944
R3596 vdd.n2054 vdd.n2053 19.3944
R3597 vdd.n2053 vdd.n2052 19.3944
R3598 vdd.n2052 vdd.n1956 19.3944
R3599 vdd.n2047 vdd.n1956 19.3944
R3600 vdd.n2047 vdd.n2046 19.3944
R3601 vdd.n2046 vdd.n2045 19.3944
R3602 vdd.n2045 vdd.n1963 19.3944
R3603 vdd.n2040 vdd.n1963 19.3944
R3604 vdd.n2040 vdd.n2039 19.3944
R3605 vdd.n2324 vdd.n2323 19.3944
R3606 vdd.n2323 vdd.n1901 19.3944
R3607 vdd.n2318 vdd.n2317 19.3944
R3608 vdd.n2100 vdd.n1905 19.3944
R3609 vdd.n2100 vdd.n1907 19.3944
R3610 vdd.n1910 vdd.n1907 19.3944
R3611 vdd.n2093 vdd.n1910 19.3944
R3612 vdd.n2093 vdd.n2092 19.3944
R3613 vdd.n2092 vdd.n2091 19.3944
R3614 vdd.n2091 vdd.n1916 19.3944
R3615 vdd.n2086 vdd.n1916 19.3944
R3616 vdd.n2086 vdd.n2085 19.3944
R3617 vdd.n2085 vdd.n2084 19.3944
R3618 vdd.n2084 vdd.n1923 19.3944
R3619 vdd.n2079 vdd.n1923 19.3944
R3620 vdd.n2079 vdd.n2078 19.3944
R3621 vdd.n1425 vdd.n1190 19.3944
R3622 vdd.n1425 vdd.n1181 19.3944
R3623 vdd.n1438 vdd.n1181 19.3944
R3624 vdd.n1438 vdd.n1179 19.3944
R3625 vdd.n1442 vdd.n1179 19.3944
R3626 vdd.n1442 vdd.n1170 19.3944
R3627 vdd.n1455 vdd.n1170 19.3944
R3628 vdd.n1455 vdd.n1168 19.3944
R3629 vdd.n1459 vdd.n1168 19.3944
R3630 vdd.n1459 vdd.n1159 19.3944
R3631 vdd.n1471 vdd.n1159 19.3944
R3632 vdd.n1471 vdd.n1157 19.3944
R3633 vdd.n1475 vdd.n1157 19.3944
R3634 vdd.n1475 vdd.n1147 19.3944
R3635 vdd.n1488 vdd.n1147 19.3944
R3636 vdd.n1488 vdd.n1145 19.3944
R3637 vdd.n1492 vdd.n1145 19.3944
R3638 vdd.n1492 vdd.n1136 19.3944
R3639 vdd.n1504 vdd.n1136 19.3944
R3640 vdd.n1504 vdd.n1134 19.3944
R3641 vdd.n1815 vdd.n1134 19.3944
R3642 vdd.n1815 vdd.n1124 19.3944
R3643 vdd.n1828 vdd.n1124 19.3944
R3644 vdd.n1828 vdd.n1122 19.3944
R3645 vdd.n1832 vdd.n1122 19.3944
R3646 vdd.n1832 vdd.n1113 19.3944
R3647 vdd.n1845 vdd.n1113 19.3944
R3648 vdd.n1845 vdd.n1111 19.3944
R3649 vdd.n1849 vdd.n1111 19.3944
R3650 vdd.n1849 vdd.n1102 19.3944
R3651 vdd.n1861 vdd.n1102 19.3944
R3652 vdd.n1861 vdd.n1100 19.3944
R3653 vdd.n1865 vdd.n1100 19.3944
R3654 vdd.n1865 vdd.n1090 19.3944
R3655 vdd.n1878 vdd.n1090 19.3944
R3656 vdd.n1878 vdd.n1088 19.3944
R3657 vdd.n1882 vdd.n1088 19.3944
R3658 vdd.n1882 vdd.n1078 19.3944
R3659 vdd.n1897 vdd.n1078 19.3944
R3660 vdd.n1897 vdd.n1076 19.3944
R3661 vdd.n2327 vdd.n1076 19.3944
R3662 vdd.n3229 vdd.n686 19.3944
R3663 vdd.n3229 vdd.n676 19.3944
R3664 vdd.n3241 vdd.n676 19.3944
R3665 vdd.n3241 vdd.n674 19.3944
R3666 vdd.n3245 vdd.n674 19.3944
R3667 vdd.n3245 vdd.n666 19.3944
R3668 vdd.n3258 vdd.n666 19.3944
R3669 vdd.n3258 vdd.n664 19.3944
R3670 vdd.n3262 vdd.n664 19.3944
R3671 vdd.n3262 vdd.n653 19.3944
R3672 vdd.n3274 vdd.n653 19.3944
R3673 vdd.n3274 vdd.n651 19.3944
R3674 vdd.n3278 vdd.n651 19.3944
R3675 vdd.n3278 vdd.n642 19.3944
R3676 vdd.n3291 vdd.n642 19.3944
R3677 vdd.n3291 vdd.n640 19.3944
R3678 vdd.n3298 vdd.n640 19.3944
R3679 vdd.n3298 vdd.n3297 19.3944
R3680 vdd.n3297 vdd.n631 19.3944
R3681 vdd.n3311 vdd.n631 19.3944
R3682 vdd.n3312 vdd.n3311 19.3944
R3683 vdd.n3312 vdd.n629 19.3944
R3684 vdd.n3316 vdd.n629 19.3944
R3685 vdd.n3318 vdd.n3316 19.3944
R3686 vdd.n3319 vdd.n3318 19.3944
R3687 vdd.n3319 vdd.n627 19.3944
R3688 vdd.n3323 vdd.n627 19.3944
R3689 vdd.n3325 vdd.n3323 19.3944
R3690 vdd.n3326 vdd.n3325 19.3944
R3691 vdd.n3326 vdd.n625 19.3944
R3692 vdd.n3330 vdd.n625 19.3944
R3693 vdd.n3333 vdd.n3330 19.3944
R3694 vdd.n3334 vdd.n3333 19.3944
R3695 vdd.n3334 vdd.n623 19.3944
R3696 vdd.n3338 vdd.n623 19.3944
R3697 vdd.n3340 vdd.n3338 19.3944
R3698 vdd.n3341 vdd.n3340 19.3944
R3699 vdd.n3341 vdd.n621 19.3944
R3700 vdd.n3345 vdd.n621 19.3944
R3701 vdd.n3347 vdd.n3345 19.3944
R3702 vdd.n3348 vdd.n3347 19.3944
R3703 vdd.n569 vdd.n438 19.3944
R3704 vdd.n575 vdd.n438 19.3944
R3705 vdd.n576 vdd.n575 19.3944
R3706 vdd.n579 vdd.n576 19.3944
R3707 vdd.n579 vdd.n436 19.3944
R3708 vdd.n585 vdd.n436 19.3944
R3709 vdd.n586 vdd.n585 19.3944
R3710 vdd.n589 vdd.n586 19.3944
R3711 vdd.n589 vdd.n434 19.3944
R3712 vdd.n595 vdd.n434 19.3944
R3713 vdd.n596 vdd.n595 19.3944
R3714 vdd.n599 vdd.n596 19.3944
R3715 vdd.n599 vdd.n432 19.3944
R3716 vdd.n605 vdd.n432 19.3944
R3717 vdd.n606 vdd.n605 19.3944
R3718 vdd.n609 vdd.n606 19.3944
R3719 vdd.n609 vdd.n430 19.3944
R3720 vdd.n615 vdd.n430 19.3944
R3721 vdd.n617 vdd.n615 19.3944
R3722 vdd.n618 vdd.n617 19.3944
R3723 vdd.n516 vdd.n515 19.3944
R3724 vdd.n519 vdd.n516 19.3944
R3725 vdd.n519 vdd.n450 19.3944
R3726 vdd.n525 vdd.n450 19.3944
R3727 vdd.n526 vdd.n525 19.3944
R3728 vdd.n529 vdd.n526 19.3944
R3729 vdd.n529 vdd.n448 19.3944
R3730 vdd.n535 vdd.n448 19.3944
R3731 vdd.n536 vdd.n535 19.3944
R3732 vdd.n539 vdd.n536 19.3944
R3733 vdd.n539 vdd.n446 19.3944
R3734 vdd.n545 vdd.n446 19.3944
R3735 vdd.n546 vdd.n545 19.3944
R3736 vdd.n549 vdd.n546 19.3944
R3737 vdd.n549 vdd.n444 19.3944
R3738 vdd.n555 vdd.n444 19.3944
R3739 vdd.n556 vdd.n555 19.3944
R3740 vdd.n559 vdd.n556 19.3944
R3741 vdd.n559 vdd.n442 19.3944
R3742 vdd.n565 vdd.n442 19.3944
R3743 vdd.n466 vdd.n465 19.3944
R3744 vdd.n469 vdd.n466 19.3944
R3745 vdd.n469 vdd.n462 19.3944
R3746 vdd.n475 vdd.n462 19.3944
R3747 vdd.n476 vdd.n475 19.3944
R3748 vdd.n479 vdd.n476 19.3944
R3749 vdd.n479 vdd.n460 19.3944
R3750 vdd.n485 vdd.n460 19.3944
R3751 vdd.n486 vdd.n485 19.3944
R3752 vdd.n489 vdd.n486 19.3944
R3753 vdd.n489 vdd.n458 19.3944
R3754 vdd.n495 vdd.n458 19.3944
R3755 vdd.n496 vdd.n495 19.3944
R3756 vdd.n499 vdd.n496 19.3944
R3757 vdd.n499 vdd.n456 19.3944
R3758 vdd.n505 vdd.n456 19.3944
R3759 vdd.n506 vdd.n505 19.3944
R3760 vdd.n509 vdd.n506 19.3944
R3761 vdd.n3233 vdd.n683 19.3944
R3762 vdd.n3233 vdd.n681 19.3944
R3763 vdd.n3237 vdd.n681 19.3944
R3764 vdd.n3237 vdd.n671 19.3944
R3765 vdd.n3250 vdd.n671 19.3944
R3766 vdd.n3250 vdd.n669 19.3944
R3767 vdd.n3254 vdd.n669 19.3944
R3768 vdd.n3254 vdd.n660 19.3944
R3769 vdd.n3266 vdd.n660 19.3944
R3770 vdd.n3266 vdd.n658 19.3944
R3771 vdd.n3270 vdd.n658 19.3944
R3772 vdd.n3270 vdd.n648 19.3944
R3773 vdd.n3283 vdd.n648 19.3944
R3774 vdd.n3283 vdd.n646 19.3944
R3775 vdd.n3287 vdd.n646 19.3944
R3776 vdd.n3287 vdd.n637 19.3944
R3777 vdd.n3302 vdd.n637 19.3944
R3778 vdd.n3302 vdd.n635 19.3944
R3779 vdd.n3306 vdd.n635 19.3944
R3780 vdd.n3306 vdd.n336 19.3944
R3781 vdd.n3397 vdd.n336 19.3944
R3782 vdd.n3397 vdd.n337 19.3944
R3783 vdd.n3391 vdd.n337 19.3944
R3784 vdd.n3391 vdd.n3390 19.3944
R3785 vdd.n3390 vdd.n3389 19.3944
R3786 vdd.n3389 vdd.n349 19.3944
R3787 vdd.n3383 vdd.n349 19.3944
R3788 vdd.n3383 vdd.n3382 19.3944
R3789 vdd.n3382 vdd.n3381 19.3944
R3790 vdd.n3381 vdd.n359 19.3944
R3791 vdd.n3375 vdd.n359 19.3944
R3792 vdd.n3375 vdd.n3374 19.3944
R3793 vdd.n3374 vdd.n3373 19.3944
R3794 vdd.n3373 vdd.n370 19.3944
R3795 vdd.n3367 vdd.n370 19.3944
R3796 vdd.n3367 vdd.n3366 19.3944
R3797 vdd.n3366 vdd.n3365 19.3944
R3798 vdd.n3365 vdd.n381 19.3944
R3799 vdd.n3359 vdd.n381 19.3944
R3800 vdd.n3359 vdd.n3358 19.3944
R3801 vdd.n3358 vdd.n3357 19.3944
R3802 vdd.n3180 vdd.n747 19.3944
R3803 vdd.n3180 vdd.n3177 19.3944
R3804 vdd.n3177 vdd.n3174 19.3944
R3805 vdd.n3174 vdd.n3173 19.3944
R3806 vdd.n3173 vdd.n3170 19.3944
R3807 vdd.n3170 vdd.n3169 19.3944
R3808 vdd.n3169 vdd.n3166 19.3944
R3809 vdd.n3166 vdd.n3165 19.3944
R3810 vdd.n3165 vdd.n3162 19.3944
R3811 vdd.n3162 vdd.n3161 19.3944
R3812 vdd.n3161 vdd.n3158 19.3944
R3813 vdd.n3158 vdd.n3157 19.3944
R3814 vdd.n3157 vdd.n3154 19.3944
R3815 vdd.n3154 vdd.n3153 19.3944
R3816 vdd.n3153 vdd.n3150 19.3944
R3817 vdd.n3150 vdd.n3149 19.3944
R3818 vdd.n3149 vdd.n3146 19.3944
R3819 vdd.n3146 vdd.n3145 19.3944
R3820 vdd.n3145 vdd.n3142 19.3944
R3821 vdd.n3142 vdd.n3141 19.3944
R3822 vdd.n3220 vdd.n3219 19.3944
R3823 vdd.n3219 vdd.n3218 19.3944
R3824 vdd.n732 vdd.n729 19.3944
R3825 vdd.n3214 vdd.n3213 19.3944
R3826 vdd.n3213 vdd.n3210 19.3944
R3827 vdd.n3210 vdd.n3209 19.3944
R3828 vdd.n3209 vdd.n3206 19.3944
R3829 vdd.n3206 vdd.n3205 19.3944
R3830 vdd.n3205 vdd.n3202 19.3944
R3831 vdd.n3202 vdd.n3201 19.3944
R3832 vdd.n3201 vdd.n3198 19.3944
R3833 vdd.n3198 vdd.n3197 19.3944
R3834 vdd.n3197 vdd.n3194 19.3944
R3835 vdd.n3194 vdd.n3193 19.3944
R3836 vdd.n3193 vdd.n3190 19.3944
R3837 vdd.n3190 vdd.n3189 19.3944
R3838 vdd.n3134 vdd.n767 19.3944
R3839 vdd.n3134 vdd.n3131 19.3944
R3840 vdd.n3131 vdd.n3128 19.3944
R3841 vdd.n3128 vdd.n3127 19.3944
R3842 vdd.n3127 vdd.n3124 19.3944
R3843 vdd.n3124 vdd.n3123 19.3944
R3844 vdd.n3123 vdd.n3120 19.3944
R3845 vdd.n3120 vdd.n3119 19.3944
R3846 vdd.n3119 vdd.n3116 19.3944
R3847 vdd.n3116 vdd.n3115 19.3944
R3848 vdd.n3115 vdd.n3112 19.3944
R3849 vdd.n3112 vdd.n3111 19.3944
R3850 vdd.n3111 vdd.n3108 19.3944
R3851 vdd.n3108 vdd.n3107 19.3944
R3852 vdd.n3107 vdd.n3104 19.3944
R3853 vdd.n3104 vdd.n3103 19.3944
R3854 vdd.n3100 vdd.n3099 19.3944
R3855 vdd.n3096 vdd.n3095 19.3944
R3856 vdd.n1357 vdd.n1353 19.0066
R3857 vdd.n2038 vdd.n1969 19.0066
R3858 vdd.n569 vdd.n566 19.0066
R3859 vdd.n3138 vdd.n767 19.0066
R3860 vdd.n2178 vdd.n2177 16.0975
R3861 vdd.n966 vdd.n965 16.0975
R3862 vdd.n1318 vdd.n1317 16.0975
R3863 vdd.n1356 vdd.n1355 16.0975
R3864 vdd.n1252 vdd.n1251 16.0975
R3865 vdd.n2334 vdd.n2333 16.0975
R3866 vdd.n1971 vdd.n1970 16.0975
R3867 vdd.n1931 vdd.n1930 16.0975
R3868 vdd.n2152 vdd.n2151 16.0975
R3869 vdd.n958 vdd.n957 16.0975
R3870 vdd.n2643 vdd.n2642 16.0975
R3871 vdd.n427 vdd.n426 16.0975
R3872 vdd.n441 vdd.n440 16.0975
R3873 vdd.n453 vdd.n452 16.0975
R3874 vdd.n769 vdd.n768 16.0975
R3875 vdd.n3185 vdd.n3184 16.0975
R3876 vdd.n833 vdd.n832 16.0975
R3877 vdd.n2640 vdd.n2639 16.0975
R3878 vdd.n689 vdd.n688 16.0975
R3879 vdd.n800 vdd.n799 16.0975
R3880 vdd.t253 vdd.n2604 15.4182
R3881 vdd.n2857 vdd.t240 15.4182
R3882 vdd.n28 vdd.n27 15.0023
R3883 vdd.n2375 vdd.n1049 14.5112
R3884 vdd.n3059 vdd.n692 14.5112
R3885 vdd.n328 vdd.n293 13.1884
R3886 vdd.n269 vdd.n234 13.1884
R3887 vdd.n226 vdd.n191 13.1884
R3888 vdd.n167 vdd.n132 13.1884
R3889 vdd.n125 vdd.n90 13.1884
R3890 vdd.n66 vdd.n31 13.1884
R3891 vdd.n1747 vdd.n1712 13.1884
R3892 vdd.n1806 vdd.n1771 13.1884
R3893 vdd.n1645 vdd.n1610 13.1884
R3894 vdd.n1704 vdd.n1669 13.1884
R3895 vdd.n1544 vdd.n1509 13.1884
R3896 vdd.n1603 vdd.n1568 13.1884
R3897 vdd.n1388 vdd.n1253 12.9944
R3898 vdd.n1392 vdd.n1253 12.9944
R3899 vdd.n2077 vdd.n1929 12.9944
R3900 vdd.n2078 vdd.n2077 12.9944
R3901 vdd.n515 vdd.n454 12.9944
R3902 vdd.n509 vdd.n454 12.9944
R3903 vdd.n3186 vdd.n747 12.9944
R3904 vdd.n3189 vdd.n3186 12.9944
R3905 vdd.n329 vdd.n291 12.8005
R3906 vdd.n324 vdd.n295 12.8005
R3907 vdd.n270 vdd.n232 12.8005
R3908 vdd.n265 vdd.n236 12.8005
R3909 vdd.n227 vdd.n189 12.8005
R3910 vdd.n222 vdd.n193 12.8005
R3911 vdd.n168 vdd.n130 12.8005
R3912 vdd.n163 vdd.n134 12.8005
R3913 vdd.n126 vdd.n88 12.8005
R3914 vdd.n121 vdd.n92 12.8005
R3915 vdd.n67 vdd.n29 12.8005
R3916 vdd.n62 vdd.n33 12.8005
R3917 vdd.n1748 vdd.n1710 12.8005
R3918 vdd.n1743 vdd.n1714 12.8005
R3919 vdd.n1807 vdd.n1769 12.8005
R3920 vdd.n1802 vdd.n1773 12.8005
R3921 vdd.n1646 vdd.n1608 12.8005
R3922 vdd.n1641 vdd.n1612 12.8005
R3923 vdd.n1705 vdd.n1667 12.8005
R3924 vdd.n1700 vdd.n1671 12.8005
R3925 vdd.n1545 vdd.n1507 12.8005
R3926 vdd.n1540 vdd.n1511 12.8005
R3927 vdd.n1604 vdd.n1566 12.8005
R3928 vdd.n1599 vdd.n1570 12.8005
R3929 vdd.n323 vdd.n296 12.0247
R3930 vdd.n264 vdd.n237 12.0247
R3931 vdd.n221 vdd.n194 12.0247
R3932 vdd.n162 vdd.n135 12.0247
R3933 vdd.n120 vdd.n93 12.0247
R3934 vdd.n61 vdd.n34 12.0247
R3935 vdd.n1742 vdd.n1715 12.0247
R3936 vdd.n1801 vdd.n1774 12.0247
R3937 vdd.n1640 vdd.n1613 12.0247
R3938 vdd.n1699 vdd.n1672 12.0247
R3939 vdd.n1539 vdd.n1512 12.0247
R3940 vdd.n1598 vdd.n1571 12.0247
R3941 vdd.n1427 vdd.n1183 11.337
R3942 vdd.n1436 vdd.n1183 11.337
R3943 vdd.n1436 vdd.n1435 11.337
R3944 vdd.n1444 vdd.n1177 11.337
R3945 vdd.n1453 vdd.n1452 11.337
R3946 vdd.n1469 vdd.n1161 11.337
R3947 vdd.n1477 vdd.n1154 11.337
R3948 vdd.n1486 vdd.n1485 11.337
R3949 vdd.n1494 vdd.n1143 11.337
R3950 vdd.n1817 vdd.n1132 11.337
R3951 vdd.n1826 vdd.n1126 11.337
R3952 vdd.n1834 vdd.n1120 11.337
R3953 vdd.n1843 vdd.n1842 11.337
R3954 vdd.n1859 vdd.n1104 11.337
R3955 vdd.n1867 vdd.n1097 11.337
R3956 vdd.n1876 vdd.n1875 11.337
R3957 vdd.n1884 vdd.n1080 11.337
R3958 vdd.n1895 vdd.n1080 11.337
R3959 vdd.n1895 vdd.n1894 11.337
R3960 vdd.n3231 vdd.n678 11.337
R3961 vdd.n3239 vdd.n678 11.337
R3962 vdd.n3239 vdd.n679 11.337
R3963 vdd.n3248 vdd.n3247 11.337
R3964 vdd.n3264 vdd.n662 11.337
R3965 vdd.n3272 vdd.n655 11.337
R3966 vdd.n3281 vdd.n3280 11.337
R3967 vdd.n3289 vdd.n644 11.337
R3968 vdd.n3308 vdd.n633 11.337
R3969 vdd.n3395 vdd.n340 11.337
R3970 vdd.n3393 vdd.n344 11.337
R3971 vdd.n3387 vdd.n3386 11.337
R3972 vdd.n3379 vdd.n361 11.337
R3973 vdd.n3378 vdd.n3377 11.337
R3974 vdd.n3371 vdd.n3370 11.337
R3975 vdd.n3369 vdd.n375 11.337
R3976 vdd.n3363 vdd.n3362 11.337
R3977 vdd.n3362 vdd.n3361 11.337
R3978 vdd.n3361 vdd.n386 11.337
R3979 vdd.n320 vdd.n319 11.249
R3980 vdd.n261 vdd.n260 11.249
R3981 vdd.n218 vdd.n217 11.249
R3982 vdd.n159 vdd.n158 11.249
R3983 vdd.n117 vdd.n116 11.249
R3984 vdd.n58 vdd.n57 11.249
R3985 vdd.n1739 vdd.n1738 11.249
R3986 vdd.n1798 vdd.n1797 11.249
R3987 vdd.n1637 vdd.n1636 11.249
R3988 vdd.n1696 vdd.n1695 11.249
R3989 vdd.n1536 vdd.n1535 11.249
R3990 vdd.n1595 vdd.n1594 11.249
R3991 vdd.n1225 vdd.t160 11.2237
R3992 vdd.n3355 vdd.t167 11.2237
R3993 vdd.n2532 vdd.t266 11.1103
R3994 vdd.n2864 vdd.t256 11.1103
R3995 vdd.t5 vdd.n1098 10.7702
R3996 vdd.n3256 vdd.t72 10.7702
R3997 vdd.n305 vdd.n304 10.7238
R3998 vdd.n246 vdd.n245 10.7238
R3999 vdd.n203 vdd.n202 10.7238
R4000 vdd.n144 vdd.n143 10.7238
R4001 vdd.n102 vdd.n101 10.7238
R4002 vdd.n43 vdd.n42 10.7238
R4003 vdd.n1724 vdd.n1723 10.7238
R4004 vdd.n1783 vdd.n1782 10.7238
R4005 vdd.n1622 vdd.n1621 10.7238
R4006 vdd.n1681 vdd.n1680 10.7238
R4007 vdd.n1521 vdd.n1520 10.7238
R4008 vdd.n1580 vdd.n1579 10.7238
R4009 vdd.n2378 vdd.n2377 10.6151
R4010 vdd.n2379 vdd.n2378 10.6151
R4011 vdd.n2379 vdd.n1035 10.6151
R4012 vdd.n2389 vdd.n1035 10.6151
R4013 vdd.n2390 vdd.n2389 10.6151
R4014 vdd.n2391 vdd.n2390 10.6151
R4015 vdd.n2391 vdd.n1022 10.6151
R4016 vdd.n2402 vdd.n1022 10.6151
R4017 vdd.n2403 vdd.n2402 10.6151
R4018 vdd.n2404 vdd.n2403 10.6151
R4019 vdd.n2404 vdd.n1010 10.6151
R4020 vdd.n2414 vdd.n1010 10.6151
R4021 vdd.n2415 vdd.n2414 10.6151
R4022 vdd.n2416 vdd.n2415 10.6151
R4023 vdd.n2416 vdd.n998 10.6151
R4024 vdd.n2426 vdd.n998 10.6151
R4025 vdd.n2427 vdd.n2426 10.6151
R4026 vdd.n2428 vdd.n2427 10.6151
R4027 vdd.n2428 vdd.n987 10.6151
R4028 vdd.n2438 vdd.n987 10.6151
R4029 vdd.n2439 vdd.n2438 10.6151
R4030 vdd.n2440 vdd.n2439 10.6151
R4031 vdd.n2440 vdd.n974 10.6151
R4032 vdd.n2452 vdd.n974 10.6151
R4033 vdd.n2453 vdd.n2452 10.6151
R4034 vdd.n2455 vdd.n2453 10.6151
R4035 vdd.n2455 vdd.n2454 10.6151
R4036 vdd.n2454 vdd.n956 10.6151
R4037 vdd.n2602 vdd.n2601 10.6151
R4038 vdd.n2601 vdd.n2600 10.6151
R4039 vdd.n2600 vdd.n2597 10.6151
R4040 vdd.n2597 vdd.n2596 10.6151
R4041 vdd.n2596 vdd.n2593 10.6151
R4042 vdd.n2593 vdd.n2592 10.6151
R4043 vdd.n2592 vdd.n2589 10.6151
R4044 vdd.n2589 vdd.n2588 10.6151
R4045 vdd.n2588 vdd.n2585 10.6151
R4046 vdd.n2585 vdd.n2584 10.6151
R4047 vdd.n2584 vdd.n2581 10.6151
R4048 vdd.n2581 vdd.n2580 10.6151
R4049 vdd.n2580 vdd.n2577 10.6151
R4050 vdd.n2577 vdd.n2576 10.6151
R4051 vdd.n2576 vdd.n2573 10.6151
R4052 vdd.n2573 vdd.n2572 10.6151
R4053 vdd.n2572 vdd.n2569 10.6151
R4054 vdd.n2569 vdd.n2568 10.6151
R4055 vdd.n2568 vdd.n2565 10.6151
R4056 vdd.n2565 vdd.n2564 10.6151
R4057 vdd.n2564 vdd.n2561 10.6151
R4058 vdd.n2561 vdd.n2560 10.6151
R4059 vdd.n2560 vdd.n2557 10.6151
R4060 vdd.n2557 vdd.n2556 10.6151
R4061 vdd.n2556 vdd.n2553 10.6151
R4062 vdd.n2553 vdd.n2552 10.6151
R4063 vdd.n2552 vdd.n2549 10.6151
R4064 vdd.n2549 vdd.n2548 10.6151
R4065 vdd.n2548 vdd.n2545 10.6151
R4066 vdd.n2545 vdd.n2544 10.6151
R4067 vdd.n2544 vdd.n2541 10.6151
R4068 vdd.n2539 vdd.n2536 10.6151
R4069 vdd.n2536 vdd.n2535 10.6151
R4070 vdd.n2278 vdd.n2277 10.6151
R4071 vdd.n2277 vdd.n2275 10.6151
R4072 vdd.n2275 vdd.n2274 10.6151
R4073 vdd.n2274 vdd.n2272 10.6151
R4074 vdd.n2272 vdd.n2271 10.6151
R4075 vdd.n2271 vdd.n2269 10.6151
R4076 vdd.n2269 vdd.n2268 10.6151
R4077 vdd.n2268 vdd.n2266 10.6151
R4078 vdd.n2266 vdd.n2265 10.6151
R4079 vdd.n2265 vdd.n2263 10.6151
R4080 vdd.n2263 vdd.n2262 10.6151
R4081 vdd.n2262 vdd.n2260 10.6151
R4082 vdd.n2260 vdd.n2259 10.6151
R4083 vdd.n2259 vdd.n2174 10.6151
R4084 vdd.n2174 vdd.n2173 10.6151
R4085 vdd.n2173 vdd.n2171 10.6151
R4086 vdd.n2171 vdd.n2170 10.6151
R4087 vdd.n2170 vdd.n2168 10.6151
R4088 vdd.n2168 vdd.n2167 10.6151
R4089 vdd.n2167 vdd.n2165 10.6151
R4090 vdd.n2165 vdd.n2164 10.6151
R4091 vdd.n2164 vdd.n2162 10.6151
R4092 vdd.n2162 vdd.n2161 10.6151
R4093 vdd.n2161 vdd.n2159 10.6151
R4094 vdd.n2159 vdd.n2158 10.6151
R4095 vdd.n2158 vdd.n2155 10.6151
R4096 vdd.n2155 vdd.n2154 10.6151
R4097 vdd.n2154 vdd.n959 10.6151
R4098 vdd.n2112 vdd.n1047 10.6151
R4099 vdd.n2113 vdd.n2112 10.6151
R4100 vdd.n2114 vdd.n2113 10.6151
R4101 vdd.n2114 vdd.n2108 10.6151
R4102 vdd.n2120 vdd.n2108 10.6151
R4103 vdd.n2121 vdd.n2120 10.6151
R4104 vdd.n2122 vdd.n2121 10.6151
R4105 vdd.n2122 vdd.n2106 10.6151
R4106 vdd.n2128 vdd.n2106 10.6151
R4107 vdd.n2129 vdd.n2128 10.6151
R4108 vdd.n2130 vdd.n2129 10.6151
R4109 vdd.n2130 vdd.n2104 10.6151
R4110 vdd.n2136 vdd.n2104 10.6151
R4111 vdd.n2137 vdd.n2136 10.6151
R4112 vdd.n2138 vdd.n2137 10.6151
R4113 vdd.n2138 vdd.n2102 10.6151
R4114 vdd.n2314 vdd.n2102 10.6151
R4115 vdd.n2314 vdd.n2313 10.6151
R4116 vdd.n2313 vdd.n2143 10.6151
R4117 vdd.n2307 vdd.n2143 10.6151
R4118 vdd.n2307 vdd.n2306 10.6151
R4119 vdd.n2306 vdd.n2305 10.6151
R4120 vdd.n2305 vdd.n2145 10.6151
R4121 vdd.n2299 vdd.n2145 10.6151
R4122 vdd.n2299 vdd.n2298 10.6151
R4123 vdd.n2298 vdd.n2297 10.6151
R4124 vdd.n2297 vdd.n2147 10.6151
R4125 vdd.n2291 vdd.n2147 10.6151
R4126 vdd.n2291 vdd.n2290 10.6151
R4127 vdd.n2290 vdd.n2289 10.6151
R4128 vdd.n2289 vdd.n2149 10.6151
R4129 vdd.n2283 vdd.n2282 10.6151
R4130 vdd.n2282 vdd.n2281 10.6151
R4131 vdd.n2787 vdd.n2786 10.6151
R4132 vdd.n2786 vdd.n2784 10.6151
R4133 vdd.n2784 vdd.n2783 10.6151
R4134 vdd.n2783 vdd.n2641 10.6151
R4135 vdd.n2730 vdd.n2641 10.6151
R4136 vdd.n2731 vdd.n2730 10.6151
R4137 vdd.n2733 vdd.n2731 10.6151
R4138 vdd.n2734 vdd.n2733 10.6151
R4139 vdd.n2736 vdd.n2734 10.6151
R4140 vdd.n2737 vdd.n2736 10.6151
R4141 vdd.n2739 vdd.n2737 10.6151
R4142 vdd.n2740 vdd.n2739 10.6151
R4143 vdd.n2742 vdd.n2740 10.6151
R4144 vdd.n2743 vdd.n2742 10.6151
R4145 vdd.n2758 vdd.n2743 10.6151
R4146 vdd.n2758 vdd.n2757 10.6151
R4147 vdd.n2757 vdd.n2756 10.6151
R4148 vdd.n2756 vdd.n2754 10.6151
R4149 vdd.n2754 vdd.n2753 10.6151
R4150 vdd.n2753 vdd.n2751 10.6151
R4151 vdd.n2751 vdd.n2750 10.6151
R4152 vdd.n2750 vdd.n2748 10.6151
R4153 vdd.n2748 vdd.n2747 10.6151
R4154 vdd.n2747 vdd.n2745 10.6151
R4155 vdd.n2745 vdd.n2744 10.6151
R4156 vdd.n2744 vdd.n836 10.6151
R4157 vdd.n2992 vdd.n836 10.6151
R4158 vdd.n2993 vdd.n2992 10.6151
R4159 vdd.n2854 vdd.n912 10.6151
R4160 vdd.n2854 vdd.n2853 10.6151
R4161 vdd.n2853 vdd.n2852 10.6151
R4162 vdd.n2852 vdd.n2850 10.6151
R4163 vdd.n2850 vdd.n2847 10.6151
R4164 vdd.n2847 vdd.n2846 10.6151
R4165 vdd.n2846 vdd.n2843 10.6151
R4166 vdd.n2843 vdd.n2842 10.6151
R4167 vdd.n2842 vdd.n2839 10.6151
R4168 vdd.n2839 vdd.n2838 10.6151
R4169 vdd.n2838 vdd.n2835 10.6151
R4170 vdd.n2835 vdd.n2834 10.6151
R4171 vdd.n2834 vdd.n2831 10.6151
R4172 vdd.n2831 vdd.n2830 10.6151
R4173 vdd.n2830 vdd.n2827 10.6151
R4174 vdd.n2827 vdd.n2826 10.6151
R4175 vdd.n2826 vdd.n2823 10.6151
R4176 vdd.n2823 vdd.n2822 10.6151
R4177 vdd.n2822 vdd.n2819 10.6151
R4178 vdd.n2819 vdd.n2818 10.6151
R4179 vdd.n2818 vdd.n2815 10.6151
R4180 vdd.n2815 vdd.n2814 10.6151
R4181 vdd.n2814 vdd.n2811 10.6151
R4182 vdd.n2811 vdd.n2810 10.6151
R4183 vdd.n2810 vdd.n2807 10.6151
R4184 vdd.n2807 vdd.n2806 10.6151
R4185 vdd.n2806 vdd.n2803 10.6151
R4186 vdd.n2803 vdd.n2802 10.6151
R4187 vdd.n2802 vdd.n2799 10.6151
R4188 vdd.n2799 vdd.n2798 10.6151
R4189 vdd.n2798 vdd.n2795 10.6151
R4190 vdd.n2793 vdd.n2790 10.6151
R4191 vdd.n2790 vdd.n2789 10.6151
R4192 vdd.n2867 vdd.n2866 10.6151
R4193 vdd.n2868 vdd.n2867 10.6151
R4194 vdd.n2868 vdd.n902 10.6151
R4195 vdd.n2878 vdd.n902 10.6151
R4196 vdd.n2879 vdd.n2878 10.6151
R4197 vdd.n2880 vdd.n2879 10.6151
R4198 vdd.n2880 vdd.n889 10.6151
R4199 vdd.n2890 vdd.n889 10.6151
R4200 vdd.n2891 vdd.n2890 10.6151
R4201 vdd.n2892 vdd.n2891 10.6151
R4202 vdd.n2892 vdd.n878 10.6151
R4203 vdd.n2902 vdd.n878 10.6151
R4204 vdd.n2903 vdd.n2902 10.6151
R4205 vdd.n2904 vdd.n2903 10.6151
R4206 vdd.n2904 vdd.n866 10.6151
R4207 vdd.n2914 vdd.n866 10.6151
R4208 vdd.n2915 vdd.n2914 10.6151
R4209 vdd.n2916 vdd.n2915 10.6151
R4210 vdd.n2916 vdd.n855 10.6151
R4211 vdd.n2928 vdd.n855 10.6151
R4212 vdd.n2929 vdd.n2928 10.6151
R4213 vdd.n2930 vdd.n2929 10.6151
R4214 vdd.n2930 vdd.n841 10.6151
R4215 vdd.n2985 vdd.n841 10.6151
R4216 vdd.n2986 vdd.n2985 10.6151
R4217 vdd.n2987 vdd.n2986 10.6151
R4218 vdd.n2987 vdd.n810 10.6151
R4219 vdd.n3057 vdd.n810 10.6151
R4220 vdd.n3056 vdd.n3055 10.6151
R4221 vdd.n3055 vdd.n811 10.6151
R4222 vdd.n812 vdd.n811 10.6151
R4223 vdd.n3048 vdd.n812 10.6151
R4224 vdd.n3048 vdd.n3047 10.6151
R4225 vdd.n3047 vdd.n3046 10.6151
R4226 vdd.n3046 vdd.n814 10.6151
R4227 vdd.n3041 vdd.n814 10.6151
R4228 vdd.n3041 vdd.n3040 10.6151
R4229 vdd.n3040 vdd.n3039 10.6151
R4230 vdd.n3039 vdd.n817 10.6151
R4231 vdd.n3034 vdd.n817 10.6151
R4232 vdd.n3034 vdd.n3033 10.6151
R4233 vdd.n3033 vdd.n3032 10.6151
R4234 vdd.n3032 vdd.n820 10.6151
R4235 vdd.n3027 vdd.n820 10.6151
R4236 vdd.n3027 vdd.n731 10.6151
R4237 vdd.n3023 vdd.n731 10.6151
R4238 vdd.n3023 vdd.n3022 10.6151
R4239 vdd.n3022 vdd.n3021 10.6151
R4240 vdd.n3021 vdd.n823 10.6151
R4241 vdd.n3016 vdd.n823 10.6151
R4242 vdd.n3016 vdd.n3015 10.6151
R4243 vdd.n3015 vdd.n3014 10.6151
R4244 vdd.n3014 vdd.n826 10.6151
R4245 vdd.n3009 vdd.n826 10.6151
R4246 vdd.n3009 vdd.n3008 10.6151
R4247 vdd.n3008 vdd.n3007 10.6151
R4248 vdd.n3007 vdd.n829 10.6151
R4249 vdd.n3002 vdd.n829 10.6151
R4250 vdd.n3002 vdd.n3001 10.6151
R4251 vdd.n2999 vdd.n834 10.6151
R4252 vdd.n2994 vdd.n834 10.6151
R4253 vdd.n2975 vdd.n2936 10.6151
R4254 vdd.n2970 vdd.n2936 10.6151
R4255 vdd.n2970 vdd.n2969 10.6151
R4256 vdd.n2969 vdd.n2968 10.6151
R4257 vdd.n2968 vdd.n2938 10.6151
R4258 vdd.n2963 vdd.n2938 10.6151
R4259 vdd.n2963 vdd.n2962 10.6151
R4260 vdd.n2962 vdd.n2961 10.6151
R4261 vdd.n2961 vdd.n2941 10.6151
R4262 vdd.n2956 vdd.n2941 10.6151
R4263 vdd.n2956 vdd.n2955 10.6151
R4264 vdd.n2955 vdd.n2954 10.6151
R4265 vdd.n2954 vdd.n2944 10.6151
R4266 vdd.n2949 vdd.n2944 10.6151
R4267 vdd.n2949 vdd.n2948 10.6151
R4268 vdd.n2948 vdd.n785 10.6151
R4269 vdd.n3092 vdd.n785 10.6151
R4270 vdd.n3092 vdd.n786 10.6151
R4271 vdd.n788 vdd.n786 10.6151
R4272 vdd.n3085 vdd.n788 10.6151
R4273 vdd.n3085 vdd.n3084 10.6151
R4274 vdd.n3084 vdd.n3083 10.6151
R4275 vdd.n3083 vdd.n790 10.6151
R4276 vdd.n3078 vdd.n790 10.6151
R4277 vdd.n3078 vdd.n3077 10.6151
R4278 vdd.n3077 vdd.n3076 10.6151
R4279 vdd.n3076 vdd.n793 10.6151
R4280 vdd.n3071 vdd.n793 10.6151
R4281 vdd.n3071 vdd.n3070 10.6151
R4282 vdd.n3070 vdd.n3069 10.6151
R4283 vdd.n3069 vdd.n796 10.6151
R4284 vdd.n3064 vdd.n3063 10.6151
R4285 vdd.n3063 vdd.n3062 10.6151
R4286 vdd.n2710 vdd.n2708 10.6151
R4287 vdd.n2711 vdd.n2710 10.6151
R4288 vdd.n2779 vdd.n2711 10.6151
R4289 vdd.n2779 vdd.n2778 10.6151
R4290 vdd.n2778 vdd.n2777 10.6151
R4291 vdd.n2777 vdd.n2775 10.6151
R4292 vdd.n2775 vdd.n2774 10.6151
R4293 vdd.n2774 vdd.n2772 10.6151
R4294 vdd.n2772 vdd.n2771 10.6151
R4295 vdd.n2771 vdd.n2769 10.6151
R4296 vdd.n2769 vdd.n2768 10.6151
R4297 vdd.n2768 vdd.n2766 10.6151
R4298 vdd.n2766 vdd.n2765 10.6151
R4299 vdd.n2765 vdd.n2763 10.6151
R4300 vdd.n2763 vdd.n2762 10.6151
R4301 vdd.n2762 vdd.n2728 10.6151
R4302 vdd.n2728 vdd.n2727 10.6151
R4303 vdd.n2727 vdd.n2725 10.6151
R4304 vdd.n2725 vdd.n2724 10.6151
R4305 vdd.n2724 vdd.n2722 10.6151
R4306 vdd.n2722 vdd.n2721 10.6151
R4307 vdd.n2721 vdd.n2719 10.6151
R4308 vdd.n2719 vdd.n2718 10.6151
R4309 vdd.n2718 vdd.n2716 10.6151
R4310 vdd.n2716 vdd.n2715 10.6151
R4311 vdd.n2715 vdd.n2713 10.6151
R4312 vdd.n2713 vdd.n2712 10.6151
R4313 vdd.n2712 vdd.n802 10.6151
R4314 vdd.n2861 vdd.n2860 10.6151
R4315 vdd.n2860 vdd.n917 10.6151
R4316 vdd.n2645 vdd.n917 10.6151
R4317 vdd.n2648 vdd.n2645 10.6151
R4318 vdd.n2649 vdd.n2648 10.6151
R4319 vdd.n2652 vdd.n2649 10.6151
R4320 vdd.n2653 vdd.n2652 10.6151
R4321 vdd.n2656 vdd.n2653 10.6151
R4322 vdd.n2657 vdd.n2656 10.6151
R4323 vdd.n2660 vdd.n2657 10.6151
R4324 vdd.n2661 vdd.n2660 10.6151
R4325 vdd.n2664 vdd.n2661 10.6151
R4326 vdd.n2665 vdd.n2664 10.6151
R4327 vdd.n2668 vdd.n2665 10.6151
R4328 vdd.n2669 vdd.n2668 10.6151
R4329 vdd.n2672 vdd.n2669 10.6151
R4330 vdd.n2673 vdd.n2672 10.6151
R4331 vdd.n2676 vdd.n2673 10.6151
R4332 vdd.n2677 vdd.n2676 10.6151
R4333 vdd.n2680 vdd.n2677 10.6151
R4334 vdd.n2681 vdd.n2680 10.6151
R4335 vdd.n2684 vdd.n2681 10.6151
R4336 vdd.n2685 vdd.n2684 10.6151
R4337 vdd.n2688 vdd.n2685 10.6151
R4338 vdd.n2689 vdd.n2688 10.6151
R4339 vdd.n2692 vdd.n2689 10.6151
R4340 vdd.n2693 vdd.n2692 10.6151
R4341 vdd.n2696 vdd.n2693 10.6151
R4342 vdd.n2697 vdd.n2696 10.6151
R4343 vdd.n2700 vdd.n2697 10.6151
R4344 vdd.n2701 vdd.n2700 10.6151
R4345 vdd.n2706 vdd.n2704 10.6151
R4346 vdd.n2707 vdd.n2706 10.6151
R4347 vdd.n2862 vdd.n907 10.6151
R4348 vdd.n2872 vdd.n907 10.6151
R4349 vdd.n2873 vdd.n2872 10.6151
R4350 vdd.n2874 vdd.n2873 10.6151
R4351 vdd.n2874 vdd.n895 10.6151
R4352 vdd.n2884 vdd.n895 10.6151
R4353 vdd.n2885 vdd.n2884 10.6151
R4354 vdd.n2886 vdd.n2885 10.6151
R4355 vdd.n2886 vdd.n884 10.6151
R4356 vdd.n2896 vdd.n884 10.6151
R4357 vdd.n2897 vdd.n2896 10.6151
R4358 vdd.n2898 vdd.n2897 10.6151
R4359 vdd.n2898 vdd.n872 10.6151
R4360 vdd.n2908 vdd.n872 10.6151
R4361 vdd.n2909 vdd.n2908 10.6151
R4362 vdd.n2910 vdd.n2909 10.6151
R4363 vdd.n2910 vdd.n861 10.6151
R4364 vdd.n2920 vdd.n861 10.6151
R4365 vdd.n2921 vdd.n2920 10.6151
R4366 vdd.n2924 vdd.n2921 10.6151
R4367 vdd.n2934 vdd.n849 10.6151
R4368 vdd.n2935 vdd.n2934 10.6151
R4369 vdd.n2981 vdd.n2935 10.6151
R4370 vdd.n2981 vdd.n2980 10.6151
R4371 vdd.n2980 vdd.n2979 10.6151
R4372 vdd.n2979 vdd.n2978 10.6151
R4373 vdd.n2978 vdd.n2976 10.6151
R4374 vdd.n2373 vdd.n1041 10.6151
R4375 vdd.n2383 vdd.n1041 10.6151
R4376 vdd.n2384 vdd.n2383 10.6151
R4377 vdd.n2385 vdd.n2384 10.6151
R4378 vdd.n2385 vdd.n1028 10.6151
R4379 vdd.n2395 vdd.n1028 10.6151
R4380 vdd.n2396 vdd.n2395 10.6151
R4381 vdd.n2398 vdd.n1016 10.6151
R4382 vdd.n2408 vdd.n1016 10.6151
R4383 vdd.n2409 vdd.n2408 10.6151
R4384 vdd.n2410 vdd.n2409 10.6151
R4385 vdd.n2410 vdd.n1004 10.6151
R4386 vdd.n2420 vdd.n1004 10.6151
R4387 vdd.n2421 vdd.n2420 10.6151
R4388 vdd.n2422 vdd.n2421 10.6151
R4389 vdd.n2422 vdd.n993 10.6151
R4390 vdd.n2432 vdd.n993 10.6151
R4391 vdd.n2433 vdd.n2432 10.6151
R4392 vdd.n2434 vdd.n2433 10.6151
R4393 vdd.n2434 vdd.n981 10.6151
R4394 vdd.n2444 vdd.n981 10.6151
R4395 vdd.n2445 vdd.n2444 10.6151
R4396 vdd.n2448 vdd.n2445 10.6151
R4397 vdd.n2448 vdd.n2447 10.6151
R4398 vdd.n2447 vdd.n2446 10.6151
R4399 vdd.n2446 vdd.n964 10.6151
R4400 vdd.n2530 vdd.n964 10.6151
R4401 vdd.n2529 vdd.n2528 10.6151
R4402 vdd.n2528 vdd.n2525 10.6151
R4403 vdd.n2525 vdd.n2524 10.6151
R4404 vdd.n2524 vdd.n2521 10.6151
R4405 vdd.n2521 vdd.n2520 10.6151
R4406 vdd.n2520 vdd.n2517 10.6151
R4407 vdd.n2517 vdd.n2516 10.6151
R4408 vdd.n2516 vdd.n2513 10.6151
R4409 vdd.n2513 vdd.n2512 10.6151
R4410 vdd.n2512 vdd.n2509 10.6151
R4411 vdd.n2509 vdd.n2508 10.6151
R4412 vdd.n2508 vdd.n2505 10.6151
R4413 vdd.n2505 vdd.n2504 10.6151
R4414 vdd.n2504 vdd.n2501 10.6151
R4415 vdd.n2501 vdd.n2500 10.6151
R4416 vdd.n2500 vdd.n2497 10.6151
R4417 vdd.n2497 vdd.n2496 10.6151
R4418 vdd.n2496 vdd.n2493 10.6151
R4419 vdd.n2493 vdd.n2492 10.6151
R4420 vdd.n2492 vdd.n2489 10.6151
R4421 vdd.n2489 vdd.n2488 10.6151
R4422 vdd.n2488 vdd.n2485 10.6151
R4423 vdd.n2485 vdd.n2484 10.6151
R4424 vdd.n2484 vdd.n2481 10.6151
R4425 vdd.n2481 vdd.n2480 10.6151
R4426 vdd.n2480 vdd.n2477 10.6151
R4427 vdd.n2477 vdd.n2476 10.6151
R4428 vdd.n2476 vdd.n2473 10.6151
R4429 vdd.n2473 vdd.n2472 10.6151
R4430 vdd.n2472 vdd.n2469 10.6151
R4431 vdd.n2469 vdd.n2468 10.6151
R4432 vdd.n2465 vdd.n2464 10.6151
R4433 vdd.n2464 vdd.n2462 10.6151
R4434 vdd.n2221 vdd.n2219 10.6151
R4435 vdd.n2222 vdd.n2221 10.6151
R4436 vdd.n2224 vdd.n2222 10.6151
R4437 vdd.n2225 vdd.n2224 10.6151
R4438 vdd.n2227 vdd.n2225 10.6151
R4439 vdd.n2228 vdd.n2227 10.6151
R4440 vdd.n2230 vdd.n2228 10.6151
R4441 vdd.n2231 vdd.n2230 10.6151
R4442 vdd.n2233 vdd.n2231 10.6151
R4443 vdd.n2234 vdd.n2233 10.6151
R4444 vdd.n2236 vdd.n2234 10.6151
R4445 vdd.n2237 vdd.n2236 10.6151
R4446 vdd.n2255 vdd.n2237 10.6151
R4447 vdd.n2255 vdd.n2254 10.6151
R4448 vdd.n2254 vdd.n2253 10.6151
R4449 vdd.n2253 vdd.n2251 10.6151
R4450 vdd.n2251 vdd.n2250 10.6151
R4451 vdd.n2250 vdd.n2248 10.6151
R4452 vdd.n2248 vdd.n2247 10.6151
R4453 vdd.n2247 vdd.n2245 10.6151
R4454 vdd.n2245 vdd.n2244 10.6151
R4455 vdd.n2244 vdd.n2242 10.6151
R4456 vdd.n2242 vdd.n2241 10.6151
R4457 vdd.n2241 vdd.n2239 10.6151
R4458 vdd.n2239 vdd.n2238 10.6151
R4459 vdd.n2238 vdd.n968 10.6151
R4460 vdd.n2460 vdd.n968 10.6151
R4461 vdd.n2461 vdd.n2460 10.6151
R4462 vdd.n2372 vdd.n2371 10.6151
R4463 vdd.n2371 vdd.n1053 10.6151
R4464 vdd.n2365 vdd.n1053 10.6151
R4465 vdd.n2365 vdd.n2364 10.6151
R4466 vdd.n2364 vdd.n2363 10.6151
R4467 vdd.n2363 vdd.n1055 10.6151
R4468 vdd.n2357 vdd.n1055 10.6151
R4469 vdd.n2357 vdd.n2356 10.6151
R4470 vdd.n2356 vdd.n2355 10.6151
R4471 vdd.n2355 vdd.n1057 10.6151
R4472 vdd.n2349 vdd.n1057 10.6151
R4473 vdd.n2349 vdd.n2348 10.6151
R4474 vdd.n2348 vdd.n2347 10.6151
R4475 vdd.n2347 vdd.n1059 10.6151
R4476 vdd.n2341 vdd.n1059 10.6151
R4477 vdd.n2341 vdd.n2340 10.6151
R4478 vdd.n2340 vdd.n2339 10.6151
R4479 vdd.n2339 vdd.n1063 10.6151
R4480 vdd.n2187 vdd.n1063 10.6151
R4481 vdd.n2188 vdd.n2187 10.6151
R4482 vdd.n2188 vdd.n2183 10.6151
R4483 vdd.n2194 vdd.n2183 10.6151
R4484 vdd.n2195 vdd.n2194 10.6151
R4485 vdd.n2196 vdd.n2195 10.6151
R4486 vdd.n2196 vdd.n2181 10.6151
R4487 vdd.n2202 vdd.n2181 10.6151
R4488 vdd.n2203 vdd.n2202 10.6151
R4489 vdd.n2204 vdd.n2203 10.6151
R4490 vdd.n2204 vdd.n2179 10.6151
R4491 vdd.n2210 vdd.n2179 10.6151
R4492 vdd.n2211 vdd.n2210 10.6151
R4493 vdd.n2213 vdd.n2175 10.6151
R4494 vdd.n2218 vdd.n2175 10.6151
R4495 vdd.n1851 vdd.t67 10.5435
R4496 vdd.n656 vdd.t99 10.5435
R4497 vdd.n316 vdd.n298 10.4732
R4498 vdd.n257 vdd.n239 10.4732
R4499 vdd.n214 vdd.n196 10.4732
R4500 vdd.n155 vdd.n137 10.4732
R4501 vdd.n113 vdd.n95 10.4732
R4502 vdd.n54 vdd.n36 10.4732
R4503 vdd.n1735 vdd.n1717 10.4732
R4504 vdd.n1794 vdd.n1776 10.4732
R4505 vdd.n1633 vdd.n1615 10.4732
R4506 vdd.n1692 vdd.n1674 10.4732
R4507 vdd.n1532 vdd.n1514 10.4732
R4508 vdd.n1591 vdd.n1573 10.4732
R4509 vdd.t76 vdd.n1825 10.3167
R4510 vdd.n3300 vdd.t16 10.3167
R4511 vdd.n1502 vdd.t115 10.09
R4512 vdd.n3394 vdd.t64 10.09
R4513 vdd.t26 vdd.n1155 9.86327
R4514 vdd.n3385 vdd.t37 9.86327
R4515 vdd.n315 vdd.n300 9.69747
R4516 vdd.n256 vdd.n241 9.69747
R4517 vdd.n213 vdd.n198 9.69747
R4518 vdd.n154 vdd.n139 9.69747
R4519 vdd.n112 vdd.n97 9.69747
R4520 vdd.n53 vdd.n38 9.69747
R4521 vdd.n1734 vdd.n1719 9.69747
R4522 vdd.n1793 vdd.n1778 9.69747
R4523 vdd.n1632 vdd.n1617 9.69747
R4524 vdd.n1691 vdd.n1676 9.69747
R4525 vdd.n1531 vdd.n1516 9.69747
R4526 vdd.n1590 vdd.n1575 9.69747
R4527 vdd.n2315 vdd.n2314 9.67831
R4528 vdd.n3216 vdd.n731 9.67831
R4529 vdd.n3093 vdd.n3092 9.67831
R4530 vdd.n2339 vdd.n2338 9.67831
R4531 vdd.n1461 vdd.t54 9.63654
R4532 vdd.n3331 vdd.t30 9.63654
R4533 vdd.n331 vdd.n330 9.45567
R4534 vdd.n272 vdd.n271 9.45567
R4535 vdd.n229 vdd.n228 9.45567
R4536 vdd.n170 vdd.n169 9.45567
R4537 vdd.n128 vdd.n127 9.45567
R4538 vdd.n69 vdd.n68 9.45567
R4539 vdd.n1750 vdd.n1749 9.45567
R4540 vdd.n1809 vdd.n1808 9.45567
R4541 vdd.n1648 vdd.n1647 9.45567
R4542 vdd.n1707 vdd.n1706 9.45567
R4543 vdd.n1547 vdd.n1546 9.45567
R4544 vdd.n1606 vdd.n1605 9.45567
R4545 vdd.n1435 vdd.t52 9.40981
R4546 vdd.n3363 vdd.t103 9.40981
R4547 vdd.n2075 vdd.n1929 9.3005
R4548 vdd.n2074 vdd.n2073 9.3005
R4549 vdd.n1935 vdd.n1934 9.3005
R4550 vdd.n2068 vdd.n1939 9.3005
R4551 vdd.n2067 vdd.n1940 9.3005
R4552 vdd.n2066 vdd.n1941 9.3005
R4553 vdd.n1945 vdd.n1942 9.3005
R4554 vdd.n2061 vdd.n1946 9.3005
R4555 vdd.n2060 vdd.n1947 9.3005
R4556 vdd.n2059 vdd.n1948 9.3005
R4557 vdd.n1952 vdd.n1949 9.3005
R4558 vdd.n2054 vdd.n1953 9.3005
R4559 vdd.n2053 vdd.n1954 9.3005
R4560 vdd.n2052 vdd.n1955 9.3005
R4561 vdd.n1959 vdd.n1956 9.3005
R4562 vdd.n2047 vdd.n1960 9.3005
R4563 vdd.n2046 vdd.n1961 9.3005
R4564 vdd.n2045 vdd.n1962 9.3005
R4565 vdd.n1966 vdd.n1963 9.3005
R4566 vdd.n2040 vdd.n1967 9.3005
R4567 vdd.n2039 vdd.n1968 9.3005
R4568 vdd.n2038 vdd.n2037 9.3005
R4569 vdd.n2036 vdd.n1969 9.3005
R4570 vdd.n2035 vdd.n2034 9.3005
R4571 vdd.n1975 vdd.n1974 9.3005
R4572 vdd.n2029 vdd.n1979 9.3005
R4573 vdd.n2028 vdd.n1980 9.3005
R4574 vdd.n2027 vdd.n1981 9.3005
R4575 vdd.n1985 vdd.n1982 9.3005
R4576 vdd.n2022 vdd.n1986 9.3005
R4577 vdd.n2021 vdd.n1987 9.3005
R4578 vdd.n2020 vdd.n1988 9.3005
R4579 vdd.n1992 vdd.n1989 9.3005
R4580 vdd.n2015 vdd.n1993 9.3005
R4581 vdd.n2014 vdd.n1994 9.3005
R4582 vdd.n2013 vdd.n1995 9.3005
R4583 vdd.n1997 vdd.n1996 9.3005
R4584 vdd.n2008 vdd.n1064 9.3005
R4585 vdd.n2077 vdd.n2076 9.3005
R4586 vdd.n2101 vdd.n2100 9.3005
R4587 vdd.n1907 vdd.n1906 9.3005
R4588 vdd.n1912 vdd.n1910 9.3005
R4589 vdd.n2093 vdd.n1913 9.3005
R4590 vdd.n2092 vdd.n1914 9.3005
R4591 vdd.n2091 vdd.n1915 9.3005
R4592 vdd.n1919 vdd.n1916 9.3005
R4593 vdd.n2086 vdd.n1920 9.3005
R4594 vdd.n2085 vdd.n1921 9.3005
R4595 vdd.n2084 vdd.n1922 9.3005
R4596 vdd.n1926 vdd.n1923 9.3005
R4597 vdd.n2079 vdd.n1927 9.3005
R4598 vdd.n2078 vdd.n1928 9.3005
R4599 vdd.n2323 vdd.n1900 9.3005
R4600 vdd.n2325 vdd.n2324 9.3005
R4601 vdd.n1815 vdd.n1814 9.3005
R4602 vdd.n1124 vdd.n1123 9.3005
R4603 vdd.n1829 vdd.n1828 9.3005
R4604 vdd.n1830 vdd.n1122 9.3005
R4605 vdd.n1832 vdd.n1831 9.3005
R4606 vdd.n1113 vdd.n1112 9.3005
R4607 vdd.n1846 vdd.n1845 9.3005
R4608 vdd.n1847 vdd.n1111 9.3005
R4609 vdd.n1849 vdd.n1848 9.3005
R4610 vdd.n1102 vdd.n1101 9.3005
R4611 vdd.n1862 vdd.n1861 9.3005
R4612 vdd.n1863 vdd.n1100 9.3005
R4613 vdd.n1865 vdd.n1864 9.3005
R4614 vdd.n1090 vdd.n1089 9.3005
R4615 vdd.n1879 vdd.n1878 9.3005
R4616 vdd.n1880 vdd.n1088 9.3005
R4617 vdd.n1882 vdd.n1881 9.3005
R4618 vdd.n1078 vdd.n1077 9.3005
R4619 vdd.n1898 vdd.n1897 9.3005
R4620 vdd.n1899 vdd.n1076 9.3005
R4621 vdd.n2327 vdd.n2326 9.3005
R4622 vdd.n307 vdd.n306 9.3005
R4623 vdd.n302 vdd.n301 9.3005
R4624 vdd.n313 vdd.n312 9.3005
R4625 vdd.n315 vdd.n314 9.3005
R4626 vdd.n298 vdd.n297 9.3005
R4627 vdd.n321 vdd.n320 9.3005
R4628 vdd.n323 vdd.n322 9.3005
R4629 vdd.n295 vdd.n292 9.3005
R4630 vdd.n330 vdd.n329 9.3005
R4631 vdd.n248 vdd.n247 9.3005
R4632 vdd.n243 vdd.n242 9.3005
R4633 vdd.n254 vdd.n253 9.3005
R4634 vdd.n256 vdd.n255 9.3005
R4635 vdd.n239 vdd.n238 9.3005
R4636 vdd.n262 vdd.n261 9.3005
R4637 vdd.n264 vdd.n263 9.3005
R4638 vdd.n236 vdd.n233 9.3005
R4639 vdd.n271 vdd.n270 9.3005
R4640 vdd.n205 vdd.n204 9.3005
R4641 vdd.n200 vdd.n199 9.3005
R4642 vdd.n211 vdd.n210 9.3005
R4643 vdd.n213 vdd.n212 9.3005
R4644 vdd.n196 vdd.n195 9.3005
R4645 vdd.n219 vdd.n218 9.3005
R4646 vdd.n221 vdd.n220 9.3005
R4647 vdd.n193 vdd.n190 9.3005
R4648 vdd.n228 vdd.n227 9.3005
R4649 vdd.n146 vdd.n145 9.3005
R4650 vdd.n141 vdd.n140 9.3005
R4651 vdd.n152 vdd.n151 9.3005
R4652 vdd.n154 vdd.n153 9.3005
R4653 vdd.n137 vdd.n136 9.3005
R4654 vdd.n160 vdd.n159 9.3005
R4655 vdd.n162 vdd.n161 9.3005
R4656 vdd.n134 vdd.n131 9.3005
R4657 vdd.n169 vdd.n168 9.3005
R4658 vdd.n104 vdd.n103 9.3005
R4659 vdd.n99 vdd.n98 9.3005
R4660 vdd.n110 vdd.n109 9.3005
R4661 vdd.n112 vdd.n111 9.3005
R4662 vdd.n95 vdd.n94 9.3005
R4663 vdd.n118 vdd.n117 9.3005
R4664 vdd.n120 vdd.n119 9.3005
R4665 vdd.n92 vdd.n89 9.3005
R4666 vdd.n127 vdd.n126 9.3005
R4667 vdd.n45 vdd.n44 9.3005
R4668 vdd.n40 vdd.n39 9.3005
R4669 vdd.n51 vdd.n50 9.3005
R4670 vdd.n53 vdd.n52 9.3005
R4671 vdd.n36 vdd.n35 9.3005
R4672 vdd.n59 vdd.n58 9.3005
R4673 vdd.n61 vdd.n60 9.3005
R4674 vdd.n33 vdd.n30 9.3005
R4675 vdd.n68 vdd.n67 9.3005
R4676 vdd.n3138 vdd.n3137 9.3005
R4677 vdd.n3141 vdd.n766 9.3005
R4678 vdd.n3142 vdd.n765 9.3005
R4679 vdd.n3145 vdd.n764 9.3005
R4680 vdd.n3146 vdd.n763 9.3005
R4681 vdd.n3149 vdd.n762 9.3005
R4682 vdd.n3150 vdd.n761 9.3005
R4683 vdd.n3153 vdd.n760 9.3005
R4684 vdd.n3154 vdd.n759 9.3005
R4685 vdd.n3157 vdd.n758 9.3005
R4686 vdd.n3158 vdd.n757 9.3005
R4687 vdd.n3161 vdd.n756 9.3005
R4688 vdd.n3162 vdd.n755 9.3005
R4689 vdd.n3165 vdd.n754 9.3005
R4690 vdd.n3166 vdd.n753 9.3005
R4691 vdd.n3169 vdd.n752 9.3005
R4692 vdd.n3170 vdd.n751 9.3005
R4693 vdd.n3173 vdd.n750 9.3005
R4694 vdd.n3174 vdd.n749 9.3005
R4695 vdd.n3177 vdd.n748 9.3005
R4696 vdd.n3181 vdd.n3180 9.3005
R4697 vdd.n3182 vdd.n747 9.3005
R4698 vdd.n3186 vdd.n3183 9.3005
R4699 vdd.n3189 vdd.n746 9.3005
R4700 vdd.n3190 vdd.n745 9.3005
R4701 vdd.n3193 vdd.n744 9.3005
R4702 vdd.n3194 vdd.n743 9.3005
R4703 vdd.n3197 vdd.n742 9.3005
R4704 vdd.n3198 vdd.n741 9.3005
R4705 vdd.n3201 vdd.n740 9.3005
R4706 vdd.n3202 vdd.n739 9.3005
R4707 vdd.n3205 vdd.n738 9.3005
R4708 vdd.n3206 vdd.n737 9.3005
R4709 vdd.n3209 vdd.n736 9.3005
R4710 vdd.n3210 vdd.n735 9.3005
R4711 vdd.n3213 vdd.n730 9.3005
R4712 vdd.n3219 vdd.n727 9.3005
R4713 vdd.n3220 vdd.n726 9.3005
R4714 vdd.n3234 vdd.n3233 9.3005
R4715 vdd.n3235 vdd.n681 9.3005
R4716 vdd.n3237 vdd.n3236 9.3005
R4717 vdd.n671 vdd.n670 9.3005
R4718 vdd.n3251 vdd.n3250 9.3005
R4719 vdd.n3252 vdd.n669 9.3005
R4720 vdd.n3254 vdd.n3253 9.3005
R4721 vdd.n660 vdd.n659 9.3005
R4722 vdd.n3267 vdd.n3266 9.3005
R4723 vdd.n3268 vdd.n658 9.3005
R4724 vdd.n3270 vdd.n3269 9.3005
R4725 vdd.n648 vdd.n647 9.3005
R4726 vdd.n3284 vdd.n3283 9.3005
R4727 vdd.n3285 vdd.n646 9.3005
R4728 vdd.n3287 vdd.n3286 9.3005
R4729 vdd.n637 vdd.n636 9.3005
R4730 vdd.n3303 vdd.n3302 9.3005
R4731 vdd.n3304 vdd.n635 9.3005
R4732 vdd.n3306 vdd.n3305 9.3005
R4733 vdd.n336 vdd.n334 9.3005
R4734 vdd.n683 vdd.n682 9.3005
R4735 vdd.n3398 vdd.n3397 9.3005
R4736 vdd.n337 vdd.n335 9.3005
R4737 vdd.n3391 vdd.n346 9.3005
R4738 vdd.n3390 vdd.n347 9.3005
R4739 vdd.n3389 vdd.n348 9.3005
R4740 vdd.n355 vdd.n349 9.3005
R4741 vdd.n3383 vdd.n356 9.3005
R4742 vdd.n3382 vdd.n357 9.3005
R4743 vdd.n3381 vdd.n358 9.3005
R4744 vdd.n366 vdd.n359 9.3005
R4745 vdd.n3375 vdd.n367 9.3005
R4746 vdd.n3374 vdd.n368 9.3005
R4747 vdd.n3373 vdd.n369 9.3005
R4748 vdd.n377 vdd.n370 9.3005
R4749 vdd.n3367 vdd.n378 9.3005
R4750 vdd.n3366 vdd.n379 9.3005
R4751 vdd.n3365 vdd.n380 9.3005
R4752 vdd.n388 vdd.n381 9.3005
R4753 vdd.n3359 vdd.n389 9.3005
R4754 vdd.n3358 vdd.n390 9.3005
R4755 vdd.n3357 vdd.n391 9.3005
R4756 vdd.n466 vdd.n463 9.3005
R4757 vdd.n470 vdd.n469 9.3005
R4758 vdd.n471 vdd.n462 9.3005
R4759 vdd.n475 vdd.n472 9.3005
R4760 vdd.n476 vdd.n461 9.3005
R4761 vdd.n480 vdd.n479 9.3005
R4762 vdd.n481 vdd.n460 9.3005
R4763 vdd.n485 vdd.n482 9.3005
R4764 vdd.n486 vdd.n459 9.3005
R4765 vdd.n490 vdd.n489 9.3005
R4766 vdd.n491 vdd.n458 9.3005
R4767 vdd.n495 vdd.n492 9.3005
R4768 vdd.n496 vdd.n457 9.3005
R4769 vdd.n500 vdd.n499 9.3005
R4770 vdd.n501 vdd.n456 9.3005
R4771 vdd.n505 vdd.n502 9.3005
R4772 vdd.n506 vdd.n455 9.3005
R4773 vdd.n510 vdd.n509 9.3005
R4774 vdd.n511 vdd.n454 9.3005
R4775 vdd.n515 vdd.n512 9.3005
R4776 vdd.n516 vdd.n451 9.3005
R4777 vdd.n520 vdd.n519 9.3005
R4778 vdd.n521 vdd.n450 9.3005
R4779 vdd.n525 vdd.n522 9.3005
R4780 vdd.n526 vdd.n449 9.3005
R4781 vdd.n530 vdd.n529 9.3005
R4782 vdd.n531 vdd.n448 9.3005
R4783 vdd.n535 vdd.n532 9.3005
R4784 vdd.n536 vdd.n447 9.3005
R4785 vdd.n540 vdd.n539 9.3005
R4786 vdd.n541 vdd.n446 9.3005
R4787 vdd.n545 vdd.n542 9.3005
R4788 vdd.n546 vdd.n445 9.3005
R4789 vdd.n550 vdd.n549 9.3005
R4790 vdd.n551 vdd.n444 9.3005
R4791 vdd.n555 vdd.n552 9.3005
R4792 vdd.n556 vdd.n443 9.3005
R4793 vdd.n560 vdd.n559 9.3005
R4794 vdd.n561 vdd.n442 9.3005
R4795 vdd.n565 vdd.n562 9.3005
R4796 vdd.n566 vdd.n439 9.3005
R4797 vdd.n570 vdd.n569 9.3005
R4798 vdd.n571 vdd.n438 9.3005
R4799 vdd.n575 vdd.n572 9.3005
R4800 vdd.n576 vdd.n437 9.3005
R4801 vdd.n580 vdd.n579 9.3005
R4802 vdd.n581 vdd.n436 9.3005
R4803 vdd.n585 vdd.n582 9.3005
R4804 vdd.n586 vdd.n435 9.3005
R4805 vdd.n590 vdd.n589 9.3005
R4806 vdd.n591 vdd.n434 9.3005
R4807 vdd.n595 vdd.n592 9.3005
R4808 vdd.n596 vdd.n433 9.3005
R4809 vdd.n600 vdd.n599 9.3005
R4810 vdd.n601 vdd.n432 9.3005
R4811 vdd.n605 vdd.n602 9.3005
R4812 vdd.n606 vdd.n431 9.3005
R4813 vdd.n610 vdd.n609 9.3005
R4814 vdd.n611 vdd.n430 9.3005
R4815 vdd.n615 vdd.n612 9.3005
R4816 vdd.n617 vdd.n429 9.3005
R4817 vdd.n619 vdd.n618 9.3005
R4818 vdd.n3351 vdd.n3350 9.3005
R4819 vdd.n465 vdd.n464 9.3005
R4820 vdd.n3229 vdd.n3228 9.3005
R4821 vdd.n676 vdd.n675 9.3005
R4822 vdd.n3242 vdd.n3241 9.3005
R4823 vdd.n3243 vdd.n674 9.3005
R4824 vdd.n3245 vdd.n3244 9.3005
R4825 vdd.n666 vdd.n665 9.3005
R4826 vdd.n3259 vdd.n3258 9.3005
R4827 vdd.n3260 vdd.n664 9.3005
R4828 vdd.n3262 vdd.n3261 9.3005
R4829 vdd.n653 vdd.n652 9.3005
R4830 vdd.n3275 vdd.n3274 9.3005
R4831 vdd.n3276 vdd.n651 9.3005
R4832 vdd.n3278 vdd.n3277 9.3005
R4833 vdd.n642 vdd.n641 9.3005
R4834 vdd.n3292 vdd.n3291 9.3005
R4835 vdd.n3293 vdd.n640 9.3005
R4836 vdd.n3298 vdd.n3294 9.3005
R4837 vdd.n3297 vdd.n3296 9.3005
R4838 vdd.n3295 vdd.n631 9.3005
R4839 vdd.n3311 vdd.n630 9.3005
R4840 vdd.n3313 vdd.n3312 9.3005
R4841 vdd.n3314 vdd.n629 9.3005
R4842 vdd.n3316 vdd.n3315 9.3005
R4843 vdd.n3318 vdd.n628 9.3005
R4844 vdd.n3320 vdd.n3319 9.3005
R4845 vdd.n3321 vdd.n627 9.3005
R4846 vdd.n3323 vdd.n3322 9.3005
R4847 vdd.n3325 vdd.n626 9.3005
R4848 vdd.n3327 vdd.n3326 9.3005
R4849 vdd.n3328 vdd.n625 9.3005
R4850 vdd.n3330 vdd.n3329 9.3005
R4851 vdd.n3333 vdd.n624 9.3005
R4852 vdd.n3335 vdd.n3334 9.3005
R4853 vdd.n3336 vdd.n623 9.3005
R4854 vdd.n3338 vdd.n3337 9.3005
R4855 vdd.n3340 vdd.n622 9.3005
R4856 vdd.n3342 vdd.n3341 9.3005
R4857 vdd.n3343 vdd.n621 9.3005
R4858 vdd.n3345 vdd.n3344 9.3005
R4859 vdd.n3347 vdd.n620 9.3005
R4860 vdd.n3349 vdd.n3348 9.3005
R4861 vdd.n3227 vdd.n686 9.3005
R4862 vdd.n3226 vdd.n3225 9.3005
R4863 vdd.n3095 vdd.n687 9.3005
R4864 vdd.n3104 vdd.n783 9.3005
R4865 vdd.n3107 vdd.n782 9.3005
R4866 vdd.n3108 vdd.n781 9.3005
R4867 vdd.n3111 vdd.n780 9.3005
R4868 vdd.n3112 vdd.n779 9.3005
R4869 vdd.n3115 vdd.n778 9.3005
R4870 vdd.n3116 vdd.n777 9.3005
R4871 vdd.n3119 vdd.n776 9.3005
R4872 vdd.n3120 vdd.n775 9.3005
R4873 vdd.n3123 vdd.n774 9.3005
R4874 vdd.n3124 vdd.n773 9.3005
R4875 vdd.n3127 vdd.n772 9.3005
R4876 vdd.n3128 vdd.n771 9.3005
R4877 vdd.n3131 vdd.n770 9.3005
R4878 vdd.n3135 vdd.n3134 9.3005
R4879 vdd.n3136 vdd.n767 9.3005
R4880 vdd.n2337 vdd.n2336 9.3005
R4881 vdd.n2332 vdd.n1067 9.3005
R4882 vdd.n1430 vdd.n1429 9.3005
R4883 vdd.n1431 vdd.n1185 9.3005
R4884 vdd.n1433 vdd.n1432 9.3005
R4885 vdd.n1175 vdd.n1174 9.3005
R4886 vdd.n1447 vdd.n1446 9.3005
R4887 vdd.n1448 vdd.n1173 9.3005
R4888 vdd.n1450 vdd.n1449 9.3005
R4889 vdd.n1165 vdd.n1164 9.3005
R4890 vdd.n1464 vdd.n1463 9.3005
R4891 vdd.n1465 vdd.n1163 9.3005
R4892 vdd.n1467 vdd.n1466 9.3005
R4893 vdd.n1152 vdd.n1151 9.3005
R4894 vdd.n1480 vdd.n1479 9.3005
R4895 vdd.n1481 vdd.n1150 9.3005
R4896 vdd.n1483 vdd.n1482 9.3005
R4897 vdd.n1141 vdd.n1140 9.3005
R4898 vdd.n1497 vdd.n1496 9.3005
R4899 vdd.n1498 vdd.n1139 9.3005
R4900 vdd.n1500 vdd.n1499 9.3005
R4901 vdd.n1130 vdd.n1129 9.3005
R4902 vdd.n1820 vdd.n1819 9.3005
R4903 vdd.n1821 vdd.n1128 9.3005
R4904 vdd.n1823 vdd.n1822 9.3005
R4905 vdd.n1118 vdd.n1117 9.3005
R4906 vdd.n1837 vdd.n1836 9.3005
R4907 vdd.n1838 vdd.n1116 9.3005
R4908 vdd.n1840 vdd.n1839 9.3005
R4909 vdd.n1108 vdd.n1107 9.3005
R4910 vdd.n1854 vdd.n1853 9.3005
R4911 vdd.n1855 vdd.n1106 9.3005
R4912 vdd.n1857 vdd.n1856 9.3005
R4913 vdd.n1095 vdd.n1094 9.3005
R4914 vdd.n1870 vdd.n1869 9.3005
R4915 vdd.n1871 vdd.n1093 9.3005
R4916 vdd.n1873 vdd.n1872 9.3005
R4917 vdd.n1085 vdd.n1084 9.3005
R4918 vdd.n1887 vdd.n1886 9.3005
R4919 vdd.n1888 vdd.n1082 9.3005
R4920 vdd.n1892 vdd.n1891 9.3005
R4921 vdd.n1890 vdd.n1083 9.3005
R4922 vdd.n1889 vdd.n1072 9.3005
R4923 vdd.n1187 vdd.n1186 9.3005
R4924 vdd.n1323 vdd.n1322 9.3005
R4925 vdd.n1324 vdd.n1313 9.3005
R4926 vdd.n1326 vdd.n1325 9.3005
R4927 vdd.n1327 vdd.n1312 9.3005
R4928 vdd.n1329 vdd.n1328 9.3005
R4929 vdd.n1330 vdd.n1307 9.3005
R4930 vdd.n1332 vdd.n1331 9.3005
R4931 vdd.n1333 vdd.n1306 9.3005
R4932 vdd.n1335 vdd.n1334 9.3005
R4933 vdd.n1336 vdd.n1301 9.3005
R4934 vdd.n1338 vdd.n1337 9.3005
R4935 vdd.n1339 vdd.n1300 9.3005
R4936 vdd.n1341 vdd.n1340 9.3005
R4937 vdd.n1342 vdd.n1295 9.3005
R4938 vdd.n1344 vdd.n1343 9.3005
R4939 vdd.n1345 vdd.n1294 9.3005
R4940 vdd.n1347 vdd.n1346 9.3005
R4941 vdd.n1348 vdd.n1289 9.3005
R4942 vdd.n1350 vdd.n1349 9.3005
R4943 vdd.n1351 vdd.n1288 9.3005
R4944 vdd.n1353 vdd.n1352 9.3005
R4945 vdd.n1357 vdd.n1284 9.3005
R4946 vdd.n1359 vdd.n1358 9.3005
R4947 vdd.n1360 vdd.n1283 9.3005
R4948 vdd.n1362 vdd.n1361 9.3005
R4949 vdd.n1363 vdd.n1278 9.3005
R4950 vdd.n1365 vdd.n1364 9.3005
R4951 vdd.n1366 vdd.n1277 9.3005
R4952 vdd.n1368 vdd.n1367 9.3005
R4953 vdd.n1369 vdd.n1272 9.3005
R4954 vdd.n1371 vdd.n1370 9.3005
R4955 vdd.n1372 vdd.n1271 9.3005
R4956 vdd.n1374 vdd.n1373 9.3005
R4957 vdd.n1375 vdd.n1266 9.3005
R4958 vdd.n1377 vdd.n1376 9.3005
R4959 vdd.n1378 vdd.n1265 9.3005
R4960 vdd.n1380 vdd.n1379 9.3005
R4961 vdd.n1381 vdd.n1260 9.3005
R4962 vdd.n1383 vdd.n1382 9.3005
R4963 vdd.n1384 vdd.n1259 9.3005
R4964 vdd.n1386 vdd.n1385 9.3005
R4965 vdd.n1387 vdd.n1254 9.3005
R4966 vdd.n1389 vdd.n1388 9.3005
R4967 vdd.n1390 vdd.n1253 9.3005
R4968 vdd.n1392 vdd.n1391 9.3005
R4969 vdd.n1393 vdd.n1246 9.3005
R4970 vdd.n1395 vdd.n1394 9.3005
R4971 vdd.n1396 vdd.n1245 9.3005
R4972 vdd.n1398 vdd.n1397 9.3005
R4973 vdd.n1399 vdd.n1240 9.3005
R4974 vdd.n1401 vdd.n1400 9.3005
R4975 vdd.n1402 vdd.n1239 9.3005
R4976 vdd.n1404 vdd.n1403 9.3005
R4977 vdd.n1405 vdd.n1234 9.3005
R4978 vdd.n1407 vdd.n1406 9.3005
R4979 vdd.n1408 vdd.n1233 9.3005
R4980 vdd.n1410 vdd.n1409 9.3005
R4981 vdd.n1411 vdd.n1228 9.3005
R4982 vdd.n1413 vdd.n1412 9.3005
R4983 vdd.n1414 vdd.n1227 9.3005
R4984 vdd.n1416 vdd.n1415 9.3005
R4985 vdd.n1192 vdd.n1191 9.3005
R4986 vdd.n1422 vdd.n1421 9.3005
R4987 vdd.n1321 vdd.n1320 9.3005
R4988 vdd.n1425 vdd.n1424 9.3005
R4989 vdd.n1181 vdd.n1180 9.3005
R4990 vdd.n1439 vdd.n1438 9.3005
R4991 vdd.n1440 vdd.n1179 9.3005
R4992 vdd.n1442 vdd.n1441 9.3005
R4993 vdd.n1170 vdd.n1169 9.3005
R4994 vdd.n1456 vdd.n1455 9.3005
R4995 vdd.n1457 vdd.n1168 9.3005
R4996 vdd.n1459 vdd.n1458 9.3005
R4997 vdd.n1159 vdd.n1158 9.3005
R4998 vdd.n1472 vdd.n1471 9.3005
R4999 vdd.n1473 vdd.n1157 9.3005
R5000 vdd.n1475 vdd.n1474 9.3005
R5001 vdd.n1147 vdd.n1146 9.3005
R5002 vdd.n1489 vdd.n1488 9.3005
R5003 vdd.n1490 vdd.n1145 9.3005
R5004 vdd.n1492 vdd.n1491 9.3005
R5005 vdd.n1136 vdd.n1135 9.3005
R5006 vdd.n1505 vdd.n1504 9.3005
R5007 vdd.n1506 vdd.n1134 9.3005
R5008 vdd.n1423 vdd.n1190 9.3005
R5009 vdd.n1726 vdd.n1725 9.3005
R5010 vdd.n1721 vdd.n1720 9.3005
R5011 vdd.n1732 vdd.n1731 9.3005
R5012 vdd.n1734 vdd.n1733 9.3005
R5013 vdd.n1717 vdd.n1716 9.3005
R5014 vdd.n1740 vdd.n1739 9.3005
R5015 vdd.n1742 vdd.n1741 9.3005
R5016 vdd.n1714 vdd.n1711 9.3005
R5017 vdd.n1749 vdd.n1748 9.3005
R5018 vdd.n1785 vdd.n1784 9.3005
R5019 vdd.n1780 vdd.n1779 9.3005
R5020 vdd.n1791 vdd.n1790 9.3005
R5021 vdd.n1793 vdd.n1792 9.3005
R5022 vdd.n1776 vdd.n1775 9.3005
R5023 vdd.n1799 vdd.n1798 9.3005
R5024 vdd.n1801 vdd.n1800 9.3005
R5025 vdd.n1773 vdd.n1770 9.3005
R5026 vdd.n1808 vdd.n1807 9.3005
R5027 vdd.n1624 vdd.n1623 9.3005
R5028 vdd.n1619 vdd.n1618 9.3005
R5029 vdd.n1630 vdd.n1629 9.3005
R5030 vdd.n1632 vdd.n1631 9.3005
R5031 vdd.n1615 vdd.n1614 9.3005
R5032 vdd.n1638 vdd.n1637 9.3005
R5033 vdd.n1640 vdd.n1639 9.3005
R5034 vdd.n1612 vdd.n1609 9.3005
R5035 vdd.n1647 vdd.n1646 9.3005
R5036 vdd.n1683 vdd.n1682 9.3005
R5037 vdd.n1678 vdd.n1677 9.3005
R5038 vdd.n1689 vdd.n1688 9.3005
R5039 vdd.n1691 vdd.n1690 9.3005
R5040 vdd.n1674 vdd.n1673 9.3005
R5041 vdd.n1697 vdd.n1696 9.3005
R5042 vdd.n1699 vdd.n1698 9.3005
R5043 vdd.n1671 vdd.n1668 9.3005
R5044 vdd.n1706 vdd.n1705 9.3005
R5045 vdd.n1523 vdd.n1522 9.3005
R5046 vdd.n1518 vdd.n1517 9.3005
R5047 vdd.n1529 vdd.n1528 9.3005
R5048 vdd.n1531 vdd.n1530 9.3005
R5049 vdd.n1514 vdd.n1513 9.3005
R5050 vdd.n1537 vdd.n1536 9.3005
R5051 vdd.n1539 vdd.n1538 9.3005
R5052 vdd.n1511 vdd.n1508 9.3005
R5053 vdd.n1546 vdd.n1545 9.3005
R5054 vdd.n1582 vdd.n1581 9.3005
R5055 vdd.n1577 vdd.n1576 9.3005
R5056 vdd.n1588 vdd.n1587 9.3005
R5057 vdd.n1590 vdd.n1589 9.3005
R5058 vdd.n1573 vdd.n1572 9.3005
R5059 vdd.n1596 vdd.n1595 9.3005
R5060 vdd.n1598 vdd.n1597 9.3005
R5061 vdd.n1570 vdd.n1567 9.3005
R5062 vdd.n1605 vdd.n1604 9.3005
R5063 vdd.n1461 vdd.t41 9.18308
R5064 vdd.n3331 vdd.t125 9.18308
R5065 vdd.n1155 vdd.t28 8.95635
R5066 vdd.n2329 vdd.t152 8.95635
R5067 vdd.n723 vdd.t145 8.95635
R5068 vdd.t24 vdd.n3385 8.95635
R5069 vdd.n312 vdd.n311 8.92171
R5070 vdd.n253 vdd.n252 8.92171
R5071 vdd.n210 vdd.n209 8.92171
R5072 vdd.n151 vdd.n150 8.92171
R5073 vdd.n109 vdd.n108 8.92171
R5074 vdd.n50 vdd.n49 8.92171
R5075 vdd.n1731 vdd.n1730 8.92171
R5076 vdd.n1790 vdd.n1789 8.92171
R5077 vdd.n1629 vdd.n1628 8.92171
R5078 vdd.n1688 vdd.n1687 8.92171
R5079 vdd.n1528 vdd.n1527 8.92171
R5080 vdd.n1587 vdd.n1586 8.92171
R5081 vdd.n231 vdd.n129 8.81535
R5082 vdd.n1709 vdd.n1607 8.81535
R5083 vdd.n1502 vdd.t43 8.72962
R5084 vdd.t7 vdd.n3394 8.72962
R5085 vdd.n1825 vdd.t59 8.50289
R5086 vdd.n3300 vdd.t3 8.50289
R5087 vdd.n28 vdd.n14 8.42249
R5088 vdd.n1851 vdd.t50 8.27616
R5089 vdd.t18 vdd.n656 8.27616
R5090 vdd.n3400 vdd.n3399 8.16225
R5091 vdd.n1813 vdd.n1812 8.16225
R5092 vdd.n308 vdd.n302 8.14595
R5093 vdd.n249 vdd.n243 8.14595
R5094 vdd.n206 vdd.n200 8.14595
R5095 vdd.n147 vdd.n141 8.14595
R5096 vdd.n105 vdd.n99 8.14595
R5097 vdd.n46 vdd.n40 8.14595
R5098 vdd.n1727 vdd.n1721 8.14595
R5099 vdd.n1786 vdd.n1780 8.14595
R5100 vdd.n1625 vdd.n1619 8.14595
R5101 vdd.n1684 vdd.n1678 8.14595
R5102 vdd.n1524 vdd.n1518 8.14595
R5103 vdd.n1583 vdd.n1577 8.14595
R5104 vdd.n2923 vdd.n849 8.11757
R5105 vdd.n2397 vdd.n2396 8.11757
R5106 vdd.n1098 vdd.t227 8.04943
R5107 vdd.n3256 vdd.t20 8.04943
R5108 vdd.n2375 vdd.n1043 7.70933
R5109 vdd.n2381 vdd.n1043 7.70933
R5110 vdd.n2387 vdd.n1037 7.70933
R5111 vdd.n2387 vdd.n1030 7.70933
R5112 vdd.n2393 vdd.n1030 7.70933
R5113 vdd.n2393 vdd.n1033 7.70933
R5114 vdd.n2400 vdd.n1018 7.70933
R5115 vdd.n2406 vdd.n1018 7.70933
R5116 vdd.n2412 vdd.n1012 7.70933
R5117 vdd.n2418 vdd.n1008 7.70933
R5118 vdd.n2424 vdd.n1002 7.70933
R5119 vdd.n2436 vdd.n989 7.70933
R5120 vdd.n2442 vdd.n983 7.70933
R5121 vdd.n2442 vdd.n976 7.70933
R5122 vdd.n2450 vdd.n976 7.70933
R5123 vdd.n2457 vdd.t268 7.70933
R5124 vdd.n2532 vdd.t268 7.70933
R5125 vdd.n2864 vdd.t235 7.70933
R5126 vdd.n2870 vdd.t235 7.70933
R5127 vdd.n2876 vdd.n897 7.70933
R5128 vdd.n2882 vdd.n897 7.70933
R5129 vdd.n2882 vdd.n900 7.70933
R5130 vdd.n2888 vdd.n893 7.70933
R5131 vdd.n2900 vdd.n880 7.70933
R5132 vdd.n2906 vdd.n874 7.70933
R5133 vdd.n2912 vdd.n870 7.70933
R5134 vdd.n2918 vdd.n857 7.70933
R5135 vdd.n2926 vdd.n857 7.70933
R5136 vdd.n2932 vdd.n851 7.70933
R5137 vdd.n2932 vdd.n843 7.70933
R5138 vdd.n2983 vdd.n843 7.70933
R5139 vdd.n2983 vdd.n846 7.70933
R5140 vdd.n2989 vdd.n805 7.70933
R5141 vdd.n3059 vdd.n805 7.70933
R5142 vdd.n307 vdd.n304 7.3702
R5143 vdd.n248 vdd.n245 7.3702
R5144 vdd.n205 vdd.n202 7.3702
R5145 vdd.n146 vdd.n143 7.3702
R5146 vdd.n104 vdd.n101 7.3702
R5147 vdd.n45 vdd.n42 7.3702
R5148 vdd.n1726 vdd.n1723 7.3702
R5149 vdd.n1785 vdd.n1782 7.3702
R5150 vdd.n1624 vdd.n1621 7.3702
R5151 vdd.n1683 vdd.n1680 7.3702
R5152 vdd.n1523 vdd.n1520 7.3702
R5153 vdd.n1582 vdd.n1579 7.3702
R5154 vdd.n1884 vdd.t61 7.1425
R5155 vdd.n679 vdd.t22 7.1425
R5156 vdd.n1358 vdd.n1357 6.98232
R5157 vdd.n2039 vdd.n2038 6.98232
R5158 vdd.n566 vdd.n565 6.98232
R5159 vdd.n3141 vdd.n3138 6.98232
R5160 vdd.t57 vdd.n1097 6.91577
R5161 vdd.n3264 vdd.t80 6.91577
R5162 vdd.n1843 vdd.t70 6.68904
R5163 vdd.n3280 vdd.t82 6.68904
R5164 vdd.t85 vdd.n1126 6.46231
R5165 vdd.n3308 vdd.t14 6.46231
R5166 vdd.n3400 vdd.n333 6.38151
R5167 vdd.n1812 vdd.n1811 6.38151
R5168 vdd.n1494 vdd.t32 6.23558
R5169 vdd.t224 vdd.n344 6.23558
R5170 vdd.t87 vdd.n1154 6.00885
R5171 vdd.n2412 vdd.t270 6.00885
R5172 vdd.n2912 vdd.t260 6.00885
R5173 vdd.n3379 vdd.t95 6.00885
R5174 vdd.n1033 vdd.t199 5.89549
R5175 vdd.t156 vdd.n851 5.89549
R5176 vdd.n308 vdd.n307 5.81868
R5177 vdd.n249 vdd.n248 5.81868
R5178 vdd.n206 vdd.n205 5.81868
R5179 vdd.n147 vdd.n146 5.81868
R5180 vdd.n105 vdd.n104 5.81868
R5181 vdd.n46 vdd.n45 5.81868
R5182 vdd.n1727 vdd.n1726 5.81868
R5183 vdd.n1786 vdd.n1785 5.81868
R5184 vdd.n1625 vdd.n1624 5.81868
R5185 vdd.n1684 vdd.n1683 5.81868
R5186 vdd.n1524 vdd.n1523 5.81868
R5187 vdd.n1583 vdd.n1582 5.81868
R5188 vdd.n1453 vdd.t39 5.78212
R5189 vdd.t195 vdd.n1037 5.78212
R5190 vdd.n2156 vdd.t180 5.78212
R5191 vdd.n2781 vdd.t188 5.78212
R5192 vdd.n846 vdd.t184 5.78212
R5193 vdd.n3370 vdd.t74 5.78212
R5194 vdd.n2540 vdd.n2539 5.77611
R5195 vdd.n2283 vdd.n2153 5.77611
R5196 vdd.n2794 vdd.n2793 5.77611
R5197 vdd.n3000 vdd.n2999 5.77611
R5198 vdd.n3064 vdd.n801 5.77611
R5199 vdd.n2704 vdd.n2644 5.77611
R5200 vdd.n2465 vdd.n967 5.77611
R5201 vdd.n2213 vdd.n2212 5.77611
R5202 vdd.n1320 vdd.n1319 5.62474
R5203 vdd.n2335 vdd.n2332 5.62474
R5204 vdd.n3351 vdd.n428 5.62474
R5205 vdd.n3225 vdd.n690 5.62474
R5206 vdd.n1177 vdd.t39 5.55539
R5207 vdd.t74 vdd.n3369 5.55539
R5208 vdd.t274 vdd.n989 5.44203
R5209 vdd.n893 vdd.t264 5.44203
R5210 vdd.n1469 vdd.t87 5.32866
R5211 vdd.t95 vdd.n3378 5.32866
R5212 vdd.n1485 vdd.t32 5.10193
R5213 vdd.t242 vdd.n1012 5.10193
R5214 vdd.n1002 vdd.t250 5.10193
R5215 vdd.t261 vdd.n880 5.10193
R5216 vdd.n870 vdd.t247 5.10193
R5217 vdd.n3387 vdd.t224 5.10193
R5218 vdd.n311 vdd.n302 5.04292
R5219 vdd.n252 vdd.n243 5.04292
R5220 vdd.n209 vdd.n200 5.04292
R5221 vdd.n150 vdd.n141 5.04292
R5222 vdd.n108 vdd.n99 5.04292
R5223 vdd.n49 vdd.n40 5.04292
R5224 vdd.n1730 vdd.n1721 5.04292
R5225 vdd.n1789 vdd.n1780 5.04292
R5226 vdd.n1628 vdd.n1619 5.04292
R5227 vdd.n1687 vdd.n1678 5.04292
R5228 vdd.n1527 vdd.n1518 5.04292
R5229 vdd.n1586 vdd.n1577 5.04292
R5230 vdd.n1817 vdd.t85 4.8752
R5231 vdd.t239 vdd.t248 4.8752
R5232 vdd.t271 vdd.t258 4.8752
R5233 vdd.t251 vdd.t232 4.8752
R5234 vdd.t272 vdd.t255 4.8752
R5235 vdd.t14 vdd.n340 4.8752
R5236 vdd.n2541 vdd.n2540 4.83952
R5237 vdd.n2153 vdd.n2149 4.83952
R5238 vdd.n2795 vdd.n2794 4.83952
R5239 vdd.n3001 vdd.n3000 4.83952
R5240 vdd.n801 vdd.n796 4.83952
R5241 vdd.n2701 vdd.n2644 4.83952
R5242 vdd.n2468 vdd.n967 4.83952
R5243 vdd.n2212 vdd.n2211 4.83952
R5244 vdd.n2007 vdd.n1065 4.74817
R5245 vdd.n2002 vdd.n1066 4.74817
R5246 vdd.n1904 vdd.n1901 4.74817
R5247 vdd.n2316 vdd.n1905 4.74817
R5248 vdd.n2318 vdd.n1904 4.74817
R5249 vdd.n2317 vdd.n2316 4.74817
R5250 vdd.n3218 vdd.n3217 4.74817
R5251 vdd.n3215 vdd.n3214 4.74817
R5252 vdd.n3215 vdd.n732 4.74817
R5253 vdd.n3217 vdd.n729 4.74817
R5254 vdd.n3100 vdd.n784 4.74817
R5255 vdd.n3096 vdd.n3094 4.74817
R5256 vdd.n3099 vdd.n3094 4.74817
R5257 vdd.n3103 vdd.n784 4.74817
R5258 vdd.n2003 vdd.n1065 4.74817
R5259 vdd.n1068 vdd.n1066 4.74817
R5260 vdd.n333 vdd.n332 4.7074
R5261 vdd.n231 vdd.n230 4.7074
R5262 vdd.n1811 vdd.n1810 4.7074
R5263 vdd.n1709 vdd.n1708 4.7074
R5264 vdd.n1120 vdd.t70 4.64847
R5265 vdd.n3289 vdd.t82 4.64847
R5266 vdd.n2418 vdd.t262 4.53511
R5267 vdd.n2906 vdd.t243 4.53511
R5268 vdd.n1859 vdd.t57 4.42174
R5269 vdd.t80 vdd.n655 4.42174
R5270 vdd.n2450 vdd.t245 4.30838
R5271 vdd.n2876 vdd.t233 4.30838
R5272 vdd.n312 vdd.n300 4.26717
R5273 vdd.n253 vdd.n241 4.26717
R5274 vdd.n210 vdd.n198 4.26717
R5275 vdd.n151 vdd.n139 4.26717
R5276 vdd.n109 vdd.n97 4.26717
R5277 vdd.n50 vdd.n38 4.26717
R5278 vdd.n1731 vdd.n1719 4.26717
R5279 vdd.n1790 vdd.n1778 4.26717
R5280 vdd.n1629 vdd.n1617 4.26717
R5281 vdd.n1688 vdd.n1676 4.26717
R5282 vdd.n1528 vdd.n1516 4.26717
R5283 vdd.n1587 vdd.n1575 4.26717
R5284 vdd.n1875 vdd.t61 4.19501
R5285 vdd.n3248 vdd.t22 4.19501
R5286 vdd.n333 vdd.n231 4.10845
R5287 vdd.n1811 vdd.n1709 4.10845
R5288 vdd.n289 vdd.t129 4.06363
R5289 vdd.n289 vdd.t131 4.06363
R5290 vdd.n287 vdd.t283 4.06363
R5291 vdd.n287 vdd.t292 4.06363
R5292 vdd.n285 vdd.t90 4.06363
R5293 vdd.n285 vdd.t140 4.06363
R5294 vdd.n283 vdd.t278 4.06363
R5295 vdd.n283 vdd.t294 4.06363
R5296 vdd.n281 vdd.t89 4.06363
R5297 vdd.n281 vdd.t13 4.06363
R5298 vdd.n279 vdd.t135 4.06363
R5299 vdd.n279 vdd.t91 4.06363
R5300 vdd.n277 vdd.t100 4.06363
R5301 vdd.n277 vdd.t117 4.06363
R5302 vdd.n275 vdd.t108 4.06363
R5303 vdd.n275 vdd.t122 4.06363
R5304 vdd.n273 vdd.t21 4.06363
R5305 vdd.n273 vdd.t229 4.06363
R5306 vdd.n187 vdd.t36 4.06363
R5307 vdd.n187 vdd.t75 4.06363
R5308 vdd.n185 vdd.t96 4.06363
R5309 vdd.n185 vdd.t287 4.06363
R5310 vdd.n183 vdd.t285 4.06363
R5311 vdd.n183 vdd.t38 4.06363
R5312 vdd.n181 vdd.t277 4.06363
R5313 vdd.n181 vdd.t225 4.06363
R5314 vdd.n179 vdd.t230 4.06363
R5315 vdd.n179 vdd.t8 4.06363
R5316 vdd.n177 vdd.t4 4.06363
R5317 vdd.n177 vdd.t17 4.06363
R5318 vdd.n175 vdd.t106 4.06363
R5319 vdd.n175 vdd.t83 4.06363
R5320 vdd.n173 vdd.t134 4.06363
R5321 vdd.n173 vdd.t34 4.06363
R5322 vdd.n171 vdd.t45 4.06363
R5323 vdd.n171 vdd.t94 4.06363
R5324 vdd.n86 vdd.t31 4.06363
R5325 vdd.n86 vdd.t97 4.06363
R5326 vdd.n84 vdd.t105 4.06363
R5327 vdd.n84 vdd.t126 4.06363
R5328 vdd.n82 vdd.t25 4.06363
R5329 vdd.n82 vdd.t286 4.06363
R5330 vdd.n80 vdd.t65 4.06363
R5331 vdd.n80 vdd.t280 4.06363
R5332 vdd.n78 vdd.t15 4.06363
R5333 vdd.n78 vdd.t12 4.06363
R5334 vdd.n76 vdd.t293 4.06363
R5335 vdd.n76 vdd.t98 4.06363
R5336 vdd.n74 vdd.t223 4.06363
R5337 vdd.n74 vdd.t119 4.06363
R5338 vdd.n72 vdd.t81 4.06363
R5339 vdd.n72 vdd.t19 4.06363
R5340 vdd.n70 vdd.t284 4.06363
R5341 vdd.n70 vdd.t73 4.06363
R5342 vdd.n1751 vdd.t276 4.06363
R5343 vdd.n1751 vdd.t290 4.06363
R5344 vdd.n1753 vdd.t289 4.06363
R5345 vdd.n1753 vdd.t101 4.06363
R5346 vdd.n1755 vdd.t78 4.06363
R5347 vdd.n1755 vdd.t68 4.06363
R5348 vdd.n1757 vdd.t84 4.06363
R5349 vdd.n1757 vdd.t220 4.06363
R5350 vdd.n1759 vdd.t128 4.06363
R5351 vdd.n1759 vdd.t110 4.06363
R5352 vdd.n1761 vdd.t69 4.06363
R5353 vdd.n1761 vdd.t127 4.06363
R5354 vdd.n1763 vdd.t27 4.06363
R5355 vdd.n1763 vdd.t29 4.06363
R5356 vdd.n1765 vdd.t42 4.06363
R5357 vdd.n1765 vdd.t279 4.06363
R5358 vdd.n1767 vdd.t40 4.06363
R5359 vdd.n1767 vdd.t130 4.06363
R5360 vdd.n1649 vdd.t6 4.06363
R5361 vdd.n1649 vdd.t228 4.06363
R5362 vdd.n1651 vdd.t102 4.06363
R5363 vdd.n1651 vdd.t58 4.06363
R5364 vdd.n1653 vdd.t92 4.06363
R5365 vdd.n1653 vdd.t114 4.06363
R5366 vdd.n1655 vdd.t288 4.06363
R5367 vdd.n1655 vdd.t60 4.06363
R5368 vdd.n1657 vdd.t133 4.06363
R5369 vdd.n1657 vdd.t109 4.06363
R5370 vdd.n1659 vdd.t33 4.06363
R5371 vdd.n1659 vdd.t132 4.06363
R5372 vdd.n1661 vdd.t120 4.06363
R5373 vdd.n1661 vdd.t121 4.06363
R5374 vdd.n1663 vdd.t111 4.06363
R5375 vdd.n1663 vdd.t88 4.06363
R5376 vdd.n1665 vdd.t113 4.06363
R5377 vdd.n1665 vdd.t55 4.06363
R5378 vdd.n1548 vdd.t281 4.06363
R5379 vdd.n1548 vdd.t231 4.06363
R5380 vdd.n1550 vdd.t51 4.06363
R5381 vdd.n1550 vdd.t221 4.06363
R5382 vdd.n1552 vdd.t71 4.06363
R5383 vdd.n1552 vdd.t222 4.06363
R5384 vdd.n1554 vdd.t77 4.06363
R5385 vdd.n1554 vdd.t295 4.06363
R5386 vdd.n1556 vdd.t44 4.06363
R5387 vdd.n1556 vdd.t86 4.06363
R5388 vdd.n1558 vdd.t56 4.06363
R5389 vdd.n1558 vdd.t116 4.06363
R5390 vdd.n1560 vdd.t226 4.06363
R5391 vdd.n1560 vdd.t79 4.06363
R5392 vdd.n1562 vdd.t124 4.06363
R5393 vdd.n1562 vdd.t93 4.06363
R5394 vdd.n1564 vdd.t123 4.06363
R5395 vdd.n1564 vdd.t112 4.06363
R5396 vdd.n26 vdd.t141 3.9605
R5397 vdd.n26 vdd.t48 3.9605
R5398 vdd.n23 vdd.t9 3.9605
R5399 vdd.n23 vdd.t10 3.9605
R5400 vdd.n21 vdd.t47 3.9605
R5401 vdd.n21 vdd.t0 3.9605
R5402 vdd.n20 vdd.t11 3.9605
R5403 vdd.n20 vdd.t138 3.9605
R5404 vdd.n15 vdd.t2 3.9605
R5405 vdd.n15 vdd.t142 3.9605
R5406 vdd.n16 vdd.t136 3.9605
R5407 vdd.n16 vdd.t137 3.9605
R5408 vdd.n18 vdd.t49 3.9605
R5409 vdd.n18 vdd.t143 3.9605
R5410 vdd.n25 vdd.t1 3.9605
R5411 vdd.n25 vdd.t139 3.9605
R5412 vdd.n7 vdd.t273 3.61217
R5413 vdd.n7 vdd.t244 3.61217
R5414 vdd.n8 vdd.t252 3.61217
R5415 vdd.n8 vdd.t265 3.61217
R5416 vdd.n10 vdd.t236 3.61217
R5417 vdd.n10 vdd.t234 3.61217
R5418 vdd.n12 vdd.t241 3.61217
R5419 vdd.n12 vdd.t257 3.61217
R5420 vdd.n5 vdd.t267 3.61217
R5421 vdd.n5 vdd.t254 3.61217
R5422 vdd.n3 vdd.t246 3.61217
R5423 vdd.n3 vdd.t269 3.61217
R5424 vdd.n1 vdd.t275 3.61217
R5425 vdd.n1 vdd.t259 3.61217
R5426 vdd.n0 vdd.t263 3.61217
R5427 vdd.n0 vdd.t249 3.61217
R5428 vdd.n316 vdd.n315 3.49141
R5429 vdd.n257 vdd.n256 3.49141
R5430 vdd.n214 vdd.n213 3.49141
R5431 vdd.n155 vdd.n154 3.49141
R5432 vdd.n113 vdd.n112 3.49141
R5433 vdd.n54 vdd.n53 3.49141
R5434 vdd.n1735 vdd.n1734 3.49141
R5435 vdd.n1794 vdd.n1793 3.49141
R5436 vdd.n1633 vdd.n1632 3.49141
R5437 vdd.n1692 vdd.n1691 3.49141
R5438 vdd.n1532 vdd.n1531 3.49141
R5439 vdd.n1591 vdd.n1590 3.49141
R5440 vdd.n2156 vdd.t245 3.40145
R5441 vdd.n2604 vdd.t266 3.40145
R5442 vdd.n2857 vdd.t256 3.40145
R5443 vdd.n2781 vdd.t233 3.40145
R5444 vdd.n1876 vdd.t227 3.28809
R5445 vdd.n3247 vdd.t20 3.28809
R5446 vdd.n2257 vdd.t262 3.17472
R5447 vdd.n2760 vdd.t243 3.17472
R5448 vdd.t50 vdd.n1104 3.06136
R5449 vdd.n3272 vdd.t18 3.06136
R5450 vdd.n1834 vdd.t59 2.83463
R5451 vdd.n644 vdd.t3 2.83463
R5452 vdd.n319 vdd.n298 2.71565
R5453 vdd.n260 vdd.n239 2.71565
R5454 vdd.n217 vdd.n196 2.71565
R5455 vdd.n158 vdd.n137 2.71565
R5456 vdd.n116 vdd.n95 2.71565
R5457 vdd.n57 vdd.n36 2.71565
R5458 vdd.n1738 vdd.n1717 2.71565
R5459 vdd.n1797 vdd.n1776 2.71565
R5460 vdd.n1636 vdd.n1615 2.71565
R5461 vdd.n1695 vdd.n1674 2.71565
R5462 vdd.n1535 vdd.n1514 2.71565
R5463 vdd.n1594 vdd.n1573 2.71565
R5464 vdd.t43 vdd.n1132 2.6079
R5465 vdd.n2406 vdd.t242 2.6079
R5466 vdd.n2430 vdd.t250 2.6079
R5467 vdd.n2894 vdd.t261 2.6079
R5468 vdd.n2918 vdd.t247 2.6079
R5469 vdd.n3395 vdd.t7 2.6079
R5470 vdd.n2924 vdd.n2923 2.49806
R5471 vdd.n2398 vdd.n2397 2.49806
R5472 vdd.n306 vdd.n305 2.4129
R5473 vdd.n247 vdd.n246 2.4129
R5474 vdd.n204 vdd.n203 2.4129
R5475 vdd.n145 vdd.n144 2.4129
R5476 vdd.n103 vdd.n102 2.4129
R5477 vdd.n44 vdd.n43 2.4129
R5478 vdd.n1725 vdd.n1724 2.4129
R5479 vdd.n1784 vdd.n1783 2.4129
R5480 vdd.n1623 vdd.n1622 2.4129
R5481 vdd.n1682 vdd.n1681 2.4129
R5482 vdd.n1522 vdd.n1521 2.4129
R5483 vdd.n1581 vdd.n1580 2.4129
R5484 vdd.n1486 vdd.t28 2.38117
R5485 vdd.n1894 vdd.t152 2.38117
R5486 vdd.n3231 vdd.t145 2.38117
R5487 vdd.n3386 vdd.t24 2.38117
R5488 vdd.n2315 vdd.n1904 2.27742
R5489 vdd.n2316 vdd.n2315 2.27742
R5490 vdd.n3216 vdd.n3215 2.27742
R5491 vdd.n3217 vdd.n3216 2.27742
R5492 vdd.n3094 vdd.n3093 2.27742
R5493 vdd.n3093 vdd.n784 2.27742
R5494 vdd.n2338 vdd.n1065 2.27742
R5495 vdd.n2338 vdd.n1066 2.27742
R5496 vdd.n2430 vdd.t274 2.2678
R5497 vdd.n2894 vdd.t264 2.2678
R5498 vdd.t41 vdd.n1161 2.15444
R5499 vdd.n3377 vdd.t125 2.15444
R5500 vdd.t258 vdd.n983 2.04107
R5501 vdd.n900 vdd.t251 2.04107
R5502 vdd.n320 vdd.n296 1.93989
R5503 vdd.n261 vdd.n237 1.93989
R5504 vdd.n218 vdd.n194 1.93989
R5505 vdd.n159 vdd.n135 1.93989
R5506 vdd.n117 vdd.n93 1.93989
R5507 vdd.n58 vdd.n34 1.93989
R5508 vdd.n1739 vdd.n1715 1.93989
R5509 vdd.n1798 vdd.n1774 1.93989
R5510 vdd.n1637 vdd.n1613 1.93989
R5511 vdd.n1696 vdd.n1672 1.93989
R5512 vdd.n1536 vdd.n1512 1.93989
R5513 vdd.n1595 vdd.n1571 1.93989
R5514 vdd.n1444 vdd.t52 1.92771
R5515 vdd.n2381 vdd.t195 1.92771
R5516 vdd.n2457 vdd.t180 1.92771
R5517 vdd.n2870 vdd.t188 1.92771
R5518 vdd.n2989 vdd.t184 1.92771
R5519 vdd.t103 vdd.n375 1.92771
R5520 vdd.n1452 vdd.t54 1.70098
R5521 vdd.n2257 vdd.t270 1.70098
R5522 vdd.n1008 vdd.t239 1.70098
R5523 vdd.t255 vdd.n874 1.70098
R5524 vdd.n2760 vdd.t260 1.70098
R5525 vdd.n3371 vdd.t30 1.70098
R5526 vdd.n1477 vdd.t26 1.47425
R5527 vdd.n361 vdd.t37 1.47425
R5528 vdd.n1143 vdd.t115 1.24752
R5529 vdd.t64 vdd.n3393 1.24752
R5530 vdd.n331 vdd.n291 1.16414
R5531 vdd.n324 vdd.n323 1.16414
R5532 vdd.n272 vdd.n232 1.16414
R5533 vdd.n265 vdd.n264 1.16414
R5534 vdd.n229 vdd.n189 1.16414
R5535 vdd.n222 vdd.n221 1.16414
R5536 vdd.n170 vdd.n130 1.16414
R5537 vdd.n163 vdd.n162 1.16414
R5538 vdd.n128 vdd.n88 1.16414
R5539 vdd.n121 vdd.n120 1.16414
R5540 vdd.n69 vdd.n29 1.16414
R5541 vdd.n62 vdd.n61 1.16414
R5542 vdd.n1750 vdd.n1710 1.16414
R5543 vdd.n1743 vdd.n1742 1.16414
R5544 vdd.n1809 vdd.n1769 1.16414
R5545 vdd.n1802 vdd.n1801 1.16414
R5546 vdd.n1648 vdd.n1608 1.16414
R5547 vdd.n1641 vdd.n1640 1.16414
R5548 vdd.n1707 vdd.n1667 1.16414
R5549 vdd.n1700 vdd.n1699 1.16414
R5550 vdd.n1547 vdd.n1507 1.16414
R5551 vdd.n1540 vdd.n1539 1.16414
R5552 vdd.n1606 vdd.n1566 1.16414
R5553 vdd.n1599 vdd.n1598 1.16414
R5554 vdd.n2424 vdd.t248 1.13415
R5555 vdd.n2900 vdd.t272 1.13415
R5556 vdd.n1826 vdd.t76 1.02079
R5557 vdd.t199 vdd.t238 1.02079
R5558 vdd.t237 vdd.t156 1.02079
R5559 vdd.t16 vdd.n633 1.02079
R5560 vdd.n1323 vdd.n1319 0.970197
R5561 vdd.n2336 vdd.n2335 0.970197
R5562 vdd.n618 vdd.n428 0.970197
R5563 vdd.n3095 vdd.n690 0.970197
R5564 vdd.n1812 vdd.n28 0.90431
R5565 vdd vdd.n3400 0.896477
R5566 vdd.n1842 vdd.t67 0.794056
R5567 vdd.n2400 vdd.t238 0.794056
R5568 vdd.n2436 vdd.t271 0.794056
R5569 vdd.n2888 vdd.t232 0.794056
R5570 vdd.n2926 vdd.t237 0.794056
R5571 vdd.n3281 vdd.t99 0.794056
R5572 vdd.n1867 vdd.t5 0.567326
R5573 vdd.t72 vdd.n662 0.567326
R5574 vdd.n2326 vdd.n2325 0.530988
R5575 vdd.n726 vdd.n682 0.530988
R5576 vdd.n464 vdd.n391 0.530988
R5577 vdd.n3350 vdd.n3349 0.530988
R5578 vdd.n3227 vdd.n3226 0.530988
R5579 vdd.n1889 vdd.n1067 0.530988
R5580 vdd.n1321 vdd.n1186 0.530988
R5581 vdd.n1423 vdd.n1422 0.530988
R5582 vdd.n4 vdd.n2 0.459552
R5583 vdd.n11 vdd.n9 0.459552
R5584 vdd.n329 vdd.n328 0.388379
R5585 vdd.n295 vdd.n293 0.388379
R5586 vdd.n270 vdd.n269 0.388379
R5587 vdd.n236 vdd.n234 0.388379
R5588 vdd.n227 vdd.n226 0.388379
R5589 vdd.n193 vdd.n191 0.388379
R5590 vdd.n168 vdd.n167 0.388379
R5591 vdd.n134 vdd.n132 0.388379
R5592 vdd.n126 vdd.n125 0.388379
R5593 vdd.n92 vdd.n90 0.388379
R5594 vdd.n67 vdd.n66 0.388379
R5595 vdd.n33 vdd.n31 0.388379
R5596 vdd.n1748 vdd.n1747 0.388379
R5597 vdd.n1714 vdd.n1712 0.388379
R5598 vdd.n1807 vdd.n1806 0.388379
R5599 vdd.n1773 vdd.n1771 0.388379
R5600 vdd.n1646 vdd.n1645 0.388379
R5601 vdd.n1612 vdd.n1610 0.388379
R5602 vdd.n1705 vdd.n1704 0.388379
R5603 vdd.n1671 vdd.n1669 0.388379
R5604 vdd.n1545 vdd.n1544 0.388379
R5605 vdd.n1511 vdd.n1509 0.388379
R5606 vdd.n1604 vdd.n1603 0.388379
R5607 vdd.n1570 vdd.n1568 0.388379
R5608 vdd.n19 vdd.n17 0.387128
R5609 vdd.n24 vdd.n22 0.387128
R5610 vdd.n6 vdd.n4 0.358259
R5611 vdd.n13 vdd.n11 0.358259
R5612 vdd.n276 vdd.n274 0.358259
R5613 vdd.n278 vdd.n276 0.358259
R5614 vdd.n280 vdd.n278 0.358259
R5615 vdd.n282 vdd.n280 0.358259
R5616 vdd.n284 vdd.n282 0.358259
R5617 vdd.n286 vdd.n284 0.358259
R5618 vdd.n288 vdd.n286 0.358259
R5619 vdd.n290 vdd.n288 0.358259
R5620 vdd.n332 vdd.n290 0.358259
R5621 vdd.n174 vdd.n172 0.358259
R5622 vdd.n176 vdd.n174 0.358259
R5623 vdd.n178 vdd.n176 0.358259
R5624 vdd.n180 vdd.n178 0.358259
R5625 vdd.n182 vdd.n180 0.358259
R5626 vdd.n184 vdd.n182 0.358259
R5627 vdd.n186 vdd.n184 0.358259
R5628 vdd.n188 vdd.n186 0.358259
R5629 vdd.n230 vdd.n188 0.358259
R5630 vdd.n73 vdd.n71 0.358259
R5631 vdd.n75 vdd.n73 0.358259
R5632 vdd.n77 vdd.n75 0.358259
R5633 vdd.n79 vdd.n77 0.358259
R5634 vdd.n81 vdd.n79 0.358259
R5635 vdd.n83 vdd.n81 0.358259
R5636 vdd.n85 vdd.n83 0.358259
R5637 vdd.n87 vdd.n85 0.358259
R5638 vdd.n129 vdd.n87 0.358259
R5639 vdd.n1810 vdd.n1768 0.358259
R5640 vdd.n1768 vdd.n1766 0.358259
R5641 vdd.n1766 vdd.n1764 0.358259
R5642 vdd.n1764 vdd.n1762 0.358259
R5643 vdd.n1762 vdd.n1760 0.358259
R5644 vdd.n1760 vdd.n1758 0.358259
R5645 vdd.n1758 vdd.n1756 0.358259
R5646 vdd.n1756 vdd.n1754 0.358259
R5647 vdd.n1754 vdd.n1752 0.358259
R5648 vdd.n1708 vdd.n1666 0.358259
R5649 vdd.n1666 vdd.n1664 0.358259
R5650 vdd.n1664 vdd.n1662 0.358259
R5651 vdd.n1662 vdd.n1660 0.358259
R5652 vdd.n1660 vdd.n1658 0.358259
R5653 vdd.n1658 vdd.n1656 0.358259
R5654 vdd.n1656 vdd.n1654 0.358259
R5655 vdd.n1654 vdd.n1652 0.358259
R5656 vdd.n1652 vdd.n1650 0.358259
R5657 vdd.n1607 vdd.n1565 0.358259
R5658 vdd.n1565 vdd.n1563 0.358259
R5659 vdd.n1563 vdd.n1561 0.358259
R5660 vdd.n1561 vdd.n1559 0.358259
R5661 vdd.n1559 vdd.n1557 0.358259
R5662 vdd.n1557 vdd.n1555 0.358259
R5663 vdd.n1555 vdd.n1553 0.358259
R5664 vdd.n1553 vdd.n1551 0.358259
R5665 vdd.n1551 vdd.n1549 0.358259
R5666 vdd.n14 vdd.n6 0.334552
R5667 vdd.n14 vdd.n13 0.334552
R5668 vdd.n27 vdd.n19 0.21707
R5669 vdd.n27 vdd.n24 0.21707
R5670 vdd.n330 vdd.n292 0.155672
R5671 vdd.n322 vdd.n292 0.155672
R5672 vdd.n322 vdd.n321 0.155672
R5673 vdd.n321 vdd.n297 0.155672
R5674 vdd.n314 vdd.n297 0.155672
R5675 vdd.n314 vdd.n313 0.155672
R5676 vdd.n313 vdd.n301 0.155672
R5677 vdd.n306 vdd.n301 0.155672
R5678 vdd.n271 vdd.n233 0.155672
R5679 vdd.n263 vdd.n233 0.155672
R5680 vdd.n263 vdd.n262 0.155672
R5681 vdd.n262 vdd.n238 0.155672
R5682 vdd.n255 vdd.n238 0.155672
R5683 vdd.n255 vdd.n254 0.155672
R5684 vdd.n254 vdd.n242 0.155672
R5685 vdd.n247 vdd.n242 0.155672
R5686 vdd.n228 vdd.n190 0.155672
R5687 vdd.n220 vdd.n190 0.155672
R5688 vdd.n220 vdd.n219 0.155672
R5689 vdd.n219 vdd.n195 0.155672
R5690 vdd.n212 vdd.n195 0.155672
R5691 vdd.n212 vdd.n211 0.155672
R5692 vdd.n211 vdd.n199 0.155672
R5693 vdd.n204 vdd.n199 0.155672
R5694 vdd.n169 vdd.n131 0.155672
R5695 vdd.n161 vdd.n131 0.155672
R5696 vdd.n161 vdd.n160 0.155672
R5697 vdd.n160 vdd.n136 0.155672
R5698 vdd.n153 vdd.n136 0.155672
R5699 vdd.n153 vdd.n152 0.155672
R5700 vdd.n152 vdd.n140 0.155672
R5701 vdd.n145 vdd.n140 0.155672
R5702 vdd.n127 vdd.n89 0.155672
R5703 vdd.n119 vdd.n89 0.155672
R5704 vdd.n119 vdd.n118 0.155672
R5705 vdd.n118 vdd.n94 0.155672
R5706 vdd.n111 vdd.n94 0.155672
R5707 vdd.n111 vdd.n110 0.155672
R5708 vdd.n110 vdd.n98 0.155672
R5709 vdd.n103 vdd.n98 0.155672
R5710 vdd.n68 vdd.n30 0.155672
R5711 vdd.n60 vdd.n30 0.155672
R5712 vdd.n60 vdd.n59 0.155672
R5713 vdd.n59 vdd.n35 0.155672
R5714 vdd.n52 vdd.n35 0.155672
R5715 vdd.n52 vdd.n51 0.155672
R5716 vdd.n51 vdd.n39 0.155672
R5717 vdd.n44 vdd.n39 0.155672
R5718 vdd.n1749 vdd.n1711 0.155672
R5719 vdd.n1741 vdd.n1711 0.155672
R5720 vdd.n1741 vdd.n1740 0.155672
R5721 vdd.n1740 vdd.n1716 0.155672
R5722 vdd.n1733 vdd.n1716 0.155672
R5723 vdd.n1733 vdd.n1732 0.155672
R5724 vdd.n1732 vdd.n1720 0.155672
R5725 vdd.n1725 vdd.n1720 0.155672
R5726 vdd.n1808 vdd.n1770 0.155672
R5727 vdd.n1800 vdd.n1770 0.155672
R5728 vdd.n1800 vdd.n1799 0.155672
R5729 vdd.n1799 vdd.n1775 0.155672
R5730 vdd.n1792 vdd.n1775 0.155672
R5731 vdd.n1792 vdd.n1791 0.155672
R5732 vdd.n1791 vdd.n1779 0.155672
R5733 vdd.n1784 vdd.n1779 0.155672
R5734 vdd.n1647 vdd.n1609 0.155672
R5735 vdd.n1639 vdd.n1609 0.155672
R5736 vdd.n1639 vdd.n1638 0.155672
R5737 vdd.n1638 vdd.n1614 0.155672
R5738 vdd.n1631 vdd.n1614 0.155672
R5739 vdd.n1631 vdd.n1630 0.155672
R5740 vdd.n1630 vdd.n1618 0.155672
R5741 vdd.n1623 vdd.n1618 0.155672
R5742 vdd.n1706 vdd.n1668 0.155672
R5743 vdd.n1698 vdd.n1668 0.155672
R5744 vdd.n1698 vdd.n1697 0.155672
R5745 vdd.n1697 vdd.n1673 0.155672
R5746 vdd.n1690 vdd.n1673 0.155672
R5747 vdd.n1690 vdd.n1689 0.155672
R5748 vdd.n1689 vdd.n1677 0.155672
R5749 vdd.n1682 vdd.n1677 0.155672
R5750 vdd.n1546 vdd.n1508 0.155672
R5751 vdd.n1538 vdd.n1508 0.155672
R5752 vdd.n1538 vdd.n1537 0.155672
R5753 vdd.n1537 vdd.n1513 0.155672
R5754 vdd.n1530 vdd.n1513 0.155672
R5755 vdd.n1530 vdd.n1529 0.155672
R5756 vdd.n1529 vdd.n1517 0.155672
R5757 vdd.n1522 vdd.n1517 0.155672
R5758 vdd.n1605 vdd.n1567 0.155672
R5759 vdd.n1597 vdd.n1567 0.155672
R5760 vdd.n1597 vdd.n1596 0.155672
R5761 vdd.n1596 vdd.n1572 0.155672
R5762 vdd.n1589 vdd.n1572 0.155672
R5763 vdd.n1589 vdd.n1588 0.155672
R5764 vdd.n1588 vdd.n1576 0.155672
R5765 vdd.n1581 vdd.n1576 0.155672
R5766 vdd.n2101 vdd.n1906 0.152939
R5767 vdd.n1912 vdd.n1906 0.152939
R5768 vdd.n1913 vdd.n1912 0.152939
R5769 vdd.n1914 vdd.n1913 0.152939
R5770 vdd.n1915 vdd.n1914 0.152939
R5771 vdd.n1919 vdd.n1915 0.152939
R5772 vdd.n1920 vdd.n1919 0.152939
R5773 vdd.n1921 vdd.n1920 0.152939
R5774 vdd.n1922 vdd.n1921 0.152939
R5775 vdd.n1926 vdd.n1922 0.152939
R5776 vdd.n1927 vdd.n1926 0.152939
R5777 vdd.n1928 vdd.n1927 0.152939
R5778 vdd.n2076 vdd.n1928 0.152939
R5779 vdd.n2076 vdd.n2075 0.152939
R5780 vdd.n2075 vdd.n2074 0.152939
R5781 vdd.n2074 vdd.n1934 0.152939
R5782 vdd.n1939 vdd.n1934 0.152939
R5783 vdd.n1940 vdd.n1939 0.152939
R5784 vdd.n1941 vdd.n1940 0.152939
R5785 vdd.n1945 vdd.n1941 0.152939
R5786 vdd.n1946 vdd.n1945 0.152939
R5787 vdd.n1947 vdd.n1946 0.152939
R5788 vdd.n1948 vdd.n1947 0.152939
R5789 vdd.n1952 vdd.n1948 0.152939
R5790 vdd.n1953 vdd.n1952 0.152939
R5791 vdd.n1954 vdd.n1953 0.152939
R5792 vdd.n1955 vdd.n1954 0.152939
R5793 vdd.n1959 vdd.n1955 0.152939
R5794 vdd.n1960 vdd.n1959 0.152939
R5795 vdd.n1961 vdd.n1960 0.152939
R5796 vdd.n1962 vdd.n1961 0.152939
R5797 vdd.n1966 vdd.n1962 0.152939
R5798 vdd.n1967 vdd.n1966 0.152939
R5799 vdd.n1968 vdd.n1967 0.152939
R5800 vdd.n2037 vdd.n1968 0.152939
R5801 vdd.n2037 vdd.n2036 0.152939
R5802 vdd.n2036 vdd.n2035 0.152939
R5803 vdd.n2035 vdd.n1974 0.152939
R5804 vdd.n1979 vdd.n1974 0.152939
R5805 vdd.n1980 vdd.n1979 0.152939
R5806 vdd.n1981 vdd.n1980 0.152939
R5807 vdd.n1985 vdd.n1981 0.152939
R5808 vdd.n1986 vdd.n1985 0.152939
R5809 vdd.n1987 vdd.n1986 0.152939
R5810 vdd.n1988 vdd.n1987 0.152939
R5811 vdd.n1992 vdd.n1988 0.152939
R5812 vdd.n1993 vdd.n1992 0.152939
R5813 vdd.n1994 vdd.n1993 0.152939
R5814 vdd.n1995 vdd.n1994 0.152939
R5815 vdd.n1996 vdd.n1995 0.152939
R5816 vdd.n1996 vdd.n1064 0.152939
R5817 vdd.n2325 vdd.n1900 0.152939
R5818 vdd.n1814 vdd.n1123 0.152939
R5819 vdd.n1829 vdd.n1123 0.152939
R5820 vdd.n1830 vdd.n1829 0.152939
R5821 vdd.n1831 vdd.n1830 0.152939
R5822 vdd.n1831 vdd.n1112 0.152939
R5823 vdd.n1846 vdd.n1112 0.152939
R5824 vdd.n1847 vdd.n1846 0.152939
R5825 vdd.n1848 vdd.n1847 0.152939
R5826 vdd.n1848 vdd.n1101 0.152939
R5827 vdd.n1862 vdd.n1101 0.152939
R5828 vdd.n1863 vdd.n1862 0.152939
R5829 vdd.n1864 vdd.n1863 0.152939
R5830 vdd.n1864 vdd.n1089 0.152939
R5831 vdd.n1879 vdd.n1089 0.152939
R5832 vdd.n1880 vdd.n1879 0.152939
R5833 vdd.n1881 vdd.n1880 0.152939
R5834 vdd.n1881 vdd.n1077 0.152939
R5835 vdd.n1898 vdd.n1077 0.152939
R5836 vdd.n1899 vdd.n1898 0.152939
R5837 vdd.n2326 vdd.n1899 0.152939
R5838 vdd.n735 vdd.n730 0.152939
R5839 vdd.n736 vdd.n735 0.152939
R5840 vdd.n737 vdd.n736 0.152939
R5841 vdd.n738 vdd.n737 0.152939
R5842 vdd.n739 vdd.n738 0.152939
R5843 vdd.n740 vdd.n739 0.152939
R5844 vdd.n741 vdd.n740 0.152939
R5845 vdd.n742 vdd.n741 0.152939
R5846 vdd.n743 vdd.n742 0.152939
R5847 vdd.n744 vdd.n743 0.152939
R5848 vdd.n745 vdd.n744 0.152939
R5849 vdd.n746 vdd.n745 0.152939
R5850 vdd.n3183 vdd.n746 0.152939
R5851 vdd.n3183 vdd.n3182 0.152939
R5852 vdd.n3182 vdd.n3181 0.152939
R5853 vdd.n3181 vdd.n748 0.152939
R5854 vdd.n749 vdd.n748 0.152939
R5855 vdd.n750 vdd.n749 0.152939
R5856 vdd.n751 vdd.n750 0.152939
R5857 vdd.n752 vdd.n751 0.152939
R5858 vdd.n753 vdd.n752 0.152939
R5859 vdd.n754 vdd.n753 0.152939
R5860 vdd.n755 vdd.n754 0.152939
R5861 vdd.n756 vdd.n755 0.152939
R5862 vdd.n757 vdd.n756 0.152939
R5863 vdd.n758 vdd.n757 0.152939
R5864 vdd.n759 vdd.n758 0.152939
R5865 vdd.n760 vdd.n759 0.152939
R5866 vdd.n761 vdd.n760 0.152939
R5867 vdd.n762 vdd.n761 0.152939
R5868 vdd.n763 vdd.n762 0.152939
R5869 vdd.n764 vdd.n763 0.152939
R5870 vdd.n765 vdd.n764 0.152939
R5871 vdd.n766 vdd.n765 0.152939
R5872 vdd.n3137 vdd.n766 0.152939
R5873 vdd.n3137 vdd.n3136 0.152939
R5874 vdd.n3136 vdd.n3135 0.152939
R5875 vdd.n3135 vdd.n770 0.152939
R5876 vdd.n771 vdd.n770 0.152939
R5877 vdd.n772 vdd.n771 0.152939
R5878 vdd.n773 vdd.n772 0.152939
R5879 vdd.n774 vdd.n773 0.152939
R5880 vdd.n775 vdd.n774 0.152939
R5881 vdd.n776 vdd.n775 0.152939
R5882 vdd.n777 vdd.n776 0.152939
R5883 vdd.n778 vdd.n777 0.152939
R5884 vdd.n779 vdd.n778 0.152939
R5885 vdd.n780 vdd.n779 0.152939
R5886 vdd.n781 vdd.n780 0.152939
R5887 vdd.n782 vdd.n781 0.152939
R5888 vdd.n783 vdd.n782 0.152939
R5889 vdd.n727 vdd.n726 0.152939
R5890 vdd.n3234 vdd.n682 0.152939
R5891 vdd.n3235 vdd.n3234 0.152939
R5892 vdd.n3236 vdd.n3235 0.152939
R5893 vdd.n3236 vdd.n670 0.152939
R5894 vdd.n3251 vdd.n670 0.152939
R5895 vdd.n3252 vdd.n3251 0.152939
R5896 vdd.n3253 vdd.n3252 0.152939
R5897 vdd.n3253 vdd.n659 0.152939
R5898 vdd.n3267 vdd.n659 0.152939
R5899 vdd.n3268 vdd.n3267 0.152939
R5900 vdd.n3269 vdd.n3268 0.152939
R5901 vdd.n3269 vdd.n647 0.152939
R5902 vdd.n3284 vdd.n647 0.152939
R5903 vdd.n3285 vdd.n3284 0.152939
R5904 vdd.n3286 vdd.n3285 0.152939
R5905 vdd.n3286 vdd.n636 0.152939
R5906 vdd.n3303 vdd.n636 0.152939
R5907 vdd.n3304 vdd.n3303 0.152939
R5908 vdd.n3305 vdd.n3304 0.152939
R5909 vdd.n3305 vdd.n334 0.152939
R5910 vdd.n3398 vdd.n335 0.152939
R5911 vdd.n346 vdd.n335 0.152939
R5912 vdd.n347 vdd.n346 0.152939
R5913 vdd.n348 vdd.n347 0.152939
R5914 vdd.n355 vdd.n348 0.152939
R5915 vdd.n356 vdd.n355 0.152939
R5916 vdd.n357 vdd.n356 0.152939
R5917 vdd.n358 vdd.n357 0.152939
R5918 vdd.n366 vdd.n358 0.152939
R5919 vdd.n367 vdd.n366 0.152939
R5920 vdd.n368 vdd.n367 0.152939
R5921 vdd.n369 vdd.n368 0.152939
R5922 vdd.n377 vdd.n369 0.152939
R5923 vdd.n378 vdd.n377 0.152939
R5924 vdd.n379 vdd.n378 0.152939
R5925 vdd.n380 vdd.n379 0.152939
R5926 vdd.n388 vdd.n380 0.152939
R5927 vdd.n389 vdd.n388 0.152939
R5928 vdd.n390 vdd.n389 0.152939
R5929 vdd.n391 vdd.n390 0.152939
R5930 vdd.n464 vdd.n463 0.152939
R5931 vdd.n470 vdd.n463 0.152939
R5932 vdd.n471 vdd.n470 0.152939
R5933 vdd.n472 vdd.n471 0.152939
R5934 vdd.n472 vdd.n461 0.152939
R5935 vdd.n480 vdd.n461 0.152939
R5936 vdd.n481 vdd.n480 0.152939
R5937 vdd.n482 vdd.n481 0.152939
R5938 vdd.n482 vdd.n459 0.152939
R5939 vdd.n490 vdd.n459 0.152939
R5940 vdd.n491 vdd.n490 0.152939
R5941 vdd.n492 vdd.n491 0.152939
R5942 vdd.n492 vdd.n457 0.152939
R5943 vdd.n500 vdd.n457 0.152939
R5944 vdd.n501 vdd.n500 0.152939
R5945 vdd.n502 vdd.n501 0.152939
R5946 vdd.n502 vdd.n455 0.152939
R5947 vdd.n510 vdd.n455 0.152939
R5948 vdd.n511 vdd.n510 0.152939
R5949 vdd.n512 vdd.n511 0.152939
R5950 vdd.n512 vdd.n451 0.152939
R5951 vdd.n520 vdd.n451 0.152939
R5952 vdd.n521 vdd.n520 0.152939
R5953 vdd.n522 vdd.n521 0.152939
R5954 vdd.n522 vdd.n449 0.152939
R5955 vdd.n530 vdd.n449 0.152939
R5956 vdd.n531 vdd.n530 0.152939
R5957 vdd.n532 vdd.n531 0.152939
R5958 vdd.n532 vdd.n447 0.152939
R5959 vdd.n540 vdd.n447 0.152939
R5960 vdd.n541 vdd.n540 0.152939
R5961 vdd.n542 vdd.n541 0.152939
R5962 vdd.n542 vdd.n445 0.152939
R5963 vdd.n550 vdd.n445 0.152939
R5964 vdd.n551 vdd.n550 0.152939
R5965 vdd.n552 vdd.n551 0.152939
R5966 vdd.n552 vdd.n443 0.152939
R5967 vdd.n560 vdd.n443 0.152939
R5968 vdd.n561 vdd.n560 0.152939
R5969 vdd.n562 vdd.n561 0.152939
R5970 vdd.n562 vdd.n439 0.152939
R5971 vdd.n570 vdd.n439 0.152939
R5972 vdd.n571 vdd.n570 0.152939
R5973 vdd.n572 vdd.n571 0.152939
R5974 vdd.n572 vdd.n437 0.152939
R5975 vdd.n580 vdd.n437 0.152939
R5976 vdd.n581 vdd.n580 0.152939
R5977 vdd.n582 vdd.n581 0.152939
R5978 vdd.n582 vdd.n435 0.152939
R5979 vdd.n590 vdd.n435 0.152939
R5980 vdd.n591 vdd.n590 0.152939
R5981 vdd.n592 vdd.n591 0.152939
R5982 vdd.n592 vdd.n433 0.152939
R5983 vdd.n600 vdd.n433 0.152939
R5984 vdd.n601 vdd.n600 0.152939
R5985 vdd.n602 vdd.n601 0.152939
R5986 vdd.n602 vdd.n431 0.152939
R5987 vdd.n610 vdd.n431 0.152939
R5988 vdd.n611 vdd.n610 0.152939
R5989 vdd.n612 vdd.n611 0.152939
R5990 vdd.n612 vdd.n429 0.152939
R5991 vdd.n619 vdd.n429 0.152939
R5992 vdd.n3350 vdd.n619 0.152939
R5993 vdd.n3228 vdd.n3227 0.152939
R5994 vdd.n3228 vdd.n675 0.152939
R5995 vdd.n3242 vdd.n675 0.152939
R5996 vdd.n3243 vdd.n3242 0.152939
R5997 vdd.n3244 vdd.n3243 0.152939
R5998 vdd.n3244 vdd.n665 0.152939
R5999 vdd.n3259 vdd.n665 0.152939
R6000 vdd.n3260 vdd.n3259 0.152939
R6001 vdd.n3261 vdd.n3260 0.152939
R6002 vdd.n3261 vdd.n652 0.152939
R6003 vdd.n3275 vdd.n652 0.152939
R6004 vdd.n3276 vdd.n3275 0.152939
R6005 vdd.n3277 vdd.n3276 0.152939
R6006 vdd.n3277 vdd.n641 0.152939
R6007 vdd.n3292 vdd.n641 0.152939
R6008 vdd.n3293 vdd.n3292 0.152939
R6009 vdd.n3294 vdd.n3293 0.152939
R6010 vdd.n3296 vdd.n3294 0.152939
R6011 vdd.n3296 vdd.n3295 0.152939
R6012 vdd.n3295 vdd.n630 0.152939
R6013 vdd.n3313 vdd.n630 0.152939
R6014 vdd.n3314 vdd.n3313 0.152939
R6015 vdd.n3315 vdd.n3314 0.152939
R6016 vdd.n3315 vdd.n628 0.152939
R6017 vdd.n3320 vdd.n628 0.152939
R6018 vdd.n3321 vdd.n3320 0.152939
R6019 vdd.n3322 vdd.n3321 0.152939
R6020 vdd.n3322 vdd.n626 0.152939
R6021 vdd.n3327 vdd.n626 0.152939
R6022 vdd.n3328 vdd.n3327 0.152939
R6023 vdd.n3329 vdd.n3328 0.152939
R6024 vdd.n3329 vdd.n624 0.152939
R6025 vdd.n3335 vdd.n624 0.152939
R6026 vdd.n3336 vdd.n3335 0.152939
R6027 vdd.n3337 vdd.n3336 0.152939
R6028 vdd.n3337 vdd.n622 0.152939
R6029 vdd.n3342 vdd.n622 0.152939
R6030 vdd.n3343 vdd.n3342 0.152939
R6031 vdd.n3344 vdd.n3343 0.152939
R6032 vdd.n3344 vdd.n620 0.152939
R6033 vdd.n3349 vdd.n620 0.152939
R6034 vdd.n3226 vdd.n687 0.152939
R6035 vdd.n2337 vdd.n1067 0.152939
R6036 vdd.n1430 vdd.n1186 0.152939
R6037 vdd.n1431 vdd.n1430 0.152939
R6038 vdd.n1432 vdd.n1431 0.152939
R6039 vdd.n1432 vdd.n1174 0.152939
R6040 vdd.n1447 vdd.n1174 0.152939
R6041 vdd.n1448 vdd.n1447 0.152939
R6042 vdd.n1449 vdd.n1448 0.152939
R6043 vdd.n1449 vdd.n1164 0.152939
R6044 vdd.n1464 vdd.n1164 0.152939
R6045 vdd.n1465 vdd.n1464 0.152939
R6046 vdd.n1466 vdd.n1465 0.152939
R6047 vdd.n1466 vdd.n1151 0.152939
R6048 vdd.n1480 vdd.n1151 0.152939
R6049 vdd.n1481 vdd.n1480 0.152939
R6050 vdd.n1482 vdd.n1481 0.152939
R6051 vdd.n1482 vdd.n1140 0.152939
R6052 vdd.n1497 vdd.n1140 0.152939
R6053 vdd.n1498 vdd.n1497 0.152939
R6054 vdd.n1499 vdd.n1498 0.152939
R6055 vdd.n1499 vdd.n1129 0.152939
R6056 vdd.n1820 vdd.n1129 0.152939
R6057 vdd.n1821 vdd.n1820 0.152939
R6058 vdd.n1822 vdd.n1821 0.152939
R6059 vdd.n1822 vdd.n1117 0.152939
R6060 vdd.n1837 vdd.n1117 0.152939
R6061 vdd.n1838 vdd.n1837 0.152939
R6062 vdd.n1839 vdd.n1838 0.152939
R6063 vdd.n1839 vdd.n1107 0.152939
R6064 vdd.n1854 vdd.n1107 0.152939
R6065 vdd.n1855 vdd.n1854 0.152939
R6066 vdd.n1856 vdd.n1855 0.152939
R6067 vdd.n1856 vdd.n1094 0.152939
R6068 vdd.n1870 vdd.n1094 0.152939
R6069 vdd.n1871 vdd.n1870 0.152939
R6070 vdd.n1872 vdd.n1871 0.152939
R6071 vdd.n1872 vdd.n1084 0.152939
R6072 vdd.n1887 vdd.n1084 0.152939
R6073 vdd.n1888 vdd.n1887 0.152939
R6074 vdd.n1891 vdd.n1888 0.152939
R6075 vdd.n1891 vdd.n1890 0.152939
R6076 vdd.n1890 vdd.n1889 0.152939
R6077 vdd.n1422 vdd.n1191 0.152939
R6078 vdd.n1415 vdd.n1191 0.152939
R6079 vdd.n1415 vdd.n1414 0.152939
R6080 vdd.n1414 vdd.n1413 0.152939
R6081 vdd.n1413 vdd.n1228 0.152939
R6082 vdd.n1409 vdd.n1228 0.152939
R6083 vdd.n1409 vdd.n1408 0.152939
R6084 vdd.n1408 vdd.n1407 0.152939
R6085 vdd.n1407 vdd.n1234 0.152939
R6086 vdd.n1403 vdd.n1234 0.152939
R6087 vdd.n1403 vdd.n1402 0.152939
R6088 vdd.n1402 vdd.n1401 0.152939
R6089 vdd.n1401 vdd.n1240 0.152939
R6090 vdd.n1397 vdd.n1240 0.152939
R6091 vdd.n1397 vdd.n1396 0.152939
R6092 vdd.n1396 vdd.n1395 0.152939
R6093 vdd.n1395 vdd.n1246 0.152939
R6094 vdd.n1391 vdd.n1246 0.152939
R6095 vdd.n1391 vdd.n1390 0.152939
R6096 vdd.n1390 vdd.n1389 0.152939
R6097 vdd.n1389 vdd.n1254 0.152939
R6098 vdd.n1385 vdd.n1254 0.152939
R6099 vdd.n1385 vdd.n1384 0.152939
R6100 vdd.n1384 vdd.n1383 0.152939
R6101 vdd.n1383 vdd.n1260 0.152939
R6102 vdd.n1379 vdd.n1260 0.152939
R6103 vdd.n1379 vdd.n1378 0.152939
R6104 vdd.n1378 vdd.n1377 0.152939
R6105 vdd.n1377 vdd.n1266 0.152939
R6106 vdd.n1373 vdd.n1266 0.152939
R6107 vdd.n1373 vdd.n1372 0.152939
R6108 vdd.n1372 vdd.n1371 0.152939
R6109 vdd.n1371 vdd.n1272 0.152939
R6110 vdd.n1367 vdd.n1272 0.152939
R6111 vdd.n1367 vdd.n1366 0.152939
R6112 vdd.n1366 vdd.n1365 0.152939
R6113 vdd.n1365 vdd.n1278 0.152939
R6114 vdd.n1361 vdd.n1278 0.152939
R6115 vdd.n1361 vdd.n1360 0.152939
R6116 vdd.n1360 vdd.n1359 0.152939
R6117 vdd.n1359 vdd.n1284 0.152939
R6118 vdd.n1352 vdd.n1284 0.152939
R6119 vdd.n1352 vdd.n1351 0.152939
R6120 vdd.n1351 vdd.n1350 0.152939
R6121 vdd.n1350 vdd.n1289 0.152939
R6122 vdd.n1346 vdd.n1289 0.152939
R6123 vdd.n1346 vdd.n1345 0.152939
R6124 vdd.n1345 vdd.n1344 0.152939
R6125 vdd.n1344 vdd.n1295 0.152939
R6126 vdd.n1340 vdd.n1295 0.152939
R6127 vdd.n1340 vdd.n1339 0.152939
R6128 vdd.n1339 vdd.n1338 0.152939
R6129 vdd.n1338 vdd.n1301 0.152939
R6130 vdd.n1334 vdd.n1301 0.152939
R6131 vdd.n1334 vdd.n1333 0.152939
R6132 vdd.n1333 vdd.n1332 0.152939
R6133 vdd.n1332 vdd.n1307 0.152939
R6134 vdd.n1328 vdd.n1307 0.152939
R6135 vdd.n1328 vdd.n1327 0.152939
R6136 vdd.n1327 vdd.n1326 0.152939
R6137 vdd.n1326 vdd.n1313 0.152939
R6138 vdd.n1322 vdd.n1313 0.152939
R6139 vdd.n1322 vdd.n1321 0.152939
R6140 vdd.n1424 vdd.n1423 0.152939
R6141 vdd.n1424 vdd.n1180 0.152939
R6142 vdd.n1439 vdd.n1180 0.152939
R6143 vdd.n1440 vdd.n1439 0.152939
R6144 vdd.n1441 vdd.n1440 0.152939
R6145 vdd.n1441 vdd.n1169 0.152939
R6146 vdd.n1456 vdd.n1169 0.152939
R6147 vdd.n1457 vdd.n1456 0.152939
R6148 vdd.n1458 vdd.n1457 0.152939
R6149 vdd.n1458 vdd.n1158 0.152939
R6150 vdd.n1472 vdd.n1158 0.152939
R6151 vdd.n1473 vdd.n1472 0.152939
R6152 vdd.n1474 vdd.n1473 0.152939
R6153 vdd.n1474 vdd.n1146 0.152939
R6154 vdd.n1489 vdd.n1146 0.152939
R6155 vdd.n1490 vdd.n1489 0.152939
R6156 vdd.n1491 vdd.n1490 0.152939
R6157 vdd.n1491 vdd.n1135 0.152939
R6158 vdd.n1505 vdd.n1135 0.152939
R6159 vdd.n1506 vdd.n1505 0.152939
R6160 vdd.n1427 vdd.t160 0.113865
R6161 vdd.t167 vdd.n386 0.113865
R6162 vdd.n2315 vdd.n1900 0.110256
R6163 vdd.n3216 vdd.n727 0.110256
R6164 vdd.n3093 vdd.n687 0.110256
R6165 vdd.n2338 vdd.n2337 0.110256
R6166 vdd.n1814 vdd.n1813 0.0695946
R6167 vdd.n3399 vdd.n334 0.0695946
R6168 vdd.n3399 vdd.n3398 0.0695946
R6169 vdd.n1813 vdd.n1506 0.0695946
R6170 vdd.n2315 vdd.n2101 0.0431829
R6171 vdd.n2338 vdd.n1064 0.0431829
R6172 vdd.n3216 vdd.n730 0.0431829
R6173 vdd.n3093 vdd.n783 0.0431829
R6174 vdd vdd.n28 0.00833333
R6175 a_n1986_8322.n17 a_n1986_8322.t15 74.6477
R6176 a_n1986_8322.n7 a_n1986_8322.t6 74.6477
R6177 a_n1986_8322.n1 a_n1986_8322.t7 74.6474
R6178 a_n1986_8322.n16 a_n1986_8322.t13 74.2899
R6179 a_n1986_8322.n15 a_n1986_8322.t16 74.2899
R6180 a_n1986_8322.n12 a_n1986_8322.t17 74.2899
R6181 a_n1986_8322.n4 a_n1986_8322.t4 74.2899
R6182 a_n1986_8322.n10 a_n1986_8322.t5 74.2899
R6183 a_n1986_8322.n14 a_n1986_8322.n13 70.6783
R6184 a_n1986_8322.n1 a_n1986_8322.n0 70.6783
R6185 a_n1986_8322.n3 a_n1986_8322.n2 70.6783
R6186 a_n1986_8322.n7 a_n1986_8322.n6 70.6783
R6187 a_n1986_8322.n9 a_n1986_8322.n8 70.6783
R6188 a_n1986_8322.n18 a_n1986_8322.n17 70.6782
R6189 a_n1986_8322.n11 a_n1986_8322.n10 22.7556
R6190 a_n1986_8322.n5 a_n1986_8322.t0 10.2757
R6191 a_n1986_8322.n12 a_n1986_8322.n11 6.2408
R6192 a_n1986_8322.n5 a_n1986_8322.n4 5.83671
R6193 a_n1986_8322.n11 a_n1986_8322.n5 5.3452
R6194 a_n1986_8322.n13 a_n1986_8322.t14 3.61217
R6195 a_n1986_8322.n13 a_n1986_8322.t20 3.61217
R6196 a_n1986_8322.n0 a_n1986_8322.t11 3.61217
R6197 a_n1986_8322.n0 a_n1986_8322.t10 3.61217
R6198 a_n1986_8322.n2 a_n1986_8322.t3 3.61217
R6199 a_n1986_8322.n2 a_n1986_8322.t8 3.61217
R6200 a_n1986_8322.n6 a_n1986_8322.t12 3.61217
R6201 a_n1986_8322.n6 a_n1986_8322.t9 3.61217
R6202 a_n1986_8322.n8 a_n1986_8322.t2 3.61217
R6203 a_n1986_8322.n8 a_n1986_8322.t1 3.61217
R6204 a_n1986_8322.t19 a_n1986_8322.n18 3.61217
R6205 a_n1986_8322.n18 a_n1986_8322.t18 3.61217
R6206 a_n1986_8322.n4 a_n1986_8322.n3 0.358259
R6207 a_n1986_8322.n3 a_n1986_8322.n1 0.358259
R6208 a_n1986_8322.n10 a_n1986_8322.n9 0.358259
R6209 a_n1986_8322.n9 a_n1986_8322.n7 0.358259
R6210 a_n1986_8322.n14 a_n1986_8322.n12 0.358259
R6211 a_n1986_8322.n15 a_n1986_8322.n14 0.358259
R6212 a_n1986_8322.n17 a_n1986_8322.n16 0.358259
R6213 a_n1986_8322.n16 a_n1986_8322.n15 0.101793
R6214 gnd.n7142 gnd.n546 965.481
R6215 gnd.n3808 gnd.n3807 939.716
R6216 gnd.n3715 gnd.n2334 766.379
R6217 gnd.n3718 gnd.n3717 766.379
R6218 gnd.n2957 gnd.n2860 766.379
R6219 gnd.n2953 gnd.n2858 766.379
R6220 gnd.n3806 gnd.n2356 756.769
R6221 gnd.n3709 gnd.n3708 756.769
R6222 gnd.n3050 gnd.n2767 756.769
R6223 gnd.n3048 gnd.n2770 756.769
R6224 gnd.n6720 gnd.n798 756.769
R6225 gnd.n7141 gnd.n547 756.769
R6226 gnd.n7353 gnd.n7352 756.769
R6227 gnd.n6543 gnd.n963 756.769
R6228 gnd.n7648 gnd.n129 751.963
R6229 gnd.n7806 gnd.n7805 751.963
R6230 gnd.n1337 gnd.n1284 751.963
R6231 gnd.n6217 gnd.n1339 751.963
R6232 gnd.n6462 gnd.n1113 751.963
R6233 gnd.n5558 gnd.n1111 751.963
R6234 gnd.n3875 gnd.n3810 751.963
R6235 gnd.n4195 gnd.n2333 751.963
R6236 gnd.n7803 gnd.n131 732.745
R6237 gnd.n199 gnd.n127 732.745
R6238 gnd.n6220 gnd.n6219 732.745
R6239 gnd.n6292 gnd.n1288 732.745
R6240 gnd.n6464 gnd.n1108 732.745
R6241 gnd.n2118 gnd.n1110 732.745
R6242 gnd.n4114 gnd.n3809 732.745
R6243 gnd.n4193 gnd.n3973 732.745
R6244 gnd.n5604 gnd.n1118 711.122
R6245 gnd.n6304 gnd.n1244 711.122
R6246 gnd.n5608 gnd.n1968 711.122
R6247 gnd.n6022 gnd.n1247 711.122
R6248 gnd.n6716 gnd.n798 585
R6249 gnd.n798 gnd.n797 585
R6250 gnd.n6715 gnd.n6714 585
R6251 gnd.n6714 gnd.n6713 585
R6252 gnd.n801 gnd.n800 585
R6253 gnd.n6712 gnd.n801 585
R6254 gnd.n6710 gnd.n6709 585
R6255 gnd.n6711 gnd.n6710 585
R6256 gnd.n6708 gnd.n803 585
R6257 gnd.n803 gnd.n802 585
R6258 gnd.n6707 gnd.n6706 585
R6259 gnd.n6706 gnd.n6705 585
R6260 gnd.n809 gnd.n808 585
R6261 gnd.n6704 gnd.n809 585
R6262 gnd.n6702 gnd.n6701 585
R6263 gnd.n6703 gnd.n6702 585
R6264 gnd.n6700 gnd.n811 585
R6265 gnd.n811 gnd.n810 585
R6266 gnd.n6699 gnd.n6698 585
R6267 gnd.n6698 gnd.n6697 585
R6268 gnd.n817 gnd.n816 585
R6269 gnd.n6696 gnd.n817 585
R6270 gnd.n6694 gnd.n6693 585
R6271 gnd.n6695 gnd.n6694 585
R6272 gnd.n6692 gnd.n819 585
R6273 gnd.n819 gnd.n818 585
R6274 gnd.n6691 gnd.n6690 585
R6275 gnd.n6690 gnd.n6689 585
R6276 gnd.n825 gnd.n824 585
R6277 gnd.n6688 gnd.n825 585
R6278 gnd.n6686 gnd.n6685 585
R6279 gnd.n6687 gnd.n6686 585
R6280 gnd.n6684 gnd.n827 585
R6281 gnd.n827 gnd.n826 585
R6282 gnd.n6683 gnd.n6682 585
R6283 gnd.n6682 gnd.n6681 585
R6284 gnd.n833 gnd.n832 585
R6285 gnd.n6680 gnd.n833 585
R6286 gnd.n6678 gnd.n6677 585
R6287 gnd.n6679 gnd.n6678 585
R6288 gnd.n6676 gnd.n835 585
R6289 gnd.n835 gnd.n834 585
R6290 gnd.n6675 gnd.n6674 585
R6291 gnd.n6674 gnd.n6673 585
R6292 gnd.n841 gnd.n840 585
R6293 gnd.n6672 gnd.n841 585
R6294 gnd.n6670 gnd.n6669 585
R6295 gnd.n6671 gnd.n6670 585
R6296 gnd.n6668 gnd.n843 585
R6297 gnd.n843 gnd.n842 585
R6298 gnd.n6667 gnd.n6666 585
R6299 gnd.n6666 gnd.n6665 585
R6300 gnd.n849 gnd.n848 585
R6301 gnd.n6664 gnd.n849 585
R6302 gnd.n6662 gnd.n6661 585
R6303 gnd.n6663 gnd.n6662 585
R6304 gnd.n6660 gnd.n851 585
R6305 gnd.n851 gnd.n850 585
R6306 gnd.n6659 gnd.n6658 585
R6307 gnd.n6658 gnd.n6657 585
R6308 gnd.n857 gnd.n856 585
R6309 gnd.n6656 gnd.n857 585
R6310 gnd.n6654 gnd.n6653 585
R6311 gnd.n6655 gnd.n6654 585
R6312 gnd.n6652 gnd.n859 585
R6313 gnd.n859 gnd.n858 585
R6314 gnd.n6651 gnd.n6650 585
R6315 gnd.n6650 gnd.n6649 585
R6316 gnd.n865 gnd.n864 585
R6317 gnd.n6648 gnd.n865 585
R6318 gnd.n6646 gnd.n6645 585
R6319 gnd.n6647 gnd.n6646 585
R6320 gnd.n6644 gnd.n867 585
R6321 gnd.n867 gnd.n866 585
R6322 gnd.n6643 gnd.n6642 585
R6323 gnd.n6642 gnd.n6641 585
R6324 gnd.n873 gnd.n872 585
R6325 gnd.n6640 gnd.n873 585
R6326 gnd.n6638 gnd.n6637 585
R6327 gnd.n6639 gnd.n6638 585
R6328 gnd.n6636 gnd.n875 585
R6329 gnd.n875 gnd.n874 585
R6330 gnd.n6635 gnd.n6634 585
R6331 gnd.n6634 gnd.n6633 585
R6332 gnd.n881 gnd.n880 585
R6333 gnd.n6632 gnd.n881 585
R6334 gnd.n6630 gnd.n6629 585
R6335 gnd.n6631 gnd.n6630 585
R6336 gnd.n6628 gnd.n883 585
R6337 gnd.n883 gnd.n882 585
R6338 gnd.n6627 gnd.n6626 585
R6339 gnd.n6626 gnd.n6625 585
R6340 gnd.n889 gnd.n888 585
R6341 gnd.n6624 gnd.n889 585
R6342 gnd.n6622 gnd.n6621 585
R6343 gnd.n6623 gnd.n6622 585
R6344 gnd.n6620 gnd.n891 585
R6345 gnd.n891 gnd.n890 585
R6346 gnd.n6619 gnd.n6618 585
R6347 gnd.n6618 gnd.n6617 585
R6348 gnd.n897 gnd.n896 585
R6349 gnd.n6616 gnd.n897 585
R6350 gnd.n6614 gnd.n6613 585
R6351 gnd.n6615 gnd.n6614 585
R6352 gnd.n6612 gnd.n899 585
R6353 gnd.n899 gnd.n898 585
R6354 gnd.n6611 gnd.n6610 585
R6355 gnd.n6610 gnd.n6609 585
R6356 gnd.n905 gnd.n904 585
R6357 gnd.n6608 gnd.n905 585
R6358 gnd.n6606 gnd.n6605 585
R6359 gnd.n6607 gnd.n6606 585
R6360 gnd.n6604 gnd.n907 585
R6361 gnd.n907 gnd.n906 585
R6362 gnd.n6603 gnd.n6602 585
R6363 gnd.n6602 gnd.n6601 585
R6364 gnd.n913 gnd.n912 585
R6365 gnd.n6600 gnd.n913 585
R6366 gnd.n6598 gnd.n6597 585
R6367 gnd.n6599 gnd.n6598 585
R6368 gnd.n6596 gnd.n915 585
R6369 gnd.n915 gnd.n914 585
R6370 gnd.n6595 gnd.n6594 585
R6371 gnd.n6594 gnd.n6593 585
R6372 gnd.n921 gnd.n920 585
R6373 gnd.n6592 gnd.n921 585
R6374 gnd.n6590 gnd.n6589 585
R6375 gnd.n6591 gnd.n6590 585
R6376 gnd.n6588 gnd.n923 585
R6377 gnd.n923 gnd.n922 585
R6378 gnd.n6587 gnd.n6586 585
R6379 gnd.n6586 gnd.n6585 585
R6380 gnd.n929 gnd.n928 585
R6381 gnd.n6584 gnd.n929 585
R6382 gnd.n6582 gnd.n6581 585
R6383 gnd.n6583 gnd.n6582 585
R6384 gnd.n6580 gnd.n931 585
R6385 gnd.n931 gnd.n930 585
R6386 gnd.n6579 gnd.n6578 585
R6387 gnd.n6578 gnd.n6577 585
R6388 gnd.n937 gnd.n936 585
R6389 gnd.n6576 gnd.n937 585
R6390 gnd.n6574 gnd.n6573 585
R6391 gnd.n6575 gnd.n6574 585
R6392 gnd.n6572 gnd.n939 585
R6393 gnd.n939 gnd.n938 585
R6394 gnd.n6571 gnd.n6570 585
R6395 gnd.n6570 gnd.n6569 585
R6396 gnd.n945 gnd.n944 585
R6397 gnd.n6568 gnd.n945 585
R6398 gnd.n6566 gnd.n6565 585
R6399 gnd.n6567 gnd.n6566 585
R6400 gnd.n6564 gnd.n947 585
R6401 gnd.n947 gnd.n946 585
R6402 gnd.n6563 gnd.n6562 585
R6403 gnd.n6562 gnd.n6561 585
R6404 gnd.n953 gnd.n952 585
R6405 gnd.n6560 gnd.n953 585
R6406 gnd.n6558 gnd.n6557 585
R6407 gnd.n6559 gnd.n6558 585
R6408 gnd.n6556 gnd.n955 585
R6409 gnd.n955 gnd.n954 585
R6410 gnd.n6555 gnd.n6554 585
R6411 gnd.n6554 gnd.n6553 585
R6412 gnd.n961 gnd.n960 585
R6413 gnd.n6552 gnd.n961 585
R6414 gnd.n6550 gnd.n6549 585
R6415 gnd.n6551 gnd.n6550 585
R6416 gnd.n6720 gnd.n6719 585
R6417 gnd.n6721 gnd.n6720 585
R6418 gnd.n796 gnd.n795 585
R6419 gnd.n6722 gnd.n796 585
R6420 gnd.n6725 gnd.n6724 585
R6421 gnd.n6724 gnd.n6723 585
R6422 gnd.n793 gnd.n792 585
R6423 gnd.n792 gnd.n791 585
R6424 gnd.n6730 gnd.n6729 585
R6425 gnd.n6731 gnd.n6730 585
R6426 gnd.n790 gnd.n789 585
R6427 gnd.n6732 gnd.n790 585
R6428 gnd.n6735 gnd.n6734 585
R6429 gnd.n6734 gnd.n6733 585
R6430 gnd.n787 gnd.n786 585
R6431 gnd.n786 gnd.n785 585
R6432 gnd.n6740 gnd.n6739 585
R6433 gnd.n6741 gnd.n6740 585
R6434 gnd.n784 gnd.n783 585
R6435 gnd.n6742 gnd.n784 585
R6436 gnd.n6745 gnd.n6744 585
R6437 gnd.n6744 gnd.n6743 585
R6438 gnd.n781 gnd.n780 585
R6439 gnd.n780 gnd.n779 585
R6440 gnd.n6750 gnd.n6749 585
R6441 gnd.n6751 gnd.n6750 585
R6442 gnd.n778 gnd.n777 585
R6443 gnd.n6752 gnd.n778 585
R6444 gnd.n6755 gnd.n6754 585
R6445 gnd.n6754 gnd.n6753 585
R6446 gnd.n775 gnd.n774 585
R6447 gnd.n774 gnd.n773 585
R6448 gnd.n6760 gnd.n6759 585
R6449 gnd.n6761 gnd.n6760 585
R6450 gnd.n772 gnd.n771 585
R6451 gnd.n6762 gnd.n772 585
R6452 gnd.n6765 gnd.n6764 585
R6453 gnd.n6764 gnd.n6763 585
R6454 gnd.n769 gnd.n768 585
R6455 gnd.n768 gnd.n767 585
R6456 gnd.n6770 gnd.n6769 585
R6457 gnd.n6771 gnd.n6770 585
R6458 gnd.n766 gnd.n765 585
R6459 gnd.n6772 gnd.n766 585
R6460 gnd.n6775 gnd.n6774 585
R6461 gnd.n6774 gnd.n6773 585
R6462 gnd.n763 gnd.n762 585
R6463 gnd.n762 gnd.n761 585
R6464 gnd.n6780 gnd.n6779 585
R6465 gnd.n6781 gnd.n6780 585
R6466 gnd.n760 gnd.n759 585
R6467 gnd.n6782 gnd.n760 585
R6468 gnd.n6785 gnd.n6784 585
R6469 gnd.n6784 gnd.n6783 585
R6470 gnd.n757 gnd.n756 585
R6471 gnd.n756 gnd.n755 585
R6472 gnd.n6790 gnd.n6789 585
R6473 gnd.n6791 gnd.n6790 585
R6474 gnd.n754 gnd.n753 585
R6475 gnd.n6792 gnd.n754 585
R6476 gnd.n6795 gnd.n6794 585
R6477 gnd.n6794 gnd.n6793 585
R6478 gnd.n751 gnd.n750 585
R6479 gnd.n750 gnd.n749 585
R6480 gnd.n6800 gnd.n6799 585
R6481 gnd.n6801 gnd.n6800 585
R6482 gnd.n748 gnd.n747 585
R6483 gnd.n6802 gnd.n748 585
R6484 gnd.n6805 gnd.n6804 585
R6485 gnd.n6804 gnd.n6803 585
R6486 gnd.n745 gnd.n744 585
R6487 gnd.n744 gnd.n743 585
R6488 gnd.n6810 gnd.n6809 585
R6489 gnd.n6811 gnd.n6810 585
R6490 gnd.n742 gnd.n741 585
R6491 gnd.n6812 gnd.n742 585
R6492 gnd.n6815 gnd.n6814 585
R6493 gnd.n6814 gnd.n6813 585
R6494 gnd.n739 gnd.n738 585
R6495 gnd.n738 gnd.n737 585
R6496 gnd.n6820 gnd.n6819 585
R6497 gnd.n6821 gnd.n6820 585
R6498 gnd.n736 gnd.n735 585
R6499 gnd.n6822 gnd.n736 585
R6500 gnd.n6825 gnd.n6824 585
R6501 gnd.n6824 gnd.n6823 585
R6502 gnd.n733 gnd.n732 585
R6503 gnd.n732 gnd.n731 585
R6504 gnd.n6830 gnd.n6829 585
R6505 gnd.n6831 gnd.n6830 585
R6506 gnd.n730 gnd.n729 585
R6507 gnd.n6832 gnd.n730 585
R6508 gnd.n6835 gnd.n6834 585
R6509 gnd.n6834 gnd.n6833 585
R6510 gnd.n727 gnd.n726 585
R6511 gnd.n726 gnd.n725 585
R6512 gnd.n6840 gnd.n6839 585
R6513 gnd.n6841 gnd.n6840 585
R6514 gnd.n724 gnd.n723 585
R6515 gnd.n6842 gnd.n724 585
R6516 gnd.n6845 gnd.n6844 585
R6517 gnd.n6844 gnd.n6843 585
R6518 gnd.n721 gnd.n720 585
R6519 gnd.n720 gnd.n719 585
R6520 gnd.n6850 gnd.n6849 585
R6521 gnd.n6851 gnd.n6850 585
R6522 gnd.n718 gnd.n717 585
R6523 gnd.n6852 gnd.n718 585
R6524 gnd.n6855 gnd.n6854 585
R6525 gnd.n6854 gnd.n6853 585
R6526 gnd.n715 gnd.n714 585
R6527 gnd.n714 gnd.n713 585
R6528 gnd.n6860 gnd.n6859 585
R6529 gnd.n6861 gnd.n6860 585
R6530 gnd.n712 gnd.n711 585
R6531 gnd.n6862 gnd.n712 585
R6532 gnd.n6865 gnd.n6864 585
R6533 gnd.n6864 gnd.n6863 585
R6534 gnd.n709 gnd.n708 585
R6535 gnd.n708 gnd.n707 585
R6536 gnd.n6870 gnd.n6869 585
R6537 gnd.n6871 gnd.n6870 585
R6538 gnd.n706 gnd.n705 585
R6539 gnd.n6872 gnd.n706 585
R6540 gnd.n6875 gnd.n6874 585
R6541 gnd.n6874 gnd.n6873 585
R6542 gnd.n703 gnd.n702 585
R6543 gnd.n702 gnd.n701 585
R6544 gnd.n6880 gnd.n6879 585
R6545 gnd.n6881 gnd.n6880 585
R6546 gnd.n700 gnd.n699 585
R6547 gnd.n6882 gnd.n700 585
R6548 gnd.n6885 gnd.n6884 585
R6549 gnd.n6884 gnd.n6883 585
R6550 gnd.n697 gnd.n696 585
R6551 gnd.n696 gnd.n695 585
R6552 gnd.n6890 gnd.n6889 585
R6553 gnd.n6891 gnd.n6890 585
R6554 gnd.n694 gnd.n693 585
R6555 gnd.n6892 gnd.n694 585
R6556 gnd.n6895 gnd.n6894 585
R6557 gnd.n6894 gnd.n6893 585
R6558 gnd.n691 gnd.n690 585
R6559 gnd.n690 gnd.n689 585
R6560 gnd.n6900 gnd.n6899 585
R6561 gnd.n6901 gnd.n6900 585
R6562 gnd.n688 gnd.n687 585
R6563 gnd.n6902 gnd.n688 585
R6564 gnd.n6905 gnd.n6904 585
R6565 gnd.n6904 gnd.n6903 585
R6566 gnd.n685 gnd.n684 585
R6567 gnd.n684 gnd.n683 585
R6568 gnd.n6910 gnd.n6909 585
R6569 gnd.n6911 gnd.n6910 585
R6570 gnd.n682 gnd.n681 585
R6571 gnd.n6912 gnd.n682 585
R6572 gnd.n6915 gnd.n6914 585
R6573 gnd.n6914 gnd.n6913 585
R6574 gnd.n679 gnd.n678 585
R6575 gnd.n678 gnd.n677 585
R6576 gnd.n6920 gnd.n6919 585
R6577 gnd.n6921 gnd.n6920 585
R6578 gnd.n676 gnd.n675 585
R6579 gnd.n6922 gnd.n676 585
R6580 gnd.n6925 gnd.n6924 585
R6581 gnd.n6924 gnd.n6923 585
R6582 gnd.n673 gnd.n672 585
R6583 gnd.n672 gnd.n671 585
R6584 gnd.n6930 gnd.n6929 585
R6585 gnd.n6931 gnd.n6930 585
R6586 gnd.n670 gnd.n669 585
R6587 gnd.n6932 gnd.n670 585
R6588 gnd.n6935 gnd.n6934 585
R6589 gnd.n6934 gnd.n6933 585
R6590 gnd.n667 gnd.n666 585
R6591 gnd.n666 gnd.n665 585
R6592 gnd.n6940 gnd.n6939 585
R6593 gnd.n6941 gnd.n6940 585
R6594 gnd.n664 gnd.n663 585
R6595 gnd.n6942 gnd.n664 585
R6596 gnd.n6945 gnd.n6944 585
R6597 gnd.n6944 gnd.n6943 585
R6598 gnd.n661 gnd.n660 585
R6599 gnd.n660 gnd.n659 585
R6600 gnd.n6950 gnd.n6949 585
R6601 gnd.n6951 gnd.n6950 585
R6602 gnd.n658 gnd.n657 585
R6603 gnd.n6952 gnd.n658 585
R6604 gnd.n6955 gnd.n6954 585
R6605 gnd.n6954 gnd.n6953 585
R6606 gnd.n655 gnd.n654 585
R6607 gnd.n654 gnd.n653 585
R6608 gnd.n6960 gnd.n6959 585
R6609 gnd.n6961 gnd.n6960 585
R6610 gnd.n652 gnd.n651 585
R6611 gnd.n6962 gnd.n652 585
R6612 gnd.n6965 gnd.n6964 585
R6613 gnd.n6964 gnd.n6963 585
R6614 gnd.n649 gnd.n648 585
R6615 gnd.n648 gnd.n647 585
R6616 gnd.n6970 gnd.n6969 585
R6617 gnd.n6971 gnd.n6970 585
R6618 gnd.n646 gnd.n645 585
R6619 gnd.n6972 gnd.n646 585
R6620 gnd.n6975 gnd.n6974 585
R6621 gnd.n6974 gnd.n6973 585
R6622 gnd.n643 gnd.n642 585
R6623 gnd.n642 gnd.n641 585
R6624 gnd.n6980 gnd.n6979 585
R6625 gnd.n6981 gnd.n6980 585
R6626 gnd.n640 gnd.n639 585
R6627 gnd.n6982 gnd.n640 585
R6628 gnd.n6985 gnd.n6984 585
R6629 gnd.n6984 gnd.n6983 585
R6630 gnd.n637 gnd.n636 585
R6631 gnd.n636 gnd.n635 585
R6632 gnd.n6990 gnd.n6989 585
R6633 gnd.n6991 gnd.n6990 585
R6634 gnd.n634 gnd.n633 585
R6635 gnd.n6992 gnd.n634 585
R6636 gnd.n6995 gnd.n6994 585
R6637 gnd.n6994 gnd.n6993 585
R6638 gnd.n631 gnd.n630 585
R6639 gnd.n630 gnd.n629 585
R6640 gnd.n7000 gnd.n6999 585
R6641 gnd.n7001 gnd.n7000 585
R6642 gnd.n628 gnd.n627 585
R6643 gnd.n7002 gnd.n628 585
R6644 gnd.n7005 gnd.n7004 585
R6645 gnd.n7004 gnd.n7003 585
R6646 gnd.n625 gnd.n624 585
R6647 gnd.n624 gnd.n623 585
R6648 gnd.n7010 gnd.n7009 585
R6649 gnd.n7011 gnd.n7010 585
R6650 gnd.n622 gnd.n621 585
R6651 gnd.n7012 gnd.n622 585
R6652 gnd.n7015 gnd.n7014 585
R6653 gnd.n7014 gnd.n7013 585
R6654 gnd.n619 gnd.n618 585
R6655 gnd.n618 gnd.n617 585
R6656 gnd.n7020 gnd.n7019 585
R6657 gnd.n7021 gnd.n7020 585
R6658 gnd.n616 gnd.n615 585
R6659 gnd.n7022 gnd.n616 585
R6660 gnd.n7025 gnd.n7024 585
R6661 gnd.n7024 gnd.n7023 585
R6662 gnd.n613 gnd.n612 585
R6663 gnd.n612 gnd.n611 585
R6664 gnd.n7030 gnd.n7029 585
R6665 gnd.n7031 gnd.n7030 585
R6666 gnd.n610 gnd.n609 585
R6667 gnd.n7032 gnd.n610 585
R6668 gnd.n7035 gnd.n7034 585
R6669 gnd.n7034 gnd.n7033 585
R6670 gnd.n607 gnd.n606 585
R6671 gnd.n606 gnd.n605 585
R6672 gnd.n7040 gnd.n7039 585
R6673 gnd.n7041 gnd.n7040 585
R6674 gnd.n604 gnd.n603 585
R6675 gnd.n7042 gnd.n604 585
R6676 gnd.n7045 gnd.n7044 585
R6677 gnd.n7044 gnd.n7043 585
R6678 gnd.n601 gnd.n600 585
R6679 gnd.n600 gnd.n599 585
R6680 gnd.n7050 gnd.n7049 585
R6681 gnd.n7051 gnd.n7050 585
R6682 gnd.n598 gnd.n597 585
R6683 gnd.n7052 gnd.n598 585
R6684 gnd.n7055 gnd.n7054 585
R6685 gnd.n7054 gnd.n7053 585
R6686 gnd.n595 gnd.n594 585
R6687 gnd.n594 gnd.n593 585
R6688 gnd.n7060 gnd.n7059 585
R6689 gnd.n7061 gnd.n7060 585
R6690 gnd.n592 gnd.n591 585
R6691 gnd.n7062 gnd.n592 585
R6692 gnd.n7065 gnd.n7064 585
R6693 gnd.n7064 gnd.n7063 585
R6694 gnd.n589 gnd.n588 585
R6695 gnd.n588 gnd.n587 585
R6696 gnd.n7070 gnd.n7069 585
R6697 gnd.n7071 gnd.n7070 585
R6698 gnd.n586 gnd.n585 585
R6699 gnd.n7072 gnd.n586 585
R6700 gnd.n7075 gnd.n7074 585
R6701 gnd.n7074 gnd.n7073 585
R6702 gnd.n583 gnd.n582 585
R6703 gnd.n582 gnd.n581 585
R6704 gnd.n7080 gnd.n7079 585
R6705 gnd.n7081 gnd.n7080 585
R6706 gnd.n580 gnd.n579 585
R6707 gnd.n7082 gnd.n580 585
R6708 gnd.n7085 gnd.n7084 585
R6709 gnd.n7084 gnd.n7083 585
R6710 gnd.n577 gnd.n576 585
R6711 gnd.n576 gnd.n575 585
R6712 gnd.n7090 gnd.n7089 585
R6713 gnd.n7091 gnd.n7090 585
R6714 gnd.n574 gnd.n573 585
R6715 gnd.n7092 gnd.n574 585
R6716 gnd.n7095 gnd.n7094 585
R6717 gnd.n7094 gnd.n7093 585
R6718 gnd.n571 gnd.n570 585
R6719 gnd.n570 gnd.n569 585
R6720 gnd.n7100 gnd.n7099 585
R6721 gnd.n7101 gnd.n7100 585
R6722 gnd.n568 gnd.n567 585
R6723 gnd.n7102 gnd.n568 585
R6724 gnd.n7105 gnd.n7104 585
R6725 gnd.n7104 gnd.n7103 585
R6726 gnd.n565 gnd.n564 585
R6727 gnd.n564 gnd.n563 585
R6728 gnd.n7110 gnd.n7109 585
R6729 gnd.n7111 gnd.n7110 585
R6730 gnd.n562 gnd.n561 585
R6731 gnd.n7112 gnd.n562 585
R6732 gnd.n7115 gnd.n7114 585
R6733 gnd.n7114 gnd.n7113 585
R6734 gnd.n559 gnd.n558 585
R6735 gnd.n558 gnd.n557 585
R6736 gnd.n7120 gnd.n7119 585
R6737 gnd.n7121 gnd.n7120 585
R6738 gnd.n556 gnd.n555 585
R6739 gnd.n7122 gnd.n556 585
R6740 gnd.n7125 gnd.n7124 585
R6741 gnd.n7124 gnd.n7123 585
R6742 gnd.n553 gnd.n552 585
R6743 gnd.n552 gnd.n551 585
R6744 gnd.n7131 gnd.n7130 585
R6745 gnd.n7132 gnd.n7131 585
R6746 gnd.n550 gnd.n549 585
R6747 gnd.n7133 gnd.n550 585
R6748 gnd.n7136 gnd.n7135 585
R6749 gnd.n7135 gnd.n7134 585
R6750 gnd.n7137 gnd.n547 585
R6751 gnd.n547 gnd.n546 585
R6752 gnd.n422 gnd.n421 585
R6753 gnd.n7344 gnd.n421 585
R6754 gnd.n7347 gnd.n7346 585
R6755 gnd.n7346 gnd.n7345 585
R6756 gnd.n425 gnd.n424 585
R6757 gnd.n7343 gnd.n425 585
R6758 gnd.n7341 gnd.n7340 585
R6759 gnd.n7342 gnd.n7341 585
R6760 gnd.n428 gnd.n427 585
R6761 gnd.n427 gnd.n426 585
R6762 gnd.n7336 gnd.n7335 585
R6763 gnd.n7335 gnd.n7334 585
R6764 gnd.n431 gnd.n430 585
R6765 gnd.n7333 gnd.n431 585
R6766 gnd.n7331 gnd.n7330 585
R6767 gnd.n7332 gnd.n7331 585
R6768 gnd.n434 gnd.n433 585
R6769 gnd.n433 gnd.n432 585
R6770 gnd.n7326 gnd.n7325 585
R6771 gnd.n7325 gnd.n7324 585
R6772 gnd.n437 gnd.n436 585
R6773 gnd.n7323 gnd.n437 585
R6774 gnd.n7321 gnd.n7320 585
R6775 gnd.n7322 gnd.n7321 585
R6776 gnd.n440 gnd.n439 585
R6777 gnd.n439 gnd.n438 585
R6778 gnd.n7316 gnd.n7315 585
R6779 gnd.n7315 gnd.n7314 585
R6780 gnd.n443 gnd.n442 585
R6781 gnd.n7313 gnd.n443 585
R6782 gnd.n7311 gnd.n7310 585
R6783 gnd.n7312 gnd.n7311 585
R6784 gnd.n446 gnd.n445 585
R6785 gnd.n445 gnd.n444 585
R6786 gnd.n7306 gnd.n7305 585
R6787 gnd.n7305 gnd.n7304 585
R6788 gnd.n449 gnd.n448 585
R6789 gnd.n7303 gnd.n449 585
R6790 gnd.n7301 gnd.n7300 585
R6791 gnd.n7302 gnd.n7301 585
R6792 gnd.n452 gnd.n451 585
R6793 gnd.n451 gnd.n450 585
R6794 gnd.n7296 gnd.n7295 585
R6795 gnd.n7295 gnd.n7294 585
R6796 gnd.n455 gnd.n454 585
R6797 gnd.n7293 gnd.n455 585
R6798 gnd.n7291 gnd.n7290 585
R6799 gnd.n7292 gnd.n7291 585
R6800 gnd.n458 gnd.n457 585
R6801 gnd.n457 gnd.n456 585
R6802 gnd.n7286 gnd.n7285 585
R6803 gnd.n7285 gnd.n7284 585
R6804 gnd.n461 gnd.n460 585
R6805 gnd.n7283 gnd.n461 585
R6806 gnd.n7281 gnd.n7280 585
R6807 gnd.n7282 gnd.n7281 585
R6808 gnd.n464 gnd.n463 585
R6809 gnd.n463 gnd.n462 585
R6810 gnd.n7276 gnd.n7275 585
R6811 gnd.n7275 gnd.n7274 585
R6812 gnd.n467 gnd.n466 585
R6813 gnd.n7273 gnd.n467 585
R6814 gnd.n7271 gnd.n7270 585
R6815 gnd.n7272 gnd.n7271 585
R6816 gnd.n470 gnd.n469 585
R6817 gnd.n469 gnd.n468 585
R6818 gnd.n7266 gnd.n7265 585
R6819 gnd.n7265 gnd.n7264 585
R6820 gnd.n473 gnd.n472 585
R6821 gnd.n7263 gnd.n473 585
R6822 gnd.n7261 gnd.n7260 585
R6823 gnd.n7262 gnd.n7261 585
R6824 gnd.n476 gnd.n475 585
R6825 gnd.n475 gnd.n474 585
R6826 gnd.n7256 gnd.n7255 585
R6827 gnd.n7255 gnd.n7254 585
R6828 gnd.n479 gnd.n478 585
R6829 gnd.n7253 gnd.n479 585
R6830 gnd.n7251 gnd.n7250 585
R6831 gnd.n7252 gnd.n7251 585
R6832 gnd.n482 gnd.n481 585
R6833 gnd.n481 gnd.n480 585
R6834 gnd.n7246 gnd.n7245 585
R6835 gnd.n7245 gnd.n7244 585
R6836 gnd.n485 gnd.n484 585
R6837 gnd.n7243 gnd.n485 585
R6838 gnd.n7241 gnd.n7240 585
R6839 gnd.n7242 gnd.n7241 585
R6840 gnd.n488 gnd.n487 585
R6841 gnd.n487 gnd.n486 585
R6842 gnd.n7236 gnd.n7235 585
R6843 gnd.n7235 gnd.n7234 585
R6844 gnd.n491 gnd.n490 585
R6845 gnd.n7233 gnd.n491 585
R6846 gnd.n7231 gnd.n7230 585
R6847 gnd.n7232 gnd.n7231 585
R6848 gnd.n494 gnd.n493 585
R6849 gnd.n493 gnd.n492 585
R6850 gnd.n7226 gnd.n7225 585
R6851 gnd.n7225 gnd.n7224 585
R6852 gnd.n497 gnd.n496 585
R6853 gnd.n7223 gnd.n497 585
R6854 gnd.n7221 gnd.n7220 585
R6855 gnd.n7222 gnd.n7221 585
R6856 gnd.n500 gnd.n499 585
R6857 gnd.n499 gnd.n498 585
R6858 gnd.n7216 gnd.n7215 585
R6859 gnd.n7215 gnd.n7214 585
R6860 gnd.n503 gnd.n502 585
R6861 gnd.n7213 gnd.n503 585
R6862 gnd.n7211 gnd.n7210 585
R6863 gnd.n7212 gnd.n7211 585
R6864 gnd.n506 gnd.n505 585
R6865 gnd.n505 gnd.n504 585
R6866 gnd.n7206 gnd.n7205 585
R6867 gnd.n7205 gnd.n7204 585
R6868 gnd.n509 gnd.n508 585
R6869 gnd.n7203 gnd.n509 585
R6870 gnd.n7201 gnd.n7200 585
R6871 gnd.n7202 gnd.n7201 585
R6872 gnd.n512 gnd.n511 585
R6873 gnd.n511 gnd.n510 585
R6874 gnd.n7196 gnd.n7195 585
R6875 gnd.n7195 gnd.n7194 585
R6876 gnd.n515 gnd.n514 585
R6877 gnd.n7193 gnd.n515 585
R6878 gnd.n7191 gnd.n7190 585
R6879 gnd.n7192 gnd.n7191 585
R6880 gnd.n518 gnd.n517 585
R6881 gnd.n517 gnd.n516 585
R6882 gnd.n7186 gnd.n7185 585
R6883 gnd.n7185 gnd.n7184 585
R6884 gnd.n521 gnd.n520 585
R6885 gnd.n7183 gnd.n521 585
R6886 gnd.n7181 gnd.n7180 585
R6887 gnd.n7182 gnd.n7181 585
R6888 gnd.n524 gnd.n523 585
R6889 gnd.n523 gnd.n522 585
R6890 gnd.n7176 gnd.n7175 585
R6891 gnd.n7175 gnd.n7174 585
R6892 gnd.n527 gnd.n526 585
R6893 gnd.n7173 gnd.n527 585
R6894 gnd.n7171 gnd.n7170 585
R6895 gnd.n7172 gnd.n7171 585
R6896 gnd.n530 gnd.n529 585
R6897 gnd.n529 gnd.n528 585
R6898 gnd.n7166 gnd.n7165 585
R6899 gnd.n7165 gnd.n7164 585
R6900 gnd.n533 gnd.n532 585
R6901 gnd.n7163 gnd.n533 585
R6902 gnd.n7161 gnd.n7160 585
R6903 gnd.n7162 gnd.n7161 585
R6904 gnd.n536 gnd.n535 585
R6905 gnd.n535 gnd.n534 585
R6906 gnd.n7156 gnd.n7155 585
R6907 gnd.n7155 gnd.n7154 585
R6908 gnd.n539 gnd.n538 585
R6909 gnd.n7153 gnd.n539 585
R6910 gnd.n7151 gnd.n7150 585
R6911 gnd.n7152 gnd.n7151 585
R6912 gnd.n542 gnd.n541 585
R6913 gnd.n541 gnd.n540 585
R6914 gnd.n7146 gnd.n7145 585
R6915 gnd.n7145 gnd.n7144 585
R6916 gnd.n545 gnd.n544 585
R6917 gnd.n7143 gnd.n545 585
R6918 gnd.n7141 gnd.n7140 585
R6919 gnd.n7142 gnd.n7141 585
R6920 gnd.n6462 gnd.n6461 585
R6921 gnd.n6463 gnd.n6462 585
R6922 gnd.n1099 gnd.n1098 585
R6923 gnd.n4568 gnd.n1099 585
R6924 gnd.n6471 gnd.n6470 585
R6925 gnd.n6470 gnd.n6469 585
R6926 gnd.n6472 gnd.n1093 585
R6927 gnd.n4528 gnd.n1093 585
R6928 gnd.n6474 gnd.n6473 585
R6929 gnd.n6475 gnd.n6474 585
R6930 gnd.n1078 gnd.n1077 585
R6931 gnd.n4519 gnd.n1078 585
R6932 gnd.n6483 gnd.n6482 585
R6933 gnd.n6482 gnd.n6481 585
R6934 gnd.n6484 gnd.n1072 585
R6935 gnd.n4511 gnd.n1072 585
R6936 gnd.n6486 gnd.n6485 585
R6937 gnd.n6487 gnd.n6486 585
R6938 gnd.n1056 gnd.n1055 585
R6939 gnd.n4446 gnd.n1056 585
R6940 gnd.n6495 gnd.n6494 585
R6941 gnd.n6494 gnd.n6493 585
R6942 gnd.n6496 gnd.n1050 585
R6943 gnd.n4434 gnd.n1050 585
R6944 gnd.n6498 gnd.n6497 585
R6945 gnd.n6499 gnd.n6498 585
R6946 gnd.n1036 gnd.n1035 585
R6947 gnd.n4457 gnd.n1036 585
R6948 gnd.n6507 gnd.n6506 585
R6949 gnd.n6506 gnd.n6505 585
R6950 gnd.n6508 gnd.n1030 585
R6951 gnd.n4426 gnd.n1030 585
R6952 gnd.n6510 gnd.n6509 585
R6953 gnd.n6511 gnd.n6510 585
R6954 gnd.n1014 gnd.n1013 585
R6955 gnd.n4393 gnd.n1014 585
R6956 gnd.n6519 gnd.n6518 585
R6957 gnd.n6518 gnd.n6517 585
R6958 gnd.n6520 gnd.n1008 585
R6959 gnd.n4385 gnd.n1008 585
R6960 gnd.n6522 gnd.n6521 585
R6961 gnd.n6523 gnd.n6522 585
R6962 gnd.n994 gnd.n993 585
R6963 gnd.n4408 gnd.n994 585
R6964 gnd.n6531 gnd.n6530 585
R6965 gnd.n6530 gnd.n6529 585
R6966 gnd.n6532 gnd.n988 585
R6967 gnd.n4377 gnd.n988 585
R6968 gnd.n6534 gnd.n6533 585
R6969 gnd.n6535 gnd.n6534 585
R6970 gnd.n989 gnd.n987 585
R6971 gnd.n4359 gnd.n987 585
R6972 gnd.n4336 gnd.n974 585
R6973 gnd.n6541 gnd.n974 585
R6974 gnd.n4338 gnd.n4337 585
R6975 gnd.n4337 gnd.n970 585
R6976 gnd.n4339 gnd.n2186 585
R6977 gnd.n4350 gnd.n2186 585
R6978 gnd.n4340 gnd.n2195 585
R6979 gnd.n2195 gnd.n2193 585
R6980 gnd.n4342 gnd.n4341 585
R6981 gnd.n4343 gnd.n4342 585
R6982 gnd.n2196 gnd.n2194 585
R6983 gnd.n2211 gnd.n2194 585
R6984 gnd.n2212 gnd.n2198 585
R6985 gnd.n4324 gnd.n2212 585
R6986 gnd.n4313 gnd.n2220 585
R6987 gnd.n2220 gnd.n2209 585
R6988 gnd.n4315 gnd.n4314 585
R6989 gnd.n4316 gnd.n4315 585
R6990 gnd.n2221 gnd.n2219 585
R6991 gnd.n2219 gnd.n2216 585
R6992 gnd.n4309 gnd.n4308 585
R6993 gnd.n4308 gnd.n4307 585
R6994 gnd.n2224 gnd.n2223 585
R6995 gnd.n2225 gnd.n2224 585
R6996 gnd.n4298 gnd.n4297 585
R6997 gnd.n4299 gnd.n4298 585
R6998 gnd.n2235 gnd.n2234 585
R6999 gnd.n2242 gnd.n2234 585
R7000 gnd.n4293 gnd.n4292 585
R7001 gnd.n4292 gnd.n4291 585
R7002 gnd.n2238 gnd.n2237 585
R7003 gnd.n2239 gnd.n2238 585
R7004 gnd.n4281 gnd.n4280 585
R7005 gnd.n4282 gnd.n4281 585
R7006 gnd.n2252 gnd.n2251 585
R7007 gnd.n2251 gnd.n2248 585
R7008 gnd.n4276 gnd.n4275 585
R7009 gnd.n4275 gnd.n4274 585
R7010 gnd.n2255 gnd.n2254 585
R7011 gnd.n2256 gnd.n2255 585
R7012 gnd.n4265 gnd.n4264 585
R7013 gnd.n4266 gnd.n4265 585
R7014 gnd.n2267 gnd.n2266 585
R7015 gnd.n2274 gnd.n2266 585
R7016 gnd.n4260 gnd.n4259 585
R7017 gnd.n4259 gnd.n4258 585
R7018 gnd.n2270 gnd.n2269 585
R7019 gnd.n2271 gnd.n2270 585
R7020 gnd.n4249 gnd.n4248 585
R7021 gnd.n4250 gnd.n4249 585
R7022 gnd.n2284 gnd.n2283 585
R7023 gnd.n2283 gnd.n2280 585
R7024 gnd.n4244 gnd.n4243 585
R7025 gnd.n4243 gnd.n4242 585
R7026 gnd.n2287 gnd.n2286 585
R7027 gnd.n2288 gnd.n2287 585
R7028 gnd.n4233 gnd.n4232 585
R7029 gnd.n4234 gnd.n4233 585
R7030 gnd.n2299 gnd.n2298 585
R7031 gnd.n2306 gnd.n2298 585
R7032 gnd.n4228 gnd.n4227 585
R7033 gnd.n4227 gnd.n4226 585
R7034 gnd.n2302 gnd.n2301 585
R7035 gnd.n2303 gnd.n2302 585
R7036 gnd.n4217 gnd.n4216 585
R7037 gnd.n4218 gnd.n4217 585
R7038 gnd.n2316 gnd.n2315 585
R7039 gnd.n2315 gnd.n2312 585
R7040 gnd.n4212 gnd.n4211 585
R7041 gnd.n4211 gnd.n4210 585
R7042 gnd.n2319 gnd.n2318 585
R7043 gnd.n2320 gnd.n2319 585
R7044 gnd.n4201 gnd.n4200 585
R7045 gnd.n4202 gnd.n4201 585
R7046 gnd.n2331 gnd.n2330 585
R7047 gnd.n3972 gnd.n2330 585
R7048 gnd.n4196 gnd.n4195 585
R7049 gnd.n4195 gnd.n4194 585
R7050 gnd.n3831 gnd.n2333 585
R7051 gnd.n3834 gnd.n3832 585
R7052 gnd.n3837 gnd.n3836 585
R7053 gnd.n3829 gnd.n3828 585
R7054 gnd.n3842 gnd.n3841 585
R7055 gnd.n3844 gnd.n3827 585
R7056 gnd.n3847 gnd.n3846 585
R7057 gnd.n3825 gnd.n3824 585
R7058 gnd.n3852 gnd.n3851 585
R7059 gnd.n3854 gnd.n3823 585
R7060 gnd.n3857 gnd.n3856 585
R7061 gnd.n3821 gnd.n3820 585
R7062 gnd.n3862 gnd.n3861 585
R7063 gnd.n3864 gnd.n3819 585
R7064 gnd.n3867 gnd.n3866 585
R7065 gnd.n3817 gnd.n3816 585
R7066 gnd.n3872 gnd.n3871 585
R7067 gnd.n3874 gnd.n3815 585
R7068 gnd.n3876 gnd.n3875 585
R7069 gnd.n3875 gnd.n3808 585
R7070 gnd.n5559 gnd.n5558 585
R7071 gnd.n2041 gnd.n2033 585
R7072 gnd.n5566 gnd.n2030 585
R7073 gnd.n5567 gnd.n2029 585
R7074 gnd.n2055 gnd.n2023 585
R7075 gnd.n5574 gnd.n2022 585
R7076 gnd.n5575 gnd.n2021 585
R7077 gnd.n2053 gnd.n2013 585
R7078 gnd.n5582 gnd.n2012 585
R7079 gnd.n5583 gnd.n2011 585
R7080 gnd.n2050 gnd.n2005 585
R7081 gnd.n5590 gnd.n2004 585
R7082 gnd.n5591 gnd.n2003 585
R7083 gnd.n2048 gnd.n1996 585
R7084 gnd.n5598 gnd.n1995 585
R7085 gnd.n5599 gnd.n1994 585
R7086 gnd.n2045 gnd.n1993 585
R7087 gnd.n2044 gnd.n2043 585
R7088 gnd.n1115 gnd.n1113 585
R7089 gnd.n5556 gnd.n1113 585
R7090 gnd.n2126 gnd.n1111 585
R7091 gnd.n6463 gnd.n1111 585
R7092 gnd.n4567 gnd.n4566 585
R7093 gnd.n4568 gnd.n4567 585
R7094 gnd.n2125 gnd.n1102 585
R7095 gnd.n6469 gnd.n1102 585
R7096 gnd.n4530 gnd.n4529 585
R7097 gnd.n4529 gnd.n4528 585
R7098 gnd.n2128 gnd.n1091 585
R7099 gnd.n6475 gnd.n1091 585
R7100 gnd.n4518 gnd.n4517 585
R7101 gnd.n4519 gnd.n4518 585
R7102 gnd.n2132 gnd.n1080 585
R7103 gnd.n6481 gnd.n1080 585
R7104 gnd.n4513 gnd.n4512 585
R7105 gnd.n4512 gnd.n4511 585
R7106 gnd.n2134 gnd.n1070 585
R7107 gnd.n6487 gnd.n1070 585
R7108 gnd.n4449 gnd.n4447 585
R7109 gnd.n4447 gnd.n4446 585
R7110 gnd.n4450 gnd.n1059 585
R7111 gnd.n6493 gnd.n1059 585
R7112 gnd.n4451 gnd.n2151 585
R7113 gnd.n4434 gnd.n2151 585
R7114 gnd.n2148 gnd.n1048 585
R7115 gnd.n6499 gnd.n1048 585
R7116 gnd.n4456 gnd.n4455 585
R7117 gnd.n4457 gnd.n4456 585
R7118 gnd.n2147 gnd.n1038 585
R7119 gnd.n6505 gnd.n1038 585
R7120 gnd.n4396 gnd.n2157 585
R7121 gnd.n4426 gnd.n2157 585
R7122 gnd.n4395 gnd.n1028 585
R7123 gnd.n6511 gnd.n1028 585
R7124 gnd.n4400 gnd.n4394 585
R7125 gnd.n4394 gnd.n4393 585
R7126 gnd.n4401 gnd.n1017 585
R7127 gnd.n6517 gnd.n1017 585
R7128 gnd.n4402 gnd.n2172 585
R7129 gnd.n4385 gnd.n2172 585
R7130 gnd.n2169 gnd.n1006 585
R7131 gnd.n6523 gnd.n1006 585
R7132 gnd.n4407 gnd.n4406 585
R7133 gnd.n4408 gnd.n4407 585
R7134 gnd.n2168 gnd.n996 585
R7135 gnd.n6529 gnd.n996 585
R7136 gnd.n4366 gnd.n4365 585
R7137 gnd.n4377 gnd.n4366 585
R7138 gnd.n2178 gnd.n985 585
R7139 gnd.n6535 gnd.n985 585
R7140 gnd.n4361 gnd.n4360 585
R7141 gnd.n4360 gnd.n4359 585
R7142 gnd.n2180 gnd.n972 585
R7143 gnd.n6541 gnd.n972 585
R7144 gnd.n3915 gnd.n3914 585
R7145 gnd.n3914 gnd.n970 585
R7146 gnd.n3918 gnd.n2185 585
R7147 gnd.n4350 gnd.n2185 585
R7148 gnd.n3919 gnd.n3913 585
R7149 gnd.n3913 gnd.n2193 585
R7150 gnd.n3920 gnd.n2191 585
R7151 gnd.n4343 gnd.n2191 585
R7152 gnd.n3911 gnd.n3910 585
R7153 gnd.n3910 gnd.n2211 585
R7154 gnd.n3924 gnd.n2210 585
R7155 gnd.n4324 gnd.n2210 585
R7156 gnd.n3926 gnd.n3925 585
R7157 gnd.n3925 gnd.n2209 585
R7158 gnd.n3927 gnd.n2218 585
R7159 gnd.n4316 gnd.n2218 585
R7160 gnd.n3929 gnd.n3928 585
R7161 gnd.n3928 gnd.n2216 585
R7162 gnd.n3930 gnd.n2227 585
R7163 gnd.n4307 gnd.n2227 585
R7164 gnd.n3932 gnd.n3931 585
R7165 gnd.n3931 gnd.n2225 585
R7166 gnd.n3933 gnd.n2233 585
R7167 gnd.n4299 gnd.n2233 585
R7168 gnd.n3935 gnd.n3934 585
R7169 gnd.n3934 gnd.n2242 585
R7170 gnd.n3936 gnd.n2241 585
R7171 gnd.n4291 gnd.n2241 585
R7172 gnd.n3938 gnd.n3937 585
R7173 gnd.n3937 gnd.n2239 585
R7174 gnd.n3939 gnd.n2250 585
R7175 gnd.n4282 gnd.n2250 585
R7176 gnd.n3941 gnd.n3940 585
R7177 gnd.n3940 gnd.n2248 585
R7178 gnd.n3942 gnd.n2258 585
R7179 gnd.n4274 gnd.n2258 585
R7180 gnd.n3944 gnd.n3943 585
R7181 gnd.n3943 gnd.n2256 585
R7182 gnd.n3945 gnd.n2265 585
R7183 gnd.n4266 gnd.n2265 585
R7184 gnd.n3947 gnd.n3946 585
R7185 gnd.n3946 gnd.n2274 585
R7186 gnd.n3948 gnd.n2273 585
R7187 gnd.n4258 gnd.n2273 585
R7188 gnd.n3950 gnd.n3949 585
R7189 gnd.n3949 gnd.n2271 585
R7190 gnd.n3951 gnd.n2282 585
R7191 gnd.n4250 gnd.n2282 585
R7192 gnd.n3953 gnd.n3952 585
R7193 gnd.n3952 gnd.n2280 585
R7194 gnd.n3954 gnd.n2290 585
R7195 gnd.n4242 gnd.n2290 585
R7196 gnd.n3956 gnd.n3955 585
R7197 gnd.n3955 gnd.n2288 585
R7198 gnd.n3957 gnd.n2297 585
R7199 gnd.n4234 gnd.n2297 585
R7200 gnd.n3959 gnd.n3958 585
R7201 gnd.n3958 gnd.n2306 585
R7202 gnd.n3960 gnd.n2305 585
R7203 gnd.n4226 gnd.n2305 585
R7204 gnd.n3962 gnd.n3961 585
R7205 gnd.n3961 gnd.n2303 585
R7206 gnd.n3963 gnd.n2314 585
R7207 gnd.n4218 gnd.n2314 585
R7208 gnd.n3965 gnd.n3964 585
R7209 gnd.n3964 gnd.n2312 585
R7210 gnd.n3966 gnd.n2322 585
R7211 gnd.n4210 gnd.n2322 585
R7212 gnd.n3968 gnd.n3967 585
R7213 gnd.n3967 gnd.n2320 585
R7214 gnd.n3969 gnd.n2329 585
R7215 gnd.n4202 gnd.n2329 585
R7216 gnd.n3971 gnd.n3970 585
R7217 gnd.n3972 gnd.n3971 585
R7218 gnd.n3811 gnd.n3810 585
R7219 gnd.n4194 gnd.n3810 585
R7220 gnd.n7708 gnd.n129 585
R7221 gnd.n7804 gnd.n129 585
R7222 gnd.n7709 gnd.n7646 585
R7223 gnd.n7646 gnd.n126 585
R7224 gnd.n7710 gnd.n207 585
R7225 gnd.n7724 gnd.n207 585
R7226 gnd.n219 gnd.n217 585
R7227 gnd.n217 gnd.n206 585
R7228 gnd.n7715 gnd.n7714 585
R7229 gnd.n7716 gnd.n7715 585
R7230 gnd.n218 gnd.n216 585
R7231 gnd.n216 gnd.n213 585
R7232 gnd.n7642 gnd.n7641 585
R7233 gnd.n7641 gnd.n7640 585
R7234 gnd.n222 gnd.n221 585
R7235 gnd.n232 gnd.n222 585
R7236 gnd.n7631 gnd.n7630 585
R7237 gnd.n7632 gnd.n7631 585
R7238 gnd.n234 gnd.n233 585
R7239 gnd.n233 gnd.n229 585
R7240 gnd.n7626 gnd.n7625 585
R7241 gnd.n7625 gnd.n7624 585
R7242 gnd.n237 gnd.n236 585
R7243 gnd.n247 gnd.n237 585
R7244 gnd.n7615 gnd.n7614 585
R7245 gnd.n7616 gnd.n7615 585
R7246 gnd.n249 gnd.n248 585
R7247 gnd.n254 gnd.n248 585
R7248 gnd.n7610 gnd.n7609 585
R7249 gnd.n7609 gnd.n7608 585
R7250 gnd.n252 gnd.n251 585
R7251 gnd.n263 gnd.n252 585
R7252 gnd.n7599 gnd.n7598 585
R7253 gnd.n7600 gnd.n7599 585
R7254 gnd.n265 gnd.n264 585
R7255 gnd.n264 gnd.n260 585
R7256 gnd.n7594 gnd.n7593 585
R7257 gnd.n7593 gnd.n7592 585
R7258 gnd.n268 gnd.n267 585
R7259 gnd.n269 gnd.n268 585
R7260 gnd.n7583 gnd.n7582 585
R7261 gnd.n7584 gnd.n7583 585
R7262 gnd.n279 gnd.n278 585
R7263 gnd.n284 gnd.n278 585
R7264 gnd.n7578 gnd.n7577 585
R7265 gnd.n7577 gnd.n7576 585
R7266 gnd.n282 gnd.n281 585
R7267 gnd.n293 gnd.n282 585
R7268 gnd.n7567 gnd.n7566 585
R7269 gnd.n7568 gnd.n7567 585
R7270 gnd.n295 gnd.n294 585
R7271 gnd.n294 gnd.n290 585
R7272 gnd.n7562 gnd.n7561 585
R7273 gnd.n7561 gnd.n7560 585
R7274 gnd.n298 gnd.n297 585
R7275 gnd.n299 gnd.n298 585
R7276 gnd.n7538 gnd.n7537 585
R7277 gnd.n7537 gnd.n7536 585
R7278 gnd.n7539 gnd.n327 585
R7279 gnd.n7532 gnd.n327 585
R7280 gnd.n333 gnd.n325 585
R7281 gnd.n334 gnd.n333 585
R7282 gnd.n7543 gnd.n324 585
R7283 gnd.n7459 gnd.n324 585
R7284 gnd.n7544 gnd.n323 585
R7285 gnd.n340 gnd.n323 585
R7286 gnd.n7545 gnd.n322 585
R7287 gnd.n7453 gnd.n322 585
R7288 gnd.n319 gnd.n317 585
R7289 gnd.n317 gnd.n315 585
R7290 gnd.n7550 gnd.n7549 585
R7291 gnd.n7551 gnd.n7550 585
R7292 gnd.n318 gnd.n316 585
R7293 gnd.n7444 gnd.n316 585
R7294 gnd.n7412 gnd.n7410 585
R7295 gnd.n7410 gnd.n350 585
R7296 gnd.n7413 gnd.n359 585
R7297 gnd.n7429 gnd.n359 585
R7298 gnd.n7414 gnd.n7409 585
R7299 gnd.n7409 gnd.n7408 585
R7300 gnd.n374 gnd.n372 585
R7301 gnd.n7392 gnd.n372 585
R7302 gnd.n7419 gnd.n7418 585
R7303 gnd.n7420 gnd.n7419 585
R7304 gnd.n373 gnd.n371 585
R7305 gnd.n7398 gnd.n371 585
R7306 gnd.n7367 gnd.n7366 585
R7307 gnd.n7366 gnd.n7365 585
R7308 gnd.n7368 gnd.n392 585
R7309 gnd.n7384 gnd.n392 585
R7310 gnd.n406 gnd.n404 585
R7311 gnd.n6143 gnd.n404 585
R7312 gnd.n7373 gnd.n7372 585
R7313 gnd.n7374 gnd.n7373 585
R7314 gnd.n405 gnd.n403 585
R7315 gnd.n6138 gnd.n403 585
R7316 gnd.n6192 gnd.n6190 585
R7317 gnd.n6190 gnd.n6189 585
R7318 gnd.n6193 gnd.n1360 585
R7319 gnd.n1373 gnd.n1360 585
R7320 gnd.n6194 gnd.n1359 585
R7321 gnd.n6181 gnd.n1359 585
R7322 gnd.n6158 gnd.n1357 585
R7323 gnd.n6159 gnd.n6158 585
R7324 gnd.n6198 gnd.n1356 585
R7325 gnd.n1398 gnd.n1356 585
R7326 gnd.n6199 gnd.n1355 585
R7327 gnd.n6121 gnd.n1355 585
R7328 gnd.n6200 gnd.n1354 585
R7329 gnd.n1407 gnd.n1354 585
R7330 gnd.n6110 gnd.n1352 585
R7331 gnd.n6111 gnd.n6110 585
R7332 gnd.n6204 gnd.n1351 585
R7333 gnd.n6098 gnd.n1351 585
R7334 gnd.n6205 gnd.n1350 585
R7335 gnd.n1414 gnd.n1350 585
R7336 gnd.n6206 gnd.n1349 585
R7337 gnd.n6084 gnd.n1349 585
R7338 gnd.n1434 gnd.n1347 585
R7339 gnd.n1435 gnd.n1434 585
R7340 gnd.n6210 gnd.n1346 585
R7341 gnd.n6074 gnd.n1346 585
R7342 gnd.n6211 gnd.n1345 585
R7343 gnd.n6062 gnd.n1345 585
R7344 gnd.n6212 gnd.n1344 585
R7345 gnd.n1452 gnd.n1344 585
R7346 gnd.n1341 gnd.n1340 585
R7347 gnd.n6053 gnd.n1340 585
R7348 gnd.n6217 gnd.n6216 585
R7349 gnd.n6218 gnd.n6217 585
R7350 gnd.n1517 gnd.n1339 585
R7351 gnd.n1522 gnd.n1521 585
R7352 gnd.n1524 gnd.n1523 585
R7353 gnd.n1527 gnd.n1526 585
R7354 gnd.n1525 gnd.n1510 585
R7355 gnd.n1541 gnd.n1540 585
R7356 gnd.n1543 gnd.n1542 585
R7357 gnd.n1546 gnd.n1545 585
R7358 gnd.n1544 gnd.n1503 585
R7359 gnd.n1560 gnd.n1559 585
R7360 gnd.n1562 gnd.n1561 585
R7361 gnd.n1565 gnd.n1564 585
R7362 gnd.n1563 gnd.n1496 585
R7363 gnd.n1578 gnd.n1577 585
R7364 gnd.n1580 gnd.n1579 585
R7365 gnd.n1489 gnd.n1488 585
R7366 gnd.n1593 gnd.n1490 585
R7367 gnd.n1594 gnd.n1485 585
R7368 gnd.n1595 gnd.n1284 585
R7369 gnd.n6294 gnd.n1284 585
R7370 gnd.n7807 gnd.n7806 585
R7371 gnd.n7679 gnd.n124 585
R7372 gnd.n7681 gnd.n7680 585
R7373 gnd.n7677 gnd.n7676 585
R7374 gnd.n7685 gnd.n7675 585
R7375 gnd.n7686 gnd.n7673 585
R7376 gnd.n7687 gnd.n7672 585
R7377 gnd.n7670 gnd.n7668 585
R7378 gnd.n7691 gnd.n7667 585
R7379 gnd.n7692 gnd.n7665 585
R7380 gnd.n7693 gnd.n7664 585
R7381 gnd.n7662 gnd.n7660 585
R7382 gnd.n7697 gnd.n7659 585
R7383 gnd.n7698 gnd.n7657 585
R7384 gnd.n7699 gnd.n7656 585
R7385 gnd.n7654 gnd.n7652 585
R7386 gnd.n7703 gnd.n7651 585
R7387 gnd.n7704 gnd.n7649 585
R7388 gnd.n7705 gnd.n7648 585
R7389 gnd.n7648 gnd.n128 585
R7390 gnd.n7805 gnd.n120 585
R7391 gnd.n7805 gnd.n7804 585
R7392 gnd.n7811 gnd.n119 585
R7393 gnd.n126 gnd.n119 585
R7394 gnd.n7812 gnd.n118 585
R7395 gnd.n7724 gnd.n118 585
R7396 gnd.n7813 gnd.n117 585
R7397 gnd.n206 gnd.n117 585
R7398 gnd.n215 gnd.n115 585
R7399 gnd.n7716 gnd.n215 585
R7400 gnd.n7817 gnd.n114 585
R7401 gnd.n213 gnd.n114 585
R7402 gnd.n7818 gnd.n113 585
R7403 gnd.n7640 gnd.n113 585
R7404 gnd.n7819 gnd.n112 585
R7405 gnd.n232 gnd.n112 585
R7406 gnd.n231 gnd.n110 585
R7407 gnd.n7632 gnd.n231 585
R7408 gnd.n7823 gnd.n109 585
R7409 gnd.n229 gnd.n109 585
R7410 gnd.n7824 gnd.n108 585
R7411 gnd.n7624 gnd.n108 585
R7412 gnd.n7825 gnd.n107 585
R7413 gnd.n247 gnd.n107 585
R7414 gnd.n246 gnd.n105 585
R7415 gnd.n7616 gnd.n246 585
R7416 gnd.n7829 gnd.n104 585
R7417 gnd.n254 gnd.n104 585
R7418 gnd.n7830 gnd.n103 585
R7419 gnd.n7608 gnd.n103 585
R7420 gnd.n7831 gnd.n102 585
R7421 gnd.n263 gnd.n102 585
R7422 gnd.n262 gnd.n100 585
R7423 gnd.n7600 gnd.n262 585
R7424 gnd.n7835 gnd.n99 585
R7425 gnd.n260 gnd.n99 585
R7426 gnd.n7836 gnd.n98 585
R7427 gnd.n7592 gnd.n98 585
R7428 gnd.n7837 gnd.n97 585
R7429 gnd.n269 gnd.n97 585
R7430 gnd.n277 gnd.n95 585
R7431 gnd.n7584 gnd.n277 585
R7432 gnd.n7841 gnd.n94 585
R7433 gnd.n284 gnd.n94 585
R7434 gnd.n7842 gnd.n93 585
R7435 gnd.n7576 gnd.n93 585
R7436 gnd.n7843 gnd.n92 585
R7437 gnd.n293 gnd.n92 585
R7438 gnd.n292 gnd.n90 585
R7439 gnd.n7568 gnd.n292 585
R7440 gnd.n7847 gnd.n89 585
R7441 gnd.n290 gnd.n89 585
R7442 gnd.n7848 gnd.n88 585
R7443 gnd.n7560 gnd.n88 585
R7444 gnd.n7849 gnd.n87 585
R7445 gnd.n299 gnd.n87 585
R7446 gnd.n329 gnd.n85 585
R7447 gnd.n7536 gnd.n329 585
R7448 gnd.n7853 gnd.n84 585
R7449 gnd.n7532 gnd.n84 585
R7450 gnd.n7854 gnd.n83 585
R7451 gnd.n334 gnd.n83 585
R7452 gnd.n7855 gnd.n82 585
R7453 gnd.n7459 gnd.n82 585
R7454 gnd.n345 gnd.n80 585
R7455 gnd.n345 gnd.n340 585
R7456 gnd.n7452 gnd.n7451 585
R7457 gnd.n7453 gnd.n7452 585
R7458 gnd.n7450 gnd.n344 585
R7459 gnd.n344 gnd.n315 585
R7460 gnd.n346 gnd.n314 585
R7461 gnd.n7551 gnd.n314 585
R7462 gnd.n7446 gnd.n7445 585
R7463 gnd.n7445 gnd.n7444 585
R7464 gnd.n349 gnd.n348 585
R7465 gnd.n350 gnd.n349 585
R7466 gnd.n380 gnd.n357 585
R7467 gnd.n7429 gnd.n357 585
R7468 gnd.n7407 gnd.n7406 585
R7469 gnd.n7408 gnd.n7407 585
R7470 gnd.n379 gnd.n378 585
R7471 gnd.n7392 gnd.n378 585
R7472 gnd.n7401 gnd.n369 585
R7473 gnd.n7420 gnd.n369 585
R7474 gnd.n7400 gnd.n7399 585
R7475 gnd.n7399 gnd.n7398 585
R7476 gnd.n383 gnd.n382 585
R7477 gnd.n7365 gnd.n383 585
R7478 gnd.n6145 gnd.n391 585
R7479 gnd.n7384 gnd.n391 585
R7480 gnd.n6146 gnd.n6144 585
R7481 gnd.n6144 gnd.n6143 585
R7482 gnd.n6140 gnd.n401 585
R7483 gnd.n7374 gnd.n401 585
R7484 gnd.n6150 gnd.n6139 585
R7485 gnd.n6139 gnd.n6138 585
R7486 gnd.n6151 gnd.n1363 585
R7487 gnd.n6189 gnd.n1363 585
R7488 gnd.n6152 gnd.n1386 585
R7489 gnd.n1386 gnd.n1373 585
R7490 gnd.n1383 gnd.n1372 585
R7491 gnd.n6181 gnd.n1372 585
R7492 gnd.n6157 gnd.n6156 585
R7493 gnd.n6159 gnd.n6157 585
R7494 gnd.n1382 gnd.n1381 585
R7495 gnd.n1398 gnd.n1381 585
R7496 gnd.n6091 gnd.n1395 585
R7497 gnd.n6121 gnd.n1395 585
R7498 gnd.n6092 gnd.n6090 585
R7499 gnd.n6090 gnd.n1407 585
R7500 gnd.n1418 gnd.n1406 585
R7501 gnd.n6111 gnd.n1406 585
R7502 gnd.n6097 gnd.n6096 585
R7503 gnd.n6098 gnd.n6097 585
R7504 gnd.n1417 gnd.n1416 585
R7505 gnd.n1416 gnd.n1414 585
R7506 gnd.n6086 gnd.n6085 585
R7507 gnd.n6085 gnd.n6084 585
R7508 gnd.n1421 gnd.n1420 585
R7509 gnd.n1435 gnd.n1421 585
R7510 gnd.n1477 gnd.n1433 585
R7511 gnd.n6074 gnd.n1433 585
R7512 gnd.n6061 gnd.n6060 585
R7513 gnd.n6062 gnd.n6061 585
R7514 gnd.n1476 gnd.n1475 585
R7515 gnd.n1475 gnd.n1452 585
R7516 gnd.n6055 gnd.n6054 585
R7517 gnd.n6054 gnd.n6053 585
R7518 gnd.n6043 gnd.n1337 585
R7519 gnd.n6218 gnd.n1337 585
R7520 gnd.n3715 gnd.n3714 585
R7521 gnd.n3716 gnd.n3715 585
R7522 gnd.n2410 gnd.n2409 585
R7523 gnd.n2416 gnd.n2409 585
R7524 gnd.n3690 gnd.n2428 585
R7525 gnd.n2428 gnd.n2415 585
R7526 gnd.n3692 gnd.n3691 585
R7527 gnd.n3693 gnd.n3692 585
R7528 gnd.n2429 gnd.n2427 585
R7529 gnd.n2427 gnd.n2423 585
R7530 gnd.n3424 gnd.n3423 585
R7531 gnd.n3423 gnd.n3422 585
R7532 gnd.n2434 gnd.n2433 585
R7533 gnd.n3393 gnd.n2434 585
R7534 gnd.n3413 gnd.n3412 585
R7535 gnd.n3412 gnd.n3411 585
R7536 gnd.n2441 gnd.n2440 585
R7537 gnd.n3399 gnd.n2441 585
R7538 gnd.n3369 gnd.n2461 585
R7539 gnd.n2461 gnd.n2460 585
R7540 gnd.n3371 gnd.n3370 585
R7541 gnd.n3372 gnd.n3371 585
R7542 gnd.n2462 gnd.n2459 585
R7543 gnd.n2470 gnd.n2459 585
R7544 gnd.n3347 gnd.n2482 585
R7545 gnd.n2482 gnd.n2469 585
R7546 gnd.n3349 gnd.n3348 585
R7547 gnd.n3350 gnd.n3349 585
R7548 gnd.n2483 gnd.n2481 585
R7549 gnd.n2481 gnd.n2477 585
R7550 gnd.n3335 gnd.n3334 585
R7551 gnd.n3334 gnd.n3333 585
R7552 gnd.n2488 gnd.n2487 585
R7553 gnd.n2498 gnd.n2488 585
R7554 gnd.n3324 gnd.n3323 585
R7555 gnd.n3323 gnd.n3322 585
R7556 gnd.n2495 gnd.n2494 585
R7557 gnd.n3310 gnd.n2495 585
R7558 gnd.n3284 gnd.n2516 585
R7559 gnd.n2516 gnd.n2505 585
R7560 gnd.n3286 gnd.n3285 585
R7561 gnd.n3287 gnd.n3286 585
R7562 gnd.n2517 gnd.n2515 585
R7563 gnd.n2525 gnd.n2515 585
R7564 gnd.n3262 gnd.n2537 585
R7565 gnd.n2537 gnd.n2524 585
R7566 gnd.n3264 gnd.n3263 585
R7567 gnd.n3265 gnd.n3264 585
R7568 gnd.n2538 gnd.n2536 585
R7569 gnd.n2536 gnd.n2532 585
R7570 gnd.n3250 gnd.n3249 585
R7571 gnd.n3249 gnd.n3248 585
R7572 gnd.n2543 gnd.n2542 585
R7573 gnd.n2552 gnd.n2543 585
R7574 gnd.n3239 gnd.n3238 585
R7575 gnd.n3238 gnd.n3237 585
R7576 gnd.n2550 gnd.n2549 585
R7577 gnd.n3225 gnd.n2550 585
R7578 gnd.n2663 gnd.n2662 585
R7579 gnd.n2663 gnd.n2559 585
R7580 gnd.n3182 gnd.n3181 585
R7581 gnd.n3181 gnd.n3180 585
R7582 gnd.n3183 gnd.n2657 585
R7583 gnd.n2668 gnd.n2657 585
R7584 gnd.n3185 gnd.n3184 585
R7585 gnd.n3186 gnd.n3185 585
R7586 gnd.n2658 gnd.n2656 585
R7587 gnd.n2681 gnd.n2656 585
R7588 gnd.n2641 gnd.n2640 585
R7589 gnd.n2644 gnd.n2641 585
R7590 gnd.n3196 gnd.n3195 585
R7591 gnd.n3195 gnd.n3194 585
R7592 gnd.n3197 gnd.n2635 585
R7593 gnd.n3156 gnd.n2635 585
R7594 gnd.n3199 gnd.n3198 585
R7595 gnd.n3200 gnd.n3199 585
R7596 gnd.n2636 gnd.n2634 585
R7597 gnd.n2695 gnd.n2634 585
R7598 gnd.n3148 gnd.n3147 585
R7599 gnd.n3147 gnd.n3146 585
R7600 gnd.n2692 gnd.n2691 585
R7601 gnd.n3130 gnd.n2692 585
R7602 gnd.n3117 gnd.n2711 585
R7603 gnd.n2711 gnd.n2710 585
R7604 gnd.n3119 gnd.n3118 585
R7605 gnd.n3120 gnd.n3119 585
R7606 gnd.n2712 gnd.n2709 585
R7607 gnd.n2718 gnd.n2709 585
R7608 gnd.n3098 gnd.n3097 585
R7609 gnd.n3099 gnd.n3098 585
R7610 gnd.n2729 gnd.n2728 585
R7611 gnd.n2728 gnd.n2724 585
R7612 gnd.n3088 gnd.n3087 585
R7613 gnd.n3089 gnd.n3088 585
R7614 gnd.n2739 gnd.n2738 585
R7615 gnd.n2744 gnd.n2738 585
R7616 gnd.n3066 gnd.n2757 585
R7617 gnd.n2757 gnd.n2743 585
R7618 gnd.n3068 gnd.n3067 585
R7619 gnd.n3069 gnd.n3068 585
R7620 gnd.n2758 gnd.n2756 585
R7621 gnd.n2756 gnd.n2752 585
R7622 gnd.n3057 gnd.n3056 585
R7623 gnd.n3058 gnd.n3057 585
R7624 gnd.n2765 gnd.n2764 585
R7625 gnd.n2769 gnd.n2764 585
R7626 gnd.n3034 gnd.n2786 585
R7627 gnd.n2786 gnd.n2768 585
R7628 gnd.n3036 gnd.n3035 585
R7629 gnd.n3037 gnd.n3036 585
R7630 gnd.n2787 gnd.n2785 585
R7631 gnd.n2785 gnd.n2776 585
R7632 gnd.n3029 gnd.n3028 585
R7633 gnd.n3028 gnd.n3027 585
R7634 gnd.n2834 gnd.n2833 585
R7635 gnd.n2835 gnd.n2834 585
R7636 gnd.n2988 gnd.n2987 585
R7637 gnd.n2989 gnd.n2988 585
R7638 gnd.n2844 gnd.n2843 585
R7639 gnd.n2843 gnd.n2842 585
R7640 gnd.n2983 gnd.n2982 585
R7641 gnd.n2982 gnd.n2981 585
R7642 gnd.n2847 gnd.n2846 585
R7643 gnd.n2848 gnd.n2847 585
R7644 gnd.n2972 gnd.n2971 585
R7645 gnd.n2973 gnd.n2972 585
R7646 gnd.n2855 gnd.n2854 585
R7647 gnd.n2964 gnd.n2854 585
R7648 gnd.n2967 gnd.n2966 585
R7649 gnd.n2966 gnd.n2965 585
R7650 gnd.n2858 gnd.n2857 585
R7651 gnd.n2859 gnd.n2858 585
R7652 gnd.n2953 gnd.n2952 585
R7653 gnd.n2951 gnd.n2877 585
R7654 gnd.n2950 gnd.n2876 585
R7655 gnd.n2955 gnd.n2876 585
R7656 gnd.n2949 gnd.n2948 585
R7657 gnd.n2947 gnd.n2946 585
R7658 gnd.n2945 gnd.n2944 585
R7659 gnd.n2943 gnd.n2942 585
R7660 gnd.n2941 gnd.n2940 585
R7661 gnd.n2939 gnd.n2938 585
R7662 gnd.n2937 gnd.n2936 585
R7663 gnd.n2935 gnd.n2934 585
R7664 gnd.n2933 gnd.n2932 585
R7665 gnd.n2931 gnd.n2930 585
R7666 gnd.n2929 gnd.n2928 585
R7667 gnd.n2927 gnd.n2926 585
R7668 gnd.n2925 gnd.n2924 585
R7669 gnd.n2923 gnd.n2922 585
R7670 gnd.n2921 gnd.n2920 585
R7671 gnd.n2919 gnd.n2918 585
R7672 gnd.n2917 gnd.n2916 585
R7673 gnd.n2915 gnd.n2914 585
R7674 gnd.n2913 gnd.n2912 585
R7675 gnd.n2911 gnd.n2910 585
R7676 gnd.n2909 gnd.n2908 585
R7677 gnd.n2907 gnd.n2906 585
R7678 gnd.n2864 gnd.n2863 585
R7679 gnd.n2958 gnd.n2957 585
R7680 gnd.n3719 gnd.n3718 585
R7681 gnd.n3721 gnd.n3720 585
R7682 gnd.n3723 gnd.n3722 585
R7683 gnd.n3725 gnd.n3724 585
R7684 gnd.n3727 gnd.n3726 585
R7685 gnd.n3729 gnd.n3728 585
R7686 gnd.n3731 gnd.n3730 585
R7687 gnd.n3733 gnd.n3732 585
R7688 gnd.n3735 gnd.n3734 585
R7689 gnd.n3737 gnd.n3736 585
R7690 gnd.n3739 gnd.n3738 585
R7691 gnd.n3741 gnd.n3740 585
R7692 gnd.n3743 gnd.n3742 585
R7693 gnd.n3745 gnd.n3744 585
R7694 gnd.n3747 gnd.n3746 585
R7695 gnd.n3749 gnd.n3748 585
R7696 gnd.n3751 gnd.n3750 585
R7697 gnd.n3753 gnd.n3752 585
R7698 gnd.n3755 gnd.n3754 585
R7699 gnd.n3757 gnd.n3756 585
R7700 gnd.n3759 gnd.n3758 585
R7701 gnd.n3761 gnd.n3760 585
R7702 gnd.n3763 gnd.n3762 585
R7703 gnd.n3765 gnd.n3764 585
R7704 gnd.n3767 gnd.n3766 585
R7705 gnd.n3768 gnd.n2376 585
R7706 gnd.n3769 gnd.n2334 585
R7707 gnd.n3807 gnd.n2334 585
R7708 gnd.n3717 gnd.n2406 585
R7709 gnd.n3717 gnd.n3716 585
R7710 gnd.n3386 gnd.n2405 585
R7711 gnd.n2416 gnd.n2405 585
R7712 gnd.n3388 gnd.n3387 585
R7713 gnd.n3387 gnd.n2415 585
R7714 gnd.n3389 gnd.n2425 585
R7715 gnd.n3693 gnd.n2425 585
R7716 gnd.n3391 gnd.n3390 585
R7717 gnd.n3390 gnd.n2423 585
R7718 gnd.n3392 gnd.n2436 585
R7719 gnd.n3422 gnd.n2436 585
R7720 gnd.n3395 gnd.n3394 585
R7721 gnd.n3394 gnd.n3393 585
R7722 gnd.n3396 gnd.n2443 585
R7723 gnd.n3411 gnd.n2443 585
R7724 gnd.n3398 gnd.n3397 585
R7725 gnd.n3399 gnd.n3398 585
R7726 gnd.n2453 gnd.n2452 585
R7727 gnd.n2460 gnd.n2452 585
R7728 gnd.n3374 gnd.n3373 585
R7729 gnd.n3373 gnd.n3372 585
R7730 gnd.n2456 gnd.n2455 585
R7731 gnd.n2470 gnd.n2456 585
R7732 gnd.n3300 gnd.n3299 585
R7733 gnd.n3299 gnd.n2469 585
R7734 gnd.n3301 gnd.n2479 585
R7735 gnd.n3350 gnd.n2479 585
R7736 gnd.n3303 gnd.n3302 585
R7737 gnd.n3302 gnd.n2477 585
R7738 gnd.n3304 gnd.n2490 585
R7739 gnd.n3333 gnd.n2490 585
R7740 gnd.n3306 gnd.n3305 585
R7741 gnd.n3305 gnd.n2498 585
R7742 gnd.n3307 gnd.n2497 585
R7743 gnd.n3322 gnd.n2497 585
R7744 gnd.n3309 gnd.n3308 585
R7745 gnd.n3310 gnd.n3309 585
R7746 gnd.n2509 gnd.n2508 585
R7747 gnd.n2508 gnd.n2505 585
R7748 gnd.n3289 gnd.n3288 585
R7749 gnd.n3288 gnd.n3287 585
R7750 gnd.n2512 gnd.n2511 585
R7751 gnd.n2525 gnd.n2512 585
R7752 gnd.n3213 gnd.n3212 585
R7753 gnd.n3212 gnd.n2524 585
R7754 gnd.n3214 gnd.n2534 585
R7755 gnd.n3265 gnd.n2534 585
R7756 gnd.n3216 gnd.n3215 585
R7757 gnd.n3215 gnd.n2532 585
R7758 gnd.n3217 gnd.n2545 585
R7759 gnd.n3248 gnd.n2545 585
R7760 gnd.n3219 gnd.n3218 585
R7761 gnd.n3218 gnd.n2552 585
R7762 gnd.n3220 gnd.n2551 585
R7763 gnd.n3237 gnd.n2551 585
R7764 gnd.n3222 gnd.n3221 585
R7765 gnd.n3225 gnd.n3222 585
R7766 gnd.n2562 gnd.n2561 585
R7767 gnd.n2561 gnd.n2559 585
R7768 gnd.n2665 gnd.n2664 585
R7769 gnd.n3180 gnd.n2664 585
R7770 gnd.n2667 gnd.n2666 585
R7771 gnd.n2668 gnd.n2667 585
R7772 gnd.n2678 gnd.n2654 585
R7773 gnd.n3186 gnd.n2654 585
R7774 gnd.n2680 gnd.n2679 585
R7775 gnd.n2681 gnd.n2680 585
R7776 gnd.n2677 gnd.n2676 585
R7777 gnd.n2677 gnd.n2644 585
R7778 gnd.n2675 gnd.n2642 585
R7779 gnd.n3194 gnd.n2642 585
R7780 gnd.n2631 gnd.n2629 585
R7781 gnd.n3156 gnd.n2631 585
R7782 gnd.n3202 gnd.n3201 585
R7783 gnd.n3201 gnd.n3200 585
R7784 gnd.n2630 gnd.n2628 585
R7785 gnd.n2695 gnd.n2630 585
R7786 gnd.n3127 gnd.n2694 585
R7787 gnd.n3146 gnd.n2694 585
R7788 gnd.n3129 gnd.n3128 585
R7789 gnd.n3130 gnd.n3129 585
R7790 gnd.n2704 gnd.n2703 585
R7791 gnd.n2710 gnd.n2703 585
R7792 gnd.n3122 gnd.n3121 585
R7793 gnd.n3121 gnd.n3120 585
R7794 gnd.n2707 gnd.n2706 585
R7795 gnd.n2718 gnd.n2707 585
R7796 gnd.n3007 gnd.n2726 585
R7797 gnd.n3099 gnd.n2726 585
R7798 gnd.n3009 gnd.n3008 585
R7799 gnd.n3008 gnd.n2724 585
R7800 gnd.n3010 gnd.n2737 585
R7801 gnd.n3089 gnd.n2737 585
R7802 gnd.n3012 gnd.n3011 585
R7803 gnd.n3012 gnd.n2744 585
R7804 gnd.n3014 gnd.n3013 585
R7805 gnd.n3013 gnd.n2743 585
R7806 gnd.n3015 gnd.n2754 585
R7807 gnd.n3069 gnd.n2754 585
R7808 gnd.n3017 gnd.n3016 585
R7809 gnd.n3016 gnd.n2752 585
R7810 gnd.n3018 gnd.n2763 585
R7811 gnd.n3058 gnd.n2763 585
R7812 gnd.n3020 gnd.n3019 585
R7813 gnd.n3020 gnd.n2769 585
R7814 gnd.n3022 gnd.n3021 585
R7815 gnd.n3021 gnd.n2768 585
R7816 gnd.n3023 gnd.n2784 585
R7817 gnd.n3037 gnd.n2784 585
R7818 gnd.n3024 gnd.n2837 585
R7819 gnd.n2837 gnd.n2776 585
R7820 gnd.n3026 gnd.n3025 585
R7821 gnd.n3027 gnd.n3026 585
R7822 gnd.n2838 gnd.n2836 585
R7823 gnd.n2836 gnd.n2835 585
R7824 gnd.n2991 gnd.n2990 585
R7825 gnd.n2990 gnd.n2989 585
R7826 gnd.n2841 gnd.n2840 585
R7827 gnd.n2842 gnd.n2841 585
R7828 gnd.n2980 gnd.n2979 585
R7829 gnd.n2981 gnd.n2980 585
R7830 gnd.n2850 gnd.n2849 585
R7831 gnd.n2849 gnd.n2848 585
R7832 gnd.n2975 gnd.n2974 585
R7833 gnd.n2974 gnd.n2973 585
R7834 gnd.n2853 gnd.n2852 585
R7835 gnd.n2964 gnd.n2853 585
R7836 gnd.n2963 gnd.n2962 585
R7837 gnd.n2965 gnd.n2963 585
R7838 gnd.n2861 gnd.n2860 585
R7839 gnd.n2860 gnd.n2859 585
R7840 gnd.n3702 gnd.n2356 585
R7841 gnd.n2408 gnd.n2356 585
R7842 gnd.n3703 gnd.n2418 585
R7843 gnd.n2418 gnd.n2407 585
R7844 gnd.n3705 gnd.n3704 585
R7845 gnd.n3706 gnd.n3705 585
R7846 gnd.n2419 gnd.n2417 585
R7847 gnd.n2426 gnd.n2417 585
R7848 gnd.n3696 gnd.n3695 585
R7849 gnd.n3695 gnd.n3694 585
R7850 gnd.n2422 gnd.n2421 585
R7851 gnd.n3421 gnd.n2422 585
R7852 gnd.n3407 gnd.n2445 585
R7853 gnd.n2445 gnd.n2435 585
R7854 gnd.n3409 gnd.n3408 585
R7855 gnd.n3410 gnd.n3409 585
R7856 gnd.n2446 gnd.n2444 585
R7857 gnd.n2444 gnd.n2442 585
R7858 gnd.n3402 gnd.n3401 585
R7859 gnd.n3401 gnd.n3400 585
R7860 gnd.n2449 gnd.n2448 585
R7861 gnd.n2458 gnd.n2449 585
R7862 gnd.n3358 gnd.n2472 585
R7863 gnd.n2472 gnd.n2457 585
R7864 gnd.n3360 gnd.n3359 585
R7865 gnd.n3361 gnd.n3360 585
R7866 gnd.n2473 gnd.n2471 585
R7867 gnd.n2480 gnd.n2471 585
R7868 gnd.n3353 gnd.n3352 585
R7869 gnd.n3352 gnd.n3351 585
R7870 gnd.n2476 gnd.n2475 585
R7871 gnd.n3332 gnd.n2476 585
R7872 gnd.n3318 gnd.n2500 585
R7873 gnd.n2500 gnd.n2489 585
R7874 gnd.n3320 gnd.n3319 585
R7875 gnd.n3321 gnd.n3320 585
R7876 gnd.n2501 gnd.n2499 585
R7877 gnd.n2499 gnd.n2496 585
R7878 gnd.n3313 gnd.n3312 585
R7879 gnd.n3312 gnd.n3311 585
R7880 gnd.n2504 gnd.n2503 585
R7881 gnd.n2514 gnd.n2504 585
R7882 gnd.n3273 gnd.n2527 585
R7883 gnd.n2527 gnd.n2513 585
R7884 gnd.n3275 gnd.n3274 585
R7885 gnd.n3276 gnd.n3275 585
R7886 gnd.n2528 gnd.n2526 585
R7887 gnd.n2535 gnd.n2526 585
R7888 gnd.n3268 gnd.n3267 585
R7889 gnd.n3267 gnd.n3266 585
R7890 gnd.n2531 gnd.n2530 585
R7891 gnd.n3247 gnd.n2531 585
R7892 gnd.n3233 gnd.n2554 585
R7893 gnd.n2554 gnd.n2544 585
R7894 gnd.n3235 gnd.n3234 585
R7895 gnd.n3236 gnd.n3235 585
R7896 gnd.n2555 gnd.n2553 585
R7897 gnd.n3224 gnd.n2553 585
R7898 gnd.n3228 gnd.n3227 585
R7899 gnd.n3227 gnd.n3226 585
R7900 gnd.n2558 gnd.n2557 585
R7901 gnd.n3179 gnd.n2558 585
R7902 gnd.n2672 gnd.n2671 585
R7903 gnd.n2673 gnd.n2672 585
R7904 gnd.n2652 gnd.n2651 585
R7905 gnd.n2655 gnd.n2652 585
R7906 gnd.n3189 gnd.n3188 585
R7907 gnd.n3188 gnd.n3187 585
R7908 gnd.n3190 gnd.n2646 585
R7909 gnd.n2682 gnd.n2646 585
R7910 gnd.n3192 gnd.n3191 585
R7911 gnd.n3193 gnd.n3192 585
R7912 gnd.n2647 gnd.n2645 585
R7913 gnd.n3157 gnd.n2645 585
R7914 gnd.n3141 gnd.n3140 585
R7915 gnd.n3140 gnd.n2633 585
R7916 gnd.n3142 gnd.n2697 585
R7917 gnd.n2697 gnd.n2632 585
R7918 gnd.n3144 gnd.n3143 585
R7919 gnd.n3145 gnd.n3144 585
R7920 gnd.n2698 gnd.n2696 585
R7921 gnd.n2696 gnd.n2693 585
R7922 gnd.n3133 gnd.n3132 585
R7923 gnd.n3132 gnd.n3131 585
R7924 gnd.n2701 gnd.n2700 585
R7925 gnd.n2708 gnd.n2701 585
R7926 gnd.n3107 gnd.n3106 585
R7927 gnd.n3108 gnd.n3107 585
R7928 gnd.n2720 gnd.n2719 585
R7929 gnd.n2727 gnd.n2719 585
R7930 gnd.n3102 gnd.n3101 585
R7931 gnd.n3101 gnd.n3100 585
R7932 gnd.n2723 gnd.n2722 585
R7933 gnd.n3090 gnd.n2723 585
R7934 gnd.n3077 gnd.n2747 585
R7935 gnd.n2747 gnd.n2746 585
R7936 gnd.n3079 gnd.n3078 585
R7937 gnd.n3080 gnd.n3079 585
R7938 gnd.n2748 gnd.n2745 585
R7939 gnd.n2755 gnd.n2745 585
R7940 gnd.n3072 gnd.n3071 585
R7941 gnd.n3071 gnd.n3070 585
R7942 gnd.n2751 gnd.n2750 585
R7943 gnd.n3059 gnd.n2751 585
R7944 gnd.n3046 gnd.n2772 585
R7945 gnd.n2772 gnd.n2771 585
R7946 gnd.n3048 gnd.n3047 585
R7947 gnd.n3049 gnd.n3048 585
R7948 gnd.n3042 gnd.n2770 585
R7949 gnd.n3041 gnd.n3040 585
R7950 gnd.n2775 gnd.n2774 585
R7951 gnd.n3038 gnd.n2775 585
R7952 gnd.n2797 gnd.n2796 585
R7953 gnd.n2800 gnd.n2799 585
R7954 gnd.n2798 gnd.n2793 585
R7955 gnd.n2805 gnd.n2804 585
R7956 gnd.n2807 gnd.n2806 585
R7957 gnd.n2810 gnd.n2809 585
R7958 gnd.n2808 gnd.n2791 585
R7959 gnd.n2815 gnd.n2814 585
R7960 gnd.n2817 gnd.n2816 585
R7961 gnd.n2820 gnd.n2819 585
R7962 gnd.n2818 gnd.n2789 585
R7963 gnd.n2825 gnd.n2824 585
R7964 gnd.n2829 gnd.n2826 585
R7965 gnd.n2830 gnd.n2767 585
R7966 gnd.n3708 gnd.n2371 585
R7967 gnd.n3775 gnd.n3774 585
R7968 gnd.n3777 gnd.n3776 585
R7969 gnd.n3779 gnd.n3778 585
R7970 gnd.n3781 gnd.n3780 585
R7971 gnd.n3783 gnd.n3782 585
R7972 gnd.n3785 gnd.n3784 585
R7973 gnd.n3787 gnd.n3786 585
R7974 gnd.n3789 gnd.n3788 585
R7975 gnd.n3791 gnd.n3790 585
R7976 gnd.n3793 gnd.n3792 585
R7977 gnd.n3795 gnd.n3794 585
R7978 gnd.n3797 gnd.n3796 585
R7979 gnd.n3800 gnd.n3799 585
R7980 gnd.n3798 gnd.n2359 585
R7981 gnd.n3804 gnd.n2357 585
R7982 gnd.n3806 gnd.n3805 585
R7983 gnd.n3807 gnd.n3806 585
R7984 gnd.n3709 gnd.n2413 585
R7985 gnd.n3709 gnd.n2408 585
R7986 gnd.n3711 gnd.n3710 585
R7987 gnd.n3710 gnd.n2407 585
R7988 gnd.n3707 gnd.n2412 585
R7989 gnd.n3707 gnd.n3706 585
R7990 gnd.n3686 gnd.n2414 585
R7991 gnd.n2426 gnd.n2414 585
R7992 gnd.n3685 gnd.n2424 585
R7993 gnd.n3694 gnd.n2424 585
R7994 gnd.n3420 gnd.n2431 585
R7995 gnd.n3421 gnd.n3420 585
R7996 gnd.n3419 gnd.n3418 585
R7997 gnd.n3419 gnd.n2435 585
R7998 gnd.n3417 gnd.n2437 585
R7999 gnd.n3410 gnd.n2437 585
R8000 gnd.n2450 gnd.n2438 585
R8001 gnd.n2450 gnd.n2442 585
R8002 gnd.n3366 gnd.n2451 585
R8003 gnd.n3400 gnd.n2451 585
R8004 gnd.n3365 gnd.n3364 585
R8005 gnd.n3364 gnd.n2458 585
R8006 gnd.n3363 gnd.n2466 585
R8007 gnd.n3363 gnd.n2457 585
R8008 gnd.n3362 gnd.n2468 585
R8009 gnd.n3362 gnd.n3361 585
R8010 gnd.n3341 gnd.n2467 585
R8011 gnd.n2480 gnd.n2467 585
R8012 gnd.n3340 gnd.n2478 585
R8013 gnd.n3351 gnd.n2478 585
R8014 gnd.n3331 gnd.n2485 585
R8015 gnd.n3332 gnd.n3331 585
R8016 gnd.n3330 gnd.n3329 585
R8017 gnd.n3330 gnd.n2489 585
R8018 gnd.n3328 gnd.n2491 585
R8019 gnd.n3321 gnd.n2491 585
R8020 gnd.n2506 gnd.n2492 585
R8021 gnd.n2506 gnd.n2496 585
R8022 gnd.n3281 gnd.n2507 585
R8023 gnd.n3311 gnd.n2507 585
R8024 gnd.n3280 gnd.n3279 585
R8025 gnd.n3279 gnd.n2514 585
R8026 gnd.n3278 gnd.n2521 585
R8027 gnd.n3278 gnd.n2513 585
R8028 gnd.n3277 gnd.n2523 585
R8029 gnd.n3277 gnd.n3276 585
R8030 gnd.n3256 gnd.n2522 585
R8031 gnd.n2535 gnd.n2522 585
R8032 gnd.n3255 gnd.n2533 585
R8033 gnd.n3266 gnd.n2533 585
R8034 gnd.n3246 gnd.n2540 585
R8035 gnd.n3247 gnd.n3246 585
R8036 gnd.n3245 gnd.n3244 585
R8037 gnd.n3245 gnd.n2544 585
R8038 gnd.n3243 gnd.n2546 585
R8039 gnd.n3236 gnd.n2546 585
R8040 gnd.n3223 gnd.n2547 585
R8041 gnd.n3224 gnd.n3223 585
R8042 gnd.n3176 gnd.n2560 585
R8043 gnd.n3226 gnd.n2560 585
R8044 gnd.n3178 gnd.n3177 585
R8045 gnd.n3179 gnd.n3178 585
R8046 gnd.n3171 gnd.n2674 585
R8047 gnd.n2674 gnd.n2673 585
R8048 gnd.n3169 gnd.n3168 585
R8049 gnd.n3168 gnd.n2655 585
R8050 gnd.n3166 gnd.n2653 585
R8051 gnd.n3187 gnd.n2653 585
R8052 gnd.n2684 gnd.n2683 585
R8053 gnd.n2683 gnd.n2682 585
R8054 gnd.n3160 gnd.n2643 585
R8055 gnd.n3193 gnd.n2643 585
R8056 gnd.n3159 gnd.n3158 585
R8057 gnd.n3158 gnd.n3157 585
R8058 gnd.n3155 gnd.n2686 585
R8059 gnd.n3155 gnd.n2633 585
R8060 gnd.n3154 gnd.n3153 585
R8061 gnd.n3154 gnd.n2632 585
R8062 gnd.n2689 gnd.n2688 585
R8063 gnd.n3145 gnd.n2688 585
R8064 gnd.n3113 gnd.n3112 585
R8065 gnd.n3112 gnd.n2693 585
R8066 gnd.n3114 gnd.n2702 585
R8067 gnd.n3131 gnd.n2702 585
R8068 gnd.n3111 gnd.n3110 585
R8069 gnd.n3110 gnd.n2708 585
R8070 gnd.n3109 gnd.n2716 585
R8071 gnd.n3109 gnd.n3108 585
R8072 gnd.n3094 gnd.n2717 585
R8073 gnd.n2727 gnd.n2717 585
R8074 gnd.n3093 gnd.n2725 585
R8075 gnd.n3100 gnd.n2725 585
R8076 gnd.n3092 gnd.n3091 585
R8077 gnd.n3091 gnd.n3090 585
R8078 gnd.n2736 gnd.n2733 585
R8079 gnd.n2746 gnd.n2736 585
R8080 gnd.n3082 gnd.n3081 585
R8081 gnd.n3081 gnd.n3080 585
R8082 gnd.n2742 gnd.n2741 585
R8083 gnd.n2755 gnd.n2742 585
R8084 gnd.n3062 gnd.n2753 585
R8085 gnd.n3070 gnd.n2753 585
R8086 gnd.n3061 gnd.n3060 585
R8087 gnd.n3060 gnd.n3059 585
R8088 gnd.n2762 gnd.n2760 585
R8089 gnd.n2771 gnd.n2762 585
R8090 gnd.n3051 gnd.n3050 585
R8091 gnd.n3050 gnd.n3049 585
R8092 gnd.n6465 gnd.n6464 585
R8093 gnd.n6464 gnd.n6463 585
R8094 gnd.n6466 gnd.n1103 585
R8095 gnd.n4568 gnd.n1103 585
R8096 gnd.n6468 gnd.n6467 585
R8097 gnd.n6469 gnd.n6468 585
R8098 gnd.n1088 gnd.n1087 585
R8099 gnd.n4528 gnd.n1088 585
R8100 gnd.n6477 gnd.n6476 585
R8101 gnd.n6476 gnd.n6475 585
R8102 gnd.n6478 gnd.n1082 585
R8103 gnd.n4519 gnd.n1082 585
R8104 gnd.n6480 gnd.n6479 585
R8105 gnd.n6481 gnd.n6480 585
R8106 gnd.n1067 gnd.n1066 585
R8107 gnd.n4511 gnd.n1067 585
R8108 gnd.n6489 gnd.n6488 585
R8109 gnd.n6488 gnd.n6487 585
R8110 gnd.n6490 gnd.n1061 585
R8111 gnd.n4446 gnd.n1061 585
R8112 gnd.n6492 gnd.n6491 585
R8113 gnd.n6493 gnd.n6492 585
R8114 gnd.n1046 gnd.n1045 585
R8115 gnd.n4434 gnd.n1046 585
R8116 gnd.n6501 gnd.n6500 585
R8117 gnd.n6500 gnd.n6499 585
R8118 gnd.n6502 gnd.n1040 585
R8119 gnd.n4457 gnd.n1040 585
R8120 gnd.n6504 gnd.n6503 585
R8121 gnd.n6505 gnd.n6504 585
R8122 gnd.n1025 gnd.n1024 585
R8123 gnd.n4426 gnd.n1025 585
R8124 gnd.n6513 gnd.n6512 585
R8125 gnd.n6512 gnd.n6511 585
R8126 gnd.n6514 gnd.n1019 585
R8127 gnd.n4393 gnd.n1019 585
R8128 gnd.n6516 gnd.n6515 585
R8129 gnd.n6517 gnd.n6516 585
R8130 gnd.n1004 gnd.n1003 585
R8131 gnd.n4385 gnd.n1004 585
R8132 gnd.n6525 gnd.n6524 585
R8133 gnd.n6524 gnd.n6523 585
R8134 gnd.n6526 gnd.n998 585
R8135 gnd.n4408 gnd.n998 585
R8136 gnd.n6528 gnd.n6527 585
R8137 gnd.n6529 gnd.n6528 585
R8138 gnd.n982 gnd.n981 585
R8139 gnd.n4377 gnd.n982 585
R8140 gnd.n6537 gnd.n6536 585
R8141 gnd.n6536 gnd.n6535 585
R8142 gnd.n6538 gnd.n976 585
R8143 gnd.n4359 gnd.n976 585
R8144 gnd.n6540 gnd.n6539 585
R8145 gnd.n6541 gnd.n6540 585
R8146 gnd.n977 gnd.n975 585
R8147 gnd.n975 gnd.n970 585
R8148 gnd.n4349 gnd.n4348 585
R8149 gnd.n4350 gnd.n4349 585
R8150 gnd.n4346 gnd.n2187 585
R8151 gnd.n2193 gnd.n2187 585
R8152 gnd.n4345 gnd.n4344 585
R8153 gnd.n4344 gnd.n4343 585
R8154 gnd.n4321 gnd.n2189 585
R8155 gnd.n2211 gnd.n2189 585
R8156 gnd.n4323 gnd.n4322 585
R8157 gnd.n4324 gnd.n4323 585
R8158 gnd.n4319 gnd.n2213 585
R8159 gnd.n2213 gnd.n2209 585
R8160 gnd.n4318 gnd.n4317 585
R8161 gnd.n4317 gnd.n4316 585
R8162 gnd.n4304 gnd.n2215 585
R8163 gnd.n2216 gnd.n2215 585
R8164 gnd.n4306 gnd.n4305 585
R8165 gnd.n4307 gnd.n4306 585
R8166 gnd.n4302 gnd.n2228 585
R8167 gnd.n2228 gnd.n2225 585
R8168 gnd.n4301 gnd.n4300 585
R8169 gnd.n4300 gnd.n4299 585
R8170 gnd.n2231 gnd.n2229 585
R8171 gnd.n2242 gnd.n2231 585
R8172 gnd.n4290 gnd.n4289 585
R8173 gnd.n4291 gnd.n4290 585
R8174 gnd.n2244 gnd.n2243 585
R8175 gnd.n2243 gnd.n2239 585
R8176 gnd.n4284 gnd.n4283 585
R8177 gnd.n4283 gnd.n4282 585
R8178 gnd.n2247 gnd.n2246 585
R8179 gnd.n2248 gnd.n2247 585
R8180 gnd.n4273 gnd.n4272 585
R8181 gnd.n4274 gnd.n4273 585
R8182 gnd.n2260 gnd.n2259 585
R8183 gnd.n2259 gnd.n2256 585
R8184 gnd.n4268 gnd.n4267 585
R8185 gnd.n4267 gnd.n4266 585
R8186 gnd.n2263 gnd.n2262 585
R8187 gnd.n2274 gnd.n2263 585
R8188 gnd.n4257 gnd.n4256 585
R8189 gnd.n4258 gnd.n4257 585
R8190 gnd.n2276 gnd.n2275 585
R8191 gnd.n2275 gnd.n2271 585
R8192 gnd.n4252 gnd.n4251 585
R8193 gnd.n4251 gnd.n4250 585
R8194 gnd.n2279 gnd.n2278 585
R8195 gnd.n2280 gnd.n2279 585
R8196 gnd.n4241 gnd.n4240 585
R8197 gnd.n4242 gnd.n4241 585
R8198 gnd.n2292 gnd.n2291 585
R8199 gnd.n2291 gnd.n2288 585
R8200 gnd.n4236 gnd.n4235 585
R8201 gnd.n4235 gnd.n4234 585
R8202 gnd.n2295 gnd.n2294 585
R8203 gnd.n2306 gnd.n2295 585
R8204 gnd.n4225 gnd.n4224 585
R8205 gnd.n4226 gnd.n4225 585
R8206 gnd.n2308 gnd.n2307 585
R8207 gnd.n2307 gnd.n2303 585
R8208 gnd.n4220 gnd.n4219 585
R8209 gnd.n4219 gnd.n4218 585
R8210 gnd.n2311 gnd.n2310 585
R8211 gnd.n2312 gnd.n2311 585
R8212 gnd.n4209 gnd.n4208 585
R8213 gnd.n4210 gnd.n4209 585
R8214 gnd.n2324 gnd.n2323 585
R8215 gnd.n2323 gnd.n2320 585
R8216 gnd.n4204 gnd.n4203 585
R8217 gnd.n4203 gnd.n4202 585
R8218 gnd.n2327 gnd.n2326 585
R8219 gnd.n3972 gnd.n2327 585
R8220 gnd.n4193 gnd.n4192 585
R8221 gnd.n4194 gnd.n4193 585
R8222 gnd.n4189 gnd.n3973 585
R8223 gnd.n4188 gnd.n4187 585
R8224 gnd.n4185 gnd.n3975 585
R8225 gnd.n4185 gnd.n3808 585
R8226 gnd.n4184 gnd.n4183 585
R8227 gnd.n4182 gnd.n4181 585
R8228 gnd.n4180 gnd.n3980 585
R8229 gnd.n4178 gnd.n4177 585
R8230 gnd.n4176 gnd.n3981 585
R8231 gnd.n4175 gnd.n4174 585
R8232 gnd.n4172 gnd.n3986 585
R8233 gnd.n4170 gnd.n4169 585
R8234 gnd.n4168 gnd.n3987 585
R8235 gnd.n4167 gnd.n4166 585
R8236 gnd.n4164 gnd.n3992 585
R8237 gnd.n4162 gnd.n4161 585
R8238 gnd.n4160 gnd.n3993 585
R8239 gnd.n4159 gnd.n4158 585
R8240 gnd.n4156 gnd.n3998 585
R8241 gnd.n4154 gnd.n4153 585
R8242 gnd.n4152 gnd.n3999 585
R8243 gnd.n4151 gnd.n4150 585
R8244 gnd.n4148 gnd.n4007 585
R8245 gnd.n4146 gnd.n4145 585
R8246 gnd.n4144 gnd.n4008 585
R8247 gnd.n4143 gnd.n4142 585
R8248 gnd.n4140 gnd.n4013 585
R8249 gnd.n4138 gnd.n4137 585
R8250 gnd.n4136 gnd.n4014 585
R8251 gnd.n4135 gnd.n4134 585
R8252 gnd.n4132 gnd.n4019 585
R8253 gnd.n4130 gnd.n4129 585
R8254 gnd.n4128 gnd.n4020 585
R8255 gnd.n4127 gnd.n4126 585
R8256 gnd.n4124 gnd.n4025 585
R8257 gnd.n4122 gnd.n4121 585
R8258 gnd.n4120 gnd.n4026 585
R8259 gnd.n4119 gnd.n4031 585
R8260 gnd.n4112 gnd.n4034 585
R8261 gnd.n4115 gnd.n4114 585
R8262 gnd.n2119 gnd.n2118 585
R8263 gnd.n4576 gnd.n4575 585
R8264 gnd.n4578 gnd.n4577 585
R8265 gnd.n4580 gnd.n4579 585
R8266 gnd.n4582 gnd.n4581 585
R8267 gnd.n4584 gnd.n4583 585
R8268 gnd.n4586 gnd.n4585 585
R8269 gnd.n4588 gnd.n4587 585
R8270 gnd.n4590 gnd.n4589 585
R8271 gnd.n4592 gnd.n4591 585
R8272 gnd.n4594 gnd.n4593 585
R8273 gnd.n4596 gnd.n4595 585
R8274 gnd.n4598 gnd.n4597 585
R8275 gnd.n4600 gnd.n4599 585
R8276 gnd.n4602 gnd.n4601 585
R8277 gnd.n4604 gnd.n4603 585
R8278 gnd.n4606 gnd.n4605 585
R8279 gnd.n4608 gnd.n4607 585
R8280 gnd.n4610 gnd.n4609 585
R8281 gnd.n4613 gnd.n4612 585
R8282 gnd.n4611 gnd.n2097 585
R8283 gnd.n5529 gnd.n5528 585
R8284 gnd.n5531 gnd.n5530 585
R8285 gnd.n5533 gnd.n5532 585
R8286 gnd.n5535 gnd.n5534 585
R8287 gnd.n5537 gnd.n5536 585
R8288 gnd.n5539 gnd.n5538 585
R8289 gnd.n5541 gnd.n5540 585
R8290 gnd.n5543 gnd.n5542 585
R8291 gnd.n5545 gnd.n5544 585
R8292 gnd.n5547 gnd.n5546 585
R8293 gnd.n5549 gnd.n5548 585
R8294 gnd.n5551 gnd.n5550 585
R8295 gnd.n5552 gnd.n2078 585
R8296 gnd.n5554 gnd.n5553 585
R8297 gnd.n2079 gnd.n2077 585
R8298 gnd.n2080 gnd.n1108 585
R8299 gnd.n5556 gnd.n1108 585
R8300 gnd.n4571 gnd.n1110 585
R8301 gnd.n6463 gnd.n1110 585
R8302 gnd.n4570 gnd.n4569 585
R8303 gnd.n4569 gnd.n4568 585
R8304 gnd.n2123 gnd.n1101 585
R8305 gnd.n6469 gnd.n1101 585
R8306 gnd.n4527 gnd.n4526 585
R8307 gnd.n4528 gnd.n4527 585
R8308 gnd.n2129 gnd.n1090 585
R8309 gnd.n6475 gnd.n1090 585
R8310 gnd.n4521 gnd.n4520 585
R8311 gnd.n4520 gnd.n4519 585
R8312 gnd.n2131 gnd.n1079 585
R8313 gnd.n6481 gnd.n1079 585
R8314 gnd.n4442 gnd.n2135 585
R8315 gnd.n4511 gnd.n2135 585
R8316 gnd.n4443 gnd.n1069 585
R8317 gnd.n6487 gnd.n1069 585
R8318 gnd.n4445 gnd.n4444 585
R8319 gnd.n4446 gnd.n4445 585
R8320 gnd.n2152 gnd.n1058 585
R8321 gnd.n6493 gnd.n1058 585
R8322 gnd.n4436 gnd.n4435 585
R8323 gnd.n4435 gnd.n4434 585
R8324 gnd.n4433 gnd.n1047 585
R8325 gnd.n6499 gnd.n1047 585
R8326 gnd.n4432 gnd.n2146 585
R8327 gnd.n4457 gnd.n2146 585
R8328 gnd.n2154 gnd.n1037 585
R8329 gnd.n6505 gnd.n1037 585
R8330 gnd.n4428 gnd.n4427 585
R8331 gnd.n4427 gnd.n4426 585
R8332 gnd.n2156 gnd.n1027 585
R8333 gnd.n6511 gnd.n1027 585
R8334 gnd.n4392 gnd.n4391 585
R8335 gnd.n4393 gnd.n4392 585
R8336 gnd.n2173 gnd.n1016 585
R8337 gnd.n6517 gnd.n1016 585
R8338 gnd.n4387 gnd.n4386 585
R8339 gnd.n4386 gnd.n4385 585
R8340 gnd.n4384 gnd.n1005 585
R8341 gnd.n6523 gnd.n1005 585
R8342 gnd.n4383 gnd.n2167 585
R8343 gnd.n4408 gnd.n2167 585
R8344 gnd.n2175 gnd.n995 585
R8345 gnd.n6529 gnd.n995 585
R8346 gnd.n4379 gnd.n4378 585
R8347 gnd.n4378 gnd.n4377 585
R8348 gnd.n2177 gnd.n984 585
R8349 gnd.n6535 gnd.n984 585
R8350 gnd.n4358 gnd.n4357 585
R8351 gnd.n4359 gnd.n4358 585
R8352 gnd.n2181 gnd.n971 585
R8353 gnd.n6541 gnd.n971 585
R8354 gnd.n4353 gnd.n4352 585
R8355 gnd.n4352 gnd.n970 585
R8356 gnd.n4351 gnd.n2183 585
R8357 gnd.n4351 gnd.n4350 585
R8358 gnd.n2204 gnd.n2184 585
R8359 gnd.n2193 gnd.n2184 585
R8360 gnd.n2205 gnd.n2190 585
R8361 gnd.n4343 gnd.n2190 585
R8362 gnd.n2208 gnd.n2206 585
R8363 gnd.n2211 gnd.n2208 585
R8364 gnd.n4326 gnd.n4325 585
R8365 gnd.n4325 gnd.n4324 585
R8366 gnd.n2207 gnd.n2201 585
R8367 gnd.n2209 gnd.n2207 585
R8368 gnd.n4066 gnd.n2217 585
R8369 gnd.n4316 gnd.n2217 585
R8370 gnd.n4068 gnd.n4067 585
R8371 gnd.n4067 gnd.n2216 585
R8372 gnd.n4069 gnd.n2226 585
R8373 gnd.n4307 gnd.n2226 585
R8374 gnd.n4071 gnd.n4070 585
R8375 gnd.n4070 gnd.n2225 585
R8376 gnd.n4072 gnd.n2232 585
R8377 gnd.n4299 gnd.n2232 585
R8378 gnd.n4074 gnd.n4073 585
R8379 gnd.n4073 gnd.n2242 585
R8380 gnd.n4075 gnd.n2240 585
R8381 gnd.n4291 gnd.n2240 585
R8382 gnd.n4077 gnd.n4076 585
R8383 gnd.n4076 gnd.n2239 585
R8384 gnd.n4078 gnd.n2249 585
R8385 gnd.n4282 gnd.n2249 585
R8386 gnd.n4080 gnd.n4079 585
R8387 gnd.n4079 gnd.n2248 585
R8388 gnd.n4081 gnd.n2257 585
R8389 gnd.n4274 gnd.n2257 585
R8390 gnd.n4083 gnd.n4082 585
R8391 gnd.n4082 gnd.n2256 585
R8392 gnd.n4084 gnd.n2264 585
R8393 gnd.n4266 gnd.n2264 585
R8394 gnd.n4086 gnd.n4085 585
R8395 gnd.n4085 gnd.n2274 585
R8396 gnd.n4087 gnd.n2272 585
R8397 gnd.n4258 gnd.n2272 585
R8398 gnd.n4089 gnd.n4088 585
R8399 gnd.n4088 gnd.n2271 585
R8400 gnd.n4090 gnd.n2281 585
R8401 gnd.n4250 gnd.n2281 585
R8402 gnd.n4092 gnd.n4091 585
R8403 gnd.n4091 gnd.n2280 585
R8404 gnd.n4093 gnd.n2289 585
R8405 gnd.n4242 gnd.n2289 585
R8406 gnd.n4095 gnd.n4094 585
R8407 gnd.n4094 gnd.n2288 585
R8408 gnd.n4096 gnd.n2296 585
R8409 gnd.n4234 gnd.n2296 585
R8410 gnd.n4098 gnd.n4097 585
R8411 gnd.n4097 gnd.n2306 585
R8412 gnd.n4099 gnd.n2304 585
R8413 gnd.n4226 gnd.n2304 585
R8414 gnd.n4101 gnd.n4100 585
R8415 gnd.n4100 gnd.n2303 585
R8416 gnd.n4102 gnd.n2313 585
R8417 gnd.n4218 gnd.n2313 585
R8418 gnd.n4104 gnd.n4103 585
R8419 gnd.n4103 gnd.n2312 585
R8420 gnd.n4105 gnd.n2321 585
R8421 gnd.n4210 gnd.n2321 585
R8422 gnd.n4107 gnd.n4106 585
R8423 gnd.n4106 gnd.n2320 585
R8424 gnd.n4108 gnd.n2328 585
R8425 gnd.n4202 gnd.n2328 585
R8426 gnd.n4109 gnd.n4036 585
R8427 gnd.n4036 gnd.n3972 585
R8428 gnd.n4110 gnd.n3809 585
R8429 gnd.n4194 gnd.n3809 585
R8430 gnd.n7803 gnd.n7802 585
R8431 gnd.n7804 gnd.n7803 585
R8432 gnd.n132 gnd.n130 585
R8433 gnd.n130 gnd.n126 585
R8434 gnd.n7723 gnd.n7722 585
R8435 gnd.n7724 gnd.n7723 585
R8436 gnd.n209 gnd.n208 585
R8437 gnd.n208 gnd.n206 585
R8438 gnd.n7718 gnd.n7717 585
R8439 gnd.n7717 gnd.n7716 585
R8440 gnd.n212 gnd.n211 585
R8441 gnd.n213 gnd.n212 585
R8442 gnd.n7639 gnd.n7638 585
R8443 gnd.n7640 gnd.n7639 585
R8444 gnd.n225 gnd.n224 585
R8445 gnd.n232 gnd.n224 585
R8446 gnd.n7634 gnd.n7633 585
R8447 gnd.n7633 gnd.n7632 585
R8448 gnd.n228 gnd.n227 585
R8449 gnd.n229 gnd.n228 585
R8450 gnd.n7623 gnd.n7622 585
R8451 gnd.n7624 gnd.n7623 585
R8452 gnd.n241 gnd.n240 585
R8453 gnd.n247 gnd.n240 585
R8454 gnd.n7618 gnd.n7617 585
R8455 gnd.n7617 gnd.n7616 585
R8456 gnd.n244 gnd.n243 585
R8457 gnd.n254 gnd.n244 585
R8458 gnd.n7607 gnd.n7606 585
R8459 gnd.n7608 gnd.n7607 585
R8460 gnd.n256 gnd.n255 585
R8461 gnd.n263 gnd.n255 585
R8462 gnd.n7602 gnd.n7601 585
R8463 gnd.n7601 gnd.n7600 585
R8464 gnd.n259 gnd.n258 585
R8465 gnd.n260 gnd.n259 585
R8466 gnd.n7591 gnd.n7590 585
R8467 gnd.n7592 gnd.n7591 585
R8468 gnd.n272 gnd.n271 585
R8469 gnd.n271 gnd.n269 585
R8470 gnd.n7586 gnd.n7585 585
R8471 gnd.n7585 gnd.n7584 585
R8472 gnd.n275 gnd.n274 585
R8473 gnd.n284 gnd.n275 585
R8474 gnd.n7575 gnd.n7574 585
R8475 gnd.n7576 gnd.n7575 585
R8476 gnd.n286 gnd.n285 585
R8477 gnd.n293 gnd.n285 585
R8478 gnd.n7570 gnd.n7569 585
R8479 gnd.n7569 gnd.n7568 585
R8480 gnd.n289 gnd.n288 585
R8481 gnd.n290 gnd.n289 585
R8482 gnd.n7559 gnd.n7558 585
R8483 gnd.n7560 gnd.n7559 585
R8484 gnd.n302 gnd.n301 585
R8485 gnd.n301 gnd.n299 585
R8486 gnd.n7535 gnd.n7534 585
R8487 gnd.n7536 gnd.n7535 585
R8488 gnd.n7533 gnd.n332 585
R8489 gnd.n7533 gnd.n7532 585
R8490 gnd.n331 gnd.n330 585
R8491 gnd.n334 gnd.n330 585
R8492 gnd.n7458 gnd.n7457 585
R8493 gnd.n7459 gnd.n7458 585
R8494 gnd.n7456 gnd.n7455 585
R8495 gnd.n7455 gnd.n340 585
R8496 gnd.n7454 gnd.n342 585
R8497 gnd.n7454 gnd.n7453 585
R8498 gnd.n341 gnd.n311 585
R8499 gnd.n315 gnd.n311 585
R8500 gnd.n7553 gnd.n7552 585
R8501 gnd.n7552 gnd.n7551 585
R8502 gnd.n7554 gnd.n310 585
R8503 gnd.n7444 gnd.n310 585
R8504 gnd.n361 gnd.n309 585
R8505 gnd.n361 gnd.n350 585
R8506 gnd.n7428 gnd.n7427 585
R8507 gnd.n7429 gnd.n7428 585
R8508 gnd.n7426 gnd.n360 585
R8509 gnd.n7408 gnd.n360 585
R8510 gnd.n366 gnd.n362 585
R8511 gnd.n7392 gnd.n366 585
R8512 gnd.n7422 gnd.n7421 585
R8513 gnd.n7421 gnd.n7420 585
R8514 gnd.n365 gnd.n364 585
R8515 gnd.n7398 gnd.n365 585
R8516 gnd.n7381 gnd.n394 585
R8517 gnd.n7365 gnd.n394 585
R8518 gnd.n7383 gnd.n7382 585
R8519 gnd.n7384 gnd.n7383 585
R8520 gnd.n395 gnd.n393 585
R8521 gnd.n6143 gnd.n393 585
R8522 gnd.n7376 gnd.n7375 585
R8523 gnd.n7375 gnd.n7374 585
R8524 gnd.n398 gnd.n397 585
R8525 gnd.n6138 gnd.n398 585
R8526 gnd.n6188 gnd.n6187 585
R8527 gnd.n6189 gnd.n6188 585
R8528 gnd.n1366 gnd.n1365 585
R8529 gnd.n1373 gnd.n1365 585
R8530 gnd.n6183 gnd.n6182 585
R8531 gnd.n6182 gnd.n6181 585
R8532 gnd.n1369 gnd.n1368 585
R8533 gnd.n6159 gnd.n1369 585
R8534 gnd.n6118 gnd.n1399 585
R8535 gnd.n1399 gnd.n1398 585
R8536 gnd.n6120 gnd.n6119 585
R8537 gnd.n6121 gnd.n6120 585
R8538 gnd.n1400 gnd.n1397 585
R8539 gnd.n1407 gnd.n1397 585
R8540 gnd.n6113 gnd.n6112 585
R8541 gnd.n6112 gnd.n6111 585
R8542 gnd.n1403 gnd.n1402 585
R8543 gnd.n6098 gnd.n1403 585
R8544 gnd.n6081 gnd.n1426 585
R8545 gnd.n1426 gnd.n1414 585
R8546 gnd.n6083 gnd.n6082 585
R8547 gnd.n6084 gnd.n6083 585
R8548 gnd.n1427 gnd.n1425 585
R8549 gnd.n1435 gnd.n1425 585
R8550 gnd.n6076 gnd.n6075 585
R8551 gnd.n6075 gnd.n6074 585
R8552 gnd.n1430 gnd.n1429 585
R8553 gnd.n6062 gnd.n1430 585
R8554 gnd.n6050 gnd.n6045 585
R8555 gnd.n6045 gnd.n1452 585
R8556 gnd.n6052 gnd.n6051 585
R8557 gnd.n6053 gnd.n6052 585
R8558 gnd.n6046 gnd.n1288 585
R8559 gnd.n6218 gnd.n1288 585
R8560 gnd.n6292 gnd.n6291 585
R8561 gnd.n6290 gnd.n1287 585
R8562 gnd.n6289 gnd.n1286 585
R8563 gnd.n6294 gnd.n1286 585
R8564 gnd.n6288 gnd.n6287 585
R8565 gnd.n6286 gnd.n6285 585
R8566 gnd.n6284 gnd.n6283 585
R8567 gnd.n6282 gnd.n6281 585
R8568 gnd.n6280 gnd.n6279 585
R8569 gnd.n6278 gnd.n6277 585
R8570 gnd.n6276 gnd.n6275 585
R8571 gnd.n6274 gnd.n6273 585
R8572 gnd.n6272 gnd.n6271 585
R8573 gnd.n6270 gnd.n6269 585
R8574 gnd.n6268 gnd.n6267 585
R8575 gnd.n6266 gnd.n6265 585
R8576 gnd.n6264 gnd.n6263 585
R8577 gnd.n6261 gnd.n6260 585
R8578 gnd.n6259 gnd.n6258 585
R8579 gnd.n6257 gnd.n6256 585
R8580 gnd.n6255 gnd.n6254 585
R8581 gnd.n6253 gnd.n6252 585
R8582 gnd.n6251 gnd.n6250 585
R8583 gnd.n6249 gnd.n6248 585
R8584 gnd.n6247 gnd.n6246 585
R8585 gnd.n6245 gnd.n6244 585
R8586 gnd.n6243 gnd.n6242 585
R8587 gnd.n6241 gnd.n6240 585
R8588 gnd.n6239 gnd.n6238 585
R8589 gnd.n6237 gnd.n6236 585
R8590 gnd.n6235 gnd.n6234 585
R8591 gnd.n6233 gnd.n6232 585
R8592 gnd.n6231 gnd.n6230 585
R8593 gnd.n6229 gnd.n6228 585
R8594 gnd.n6227 gnd.n6226 585
R8595 gnd.n6225 gnd.n1328 585
R8596 gnd.n1332 gnd.n1329 585
R8597 gnd.n6221 gnd.n6220 585
R8598 gnd.n200 gnd.n199 585
R8599 gnd.n7732 gnd.n195 585
R8600 gnd.n7734 gnd.n7733 585
R8601 gnd.n7736 gnd.n193 585
R8602 gnd.n7738 gnd.n7737 585
R8603 gnd.n7739 gnd.n188 585
R8604 gnd.n7741 gnd.n7740 585
R8605 gnd.n7743 gnd.n186 585
R8606 gnd.n7745 gnd.n7744 585
R8607 gnd.n7746 gnd.n181 585
R8608 gnd.n7748 gnd.n7747 585
R8609 gnd.n7750 gnd.n179 585
R8610 gnd.n7752 gnd.n7751 585
R8611 gnd.n7753 gnd.n174 585
R8612 gnd.n7755 gnd.n7754 585
R8613 gnd.n7757 gnd.n172 585
R8614 gnd.n7759 gnd.n7758 585
R8615 gnd.n7760 gnd.n167 585
R8616 gnd.n7762 gnd.n7761 585
R8617 gnd.n7764 gnd.n165 585
R8618 gnd.n7766 gnd.n7765 585
R8619 gnd.n7770 gnd.n160 585
R8620 gnd.n7772 gnd.n7771 585
R8621 gnd.n7774 gnd.n158 585
R8622 gnd.n7776 gnd.n7775 585
R8623 gnd.n7777 gnd.n153 585
R8624 gnd.n7779 gnd.n7778 585
R8625 gnd.n7781 gnd.n151 585
R8626 gnd.n7783 gnd.n7782 585
R8627 gnd.n7784 gnd.n146 585
R8628 gnd.n7786 gnd.n7785 585
R8629 gnd.n7788 gnd.n144 585
R8630 gnd.n7790 gnd.n7789 585
R8631 gnd.n7791 gnd.n139 585
R8632 gnd.n7793 gnd.n7792 585
R8633 gnd.n7795 gnd.n137 585
R8634 gnd.n7797 gnd.n7796 585
R8635 gnd.n7798 gnd.n135 585
R8636 gnd.n7799 gnd.n131 585
R8637 gnd.n131 gnd.n128 585
R8638 gnd.n7728 gnd.n127 585
R8639 gnd.n7804 gnd.n127 585
R8640 gnd.n7727 gnd.n7726 585
R8641 gnd.n7726 gnd.n126 585
R8642 gnd.n7725 gnd.n204 585
R8643 gnd.n7725 gnd.n7724 585
R8644 gnd.n7492 gnd.n205 585
R8645 gnd.n206 gnd.n205 585
R8646 gnd.n7493 gnd.n214 585
R8647 gnd.n7716 gnd.n214 585
R8648 gnd.n7495 gnd.n7494 585
R8649 gnd.n7494 gnd.n213 585
R8650 gnd.n7496 gnd.n223 585
R8651 gnd.n7640 gnd.n223 585
R8652 gnd.n7498 gnd.n7497 585
R8653 gnd.n7497 gnd.n232 585
R8654 gnd.n7499 gnd.n230 585
R8655 gnd.n7632 gnd.n230 585
R8656 gnd.n7501 gnd.n7500 585
R8657 gnd.n7500 gnd.n229 585
R8658 gnd.n7502 gnd.n239 585
R8659 gnd.n7624 gnd.n239 585
R8660 gnd.n7504 gnd.n7503 585
R8661 gnd.n7503 gnd.n247 585
R8662 gnd.n7505 gnd.n245 585
R8663 gnd.n7616 gnd.n245 585
R8664 gnd.n7507 gnd.n7506 585
R8665 gnd.n7506 gnd.n254 585
R8666 gnd.n7508 gnd.n253 585
R8667 gnd.n7608 gnd.n253 585
R8668 gnd.n7510 gnd.n7509 585
R8669 gnd.n7509 gnd.n263 585
R8670 gnd.n7511 gnd.n261 585
R8671 gnd.n7600 gnd.n261 585
R8672 gnd.n7513 gnd.n7512 585
R8673 gnd.n7512 gnd.n260 585
R8674 gnd.n7514 gnd.n270 585
R8675 gnd.n7592 gnd.n270 585
R8676 gnd.n7516 gnd.n7515 585
R8677 gnd.n7515 gnd.n269 585
R8678 gnd.n7517 gnd.n276 585
R8679 gnd.n7584 gnd.n276 585
R8680 gnd.n7519 gnd.n7518 585
R8681 gnd.n7518 gnd.n284 585
R8682 gnd.n7520 gnd.n283 585
R8683 gnd.n7576 gnd.n283 585
R8684 gnd.n7522 gnd.n7521 585
R8685 gnd.n7521 gnd.n293 585
R8686 gnd.n7523 gnd.n291 585
R8687 gnd.n7568 gnd.n291 585
R8688 gnd.n7525 gnd.n7524 585
R8689 gnd.n7524 gnd.n290 585
R8690 gnd.n7526 gnd.n300 585
R8691 gnd.n7560 gnd.n300 585
R8692 gnd.n7528 gnd.n7527 585
R8693 gnd.n7527 gnd.n299 585
R8694 gnd.n7529 gnd.n328 585
R8695 gnd.n7536 gnd.n328 585
R8696 gnd.n7531 gnd.n7530 585
R8697 gnd.n7532 gnd.n7531 585
R8698 gnd.n336 gnd.n335 585
R8699 gnd.n335 gnd.n334 585
R8700 gnd.n7461 gnd.n7460 585
R8701 gnd.n7460 gnd.n7459 585
R8702 gnd.n339 gnd.n338 585
R8703 gnd.n340 gnd.n339 585
R8704 gnd.n7438 gnd.n343 585
R8705 gnd.n7453 gnd.n343 585
R8706 gnd.n7440 gnd.n7439 585
R8707 gnd.n7439 gnd.n315 585
R8708 gnd.n7441 gnd.n313 585
R8709 gnd.n7551 gnd.n313 585
R8710 gnd.n7443 gnd.n7442 585
R8711 gnd.n7444 gnd.n7443 585
R8712 gnd.n352 gnd.n351 585
R8713 gnd.n351 gnd.n350 585
R8714 gnd.n7431 gnd.n7430 585
R8715 gnd.n7430 gnd.n7429 585
R8716 gnd.n355 gnd.n354 585
R8717 gnd.n7408 gnd.n355 585
R8718 gnd.n7394 gnd.n7393 585
R8719 gnd.n7393 gnd.n7392 585
R8720 gnd.n7395 gnd.n368 585
R8721 gnd.n7420 gnd.n368 585
R8722 gnd.n7397 gnd.n7396 585
R8723 gnd.n7398 gnd.n7397 585
R8724 gnd.n386 gnd.n385 585
R8725 gnd.n7365 gnd.n385 585
R8726 gnd.n7386 gnd.n7385 585
R8727 gnd.n7385 gnd.n7384 585
R8728 gnd.n389 gnd.n388 585
R8729 gnd.n6143 gnd.n389 585
R8730 gnd.n6135 gnd.n400 585
R8731 gnd.n7374 gnd.n400 585
R8732 gnd.n6137 gnd.n6136 585
R8733 gnd.n6138 gnd.n6137 585
R8734 gnd.n1387 gnd.n1362 585
R8735 gnd.n6189 gnd.n1362 585
R8736 gnd.n6130 gnd.n6129 585
R8737 gnd.n6129 gnd.n1373 585
R8738 gnd.n6128 gnd.n1371 585
R8739 gnd.n6181 gnd.n1371 585
R8740 gnd.n6127 gnd.n1380 585
R8741 gnd.n6159 gnd.n1380 585
R8742 gnd.n1393 gnd.n1389 585
R8743 gnd.n1398 gnd.n1393 585
R8744 gnd.n6123 gnd.n6122 585
R8745 gnd.n6122 gnd.n6121 585
R8746 gnd.n1392 gnd.n1391 585
R8747 gnd.n1407 gnd.n1392 585
R8748 gnd.n1465 gnd.n1405 585
R8749 gnd.n6111 gnd.n1405 585
R8750 gnd.n1466 gnd.n1415 585
R8751 gnd.n6098 gnd.n1415 585
R8752 gnd.n1468 gnd.n1467 585
R8753 gnd.n1467 gnd.n1414 585
R8754 gnd.n1469 gnd.n1423 585
R8755 gnd.n6084 gnd.n1423 585
R8756 gnd.n1471 gnd.n1470 585
R8757 gnd.n1470 gnd.n1435 585
R8758 gnd.n1472 gnd.n1432 585
R8759 gnd.n6074 gnd.n1432 585
R8760 gnd.n1474 gnd.n1473 585
R8761 gnd.n6062 gnd.n1474 585
R8762 gnd.n1454 gnd.n1453 585
R8763 gnd.n1453 gnd.n1452 585
R8764 gnd.n1455 gnd.n1334 585
R8765 gnd.n6053 gnd.n1334 585
R8766 gnd.n6219 gnd.n1335 585
R8767 gnd.n6219 gnd.n6218 585
R8768 gnd.n5195 gnd.n5194 585
R8769 gnd.n5196 gnd.n5195 585
R8770 gnd.n5005 gnd.n5001 585
R8771 gnd.n5001 gnd.n1662 585
R8772 gnd.n5004 gnd.n5003 585
R8773 gnd.n5003 gnd.n1660 585
R8774 gnd.n4995 gnd.n4994 585
R8775 gnd.n5204 gnd.n4995 585
R8776 gnd.n5207 gnd.n5206 585
R8777 gnd.n5206 gnd.n5205 585
R8778 gnd.n5208 gnd.n4991 585
R8779 gnd.n4991 gnd.n4990 585
R8780 gnd.n5210 gnd.n5209 585
R8781 gnd.n5211 gnd.n5210 585
R8782 gnd.n4993 gnd.n4989 585
R8783 gnd.n4989 gnd.n1674 585
R8784 gnd.n4992 gnd.n4979 585
R8785 gnd.n5217 gnd.n4979 585
R8786 gnd.n5220 gnd.n4978 585
R8787 gnd.n5220 gnd.n5219 585
R8788 gnd.n5222 gnd.n5221 585
R8789 gnd.n5221 gnd.n1680 585
R8790 gnd.n5223 gnd.n4963 585
R8791 gnd.n4963 gnd.n4962 585
R8792 gnd.n5225 gnd.n5224 585
R8793 gnd.n5226 gnd.n5225 585
R8794 gnd.n4977 gnd.n4960 585
R8795 gnd.n4960 gnd.n1688 585
R8796 gnd.n4976 gnd.n4975 585
R8797 gnd.n4975 gnd.n1686 585
R8798 gnd.n4974 gnd.n4964 585
R8799 gnd.n4974 gnd.n4973 585
R8800 gnd.n4971 gnd.n4970 585
R8801 gnd.n4971 gnd.n1695 585
R8802 gnd.n4969 gnd.n4965 585
R8803 gnd.n4965 gnd.n1694 585
R8804 gnd.n4968 gnd.n4967 585
R8805 gnd.n4967 gnd.n1704 585
R8806 gnd.n4966 gnd.n4947 585
R8807 gnd.n4947 gnd.n1701 585
R8808 gnd.n5241 gnd.n4948 585
R8809 gnd.n5241 gnd.n5240 585
R8810 gnd.n5242 gnd.n4946 585
R8811 gnd.n5242 gnd.n1711 585
R8812 gnd.n5244 gnd.n5243 585
R8813 gnd.n5243 gnd.n1710 585
R8814 gnd.n5245 gnd.n4944 585
R8815 gnd.n4944 gnd.n4943 585
R8816 gnd.n5247 gnd.n5246 585
R8817 gnd.n5248 gnd.n5247 585
R8818 gnd.n4945 gnd.n4934 585
R8819 gnd.n4934 gnd.n1717 585
R8820 gnd.n5255 gnd.n4933 585
R8821 gnd.n5255 gnd.n5254 585
R8822 gnd.n5257 gnd.n5256 585
R8823 gnd.n5256 gnd.n1725 585
R8824 gnd.n5258 gnd.n4929 585
R8825 gnd.n4929 gnd.n1724 585
R8826 gnd.n5260 gnd.n5259 585
R8827 gnd.n5261 gnd.n5260 585
R8828 gnd.n4932 gnd.n4928 585
R8829 gnd.n4928 gnd.n1733 585
R8830 gnd.n4931 gnd.n4930 585
R8831 gnd.n4930 gnd.n1731 585
R8832 gnd.n4920 gnd.n4919 585
R8833 gnd.n5268 gnd.n4920 585
R8834 gnd.n5272 gnd.n5271 585
R8835 gnd.n5271 gnd.n5270 585
R8836 gnd.n5273 gnd.n4916 585
R8837 gnd.n4916 gnd.n1739 585
R8838 gnd.n5275 gnd.n5274 585
R8839 gnd.n5276 gnd.n5275 585
R8840 gnd.n4918 gnd.n4915 585
R8841 gnd.n4915 gnd.n1747 585
R8842 gnd.n4917 gnd.n4906 585
R8843 gnd.n4906 gnd.n1745 585
R8844 gnd.n5284 gnd.n4905 585
R8845 gnd.n5284 gnd.n5283 585
R8846 gnd.n5286 gnd.n5285 585
R8847 gnd.n5285 gnd.n1754 585
R8848 gnd.n5287 gnd.n4902 585
R8849 gnd.n4902 gnd.n1753 585
R8850 gnd.n5289 gnd.n5288 585
R8851 gnd.n5290 gnd.n5289 585
R8852 gnd.n4904 gnd.n4901 585
R8853 gnd.n4901 gnd.n1762 585
R8854 gnd.n4903 gnd.n4893 585
R8855 gnd.n4893 gnd.n1760 585
R8856 gnd.n5299 gnd.n4892 585
R8857 gnd.n5299 gnd.n5298 585
R8858 gnd.n5301 gnd.n5300 585
R8859 gnd.n5300 gnd.n1769 585
R8860 gnd.n5302 gnd.n4889 585
R8861 gnd.n4889 gnd.n1768 585
R8862 gnd.n5304 gnd.n5303 585
R8863 gnd.n5305 gnd.n5304 585
R8864 gnd.n4891 gnd.n4888 585
R8865 gnd.n4888 gnd.n1777 585
R8866 gnd.n4890 gnd.n4880 585
R8867 gnd.n4880 gnd.n1775 585
R8868 gnd.n5314 gnd.n4879 585
R8869 gnd.n5314 gnd.n5313 585
R8870 gnd.n5316 gnd.n5315 585
R8871 gnd.n5315 gnd.n1783 585
R8872 gnd.n5317 gnd.n4876 585
R8873 gnd.n4876 gnd.n4875 585
R8874 gnd.n5319 gnd.n5318 585
R8875 gnd.n5320 gnd.n5319 585
R8876 gnd.n4878 gnd.n4874 585
R8877 gnd.n4874 gnd.n1791 585
R8878 gnd.n4877 gnd.n4866 585
R8879 gnd.n4866 gnd.n1789 585
R8880 gnd.n5329 gnd.n4865 585
R8881 gnd.n5329 gnd.n5328 585
R8882 gnd.n5331 gnd.n5330 585
R8883 gnd.n5330 gnd.n1798 585
R8884 gnd.n5332 gnd.n4862 585
R8885 gnd.n4862 gnd.n1797 585
R8886 gnd.n5334 gnd.n5333 585
R8887 gnd.n5335 gnd.n5334 585
R8888 gnd.n4864 gnd.n4861 585
R8889 gnd.n4861 gnd.n1806 585
R8890 gnd.n4863 gnd.n4841 585
R8891 gnd.n4841 gnd.n1804 585
R8892 gnd.n5344 gnd.n4842 585
R8893 gnd.n5344 gnd.n5343 585
R8894 gnd.n5345 gnd.n4840 585
R8895 gnd.n5345 gnd.n1813 585
R8896 gnd.n5347 gnd.n5346 585
R8897 gnd.n5346 gnd.n1812 585
R8898 gnd.n5348 gnd.n4839 585
R8899 gnd.n4853 gnd.n4839 585
R8900 gnd.n5350 gnd.n5349 585
R8901 gnd.n5350 gnd.n1821 585
R8902 gnd.n5351 gnd.n4838 585
R8903 gnd.n5351 gnd.n1819 585
R8904 gnd.n5353 gnd.n5352 585
R8905 gnd.n5352 gnd.n1829 585
R8906 gnd.n5354 gnd.n4835 585
R8907 gnd.n4835 gnd.n1827 585
R8908 gnd.n5356 gnd.n5355 585
R8909 gnd.n5357 gnd.n5356 585
R8910 gnd.n4837 gnd.n4834 585
R8911 gnd.n4834 gnd.n1836 585
R8912 gnd.n4836 gnd.n4823 585
R8913 gnd.n5363 gnd.n4823 585
R8914 gnd.n5365 gnd.n4822 585
R8915 gnd.n5365 gnd.n5364 585
R8916 gnd.n5367 gnd.n5366 585
R8917 gnd.n5366 gnd.n1843 585
R8918 gnd.n5368 gnd.n4818 585
R8919 gnd.n4818 gnd.n1842 585
R8920 gnd.n5370 gnd.n5369 585
R8921 gnd.n5371 gnd.n5370 585
R8922 gnd.n4821 gnd.n4817 585
R8923 gnd.n4817 gnd.n1851 585
R8924 gnd.n4820 gnd.n4819 585
R8925 gnd.n4819 gnd.n1849 585
R8926 gnd.n4810 gnd.n4809 585
R8927 gnd.n5378 gnd.n4810 585
R8928 gnd.n5382 gnd.n5381 585
R8929 gnd.n5381 gnd.n5380 585
R8930 gnd.n5383 gnd.n4806 585
R8931 gnd.n4806 gnd.n1857 585
R8932 gnd.n5385 gnd.n5384 585
R8933 gnd.n5386 gnd.n5385 585
R8934 gnd.n4808 gnd.n4805 585
R8935 gnd.n4805 gnd.n1864 585
R8936 gnd.n4807 gnd.n4794 585
R8937 gnd.n5392 gnd.n4794 585
R8938 gnd.n5394 gnd.n4793 585
R8939 gnd.n5394 gnd.n5393 585
R8940 gnd.n5396 gnd.n5395 585
R8941 gnd.n5395 gnd.n1871 585
R8942 gnd.n5397 gnd.n4789 585
R8943 gnd.n4789 gnd.n1870 585
R8944 gnd.n5399 gnd.n5398 585
R8945 gnd.n5400 gnd.n5399 585
R8946 gnd.n4792 gnd.n4788 585
R8947 gnd.n4788 gnd.n1879 585
R8948 gnd.n4791 gnd.n4790 585
R8949 gnd.n4790 gnd.n1877 585
R8950 gnd.n4780 gnd.n4779 585
R8951 gnd.n5407 gnd.n4780 585
R8952 gnd.n5411 gnd.n5410 585
R8953 gnd.n5410 gnd.n5409 585
R8954 gnd.n5412 gnd.n4775 585
R8955 gnd.n4775 gnd.n1885 585
R8956 gnd.n5414 gnd.n5413 585
R8957 gnd.n5415 gnd.n5414 585
R8958 gnd.n4778 gnd.n4774 585
R8959 gnd.n4774 gnd.n1893 585
R8960 gnd.n4777 gnd.n4776 585
R8961 gnd.n4776 gnd.n1891 585
R8962 gnd.n4766 gnd.n4765 585
R8963 gnd.n5423 gnd.n4766 585
R8964 gnd.n5426 gnd.n5425 585
R8965 gnd.n5425 gnd.n5424 585
R8966 gnd.n5427 gnd.n4762 585
R8967 gnd.n4762 gnd.n1899 585
R8968 gnd.n5429 gnd.n5428 585
R8969 gnd.n5430 gnd.n5429 585
R8970 gnd.n4764 gnd.n4761 585
R8971 gnd.n4761 gnd.n1907 585
R8972 gnd.n4763 gnd.n4753 585
R8973 gnd.n4753 gnd.n1905 585
R8974 gnd.n5439 gnd.n4752 585
R8975 gnd.n5439 gnd.n5438 585
R8976 gnd.n5441 gnd.n5440 585
R8977 gnd.n5440 gnd.n1914 585
R8978 gnd.n5442 gnd.n4750 585
R8979 gnd.n4750 gnd.n1913 585
R8980 gnd.n5444 gnd.n5443 585
R8981 gnd.n5445 gnd.n5444 585
R8982 gnd.n4751 gnd.n4749 585
R8983 gnd.n4749 gnd.n1922 585
R8984 gnd.n4677 gnd.n4676 585
R8985 gnd.n4677 gnd.n1920 585
R8986 gnd.n5455 gnd.n5454 585
R8987 gnd.n5454 gnd.n5453 585
R8988 gnd.n5456 gnd.n4655 585
R8989 gnd.n4655 gnd.n1928 585
R8990 gnd.n5521 gnd.n5520 585
R8991 gnd.n5519 gnd.n4654 585
R8992 gnd.n5518 gnd.n4653 585
R8993 gnd.n5523 gnd.n4653 585
R8994 gnd.n5517 gnd.n5516 585
R8995 gnd.n5515 gnd.n5514 585
R8996 gnd.n5513 gnd.n5512 585
R8997 gnd.n5511 gnd.n5510 585
R8998 gnd.n5509 gnd.n5508 585
R8999 gnd.n5507 gnd.n5506 585
R9000 gnd.n5505 gnd.n5504 585
R9001 gnd.n5503 gnd.n5502 585
R9002 gnd.n5501 gnd.n5500 585
R9003 gnd.n5499 gnd.n5498 585
R9004 gnd.n5497 gnd.n5496 585
R9005 gnd.n5495 gnd.n5494 585
R9006 gnd.n5493 gnd.n5492 585
R9007 gnd.n5491 gnd.n5490 585
R9008 gnd.n5489 gnd.n5488 585
R9009 gnd.n5487 gnd.n5486 585
R9010 gnd.n5485 gnd.n5484 585
R9011 gnd.n5483 gnd.n5482 585
R9012 gnd.n5481 gnd.n5480 585
R9013 gnd.n5479 gnd.n5478 585
R9014 gnd.n5477 gnd.n5476 585
R9015 gnd.n5475 gnd.n5474 585
R9016 gnd.n5473 gnd.n5472 585
R9017 gnd.n5471 gnd.n5470 585
R9018 gnd.n5469 gnd.n5468 585
R9019 gnd.n5467 gnd.n5466 585
R9020 gnd.n5465 gnd.n5464 585
R9021 gnd.n5463 gnd.n5462 585
R9022 gnd.n5461 gnd.n4618 585
R9023 gnd.n5526 gnd.n5525 585
R9024 gnd.n4620 gnd.n4617 585
R9025 gnd.n4683 gnd.n4682 585
R9026 gnd.n4685 gnd.n4684 585
R9027 gnd.n4688 gnd.n4687 585
R9028 gnd.n4690 gnd.n4689 585
R9029 gnd.n4692 gnd.n4691 585
R9030 gnd.n4694 gnd.n4693 585
R9031 gnd.n4696 gnd.n4695 585
R9032 gnd.n4698 gnd.n4697 585
R9033 gnd.n4700 gnd.n4699 585
R9034 gnd.n4702 gnd.n4701 585
R9035 gnd.n4704 gnd.n4703 585
R9036 gnd.n4706 gnd.n4705 585
R9037 gnd.n4708 gnd.n4707 585
R9038 gnd.n4710 gnd.n4709 585
R9039 gnd.n4712 gnd.n4711 585
R9040 gnd.n4714 gnd.n4713 585
R9041 gnd.n4716 gnd.n4715 585
R9042 gnd.n4718 gnd.n4717 585
R9043 gnd.n4720 gnd.n4719 585
R9044 gnd.n4722 gnd.n4721 585
R9045 gnd.n4724 gnd.n4723 585
R9046 gnd.n4726 gnd.n4725 585
R9047 gnd.n4728 gnd.n4727 585
R9048 gnd.n4730 gnd.n4729 585
R9049 gnd.n4732 gnd.n4731 585
R9050 gnd.n4734 gnd.n4733 585
R9051 gnd.n4736 gnd.n4735 585
R9052 gnd.n4738 gnd.n4737 585
R9053 gnd.n4740 gnd.n4739 585
R9054 gnd.n4742 gnd.n4741 585
R9055 gnd.n4744 gnd.n4743 585
R9056 gnd.n5076 gnd.n5000 585
R9057 gnd.n5077 gnd.n5075 585
R9058 gnd.n5079 gnd.n5078 585
R9059 gnd.n5081 gnd.n5072 585
R9060 gnd.n5083 gnd.n5082 585
R9061 gnd.n5084 gnd.n5071 585
R9062 gnd.n5086 gnd.n5085 585
R9063 gnd.n5088 gnd.n5069 585
R9064 gnd.n5090 gnd.n5089 585
R9065 gnd.n5091 gnd.n5068 585
R9066 gnd.n5093 gnd.n5092 585
R9067 gnd.n5095 gnd.n5066 585
R9068 gnd.n5097 gnd.n5096 585
R9069 gnd.n5098 gnd.n5065 585
R9070 gnd.n5100 gnd.n5099 585
R9071 gnd.n5102 gnd.n5063 585
R9072 gnd.n5104 gnd.n5103 585
R9073 gnd.n5105 gnd.n5062 585
R9074 gnd.n5107 gnd.n5106 585
R9075 gnd.n5109 gnd.n5060 585
R9076 gnd.n5111 gnd.n5110 585
R9077 gnd.n5112 gnd.n5059 585
R9078 gnd.n5114 gnd.n5113 585
R9079 gnd.n5116 gnd.n5057 585
R9080 gnd.n5118 gnd.n5117 585
R9081 gnd.n5119 gnd.n5056 585
R9082 gnd.n5121 gnd.n5120 585
R9083 gnd.n5123 gnd.n5054 585
R9084 gnd.n5125 gnd.n5124 585
R9085 gnd.n5127 gnd.n5051 585
R9086 gnd.n5129 gnd.n5128 585
R9087 gnd.n5131 gnd.n5050 585
R9088 gnd.n5132 gnd.n1654 585
R9089 gnd.n5135 gnd.n1305 585
R9090 gnd.n5137 gnd.n5136 585
R9091 gnd.n5139 gnd.n5048 585
R9092 gnd.n5141 gnd.n5140 585
R9093 gnd.n5143 gnd.n5045 585
R9094 gnd.n5145 gnd.n5144 585
R9095 gnd.n5147 gnd.n5043 585
R9096 gnd.n5149 gnd.n5148 585
R9097 gnd.n5150 gnd.n5042 585
R9098 gnd.n5152 gnd.n5151 585
R9099 gnd.n5154 gnd.n5040 585
R9100 gnd.n5156 gnd.n5155 585
R9101 gnd.n5157 gnd.n5039 585
R9102 gnd.n5159 gnd.n5158 585
R9103 gnd.n5161 gnd.n5037 585
R9104 gnd.n5163 gnd.n5162 585
R9105 gnd.n5164 gnd.n5036 585
R9106 gnd.n5166 gnd.n5165 585
R9107 gnd.n5168 gnd.n5034 585
R9108 gnd.n5170 gnd.n5169 585
R9109 gnd.n5171 gnd.n5033 585
R9110 gnd.n5173 gnd.n5172 585
R9111 gnd.n5175 gnd.n5031 585
R9112 gnd.n5177 gnd.n5176 585
R9113 gnd.n5178 gnd.n5030 585
R9114 gnd.n5180 gnd.n5179 585
R9115 gnd.n5182 gnd.n5028 585
R9116 gnd.n5184 gnd.n5183 585
R9117 gnd.n5185 gnd.n5027 585
R9118 gnd.n5187 gnd.n5186 585
R9119 gnd.n5189 gnd.n5025 585
R9120 gnd.n5191 gnd.n5190 585
R9121 gnd.n5192 gnd.n5002 585
R9122 gnd.n5197 gnd.n4999 585
R9123 gnd.n5197 gnd.n5196 585
R9124 gnd.n5199 gnd.n5198 585
R9125 gnd.n5198 gnd.n1662 585
R9126 gnd.n5200 gnd.n4997 585
R9127 gnd.n4997 gnd.n1660 585
R9128 gnd.n5202 gnd.n5201 585
R9129 gnd.n5204 gnd.n5202 585
R9130 gnd.n4998 gnd.n4996 585
R9131 gnd.n5205 gnd.n4996 585
R9132 gnd.n4987 gnd.n4986 585
R9133 gnd.n4990 gnd.n4987 585
R9134 gnd.n5213 gnd.n5212 585
R9135 gnd.n5212 gnd.n5211 585
R9136 gnd.n5214 gnd.n4981 585
R9137 gnd.n4981 gnd.n1674 585
R9138 gnd.n5216 gnd.n5215 585
R9139 gnd.n5217 gnd.n5216 585
R9140 gnd.n4985 gnd.n4980 585
R9141 gnd.n5219 gnd.n4980 585
R9142 gnd.n4984 gnd.n4983 585
R9143 gnd.n4983 gnd.n1680 585
R9144 gnd.n4982 gnd.n4958 585
R9145 gnd.n4962 gnd.n4958 585
R9146 gnd.n5227 gnd.n4959 585
R9147 gnd.n5227 gnd.n5226 585
R9148 gnd.n5228 gnd.n4957 585
R9149 gnd.n5228 gnd.n1688 585
R9150 gnd.n5230 gnd.n5229 585
R9151 gnd.n5229 gnd.n1686 585
R9152 gnd.n5231 gnd.n4956 585
R9153 gnd.n4973 gnd.n4956 585
R9154 gnd.n5233 gnd.n5232 585
R9155 gnd.n5233 gnd.n1695 585
R9156 gnd.n5234 gnd.n4955 585
R9157 gnd.n5234 gnd.n1694 585
R9158 gnd.n5236 gnd.n5235 585
R9159 gnd.n5235 gnd.n1704 585
R9160 gnd.n5237 gnd.n4951 585
R9161 gnd.n4951 gnd.n1701 585
R9162 gnd.n5239 gnd.n5238 585
R9163 gnd.n5240 gnd.n5239 585
R9164 gnd.n4954 gnd.n4950 585
R9165 gnd.n4950 gnd.n1711 585
R9166 gnd.n4953 gnd.n4952 585
R9167 gnd.n4952 gnd.n1710 585
R9168 gnd.n4941 gnd.n4940 585
R9169 gnd.n4943 gnd.n4941 585
R9170 gnd.n5250 gnd.n5249 585
R9171 gnd.n5249 gnd.n5248 585
R9172 gnd.n5251 gnd.n4937 585
R9173 gnd.n4937 gnd.n1717 585
R9174 gnd.n5253 gnd.n5252 585
R9175 gnd.n5254 gnd.n5253 585
R9176 gnd.n4939 gnd.n4936 585
R9177 gnd.n4936 gnd.n1725 585
R9178 gnd.n4938 gnd.n4926 585
R9179 gnd.n4926 gnd.n1724 585
R9180 gnd.n5262 gnd.n4925 585
R9181 gnd.n5262 gnd.n5261 585
R9182 gnd.n5264 gnd.n5263 585
R9183 gnd.n5263 gnd.n1733 585
R9184 gnd.n5265 gnd.n4922 585
R9185 gnd.n4922 gnd.n1731 585
R9186 gnd.n5267 gnd.n5266 585
R9187 gnd.n5268 gnd.n5267 585
R9188 gnd.n4924 gnd.n4921 585
R9189 gnd.n5270 gnd.n4921 585
R9190 gnd.n4923 gnd.n4913 585
R9191 gnd.n4913 gnd.n1739 585
R9192 gnd.n5277 gnd.n4912 585
R9193 gnd.n5277 gnd.n5276 585
R9194 gnd.n5279 gnd.n5278 585
R9195 gnd.n5278 gnd.n1747 585
R9196 gnd.n5280 gnd.n4909 585
R9197 gnd.n4909 gnd.n1745 585
R9198 gnd.n5282 gnd.n5281 585
R9199 gnd.n5283 gnd.n5282 585
R9200 gnd.n4911 gnd.n4908 585
R9201 gnd.n4908 gnd.n1754 585
R9202 gnd.n4910 gnd.n4899 585
R9203 gnd.n4899 gnd.n1753 585
R9204 gnd.n5291 gnd.n4898 585
R9205 gnd.n5291 gnd.n5290 585
R9206 gnd.n5293 gnd.n5292 585
R9207 gnd.n5292 gnd.n1762 585
R9208 gnd.n5294 gnd.n4895 585
R9209 gnd.n4895 gnd.n1760 585
R9210 gnd.n5296 gnd.n5295 585
R9211 gnd.n5298 gnd.n5296 585
R9212 gnd.n4897 gnd.n4894 585
R9213 gnd.n4894 gnd.n1769 585
R9214 gnd.n4896 gnd.n4886 585
R9215 gnd.n4886 gnd.n1768 585
R9216 gnd.n5306 gnd.n4885 585
R9217 gnd.n5306 gnd.n5305 585
R9218 gnd.n5308 gnd.n5307 585
R9219 gnd.n5307 gnd.n1777 585
R9220 gnd.n5309 gnd.n4882 585
R9221 gnd.n4882 gnd.n1775 585
R9222 gnd.n5311 gnd.n5310 585
R9223 gnd.n5313 gnd.n5311 585
R9224 gnd.n4884 gnd.n4881 585
R9225 gnd.n4881 gnd.n1783 585
R9226 gnd.n4883 gnd.n4872 585
R9227 gnd.n4875 gnd.n4872 585
R9228 gnd.n5321 gnd.n4871 585
R9229 gnd.n5321 gnd.n5320 585
R9230 gnd.n5323 gnd.n5322 585
R9231 gnd.n5322 gnd.n1791 585
R9232 gnd.n5324 gnd.n4868 585
R9233 gnd.n4868 gnd.n1789 585
R9234 gnd.n5326 gnd.n5325 585
R9235 gnd.n5328 gnd.n5326 585
R9236 gnd.n4870 gnd.n4867 585
R9237 gnd.n4867 gnd.n1798 585
R9238 gnd.n4869 gnd.n4859 585
R9239 gnd.n4859 gnd.n1797 585
R9240 gnd.n5336 gnd.n4858 585
R9241 gnd.n5336 gnd.n5335 585
R9242 gnd.n5338 gnd.n5337 585
R9243 gnd.n5337 gnd.n1806 585
R9244 gnd.n5339 gnd.n4844 585
R9245 gnd.n4844 gnd.n1804 585
R9246 gnd.n5341 gnd.n5340 585
R9247 gnd.n5343 gnd.n5341 585
R9248 gnd.n4857 gnd.n4843 585
R9249 gnd.n4843 gnd.n1813 585
R9250 gnd.n4856 gnd.n4855 585
R9251 gnd.n4855 gnd.n1812 585
R9252 gnd.n4854 gnd.n4845 585
R9253 gnd.n4854 gnd.n4853 585
R9254 gnd.n4851 gnd.n4850 585
R9255 gnd.n4851 gnd.n1821 585
R9256 gnd.n4849 gnd.n4846 585
R9257 gnd.n4846 gnd.n1819 585
R9258 gnd.n4848 gnd.n4847 585
R9259 gnd.n4847 gnd.n1829 585
R9260 gnd.n4832 gnd.n4831 585
R9261 gnd.n4832 gnd.n1827 585
R9262 gnd.n5359 gnd.n5358 585
R9263 gnd.n5358 gnd.n5357 585
R9264 gnd.n5360 gnd.n4826 585
R9265 gnd.n4826 gnd.n1836 585
R9266 gnd.n5362 gnd.n5361 585
R9267 gnd.n5363 gnd.n5362 585
R9268 gnd.n4830 gnd.n4825 585
R9269 gnd.n5364 gnd.n4825 585
R9270 gnd.n4829 gnd.n4828 585
R9271 gnd.n4828 gnd.n1843 585
R9272 gnd.n4827 gnd.n4815 585
R9273 gnd.n4815 gnd.n1842 585
R9274 gnd.n5372 gnd.n4814 585
R9275 gnd.n5372 gnd.n5371 585
R9276 gnd.n5374 gnd.n5373 585
R9277 gnd.n5373 gnd.n1851 585
R9278 gnd.n5375 gnd.n4812 585
R9279 gnd.n4812 gnd.n1849 585
R9280 gnd.n5377 gnd.n5376 585
R9281 gnd.n5378 gnd.n5377 585
R9282 gnd.n4813 gnd.n4811 585
R9283 gnd.n5380 gnd.n4811 585
R9284 gnd.n4803 gnd.n4802 585
R9285 gnd.n4803 gnd.n1857 585
R9286 gnd.n5388 gnd.n5387 585
R9287 gnd.n5387 gnd.n5386 585
R9288 gnd.n5389 gnd.n4797 585
R9289 gnd.n4797 gnd.n1864 585
R9290 gnd.n5391 gnd.n5390 585
R9291 gnd.n5392 gnd.n5391 585
R9292 gnd.n4801 gnd.n4796 585
R9293 gnd.n5393 gnd.n4796 585
R9294 gnd.n4800 gnd.n4799 585
R9295 gnd.n4799 gnd.n1871 585
R9296 gnd.n4798 gnd.n4786 585
R9297 gnd.n4786 gnd.n1870 585
R9298 gnd.n5401 gnd.n4785 585
R9299 gnd.n5401 gnd.n5400 585
R9300 gnd.n5403 gnd.n5402 585
R9301 gnd.n5402 gnd.n1879 585
R9302 gnd.n5404 gnd.n4782 585
R9303 gnd.n4782 gnd.n1877 585
R9304 gnd.n5406 gnd.n5405 585
R9305 gnd.n5407 gnd.n5406 585
R9306 gnd.n4784 gnd.n4781 585
R9307 gnd.n5409 gnd.n4781 585
R9308 gnd.n4783 gnd.n4772 585
R9309 gnd.n4772 gnd.n1885 585
R9310 gnd.n5416 gnd.n4771 585
R9311 gnd.n5416 gnd.n5415 585
R9312 gnd.n5418 gnd.n5417 585
R9313 gnd.n5417 gnd.n1893 585
R9314 gnd.n5419 gnd.n4768 585
R9315 gnd.n4768 gnd.n1891 585
R9316 gnd.n5421 gnd.n5420 585
R9317 gnd.n5423 gnd.n5421 585
R9318 gnd.n4770 gnd.n4767 585
R9319 gnd.n5424 gnd.n4767 585
R9320 gnd.n4769 gnd.n4759 585
R9321 gnd.n4759 gnd.n1899 585
R9322 gnd.n5431 gnd.n4758 585
R9323 gnd.n5431 gnd.n5430 585
R9324 gnd.n5433 gnd.n5432 585
R9325 gnd.n5432 gnd.n1907 585
R9326 gnd.n5434 gnd.n4755 585
R9327 gnd.n4755 gnd.n1905 585
R9328 gnd.n5436 gnd.n5435 585
R9329 gnd.n5438 gnd.n5436 585
R9330 gnd.n4757 gnd.n4754 585
R9331 gnd.n4754 gnd.n1914 585
R9332 gnd.n4756 gnd.n4747 585
R9333 gnd.n4747 gnd.n1913 585
R9334 gnd.n5446 gnd.n4746 585
R9335 gnd.n5446 gnd.n5445 585
R9336 gnd.n5448 gnd.n5447 585
R9337 gnd.n5447 gnd.n1922 585
R9338 gnd.n5449 gnd.n4679 585
R9339 gnd.n4679 gnd.n1920 585
R9340 gnd.n5451 gnd.n5450 585
R9341 gnd.n5453 gnd.n5451 585
R9342 gnd.n4745 gnd.n4678 585
R9343 gnd.n4678 gnd.n1928 585
R9344 gnd.n6548 gnd.n963 585
R9345 gnd.n2192 gnd.n963 585
R9346 gnd.n7352 gnd.n7351 585
R9347 gnd.n7352 gnd.n312 585
R9348 gnd.n7354 gnd.n7353 585
R9349 gnd.n7353 gnd.n358 585
R9350 gnd.n7355 gnd.n416 585
R9351 gnd.n416 gnd.n356 585
R9352 gnd.n7357 gnd.n7356 585
R9353 gnd.n7357 gnd.n377 585
R9354 gnd.n7358 gnd.n415 585
R9355 gnd.n7358 gnd.n370 585
R9356 gnd.n7360 gnd.n7359 585
R9357 gnd.n7359 gnd.n367 585
R9358 gnd.n7361 gnd.n410 585
R9359 gnd.n410 gnd.n384 585
R9360 gnd.n7363 gnd.n7362 585
R9361 gnd.n7364 gnd.n7363 585
R9362 gnd.n411 gnd.n409 585
R9363 gnd.n409 gnd.n390 585
R9364 gnd.n6173 gnd.n6172 585
R9365 gnd.n6173 gnd.n402 585
R9366 gnd.n6174 gnd.n6168 585
R9367 gnd.n6174 gnd.n399 585
R9368 gnd.n6176 gnd.n6175 585
R9369 gnd.n6175 gnd.n1364 585
R9370 gnd.n6177 gnd.n1375 585
R9371 gnd.n1375 gnd.n1361 585
R9372 gnd.n6179 gnd.n6178 585
R9373 gnd.n6180 gnd.n6179 585
R9374 gnd.n1376 gnd.n1374 585
R9375 gnd.n1374 gnd.n1370 585
R9376 gnd.n6162 gnd.n6161 585
R9377 gnd.n6161 gnd.n6160 585
R9378 gnd.n1379 gnd.n1378 585
R9379 gnd.n1396 gnd.n1379 585
R9380 gnd.n6106 gnd.n1409 585
R9381 gnd.n1409 gnd.n1394 585
R9382 gnd.n6108 gnd.n6107 585
R9383 gnd.n6109 gnd.n6108 585
R9384 gnd.n1410 gnd.n1408 585
R9385 gnd.n1408 gnd.n1404 585
R9386 gnd.n6101 gnd.n6100 585
R9387 gnd.n6100 gnd.n6099 585
R9388 gnd.n1413 gnd.n1412 585
R9389 gnd.n1424 gnd.n1413 585
R9390 gnd.n6070 gnd.n1437 585
R9391 gnd.n1437 gnd.n1422 585
R9392 gnd.n6072 gnd.n6071 585
R9393 gnd.n6073 gnd.n6072 585
R9394 gnd.n1438 gnd.n1436 585
R9395 gnd.n1436 gnd.n1431 585
R9396 gnd.n6065 gnd.n6064 585
R9397 gnd.n6064 gnd.n6063 585
R9398 gnd.n1451 gnd.n1440 585
R9399 gnd.n6044 gnd.n1451 585
R9400 gnd.n1450 gnd.n1449 585
R9401 gnd.n1450 gnd.n1338 585
R9402 gnd.n1442 gnd.n1441 585
R9403 gnd.n1441 gnd.n1336 585
R9404 gnd.n1445 gnd.n1444 585
R9405 gnd.n1444 gnd.n1285 585
R9406 gnd.n1255 gnd.n1254 585
R9407 gnd.n6295 gnd.n1255 585
R9408 gnd.n6298 gnd.n6297 585
R9409 gnd.n6297 gnd.n6296 585
R9410 gnd.n6299 gnd.n1249 585
R9411 gnd.n1256 gnd.n1249 585
R9412 gnd.n6301 gnd.n6300 585
R9413 gnd.n6302 gnd.n6301 585
R9414 gnd.n1250 gnd.n1246 585
R9415 gnd.n6303 gnd.n1246 585
R9416 gnd.n6009 gnd.n1621 585
R9417 gnd.n1621 gnd.n1245 585
R9418 gnd.n6011 gnd.n6010 585
R9419 gnd.n6012 gnd.n6011 585
R9420 gnd.n1622 gnd.n1620 585
R9421 gnd.n1620 gnd.n1618 585
R9422 gnd.n6003 gnd.n6002 585
R9423 gnd.n6002 gnd.n6001 585
R9424 gnd.n1625 gnd.n1624 585
R9425 gnd.n1626 gnd.n1625 585
R9426 gnd.n5990 gnd.n5989 585
R9427 gnd.n5991 gnd.n5990 585
R9428 gnd.n1635 gnd.n1634 585
R9429 gnd.n1640 gnd.n1634 585
R9430 gnd.n5985 gnd.n5984 585
R9431 gnd.n5984 gnd.n5983 585
R9432 gnd.n1638 gnd.n1637 585
R9433 gnd.n1639 gnd.n1638 585
R9434 gnd.n5974 gnd.n5973 585
R9435 gnd.n5975 gnd.n5974 585
R9436 gnd.n1649 gnd.n1648 585
R9437 gnd.n1648 gnd.n1646 585
R9438 gnd.n5969 gnd.n5968 585
R9439 gnd.n5968 gnd.n5967 585
R9440 gnd.n1652 gnd.n1651 585
R9441 gnd.n1653 gnd.n1652 585
R9442 gnd.n5958 gnd.n5957 585
R9443 gnd.n5959 gnd.n5958 585
R9444 gnd.n1664 gnd.n1663 585
R9445 gnd.n5203 gnd.n1663 585
R9446 gnd.n5953 gnd.n5952 585
R9447 gnd.n5952 gnd.n5951 585
R9448 gnd.n1667 gnd.n1666 585
R9449 gnd.n4988 gnd.n1667 585
R9450 gnd.n5942 gnd.n5941 585
R9451 gnd.n5943 gnd.n5942 585
R9452 gnd.n1676 gnd.n1675 585
R9453 gnd.n5218 gnd.n1675 585
R9454 gnd.n5937 gnd.n5936 585
R9455 gnd.n5936 gnd.n5935 585
R9456 gnd.n1679 gnd.n1678 585
R9457 gnd.n4961 gnd.n1679 585
R9458 gnd.n5926 gnd.n5925 585
R9459 gnd.n5927 gnd.n5926 585
R9460 gnd.n1690 gnd.n1689 585
R9461 gnd.n4972 gnd.n1689 585
R9462 gnd.n5921 gnd.n5920 585
R9463 gnd.n5920 gnd.n5919 585
R9464 gnd.n1693 gnd.n1692 585
R9465 gnd.n1703 gnd.n1693 585
R9466 gnd.n5910 gnd.n5909 585
R9467 gnd.n5911 gnd.n5910 585
R9468 gnd.n1706 gnd.n1705 585
R9469 gnd.n4949 gnd.n1705 585
R9470 gnd.n5905 gnd.n5904 585
R9471 gnd.n5904 gnd.n5903 585
R9472 gnd.n1709 gnd.n1708 585
R9473 gnd.n4942 gnd.n1709 585
R9474 gnd.n5894 gnd.n5893 585
R9475 gnd.n5895 gnd.n5894 585
R9476 gnd.n1720 gnd.n1719 585
R9477 gnd.n4935 gnd.n1719 585
R9478 gnd.n5889 gnd.n5888 585
R9479 gnd.n5888 gnd.n5887 585
R9480 gnd.n1723 gnd.n1722 585
R9481 gnd.n4927 gnd.n1723 585
R9482 gnd.n5878 gnd.n5877 585
R9483 gnd.n5879 gnd.n5878 585
R9484 gnd.n1735 gnd.n1734 585
R9485 gnd.n5269 gnd.n1734 585
R9486 gnd.n5873 gnd.n5872 585
R9487 gnd.n5872 gnd.n5871 585
R9488 gnd.n1738 gnd.n1737 585
R9489 gnd.n4914 gnd.n1738 585
R9490 gnd.n5862 gnd.n5861 585
R9491 gnd.n5863 gnd.n5862 585
R9492 gnd.n1749 gnd.n1748 585
R9493 gnd.n4907 gnd.n1748 585
R9494 gnd.n5857 gnd.n5856 585
R9495 gnd.n5856 gnd.n5855 585
R9496 gnd.n1752 gnd.n1751 585
R9497 gnd.n4900 gnd.n1752 585
R9498 gnd.n5846 gnd.n5845 585
R9499 gnd.n5847 gnd.n5846 585
R9500 gnd.n1764 gnd.n1763 585
R9501 gnd.n5297 gnd.n1763 585
R9502 gnd.n5841 gnd.n5840 585
R9503 gnd.n5840 gnd.n5839 585
R9504 gnd.n1767 gnd.n1766 585
R9505 gnd.n4887 gnd.n1767 585
R9506 gnd.n5830 gnd.n5829 585
R9507 gnd.n5831 gnd.n5830 585
R9508 gnd.n1779 gnd.n1778 585
R9509 gnd.n5312 gnd.n1778 585
R9510 gnd.n5825 gnd.n5824 585
R9511 gnd.n5824 gnd.n5823 585
R9512 gnd.n1782 gnd.n1781 585
R9513 gnd.n4873 gnd.n1782 585
R9514 gnd.n5814 gnd.n5813 585
R9515 gnd.n5815 gnd.n5814 585
R9516 gnd.n1793 gnd.n1792 585
R9517 gnd.n5327 gnd.n1792 585
R9518 gnd.n5809 gnd.n5808 585
R9519 gnd.n5808 gnd.n5807 585
R9520 gnd.n1796 gnd.n1795 585
R9521 gnd.n4860 gnd.n1796 585
R9522 gnd.n5798 gnd.n5797 585
R9523 gnd.n5799 gnd.n5798 585
R9524 gnd.n1808 gnd.n1807 585
R9525 gnd.n5342 gnd.n1807 585
R9526 gnd.n5793 gnd.n5792 585
R9527 gnd.n5792 gnd.n5791 585
R9528 gnd.n1811 gnd.n1810 585
R9529 gnd.n4852 gnd.n1811 585
R9530 gnd.n5782 gnd.n5781 585
R9531 gnd.n5783 gnd.n5782 585
R9532 gnd.n1823 gnd.n1822 585
R9533 gnd.n1828 gnd.n1822 585
R9534 gnd.n5777 gnd.n5776 585
R9535 gnd.n5776 gnd.n5775 585
R9536 gnd.n1826 gnd.n1825 585
R9537 gnd.n4833 gnd.n1826 585
R9538 gnd.n5766 gnd.n5765 585
R9539 gnd.n5767 gnd.n5766 585
R9540 gnd.n1838 gnd.n1837 585
R9541 gnd.n4824 gnd.n1837 585
R9542 gnd.n5761 gnd.n5760 585
R9543 gnd.n5760 gnd.n5759 585
R9544 gnd.n1841 gnd.n1840 585
R9545 gnd.n4816 gnd.n1841 585
R9546 gnd.n5750 gnd.n5749 585
R9547 gnd.n5751 gnd.n5750 585
R9548 gnd.n1853 gnd.n1852 585
R9549 gnd.n5379 gnd.n1852 585
R9550 gnd.n5745 gnd.n5744 585
R9551 gnd.n5744 gnd.n5743 585
R9552 gnd.n1856 gnd.n1855 585
R9553 gnd.n4804 gnd.n1856 585
R9554 gnd.n5734 gnd.n5733 585
R9555 gnd.n5735 gnd.n5734 585
R9556 gnd.n1866 gnd.n1865 585
R9557 gnd.n4795 gnd.n1865 585
R9558 gnd.n5729 gnd.n5728 585
R9559 gnd.n5728 gnd.n5727 585
R9560 gnd.n1869 gnd.n1868 585
R9561 gnd.n4787 gnd.n1869 585
R9562 gnd.n5718 gnd.n5717 585
R9563 gnd.n5719 gnd.n5718 585
R9564 gnd.n1881 gnd.n1880 585
R9565 gnd.n5408 gnd.n1880 585
R9566 gnd.n5713 gnd.n5712 585
R9567 gnd.n5712 gnd.n5711 585
R9568 gnd.n1884 gnd.n1883 585
R9569 gnd.n4773 gnd.n1884 585
R9570 gnd.n5702 gnd.n5701 585
R9571 gnd.n5703 gnd.n5702 585
R9572 gnd.n1895 gnd.n1894 585
R9573 gnd.n5422 gnd.n1894 585
R9574 gnd.n5697 gnd.n5696 585
R9575 gnd.n5696 gnd.n5695 585
R9576 gnd.n1898 gnd.n1897 585
R9577 gnd.n4760 gnd.n1898 585
R9578 gnd.n5686 gnd.n5685 585
R9579 gnd.n5687 gnd.n5686 585
R9580 gnd.n1909 gnd.n1908 585
R9581 gnd.n5437 gnd.n1908 585
R9582 gnd.n5681 gnd.n5680 585
R9583 gnd.n5680 gnd.n5679 585
R9584 gnd.n1912 gnd.n1911 585
R9585 gnd.n4748 gnd.n1912 585
R9586 gnd.n5670 gnd.n5669 585
R9587 gnd.n5671 gnd.n5670 585
R9588 gnd.n1924 gnd.n1923 585
R9589 gnd.n5452 gnd.n1923 585
R9590 gnd.n5665 gnd.n5664 585
R9591 gnd.n5664 gnd.n5663 585
R9592 gnd.n1927 gnd.n1926 585
R9593 gnd.n4652 gnd.n1927 585
R9594 gnd.n5654 gnd.n5653 585
R9595 gnd.n5655 gnd.n5654 585
R9596 gnd.n1937 gnd.n1936 585
R9597 gnd.n1936 gnd.n1934 585
R9598 gnd.n5649 gnd.n5648 585
R9599 gnd.n5648 gnd.n5647 585
R9600 gnd.n1940 gnd.n1939 585
R9601 gnd.n1941 gnd.n1940 585
R9602 gnd.n5638 gnd.n5637 585
R9603 gnd.n5639 gnd.n5638 585
R9604 gnd.n1949 gnd.n1948 585
R9605 gnd.n1954 gnd.n1948 585
R9606 gnd.n5633 gnd.n5632 585
R9607 gnd.n5632 gnd.n5631 585
R9608 gnd.n1952 gnd.n1951 585
R9609 gnd.n1953 gnd.n1952 585
R9610 gnd.n5622 gnd.n5621 585
R9611 gnd.n5623 gnd.n5622 585
R9612 gnd.n1963 gnd.n1962 585
R9613 gnd.n1962 gnd.n1960 585
R9614 gnd.n5617 gnd.n5616 585
R9615 gnd.n5616 gnd.n5615 585
R9616 gnd.n1966 gnd.n1965 585
R9617 gnd.n1967 gnd.n1966 585
R9618 gnd.n4490 gnd.n4489 585
R9619 gnd.n4490 gnd.n1986 585
R9620 gnd.n4491 gnd.n4486 585
R9621 gnd.n4491 gnd.n1973 585
R9622 gnd.n4494 gnd.n4493 585
R9623 gnd.n4493 gnd.n4492 585
R9624 gnd.n4495 gnd.n4481 585
R9625 gnd.n4481 gnd.n2058 585
R9626 gnd.n4497 gnd.n4496 585
R9627 gnd.n4497 gnd.n2042 585
R9628 gnd.n4498 gnd.n4480 585
R9629 gnd.n4498 gnd.n1112 585
R9630 gnd.n4500 gnd.n4499 585
R9631 gnd.n4499 gnd.n1109 585
R9632 gnd.n4501 gnd.n4475 585
R9633 gnd.n4475 gnd.n2124 585
R9634 gnd.n4503 gnd.n4502 585
R9635 gnd.n4503 gnd.n1100 585
R9636 gnd.n4504 gnd.n4474 585
R9637 gnd.n4504 gnd.n1092 585
R9638 gnd.n4506 gnd.n4505 585
R9639 gnd.n4505 gnd.n1089 585
R9640 gnd.n4507 gnd.n2137 585
R9641 gnd.n2137 gnd.n1081 585
R9642 gnd.n4509 gnd.n4508 585
R9643 gnd.n4510 gnd.n4509 585
R9644 gnd.n2138 gnd.n2136 585
R9645 gnd.n2136 gnd.n1071 585
R9646 gnd.n4468 gnd.n4467 585
R9647 gnd.n4467 gnd.n1068 585
R9648 gnd.n4466 gnd.n2140 585
R9649 gnd.n4466 gnd.n1060 585
R9650 gnd.n4465 gnd.n4464 585
R9651 gnd.n4465 gnd.n1057 585
R9652 gnd.n2142 gnd.n2141 585
R9653 gnd.n2141 gnd.n1049 585
R9654 gnd.n4460 gnd.n4459 585
R9655 gnd.n4459 gnd.n4458 585
R9656 gnd.n2145 gnd.n2144 585
R9657 gnd.n2145 gnd.n1039 585
R9658 gnd.n4424 gnd.n4423 585
R9659 gnd.n4425 gnd.n4424 585
R9660 gnd.n2159 gnd.n2158 585
R9661 gnd.n2158 gnd.n1029 585
R9662 gnd.n4419 gnd.n4418 585
R9663 gnd.n4418 gnd.n1026 585
R9664 gnd.n4417 gnd.n2161 585
R9665 gnd.n4417 gnd.n1018 585
R9666 gnd.n4416 gnd.n4415 585
R9667 gnd.n4416 gnd.n1015 585
R9668 gnd.n2163 gnd.n2162 585
R9669 gnd.n2162 gnd.n1007 585
R9670 gnd.n4411 gnd.n4410 585
R9671 gnd.n4410 gnd.n4409 585
R9672 gnd.n2166 gnd.n2165 585
R9673 gnd.n2166 gnd.n997 585
R9674 gnd.n4375 gnd.n4374 585
R9675 gnd.n4376 gnd.n4375 585
R9676 gnd.n4368 gnd.n4367 585
R9677 gnd.n4367 gnd.n986 585
R9678 gnd.n4370 gnd.n4369 585
R9679 gnd.n4369 gnd.n983 585
R9680 gnd.n969 gnd.n968 585
R9681 gnd.n973 gnd.n969 585
R9682 gnd.n6544 gnd.n6543 585
R9683 gnd.n6543 gnd.n6542 585
R9684 gnd.n6305 gnd.n6304 585
R9685 gnd.n6304 gnd.n6303 585
R9686 gnd.n6306 gnd.n1243 585
R9687 gnd.n1245 gnd.n1243 585
R9688 gnd.n1619 gnd.n1241 585
R9689 gnd.n6012 gnd.n1619 585
R9690 gnd.n6310 gnd.n1240 585
R9691 gnd.n1618 gnd.n1240 585
R9692 gnd.n6311 gnd.n1239 585
R9693 gnd.n6001 gnd.n1239 585
R9694 gnd.n6312 gnd.n1238 585
R9695 gnd.n1626 gnd.n1238 585
R9696 gnd.n1633 gnd.n1236 585
R9697 gnd.n5991 gnd.n1633 585
R9698 gnd.n6316 gnd.n1235 585
R9699 gnd.n1640 gnd.n1235 585
R9700 gnd.n6317 gnd.n1234 585
R9701 gnd.n5983 gnd.n1234 585
R9702 gnd.n6318 gnd.n1233 585
R9703 gnd.n1639 gnd.n1233 585
R9704 gnd.n1647 gnd.n1231 585
R9705 gnd.n5975 gnd.n1647 585
R9706 gnd.n6322 gnd.n1230 585
R9707 gnd.n1646 gnd.n1230 585
R9708 gnd.n6323 gnd.n1229 585
R9709 gnd.n5967 gnd.n1229 585
R9710 gnd.n6324 gnd.n1228 585
R9711 gnd.n1653 gnd.n1228 585
R9712 gnd.n1661 gnd.n1226 585
R9713 gnd.n5959 gnd.n1661 585
R9714 gnd.n6328 gnd.n1225 585
R9715 gnd.n5203 gnd.n1225 585
R9716 gnd.n6329 gnd.n1224 585
R9717 gnd.n5951 gnd.n1224 585
R9718 gnd.n6330 gnd.n1223 585
R9719 gnd.n4988 gnd.n1223 585
R9720 gnd.n1673 gnd.n1221 585
R9721 gnd.n5943 gnd.n1673 585
R9722 gnd.n6334 gnd.n1220 585
R9723 gnd.n5218 gnd.n1220 585
R9724 gnd.n6335 gnd.n1219 585
R9725 gnd.n5935 gnd.n1219 585
R9726 gnd.n6336 gnd.n1218 585
R9727 gnd.n4961 gnd.n1218 585
R9728 gnd.n1687 gnd.n1216 585
R9729 gnd.n5927 gnd.n1687 585
R9730 gnd.n6340 gnd.n1215 585
R9731 gnd.n4972 gnd.n1215 585
R9732 gnd.n6341 gnd.n1214 585
R9733 gnd.n5919 gnd.n1214 585
R9734 gnd.n6342 gnd.n1213 585
R9735 gnd.n1703 gnd.n1213 585
R9736 gnd.n1702 gnd.n1211 585
R9737 gnd.n5911 gnd.n1702 585
R9738 gnd.n6346 gnd.n1210 585
R9739 gnd.n4949 gnd.n1210 585
R9740 gnd.n6347 gnd.n1209 585
R9741 gnd.n5903 gnd.n1209 585
R9742 gnd.n6348 gnd.n1208 585
R9743 gnd.n4942 gnd.n1208 585
R9744 gnd.n1718 gnd.n1206 585
R9745 gnd.n5895 gnd.n1718 585
R9746 gnd.n6352 gnd.n1205 585
R9747 gnd.n4935 gnd.n1205 585
R9748 gnd.n6353 gnd.n1204 585
R9749 gnd.n5887 gnd.n1204 585
R9750 gnd.n6354 gnd.n1203 585
R9751 gnd.n4927 gnd.n1203 585
R9752 gnd.n1732 gnd.n1201 585
R9753 gnd.n5879 gnd.n1732 585
R9754 gnd.n6358 gnd.n1200 585
R9755 gnd.n5269 gnd.n1200 585
R9756 gnd.n6359 gnd.n1199 585
R9757 gnd.n5871 gnd.n1199 585
R9758 gnd.n6360 gnd.n1198 585
R9759 gnd.n4914 gnd.n1198 585
R9760 gnd.n1746 gnd.n1196 585
R9761 gnd.n5863 gnd.n1746 585
R9762 gnd.n6364 gnd.n1195 585
R9763 gnd.n4907 gnd.n1195 585
R9764 gnd.n6365 gnd.n1194 585
R9765 gnd.n5855 gnd.n1194 585
R9766 gnd.n6366 gnd.n1193 585
R9767 gnd.n4900 gnd.n1193 585
R9768 gnd.n1761 gnd.n1191 585
R9769 gnd.n5847 gnd.n1761 585
R9770 gnd.n6370 gnd.n1190 585
R9771 gnd.n5297 gnd.n1190 585
R9772 gnd.n6371 gnd.n1189 585
R9773 gnd.n5839 gnd.n1189 585
R9774 gnd.n6372 gnd.n1188 585
R9775 gnd.n4887 gnd.n1188 585
R9776 gnd.n1776 gnd.n1186 585
R9777 gnd.n5831 gnd.n1776 585
R9778 gnd.n6376 gnd.n1185 585
R9779 gnd.n5312 gnd.n1185 585
R9780 gnd.n6377 gnd.n1184 585
R9781 gnd.n5823 gnd.n1184 585
R9782 gnd.n6378 gnd.n1183 585
R9783 gnd.n4873 gnd.n1183 585
R9784 gnd.n1790 gnd.n1181 585
R9785 gnd.n5815 gnd.n1790 585
R9786 gnd.n6382 gnd.n1180 585
R9787 gnd.n5327 gnd.n1180 585
R9788 gnd.n6383 gnd.n1179 585
R9789 gnd.n5807 gnd.n1179 585
R9790 gnd.n6384 gnd.n1178 585
R9791 gnd.n4860 gnd.n1178 585
R9792 gnd.n1805 gnd.n1176 585
R9793 gnd.n5799 gnd.n1805 585
R9794 gnd.n6388 gnd.n1175 585
R9795 gnd.n5342 gnd.n1175 585
R9796 gnd.n6389 gnd.n1174 585
R9797 gnd.n5791 gnd.n1174 585
R9798 gnd.n6390 gnd.n1173 585
R9799 gnd.n4852 gnd.n1173 585
R9800 gnd.n1820 gnd.n1171 585
R9801 gnd.n5783 gnd.n1820 585
R9802 gnd.n6394 gnd.n1170 585
R9803 gnd.n1828 gnd.n1170 585
R9804 gnd.n6395 gnd.n1169 585
R9805 gnd.n5775 gnd.n1169 585
R9806 gnd.n6396 gnd.n1168 585
R9807 gnd.n4833 gnd.n1168 585
R9808 gnd.n1835 gnd.n1166 585
R9809 gnd.n5767 gnd.n1835 585
R9810 gnd.n6400 gnd.n1165 585
R9811 gnd.n4824 gnd.n1165 585
R9812 gnd.n6401 gnd.n1164 585
R9813 gnd.n5759 gnd.n1164 585
R9814 gnd.n6402 gnd.n1163 585
R9815 gnd.n4816 gnd.n1163 585
R9816 gnd.n1850 gnd.n1161 585
R9817 gnd.n5751 gnd.n1850 585
R9818 gnd.n6406 gnd.n1160 585
R9819 gnd.n5379 gnd.n1160 585
R9820 gnd.n6407 gnd.n1159 585
R9821 gnd.n5743 gnd.n1159 585
R9822 gnd.n6408 gnd.n1158 585
R9823 gnd.n4804 gnd.n1158 585
R9824 gnd.n1863 gnd.n1156 585
R9825 gnd.n5735 gnd.n1863 585
R9826 gnd.n6412 gnd.n1155 585
R9827 gnd.n4795 gnd.n1155 585
R9828 gnd.n6413 gnd.n1154 585
R9829 gnd.n5727 gnd.n1154 585
R9830 gnd.n6414 gnd.n1153 585
R9831 gnd.n4787 gnd.n1153 585
R9832 gnd.n1878 gnd.n1151 585
R9833 gnd.n5719 gnd.n1878 585
R9834 gnd.n6418 gnd.n1150 585
R9835 gnd.n5408 gnd.n1150 585
R9836 gnd.n6419 gnd.n1149 585
R9837 gnd.n5711 gnd.n1149 585
R9838 gnd.n6420 gnd.n1148 585
R9839 gnd.n4773 gnd.n1148 585
R9840 gnd.n1892 gnd.n1146 585
R9841 gnd.n5703 gnd.n1892 585
R9842 gnd.n6424 gnd.n1145 585
R9843 gnd.n5422 gnd.n1145 585
R9844 gnd.n6425 gnd.n1144 585
R9845 gnd.n5695 gnd.n1144 585
R9846 gnd.n6426 gnd.n1143 585
R9847 gnd.n4760 gnd.n1143 585
R9848 gnd.n1906 gnd.n1141 585
R9849 gnd.n5687 gnd.n1906 585
R9850 gnd.n6430 gnd.n1140 585
R9851 gnd.n5437 gnd.n1140 585
R9852 gnd.n6431 gnd.n1139 585
R9853 gnd.n5679 gnd.n1139 585
R9854 gnd.n6432 gnd.n1138 585
R9855 gnd.n4748 gnd.n1138 585
R9856 gnd.n1921 gnd.n1136 585
R9857 gnd.n5671 gnd.n1921 585
R9858 gnd.n6436 gnd.n1135 585
R9859 gnd.n5452 gnd.n1135 585
R9860 gnd.n6437 gnd.n1134 585
R9861 gnd.n5663 gnd.n1134 585
R9862 gnd.n6438 gnd.n1133 585
R9863 gnd.n4652 gnd.n1133 585
R9864 gnd.n1935 gnd.n1131 585
R9865 gnd.n5655 gnd.n1935 585
R9866 gnd.n6442 gnd.n1130 585
R9867 gnd.n1934 gnd.n1130 585
R9868 gnd.n6443 gnd.n1129 585
R9869 gnd.n5647 gnd.n1129 585
R9870 gnd.n6444 gnd.n1128 585
R9871 gnd.n1941 gnd.n1128 585
R9872 gnd.n1947 gnd.n1126 585
R9873 gnd.n5639 gnd.n1947 585
R9874 gnd.n6448 gnd.n1125 585
R9875 gnd.n1954 gnd.n1125 585
R9876 gnd.n6449 gnd.n1124 585
R9877 gnd.n5631 gnd.n1124 585
R9878 gnd.n6450 gnd.n1123 585
R9879 gnd.n1953 gnd.n1123 585
R9880 gnd.n1961 gnd.n1121 585
R9881 gnd.n5623 gnd.n1961 585
R9882 gnd.n6454 gnd.n1120 585
R9883 gnd.n1960 gnd.n1120 585
R9884 gnd.n6455 gnd.n1119 585
R9885 gnd.n5615 gnd.n1119 585
R9886 gnd.n6456 gnd.n1118 585
R9887 gnd.n1967 gnd.n1118 585
R9888 gnd.n5604 gnd.n5603 585
R9889 gnd.n5602 gnd.n1988 585
R9890 gnd.n1990 gnd.n1987 585
R9891 gnd.n5606 gnd.n1987 585
R9892 gnd.n5595 gnd.n1998 585
R9893 gnd.n5594 gnd.n1999 585
R9894 gnd.n2001 gnd.n2000 585
R9895 gnd.n5587 gnd.n2007 585
R9896 gnd.n5586 gnd.n2008 585
R9897 gnd.n2015 gnd.n2009 585
R9898 gnd.n5579 gnd.n2016 585
R9899 gnd.n5578 gnd.n2017 585
R9900 gnd.n2019 gnd.n2018 585
R9901 gnd.n5571 gnd.n2025 585
R9902 gnd.n5570 gnd.n2026 585
R9903 gnd.n2035 gnd.n2027 585
R9904 gnd.n5563 gnd.n2036 585
R9905 gnd.n5562 gnd.n2037 585
R9906 gnd.n2039 gnd.n2038 585
R9907 gnd.n4561 gnd.n4534 585
R9908 gnd.n4560 gnd.n4535 585
R9909 gnd.n4559 gnd.n4536 585
R9910 gnd.n4538 gnd.n4537 585
R9911 gnd.n4555 gnd.n4540 585
R9912 gnd.n4554 gnd.n4541 585
R9913 gnd.n4553 gnd.n4542 585
R9914 gnd.n4550 gnd.n4547 585
R9915 gnd.n4549 gnd.n4548 585
R9916 gnd.n1972 gnd.n1971 585
R9917 gnd.n5609 gnd.n5608 585
R9918 gnd.n6016 gnd.n1247 585
R9919 gnd.n6303 gnd.n1247 585
R9920 gnd.n6015 gnd.n6014 585
R9921 gnd.n6014 gnd.n1245 585
R9922 gnd.n6013 gnd.n1616 585
R9923 gnd.n6013 gnd.n6012 585
R9924 gnd.n1629 gnd.n1617 585
R9925 gnd.n1618 gnd.n1617 585
R9926 gnd.n6000 gnd.n5999 585
R9927 gnd.n6001 gnd.n6000 585
R9928 gnd.n1628 gnd.n1627 585
R9929 gnd.n1627 gnd.n1626 585
R9930 gnd.n5993 gnd.n5992 585
R9931 gnd.n5992 gnd.n5991 585
R9932 gnd.n1632 gnd.n1631 585
R9933 gnd.n1640 gnd.n1632 585
R9934 gnd.n5982 gnd.n5981 585
R9935 gnd.n5983 gnd.n5982 585
R9936 gnd.n1642 gnd.n1641 585
R9937 gnd.n1641 gnd.n1639 585
R9938 gnd.n5977 gnd.n5976 585
R9939 gnd.n5976 gnd.n5975 585
R9940 gnd.n1645 gnd.n1644 585
R9941 gnd.n1646 gnd.n1645 585
R9942 gnd.n5966 gnd.n5965 585
R9943 gnd.n5967 gnd.n5966 585
R9944 gnd.n1656 gnd.n1655 585
R9945 gnd.n1655 gnd.n1653 585
R9946 gnd.n5961 gnd.n5960 585
R9947 gnd.n5960 gnd.n5959 585
R9948 gnd.n1659 gnd.n1658 585
R9949 gnd.n5203 gnd.n1659 585
R9950 gnd.n5950 gnd.n5949 585
R9951 gnd.n5951 gnd.n5950 585
R9952 gnd.n1669 gnd.n1668 585
R9953 gnd.n4988 gnd.n1668 585
R9954 gnd.n5945 gnd.n5944 585
R9955 gnd.n5944 gnd.n5943 585
R9956 gnd.n1672 gnd.n1671 585
R9957 gnd.n5218 gnd.n1672 585
R9958 gnd.n5934 gnd.n5933 585
R9959 gnd.n5935 gnd.n5934 585
R9960 gnd.n1682 gnd.n1681 585
R9961 gnd.n4961 gnd.n1681 585
R9962 gnd.n5929 gnd.n5928 585
R9963 gnd.n5928 gnd.n5927 585
R9964 gnd.n1685 gnd.n1684 585
R9965 gnd.n4972 gnd.n1685 585
R9966 gnd.n5918 gnd.n5917 585
R9967 gnd.n5919 gnd.n5918 585
R9968 gnd.n1697 gnd.n1696 585
R9969 gnd.n1703 gnd.n1696 585
R9970 gnd.n5913 gnd.n5912 585
R9971 gnd.n5912 gnd.n5911 585
R9972 gnd.n1700 gnd.n1699 585
R9973 gnd.n4949 gnd.n1700 585
R9974 gnd.n5902 gnd.n5901 585
R9975 gnd.n5903 gnd.n5902 585
R9976 gnd.n1713 gnd.n1712 585
R9977 gnd.n4942 gnd.n1712 585
R9978 gnd.n5897 gnd.n5896 585
R9979 gnd.n5896 gnd.n5895 585
R9980 gnd.n1716 gnd.n1715 585
R9981 gnd.n4935 gnd.n1716 585
R9982 gnd.n5886 gnd.n5885 585
R9983 gnd.n5887 gnd.n5886 585
R9984 gnd.n1727 gnd.n1726 585
R9985 gnd.n4927 gnd.n1726 585
R9986 gnd.n5881 gnd.n5880 585
R9987 gnd.n5880 gnd.n5879 585
R9988 gnd.n1730 gnd.n1729 585
R9989 gnd.n5269 gnd.n1730 585
R9990 gnd.n5870 gnd.n5869 585
R9991 gnd.n5871 gnd.n5870 585
R9992 gnd.n1741 gnd.n1740 585
R9993 gnd.n4914 gnd.n1740 585
R9994 gnd.n5865 gnd.n5864 585
R9995 gnd.n5864 gnd.n5863 585
R9996 gnd.n1744 gnd.n1743 585
R9997 gnd.n4907 gnd.n1744 585
R9998 gnd.n5854 gnd.n5853 585
R9999 gnd.n5855 gnd.n5854 585
R10000 gnd.n1756 gnd.n1755 585
R10001 gnd.n4900 gnd.n1755 585
R10002 gnd.n5849 gnd.n5848 585
R10003 gnd.n5848 gnd.n5847 585
R10004 gnd.n1759 gnd.n1758 585
R10005 gnd.n5297 gnd.n1759 585
R10006 gnd.n5838 gnd.n5837 585
R10007 gnd.n5839 gnd.n5838 585
R10008 gnd.n1771 gnd.n1770 585
R10009 gnd.n4887 gnd.n1770 585
R10010 gnd.n5833 gnd.n5832 585
R10011 gnd.n5832 gnd.n5831 585
R10012 gnd.n1774 gnd.n1773 585
R10013 gnd.n5312 gnd.n1774 585
R10014 gnd.n5822 gnd.n5821 585
R10015 gnd.n5823 gnd.n5822 585
R10016 gnd.n1785 gnd.n1784 585
R10017 gnd.n4873 gnd.n1784 585
R10018 gnd.n5817 gnd.n5816 585
R10019 gnd.n5816 gnd.n5815 585
R10020 gnd.n1788 gnd.n1787 585
R10021 gnd.n5327 gnd.n1788 585
R10022 gnd.n5806 gnd.n5805 585
R10023 gnd.n5807 gnd.n5806 585
R10024 gnd.n1800 gnd.n1799 585
R10025 gnd.n4860 gnd.n1799 585
R10026 gnd.n5801 gnd.n5800 585
R10027 gnd.n5800 gnd.n5799 585
R10028 gnd.n1803 gnd.n1802 585
R10029 gnd.n5342 gnd.n1803 585
R10030 gnd.n5790 gnd.n5789 585
R10031 gnd.n5791 gnd.n5790 585
R10032 gnd.n1815 gnd.n1814 585
R10033 gnd.n4852 gnd.n1814 585
R10034 gnd.n5785 gnd.n5784 585
R10035 gnd.n5784 gnd.n5783 585
R10036 gnd.n1818 gnd.n1817 585
R10037 gnd.n1828 gnd.n1818 585
R10038 gnd.n5774 gnd.n5773 585
R10039 gnd.n5775 gnd.n5774 585
R10040 gnd.n1831 gnd.n1830 585
R10041 gnd.n4833 gnd.n1830 585
R10042 gnd.n5769 gnd.n5768 585
R10043 gnd.n5768 gnd.n5767 585
R10044 gnd.n1834 gnd.n1833 585
R10045 gnd.n4824 gnd.n1834 585
R10046 gnd.n5758 gnd.n5757 585
R10047 gnd.n5759 gnd.n5758 585
R10048 gnd.n1845 gnd.n1844 585
R10049 gnd.n4816 gnd.n1844 585
R10050 gnd.n5753 gnd.n5752 585
R10051 gnd.n5752 gnd.n5751 585
R10052 gnd.n1848 gnd.n1847 585
R10053 gnd.n5379 gnd.n1848 585
R10054 gnd.n5742 gnd.n5741 585
R10055 gnd.n5743 gnd.n5742 585
R10056 gnd.n1859 gnd.n1858 585
R10057 gnd.n4804 gnd.n1858 585
R10058 gnd.n5737 gnd.n5736 585
R10059 gnd.n5736 gnd.n5735 585
R10060 gnd.n1862 gnd.n1861 585
R10061 gnd.n4795 gnd.n1862 585
R10062 gnd.n5726 gnd.n5725 585
R10063 gnd.n5727 gnd.n5726 585
R10064 gnd.n1873 gnd.n1872 585
R10065 gnd.n4787 gnd.n1872 585
R10066 gnd.n5721 gnd.n5720 585
R10067 gnd.n5720 gnd.n5719 585
R10068 gnd.n1876 gnd.n1875 585
R10069 gnd.n5408 gnd.n1876 585
R10070 gnd.n5710 gnd.n5709 585
R10071 gnd.n5711 gnd.n5710 585
R10072 gnd.n1887 gnd.n1886 585
R10073 gnd.n4773 gnd.n1886 585
R10074 gnd.n5705 gnd.n5704 585
R10075 gnd.n5704 gnd.n5703 585
R10076 gnd.n1890 gnd.n1889 585
R10077 gnd.n5422 gnd.n1890 585
R10078 gnd.n5694 gnd.n5693 585
R10079 gnd.n5695 gnd.n5694 585
R10080 gnd.n1901 gnd.n1900 585
R10081 gnd.n4760 gnd.n1900 585
R10082 gnd.n5689 gnd.n5688 585
R10083 gnd.n5688 gnd.n5687 585
R10084 gnd.n1904 gnd.n1903 585
R10085 gnd.n5437 gnd.n1904 585
R10086 gnd.n5678 gnd.n5677 585
R10087 gnd.n5679 gnd.n5678 585
R10088 gnd.n1916 gnd.n1915 585
R10089 gnd.n4748 gnd.n1915 585
R10090 gnd.n5673 gnd.n5672 585
R10091 gnd.n5672 gnd.n5671 585
R10092 gnd.n1919 gnd.n1918 585
R10093 gnd.n5452 gnd.n1919 585
R10094 gnd.n5662 gnd.n5661 585
R10095 gnd.n5663 gnd.n5662 585
R10096 gnd.n1930 gnd.n1929 585
R10097 gnd.n4652 gnd.n1929 585
R10098 gnd.n5657 gnd.n5656 585
R10099 gnd.n5656 gnd.n5655 585
R10100 gnd.n1933 gnd.n1932 585
R10101 gnd.n1934 gnd.n1933 585
R10102 gnd.n5646 gnd.n5645 585
R10103 gnd.n5647 gnd.n5646 585
R10104 gnd.n1943 gnd.n1942 585
R10105 gnd.n1942 gnd.n1941 585
R10106 gnd.n5641 gnd.n5640 585
R10107 gnd.n5640 gnd.n5639 585
R10108 gnd.n1946 gnd.n1945 585
R10109 gnd.n1954 gnd.n1946 585
R10110 gnd.n5630 gnd.n5629 585
R10111 gnd.n5631 gnd.n5630 585
R10112 gnd.n1956 gnd.n1955 585
R10113 gnd.n1955 gnd.n1953 585
R10114 gnd.n5625 gnd.n5624 585
R10115 gnd.n5624 gnd.n5623 585
R10116 gnd.n1959 gnd.n1958 585
R10117 gnd.n1960 gnd.n1959 585
R10118 gnd.n5614 gnd.n5613 585
R10119 gnd.n5615 gnd.n5614 585
R10120 gnd.n1969 gnd.n1968 585
R10121 gnd.n1968 gnd.n1967 585
R10122 gnd.n6023 gnd.n6022 585
R10123 gnd.n6022 gnd.n1248 585
R10124 gnd.n6024 gnd.n6021 585
R10125 gnd.n6019 gnd.n1614 585
R10126 gnd.n6028 gnd.n1613 585
R10127 gnd.n6032 gnd.n1611 585
R10128 gnd.n6033 gnd.n1610 585
R10129 gnd.n1608 gnd.n1606 585
R10130 gnd.n6037 gnd.n1605 585
R10131 gnd.n6038 gnd.n1603 585
R10132 gnd.n6039 gnd.n1602 585
R10133 gnd.n1600 gnd.n1480 585
R10134 gnd.n1599 gnd.n1598 585
R10135 gnd.n1588 gnd.n1482 585
R10136 gnd.n1590 gnd.n1589 585
R10137 gnd.n1586 gnd.n1492 585
R10138 gnd.n1585 gnd.n1584 585
R10139 gnd.n1572 gnd.n1494 585
R10140 gnd.n1574 gnd.n1573 585
R10141 gnd.n1570 gnd.n1498 585
R10142 gnd.n1569 gnd.n1568 585
R10143 gnd.n1553 gnd.n1500 585
R10144 gnd.n1555 gnd.n1554 585
R10145 gnd.n1551 gnd.n1505 585
R10146 gnd.n1550 gnd.n1549 585
R10147 gnd.n1534 gnd.n1507 585
R10148 gnd.n1536 gnd.n1535 585
R10149 gnd.n1532 gnd.n1512 585
R10150 gnd.n1531 gnd.n1530 585
R10151 gnd.n1514 gnd.n1244 585
R10152 gnd.n5195 gnd.n5002 506.916
R10153 gnd.n5197 gnd.n5000 506.916
R10154 gnd.n4743 gnd.n4678 506.916
R10155 gnd.n5521 gnd.n4655 506.916
R10156 gnd.n6721 gnd.n797 440.005
R10157 gnd.n4680 gnd.t282 389.64
R10158 gnd.n5052 gnd.t230 389.64
R10159 gnd.n5458 gnd.t234 389.64
R10160 gnd.n5046 gnd.t268 389.64
R10161 gnd.n4543 gnd.t248 371.625
R10162 gnd.n122 gnd.t256 371.625
R10163 gnd.n1486 gnd.t271 371.625
R10164 gnd.n2031 gnd.t291 371.625
R10165 gnd.n1308 gnd.t241 371.625
R10166 gnd.n1330 gnd.t223 371.625
R10167 gnd.n201 gnd.t285 371.625
R10168 gnd.n7767 gnd.t202 371.625
R10169 gnd.n4000 gnd.t300 371.625
R10170 gnd.n4032 gnd.t278 371.625
R10171 gnd.n3813 gnd.t297 371.625
R10172 gnd.n2120 gnd.t294 371.625
R10173 gnd.n2098 gnd.t216 371.625
R10174 gnd.n6029 gnd.t212 371.625
R10175 gnd.n2827 gnd.t303 323.425
R10176 gnd.n2372 gnd.t244 323.425
R10177 gnd.n3675 gnd.n3649 289.615
R10178 gnd.n3643 gnd.n3617 289.615
R10179 gnd.n3611 gnd.n3585 289.615
R10180 gnd.n3580 gnd.n3554 289.615
R10181 gnd.n3548 gnd.n3522 289.615
R10182 gnd.n3516 gnd.n3490 289.615
R10183 gnd.n3484 gnd.n3458 289.615
R10184 gnd.n3453 gnd.n3427 289.615
R10185 gnd.n2901 gnd.t274 279.217
R10186 gnd.n2398 gnd.t252 279.217
R10187 gnd.n4662 gnd.t264 260.649
R10188 gnd.n5017 gnd.t267 260.649
R10189 gnd.n5523 gnd.n5522 256.663
R10190 gnd.n5523 gnd.n4621 256.663
R10191 gnd.n5523 gnd.n4622 256.663
R10192 gnd.n5523 gnd.n4623 256.663
R10193 gnd.n5523 gnd.n4624 256.663
R10194 gnd.n5523 gnd.n4625 256.663
R10195 gnd.n5523 gnd.n4626 256.663
R10196 gnd.n5523 gnd.n4627 256.663
R10197 gnd.n5523 gnd.n4628 256.663
R10198 gnd.n5523 gnd.n4629 256.663
R10199 gnd.n5523 gnd.n4630 256.663
R10200 gnd.n5523 gnd.n4631 256.663
R10201 gnd.n5523 gnd.n4632 256.663
R10202 gnd.n5523 gnd.n4633 256.663
R10203 gnd.n5523 gnd.n4634 256.663
R10204 gnd.n5523 gnd.n4635 256.663
R10205 gnd.n5526 gnd.n4619 256.663
R10206 gnd.n5524 gnd.n5523 256.663
R10207 gnd.n5523 gnd.n4636 256.663
R10208 gnd.n5523 gnd.n4637 256.663
R10209 gnd.n5523 gnd.n4638 256.663
R10210 gnd.n5523 gnd.n4639 256.663
R10211 gnd.n5523 gnd.n4640 256.663
R10212 gnd.n5523 gnd.n4641 256.663
R10213 gnd.n5523 gnd.n4642 256.663
R10214 gnd.n5523 gnd.n4643 256.663
R10215 gnd.n5523 gnd.n4644 256.663
R10216 gnd.n5523 gnd.n4645 256.663
R10217 gnd.n5523 gnd.n4646 256.663
R10218 gnd.n5523 gnd.n4647 256.663
R10219 gnd.n5523 gnd.n4648 256.663
R10220 gnd.n5523 gnd.n4649 256.663
R10221 gnd.n5523 gnd.n4650 256.663
R10222 gnd.n5523 gnd.n4651 256.663
R10223 gnd.n5074 gnd.n1654 256.663
R10224 gnd.n5080 gnd.n1654 256.663
R10225 gnd.n5073 gnd.n1654 256.663
R10226 gnd.n5087 gnd.n1654 256.663
R10227 gnd.n5070 gnd.n1654 256.663
R10228 gnd.n5094 gnd.n1654 256.663
R10229 gnd.n5067 gnd.n1654 256.663
R10230 gnd.n5101 gnd.n1654 256.663
R10231 gnd.n5064 gnd.n1654 256.663
R10232 gnd.n5108 gnd.n1654 256.663
R10233 gnd.n5061 gnd.n1654 256.663
R10234 gnd.n5115 gnd.n1654 256.663
R10235 gnd.n5058 gnd.n1654 256.663
R10236 gnd.n5122 gnd.n1654 256.663
R10237 gnd.n5055 gnd.n1654 256.663
R10238 gnd.n5130 gnd.n1654 256.663
R10239 gnd.n5133 gnd.n1305 256.663
R10240 gnd.n5134 gnd.n1654 256.663
R10241 gnd.n5138 gnd.n1654 256.663
R10242 gnd.n5049 gnd.n1654 256.663
R10243 gnd.n5146 gnd.n1654 256.663
R10244 gnd.n5044 gnd.n1654 256.663
R10245 gnd.n5153 gnd.n1654 256.663
R10246 gnd.n5041 gnd.n1654 256.663
R10247 gnd.n5160 gnd.n1654 256.663
R10248 gnd.n5038 gnd.n1654 256.663
R10249 gnd.n5167 gnd.n1654 256.663
R10250 gnd.n5035 gnd.n1654 256.663
R10251 gnd.n5174 gnd.n1654 256.663
R10252 gnd.n5032 gnd.n1654 256.663
R10253 gnd.n5181 gnd.n1654 256.663
R10254 gnd.n5029 gnd.n1654 256.663
R10255 gnd.n5188 gnd.n1654 256.663
R10256 gnd.n5026 gnd.n1654 256.663
R10257 gnd.n3833 gnd.n3808 242.672
R10258 gnd.n3835 gnd.n3808 242.672
R10259 gnd.n3843 gnd.n3808 242.672
R10260 gnd.n3845 gnd.n3808 242.672
R10261 gnd.n3853 gnd.n3808 242.672
R10262 gnd.n3855 gnd.n3808 242.672
R10263 gnd.n3863 gnd.n3808 242.672
R10264 gnd.n3865 gnd.n3808 242.672
R10265 gnd.n3873 gnd.n3808 242.672
R10266 gnd.n5557 gnd.n5556 242.672
R10267 gnd.n5556 gnd.n2057 242.672
R10268 gnd.n5556 gnd.n2056 242.672
R10269 gnd.n5556 gnd.n2054 242.672
R10270 gnd.n5556 gnd.n2052 242.672
R10271 gnd.n5556 gnd.n2051 242.672
R10272 gnd.n5556 gnd.n2049 242.672
R10273 gnd.n5556 gnd.n2047 242.672
R10274 gnd.n5556 gnd.n2046 242.672
R10275 gnd.n6294 gnd.n1275 242.672
R10276 gnd.n6294 gnd.n1276 242.672
R10277 gnd.n6294 gnd.n1277 242.672
R10278 gnd.n6294 gnd.n1278 242.672
R10279 gnd.n6294 gnd.n1279 242.672
R10280 gnd.n6294 gnd.n1280 242.672
R10281 gnd.n6294 gnd.n1281 242.672
R10282 gnd.n6294 gnd.n1282 242.672
R10283 gnd.n6294 gnd.n1283 242.672
R10284 gnd.n128 gnd.n125 242.672
R10285 gnd.n7678 gnd.n128 242.672
R10286 gnd.n7674 gnd.n128 242.672
R10287 gnd.n7671 gnd.n128 242.672
R10288 gnd.n7666 gnd.n128 242.672
R10289 gnd.n7663 gnd.n128 242.672
R10290 gnd.n7658 gnd.n128 242.672
R10291 gnd.n7655 gnd.n128 242.672
R10292 gnd.n7650 gnd.n128 242.672
R10293 gnd.n2955 gnd.n2954 242.672
R10294 gnd.n2955 gnd.n2865 242.672
R10295 gnd.n2955 gnd.n2866 242.672
R10296 gnd.n2955 gnd.n2867 242.672
R10297 gnd.n2955 gnd.n2868 242.672
R10298 gnd.n2955 gnd.n2869 242.672
R10299 gnd.n2955 gnd.n2870 242.672
R10300 gnd.n2955 gnd.n2871 242.672
R10301 gnd.n2955 gnd.n2872 242.672
R10302 gnd.n2955 gnd.n2873 242.672
R10303 gnd.n2955 gnd.n2874 242.672
R10304 gnd.n2955 gnd.n2875 242.672
R10305 gnd.n2956 gnd.n2955 242.672
R10306 gnd.n3807 gnd.n2347 242.672
R10307 gnd.n3807 gnd.n2346 242.672
R10308 gnd.n3807 gnd.n2345 242.672
R10309 gnd.n3807 gnd.n2344 242.672
R10310 gnd.n3807 gnd.n2343 242.672
R10311 gnd.n3807 gnd.n2342 242.672
R10312 gnd.n3807 gnd.n2341 242.672
R10313 gnd.n3807 gnd.n2340 242.672
R10314 gnd.n3807 gnd.n2339 242.672
R10315 gnd.n3807 gnd.n2338 242.672
R10316 gnd.n3807 gnd.n2337 242.672
R10317 gnd.n3807 gnd.n2336 242.672
R10318 gnd.n3807 gnd.n2335 242.672
R10319 gnd.n3039 gnd.n3038 242.672
R10320 gnd.n3038 gnd.n2777 242.672
R10321 gnd.n3038 gnd.n2778 242.672
R10322 gnd.n3038 gnd.n2779 242.672
R10323 gnd.n3038 gnd.n2780 242.672
R10324 gnd.n3038 gnd.n2781 242.672
R10325 gnd.n3038 gnd.n2782 242.672
R10326 gnd.n3038 gnd.n2783 242.672
R10327 gnd.n3807 gnd.n2348 242.672
R10328 gnd.n3807 gnd.n2349 242.672
R10329 gnd.n3807 gnd.n2350 242.672
R10330 gnd.n3807 gnd.n2351 242.672
R10331 gnd.n3807 gnd.n2352 242.672
R10332 gnd.n3807 gnd.n2353 242.672
R10333 gnd.n3807 gnd.n2354 242.672
R10334 gnd.n3807 gnd.n2355 242.672
R10335 gnd.n4186 gnd.n3808 242.672
R10336 gnd.n3976 gnd.n3808 242.672
R10337 gnd.n4179 gnd.n3808 242.672
R10338 gnd.n4173 gnd.n3808 242.672
R10339 gnd.n4171 gnd.n3808 242.672
R10340 gnd.n4165 gnd.n3808 242.672
R10341 gnd.n4163 gnd.n3808 242.672
R10342 gnd.n4157 gnd.n3808 242.672
R10343 gnd.n4155 gnd.n3808 242.672
R10344 gnd.n4149 gnd.n3808 242.672
R10345 gnd.n4147 gnd.n3808 242.672
R10346 gnd.n4141 gnd.n3808 242.672
R10347 gnd.n4139 gnd.n3808 242.672
R10348 gnd.n4133 gnd.n3808 242.672
R10349 gnd.n4131 gnd.n3808 242.672
R10350 gnd.n4125 gnd.n3808 242.672
R10351 gnd.n4123 gnd.n3808 242.672
R10352 gnd.n4030 gnd.n3808 242.672
R10353 gnd.n4113 gnd.n3808 242.672
R10354 gnd.n5556 gnd.n2059 242.672
R10355 gnd.n5556 gnd.n2060 242.672
R10356 gnd.n5556 gnd.n2061 242.672
R10357 gnd.n5556 gnd.n2062 242.672
R10358 gnd.n5556 gnd.n2063 242.672
R10359 gnd.n5556 gnd.n2064 242.672
R10360 gnd.n5556 gnd.n2065 242.672
R10361 gnd.n5556 gnd.n2066 242.672
R10362 gnd.n5556 gnd.n2067 242.672
R10363 gnd.n5556 gnd.n2068 242.672
R10364 gnd.n5556 gnd.n2069 242.672
R10365 gnd.n5527 gnd.n2100 242.672
R10366 gnd.n5556 gnd.n2070 242.672
R10367 gnd.n5556 gnd.n2071 242.672
R10368 gnd.n5556 gnd.n2072 242.672
R10369 gnd.n5556 gnd.n2073 242.672
R10370 gnd.n5556 gnd.n2074 242.672
R10371 gnd.n5556 gnd.n2075 242.672
R10372 gnd.n5556 gnd.n2076 242.672
R10373 gnd.n5556 gnd.n5555 242.672
R10374 gnd.n6294 gnd.n6293 242.672
R10375 gnd.n6294 gnd.n1257 242.672
R10376 gnd.n6294 gnd.n1258 242.672
R10377 gnd.n6294 gnd.n1259 242.672
R10378 gnd.n6294 gnd.n1260 242.672
R10379 gnd.n6294 gnd.n1261 242.672
R10380 gnd.n6294 gnd.n1262 242.672
R10381 gnd.n6294 gnd.n1263 242.672
R10382 gnd.n6262 gnd.n1306 242.672
R10383 gnd.n6294 gnd.n1264 242.672
R10384 gnd.n6294 gnd.n1265 242.672
R10385 gnd.n6294 gnd.n1266 242.672
R10386 gnd.n6294 gnd.n1267 242.672
R10387 gnd.n6294 gnd.n1268 242.672
R10388 gnd.n6294 gnd.n1269 242.672
R10389 gnd.n6294 gnd.n1270 242.672
R10390 gnd.n6294 gnd.n1271 242.672
R10391 gnd.n6294 gnd.n1272 242.672
R10392 gnd.n6294 gnd.n1273 242.672
R10393 gnd.n6294 gnd.n1274 242.672
R10394 gnd.n198 gnd.n128 242.672
R10395 gnd.n7735 gnd.n128 242.672
R10396 gnd.n194 gnd.n128 242.672
R10397 gnd.n7742 gnd.n128 242.672
R10398 gnd.n187 gnd.n128 242.672
R10399 gnd.n7749 gnd.n128 242.672
R10400 gnd.n180 gnd.n128 242.672
R10401 gnd.n7756 gnd.n128 242.672
R10402 gnd.n173 gnd.n128 242.672
R10403 gnd.n7763 gnd.n128 242.672
R10404 gnd.n166 gnd.n128 242.672
R10405 gnd.n7773 gnd.n128 242.672
R10406 gnd.n159 gnd.n128 242.672
R10407 gnd.n7780 gnd.n128 242.672
R10408 gnd.n152 gnd.n128 242.672
R10409 gnd.n7787 gnd.n128 242.672
R10410 gnd.n145 gnd.n128 242.672
R10411 gnd.n7794 gnd.n128 242.672
R10412 gnd.n138 gnd.n128 242.672
R10413 gnd.n5606 gnd.n5605 242.672
R10414 gnd.n5606 gnd.n1974 242.672
R10415 gnd.n5606 gnd.n1975 242.672
R10416 gnd.n5606 gnd.n1976 242.672
R10417 gnd.n5606 gnd.n1977 242.672
R10418 gnd.n5606 gnd.n1978 242.672
R10419 gnd.n5606 gnd.n1979 242.672
R10420 gnd.n5606 gnd.n1980 242.672
R10421 gnd.n5606 gnd.n1981 242.672
R10422 gnd.n5606 gnd.n1982 242.672
R10423 gnd.n5606 gnd.n1983 242.672
R10424 gnd.n5606 gnd.n1984 242.672
R10425 gnd.n5606 gnd.n1985 242.672
R10426 gnd.n5607 gnd.n5606 242.672
R10427 gnd.n6020 gnd.n1248 242.672
R10428 gnd.n1612 gnd.n1248 242.672
R10429 gnd.n1609 gnd.n1248 242.672
R10430 gnd.n1604 gnd.n1248 242.672
R10431 gnd.n1601 gnd.n1248 242.672
R10432 gnd.n1481 gnd.n1248 242.672
R10433 gnd.n1587 gnd.n1248 242.672
R10434 gnd.n1493 gnd.n1248 242.672
R10435 gnd.n1571 gnd.n1248 242.672
R10436 gnd.n1499 gnd.n1248 242.672
R10437 gnd.n1552 gnd.n1248 242.672
R10438 gnd.n1506 gnd.n1248 242.672
R10439 gnd.n1533 gnd.n1248 242.672
R10440 gnd.n1513 gnd.n1248 242.672
R10441 gnd.n135 gnd.n131 240.244
R10442 gnd.n7796 gnd.n7795 240.244
R10443 gnd.n7793 gnd.n139 240.244
R10444 gnd.n7789 gnd.n7788 240.244
R10445 gnd.n7786 gnd.n146 240.244
R10446 gnd.n7782 gnd.n7781 240.244
R10447 gnd.n7779 gnd.n153 240.244
R10448 gnd.n7775 gnd.n7774 240.244
R10449 gnd.n7772 gnd.n160 240.244
R10450 gnd.n7765 gnd.n7764 240.244
R10451 gnd.n7762 gnd.n167 240.244
R10452 gnd.n7758 gnd.n7757 240.244
R10453 gnd.n7755 gnd.n174 240.244
R10454 gnd.n7751 gnd.n7750 240.244
R10455 gnd.n7748 gnd.n181 240.244
R10456 gnd.n7744 gnd.n7743 240.244
R10457 gnd.n7741 gnd.n188 240.244
R10458 gnd.n7737 gnd.n7736 240.244
R10459 gnd.n7734 gnd.n195 240.244
R10460 gnd.n6219 gnd.n1334 240.244
R10461 gnd.n1453 gnd.n1334 240.244
R10462 gnd.n1474 gnd.n1453 240.244
R10463 gnd.n1474 gnd.n1432 240.244
R10464 gnd.n1470 gnd.n1432 240.244
R10465 gnd.n1470 gnd.n1423 240.244
R10466 gnd.n1467 gnd.n1423 240.244
R10467 gnd.n1467 gnd.n1415 240.244
R10468 gnd.n1415 gnd.n1405 240.244
R10469 gnd.n1405 gnd.n1392 240.244
R10470 gnd.n6122 gnd.n1392 240.244
R10471 gnd.n6122 gnd.n1393 240.244
R10472 gnd.n1393 gnd.n1380 240.244
R10473 gnd.n1380 gnd.n1371 240.244
R10474 gnd.n6129 gnd.n1371 240.244
R10475 gnd.n6129 gnd.n1362 240.244
R10476 gnd.n6137 gnd.n1362 240.244
R10477 gnd.n6137 gnd.n400 240.244
R10478 gnd.n400 gnd.n389 240.244
R10479 gnd.n7385 gnd.n389 240.244
R10480 gnd.n7385 gnd.n385 240.244
R10481 gnd.n7397 gnd.n385 240.244
R10482 gnd.n7397 gnd.n368 240.244
R10483 gnd.n7393 gnd.n368 240.244
R10484 gnd.n7393 gnd.n355 240.244
R10485 gnd.n7430 gnd.n355 240.244
R10486 gnd.n7430 gnd.n351 240.244
R10487 gnd.n7443 gnd.n351 240.244
R10488 gnd.n7443 gnd.n313 240.244
R10489 gnd.n7439 gnd.n313 240.244
R10490 gnd.n7439 gnd.n343 240.244
R10491 gnd.n343 gnd.n339 240.244
R10492 gnd.n7460 gnd.n339 240.244
R10493 gnd.n7460 gnd.n335 240.244
R10494 gnd.n7531 gnd.n335 240.244
R10495 gnd.n7531 gnd.n328 240.244
R10496 gnd.n7527 gnd.n328 240.244
R10497 gnd.n7527 gnd.n300 240.244
R10498 gnd.n7524 gnd.n300 240.244
R10499 gnd.n7524 gnd.n291 240.244
R10500 gnd.n7521 gnd.n291 240.244
R10501 gnd.n7521 gnd.n283 240.244
R10502 gnd.n7518 gnd.n283 240.244
R10503 gnd.n7518 gnd.n276 240.244
R10504 gnd.n7515 gnd.n276 240.244
R10505 gnd.n7515 gnd.n270 240.244
R10506 gnd.n7512 gnd.n270 240.244
R10507 gnd.n7512 gnd.n261 240.244
R10508 gnd.n7509 gnd.n261 240.244
R10509 gnd.n7509 gnd.n253 240.244
R10510 gnd.n7506 gnd.n253 240.244
R10511 gnd.n7506 gnd.n245 240.244
R10512 gnd.n7503 gnd.n245 240.244
R10513 gnd.n7503 gnd.n239 240.244
R10514 gnd.n7500 gnd.n239 240.244
R10515 gnd.n7500 gnd.n230 240.244
R10516 gnd.n7497 gnd.n230 240.244
R10517 gnd.n7497 gnd.n223 240.244
R10518 gnd.n7494 gnd.n223 240.244
R10519 gnd.n7494 gnd.n214 240.244
R10520 gnd.n214 gnd.n205 240.244
R10521 gnd.n7725 gnd.n205 240.244
R10522 gnd.n7726 gnd.n7725 240.244
R10523 gnd.n7726 gnd.n127 240.244
R10524 gnd.n1287 gnd.n1286 240.244
R10525 gnd.n6287 gnd.n1286 240.244
R10526 gnd.n6285 gnd.n6284 240.244
R10527 gnd.n6281 gnd.n6280 240.244
R10528 gnd.n6277 gnd.n6276 240.244
R10529 gnd.n6273 gnd.n6272 240.244
R10530 gnd.n6269 gnd.n6268 240.244
R10531 gnd.n6265 gnd.n6264 240.244
R10532 gnd.n6260 gnd.n6259 240.244
R10533 gnd.n6256 gnd.n6255 240.244
R10534 gnd.n6252 gnd.n6251 240.244
R10535 gnd.n6248 gnd.n6247 240.244
R10536 gnd.n6244 gnd.n6243 240.244
R10537 gnd.n6240 gnd.n6239 240.244
R10538 gnd.n6236 gnd.n6235 240.244
R10539 gnd.n6232 gnd.n6231 240.244
R10540 gnd.n6228 gnd.n6227 240.244
R10541 gnd.n1329 gnd.n1328 240.244
R10542 gnd.n6052 gnd.n1288 240.244
R10543 gnd.n6052 gnd.n6045 240.244
R10544 gnd.n6045 gnd.n1430 240.244
R10545 gnd.n6075 gnd.n1430 240.244
R10546 gnd.n6075 gnd.n1425 240.244
R10547 gnd.n6083 gnd.n1425 240.244
R10548 gnd.n6083 gnd.n1426 240.244
R10549 gnd.n1426 gnd.n1403 240.244
R10550 gnd.n6112 gnd.n1403 240.244
R10551 gnd.n6112 gnd.n1397 240.244
R10552 gnd.n6120 gnd.n1397 240.244
R10553 gnd.n6120 gnd.n1399 240.244
R10554 gnd.n1399 gnd.n1369 240.244
R10555 gnd.n6182 gnd.n1369 240.244
R10556 gnd.n6182 gnd.n1365 240.244
R10557 gnd.n6188 gnd.n1365 240.244
R10558 gnd.n6188 gnd.n398 240.244
R10559 gnd.n7375 gnd.n398 240.244
R10560 gnd.n7375 gnd.n393 240.244
R10561 gnd.n7383 gnd.n393 240.244
R10562 gnd.n7383 gnd.n394 240.244
R10563 gnd.n394 gnd.n365 240.244
R10564 gnd.n7421 gnd.n365 240.244
R10565 gnd.n7421 gnd.n366 240.244
R10566 gnd.n366 gnd.n360 240.244
R10567 gnd.n7428 gnd.n360 240.244
R10568 gnd.n7428 gnd.n361 240.244
R10569 gnd.n361 gnd.n310 240.244
R10570 gnd.n7552 gnd.n310 240.244
R10571 gnd.n7552 gnd.n311 240.244
R10572 gnd.n7454 gnd.n311 240.244
R10573 gnd.n7455 gnd.n7454 240.244
R10574 gnd.n7458 gnd.n7455 240.244
R10575 gnd.n7458 gnd.n330 240.244
R10576 gnd.n7533 gnd.n330 240.244
R10577 gnd.n7535 gnd.n7533 240.244
R10578 gnd.n7535 gnd.n301 240.244
R10579 gnd.n7559 gnd.n301 240.244
R10580 gnd.n7559 gnd.n289 240.244
R10581 gnd.n7569 gnd.n289 240.244
R10582 gnd.n7569 gnd.n285 240.244
R10583 gnd.n7575 gnd.n285 240.244
R10584 gnd.n7575 gnd.n275 240.244
R10585 gnd.n7585 gnd.n275 240.244
R10586 gnd.n7585 gnd.n271 240.244
R10587 gnd.n7591 gnd.n271 240.244
R10588 gnd.n7591 gnd.n259 240.244
R10589 gnd.n7601 gnd.n259 240.244
R10590 gnd.n7601 gnd.n255 240.244
R10591 gnd.n7607 gnd.n255 240.244
R10592 gnd.n7607 gnd.n244 240.244
R10593 gnd.n7617 gnd.n244 240.244
R10594 gnd.n7617 gnd.n240 240.244
R10595 gnd.n7623 gnd.n240 240.244
R10596 gnd.n7623 gnd.n228 240.244
R10597 gnd.n7633 gnd.n228 240.244
R10598 gnd.n7633 gnd.n224 240.244
R10599 gnd.n7639 gnd.n224 240.244
R10600 gnd.n7639 gnd.n212 240.244
R10601 gnd.n7717 gnd.n212 240.244
R10602 gnd.n7717 gnd.n208 240.244
R10603 gnd.n7723 gnd.n208 240.244
R10604 gnd.n7723 gnd.n130 240.244
R10605 gnd.n7803 gnd.n130 240.244
R10606 gnd.n2077 gnd.n1108 240.244
R10607 gnd.n5554 gnd.n2078 240.244
R10608 gnd.n5550 gnd.n5549 240.244
R10609 gnd.n5546 gnd.n5545 240.244
R10610 gnd.n5542 gnd.n5541 240.244
R10611 gnd.n5538 gnd.n5537 240.244
R10612 gnd.n5534 gnd.n5533 240.244
R10613 gnd.n5530 gnd.n5529 240.244
R10614 gnd.n4612 gnd.n4611 240.244
R10615 gnd.n4609 gnd.n4608 240.244
R10616 gnd.n4605 gnd.n4604 240.244
R10617 gnd.n4601 gnd.n4600 240.244
R10618 gnd.n4597 gnd.n4596 240.244
R10619 gnd.n4593 gnd.n4592 240.244
R10620 gnd.n4589 gnd.n4588 240.244
R10621 gnd.n4585 gnd.n4584 240.244
R10622 gnd.n4581 gnd.n4580 240.244
R10623 gnd.n4577 gnd.n4576 240.244
R10624 gnd.n4036 gnd.n3809 240.244
R10625 gnd.n4036 gnd.n2328 240.244
R10626 gnd.n4106 gnd.n2328 240.244
R10627 gnd.n4106 gnd.n2321 240.244
R10628 gnd.n4103 gnd.n2321 240.244
R10629 gnd.n4103 gnd.n2313 240.244
R10630 gnd.n4100 gnd.n2313 240.244
R10631 gnd.n4100 gnd.n2304 240.244
R10632 gnd.n4097 gnd.n2304 240.244
R10633 gnd.n4097 gnd.n2296 240.244
R10634 gnd.n4094 gnd.n2296 240.244
R10635 gnd.n4094 gnd.n2289 240.244
R10636 gnd.n4091 gnd.n2289 240.244
R10637 gnd.n4091 gnd.n2281 240.244
R10638 gnd.n4088 gnd.n2281 240.244
R10639 gnd.n4088 gnd.n2272 240.244
R10640 gnd.n4085 gnd.n2272 240.244
R10641 gnd.n4085 gnd.n2264 240.244
R10642 gnd.n4082 gnd.n2264 240.244
R10643 gnd.n4082 gnd.n2257 240.244
R10644 gnd.n4079 gnd.n2257 240.244
R10645 gnd.n4079 gnd.n2249 240.244
R10646 gnd.n4076 gnd.n2249 240.244
R10647 gnd.n4076 gnd.n2240 240.244
R10648 gnd.n4073 gnd.n2240 240.244
R10649 gnd.n4073 gnd.n2232 240.244
R10650 gnd.n4070 gnd.n2232 240.244
R10651 gnd.n4070 gnd.n2226 240.244
R10652 gnd.n4067 gnd.n2226 240.244
R10653 gnd.n4067 gnd.n2217 240.244
R10654 gnd.n2217 gnd.n2207 240.244
R10655 gnd.n4325 gnd.n2207 240.244
R10656 gnd.n4325 gnd.n2208 240.244
R10657 gnd.n2208 gnd.n2190 240.244
R10658 gnd.n2190 gnd.n2184 240.244
R10659 gnd.n4351 gnd.n2184 240.244
R10660 gnd.n4352 gnd.n4351 240.244
R10661 gnd.n4352 gnd.n971 240.244
R10662 gnd.n4358 gnd.n971 240.244
R10663 gnd.n4358 gnd.n984 240.244
R10664 gnd.n4378 gnd.n984 240.244
R10665 gnd.n4378 gnd.n995 240.244
R10666 gnd.n2167 gnd.n995 240.244
R10667 gnd.n2167 gnd.n1005 240.244
R10668 gnd.n4386 gnd.n1005 240.244
R10669 gnd.n4386 gnd.n1016 240.244
R10670 gnd.n4392 gnd.n1016 240.244
R10671 gnd.n4392 gnd.n1027 240.244
R10672 gnd.n4427 gnd.n1027 240.244
R10673 gnd.n4427 gnd.n1037 240.244
R10674 gnd.n2146 gnd.n1037 240.244
R10675 gnd.n2146 gnd.n1047 240.244
R10676 gnd.n4435 gnd.n1047 240.244
R10677 gnd.n4435 gnd.n1058 240.244
R10678 gnd.n4445 gnd.n1058 240.244
R10679 gnd.n4445 gnd.n1069 240.244
R10680 gnd.n2135 gnd.n1069 240.244
R10681 gnd.n2135 gnd.n1079 240.244
R10682 gnd.n4520 gnd.n1079 240.244
R10683 gnd.n4520 gnd.n1090 240.244
R10684 gnd.n4527 gnd.n1090 240.244
R10685 gnd.n4527 gnd.n1101 240.244
R10686 gnd.n4569 gnd.n1101 240.244
R10687 gnd.n4569 gnd.n1110 240.244
R10688 gnd.n4187 gnd.n4185 240.244
R10689 gnd.n4185 gnd.n4184 240.244
R10690 gnd.n4181 gnd.n4180 240.244
R10691 gnd.n4178 gnd.n3981 240.244
R10692 gnd.n4174 gnd.n4172 240.244
R10693 gnd.n4170 gnd.n3987 240.244
R10694 gnd.n4166 gnd.n4164 240.244
R10695 gnd.n4162 gnd.n3993 240.244
R10696 gnd.n4158 gnd.n4156 240.244
R10697 gnd.n4154 gnd.n3999 240.244
R10698 gnd.n4150 gnd.n4148 240.244
R10699 gnd.n4146 gnd.n4008 240.244
R10700 gnd.n4142 gnd.n4140 240.244
R10701 gnd.n4138 gnd.n4014 240.244
R10702 gnd.n4134 gnd.n4132 240.244
R10703 gnd.n4130 gnd.n4020 240.244
R10704 gnd.n4126 gnd.n4124 240.244
R10705 gnd.n4122 gnd.n4026 240.244
R10706 gnd.n4112 gnd.n4031 240.244
R10707 gnd.n4193 gnd.n2327 240.244
R10708 gnd.n4203 gnd.n2327 240.244
R10709 gnd.n4203 gnd.n2323 240.244
R10710 gnd.n4209 gnd.n2323 240.244
R10711 gnd.n4209 gnd.n2311 240.244
R10712 gnd.n4219 gnd.n2311 240.244
R10713 gnd.n4219 gnd.n2307 240.244
R10714 gnd.n4225 gnd.n2307 240.244
R10715 gnd.n4225 gnd.n2295 240.244
R10716 gnd.n4235 gnd.n2295 240.244
R10717 gnd.n4235 gnd.n2291 240.244
R10718 gnd.n4241 gnd.n2291 240.244
R10719 gnd.n4241 gnd.n2279 240.244
R10720 gnd.n4251 gnd.n2279 240.244
R10721 gnd.n4251 gnd.n2275 240.244
R10722 gnd.n4257 gnd.n2275 240.244
R10723 gnd.n4257 gnd.n2263 240.244
R10724 gnd.n4267 gnd.n2263 240.244
R10725 gnd.n4267 gnd.n2259 240.244
R10726 gnd.n4273 gnd.n2259 240.244
R10727 gnd.n4273 gnd.n2247 240.244
R10728 gnd.n4283 gnd.n2247 240.244
R10729 gnd.n4283 gnd.n2243 240.244
R10730 gnd.n4290 gnd.n2243 240.244
R10731 gnd.n4290 gnd.n2231 240.244
R10732 gnd.n4300 gnd.n2231 240.244
R10733 gnd.n4300 gnd.n2228 240.244
R10734 gnd.n4306 gnd.n2228 240.244
R10735 gnd.n4306 gnd.n2215 240.244
R10736 gnd.n4317 gnd.n2215 240.244
R10737 gnd.n4317 gnd.n2213 240.244
R10738 gnd.n4323 gnd.n2213 240.244
R10739 gnd.n4323 gnd.n2189 240.244
R10740 gnd.n4344 gnd.n2189 240.244
R10741 gnd.n4344 gnd.n2187 240.244
R10742 gnd.n4349 gnd.n2187 240.244
R10743 gnd.n4349 gnd.n975 240.244
R10744 gnd.n6540 gnd.n975 240.244
R10745 gnd.n6540 gnd.n976 240.244
R10746 gnd.n6536 gnd.n976 240.244
R10747 gnd.n6536 gnd.n982 240.244
R10748 gnd.n6528 gnd.n982 240.244
R10749 gnd.n6528 gnd.n998 240.244
R10750 gnd.n6524 gnd.n998 240.244
R10751 gnd.n6524 gnd.n1004 240.244
R10752 gnd.n6516 gnd.n1004 240.244
R10753 gnd.n6516 gnd.n1019 240.244
R10754 gnd.n6512 gnd.n1019 240.244
R10755 gnd.n6512 gnd.n1025 240.244
R10756 gnd.n6504 gnd.n1025 240.244
R10757 gnd.n6504 gnd.n1040 240.244
R10758 gnd.n6500 gnd.n1040 240.244
R10759 gnd.n6500 gnd.n1046 240.244
R10760 gnd.n6492 gnd.n1046 240.244
R10761 gnd.n6492 gnd.n1061 240.244
R10762 gnd.n6488 gnd.n1061 240.244
R10763 gnd.n6488 gnd.n1067 240.244
R10764 gnd.n6480 gnd.n1067 240.244
R10765 gnd.n6480 gnd.n1082 240.244
R10766 gnd.n6476 gnd.n1082 240.244
R10767 gnd.n6476 gnd.n1088 240.244
R10768 gnd.n6468 gnd.n1088 240.244
R10769 gnd.n6468 gnd.n1103 240.244
R10770 gnd.n6464 gnd.n1103 240.244
R10771 gnd.n3806 gnd.n2357 240.244
R10772 gnd.n3799 gnd.n3798 240.244
R10773 gnd.n3796 gnd.n3795 240.244
R10774 gnd.n3792 gnd.n3791 240.244
R10775 gnd.n3788 gnd.n3787 240.244
R10776 gnd.n3784 gnd.n3783 240.244
R10777 gnd.n3780 gnd.n3779 240.244
R10778 gnd.n3776 gnd.n3775 240.244
R10779 gnd.n3050 gnd.n2762 240.244
R10780 gnd.n3060 gnd.n2762 240.244
R10781 gnd.n3060 gnd.n2753 240.244
R10782 gnd.n2753 gnd.n2742 240.244
R10783 gnd.n3081 gnd.n2742 240.244
R10784 gnd.n3081 gnd.n2736 240.244
R10785 gnd.n3091 gnd.n2736 240.244
R10786 gnd.n3091 gnd.n2725 240.244
R10787 gnd.n2725 gnd.n2717 240.244
R10788 gnd.n3109 gnd.n2717 240.244
R10789 gnd.n3110 gnd.n3109 240.244
R10790 gnd.n3110 gnd.n2702 240.244
R10791 gnd.n3112 gnd.n2702 240.244
R10792 gnd.n3112 gnd.n2688 240.244
R10793 gnd.n3154 gnd.n2688 240.244
R10794 gnd.n3155 gnd.n3154 240.244
R10795 gnd.n3158 gnd.n3155 240.244
R10796 gnd.n3158 gnd.n2643 240.244
R10797 gnd.n2683 gnd.n2643 240.244
R10798 gnd.n2683 gnd.n2653 240.244
R10799 gnd.n3168 gnd.n2653 240.244
R10800 gnd.n3168 gnd.n2674 240.244
R10801 gnd.n3178 gnd.n2674 240.244
R10802 gnd.n3178 gnd.n2560 240.244
R10803 gnd.n3223 gnd.n2560 240.244
R10804 gnd.n3223 gnd.n2546 240.244
R10805 gnd.n3245 gnd.n2546 240.244
R10806 gnd.n3246 gnd.n3245 240.244
R10807 gnd.n3246 gnd.n2533 240.244
R10808 gnd.n2533 gnd.n2522 240.244
R10809 gnd.n3277 gnd.n2522 240.244
R10810 gnd.n3278 gnd.n3277 240.244
R10811 gnd.n3279 gnd.n3278 240.244
R10812 gnd.n3279 gnd.n2507 240.244
R10813 gnd.n2507 gnd.n2506 240.244
R10814 gnd.n2506 gnd.n2491 240.244
R10815 gnd.n3330 gnd.n2491 240.244
R10816 gnd.n3331 gnd.n3330 240.244
R10817 gnd.n3331 gnd.n2478 240.244
R10818 gnd.n2478 gnd.n2467 240.244
R10819 gnd.n3362 gnd.n2467 240.244
R10820 gnd.n3363 gnd.n3362 240.244
R10821 gnd.n3364 gnd.n3363 240.244
R10822 gnd.n3364 gnd.n2451 240.244
R10823 gnd.n2451 gnd.n2450 240.244
R10824 gnd.n2450 gnd.n2437 240.244
R10825 gnd.n3419 gnd.n2437 240.244
R10826 gnd.n3420 gnd.n3419 240.244
R10827 gnd.n3420 gnd.n2424 240.244
R10828 gnd.n2424 gnd.n2414 240.244
R10829 gnd.n3707 gnd.n2414 240.244
R10830 gnd.n3710 gnd.n3707 240.244
R10831 gnd.n3710 gnd.n3709 240.244
R10832 gnd.n3040 gnd.n2775 240.244
R10833 gnd.n2796 gnd.n2775 240.244
R10834 gnd.n2799 gnd.n2798 240.244
R10835 gnd.n2806 gnd.n2805 240.244
R10836 gnd.n2809 gnd.n2808 240.244
R10837 gnd.n2816 gnd.n2815 240.244
R10838 gnd.n2819 gnd.n2818 240.244
R10839 gnd.n2826 gnd.n2825 240.244
R10840 gnd.n3048 gnd.n2772 240.244
R10841 gnd.n2772 gnd.n2751 240.244
R10842 gnd.n3071 gnd.n2751 240.244
R10843 gnd.n3071 gnd.n2745 240.244
R10844 gnd.n3079 gnd.n2745 240.244
R10845 gnd.n3079 gnd.n2747 240.244
R10846 gnd.n2747 gnd.n2723 240.244
R10847 gnd.n3101 gnd.n2723 240.244
R10848 gnd.n3101 gnd.n2719 240.244
R10849 gnd.n3107 gnd.n2719 240.244
R10850 gnd.n3107 gnd.n2701 240.244
R10851 gnd.n3132 gnd.n2701 240.244
R10852 gnd.n3132 gnd.n2696 240.244
R10853 gnd.n3144 gnd.n2696 240.244
R10854 gnd.n3144 gnd.n2697 240.244
R10855 gnd.n3140 gnd.n2697 240.244
R10856 gnd.n3140 gnd.n2645 240.244
R10857 gnd.n3192 gnd.n2645 240.244
R10858 gnd.n3192 gnd.n2646 240.244
R10859 gnd.n3188 gnd.n2646 240.244
R10860 gnd.n3188 gnd.n2652 240.244
R10861 gnd.n2672 gnd.n2652 240.244
R10862 gnd.n2672 gnd.n2558 240.244
R10863 gnd.n3227 gnd.n2558 240.244
R10864 gnd.n3227 gnd.n2553 240.244
R10865 gnd.n3235 gnd.n2553 240.244
R10866 gnd.n3235 gnd.n2554 240.244
R10867 gnd.n2554 gnd.n2531 240.244
R10868 gnd.n3267 gnd.n2531 240.244
R10869 gnd.n3267 gnd.n2526 240.244
R10870 gnd.n3275 gnd.n2526 240.244
R10871 gnd.n3275 gnd.n2527 240.244
R10872 gnd.n2527 gnd.n2504 240.244
R10873 gnd.n3312 gnd.n2504 240.244
R10874 gnd.n3312 gnd.n2499 240.244
R10875 gnd.n3320 gnd.n2499 240.244
R10876 gnd.n3320 gnd.n2500 240.244
R10877 gnd.n2500 gnd.n2476 240.244
R10878 gnd.n3352 gnd.n2476 240.244
R10879 gnd.n3352 gnd.n2471 240.244
R10880 gnd.n3360 gnd.n2471 240.244
R10881 gnd.n3360 gnd.n2472 240.244
R10882 gnd.n2472 gnd.n2449 240.244
R10883 gnd.n3401 gnd.n2449 240.244
R10884 gnd.n3401 gnd.n2444 240.244
R10885 gnd.n3409 gnd.n2444 240.244
R10886 gnd.n3409 gnd.n2445 240.244
R10887 gnd.n2445 gnd.n2422 240.244
R10888 gnd.n3695 gnd.n2422 240.244
R10889 gnd.n3695 gnd.n2417 240.244
R10890 gnd.n3705 gnd.n2417 240.244
R10891 gnd.n3705 gnd.n2418 240.244
R10892 gnd.n2418 gnd.n2356 240.244
R10893 gnd.n2376 gnd.n2334 240.244
R10894 gnd.n3766 gnd.n3765 240.244
R10895 gnd.n3762 gnd.n3761 240.244
R10896 gnd.n3758 gnd.n3757 240.244
R10897 gnd.n3754 gnd.n3753 240.244
R10898 gnd.n3750 gnd.n3749 240.244
R10899 gnd.n3746 gnd.n3745 240.244
R10900 gnd.n3742 gnd.n3741 240.244
R10901 gnd.n3738 gnd.n3737 240.244
R10902 gnd.n3734 gnd.n3733 240.244
R10903 gnd.n3730 gnd.n3729 240.244
R10904 gnd.n3726 gnd.n3725 240.244
R10905 gnd.n3722 gnd.n3721 240.244
R10906 gnd.n2963 gnd.n2860 240.244
R10907 gnd.n2963 gnd.n2853 240.244
R10908 gnd.n2974 gnd.n2853 240.244
R10909 gnd.n2974 gnd.n2849 240.244
R10910 gnd.n2980 gnd.n2849 240.244
R10911 gnd.n2980 gnd.n2841 240.244
R10912 gnd.n2990 gnd.n2841 240.244
R10913 gnd.n2990 gnd.n2836 240.244
R10914 gnd.n3026 gnd.n2836 240.244
R10915 gnd.n3026 gnd.n2837 240.244
R10916 gnd.n2837 gnd.n2784 240.244
R10917 gnd.n3021 gnd.n2784 240.244
R10918 gnd.n3021 gnd.n3020 240.244
R10919 gnd.n3020 gnd.n2763 240.244
R10920 gnd.n3016 gnd.n2763 240.244
R10921 gnd.n3016 gnd.n2754 240.244
R10922 gnd.n3013 gnd.n2754 240.244
R10923 gnd.n3013 gnd.n3012 240.244
R10924 gnd.n3012 gnd.n2737 240.244
R10925 gnd.n3008 gnd.n2737 240.244
R10926 gnd.n3008 gnd.n2726 240.244
R10927 gnd.n2726 gnd.n2707 240.244
R10928 gnd.n3121 gnd.n2707 240.244
R10929 gnd.n3121 gnd.n2703 240.244
R10930 gnd.n3129 gnd.n2703 240.244
R10931 gnd.n3129 gnd.n2694 240.244
R10932 gnd.n2694 gnd.n2630 240.244
R10933 gnd.n3201 gnd.n2630 240.244
R10934 gnd.n3201 gnd.n2631 240.244
R10935 gnd.n2642 gnd.n2631 240.244
R10936 gnd.n2677 gnd.n2642 240.244
R10937 gnd.n2680 gnd.n2677 240.244
R10938 gnd.n2680 gnd.n2654 240.244
R10939 gnd.n2667 gnd.n2654 240.244
R10940 gnd.n2667 gnd.n2664 240.244
R10941 gnd.n2664 gnd.n2561 240.244
R10942 gnd.n3222 gnd.n2561 240.244
R10943 gnd.n3222 gnd.n2551 240.244
R10944 gnd.n3218 gnd.n2551 240.244
R10945 gnd.n3218 gnd.n2545 240.244
R10946 gnd.n3215 gnd.n2545 240.244
R10947 gnd.n3215 gnd.n2534 240.244
R10948 gnd.n3212 gnd.n2534 240.244
R10949 gnd.n3212 gnd.n2512 240.244
R10950 gnd.n3288 gnd.n2512 240.244
R10951 gnd.n3288 gnd.n2508 240.244
R10952 gnd.n3309 gnd.n2508 240.244
R10953 gnd.n3309 gnd.n2497 240.244
R10954 gnd.n3305 gnd.n2497 240.244
R10955 gnd.n3305 gnd.n2490 240.244
R10956 gnd.n3302 gnd.n2490 240.244
R10957 gnd.n3302 gnd.n2479 240.244
R10958 gnd.n3299 gnd.n2479 240.244
R10959 gnd.n3299 gnd.n2456 240.244
R10960 gnd.n3373 gnd.n2456 240.244
R10961 gnd.n3373 gnd.n2452 240.244
R10962 gnd.n3398 gnd.n2452 240.244
R10963 gnd.n3398 gnd.n2443 240.244
R10964 gnd.n3394 gnd.n2443 240.244
R10965 gnd.n3394 gnd.n2436 240.244
R10966 gnd.n3390 gnd.n2436 240.244
R10967 gnd.n3390 gnd.n2425 240.244
R10968 gnd.n3387 gnd.n2425 240.244
R10969 gnd.n3387 gnd.n2405 240.244
R10970 gnd.n3717 gnd.n2405 240.244
R10971 gnd.n2877 gnd.n2876 240.244
R10972 gnd.n2948 gnd.n2876 240.244
R10973 gnd.n2946 gnd.n2945 240.244
R10974 gnd.n2942 gnd.n2941 240.244
R10975 gnd.n2938 gnd.n2937 240.244
R10976 gnd.n2934 gnd.n2933 240.244
R10977 gnd.n2930 gnd.n2929 240.244
R10978 gnd.n2926 gnd.n2925 240.244
R10979 gnd.n2922 gnd.n2921 240.244
R10980 gnd.n2918 gnd.n2917 240.244
R10981 gnd.n2914 gnd.n2913 240.244
R10982 gnd.n2910 gnd.n2909 240.244
R10983 gnd.n2906 gnd.n2864 240.244
R10984 gnd.n2966 gnd.n2858 240.244
R10985 gnd.n2966 gnd.n2854 240.244
R10986 gnd.n2972 gnd.n2854 240.244
R10987 gnd.n2972 gnd.n2847 240.244
R10988 gnd.n2982 gnd.n2847 240.244
R10989 gnd.n2982 gnd.n2843 240.244
R10990 gnd.n2988 gnd.n2843 240.244
R10991 gnd.n2988 gnd.n2834 240.244
R10992 gnd.n3028 gnd.n2834 240.244
R10993 gnd.n3028 gnd.n2785 240.244
R10994 gnd.n3036 gnd.n2785 240.244
R10995 gnd.n3036 gnd.n2786 240.244
R10996 gnd.n2786 gnd.n2764 240.244
R10997 gnd.n3057 gnd.n2764 240.244
R10998 gnd.n3057 gnd.n2756 240.244
R10999 gnd.n3068 gnd.n2756 240.244
R11000 gnd.n3068 gnd.n2757 240.244
R11001 gnd.n2757 gnd.n2738 240.244
R11002 gnd.n3088 gnd.n2738 240.244
R11003 gnd.n3088 gnd.n2728 240.244
R11004 gnd.n3098 gnd.n2728 240.244
R11005 gnd.n3098 gnd.n2709 240.244
R11006 gnd.n3119 gnd.n2709 240.244
R11007 gnd.n3119 gnd.n2711 240.244
R11008 gnd.n2711 gnd.n2692 240.244
R11009 gnd.n3147 gnd.n2692 240.244
R11010 gnd.n3147 gnd.n2634 240.244
R11011 gnd.n3199 gnd.n2634 240.244
R11012 gnd.n3199 gnd.n2635 240.244
R11013 gnd.n3195 gnd.n2635 240.244
R11014 gnd.n3195 gnd.n2641 240.244
R11015 gnd.n2656 gnd.n2641 240.244
R11016 gnd.n3185 gnd.n2656 240.244
R11017 gnd.n3185 gnd.n2657 240.244
R11018 gnd.n3181 gnd.n2657 240.244
R11019 gnd.n3181 gnd.n2663 240.244
R11020 gnd.n2663 gnd.n2550 240.244
R11021 gnd.n3238 gnd.n2550 240.244
R11022 gnd.n3238 gnd.n2543 240.244
R11023 gnd.n3249 gnd.n2543 240.244
R11024 gnd.n3249 gnd.n2536 240.244
R11025 gnd.n3264 gnd.n2536 240.244
R11026 gnd.n3264 gnd.n2537 240.244
R11027 gnd.n2537 gnd.n2515 240.244
R11028 gnd.n3286 gnd.n2515 240.244
R11029 gnd.n3286 gnd.n2516 240.244
R11030 gnd.n2516 gnd.n2495 240.244
R11031 gnd.n3323 gnd.n2495 240.244
R11032 gnd.n3323 gnd.n2488 240.244
R11033 gnd.n3334 gnd.n2488 240.244
R11034 gnd.n3334 gnd.n2481 240.244
R11035 gnd.n3349 gnd.n2481 240.244
R11036 gnd.n3349 gnd.n2482 240.244
R11037 gnd.n2482 gnd.n2459 240.244
R11038 gnd.n3371 gnd.n2459 240.244
R11039 gnd.n3371 gnd.n2461 240.244
R11040 gnd.n2461 gnd.n2441 240.244
R11041 gnd.n3412 gnd.n2441 240.244
R11042 gnd.n3412 gnd.n2434 240.244
R11043 gnd.n3423 gnd.n2434 240.244
R11044 gnd.n3423 gnd.n2427 240.244
R11045 gnd.n3692 gnd.n2427 240.244
R11046 gnd.n3692 gnd.n2428 240.244
R11047 gnd.n2428 gnd.n2409 240.244
R11048 gnd.n3715 gnd.n2409 240.244
R11049 gnd.n7649 gnd.n7648 240.244
R11050 gnd.n7654 gnd.n7651 240.244
R11051 gnd.n7657 gnd.n7656 240.244
R11052 gnd.n7662 gnd.n7659 240.244
R11053 gnd.n7665 gnd.n7664 240.244
R11054 gnd.n7670 gnd.n7667 240.244
R11055 gnd.n7673 gnd.n7672 240.244
R11056 gnd.n7677 gnd.n7675 240.244
R11057 gnd.n7680 gnd.n7679 240.244
R11058 gnd.n6054 gnd.n1337 240.244
R11059 gnd.n6054 gnd.n1475 240.244
R11060 gnd.n6061 gnd.n1475 240.244
R11061 gnd.n6061 gnd.n1433 240.244
R11062 gnd.n1433 gnd.n1421 240.244
R11063 gnd.n6085 gnd.n1421 240.244
R11064 gnd.n6085 gnd.n1416 240.244
R11065 gnd.n6097 gnd.n1416 240.244
R11066 gnd.n6097 gnd.n1406 240.244
R11067 gnd.n6090 gnd.n1406 240.244
R11068 gnd.n6090 gnd.n1395 240.244
R11069 gnd.n1395 gnd.n1381 240.244
R11070 gnd.n6157 gnd.n1381 240.244
R11071 gnd.n6157 gnd.n1372 240.244
R11072 gnd.n1386 gnd.n1372 240.244
R11073 gnd.n1386 gnd.n1363 240.244
R11074 gnd.n6139 gnd.n1363 240.244
R11075 gnd.n6139 gnd.n401 240.244
R11076 gnd.n6144 gnd.n401 240.244
R11077 gnd.n6144 gnd.n391 240.244
R11078 gnd.n391 gnd.n383 240.244
R11079 gnd.n7399 gnd.n383 240.244
R11080 gnd.n7399 gnd.n369 240.244
R11081 gnd.n378 gnd.n369 240.244
R11082 gnd.n7407 gnd.n378 240.244
R11083 gnd.n7407 gnd.n357 240.244
R11084 gnd.n357 gnd.n349 240.244
R11085 gnd.n7445 gnd.n349 240.244
R11086 gnd.n7445 gnd.n314 240.244
R11087 gnd.n344 gnd.n314 240.244
R11088 gnd.n7452 gnd.n344 240.244
R11089 gnd.n7452 gnd.n345 240.244
R11090 gnd.n345 gnd.n82 240.244
R11091 gnd.n83 gnd.n82 240.244
R11092 gnd.n84 gnd.n83 240.244
R11093 gnd.n329 gnd.n84 240.244
R11094 gnd.n329 gnd.n87 240.244
R11095 gnd.n88 gnd.n87 240.244
R11096 gnd.n89 gnd.n88 240.244
R11097 gnd.n292 gnd.n89 240.244
R11098 gnd.n292 gnd.n92 240.244
R11099 gnd.n93 gnd.n92 240.244
R11100 gnd.n94 gnd.n93 240.244
R11101 gnd.n277 gnd.n94 240.244
R11102 gnd.n277 gnd.n97 240.244
R11103 gnd.n98 gnd.n97 240.244
R11104 gnd.n99 gnd.n98 240.244
R11105 gnd.n262 gnd.n99 240.244
R11106 gnd.n262 gnd.n102 240.244
R11107 gnd.n103 gnd.n102 240.244
R11108 gnd.n104 gnd.n103 240.244
R11109 gnd.n246 gnd.n104 240.244
R11110 gnd.n246 gnd.n107 240.244
R11111 gnd.n108 gnd.n107 240.244
R11112 gnd.n109 gnd.n108 240.244
R11113 gnd.n231 gnd.n109 240.244
R11114 gnd.n231 gnd.n112 240.244
R11115 gnd.n113 gnd.n112 240.244
R11116 gnd.n114 gnd.n113 240.244
R11117 gnd.n215 gnd.n114 240.244
R11118 gnd.n215 gnd.n117 240.244
R11119 gnd.n118 gnd.n117 240.244
R11120 gnd.n119 gnd.n118 240.244
R11121 gnd.n7805 gnd.n119 240.244
R11122 gnd.n1523 gnd.n1522 240.244
R11123 gnd.n1526 gnd.n1525 240.244
R11124 gnd.n1542 gnd.n1541 240.244
R11125 gnd.n1545 gnd.n1544 240.244
R11126 gnd.n1561 gnd.n1560 240.244
R11127 gnd.n1564 gnd.n1563 240.244
R11128 gnd.n1579 gnd.n1578 240.244
R11129 gnd.n1490 gnd.n1489 240.244
R11130 gnd.n1485 gnd.n1284 240.244
R11131 gnd.n6217 gnd.n1340 240.244
R11132 gnd.n1344 gnd.n1340 240.244
R11133 gnd.n1345 gnd.n1344 240.244
R11134 gnd.n1346 gnd.n1345 240.244
R11135 gnd.n1434 gnd.n1346 240.244
R11136 gnd.n1434 gnd.n1349 240.244
R11137 gnd.n1350 gnd.n1349 240.244
R11138 gnd.n1351 gnd.n1350 240.244
R11139 gnd.n6110 gnd.n1351 240.244
R11140 gnd.n6110 gnd.n1354 240.244
R11141 gnd.n1355 gnd.n1354 240.244
R11142 gnd.n1356 gnd.n1355 240.244
R11143 gnd.n6158 gnd.n1356 240.244
R11144 gnd.n6158 gnd.n1359 240.244
R11145 gnd.n1360 gnd.n1359 240.244
R11146 gnd.n6190 gnd.n1360 240.244
R11147 gnd.n6190 gnd.n403 240.244
R11148 gnd.n7373 gnd.n403 240.244
R11149 gnd.n7373 gnd.n404 240.244
R11150 gnd.n404 gnd.n392 240.244
R11151 gnd.n7366 gnd.n392 240.244
R11152 gnd.n7366 gnd.n371 240.244
R11153 gnd.n7419 gnd.n371 240.244
R11154 gnd.n7419 gnd.n372 240.244
R11155 gnd.n7409 gnd.n372 240.244
R11156 gnd.n7409 gnd.n359 240.244
R11157 gnd.n7410 gnd.n359 240.244
R11158 gnd.n7410 gnd.n316 240.244
R11159 gnd.n7550 gnd.n316 240.244
R11160 gnd.n7550 gnd.n317 240.244
R11161 gnd.n322 gnd.n317 240.244
R11162 gnd.n323 gnd.n322 240.244
R11163 gnd.n324 gnd.n323 240.244
R11164 gnd.n333 gnd.n324 240.244
R11165 gnd.n333 gnd.n327 240.244
R11166 gnd.n7537 gnd.n327 240.244
R11167 gnd.n7537 gnd.n298 240.244
R11168 gnd.n7561 gnd.n298 240.244
R11169 gnd.n7561 gnd.n294 240.244
R11170 gnd.n7567 gnd.n294 240.244
R11171 gnd.n7567 gnd.n282 240.244
R11172 gnd.n7577 gnd.n282 240.244
R11173 gnd.n7577 gnd.n278 240.244
R11174 gnd.n7583 gnd.n278 240.244
R11175 gnd.n7583 gnd.n268 240.244
R11176 gnd.n7593 gnd.n268 240.244
R11177 gnd.n7593 gnd.n264 240.244
R11178 gnd.n7599 gnd.n264 240.244
R11179 gnd.n7599 gnd.n252 240.244
R11180 gnd.n7609 gnd.n252 240.244
R11181 gnd.n7609 gnd.n248 240.244
R11182 gnd.n7615 gnd.n248 240.244
R11183 gnd.n7615 gnd.n237 240.244
R11184 gnd.n7625 gnd.n237 240.244
R11185 gnd.n7625 gnd.n233 240.244
R11186 gnd.n7631 gnd.n233 240.244
R11187 gnd.n7631 gnd.n222 240.244
R11188 gnd.n7641 gnd.n222 240.244
R11189 gnd.n7641 gnd.n216 240.244
R11190 gnd.n7715 gnd.n216 240.244
R11191 gnd.n7715 gnd.n217 240.244
R11192 gnd.n217 gnd.n207 240.244
R11193 gnd.n7646 gnd.n207 240.244
R11194 gnd.n7646 gnd.n129 240.244
R11195 gnd.n2044 gnd.n1113 240.244
R11196 gnd.n2045 gnd.n1994 240.244
R11197 gnd.n2048 gnd.n1995 240.244
R11198 gnd.n2004 gnd.n2003 240.244
R11199 gnd.n2050 gnd.n2011 240.244
R11200 gnd.n2053 gnd.n2012 240.244
R11201 gnd.n2022 gnd.n2021 240.244
R11202 gnd.n2055 gnd.n2029 240.244
R11203 gnd.n2041 gnd.n2030 240.244
R11204 gnd.n3971 gnd.n3810 240.244
R11205 gnd.n3971 gnd.n2329 240.244
R11206 gnd.n3967 gnd.n2329 240.244
R11207 gnd.n3967 gnd.n2322 240.244
R11208 gnd.n3964 gnd.n2322 240.244
R11209 gnd.n3964 gnd.n2314 240.244
R11210 gnd.n3961 gnd.n2314 240.244
R11211 gnd.n3961 gnd.n2305 240.244
R11212 gnd.n3958 gnd.n2305 240.244
R11213 gnd.n3958 gnd.n2297 240.244
R11214 gnd.n3955 gnd.n2297 240.244
R11215 gnd.n3955 gnd.n2290 240.244
R11216 gnd.n3952 gnd.n2290 240.244
R11217 gnd.n3952 gnd.n2282 240.244
R11218 gnd.n3949 gnd.n2282 240.244
R11219 gnd.n3949 gnd.n2273 240.244
R11220 gnd.n3946 gnd.n2273 240.244
R11221 gnd.n3946 gnd.n2265 240.244
R11222 gnd.n3943 gnd.n2265 240.244
R11223 gnd.n3943 gnd.n2258 240.244
R11224 gnd.n3940 gnd.n2258 240.244
R11225 gnd.n3940 gnd.n2250 240.244
R11226 gnd.n3937 gnd.n2250 240.244
R11227 gnd.n3937 gnd.n2241 240.244
R11228 gnd.n3934 gnd.n2241 240.244
R11229 gnd.n3934 gnd.n2233 240.244
R11230 gnd.n3931 gnd.n2233 240.244
R11231 gnd.n3931 gnd.n2227 240.244
R11232 gnd.n3928 gnd.n2227 240.244
R11233 gnd.n3928 gnd.n2218 240.244
R11234 gnd.n3925 gnd.n2218 240.244
R11235 gnd.n3925 gnd.n2210 240.244
R11236 gnd.n3910 gnd.n2210 240.244
R11237 gnd.n3910 gnd.n2191 240.244
R11238 gnd.n3913 gnd.n2191 240.244
R11239 gnd.n3913 gnd.n2185 240.244
R11240 gnd.n3914 gnd.n2185 240.244
R11241 gnd.n3914 gnd.n972 240.244
R11242 gnd.n4360 gnd.n972 240.244
R11243 gnd.n4360 gnd.n985 240.244
R11244 gnd.n4366 gnd.n985 240.244
R11245 gnd.n4366 gnd.n996 240.244
R11246 gnd.n4407 gnd.n996 240.244
R11247 gnd.n4407 gnd.n1006 240.244
R11248 gnd.n2172 gnd.n1006 240.244
R11249 gnd.n2172 gnd.n1017 240.244
R11250 gnd.n4394 gnd.n1017 240.244
R11251 gnd.n4394 gnd.n1028 240.244
R11252 gnd.n2157 gnd.n1028 240.244
R11253 gnd.n2157 gnd.n1038 240.244
R11254 gnd.n4456 gnd.n1038 240.244
R11255 gnd.n4456 gnd.n1048 240.244
R11256 gnd.n2151 gnd.n1048 240.244
R11257 gnd.n2151 gnd.n1059 240.244
R11258 gnd.n4447 gnd.n1059 240.244
R11259 gnd.n4447 gnd.n1070 240.244
R11260 gnd.n4512 gnd.n1070 240.244
R11261 gnd.n4512 gnd.n1080 240.244
R11262 gnd.n4518 gnd.n1080 240.244
R11263 gnd.n4518 gnd.n1091 240.244
R11264 gnd.n4529 gnd.n1091 240.244
R11265 gnd.n4529 gnd.n1102 240.244
R11266 gnd.n4567 gnd.n1102 240.244
R11267 gnd.n4567 gnd.n1111 240.244
R11268 gnd.n3836 gnd.n3834 240.244
R11269 gnd.n3842 gnd.n3828 240.244
R11270 gnd.n3846 gnd.n3844 240.244
R11271 gnd.n3852 gnd.n3824 240.244
R11272 gnd.n3856 gnd.n3854 240.244
R11273 gnd.n3862 gnd.n3820 240.244
R11274 gnd.n3866 gnd.n3864 240.244
R11275 gnd.n3872 gnd.n3816 240.244
R11276 gnd.n3875 gnd.n3874 240.244
R11277 gnd.n4195 gnd.n2330 240.244
R11278 gnd.n4201 gnd.n2330 240.244
R11279 gnd.n4201 gnd.n2319 240.244
R11280 gnd.n4211 gnd.n2319 240.244
R11281 gnd.n4211 gnd.n2315 240.244
R11282 gnd.n4217 gnd.n2315 240.244
R11283 gnd.n4217 gnd.n2302 240.244
R11284 gnd.n4227 gnd.n2302 240.244
R11285 gnd.n4227 gnd.n2298 240.244
R11286 gnd.n4233 gnd.n2298 240.244
R11287 gnd.n4233 gnd.n2287 240.244
R11288 gnd.n4243 gnd.n2287 240.244
R11289 gnd.n4243 gnd.n2283 240.244
R11290 gnd.n4249 gnd.n2283 240.244
R11291 gnd.n4249 gnd.n2270 240.244
R11292 gnd.n4259 gnd.n2270 240.244
R11293 gnd.n4259 gnd.n2266 240.244
R11294 gnd.n4265 gnd.n2266 240.244
R11295 gnd.n4265 gnd.n2255 240.244
R11296 gnd.n4275 gnd.n2255 240.244
R11297 gnd.n4275 gnd.n2251 240.244
R11298 gnd.n4281 gnd.n2251 240.244
R11299 gnd.n4281 gnd.n2238 240.244
R11300 gnd.n4292 gnd.n2238 240.244
R11301 gnd.n4292 gnd.n2234 240.244
R11302 gnd.n4298 gnd.n2234 240.244
R11303 gnd.n4298 gnd.n2224 240.244
R11304 gnd.n4308 gnd.n2224 240.244
R11305 gnd.n4308 gnd.n2219 240.244
R11306 gnd.n4315 gnd.n2219 240.244
R11307 gnd.n4315 gnd.n2220 240.244
R11308 gnd.n2220 gnd.n2212 240.244
R11309 gnd.n2212 gnd.n2194 240.244
R11310 gnd.n4342 gnd.n2194 240.244
R11311 gnd.n4342 gnd.n2195 240.244
R11312 gnd.n2195 gnd.n2186 240.244
R11313 gnd.n4337 gnd.n2186 240.244
R11314 gnd.n4337 gnd.n974 240.244
R11315 gnd.n987 gnd.n974 240.244
R11316 gnd.n6534 gnd.n987 240.244
R11317 gnd.n6534 gnd.n988 240.244
R11318 gnd.n6530 gnd.n988 240.244
R11319 gnd.n6530 gnd.n994 240.244
R11320 gnd.n6522 gnd.n994 240.244
R11321 gnd.n6522 gnd.n1008 240.244
R11322 gnd.n6518 gnd.n1008 240.244
R11323 gnd.n6518 gnd.n1014 240.244
R11324 gnd.n6510 gnd.n1014 240.244
R11325 gnd.n6510 gnd.n1030 240.244
R11326 gnd.n6506 gnd.n1030 240.244
R11327 gnd.n6506 gnd.n1036 240.244
R11328 gnd.n6498 gnd.n1036 240.244
R11329 gnd.n6498 gnd.n1050 240.244
R11330 gnd.n6494 gnd.n1050 240.244
R11331 gnd.n6494 gnd.n1056 240.244
R11332 gnd.n6486 gnd.n1056 240.244
R11333 gnd.n6486 gnd.n1072 240.244
R11334 gnd.n6482 gnd.n1072 240.244
R11335 gnd.n6482 gnd.n1078 240.244
R11336 gnd.n6474 gnd.n1078 240.244
R11337 gnd.n6474 gnd.n1093 240.244
R11338 gnd.n6470 gnd.n1093 240.244
R11339 gnd.n6470 gnd.n1099 240.244
R11340 gnd.n6462 gnd.n1099 240.244
R11341 gnd.n6720 gnd.n796 240.244
R11342 gnd.n6724 gnd.n796 240.244
R11343 gnd.n6724 gnd.n792 240.244
R11344 gnd.n6730 gnd.n792 240.244
R11345 gnd.n6730 gnd.n790 240.244
R11346 gnd.n6734 gnd.n790 240.244
R11347 gnd.n6734 gnd.n786 240.244
R11348 gnd.n6740 gnd.n786 240.244
R11349 gnd.n6740 gnd.n784 240.244
R11350 gnd.n6744 gnd.n784 240.244
R11351 gnd.n6744 gnd.n780 240.244
R11352 gnd.n6750 gnd.n780 240.244
R11353 gnd.n6750 gnd.n778 240.244
R11354 gnd.n6754 gnd.n778 240.244
R11355 gnd.n6754 gnd.n774 240.244
R11356 gnd.n6760 gnd.n774 240.244
R11357 gnd.n6760 gnd.n772 240.244
R11358 gnd.n6764 gnd.n772 240.244
R11359 gnd.n6764 gnd.n768 240.244
R11360 gnd.n6770 gnd.n768 240.244
R11361 gnd.n6770 gnd.n766 240.244
R11362 gnd.n6774 gnd.n766 240.244
R11363 gnd.n6774 gnd.n762 240.244
R11364 gnd.n6780 gnd.n762 240.244
R11365 gnd.n6780 gnd.n760 240.244
R11366 gnd.n6784 gnd.n760 240.244
R11367 gnd.n6784 gnd.n756 240.244
R11368 gnd.n6790 gnd.n756 240.244
R11369 gnd.n6790 gnd.n754 240.244
R11370 gnd.n6794 gnd.n754 240.244
R11371 gnd.n6794 gnd.n750 240.244
R11372 gnd.n6800 gnd.n750 240.244
R11373 gnd.n6800 gnd.n748 240.244
R11374 gnd.n6804 gnd.n748 240.244
R11375 gnd.n6804 gnd.n744 240.244
R11376 gnd.n6810 gnd.n744 240.244
R11377 gnd.n6810 gnd.n742 240.244
R11378 gnd.n6814 gnd.n742 240.244
R11379 gnd.n6814 gnd.n738 240.244
R11380 gnd.n6820 gnd.n738 240.244
R11381 gnd.n6820 gnd.n736 240.244
R11382 gnd.n6824 gnd.n736 240.244
R11383 gnd.n6824 gnd.n732 240.244
R11384 gnd.n6830 gnd.n732 240.244
R11385 gnd.n6830 gnd.n730 240.244
R11386 gnd.n6834 gnd.n730 240.244
R11387 gnd.n6834 gnd.n726 240.244
R11388 gnd.n6840 gnd.n726 240.244
R11389 gnd.n6840 gnd.n724 240.244
R11390 gnd.n6844 gnd.n724 240.244
R11391 gnd.n6844 gnd.n720 240.244
R11392 gnd.n6850 gnd.n720 240.244
R11393 gnd.n6850 gnd.n718 240.244
R11394 gnd.n6854 gnd.n718 240.244
R11395 gnd.n6854 gnd.n714 240.244
R11396 gnd.n6860 gnd.n714 240.244
R11397 gnd.n6860 gnd.n712 240.244
R11398 gnd.n6864 gnd.n712 240.244
R11399 gnd.n6864 gnd.n708 240.244
R11400 gnd.n6870 gnd.n708 240.244
R11401 gnd.n6870 gnd.n706 240.244
R11402 gnd.n6874 gnd.n706 240.244
R11403 gnd.n6874 gnd.n702 240.244
R11404 gnd.n6880 gnd.n702 240.244
R11405 gnd.n6880 gnd.n700 240.244
R11406 gnd.n6884 gnd.n700 240.244
R11407 gnd.n6884 gnd.n696 240.244
R11408 gnd.n6890 gnd.n696 240.244
R11409 gnd.n6890 gnd.n694 240.244
R11410 gnd.n6894 gnd.n694 240.244
R11411 gnd.n6894 gnd.n690 240.244
R11412 gnd.n6900 gnd.n690 240.244
R11413 gnd.n6900 gnd.n688 240.244
R11414 gnd.n6904 gnd.n688 240.244
R11415 gnd.n6904 gnd.n684 240.244
R11416 gnd.n6910 gnd.n684 240.244
R11417 gnd.n6910 gnd.n682 240.244
R11418 gnd.n6914 gnd.n682 240.244
R11419 gnd.n6914 gnd.n678 240.244
R11420 gnd.n6920 gnd.n678 240.244
R11421 gnd.n6920 gnd.n676 240.244
R11422 gnd.n6924 gnd.n676 240.244
R11423 gnd.n6924 gnd.n672 240.244
R11424 gnd.n6930 gnd.n672 240.244
R11425 gnd.n6930 gnd.n670 240.244
R11426 gnd.n6934 gnd.n670 240.244
R11427 gnd.n6934 gnd.n666 240.244
R11428 gnd.n6940 gnd.n666 240.244
R11429 gnd.n6940 gnd.n664 240.244
R11430 gnd.n6944 gnd.n664 240.244
R11431 gnd.n6944 gnd.n660 240.244
R11432 gnd.n6950 gnd.n660 240.244
R11433 gnd.n6950 gnd.n658 240.244
R11434 gnd.n6954 gnd.n658 240.244
R11435 gnd.n6954 gnd.n654 240.244
R11436 gnd.n6960 gnd.n654 240.244
R11437 gnd.n6960 gnd.n652 240.244
R11438 gnd.n6964 gnd.n652 240.244
R11439 gnd.n6964 gnd.n648 240.244
R11440 gnd.n6970 gnd.n648 240.244
R11441 gnd.n6970 gnd.n646 240.244
R11442 gnd.n6974 gnd.n646 240.244
R11443 gnd.n6974 gnd.n642 240.244
R11444 gnd.n6980 gnd.n642 240.244
R11445 gnd.n6980 gnd.n640 240.244
R11446 gnd.n6984 gnd.n640 240.244
R11447 gnd.n6984 gnd.n636 240.244
R11448 gnd.n6990 gnd.n636 240.244
R11449 gnd.n6990 gnd.n634 240.244
R11450 gnd.n6994 gnd.n634 240.244
R11451 gnd.n6994 gnd.n630 240.244
R11452 gnd.n7000 gnd.n630 240.244
R11453 gnd.n7000 gnd.n628 240.244
R11454 gnd.n7004 gnd.n628 240.244
R11455 gnd.n7004 gnd.n624 240.244
R11456 gnd.n7010 gnd.n624 240.244
R11457 gnd.n7010 gnd.n622 240.244
R11458 gnd.n7014 gnd.n622 240.244
R11459 gnd.n7014 gnd.n618 240.244
R11460 gnd.n7020 gnd.n618 240.244
R11461 gnd.n7020 gnd.n616 240.244
R11462 gnd.n7024 gnd.n616 240.244
R11463 gnd.n7024 gnd.n612 240.244
R11464 gnd.n7030 gnd.n612 240.244
R11465 gnd.n7030 gnd.n610 240.244
R11466 gnd.n7034 gnd.n610 240.244
R11467 gnd.n7034 gnd.n606 240.244
R11468 gnd.n7040 gnd.n606 240.244
R11469 gnd.n7040 gnd.n604 240.244
R11470 gnd.n7044 gnd.n604 240.244
R11471 gnd.n7044 gnd.n600 240.244
R11472 gnd.n7050 gnd.n600 240.244
R11473 gnd.n7050 gnd.n598 240.244
R11474 gnd.n7054 gnd.n598 240.244
R11475 gnd.n7054 gnd.n594 240.244
R11476 gnd.n7060 gnd.n594 240.244
R11477 gnd.n7060 gnd.n592 240.244
R11478 gnd.n7064 gnd.n592 240.244
R11479 gnd.n7064 gnd.n588 240.244
R11480 gnd.n7070 gnd.n588 240.244
R11481 gnd.n7070 gnd.n586 240.244
R11482 gnd.n7074 gnd.n586 240.244
R11483 gnd.n7074 gnd.n582 240.244
R11484 gnd.n7080 gnd.n582 240.244
R11485 gnd.n7080 gnd.n580 240.244
R11486 gnd.n7084 gnd.n580 240.244
R11487 gnd.n7084 gnd.n576 240.244
R11488 gnd.n7090 gnd.n576 240.244
R11489 gnd.n7090 gnd.n574 240.244
R11490 gnd.n7094 gnd.n574 240.244
R11491 gnd.n7094 gnd.n570 240.244
R11492 gnd.n7100 gnd.n570 240.244
R11493 gnd.n7100 gnd.n568 240.244
R11494 gnd.n7104 gnd.n568 240.244
R11495 gnd.n7104 gnd.n564 240.244
R11496 gnd.n7110 gnd.n564 240.244
R11497 gnd.n7110 gnd.n562 240.244
R11498 gnd.n7114 gnd.n562 240.244
R11499 gnd.n7114 gnd.n558 240.244
R11500 gnd.n7120 gnd.n558 240.244
R11501 gnd.n7120 gnd.n556 240.244
R11502 gnd.n7124 gnd.n556 240.244
R11503 gnd.n7124 gnd.n552 240.244
R11504 gnd.n7131 gnd.n552 240.244
R11505 gnd.n7131 gnd.n550 240.244
R11506 gnd.n7135 gnd.n550 240.244
R11507 gnd.n7135 gnd.n547 240.244
R11508 gnd.n7141 gnd.n545 240.244
R11509 gnd.n7145 gnd.n545 240.244
R11510 gnd.n7145 gnd.n541 240.244
R11511 gnd.n7151 gnd.n541 240.244
R11512 gnd.n7151 gnd.n539 240.244
R11513 gnd.n7155 gnd.n539 240.244
R11514 gnd.n7155 gnd.n535 240.244
R11515 gnd.n7161 gnd.n535 240.244
R11516 gnd.n7161 gnd.n533 240.244
R11517 gnd.n7165 gnd.n533 240.244
R11518 gnd.n7165 gnd.n529 240.244
R11519 gnd.n7171 gnd.n529 240.244
R11520 gnd.n7171 gnd.n527 240.244
R11521 gnd.n7175 gnd.n527 240.244
R11522 gnd.n7175 gnd.n523 240.244
R11523 gnd.n7181 gnd.n523 240.244
R11524 gnd.n7181 gnd.n521 240.244
R11525 gnd.n7185 gnd.n521 240.244
R11526 gnd.n7185 gnd.n517 240.244
R11527 gnd.n7191 gnd.n517 240.244
R11528 gnd.n7191 gnd.n515 240.244
R11529 gnd.n7195 gnd.n515 240.244
R11530 gnd.n7195 gnd.n511 240.244
R11531 gnd.n7201 gnd.n511 240.244
R11532 gnd.n7201 gnd.n509 240.244
R11533 gnd.n7205 gnd.n509 240.244
R11534 gnd.n7205 gnd.n505 240.244
R11535 gnd.n7211 gnd.n505 240.244
R11536 gnd.n7211 gnd.n503 240.244
R11537 gnd.n7215 gnd.n503 240.244
R11538 gnd.n7215 gnd.n499 240.244
R11539 gnd.n7221 gnd.n499 240.244
R11540 gnd.n7221 gnd.n497 240.244
R11541 gnd.n7225 gnd.n497 240.244
R11542 gnd.n7225 gnd.n493 240.244
R11543 gnd.n7231 gnd.n493 240.244
R11544 gnd.n7231 gnd.n491 240.244
R11545 gnd.n7235 gnd.n491 240.244
R11546 gnd.n7235 gnd.n487 240.244
R11547 gnd.n7241 gnd.n487 240.244
R11548 gnd.n7241 gnd.n485 240.244
R11549 gnd.n7245 gnd.n485 240.244
R11550 gnd.n7245 gnd.n481 240.244
R11551 gnd.n7251 gnd.n481 240.244
R11552 gnd.n7251 gnd.n479 240.244
R11553 gnd.n7255 gnd.n479 240.244
R11554 gnd.n7255 gnd.n475 240.244
R11555 gnd.n7261 gnd.n475 240.244
R11556 gnd.n7261 gnd.n473 240.244
R11557 gnd.n7265 gnd.n473 240.244
R11558 gnd.n7265 gnd.n469 240.244
R11559 gnd.n7271 gnd.n469 240.244
R11560 gnd.n7271 gnd.n467 240.244
R11561 gnd.n7275 gnd.n467 240.244
R11562 gnd.n7275 gnd.n463 240.244
R11563 gnd.n7281 gnd.n463 240.244
R11564 gnd.n7281 gnd.n461 240.244
R11565 gnd.n7285 gnd.n461 240.244
R11566 gnd.n7285 gnd.n457 240.244
R11567 gnd.n7291 gnd.n457 240.244
R11568 gnd.n7291 gnd.n455 240.244
R11569 gnd.n7295 gnd.n455 240.244
R11570 gnd.n7295 gnd.n451 240.244
R11571 gnd.n7301 gnd.n451 240.244
R11572 gnd.n7301 gnd.n449 240.244
R11573 gnd.n7305 gnd.n449 240.244
R11574 gnd.n7305 gnd.n445 240.244
R11575 gnd.n7311 gnd.n445 240.244
R11576 gnd.n7311 gnd.n443 240.244
R11577 gnd.n7315 gnd.n443 240.244
R11578 gnd.n7315 gnd.n439 240.244
R11579 gnd.n7321 gnd.n439 240.244
R11580 gnd.n7321 gnd.n437 240.244
R11581 gnd.n7325 gnd.n437 240.244
R11582 gnd.n7325 gnd.n433 240.244
R11583 gnd.n7331 gnd.n433 240.244
R11584 gnd.n7331 gnd.n431 240.244
R11585 gnd.n7335 gnd.n431 240.244
R11586 gnd.n7335 gnd.n427 240.244
R11587 gnd.n7341 gnd.n427 240.244
R11588 gnd.n7341 gnd.n425 240.244
R11589 gnd.n7346 gnd.n425 240.244
R11590 gnd.n7346 gnd.n421 240.244
R11591 gnd.n7352 gnd.n421 240.244
R11592 gnd.n6543 gnd.n969 240.244
R11593 gnd.n4369 gnd.n969 240.244
R11594 gnd.n4369 gnd.n4367 240.244
R11595 gnd.n4375 gnd.n4367 240.244
R11596 gnd.n4375 gnd.n2166 240.244
R11597 gnd.n4410 gnd.n2166 240.244
R11598 gnd.n4410 gnd.n2162 240.244
R11599 gnd.n4416 gnd.n2162 240.244
R11600 gnd.n4417 gnd.n4416 240.244
R11601 gnd.n4418 gnd.n4417 240.244
R11602 gnd.n4418 gnd.n2158 240.244
R11603 gnd.n4424 gnd.n2158 240.244
R11604 gnd.n4424 gnd.n2145 240.244
R11605 gnd.n4459 gnd.n2145 240.244
R11606 gnd.n4459 gnd.n2141 240.244
R11607 gnd.n4465 gnd.n2141 240.244
R11608 gnd.n4466 gnd.n4465 240.244
R11609 gnd.n4467 gnd.n4466 240.244
R11610 gnd.n4467 gnd.n2136 240.244
R11611 gnd.n4509 gnd.n2136 240.244
R11612 gnd.n4509 gnd.n2137 240.244
R11613 gnd.n4505 gnd.n2137 240.244
R11614 gnd.n4505 gnd.n4504 240.244
R11615 gnd.n4504 gnd.n4503 240.244
R11616 gnd.n4503 gnd.n4475 240.244
R11617 gnd.n4499 gnd.n4475 240.244
R11618 gnd.n4499 gnd.n4498 240.244
R11619 gnd.n4498 gnd.n4497 240.244
R11620 gnd.n4497 gnd.n4481 240.244
R11621 gnd.n4493 gnd.n4481 240.244
R11622 gnd.n4493 gnd.n4491 240.244
R11623 gnd.n4491 gnd.n4490 240.244
R11624 gnd.n4490 gnd.n1966 240.244
R11625 gnd.n5616 gnd.n1966 240.244
R11626 gnd.n5616 gnd.n1962 240.244
R11627 gnd.n5622 gnd.n1962 240.244
R11628 gnd.n5622 gnd.n1952 240.244
R11629 gnd.n5632 gnd.n1952 240.244
R11630 gnd.n5632 gnd.n1948 240.244
R11631 gnd.n5638 gnd.n1948 240.244
R11632 gnd.n5638 gnd.n1940 240.244
R11633 gnd.n5648 gnd.n1940 240.244
R11634 gnd.n5648 gnd.n1936 240.244
R11635 gnd.n5654 gnd.n1936 240.244
R11636 gnd.n5654 gnd.n1927 240.244
R11637 gnd.n5664 gnd.n1927 240.244
R11638 gnd.n5664 gnd.n1923 240.244
R11639 gnd.n5670 gnd.n1923 240.244
R11640 gnd.n5670 gnd.n1912 240.244
R11641 gnd.n5680 gnd.n1912 240.244
R11642 gnd.n5680 gnd.n1908 240.244
R11643 gnd.n5686 gnd.n1908 240.244
R11644 gnd.n5686 gnd.n1898 240.244
R11645 gnd.n5696 gnd.n1898 240.244
R11646 gnd.n5696 gnd.n1894 240.244
R11647 gnd.n5702 gnd.n1894 240.244
R11648 gnd.n5702 gnd.n1884 240.244
R11649 gnd.n5712 gnd.n1884 240.244
R11650 gnd.n5712 gnd.n1880 240.244
R11651 gnd.n5718 gnd.n1880 240.244
R11652 gnd.n5718 gnd.n1869 240.244
R11653 gnd.n5728 gnd.n1869 240.244
R11654 gnd.n5728 gnd.n1865 240.244
R11655 gnd.n5734 gnd.n1865 240.244
R11656 gnd.n5734 gnd.n1856 240.244
R11657 gnd.n5744 gnd.n1856 240.244
R11658 gnd.n5744 gnd.n1852 240.244
R11659 gnd.n5750 gnd.n1852 240.244
R11660 gnd.n5750 gnd.n1841 240.244
R11661 gnd.n5760 gnd.n1841 240.244
R11662 gnd.n5760 gnd.n1837 240.244
R11663 gnd.n5766 gnd.n1837 240.244
R11664 gnd.n5766 gnd.n1826 240.244
R11665 gnd.n5776 gnd.n1826 240.244
R11666 gnd.n5776 gnd.n1822 240.244
R11667 gnd.n5782 gnd.n1822 240.244
R11668 gnd.n5782 gnd.n1811 240.244
R11669 gnd.n5792 gnd.n1811 240.244
R11670 gnd.n5792 gnd.n1807 240.244
R11671 gnd.n5798 gnd.n1807 240.244
R11672 gnd.n5798 gnd.n1796 240.244
R11673 gnd.n5808 gnd.n1796 240.244
R11674 gnd.n5808 gnd.n1792 240.244
R11675 gnd.n5814 gnd.n1792 240.244
R11676 gnd.n5814 gnd.n1782 240.244
R11677 gnd.n5824 gnd.n1782 240.244
R11678 gnd.n5824 gnd.n1778 240.244
R11679 gnd.n5830 gnd.n1778 240.244
R11680 gnd.n5830 gnd.n1767 240.244
R11681 gnd.n5840 gnd.n1767 240.244
R11682 gnd.n5840 gnd.n1763 240.244
R11683 gnd.n5846 gnd.n1763 240.244
R11684 gnd.n5846 gnd.n1752 240.244
R11685 gnd.n5856 gnd.n1752 240.244
R11686 gnd.n5856 gnd.n1748 240.244
R11687 gnd.n5862 gnd.n1748 240.244
R11688 gnd.n5862 gnd.n1738 240.244
R11689 gnd.n5872 gnd.n1738 240.244
R11690 gnd.n5872 gnd.n1734 240.244
R11691 gnd.n5878 gnd.n1734 240.244
R11692 gnd.n5878 gnd.n1723 240.244
R11693 gnd.n5888 gnd.n1723 240.244
R11694 gnd.n5888 gnd.n1719 240.244
R11695 gnd.n5894 gnd.n1719 240.244
R11696 gnd.n5894 gnd.n1709 240.244
R11697 gnd.n5904 gnd.n1709 240.244
R11698 gnd.n5904 gnd.n1705 240.244
R11699 gnd.n5910 gnd.n1705 240.244
R11700 gnd.n5910 gnd.n1693 240.244
R11701 gnd.n5920 gnd.n1693 240.244
R11702 gnd.n5920 gnd.n1689 240.244
R11703 gnd.n5926 gnd.n1689 240.244
R11704 gnd.n5926 gnd.n1679 240.244
R11705 gnd.n5936 gnd.n1679 240.244
R11706 gnd.n5936 gnd.n1675 240.244
R11707 gnd.n5942 gnd.n1675 240.244
R11708 gnd.n5942 gnd.n1667 240.244
R11709 gnd.n5952 gnd.n1667 240.244
R11710 gnd.n5952 gnd.n1663 240.244
R11711 gnd.n5958 gnd.n1663 240.244
R11712 gnd.n5958 gnd.n1652 240.244
R11713 gnd.n5968 gnd.n1652 240.244
R11714 gnd.n5968 gnd.n1648 240.244
R11715 gnd.n5974 gnd.n1648 240.244
R11716 gnd.n5974 gnd.n1638 240.244
R11717 gnd.n5984 gnd.n1638 240.244
R11718 gnd.n5984 gnd.n1634 240.244
R11719 gnd.n5990 gnd.n1634 240.244
R11720 gnd.n5990 gnd.n1625 240.244
R11721 gnd.n6002 gnd.n1625 240.244
R11722 gnd.n6002 gnd.n1620 240.244
R11723 gnd.n6011 gnd.n1620 240.244
R11724 gnd.n6011 gnd.n1621 240.244
R11725 gnd.n1621 gnd.n1246 240.244
R11726 gnd.n6301 gnd.n1246 240.244
R11727 gnd.n6301 gnd.n1249 240.244
R11728 gnd.n6297 gnd.n1249 240.244
R11729 gnd.n6297 gnd.n1255 240.244
R11730 gnd.n1444 gnd.n1255 240.244
R11731 gnd.n1444 gnd.n1441 240.244
R11732 gnd.n1450 gnd.n1441 240.244
R11733 gnd.n1451 gnd.n1450 240.244
R11734 gnd.n6064 gnd.n1451 240.244
R11735 gnd.n6064 gnd.n1436 240.244
R11736 gnd.n6072 gnd.n1436 240.244
R11737 gnd.n6072 gnd.n1437 240.244
R11738 gnd.n1437 gnd.n1413 240.244
R11739 gnd.n6100 gnd.n1413 240.244
R11740 gnd.n6100 gnd.n1408 240.244
R11741 gnd.n6108 gnd.n1408 240.244
R11742 gnd.n6108 gnd.n1409 240.244
R11743 gnd.n1409 gnd.n1379 240.244
R11744 gnd.n6161 gnd.n1379 240.244
R11745 gnd.n6161 gnd.n1374 240.244
R11746 gnd.n6179 gnd.n1374 240.244
R11747 gnd.n6179 gnd.n1375 240.244
R11748 gnd.n6175 gnd.n1375 240.244
R11749 gnd.n6175 gnd.n6174 240.244
R11750 gnd.n6174 gnd.n6173 240.244
R11751 gnd.n6173 gnd.n409 240.244
R11752 gnd.n7363 gnd.n409 240.244
R11753 gnd.n7363 gnd.n410 240.244
R11754 gnd.n7359 gnd.n410 240.244
R11755 gnd.n7359 gnd.n7358 240.244
R11756 gnd.n7358 gnd.n7357 240.244
R11757 gnd.n7357 gnd.n416 240.244
R11758 gnd.n7353 gnd.n416 240.244
R11759 gnd.n6714 gnd.n798 240.244
R11760 gnd.n6714 gnd.n801 240.244
R11761 gnd.n6710 gnd.n801 240.244
R11762 gnd.n6710 gnd.n803 240.244
R11763 gnd.n6706 gnd.n803 240.244
R11764 gnd.n6706 gnd.n809 240.244
R11765 gnd.n6702 gnd.n809 240.244
R11766 gnd.n6702 gnd.n811 240.244
R11767 gnd.n6698 gnd.n811 240.244
R11768 gnd.n6698 gnd.n817 240.244
R11769 gnd.n6694 gnd.n817 240.244
R11770 gnd.n6694 gnd.n819 240.244
R11771 gnd.n6690 gnd.n819 240.244
R11772 gnd.n6690 gnd.n825 240.244
R11773 gnd.n6686 gnd.n825 240.244
R11774 gnd.n6686 gnd.n827 240.244
R11775 gnd.n6682 gnd.n827 240.244
R11776 gnd.n6682 gnd.n833 240.244
R11777 gnd.n6678 gnd.n833 240.244
R11778 gnd.n6678 gnd.n835 240.244
R11779 gnd.n6674 gnd.n835 240.244
R11780 gnd.n6674 gnd.n841 240.244
R11781 gnd.n6670 gnd.n841 240.244
R11782 gnd.n6670 gnd.n843 240.244
R11783 gnd.n6666 gnd.n843 240.244
R11784 gnd.n6666 gnd.n849 240.244
R11785 gnd.n6662 gnd.n849 240.244
R11786 gnd.n6662 gnd.n851 240.244
R11787 gnd.n6658 gnd.n851 240.244
R11788 gnd.n6658 gnd.n857 240.244
R11789 gnd.n6654 gnd.n857 240.244
R11790 gnd.n6654 gnd.n859 240.244
R11791 gnd.n6650 gnd.n859 240.244
R11792 gnd.n6650 gnd.n865 240.244
R11793 gnd.n6646 gnd.n865 240.244
R11794 gnd.n6646 gnd.n867 240.244
R11795 gnd.n6642 gnd.n867 240.244
R11796 gnd.n6642 gnd.n873 240.244
R11797 gnd.n6638 gnd.n873 240.244
R11798 gnd.n6638 gnd.n875 240.244
R11799 gnd.n6634 gnd.n875 240.244
R11800 gnd.n6634 gnd.n881 240.244
R11801 gnd.n6630 gnd.n881 240.244
R11802 gnd.n6630 gnd.n883 240.244
R11803 gnd.n6626 gnd.n883 240.244
R11804 gnd.n6626 gnd.n889 240.244
R11805 gnd.n6622 gnd.n889 240.244
R11806 gnd.n6622 gnd.n891 240.244
R11807 gnd.n6618 gnd.n891 240.244
R11808 gnd.n6618 gnd.n897 240.244
R11809 gnd.n6614 gnd.n897 240.244
R11810 gnd.n6614 gnd.n899 240.244
R11811 gnd.n6610 gnd.n899 240.244
R11812 gnd.n6610 gnd.n905 240.244
R11813 gnd.n6606 gnd.n905 240.244
R11814 gnd.n6606 gnd.n907 240.244
R11815 gnd.n6602 gnd.n907 240.244
R11816 gnd.n6602 gnd.n913 240.244
R11817 gnd.n6598 gnd.n913 240.244
R11818 gnd.n6598 gnd.n915 240.244
R11819 gnd.n6594 gnd.n915 240.244
R11820 gnd.n6594 gnd.n921 240.244
R11821 gnd.n6590 gnd.n921 240.244
R11822 gnd.n6590 gnd.n923 240.244
R11823 gnd.n6586 gnd.n923 240.244
R11824 gnd.n6586 gnd.n929 240.244
R11825 gnd.n6582 gnd.n929 240.244
R11826 gnd.n6582 gnd.n931 240.244
R11827 gnd.n6578 gnd.n931 240.244
R11828 gnd.n6578 gnd.n937 240.244
R11829 gnd.n6574 gnd.n937 240.244
R11830 gnd.n6574 gnd.n939 240.244
R11831 gnd.n6570 gnd.n939 240.244
R11832 gnd.n6570 gnd.n945 240.244
R11833 gnd.n6566 gnd.n945 240.244
R11834 gnd.n6566 gnd.n947 240.244
R11835 gnd.n6562 gnd.n947 240.244
R11836 gnd.n6562 gnd.n953 240.244
R11837 gnd.n6558 gnd.n953 240.244
R11838 gnd.n6558 gnd.n955 240.244
R11839 gnd.n6554 gnd.n955 240.244
R11840 gnd.n6554 gnd.n961 240.244
R11841 gnd.n6550 gnd.n961 240.244
R11842 gnd.n6550 gnd.n963 240.244
R11843 gnd.n1119 gnd.n1118 240.244
R11844 gnd.n1120 gnd.n1119 240.244
R11845 gnd.n1961 gnd.n1120 240.244
R11846 gnd.n1961 gnd.n1123 240.244
R11847 gnd.n1124 gnd.n1123 240.244
R11848 gnd.n1125 gnd.n1124 240.244
R11849 gnd.n1947 gnd.n1125 240.244
R11850 gnd.n1947 gnd.n1128 240.244
R11851 gnd.n1129 gnd.n1128 240.244
R11852 gnd.n1130 gnd.n1129 240.244
R11853 gnd.n1935 gnd.n1130 240.244
R11854 gnd.n1935 gnd.n1133 240.244
R11855 gnd.n1134 gnd.n1133 240.244
R11856 gnd.n1135 gnd.n1134 240.244
R11857 gnd.n1921 gnd.n1135 240.244
R11858 gnd.n1921 gnd.n1138 240.244
R11859 gnd.n1139 gnd.n1138 240.244
R11860 gnd.n1140 gnd.n1139 240.244
R11861 gnd.n1906 gnd.n1140 240.244
R11862 gnd.n1906 gnd.n1143 240.244
R11863 gnd.n1144 gnd.n1143 240.244
R11864 gnd.n1145 gnd.n1144 240.244
R11865 gnd.n1892 gnd.n1145 240.244
R11866 gnd.n1892 gnd.n1148 240.244
R11867 gnd.n1149 gnd.n1148 240.244
R11868 gnd.n1150 gnd.n1149 240.244
R11869 gnd.n1878 gnd.n1150 240.244
R11870 gnd.n1878 gnd.n1153 240.244
R11871 gnd.n1154 gnd.n1153 240.244
R11872 gnd.n1155 gnd.n1154 240.244
R11873 gnd.n1863 gnd.n1155 240.244
R11874 gnd.n1863 gnd.n1158 240.244
R11875 gnd.n1159 gnd.n1158 240.244
R11876 gnd.n1160 gnd.n1159 240.244
R11877 gnd.n1850 gnd.n1160 240.244
R11878 gnd.n1850 gnd.n1163 240.244
R11879 gnd.n1164 gnd.n1163 240.244
R11880 gnd.n1165 gnd.n1164 240.244
R11881 gnd.n1835 gnd.n1165 240.244
R11882 gnd.n1835 gnd.n1168 240.244
R11883 gnd.n1169 gnd.n1168 240.244
R11884 gnd.n1170 gnd.n1169 240.244
R11885 gnd.n1820 gnd.n1170 240.244
R11886 gnd.n1820 gnd.n1173 240.244
R11887 gnd.n1174 gnd.n1173 240.244
R11888 gnd.n1175 gnd.n1174 240.244
R11889 gnd.n1805 gnd.n1175 240.244
R11890 gnd.n1805 gnd.n1178 240.244
R11891 gnd.n1179 gnd.n1178 240.244
R11892 gnd.n1180 gnd.n1179 240.244
R11893 gnd.n1790 gnd.n1180 240.244
R11894 gnd.n1790 gnd.n1183 240.244
R11895 gnd.n1184 gnd.n1183 240.244
R11896 gnd.n1185 gnd.n1184 240.244
R11897 gnd.n1776 gnd.n1185 240.244
R11898 gnd.n1776 gnd.n1188 240.244
R11899 gnd.n1189 gnd.n1188 240.244
R11900 gnd.n1190 gnd.n1189 240.244
R11901 gnd.n1761 gnd.n1190 240.244
R11902 gnd.n1761 gnd.n1193 240.244
R11903 gnd.n1194 gnd.n1193 240.244
R11904 gnd.n1195 gnd.n1194 240.244
R11905 gnd.n1746 gnd.n1195 240.244
R11906 gnd.n1746 gnd.n1198 240.244
R11907 gnd.n1199 gnd.n1198 240.244
R11908 gnd.n1200 gnd.n1199 240.244
R11909 gnd.n1732 gnd.n1200 240.244
R11910 gnd.n1732 gnd.n1203 240.244
R11911 gnd.n1204 gnd.n1203 240.244
R11912 gnd.n1205 gnd.n1204 240.244
R11913 gnd.n1718 gnd.n1205 240.244
R11914 gnd.n1718 gnd.n1208 240.244
R11915 gnd.n1209 gnd.n1208 240.244
R11916 gnd.n1210 gnd.n1209 240.244
R11917 gnd.n1702 gnd.n1210 240.244
R11918 gnd.n1702 gnd.n1213 240.244
R11919 gnd.n1214 gnd.n1213 240.244
R11920 gnd.n1215 gnd.n1214 240.244
R11921 gnd.n1687 gnd.n1215 240.244
R11922 gnd.n1687 gnd.n1218 240.244
R11923 gnd.n1219 gnd.n1218 240.244
R11924 gnd.n1220 gnd.n1219 240.244
R11925 gnd.n1673 gnd.n1220 240.244
R11926 gnd.n1673 gnd.n1223 240.244
R11927 gnd.n1224 gnd.n1223 240.244
R11928 gnd.n1225 gnd.n1224 240.244
R11929 gnd.n1661 gnd.n1225 240.244
R11930 gnd.n1661 gnd.n1228 240.244
R11931 gnd.n1229 gnd.n1228 240.244
R11932 gnd.n1230 gnd.n1229 240.244
R11933 gnd.n1647 gnd.n1230 240.244
R11934 gnd.n1647 gnd.n1233 240.244
R11935 gnd.n1234 gnd.n1233 240.244
R11936 gnd.n1235 gnd.n1234 240.244
R11937 gnd.n1633 gnd.n1235 240.244
R11938 gnd.n1633 gnd.n1238 240.244
R11939 gnd.n1239 gnd.n1238 240.244
R11940 gnd.n1240 gnd.n1239 240.244
R11941 gnd.n1619 gnd.n1240 240.244
R11942 gnd.n1619 gnd.n1243 240.244
R11943 gnd.n6304 gnd.n1243 240.244
R11944 gnd.n1988 gnd.n1987 240.244
R11945 gnd.n1998 gnd.n1987 240.244
R11946 gnd.n2000 gnd.n1999 240.244
R11947 gnd.n2008 gnd.n2007 240.244
R11948 gnd.n2016 gnd.n2015 240.244
R11949 gnd.n2018 gnd.n2017 240.244
R11950 gnd.n2026 gnd.n2025 240.244
R11951 gnd.n2036 gnd.n2035 240.244
R11952 gnd.n2038 gnd.n2037 240.244
R11953 gnd.n4535 gnd.n4534 240.244
R11954 gnd.n4537 gnd.n4536 240.244
R11955 gnd.n4541 gnd.n4540 240.244
R11956 gnd.n4547 gnd.n4542 240.244
R11957 gnd.n4548 gnd.n1972 240.244
R11958 gnd.n5614 gnd.n1968 240.244
R11959 gnd.n5614 gnd.n1959 240.244
R11960 gnd.n5624 gnd.n1959 240.244
R11961 gnd.n5624 gnd.n1955 240.244
R11962 gnd.n5630 gnd.n1955 240.244
R11963 gnd.n5630 gnd.n1946 240.244
R11964 gnd.n5640 gnd.n1946 240.244
R11965 gnd.n5640 gnd.n1942 240.244
R11966 gnd.n5646 gnd.n1942 240.244
R11967 gnd.n5646 gnd.n1933 240.244
R11968 gnd.n5656 gnd.n1933 240.244
R11969 gnd.n5656 gnd.n1929 240.244
R11970 gnd.n5662 gnd.n1929 240.244
R11971 gnd.n5662 gnd.n1919 240.244
R11972 gnd.n5672 gnd.n1919 240.244
R11973 gnd.n5672 gnd.n1915 240.244
R11974 gnd.n5678 gnd.n1915 240.244
R11975 gnd.n5678 gnd.n1904 240.244
R11976 gnd.n5688 gnd.n1904 240.244
R11977 gnd.n5688 gnd.n1900 240.244
R11978 gnd.n5694 gnd.n1900 240.244
R11979 gnd.n5694 gnd.n1890 240.244
R11980 gnd.n5704 gnd.n1890 240.244
R11981 gnd.n5704 gnd.n1886 240.244
R11982 gnd.n5710 gnd.n1886 240.244
R11983 gnd.n5710 gnd.n1876 240.244
R11984 gnd.n5720 gnd.n1876 240.244
R11985 gnd.n5720 gnd.n1872 240.244
R11986 gnd.n5726 gnd.n1872 240.244
R11987 gnd.n5726 gnd.n1862 240.244
R11988 gnd.n5736 gnd.n1862 240.244
R11989 gnd.n5736 gnd.n1858 240.244
R11990 gnd.n5742 gnd.n1858 240.244
R11991 gnd.n5742 gnd.n1848 240.244
R11992 gnd.n5752 gnd.n1848 240.244
R11993 gnd.n5752 gnd.n1844 240.244
R11994 gnd.n5758 gnd.n1844 240.244
R11995 gnd.n5758 gnd.n1834 240.244
R11996 gnd.n5768 gnd.n1834 240.244
R11997 gnd.n5768 gnd.n1830 240.244
R11998 gnd.n5774 gnd.n1830 240.244
R11999 gnd.n5774 gnd.n1818 240.244
R12000 gnd.n5784 gnd.n1818 240.244
R12001 gnd.n5784 gnd.n1814 240.244
R12002 gnd.n5790 gnd.n1814 240.244
R12003 gnd.n5790 gnd.n1803 240.244
R12004 gnd.n5800 gnd.n1803 240.244
R12005 gnd.n5800 gnd.n1799 240.244
R12006 gnd.n5806 gnd.n1799 240.244
R12007 gnd.n5806 gnd.n1788 240.244
R12008 gnd.n5816 gnd.n1788 240.244
R12009 gnd.n5816 gnd.n1784 240.244
R12010 gnd.n5822 gnd.n1784 240.244
R12011 gnd.n5822 gnd.n1774 240.244
R12012 gnd.n5832 gnd.n1774 240.244
R12013 gnd.n5832 gnd.n1770 240.244
R12014 gnd.n5838 gnd.n1770 240.244
R12015 gnd.n5838 gnd.n1759 240.244
R12016 gnd.n5848 gnd.n1759 240.244
R12017 gnd.n5848 gnd.n1755 240.244
R12018 gnd.n5854 gnd.n1755 240.244
R12019 gnd.n5854 gnd.n1744 240.244
R12020 gnd.n5864 gnd.n1744 240.244
R12021 gnd.n5864 gnd.n1740 240.244
R12022 gnd.n5870 gnd.n1740 240.244
R12023 gnd.n5870 gnd.n1730 240.244
R12024 gnd.n5880 gnd.n1730 240.244
R12025 gnd.n5880 gnd.n1726 240.244
R12026 gnd.n5886 gnd.n1726 240.244
R12027 gnd.n5886 gnd.n1716 240.244
R12028 gnd.n5896 gnd.n1716 240.244
R12029 gnd.n5896 gnd.n1712 240.244
R12030 gnd.n5902 gnd.n1712 240.244
R12031 gnd.n5902 gnd.n1700 240.244
R12032 gnd.n5912 gnd.n1700 240.244
R12033 gnd.n5912 gnd.n1696 240.244
R12034 gnd.n5918 gnd.n1696 240.244
R12035 gnd.n5918 gnd.n1685 240.244
R12036 gnd.n5928 gnd.n1685 240.244
R12037 gnd.n5928 gnd.n1681 240.244
R12038 gnd.n5934 gnd.n1681 240.244
R12039 gnd.n5934 gnd.n1672 240.244
R12040 gnd.n5944 gnd.n1672 240.244
R12041 gnd.n5944 gnd.n1668 240.244
R12042 gnd.n5950 gnd.n1668 240.244
R12043 gnd.n5950 gnd.n1659 240.244
R12044 gnd.n5960 gnd.n1659 240.244
R12045 gnd.n5960 gnd.n1655 240.244
R12046 gnd.n5966 gnd.n1655 240.244
R12047 gnd.n5966 gnd.n1645 240.244
R12048 gnd.n5976 gnd.n1645 240.244
R12049 gnd.n5976 gnd.n1641 240.244
R12050 gnd.n5982 gnd.n1641 240.244
R12051 gnd.n5982 gnd.n1632 240.244
R12052 gnd.n5992 gnd.n1632 240.244
R12053 gnd.n5992 gnd.n1627 240.244
R12054 gnd.n6000 gnd.n1627 240.244
R12055 gnd.n6000 gnd.n1617 240.244
R12056 gnd.n6013 gnd.n1617 240.244
R12057 gnd.n6014 gnd.n6013 240.244
R12058 gnd.n6014 gnd.n1247 240.244
R12059 gnd.n1532 gnd.n1531 240.244
R12060 gnd.n1535 gnd.n1534 240.244
R12061 gnd.n1551 gnd.n1550 240.244
R12062 gnd.n1554 gnd.n1553 240.244
R12063 gnd.n1570 gnd.n1569 240.244
R12064 gnd.n1573 gnd.n1572 240.244
R12065 gnd.n1586 gnd.n1585 240.244
R12066 gnd.n1589 gnd.n1588 240.244
R12067 gnd.n1600 gnd.n1599 240.244
R12068 gnd.n1603 gnd.n1602 240.244
R12069 gnd.n1608 gnd.n1605 240.244
R12070 gnd.n1611 gnd.n1610 240.244
R12071 gnd.n6019 gnd.n1613 240.244
R12072 gnd.n6022 gnd.n6021 240.244
R12073 gnd.n4662 gnd.n4661 240.132
R12074 gnd.n5017 gnd.n5016 240.132
R12075 gnd.n6722 gnd.n6721 225.874
R12076 gnd.n6723 gnd.n6722 225.874
R12077 gnd.n6723 gnd.n791 225.874
R12078 gnd.n6731 gnd.n791 225.874
R12079 gnd.n6732 gnd.n6731 225.874
R12080 gnd.n6733 gnd.n6732 225.874
R12081 gnd.n6733 gnd.n785 225.874
R12082 gnd.n6741 gnd.n785 225.874
R12083 gnd.n6742 gnd.n6741 225.874
R12084 gnd.n6743 gnd.n6742 225.874
R12085 gnd.n6743 gnd.n779 225.874
R12086 gnd.n6751 gnd.n779 225.874
R12087 gnd.n6752 gnd.n6751 225.874
R12088 gnd.n6753 gnd.n6752 225.874
R12089 gnd.n6753 gnd.n773 225.874
R12090 gnd.n6761 gnd.n773 225.874
R12091 gnd.n6762 gnd.n6761 225.874
R12092 gnd.n6763 gnd.n6762 225.874
R12093 gnd.n6763 gnd.n767 225.874
R12094 gnd.n6771 gnd.n767 225.874
R12095 gnd.n6772 gnd.n6771 225.874
R12096 gnd.n6773 gnd.n6772 225.874
R12097 gnd.n6773 gnd.n761 225.874
R12098 gnd.n6781 gnd.n761 225.874
R12099 gnd.n6782 gnd.n6781 225.874
R12100 gnd.n6783 gnd.n6782 225.874
R12101 gnd.n6783 gnd.n755 225.874
R12102 gnd.n6791 gnd.n755 225.874
R12103 gnd.n6792 gnd.n6791 225.874
R12104 gnd.n6793 gnd.n6792 225.874
R12105 gnd.n6793 gnd.n749 225.874
R12106 gnd.n6801 gnd.n749 225.874
R12107 gnd.n6802 gnd.n6801 225.874
R12108 gnd.n6803 gnd.n6802 225.874
R12109 gnd.n6803 gnd.n743 225.874
R12110 gnd.n6811 gnd.n743 225.874
R12111 gnd.n6812 gnd.n6811 225.874
R12112 gnd.n6813 gnd.n6812 225.874
R12113 gnd.n6813 gnd.n737 225.874
R12114 gnd.n6821 gnd.n737 225.874
R12115 gnd.n6822 gnd.n6821 225.874
R12116 gnd.n6823 gnd.n6822 225.874
R12117 gnd.n6823 gnd.n731 225.874
R12118 gnd.n6831 gnd.n731 225.874
R12119 gnd.n6832 gnd.n6831 225.874
R12120 gnd.n6833 gnd.n6832 225.874
R12121 gnd.n6833 gnd.n725 225.874
R12122 gnd.n6841 gnd.n725 225.874
R12123 gnd.n6842 gnd.n6841 225.874
R12124 gnd.n6843 gnd.n6842 225.874
R12125 gnd.n6843 gnd.n719 225.874
R12126 gnd.n6851 gnd.n719 225.874
R12127 gnd.n6852 gnd.n6851 225.874
R12128 gnd.n6853 gnd.n6852 225.874
R12129 gnd.n6853 gnd.n713 225.874
R12130 gnd.n6861 gnd.n713 225.874
R12131 gnd.n6862 gnd.n6861 225.874
R12132 gnd.n6863 gnd.n6862 225.874
R12133 gnd.n6863 gnd.n707 225.874
R12134 gnd.n6871 gnd.n707 225.874
R12135 gnd.n6872 gnd.n6871 225.874
R12136 gnd.n6873 gnd.n6872 225.874
R12137 gnd.n6873 gnd.n701 225.874
R12138 gnd.n6881 gnd.n701 225.874
R12139 gnd.n6882 gnd.n6881 225.874
R12140 gnd.n6883 gnd.n6882 225.874
R12141 gnd.n6883 gnd.n695 225.874
R12142 gnd.n6891 gnd.n695 225.874
R12143 gnd.n6892 gnd.n6891 225.874
R12144 gnd.n6893 gnd.n6892 225.874
R12145 gnd.n6893 gnd.n689 225.874
R12146 gnd.n6901 gnd.n689 225.874
R12147 gnd.n6902 gnd.n6901 225.874
R12148 gnd.n6903 gnd.n6902 225.874
R12149 gnd.n6903 gnd.n683 225.874
R12150 gnd.n6911 gnd.n683 225.874
R12151 gnd.n6912 gnd.n6911 225.874
R12152 gnd.n6913 gnd.n6912 225.874
R12153 gnd.n6913 gnd.n677 225.874
R12154 gnd.n6921 gnd.n677 225.874
R12155 gnd.n6922 gnd.n6921 225.874
R12156 gnd.n6923 gnd.n6922 225.874
R12157 gnd.n6923 gnd.n671 225.874
R12158 gnd.n6931 gnd.n671 225.874
R12159 gnd.n6932 gnd.n6931 225.874
R12160 gnd.n6933 gnd.n6932 225.874
R12161 gnd.n6933 gnd.n665 225.874
R12162 gnd.n6941 gnd.n665 225.874
R12163 gnd.n6942 gnd.n6941 225.874
R12164 gnd.n6943 gnd.n6942 225.874
R12165 gnd.n6943 gnd.n659 225.874
R12166 gnd.n6951 gnd.n659 225.874
R12167 gnd.n6952 gnd.n6951 225.874
R12168 gnd.n6953 gnd.n6952 225.874
R12169 gnd.n6953 gnd.n653 225.874
R12170 gnd.n6961 gnd.n653 225.874
R12171 gnd.n6962 gnd.n6961 225.874
R12172 gnd.n6963 gnd.n6962 225.874
R12173 gnd.n6963 gnd.n647 225.874
R12174 gnd.n6971 gnd.n647 225.874
R12175 gnd.n6972 gnd.n6971 225.874
R12176 gnd.n6973 gnd.n6972 225.874
R12177 gnd.n6973 gnd.n641 225.874
R12178 gnd.n6981 gnd.n641 225.874
R12179 gnd.n6982 gnd.n6981 225.874
R12180 gnd.n6983 gnd.n6982 225.874
R12181 gnd.n6983 gnd.n635 225.874
R12182 gnd.n6991 gnd.n635 225.874
R12183 gnd.n6992 gnd.n6991 225.874
R12184 gnd.n6993 gnd.n6992 225.874
R12185 gnd.n6993 gnd.n629 225.874
R12186 gnd.n7001 gnd.n629 225.874
R12187 gnd.n7002 gnd.n7001 225.874
R12188 gnd.n7003 gnd.n7002 225.874
R12189 gnd.n7003 gnd.n623 225.874
R12190 gnd.n7011 gnd.n623 225.874
R12191 gnd.n7012 gnd.n7011 225.874
R12192 gnd.n7013 gnd.n7012 225.874
R12193 gnd.n7013 gnd.n617 225.874
R12194 gnd.n7021 gnd.n617 225.874
R12195 gnd.n7022 gnd.n7021 225.874
R12196 gnd.n7023 gnd.n7022 225.874
R12197 gnd.n7023 gnd.n611 225.874
R12198 gnd.n7031 gnd.n611 225.874
R12199 gnd.n7032 gnd.n7031 225.874
R12200 gnd.n7033 gnd.n7032 225.874
R12201 gnd.n7033 gnd.n605 225.874
R12202 gnd.n7041 gnd.n605 225.874
R12203 gnd.n7042 gnd.n7041 225.874
R12204 gnd.n7043 gnd.n7042 225.874
R12205 gnd.n7043 gnd.n599 225.874
R12206 gnd.n7051 gnd.n599 225.874
R12207 gnd.n7052 gnd.n7051 225.874
R12208 gnd.n7053 gnd.n7052 225.874
R12209 gnd.n7053 gnd.n593 225.874
R12210 gnd.n7061 gnd.n593 225.874
R12211 gnd.n7062 gnd.n7061 225.874
R12212 gnd.n7063 gnd.n7062 225.874
R12213 gnd.n7063 gnd.n587 225.874
R12214 gnd.n7071 gnd.n587 225.874
R12215 gnd.n7072 gnd.n7071 225.874
R12216 gnd.n7073 gnd.n7072 225.874
R12217 gnd.n7073 gnd.n581 225.874
R12218 gnd.n7081 gnd.n581 225.874
R12219 gnd.n7082 gnd.n7081 225.874
R12220 gnd.n7083 gnd.n7082 225.874
R12221 gnd.n7083 gnd.n575 225.874
R12222 gnd.n7091 gnd.n575 225.874
R12223 gnd.n7092 gnd.n7091 225.874
R12224 gnd.n7093 gnd.n7092 225.874
R12225 gnd.n7093 gnd.n569 225.874
R12226 gnd.n7101 gnd.n569 225.874
R12227 gnd.n7102 gnd.n7101 225.874
R12228 gnd.n7103 gnd.n7102 225.874
R12229 gnd.n7103 gnd.n563 225.874
R12230 gnd.n7111 gnd.n563 225.874
R12231 gnd.n7112 gnd.n7111 225.874
R12232 gnd.n7113 gnd.n7112 225.874
R12233 gnd.n7113 gnd.n557 225.874
R12234 gnd.n7121 gnd.n557 225.874
R12235 gnd.n7122 gnd.n7121 225.874
R12236 gnd.n7123 gnd.n7122 225.874
R12237 gnd.n7123 gnd.n551 225.874
R12238 gnd.n7132 gnd.n551 225.874
R12239 gnd.n7133 gnd.n7132 225.874
R12240 gnd.n7134 gnd.n7133 225.874
R12241 gnd.n7134 gnd.n546 225.874
R12242 gnd.n2901 gnd.t277 224.174
R12243 gnd.n2398 gnd.t254 224.174
R12244 gnd.n1306 gnd.n1263 199.319
R12245 gnd.n1306 gnd.n1264 199.319
R12246 gnd.n2100 gnd.n2070 199.319
R12247 gnd.n2100 gnd.n2069 199.319
R12248 gnd.n4663 gnd.n4660 186.49
R12249 gnd.n5018 gnd.n5015 186.49
R12250 gnd.n3676 gnd.n3675 185
R12251 gnd.n3674 gnd.n3673 185
R12252 gnd.n3653 gnd.n3652 185
R12253 gnd.n3668 gnd.n3667 185
R12254 gnd.n3666 gnd.n3665 185
R12255 gnd.n3657 gnd.n3656 185
R12256 gnd.n3660 gnd.n3659 185
R12257 gnd.n3644 gnd.n3643 185
R12258 gnd.n3642 gnd.n3641 185
R12259 gnd.n3621 gnd.n3620 185
R12260 gnd.n3636 gnd.n3635 185
R12261 gnd.n3634 gnd.n3633 185
R12262 gnd.n3625 gnd.n3624 185
R12263 gnd.n3628 gnd.n3627 185
R12264 gnd.n3612 gnd.n3611 185
R12265 gnd.n3610 gnd.n3609 185
R12266 gnd.n3589 gnd.n3588 185
R12267 gnd.n3604 gnd.n3603 185
R12268 gnd.n3602 gnd.n3601 185
R12269 gnd.n3593 gnd.n3592 185
R12270 gnd.n3596 gnd.n3595 185
R12271 gnd.n3581 gnd.n3580 185
R12272 gnd.n3579 gnd.n3578 185
R12273 gnd.n3558 gnd.n3557 185
R12274 gnd.n3573 gnd.n3572 185
R12275 gnd.n3571 gnd.n3570 185
R12276 gnd.n3562 gnd.n3561 185
R12277 gnd.n3565 gnd.n3564 185
R12278 gnd.n3549 gnd.n3548 185
R12279 gnd.n3547 gnd.n3546 185
R12280 gnd.n3526 gnd.n3525 185
R12281 gnd.n3541 gnd.n3540 185
R12282 gnd.n3539 gnd.n3538 185
R12283 gnd.n3530 gnd.n3529 185
R12284 gnd.n3533 gnd.n3532 185
R12285 gnd.n3517 gnd.n3516 185
R12286 gnd.n3515 gnd.n3514 185
R12287 gnd.n3494 gnd.n3493 185
R12288 gnd.n3509 gnd.n3508 185
R12289 gnd.n3507 gnd.n3506 185
R12290 gnd.n3498 gnd.n3497 185
R12291 gnd.n3501 gnd.n3500 185
R12292 gnd.n3485 gnd.n3484 185
R12293 gnd.n3483 gnd.n3482 185
R12294 gnd.n3462 gnd.n3461 185
R12295 gnd.n3477 gnd.n3476 185
R12296 gnd.n3475 gnd.n3474 185
R12297 gnd.n3466 gnd.n3465 185
R12298 gnd.n3469 gnd.n3468 185
R12299 gnd.n3454 gnd.n3453 185
R12300 gnd.n3452 gnd.n3451 185
R12301 gnd.n3431 gnd.n3430 185
R12302 gnd.n3446 gnd.n3445 185
R12303 gnd.n3444 gnd.n3443 185
R12304 gnd.n3435 gnd.n3434 185
R12305 gnd.n3438 gnd.n3437 185
R12306 gnd.n2902 gnd.t276 178.987
R12307 gnd.n2399 gnd.t255 178.987
R12308 gnd.n1 gnd.t312 170.774
R12309 gnd.n9 gnd.t61 170.103
R12310 gnd.n8 gnd.t357 170.103
R12311 gnd.n7 gnd.t27 170.103
R12312 gnd.n6 gnd.t159 170.103
R12313 gnd.n5 gnd.t31 170.103
R12314 gnd.n4 gnd.t359 170.103
R12315 gnd.n3 gnd.t130 170.103
R12316 gnd.n2 gnd.t85 170.103
R12317 gnd.n1 gnd.t350 170.103
R12318 gnd.n5190 gnd.n5189 163.367
R12319 gnd.n5187 gnd.n5027 163.367
R12320 gnd.n5183 gnd.n5182 163.367
R12321 gnd.n5180 gnd.n5030 163.367
R12322 gnd.n5176 gnd.n5175 163.367
R12323 gnd.n5173 gnd.n5033 163.367
R12324 gnd.n5169 gnd.n5168 163.367
R12325 gnd.n5166 gnd.n5036 163.367
R12326 gnd.n5162 gnd.n5161 163.367
R12327 gnd.n5159 gnd.n5039 163.367
R12328 gnd.n5155 gnd.n5154 163.367
R12329 gnd.n5152 gnd.n5042 163.367
R12330 gnd.n5148 gnd.n5147 163.367
R12331 gnd.n5145 gnd.n5045 163.367
R12332 gnd.n5140 gnd.n5139 163.367
R12333 gnd.n5137 gnd.n5135 163.367
R12334 gnd.n5132 gnd.n5131 163.367
R12335 gnd.n5129 gnd.n5051 163.367
R12336 gnd.n5124 gnd.n5123 163.367
R12337 gnd.n5121 gnd.n5056 163.367
R12338 gnd.n5117 gnd.n5116 163.367
R12339 gnd.n5114 gnd.n5059 163.367
R12340 gnd.n5110 gnd.n5109 163.367
R12341 gnd.n5107 gnd.n5062 163.367
R12342 gnd.n5103 gnd.n5102 163.367
R12343 gnd.n5100 gnd.n5065 163.367
R12344 gnd.n5096 gnd.n5095 163.367
R12345 gnd.n5093 gnd.n5068 163.367
R12346 gnd.n5089 gnd.n5088 163.367
R12347 gnd.n5086 gnd.n5071 163.367
R12348 gnd.n5082 gnd.n5081 163.367
R12349 gnd.n5079 gnd.n5075 163.367
R12350 gnd.n5451 gnd.n4678 163.367
R12351 gnd.n5451 gnd.n4679 163.367
R12352 gnd.n5447 gnd.n4679 163.367
R12353 gnd.n5447 gnd.n5446 163.367
R12354 gnd.n5446 gnd.n4747 163.367
R12355 gnd.n4754 gnd.n4747 163.367
R12356 gnd.n5436 gnd.n4754 163.367
R12357 gnd.n5436 gnd.n4755 163.367
R12358 gnd.n5432 gnd.n4755 163.367
R12359 gnd.n5432 gnd.n5431 163.367
R12360 gnd.n5431 gnd.n4759 163.367
R12361 gnd.n4767 gnd.n4759 163.367
R12362 gnd.n5421 gnd.n4767 163.367
R12363 gnd.n5421 gnd.n4768 163.367
R12364 gnd.n5417 gnd.n4768 163.367
R12365 gnd.n5417 gnd.n5416 163.367
R12366 gnd.n5416 gnd.n4772 163.367
R12367 gnd.n4781 gnd.n4772 163.367
R12368 gnd.n5406 gnd.n4781 163.367
R12369 gnd.n5406 gnd.n4782 163.367
R12370 gnd.n5402 gnd.n4782 163.367
R12371 gnd.n5402 gnd.n5401 163.367
R12372 gnd.n5401 gnd.n4786 163.367
R12373 gnd.n4799 gnd.n4786 163.367
R12374 gnd.n4799 gnd.n4796 163.367
R12375 gnd.n5391 gnd.n4796 163.367
R12376 gnd.n5391 gnd.n4797 163.367
R12377 gnd.n5387 gnd.n4797 163.367
R12378 gnd.n5387 gnd.n4803 163.367
R12379 gnd.n4811 gnd.n4803 163.367
R12380 gnd.n5377 gnd.n4811 163.367
R12381 gnd.n5377 gnd.n4812 163.367
R12382 gnd.n5373 gnd.n4812 163.367
R12383 gnd.n5373 gnd.n5372 163.367
R12384 gnd.n5372 gnd.n4815 163.367
R12385 gnd.n4828 gnd.n4815 163.367
R12386 gnd.n4828 gnd.n4825 163.367
R12387 gnd.n5362 gnd.n4825 163.367
R12388 gnd.n5362 gnd.n4826 163.367
R12389 gnd.n5358 gnd.n4826 163.367
R12390 gnd.n5358 gnd.n4832 163.367
R12391 gnd.n4847 gnd.n4832 163.367
R12392 gnd.n4847 gnd.n4846 163.367
R12393 gnd.n4851 gnd.n4846 163.367
R12394 gnd.n4854 gnd.n4851 163.367
R12395 gnd.n4855 gnd.n4854 163.367
R12396 gnd.n4855 gnd.n4843 163.367
R12397 gnd.n5341 gnd.n4843 163.367
R12398 gnd.n5341 gnd.n4844 163.367
R12399 gnd.n5337 gnd.n4844 163.367
R12400 gnd.n5337 gnd.n5336 163.367
R12401 gnd.n5336 gnd.n4859 163.367
R12402 gnd.n4867 gnd.n4859 163.367
R12403 gnd.n5326 gnd.n4867 163.367
R12404 gnd.n5326 gnd.n4868 163.367
R12405 gnd.n5322 gnd.n4868 163.367
R12406 gnd.n5322 gnd.n5321 163.367
R12407 gnd.n5321 gnd.n4872 163.367
R12408 gnd.n4881 gnd.n4872 163.367
R12409 gnd.n5311 gnd.n4881 163.367
R12410 gnd.n5311 gnd.n4882 163.367
R12411 gnd.n5307 gnd.n4882 163.367
R12412 gnd.n5307 gnd.n5306 163.367
R12413 gnd.n5306 gnd.n4886 163.367
R12414 gnd.n4894 gnd.n4886 163.367
R12415 gnd.n5296 gnd.n4894 163.367
R12416 gnd.n5296 gnd.n4895 163.367
R12417 gnd.n5292 gnd.n4895 163.367
R12418 gnd.n5292 gnd.n5291 163.367
R12419 gnd.n5291 gnd.n4899 163.367
R12420 gnd.n4908 gnd.n4899 163.367
R12421 gnd.n5282 gnd.n4908 163.367
R12422 gnd.n5282 gnd.n4909 163.367
R12423 gnd.n5278 gnd.n4909 163.367
R12424 gnd.n5278 gnd.n5277 163.367
R12425 gnd.n5277 gnd.n4913 163.367
R12426 gnd.n4921 gnd.n4913 163.367
R12427 gnd.n5267 gnd.n4921 163.367
R12428 gnd.n5267 gnd.n4922 163.367
R12429 gnd.n5263 gnd.n4922 163.367
R12430 gnd.n5263 gnd.n5262 163.367
R12431 gnd.n5262 gnd.n4926 163.367
R12432 gnd.n4936 gnd.n4926 163.367
R12433 gnd.n5253 gnd.n4936 163.367
R12434 gnd.n5253 gnd.n4937 163.367
R12435 gnd.n5249 gnd.n4937 163.367
R12436 gnd.n5249 gnd.n4941 163.367
R12437 gnd.n4952 gnd.n4941 163.367
R12438 gnd.n4952 gnd.n4950 163.367
R12439 gnd.n5239 gnd.n4950 163.367
R12440 gnd.n5239 gnd.n4951 163.367
R12441 gnd.n5235 gnd.n4951 163.367
R12442 gnd.n5235 gnd.n5234 163.367
R12443 gnd.n5234 gnd.n5233 163.367
R12444 gnd.n5233 gnd.n4956 163.367
R12445 gnd.n5229 gnd.n4956 163.367
R12446 gnd.n5229 gnd.n5228 163.367
R12447 gnd.n5228 gnd.n5227 163.367
R12448 gnd.n5227 gnd.n4958 163.367
R12449 gnd.n4983 gnd.n4958 163.367
R12450 gnd.n4983 gnd.n4980 163.367
R12451 gnd.n5216 gnd.n4980 163.367
R12452 gnd.n5216 gnd.n4981 163.367
R12453 gnd.n5212 gnd.n4981 163.367
R12454 gnd.n5212 gnd.n4987 163.367
R12455 gnd.n4996 gnd.n4987 163.367
R12456 gnd.n5202 gnd.n4996 163.367
R12457 gnd.n5202 gnd.n4997 163.367
R12458 gnd.n5198 gnd.n4997 163.367
R12459 gnd.n5198 gnd.n5197 163.367
R12460 gnd.n4654 gnd.n4653 163.367
R12461 gnd.n5516 gnd.n4653 163.367
R12462 gnd.n5514 gnd.n5513 163.367
R12463 gnd.n5510 gnd.n5509 163.367
R12464 gnd.n5506 gnd.n5505 163.367
R12465 gnd.n5502 gnd.n5501 163.367
R12466 gnd.n5498 gnd.n5497 163.367
R12467 gnd.n5494 gnd.n5493 163.367
R12468 gnd.n5490 gnd.n5489 163.367
R12469 gnd.n5486 gnd.n5485 163.367
R12470 gnd.n5482 gnd.n5481 163.367
R12471 gnd.n5478 gnd.n5477 163.367
R12472 gnd.n5474 gnd.n5473 163.367
R12473 gnd.n5470 gnd.n5469 163.367
R12474 gnd.n5466 gnd.n5465 163.367
R12475 gnd.n5462 gnd.n5461 163.367
R12476 gnd.n5525 gnd.n4620 163.367
R12477 gnd.n4684 gnd.n4683 163.367
R12478 gnd.n4689 gnd.n4688 163.367
R12479 gnd.n4693 gnd.n4692 163.367
R12480 gnd.n4697 gnd.n4696 163.367
R12481 gnd.n4701 gnd.n4700 163.367
R12482 gnd.n4705 gnd.n4704 163.367
R12483 gnd.n4709 gnd.n4708 163.367
R12484 gnd.n4713 gnd.n4712 163.367
R12485 gnd.n4717 gnd.n4716 163.367
R12486 gnd.n4721 gnd.n4720 163.367
R12487 gnd.n4725 gnd.n4724 163.367
R12488 gnd.n4729 gnd.n4728 163.367
R12489 gnd.n4733 gnd.n4732 163.367
R12490 gnd.n4737 gnd.n4736 163.367
R12491 gnd.n4741 gnd.n4740 163.367
R12492 gnd.n5454 gnd.n4655 163.367
R12493 gnd.n5454 gnd.n4677 163.367
R12494 gnd.n4749 gnd.n4677 163.367
R12495 gnd.n5444 gnd.n4749 163.367
R12496 gnd.n5444 gnd.n4750 163.367
R12497 gnd.n5440 gnd.n4750 163.367
R12498 gnd.n5440 gnd.n5439 163.367
R12499 gnd.n5439 gnd.n4753 163.367
R12500 gnd.n4761 gnd.n4753 163.367
R12501 gnd.n5429 gnd.n4761 163.367
R12502 gnd.n5429 gnd.n4762 163.367
R12503 gnd.n5425 gnd.n4762 163.367
R12504 gnd.n5425 gnd.n4766 163.367
R12505 gnd.n4776 gnd.n4766 163.367
R12506 gnd.n4776 gnd.n4774 163.367
R12507 gnd.n5414 gnd.n4774 163.367
R12508 gnd.n5414 gnd.n4775 163.367
R12509 gnd.n5410 gnd.n4775 163.367
R12510 gnd.n5410 gnd.n4780 163.367
R12511 gnd.n4790 gnd.n4780 163.367
R12512 gnd.n4790 gnd.n4788 163.367
R12513 gnd.n5399 gnd.n4788 163.367
R12514 gnd.n5399 gnd.n4789 163.367
R12515 gnd.n5395 gnd.n4789 163.367
R12516 gnd.n5395 gnd.n5394 163.367
R12517 gnd.n5394 gnd.n4794 163.367
R12518 gnd.n4805 gnd.n4794 163.367
R12519 gnd.n5385 gnd.n4805 163.367
R12520 gnd.n5385 gnd.n4806 163.367
R12521 gnd.n5381 gnd.n4806 163.367
R12522 gnd.n5381 gnd.n4810 163.367
R12523 gnd.n4819 gnd.n4810 163.367
R12524 gnd.n4819 gnd.n4817 163.367
R12525 gnd.n5370 gnd.n4817 163.367
R12526 gnd.n5370 gnd.n4818 163.367
R12527 gnd.n5366 gnd.n4818 163.367
R12528 gnd.n5366 gnd.n5365 163.367
R12529 gnd.n5365 gnd.n4823 163.367
R12530 gnd.n4834 gnd.n4823 163.367
R12531 gnd.n5356 gnd.n4834 163.367
R12532 gnd.n5356 gnd.n4835 163.367
R12533 gnd.n5352 gnd.n4835 163.367
R12534 gnd.n5352 gnd.n5351 163.367
R12535 gnd.n5351 gnd.n5350 163.367
R12536 gnd.n5350 gnd.n4839 163.367
R12537 gnd.n5346 gnd.n4839 163.367
R12538 gnd.n5346 gnd.n5345 163.367
R12539 gnd.n5345 gnd.n5344 163.367
R12540 gnd.n5344 gnd.n4841 163.367
R12541 gnd.n4861 gnd.n4841 163.367
R12542 gnd.n5334 gnd.n4861 163.367
R12543 gnd.n5334 gnd.n4862 163.367
R12544 gnd.n5330 gnd.n4862 163.367
R12545 gnd.n5330 gnd.n5329 163.367
R12546 gnd.n5329 gnd.n4866 163.367
R12547 gnd.n4874 gnd.n4866 163.367
R12548 gnd.n5319 gnd.n4874 163.367
R12549 gnd.n5319 gnd.n4876 163.367
R12550 gnd.n5315 gnd.n4876 163.367
R12551 gnd.n5315 gnd.n5314 163.367
R12552 gnd.n5314 gnd.n4880 163.367
R12553 gnd.n4888 gnd.n4880 163.367
R12554 gnd.n5304 gnd.n4888 163.367
R12555 gnd.n5304 gnd.n4889 163.367
R12556 gnd.n5300 gnd.n4889 163.367
R12557 gnd.n5300 gnd.n5299 163.367
R12558 gnd.n5299 gnd.n4893 163.367
R12559 gnd.n4901 gnd.n4893 163.367
R12560 gnd.n5289 gnd.n4901 163.367
R12561 gnd.n5289 gnd.n4902 163.367
R12562 gnd.n5285 gnd.n4902 163.367
R12563 gnd.n5285 gnd.n5284 163.367
R12564 gnd.n5284 gnd.n4906 163.367
R12565 gnd.n4915 gnd.n4906 163.367
R12566 gnd.n5275 gnd.n4915 163.367
R12567 gnd.n5275 gnd.n4916 163.367
R12568 gnd.n5271 gnd.n4916 163.367
R12569 gnd.n5271 gnd.n4920 163.367
R12570 gnd.n4930 gnd.n4920 163.367
R12571 gnd.n4930 gnd.n4928 163.367
R12572 gnd.n5260 gnd.n4928 163.367
R12573 gnd.n5260 gnd.n4929 163.367
R12574 gnd.n5256 gnd.n4929 163.367
R12575 gnd.n5256 gnd.n5255 163.367
R12576 gnd.n5255 gnd.n4934 163.367
R12577 gnd.n5247 gnd.n4934 163.367
R12578 gnd.n5247 gnd.n4944 163.367
R12579 gnd.n5243 gnd.n4944 163.367
R12580 gnd.n5243 gnd.n5242 163.367
R12581 gnd.n5242 gnd.n5241 163.367
R12582 gnd.n5241 gnd.n4947 163.367
R12583 gnd.n4967 gnd.n4947 163.367
R12584 gnd.n4967 gnd.n4965 163.367
R12585 gnd.n4971 gnd.n4965 163.367
R12586 gnd.n4974 gnd.n4971 163.367
R12587 gnd.n4975 gnd.n4974 163.367
R12588 gnd.n4975 gnd.n4960 163.367
R12589 gnd.n5225 gnd.n4960 163.367
R12590 gnd.n5225 gnd.n4963 163.367
R12591 gnd.n5221 gnd.n4963 163.367
R12592 gnd.n5221 gnd.n5220 163.367
R12593 gnd.n5220 gnd.n4979 163.367
R12594 gnd.n4989 gnd.n4979 163.367
R12595 gnd.n5210 gnd.n4989 163.367
R12596 gnd.n5210 gnd.n4991 163.367
R12597 gnd.n5206 gnd.n4991 163.367
R12598 gnd.n5206 gnd.n4995 163.367
R12599 gnd.n5003 gnd.n4995 163.367
R12600 gnd.n5003 gnd.n5001 163.367
R12601 gnd.n5195 gnd.n5001 163.367
R12602 gnd.n5024 gnd.n5023 156.462
R12603 gnd.n3616 gnd.n3584 153.042
R12604 gnd.n3680 gnd.n3679 152.079
R12605 gnd.n3648 gnd.n3647 152.079
R12606 gnd.n3616 gnd.n3615 152.079
R12607 gnd.n4668 gnd.n4667 152
R12608 gnd.n4669 gnd.n4658 152
R12609 gnd.n4671 gnd.n4670 152
R12610 gnd.n4673 gnd.n4656 152
R12611 gnd.n4675 gnd.n4674 152
R12612 gnd.n5022 gnd.n5006 152
R12613 gnd.n5014 gnd.n5007 152
R12614 gnd.n5013 gnd.n5012 152
R12615 gnd.n5011 gnd.n5008 152
R12616 gnd.n5009 gnd.t265 150.546
R12617 gnd.t126 gnd.n3658 147.661
R12618 gnd.t95 gnd.n3626 147.661
R12619 gnd.t25 gnd.n3594 147.661
R12620 gnd.t163 gnd.n3563 147.661
R12621 gnd.t320 gnd.n3531 147.661
R12622 gnd.t17 gnd.n3499 147.661
R12623 gnd.t167 gnd.n3467 147.661
R12624 gnd.t180 gnd.n3436 147.661
R12625 gnd.n5134 gnd.n5133 143.351
R12626 gnd.n4635 gnd.n4619 143.351
R12627 gnd.n5524 gnd.n4619 143.351
R12628 gnd.n4665 gnd.t209 130.484
R12629 gnd.n4674 gnd.t262 126.766
R12630 gnd.n4672 gnd.t206 126.766
R12631 gnd.n4658 gnd.t227 126.766
R12632 gnd.n4666 gnd.t288 126.766
R12633 gnd.n5010 gnd.t259 126.766
R12634 gnd.n5012 gnd.t199 126.766
R12635 gnd.n5021 gnd.t238 126.766
R12636 gnd.n5023 gnd.t220 126.766
R12637 gnd.n6262 gnd.n1305 104.897
R12638 gnd.n5527 gnd.n5526 104.897
R12639 gnd.n3675 gnd.n3674 104.615
R12640 gnd.n3674 gnd.n3652 104.615
R12641 gnd.n3667 gnd.n3652 104.615
R12642 gnd.n3667 gnd.n3666 104.615
R12643 gnd.n3666 gnd.n3656 104.615
R12644 gnd.n3659 gnd.n3656 104.615
R12645 gnd.n3643 gnd.n3642 104.615
R12646 gnd.n3642 gnd.n3620 104.615
R12647 gnd.n3635 gnd.n3620 104.615
R12648 gnd.n3635 gnd.n3634 104.615
R12649 gnd.n3634 gnd.n3624 104.615
R12650 gnd.n3627 gnd.n3624 104.615
R12651 gnd.n3611 gnd.n3610 104.615
R12652 gnd.n3610 gnd.n3588 104.615
R12653 gnd.n3603 gnd.n3588 104.615
R12654 gnd.n3603 gnd.n3602 104.615
R12655 gnd.n3602 gnd.n3592 104.615
R12656 gnd.n3595 gnd.n3592 104.615
R12657 gnd.n3580 gnd.n3579 104.615
R12658 gnd.n3579 gnd.n3557 104.615
R12659 gnd.n3572 gnd.n3557 104.615
R12660 gnd.n3572 gnd.n3571 104.615
R12661 gnd.n3571 gnd.n3561 104.615
R12662 gnd.n3564 gnd.n3561 104.615
R12663 gnd.n3548 gnd.n3547 104.615
R12664 gnd.n3547 gnd.n3525 104.615
R12665 gnd.n3540 gnd.n3525 104.615
R12666 gnd.n3540 gnd.n3539 104.615
R12667 gnd.n3539 gnd.n3529 104.615
R12668 gnd.n3532 gnd.n3529 104.615
R12669 gnd.n3516 gnd.n3515 104.615
R12670 gnd.n3515 gnd.n3493 104.615
R12671 gnd.n3508 gnd.n3493 104.615
R12672 gnd.n3508 gnd.n3507 104.615
R12673 gnd.n3507 gnd.n3497 104.615
R12674 gnd.n3500 gnd.n3497 104.615
R12675 gnd.n3484 gnd.n3483 104.615
R12676 gnd.n3483 gnd.n3461 104.615
R12677 gnd.n3476 gnd.n3461 104.615
R12678 gnd.n3476 gnd.n3475 104.615
R12679 gnd.n3475 gnd.n3465 104.615
R12680 gnd.n3468 gnd.n3465 104.615
R12681 gnd.n3453 gnd.n3452 104.615
R12682 gnd.n3452 gnd.n3430 104.615
R12683 gnd.n3445 gnd.n3430 104.615
R12684 gnd.n3445 gnd.n3444 104.615
R12685 gnd.n3444 gnd.n3434 104.615
R12686 gnd.n3437 gnd.n3434 104.615
R12687 gnd.n2827 gnd.t306 100.632
R12688 gnd.n2372 gnd.t246 100.632
R12689 gnd.n7796 gnd.n138 99.6594
R12690 gnd.n7794 gnd.n7793 99.6594
R12691 gnd.n7789 gnd.n145 99.6594
R12692 gnd.n7787 gnd.n7786 99.6594
R12693 gnd.n7782 gnd.n152 99.6594
R12694 gnd.n7780 gnd.n7779 99.6594
R12695 gnd.n7775 gnd.n159 99.6594
R12696 gnd.n7773 gnd.n7772 99.6594
R12697 gnd.n7765 gnd.n166 99.6594
R12698 gnd.n7763 gnd.n7762 99.6594
R12699 gnd.n7758 gnd.n173 99.6594
R12700 gnd.n7756 gnd.n7755 99.6594
R12701 gnd.n7751 gnd.n180 99.6594
R12702 gnd.n7749 gnd.n7748 99.6594
R12703 gnd.n7744 gnd.n187 99.6594
R12704 gnd.n7742 gnd.n7741 99.6594
R12705 gnd.n7737 gnd.n194 99.6594
R12706 gnd.n7735 gnd.n7734 99.6594
R12707 gnd.n199 gnd.n198 99.6594
R12708 gnd.n6293 gnd.n6292 99.6594
R12709 gnd.n6287 gnd.n1257 99.6594
R12710 gnd.n6284 gnd.n1258 99.6594
R12711 gnd.n6280 gnd.n1259 99.6594
R12712 gnd.n6276 gnd.n1260 99.6594
R12713 gnd.n6272 gnd.n1261 99.6594
R12714 gnd.n6268 gnd.n1262 99.6594
R12715 gnd.n6264 gnd.n1263 99.6594
R12716 gnd.n6259 gnd.n1265 99.6594
R12717 gnd.n6255 gnd.n1266 99.6594
R12718 gnd.n6251 gnd.n1267 99.6594
R12719 gnd.n6247 gnd.n1268 99.6594
R12720 gnd.n6243 gnd.n1269 99.6594
R12721 gnd.n6239 gnd.n1270 99.6594
R12722 gnd.n6235 gnd.n1271 99.6594
R12723 gnd.n6231 gnd.n1272 99.6594
R12724 gnd.n6227 gnd.n1273 99.6594
R12725 gnd.n1329 gnd.n1274 99.6594
R12726 gnd.n5555 gnd.n5554 99.6594
R12727 gnd.n5550 gnd.n2076 99.6594
R12728 gnd.n5546 gnd.n2075 99.6594
R12729 gnd.n5542 gnd.n2074 99.6594
R12730 gnd.n5538 gnd.n2073 99.6594
R12731 gnd.n5534 gnd.n2072 99.6594
R12732 gnd.n5530 gnd.n2071 99.6594
R12733 gnd.n4611 gnd.n2069 99.6594
R12734 gnd.n4609 gnd.n2068 99.6594
R12735 gnd.n4605 gnd.n2067 99.6594
R12736 gnd.n4601 gnd.n2066 99.6594
R12737 gnd.n4597 gnd.n2065 99.6594
R12738 gnd.n4593 gnd.n2064 99.6594
R12739 gnd.n4589 gnd.n2063 99.6594
R12740 gnd.n4585 gnd.n2062 99.6594
R12741 gnd.n4581 gnd.n2061 99.6594
R12742 gnd.n4577 gnd.n2060 99.6594
R12743 gnd.n2118 gnd.n2059 99.6594
R12744 gnd.n4186 gnd.n3973 99.6594
R12745 gnd.n4184 gnd.n3976 99.6594
R12746 gnd.n4180 gnd.n4179 99.6594
R12747 gnd.n4173 gnd.n3981 99.6594
R12748 gnd.n4172 gnd.n4171 99.6594
R12749 gnd.n4165 gnd.n3987 99.6594
R12750 gnd.n4164 gnd.n4163 99.6594
R12751 gnd.n4157 gnd.n3993 99.6594
R12752 gnd.n4156 gnd.n4155 99.6594
R12753 gnd.n4149 gnd.n3999 99.6594
R12754 gnd.n4148 gnd.n4147 99.6594
R12755 gnd.n4141 gnd.n4008 99.6594
R12756 gnd.n4140 gnd.n4139 99.6594
R12757 gnd.n4133 gnd.n4014 99.6594
R12758 gnd.n4132 gnd.n4131 99.6594
R12759 gnd.n4125 gnd.n4020 99.6594
R12760 gnd.n4124 gnd.n4123 99.6594
R12761 gnd.n4030 gnd.n4026 99.6594
R12762 gnd.n4113 gnd.n4112 99.6594
R12763 gnd.n3798 gnd.n2355 99.6594
R12764 gnd.n3796 gnd.n2354 99.6594
R12765 gnd.n3792 gnd.n2353 99.6594
R12766 gnd.n3788 gnd.n2352 99.6594
R12767 gnd.n3784 gnd.n2351 99.6594
R12768 gnd.n3780 gnd.n2350 99.6594
R12769 gnd.n3776 gnd.n2349 99.6594
R12770 gnd.n3708 gnd.n2348 99.6594
R12771 gnd.n3039 gnd.n2770 99.6594
R12772 gnd.n2796 gnd.n2777 99.6594
R12773 gnd.n2798 gnd.n2778 99.6594
R12774 gnd.n2806 gnd.n2779 99.6594
R12775 gnd.n2808 gnd.n2780 99.6594
R12776 gnd.n2816 gnd.n2781 99.6594
R12777 gnd.n2818 gnd.n2782 99.6594
R12778 gnd.n2826 gnd.n2783 99.6594
R12779 gnd.n3766 gnd.n2335 99.6594
R12780 gnd.n3762 gnd.n2336 99.6594
R12781 gnd.n3758 gnd.n2337 99.6594
R12782 gnd.n3754 gnd.n2338 99.6594
R12783 gnd.n3750 gnd.n2339 99.6594
R12784 gnd.n3746 gnd.n2340 99.6594
R12785 gnd.n3742 gnd.n2341 99.6594
R12786 gnd.n3738 gnd.n2342 99.6594
R12787 gnd.n3734 gnd.n2343 99.6594
R12788 gnd.n3730 gnd.n2344 99.6594
R12789 gnd.n3726 gnd.n2345 99.6594
R12790 gnd.n3722 gnd.n2346 99.6594
R12791 gnd.n3718 gnd.n2347 99.6594
R12792 gnd.n2954 gnd.n2953 99.6594
R12793 gnd.n2948 gnd.n2865 99.6594
R12794 gnd.n2945 gnd.n2866 99.6594
R12795 gnd.n2941 gnd.n2867 99.6594
R12796 gnd.n2937 gnd.n2868 99.6594
R12797 gnd.n2933 gnd.n2869 99.6594
R12798 gnd.n2929 gnd.n2870 99.6594
R12799 gnd.n2925 gnd.n2871 99.6594
R12800 gnd.n2921 gnd.n2872 99.6594
R12801 gnd.n2917 gnd.n2873 99.6594
R12802 gnd.n2913 gnd.n2874 99.6594
R12803 gnd.n2909 gnd.n2875 99.6594
R12804 gnd.n2956 gnd.n2864 99.6594
R12805 gnd.n7651 gnd.n7650 99.6594
R12806 gnd.n7656 gnd.n7655 99.6594
R12807 gnd.n7659 gnd.n7658 99.6594
R12808 gnd.n7664 gnd.n7663 99.6594
R12809 gnd.n7667 gnd.n7666 99.6594
R12810 gnd.n7672 gnd.n7671 99.6594
R12811 gnd.n7675 gnd.n7674 99.6594
R12812 gnd.n7680 gnd.n7678 99.6594
R12813 gnd.n7806 gnd.n125 99.6594
R12814 gnd.n1339 gnd.n1275 99.6594
R12815 gnd.n1523 gnd.n1276 99.6594
R12816 gnd.n1525 gnd.n1277 99.6594
R12817 gnd.n1542 gnd.n1278 99.6594
R12818 gnd.n1544 gnd.n1279 99.6594
R12819 gnd.n1561 gnd.n1280 99.6594
R12820 gnd.n1563 gnd.n1281 99.6594
R12821 gnd.n1579 gnd.n1282 99.6594
R12822 gnd.n1490 gnd.n1283 99.6594
R12823 gnd.n2046 gnd.n2045 99.6594
R12824 gnd.n2047 gnd.n1995 99.6594
R12825 gnd.n2049 gnd.n2003 99.6594
R12826 gnd.n2051 gnd.n2050 99.6594
R12827 gnd.n2052 gnd.n2012 99.6594
R12828 gnd.n2054 gnd.n2021 99.6594
R12829 gnd.n2056 gnd.n2055 99.6594
R12830 gnd.n2057 gnd.n2030 99.6594
R12831 gnd.n5558 gnd.n5557 99.6594
R12832 gnd.n3833 gnd.n2333 99.6594
R12833 gnd.n3836 gnd.n3835 99.6594
R12834 gnd.n3843 gnd.n3842 99.6594
R12835 gnd.n3846 gnd.n3845 99.6594
R12836 gnd.n3853 gnd.n3852 99.6594
R12837 gnd.n3856 gnd.n3855 99.6594
R12838 gnd.n3863 gnd.n3862 99.6594
R12839 gnd.n3866 gnd.n3865 99.6594
R12840 gnd.n3873 gnd.n3872 99.6594
R12841 gnd.n3834 gnd.n3833 99.6594
R12842 gnd.n3835 gnd.n3828 99.6594
R12843 gnd.n3844 gnd.n3843 99.6594
R12844 gnd.n3845 gnd.n3824 99.6594
R12845 gnd.n3854 gnd.n3853 99.6594
R12846 gnd.n3855 gnd.n3820 99.6594
R12847 gnd.n3864 gnd.n3863 99.6594
R12848 gnd.n3865 gnd.n3816 99.6594
R12849 gnd.n3874 gnd.n3873 99.6594
R12850 gnd.n5557 gnd.n2041 99.6594
R12851 gnd.n2057 gnd.n2029 99.6594
R12852 gnd.n2056 gnd.n2022 99.6594
R12853 gnd.n2054 gnd.n2053 99.6594
R12854 gnd.n2052 gnd.n2011 99.6594
R12855 gnd.n2051 gnd.n2004 99.6594
R12856 gnd.n2049 gnd.n2048 99.6594
R12857 gnd.n2047 gnd.n1994 99.6594
R12858 gnd.n2046 gnd.n2044 99.6594
R12859 gnd.n1522 gnd.n1275 99.6594
R12860 gnd.n1526 gnd.n1276 99.6594
R12861 gnd.n1541 gnd.n1277 99.6594
R12862 gnd.n1545 gnd.n1278 99.6594
R12863 gnd.n1560 gnd.n1279 99.6594
R12864 gnd.n1564 gnd.n1280 99.6594
R12865 gnd.n1578 gnd.n1281 99.6594
R12866 gnd.n1489 gnd.n1282 99.6594
R12867 gnd.n1485 gnd.n1283 99.6594
R12868 gnd.n7679 gnd.n125 99.6594
R12869 gnd.n7678 gnd.n7677 99.6594
R12870 gnd.n7674 gnd.n7673 99.6594
R12871 gnd.n7671 gnd.n7670 99.6594
R12872 gnd.n7666 gnd.n7665 99.6594
R12873 gnd.n7663 gnd.n7662 99.6594
R12874 gnd.n7658 gnd.n7657 99.6594
R12875 gnd.n7655 gnd.n7654 99.6594
R12876 gnd.n7650 gnd.n7649 99.6594
R12877 gnd.n2954 gnd.n2877 99.6594
R12878 gnd.n2946 gnd.n2865 99.6594
R12879 gnd.n2942 gnd.n2866 99.6594
R12880 gnd.n2938 gnd.n2867 99.6594
R12881 gnd.n2934 gnd.n2868 99.6594
R12882 gnd.n2930 gnd.n2869 99.6594
R12883 gnd.n2926 gnd.n2870 99.6594
R12884 gnd.n2922 gnd.n2871 99.6594
R12885 gnd.n2918 gnd.n2872 99.6594
R12886 gnd.n2914 gnd.n2873 99.6594
R12887 gnd.n2910 gnd.n2874 99.6594
R12888 gnd.n2906 gnd.n2875 99.6594
R12889 gnd.n2957 gnd.n2956 99.6594
R12890 gnd.n3721 gnd.n2347 99.6594
R12891 gnd.n3725 gnd.n2346 99.6594
R12892 gnd.n3729 gnd.n2345 99.6594
R12893 gnd.n3733 gnd.n2344 99.6594
R12894 gnd.n3737 gnd.n2343 99.6594
R12895 gnd.n3741 gnd.n2342 99.6594
R12896 gnd.n3745 gnd.n2341 99.6594
R12897 gnd.n3749 gnd.n2340 99.6594
R12898 gnd.n3753 gnd.n2339 99.6594
R12899 gnd.n3757 gnd.n2338 99.6594
R12900 gnd.n3761 gnd.n2337 99.6594
R12901 gnd.n3765 gnd.n2336 99.6594
R12902 gnd.n2376 gnd.n2335 99.6594
R12903 gnd.n3040 gnd.n3039 99.6594
R12904 gnd.n2799 gnd.n2777 99.6594
R12905 gnd.n2805 gnd.n2778 99.6594
R12906 gnd.n2809 gnd.n2779 99.6594
R12907 gnd.n2815 gnd.n2780 99.6594
R12908 gnd.n2819 gnd.n2781 99.6594
R12909 gnd.n2825 gnd.n2782 99.6594
R12910 gnd.n2783 gnd.n2767 99.6594
R12911 gnd.n3775 gnd.n2348 99.6594
R12912 gnd.n3779 gnd.n2349 99.6594
R12913 gnd.n3783 gnd.n2350 99.6594
R12914 gnd.n3787 gnd.n2351 99.6594
R12915 gnd.n3791 gnd.n2352 99.6594
R12916 gnd.n3795 gnd.n2353 99.6594
R12917 gnd.n3799 gnd.n2354 99.6594
R12918 gnd.n2357 gnd.n2355 99.6594
R12919 gnd.n4187 gnd.n4186 99.6594
R12920 gnd.n4181 gnd.n3976 99.6594
R12921 gnd.n4179 gnd.n4178 99.6594
R12922 gnd.n4174 gnd.n4173 99.6594
R12923 gnd.n4171 gnd.n4170 99.6594
R12924 gnd.n4166 gnd.n4165 99.6594
R12925 gnd.n4163 gnd.n4162 99.6594
R12926 gnd.n4158 gnd.n4157 99.6594
R12927 gnd.n4155 gnd.n4154 99.6594
R12928 gnd.n4150 gnd.n4149 99.6594
R12929 gnd.n4147 gnd.n4146 99.6594
R12930 gnd.n4142 gnd.n4141 99.6594
R12931 gnd.n4139 gnd.n4138 99.6594
R12932 gnd.n4134 gnd.n4133 99.6594
R12933 gnd.n4131 gnd.n4130 99.6594
R12934 gnd.n4126 gnd.n4125 99.6594
R12935 gnd.n4123 gnd.n4122 99.6594
R12936 gnd.n4031 gnd.n4030 99.6594
R12937 gnd.n4114 gnd.n4113 99.6594
R12938 gnd.n4576 gnd.n2059 99.6594
R12939 gnd.n4580 gnd.n2060 99.6594
R12940 gnd.n4584 gnd.n2061 99.6594
R12941 gnd.n4588 gnd.n2062 99.6594
R12942 gnd.n4592 gnd.n2063 99.6594
R12943 gnd.n4596 gnd.n2064 99.6594
R12944 gnd.n4600 gnd.n2065 99.6594
R12945 gnd.n4604 gnd.n2066 99.6594
R12946 gnd.n4608 gnd.n2067 99.6594
R12947 gnd.n4612 gnd.n2068 99.6594
R12948 gnd.n5529 gnd.n2070 99.6594
R12949 gnd.n5533 gnd.n2071 99.6594
R12950 gnd.n5537 gnd.n2072 99.6594
R12951 gnd.n5541 gnd.n2073 99.6594
R12952 gnd.n5545 gnd.n2074 99.6594
R12953 gnd.n5549 gnd.n2075 99.6594
R12954 gnd.n2078 gnd.n2076 99.6594
R12955 gnd.n5555 gnd.n2077 99.6594
R12956 gnd.n6293 gnd.n1287 99.6594
R12957 gnd.n6285 gnd.n1257 99.6594
R12958 gnd.n6281 gnd.n1258 99.6594
R12959 gnd.n6277 gnd.n1259 99.6594
R12960 gnd.n6273 gnd.n1260 99.6594
R12961 gnd.n6269 gnd.n1261 99.6594
R12962 gnd.n6265 gnd.n1262 99.6594
R12963 gnd.n6260 gnd.n1264 99.6594
R12964 gnd.n6256 gnd.n1265 99.6594
R12965 gnd.n6252 gnd.n1266 99.6594
R12966 gnd.n6248 gnd.n1267 99.6594
R12967 gnd.n6244 gnd.n1268 99.6594
R12968 gnd.n6240 gnd.n1269 99.6594
R12969 gnd.n6236 gnd.n1270 99.6594
R12970 gnd.n6232 gnd.n1271 99.6594
R12971 gnd.n6228 gnd.n1272 99.6594
R12972 gnd.n1328 gnd.n1273 99.6594
R12973 gnd.n6220 gnd.n1274 99.6594
R12974 gnd.n198 gnd.n195 99.6594
R12975 gnd.n7736 gnd.n7735 99.6594
R12976 gnd.n194 gnd.n188 99.6594
R12977 gnd.n7743 gnd.n7742 99.6594
R12978 gnd.n187 gnd.n181 99.6594
R12979 gnd.n7750 gnd.n7749 99.6594
R12980 gnd.n180 gnd.n174 99.6594
R12981 gnd.n7757 gnd.n7756 99.6594
R12982 gnd.n173 gnd.n167 99.6594
R12983 gnd.n7764 gnd.n7763 99.6594
R12984 gnd.n166 gnd.n160 99.6594
R12985 gnd.n7774 gnd.n7773 99.6594
R12986 gnd.n159 gnd.n153 99.6594
R12987 gnd.n7781 gnd.n7780 99.6594
R12988 gnd.n152 gnd.n146 99.6594
R12989 gnd.n7788 gnd.n7787 99.6594
R12990 gnd.n145 gnd.n139 99.6594
R12991 gnd.n7795 gnd.n7794 99.6594
R12992 gnd.n138 gnd.n135 99.6594
R12993 gnd.n5605 gnd.n5604 99.6594
R12994 gnd.n1998 gnd.n1974 99.6594
R12995 gnd.n2000 gnd.n1975 99.6594
R12996 gnd.n2008 gnd.n1976 99.6594
R12997 gnd.n2016 gnd.n1977 99.6594
R12998 gnd.n2018 gnd.n1978 99.6594
R12999 gnd.n2026 gnd.n1979 99.6594
R13000 gnd.n2036 gnd.n1980 99.6594
R13001 gnd.n2038 gnd.n1981 99.6594
R13002 gnd.n4535 gnd.n1982 99.6594
R13003 gnd.n4537 gnd.n1983 99.6594
R13004 gnd.n4541 gnd.n1984 99.6594
R13005 gnd.n4547 gnd.n1985 99.6594
R13006 gnd.n5607 gnd.n1972 99.6594
R13007 gnd.n5605 gnd.n1988 99.6594
R13008 gnd.n1999 gnd.n1974 99.6594
R13009 gnd.n2007 gnd.n1975 99.6594
R13010 gnd.n2015 gnd.n1976 99.6594
R13011 gnd.n2017 gnd.n1977 99.6594
R13012 gnd.n2025 gnd.n1978 99.6594
R13013 gnd.n2035 gnd.n1979 99.6594
R13014 gnd.n2037 gnd.n1980 99.6594
R13015 gnd.n4534 gnd.n1981 99.6594
R13016 gnd.n4536 gnd.n1982 99.6594
R13017 gnd.n4540 gnd.n1983 99.6594
R13018 gnd.n4542 gnd.n1984 99.6594
R13019 gnd.n4548 gnd.n1985 99.6594
R13020 gnd.n5608 gnd.n5607 99.6594
R13021 gnd.n1531 gnd.n1513 99.6594
R13022 gnd.n1535 gnd.n1533 99.6594
R13023 gnd.n1550 gnd.n1506 99.6594
R13024 gnd.n1554 gnd.n1552 99.6594
R13025 gnd.n1569 gnd.n1499 99.6594
R13026 gnd.n1573 gnd.n1571 99.6594
R13027 gnd.n1585 gnd.n1493 99.6594
R13028 gnd.n1589 gnd.n1587 99.6594
R13029 gnd.n1599 gnd.n1481 99.6594
R13030 gnd.n1602 gnd.n1601 99.6594
R13031 gnd.n1605 gnd.n1604 99.6594
R13032 gnd.n1610 gnd.n1609 99.6594
R13033 gnd.n1613 gnd.n1612 99.6594
R13034 gnd.n6021 gnd.n6020 99.6594
R13035 gnd.n6020 gnd.n6019 99.6594
R13036 gnd.n1612 gnd.n1611 99.6594
R13037 gnd.n1609 gnd.n1608 99.6594
R13038 gnd.n1604 gnd.n1603 99.6594
R13039 gnd.n1601 gnd.n1600 99.6594
R13040 gnd.n1588 gnd.n1481 99.6594
R13041 gnd.n1587 gnd.n1586 99.6594
R13042 gnd.n1572 gnd.n1493 99.6594
R13043 gnd.n1571 gnd.n1570 99.6594
R13044 gnd.n1553 gnd.n1499 99.6594
R13045 gnd.n1552 gnd.n1551 99.6594
R13046 gnd.n1534 gnd.n1506 99.6594
R13047 gnd.n1533 gnd.n1532 99.6594
R13048 gnd.n1513 gnd.n1244 99.6594
R13049 gnd.n4543 gnd.t251 98.63
R13050 gnd.n122 gnd.t257 98.63
R13051 gnd.n1486 gnd.t273 98.63
R13052 gnd.n2031 gnd.t292 98.63
R13053 gnd.n1308 gnd.t243 98.63
R13054 gnd.n1330 gnd.t226 98.63
R13055 gnd.n201 gnd.t286 98.63
R13056 gnd.n7767 gnd.t204 98.63
R13057 gnd.n4000 gnd.t302 98.63
R13058 gnd.n4032 gnd.t281 98.63
R13059 gnd.n3813 gnd.t299 98.63
R13060 gnd.n2120 gnd.t295 98.63
R13061 gnd.n2098 gnd.t218 98.63
R13062 gnd.n6029 gnd.t214 98.63
R13063 gnd.n4680 gnd.t284 96.6984
R13064 gnd.n5052 gnd.t232 96.6984
R13065 gnd.n5458 gnd.t237 96.6906
R13066 gnd.n5046 gnd.t269 96.6906
R13067 gnd.n7143 gnd.n7142 84.8607
R13068 gnd.n7144 gnd.n7143 84.8607
R13069 gnd.n7144 gnd.n540 84.8607
R13070 gnd.n7152 gnd.n540 84.8607
R13071 gnd.n7153 gnd.n7152 84.8607
R13072 gnd.n7154 gnd.n7153 84.8607
R13073 gnd.n7154 gnd.n534 84.8607
R13074 gnd.n7162 gnd.n534 84.8607
R13075 gnd.n7163 gnd.n7162 84.8607
R13076 gnd.n7164 gnd.n7163 84.8607
R13077 gnd.n7164 gnd.n528 84.8607
R13078 gnd.n7172 gnd.n528 84.8607
R13079 gnd.n7173 gnd.n7172 84.8607
R13080 gnd.n7174 gnd.n7173 84.8607
R13081 gnd.n7174 gnd.n522 84.8607
R13082 gnd.n7182 gnd.n522 84.8607
R13083 gnd.n7183 gnd.n7182 84.8607
R13084 gnd.n7184 gnd.n7183 84.8607
R13085 gnd.n7184 gnd.n516 84.8607
R13086 gnd.n7192 gnd.n516 84.8607
R13087 gnd.n7193 gnd.n7192 84.8607
R13088 gnd.n7194 gnd.n7193 84.8607
R13089 gnd.n7194 gnd.n510 84.8607
R13090 gnd.n7202 gnd.n510 84.8607
R13091 gnd.n7203 gnd.n7202 84.8607
R13092 gnd.n7204 gnd.n7203 84.8607
R13093 gnd.n7204 gnd.n504 84.8607
R13094 gnd.n7212 gnd.n504 84.8607
R13095 gnd.n7213 gnd.n7212 84.8607
R13096 gnd.n7214 gnd.n7213 84.8607
R13097 gnd.n7214 gnd.n498 84.8607
R13098 gnd.n7222 gnd.n498 84.8607
R13099 gnd.n7223 gnd.n7222 84.8607
R13100 gnd.n7224 gnd.n7223 84.8607
R13101 gnd.n7224 gnd.n492 84.8607
R13102 gnd.n7232 gnd.n492 84.8607
R13103 gnd.n7233 gnd.n7232 84.8607
R13104 gnd.n7234 gnd.n7233 84.8607
R13105 gnd.n7234 gnd.n486 84.8607
R13106 gnd.n7242 gnd.n486 84.8607
R13107 gnd.n7243 gnd.n7242 84.8607
R13108 gnd.n7244 gnd.n7243 84.8607
R13109 gnd.n7244 gnd.n480 84.8607
R13110 gnd.n7252 gnd.n480 84.8607
R13111 gnd.n7253 gnd.n7252 84.8607
R13112 gnd.n7254 gnd.n7253 84.8607
R13113 gnd.n7254 gnd.n474 84.8607
R13114 gnd.n7262 gnd.n474 84.8607
R13115 gnd.n7263 gnd.n7262 84.8607
R13116 gnd.n7264 gnd.n7263 84.8607
R13117 gnd.n7264 gnd.n468 84.8607
R13118 gnd.n7272 gnd.n468 84.8607
R13119 gnd.n7273 gnd.n7272 84.8607
R13120 gnd.n7274 gnd.n7273 84.8607
R13121 gnd.n7274 gnd.n462 84.8607
R13122 gnd.n7282 gnd.n462 84.8607
R13123 gnd.n7283 gnd.n7282 84.8607
R13124 gnd.n7284 gnd.n7283 84.8607
R13125 gnd.n7284 gnd.n456 84.8607
R13126 gnd.n7292 gnd.n456 84.8607
R13127 gnd.n7293 gnd.n7292 84.8607
R13128 gnd.n7294 gnd.n7293 84.8607
R13129 gnd.n7294 gnd.n450 84.8607
R13130 gnd.n7302 gnd.n450 84.8607
R13131 gnd.n7303 gnd.n7302 84.8607
R13132 gnd.n7304 gnd.n7303 84.8607
R13133 gnd.n7304 gnd.n444 84.8607
R13134 gnd.n7312 gnd.n444 84.8607
R13135 gnd.n7313 gnd.n7312 84.8607
R13136 gnd.n7314 gnd.n7313 84.8607
R13137 gnd.n7314 gnd.n438 84.8607
R13138 gnd.n7322 gnd.n438 84.8607
R13139 gnd.n7323 gnd.n7322 84.8607
R13140 gnd.n7324 gnd.n7323 84.8607
R13141 gnd.n7324 gnd.n432 84.8607
R13142 gnd.n7332 gnd.n432 84.8607
R13143 gnd.n7333 gnd.n7332 84.8607
R13144 gnd.n7334 gnd.n7333 84.8607
R13145 gnd.n7334 gnd.n426 84.8607
R13146 gnd.n7342 gnd.n426 84.8607
R13147 gnd.n7343 gnd.n7342 84.8607
R13148 gnd.n7345 gnd.n7343 84.8607
R13149 gnd.n7345 gnd.n7344 84.8607
R13150 gnd.n4665 gnd.n4664 81.8399
R13151 gnd.n2828 gnd.t305 74.8376
R13152 gnd.n2373 gnd.t247 74.8376
R13153 gnd.n4681 gnd.t283 72.8438
R13154 gnd.n5053 gnd.t233 72.8438
R13155 gnd.n4666 gnd.n4659 72.8411
R13156 gnd.n4672 gnd.n4657 72.8411
R13157 gnd.n5021 gnd.n5020 72.8411
R13158 gnd.n4544 gnd.t250 72.836
R13159 gnd.n5459 gnd.t236 72.836
R13160 gnd.n5047 gnd.t270 72.836
R13161 gnd.n123 gnd.t258 72.836
R13162 gnd.n1487 gnd.t272 72.836
R13163 gnd.n2032 gnd.t293 72.836
R13164 gnd.n1309 gnd.t242 72.836
R13165 gnd.n1331 gnd.t225 72.836
R13166 gnd.n202 gnd.t287 72.836
R13167 gnd.n7768 gnd.t205 72.836
R13168 gnd.n4001 gnd.t301 72.836
R13169 gnd.n4033 gnd.t280 72.836
R13170 gnd.n3814 gnd.t298 72.836
R13171 gnd.n2121 gnd.t296 72.836
R13172 gnd.n2099 gnd.t219 72.836
R13173 gnd.n6030 gnd.t215 72.836
R13174 gnd.n5190 gnd.n5026 71.676
R13175 gnd.n5188 gnd.n5187 71.676
R13176 gnd.n5183 gnd.n5029 71.676
R13177 gnd.n5181 gnd.n5180 71.676
R13178 gnd.n5176 gnd.n5032 71.676
R13179 gnd.n5174 gnd.n5173 71.676
R13180 gnd.n5169 gnd.n5035 71.676
R13181 gnd.n5167 gnd.n5166 71.676
R13182 gnd.n5162 gnd.n5038 71.676
R13183 gnd.n5160 gnd.n5159 71.676
R13184 gnd.n5155 gnd.n5041 71.676
R13185 gnd.n5153 gnd.n5152 71.676
R13186 gnd.n5148 gnd.n5044 71.676
R13187 gnd.n5146 gnd.n5145 71.676
R13188 gnd.n5140 gnd.n5049 71.676
R13189 gnd.n5138 gnd.n5137 71.676
R13190 gnd.n5133 gnd.n5132 71.676
R13191 gnd.n5130 gnd.n5129 71.676
R13192 gnd.n5124 gnd.n5055 71.676
R13193 gnd.n5122 gnd.n5121 71.676
R13194 gnd.n5117 gnd.n5058 71.676
R13195 gnd.n5115 gnd.n5114 71.676
R13196 gnd.n5110 gnd.n5061 71.676
R13197 gnd.n5108 gnd.n5107 71.676
R13198 gnd.n5103 gnd.n5064 71.676
R13199 gnd.n5101 gnd.n5100 71.676
R13200 gnd.n5096 gnd.n5067 71.676
R13201 gnd.n5094 gnd.n5093 71.676
R13202 gnd.n5089 gnd.n5070 71.676
R13203 gnd.n5087 gnd.n5086 71.676
R13204 gnd.n5082 gnd.n5073 71.676
R13205 gnd.n5080 gnd.n5079 71.676
R13206 gnd.n5074 gnd.n5000 71.676
R13207 gnd.n5522 gnd.n5521 71.676
R13208 gnd.n5516 gnd.n4621 71.676
R13209 gnd.n5513 gnd.n4622 71.676
R13210 gnd.n5509 gnd.n4623 71.676
R13211 gnd.n5505 gnd.n4624 71.676
R13212 gnd.n5501 gnd.n4625 71.676
R13213 gnd.n5497 gnd.n4626 71.676
R13214 gnd.n5493 gnd.n4627 71.676
R13215 gnd.n5489 gnd.n4628 71.676
R13216 gnd.n5485 gnd.n4629 71.676
R13217 gnd.n5481 gnd.n4630 71.676
R13218 gnd.n5477 gnd.n4631 71.676
R13219 gnd.n5473 gnd.n4632 71.676
R13220 gnd.n5469 gnd.n4633 71.676
R13221 gnd.n5465 gnd.n4634 71.676
R13222 gnd.n5461 gnd.n4635 71.676
R13223 gnd.n4636 gnd.n4620 71.676
R13224 gnd.n4684 gnd.n4637 71.676
R13225 gnd.n4689 gnd.n4638 71.676
R13226 gnd.n4693 gnd.n4639 71.676
R13227 gnd.n4697 gnd.n4640 71.676
R13228 gnd.n4701 gnd.n4641 71.676
R13229 gnd.n4705 gnd.n4642 71.676
R13230 gnd.n4709 gnd.n4643 71.676
R13231 gnd.n4713 gnd.n4644 71.676
R13232 gnd.n4717 gnd.n4645 71.676
R13233 gnd.n4721 gnd.n4646 71.676
R13234 gnd.n4725 gnd.n4647 71.676
R13235 gnd.n4729 gnd.n4648 71.676
R13236 gnd.n4733 gnd.n4649 71.676
R13237 gnd.n4737 gnd.n4650 71.676
R13238 gnd.n4741 gnd.n4651 71.676
R13239 gnd.n5522 gnd.n4654 71.676
R13240 gnd.n5514 gnd.n4621 71.676
R13241 gnd.n5510 gnd.n4622 71.676
R13242 gnd.n5506 gnd.n4623 71.676
R13243 gnd.n5502 gnd.n4624 71.676
R13244 gnd.n5498 gnd.n4625 71.676
R13245 gnd.n5494 gnd.n4626 71.676
R13246 gnd.n5490 gnd.n4627 71.676
R13247 gnd.n5486 gnd.n4628 71.676
R13248 gnd.n5482 gnd.n4629 71.676
R13249 gnd.n5478 gnd.n4630 71.676
R13250 gnd.n5474 gnd.n4631 71.676
R13251 gnd.n5470 gnd.n4632 71.676
R13252 gnd.n5466 gnd.n4633 71.676
R13253 gnd.n5462 gnd.n4634 71.676
R13254 gnd.n5525 gnd.n5524 71.676
R13255 gnd.n4683 gnd.n4636 71.676
R13256 gnd.n4688 gnd.n4637 71.676
R13257 gnd.n4692 gnd.n4638 71.676
R13258 gnd.n4696 gnd.n4639 71.676
R13259 gnd.n4700 gnd.n4640 71.676
R13260 gnd.n4704 gnd.n4641 71.676
R13261 gnd.n4708 gnd.n4642 71.676
R13262 gnd.n4712 gnd.n4643 71.676
R13263 gnd.n4716 gnd.n4644 71.676
R13264 gnd.n4720 gnd.n4645 71.676
R13265 gnd.n4724 gnd.n4646 71.676
R13266 gnd.n4728 gnd.n4647 71.676
R13267 gnd.n4732 gnd.n4648 71.676
R13268 gnd.n4736 gnd.n4649 71.676
R13269 gnd.n4740 gnd.n4650 71.676
R13270 gnd.n4743 gnd.n4651 71.676
R13271 gnd.n5075 gnd.n5074 71.676
R13272 gnd.n5081 gnd.n5080 71.676
R13273 gnd.n5073 gnd.n5071 71.676
R13274 gnd.n5088 gnd.n5087 71.676
R13275 gnd.n5070 gnd.n5068 71.676
R13276 gnd.n5095 gnd.n5094 71.676
R13277 gnd.n5067 gnd.n5065 71.676
R13278 gnd.n5102 gnd.n5101 71.676
R13279 gnd.n5064 gnd.n5062 71.676
R13280 gnd.n5109 gnd.n5108 71.676
R13281 gnd.n5061 gnd.n5059 71.676
R13282 gnd.n5116 gnd.n5115 71.676
R13283 gnd.n5058 gnd.n5056 71.676
R13284 gnd.n5123 gnd.n5122 71.676
R13285 gnd.n5055 gnd.n5051 71.676
R13286 gnd.n5131 gnd.n5130 71.676
R13287 gnd.n5135 gnd.n5134 71.676
R13288 gnd.n5139 gnd.n5138 71.676
R13289 gnd.n5049 gnd.n5045 71.676
R13290 gnd.n5147 gnd.n5146 71.676
R13291 gnd.n5044 gnd.n5042 71.676
R13292 gnd.n5154 gnd.n5153 71.676
R13293 gnd.n5041 gnd.n5039 71.676
R13294 gnd.n5161 gnd.n5160 71.676
R13295 gnd.n5038 gnd.n5036 71.676
R13296 gnd.n5168 gnd.n5167 71.676
R13297 gnd.n5035 gnd.n5033 71.676
R13298 gnd.n5175 gnd.n5174 71.676
R13299 gnd.n5032 gnd.n5030 71.676
R13300 gnd.n5182 gnd.n5181 71.676
R13301 gnd.n5029 gnd.n5027 71.676
R13302 gnd.n5189 gnd.n5188 71.676
R13303 gnd.n5026 gnd.n5002 71.676
R13304 gnd.n10 gnd.t59 69.1507
R13305 gnd.n18 gnd.t308 68.4792
R13306 gnd.n17 gnd.t363 68.4792
R13307 gnd.n16 gnd.t1 68.4792
R13308 gnd.n15 gnd.t133 68.4792
R13309 gnd.n14 gnd.t310 68.4792
R13310 gnd.n13 gnd.t338 68.4792
R13311 gnd.n12 gnd.t3 68.4792
R13312 gnd.n11 gnd.t340 68.4792
R13313 gnd.n10 gnd.t195 68.4792
R13314 gnd.n2955 gnd.n2859 64.369
R13315 gnd.n4686 gnd.n4681 59.5399
R13316 gnd.n5126 gnd.n5053 59.5399
R13317 gnd.n5460 gnd.n5459 59.5399
R13318 gnd.n5142 gnd.n5047 59.5399
R13319 gnd.n5457 gnd.n4675 59.1804
R13320 gnd.n2606 gnd.t112 56.607
R13321 gnd.n60 gnd.t10 56.607
R13322 gnd.n2567 gnd.t361 56.407
R13323 gnd.n2586 gnd.t173 56.407
R13324 gnd.n21 gnd.t140 56.407
R13325 gnd.n40 gnd.t170 56.407
R13326 gnd.n2623 gnd.t314 55.8337
R13327 gnd.n2584 gnd.t343 55.8337
R13328 gnd.n2603 gnd.t175 55.8337
R13329 gnd.n77 gnd.t152 55.8337
R13330 gnd.n38 gnd.t347 55.8337
R13331 gnd.n57 gnd.t165 55.8337
R13332 gnd.n4663 gnd.n4662 54.358
R13333 gnd.n5018 gnd.n5017 54.358
R13334 gnd.n2606 gnd.n2605 53.0052
R13335 gnd.n2608 gnd.n2607 53.0052
R13336 gnd.n2610 gnd.n2609 53.0052
R13337 gnd.n2612 gnd.n2611 53.0052
R13338 gnd.n2614 gnd.n2613 53.0052
R13339 gnd.n2616 gnd.n2615 53.0052
R13340 gnd.n2618 gnd.n2617 53.0052
R13341 gnd.n2620 gnd.n2619 53.0052
R13342 gnd.n2622 gnd.n2621 53.0052
R13343 gnd.n2567 gnd.n2566 53.0052
R13344 gnd.n2569 gnd.n2568 53.0052
R13345 gnd.n2571 gnd.n2570 53.0052
R13346 gnd.n2573 gnd.n2572 53.0052
R13347 gnd.n2575 gnd.n2574 53.0052
R13348 gnd.n2577 gnd.n2576 53.0052
R13349 gnd.n2579 gnd.n2578 53.0052
R13350 gnd.n2581 gnd.n2580 53.0052
R13351 gnd.n2583 gnd.n2582 53.0052
R13352 gnd.n2586 gnd.n2585 53.0052
R13353 gnd.n2588 gnd.n2587 53.0052
R13354 gnd.n2590 gnd.n2589 53.0052
R13355 gnd.n2592 gnd.n2591 53.0052
R13356 gnd.n2594 gnd.n2593 53.0052
R13357 gnd.n2596 gnd.n2595 53.0052
R13358 gnd.n2598 gnd.n2597 53.0052
R13359 gnd.n2600 gnd.n2599 53.0052
R13360 gnd.n2602 gnd.n2601 53.0052
R13361 gnd.n76 gnd.n75 53.0052
R13362 gnd.n74 gnd.n73 53.0052
R13363 gnd.n72 gnd.n71 53.0052
R13364 gnd.n70 gnd.n69 53.0052
R13365 gnd.n68 gnd.n67 53.0052
R13366 gnd.n66 gnd.n65 53.0052
R13367 gnd.n64 gnd.n63 53.0052
R13368 gnd.n62 gnd.n61 53.0052
R13369 gnd.n60 gnd.n59 53.0052
R13370 gnd.n37 gnd.n36 53.0052
R13371 gnd.n35 gnd.n34 53.0052
R13372 gnd.n33 gnd.n32 53.0052
R13373 gnd.n31 gnd.n30 53.0052
R13374 gnd.n29 gnd.n28 53.0052
R13375 gnd.n27 gnd.n26 53.0052
R13376 gnd.n25 gnd.n24 53.0052
R13377 gnd.n23 gnd.n22 53.0052
R13378 gnd.n21 gnd.n20 53.0052
R13379 gnd.n56 gnd.n55 53.0052
R13380 gnd.n54 gnd.n53 53.0052
R13381 gnd.n52 gnd.n51 53.0052
R13382 gnd.n50 gnd.n49 53.0052
R13383 gnd.n48 gnd.n47 53.0052
R13384 gnd.n46 gnd.n45 53.0052
R13385 gnd.n44 gnd.n43 53.0052
R13386 gnd.n42 gnd.n41 53.0052
R13387 gnd.n40 gnd.n39 53.0052
R13388 gnd.n5009 gnd.n5008 52.4801
R13389 gnd.n3659 gnd.t126 52.3082
R13390 gnd.n3627 gnd.t95 52.3082
R13391 gnd.n3595 gnd.t25 52.3082
R13392 gnd.n3564 gnd.t163 52.3082
R13393 gnd.n3532 gnd.t320 52.3082
R13394 gnd.n3500 gnd.t17 52.3082
R13395 gnd.n3468 gnd.t167 52.3082
R13396 gnd.n3437 gnd.t180 52.3082
R13397 gnd.n4194 gnd.n3808 51.6227
R13398 gnd.n7804 gnd.n128 51.6227
R13399 gnd.n3489 gnd.n3457 51.4173
R13400 gnd.n7344 gnd.n238 50.9166
R13401 gnd.n3553 gnd.n3552 50.455
R13402 gnd.n3521 gnd.n3520 50.455
R13403 gnd.n3489 gnd.n3488 50.455
R13404 gnd.n2902 gnd.n2901 45.1884
R13405 gnd.n2399 gnd.n2398 45.1884
R13406 gnd.n5193 gnd.n5024 44.3322
R13407 gnd.n4666 gnd.n4665 44.3189
R13408 gnd.n4545 gnd.n4544 42.4732
R13409 gnd.n6031 gnd.n6030 42.4732
R13410 gnd.n2903 gnd.n2902 42.2793
R13411 gnd.n2400 gnd.n2399 42.2793
R13412 gnd.n2829 gnd.n2828 42.2793
R13413 gnd.n3774 gnd.n2373 42.2793
R13414 gnd.n124 gnd.n123 42.2793
R13415 gnd.n1594 gnd.n1487 42.2793
R13416 gnd.n2033 gnd.n2032 42.2793
R13417 gnd.n1332 gnd.n1331 42.2793
R13418 gnd.n7732 gnd.n202 42.2793
R13419 gnd.n7769 gnd.n7768 42.2793
R13420 gnd.n4002 gnd.n4001 42.2793
R13421 gnd.n4034 gnd.n4033 42.2793
R13422 gnd.n3815 gnd.n3814 42.2793
R13423 gnd.n4575 gnd.n2121 42.2793
R13424 gnd.n4664 gnd.n4663 41.6274
R13425 gnd.n5019 gnd.n5018 41.6274
R13426 gnd.n4673 gnd.n4672 40.8975
R13427 gnd.n5022 gnd.n5021 40.8975
R13428 gnd.n6262 gnd.n1309 36.9518
R13429 gnd.n5527 gnd.n2099 36.9518
R13430 gnd.n4672 gnd.n4671 35.055
R13431 gnd.n4667 gnd.n4666 35.055
R13432 gnd.n5011 gnd.n5010 35.055
R13433 gnd.n5021 gnd.n5007 35.055
R13434 gnd.n5076 gnd.n4999 32.9371
R13435 gnd.n4745 gnd.n4744 32.9371
R13436 gnd.n6713 gnd.n797 31.9958
R13437 gnd.n6713 gnd.n6712 31.9958
R13438 gnd.n6712 gnd.n6711 31.9958
R13439 gnd.n6711 gnd.n802 31.9958
R13440 gnd.n6705 gnd.n802 31.9958
R13441 gnd.n6705 gnd.n6704 31.9958
R13442 gnd.n6704 gnd.n6703 31.9958
R13443 gnd.n6703 gnd.n810 31.9958
R13444 gnd.n6697 gnd.n810 31.9958
R13445 gnd.n6697 gnd.n6696 31.9958
R13446 gnd.n6696 gnd.n6695 31.9958
R13447 gnd.n6695 gnd.n818 31.9958
R13448 gnd.n6689 gnd.n818 31.9958
R13449 gnd.n6689 gnd.n6688 31.9958
R13450 gnd.n6688 gnd.n6687 31.9958
R13451 gnd.n6687 gnd.n826 31.9958
R13452 gnd.n6681 gnd.n826 31.9958
R13453 gnd.n6681 gnd.n6680 31.9958
R13454 gnd.n6680 gnd.n6679 31.9958
R13455 gnd.n6679 gnd.n834 31.9958
R13456 gnd.n6673 gnd.n834 31.9958
R13457 gnd.n6673 gnd.n6672 31.9958
R13458 gnd.n6672 gnd.n6671 31.9958
R13459 gnd.n6671 gnd.n842 31.9958
R13460 gnd.n6665 gnd.n842 31.9958
R13461 gnd.n6665 gnd.n6664 31.9958
R13462 gnd.n6664 gnd.n6663 31.9958
R13463 gnd.n6663 gnd.n850 31.9958
R13464 gnd.n6657 gnd.n850 31.9958
R13465 gnd.n6657 gnd.n6656 31.9958
R13466 gnd.n6656 gnd.n6655 31.9958
R13467 gnd.n6655 gnd.n858 31.9958
R13468 gnd.n6649 gnd.n858 31.9958
R13469 gnd.n6649 gnd.n6648 31.9958
R13470 gnd.n6648 gnd.n6647 31.9958
R13471 gnd.n6647 gnd.n866 31.9958
R13472 gnd.n6641 gnd.n866 31.9958
R13473 gnd.n6641 gnd.n6640 31.9958
R13474 gnd.n6640 gnd.n6639 31.9958
R13475 gnd.n6639 gnd.n874 31.9958
R13476 gnd.n6633 gnd.n874 31.9958
R13477 gnd.n6633 gnd.n6632 31.9958
R13478 gnd.n6632 gnd.n6631 31.9958
R13479 gnd.n6631 gnd.n882 31.9958
R13480 gnd.n6625 gnd.n882 31.9958
R13481 gnd.n6625 gnd.n6624 31.9958
R13482 gnd.n6624 gnd.n6623 31.9958
R13483 gnd.n6623 gnd.n890 31.9958
R13484 gnd.n6617 gnd.n890 31.9958
R13485 gnd.n6617 gnd.n6616 31.9958
R13486 gnd.n6616 gnd.n6615 31.9958
R13487 gnd.n6615 gnd.n898 31.9958
R13488 gnd.n6609 gnd.n898 31.9958
R13489 gnd.n6609 gnd.n6608 31.9958
R13490 gnd.n6608 gnd.n6607 31.9958
R13491 gnd.n6607 gnd.n906 31.9958
R13492 gnd.n6601 gnd.n906 31.9958
R13493 gnd.n6601 gnd.n6600 31.9958
R13494 gnd.n6600 gnd.n6599 31.9958
R13495 gnd.n6599 gnd.n914 31.9958
R13496 gnd.n6593 gnd.n914 31.9958
R13497 gnd.n6593 gnd.n6592 31.9958
R13498 gnd.n6592 gnd.n6591 31.9958
R13499 gnd.n6591 gnd.n922 31.9958
R13500 gnd.n6585 gnd.n922 31.9958
R13501 gnd.n6585 gnd.n6584 31.9958
R13502 gnd.n6584 gnd.n6583 31.9958
R13503 gnd.n6583 gnd.n930 31.9958
R13504 gnd.n6577 gnd.n930 31.9958
R13505 gnd.n6577 gnd.n6576 31.9958
R13506 gnd.n6576 gnd.n6575 31.9958
R13507 gnd.n6575 gnd.n938 31.9958
R13508 gnd.n6569 gnd.n938 31.9958
R13509 gnd.n6569 gnd.n6568 31.9958
R13510 gnd.n6568 gnd.n6567 31.9958
R13511 gnd.n6567 gnd.n946 31.9958
R13512 gnd.n6561 gnd.n946 31.9958
R13513 gnd.n6561 gnd.n6560 31.9958
R13514 gnd.n6560 gnd.n6559 31.9958
R13515 gnd.n6559 gnd.n954 31.9958
R13516 gnd.n6553 gnd.n954 31.9958
R13517 gnd.n6553 gnd.n6552 31.9958
R13518 gnd.n6552 gnd.n6551 31.9958
R13519 gnd.n2965 gnd.n2859 31.8661
R13520 gnd.n2965 gnd.n2964 31.8661
R13521 gnd.n2973 gnd.n2848 31.8661
R13522 gnd.n2981 gnd.n2848 31.8661
R13523 gnd.n2981 gnd.n2842 31.8661
R13524 gnd.n2989 gnd.n2842 31.8661
R13525 gnd.n2989 gnd.n2835 31.8661
R13526 gnd.n3027 gnd.n2835 31.8661
R13527 gnd.n3037 gnd.n2768 31.8661
R13528 gnd.n4194 gnd.n3972 31.8661
R13529 gnd.n4202 gnd.n2320 31.8661
R13530 gnd.n4210 gnd.n2320 31.8661
R13531 gnd.n4210 gnd.n2312 31.8661
R13532 gnd.n4218 gnd.n2312 31.8661
R13533 gnd.n4226 gnd.n2303 31.8661
R13534 gnd.n4226 gnd.n2306 31.8661
R13535 gnd.n4234 gnd.n2288 31.8661
R13536 gnd.n4242 gnd.n2288 31.8661
R13537 gnd.n4250 gnd.n2280 31.8661
R13538 gnd.n4258 gnd.n2271 31.8661
R13539 gnd.n4258 gnd.n2274 31.8661
R13540 gnd.n4266 gnd.n2256 31.8661
R13541 gnd.n4274 gnd.n2256 31.8661
R13542 gnd.n4282 gnd.n2248 31.8661
R13543 gnd.n4291 gnd.n2239 31.8661
R13544 gnd.n4291 gnd.n2242 31.8661
R13545 gnd.n4299 gnd.n2225 31.8661
R13546 gnd.n4307 gnd.n2225 31.8661
R13547 gnd.n4316 gnd.n2216 31.8661
R13548 gnd.n4324 gnd.n2209 31.8661
R13549 gnd.n4324 gnd.n2211 31.8661
R13550 gnd.n4343 gnd.n2193 31.8661
R13551 gnd.n4350 gnd.n970 31.8661
R13552 gnd.n2042 gnd.n1112 31.8661
R13553 gnd.n4492 gnd.n2058 31.8661
R13554 gnd.n4492 gnd.n1973 31.8661
R13555 gnd.n1986 gnd.n1967 31.8661
R13556 gnd.n5615 gnd.n1967 31.8661
R13557 gnd.n5623 gnd.n1960 31.8661
R13558 gnd.n5623 gnd.n1953 31.8661
R13559 gnd.n5631 gnd.n1953 31.8661
R13560 gnd.n5631 gnd.n1954 31.8661
R13561 gnd.n5639 gnd.n1941 31.8661
R13562 gnd.n5647 gnd.n1941 31.8661
R13563 gnd.n5647 gnd.n1934 31.8661
R13564 gnd.n5655 gnd.n1934 31.8661
R13565 gnd.n5967 gnd.n1653 31.8661
R13566 gnd.n5975 gnd.n1646 31.8661
R13567 gnd.n5975 gnd.n1639 31.8661
R13568 gnd.n5983 gnd.n1639 31.8661
R13569 gnd.n5983 gnd.n1640 31.8661
R13570 gnd.n5991 gnd.n1626 31.8661
R13571 gnd.n6001 gnd.n1626 31.8661
R13572 gnd.n6001 gnd.n1618 31.8661
R13573 gnd.n6012 gnd.n1618 31.8661
R13574 gnd.n6303 gnd.n1245 31.8661
R13575 gnd.n6303 gnd.n6302 31.8661
R13576 gnd.n6296 gnd.n1256 31.8661
R13577 gnd.n6296 gnd.n6295 31.8661
R13578 gnd.n1336 gnd.n1285 31.8661
R13579 gnd.n7444 gnd.n350 31.8661
R13580 gnd.n7551 gnd.n315 31.8661
R13581 gnd.n7453 gnd.n340 31.8661
R13582 gnd.n7459 gnd.n340 31.8661
R13583 gnd.n7532 gnd.n334 31.8661
R13584 gnd.n7536 gnd.n299 31.8661
R13585 gnd.n7560 gnd.n299 31.8661
R13586 gnd.n7568 gnd.n290 31.8661
R13587 gnd.n7568 gnd.n293 31.8661
R13588 gnd.n7576 gnd.n284 31.8661
R13589 gnd.n7584 gnd.n269 31.8661
R13590 gnd.n7592 gnd.n269 31.8661
R13591 gnd.n7600 gnd.n260 31.8661
R13592 gnd.n7600 gnd.n263 31.8661
R13593 gnd.n7608 gnd.n254 31.8661
R13594 gnd.n7616 gnd.n247 31.8661
R13595 gnd.n7632 gnd.n229 31.8661
R13596 gnd.n7632 gnd.n232 31.8661
R13597 gnd.n7640 gnd.n213 31.8661
R13598 gnd.n7716 gnd.n213 31.8661
R13599 gnd.n7716 gnd.n206 31.8661
R13600 gnd.n7724 gnd.n206 31.8661
R13601 gnd.n7804 gnd.n126 31.8661
R13602 gnd.t11 gnd.n2216 31.5474
R13603 gnd.n7532 gnd.t107 31.5474
R13604 gnd.t186 gnd.n2248 30.9101
R13605 gnd.n284 gnd.t65 30.9101
R13606 gnd.n3807 gnd.n962 30.2728
R13607 gnd.t52 gnd.n2280 30.2728
R13608 gnd.n254 gnd.t20 30.2728
R13609 gnd.n3972 gnd.t279 28.3609
R13610 gnd.t203 gnd.n126 28.3609
R13611 gnd.n2408 gnd.n962 27.0862
R13612 gnd.n4544 gnd.n4543 25.7944
R13613 gnd.n2828 gnd.n2827 25.7944
R13614 gnd.n2373 gnd.n2372 25.7944
R13615 gnd.n123 gnd.n122 25.7944
R13616 gnd.n1487 gnd.n1486 25.7944
R13617 gnd.n2032 gnd.n2031 25.7944
R13618 gnd.n1309 gnd.n1308 25.7944
R13619 gnd.n1331 gnd.n1330 25.7944
R13620 gnd.n202 gnd.n201 25.7944
R13621 gnd.n7768 gnd.n7767 25.7944
R13622 gnd.n4001 gnd.n4000 25.7944
R13623 gnd.n4033 gnd.n4032 25.7944
R13624 gnd.n3814 gnd.n3813 25.7944
R13625 gnd.n2121 gnd.n2120 25.7944
R13626 gnd.n2099 gnd.n2098 25.7944
R13627 gnd.n6030 gnd.n6029 25.7944
R13628 gnd.n3049 gnd.n2769 24.8557
R13629 gnd.n3059 gnd.n2752 24.8557
R13630 gnd.n2755 gnd.n2743 24.8557
R13631 gnd.n3080 gnd.n2744 24.8557
R13632 gnd.n3090 gnd.n2724 24.8557
R13633 gnd.n3100 gnd.n3099 24.8557
R13634 gnd.n2710 gnd.n2708 24.8557
R13635 gnd.n3131 gnd.n3130 24.8557
R13636 gnd.n3146 gnd.n2693 24.8557
R13637 gnd.n3200 gnd.n2632 24.8557
R13638 gnd.n3156 gnd.n2633 24.8557
R13639 gnd.n3193 gnd.n2644 24.8557
R13640 gnd.n2682 gnd.n2681 24.8557
R13641 gnd.n3187 gnd.n3186 24.8557
R13642 gnd.n2668 gnd.n2655 24.8557
R13643 gnd.n3226 gnd.n3225 24.8557
R13644 gnd.n3236 gnd.n2552 24.8557
R13645 gnd.n3248 gnd.n2544 24.8557
R13646 gnd.n3247 gnd.n2532 24.8557
R13647 gnd.n3266 gnd.n3265 24.8557
R13648 gnd.n3276 gnd.n2525 24.8557
R13649 gnd.n3287 gnd.n2513 24.8557
R13650 gnd.n3311 gnd.n3310 24.8557
R13651 gnd.n3322 gnd.n2496 24.8557
R13652 gnd.n3321 gnd.n2498 24.8557
R13653 gnd.n3333 gnd.n2489 24.8557
R13654 gnd.n3351 gnd.n3350 24.8557
R13655 gnd.n2480 gnd.n2469 24.8557
R13656 gnd.n3372 gnd.n2457 24.8557
R13657 gnd.n3400 gnd.n3399 24.8557
R13658 gnd.n3411 gnd.n2442 24.8557
R13659 gnd.n3422 gnd.n2435 24.8557
R13660 gnd.n3421 gnd.n2423 24.8557
R13661 gnd.n3694 gnd.n3693 24.8557
R13662 gnd.n3716 gnd.n2407 24.8557
R13663 gnd.n5615 gnd.t249 24.537
R13664 gnd.t213 gnd.n1245 24.537
R13665 gnd.n7624 gnd.n238 24.537
R13666 gnd.n6542 gnd.n6541 24.2183
R13667 gnd.n6535 gnd.n983 24.2183
R13668 gnd.n4377 gnd.n986 24.2183
R13669 gnd.n4408 gnd.n997 24.2183
R13670 gnd.n4385 gnd.n1007 24.2183
R13671 gnd.n6517 gnd.n1015 24.2183
R13672 gnd.n6511 gnd.n1026 24.2183
R13673 gnd.n4426 gnd.n1029 24.2183
R13674 gnd.n4457 gnd.n1039 24.2183
R13675 gnd.n4434 gnd.n1049 24.2183
R13676 gnd.n6493 gnd.n1057 24.2183
R13677 gnd.n6487 gnd.n1068 24.2183
R13678 gnd.n4511 gnd.n1071 24.2183
R13679 gnd.n4519 gnd.n1081 24.2183
R13680 gnd.n6475 gnd.n1089 24.2183
R13681 gnd.n4528 gnd.n1092 24.2183
R13682 gnd.n6469 gnd.n1100 24.2183
R13683 gnd.n4568 gnd.n2124 24.2183
R13684 gnd.n6463 gnd.n1109 24.2183
R13685 gnd.n4652 gnd.t263 24.2183
R13686 gnd.n6218 gnd.n1338 24.2183
R13687 gnd.n6053 gnd.n6044 24.2183
R13688 gnd.n6063 gnd.n1452 24.2183
R13689 gnd.n6062 gnd.n1431 24.2183
R13690 gnd.n6074 gnd.n6073 24.2183
R13691 gnd.n1435 gnd.n1422 24.2183
R13692 gnd.n6099 gnd.n1414 24.2183
R13693 gnd.n6098 gnd.n1404 24.2183
R13694 gnd.n1407 gnd.n1394 24.2183
R13695 gnd.n6121 gnd.n1396 24.2183
R13696 gnd.n6159 gnd.n1370 24.2183
R13697 gnd.n1373 gnd.n1361 24.2183
R13698 gnd.n6189 gnd.n1364 24.2183
R13699 gnd.n7374 gnd.n402 24.2183
R13700 gnd.n6143 gnd.n390 24.2183
R13701 gnd.n7365 gnd.n384 24.2183
R13702 gnd.n7420 gnd.n370 24.2183
R13703 gnd.n7392 gnd.n377 24.2183
R13704 gnd.n7429 gnd.n358 24.2183
R13705 gnd.n5606 gnd.n1986 23.8997
R13706 gnd.n6302 gnd.n1248 23.8997
R13707 gnd.n4681 gnd.n4680 23.855
R13708 gnd.n5053 gnd.n5052 23.855
R13709 gnd.n5459 gnd.n5458 23.855
R13710 gnd.n5047 gnd.n5046 23.855
R13711 gnd.n3070 gnd.t179 23.2624
R13712 gnd.n4218 gnd.t174 23.2624
R13713 gnd.n4409 gnd.t97 23.2624
R13714 gnd.n6481 gnd.t111 23.2624
R13715 gnd.n6084 gnd.t9 23.2624
R13716 gnd.n7364 gnd.t105 23.2624
R13717 gnd.n7640 gnd.t151 23.2624
R13718 gnd.n2771 gnd.t304 22.6251
R13719 gnd.n4250 gnd.t70 22.6251
R13720 gnd.n6505 gnd.t54 22.6251
R13721 gnd.n4458 gnd.t42 22.6251
R13722 gnd.n6160 gnd.t7 22.6251
R13723 gnd.n6181 gnd.t113 22.6251
R13724 gnd.n7608 gnd.t67 22.6251
R13725 gnd.n2192 gnd.t49 22.3064
R13726 gnd.t18 gnd.n312 22.3064
R13727 gnd.n4282 gnd.t100 21.9878
R13728 gnd.n6529 gnd.t149 21.9878
R13729 gnd.n7398 gnd.t117 21.9878
R13730 gnd.n7576 gnd.t188 21.9878
R13731 gnd.n5453 gnd.n1928 21.6691
R13732 gnd.n5445 gnd.n1922 21.6691
R13733 gnd.n5424 gnd.n5423 21.6691
R13734 gnd.n5393 gnd.n5392 21.6691
R13735 gnd.n5386 gnd.n1857 21.6691
R13736 gnd.n5371 gnd.n1842 21.6691
R13737 gnd.n5335 gnd.n1806 21.6691
R13738 gnd.n5328 gnd.n1798 21.6691
R13739 gnd.n5320 gnd.n1791 21.6691
R13740 gnd.n5313 gnd.n1783 21.6691
R13741 gnd.n5276 gnd.n1739 21.6691
R13742 gnd.n5261 gnd.n1724 21.6691
R13743 gnd.n5254 gnd.n1717 21.6691
R13744 gnd.n5226 gnd.n1688 21.6691
R13745 gnd.n5219 gnd.n1680 21.6691
R13746 gnd.n5211 gnd.n1674 21.6691
R13747 gnd.n5205 gnd.n5204 21.6691
R13748 gnd.t162 gnd.n2776 21.3504
R13749 gnd.n4316 gnd.t36 21.3504
R13750 gnd.n4343 gnd.t86 21.3504
R13751 gnd.t79 gnd.n315 21.3504
R13752 gnd.t147 gnd.n334 21.3504
R13753 gnd.n4773 gnd.n1885 21.0318
R13754 gnd.n5409 gnd.n5408 21.0318
R13755 gnd.t197 gnd.n1877 21.0318
R13756 gnd.n5775 gnd.n1829 21.0318
R13757 gnd.n5783 gnd.n1819 21.0318
R13758 gnd.t83 gnd.n1813 21.0318
R13759 gnd.n5305 gnd.t29 21.0318
R13760 gnd.n5297 gnd.n1760 21.0318
R13761 gnd.n4900 gnd.n1762 21.0318
R13762 gnd.n5240 gnd.t131 21.0318
R13763 gnd.n5911 gnd.n1704 21.0318
R13764 gnd.n5919 gnd.n1694 21.0318
R13765 gnd.n5457 gnd.n5456 20.7615
R13766 gnd.n5194 gnd.n5193 20.7615
R13767 gnd.t331 gnd.n2470 20.7131
R13768 gnd.n4299 gnd.t102 20.7131
R13769 gnd.n7560 gnd.t192 20.7131
R13770 gnd.t124 gnd.n2505 20.0758
R13771 gnd.n4266 gnd.t22 20.0758
R13772 gnd.n7592 gnd.t109 20.0758
R13773 gnd.n4660 gnd.t290 19.8005
R13774 gnd.n4660 gnd.t211 19.8005
R13775 gnd.n4661 gnd.t208 19.8005
R13776 gnd.n4661 gnd.t229 19.8005
R13777 gnd.n5015 gnd.t240 19.8005
R13778 gnd.n5015 gnd.t222 19.8005
R13779 gnd.n5016 gnd.t261 19.8005
R13780 gnd.n5016 gnd.t201 19.8005
R13781 gnd.n5556 gnd.n2058 19.7572
R13782 gnd.n5422 gnd.n1891 19.7572
R13783 gnd.n4787 gnd.n1879 19.7572
R13784 gnd.n5767 gnd.n1836 19.7572
R13785 gnd.n5791 gnd.n1812 19.7572
R13786 gnd.n4887 gnd.n1768 19.7572
R13787 gnd.n4907 gnd.n1754 19.7572
R13788 gnd.n5903 gnd.n1711 19.7572
R13789 gnd.n5927 gnd.n1686 19.7572
R13790 gnd.n6295 gnd.n6294 19.7572
R13791 gnd.n4657 gnd.n4656 19.5087
R13792 gnd.n4670 gnd.n4657 19.5087
R13793 gnd.n4668 gnd.n4659 19.5087
R13794 gnd.n5020 gnd.n5014 19.5087
R13795 gnd.n3237 gnd.t333 19.4385
R13796 gnd.n4234 gnd.t156 19.4385
R13797 gnd.n1954 gnd.t311 19.4385
R13798 gnd.n5991 gnd.t307 19.4385
R13799 gnd.n7624 gnd.t119 19.4385
R13800 gnd.n5613 gnd.n1969 19.3944
R13801 gnd.n5613 gnd.n1958 19.3944
R13802 gnd.n5625 gnd.n1958 19.3944
R13803 gnd.n5625 gnd.n1956 19.3944
R13804 gnd.n5629 gnd.n1956 19.3944
R13805 gnd.n5629 gnd.n1945 19.3944
R13806 gnd.n5641 gnd.n1945 19.3944
R13807 gnd.n5641 gnd.n1943 19.3944
R13808 gnd.n5645 gnd.n1943 19.3944
R13809 gnd.n5645 gnd.n1932 19.3944
R13810 gnd.n5657 gnd.n1932 19.3944
R13811 gnd.n5657 gnd.n1930 19.3944
R13812 gnd.n5661 gnd.n1930 19.3944
R13813 gnd.n5661 gnd.n1918 19.3944
R13814 gnd.n5673 gnd.n1918 19.3944
R13815 gnd.n5673 gnd.n1916 19.3944
R13816 gnd.n5677 gnd.n1916 19.3944
R13817 gnd.n5677 gnd.n1903 19.3944
R13818 gnd.n5689 gnd.n1903 19.3944
R13819 gnd.n5689 gnd.n1901 19.3944
R13820 gnd.n5693 gnd.n1901 19.3944
R13821 gnd.n5693 gnd.n1889 19.3944
R13822 gnd.n5705 gnd.n1889 19.3944
R13823 gnd.n5705 gnd.n1887 19.3944
R13824 gnd.n5709 gnd.n1887 19.3944
R13825 gnd.n5709 gnd.n1875 19.3944
R13826 gnd.n5721 gnd.n1875 19.3944
R13827 gnd.n5721 gnd.n1873 19.3944
R13828 gnd.n5725 gnd.n1873 19.3944
R13829 gnd.n5725 gnd.n1861 19.3944
R13830 gnd.n5737 gnd.n1861 19.3944
R13831 gnd.n5737 gnd.n1859 19.3944
R13832 gnd.n5741 gnd.n1859 19.3944
R13833 gnd.n5741 gnd.n1847 19.3944
R13834 gnd.n5753 gnd.n1847 19.3944
R13835 gnd.n5753 gnd.n1845 19.3944
R13836 gnd.n5757 gnd.n1845 19.3944
R13837 gnd.n5757 gnd.n1833 19.3944
R13838 gnd.n5769 gnd.n1833 19.3944
R13839 gnd.n5769 gnd.n1831 19.3944
R13840 gnd.n5773 gnd.n1831 19.3944
R13841 gnd.n5773 gnd.n1817 19.3944
R13842 gnd.n5785 gnd.n1817 19.3944
R13843 gnd.n5785 gnd.n1815 19.3944
R13844 gnd.n5789 gnd.n1815 19.3944
R13845 gnd.n5789 gnd.n1802 19.3944
R13846 gnd.n5801 gnd.n1802 19.3944
R13847 gnd.n5801 gnd.n1800 19.3944
R13848 gnd.n5805 gnd.n1800 19.3944
R13849 gnd.n5805 gnd.n1787 19.3944
R13850 gnd.n5817 gnd.n1787 19.3944
R13851 gnd.n5817 gnd.n1785 19.3944
R13852 gnd.n5821 gnd.n1785 19.3944
R13853 gnd.n5821 gnd.n1773 19.3944
R13854 gnd.n5833 gnd.n1773 19.3944
R13855 gnd.n5833 gnd.n1771 19.3944
R13856 gnd.n5837 gnd.n1771 19.3944
R13857 gnd.n5837 gnd.n1758 19.3944
R13858 gnd.n5849 gnd.n1758 19.3944
R13859 gnd.n5849 gnd.n1756 19.3944
R13860 gnd.n5853 gnd.n1756 19.3944
R13861 gnd.n5853 gnd.n1743 19.3944
R13862 gnd.n5865 gnd.n1743 19.3944
R13863 gnd.n5865 gnd.n1741 19.3944
R13864 gnd.n5869 gnd.n1741 19.3944
R13865 gnd.n5869 gnd.n1729 19.3944
R13866 gnd.n5881 gnd.n1729 19.3944
R13867 gnd.n5881 gnd.n1727 19.3944
R13868 gnd.n5885 gnd.n1727 19.3944
R13869 gnd.n5885 gnd.n1715 19.3944
R13870 gnd.n5897 gnd.n1715 19.3944
R13871 gnd.n5897 gnd.n1713 19.3944
R13872 gnd.n5901 gnd.n1713 19.3944
R13873 gnd.n5901 gnd.n1699 19.3944
R13874 gnd.n5913 gnd.n1699 19.3944
R13875 gnd.n5913 gnd.n1697 19.3944
R13876 gnd.n5917 gnd.n1697 19.3944
R13877 gnd.n5917 gnd.n1684 19.3944
R13878 gnd.n5929 gnd.n1684 19.3944
R13879 gnd.n5929 gnd.n1682 19.3944
R13880 gnd.n5933 gnd.n1682 19.3944
R13881 gnd.n5933 gnd.n1671 19.3944
R13882 gnd.n5945 gnd.n1671 19.3944
R13883 gnd.n5945 gnd.n1669 19.3944
R13884 gnd.n5949 gnd.n1669 19.3944
R13885 gnd.n5949 gnd.n1658 19.3944
R13886 gnd.n5961 gnd.n1658 19.3944
R13887 gnd.n5961 gnd.n1656 19.3944
R13888 gnd.n5965 gnd.n1656 19.3944
R13889 gnd.n5965 gnd.n1644 19.3944
R13890 gnd.n5977 gnd.n1644 19.3944
R13891 gnd.n5977 gnd.n1642 19.3944
R13892 gnd.n5981 gnd.n1642 19.3944
R13893 gnd.n5981 gnd.n1631 19.3944
R13894 gnd.n5993 gnd.n1631 19.3944
R13895 gnd.n5993 gnd.n1628 19.3944
R13896 gnd.n5999 gnd.n1628 19.3944
R13897 gnd.n5999 gnd.n1629 19.3944
R13898 gnd.n1629 gnd.n1616 19.3944
R13899 gnd.n6015 gnd.n1616 19.3944
R13900 gnd.n6016 gnd.n6015 19.3944
R13901 gnd.n4550 gnd.n4549 19.3944
R13902 gnd.n4549 gnd.n1971 19.3944
R13903 gnd.n5609 gnd.n1971 19.3944
R13904 gnd.n5603 gnd.n5602 19.3944
R13905 gnd.n5602 gnd.n1990 19.3944
R13906 gnd.n5595 gnd.n1990 19.3944
R13907 gnd.n5595 gnd.n5594 19.3944
R13908 gnd.n5594 gnd.n2001 19.3944
R13909 gnd.n5587 gnd.n2001 19.3944
R13910 gnd.n5587 gnd.n5586 19.3944
R13911 gnd.n5586 gnd.n2009 19.3944
R13912 gnd.n5579 gnd.n2009 19.3944
R13913 gnd.n5579 gnd.n5578 19.3944
R13914 gnd.n5578 gnd.n2019 19.3944
R13915 gnd.n5571 gnd.n2019 19.3944
R13916 gnd.n5571 gnd.n5570 19.3944
R13917 gnd.n5570 gnd.n2027 19.3944
R13918 gnd.n5563 gnd.n2027 19.3944
R13919 gnd.n5563 gnd.n5562 19.3944
R13920 gnd.n5562 gnd.n2039 19.3944
R13921 gnd.n4561 gnd.n2039 19.3944
R13922 gnd.n4561 gnd.n4560 19.3944
R13923 gnd.n4560 gnd.n4559 19.3944
R13924 gnd.n4559 gnd.n4538 19.3944
R13925 gnd.n4555 gnd.n4538 19.3944
R13926 gnd.n4555 gnd.n4554 19.3944
R13927 gnd.n4554 gnd.n4553 19.3944
R13928 gnd.n2952 gnd.n2951 19.3944
R13929 gnd.n2951 gnd.n2950 19.3944
R13930 gnd.n2950 gnd.n2949 19.3944
R13931 gnd.n2949 gnd.n2947 19.3944
R13932 gnd.n2947 gnd.n2944 19.3944
R13933 gnd.n2944 gnd.n2943 19.3944
R13934 gnd.n2943 gnd.n2940 19.3944
R13935 gnd.n2940 gnd.n2939 19.3944
R13936 gnd.n2939 gnd.n2936 19.3944
R13937 gnd.n2936 gnd.n2935 19.3944
R13938 gnd.n2935 gnd.n2932 19.3944
R13939 gnd.n2932 gnd.n2931 19.3944
R13940 gnd.n2931 gnd.n2928 19.3944
R13941 gnd.n2928 gnd.n2927 19.3944
R13942 gnd.n2927 gnd.n2924 19.3944
R13943 gnd.n2924 gnd.n2923 19.3944
R13944 gnd.n2923 gnd.n2920 19.3944
R13945 gnd.n2920 gnd.n2919 19.3944
R13946 gnd.n2919 gnd.n2916 19.3944
R13947 gnd.n2916 gnd.n2915 19.3944
R13948 gnd.n2915 gnd.n2912 19.3944
R13949 gnd.n2912 gnd.n2911 19.3944
R13950 gnd.n2908 gnd.n2907 19.3944
R13951 gnd.n2907 gnd.n2863 19.3944
R13952 gnd.n2958 gnd.n2863 19.3944
R13953 gnd.n3724 gnd.n3723 19.3944
R13954 gnd.n3723 gnd.n3720 19.3944
R13955 gnd.n3720 gnd.n3719 19.3944
R13956 gnd.n3769 gnd.n3768 19.3944
R13957 gnd.n3768 gnd.n3767 19.3944
R13958 gnd.n3767 gnd.n3764 19.3944
R13959 gnd.n3764 gnd.n3763 19.3944
R13960 gnd.n3763 gnd.n3760 19.3944
R13961 gnd.n3760 gnd.n3759 19.3944
R13962 gnd.n3759 gnd.n3756 19.3944
R13963 gnd.n3756 gnd.n3755 19.3944
R13964 gnd.n3755 gnd.n3752 19.3944
R13965 gnd.n3752 gnd.n3751 19.3944
R13966 gnd.n3751 gnd.n3748 19.3944
R13967 gnd.n3748 gnd.n3747 19.3944
R13968 gnd.n3747 gnd.n3744 19.3944
R13969 gnd.n3744 gnd.n3743 19.3944
R13970 gnd.n3743 gnd.n3740 19.3944
R13971 gnd.n3740 gnd.n3739 19.3944
R13972 gnd.n3739 gnd.n3736 19.3944
R13973 gnd.n3736 gnd.n3735 19.3944
R13974 gnd.n3735 gnd.n3732 19.3944
R13975 gnd.n3732 gnd.n3731 19.3944
R13976 gnd.n3731 gnd.n3728 19.3944
R13977 gnd.n3728 gnd.n3727 19.3944
R13978 gnd.n3051 gnd.n2760 19.3944
R13979 gnd.n3061 gnd.n2760 19.3944
R13980 gnd.n3062 gnd.n3061 19.3944
R13981 gnd.n3062 gnd.n2741 19.3944
R13982 gnd.n3082 gnd.n2741 19.3944
R13983 gnd.n3082 gnd.n2733 19.3944
R13984 gnd.n3092 gnd.n2733 19.3944
R13985 gnd.n3093 gnd.n3092 19.3944
R13986 gnd.n3094 gnd.n3093 19.3944
R13987 gnd.n3094 gnd.n2716 19.3944
R13988 gnd.n3111 gnd.n2716 19.3944
R13989 gnd.n3114 gnd.n3111 19.3944
R13990 gnd.n3114 gnd.n3113 19.3944
R13991 gnd.n3113 gnd.n2689 19.3944
R13992 gnd.n3153 gnd.n2689 19.3944
R13993 gnd.n3153 gnd.n2686 19.3944
R13994 gnd.n3159 gnd.n2686 19.3944
R13995 gnd.n3160 gnd.n3159 19.3944
R13996 gnd.n3160 gnd.n2684 19.3944
R13997 gnd.n3166 gnd.n2684 19.3944
R13998 gnd.n3169 gnd.n3166 19.3944
R13999 gnd.n3171 gnd.n3169 19.3944
R14000 gnd.n3177 gnd.n3171 19.3944
R14001 gnd.n3177 gnd.n3176 19.3944
R14002 gnd.n3176 gnd.n2547 19.3944
R14003 gnd.n3243 gnd.n2547 19.3944
R14004 gnd.n3244 gnd.n3243 19.3944
R14005 gnd.n3244 gnd.n2540 19.3944
R14006 gnd.n3255 gnd.n2540 19.3944
R14007 gnd.n3256 gnd.n3255 19.3944
R14008 gnd.n3256 gnd.n2523 19.3944
R14009 gnd.n2523 gnd.n2521 19.3944
R14010 gnd.n3280 gnd.n2521 19.3944
R14011 gnd.n3281 gnd.n3280 19.3944
R14012 gnd.n3281 gnd.n2492 19.3944
R14013 gnd.n3328 gnd.n2492 19.3944
R14014 gnd.n3329 gnd.n3328 19.3944
R14015 gnd.n3329 gnd.n2485 19.3944
R14016 gnd.n3340 gnd.n2485 19.3944
R14017 gnd.n3341 gnd.n3340 19.3944
R14018 gnd.n3341 gnd.n2468 19.3944
R14019 gnd.n2468 gnd.n2466 19.3944
R14020 gnd.n3365 gnd.n2466 19.3944
R14021 gnd.n3366 gnd.n3365 19.3944
R14022 gnd.n3366 gnd.n2438 19.3944
R14023 gnd.n3417 gnd.n2438 19.3944
R14024 gnd.n3418 gnd.n3417 19.3944
R14025 gnd.n3418 gnd.n2431 19.3944
R14026 gnd.n3685 gnd.n2431 19.3944
R14027 gnd.n3686 gnd.n3685 19.3944
R14028 gnd.n3686 gnd.n2412 19.3944
R14029 gnd.n3711 gnd.n2412 19.3944
R14030 gnd.n3711 gnd.n2413 19.3944
R14031 gnd.n3042 gnd.n3041 19.3944
R14032 gnd.n3041 gnd.n2774 19.3944
R14033 gnd.n2797 gnd.n2774 19.3944
R14034 gnd.n2800 gnd.n2797 19.3944
R14035 gnd.n2800 gnd.n2793 19.3944
R14036 gnd.n2804 gnd.n2793 19.3944
R14037 gnd.n2807 gnd.n2804 19.3944
R14038 gnd.n2810 gnd.n2807 19.3944
R14039 gnd.n2810 gnd.n2791 19.3944
R14040 gnd.n2814 gnd.n2791 19.3944
R14041 gnd.n2817 gnd.n2814 19.3944
R14042 gnd.n2820 gnd.n2817 19.3944
R14043 gnd.n2820 gnd.n2789 19.3944
R14044 gnd.n2824 gnd.n2789 19.3944
R14045 gnd.n3047 gnd.n3046 19.3944
R14046 gnd.n3046 gnd.n2750 19.3944
R14047 gnd.n3072 gnd.n2750 19.3944
R14048 gnd.n3072 gnd.n2748 19.3944
R14049 gnd.n3078 gnd.n2748 19.3944
R14050 gnd.n3078 gnd.n3077 19.3944
R14051 gnd.n3077 gnd.n2722 19.3944
R14052 gnd.n3102 gnd.n2722 19.3944
R14053 gnd.n3102 gnd.n2720 19.3944
R14054 gnd.n3106 gnd.n2720 19.3944
R14055 gnd.n3106 gnd.n2700 19.3944
R14056 gnd.n3133 gnd.n2700 19.3944
R14057 gnd.n3133 gnd.n2698 19.3944
R14058 gnd.n3143 gnd.n2698 19.3944
R14059 gnd.n3143 gnd.n3142 19.3944
R14060 gnd.n3142 gnd.n3141 19.3944
R14061 gnd.n3141 gnd.n2647 19.3944
R14062 gnd.n3191 gnd.n2647 19.3944
R14063 gnd.n3191 gnd.n3190 19.3944
R14064 gnd.n3190 gnd.n3189 19.3944
R14065 gnd.n3189 gnd.n2651 19.3944
R14066 gnd.n2671 gnd.n2651 19.3944
R14067 gnd.n2671 gnd.n2557 19.3944
R14068 gnd.n3228 gnd.n2557 19.3944
R14069 gnd.n3228 gnd.n2555 19.3944
R14070 gnd.n3234 gnd.n2555 19.3944
R14071 gnd.n3234 gnd.n3233 19.3944
R14072 gnd.n3233 gnd.n2530 19.3944
R14073 gnd.n3268 gnd.n2530 19.3944
R14074 gnd.n3268 gnd.n2528 19.3944
R14075 gnd.n3274 gnd.n2528 19.3944
R14076 gnd.n3274 gnd.n3273 19.3944
R14077 gnd.n3273 gnd.n2503 19.3944
R14078 gnd.n3313 gnd.n2503 19.3944
R14079 gnd.n3313 gnd.n2501 19.3944
R14080 gnd.n3319 gnd.n2501 19.3944
R14081 gnd.n3319 gnd.n3318 19.3944
R14082 gnd.n3318 gnd.n2475 19.3944
R14083 gnd.n3353 gnd.n2475 19.3944
R14084 gnd.n3353 gnd.n2473 19.3944
R14085 gnd.n3359 gnd.n2473 19.3944
R14086 gnd.n3359 gnd.n3358 19.3944
R14087 gnd.n3358 gnd.n2448 19.3944
R14088 gnd.n3402 gnd.n2448 19.3944
R14089 gnd.n3402 gnd.n2446 19.3944
R14090 gnd.n3408 gnd.n2446 19.3944
R14091 gnd.n3408 gnd.n3407 19.3944
R14092 gnd.n3407 gnd.n2421 19.3944
R14093 gnd.n3696 gnd.n2421 19.3944
R14094 gnd.n3696 gnd.n2419 19.3944
R14095 gnd.n3704 gnd.n2419 19.3944
R14096 gnd.n3704 gnd.n3703 19.3944
R14097 gnd.n3703 gnd.n3702 19.3944
R14098 gnd.n3805 gnd.n3804 19.3944
R14099 gnd.n3804 gnd.n2359 19.3944
R14100 gnd.n3800 gnd.n2359 19.3944
R14101 gnd.n3800 gnd.n3797 19.3944
R14102 gnd.n3797 gnd.n3794 19.3944
R14103 gnd.n3794 gnd.n3793 19.3944
R14104 gnd.n3793 gnd.n3790 19.3944
R14105 gnd.n3790 gnd.n3789 19.3944
R14106 gnd.n3789 gnd.n3786 19.3944
R14107 gnd.n3786 gnd.n3785 19.3944
R14108 gnd.n3785 gnd.n3782 19.3944
R14109 gnd.n3782 gnd.n3781 19.3944
R14110 gnd.n3781 gnd.n3778 19.3944
R14111 gnd.n3778 gnd.n3777 19.3944
R14112 gnd.n2962 gnd.n2861 19.3944
R14113 gnd.n2962 gnd.n2852 19.3944
R14114 gnd.n2975 gnd.n2852 19.3944
R14115 gnd.n2975 gnd.n2850 19.3944
R14116 gnd.n2979 gnd.n2850 19.3944
R14117 gnd.n2979 gnd.n2840 19.3944
R14118 gnd.n2991 gnd.n2840 19.3944
R14119 gnd.n2991 gnd.n2838 19.3944
R14120 gnd.n3025 gnd.n2838 19.3944
R14121 gnd.n3025 gnd.n3024 19.3944
R14122 gnd.n3024 gnd.n3023 19.3944
R14123 gnd.n3023 gnd.n3022 19.3944
R14124 gnd.n3022 gnd.n3019 19.3944
R14125 gnd.n3019 gnd.n3018 19.3944
R14126 gnd.n3018 gnd.n3017 19.3944
R14127 gnd.n3017 gnd.n3015 19.3944
R14128 gnd.n3015 gnd.n3014 19.3944
R14129 gnd.n3014 gnd.n3011 19.3944
R14130 gnd.n3011 gnd.n3010 19.3944
R14131 gnd.n3010 gnd.n3009 19.3944
R14132 gnd.n3009 gnd.n3007 19.3944
R14133 gnd.n3007 gnd.n2706 19.3944
R14134 gnd.n3122 gnd.n2706 19.3944
R14135 gnd.n3122 gnd.n2704 19.3944
R14136 gnd.n3128 gnd.n2704 19.3944
R14137 gnd.n3128 gnd.n3127 19.3944
R14138 gnd.n3127 gnd.n2628 19.3944
R14139 gnd.n3202 gnd.n2628 19.3944
R14140 gnd.n3202 gnd.n2629 19.3944
R14141 gnd.n2676 gnd.n2675 19.3944
R14142 gnd.n2679 gnd.n2678 19.3944
R14143 gnd.n2666 gnd.n2665 19.3944
R14144 gnd.n3221 gnd.n2562 19.3944
R14145 gnd.n3221 gnd.n3220 19.3944
R14146 gnd.n3220 gnd.n3219 19.3944
R14147 gnd.n3219 gnd.n3217 19.3944
R14148 gnd.n3217 gnd.n3216 19.3944
R14149 gnd.n3216 gnd.n3214 19.3944
R14150 gnd.n3214 gnd.n3213 19.3944
R14151 gnd.n3213 gnd.n2511 19.3944
R14152 gnd.n3289 gnd.n2511 19.3944
R14153 gnd.n3289 gnd.n2509 19.3944
R14154 gnd.n3308 gnd.n2509 19.3944
R14155 gnd.n3308 gnd.n3307 19.3944
R14156 gnd.n3307 gnd.n3306 19.3944
R14157 gnd.n3306 gnd.n3304 19.3944
R14158 gnd.n3304 gnd.n3303 19.3944
R14159 gnd.n3303 gnd.n3301 19.3944
R14160 gnd.n3301 gnd.n3300 19.3944
R14161 gnd.n3300 gnd.n2455 19.3944
R14162 gnd.n3374 gnd.n2455 19.3944
R14163 gnd.n3374 gnd.n2453 19.3944
R14164 gnd.n3397 gnd.n2453 19.3944
R14165 gnd.n3397 gnd.n3396 19.3944
R14166 gnd.n3396 gnd.n3395 19.3944
R14167 gnd.n3395 gnd.n3392 19.3944
R14168 gnd.n3392 gnd.n3391 19.3944
R14169 gnd.n3391 gnd.n3389 19.3944
R14170 gnd.n3389 gnd.n3388 19.3944
R14171 gnd.n3388 gnd.n3386 19.3944
R14172 gnd.n3386 gnd.n2406 19.3944
R14173 gnd.n2967 gnd.n2857 19.3944
R14174 gnd.n2967 gnd.n2855 19.3944
R14175 gnd.n2971 gnd.n2855 19.3944
R14176 gnd.n2971 gnd.n2846 19.3944
R14177 gnd.n2983 gnd.n2846 19.3944
R14178 gnd.n2983 gnd.n2844 19.3944
R14179 gnd.n2987 gnd.n2844 19.3944
R14180 gnd.n2987 gnd.n2833 19.3944
R14181 gnd.n3029 gnd.n2833 19.3944
R14182 gnd.n3029 gnd.n2787 19.3944
R14183 gnd.n3035 gnd.n2787 19.3944
R14184 gnd.n3035 gnd.n3034 19.3944
R14185 gnd.n3034 gnd.n2765 19.3944
R14186 gnd.n3056 gnd.n2765 19.3944
R14187 gnd.n3056 gnd.n2758 19.3944
R14188 gnd.n3067 gnd.n2758 19.3944
R14189 gnd.n3067 gnd.n3066 19.3944
R14190 gnd.n3066 gnd.n2739 19.3944
R14191 gnd.n3087 gnd.n2739 19.3944
R14192 gnd.n3087 gnd.n2729 19.3944
R14193 gnd.n3097 gnd.n2729 19.3944
R14194 gnd.n3097 gnd.n2712 19.3944
R14195 gnd.n3118 gnd.n2712 19.3944
R14196 gnd.n3118 gnd.n3117 19.3944
R14197 gnd.n3117 gnd.n2691 19.3944
R14198 gnd.n3148 gnd.n2691 19.3944
R14199 gnd.n3148 gnd.n2636 19.3944
R14200 gnd.n3198 gnd.n2636 19.3944
R14201 gnd.n3198 gnd.n3197 19.3944
R14202 gnd.n3197 gnd.n3196 19.3944
R14203 gnd.n3196 gnd.n2640 19.3944
R14204 gnd.n2658 gnd.n2640 19.3944
R14205 gnd.n3184 gnd.n2658 19.3944
R14206 gnd.n3184 gnd.n3183 19.3944
R14207 gnd.n3183 gnd.n3182 19.3944
R14208 gnd.n3182 gnd.n2662 19.3944
R14209 gnd.n2662 gnd.n2549 19.3944
R14210 gnd.n3239 gnd.n2549 19.3944
R14211 gnd.n3239 gnd.n2542 19.3944
R14212 gnd.n3250 gnd.n2542 19.3944
R14213 gnd.n3250 gnd.n2538 19.3944
R14214 gnd.n3263 gnd.n2538 19.3944
R14215 gnd.n3263 gnd.n3262 19.3944
R14216 gnd.n3262 gnd.n2517 19.3944
R14217 gnd.n3285 gnd.n2517 19.3944
R14218 gnd.n3285 gnd.n3284 19.3944
R14219 gnd.n3284 gnd.n2494 19.3944
R14220 gnd.n3324 gnd.n2494 19.3944
R14221 gnd.n3324 gnd.n2487 19.3944
R14222 gnd.n3335 gnd.n2487 19.3944
R14223 gnd.n3335 gnd.n2483 19.3944
R14224 gnd.n3348 gnd.n2483 19.3944
R14225 gnd.n3348 gnd.n3347 19.3944
R14226 gnd.n3347 gnd.n2462 19.3944
R14227 gnd.n3370 gnd.n2462 19.3944
R14228 gnd.n3370 gnd.n3369 19.3944
R14229 gnd.n3369 gnd.n2440 19.3944
R14230 gnd.n3413 gnd.n2440 19.3944
R14231 gnd.n3413 gnd.n2433 19.3944
R14232 gnd.n3424 gnd.n2433 19.3944
R14233 gnd.n3424 gnd.n2429 19.3944
R14234 gnd.n3691 gnd.n2429 19.3944
R14235 gnd.n3691 gnd.n3690 19.3944
R14236 gnd.n3690 gnd.n2410 19.3944
R14237 gnd.n3714 gnd.n2410 19.3944
R14238 gnd.n6055 gnd.n6043 19.3944
R14239 gnd.n6055 gnd.n1476 19.3944
R14240 gnd.n6060 gnd.n1476 19.3944
R14241 gnd.n6060 gnd.n1477 19.3944
R14242 gnd.n1477 gnd.n1420 19.3944
R14243 gnd.n6086 gnd.n1420 19.3944
R14244 gnd.n6086 gnd.n1417 19.3944
R14245 gnd.n6096 gnd.n1417 19.3944
R14246 gnd.n6096 gnd.n1418 19.3944
R14247 gnd.n6092 gnd.n1418 19.3944
R14248 gnd.n6092 gnd.n6091 19.3944
R14249 gnd.n6091 gnd.n1382 19.3944
R14250 gnd.n6156 gnd.n1382 19.3944
R14251 gnd.n6156 gnd.n1383 19.3944
R14252 gnd.n6152 gnd.n1383 19.3944
R14253 gnd.n6152 gnd.n6151 19.3944
R14254 gnd.n6151 gnd.n6150 19.3944
R14255 gnd.n6150 gnd.n6140 19.3944
R14256 gnd.n6146 gnd.n6140 19.3944
R14257 gnd.n6146 gnd.n6145 19.3944
R14258 gnd.n6145 gnd.n382 19.3944
R14259 gnd.n7400 gnd.n382 19.3944
R14260 gnd.n7401 gnd.n7400 19.3944
R14261 gnd.n7401 gnd.n379 19.3944
R14262 gnd.n7406 gnd.n379 19.3944
R14263 gnd.n7406 gnd.n380 19.3944
R14264 gnd.n380 gnd.n348 19.3944
R14265 gnd.n7446 gnd.n348 19.3944
R14266 gnd.n7446 gnd.n346 19.3944
R14267 gnd.n7450 gnd.n346 19.3944
R14268 gnd.n7451 gnd.n7450 19.3944
R14269 gnd.n7451 gnd.n80 19.3944
R14270 gnd.n7855 gnd.n80 19.3944
R14271 gnd.n7855 gnd.n7854 19.3944
R14272 gnd.n7854 gnd.n7853 19.3944
R14273 gnd.n7853 gnd.n85 19.3944
R14274 gnd.n7849 gnd.n85 19.3944
R14275 gnd.n7849 gnd.n7848 19.3944
R14276 gnd.n7848 gnd.n7847 19.3944
R14277 gnd.n7847 gnd.n90 19.3944
R14278 gnd.n7843 gnd.n90 19.3944
R14279 gnd.n7843 gnd.n7842 19.3944
R14280 gnd.n7842 gnd.n7841 19.3944
R14281 gnd.n7841 gnd.n95 19.3944
R14282 gnd.n7837 gnd.n95 19.3944
R14283 gnd.n7837 gnd.n7836 19.3944
R14284 gnd.n7836 gnd.n7835 19.3944
R14285 gnd.n7835 gnd.n100 19.3944
R14286 gnd.n7831 gnd.n100 19.3944
R14287 gnd.n7831 gnd.n7830 19.3944
R14288 gnd.n7830 gnd.n7829 19.3944
R14289 gnd.n7829 gnd.n105 19.3944
R14290 gnd.n7825 gnd.n105 19.3944
R14291 gnd.n7825 gnd.n7824 19.3944
R14292 gnd.n7824 gnd.n7823 19.3944
R14293 gnd.n7823 gnd.n110 19.3944
R14294 gnd.n7819 gnd.n110 19.3944
R14295 gnd.n7819 gnd.n7818 19.3944
R14296 gnd.n7818 gnd.n7817 19.3944
R14297 gnd.n7817 gnd.n115 19.3944
R14298 gnd.n7813 gnd.n115 19.3944
R14299 gnd.n7813 gnd.n7812 19.3944
R14300 gnd.n7812 gnd.n7811 19.3944
R14301 gnd.n7811 gnd.n120 19.3944
R14302 gnd.n7705 gnd.n7704 19.3944
R14303 gnd.n7704 gnd.n7703 19.3944
R14304 gnd.n7703 gnd.n7652 19.3944
R14305 gnd.n7699 gnd.n7652 19.3944
R14306 gnd.n7699 gnd.n7698 19.3944
R14307 gnd.n7698 gnd.n7697 19.3944
R14308 gnd.n7697 gnd.n7660 19.3944
R14309 gnd.n7693 gnd.n7660 19.3944
R14310 gnd.n7693 gnd.n7692 19.3944
R14311 gnd.n7692 gnd.n7691 19.3944
R14312 gnd.n7691 gnd.n7668 19.3944
R14313 gnd.n7687 gnd.n7668 19.3944
R14314 gnd.n7687 gnd.n7686 19.3944
R14315 gnd.n7686 gnd.n7685 19.3944
R14316 gnd.n7685 gnd.n7676 19.3944
R14317 gnd.n7681 gnd.n7676 19.3944
R14318 gnd.n1521 gnd.n1517 19.3944
R14319 gnd.n1524 gnd.n1521 19.3944
R14320 gnd.n1527 gnd.n1524 19.3944
R14321 gnd.n1527 gnd.n1510 19.3944
R14322 gnd.n1540 gnd.n1510 19.3944
R14323 gnd.n1543 gnd.n1540 19.3944
R14324 gnd.n1546 gnd.n1543 19.3944
R14325 gnd.n1546 gnd.n1503 19.3944
R14326 gnd.n1559 gnd.n1503 19.3944
R14327 gnd.n1562 gnd.n1559 19.3944
R14328 gnd.n1565 gnd.n1562 19.3944
R14329 gnd.n1565 gnd.n1496 19.3944
R14330 gnd.n1577 gnd.n1496 19.3944
R14331 gnd.n1580 gnd.n1577 19.3944
R14332 gnd.n1580 gnd.n1488 19.3944
R14333 gnd.n1593 gnd.n1488 19.3944
R14334 gnd.n6216 gnd.n1341 19.3944
R14335 gnd.n6212 gnd.n1341 19.3944
R14336 gnd.n6212 gnd.n6211 19.3944
R14337 gnd.n6211 gnd.n6210 19.3944
R14338 gnd.n6210 gnd.n1347 19.3944
R14339 gnd.n6206 gnd.n1347 19.3944
R14340 gnd.n6206 gnd.n6205 19.3944
R14341 gnd.n6205 gnd.n6204 19.3944
R14342 gnd.n6204 gnd.n1352 19.3944
R14343 gnd.n6200 gnd.n1352 19.3944
R14344 gnd.n6200 gnd.n6199 19.3944
R14345 gnd.n6199 gnd.n6198 19.3944
R14346 gnd.n6198 gnd.n1357 19.3944
R14347 gnd.n6194 gnd.n1357 19.3944
R14348 gnd.n6194 gnd.n6193 19.3944
R14349 gnd.n6193 gnd.n6192 19.3944
R14350 gnd.n6192 gnd.n405 19.3944
R14351 gnd.n7372 gnd.n405 19.3944
R14352 gnd.n7372 gnd.n406 19.3944
R14353 gnd.n7368 gnd.n406 19.3944
R14354 gnd.n7368 gnd.n7367 19.3944
R14355 gnd.n7367 gnd.n373 19.3944
R14356 gnd.n7418 gnd.n373 19.3944
R14357 gnd.n7418 gnd.n374 19.3944
R14358 gnd.n7414 gnd.n374 19.3944
R14359 gnd.n7414 gnd.n7413 19.3944
R14360 gnd.n7413 gnd.n7412 19.3944
R14361 gnd.n7412 gnd.n318 19.3944
R14362 gnd.n7549 gnd.n318 19.3944
R14363 gnd.n7549 gnd.n319 19.3944
R14364 gnd.n7545 gnd.n319 19.3944
R14365 gnd.n7545 gnd.n7544 19.3944
R14366 gnd.n7544 gnd.n7543 19.3944
R14367 gnd.n7543 gnd.n325 19.3944
R14368 gnd.n7539 gnd.n325 19.3944
R14369 gnd.n7539 gnd.n7538 19.3944
R14370 gnd.n7538 gnd.n297 19.3944
R14371 gnd.n7562 gnd.n297 19.3944
R14372 gnd.n7562 gnd.n295 19.3944
R14373 gnd.n7566 gnd.n295 19.3944
R14374 gnd.n7566 gnd.n281 19.3944
R14375 gnd.n7578 gnd.n281 19.3944
R14376 gnd.n7578 gnd.n279 19.3944
R14377 gnd.n7582 gnd.n279 19.3944
R14378 gnd.n7582 gnd.n267 19.3944
R14379 gnd.n7594 gnd.n267 19.3944
R14380 gnd.n7594 gnd.n265 19.3944
R14381 gnd.n7598 gnd.n265 19.3944
R14382 gnd.n7598 gnd.n251 19.3944
R14383 gnd.n7610 gnd.n251 19.3944
R14384 gnd.n7610 gnd.n249 19.3944
R14385 gnd.n7614 gnd.n249 19.3944
R14386 gnd.n7614 gnd.n236 19.3944
R14387 gnd.n7626 gnd.n236 19.3944
R14388 gnd.n7626 gnd.n234 19.3944
R14389 gnd.n7630 gnd.n234 19.3944
R14390 gnd.n7630 gnd.n221 19.3944
R14391 gnd.n7642 gnd.n221 19.3944
R14392 gnd.n7642 gnd.n218 19.3944
R14393 gnd.n7714 gnd.n218 19.3944
R14394 gnd.n7714 gnd.n219 19.3944
R14395 gnd.n7710 gnd.n219 19.3944
R14396 gnd.n7710 gnd.n7709 19.3944
R14397 gnd.n7709 gnd.n7708 19.3944
R14398 gnd.n2043 gnd.n1115 19.3944
R14399 gnd.n2043 gnd.n1993 19.3944
R14400 gnd.n5599 gnd.n1993 19.3944
R14401 gnd.n5599 gnd.n5598 19.3944
R14402 gnd.n5598 gnd.n1996 19.3944
R14403 gnd.n5591 gnd.n1996 19.3944
R14404 gnd.n5591 gnd.n5590 19.3944
R14405 gnd.n5590 gnd.n2005 19.3944
R14406 gnd.n5583 gnd.n2005 19.3944
R14407 gnd.n5583 gnd.n5582 19.3944
R14408 gnd.n5582 gnd.n2013 19.3944
R14409 gnd.n5575 gnd.n2013 19.3944
R14410 gnd.n5575 gnd.n5574 19.3944
R14411 gnd.n5574 gnd.n2023 19.3944
R14412 gnd.n5567 gnd.n2023 19.3944
R14413 gnd.n5567 gnd.n5566 19.3944
R14414 gnd.n6544 gnd.n968 19.3944
R14415 gnd.n4370 gnd.n968 19.3944
R14416 gnd.n4370 gnd.n4368 19.3944
R14417 gnd.n4374 gnd.n4368 19.3944
R14418 gnd.n4374 gnd.n2165 19.3944
R14419 gnd.n4411 gnd.n2165 19.3944
R14420 gnd.n4411 gnd.n2163 19.3944
R14421 gnd.n4415 gnd.n2163 19.3944
R14422 gnd.n4415 gnd.n2161 19.3944
R14423 gnd.n4419 gnd.n2161 19.3944
R14424 gnd.n4419 gnd.n2159 19.3944
R14425 gnd.n4423 gnd.n2159 19.3944
R14426 gnd.n4423 gnd.n2144 19.3944
R14427 gnd.n4460 gnd.n2144 19.3944
R14428 gnd.n4460 gnd.n2142 19.3944
R14429 gnd.n4464 gnd.n2142 19.3944
R14430 gnd.n4464 gnd.n2140 19.3944
R14431 gnd.n4468 gnd.n2140 19.3944
R14432 gnd.n4468 gnd.n2138 19.3944
R14433 gnd.n4508 gnd.n2138 19.3944
R14434 gnd.n4508 gnd.n4507 19.3944
R14435 gnd.n4507 gnd.n4506 19.3944
R14436 gnd.n4506 gnd.n4474 19.3944
R14437 gnd.n4502 gnd.n4474 19.3944
R14438 gnd.n4502 gnd.n4501 19.3944
R14439 gnd.n4501 gnd.n4500 19.3944
R14440 gnd.n4500 gnd.n4480 19.3944
R14441 gnd.n4496 gnd.n4480 19.3944
R14442 gnd.n4496 gnd.n4495 19.3944
R14443 gnd.n4495 gnd.n4494 19.3944
R14444 gnd.n4494 gnd.n4486 19.3944
R14445 gnd.n4489 gnd.n4486 19.3944
R14446 gnd.n4489 gnd.n1965 19.3944
R14447 gnd.n5617 gnd.n1965 19.3944
R14448 gnd.n5617 gnd.n1963 19.3944
R14449 gnd.n5621 gnd.n1963 19.3944
R14450 gnd.n5621 gnd.n1951 19.3944
R14451 gnd.n5633 gnd.n1951 19.3944
R14452 gnd.n5633 gnd.n1949 19.3944
R14453 gnd.n5637 gnd.n1949 19.3944
R14454 gnd.n5637 gnd.n1939 19.3944
R14455 gnd.n5649 gnd.n1939 19.3944
R14456 gnd.n5649 gnd.n1937 19.3944
R14457 gnd.n5653 gnd.n1937 19.3944
R14458 gnd.n5653 gnd.n1926 19.3944
R14459 gnd.n5665 gnd.n1926 19.3944
R14460 gnd.n5665 gnd.n1924 19.3944
R14461 gnd.n5669 gnd.n1924 19.3944
R14462 gnd.n5669 gnd.n1911 19.3944
R14463 gnd.n5681 gnd.n1911 19.3944
R14464 gnd.n5681 gnd.n1909 19.3944
R14465 gnd.n5685 gnd.n1909 19.3944
R14466 gnd.n5685 gnd.n1897 19.3944
R14467 gnd.n5697 gnd.n1897 19.3944
R14468 gnd.n5697 gnd.n1895 19.3944
R14469 gnd.n5701 gnd.n1895 19.3944
R14470 gnd.n5701 gnd.n1883 19.3944
R14471 gnd.n5713 gnd.n1883 19.3944
R14472 gnd.n5713 gnd.n1881 19.3944
R14473 gnd.n5717 gnd.n1881 19.3944
R14474 gnd.n5717 gnd.n1868 19.3944
R14475 gnd.n5729 gnd.n1868 19.3944
R14476 gnd.n5729 gnd.n1866 19.3944
R14477 gnd.n5733 gnd.n1866 19.3944
R14478 gnd.n5733 gnd.n1855 19.3944
R14479 gnd.n5745 gnd.n1855 19.3944
R14480 gnd.n5745 gnd.n1853 19.3944
R14481 gnd.n5749 gnd.n1853 19.3944
R14482 gnd.n5749 gnd.n1840 19.3944
R14483 gnd.n5761 gnd.n1840 19.3944
R14484 gnd.n5761 gnd.n1838 19.3944
R14485 gnd.n5765 gnd.n1838 19.3944
R14486 gnd.n5765 gnd.n1825 19.3944
R14487 gnd.n5777 gnd.n1825 19.3944
R14488 gnd.n5777 gnd.n1823 19.3944
R14489 gnd.n5781 gnd.n1823 19.3944
R14490 gnd.n5781 gnd.n1810 19.3944
R14491 gnd.n5793 gnd.n1810 19.3944
R14492 gnd.n5793 gnd.n1808 19.3944
R14493 gnd.n5797 gnd.n1808 19.3944
R14494 gnd.n5797 gnd.n1795 19.3944
R14495 gnd.n5809 gnd.n1795 19.3944
R14496 gnd.n5809 gnd.n1793 19.3944
R14497 gnd.n5813 gnd.n1793 19.3944
R14498 gnd.n5813 gnd.n1781 19.3944
R14499 gnd.n5825 gnd.n1781 19.3944
R14500 gnd.n5825 gnd.n1779 19.3944
R14501 gnd.n5829 gnd.n1779 19.3944
R14502 gnd.n5829 gnd.n1766 19.3944
R14503 gnd.n5841 gnd.n1766 19.3944
R14504 gnd.n5841 gnd.n1764 19.3944
R14505 gnd.n5845 gnd.n1764 19.3944
R14506 gnd.n5845 gnd.n1751 19.3944
R14507 gnd.n5857 gnd.n1751 19.3944
R14508 gnd.n5857 gnd.n1749 19.3944
R14509 gnd.n5861 gnd.n1749 19.3944
R14510 gnd.n5861 gnd.n1737 19.3944
R14511 gnd.n5873 gnd.n1737 19.3944
R14512 gnd.n5873 gnd.n1735 19.3944
R14513 gnd.n5877 gnd.n1735 19.3944
R14514 gnd.n5877 gnd.n1722 19.3944
R14515 gnd.n5889 gnd.n1722 19.3944
R14516 gnd.n5889 gnd.n1720 19.3944
R14517 gnd.n5893 gnd.n1720 19.3944
R14518 gnd.n5893 gnd.n1708 19.3944
R14519 gnd.n5905 gnd.n1708 19.3944
R14520 gnd.n5905 gnd.n1706 19.3944
R14521 gnd.n5909 gnd.n1706 19.3944
R14522 gnd.n5909 gnd.n1692 19.3944
R14523 gnd.n5921 gnd.n1692 19.3944
R14524 gnd.n5921 gnd.n1690 19.3944
R14525 gnd.n5925 gnd.n1690 19.3944
R14526 gnd.n5925 gnd.n1678 19.3944
R14527 gnd.n5937 gnd.n1678 19.3944
R14528 gnd.n5937 gnd.n1676 19.3944
R14529 gnd.n5941 gnd.n1676 19.3944
R14530 gnd.n5941 gnd.n1666 19.3944
R14531 gnd.n5953 gnd.n1666 19.3944
R14532 gnd.n5953 gnd.n1664 19.3944
R14533 gnd.n5957 gnd.n1664 19.3944
R14534 gnd.n5957 gnd.n1651 19.3944
R14535 gnd.n5969 gnd.n1651 19.3944
R14536 gnd.n5969 gnd.n1649 19.3944
R14537 gnd.n5973 gnd.n1649 19.3944
R14538 gnd.n5973 gnd.n1637 19.3944
R14539 gnd.n5985 gnd.n1637 19.3944
R14540 gnd.n5985 gnd.n1635 19.3944
R14541 gnd.n5989 gnd.n1635 19.3944
R14542 gnd.n5989 gnd.n1624 19.3944
R14543 gnd.n6003 gnd.n1624 19.3944
R14544 gnd.n6003 gnd.n1622 19.3944
R14545 gnd.n6010 gnd.n1622 19.3944
R14546 gnd.n6010 gnd.n6009 19.3944
R14547 gnd.n6009 gnd.n1250 19.3944
R14548 gnd.n6300 gnd.n1250 19.3944
R14549 gnd.n6300 gnd.n6299 19.3944
R14550 gnd.n6299 gnd.n6298 19.3944
R14551 gnd.n6298 gnd.n1254 19.3944
R14552 gnd.n1445 gnd.n1254 19.3944
R14553 gnd.n1445 gnd.n1442 19.3944
R14554 gnd.n1449 gnd.n1442 19.3944
R14555 gnd.n1449 gnd.n1440 19.3944
R14556 gnd.n6065 gnd.n1440 19.3944
R14557 gnd.n6065 gnd.n1438 19.3944
R14558 gnd.n6071 gnd.n1438 19.3944
R14559 gnd.n6071 gnd.n6070 19.3944
R14560 gnd.n6070 gnd.n1412 19.3944
R14561 gnd.n6101 gnd.n1412 19.3944
R14562 gnd.n6101 gnd.n1410 19.3944
R14563 gnd.n6107 gnd.n1410 19.3944
R14564 gnd.n6107 gnd.n6106 19.3944
R14565 gnd.n6106 gnd.n1378 19.3944
R14566 gnd.n6162 gnd.n1378 19.3944
R14567 gnd.n6162 gnd.n1376 19.3944
R14568 gnd.n6178 gnd.n1376 19.3944
R14569 gnd.n6178 gnd.n6177 19.3944
R14570 gnd.n6177 gnd.n6176 19.3944
R14571 gnd.n6176 gnd.n6168 19.3944
R14572 gnd.n6172 gnd.n6168 19.3944
R14573 gnd.n6172 gnd.n411 19.3944
R14574 gnd.n7362 gnd.n411 19.3944
R14575 gnd.n7362 gnd.n7361 19.3944
R14576 gnd.n7361 gnd.n7360 19.3944
R14577 gnd.n7360 gnd.n415 19.3944
R14578 gnd.n7356 gnd.n415 19.3944
R14579 gnd.n7356 gnd.n7355 19.3944
R14580 gnd.n7355 gnd.n7354 19.3944
R14581 gnd.n7140 gnd.n544 19.3944
R14582 gnd.n7146 gnd.n544 19.3944
R14583 gnd.n7146 gnd.n542 19.3944
R14584 gnd.n7150 gnd.n542 19.3944
R14585 gnd.n7150 gnd.n538 19.3944
R14586 gnd.n7156 gnd.n538 19.3944
R14587 gnd.n7156 gnd.n536 19.3944
R14588 gnd.n7160 gnd.n536 19.3944
R14589 gnd.n7160 gnd.n532 19.3944
R14590 gnd.n7166 gnd.n532 19.3944
R14591 gnd.n7166 gnd.n530 19.3944
R14592 gnd.n7170 gnd.n530 19.3944
R14593 gnd.n7170 gnd.n526 19.3944
R14594 gnd.n7176 gnd.n526 19.3944
R14595 gnd.n7176 gnd.n524 19.3944
R14596 gnd.n7180 gnd.n524 19.3944
R14597 gnd.n7180 gnd.n520 19.3944
R14598 gnd.n7186 gnd.n520 19.3944
R14599 gnd.n7186 gnd.n518 19.3944
R14600 gnd.n7190 gnd.n518 19.3944
R14601 gnd.n7190 gnd.n514 19.3944
R14602 gnd.n7196 gnd.n514 19.3944
R14603 gnd.n7196 gnd.n512 19.3944
R14604 gnd.n7200 gnd.n512 19.3944
R14605 gnd.n7200 gnd.n508 19.3944
R14606 gnd.n7206 gnd.n508 19.3944
R14607 gnd.n7206 gnd.n506 19.3944
R14608 gnd.n7210 gnd.n506 19.3944
R14609 gnd.n7210 gnd.n502 19.3944
R14610 gnd.n7216 gnd.n502 19.3944
R14611 gnd.n7216 gnd.n500 19.3944
R14612 gnd.n7220 gnd.n500 19.3944
R14613 gnd.n7220 gnd.n496 19.3944
R14614 gnd.n7226 gnd.n496 19.3944
R14615 gnd.n7226 gnd.n494 19.3944
R14616 gnd.n7230 gnd.n494 19.3944
R14617 gnd.n7230 gnd.n490 19.3944
R14618 gnd.n7236 gnd.n490 19.3944
R14619 gnd.n7236 gnd.n488 19.3944
R14620 gnd.n7240 gnd.n488 19.3944
R14621 gnd.n7240 gnd.n484 19.3944
R14622 gnd.n7246 gnd.n484 19.3944
R14623 gnd.n7246 gnd.n482 19.3944
R14624 gnd.n7250 gnd.n482 19.3944
R14625 gnd.n7250 gnd.n478 19.3944
R14626 gnd.n7256 gnd.n478 19.3944
R14627 gnd.n7256 gnd.n476 19.3944
R14628 gnd.n7260 gnd.n476 19.3944
R14629 gnd.n7260 gnd.n472 19.3944
R14630 gnd.n7266 gnd.n472 19.3944
R14631 gnd.n7266 gnd.n470 19.3944
R14632 gnd.n7270 gnd.n470 19.3944
R14633 gnd.n7270 gnd.n466 19.3944
R14634 gnd.n7276 gnd.n466 19.3944
R14635 gnd.n7276 gnd.n464 19.3944
R14636 gnd.n7280 gnd.n464 19.3944
R14637 gnd.n7280 gnd.n460 19.3944
R14638 gnd.n7286 gnd.n460 19.3944
R14639 gnd.n7286 gnd.n458 19.3944
R14640 gnd.n7290 gnd.n458 19.3944
R14641 gnd.n7290 gnd.n454 19.3944
R14642 gnd.n7296 gnd.n454 19.3944
R14643 gnd.n7296 gnd.n452 19.3944
R14644 gnd.n7300 gnd.n452 19.3944
R14645 gnd.n7300 gnd.n448 19.3944
R14646 gnd.n7306 gnd.n448 19.3944
R14647 gnd.n7306 gnd.n446 19.3944
R14648 gnd.n7310 gnd.n446 19.3944
R14649 gnd.n7310 gnd.n442 19.3944
R14650 gnd.n7316 gnd.n442 19.3944
R14651 gnd.n7316 gnd.n440 19.3944
R14652 gnd.n7320 gnd.n440 19.3944
R14653 gnd.n7320 gnd.n436 19.3944
R14654 gnd.n7326 gnd.n436 19.3944
R14655 gnd.n7326 gnd.n434 19.3944
R14656 gnd.n7330 gnd.n434 19.3944
R14657 gnd.n7330 gnd.n430 19.3944
R14658 gnd.n7336 gnd.n430 19.3944
R14659 gnd.n7336 gnd.n428 19.3944
R14660 gnd.n7340 gnd.n428 19.3944
R14661 gnd.n7340 gnd.n424 19.3944
R14662 gnd.n7347 gnd.n424 19.3944
R14663 gnd.n7347 gnd.n422 19.3944
R14664 gnd.n7351 gnd.n422 19.3944
R14665 gnd.n6719 gnd.n795 19.3944
R14666 gnd.n6725 gnd.n795 19.3944
R14667 gnd.n6725 gnd.n793 19.3944
R14668 gnd.n6729 gnd.n793 19.3944
R14669 gnd.n6729 gnd.n789 19.3944
R14670 gnd.n6735 gnd.n789 19.3944
R14671 gnd.n6735 gnd.n787 19.3944
R14672 gnd.n6739 gnd.n787 19.3944
R14673 gnd.n6739 gnd.n783 19.3944
R14674 gnd.n6745 gnd.n783 19.3944
R14675 gnd.n6745 gnd.n781 19.3944
R14676 gnd.n6749 gnd.n781 19.3944
R14677 gnd.n6749 gnd.n777 19.3944
R14678 gnd.n6755 gnd.n777 19.3944
R14679 gnd.n6755 gnd.n775 19.3944
R14680 gnd.n6759 gnd.n775 19.3944
R14681 gnd.n6759 gnd.n771 19.3944
R14682 gnd.n6765 gnd.n771 19.3944
R14683 gnd.n6765 gnd.n769 19.3944
R14684 gnd.n6769 gnd.n769 19.3944
R14685 gnd.n6769 gnd.n765 19.3944
R14686 gnd.n6775 gnd.n765 19.3944
R14687 gnd.n6775 gnd.n763 19.3944
R14688 gnd.n6779 gnd.n763 19.3944
R14689 gnd.n6779 gnd.n759 19.3944
R14690 gnd.n6785 gnd.n759 19.3944
R14691 gnd.n6785 gnd.n757 19.3944
R14692 gnd.n6789 gnd.n757 19.3944
R14693 gnd.n6789 gnd.n753 19.3944
R14694 gnd.n6795 gnd.n753 19.3944
R14695 gnd.n6795 gnd.n751 19.3944
R14696 gnd.n6799 gnd.n751 19.3944
R14697 gnd.n6799 gnd.n747 19.3944
R14698 gnd.n6805 gnd.n747 19.3944
R14699 gnd.n6805 gnd.n745 19.3944
R14700 gnd.n6809 gnd.n745 19.3944
R14701 gnd.n6809 gnd.n741 19.3944
R14702 gnd.n6815 gnd.n741 19.3944
R14703 gnd.n6815 gnd.n739 19.3944
R14704 gnd.n6819 gnd.n739 19.3944
R14705 gnd.n6819 gnd.n735 19.3944
R14706 gnd.n6825 gnd.n735 19.3944
R14707 gnd.n6825 gnd.n733 19.3944
R14708 gnd.n6829 gnd.n733 19.3944
R14709 gnd.n6829 gnd.n729 19.3944
R14710 gnd.n6835 gnd.n729 19.3944
R14711 gnd.n6835 gnd.n727 19.3944
R14712 gnd.n6839 gnd.n727 19.3944
R14713 gnd.n6839 gnd.n723 19.3944
R14714 gnd.n6845 gnd.n723 19.3944
R14715 gnd.n6845 gnd.n721 19.3944
R14716 gnd.n6849 gnd.n721 19.3944
R14717 gnd.n6849 gnd.n717 19.3944
R14718 gnd.n6855 gnd.n717 19.3944
R14719 gnd.n6855 gnd.n715 19.3944
R14720 gnd.n6859 gnd.n715 19.3944
R14721 gnd.n6859 gnd.n711 19.3944
R14722 gnd.n6865 gnd.n711 19.3944
R14723 gnd.n6865 gnd.n709 19.3944
R14724 gnd.n6869 gnd.n709 19.3944
R14725 gnd.n6869 gnd.n705 19.3944
R14726 gnd.n6875 gnd.n705 19.3944
R14727 gnd.n6875 gnd.n703 19.3944
R14728 gnd.n6879 gnd.n703 19.3944
R14729 gnd.n6879 gnd.n699 19.3944
R14730 gnd.n6885 gnd.n699 19.3944
R14731 gnd.n6885 gnd.n697 19.3944
R14732 gnd.n6889 gnd.n697 19.3944
R14733 gnd.n6889 gnd.n693 19.3944
R14734 gnd.n6895 gnd.n693 19.3944
R14735 gnd.n6895 gnd.n691 19.3944
R14736 gnd.n6899 gnd.n691 19.3944
R14737 gnd.n6899 gnd.n687 19.3944
R14738 gnd.n6905 gnd.n687 19.3944
R14739 gnd.n6905 gnd.n685 19.3944
R14740 gnd.n6909 gnd.n685 19.3944
R14741 gnd.n6909 gnd.n681 19.3944
R14742 gnd.n6915 gnd.n681 19.3944
R14743 gnd.n6915 gnd.n679 19.3944
R14744 gnd.n6919 gnd.n679 19.3944
R14745 gnd.n6919 gnd.n675 19.3944
R14746 gnd.n6925 gnd.n675 19.3944
R14747 gnd.n6925 gnd.n673 19.3944
R14748 gnd.n6929 gnd.n673 19.3944
R14749 gnd.n6929 gnd.n669 19.3944
R14750 gnd.n6935 gnd.n669 19.3944
R14751 gnd.n6935 gnd.n667 19.3944
R14752 gnd.n6939 gnd.n667 19.3944
R14753 gnd.n6939 gnd.n663 19.3944
R14754 gnd.n6945 gnd.n663 19.3944
R14755 gnd.n6945 gnd.n661 19.3944
R14756 gnd.n6949 gnd.n661 19.3944
R14757 gnd.n6949 gnd.n657 19.3944
R14758 gnd.n6955 gnd.n657 19.3944
R14759 gnd.n6955 gnd.n655 19.3944
R14760 gnd.n6959 gnd.n655 19.3944
R14761 gnd.n6959 gnd.n651 19.3944
R14762 gnd.n6965 gnd.n651 19.3944
R14763 gnd.n6965 gnd.n649 19.3944
R14764 gnd.n6969 gnd.n649 19.3944
R14765 gnd.n6969 gnd.n645 19.3944
R14766 gnd.n6975 gnd.n645 19.3944
R14767 gnd.n6975 gnd.n643 19.3944
R14768 gnd.n6979 gnd.n643 19.3944
R14769 gnd.n6979 gnd.n639 19.3944
R14770 gnd.n6985 gnd.n639 19.3944
R14771 gnd.n6985 gnd.n637 19.3944
R14772 gnd.n6989 gnd.n637 19.3944
R14773 gnd.n6989 gnd.n633 19.3944
R14774 gnd.n6995 gnd.n633 19.3944
R14775 gnd.n6995 gnd.n631 19.3944
R14776 gnd.n6999 gnd.n631 19.3944
R14777 gnd.n6999 gnd.n627 19.3944
R14778 gnd.n7005 gnd.n627 19.3944
R14779 gnd.n7005 gnd.n625 19.3944
R14780 gnd.n7009 gnd.n625 19.3944
R14781 gnd.n7009 gnd.n621 19.3944
R14782 gnd.n7015 gnd.n621 19.3944
R14783 gnd.n7015 gnd.n619 19.3944
R14784 gnd.n7019 gnd.n619 19.3944
R14785 gnd.n7019 gnd.n615 19.3944
R14786 gnd.n7025 gnd.n615 19.3944
R14787 gnd.n7025 gnd.n613 19.3944
R14788 gnd.n7029 gnd.n613 19.3944
R14789 gnd.n7029 gnd.n609 19.3944
R14790 gnd.n7035 gnd.n609 19.3944
R14791 gnd.n7035 gnd.n607 19.3944
R14792 gnd.n7039 gnd.n607 19.3944
R14793 gnd.n7039 gnd.n603 19.3944
R14794 gnd.n7045 gnd.n603 19.3944
R14795 gnd.n7045 gnd.n601 19.3944
R14796 gnd.n7049 gnd.n601 19.3944
R14797 gnd.n7049 gnd.n597 19.3944
R14798 gnd.n7055 gnd.n597 19.3944
R14799 gnd.n7055 gnd.n595 19.3944
R14800 gnd.n7059 gnd.n595 19.3944
R14801 gnd.n7059 gnd.n591 19.3944
R14802 gnd.n7065 gnd.n591 19.3944
R14803 gnd.n7065 gnd.n589 19.3944
R14804 gnd.n7069 gnd.n589 19.3944
R14805 gnd.n7069 gnd.n585 19.3944
R14806 gnd.n7075 gnd.n585 19.3944
R14807 gnd.n7075 gnd.n583 19.3944
R14808 gnd.n7079 gnd.n583 19.3944
R14809 gnd.n7079 gnd.n579 19.3944
R14810 gnd.n7085 gnd.n579 19.3944
R14811 gnd.n7085 gnd.n577 19.3944
R14812 gnd.n7089 gnd.n577 19.3944
R14813 gnd.n7089 gnd.n573 19.3944
R14814 gnd.n7095 gnd.n573 19.3944
R14815 gnd.n7095 gnd.n571 19.3944
R14816 gnd.n7099 gnd.n571 19.3944
R14817 gnd.n7099 gnd.n567 19.3944
R14818 gnd.n7105 gnd.n567 19.3944
R14819 gnd.n7105 gnd.n565 19.3944
R14820 gnd.n7109 gnd.n565 19.3944
R14821 gnd.n7109 gnd.n561 19.3944
R14822 gnd.n7115 gnd.n561 19.3944
R14823 gnd.n7115 gnd.n559 19.3944
R14824 gnd.n7119 gnd.n559 19.3944
R14825 gnd.n7119 gnd.n555 19.3944
R14826 gnd.n7125 gnd.n555 19.3944
R14827 gnd.n7125 gnd.n553 19.3944
R14828 gnd.n7130 gnd.n553 19.3944
R14829 gnd.n7130 gnd.n549 19.3944
R14830 gnd.n7136 gnd.n549 19.3944
R14831 gnd.n7137 gnd.n7136 19.3944
R14832 gnd.n6291 gnd.n6290 19.3944
R14833 gnd.n6290 gnd.n6289 19.3944
R14834 gnd.n6289 gnd.n6288 19.3944
R14835 gnd.n6288 gnd.n6286 19.3944
R14836 gnd.n6286 gnd.n6283 19.3944
R14837 gnd.n6283 gnd.n6282 19.3944
R14838 gnd.n6282 gnd.n6279 19.3944
R14839 gnd.n6279 gnd.n6278 19.3944
R14840 gnd.n6278 gnd.n6275 19.3944
R14841 gnd.n6275 gnd.n6274 19.3944
R14842 gnd.n6274 gnd.n6271 19.3944
R14843 gnd.n6271 gnd.n6270 19.3944
R14844 gnd.n6270 gnd.n6267 19.3944
R14845 gnd.n6267 gnd.n6266 19.3944
R14846 gnd.n6266 gnd.n6263 19.3944
R14847 gnd.n6261 gnd.n6258 19.3944
R14848 gnd.n6258 gnd.n6257 19.3944
R14849 gnd.n6257 gnd.n6254 19.3944
R14850 gnd.n6254 gnd.n6253 19.3944
R14851 gnd.n6253 gnd.n6250 19.3944
R14852 gnd.n6250 gnd.n6249 19.3944
R14853 gnd.n6249 gnd.n6246 19.3944
R14854 gnd.n6246 gnd.n6245 19.3944
R14855 gnd.n6245 gnd.n6242 19.3944
R14856 gnd.n6242 gnd.n6241 19.3944
R14857 gnd.n6241 gnd.n6238 19.3944
R14858 gnd.n6238 gnd.n6237 19.3944
R14859 gnd.n6237 gnd.n6234 19.3944
R14860 gnd.n6234 gnd.n6233 19.3944
R14861 gnd.n6233 gnd.n6230 19.3944
R14862 gnd.n6230 gnd.n6229 19.3944
R14863 gnd.n6229 gnd.n6226 19.3944
R14864 gnd.n6226 gnd.n6225 19.3944
R14865 gnd.n1455 gnd.n1335 19.3944
R14866 gnd.n1455 gnd.n1454 19.3944
R14867 gnd.n1473 gnd.n1454 19.3944
R14868 gnd.n1473 gnd.n1472 19.3944
R14869 gnd.n1472 gnd.n1471 19.3944
R14870 gnd.n1471 gnd.n1469 19.3944
R14871 gnd.n1469 gnd.n1468 19.3944
R14872 gnd.n1468 gnd.n1466 19.3944
R14873 gnd.n1466 gnd.n1465 19.3944
R14874 gnd.n1465 gnd.n1391 19.3944
R14875 gnd.n6123 gnd.n1391 19.3944
R14876 gnd.n6123 gnd.n1389 19.3944
R14877 gnd.n6127 gnd.n1389 19.3944
R14878 gnd.n6128 gnd.n6127 19.3944
R14879 gnd.n6130 gnd.n6128 19.3944
R14880 gnd.n6130 gnd.n1387 19.3944
R14881 gnd.n6136 gnd.n1387 19.3944
R14882 gnd.n6136 gnd.n6135 19.3944
R14883 gnd.n6135 gnd.n388 19.3944
R14884 gnd.n7386 gnd.n388 19.3944
R14885 gnd.n7386 gnd.n386 19.3944
R14886 gnd.n7396 gnd.n386 19.3944
R14887 gnd.n7396 gnd.n7395 19.3944
R14888 gnd.n7395 gnd.n7394 19.3944
R14889 gnd.n7394 gnd.n354 19.3944
R14890 gnd.n7431 gnd.n354 19.3944
R14891 gnd.n7431 gnd.n352 19.3944
R14892 gnd.n7442 gnd.n352 19.3944
R14893 gnd.n7442 gnd.n7441 19.3944
R14894 gnd.n7441 gnd.n7440 19.3944
R14895 gnd.n7440 gnd.n7438 19.3944
R14896 gnd.n7438 gnd.n338 19.3944
R14897 gnd.n7461 gnd.n338 19.3944
R14898 gnd.n7461 gnd.n336 19.3944
R14899 gnd.n7530 gnd.n336 19.3944
R14900 gnd.n7530 gnd.n7529 19.3944
R14901 gnd.n7529 gnd.n7528 19.3944
R14902 gnd.n7528 gnd.n7526 19.3944
R14903 gnd.n7526 gnd.n7525 19.3944
R14904 gnd.n7525 gnd.n7523 19.3944
R14905 gnd.n7523 gnd.n7522 19.3944
R14906 gnd.n7522 gnd.n7520 19.3944
R14907 gnd.n7520 gnd.n7519 19.3944
R14908 gnd.n7519 gnd.n7517 19.3944
R14909 gnd.n7517 gnd.n7516 19.3944
R14910 gnd.n7516 gnd.n7514 19.3944
R14911 gnd.n7514 gnd.n7513 19.3944
R14912 gnd.n7513 gnd.n7511 19.3944
R14913 gnd.n7511 gnd.n7510 19.3944
R14914 gnd.n7510 gnd.n7508 19.3944
R14915 gnd.n7508 gnd.n7507 19.3944
R14916 gnd.n7507 gnd.n7505 19.3944
R14917 gnd.n7505 gnd.n7504 19.3944
R14918 gnd.n7504 gnd.n7502 19.3944
R14919 gnd.n7502 gnd.n7501 19.3944
R14920 gnd.n7501 gnd.n7499 19.3944
R14921 gnd.n7499 gnd.n7498 19.3944
R14922 gnd.n7498 gnd.n7496 19.3944
R14923 gnd.n7496 gnd.n7495 19.3944
R14924 gnd.n7495 gnd.n7493 19.3944
R14925 gnd.n7493 gnd.n7492 19.3944
R14926 gnd.n7492 gnd.n204 19.3944
R14927 gnd.n7727 gnd.n204 19.3944
R14928 gnd.n7728 gnd.n7727 19.3944
R14929 gnd.n7766 gnd.n165 19.3944
R14930 gnd.n7761 gnd.n165 19.3944
R14931 gnd.n7761 gnd.n7760 19.3944
R14932 gnd.n7760 gnd.n7759 19.3944
R14933 gnd.n7759 gnd.n172 19.3944
R14934 gnd.n7754 gnd.n172 19.3944
R14935 gnd.n7754 gnd.n7753 19.3944
R14936 gnd.n7753 gnd.n7752 19.3944
R14937 gnd.n7752 gnd.n179 19.3944
R14938 gnd.n7747 gnd.n179 19.3944
R14939 gnd.n7747 gnd.n7746 19.3944
R14940 gnd.n7746 gnd.n7745 19.3944
R14941 gnd.n7745 gnd.n186 19.3944
R14942 gnd.n7740 gnd.n186 19.3944
R14943 gnd.n7740 gnd.n7739 19.3944
R14944 gnd.n7739 gnd.n7738 19.3944
R14945 gnd.n7738 gnd.n193 19.3944
R14946 gnd.n7733 gnd.n193 19.3944
R14947 gnd.n7799 gnd.n7798 19.3944
R14948 gnd.n7798 gnd.n7797 19.3944
R14949 gnd.n7797 gnd.n137 19.3944
R14950 gnd.n7792 gnd.n137 19.3944
R14951 gnd.n7792 gnd.n7791 19.3944
R14952 gnd.n7791 gnd.n7790 19.3944
R14953 gnd.n7790 gnd.n144 19.3944
R14954 gnd.n7785 gnd.n144 19.3944
R14955 gnd.n7785 gnd.n7784 19.3944
R14956 gnd.n7784 gnd.n7783 19.3944
R14957 gnd.n7783 gnd.n151 19.3944
R14958 gnd.n7778 gnd.n151 19.3944
R14959 gnd.n7778 gnd.n7777 19.3944
R14960 gnd.n7777 gnd.n7776 19.3944
R14961 gnd.n7776 gnd.n158 19.3944
R14962 gnd.n7771 gnd.n158 19.3944
R14963 gnd.n7771 gnd.n7770 19.3944
R14964 gnd.n6051 gnd.n6046 19.3944
R14965 gnd.n6051 gnd.n6050 19.3944
R14966 gnd.n6050 gnd.n1429 19.3944
R14967 gnd.n6076 gnd.n1429 19.3944
R14968 gnd.n6076 gnd.n1427 19.3944
R14969 gnd.n6082 gnd.n1427 19.3944
R14970 gnd.n6082 gnd.n6081 19.3944
R14971 gnd.n6081 gnd.n1402 19.3944
R14972 gnd.n6113 gnd.n1402 19.3944
R14973 gnd.n6113 gnd.n1400 19.3944
R14974 gnd.n6119 gnd.n1400 19.3944
R14975 gnd.n6119 gnd.n6118 19.3944
R14976 gnd.n6118 gnd.n1368 19.3944
R14977 gnd.n6183 gnd.n1368 19.3944
R14978 gnd.n6183 gnd.n1366 19.3944
R14979 gnd.n6187 gnd.n1366 19.3944
R14980 gnd.n6187 gnd.n397 19.3944
R14981 gnd.n7376 gnd.n397 19.3944
R14982 gnd.n7376 gnd.n395 19.3944
R14983 gnd.n7382 gnd.n395 19.3944
R14984 gnd.n7382 gnd.n7381 19.3944
R14985 gnd.n7381 gnd.n364 19.3944
R14986 gnd.n7422 gnd.n364 19.3944
R14987 gnd.n7422 gnd.n362 19.3944
R14988 gnd.n7426 gnd.n362 19.3944
R14989 gnd.n7427 gnd.n7426 19.3944
R14990 gnd.n7427 gnd.n309 19.3944
R14991 gnd.n7554 gnd.n7553 19.3944
R14992 gnd.n342 gnd.n341 19.3944
R14993 gnd.n7457 gnd.n7456 19.3944
R14994 gnd.n332 gnd.n331 19.3944
R14995 gnd.n7534 gnd.n302 19.3944
R14996 gnd.n7558 gnd.n302 19.3944
R14997 gnd.n7558 gnd.n288 19.3944
R14998 gnd.n7570 gnd.n288 19.3944
R14999 gnd.n7570 gnd.n286 19.3944
R15000 gnd.n7574 gnd.n286 19.3944
R15001 gnd.n7574 gnd.n274 19.3944
R15002 gnd.n7586 gnd.n274 19.3944
R15003 gnd.n7586 gnd.n272 19.3944
R15004 gnd.n7590 gnd.n272 19.3944
R15005 gnd.n7590 gnd.n258 19.3944
R15006 gnd.n7602 gnd.n258 19.3944
R15007 gnd.n7602 gnd.n256 19.3944
R15008 gnd.n7606 gnd.n256 19.3944
R15009 gnd.n7606 gnd.n243 19.3944
R15010 gnd.n7618 gnd.n243 19.3944
R15011 gnd.n7618 gnd.n241 19.3944
R15012 gnd.n7622 gnd.n241 19.3944
R15013 gnd.n7622 gnd.n227 19.3944
R15014 gnd.n7634 gnd.n227 19.3944
R15015 gnd.n7634 gnd.n225 19.3944
R15016 gnd.n7638 gnd.n225 19.3944
R15017 gnd.n7638 gnd.n211 19.3944
R15018 gnd.n7718 gnd.n211 19.3944
R15019 gnd.n7718 gnd.n209 19.3944
R15020 gnd.n7722 gnd.n209 19.3944
R15021 gnd.n7722 gnd.n132 19.3944
R15022 gnd.n7802 gnd.n132 19.3944
R15023 gnd.n4189 gnd.n4188 19.3944
R15024 gnd.n4188 gnd.n3975 19.3944
R15025 gnd.n4183 gnd.n3975 19.3944
R15026 gnd.n4183 gnd.n4182 19.3944
R15027 gnd.n4182 gnd.n3980 19.3944
R15028 gnd.n4177 gnd.n3980 19.3944
R15029 gnd.n4177 gnd.n4176 19.3944
R15030 gnd.n4176 gnd.n4175 19.3944
R15031 gnd.n4175 gnd.n3986 19.3944
R15032 gnd.n4169 gnd.n3986 19.3944
R15033 gnd.n4169 gnd.n4168 19.3944
R15034 gnd.n4168 gnd.n4167 19.3944
R15035 gnd.n4167 gnd.n3992 19.3944
R15036 gnd.n4161 gnd.n3992 19.3944
R15037 gnd.n4161 gnd.n4160 19.3944
R15038 gnd.n4160 gnd.n4159 19.3944
R15039 gnd.n4159 gnd.n3998 19.3944
R15040 gnd.n4153 gnd.n4152 19.3944
R15041 gnd.n4152 gnd.n4151 19.3944
R15042 gnd.n4151 gnd.n4007 19.3944
R15043 gnd.n4145 gnd.n4007 19.3944
R15044 gnd.n4145 gnd.n4144 19.3944
R15045 gnd.n4144 gnd.n4143 19.3944
R15046 gnd.n4143 gnd.n4013 19.3944
R15047 gnd.n4137 gnd.n4013 19.3944
R15048 gnd.n4137 gnd.n4136 19.3944
R15049 gnd.n4136 gnd.n4135 19.3944
R15050 gnd.n4135 gnd.n4019 19.3944
R15051 gnd.n4129 gnd.n4019 19.3944
R15052 gnd.n4129 gnd.n4128 19.3944
R15053 gnd.n4128 gnd.n4127 19.3944
R15054 gnd.n4127 gnd.n4025 19.3944
R15055 gnd.n4121 gnd.n4025 19.3944
R15056 gnd.n4121 gnd.n4120 19.3944
R15057 gnd.n4120 gnd.n4119 19.3944
R15058 gnd.n4196 gnd.n2331 19.3944
R15059 gnd.n4200 gnd.n2331 19.3944
R15060 gnd.n4200 gnd.n2318 19.3944
R15061 gnd.n4212 gnd.n2318 19.3944
R15062 gnd.n4212 gnd.n2316 19.3944
R15063 gnd.n4216 gnd.n2316 19.3944
R15064 gnd.n4216 gnd.n2301 19.3944
R15065 gnd.n4228 gnd.n2301 19.3944
R15066 gnd.n4228 gnd.n2299 19.3944
R15067 gnd.n4232 gnd.n2299 19.3944
R15068 gnd.n4232 gnd.n2286 19.3944
R15069 gnd.n4244 gnd.n2286 19.3944
R15070 gnd.n4244 gnd.n2284 19.3944
R15071 gnd.n4248 gnd.n2284 19.3944
R15072 gnd.n4248 gnd.n2269 19.3944
R15073 gnd.n4260 gnd.n2269 19.3944
R15074 gnd.n4260 gnd.n2267 19.3944
R15075 gnd.n4264 gnd.n2267 19.3944
R15076 gnd.n4264 gnd.n2254 19.3944
R15077 gnd.n4276 gnd.n2254 19.3944
R15078 gnd.n4276 gnd.n2252 19.3944
R15079 gnd.n4280 gnd.n2252 19.3944
R15080 gnd.n4280 gnd.n2237 19.3944
R15081 gnd.n4293 gnd.n2237 19.3944
R15082 gnd.n4293 gnd.n2235 19.3944
R15083 gnd.n4297 gnd.n2235 19.3944
R15084 gnd.n4297 gnd.n2223 19.3944
R15085 gnd.n4309 gnd.n2223 19.3944
R15086 gnd.n4309 gnd.n2221 19.3944
R15087 gnd.n4314 gnd.n2221 19.3944
R15088 gnd.n4314 gnd.n4313 19.3944
R15089 gnd.n4313 gnd.n2198 19.3944
R15090 gnd.n2198 gnd.n2196 19.3944
R15091 gnd.n4341 gnd.n2196 19.3944
R15092 gnd.n4341 gnd.n4340 19.3944
R15093 gnd.n4340 gnd.n4339 19.3944
R15094 gnd.n4339 gnd.n4338 19.3944
R15095 gnd.n4338 gnd.n4336 19.3944
R15096 gnd.n4336 gnd.n989 19.3944
R15097 gnd.n6533 gnd.n989 19.3944
R15098 gnd.n6533 gnd.n6532 19.3944
R15099 gnd.n6532 gnd.n6531 19.3944
R15100 gnd.n6531 gnd.n993 19.3944
R15101 gnd.n6521 gnd.n993 19.3944
R15102 gnd.n6521 gnd.n6520 19.3944
R15103 gnd.n6520 gnd.n6519 19.3944
R15104 gnd.n6519 gnd.n1013 19.3944
R15105 gnd.n6509 gnd.n1013 19.3944
R15106 gnd.n6509 gnd.n6508 19.3944
R15107 gnd.n6508 gnd.n6507 19.3944
R15108 gnd.n6507 gnd.n1035 19.3944
R15109 gnd.n6497 gnd.n1035 19.3944
R15110 gnd.n6497 gnd.n6496 19.3944
R15111 gnd.n6496 gnd.n6495 19.3944
R15112 gnd.n6495 gnd.n1055 19.3944
R15113 gnd.n6485 gnd.n1055 19.3944
R15114 gnd.n6485 gnd.n6484 19.3944
R15115 gnd.n6484 gnd.n6483 19.3944
R15116 gnd.n6483 gnd.n1077 19.3944
R15117 gnd.n6473 gnd.n1077 19.3944
R15118 gnd.n6473 gnd.n6472 19.3944
R15119 gnd.n6472 gnd.n6471 19.3944
R15120 gnd.n6471 gnd.n1098 19.3944
R15121 gnd.n6461 gnd.n1098 19.3944
R15122 gnd.n3832 gnd.n3831 19.3944
R15123 gnd.n3837 gnd.n3832 19.3944
R15124 gnd.n3837 gnd.n3829 19.3944
R15125 gnd.n3841 gnd.n3829 19.3944
R15126 gnd.n3841 gnd.n3827 19.3944
R15127 gnd.n3847 gnd.n3827 19.3944
R15128 gnd.n3847 gnd.n3825 19.3944
R15129 gnd.n3851 gnd.n3825 19.3944
R15130 gnd.n3851 gnd.n3823 19.3944
R15131 gnd.n3857 gnd.n3823 19.3944
R15132 gnd.n3857 gnd.n3821 19.3944
R15133 gnd.n3861 gnd.n3821 19.3944
R15134 gnd.n3861 gnd.n3819 19.3944
R15135 gnd.n3867 gnd.n3819 19.3944
R15136 gnd.n3867 gnd.n3817 19.3944
R15137 gnd.n3871 gnd.n3817 19.3944
R15138 gnd.n3970 gnd.n3811 19.3944
R15139 gnd.n3970 gnd.n3969 19.3944
R15140 gnd.n3969 gnd.n3968 19.3944
R15141 gnd.n3968 gnd.n3966 19.3944
R15142 gnd.n3966 gnd.n3965 19.3944
R15143 gnd.n3965 gnd.n3963 19.3944
R15144 gnd.n3963 gnd.n3962 19.3944
R15145 gnd.n3962 gnd.n3960 19.3944
R15146 gnd.n3960 gnd.n3959 19.3944
R15147 gnd.n3959 gnd.n3957 19.3944
R15148 gnd.n3957 gnd.n3956 19.3944
R15149 gnd.n3956 gnd.n3954 19.3944
R15150 gnd.n3954 gnd.n3953 19.3944
R15151 gnd.n3953 gnd.n3951 19.3944
R15152 gnd.n3951 gnd.n3950 19.3944
R15153 gnd.n3950 gnd.n3948 19.3944
R15154 gnd.n3948 gnd.n3947 19.3944
R15155 gnd.n3947 gnd.n3945 19.3944
R15156 gnd.n3945 gnd.n3944 19.3944
R15157 gnd.n3944 gnd.n3942 19.3944
R15158 gnd.n3942 gnd.n3941 19.3944
R15159 gnd.n3941 gnd.n3939 19.3944
R15160 gnd.n3939 gnd.n3938 19.3944
R15161 gnd.n3938 gnd.n3936 19.3944
R15162 gnd.n3936 gnd.n3935 19.3944
R15163 gnd.n3935 gnd.n3933 19.3944
R15164 gnd.n3933 gnd.n3932 19.3944
R15165 gnd.n3932 gnd.n3930 19.3944
R15166 gnd.n3930 gnd.n3929 19.3944
R15167 gnd.n3929 gnd.n3927 19.3944
R15168 gnd.n3927 gnd.n3926 19.3944
R15169 gnd.n3926 gnd.n3924 19.3944
R15170 gnd.n3924 gnd.n3911 19.3944
R15171 gnd.n3920 gnd.n3911 19.3944
R15172 gnd.n3920 gnd.n3919 19.3944
R15173 gnd.n3919 gnd.n3918 19.3944
R15174 gnd.n3918 gnd.n3915 19.3944
R15175 gnd.n3915 gnd.n2180 19.3944
R15176 gnd.n4361 gnd.n2180 19.3944
R15177 gnd.n4361 gnd.n2178 19.3944
R15178 gnd.n4365 gnd.n2178 19.3944
R15179 gnd.n4365 gnd.n2168 19.3944
R15180 gnd.n4406 gnd.n2168 19.3944
R15181 gnd.n4406 gnd.n2169 19.3944
R15182 gnd.n4402 gnd.n2169 19.3944
R15183 gnd.n4402 gnd.n4401 19.3944
R15184 gnd.n4401 gnd.n4400 19.3944
R15185 gnd.n4400 gnd.n4395 19.3944
R15186 gnd.n4396 gnd.n4395 19.3944
R15187 gnd.n4396 gnd.n2147 19.3944
R15188 gnd.n4455 gnd.n2147 19.3944
R15189 gnd.n4455 gnd.n2148 19.3944
R15190 gnd.n4451 gnd.n2148 19.3944
R15191 gnd.n4451 gnd.n4450 19.3944
R15192 gnd.n4450 gnd.n4449 19.3944
R15193 gnd.n4449 gnd.n2134 19.3944
R15194 gnd.n4513 gnd.n2134 19.3944
R15195 gnd.n4513 gnd.n2132 19.3944
R15196 gnd.n4517 gnd.n2132 19.3944
R15197 gnd.n4517 gnd.n2128 19.3944
R15198 gnd.n4530 gnd.n2128 19.3944
R15199 gnd.n4530 gnd.n2125 19.3944
R15200 gnd.n4566 gnd.n2125 19.3944
R15201 gnd.n4566 gnd.n2126 19.3944
R15202 gnd.n4110 gnd.n4109 19.3944
R15203 gnd.n4109 gnd.n4108 19.3944
R15204 gnd.n4108 gnd.n4107 19.3944
R15205 gnd.n4107 gnd.n4105 19.3944
R15206 gnd.n4105 gnd.n4104 19.3944
R15207 gnd.n4104 gnd.n4102 19.3944
R15208 gnd.n4102 gnd.n4101 19.3944
R15209 gnd.n4101 gnd.n4099 19.3944
R15210 gnd.n4099 gnd.n4098 19.3944
R15211 gnd.n4098 gnd.n4096 19.3944
R15212 gnd.n4096 gnd.n4095 19.3944
R15213 gnd.n4095 gnd.n4093 19.3944
R15214 gnd.n4093 gnd.n4092 19.3944
R15215 gnd.n4092 gnd.n4090 19.3944
R15216 gnd.n4090 gnd.n4089 19.3944
R15217 gnd.n4089 gnd.n4087 19.3944
R15218 gnd.n4087 gnd.n4086 19.3944
R15219 gnd.n4086 gnd.n4084 19.3944
R15220 gnd.n4084 gnd.n4083 19.3944
R15221 gnd.n4083 gnd.n4081 19.3944
R15222 gnd.n4081 gnd.n4080 19.3944
R15223 gnd.n4080 gnd.n4078 19.3944
R15224 gnd.n4078 gnd.n4077 19.3944
R15225 gnd.n4077 gnd.n4075 19.3944
R15226 gnd.n4075 gnd.n4074 19.3944
R15227 gnd.n4074 gnd.n4072 19.3944
R15228 gnd.n4072 gnd.n4071 19.3944
R15229 gnd.n4071 gnd.n4069 19.3944
R15230 gnd.n4069 gnd.n4068 19.3944
R15231 gnd.n4068 gnd.n4066 19.3944
R15232 gnd.n4066 gnd.n2201 19.3944
R15233 gnd.n4326 gnd.n2201 19.3944
R15234 gnd.n4326 gnd.n2206 19.3944
R15235 gnd.n2206 gnd.n2205 19.3944
R15236 gnd.n2205 gnd.n2204 19.3944
R15237 gnd.n2204 gnd.n2183 19.3944
R15238 gnd.n4353 gnd.n2183 19.3944
R15239 gnd.n4353 gnd.n2181 19.3944
R15240 gnd.n4357 gnd.n2181 19.3944
R15241 gnd.n4357 gnd.n2177 19.3944
R15242 gnd.n4379 gnd.n2177 19.3944
R15243 gnd.n4379 gnd.n2175 19.3944
R15244 gnd.n4383 gnd.n2175 19.3944
R15245 gnd.n4384 gnd.n4383 19.3944
R15246 gnd.n4387 gnd.n4384 19.3944
R15247 gnd.n4387 gnd.n2173 19.3944
R15248 gnd.n4391 gnd.n2173 19.3944
R15249 gnd.n4391 gnd.n2156 19.3944
R15250 gnd.n4428 gnd.n2156 19.3944
R15251 gnd.n4428 gnd.n2154 19.3944
R15252 gnd.n4432 gnd.n2154 19.3944
R15253 gnd.n4433 gnd.n4432 19.3944
R15254 gnd.n4436 gnd.n4433 19.3944
R15255 gnd.n4436 gnd.n2152 19.3944
R15256 gnd.n4444 gnd.n2152 19.3944
R15257 gnd.n4444 gnd.n4443 19.3944
R15258 gnd.n4443 gnd.n4442 19.3944
R15259 gnd.n4442 gnd.n2131 19.3944
R15260 gnd.n4521 gnd.n2131 19.3944
R15261 gnd.n4521 gnd.n2129 19.3944
R15262 gnd.n4526 gnd.n2129 19.3944
R15263 gnd.n4526 gnd.n2123 19.3944
R15264 gnd.n4570 gnd.n2123 19.3944
R15265 gnd.n4571 gnd.n4570 19.3944
R15266 gnd.n4613 gnd.n2097 19.3944
R15267 gnd.n4613 gnd.n4610 19.3944
R15268 gnd.n4610 gnd.n4607 19.3944
R15269 gnd.n4607 gnd.n4606 19.3944
R15270 gnd.n4606 gnd.n4603 19.3944
R15271 gnd.n4603 gnd.n4602 19.3944
R15272 gnd.n4602 gnd.n4599 19.3944
R15273 gnd.n4599 gnd.n4598 19.3944
R15274 gnd.n4598 gnd.n4595 19.3944
R15275 gnd.n4595 gnd.n4594 19.3944
R15276 gnd.n4594 gnd.n4591 19.3944
R15277 gnd.n4591 gnd.n4590 19.3944
R15278 gnd.n4590 gnd.n4587 19.3944
R15279 gnd.n4587 gnd.n4586 19.3944
R15280 gnd.n4586 gnd.n4583 19.3944
R15281 gnd.n4583 gnd.n4582 19.3944
R15282 gnd.n4582 gnd.n4579 19.3944
R15283 gnd.n4579 gnd.n4578 19.3944
R15284 gnd.n2080 gnd.n2079 19.3944
R15285 gnd.n5553 gnd.n2079 19.3944
R15286 gnd.n5553 gnd.n5552 19.3944
R15287 gnd.n5552 gnd.n5551 19.3944
R15288 gnd.n5551 gnd.n5548 19.3944
R15289 gnd.n5548 gnd.n5547 19.3944
R15290 gnd.n5547 gnd.n5544 19.3944
R15291 gnd.n5544 gnd.n5543 19.3944
R15292 gnd.n5543 gnd.n5540 19.3944
R15293 gnd.n5540 gnd.n5539 19.3944
R15294 gnd.n5539 gnd.n5536 19.3944
R15295 gnd.n5536 gnd.n5535 19.3944
R15296 gnd.n5535 gnd.n5532 19.3944
R15297 gnd.n5532 gnd.n5531 19.3944
R15298 gnd.n5531 gnd.n5528 19.3944
R15299 gnd.n4192 gnd.n2326 19.3944
R15300 gnd.n4204 gnd.n2326 19.3944
R15301 gnd.n4204 gnd.n2324 19.3944
R15302 gnd.n4208 gnd.n2324 19.3944
R15303 gnd.n4208 gnd.n2310 19.3944
R15304 gnd.n4220 gnd.n2310 19.3944
R15305 gnd.n4220 gnd.n2308 19.3944
R15306 gnd.n4224 gnd.n2308 19.3944
R15307 gnd.n4224 gnd.n2294 19.3944
R15308 gnd.n4236 gnd.n2294 19.3944
R15309 gnd.n4236 gnd.n2292 19.3944
R15310 gnd.n4240 gnd.n2292 19.3944
R15311 gnd.n4240 gnd.n2278 19.3944
R15312 gnd.n4252 gnd.n2278 19.3944
R15313 gnd.n4252 gnd.n2276 19.3944
R15314 gnd.n4256 gnd.n2276 19.3944
R15315 gnd.n4256 gnd.n2262 19.3944
R15316 gnd.n4268 gnd.n2262 19.3944
R15317 gnd.n4268 gnd.n2260 19.3944
R15318 gnd.n4272 gnd.n2260 19.3944
R15319 gnd.n4272 gnd.n2246 19.3944
R15320 gnd.n4284 gnd.n2246 19.3944
R15321 gnd.n4284 gnd.n2244 19.3944
R15322 gnd.n4289 gnd.n2244 19.3944
R15323 gnd.n4289 gnd.n2229 19.3944
R15324 gnd.n4301 gnd.n2229 19.3944
R15325 gnd.n4302 gnd.n4301 19.3944
R15326 gnd.n4305 gnd.n4304 19.3944
R15327 gnd.n4319 gnd.n4318 19.3944
R15328 gnd.n4322 gnd.n4321 19.3944
R15329 gnd.n4346 gnd.n4345 19.3944
R15330 gnd.n4348 gnd.n977 19.3944
R15331 gnd.n6539 gnd.n977 19.3944
R15332 gnd.n6539 gnd.n6538 19.3944
R15333 gnd.n6538 gnd.n6537 19.3944
R15334 gnd.n6537 gnd.n981 19.3944
R15335 gnd.n6527 gnd.n981 19.3944
R15336 gnd.n6527 gnd.n6526 19.3944
R15337 gnd.n6526 gnd.n6525 19.3944
R15338 gnd.n6525 gnd.n1003 19.3944
R15339 gnd.n6515 gnd.n1003 19.3944
R15340 gnd.n6515 gnd.n6514 19.3944
R15341 gnd.n6514 gnd.n6513 19.3944
R15342 gnd.n6513 gnd.n1024 19.3944
R15343 gnd.n6503 gnd.n1024 19.3944
R15344 gnd.n6503 gnd.n6502 19.3944
R15345 gnd.n6502 gnd.n6501 19.3944
R15346 gnd.n6501 gnd.n1045 19.3944
R15347 gnd.n6491 gnd.n1045 19.3944
R15348 gnd.n6491 gnd.n6490 19.3944
R15349 gnd.n6490 gnd.n6489 19.3944
R15350 gnd.n6489 gnd.n1066 19.3944
R15351 gnd.n6479 gnd.n1066 19.3944
R15352 gnd.n6479 gnd.n6478 19.3944
R15353 gnd.n6478 gnd.n6477 19.3944
R15354 gnd.n6477 gnd.n1087 19.3944
R15355 gnd.n6467 gnd.n1087 19.3944
R15356 gnd.n6467 gnd.n6466 19.3944
R15357 gnd.n6466 gnd.n6465 19.3944
R15358 gnd.n6716 gnd.n6715 19.3944
R15359 gnd.n6715 gnd.n800 19.3944
R15360 gnd.n6709 gnd.n800 19.3944
R15361 gnd.n6709 gnd.n6708 19.3944
R15362 gnd.n6708 gnd.n6707 19.3944
R15363 gnd.n6707 gnd.n808 19.3944
R15364 gnd.n6701 gnd.n808 19.3944
R15365 gnd.n6701 gnd.n6700 19.3944
R15366 gnd.n6700 gnd.n6699 19.3944
R15367 gnd.n6699 gnd.n816 19.3944
R15368 gnd.n6693 gnd.n816 19.3944
R15369 gnd.n6693 gnd.n6692 19.3944
R15370 gnd.n6692 gnd.n6691 19.3944
R15371 gnd.n6691 gnd.n824 19.3944
R15372 gnd.n6685 gnd.n824 19.3944
R15373 gnd.n6685 gnd.n6684 19.3944
R15374 gnd.n6684 gnd.n6683 19.3944
R15375 gnd.n6683 gnd.n832 19.3944
R15376 gnd.n6677 gnd.n832 19.3944
R15377 gnd.n6677 gnd.n6676 19.3944
R15378 gnd.n6676 gnd.n6675 19.3944
R15379 gnd.n6675 gnd.n840 19.3944
R15380 gnd.n6669 gnd.n840 19.3944
R15381 gnd.n6669 gnd.n6668 19.3944
R15382 gnd.n6668 gnd.n6667 19.3944
R15383 gnd.n6667 gnd.n848 19.3944
R15384 gnd.n6661 gnd.n848 19.3944
R15385 gnd.n6661 gnd.n6660 19.3944
R15386 gnd.n6660 gnd.n6659 19.3944
R15387 gnd.n6659 gnd.n856 19.3944
R15388 gnd.n6653 gnd.n856 19.3944
R15389 gnd.n6653 gnd.n6652 19.3944
R15390 gnd.n6652 gnd.n6651 19.3944
R15391 gnd.n6651 gnd.n864 19.3944
R15392 gnd.n6645 gnd.n864 19.3944
R15393 gnd.n6645 gnd.n6644 19.3944
R15394 gnd.n6644 gnd.n6643 19.3944
R15395 gnd.n6643 gnd.n872 19.3944
R15396 gnd.n6637 gnd.n872 19.3944
R15397 gnd.n6637 gnd.n6636 19.3944
R15398 gnd.n6636 gnd.n6635 19.3944
R15399 gnd.n6635 gnd.n880 19.3944
R15400 gnd.n6629 gnd.n880 19.3944
R15401 gnd.n6629 gnd.n6628 19.3944
R15402 gnd.n6628 gnd.n6627 19.3944
R15403 gnd.n6627 gnd.n888 19.3944
R15404 gnd.n6621 gnd.n888 19.3944
R15405 gnd.n6621 gnd.n6620 19.3944
R15406 gnd.n6620 gnd.n6619 19.3944
R15407 gnd.n6619 gnd.n896 19.3944
R15408 gnd.n6613 gnd.n896 19.3944
R15409 gnd.n6613 gnd.n6612 19.3944
R15410 gnd.n6612 gnd.n6611 19.3944
R15411 gnd.n6611 gnd.n904 19.3944
R15412 gnd.n6605 gnd.n904 19.3944
R15413 gnd.n6605 gnd.n6604 19.3944
R15414 gnd.n6604 gnd.n6603 19.3944
R15415 gnd.n6603 gnd.n912 19.3944
R15416 gnd.n6597 gnd.n912 19.3944
R15417 gnd.n6597 gnd.n6596 19.3944
R15418 gnd.n6596 gnd.n6595 19.3944
R15419 gnd.n6595 gnd.n920 19.3944
R15420 gnd.n6589 gnd.n920 19.3944
R15421 gnd.n6589 gnd.n6588 19.3944
R15422 gnd.n6588 gnd.n6587 19.3944
R15423 gnd.n6587 gnd.n928 19.3944
R15424 gnd.n6581 gnd.n928 19.3944
R15425 gnd.n6581 gnd.n6580 19.3944
R15426 gnd.n6580 gnd.n6579 19.3944
R15427 gnd.n6579 gnd.n936 19.3944
R15428 gnd.n6573 gnd.n936 19.3944
R15429 gnd.n6573 gnd.n6572 19.3944
R15430 gnd.n6572 gnd.n6571 19.3944
R15431 gnd.n6571 gnd.n944 19.3944
R15432 gnd.n6565 gnd.n944 19.3944
R15433 gnd.n6565 gnd.n6564 19.3944
R15434 gnd.n6564 gnd.n6563 19.3944
R15435 gnd.n6563 gnd.n952 19.3944
R15436 gnd.n6557 gnd.n952 19.3944
R15437 gnd.n6557 gnd.n6556 19.3944
R15438 gnd.n6556 gnd.n6555 19.3944
R15439 gnd.n6555 gnd.n960 19.3944
R15440 gnd.n6549 gnd.n960 19.3944
R15441 gnd.n6549 gnd.n6548 19.3944
R15442 gnd.n6456 gnd.n6455 19.3944
R15443 gnd.n6455 gnd.n6454 19.3944
R15444 gnd.n6454 gnd.n1121 19.3944
R15445 gnd.n6450 gnd.n1121 19.3944
R15446 gnd.n6450 gnd.n6449 19.3944
R15447 gnd.n6449 gnd.n6448 19.3944
R15448 gnd.n6448 gnd.n1126 19.3944
R15449 gnd.n6444 gnd.n1126 19.3944
R15450 gnd.n6444 gnd.n6443 19.3944
R15451 gnd.n6443 gnd.n6442 19.3944
R15452 gnd.n6442 gnd.n1131 19.3944
R15453 gnd.n6438 gnd.n1131 19.3944
R15454 gnd.n6438 gnd.n6437 19.3944
R15455 gnd.n6437 gnd.n6436 19.3944
R15456 gnd.n6436 gnd.n1136 19.3944
R15457 gnd.n6432 gnd.n1136 19.3944
R15458 gnd.n6432 gnd.n6431 19.3944
R15459 gnd.n6431 gnd.n6430 19.3944
R15460 gnd.n6430 gnd.n1141 19.3944
R15461 gnd.n6426 gnd.n1141 19.3944
R15462 gnd.n6426 gnd.n6425 19.3944
R15463 gnd.n6425 gnd.n6424 19.3944
R15464 gnd.n6424 gnd.n1146 19.3944
R15465 gnd.n6420 gnd.n1146 19.3944
R15466 gnd.n6420 gnd.n6419 19.3944
R15467 gnd.n6419 gnd.n6418 19.3944
R15468 gnd.n6418 gnd.n1151 19.3944
R15469 gnd.n6414 gnd.n1151 19.3944
R15470 gnd.n6414 gnd.n6413 19.3944
R15471 gnd.n6413 gnd.n6412 19.3944
R15472 gnd.n6412 gnd.n1156 19.3944
R15473 gnd.n6408 gnd.n1156 19.3944
R15474 gnd.n6408 gnd.n6407 19.3944
R15475 gnd.n6407 gnd.n6406 19.3944
R15476 gnd.n6406 gnd.n1161 19.3944
R15477 gnd.n6402 gnd.n1161 19.3944
R15478 gnd.n6402 gnd.n6401 19.3944
R15479 gnd.n6401 gnd.n6400 19.3944
R15480 gnd.n6400 gnd.n1166 19.3944
R15481 gnd.n6396 gnd.n1166 19.3944
R15482 gnd.n6396 gnd.n6395 19.3944
R15483 gnd.n6395 gnd.n6394 19.3944
R15484 gnd.n6394 gnd.n1171 19.3944
R15485 gnd.n6390 gnd.n1171 19.3944
R15486 gnd.n6390 gnd.n6389 19.3944
R15487 gnd.n6389 gnd.n6388 19.3944
R15488 gnd.n6388 gnd.n1176 19.3944
R15489 gnd.n6384 gnd.n1176 19.3944
R15490 gnd.n6384 gnd.n6383 19.3944
R15491 gnd.n6383 gnd.n6382 19.3944
R15492 gnd.n6382 gnd.n1181 19.3944
R15493 gnd.n6378 gnd.n1181 19.3944
R15494 gnd.n6378 gnd.n6377 19.3944
R15495 gnd.n6377 gnd.n6376 19.3944
R15496 gnd.n6376 gnd.n1186 19.3944
R15497 gnd.n6372 gnd.n1186 19.3944
R15498 gnd.n6372 gnd.n6371 19.3944
R15499 gnd.n6371 gnd.n6370 19.3944
R15500 gnd.n6370 gnd.n1191 19.3944
R15501 gnd.n6366 gnd.n1191 19.3944
R15502 gnd.n6366 gnd.n6365 19.3944
R15503 gnd.n6365 gnd.n6364 19.3944
R15504 gnd.n6364 gnd.n1196 19.3944
R15505 gnd.n6360 gnd.n1196 19.3944
R15506 gnd.n6360 gnd.n6359 19.3944
R15507 gnd.n6359 gnd.n6358 19.3944
R15508 gnd.n6358 gnd.n1201 19.3944
R15509 gnd.n6354 gnd.n1201 19.3944
R15510 gnd.n6354 gnd.n6353 19.3944
R15511 gnd.n6353 gnd.n6352 19.3944
R15512 gnd.n6352 gnd.n1206 19.3944
R15513 gnd.n6348 gnd.n1206 19.3944
R15514 gnd.n6348 gnd.n6347 19.3944
R15515 gnd.n6347 gnd.n6346 19.3944
R15516 gnd.n6346 gnd.n1211 19.3944
R15517 gnd.n6342 gnd.n1211 19.3944
R15518 gnd.n6342 gnd.n6341 19.3944
R15519 gnd.n6341 gnd.n6340 19.3944
R15520 gnd.n6340 gnd.n1216 19.3944
R15521 gnd.n6336 gnd.n1216 19.3944
R15522 gnd.n6336 gnd.n6335 19.3944
R15523 gnd.n6335 gnd.n6334 19.3944
R15524 gnd.n6334 gnd.n1221 19.3944
R15525 gnd.n6330 gnd.n1221 19.3944
R15526 gnd.n6330 gnd.n6329 19.3944
R15527 gnd.n6329 gnd.n6328 19.3944
R15528 gnd.n6328 gnd.n1226 19.3944
R15529 gnd.n6324 gnd.n1226 19.3944
R15530 gnd.n6324 gnd.n6323 19.3944
R15531 gnd.n6323 gnd.n6322 19.3944
R15532 gnd.n6322 gnd.n1231 19.3944
R15533 gnd.n6318 gnd.n1231 19.3944
R15534 gnd.n6318 gnd.n6317 19.3944
R15535 gnd.n6317 gnd.n6316 19.3944
R15536 gnd.n6316 gnd.n1236 19.3944
R15537 gnd.n6312 gnd.n1236 19.3944
R15538 gnd.n6312 gnd.n6311 19.3944
R15539 gnd.n6311 gnd.n6310 19.3944
R15540 gnd.n6310 gnd.n1241 19.3944
R15541 gnd.n6306 gnd.n1241 19.3944
R15542 gnd.n6306 gnd.n6305 19.3944
R15543 gnd.n6028 gnd.n1614 19.3944
R15544 gnd.n6024 gnd.n1614 19.3944
R15545 gnd.n6024 gnd.n6023 19.3944
R15546 gnd.n1530 gnd.n1514 19.3944
R15547 gnd.n1530 gnd.n1512 19.3944
R15548 gnd.n1536 gnd.n1512 19.3944
R15549 gnd.n1536 gnd.n1507 19.3944
R15550 gnd.n1549 gnd.n1507 19.3944
R15551 gnd.n1549 gnd.n1505 19.3944
R15552 gnd.n1555 gnd.n1505 19.3944
R15553 gnd.n1555 gnd.n1500 19.3944
R15554 gnd.n1568 gnd.n1500 19.3944
R15555 gnd.n1568 gnd.n1498 19.3944
R15556 gnd.n1574 gnd.n1498 19.3944
R15557 gnd.n1574 gnd.n1494 19.3944
R15558 gnd.n1584 gnd.n1494 19.3944
R15559 gnd.n1584 gnd.n1492 19.3944
R15560 gnd.n1590 gnd.n1492 19.3944
R15561 gnd.n1590 gnd.n1482 19.3944
R15562 gnd.n1598 gnd.n1482 19.3944
R15563 gnd.n1598 gnd.n1480 19.3944
R15564 gnd.n6039 gnd.n1480 19.3944
R15565 gnd.n6039 gnd.n6038 19.3944
R15566 gnd.n6038 gnd.n6037 19.3944
R15567 gnd.n6037 gnd.n1606 19.3944
R15568 gnd.n6033 gnd.n1606 19.3944
R15569 gnd.n6033 gnd.n6032 19.3944
R15570 gnd.n6551 gnd.n962 19.1977
R15571 gnd.t77 gnd.n5363 19.1199
R15572 gnd.n5283 gnd.t32 19.1199
R15573 gnd.n3194 gnd.t44 18.8012
R15574 gnd.n3179 gnd.t94 18.8012
R15575 gnd.n3038 gnd.n3037 18.4825
R15576 gnd.n5759 gnd.n1843 18.4825
R15577 gnd.n5799 gnd.n1804 18.4825
R15578 gnd.n5312 gnd.n1775 18.4825
R15579 gnd.n4914 gnd.n1747 18.4825
R15580 gnd.n6263 gnd.n6262 18.4247
R15581 gnd.n5528 gnd.n5527 18.4247
R15582 gnd.n7681 gnd.n124 18.2308
R15583 gnd.n1594 gnd.n1593 18.2308
R15584 gnd.n5566 gnd.n2033 18.2308
R15585 gnd.n3871 gnd.n3815 18.2308
R15586 gnd.t332 gnd.n2718 18.1639
R15587 gnd.t289 gnd.n1914 17.8452
R15588 gnd.n2746 gnd.t46 17.5266
R15589 gnd.n5523 gnd.t58 17.2079
R15590 gnd.n5671 gnd.n1920 17.2079
R15591 gnd.n5437 gnd.n1905 17.2079
R15592 gnd.n4804 gnd.n1864 17.2079
R15593 gnd.n5751 gnd.n1851 17.2079
R15594 gnd.n5807 gnd.n1797 17.2079
R15595 gnd.n4875 gnd.n4873 17.2079
R15596 gnd.n5270 gnd.n5269 17.2079
R15597 gnd.n5887 gnd.n1725 17.2079
R15598 gnd.n3145 gnd.t13 16.8893
R15599 gnd.t129 gnd.n1849 16.8893
R15600 gnd.n5268 gnd.t132 16.8893
R15601 gnd.n2973 gnd.t275 16.2519
R15602 gnd.n2673 gnd.t14 16.2519
R15603 gnd.n5679 gnd.n1913 15.9333
R15604 gnd.n5430 gnd.t210 15.9333
R15605 gnd.n5380 gnd.n5379 15.9333
R15606 gnd.n5357 gnd.t198 15.9333
R15607 gnd.n5327 gnd.n1789 15.9333
R15608 gnd.n5815 gnd.n1789 15.9333
R15609 gnd.t28 gnd.n1753 15.9333
R15610 gnd.n5879 gnd.n1733 15.9333
R15611 gnd.t239 gnd.n1662 15.9333
R15612 gnd.n3660 gnd.n3658 15.6674
R15613 gnd.n3628 gnd.n3626 15.6674
R15614 gnd.n3596 gnd.n3594 15.6674
R15615 gnd.n3565 gnd.n3563 15.6674
R15616 gnd.n3533 gnd.n3531 15.6674
R15617 gnd.n3501 gnd.n3499 15.6674
R15618 gnd.n3469 gnd.n3467 15.6674
R15619 gnd.n3438 gnd.n3436 15.6674
R15620 gnd.n2964 gnd.t275 15.6146
R15621 gnd.t253 gnd.n2415 15.6146
R15622 gnd.t245 gnd.n2416 15.6146
R15623 gnd.n5951 gnd.t231 15.296
R15624 gnd.t200 gnd.n1660 15.296
R15625 gnd.n5010 gnd.n5009 15.0827
R15626 gnd.n4664 gnd.n4659 15.0481
R15627 gnd.n5020 gnd.n5019 15.0481
R15628 gnd.n3332 gnd.t330 14.9773
R15629 gnd.n4760 gnd.t194 14.9773
R15630 gnd.n5935 gnd.t356 14.9773
R15631 gnd.n5687 gnd.n1905 14.6587
R15632 gnd.n5735 gnd.n1864 14.6587
R15633 gnd.n4935 gnd.n1725 14.6587
R15634 gnd.n5218 gnd.n5217 14.6587
R15635 gnd.n5959 gnd.n1660 14.6587
R15636 gnd.t319 gnd.n2458 14.34
R15637 gnd.n3410 gnd.t335 14.34
R15638 gnd.n5400 gnd.t160 14.0214
R15639 gnd.t6 gnd.n1710 14.0214
R15640 gnd.n3120 gnd.t24 13.7027
R15641 gnd.n2830 gnd.n2829 13.5763
R15642 gnd.n3774 gnd.n2371 13.5763
R15643 gnd.n6225 gnd.n1332 13.5763
R15644 gnd.n7733 gnd.n7732 13.5763
R15645 gnd.n4119 gnd.n4034 13.5763
R15646 gnd.n4578 gnd.n4575 13.5763
R15647 gnd.n3038 gnd.n2776 13.384
R15648 gnd.n5452 gnd.t207 13.384
R15649 gnd.n5695 gnd.n1899 13.384
R15650 gnd.n5727 gnd.n1871 13.384
R15651 gnd.n5743 gnd.t196 13.384
R15652 gnd.n4824 gnd.n1843 13.384
R15653 gnd.n5342 gnd.n1804 13.384
R15654 gnd.n5831 gnd.n1775 13.384
R15655 gnd.n5863 gnd.n1747 13.384
R15656 gnd.n4927 gnd.t4 13.384
R15657 gnd.n5248 gnd.n4942 13.384
R15658 gnd.n4962 gnd.n4961 13.384
R15659 gnd.n4675 gnd.n4656 13.1884
R15660 gnd.n4670 gnd.n4669 13.1884
R15661 gnd.n4669 gnd.n4668 13.1884
R15662 gnd.n5013 gnd.n5008 13.1884
R15663 gnd.n5014 gnd.n5013 13.1884
R15664 gnd.n4671 gnd.n4658 13.146
R15665 gnd.n4667 gnd.n4658 13.146
R15666 gnd.n5012 gnd.n5011 13.146
R15667 gnd.n5012 gnd.n5007 13.146
R15668 gnd.t40 gnd.n973 13.0654
R15669 gnd.t38 gnd.n356 13.0654
R15670 gnd.n3661 gnd.n3657 12.8005
R15671 gnd.n3629 gnd.n3625 12.8005
R15672 gnd.n3597 gnd.n3593 12.8005
R15673 gnd.n3566 gnd.n3562 12.8005
R15674 gnd.n3534 gnd.n3530 12.8005
R15675 gnd.n3502 gnd.n3498 12.8005
R15676 gnd.n3470 gnd.n3466 12.8005
R15677 gnd.n3439 gnd.n3435 12.8005
R15678 gnd.t228 gnd.t235 12.7467
R15679 gnd.n5415 gnd.t78 12.7467
R15680 gnd.t327 gnd.n1695 12.7467
R15681 gnd.t260 gnd.n4988 12.7467
R15682 gnd.n2306 gnd.t156 12.4281
R15683 gnd.t34 gnd.n1018 12.4281
R15684 gnd.n4446 gnd.t88 12.4281
R15685 gnd.n5639 gnd.t311 12.4281
R15686 gnd.t221 gnd.t60 12.4281
R15687 gnd.n1640 gnd.t307 12.4281
R15688 gnd.n6111 gnd.t81 12.4281
R15689 gnd.t56 gnd.n399 12.4281
R15690 gnd.t119 gnd.n229 12.4281
R15691 gnd.n2829 gnd.n2824 12.4126
R15692 gnd.n3777 gnd.n3774 12.4126
R15693 gnd.n6221 gnd.n1332 12.4126
R15694 gnd.n7732 gnd.n200 12.4126
R15695 gnd.n4115 gnd.n4034 12.4126
R15696 gnd.n4575 gnd.n2119 12.4126
R15697 gnd.n5520 gnd.n5457 12.1761
R15698 gnd.n5193 gnd.n5192 12.1761
R15699 gnd.n5556 gnd.n2042 12.1094
R15700 gnd.n5703 gnd.n1891 12.1094
R15701 gnd.n5719 gnd.n1879 12.1094
R15702 gnd.n4833 gnd.n1836 12.1094
R15703 gnd.n4852 gnd.n1812 12.1094
R15704 gnd.n5839 gnd.n1768 12.1094
R15705 gnd.n5855 gnd.n1754 12.1094
R15706 gnd.n4949 gnd.n1711 12.1094
R15707 gnd.n4972 gnd.n1686 12.1094
R15708 gnd.n6294 gnd.n1285 12.1094
R15709 gnd.n3665 gnd.n3664 12.0247
R15710 gnd.n3633 gnd.n3632 12.0247
R15711 gnd.n3601 gnd.n3600 12.0247
R15712 gnd.n3570 gnd.n3569 12.0247
R15713 gnd.n3538 gnd.n3537 12.0247
R15714 gnd.n3506 gnd.n3505 12.0247
R15715 gnd.n3474 gnd.n3473 12.0247
R15716 gnd.n3443 gnd.n3442 12.0247
R15717 gnd.n2274 gnd.t22 11.7908
R15718 gnd.n4393 gnd.t34 11.7908
R15719 gnd.t88 gnd.n1060 11.7908
R15720 gnd.t81 gnd.n6109 11.7908
R15721 gnd.n6138 gnd.t56 11.7908
R15722 gnd.t109 gnd.n260 11.7908
R15723 gnd.n3668 gnd.n3655 11.249
R15724 gnd.n3636 gnd.n3623 11.249
R15725 gnd.n3604 gnd.n3591 11.249
R15726 gnd.n3573 gnd.n3560 11.249
R15727 gnd.n3541 gnd.n3528 11.249
R15728 gnd.n3509 gnd.n3496 11.249
R15729 gnd.n3477 gnd.n3464 11.249
R15730 gnd.n3446 gnd.n3433 11.249
R15731 gnd.n3108 gnd.t24 11.1535
R15732 gnd.n2242 gnd.t102 11.1535
R15733 gnd.n4359 gnd.t40 11.1535
R15734 gnd.n7408 gnd.t38 11.1535
R15735 gnd.t192 gnd.n290 11.1535
R15736 gnd.n5711 gnd.n1885 10.8348
R15737 gnd.t161 gnd.n1851 10.8348
R15738 gnd.n1829 gnd.n1828 10.8348
R15739 gnd.n1828 gnd.n1819 10.8348
R15740 gnd.n5847 gnd.n1760 10.8348
R15741 gnd.n5847 gnd.n1762 10.8348
R15742 gnd.n5270 gnd.t115 10.8348
R15743 gnd.n1703 gnd.n1694 10.8348
R15744 gnd.n5128 gnd.n5050 10.6151
R15745 gnd.n5128 gnd.n5127 10.6151
R15746 gnd.n5125 gnd.n5054 10.6151
R15747 gnd.n5120 gnd.n5054 10.6151
R15748 gnd.n5120 gnd.n5119 10.6151
R15749 gnd.n5119 gnd.n5118 10.6151
R15750 gnd.n5118 gnd.n5057 10.6151
R15751 gnd.n5113 gnd.n5057 10.6151
R15752 gnd.n5113 gnd.n5112 10.6151
R15753 gnd.n5112 gnd.n5111 10.6151
R15754 gnd.n5111 gnd.n5060 10.6151
R15755 gnd.n5106 gnd.n5060 10.6151
R15756 gnd.n5106 gnd.n5105 10.6151
R15757 gnd.n5105 gnd.n5104 10.6151
R15758 gnd.n5104 gnd.n5063 10.6151
R15759 gnd.n5099 gnd.n5063 10.6151
R15760 gnd.n5099 gnd.n5098 10.6151
R15761 gnd.n5098 gnd.n5097 10.6151
R15762 gnd.n5097 gnd.n5066 10.6151
R15763 gnd.n5092 gnd.n5066 10.6151
R15764 gnd.n5092 gnd.n5091 10.6151
R15765 gnd.n5091 gnd.n5090 10.6151
R15766 gnd.n5090 gnd.n5069 10.6151
R15767 gnd.n5085 gnd.n5069 10.6151
R15768 gnd.n5085 gnd.n5084 10.6151
R15769 gnd.n5084 gnd.n5083 10.6151
R15770 gnd.n5083 gnd.n5072 10.6151
R15771 gnd.n5078 gnd.n5072 10.6151
R15772 gnd.n5078 gnd.n5077 10.6151
R15773 gnd.n5077 gnd.n5076 10.6151
R15774 gnd.n5450 gnd.n4745 10.6151
R15775 gnd.n5450 gnd.n5449 10.6151
R15776 gnd.n5449 gnd.n5448 10.6151
R15777 gnd.n5448 gnd.n4746 10.6151
R15778 gnd.n4756 gnd.n4746 10.6151
R15779 gnd.n4757 gnd.n4756 10.6151
R15780 gnd.n5435 gnd.n4757 10.6151
R15781 gnd.n5435 gnd.n5434 10.6151
R15782 gnd.n5434 gnd.n5433 10.6151
R15783 gnd.n5433 gnd.n4758 10.6151
R15784 gnd.n4769 gnd.n4758 10.6151
R15785 gnd.n4770 gnd.n4769 10.6151
R15786 gnd.n5420 gnd.n4770 10.6151
R15787 gnd.n5420 gnd.n5419 10.6151
R15788 gnd.n5419 gnd.n5418 10.6151
R15789 gnd.n5418 gnd.n4771 10.6151
R15790 gnd.n4783 gnd.n4771 10.6151
R15791 gnd.n4784 gnd.n4783 10.6151
R15792 gnd.n5405 gnd.n4784 10.6151
R15793 gnd.n5405 gnd.n5404 10.6151
R15794 gnd.n5404 gnd.n5403 10.6151
R15795 gnd.n5403 gnd.n4785 10.6151
R15796 gnd.n4798 gnd.n4785 10.6151
R15797 gnd.n4800 gnd.n4798 10.6151
R15798 gnd.n4801 gnd.n4800 10.6151
R15799 gnd.n5390 gnd.n4801 10.6151
R15800 gnd.n5390 gnd.n5389 10.6151
R15801 gnd.n5389 gnd.n5388 10.6151
R15802 gnd.n5388 gnd.n4802 10.6151
R15803 gnd.n4813 gnd.n4802 10.6151
R15804 gnd.n5376 gnd.n4813 10.6151
R15805 gnd.n5376 gnd.n5375 10.6151
R15806 gnd.n5375 gnd.n5374 10.6151
R15807 gnd.n5374 gnd.n4814 10.6151
R15808 gnd.n4827 gnd.n4814 10.6151
R15809 gnd.n4829 gnd.n4827 10.6151
R15810 gnd.n4830 gnd.n4829 10.6151
R15811 gnd.n5361 gnd.n4830 10.6151
R15812 gnd.n5361 gnd.n5360 10.6151
R15813 gnd.n5360 gnd.n5359 10.6151
R15814 gnd.n5359 gnd.n4831 10.6151
R15815 gnd.n4848 gnd.n4831 10.6151
R15816 gnd.n4849 gnd.n4848 10.6151
R15817 gnd.n4850 gnd.n4849 10.6151
R15818 gnd.n4850 gnd.n4845 10.6151
R15819 gnd.n4856 gnd.n4845 10.6151
R15820 gnd.n4857 gnd.n4856 10.6151
R15821 gnd.n5340 gnd.n4857 10.6151
R15822 gnd.n5340 gnd.n5339 10.6151
R15823 gnd.n5339 gnd.n5338 10.6151
R15824 gnd.n5338 gnd.n4858 10.6151
R15825 gnd.n4869 gnd.n4858 10.6151
R15826 gnd.n4870 gnd.n4869 10.6151
R15827 gnd.n5325 gnd.n4870 10.6151
R15828 gnd.n5325 gnd.n5324 10.6151
R15829 gnd.n5324 gnd.n5323 10.6151
R15830 gnd.n5323 gnd.n4871 10.6151
R15831 gnd.n4883 gnd.n4871 10.6151
R15832 gnd.n4884 gnd.n4883 10.6151
R15833 gnd.n5310 gnd.n4884 10.6151
R15834 gnd.n5310 gnd.n5309 10.6151
R15835 gnd.n5309 gnd.n5308 10.6151
R15836 gnd.n5308 gnd.n4885 10.6151
R15837 gnd.n4896 gnd.n4885 10.6151
R15838 gnd.n4897 gnd.n4896 10.6151
R15839 gnd.n5295 gnd.n4897 10.6151
R15840 gnd.n5295 gnd.n5294 10.6151
R15841 gnd.n5294 gnd.n5293 10.6151
R15842 gnd.n5293 gnd.n4898 10.6151
R15843 gnd.n4910 gnd.n4898 10.6151
R15844 gnd.n4911 gnd.n4910 10.6151
R15845 gnd.n5281 gnd.n4911 10.6151
R15846 gnd.n5281 gnd.n5280 10.6151
R15847 gnd.n5280 gnd.n5279 10.6151
R15848 gnd.n5279 gnd.n4912 10.6151
R15849 gnd.n4923 gnd.n4912 10.6151
R15850 gnd.n4924 gnd.n4923 10.6151
R15851 gnd.n5266 gnd.n4924 10.6151
R15852 gnd.n5266 gnd.n5265 10.6151
R15853 gnd.n5265 gnd.n5264 10.6151
R15854 gnd.n5264 gnd.n4925 10.6151
R15855 gnd.n4938 gnd.n4925 10.6151
R15856 gnd.n4939 gnd.n4938 10.6151
R15857 gnd.n5252 gnd.n4939 10.6151
R15858 gnd.n5252 gnd.n5251 10.6151
R15859 gnd.n5251 gnd.n5250 10.6151
R15860 gnd.n5250 gnd.n4940 10.6151
R15861 gnd.n4953 gnd.n4940 10.6151
R15862 gnd.n4954 gnd.n4953 10.6151
R15863 gnd.n5238 gnd.n4954 10.6151
R15864 gnd.n5238 gnd.n5237 10.6151
R15865 gnd.n5237 gnd.n5236 10.6151
R15866 gnd.n5236 gnd.n4955 10.6151
R15867 gnd.n5232 gnd.n4955 10.6151
R15868 gnd.n5232 gnd.n5231 10.6151
R15869 gnd.n5231 gnd.n5230 10.6151
R15870 gnd.n5230 gnd.n4957 10.6151
R15871 gnd.n4959 gnd.n4957 10.6151
R15872 gnd.n4982 gnd.n4959 10.6151
R15873 gnd.n4984 gnd.n4982 10.6151
R15874 gnd.n4985 gnd.n4984 10.6151
R15875 gnd.n5215 gnd.n4985 10.6151
R15876 gnd.n5215 gnd.n5214 10.6151
R15877 gnd.n5214 gnd.n5213 10.6151
R15878 gnd.n5213 gnd.n4986 10.6151
R15879 gnd.n4998 gnd.n4986 10.6151
R15880 gnd.n5201 gnd.n4998 10.6151
R15881 gnd.n5201 gnd.n5200 10.6151
R15882 gnd.n5200 gnd.n5199 10.6151
R15883 gnd.n5199 gnd.n4999 10.6151
R15884 gnd.n4682 gnd.n4617 10.6151
R15885 gnd.n4685 gnd.n4682 10.6151
R15886 gnd.n4690 gnd.n4687 10.6151
R15887 gnd.n4691 gnd.n4690 10.6151
R15888 gnd.n4694 gnd.n4691 10.6151
R15889 gnd.n4695 gnd.n4694 10.6151
R15890 gnd.n4698 gnd.n4695 10.6151
R15891 gnd.n4699 gnd.n4698 10.6151
R15892 gnd.n4702 gnd.n4699 10.6151
R15893 gnd.n4703 gnd.n4702 10.6151
R15894 gnd.n4706 gnd.n4703 10.6151
R15895 gnd.n4707 gnd.n4706 10.6151
R15896 gnd.n4710 gnd.n4707 10.6151
R15897 gnd.n4711 gnd.n4710 10.6151
R15898 gnd.n4714 gnd.n4711 10.6151
R15899 gnd.n4715 gnd.n4714 10.6151
R15900 gnd.n4718 gnd.n4715 10.6151
R15901 gnd.n4719 gnd.n4718 10.6151
R15902 gnd.n4722 gnd.n4719 10.6151
R15903 gnd.n4723 gnd.n4722 10.6151
R15904 gnd.n4726 gnd.n4723 10.6151
R15905 gnd.n4727 gnd.n4726 10.6151
R15906 gnd.n4730 gnd.n4727 10.6151
R15907 gnd.n4731 gnd.n4730 10.6151
R15908 gnd.n4734 gnd.n4731 10.6151
R15909 gnd.n4735 gnd.n4734 10.6151
R15910 gnd.n4738 gnd.n4735 10.6151
R15911 gnd.n4739 gnd.n4738 10.6151
R15912 gnd.n4742 gnd.n4739 10.6151
R15913 gnd.n4744 gnd.n4742 10.6151
R15914 gnd.n5520 gnd.n5519 10.6151
R15915 gnd.n5519 gnd.n5518 10.6151
R15916 gnd.n5518 gnd.n5517 10.6151
R15917 gnd.n5517 gnd.n5515 10.6151
R15918 gnd.n5515 gnd.n5512 10.6151
R15919 gnd.n5512 gnd.n5511 10.6151
R15920 gnd.n5511 gnd.n5508 10.6151
R15921 gnd.n5508 gnd.n5507 10.6151
R15922 gnd.n5507 gnd.n5504 10.6151
R15923 gnd.n5504 gnd.n5503 10.6151
R15924 gnd.n5503 gnd.n5500 10.6151
R15925 gnd.n5500 gnd.n5499 10.6151
R15926 gnd.n5499 gnd.n5496 10.6151
R15927 gnd.n5496 gnd.n5495 10.6151
R15928 gnd.n5495 gnd.n5492 10.6151
R15929 gnd.n5492 gnd.n5491 10.6151
R15930 gnd.n5491 gnd.n5488 10.6151
R15931 gnd.n5488 gnd.n5487 10.6151
R15932 gnd.n5487 gnd.n5484 10.6151
R15933 gnd.n5484 gnd.n5483 10.6151
R15934 gnd.n5483 gnd.n5480 10.6151
R15935 gnd.n5480 gnd.n5479 10.6151
R15936 gnd.n5479 gnd.n5476 10.6151
R15937 gnd.n5476 gnd.n5475 10.6151
R15938 gnd.n5475 gnd.n5472 10.6151
R15939 gnd.n5472 gnd.n5471 10.6151
R15940 gnd.n5471 gnd.n5468 10.6151
R15941 gnd.n5468 gnd.n5467 10.6151
R15942 gnd.n5464 gnd.n5463 10.6151
R15943 gnd.n5463 gnd.n4618 10.6151
R15944 gnd.n5192 gnd.n5191 10.6151
R15945 gnd.n5191 gnd.n5025 10.6151
R15946 gnd.n5186 gnd.n5025 10.6151
R15947 gnd.n5186 gnd.n5185 10.6151
R15948 gnd.n5185 gnd.n5184 10.6151
R15949 gnd.n5184 gnd.n5028 10.6151
R15950 gnd.n5179 gnd.n5028 10.6151
R15951 gnd.n5179 gnd.n5178 10.6151
R15952 gnd.n5178 gnd.n5177 10.6151
R15953 gnd.n5177 gnd.n5031 10.6151
R15954 gnd.n5172 gnd.n5031 10.6151
R15955 gnd.n5172 gnd.n5171 10.6151
R15956 gnd.n5171 gnd.n5170 10.6151
R15957 gnd.n5170 gnd.n5034 10.6151
R15958 gnd.n5165 gnd.n5034 10.6151
R15959 gnd.n5165 gnd.n5164 10.6151
R15960 gnd.n5164 gnd.n5163 10.6151
R15961 gnd.n5163 gnd.n5037 10.6151
R15962 gnd.n5158 gnd.n5037 10.6151
R15963 gnd.n5158 gnd.n5157 10.6151
R15964 gnd.n5157 gnd.n5156 10.6151
R15965 gnd.n5156 gnd.n5040 10.6151
R15966 gnd.n5151 gnd.n5040 10.6151
R15967 gnd.n5151 gnd.n5150 10.6151
R15968 gnd.n5150 gnd.n5149 10.6151
R15969 gnd.n5149 gnd.n5043 10.6151
R15970 gnd.n5144 gnd.n5043 10.6151
R15971 gnd.n5144 gnd.n5143 10.6151
R15972 gnd.n5141 gnd.n5048 10.6151
R15973 gnd.n5136 gnd.n5048 10.6151
R15974 gnd.n5456 gnd.n5455 10.6151
R15975 gnd.n5455 gnd.n4676 10.6151
R15976 gnd.n4751 gnd.n4676 10.6151
R15977 gnd.n5443 gnd.n4751 10.6151
R15978 gnd.n5443 gnd.n5442 10.6151
R15979 gnd.n5442 gnd.n5441 10.6151
R15980 gnd.n5441 gnd.n4752 10.6151
R15981 gnd.n4763 gnd.n4752 10.6151
R15982 gnd.n4764 gnd.n4763 10.6151
R15983 gnd.n5428 gnd.n4764 10.6151
R15984 gnd.n5428 gnd.n5427 10.6151
R15985 gnd.n5427 gnd.n5426 10.6151
R15986 gnd.n5426 gnd.n4765 10.6151
R15987 gnd.n4777 gnd.n4765 10.6151
R15988 gnd.n4778 gnd.n4777 10.6151
R15989 gnd.n5413 gnd.n4778 10.6151
R15990 gnd.n5413 gnd.n5412 10.6151
R15991 gnd.n5412 gnd.n5411 10.6151
R15992 gnd.n5411 gnd.n4779 10.6151
R15993 gnd.n4791 gnd.n4779 10.6151
R15994 gnd.n4792 gnd.n4791 10.6151
R15995 gnd.n5398 gnd.n4792 10.6151
R15996 gnd.n5398 gnd.n5397 10.6151
R15997 gnd.n5397 gnd.n5396 10.6151
R15998 gnd.n5396 gnd.n4793 10.6151
R15999 gnd.n4807 gnd.n4793 10.6151
R16000 gnd.n4808 gnd.n4807 10.6151
R16001 gnd.n5384 gnd.n4808 10.6151
R16002 gnd.n5384 gnd.n5383 10.6151
R16003 gnd.n5383 gnd.n5382 10.6151
R16004 gnd.n5382 gnd.n4809 10.6151
R16005 gnd.n4820 gnd.n4809 10.6151
R16006 gnd.n4821 gnd.n4820 10.6151
R16007 gnd.n5369 gnd.n4821 10.6151
R16008 gnd.n5369 gnd.n5368 10.6151
R16009 gnd.n5368 gnd.n5367 10.6151
R16010 gnd.n5367 gnd.n4822 10.6151
R16011 gnd.n4836 gnd.n4822 10.6151
R16012 gnd.n4837 gnd.n4836 10.6151
R16013 gnd.n5355 gnd.n4837 10.6151
R16014 gnd.n5355 gnd.n5354 10.6151
R16015 gnd.n5354 gnd.n5353 10.6151
R16016 gnd.n5353 gnd.n4838 10.6151
R16017 gnd.n5349 gnd.n4838 10.6151
R16018 gnd.n5349 gnd.n5348 10.6151
R16019 gnd.n5348 gnd.n5347 10.6151
R16020 gnd.n5347 gnd.n4840 10.6151
R16021 gnd.n4842 gnd.n4840 10.6151
R16022 gnd.n4863 gnd.n4842 10.6151
R16023 gnd.n4864 gnd.n4863 10.6151
R16024 gnd.n5333 gnd.n4864 10.6151
R16025 gnd.n5333 gnd.n5332 10.6151
R16026 gnd.n5332 gnd.n5331 10.6151
R16027 gnd.n5331 gnd.n4865 10.6151
R16028 gnd.n4877 gnd.n4865 10.6151
R16029 gnd.n4878 gnd.n4877 10.6151
R16030 gnd.n5318 gnd.n4878 10.6151
R16031 gnd.n5318 gnd.n5317 10.6151
R16032 gnd.n5317 gnd.n5316 10.6151
R16033 gnd.n5316 gnd.n4879 10.6151
R16034 gnd.n4890 gnd.n4879 10.6151
R16035 gnd.n4891 gnd.n4890 10.6151
R16036 gnd.n5303 gnd.n4891 10.6151
R16037 gnd.n5303 gnd.n5302 10.6151
R16038 gnd.n5302 gnd.n5301 10.6151
R16039 gnd.n5301 gnd.n4892 10.6151
R16040 gnd.n4903 gnd.n4892 10.6151
R16041 gnd.n4904 gnd.n4903 10.6151
R16042 gnd.n5288 gnd.n4904 10.6151
R16043 gnd.n5288 gnd.n5287 10.6151
R16044 gnd.n5287 gnd.n5286 10.6151
R16045 gnd.n5286 gnd.n4905 10.6151
R16046 gnd.n4917 gnd.n4905 10.6151
R16047 gnd.n4918 gnd.n4917 10.6151
R16048 gnd.n5274 gnd.n4918 10.6151
R16049 gnd.n5274 gnd.n5273 10.6151
R16050 gnd.n5273 gnd.n5272 10.6151
R16051 gnd.n5272 gnd.n4919 10.6151
R16052 gnd.n4931 gnd.n4919 10.6151
R16053 gnd.n4932 gnd.n4931 10.6151
R16054 gnd.n5259 gnd.n4932 10.6151
R16055 gnd.n5259 gnd.n5258 10.6151
R16056 gnd.n5258 gnd.n5257 10.6151
R16057 gnd.n5257 gnd.n4933 10.6151
R16058 gnd.n4945 gnd.n4933 10.6151
R16059 gnd.n5246 gnd.n4945 10.6151
R16060 gnd.n5246 gnd.n5245 10.6151
R16061 gnd.n5245 gnd.n5244 10.6151
R16062 gnd.n5244 gnd.n4946 10.6151
R16063 gnd.n4948 gnd.n4946 10.6151
R16064 gnd.n4966 gnd.n4948 10.6151
R16065 gnd.n4968 gnd.n4966 10.6151
R16066 gnd.n4969 gnd.n4968 10.6151
R16067 gnd.n4970 gnd.n4969 10.6151
R16068 gnd.n4970 gnd.n4964 10.6151
R16069 gnd.n4976 gnd.n4964 10.6151
R16070 gnd.n4977 gnd.n4976 10.6151
R16071 gnd.n5224 gnd.n4977 10.6151
R16072 gnd.n5224 gnd.n5223 10.6151
R16073 gnd.n5223 gnd.n5222 10.6151
R16074 gnd.n5222 gnd.n4978 10.6151
R16075 gnd.n4992 gnd.n4978 10.6151
R16076 gnd.n4993 gnd.n4992 10.6151
R16077 gnd.n5209 gnd.n4993 10.6151
R16078 gnd.n5209 gnd.n5208 10.6151
R16079 gnd.n5208 gnd.n5207 10.6151
R16080 gnd.n5207 gnd.n4994 10.6151
R16081 gnd.n5004 gnd.n4994 10.6151
R16082 gnd.n5005 gnd.n5004 10.6151
R16083 gnd.n5194 gnd.n5005 10.6151
R16084 gnd.n3027 gnd.t162 10.5161
R16085 gnd.n2460 gnd.t319 10.5161
R16086 gnd.n3393 gnd.t335 10.5161
R16087 gnd.t36 gnd.n2209 10.5161
R16088 gnd.n2211 gnd.t86 10.5161
R16089 gnd.n7453 gnd.t79 10.5161
R16090 gnd.n7459 gnd.t147 10.5161
R16091 gnd.n3669 gnd.n3653 10.4732
R16092 gnd.n3637 gnd.n3621 10.4732
R16093 gnd.n3605 gnd.n3589 10.4732
R16094 gnd.n3574 gnd.n3558 10.4732
R16095 gnd.n3542 gnd.n3526 10.4732
R16096 gnd.n3510 gnd.n3494 10.4732
R16097 gnd.n3478 gnd.n3462 10.4732
R16098 gnd.n3447 gnd.n3431 10.4732
R16099 gnd.t330 gnd.n2477 9.87883
R16100 gnd.t100 gnd.n2239 9.87883
R16101 gnd.t358 gnd.t164 9.87883
R16102 gnd.t33 gnd.t309 9.87883
R16103 gnd.n293 gnd.t188 9.87883
R16104 gnd.n7858 gnd.n78 9.81789
R16105 gnd.n3673 gnd.n3672 9.69747
R16106 gnd.n3641 gnd.n3640 9.69747
R16107 gnd.n3609 gnd.n3608 9.69747
R16108 gnd.n3578 gnd.n3577 9.69747
R16109 gnd.n3546 gnd.n3545 9.69747
R16110 gnd.n3514 gnd.n3513 9.69747
R16111 gnd.n3482 gnd.n3481 9.69747
R16112 gnd.n3451 gnd.n3450 9.69747
R16113 gnd.n5703 gnd.n1893 9.56018
R16114 gnd.n5719 gnd.n1877 9.56018
R16115 gnd.n5357 gnd.n4833 9.56018
R16116 gnd.n4853 gnd.n4852 9.56018
R16117 gnd.n5839 gnd.n1769 9.56018
R16118 gnd.n5855 gnd.n1753 9.56018
R16119 gnd.n5240 gnd.n4949 9.56018
R16120 gnd.n4973 gnd.n4972 9.56018
R16121 gnd.n6459 gnd.n1115 9.45751
R16122 gnd.n1517 gnd.n1342 9.45599
R16123 gnd.n3679 gnd.n3678 9.45567
R16124 gnd.n3647 gnd.n3646 9.45567
R16125 gnd.n3615 gnd.n3614 9.45567
R16126 gnd.n3584 gnd.n3583 9.45567
R16127 gnd.n3552 gnd.n3551 9.45567
R16128 gnd.n3520 gnd.n3519 9.45567
R16129 gnd.n3488 gnd.n3487 9.45567
R16130 gnd.n3457 gnd.n3456 9.45567
R16131 gnd.n2625 gnd.n2624 9.39724
R16132 gnd.n3678 gnd.n3677 9.3005
R16133 gnd.n3651 gnd.n3650 9.3005
R16134 gnd.n3672 gnd.n3671 9.3005
R16135 gnd.n3670 gnd.n3669 9.3005
R16136 gnd.n3655 gnd.n3654 9.3005
R16137 gnd.n3664 gnd.n3663 9.3005
R16138 gnd.n3662 gnd.n3661 9.3005
R16139 gnd.n3646 gnd.n3645 9.3005
R16140 gnd.n3619 gnd.n3618 9.3005
R16141 gnd.n3640 gnd.n3639 9.3005
R16142 gnd.n3638 gnd.n3637 9.3005
R16143 gnd.n3623 gnd.n3622 9.3005
R16144 gnd.n3632 gnd.n3631 9.3005
R16145 gnd.n3630 gnd.n3629 9.3005
R16146 gnd.n3614 gnd.n3613 9.3005
R16147 gnd.n3587 gnd.n3586 9.3005
R16148 gnd.n3608 gnd.n3607 9.3005
R16149 gnd.n3606 gnd.n3605 9.3005
R16150 gnd.n3591 gnd.n3590 9.3005
R16151 gnd.n3600 gnd.n3599 9.3005
R16152 gnd.n3598 gnd.n3597 9.3005
R16153 gnd.n3583 gnd.n3582 9.3005
R16154 gnd.n3556 gnd.n3555 9.3005
R16155 gnd.n3577 gnd.n3576 9.3005
R16156 gnd.n3575 gnd.n3574 9.3005
R16157 gnd.n3560 gnd.n3559 9.3005
R16158 gnd.n3569 gnd.n3568 9.3005
R16159 gnd.n3567 gnd.n3566 9.3005
R16160 gnd.n3551 gnd.n3550 9.3005
R16161 gnd.n3524 gnd.n3523 9.3005
R16162 gnd.n3545 gnd.n3544 9.3005
R16163 gnd.n3543 gnd.n3542 9.3005
R16164 gnd.n3528 gnd.n3527 9.3005
R16165 gnd.n3537 gnd.n3536 9.3005
R16166 gnd.n3535 gnd.n3534 9.3005
R16167 gnd.n3519 gnd.n3518 9.3005
R16168 gnd.n3492 gnd.n3491 9.3005
R16169 gnd.n3513 gnd.n3512 9.3005
R16170 gnd.n3511 gnd.n3510 9.3005
R16171 gnd.n3496 gnd.n3495 9.3005
R16172 gnd.n3505 gnd.n3504 9.3005
R16173 gnd.n3503 gnd.n3502 9.3005
R16174 gnd.n3487 gnd.n3486 9.3005
R16175 gnd.n3460 gnd.n3459 9.3005
R16176 gnd.n3481 gnd.n3480 9.3005
R16177 gnd.n3479 gnd.n3478 9.3005
R16178 gnd.n3464 gnd.n3463 9.3005
R16179 gnd.n3473 gnd.n3472 9.3005
R16180 gnd.n3471 gnd.n3470 9.3005
R16181 gnd.n3456 gnd.n3455 9.3005
R16182 gnd.n3429 gnd.n3428 9.3005
R16183 gnd.n3450 gnd.n3449 9.3005
R16184 gnd.n3448 gnd.n3447 9.3005
R16185 gnd.n3433 gnd.n3432 9.3005
R16186 gnd.n3442 gnd.n3441 9.3005
R16187 gnd.n3440 gnd.n3439 9.3005
R16188 gnd.n3804 gnd.n3803 9.3005
R16189 gnd.n3802 gnd.n2359 9.3005
R16190 gnd.n3801 gnd.n3800 9.3005
R16191 gnd.n3797 gnd.n2360 9.3005
R16192 gnd.n3794 gnd.n2361 9.3005
R16193 gnd.n3793 gnd.n2362 9.3005
R16194 gnd.n3790 gnd.n2363 9.3005
R16195 gnd.n3789 gnd.n2364 9.3005
R16196 gnd.n3786 gnd.n2365 9.3005
R16197 gnd.n3785 gnd.n2366 9.3005
R16198 gnd.n3782 gnd.n2367 9.3005
R16199 gnd.n3781 gnd.n2368 9.3005
R16200 gnd.n3778 gnd.n2369 9.3005
R16201 gnd.n3777 gnd.n2370 9.3005
R16202 gnd.n3774 gnd.n3773 9.3005
R16203 gnd.n3772 gnd.n2371 9.3005
R16204 gnd.n3805 gnd.n2358 9.3005
R16205 gnd.n3046 gnd.n3045 9.3005
R16206 gnd.n2750 gnd.n2749 9.3005
R16207 gnd.n3073 gnd.n3072 9.3005
R16208 gnd.n3074 gnd.n2748 9.3005
R16209 gnd.n3078 gnd.n3075 9.3005
R16210 gnd.n3077 gnd.n3076 9.3005
R16211 gnd.n2722 gnd.n2721 9.3005
R16212 gnd.n3103 gnd.n3102 9.3005
R16213 gnd.n3104 gnd.n2720 9.3005
R16214 gnd.n3106 gnd.n3105 9.3005
R16215 gnd.n2700 gnd.n2699 9.3005
R16216 gnd.n3134 gnd.n3133 9.3005
R16217 gnd.n3135 gnd.n2698 9.3005
R16218 gnd.n3143 gnd.n3136 9.3005
R16219 gnd.n3142 gnd.n3137 9.3005
R16220 gnd.n3141 gnd.n3139 9.3005
R16221 gnd.n3138 gnd.n2647 9.3005
R16222 gnd.n3191 gnd.n2648 9.3005
R16223 gnd.n3190 gnd.n2649 9.3005
R16224 gnd.n3189 gnd.n2650 9.3005
R16225 gnd.n2669 gnd.n2651 9.3005
R16226 gnd.n2671 gnd.n2670 9.3005
R16227 gnd.n2557 gnd.n2556 9.3005
R16228 gnd.n3229 gnd.n3228 9.3005
R16229 gnd.n3230 gnd.n2555 9.3005
R16230 gnd.n3234 gnd.n3231 9.3005
R16231 gnd.n3233 gnd.n3232 9.3005
R16232 gnd.n2530 gnd.n2529 9.3005
R16233 gnd.n3269 gnd.n3268 9.3005
R16234 gnd.n3270 gnd.n2528 9.3005
R16235 gnd.n3274 gnd.n3271 9.3005
R16236 gnd.n3273 gnd.n3272 9.3005
R16237 gnd.n2503 gnd.n2502 9.3005
R16238 gnd.n3314 gnd.n3313 9.3005
R16239 gnd.n3315 gnd.n2501 9.3005
R16240 gnd.n3319 gnd.n3316 9.3005
R16241 gnd.n3318 gnd.n3317 9.3005
R16242 gnd.n2475 gnd.n2474 9.3005
R16243 gnd.n3354 gnd.n3353 9.3005
R16244 gnd.n3355 gnd.n2473 9.3005
R16245 gnd.n3359 gnd.n3356 9.3005
R16246 gnd.n3358 gnd.n3357 9.3005
R16247 gnd.n2448 gnd.n2447 9.3005
R16248 gnd.n3403 gnd.n3402 9.3005
R16249 gnd.n3404 gnd.n2446 9.3005
R16250 gnd.n3408 gnd.n3405 9.3005
R16251 gnd.n3407 gnd.n3406 9.3005
R16252 gnd.n2421 gnd.n2420 9.3005
R16253 gnd.n3697 gnd.n3696 9.3005
R16254 gnd.n3698 gnd.n2419 9.3005
R16255 gnd.n3704 gnd.n3699 9.3005
R16256 gnd.n3703 gnd.n3700 9.3005
R16257 gnd.n3702 gnd.n3701 9.3005
R16258 gnd.n3047 gnd.n3044 9.3005
R16259 gnd.n2829 gnd.n2788 9.3005
R16260 gnd.n2824 gnd.n2823 9.3005
R16261 gnd.n2822 gnd.n2789 9.3005
R16262 gnd.n2821 gnd.n2820 9.3005
R16263 gnd.n2817 gnd.n2790 9.3005
R16264 gnd.n2814 gnd.n2813 9.3005
R16265 gnd.n2812 gnd.n2791 9.3005
R16266 gnd.n2811 gnd.n2810 9.3005
R16267 gnd.n2807 gnd.n2792 9.3005
R16268 gnd.n2804 gnd.n2803 9.3005
R16269 gnd.n2802 gnd.n2793 9.3005
R16270 gnd.n2801 gnd.n2800 9.3005
R16271 gnd.n2797 gnd.n2795 9.3005
R16272 gnd.n2794 gnd.n2774 9.3005
R16273 gnd.n3041 gnd.n2773 9.3005
R16274 gnd.n3043 gnd.n3042 9.3005
R16275 gnd.n2831 gnd.n2830 9.3005
R16276 gnd.n3054 gnd.n2760 9.3005
R16277 gnd.n3061 gnd.n2761 9.3005
R16278 gnd.n3063 gnd.n3062 9.3005
R16279 gnd.n3064 gnd.n2741 9.3005
R16280 gnd.n3083 gnd.n3082 9.3005
R16281 gnd.n3085 gnd.n2733 9.3005
R16282 gnd.n3092 gnd.n2735 9.3005
R16283 gnd.n3093 gnd.n2730 9.3005
R16284 gnd.n3095 gnd.n3094 9.3005
R16285 gnd.n2731 gnd.n2716 9.3005
R16286 gnd.n3111 gnd.n2714 9.3005
R16287 gnd.n3115 gnd.n3114 9.3005
R16288 gnd.n3113 gnd.n2690 9.3005
R16289 gnd.n3150 gnd.n2689 9.3005
R16290 gnd.n3153 gnd.n3152 9.3005
R16291 gnd.n2686 gnd.n2685 9.3005
R16292 gnd.n3159 gnd.n2687 9.3005
R16293 gnd.n3161 gnd.n3160 9.3005
R16294 gnd.n3163 gnd.n2684 9.3005
R16295 gnd.n3166 gnd.n3165 9.3005
R16296 gnd.n3169 gnd.n3167 9.3005
R16297 gnd.n3171 gnd.n3170 9.3005
R16298 gnd.n3177 gnd.n3172 9.3005
R16299 gnd.n3176 gnd.n3175 9.3005
R16300 gnd.n2548 gnd.n2547 9.3005
R16301 gnd.n3243 gnd.n3242 9.3005
R16302 gnd.n3244 gnd.n2541 9.3005
R16303 gnd.n3252 gnd.n2540 9.3005
R16304 gnd.n3255 gnd.n3254 9.3005
R16305 gnd.n3257 gnd.n3256 9.3005
R16306 gnd.n3260 gnd.n2523 9.3005
R16307 gnd.n3258 gnd.n2521 9.3005
R16308 gnd.n3280 gnd.n2519 9.3005
R16309 gnd.n3282 gnd.n3281 9.3005
R16310 gnd.n2493 gnd.n2492 9.3005
R16311 gnd.n3328 gnd.n3327 9.3005
R16312 gnd.n3329 gnd.n2486 9.3005
R16313 gnd.n3337 gnd.n2485 9.3005
R16314 gnd.n3340 gnd.n3339 9.3005
R16315 gnd.n3342 gnd.n3341 9.3005
R16316 gnd.n3345 gnd.n2468 9.3005
R16317 gnd.n3343 gnd.n2466 9.3005
R16318 gnd.n3365 gnd.n2464 9.3005
R16319 gnd.n3367 gnd.n3366 9.3005
R16320 gnd.n2439 gnd.n2438 9.3005
R16321 gnd.n3417 gnd.n3416 9.3005
R16322 gnd.n3418 gnd.n2432 9.3005
R16323 gnd.n3426 gnd.n2431 9.3005
R16324 gnd.n3685 gnd.n3684 9.3005
R16325 gnd.n3687 gnd.n3686 9.3005
R16326 gnd.n3688 gnd.n2412 9.3005
R16327 gnd.n3712 gnd.n3711 9.3005
R16328 gnd.n2413 gnd.n2374 9.3005
R16329 gnd.n3052 gnd.n3051 9.3005
R16330 gnd.n3768 gnd.n2375 9.3005
R16331 gnd.n3767 gnd.n2377 9.3005
R16332 gnd.n3764 gnd.n2378 9.3005
R16333 gnd.n3763 gnd.n2379 9.3005
R16334 gnd.n3760 gnd.n2380 9.3005
R16335 gnd.n3759 gnd.n2381 9.3005
R16336 gnd.n3756 gnd.n2382 9.3005
R16337 gnd.n3755 gnd.n2383 9.3005
R16338 gnd.n3752 gnd.n2384 9.3005
R16339 gnd.n3751 gnd.n2385 9.3005
R16340 gnd.n3748 gnd.n2386 9.3005
R16341 gnd.n3747 gnd.n2387 9.3005
R16342 gnd.n3744 gnd.n2388 9.3005
R16343 gnd.n3743 gnd.n2389 9.3005
R16344 gnd.n3740 gnd.n2390 9.3005
R16345 gnd.n3739 gnd.n2391 9.3005
R16346 gnd.n3736 gnd.n2392 9.3005
R16347 gnd.n3735 gnd.n2393 9.3005
R16348 gnd.n3732 gnd.n2394 9.3005
R16349 gnd.n3731 gnd.n2395 9.3005
R16350 gnd.n3728 gnd.n2396 9.3005
R16351 gnd.n3727 gnd.n2397 9.3005
R16352 gnd.n3724 gnd.n2401 9.3005
R16353 gnd.n3723 gnd.n2402 9.3005
R16354 gnd.n3720 gnd.n2403 9.3005
R16355 gnd.n3719 gnd.n2404 9.3005
R16356 gnd.n3770 gnd.n3769 9.3005
R16357 gnd.n3221 gnd.n3205 9.3005
R16358 gnd.n3220 gnd.n3206 9.3005
R16359 gnd.n3219 gnd.n3207 9.3005
R16360 gnd.n3217 gnd.n3208 9.3005
R16361 gnd.n3216 gnd.n3209 9.3005
R16362 gnd.n3214 gnd.n3210 9.3005
R16363 gnd.n3213 gnd.n3211 9.3005
R16364 gnd.n2511 gnd.n2510 9.3005
R16365 gnd.n3290 gnd.n3289 9.3005
R16366 gnd.n3291 gnd.n2509 9.3005
R16367 gnd.n3308 gnd.n3292 9.3005
R16368 gnd.n3307 gnd.n3293 9.3005
R16369 gnd.n3306 gnd.n3294 9.3005
R16370 gnd.n3304 gnd.n3295 9.3005
R16371 gnd.n3303 gnd.n3296 9.3005
R16372 gnd.n3301 gnd.n3297 9.3005
R16373 gnd.n3300 gnd.n3298 9.3005
R16374 gnd.n2455 gnd.n2454 9.3005
R16375 gnd.n3375 gnd.n3374 9.3005
R16376 gnd.n3376 gnd.n2453 9.3005
R16377 gnd.n3397 gnd.n3377 9.3005
R16378 gnd.n3396 gnd.n3378 9.3005
R16379 gnd.n3395 gnd.n3379 9.3005
R16380 gnd.n3392 gnd.n3380 9.3005
R16381 gnd.n3391 gnd.n3381 9.3005
R16382 gnd.n3389 gnd.n3382 9.3005
R16383 gnd.n3388 gnd.n3383 9.3005
R16384 gnd.n3386 gnd.n3385 9.3005
R16385 gnd.n3384 gnd.n2406 9.3005
R16386 gnd.n2962 gnd.n2961 9.3005
R16387 gnd.n2852 gnd.n2851 9.3005
R16388 gnd.n2976 gnd.n2975 9.3005
R16389 gnd.n2977 gnd.n2850 9.3005
R16390 gnd.n2979 gnd.n2978 9.3005
R16391 gnd.n2840 gnd.n2839 9.3005
R16392 gnd.n2992 gnd.n2991 9.3005
R16393 gnd.n2993 gnd.n2838 9.3005
R16394 gnd.n3025 gnd.n2994 9.3005
R16395 gnd.n3024 gnd.n2995 9.3005
R16396 gnd.n3023 gnd.n2996 9.3005
R16397 gnd.n3022 gnd.n2997 9.3005
R16398 gnd.n3019 gnd.n2998 9.3005
R16399 gnd.n3018 gnd.n2999 9.3005
R16400 gnd.n3017 gnd.n3000 9.3005
R16401 gnd.n3015 gnd.n3001 9.3005
R16402 gnd.n3014 gnd.n3002 9.3005
R16403 gnd.n3011 gnd.n3003 9.3005
R16404 gnd.n3010 gnd.n3004 9.3005
R16405 gnd.n3009 gnd.n3005 9.3005
R16406 gnd.n3007 gnd.n3006 9.3005
R16407 gnd.n2706 gnd.n2705 9.3005
R16408 gnd.n3123 gnd.n3122 9.3005
R16409 gnd.n3124 gnd.n2704 9.3005
R16410 gnd.n3128 gnd.n3125 9.3005
R16411 gnd.n3127 gnd.n3126 9.3005
R16412 gnd.n2628 gnd.n2627 9.3005
R16413 gnd.n3203 gnd.n3202 9.3005
R16414 gnd.n2960 gnd.n2861 9.3005
R16415 gnd.n2863 gnd.n2862 9.3005
R16416 gnd.n2907 gnd.n2905 9.3005
R16417 gnd.n2908 gnd.n2904 9.3005
R16418 gnd.n2911 gnd.n2900 9.3005
R16419 gnd.n2912 gnd.n2899 9.3005
R16420 gnd.n2915 gnd.n2898 9.3005
R16421 gnd.n2916 gnd.n2897 9.3005
R16422 gnd.n2919 gnd.n2896 9.3005
R16423 gnd.n2920 gnd.n2895 9.3005
R16424 gnd.n2923 gnd.n2894 9.3005
R16425 gnd.n2924 gnd.n2893 9.3005
R16426 gnd.n2927 gnd.n2892 9.3005
R16427 gnd.n2928 gnd.n2891 9.3005
R16428 gnd.n2931 gnd.n2890 9.3005
R16429 gnd.n2932 gnd.n2889 9.3005
R16430 gnd.n2935 gnd.n2888 9.3005
R16431 gnd.n2936 gnd.n2887 9.3005
R16432 gnd.n2939 gnd.n2886 9.3005
R16433 gnd.n2940 gnd.n2885 9.3005
R16434 gnd.n2943 gnd.n2884 9.3005
R16435 gnd.n2944 gnd.n2883 9.3005
R16436 gnd.n2947 gnd.n2882 9.3005
R16437 gnd.n2949 gnd.n2881 9.3005
R16438 gnd.n2950 gnd.n2880 9.3005
R16439 gnd.n2951 gnd.n2879 9.3005
R16440 gnd.n2952 gnd.n2878 9.3005
R16441 gnd.n2959 gnd.n2958 9.3005
R16442 gnd.n2968 gnd.n2967 9.3005
R16443 gnd.n2969 gnd.n2855 9.3005
R16444 gnd.n2971 gnd.n2970 9.3005
R16445 gnd.n2846 gnd.n2845 9.3005
R16446 gnd.n2984 gnd.n2983 9.3005
R16447 gnd.n2985 gnd.n2844 9.3005
R16448 gnd.n2987 gnd.n2986 9.3005
R16449 gnd.n2833 gnd.n2832 9.3005
R16450 gnd.n3030 gnd.n3029 9.3005
R16451 gnd.n3031 gnd.n2787 9.3005
R16452 gnd.n3035 gnd.n3033 9.3005
R16453 gnd.n3034 gnd.n2766 9.3005
R16454 gnd.n3053 gnd.n2765 9.3005
R16455 gnd.n3056 gnd.n3055 9.3005
R16456 gnd.n2759 gnd.n2758 9.3005
R16457 gnd.n3067 gnd.n3065 9.3005
R16458 gnd.n3066 gnd.n2740 9.3005
R16459 gnd.n3084 gnd.n2739 9.3005
R16460 gnd.n3087 gnd.n3086 9.3005
R16461 gnd.n2734 gnd.n2729 9.3005
R16462 gnd.n3097 gnd.n3096 9.3005
R16463 gnd.n2732 gnd.n2712 9.3005
R16464 gnd.n3118 gnd.n2713 9.3005
R16465 gnd.n3117 gnd.n3116 9.3005
R16466 gnd.n2715 gnd.n2691 9.3005
R16467 gnd.n3149 gnd.n3148 9.3005
R16468 gnd.n3151 gnd.n2636 9.3005
R16469 gnd.n3198 gnd.n2637 9.3005
R16470 gnd.n3197 gnd.n2638 9.3005
R16471 gnd.n3196 gnd.n2639 9.3005
R16472 gnd.n3162 gnd.n2640 9.3005
R16473 gnd.n3164 gnd.n2658 9.3005
R16474 gnd.n3184 gnd.n2659 9.3005
R16475 gnd.n3183 gnd.n2660 9.3005
R16476 gnd.n3182 gnd.n2661 9.3005
R16477 gnd.n3173 gnd.n2662 9.3005
R16478 gnd.n3174 gnd.n2549 9.3005
R16479 gnd.n3240 gnd.n3239 9.3005
R16480 gnd.n3241 gnd.n2542 9.3005
R16481 gnd.n3251 gnd.n3250 9.3005
R16482 gnd.n3253 gnd.n2538 9.3005
R16483 gnd.n3263 gnd.n2539 9.3005
R16484 gnd.n3262 gnd.n3261 9.3005
R16485 gnd.n3259 gnd.n2517 9.3005
R16486 gnd.n3285 gnd.n2518 9.3005
R16487 gnd.n3284 gnd.n3283 9.3005
R16488 gnd.n2520 gnd.n2494 9.3005
R16489 gnd.n3325 gnd.n3324 9.3005
R16490 gnd.n3326 gnd.n2487 9.3005
R16491 gnd.n3336 gnd.n3335 9.3005
R16492 gnd.n3338 gnd.n2483 9.3005
R16493 gnd.n3348 gnd.n2484 9.3005
R16494 gnd.n3347 gnd.n3346 9.3005
R16495 gnd.n3344 gnd.n2462 9.3005
R16496 gnd.n3370 gnd.n2463 9.3005
R16497 gnd.n3369 gnd.n3368 9.3005
R16498 gnd.n2465 gnd.n2440 9.3005
R16499 gnd.n3414 gnd.n3413 9.3005
R16500 gnd.n3415 gnd.n2433 9.3005
R16501 gnd.n3425 gnd.n3424 9.3005
R16502 gnd.n3683 gnd.n2429 9.3005
R16503 gnd.n3691 gnd.n2430 9.3005
R16504 gnd.n3690 gnd.n3689 9.3005
R16505 gnd.n2411 gnd.n2410 9.3005
R16506 gnd.n3714 gnd.n3713 9.3005
R16507 gnd.n2857 gnd.n2856 9.3005
R16508 gnd.n6719 gnd.n6718 9.3005
R16509 gnd.n795 gnd.n794 9.3005
R16510 gnd.n6726 gnd.n6725 9.3005
R16511 gnd.n6727 gnd.n793 9.3005
R16512 gnd.n6729 gnd.n6728 9.3005
R16513 gnd.n789 gnd.n788 9.3005
R16514 gnd.n6736 gnd.n6735 9.3005
R16515 gnd.n6737 gnd.n787 9.3005
R16516 gnd.n6739 gnd.n6738 9.3005
R16517 gnd.n783 gnd.n782 9.3005
R16518 gnd.n6746 gnd.n6745 9.3005
R16519 gnd.n6747 gnd.n781 9.3005
R16520 gnd.n6749 gnd.n6748 9.3005
R16521 gnd.n777 gnd.n776 9.3005
R16522 gnd.n6756 gnd.n6755 9.3005
R16523 gnd.n6757 gnd.n775 9.3005
R16524 gnd.n6759 gnd.n6758 9.3005
R16525 gnd.n771 gnd.n770 9.3005
R16526 gnd.n6766 gnd.n6765 9.3005
R16527 gnd.n6767 gnd.n769 9.3005
R16528 gnd.n6769 gnd.n6768 9.3005
R16529 gnd.n765 gnd.n764 9.3005
R16530 gnd.n6776 gnd.n6775 9.3005
R16531 gnd.n6777 gnd.n763 9.3005
R16532 gnd.n6779 gnd.n6778 9.3005
R16533 gnd.n759 gnd.n758 9.3005
R16534 gnd.n6786 gnd.n6785 9.3005
R16535 gnd.n6787 gnd.n757 9.3005
R16536 gnd.n6789 gnd.n6788 9.3005
R16537 gnd.n753 gnd.n752 9.3005
R16538 gnd.n6796 gnd.n6795 9.3005
R16539 gnd.n6797 gnd.n751 9.3005
R16540 gnd.n6799 gnd.n6798 9.3005
R16541 gnd.n747 gnd.n746 9.3005
R16542 gnd.n6806 gnd.n6805 9.3005
R16543 gnd.n6807 gnd.n745 9.3005
R16544 gnd.n6809 gnd.n6808 9.3005
R16545 gnd.n741 gnd.n740 9.3005
R16546 gnd.n6816 gnd.n6815 9.3005
R16547 gnd.n6817 gnd.n739 9.3005
R16548 gnd.n6819 gnd.n6818 9.3005
R16549 gnd.n735 gnd.n734 9.3005
R16550 gnd.n6826 gnd.n6825 9.3005
R16551 gnd.n6827 gnd.n733 9.3005
R16552 gnd.n6829 gnd.n6828 9.3005
R16553 gnd.n729 gnd.n728 9.3005
R16554 gnd.n6836 gnd.n6835 9.3005
R16555 gnd.n6837 gnd.n727 9.3005
R16556 gnd.n6839 gnd.n6838 9.3005
R16557 gnd.n723 gnd.n722 9.3005
R16558 gnd.n6846 gnd.n6845 9.3005
R16559 gnd.n6847 gnd.n721 9.3005
R16560 gnd.n6849 gnd.n6848 9.3005
R16561 gnd.n717 gnd.n716 9.3005
R16562 gnd.n6856 gnd.n6855 9.3005
R16563 gnd.n6857 gnd.n715 9.3005
R16564 gnd.n6859 gnd.n6858 9.3005
R16565 gnd.n711 gnd.n710 9.3005
R16566 gnd.n6866 gnd.n6865 9.3005
R16567 gnd.n6867 gnd.n709 9.3005
R16568 gnd.n6869 gnd.n6868 9.3005
R16569 gnd.n705 gnd.n704 9.3005
R16570 gnd.n6876 gnd.n6875 9.3005
R16571 gnd.n6877 gnd.n703 9.3005
R16572 gnd.n6879 gnd.n6878 9.3005
R16573 gnd.n699 gnd.n698 9.3005
R16574 gnd.n6886 gnd.n6885 9.3005
R16575 gnd.n6887 gnd.n697 9.3005
R16576 gnd.n6889 gnd.n6888 9.3005
R16577 gnd.n693 gnd.n692 9.3005
R16578 gnd.n6896 gnd.n6895 9.3005
R16579 gnd.n6897 gnd.n691 9.3005
R16580 gnd.n6899 gnd.n6898 9.3005
R16581 gnd.n687 gnd.n686 9.3005
R16582 gnd.n6906 gnd.n6905 9.3005
R16583 gnd.n6907 gnd.n685 9.3005
R16584 gnd.n6909 gnd.n6908 9.3005
R16585 gnd.n681 gnd.n680 9.3005
R16586 gnd.n6916 gnd.n6915 9.3005
R16587 gnd.n6917 gnd.n679 9.3005
R16588 gnd.n6919 gnd.n6918 9.3005
R16589 gnd.n675 gnd.n674 9.3005
R16590 gnd.n6926 gnd.n6925 9.3005
R16591 gnd.n6927 gnd.n673 9.3005
R16592 gnd.n6929 gnd.n6928 9.3005
R16593 gnd.n669 gnd.n668 9.3005
R16594 gnd.n6936 gnd.n6935 9.3005
R16595 gnd.n6937 gnd.n667 9.3005
R16596 gnd.n6939 gnd.n6938 9.3005
R16597 gnd.n663 gnd.n662 9.3005
R16598 gnd.n6946 gnd.n6945 9.3005
R16599 gnd.n6947 gnd.n661 9.3005
R16600 gnd.n6949 gnd.n6948 9.3005
R16601 gnd.n657 gnd.n656 9.3005
R16602 gnd.n6956 gnd.n6955 9.3005
R16603 gnd.n6957 gnd.n655 9.3005
R16604 gnd.n6959 gnd.n6958 9.3005
R16605 gnd.n651 gnd.n650 9.3005
R16606 gnd.n6966 gnd.n6965 9.3005
R16607 gnd.n6967 gnd.n649 9.3005
R16608 gnd.n6969 gnd.n6968 9.3005
R16609 gnd.n645 gnd.n644 9.3005
R16610 gnd.n6976 gnd.n6975 9.3005
R16611 gnd.n6977 gnd.n643 9.3005
R16612 gnd.n6979 gnd.n6978 9.3005
R16613 gnd.n639 gnd.n638 9.3005
R16614 gnd.n6986 gnd.n6985 9.3005
R16615 gnd.n6987 gnd.n637 9.3005
R16616 gnd.n6989 gnd.n6988 9.3005
R16617 gnd.n633 gnd.n632 9.3005
R16618 gnd.n6996 gnd.n6995 9.3005
R16619 gnd.n6997 gnd.n631 9.3005
R16620 gnd.n6999 gnd.n6998 9.3005
R16621 gnd.n627 gnd.n626 9.3005
R16622 gnd.n7006 gnd.n7005 9.3005
R16623 gnd.n7007 gnd.n625 9.3005
R16624 gnd.n7009 gnd.n7008 9.3005
R16625 gnd.n621 gnd.n620 9.3005
R16626 gnd.n7016 gnd.n7015 9.3005
R16627 gnd.n7017 gnd.n619 9.3005
R16628 gnd.n7019 gnd.n7018 9.3005
R16629 gnd.n615 gnd.n614 9.3005
R16630 gnd.n7026 gnd.n7025 9.3005
R16631 gnd.n7027 gnd.n613 9.3005
R16632 gnd.n7029 gnd.n7028 9.3005
R16633 gnd.n609 gnd.n608 9.3005
R16634 gnd.n7036 gnd.n7035 9.3005
R16635 gnd.n7037 gnd.n607 9.3005
R16636 gnd.n7039 gnd.n7038 9.3005
R16637 gnd.n603 gnd.n602 9.3005
R16638 gnd.n7046 gnd.n7045 9.3005
R16639 gnd.n7047 gnd.n601 9.3005
R16640 gnd.n7049 gnd.n7048 9.3005
R16641 gnd.n597 gnd.n596 9.3005
R16642 gnd.n7056 gnd.n7055 9.3005
R16643 gnd.n7057 gnd.n595 9.3005
R16644 gnd.n7059 gnd.n7058 9.3005
R16645 gnd.n591 gnd.n590 9.3005
R16646 gnd.n7066 gnd.n7065 9.3005
R16647 gnd.n7067 gnd.n589 9.3005
R16648 gnd.n7069 gnd.n7068 9.3005
R16649 gnd.n585 gnd.n584 9.3005
R16650 gnd.n7076 gnd.n7075 9.3005
R16651 gnd.n7077 gnd.n583 9.3005
R16652 gnd.n7079 gnd.n7078 9.3005
R16653 gnd.n579 gnd.n578 9.3005
R16654 gnd.n7086 gnd.n7085 9.3005
R16655 gnd.n7087 gnd.n577 9.3005
R16656 gnd.n7089 gnd.n7088 9.3005
R16657 gnd.n573 gnd.n572 9.3005
R16658 gnd.n7096 gnd.n7095 9.3005
R16659 gnd.n7097 gnd.n571 9.3005
R16660 gnd.n7099 gnd.n7098 9.3005
R16661 gnd.n567 gnd.n566 9.3005
R16662 gnd.n7106 gnd.n7105 9.3005
R16663 gnd.n7107 gnd.n565 9.3005
R16664 gnd.n7109 gnd.n7108 9.3005
R16665 gnd.n561 gnd.n560 9.3005
R16666 gnd.n7116 gnd.n7115 9.3005
R16667 gnd.n7117 gnd.n559 9.3005
R16668 gnd.n7119 gnd.n7118 9.3005
R16669 gnd.n555 gnd.n554 9.3005
R16670 gnd.n7126 gnd.n7125 9.3005
R16671 gnd.n7127 gnd.n553 9.3005
R16672 gnd.n7130 gnd.n7129 9.3005
R16673 gnd.n7128 gnd.n549 9.3005
R16674 gnd.n7136 gnd.n548 9.3005
R16675 gnd.n7138 gnd.n7137 9.3005
R16676 gnd.n544 gnd.n543 9.3005
R16677 gnd.n7147 gnd.n7146 9.3005
R16678 gnd.n7148 gnd.n542 9.3005
R16679 gnd.n7150 gnd.n7149 9.3005
R16680 gnd.n538 gnd.n537 9.3005
R16681 gnd.n7157 gnd.n7156 9.3005
R16682 gnd.n7158 gnd.n536 9.3005
R16683 gnd.n7160 gnd.n7159 9.3005
R16684 gnd.n532 gnd.n531 9.3005
R16685 gnd.n7167 gnd.n7166 9.3005
R16686 gnd.n7168 gnd.n530 9.3005
R16687 gnd.n7170 gnd.n7169 9.3005
R16688 gnd.n526 gnd.n525 9.3005
R16689 gnd.n7177 gnd.n7176 9.3005
R16690 gnd.n7178 gnd.n524 9.3005
R16691 gnd.n7180 gnd.n7179 9.3005
R16692 gnd.n520 gnd.n519 9.3005
R16693 gnd.n7187 gnd.n7186 9.3005
R16694 gnd.n7188 gnd.n518 9.3005
R16695 gnd.n7190 gnd.n7189 9.3005
R16696 gnd.n514 gnd.n513 9.3005
R16697 gnd.n7197 gnd.n7196 9.3005
R16698 gnd.n7198 gnd.n512 9.3005
R16699 gnd.n7200 gnd.n7199 9.3005
R16700 gnd.n508 gnd.n507 9.3005
R16701 gnd.n7207 gnd.n7206 9.3005
R16702 gnd.n7208 gnd.n506 9.3005
R16703 gnd.n7210 gnd.n7209 9.3005
R16704 gnd.n502 gnd.n501 9.3005
R16705 gnd.n7217 gnd.n7216 9.3005
R16706 gnd.n7218 gnd.n500 9.3005
R16707 gnd.n7220 gnd.n7219 9.3005
R16708 gnd.n496 gnd.n495 9.3005
R16709 gnd.n7227 gnd.n7226 9.3005
R16710 gnd.n7228 gnd.n494 9.3005
R16711 gnd.n7230 gnd.n7229 9.3005
R16712 gnd.n490 gnd.n489 9.3005
R16713 gnd.n7237 gnd.n7236 9.3005
R16714 gnd.n7238 gnd.n488 9.3005
R16715 gnd.n7240 gnd.n7239 9.3005
R16716 gnd.n484 gnd.n483 9.3005
R16717 gnd.n7247 gnd.n7246 9.3005
R16718 gnd.n7248 gnd.n482 9.3005
R16719 gnd.n7250 gnd.n7249 9.3005
R16720 gnd.n478 gnd.n477 9.3005
R16721 gnd.n7257 gnd.n7256 9.3005
R16722 gnd.n7258 gnd.n476 9.3005
R16723 gnd.n7260 gnd.n7259 9.3005
R16724 gnd.n472 gnd.n471 9.3005
R16725 gnd.n7267 gnd.n7266 9.3005
R16726 gnd.n7268 gnd.n470 9.3005
R16727 gnd.n7270 gnd.n7269 9.3005
R16728 gnd.n466 gnd.n465 9.3005
R16729 gnd.n7277 gnd.n7276 9.3005
R16730 gnd.n7278 gnd.n464 9.3005
R16731 gnd.n7280 gnd.n7279 9.3005
R16732 gnd.n460 gnd.n459 9.3005
R16733 gnd.n7287 gnd.n7286 9.3005
R16734 gnd.n7288 gnd.n458 9.3005
R16735 gnd.n7290 gnd.n7289 9.3005
R16736 gnd.n454 gnd.n453 9.3005
R16737 gnd.n7297 gnd.n7296 9.3005
R16738 gnd.n7298 gnd.n452 9.3005
R16739 gnd.n7300 gnd.n7299 9.3005
R16740 gnd.n448 gnd.n447 9.3005
R16741 gnd.n7307 gnd.n7306 9.3005
R16742 gnd.n7308 gnd.n446 9.3005
R16743 gnd.n7310 gnd.n7309 9.3005
R16744 gnd.n442 gnd.n441 9.3005
R16745 gnd.n7317 gnd.n7316 9.3005
R16746 gnd.n7318 gnd.n440 9.3005
R16747 gnd.n7320 gnd.n7319 9.3005
R16748 gnd.n436 gnd.n435 9.3005
R16749 gnd.n7327 gnd.n7326 9.3005
R16750 gnd.n7328 gnd.n434 9.3005
R16751 gnd.n7330 gnd.n7329 9.3005
R16752 gnd.n430 gnd.n429 9.3005
R16753 gnd.n7337 gnd.n7336 9.3005
R16754 gnd.n7338 gnd.n428 9.3005
R16755 gnd.n7340 gnd.n7339 9.3005
R16756 gnd.n424 gnd.n423 9.3005
R16757 gnd.n7348 gnd.n7347 9.3005
R16758 gnd.n7349 gnd.n422 9.3005
R16759 gnd.n7351 gnd.n7350 9.3005
R16760 gnd.n7140 gnd.n7139 9.3005
R16761 gnd.n7798 gnd.n134 9.3005
R16762 gnd.n7797 gnd.n136 9.3005
R16763 gnd.n140 gnd.n137 9.3005
R16764 gnd.n7792 gnd.n141 9.3005
R16765 gnd.n7791 gnd.n142 9.3005
R16766 gnd.n7790 gnd.n143 9.3005
R16767 gnd.n147 gnd.n144 9.3005
R16768 gnd.n7785 gnd.n148 9.3005
R16769 gnd.n7784 gnd.n149 9.3005
R16770 gnd.n7783 gnd.n150 9.3005
R16771 gnd.n154 gnd.n151 9.3005
R16772 gnd.n7778 gnd.n155 9.3005
R16773 gnd.n7777 gnd.n156 9.3005
R16774 gnd.n7776 gnd.n157 9.3005
R16775 gnd.n161 gnd.n158 9.3005
R16776 gnd.n7771 gnd.n162 9.3005
R16777 gnd.n7770 gnd.n163 9.3005
R16778 gnd.n7766 gnd.n164 9.3005
R16779 gnd.n168 gnd.n165 9.3005
R16780 gnd.n7761 gnd.n169 9.3005
R16781 gnd.n7760 gnd.n170 9.3005
R16782 gnd.n7759 gnd.n171 9.3005
R16783 gnd.n175 gnd.n172 9.3005
R16784 gnd.n7754 gnd.n176 9.3005
R16785 gnd.n7753 gnd.n177 9.3005
R16786 gnd.n7752 gnd.n178 9.3005
R16787 gnd.n182 gnd.n179 9.3005
R16788 gnd.n7747 gnd.n183 9.3005
R16789 gnd.n7746 gnd.n184 9.3005
R16790 gnd.n7745 gnd.n185 9.3005
R16791 gnd.n189 gnd.n186 9.3005
R16792 gnd.n7740 gnd.n190 9.3005
R16793 gnd.n7739 gnd.n191 9.3005
R16794 gnd.n7738 gnd.n192 9.3005
R16795 gnd.n196 gnd.n193 9.3005
R16796 gnd.n7733 gnd.n197 9.3005
R16797 gnd.n7732 gnd.n7731 9.3005
R16798 gnd.n7730 gnd.n200 9.3005
R16799 gnd.n7800 gnd.n7799 9.3005
R16800 gnd.n1456 gnd.n1455 9.3005
R16801 gnd.n1457 gnd.n1454 9.3005
R16802 gnd.n1473 gnd.n1458 9.3005
R16803 gnd.n1472 gnd.n1459 9.3005
R16804 gnd.n1471 gnd.n1460 9.3005
R16805 gnd.n1469 gnd.n1461 9.3005
R16806 gnd.n1468 gnd.n1462 9.3005
R16807 gnd.n1466 gnd.n1463 9.3005
R16808 gnd.n1465 gnd.n1464 9.3005
R16809 gnd.n1391 gnd.n1390 9.3005
R16810 gnd.n6124 gnd.n6123 9.3005
R16811 gnd.n6125 gnd.n1389 9.3005
R16812 gnd.n6127 gnd.n6126 9.3005
R16813 gnd.n6128 gnd.n1388 9.3005
R16814 gnd.n6131 gnd.n6130 9.3005
R16815 gnd.n6132 gnd.n1387 9.3005
R16816 gnd.n6136 gnd.n6133 9.3005
R16817 gnd.n6135 gnd.n6134 9.3005
R16818 gnd.n388 gnd.n387 9.3005
R16819 gnd.n7387 gnd.n7386 9.3005
R16820 gnd.n7388 gnd.n386 9.3005
R16821 gnd.n7396 gnd.n7389 9.3005
R16822 gnd.n7395 gnd.n7390 9.3005
R16823 gnd.n7394 gnd.n7391 9.3005
R16824 gnd.n354 gnd.n353 9.3005
R16825 gnd.n7432 gnd.n7431 9.3005
R16826 gnd.n7433 gnd.n352 9.3005
R16827 gnd.n7442 gnd.n7434 9.3005
R16828 gnd.n7441 gnd.n7435 9.3005
R16829 gnd.n7440 gnd.n7436 9.3005
R16830 gnd.n7438 gnd.n7437 9.3005
R16831 gnd.n338 gnd.n337 9.3005
R16832 gnd.n7462 gnd.n7461 9.3005
R16833 gnd.n7463 gnd.n336 9.3005
R16834 gnd.n7530 gnd.n7464 9.3005
R16835 gnd.n7529 gnd.n7465 9.3005
R16836 gnd.n7528 gnd.n7466 9.3005
R16837 gnd.n7526 gnd.n7467 9.3005
R16838 gnd.n7525 gnd.n7468 9.3005
R16839 gnd.n7523 gnd.n7469 9.3005
R16840 gnd.n7522 gnd.n7470 9.3005
R16841 gnd.n7520 gnd.n7471 9.3005
R16842 gnd.n7519 gnd.n7472 9.3005
R16843 gnd.n7517 gnd.n7473 9.3005
R16844 gnd.n7516 gnd.n7474 9.3005
R16845 gnd.n7514 gnd.n7475 9.3005
R16846 gnd.n7513 gnd.n7476 9.3005
R16847 gnd.n7511 gnd.n7477 9.3005
R16848 gnd.n7510 gnd.n7478 9.3005
R16849 gnd.n7508 gnd.n7479 9.3005
R16850 gnd.n7507 gnd.n7480 9.3005
R16851 gnd.n7505 gnd.n7481 9.3005
R16852 gnd.n7504 gnd.n7482 9.3005
R16853 gnd.n7502 gnd.n7483 9.3005
R16854 gnd.n7501 gnd.n7484 9.3005
R16855 gnd.n7499 gnd.n7485 9.3005
R16856 gnd.n7498 gnd.n7486 9.3005
R16857 gnd.n7496 gnd.n7487 9.3005
R16858 gnd.n7495 gnd.n7488 9.3005
R16859 gnd.n7493 gnd.n7489 9.3005
R16860 gnd.n7492 gnd.n7491 9.3005
R16861 gnd.n7490 gnd.n204 9.3005
R16862 gnd.n7727 gnd.n203 9.3005
R16863 gnd.n7729 gnd.n7728 9.3005
R16864 gnd.n1335 gnd.n1333 9.3005
R16865 gnd.n6225 gnd.n6224 9.3005
R16866 gnd.n6226 gnd.n1327 9.3005
R16867 gnd.n6229 gnd.n1326 9.3005
R16868 gnd.n6230 gnd.n1325 9.3005
R16869 gnd.n6233 gnd.n1324 9.3005
R16870 gnd.n6234 gnd.n1323 9.3005
R16871 gnd.n6237 gnd.n1322 9.3005
R16872 gnd.n6238 gnd.n1321 9.3005
R16873 gnd.n6241 gnd.n1320 9.3005
R16874 gnd.n6242 gnd.n1319 9.3005
R16875 gnd.n6245 gnd.n1318 9.3005
R16876 gnd.n6246 gnd.n1317 9.3005
R16877 gnd.n6249 gnd.n1316 9.3005
R16878 gnd.n6250 gnd.n1315 9.3005
R16879 gnd.n6253 gnd.n1314 9.3005
R16880 gnd.n6254 gnd.n1313 9.3005
R16881 gnd.n6257 gnd.n1312 9.3005
R16882 gnd.n6258 gnd.n1311 9.3005
R16883 gnd.n6261 gnd.n1310 9.3005
R16884 gnd.n6263 gnd.n1304 9.3005
R16885 gnd.n6266 gnd.n1303 9.3005
R16886 gnd.n6267 gnd.n1302 9.3005
R16887 gnd.n6270 gnd.n1301 9.3005
R16888 gnd.n6271 gnd.n1300 9.3005
R16889 gnd.n6274 gnd.n1299 9.3005
R16890 gnd.n6275 gnd.n1298 9.3005
R16891 gnd.n6278 gnd.n1297 9.3005
R16892 gnd.n6279 gnd.n1296 9.3005
R16893 gnd.n6282 gnd.n1295 9.3005
R16894 gnd.n6283 gnd.n1294 9.3005
R16895 gnd.n6286 gnd.n1293 9.3005
R16896 gnd.n6288 gnd.n1292 9.3005
R16897 gnd.n6289 gnd.n1291 9.3005
R16898 gnd.n6290 gnd.n1290 9.3005
R16899 gnd.n6291 gnd.n1289 9.3005
R16900 gnd.n6223 gnd.n1332 9.3005
R16901 gnd.n6222 gnd.n6221 9.3005
R16902 gnd.n6051 gnd.n6048 9.3005
R16903 gnd.n6050 gnd.n6049 9.3005
R16904 gnd.n1429 gnd.n1428 9.3005
R16905 gnd.n6077 gnd.n6076 9.3005
R16906 gnd.n6078 gnd.n1427 9.3005
R16907 gnd.n6082 gnd.n6079 9.3005
R16908 gnd.n6081 gnd.n6080 9.3005
R16909 gnd.n1402 gnd.n1401 9.3005
R16910 gnd.n6114 gnd.n6113 9.3005
R16911 gnd.n6115 gnd.n1400 9.3005
R16912 gnd.n6119 gnd.n6116 9.3005
R16913 gnd.n6118 gnd.n6117 9.3005
R16914 gnd.n1368 gnd.n1367 9.3005
R16915 gnd.n6184 gnd.n6183 9.3005
R16916 gnd.n6185 gnd.n1366 9.3005
R16917 gnd.n6187 gnd.n6186 9.3005
R16918 gnd.n397 gnd.n396 9.3005
R16919 gnd.n7377 gnd.n7376 9.3005
R16920 gnd.n7378 gnd.n395 9.3005
R16921 gnd.n7382 gnd.n7379 9.3005
R16922 gnd.n7381 gnd.n7380 9.3005
R16923 gnd.n364 gnd.n363 9.3005
R16924 gnd.n7423 gnd.n7422 9.3005
R16925 gnd.n7424 gnd.n362 9.3005
R16926 gnd.n7426 gnd.n7425 9.3005
R16927 gnd.n7427 gnd.n303 9.3005
R16928 gnd.n7558 gnd.n7557 9.3005
R16929 gnd.n288 gnd.n287 9.3005
R16930 gnd.n7571 gnd.n7570 9.3005
R16931 gnd.n7572 gnd.n286 9.3005
R16932 gnd.n7574 gnd.n7573 9.3005
R16933 gnd.n274 gnd.n273 9.3005
R16934 gnd.n7587 gnd.n7586 9.3005
R16935 gnd.n7588 gnd.n272 9.3005
R16936 gnd.n7590 gnd.n7589 9.3005
R16937 gnd.n258 gnd.n257 9.3005
R16938 gnd.n7603 gnd.n7602 9.3005
R16939 gnd.n7604 gnd.n256 9.3005
R16940 gnd.n7606 gnd.n7605 9.3005
R16941 gnd.n243 gnd.n242 9.3005
R16942 gnd.n7619 gnd.n7618 9.3005
R16943 gnd.n7620 gnd.n241 9.3005
R16944 gnd.n7622 gnd.n7621 9.3005
R16945 gnd.n227 gnd.n226 9.3005
R16946 gnd.n7635 gnd.n7634 9.3005
R16947 gnd.n7636 gnd.n225 9.3005
R16948 gnd.n7638 gnd.n7637 9.3005
R16949 gnd.n211 gnd.n210 9.3005
R16950 gnd.n7719 gnd.n7718 9.3005
R16951 gnd.n7720 gnd.n209 9.3005
R16952 gnd.n7722 gnd.n7721 9.3005
R16953 gnd.n133 gnd.n132 9.3005
R16954 gnd.n7802 gnd.n7801 9.3005
R16955 gnd.n6047 gnd.n6046 9.3005
R16956 gnd.n7556 gnd.n302 9.3005
R16957 gnd.n968 gnd.n967 9.3005
R16958 gnd.n4371 gnd.n4370 9.3005
R16959 gnd.n4372 gnd.n4368 9.3005
R16960 gnd.n4374 gnd.n4373 9.3005
R16961 gnd.n2165 gnd.n2164 9.3005
R16962 gnd.n4412 gnd.n4411 9.3005
R16963 gnd.n4413 gnd.n2163 9.3005
R16964 gnd.n4415 gnd.n4414 9.3005
R16965 gnd.n2161 gnd.n2160 9.3005
R16966 gnd.n4420 gnd.n4419 9.3005
R16967 gnd.n4421 gnd.n2159 9.3005
R16968 gnd.n4423 gnd.n4422 9.3005
R16969 gnd.n2144 gnd.n2143 9.3005
R16970 gnd.n4461 gnd.n4460 9.3005
R16971 gnd.n4462 gnd.n2142 9.3005
R16972 gnd.n4464 gnd.n4463 9.3005
R16973 gnd.n2140 gnd.n2139 9.3005
R16974 gnd.n4469 gnd.n4468 9.3005
R16975 gnd.n4470 gnd.n2138 9.3005
R16976 gnd.n4508 gnd.n4471 9.3005
R16977 gnd.n4507 gnd.n4472 9.3005
R16978 gnd.n4506 gnd.n4473 9.3005
R16979 gnd.n4476 gnd.n4474 9.3005
R16980 gnd.n4502 gnd.n4477 9.3005
R16981 gnd.n4501 gnd.n4478 9.3005
R16982 gnd.n4500 gnd.n4479 9.3005
R16983 gnd.n4482 gnd.n4480 9.3005
R16984 gnd.n4496 gnd.n4483 9.3005
R16985 gnd.n4495 gnd.n4484 9.3005
R16986 gnd.n4494 gnd.n4485 9.3005
R16987 gnd.n4487 gnd.n4486 9.3005
R16988 gnd.n4489 gnd.n4488 9.3005
R16989 gnd.n1965 gnd.n1964 9.3005
R16990 gnd.n5618 gnd.n5617 9.3005
R16991 gnd.n5619 gnd.n1963 9.3005
R16992 gnd.n5621 gnd.n5620 9.3005
R16993 gnd.n1951 gnd.n1950 9.3005
R16994 gnd.n5634 gnd.n5633 9.3005
R16995 gnd.n5635 gnd.n1949 9.3005
R16996 gnd.n5637 gnd.n5636 9.3005
R16997 gnd.n1939 gnd.n1938 9.3005
R16998 gnd.n5650 gnd.n5649 9.3005
R16999 gnd.n5651 gnd.n1937 9.3005
R17000 gnd.n5653 gnd.n5652 9.3005
R17001 gnd.n1926 gnd.n1925 9.3005
R17002 gnd.n5666 gnd.n5665 9.3005
R17003 gnd.n5667 gnd.n1924 9.3005
R17004 gnd.n5669 gnd.n5668 9.3005
R17005 gnd.n1911 gnd.n1910 9.3005
R17006 gnd.n5682 gnd.n5681 9.3005
R17007 gnd.n5683 gnd.n1909 9.3005
R17008 gnd.n5685 gnd.n5684 9.3005
R17009 gnd.n1897 gnd.n1896 9.3005
R17010 gnd.n5698 gnd.n5697 9.3005
R17011 gnd.n5699 gnd.n1895 9.3005
R17012 gnd.n5701 gnd.n5700 9.3005
R17013 gnd.n1883 gnd.n1882 9.3005
R17014 gnd.n5714 gnd.n5713 9.3005
R17015 gnd.n5715 gnd.n1881 9.3005
R17016 gnd.n5717 gnd.n5716 9.3005
R17017 gnd.n1868 gnd.n1867 9.3005
R17018 gnd.n5730 gnd.n5729 9.3005
R17019 gnd.n5731 gnd.n1866 9.3005
R17020 gnd.n5733 gnd.n5732 9.3005
R17021 gnd.n1855 gnd.n1854 9.3005
R17022 gnd.n5746 gnd.n5745 9.3005
R17023 gnd.n5747 gnd.n1853 9.3005
R17024 gnd.n5749 gnd.n5748 9.3005
R17025 gnd.n1840 gnd.n1839 9.3005
R17026 gnd.n5762 gnd.n5761 9.3005
R17027 gnd.n5763 gnd.n1838 9.3005
R17028 gnd.n5765 gnd.n5764 9.3005
R17029 gnd.n1825 gnd.n1824 9.3005
R17030 gnd.n5778 gnd.n5777 9.3005
R17031 gnd.n5779 gnd.n1823 9.3005
R17032 gnd.n5781 gnd.n5780 9.3005
R17033 gnd.n1810 gnd.n1809 9.3005
R17034 gnd.n5794 gnd.n5793 9.3005
R17035 gnd.n5795 gnd.n1808 9.3005
R17036 gnd.n5797 gnd.n5796 9.3005
R17037 gnd.n1795 gnd.n1794 9.3005
R17038 gnd.n5810 gnd.n5809 9.3005
R17039 gnd.n5811 gnd.n1793 9.3005
R17040 gnd.n5813 gnd.n5812 9.3005
R17041 gnd.n1781 gnd.n1780 9.3005
R17042 gnd.n5826 gnd.n5825 9.3005
R17043 gnd.n5827 gnd.n1779 9.3005
R17044 gnd.n5829 gnd.n5828 9.3005
R17045 gnd.n1766 gnd.n1765 9.3005
R17046 gnd.n5842 gnd.n5841 9.3005
R17047 gnd.n5843 gnd.n1764 9.3005
R17048 gnd.n5845 gnd.n5844 9.3005
R17049 gnd.n1751 gnd.n1750 9.3005
R17050 gnd.n5858 gnd.n5857 9.3005
R17051 gnd.n5859 gnd.n1749 9.3005
R17052 gnd.n5861 gnd.n5860 9.3005
R17053 gnd.n1737 gnd.n1736 9.3005
R17054 gnd.n5874 gnd.n5873 9.3005
R17055 gnd.n5875 gnd.n1735 9.3005
R17056 gnd.n5877 gnd.n5876 9.3005
R17057 gnd.n1722 gnd.n1721 9.3005
R17058 gnd.n5890 gnd.n5889 9.3005
R17059 gnd.n5891 gnd.n1720 9.3005
R17060 gnd.n5893 gnd.n5892 9.3005
R17061 gnd.n1708 gnd.n1707 9.3005
R17062 gnd.n5906 gnd.n5905 9.3005
R17063 gnd.n5907 gnd.n1706 9.3005
R17064 gnd.n5909 gnd.n5908 9.3005
R17065 gnd.n1692 gnd.n1691 9.3005
R17066 gnd.n5922 gnd.n5921 9.3005
R17067 gnd.n5923 gnd.n1690 9.3005
R17068 gnd.n5925 gnd.n5924 9.3005
R17069 gnd.n1678 gnd.n1677 9.3005
R17070 gnd.n5938 gnd.n5937 9.3005
R17071 gnd.n5939 gnd.n1676 9.3005
R17072 gnd.n5941 gnd.n5940 9.3005
R17073 gnd.n1666 gnd.n1665 9.3005
R17074 gnd.n5954 gnd.n5953 9.3005
R17075 gnd.n5955 gnd.n1664 9.3005
R17076 gnd.n5957 gnd.n5956 9.3005
R17077 gnd.n1651 gnd.n1650 9.3005
R17078 gnd.n5970 gnd.n5969 9.3005
R17079 gnd.n5971 gnd.n1649 9.3005
R17080 gnd.n5973 gnd.n5972 9.3005
R17081 gnd.n1637 gnd.n1636 9.3005
R17082 gnd.n5986 gnd.n5985 9.3005
R17083 gnd.n5987 gnd.n1635 9.3005
R17084 gnd.n5989 gnd.n5988 9.3005
R17085 gnd.n1624 gnd.n1623 9.3005
R17086 gnd.n6004 gnd.n6003 9.3005
R17087 gnd.n6005 gnd.n1622 9.3005
R17088 gnd.n6010 gnd.n6006 9.3005
R17089 gnd.n6009 gnd.n6008 9.3005
R17090 gnd.n6007 gnd.n1250 9.3005
R17091 gnd.n6300 gnd.n1251 9.3005
R17092 gnd.n6299 gnd.n1252 9.3005
R17093 gnd.n6298 gnd.n1253 9.3005
R17094 gnd.n1443 gnd.n1254 9.3005
R17095 gnd.n1446 gnd.n1445 9.3005
R17096 gnd.n1447 gnd.n1442 9.3005
R17097 gnd.n1449 gnd.n1448 9.3005
R17098 gnd.n1440 gnd.n1439 9.3005
R17099 gnd.n6066 gnd.n6065 9.3005
R17100 gnd.n6067 gnd.n1438 9.3005
R17101 gnd.n6071 gnd.n6068 9.3005
R17102 gnd.n6070 gnd.n6069 9.3005
R17103 gnd.n1412 gnd.n1411 9.3005
R17104 gnd.n6102 gnd.n6101 9.3005
R17105 gnd.n6103 gnd.n1410 9.3005
R17106 gnd.n6107 gnd.n6104 9.3005
R17107 gnd.n6106 gnd.n6105 9.3005
R17108 gnd.n1378 gnd.n1377 9.3005
R17109 gnd.n6163 gnd.n6162 9.3005
R17110 gnd.n6164 gnd.n1376 9.3005
R17111 gnd.n6178 gnd.n6165 9.3005
R17112 gnd.n6177 gnd.n6166 9.3005
R17113 gnd.n6176 gnd.n6167 9.3005
R17114 gnd.n6169 gnd.n6168 9.3005
R17115 gnd.n6172 gnd.n6171 9.3005
R17116 gnd.n6170 gnd.n411 9.3005
R17117 gnd.n7362 gnd.n412 9.3005
R17118 gnd.n7361 gnd.n413 9.3005
R17119 gnd.n7360 gnd.n414 9.3005
R17120 gnd.n417 gnd.n415 9.3005
R17121 gnd.n7356 gnd.n418 9.3005
R17122 gnd.n7355 gnd.n419 9.3005
R17123 gnd.n7354 gnd.n420 9.3005
R17124 gnd.n6545 gnd.n6544 9.3005
R17125 gnd.n3924 gnd.n3923 9.3005
R17126 gnd.n3970 gnd.n3879 9.3005
R17127 gnd.n3969 gnd.n3880 9.3005
R17128 gnd.n3968 gnd.n3881 9.3005
R17129 gnd.n3966 gnd.n3882 9.3005
R17130 gnd.n3965 gnd.n3883 9.3005
R17131 gnd.n3963 gnd.n3884 9.3005
R17132 gnd.n3962 gnd.n3885 9.3005
R17133 gnd.n3960 gnd.n3886 9.3005
R17134 gnd.n3959 gnd.n3887 9.3005
R17135 gnd.n3957 gnd.n3888 9.3005
R17136 gnd.n3956 gnd.n3889 9.3005
R17137 gnd.n3954 gnd.n3890 9.3005
R17138 gnd.n3953 gnd.n3891 9.3005
R17139 gnd.n3951 gnd.n3892 9.3005
R17140 gnd.n3950 gnd.n3893 9.3005
R17141 gnd.n3948 gnd.n3894 9.3005
R17142 gnd.n3947 gnd.n3895 9.3005
R17143 gnd.n3945 gnd.n3896 9.3005
R17144 gnd.n3944 gnd.n3897 9.3005
R17145 gnd.n3942 gnd.n3898 9.3005
R17146 gnd.n3941 gnd.n3899 9.3005
R17147 gnd.n3939 gnd.n3900 9.3005
R17148 gnd.n3938 gnd.n3901 9.3005
R17149 gnd.n3936 gnd.n3902 9.3005
R17150 gnd.n3935 gnd.n3903 9.3005
R17151 gnd.n3933 gnd.n3904 9.3005
R17152 gnd.n3932 gnd.n3905 9.3005
R17153 gnd.n3930 gnd.n3906 9.3005
R17154 gnd.n3929 gnd.n3907 9.3005
R17155 gnd.n3927 gnd.n3908 9.3005
R17156 gnd.n3926 gnd.n3909 9.3005
R17157 gnd.n3878 gnd.n3811 9.3005
R17158 gnd.n3871 gnd.n3870 9.3005
R17159 gnd.n3869 gnd.n3817 9.3005
R17160 gnd.n3868 gnd.n3867 9.3005
R17161 gnd.n3819 gnd.n3818 9.3005
R17162 gnd.n3861 gnd.n3860 9.3005
R17163 gnd.n3859 gnd.n3821 9.3005
R17164 gnd.n3858 gnd.n3857 9.3005
R17165 gnd.n3823 gnd.n3822 9.3005
R17166 gnd.n3851 gnd.n3850 9.3005
R17167 gnd.n3849 gnd.n3825 9.3005
R17168 gnd.n3848 gnd.n3847 9.3005
R17169 gnd.n3827 gnd.n3826 9.3005
R17170 gnd.n3841 gnd.n3840 9.3005
R17171 gnd.n3839 gnd.n3829 9.3005
R17172 gnd.n3838 gnd.n3837 9.3005
R17173 gnd.n3832 gnd.n3830 9.3005
R17174 gnd.n3831 gnd.n2332 9.3005
R17175 gnd.n3815 gnd.n3812 9.3005
R17176 gnd.n3877 gnd.n3876 9.3005
R17177 gnd.n4198 gnd.n2331 9.3005
R17178 gnd.n4200 gnd.n4199 9.3005
R17179 gnd.n2318 gnd.n2317 9.3005
R17180 gnd.n4213 gnd.n4212 9.3005
R17181 gnd.n4214 gnd.n2316 9.3005
R17182 gnd.n4216 gnd.n4215 9.3005
R17183 gnd.n2301 gnd.n2300 9.3005
R17184 gnd.n4229 gnd.n4228 9.3005
R17185 gnd.n4230 gnd.n2299 9.3005
R17186 gnd.n4232 gnd.n4231 9.3005
R17187 gnd.n2286 gnd.n2285 9.3005
R17188 gnd.n4245 gnd.n4244 9.3005
R17189 gnd.n4246 gnd.n2284 9.3005
R17190 gnd.n4248 gnd.n4247 9.3005
R17191 gnd.n2269 gnd.n2268 9.3005
R17192 gnd.n4261 gnd.n4260 9.3005
R17193 gnd.n4262 gnd.n2267 9.3005
R17194 gnd.n4264 gnd.n4263 9.3005
R17195 gnd.n2254 gnd.n2253 9.3005
R17196 gnd.n4277 gnd.n4276 9.3005
R17197 gnd.n4278 gnd.n2252 9.3005
R17198 gnd.n4280 gnd.n4279 9.3005
R17199 gnd.n2237 gnd.n2236 9.3005
R17200 gnd.n4294 gnd.n4293 9.3005
R17201 gnd.n4295 gnd.n2235 9.3005
R17202 gnd.n4297 gnd.n4296 9.3005
R17203 gnd.n2223 gnd.n2222 9.3005
R17204 gnd.n4310 gnd.n4309 9.3005
R17205 gnd.n4311 gnd.n2221 9.3005
R17206 gnd.n4314 gnd.n4312 9.3005
R17207 gnd.n4313 gnd.n2197 9.3005
R17208 gnd.n4328 gnd.n2198 9.3005
R17209 gnd.n4329 gnd.n2196 9.3005
R17210 gnd.n4341 gnd.n4330 9.3005
R17211 gnd.n4340 gnd.n4331 9.3005
R17212 gnd.n4339 gnd.n4332 9.3005
R17213 gnd.n4338 gnd.n4333 9.3005
R17214 gnd.n4336 gnd.n4335 9.3005
R17215 gnd.n4334 gnd.n989 9.3005
R17216 gnd.n6533 gnd.n990 9.3005
R17217 gnd.n6532 gnd.n991 9.3005
R17218 gnd.n6531 gnd.n992 9.3005
R17219 gnd.n1009 gnd.n993 9.3005
R17220 gnd.n6521 gnd.n1010 9.3005
R17221 gnd.n6520 gnd.n1011 9.3005
R17222 gnd.n6519 gnd.n1012 9.3005
R17223 gnd.n1031 gnd.n1013 9.3005
R17224 gnd.n6509 gnd.n1032 9.3005
R17225 gnd.n6508 gnd.n1033 9.3005
R17226 gnd.n6507 gnd.n1034 9.3005
R17227 gnd.n1051 gnd.n1035 9.3005
R17228 gnd.n6497 gnd.n1052 9.3005
R17229 gnd.n6496 gnd.n1053 9.3005
R17230 gnd.n6495 gnd.n1054 9.3005
R17231 gnd.n1073 gnd.n1055 9.3005
R17232 gnd.n6485 gnd.n1074 9.3005
R17233 gnd.n6484 gnd.n1075 9.3005
R17234 gnd.n6483 gnd.n1076 9.3005
R17235 gnd.n1094 gnd.n1077 9.3005
R17236 gnd.n6473 gnd.n1095 9.3005
R17237 gnd.n6472 gnd.n1096 9.3005
R17238 gnd.n6471 gnd.n1097 9.3005
R17239 gnd.n1114 gnd.n1098 9.3005
R17240 gnd.n6461 gnd.n6460 9.3005
R17241 gnd.n4197 gnd.n4196 9.3005
R17242 gnd.n5528 gnd.n2096 9.3005
R17243 gnd.n5531 gnd.n2095 9.3005
R17244 gnd.n5532 gnd.n2094 9.3005
R17245 gnd.n5535 gnd.n2093 9.3005
R17246 gnd.n5536 gnd.n2092 9.3005
R17247 gnd.n5539 gnd.n2091 9.3005
R17248 gnd.n5540 gnd.n2090 9.3005
R17249 gnd.n5543 gnd.n2089 9.3005
R17250 gnd.n5544 gnd.n2088 9.3005
R17251 gnd.n5547 gnd.n2087 9.3005
R17252 gnd.n5548 gnd.n2086 9.3005
R17253 gnd.n5551 gnd.n2085 9.3005
R17254 gnd.n5552 gnd.n2084 9.3005
R17255 gnd.n5553 gnd.n2083 9.3005
R17256 gnd.n2082 gnd.n2079 9.3005
R17257 gnd.n2081 gnd.n2080 9.3005
R17258 gnd.n4614 gnd.n4613 9.3005
R17259 gnd.n4610 gnd.n2101 9.3005
R17260 gnd.n4607 gnd.n2102 9.3005
R17261 gnd.n4606 gnd.n2103 9.3005
R17262 gnd.n4603 gnd.n2104 9.3005
R17263 gnd.n4602 gnd.n2105 9.3005
R17264 gnd.n4599 gnd.n2106 9.3005
R17265 gnd.n4598 gnd.n2107 9.3005
R17266 gnd.n4595 gnd.n2108 9.3005
R17267 gnd.n4594 gnd.n2109 9.3005
R17268 gnd.n4591 gnd.n2110 9.3005
R17269 gnd.n4590 gnd.n2111 9.3005
R17270 gnd.n4587 gnd.n2112 9.3005
R17271 gnd.n4586 gnd.n2113 9.3005
R17272 gnd.n4583 gnd.n2114 9.3005
R17273 gnd.n4582 gnd.n2115 9.3005
R17274 gnd.n4579 gnd.n2116 9.3005
R17275 gnd.n4578 gnd.n2117 9.3005
R17276 gnd.n4575 gnd.n4574 9.3005
R17277 gnd.n4573 gnd.n2119 9.3005
R17278 gnd.n4615 gnd.n2097 9.3005
R17279 gnd.n4109 gnd.n4035 9.3005
R17280 gnd.n4108 gnd.n4037 9.3005
R17281 gnd.n4107 gnd.n4038 9.3005
R17282 gnd.n4105 gnd.n4039 9.3005
R17283 gnd.n4104 gnd.n4040 9.3005
R17284 gnd.n4102 gnd.n4041 9.3005
R17285 gnd.n4101 gnd.n4042 9.3005
R17286 gnd.n4099 gnd.n4043 9.3005
R17287 gnd.n4098 gnd.n4044 9.3005
R17288 gnd.n4096 gnd.n4045 9.3005
R17289 gnd.n4095 gnd.n4046 9.3005
R17290 gnd.n4093 gnd.n4047 9.3005
R17291 gnd.n4092 gnd.n4048 9.3005
R17292 gnd.n4090 gnd.n4049 9.3005
R17293 gnd.n4089 gnd.n4050 9.3005
R17294 gnd.n4087 gnd.n4051 9.3005
R17295 gnd.n4086 gnd.n4052 9.3005
R17296 gnd.n4084 gnd.n4053 9.3005
R17297 gnd.n4083 gnd.n4054 9.3005
R17298 gnd.n4081 gnd.n4055 9.3005
R17299 gnd.n4080 gnd.n4056 9.3005
R17300 gnd.n4078 gnd.n4057 9.3005
R17301 gnd.n4077 gnd.n4058 9.3005
R17302 gnd.n4075 gnd.n4059 9.3005
R17303 gnd.n4074 gnd.n4060 9.3005
R17304 gnd.n4072 gnd.n4061 9.3005
R17305 gnd.n4071 gnd.n4062 9.3005
R17306 gnd.n4069 gnd.n4063 9.3005
R17307 gnd.n4068 gnd.n4064 9.3005
R17308 gnd.n4066 gnd.n4065 9.3005
R17309 gnd.n2201 gnd.n2199 9.3005
R17310 gnd.n4327 gnd.n4326 9.3005
R17311 gnd.n2206 gnd.n2200 9.3005
R17312 gnd.n2205 gnd.n2202 9.3005
R17313 gnd.n2204 gnd.n2203 9.3005
R17314 gnd.n2183 gnd.n2182 9.3005
R17315 gnd.n4354 gnd.n4353 9.3005
R17316 gnd.n4355 gnd.n2181 9.3005
R17317 gnd.n4357 gnd.n4356 9.3005
R17318 gnd.n2177 gnd.n2176 9.3005
R17319 gnd.n4380 gnd.n4379 9.3005
R17320 gnd.n4381 gnd.n2175 9.3005
R17321 gnd.n4383 gnd.n4382 9.3005
R17322 gnd.n4384 gnd.n2174 9.3005
R17323 gnd.n4388 gnd.n4387 9.3005
R17324 gnd.n4389 gnd.n2173 9.3005
R17325 gnd.n4391 gnd.n4390 9.3005
R17326 gnd.n2156 gnd.n2155 9.3005
R17327 gnd.n4429 gnd.n4428 9.3005
R17328 gnd.n4430 gnd.n2154 9.3005
R17329 gnd.n4432 gnd.n4431 9.3005
R17330 gnd.n4433 gnd.n2153 9.3005
R17331 gnd.n4437 gnd.n4436 9.3005
R17332 gnd.n4438 gnd.n2152 9.3005
R17333 gnd.n4444 gnd.n4439 9.3005
R17334 gnd.n4443 gnd.n4440 9.3005
R17335 gnd.n4442 gnd.n4441 9.3005
R17336 gnd.n2131 gnd.n2130 9.3005
R17337 gnd.n4522 gnd.n4521 9.3005
R17338 gnd.n4523 gnd.n2129 9.3005
R17339 gnd.n4526 gnd.n4525 9.3005
R17340 gnd.n4524 gnd.n2123 9.3005
R17341 gnd.n4570 gnd.n2122 9.3005
R17342 gnd.n4572 gnd.n4571 9.3005
R17343 gnd.n4111 gnd.n4110 9.3005
R17344 gnd.n4119 gnd.n4118 9.3005
R17345 gnd.n4120 gnd.n4029 9.3005
R17346 gnd.n4121 gnd.n4028 9.3005
R17347 gnd.n4027 gnd.n4025 9.3005
R17348 gnd.n4127 gnd.n4024 9.3005
R17349 gnd.n4128 gnd.n4023 9.3005
R17350 gnd.n4129 gnd.n4022 9.3005
R17351 gnd.n4021 gnd.n4019 9.3005
R17352 gnd.n4135 gnd.n4018 9.3005
R17353 gnd.n4136 gnd.n4017 9.3005
R17354 gnd.n4137 gnd.n4016 9.3005
R17355 gnd.n4015 gnd.n4013 9.3005
R17356 gnd.n4143 gnd.n4012 9.3005
R17357 gnd.n4144 gnd.n4011 9.3005
R17358 gnd.n4145 gnd.n4010 9.3005
R17359 gnd.n4009 gnd.n4007 9.3005
R17360 gnd.n4151 gnd.n4006 9.3005
R17361 gnd.n4152 gnd.n4005 9.3005
R17362 gnd.n4153 gnd.n4004 9.3005
R17363 gnd.n4003 gnd.n3998 9.3005
R17364 gnd.n4159 gnd.n3997 9.3005
R17365 gnd.n4160 gnd.n3996 9.3005
R17366 gnd.n4161 gnd.n3995 9.3005
R17367 gnd.n3994 gnd.n3992 9.3005
R17368 gnd.n4167 gnd.n3991 9.3005
R17369 gnd.n4168 gnd.n3990 9.3005
R17370 gnd.n4169 gnd.n3989 9.3005
R17371 gnd.n3988 gnd.n3986 9.3005
R17372 gnd.n4175 gnd.n3985 9.3005
R17373 gnd.n4176 gnd.n3984 9.3005
R17374 gnd.n4177 gnd.n3983 9.3005
R17375 gnd.n3982 gnd.n3980 9.3005
R17376 gnd.n4182 gnd.n3979 9.3005
R17377 gnd.n4183 gnd.n3978 9.3005
R17378 gnd.n3977 gnd.n3975 9.3005
R17379 gnd.n4188 gnd.n3974 9.3005
R17380 gnd.n4190 gnd.n4189 9.3005
R17381 gnd.n4117 gnd.n4034 9.3005
R17382 gnd.n4116 gnd.n4115 9.3005
R17383 gnd.n2326 gnd.n2325 9.3005
R17384 gnd.n4205 gnd.n4204 9.3005
R17385 gnd.n4206 gnd.n2324 9.3005
R17386 gnd.n4208 gnd.n4207 9.3005
R17387 gnd.n2310 gnd.n2309 9.3005
R17388 gnd.n4221 gnd.n4220 9.3005
R17389 gnd.n4222 gnd.n2308 9.3005
R17390 gnd.n4224 gnd.n4223 9.3005
R17391 gnd.n2294 gnd.n2293 9.3005
R17392 gnd.n4237 gnd.n4236 9.3005
R17393 gnd.n4238 gnd.n2292 9.3005
R17394 gnd.n4240 gnd.n4239 9.3005
R17395 gnd.n2278 gnd.n2277 9.3005
R17396 gnd.n4253 gnd.n4252 9.3005
R17397 gnd.n4254 gnd.n2276 9.3005
R17398 gnd.n4256 gnd.n4255 9.3005
R17399 gnd.n2262 gnd.n2261 9.3005
R17400 gnd.n4269 gnd.n4268 9.3005
R17401 gnd.n4270 gnd.n2260 9.3005
R17402 gnd.n4272 gnd.n4271 9.3005
R17403 gnd.n2246 gnd.n2245 9.3005
R17404 gnd.n4285 gnd.n4284 9.3005
R17405 gnd.n4286 gnd.n2244 9.3005
R17406 gnd.n4289 gnd.n4288 9.3005
R17407 gnd.n4287 gnd.n2229 9.3005
R17408 gnd.n4301 gnd.n2230 9.3005
R17409 gnd.n6539 gnd.n978 9.3005
R17410 gnd.n6538 gnd.n979 9.3005
R17411 gnd.n6537 gnd.n980 9.3005
R17412 gnd.n999 gnd.n981 9.3005
R17413 gnd.n6527 gnd.n1000 9.3005
R17414 gnd.n6526 gnd.n1001 9.3005
R17415 gnd.n6525 gnd.n1002 9.3005
R17416 gnd.n1020 gnd.n1003 9.3005
R17417 gnd.n6515 gnd.n1021 9.3005
R17418 gnd.n6514 gnd.n1022 9.3005
R17419 gnd.n6513 gnd.n1023 9.3005
R17420 gnd.n1041 gnd.n1024 9.3005
R17421 gnd.n6503 gnd.n1042 9.3005
R17422 gnd.n6502 gnd.n1043 9.3005
R17423 gnd.n6501 gnd.n1044 9.3005
R17424 gnd.n1062 gnd.n1045 9.3005
R17425 gnd.n6491 gnd.n1063 9.3005
R17426 gnd.n6490 gnd.n1064 9.3005
R17427 gnd.n6489 gnd.n1065 9.3005
R17428 gnd.n1083 gnd.n1066 9.3005
R17429 gnd.n6479 gnd.n1084 9.3005
R17430 gnd.n6478 gnd.n1085 9.3005
R17431 gnd.n6477 gnd.n1086 9.3005
R17432 gnd.n1104 gnd.n1087 9.3005
R17433 gnd.n6467 gnd.n1105 9.3005
R17434 gnd.n6466 gnd.n1106 9.3005
R17435 gnd.n6465 gnd.n1107 9.3005
R17436 gnd.n4192 gnd.n4191 9.3005
R17437 gnd.n977 gnd.n966 9.3005
R17438 gnd.n6549 gnd.n965 9.3005
R17439 gnd.n964 gnd.n960 9.3005
R17440 gnd.n6555 gnd.n959 9.3005
R17441 gnd.n6556 gnd.n958 9.3005
R17442 gnd.n6557 gnd.n957 9.3005
R17443 gnd.n956 gnd.n952 9.3005
R17444 gnd.n6563 gnd.n951 9.3005
R17445 gnd.n6564 gnd.n950 9.3005
R17446 gnd.n6565 gnd.n949 9.3005
R17447 gnd.n948 gnd.n944 9.3005
R17448 gnd.n6571 gnd.n943 9.3005
R17449 gnd.n6572 gnd.n942 9.3005
R17450 gnd.n6573 gnd.n941 9.3005
R17451 gnd.n940 gnd.n936 9.3005
R17452 gnd.n6579 gnd.n935 9.3005
R17453 gnd.n6580 gnd.n934 9.3005
R17454 gnd.n6581 gnd.n933 9.3005
R17455 gnd.n932 gnd.n928 9.3005
R17456 gnd.n6587 gnd.n927 9.3005
R17457 gnd.n6588 gnd.n926 9.3005
R17458 gnd.n6589 gnd.n925 9.3005
R17459 gnd.n924 gnd.n920 9.3005
R17460 gnd.n6595 gnd.n919 9.3005
R17461 gnd.n6596 gnd.n918 9.3005
R17462 gnd.n6597 gnd.n917 9.3005
R17463 gnd.n916 gnd.n912 9.3005
R17464 gnd.n6603 gnd.n911 9.3005
R17465 gnd.n6604 gnd.n910 9.3005
R17466 gnd.n6605 gnd.n909 9.3005
R17467 gnd.n908 gnd.n904 9.3005
R17468 gnd.n6611 gnd.n903 9.3005
R17469 gnd.n6612 gnd.n902 9.3005
R17470 gnd.n6613 gnd.n901 9.3005
R17471 gnd.n900 gnd.n896 9.3005
R17472 gnd.n6619 gnd.n895 9.3005
R17473 gnd.n6620 gnd.n894 9.3005
R17474 gnd.n6621 gnd.n893 9.3005
R17475 gnd.n892 gnd.n888 9.3005
R17476 gnd.n6627 gnd.n887 9.3005
R17477 gnd.n6628 gnd.n886 9.3005
R17478 gnd.n6629 gnd.n885 9.3005
R17479 gnd.n884 gnd.n880 9.3005
R17480 gnd.n6635 gnd.n879 9.3005
R17481 gnd.n6636 gnd.n878 9.3005
R17482 gnd.n6637 gnd.n877 9.3005
R17483 gnd.n876 gnd.n872 9.3005
R17484 gnd.n6643 gnd.n871 9.3005
R17485 gnd.n6644 gnd.n870 9.3005
R17486 gnd.n6645 gnd.n869 9.3005
R17487 gnd.n868 gnd.n864 9.3005
R17488 gnd.n6651 gnd.n863 9.3005
R17489 gnd.n6652 gnd.n862 9.3005
R17490 gnd.n6653 gnd.n861 9.3005
R17491 gnd.n860 gnd.n856 9.3005
R17492 gnd.n6659 gnd.n855 9.3005
R17493 gnd.n6660 gnd.n854 9.3005
R17494 gnd.n6661 gnd.n853 9.3005
R17495 gnd.n852 gnd.n848 9.3005
R17496 gnd.n6667 gnd.n847 9.3005
R17497 gnd.n6668 gnd.n846 9.3005
R17498 gnd.n6669 gnd.n845 9.3005
R17499 gnd.n844 gnd.n840 9.3005
R17500 gnd.n6675 gnd.n839 9.3005
R17501 gnd.n6676 gnd.n838 9.3005
R17502 gnd.n6677 gnd.n837 9.3005
R17503 gnd.n836 gnd.n832 9.3005
R17504 gnd.n6683 gnd.n831 9.3005
R17505 gnd.n6684 gnd.n830 9.3005
R17506 gnd.n6685 gnd.n829 9.3005
R17507 gnd.n828 gnd.n824 9.3005
R17508 gnd.n6691 gnd.n823 9.3005
R17509 gnd.n6692 gnd.n822 9.3005
R17510 gnd.n6693 gnd.n821 9.3005
R17511 gnd.n820 gnd.n816 9.3005
R17512 gnd.n6699 gnd.n815 9.3005
R17513 gnd.n6700 gnd.n814 9.3005
R17514 gnd.n6701 gnd.n813 9.3005
R17515 gnd.n812 gnd.n808 9.3005
R17516 gnd.n6707 gnd.n807 9.3005
R17517 gnd.n6708 gnd.n806 9.3005
R17518 gnd.n6709 gnd.n805 9.3005
R17519 gnd.n804 gnd.n800 9.3005
R17520 gnd.n6715 gnd.n799 9.3005
R17521 gnd.n6717 gnd.n6716 9.3005
R17522 gnd.n6548 gnd.n6547 9.3005
R17523 gnd.n1530 gnd.n1529 9.3005
R17524 gnd.n1516 gnd.n1512 9.3005
R17525 gnd.n1537 gnd.n1536 9.3005
R17526 gnd.n1538 gnd.n1507 9.3005
R17527 gnd.n1549 gnd.n1548 9.3005
R17528 gnd.n1509 gnd.n1505 9.3005
R17529 gnd.n1556 gnd.n1555 9.3005
R17530 gnd.n1557 gnd.n1500 9.3005
R17531 gnd.n1568 gnd.n1567 9.3005
R17532 gnd.n1502 gnd.n1498 9.3005
R17533 gnd.n1575 gnd.n1574 9.3005
R17534 gnd.n1495 gnd.n1494 9.3005
R17535 gnd.n1584 gnd.n1583 9.3005
R17536 gnd.n1492 gnd.n1491 9.3005
R17537 gnd.n1591 gnd.n1590 9.3005
R17538 gnd.n1483 gnd.n1482 9.3005
R17539 gnd.n1598 gnd.n1597 9.3005
R17540 gnd.n1480 gnd.n1478 9.3005
R17541 gnd.n1519 gnd.n1514 9.3005
R17542 gnd.n1593 gnd.n1592 9.3005
R17543 gnd.n1582 gnd.n1488 9.3005
R17544 gnd.n1581 gnd.n1580 9.3005
R17545 gnd.n1577 gnd.n1576 9.3005
R17546 gnd.n1497 gnd.n1496 9.3005
R17547 gnd.n1566 gnd.n1565 9.3005
R17548 gnd.n1562 gnd.n1501 9.3005
R17549 gnd.n1559 gnd.n1558 9.3005
R17550 gnd.n1504 gnd.n1503 9.3005
R17551 gnd.n1547 gnd.n1546 9.3005
R17552 gnd.n1543 gnd.n1508 9.3005
R17553 gnd.n1540 gnd.n1539 9.3005
R17554 gnd.n1511 gnd.n1510 9.3005
R17555 gnd.n1528 gnd.n1527 9.3005
R17556 gnd.n1524 gnd.n1515 9.3005
R17557 gnd.n1521 gnd.n1520 9.3005
R17558 gnd.n1594 gnd.n1484 9.3005
R17559 gnd.n1596 gnd.n1595 9.3005
R17560 gnd.n6040 gnd.n6039 9.3005
R17561 gnd.n6038 gnd.n1479 9.3005
R17562 gnd.n6037 gnd.n6036 9.3005
R17563 gnd.n6035 gnd.n1606 9.3005
R17564 gnd.n6034 gnd.n6033 9.3005
R17565 gnd.n6032 gnd.n1607 9.3005
R17566 gnd.n6028 gnd.n6027 9.3005
R17567 gnd.n6026 gnd.n1614 9.3005
R17568 gnd.n6025 gnd.n6024 9.3005
R17569 gnd.n6023 gnd.n6018 9.3005
R17570 gnd.n5613 gnd.n5612 9.3005
R17571 gnd.n1958 gnd.n1957 9.3005
R17572 gnd.n5626 gnd.n5625 9.3005
R17573 gnd.n5627 gnd.n1956 9.3005
R17574 gnd.n5629 gnd.n5628 9.3005
R17575 gnd.n1945 gnd.n1944 9.3005
R17576 gnd.n5642 gnd.n5641 9.3005
R17577 gnd.n5643 gnd.n1943 9.3005
R17578 gnd.n5645 gnd.n5644 9.3005
R17579 gnd.n1932 gnd.n1931 9.3005
R17580 gnd.n5658 gnd.n5657 9.3005
R17581 gnd.n5659 gnd.n1930 9.3005
R17582 gnd.n5661 gnd.n5660 9.3005
R17583 gnd.n1918 gnd.n1917 9.3005
R17584 gnd.n5674 gnd.n5673 9.3005
R17585 gnd.n5675 gnd.n1916 9.3005
R17586 gnd.n5677 gnd.n5676 9.3005
R17587 gnd.n1903 gnd.n1902 9.3005
R17588 gnd.n5690 gnd.n5689 9.3005
R17589 gnd.n5691 gnd.n1901 9.3005
R17590 gnd.n5693 gnd.n5692 9.3005
R17591 gnd.n1889 gnd.n1888 9.3005
R17592 gnd.n5706 gnd.n5705 9.3005
R17593 gnd.n5707 gnd.n1887 9.3005
R17594 gnd.n5709 gnd.n5708 9.3005
R17595 gnd.n1875 gnd.n1874 9.3005
R17596 gnd.n5722 gnd.n5721 9.3005
R17597 gnd.n5723 gnd.n1873 9.3005
R17598 gnd.n5725 gnd.n5724 9.3005
R17599 gnd.n1861 gnd.n1860 9.3005
R17600 gnd.n5738 gnd.n5737 9.3005
R17601 gnd.n5739 gnd.n1859 9.3005
R17602 gnd.n5741 gnd.n5740 9.3005
R17603 gnd.n1847 gnd.n1846 9.3005
R17604 gnd.n5754 gnd.n5753 9.3005
R17605 gnd.n5755 gnd.n1845 9.3005
R17606 gnd.n5757 gnd.n5756 9.3005
R17607 gnd.n1833 gnd.n1832 9.3005
R17608 gnd.n5770 gnd.n5769 9.3005
R17609 gnd.n5771 gnd.n1831 9.3005
R17610 gnd.n5773 gnd.n5772 9.3005
R17611 gnd.n1817 gnd.n1816 9.3005
R17612 gnd.n5786 gnd.n5785 9.3005
R17613 gnd.n5787 gnd.n1815 9.3005
R17614 gnd.n5789 gnd.n5788 9.3005
R17615 gnd.n1802 gnd.n1801 9.3005
R17616 gnd.n5802 gnd.n5801 9.3005
R17617 gnd.n5803 gnd.n1800 9.3005
R17618 gnd.n5805 gnd.n5804 9.3005
R17619 gnd.n1787 gnd.n1786 9.3005
R17620 gnd.n5818 gnd.n5817 9.3005
R17621 gnd.n5819 gnd.n1785 9.3005
R17622 gnd.n5821 gnd.n5820 9.3005
R17623 gnd.n1773 gnd.n1772 9.3005
R17624 gnd.n5834 gnd.n5833 9.3005
R17625 gnd.n5835 gnd.n1771 9.3005
R17626 gnd.n5837 gnd.n5836 9.3005
R17627 gnd.n1758 gnd.n1757 9.3005
R17628 gnd.n5850 gnd.n5849 9.3005
R17629 gnd.n5851 gnd.n1756 9.3005
R17630 gnd.n5853 gnd.n5852 9.3005
R17631 gnd.n1743 gnd.n1742 9.3005
R17632 gnd.n5866 gnd.n5865 9.3005
R17633 gnd.n5867 gnd.n1741 9.3005
R17634 gnd.n5869 gnd.n5868 9.3005
R17635 gnd.n1729 gnd.n1728 9.3005
R17636 gnd.n5882 gnd.n5881 9.3005
R17637 gnd.n5883 gnd.n1727 9.3005
R17638 gnd.n5885 gnd.n5884 9.3005
R17639 gnd.n1715 gnd.n1714 9.3005
R17640 gnd.n5898 gnd.n5897 9.3005
R17641 gnd.n5899 gnd.n1713 9.3005
R17642 gnd.n5901 gnd.n5900 9.3005
R17643 gnd.n1699 gnd.n1698 9.3005
R17644 gnd.n5914 gnd.n5913 9.3005
R17645 gnd.n5915 gnd.n1697 9.3005
R17646 gnd.n5917 gnd.n5916 9.3005
R17647 gnd.n1684 gnd.n1683 9.3005
R17648 gnd.n5930 gnd.n5929 9.3005
R17649 gnd.n5931 gnd.n1682 9.3005
R17650 gnd.n5933 gnd.n5932 9.3005
R17651 gnd.n1671 gnd.n1670 9.3005
R17652 gnd.n5946 gnd.n5945 9.3005
R17653 gnd.n5947 gnd.n1669 9.3005
R17654 gnd.n5949 gnd.n5948 9.3005
R17655 gnd.n1658 gnd.n1657 9.3005
R17656 gnd.n5962 gnd.n5961 9.3005
R17657 gnd.n5963 gnd.n1656 9.3005
R17658 gnd.n5965 gnd.n5964 9.3005
R17659 gnd.n1644 gnd.n1643 9.3005
R17660 gnd.n5978 gnd.n5977 9.3005
R17661 gnd.n5979 gnd.n1642 9.3005
R17662 gnd.n5981 gnd.n5980 9.3005
R17663 gnd.n1631 gnd.n1630 9.3005
R17664 gnd.n5994 gnd.n5993 9.3005
R17665 gnd.n5995 gnd.n1628 9.3005
R17666 gnd.n5999 gnd.n5998 9.3005
R17667 gnd.n5997 gnd.n1629 9.3005
R17668 gnd.n5996 gnd.n1616 9.3005
R17669 gnd.n6015 gnd.n1615 9.3005
R17670 gnd.n6017 gnd.n6016 9.3005
R17671 gnd.n5611 gnd.n1969 9.3005
R17672 gnd.n1971 gnd.n1970 9.3005
R17673 gnd.n4549 gnd.n4546 9.3005
R17674 gnd.n4551 gnd.n4550 9.3005
R17675 gnd.n4553 gnd.n4552 9.3005
R17676 gnd.n4554 gnd.n4539 9.3005
R17677 gnd.n4556 gnd.n4555 9.3005
R17678 gnd.n4557 gnd.n4538 9.3005
R17679 gnd.n4559 gnd.n4558 9.3005
R17680 gnd.n4560 gnd.n4533 9.3005
R17681 gnd.n5610 gnd.n5609 9.3005
R17682 gnd.n3922 gnd.n3911 9.3005
R17683 gnd.n3921 gnd.n3920 9.3005
R17684 gnd.n3919 gnd.n3912 9.3005
R17685 gnd.n3918 gnd.n3917 9.3005
R17686 gnd.n3916 gnd.n3915 9.3005
R17687 gnd.n2180 gnd.n2179 9.3005
R17688 gnd.n4362 gnd.n4361 9.3005
R17689 gnd.n4363 gnd.n2178 9.3005
R17690 gnd.n4365 gnd.n4364 9.3005
R17691 gnd.n2170 gnd.n2168 9.3005
R17692 gnd.n4406 gnd.n4405 9.3005
R17693 gnd.n4404 gnd.n2169 9.3005
R17694 gnd.n4403 gnd.n4402 9.3005
R17695 gnd.n4401 gnd.n2171 9.3005
R17696 gnd.n4400 gnd.n4399 9.3005
R17697 gnd.n4398 gnd.n4395 9.3005
R17698 gnd.n4397 gnd.n4396 9.3005
R17699 gnd.n2149 gnd.n2147 9.3005
R17700 gnd.n4455 gnd.n4454 9.3005
R17701 gnd.n4453 gnd.n2148 9.3005
R17702 gnd.n4452 gnd.n4451 9.3005
R17703 gnd.n4450 gnd.n2150 9.3005
R17704 gnd.n4449 gnd.n4448 9.3005
R17705 gnd.n2134 gnd.n2133 9.3005
R17706 gnd.n4514 gnd.n4513 9.3005
R17707 gnd.n4515 gnd.n2132 9.3005
R17708 gnd.n4517 gnd.n4516 9.3005
R17709 gnd.n2128 gnd.n2127 9.3005
R17710 gnd.n4531 gnd.n4530 9.3005
R17711 gnd.n4532 gnd.n2125 9.3005
R17712 gnd.n4566 gnd.n4565 9.3005
R17713 gnd.n4564 gnd.n2126 9.3005
R17714 gnd.n4562 gnd.n4561 9.3005
R17715 gnd.n2040 gnd.n2039 9.3005
R17716 gnd.n5562 gnd.n5561 9.3005
R17717 gnd.n5564 gnd.n5563 9.3005
R17718 gnd.n2028 gnd.n2027 9.3005
R17719 gnd.n5570 gnd.n5569 9.3005
R17720 gnd.n5572 gnd.n5571 9.3005
R17721 gnd.n2020 gnd.n2019 9.3005
R17722 gnd.n5578 gnd.n5577 9.3005
R17723 gnd.n5580 gnd.n5579 9.3005
R17724 gnd.n2010 gnd.n2009 9.3005
R17725 gnd.n5586 gnd.n5585 9.3005
R17726 gnd.n5588 gnd.n5587 9.3005
R17727 gnd.n2002 gnd.n2001 9.3005
R17728 gnd.n5594 gnd.n5593 9.3005
R17729 gnd.n5596 gnd.n5595 9.3005
R17730 gnd.n1992 gnd.n1990 9.3005
R17731 gnd.n5602 gnd.n5601 9.3005
R17732 gnd.n5603 gnd.n1989 9.3005
R17733 gnd.n2043 gnd.n1116 9.3005
R17734 gnd.n1993 gnd.n1991 9.3005
R17735 gnd.n5600 gnd.n5599 9.3005
R17736 gnd.n5598 gnd.n5597 9.3005
R17737 gnd.n1997 gnd.n1996 9.3005
R17738 gnd.n5592 gnd.n5591 9.3005
R17739 gnd.n5590 gnd.n5589 9.3005
R17740 gnd.n2006 gnd.n2005 9.3005
R17741 gnd.n5584 gnd.n5583 9.3005
R17742 gnd.n5582 gnd.n5581 9.3005
R17743 gnd.n2014 gnd.n2013 9.3005
R17744 gnd.n5576 gnd.n5575 9.3005
R17745 gnd.n5574 gnd.n5573 9.3005
R17746 gnd.n2024 gnd.n2023 9.3005
R17747 gnd.n5568 gnd.n5567 9.3005
R17748 gnd.n5566 gnd.n5565 9.3005
R17749 gnd.n2034 gnd.n2033 9.3005
R17750 gnd.n5560 gnd.n5559 9.3005
R17751 gnd.n6455 gnd.n1117 9.3005
R17752 gnd.n6454 gnd.n6453 9.3005
R17753 gnd.n6452 gnd.n1121 9.3005
R17754 gnd.n6451 gnd.n6450 9.3005
R17755 gnd.n6449 gnd.n1122 9.3005
R17756 gnd.n6448 gnd.n6447 9.3005
R17757 gnd.n6446 gnd.n1126 9.3005
R17758 gnd.n6445 gnd.n6444 9.3005
R17759 gnd.n6443 gnd.n1127 9.3005
R17760 gnd.n6442 gnd.n6441 9.3005
R17761 gnd.n6440 gnd.n1131 9.3005
R17762 gnd.n6439 gnd.n6438 9.3005
R17763 gnd.n6437 gnd.n1132 9.3005
R17764 gnd.n6436 gnd.n6435 9.3005
R17765 gnd.n6434 gnd.n1136 9.3005
R17766 gnd.n6433 gnd.n6432 9.3005
R17767 gnd.n6431 gnd.n1137 9.3005
R17768 gnd.n6430 gnd.n6429 9.3005
R17769 gnd.n6428 gnd.n1141 9.3005
R17770 gnd.n6427 gnd.n6426 9.3005
R17771 gnd.n6425 gnd.n1142 9.3005
R17772 gnd.n6424 gnd.n6423 9.3005
R17773 gnd.n6422 gnd.n1146 9.3005
R17774 gnd.n6421 gnd.n6420 9.3005
R17775 gnd.n6419 gnd.n1147 9.3005
R17776 gnd.n6418 gnd.n6417 9.3005
R17777 gnd.n6416 gnd.n1151 9.3005
R17778 gnd.n6415 gnd.n6414 9.3005
R17779 gnd.n6413 gnd.n1152 9.3005
R17780 gnd.n6412 gnd.n6411 9.3005
R17781 gnd.n6410 gnd.n1156 9.3005
R17782 gnd.n6409 gnd.n6408 9.3005
R17783 gnd.n6407 gnd.n1157 9.3005
R17784 gnd.n6406 gnd.n6405 9.3005
R17785 gnd.n6404 gnd.n1161 9.3005
R17786 gnd.n6403 gnd.n6402 9.3005
R17787 gnd.n6401 gnd.n1162 9.3005
R17788 gnd.n6400 gnd.n6399 9.3005
R17789 gnd.n6398 gnd.n1166 9.3005
R17790 gnd.n6397 gnd.n6396 9.3005
R17791 gnd.n6395 gnd.n1167 9.3005
R17792 gnd.n6394 gnd.n6393 9.3005
R17793 gnd.n6392 gnd.n1171 9.3005
R17794 gnd.n6391 gnd.n6390 9.3005
R17795 gnd.n6389 gnd.n1172 9.3005
R17796 gnd.n6388 gnd.n6387 9.3005
R17797 gnd.n6386 gnd.n1176 9.3005
R17798 gnd.n6385 gnd.n6384 9.3005
R17799 gnd.n6383 gnd.n1177 9.3005
R17800 gnd.n6382 gnd.n6381 9.3005
R17801 gnd.n6380 gnd.n1181 9.3005
R17802 gnd.n6379 gnd.n6378 9.3005
R17803 gnd.n6377 gnd.n1182 9.3005
R17804 gnd.n6376 gnd.n6375 9.3005
R17805 gnd.n6374 gnd.n1186 9.3005
R17806 gnd.n6373 gnd.n6372 9.3005
R17807 gnd.n6371 gnd.n1187 9.3005
R17808 gnd.n6370 gnd.n6369 9.3005
R17809 gnd.n6368 gnd.n1191 9.3005
R17810 gnd.n6367 gnd.n6366 9.3005
R17811 gnd.n6365 gnd.n1192 9.3005
R17812 gnd.n6364 gnd.n6363 9.3005
R17813 gnd.n6362 gnd.n1196 9.3005
R17814 gnd.n6361 gnd.n6360 9.3005
R17815 gnd.n6359 gnd.n1197 9.3005
R17816 gnd.n6358 gnd.n6357 9.3005
R17817 gnd.n6356 gnd.n1201 9.3005
R17818 gnd.n6355 gnd.n6354 9.3005
R17819 gnd.n6353 gnd.n1202 9.3005
R17820 gnd.n6352 gnd.n6351 9.3005
R17821 gnd.n6350 gnd.n1206 9.3005
R17822 gnd.n6349 gnd.n6348 9.3005
R17823 gnd.n6347 gnd.n1207 9.3005
R17824 gnd.n6346 gnd.n6345 9.3005
R17825 gnd.n6344 gnd.n1211 9.3005
R17826 gnd.n6343 gnd.n6342 9.3005
R17827 gnd.n6341 gnd.n1212 9.3005
R17828 gnd.n6340 gnd.n6339 9.3005
R17829 gnd.n6338 gnd.n1216 9.3005
R17830 gnd.n6337 gnd.n6336 9.3005
R17831 gnd.n6335 gnd.n1217 9.3005
R17832 gnd.n6334 gnd.n6333 9.3005
R17833 gnd.n6332 gnd.n1221 9.3005
R17834 gnd.n6331 gnd.n6330 9.3005
R17835 gnd.n6329 gnd.n1222 9.3005
R17836 gnd.n6328 gnd.n6327 9.3005
R17837 gnd.n6326 gnd.n1226 9.3005
R17838 gnd.n6325 gnd.n6324 9.3005
R17839 gnd.n6323 gnd.n1227 9.3005
R17840 gnd.n6322 gnd.n6321 9.3005
R17841 gnd.n6320 gnd.n1231 9.3005
R17842 gnd.n6319 gnd.n6318 9.3005
R17843 gnd.n6317 gnd.n1232 9.3005
R17844 gnd.n6316 gnd.n6315 9.3005
R17845 gnd.n6314 gnd.n1236 9.3005
R17846 gnd.n6313 gnd.n6312 9.3005
R17847 gnd.n6311 gnd.n1237 9.3005
R17848 gnd.n6310 gnd.n6309 9.3005
R17849 gnd.n6308 gnd.n1241 9.3005
R17850 gnd.n6307 gnd.n6306 9.3005
R17851 gnd.n6305 gnd.n1242 9.3005
R17852 gnd.n6457 gnd.n6456 9.3005
R17853 gnd.n6214 gnd.n1341 9.3005
R17854 gnd.n6213 gnd.n6212 9.3005
R17855 gnd.n6211 gnd.n1343 9.3005
R17856 gnd.n6210 gnd.n6209 9.3005
R17857 gnd.n6208 gnd.n1347 9.3005
R17858 gnd.n6207 gnd.n6206 9.3005
R17859 gnd.n6205 gnd.n1348 9.3005
R17860 gnd.n6204 gnd.n6203 9.3005
R17861 gnd.n6202 gnd.n1352 9.3005
R17862 gnd.n6201 gnd.n6200 9.3005
R17863 gnd.n6199 gnd.n1353 9.3005
R17864 gnd.n6198 gnd.n6197 9.3005
R17865 gnd.n6196 gnd.n1357 9.3005
R17866 gnd.n6195 gnd.n6194 9.3005
R17867 gnd.n6193 gnd.n1358 9.3005
R17868 gnd.n6192 gnd.n6191 9.3005
R17869 gnd.n407 gnd.n405 9.3005
R17870 gnd.n7372 gnd.n7371 9.3005
R17871 gnd.n7370 gnd.n406 9.3005
R17872 gnd.n7369 gnd.n7368 9.3005
R17873 gnd.n7367 gnd.n408 9.3005
R17874 gnd.n375 gnd.n373 9.3005
R17875 gnd.n7418 gnd.n7417 9.3005
R17876 gnd.n7416 gnd.n374 9.3005
R17877 gnd.n7415 gnd.n7414 9.3005
R17878 gnd.n7413 gnd.n376 9.3005
R17879 gnd.n7412 gnd.n7411 9.3005
R17880 gnd.n320 gnd.n318 9.3005
R17881 gnd.n7549 gnd.n7548 9.3005
R17882 gnd.n7547 gnd.n319 9.3005
R17883 gnd.n7546 gnd.n7545 9.3005
R17884 gnd.n7544 gnd.n321 9.3005
R17885 gnd.n7543 gnd.n7542 9.3005
R17886 gnd.n7541 gnd.n325 9.3005
R17887 gnd.n7540 gnd.n7539 9.3005
R17888 gnd.n7538 gnd.n326 9.3005
R17889 gnd.n297 gnd.n296 9.3005
R17890 gnd.n7563 gnd.n7562 9.3005
R17891 gnd.n7564 gnd.n295 9.3005
R17892 gnd.n7566 gnd.n7565 9.3005
R17893 gnd.n281 gnd.n280 9.3005
R17894 gnd.n7579 gnd.n7578 9.3005
R17895 gnd.n7580 gnd.n279 9.3005
R17896 gnd.n7582 gnd.n7581 9.3005
R17897 gnd.n267 gnd.n266 9.3005
R17898 gnd.n7595 gnd.n7594 9.3005
R17899 gnd.n7596 gnd.n265 9.3005
R17900 gnd.n7598 gnd.n7597 9.3005
R17901 gnd.n251 gnd.n250 9.3005
R17902 gnd.n7611 gnd.n7610 9.3005
R17903 gnd.n7612 gnd.n249 9.3005
R17904 gnd.n7614 gnd.n7613 9.3005
R17905 gnd.n236 gnd.n235 9.3005
R17906 gnd.n7627 gnd.n7626 9.3005
R17907 gnd.n7628 gnd.n234 9.3005
R17908 gnd.n7630 gnd.n7629 9.3005
R17909 gnd.n221 gnd.n220 9.3005
R17910 gnd.n7643 gnd.n7642 9.3005
R17911 gnd.n7644 gnd.n218 9.3005
R17912 gnd.n7714 gnd.n7713 9.3005
R17913 gnd.n7712 gnd.n219 9.3005
R17914 gnd.n7711 gnd.n7710 9.3005
R17915 gnd.n7709 gnd.n7645 9.3005
R17916 gnd.n7708 gnd.n7707 9.3005
R17917 gnd.n6216 gnd.n6215 9.3005
R17918 gnd.n7704 gnd.n7647 9.3005
R17919 gnd.n7703 gnd.n7702 9.3005
R17920 gnd.n7701 gnd.n7652 9.3005
R17921 gnd.n7700 gnd.n7699 9.3005
R17922 gnd.n7698 gnd.n7653 9.3005
R17923 gnd.n7697 gnd.n7696 9.3005
R17924 gnd.n7695 gnd.n7660 9.3005
R17925 gnd.n7694 gnd.n7693 9.3005
R17926 gnd.n7692 gnd.n7661 9.3005
R17927 gnd.n7691 gnd.n7690 9.3005
R17928 gnd.n7689 gnd.n7668 9.3005
R17929 gnd.n7688 gnd.n7687 9.3005
R17930 gnd.n7686 gnd.n7669 9.3005
R17931 gnd.n7685 gnd.n7684 9.3005
R17932 gnd.n7683 gnd.n7676 9.3005
R17933 gnd.n7682 gnd.n7681 9.3005
R17934 gnd.n124 gnd.n121 9.3005
R17935 gnd.n7808 gnd.n7807 9.3005
R17936 gnd.n7706 gnd.n7705 9.3005
R17937 gnd.n6056 gnd.n6055 9.3005
R17938 gnd.n6057 gnd.n1476 9.3005
R17939 gnd.n6060 gnd.n6059 9.3005
R17940 gnd.n6058 gnd.n1477 9.3005
R17941 gnd.n1420 gnd.n1419 9.3005
R17942 gnd.n6087 gnd.n6086 9.3005
R17943 gnd.n6088 gnd.n1417 9.3005
R17944 gnd.n6096 gnd.n6095 9.3005
R17945 gnd.n6094 gnd.n1418 9.3005
R17946 gnd.n6093 gnd.n6092 9.3005
R17947 gnd.n6091 gnd.n6089 9.3005
R17948 gnd.n1384 gnd.n1382 9.3005
R17949 gnd.n6156 gnd.n6155 9.3005
R17950 gnd.n6154 gnd.n1383 9.3005
R17951 gnd.n6153 gnd.n6152 9.3005
R17952 gnd.n6151 gnd.n1385 9.3005
R17953 gnd.n6150 gnd.n6149 9.3005
R17954 gnd.n6148 gnd.n6140 9.3005
R17955 gnd.n6147 gnd.n6146 9.3005
R17956 gnd.n6145 gnd.n6142 9.3005
R17957 gnd.n6141 gnd.n382 9.3005
R17958 gnd.n7400 gnd.n381 9.3005
R17959 gnd.n7402 gnd.n7401 9.3005
R17960 gnd.n7403 gnd.n379 9.3005
R17961 gnd.n7406 gnd.n7405 9.3005
R17962 gnd.n7404 gnd.n380 9.3005
R17963 gnd.n348 gnd.n347 9.3005
R17964 gnd.n7447 gnd.n7446 9.3005
R17965 gnd.n7448 gnd.n346 9.3005
R17966 gnd.n7450 gnd.n7449 9.3005
R17967 gnd.n7451 gnd.n79 9.3005
R17968 gnd.n7857 gnd.n80 9.3005
R17969 gnd.n7856 gnd.n7855 9.3005
R17970 gnd.n7854 gnd.n81 9.3005
R17971 gnd.n7853 gnd.n7852 9.3005
R17972 gnd.n7851 gnd.n85 9.3005
R17973 gnd.n7850 gnd.n7849 9.3005
R17974 gnd.n7848 gnd.n86 9.3005
R17975 gnd.n7847 gnd.n7846 9.3005
R17976 gnd.n7845 gnd.n90 9.3005
R17977 gnd.n7844 gnd.n7843 9.3005
R17978 gnd.n7842 gnd.n91 9.3005
R17979 gnd.n7841 gnd.n7840 9.3005
R17980 gnd.n7839 gnd.n95 9.3005
R17981 gnd.n7838 gnd.n7837 9.3005
R17982 gnd.n7836 gnd.n96 9.3005
R17983 gnd.n7835 gnd.n7834 9.3005
R17984 gnd.n7833 gnd.n100 9.3005
R17985 gnd.n7832 gnd.n7831 9.3005
R17986 gnd.n7830 gnd.n101 9.3005
R17987 gnd.n7829 gnd.n7828 9.3005
R17988 gnd.n7827 gnd.n105 9.3005
R17989 gnd.n7826 gnd.n7825 9.3005
R17990 gnd.n7824 gnd.n106 9.3005
R17991 gnd.n7823 gnd.n7822 9.3005
R17992 gnd.n7821 gnd.n110 9.3005
R17993 gnd.n7820 gnd.n7819 9.3005
R17994 gnd.n7818 gnd.n111 9.3005
R17995 gnd.n7817 gnd.n7816 9.3005
R17996 gnd.n7815 gnd.n115 9.3005
R17997 gnd.n7814 gnd.n7813 9.3005
R17998 gnd.n7812 gnd.n116 9.3005
R17999 gnd.n7811 gnd.n7810 9.3005
R18000 gnd.n7809 gnd.n120 9.3005
R18001 gnd.n6043 gnd.n6042 9.3005
R18002 gnd.t123 gnd.n2524 9.24152
R18003 gnd.n2426 gnd.t253 9.24152
R18004 gnd.n3706 gnd.t245 9.24152
R18005 gnd.t70 gnd.n2271 9.24152
R18006 gnd.n2193 gnd.n2192 9.24152
R18007 gnd.t339 gnd.n1871 9.24152
R18008 gnd.n4795 gnd.t339 9.24152
R18009 gnd.n5895 gnd.t26 9.24152
R18010 gnd.n5248 gnd.t26 9.24152
R18011 gnd.n7551 gnd.n312 9.24152
R18012 gnd.n263 gnd.t67 9.24152
R18013 gnd.t16 gnd.t123 8.92286
R18014 gnd.t78 gnd.n1893 8.92286
R18015 gnd.n4973 gnd.t327 8.92286
R18016 gnd.n5217 gnd.t266 8.92286
R18017 gnd.n3676 gnd.n3651 8.92171
R18018 gnd.n3644 gnd.n3619 8.92171
R18019 gnd.n3612 gnd.n3587 8.92171
R18020 gnd.n3581 gnd.n3556 8.92171
R18021 gnd.n3549 gnd.n3524 8.92171
R18022 gnd.n3517 gnd.n3492 8.92171
R18023 gnd.n3485 gnd.n3460 8.92171
R18024 gnd.n3454 gnd.n3429 8.92171
R18025 gnd.n5024 gnd.n5006 8.72777
R18026 gnd.n3180 gnd.t14 8.60421
R18027 gnd.t174 gnd.n2303 8.60421
R18028 gnd.t337 gnd.n1797 8.60421
R18029 gnd.n4875 gnd.t30 8.60421
R18030 gnd.n232 gnd.t151 8.60421
R18031 gnd.n2604 gnd.n2584 8.43467
R18032 gnd.n58 gnd.n38 8.43467
R18033 gnd.n3923 gnd.n0 8.41456
R18034 gnd.n7858 gnd.n7857 8.41456
R18035 gnd.n5727 gnd.n1870 8.28555
R18036 gnd.n5364 gnd.n4824 8.28555
R18037 gnd.n5343 gnd.n5342 8.28555
R18038 gnd.n5831 gnd.n1777 8.28555
R18039 gnd.n5863 gnd.n1745 8.28555
R18040 gnd.n4943 gnd.n4942 8.28555
R18041 gnd.n5943 gnd.t266 8.28555
R18042 gnd.n3677 gnd.n3649 8.14595
R18043 gnd.n3645 gnd.n3617 8.14595
R18044 gnd.n3613 gnd.n3585 8.14595
R18045 gnd.n3582 gnd.n3554 8.14595
R18046 gnd.n3550 gnd.n3522 8.14595
R18047 gnd.n3518 gnd.n3490 8.14595
R18048 gnd.n3486 gnd.n3458 8.14595
R18049 gnd.n3455 gnd.n3427 8.14595
R18050 gnd.n3682 gnd.n3681 7.97301
R18051 gnd.t13 gnd.n2695 7.9669
R18052 gnd.n5606 gnd.n1973 7.9669
R18053 gnd.n5409 gnd.t84 7.9669
R18054 gnd.n1704 gnd.t0 7.9669
R18055 gnd.n1256 gnd.n1248 7.9669
R18056 gnd.n7807 gnd.n124 7.75808
R18057 gnd.n1595 gnd.n1594 7.75808
R18058 gnd.n5559 gnd.n2033 7.75808
R18059 gnd.n3876 gnd.n3815 7.75808
R18060 gnd.n6542 gnd.n970 7.64824
R18061 gnd.n6541 gnd.n973 7.64824
R18062 gnd.n4359 gnd.n983 7.64824
R18063 gnd.n6535 gnd.n986 7.64824
R18064 gnd.n4377 gnd.n4376 7.64824
R18065 gnd.n6529 gnd.n997 7.64824
R18066 gnd.n4409 gnd.n4408 7.64824
R18067 gnd.n6523 gnd.n1007 7.64824
R18068 gnd.n4385 gnd.n1015 7.64824
R18069 gnd.n6517 gnd.n1018 7.64824
R18070 gnd.n4393 gnd.n1026 7.64824
R18071 gnd.n6511 gnd.n1029 7.64824
R18072 gnd.n4426 gnd.n4425 7.64824
R18073 gnd.n6505 gnd.n1039 7.64824
R18074 gnd.n4458 gnd.n4457 7.64824
R18075 gnd.n6499 gnd.n1049 7.64824
R18076 gnd.n4434 gnd.n1057 7.64824
R18077 gnd.n6493 gnd.n1060 7.64824
R18078 gnd.n4446 gnd.n1068 7.64824
R18079 gnd.n6487 gnd.n1071 7.64824
R18080 gnd.n4511 gnd.n4510 7.64824
R18081 gnd.n6481 gnd.n1081 7.64824
R18082 gnd.n4519 gnd.n1089 7.64824
R18083 gnd.n6475 gnd.n1092 7.64824
R18084 gnd.n4528 gnd.n1100 7.64824
R18085 gnd.n4568 gnd.n1109 7.64824
R18086 gnd.n6463 gnd.n1112 7.64824
R18087 gnd.n5663 gnd.t263 7.64824
R18088 gnd.t160 gnd.n1870 7.64824
R18089 gnd.t164 gnd.n1821 7.64824
R18090 gnd.n5298 gnd.t33 7.64824
R18091 gnd.n4943 gnd.t6 7.64824
R18092 gnd.n6218 gnd.n1336 7.64824
R18093 gnd.n6053 gnd.n1338 7.64824
R18094 gnd.n6063 gnd.n6062 7.64824
R18095 gnd.n6074 gnd.n1431 7.64824
R18096 gnd.n6073 gnd.n1435 7.64824
R18097 gnd.n6084 gnd.n1422 7.64824
R18098 gnd.n1424 gnd.n1414 7.64824
R18099 gnd.n6099 gnd.n6098 7.64824
R18100 gnd.n6111 gnd.n1404 7.64824
R18101 gnd.n6109 gnd.n1407 7.64824
R18102 gnd.n6121 gnd.n1394 7.64824
R18103 gnd.n1398 gnd.n1396 7.64824
R18104 gnd.n6160 gnd.n6159 7.64824
R18105 gnd.n6181 gnd.n1370 7.64824
R18106 gnd.n6180 gnd.n1373 7.64824
R18107 gnd.n6189 gnd.n1361 7.64824
R18108 gnd.n6138 gnd.n1364 7.64824
R18109 gnd.n7374 gnd.n399 7.64824
R18110 gnd.n6143 gnd.n402 7.64824
R18111 gnd.n7384 gnd.n390 7.64824
R18112 gnd.n7365 gnd.n7364 7.64824
R18113 gnd.n7398 gnd.n384 7.64824
R18114 gnd.n7420 gnd.n367 7.64824
R18115 gnd.n7392 gnd.n370 7.64824
R18116 gnd.n7408 gnd.n377 7.64824
R18117 gnd.n7429 gnd.n356 7.64824
R18118 gnd.n358 gnd.n350 7.64824
R18119 gnd.n3089 gnd.t46 7.32958
R18120 gnd.t249 gnd.n1960 7.32958
R18121 gnd.n5655 gnd.t58 7.32958
R18122 gnd.n5523 gnd.n4652 7.32958
R18123 gnd.n5967 gnd.n1654 7.32958
R18124 gnd.t60 gnd.n1646 7.32958
R18125 gnd.n6012 gnd.t213 7.32958
R18126 gnd.n247 gnd.n238 7.32958
R18127 gnd.n4674 gnd.n4673 7.30353
R18128 gnd.n5023 gnd.n5022 7.30353
R18129 gnd.n3049 gnd.n2768 7.01093
R18130 gnd.n2771 gnd.n2769 7.01093
R18131 gnd.n3059 gnd.n3058 7.01093
R18132 gnd.n3070 gnd.n2752 7.01093
R18133 gnd.n3069 gnd.n2755 7.01093
R18134 gnd.n3080 gnd.n2743 7.01093
R18135 gnd.n2746 gnd.n2744 7.01093
R18136 gnd.n3090 gnd.n3089 7.01093
R18137 gnd.n3100 gnd.n2724 7.01093
R18138 gnd.n3099 gnd.n2727 7.01093
R18139 gnd.n3108 gnd.n2718 7.01093
R18140 gnd.n3120 gnd.n2708 7.01093
R18141 gnd.n3130 gnd.n2693 7.01093
R18142 gnd.n3146 gnd.n3145 7.01093
R18143 gnd.n2695 gnd.n2632 7.01093
R18144 gnd.n3200 gnd.n2633 7.01093
R18145 gnd.n3194 gnd.n3193 7.01093
R18146 gnd.n2682 gnd.n2644 7.01093
R18147 gnd.n3186 gnd.n2655 7.01093
R18148 gnd.n2673 gnd.n2668 7.01093
R18149 gnd.n3180 gnd.n3179 7.01093
R18150 gnd.n3226 gnd.n2559 7.01093
R18151 gnd.n3225 gnd.n3224 7.01093
R18152 gnd.n3237 gnd.n3236 7.01093
R18153 gnd.n2552 gnd.n2544 7.01093
R18154 gnd.n3266 gnd.n2532 7.01093
R18155 gnd.n3265 gnd.n2535 7.01093
R18156 gnd.n3276 gnd.n2524 7.01093
R18157 gnd.n2525 gnd.n2513 7.01093
R18158 gnd.n3287 gnd.n2514 7.01093
R18159 gnd.n3311 gnd.n2505 7.01093
R18160 gnd.n3310 gnd.n2496 7.01093
R18161 gnd.n3333 gnd.n3332 7.01093
R18162 gnd.n3351 gnd.n2477 7.01093
R18163 gnd.n3350 gnd.n2480 7.01093
R18164 gnd.n3361 gnd.n2469 7.01093
R18165 gnd.n2470 gnd.n2457 7.01093
R18166 gnd.n3372 gnd.n2458 7.01093
R18167 gnd.n3399 gnd.n2442 7.01093
R18168 gnd.n3411 gnd.n3410 7.01093
R18169 gnd.n3393 gnd.n2435 7.01093
R18170 gnd.n3422 gnd.n3421 7.01093
R18171 gnd.n3694 gnd.n2423 7.01093
R18172 gnd.n3693 gnd.n2426 7.01093
R18173 gnd.n3706 gnd.n2415 7.01093
R18174 gnd.n2416 gnd.n2407 7.01093
R18175 gnd.n3716 gnd.n2408 7.01093
R18176 gnd.n5453 gnd.n5452 7.01093
R18177 gnd.n5687 gnd.n1907 7.01093
R18178 gnd.n5371 gnd.n4816 7.01093
R18179 gnd.n5335 gnd.n4860 7.01093
R18180 gnd.n5823 gnd.n1783 7.01093
R18181 gnd.n5871 gnd.n1739 7.01093
R18182 gnd.n5219 gnd.n5218 7.01093
R18183 gnd.n5959 gnd.n1662 7.01093
R18184 gnd.n2727 gnd.t332 6.69227
R18185 gnd.n2535 gnd.t16 6.69227
R18186 gnd.n3400 gnd.t15 6.69227
R18187 gnd.n5127 gnd.n5126 6.5566
R18188 gnd.n4686 gnd.n4685 6.5566
R18189 gnd.n5464 gnd.n5460 6.5566
R18190 gnd.n5142 gnd.n5141 6.5566
R18191 gnd.n4550 gnd.n4545 6.20656
R18192 gnd.n7769 gnd.n7766 6.20656
R18193 gnd.n4153 gnd.n4002 6.20656
R18194 gnd.n6031 gnd.n6028 6.20656
R18195 gnd.t166 gnd.n3156 6.05496
R18196 gnd.n3157 gnd.t44 6.05496
R18197 gnd.t94 gnd.n2559 6.05496
R18198 gnd.t336 gnd.n3321 6.05496
R18199 gnd.n3679 gnd.n3649 5.81868
R18200 gnd.n3647 gnd.n3617 5.81868
R18201 gnd.n3615 gnd.n3585 5.81868
R18202 gnd.n3584 gnd.n3554 5.81868
R18203 gnd.n3552 gnd.n3522 5.81868
R18204 gnd.n3520 gnd.n3490 5.81868
R18205 gnd.n3488 gnd.n3458 5.81868
R18206 gnd.n3457 gnd.n3427 5.81868
R18207 gnd.n5679 gnd.n1914 5.73631
R18208 gnd.t210 gnd.n1907 5.73631
R18209 gnd.n5392 gnd.t116 5.73631
R18210 gnd.n5743 gnd.n1857 5.73631
R18211 gnd.n5379 gnd.n5378 5.73631
R18212 gnd.t198 gnd.n1827 5.73631
R18213 gnd.n4860 gnd.t5 5.73631
R18214 gnd.n5328 gnd.n5327 5.73631
R18215 gnd.n5815 gnd.n1791 5.73631
R18216 gnd.n5823 gnd.t313 5.73631
R18217 gnd.n5290 gnd.t28 5.73631
R18218 gnd.n5879 gnd.n1731 5.73631
R18219 gnd.n5261 gnd.n4927 5.73631
R18220 gnd.n5254 gnd.t96 5.73631
R18221 gnd.n5211 gnd.n4988 5.73631
R18222 gnd.n5196 gnd.t239 5.73631
R18223 gnd.n5050 gnd.n1305 5.62001
R18224 gnd.n5526 gnd.n4617 5.62001
R18225 gnd.n5526 gnd.n4618 5.62001
R18226 gnd.n5136 gnd.n1305 5.62001
R18227 gnd.n2908 gnd.n2903 5.4308
R18228 gnd.n3724 gnd.n2400 5.4308
R18229 gnd.n3224 gnd.t333 5.41765
R18230 gnd.t334 gnd.n3247 5.41765
R18231 gnd.t125 gnd.n2489 5.41765
R18232 gnd.n3677 gnd.n3676 5.04292
R18233 gnd.n3645 gnd.n3644 5.04292
R18234 gnd.n3613 gnd.n3612 5.04292
R18235 gnd.n3582 gnd.n3581 5.04292
R18236 gnd.n3550 gnd.n3549 5.04292
R18237 gnd.n3518 gnd.n3517 5.04292
R18238 gnd.n3486 gnd.n3485 5.04292
R18239 gnd.n3455 gnd.n3454 5.04292
R18240 gnd.n2624 gnd.n2623 4.82753
R18241 gnd.n78 gnd.n77 4.82753
R18242 gnd.n3187 gnd.t45 4.78034
R18243 gnd.n2514 gnd.t124 4.78034
R18244 gnd.t349 gnd.n4748 4.78034
R18245 gnd.n5378 gnd.t129 4.78034
R18246 gnd.t132 gnd.n1731 4.78034
R18247 gnd.n5951 gnd.t362 4.78034
R18248 gnd.n1654 gnd.t221 4.78034
R18249 gnd.n2629 gnd.n2626 4.74817
R18250 gnd.n2679 gnd.n2565 4.74817
R18251 gnd.n2666 gnd.n2564 4.74817
R18252 gnd.n2563 gnd.n2562 4.74817
R18253 gnd.n2675 gnd.n2626 4.74817
R18254 gnd.n2676 gnd.n2565 4.74817
R18255 gnd.n2678 gnd.n2564 4.74817
R18256 gnd.n2665 gnd.n2563 4.74817
R18257 gnd.n7555 gnd.n7554 4.74817
R18258 gnd.n341 gnd.n308 4.74817
R18259 gnd.n7456 gnd.n307 4.74817
R18260 gnd.n331 gnd.n306 4.74817
R18261 gnd.n7534 gnd.n305 4.74817
R18262 gnd.n7555 gnd.n309 4.74817
R18263 gnd.n7553 gnd.n308 4.74817
R18264 gnd.n342 gnd.n307 4.74817
R18265 gnd.n7457 gnd.n306 4.74817
R18266 gnd.n332 gnd.n305 4.74817
R18267 gnd.n4305 gnd.n4303 4.74817
R18268 gnd.n4318 gnd.n2214 4.74817
R18269 gnd.n4322 gnd.n4320 4.74817
R18270 gnd.n4345 gnd.n2188 4.74817
R18271 gnd.n4348 gnd.n4347 4.74817
R18272 gnd.n4303 gnd.n4302 4.74817
R18273 gnd.n4304 gnd.n2214 4.74817
R18274 gnd.n4320 gnd.n4319 4.74817
R18275 gnd.n4321 gnd.n2188 4.74817
R18276 gnd.n4347 gnd.n4346 4.74817
R18277 gnd.n2604 gnd.n2603 4.7074
R18278 gnd.n58 gnd.n57 4.7074
R18279 gnd.n2624 gnd.n2604 4.65959
R18280 gnd.n78 gnd.n58 4.65959
R18281 gnd.n6262 gnd.n1307 4.6132
R18282 gnd.n5527 gnd.n4616 4.6132
R18283 gnd.n5671 gnd.n1922 4.46168
R18284 gnd.n5438 gnd.n5437 4.46168
R18285 gnd.n5424 gnd.t62 4.46168
R18286 gnd.n5386 gnd.n4804 4.46168
R18287 gnd.n5751 gnd.n1849 4.46168
R18288 gnd.n5807 gnd.n1798 4.46168
R18289 gnd.n5320 gnd.n4873 4.46168
R18290 gnd.n5269 gnd.n5268 4.46168
R18291 gnd.n5887 gnd.n1724 4.46168
R18292 gnd.n5226 gnd.t127 4.46168
R18293 gnd.n5943 gnd.n1674 4.46168
R18294 gnd.n5204 gnd.n5203 4.46168
R18295 gnd.n5019 gnd.n5006 4.46111
R18296 gnd.n3662 gnd.n3658 4.38594
R18297 gnd.n3630 gnd.n3626 4.38594
R18298 gnd.n3598 gnd.n3594 4.38594
R18299 gnd.n3567 gnd.n3563 4.38594
R18300 gnd.n3535 gnd.n3531 4.38594
R18301 gnd.n3503 gnd.n3499 4.38594
R18302 gnd.n3471 gnd.n3467 4.38594
R18303 gnd.n3440 gnd.n3436 4.38594
R18304 gnd.n3673 gnd.n3651 4.26717
R18305 gnd.n3641 gnd.n3619 4.26717
R18306 gnd.n3609 gnd.n3587 4.26717
R18307 gnd.n3578 gnd.n3556 4.26717
R18308 gnd.n3546 gnd.n3524 4.26717
R18309 gnd.n3514 gnd.n3492 4.26717
R18310 gnd.n3482 gnd.n3460 4.26717
R18311 gnd.n3451 gnd.n3429 4.26717
R18312 gnd.n3131 gnd.t122 4.14303
R18313 gnd.n3361 gnd.t331 4.14303
R18314 gnd.n2124 gnd.t217 4.14303
R18315 gnd.n4853 gnd.t358 4.14303
R18316 gnd.t309 gnd.n1769 4.14303
R18317 gnd.n6044 gnd.t224 4.14303
R18318 gnd.n3681 gnd.n3680 4.08274
R18319 gnd.n5126 gnd.n5125 4.05904
R18320 gnd.n4687 gnd.n4686 4.05904
R18321 gnd.n5467 gnd.n5460 4.05904
R18322 gnd.n5143 gnd.n5142 4.05904
R18323 gnd.n19 gnd.n9 3.99943
R18324 gnd.n5438 gnd.t289 3.82437
R18325 gnd.n5695 gnd.t62 3.82437
R18326 gnd.n4816 gnd.t161 3.82437
R18327 gnd.n5871 gnd.t115 3.82437
R18328 gnd.n4961 gnd.t127 3.82437
R18329 gnd.n3681 gnd.n3553 3.70378
R18330 gnd.n3204 gnd.n2625 3.65935
R18331 gnd.n19 gnd.n18 3.60163
R18332 gnd.n4202 gnd.t279 3.50571
R18333 gnd.n6469 gnd.t217 3.50571
R18334 gnd.t194 gnd.n1899 3.50571
R18335 gnd.n4962 gnd.t356 3.50571
R18336 gnd.t224 gnd.n1452 3.50571
R18337 gnd.n7724 gnd.t203 3.50571
R18338 gnd.n3672 gnd.n3653 3.49141
R18339 gnd.n3640 gnd.n3621 3.49141
R18340 gnd.n3608 gnd.n3589 3.49141
R18341 gnd.n3577 gnd.n3558 3.49141
R18342 gnd.n3545 gnd.n3526 3.49141
R18343 gnd.n3513 gnd.n3494 3.49141
R18344 gnd.n3481 gnd.n3462 3.49141
R18345 gnd.n3450 gnd.n3431 3.49141
R18346 gnd.n5663 gnd.n1928 3.18706
R18347 gnd.n5430 gnd.n4760 3.18706
R18348 gnd.n5393 gnd.n4795 3.18706
R18349 gnd.n5759 gnd.n1842 3.18706
R18350 gnd.n5799 gnd.n1806 3.18706
R18351 gnd.n5313 gnd.n5312 3.18706
R18352 gnd.n5276 gnd.n4914 3.18706
R18353 gnd.n5895 gnd.n1717 3.18706
R18354 gnd.n5935 gnd.n1680 3.18706
R18355 gnd.n4990 gnd.t260 3.18706
R18356 gnd.n5196 gnd.n1653 3.18706
R18357 gnd.n2710 gnd.t122 2.8684
R18358 gnd.n5711 gnd.t84 2.8684
R18359 gnd.t0 gnd.n1703 2.8684
R18360 gnd.n2605 gnd.t43 2.82907
R18361 gnd.n2605 gnd.t91 2.82907
R18362 gnd.n2607 gnd.t178 2.82907
R18363 gnd.n2607 gnd.t69 2.82907
R18364 gnd.n2609 gnd.t191 2.82907
R18365 gnd.n2609 gnd.t316 2.82907
R18366 gnd.n2611 gnd.t93 2.82907
R18367 gnd.n2611 gnd.t41 2.82907
R18368 gnd.n2613 gnd.t47 2.82907
R18369 gnd.n2613 gnd.t329 2.82907
R18370 gnd.n2615 gnd.t121 2.82907
R18371 gnd.n2615 gnd.t12 2.82907
R18372 gnd.n2617 gnd.t190 2.82907
R18373 gnd.n2617 gnd.t155 2.82907
R18374 gnd.n2619 gnd.t71 2.82907
R18375 gnd.n2619 gnd.t23 2.82907
R18376 gnd.n2621 gnd.t157 2.82907
R18377 gnd.n2621 gnd.t348 2.82907
R18378 gnd.n2566 gnd.t182 2.82907
R18379 gnd.n2566 gnd.t136 2.82907
R18380 gnd.n2568 gnd.t35 2.82907
R18381 gnd.n2568 gnd.t74 2.82907
R18382 gnd.n2570 gnd.t354 2.82907
R18383 gnd.n2570 gnd.t98 2.82907
R18384 gnd.n2572 gnd.t137 2.82907
R18385 gnd.n2572 gnd.t144 2.82907
R18386 gnd.n2574 gnd.t90 2.82907
R18387 gnd.n2574 gnd.t87 2.82907
R18388 gnd.n2576 gnd.t168 2.82907
R18389 gnd.n2576 gnd.t104 2.82907
R18390 gnd.n2578 gnd.t187 2.82907
R18391 gnd.n2578 gnd.t101 2.82907
R18392 gnd.n2580 gnd.t172 2.82907
R18393 gnd.n2580 gnd.t143 2.82907
R18394 gnd.n2582 gnd.t185 2.82907
R18395 gnd.n2582 gnd.t53 2.82907
R18396 gnd.n2585 gnd.t176 2.82907
R18397 gnd.n2585 gnd.t89 2.82907
R18398 gnd.n2587 gnd.t134 2.82907
R18399 gnd.n2587 gnd.t55 2.82907
R18400 gnd.n2589 gnd.t150 2.82907
R18401 gnd.n2589 gnd.t353 2.82907
R18402 gnd.n2591 gnd.t50 2.82907
R18403 gnd.n2591 gnd.t73 2.82907
R18404 gnd.n2593 gnd.t37 2.82907
R18405 gnd.n2593 gnd.t177 2.82907
R18406 gnd.n2595 gnd.t103 2.82907
R18407 gnd.n2595 gnd.t99 2.82907
R18408 gnd.n2597 gnd.t341 2.82907
R18409 gnd.n2597 gnd.t181 2.82907
R18410 gnd.n2599 gnd.t72 2.82907
R18411 gnd.n2599 gnd.t64 2.82907
R18412 gnd.n2601 gnd.t345 2.82907
R18413 gnd.n2601 gnd.t63 2.82907
R18414 gnd.n75 gnd.t318 2.82907
R18415 gnd.n75 gnd.t324 2.82907
R18416 gnd.n73 gnd.t110 2.82907
R18417 gnd.n73 gnd.t76 2.82907
R18418 gnd.n71 gnd.t189 2.82907
R18419 gnd.n71 gnd.t315 2.82907
R18420 gnd.n69 gnd.t108 2.82907
R18421 gnd.n69 gnd.t193 2.82907
R18422 gnd.n67 gnd.t325 2.82907
R18423 gnd.n67 gnd.t355 2.82907
R18424 gnd.n65 gnd.t326 2.82907
R18425 gnd.n65 gnd.t317 2.82907
R18426 gnd.n63 gnd.t328 2.82907
R18427 gnd.n63 gnd.t153 2.82907
R18428 gnd.n61 gnd.t114 2.82907
R18429 gnd.n61 gnd.t92 2.82907
R18430 gnd.n59 gnd.t154 2.82907
R18431 gnd.n59 gnd.t48 2.82907
R18432 gnd.n36 gnd.t21 2.82907
R18433 gnd.n36 gnd.t120 2.82907
R18434 gnd.n34 gnd.t184 2.82907
R18435 gnd.n34 gnd.t68 2.82907
R18436 gnd.n32 gnd.t352 2.82907
R18437 gnd.n32 gnd.t146 2.82907
R18438 gnd.n30 gnd.t342 2.82907
R18439 gnd.n30 gnd.t346 2.82907
R18440 gnd.n28 gnd.t351 2.82907
R18441 gnd.n28 gnd.t171 2.82907
R18442 gnd.n26 gnd.t39 2.82907
R18443 gnd.n26 gnd.t323 2.82907
R18444 gnd.n24 gnd.t106 2.82907
R18445 gnd.n24 gnd.t118 2.82907
R18446 gnd.n22 gnd.t183 2.82907
R18447 gnd.n22 gnd.t75 2.82907
R18448 gnd.n20 gnd.t322 2.82907
R18449 gnd.n20 gnd.t8 2.82907
R18450 gnd.n55 gnd.t135 2.82907
R18451 gnd.n55 gnd.t142 2.82907
R18452 gnd.n53 gnd.t169 2.82907
R18453 gnd.n53 gnd.t138 2.82907
R18454 gnd.n51 gnd.t360 2.82907
R18455 gnd.n51 gnd.t66 2.82907
R18456 gnd.n49 gnd.t139 2.82907
R18457 gnd.n49 gnd.t321 2.82907
R18458 gnd.n47 gnd.t80 2.82907
R18459 gnd.n47 gnd.t148 2.82907
R18460 gnd.n45 gnd.t145 2.82907
R18461 gnd.n45 gnd.t19 2.82907
R18462 gnd.n43 gnd.t128 2.82907
R18463 gnd.n43 gnd.t141 2.82907
R18464 gnd.n41 gnd.t344 2.82907
R18465 gnd.n41 gnd.t57 2.82907
R18466 gnd.n39 gnd.t82 2.82907
R18467 gnd.n39 gnd.t51 2.82907
R18468 gnd.n3669 gnd.n3668 2.71565
R18469 gnd.n3637 gnd.n3636 2.71565
R18470 gnd.n3605 gnd.n3604 2.71565
R18471 gnd.n3574 gnd.n3573 2.71565
R18472 gnd.n3542 gnd.n3541 2.71565
R18473 gnd.n3510 gnd.n3509 2.71565
R18474 gnd.n3478 gnd.n3477 2.71565
R18475 gnd.n3447 gnd.n3446 2.71565
R18476 gnd.n4748 gnd.t228 2.54975
R18477 gnd.n5380 gnd.t196 2.54975
R18478 gnd.n5364 gnd.t77 2.54975
R18479 gnd.t32 gnd.n1745 2.54975
R18480 gnd.t4 gnd.n1733 2.54975
R18481 gnd.n3204 gnd.n2626 2.27742
R18482 gnd.n3204 gnd.n2565 2.27742
R18483 gnd.n3204 gnd.n2564 2.27742
R18484 gnd.n3204 gnd.n2563 2.27742
R18485 gnd.n7556 gnd.n7555 2.27742
R18486 gnd.n7556 gnd.n308 2.27742
R18487 gnd.n7556 gnd.n307 2.27742
R18488 gnd.n7556 gnd.n306 2.27742
R18489 gnd.n7556 gnd.n305 2.27742
R18490 gnd.n4303 gnd.n966 2.27742
R18491 gnd.n2214 gnd.n966 2.27742
R18492 gnd.n4320 gnd.n966 2.27742
R18493 gnd.n2188 gnd.n966 2.27742
R18494 gnd.n4347 gnd.n966 2.27742
R18495 gnd.n3058 gnd.t304 2.23109
R18496 gnd.n2681 gnd.t45 2.23109
R18497 gnd.n4376 gnd.t149 2.23109
R18498 gnd.t117 gnd.n367 2.23109
R18499 gnd.n3665 gnd.n3655 1.93989
R18500 gnd.n3633 gnd.n3623 1.93989
R18501 gnd.n3601 gnd.n3591 1.93989
R18502 gnd.n3570 gnd.n3560 1.93989
R18503 gnd.n3538 gnd.n3528 1.93989
R18504 gnd.n3506 gnd.n3496 1.93989
R18505 gnd.n3474 gnd.n3464 1.93989
R18506 gnd.n3443 gnd.n3433 1.93989
R18507 gnd.n5423 gnd.n5422 1.91244
R18508 gnd.n5400 gnd.n4787 1.91244
R18509 gnd.n5791 gnd.n1813 1.91244
R18510 gnd.n5305 gnd.n4887 1.91244
R18511 gnd.n5903 gnd.n1710 1.91244
R18512 gnd.n5927 gnd.n1688 1.91244
R18513 gnd.n5203 gnd.t200 1.91244
R18514 gnd.t179 gnd.n3069 1.59378
R18515 gnd.n3248 gnd.t334 1.59378
R18516 gnd.n2498 gnd.t125 1.59378
R18517 gnd.n4242 gnd.t52 1.59378
R18518 gnd.n4425 gnd.t54 1.59378
R18519 gnd.n6499 gnd.t42 1.59378
R18520 gnd.n5767 gnd.t2 1.59378
R18521 gnd.t158 gnd.n4907 1.59378
R18522 gnd.n1398 gnd.t7 1.59378
R18523 gnd.t113 gnd.n6180 1.59378
R18524 gnd.n7616 gnd.t20 1.59378
R18525 gnd.t207 gnd.n1920 1.27512
R18526 gnd.n5735 gnd.t116 1.27512
R18527 gnd.t96 gnd.n4935 1.27512
R18528 gnd.n2911 gnd.n2903 1.16414
R18529 gnd.n3727 gnd.n2400 1.16414
R18530 gnd.n3664 gnd.n3657 1.16414
R18531 gnd.n3632 gnd.n3625 1.16414
R18532 gnd.n3600 gnd.n3593 1.16414
R18533 gnd.n3569 gnd.n3562 1.16414
R18534 gnd.n3537 gnd.n3530 1.16414
R18535 gnd.n3505 gnd.n3498 1.16414
R18536 gnd.n3473 gnd.n3466 1.16414
R18537 gnd.n3442 gnd.n3435 1.16414
R18538 gnd.n6262 gnd.n6261 0.970197
R18539 gnd.n5527 gnd.n2097 0.970197
R18540 gnd.n3648 gnd.n3616 0.962709
R18541 gnd.n3680 gnd.n3648 0.962709
R18542 gnd.n3521 gnd.n3489 0.962709
R18543 gnd.n3553 gnd.n3521 0.962709
R18544 gnd.n3157 gnd.t166 0.956468
R18545 gnd.n3322 gnd.t336 0.956468
R18546 gnd.n4274 gnd.t186 0.956468
R18547 gnd.n6523 gnd.t97 0.956468
R18548 gnd.n4510 gnd.t111 0.956468
R18549 gnd.n5445 gnd.t349 0.956468
R18550 gnd.n5205 gnd.t362 0.956468
R18551 gnd.t9 gnd.n1424 0.956468
R18552 gnd.n7384 gnd.t105 0.956468
R18553 gnd.n7584 gnd.t65 0.956468
R18554 gnd.n2616 gnd.n2614 0.773756
R18555 gnd.n70 gnd.n68 0.773756
R18556 gnd.n2623 gnd.n2622 0.773756
R18557 gnd.n2622 gnd.n2620 0.773756
R18558 gnd.n2620 gnd.n2618 0.773756
R18559 gnd.n2618 gnd.n2616 0.773756
R18560 gnd.n2614 gnd.n2612 0.773756
R18561 gnd.n2612 gnd.n2610 0.773756
R18562 gnd.n2610 gnd.n2608 0.773756
R18563 gnd.n2608 gnd.n2606 0.773756
R18564 gnd.n62 gnd.n60 0.773756
R18565 gnd.n64 gnd.n62 0.773756
R18566 gnd.n66 gnd.n64 0.773756
R18567 gnd.n68 gnd.n66 0.773756
R18568 gnd.n72 gnd.n70 0.773756
R18569 gnd.n74 gnd.n72 0.773756
R18570 gnd.n76 gnd.n74 0.773756
R18571 gnd.n77 gnd.n76 0.773756
R18572 gnd gnd.n0 0.70738
R18573 gnd.n2 gnd.n1 0.672012
R18574 gnd.n3 gnd.n2 0.672012
R18575 gnd.n4 gnd.n3 0.672012
R18576 gnd.n5 gnd.n4 0.672012
R18577 gnd.n6 gnd.n5 0.672012
R18578 gnd.n7 gnd.n6 0.672012
R18579 gnd.n8 gnd.n7 0.672012
R18580 gnd.n9 gnd.n8 0.672012
R18581 gnd.n11 gnd.n10 0.672012
R18582 gnd.n12 gnd.n11 0.672012
R18583 gnd.n13 gnd.n12 0.672012
R18584 gnd.n14 gnd.n13 0.672012
R18585 gnd.n15 gnd.n14 0.672012
R18586 gnd.n16 gnd.n15 0.672012
R18587 gnd.n17 gnd.n16 0.672012
R18588 gnd.n18 gnd.n17 0.672012
R18589 gnd.t235 gnd.n1913 0.637812
R18590 gnd.n5415 gnd.n4773 0.637812
R18591 gnd.n5408 gnd.n5407 0.637812
R18592 gnd.n5407 gnd.t197 0.637812
R18593 gnd.n5775 gnd.n1827 0.637812
R18594 gnd.n5783 gnd.n1821 0.637812
R18595 gnd.n5343 gnd.t83 0.637812
R18596 gnd.t29 gnd.n1777 0.637812
R18597 gnd.n5298 gnd.n5297 0.637812
R18598 gnd.n5290 gnd.n4900 0.637812
R18599 gnd.t131 gnd.n1701 0.637812
R18600 gnd.n5911 gnd.n1701 0.637812
R18601 gnd.n5919 gnd.n1695 0.637812
R18602 gnd.n4990 gnd.t231 0.637812
R18603 gnd.n7859 gnd.n7858 0.637193
R18604 gnd.n2584 gnd.n2583 0.573776
R18605 gnd.n2583 gnd.n2581 0.573776
R18606 gnd.n2581 gnd.n2579 0.573776
R18607 gnd.n2579 gnd.n2577 0.573776
R18608 gnd.n2577 gnd.n2575 0.573776
R18609 gnd.n2575 gnd.n2573 0.573776
R18610 gnd.n2573 gnd.n2571 0.573776
R18611 gnd.n2571 gnd.n2569 0.573776
R18612 gnd.n2569 gnd.n2567 0.573776
R18613 gnd.n2603 gnd.n2602 0.573776
R18614 gnd.n2602 gnd.n2600 0.573776
R18615 gnd.n2600 gnd.n2598 0.573776
R18616 gnd.n2598 gnd.n2596 0.573776
R18617 gnd.n2596 gnd.n2594 0.573776
R18618 gnd.n2594 gnd.n2592 0.573776
R18619 gnd.n2592 gnd.n2590 0.573776
R18620 gnd.n2590 gnd.n2588 0.573776
R18621 gnd.n2588 gnd.n2586 0.573776
R18622 gnd.n23 gnd.n21 0.573776
R18623 gnd.n25 gnd.n23 0.573776
R18624 gnd.n27 gnd.n25 0.573776
R18625 gnd.n29 gnd.n27 0.573776
R18626 gnd.n31 gnd.n29 0.573776
R18627 gnd.n33 gnd.n31 0.573776
R18628 gnd.n35 gnd.n33 0.573776
R18629 gnd.n37 gnd.n35 0.573776
R18630 gnd.n38 gnd.n37 0.573776
R18631 gnd.n42 gnd.n40 0.573776
R18632 gnd.n44 gnd.n42 0.573776
R18633 gnd.n46 gnd.n44 0.573776
R18634 gnd.n48 gnd.n46 0.573776
R18635 gnd.n50 gnd.n48 0.573776
R18636 gnd.n52 gnd.n50 0.573776
R18637 gnd.n54 gnd.n52 0.573776
R18638 gnd.n56 gnd.n54 0.573776
R18639 gnd.n57 gnd.n56 0.573776
R18640 gnd.n7556 gnd.n304 0.5435
R18641 gnd.n6546 gnd.n966 0.5435
R18642 gnd.n3384 gnd.n2404 0.486781
R18643 gnd.n1518 gnd.n1242 0.486781
R18644 gnd.n2960 gnd.n2959 0.48678
R18645 gnd.n6458 gnd.n6457 0.485256
R18646 gnd.n3701 gnd.n2358 0.480683
R18647 gnd.n3044 gnd.n3043 0.480683
R18648 gnd.n6718 gnd.n6717 0.480683
R18649 gnd.n7139 gnd.n7138 0.480683
R18650 gnd.n3878 gnd.n3877 0.477634
R18651 gnd.n4197 gnd.n2332 0.477634
R18652 gnd.n7707 gnd.n7706 0.477634
R18653 gnd.n7809 gnd.n7808 0.477634
R18654 gnd.n7801 gnd.n7800 0.465439
R18655 gnd.n7730 gnd.n7729 0.465439
R18656 gnd.n6222 gnd.n1333 0.465439
R18657 gnd.n6047 gnd.n1289 0.465439
R18658 gnd.n2081 gnd.n1107 0.465439
R18659 gnd.n4573 gnd.n4572 0.465439
R18660 gnd.n4116 gnd.n4111 0.465439
R18661 gnd.n4191 gnd.n4190 0.465439
R18662 gnd.n6018 gnd.n6017 0.451719
R18663 gnd.n5611 gnd.n5610 0.451719
R18664 gnd.n4553 gnd.n4545 0.388379
R18665 gnd.n3661 gnd.n3660 0.388379
R18666 gnd.n3629 gnd.n3628 0.388379
R18667 gnd.n3597 gnd.n3596 0.388379
R18668 gnd.n3566 gnd.n3565 0.388379
R18669 gnd.n3534 gnd.n3533 0.388379
R18670 gnd.n3502 gnd.n3501 0.388379
R18671 gnd.n3470 gnd.n3469 0.388379
R18672 gnd.n3439 gnd.n3438 0.388379
R18673 gnd.n7770 gnd.n7769 0.388379
R18674 gnd.n4002 gnd.n3998 0.388379
R18675 gnd.n6032 gnd.n6031 0.388379
R18676 gnd.n6460 gnd.n6459 0.378829
R18677 gnd.n6215 gnd.n1342 0.377553
R18678 gnd.n7859 gnd.n19 0.374463
R18679 gnd gnd.n7859 0.367492
R18680 gnd.n2460 gnd.t15 0.319156
R18681 gnd.n4307 gnd.t11 0.319156
R18682 gnd.n4350 gnd.t49 0.319156
R18683 gnd.n5363 gnd.t2 0.319156
R18684 gnd.t5 gnd.t337 0.319156
R18685 gnd.t30 gnd.t313 0.319156
R18686 gnd.n5283 gnd.t158 0.319156
R18687 gnd.n7444 gnd.t18 0.319156
R18688 gnd.n7536 gnd.t107 0.319156
R18689 gnd.n2878 gnd.n2856 0.311721
R18690 gnd.n7350 gnd.n304 0.282512
R18691 gnd.n6547 gnd.n6546 0.282512
R18692 gnd.n3772 gnd.n3771 0.268793
R18693 gnd.n4564 gnd.n4563 0.247451
R18694 gnd.n6042 gnd.n6041 0.247451
R18695 gnd.n3771 gnd.n3770 0.241354
R18696 gnd.n1307 gnd.n1304 0.229039
R18697 gnd.n1310 gnd.n1307 0.229039
R18698 gnd.n4616 gnd.n2096 0.229039
R18699 gnd.n4616 gnd.n4615 0.229039
R18700 gnd.n2625 gnd.n0 0.210825
R18701 gnd.n3032 gnd.n2831 0.206293
R18702 gnd.n420 gnd.n304 0.198671
R18703 gnd.n6546 gnd.n6545 0.198671
R18704 gnd.n3678 gnd.n3650 0.155672
R18705 gnd.n3671 gnd.n3650 0.155672
R18706 gnd.n3671 gnd.n3670 0.155672
R18707 gnd.n3670 gnd.n3654 0.155672
R18708 gnd.n3663 gnd.n3654 0.155672
R18709 gnd.n3663 gnd.n3662 0.155672
R18710 gnd.n3646 gnd.n3618 0.155672
R18711 gnd.n3639 gnd.n3618 0.155672
R18712 gnd.n3639 gnd.n3638 0.155672
R18713 gnd.n3638 gnd.n3622 0.155672
R18714 gnd.n3631 gnd.n3622 0.155672
R18715 gnd.n3631 gnd.n3630 0.155672
R18716 gnd.n3614 gnd.n3586 0.155672
R18717 gnd.n3607 gnd.n3586 0.155672
R18718 gnd.n3607 gnd.n3606 0.155672
R18719 gnd.n3606 gnd.n3590 0.155672
R18720 gnd.n3599 gnd.n3590 0.155672
R18721 gnd.n3599 gnd.n3598 0.155672
R18722 gnd.n3583 gnd.n3555 0.155672
R18723 gnd.n3576 gnd.n3555 0.155672
R18724 gnd.n3576 gnd.n3575 0.155672
R18725 gnd.n3575 gnd.n3559 0.155672
R18726 gnd.n3568 gnd.n3559 0.155672
R18727 gnd.n3568 gnd.n3567 0.155672
R18728 gnd.n3551 gnd.n3523 0.155672
R18729 gnd.n3544 gnd.n3523 0.155672
R18730 gnd.n3544 gnd.n3543 0.155672
R18731 gnd.n3543 gnd.n3527 0.155672
R18732 gnd.n3536 gnd.n3527 0.155672
R18733 gnd.n3536 gnd.n3535 0.155672
R18734 gnd.n3519 gnd.n3491 0.155672
R18735 gnd.n3512 gnd.n3491 0.155672
R18736 gnd.n3512 gnd.n3511 0.155672
R18737 gnd.n3511 gnd.n3495 0.155672
R18738 gnd.n3504 gnd.n3495 0.155672
R18739 gnd.n3504 gnd.n3503 0.155672
R18740 gnd.n3487 gnd.n3459 0.155672
R18741 gnd.n3480 gnd.n3459 0.155672
R18742 gnd.n3480 gnd.n3479 0.155672
R18743 gnd.n3479 gnd.n3463 0.155672
R18744 gnd.n3472 gnd.n3463 0.155672
R18745 gnd.n3472 gnd.n3471 0.155672
R18746 gnd.n3456 gnd.n3428 0.155672
R18747 gnd.n3449 gnd.n3428 0.155672
R18748 gnd.n3449 gnd.n3448 0.155672
R18749 gnd.n3448 gnd.n3432 0.155672
R18750 gnd.n3441 gnd.n3432 0.155672
R18751 gnd.n3441 gnd.n3440 0.155672
R18752 gnd.n3803 gnd.n2358 0.152939
R18753 gnd.n3803 gnd.n3802 0.152939
R18754 gnd.n3802 gnd.n3801 0.152939
R18755 gnd.n3801 gnd.n2360 0.152939
R18756 gnd.n2361 gnd.n2360 0.152939
R18757 gnd.n2362 gnd.n2361 0.152939
R18758 gnd.n2363 gnd.n2362 0.152939
R18759 gnd.n2364 gnd.n2363 0.152939
R18760 gnd.n2365 gnd.n2364 0.152939
R18761 gnd.n2366 gnd.n2365 0.152939
R18762 gnd.n2367 gnd.n2366 0.152939
R18763 gnd.n2368 gnd.n2367 0.152939
R18764 gnd.n2369 gnd.n2368 0.152939
R18765 gnd.n2370 gnd.n2369 0.152939
R18766 gnd.n3773 gnd.n2370 0.152939
R18767 gnd.n3773 gnd.n3772 0.152939
R18768 gnd.n3045 gnd.n3044 0.152939
R18769 gnd.n3045 gnd.n2749 0.152939
R18770 gnd.n3073 gnd.n2749 0.152939
R18771 gnd.n3074 gnd.n3073 0.152939
R18772 gnd.n3075 gnd.n3074 0.152939
R18773 gnd.n3076 gnd.n3075 0.152939
R18774 gnd.n3076 gnd.n2721 0.152939
R18775 gnd.n3103 gnd.n2721 0.152939
R18776 gnd.n3104 gnd.n3103 0.152939
R18777 gnd.n3105 gnd.n3104 0.152939
R18778 gnd.n3105 gnd.n2699 0.152939
R18779 gnd.n3134 gnd.n2699 0.152939
R18780 gnd.n3135 gnd.n3134 0.152939
R18781 gnd.n3136 gnd.n3135 0.152939
R18782 gnd.n3137 gnd.n3136 0.152939
R18783 gnd.n3139 gnd.n3137 0.152939
R18784 gnd.n3139 gnd.n3138 0.152939
R18785 gnd.n3138 gnd.n2648 0.152939
R18786 gnd.n2649 gnd.n2648 0.152939
R18787 gnd.n2650 gnd.n2649 0.152939
R18788 gnd.n2669 gnd.n2650 0.152939
R18789 gnd.n2670 gnd.n2669 0.152939
R18790 gnd.n2670 gnd.n2556 0.152939
R18791 gnd.n3229 gnd.n2556 0.152939
R18792 gnd.n3230 gnd.n3229 0.152939
R18793 gnd.n3231 gnd.n3230 0.152939
R18794 gnd.n3232 gnd.n3231 0.152939
R18795 gnd.n3232 gnd.n2529 0.152939
R18796 gnd.n3269 gnd.n2529 0.152939
R18797 gnd.n3270 gnd.n3269 0.152939
R18798 gnd.n3271 gnd.n3270 0.152939
R18799 gnd.n3272 gnd.n3271 0.152939
R18800 gnd.n3272 gnd.n2502 0.152939
R18801 gnd.n3314 gnd.n2502 0.152939
R18802 gnd.n3315 gnd.n3314 0.152939
R18803 gnd.n3316 gnd.n3315 0.152939
R18804 gnd.n3317 gnd.n3316 0.152939
R18805 gnd.n3317 gnd.n2474 0.152939
R18806 gnd.n3354 gnd.n2474 0.152939
R18807 gnd.n3355 gnd.n3354 0.152939
R18808 gnd.n3356 gnd.n3355 0.152939
R18809 gnd.n3357 gnd.n3356 0.152939
R18810 gnd.n3357 gnd.n2447 0.152939
R18811 gnd.n3403 gnd.n2447 0.152939
R18812 gnd.n3404 gnd.n3403 0.152939
R18813 gnd.n3405 gnd.n3404 0.152939
R18814 gnd.n3406 gnd.n3405 0.152939
R18815 gnd.n3406 gnd.n2420 0.152939
R18816 gnd.n3697 gnd.n2420 0.152939
R18817 gnd.n3698 gnd.n3697 0.152939
R18818 gnd.n3699 gnd.n3698 0.152939
R18819 gnd.n3700 gnd.n3699 0.152939
R18820 gnd.n3701 gnd.n3700 0.152939
R18821 gnd.n3043 gnd.n2773 0.152939
R18822 gnd.n2794 gnd.n2773 0.152939
R18823 gnd.n2795 gnd.n2794 0.152939
R18824 gnd.n2801 gnd.n2795 0.152939
R18825 gnd.n2802 gnd.n2801 0.152939
R18826 gnd.n2803 gnd.n2802 0.152939
R18827 gnd.n2803 gnd.n2792 0.152939
R18828 gnd.n2811 gnd.n2792 0.152939
R18829 gnd.n2812 gnd.n2811 0.152939
R18830 gnd.n2813 gnd.n2812 0.152939
R18831 gnd.n2813 gnd.n2790 0.152939
R18832 gnd.n2821 gnd.n2790 0.152939
R18833 gnd.n2822 gnd.n2821 0.152939
R18834 gnd.n2823 gnd.n2822 0.152939
R18835 gnd.n2823 gnd.n2788 0.152939
R18836 gnd.n2831 gnd.n2788 0.152939
R18837 gnd.n3770 gnd.n2375 0.152939
R18838 gnd.n2377 gnd.n2375 0.152939
R18839 gnd.n2378 gnd.n2377 0.152939
R18840 gnd.n2379 gnd.n2378 0.152939
R18841 gnd.n2380 gnd.n2379 0.152939
R18842 gnd.n2381 gnd.n2380 0.152939
R18843 gnd.n2382 gnd.n2381 0.152939
R18844 gnd.n2383 gnd.n2382 0.152939
R18845 gnd.n2384 gnd.n2383 0.152939
R18846 gnd.n2385 gnd.n2384 0.152939
R18847 gnd.n2386 gnd.n2385 0.152939
R18848 gnd.n2387 gnd.n2386 0.152939
R18849 gnd.n2388 gnd.n2387 0.152939
R18850 gnd.n2389 gnd.n2388 0.152939
R18851 gnd.n2390 gnd.n2389 0.152939
R18852 gnd.n2391 gnd.n2390 0.152939
R18853 gnd.n2392 gnd.n2391 0.152939
R18854 gnd.n2393 gnd.n2392 0.152939
R18855 gnd.n2394 gnd.n2393 0.152939
R18856 gnd.n2395 gnd.n2394 0.152939
R18857 gnd.n2396 gnd.n2395 0.152939
R18858 gnd.n2397 gnd.n2396 0.152939
R18859 gnd.n2401 gnd.n2397 0.152939
R18860 gnd.n2402 gnd.n2401 0.152939
R18861 gnd.n2403 gnd.n2402 0.152939
R18862 gnd.n2404 gnd.n2403 0.152939
R18863 gnd.n3206 gnd.n3205 0.152939
R18864 gnd.n3207 gnd.n3206 0.152939
R18865 gnd.n3208 gnd.n3207 0.152939
R18866 gnd.n3209 gnd.n3208 0.152939
R18867 gnd.n3210 gnd.n3209 0.152939
R18868 gnd.n3211 gnd.n3210 0.152939
R18869 gnd.n3211 gnd.n2510 0.152939
R18870 gnd.n3290 gnd.n2510 0.152939
R18871 gnd.n3291 gnd.n3290 0.152939
R18872 gnd.n3292 gnd.n3291 0.152939
R18873 gnd.n3293 gnd.n3292 0.152939
R18874 gnd.n3294 gnd.n3293 0.152939
R18875 gnd.n3295 gnd.n3294 0.152939
R18876 gnd.n3296 gnd.n3295 0.152939
R18877 gnd.n3297 gnd.n3296 0.152939
R18878 gnd.n3298 gnd.n3297 0.152939
R18879 gnd.n3298 gnd.n2454 0.152939
R18880 gnd.n3375 gnd.n2454 0.152939
R18881 gnd.n3376 gnd.n3375 0.152939
R18882 gnd.n3377 gnd.n3376 0.152939
R18883 gnd.n3378 gnd.n3377 0.152939
R18884 gnd.n3379 gnd.n3378 0.152939
R18885 gnd.n3380 gnd.n3379 0.152939
R18886 gnd.n3381 gnd.n3380 0.152939
R18887 gnd.n3382 gnd.n3381 0.152939
R18888 gnd.n3383 gnd.n3382 0.152939
R18889 gnd.n3385 gnd.n3383 0.152939
R18890 gnd.n3385 gnd.n3384 0.152939
R18891 gnd.n2961 gnd.n2960 0.152939
R18892 gnd.n2961 gnd.n2851 0.152939
R18893 gnd.n2976 gnd.n2851 0.152939
R18894 gnd.n2977 gnd.n2976 0.152939
R18895 gnd.n2978 gnd.n2977 0.152939
R18896 gnd.n2978 gnd.n2839 0.152939
R18897 gnd.n2992 gnd.n2839 0.152939
R18898 gnd.n2993 gnd.n2992 0.152939
R18899 gnd.n2994 gnd.n2993 0.152939
R18900 gnd.n2995 gnd.n2994 0.152939
R18901 gnd.n2996 gnd.n2995 0.152939
R18902 gnd.n2997 gnd.n2996 0.152939
R18903 gnd.n2998 gnd.n2997 0.152939
R18904 gnd.n2999 gnd.n2998 0.152939
R18905 gnd.n3000 gnd.n2999 0.152939
R18906 gnd.n3001 gnd.n3000 0.152939
R18907 gnd.n3002 gnd.n3001 0.152939
R18908 gnd.n3003 gnd.n3002 0.152939
R18909 gnd.n3004 gnd.n3003 0.152939
R18910 gnd.n3005 gnd.n3004 0.152939
R18911 gnd.n3006 gnd.n3005 0.152939
R18912 gnd.n3006 gnd.n2705 0.152939
R18913 gnd.n3123 gnd.n2705 0.152939
R18914 gnd.n3124 gnd.n3123 0.152939
R18915 gnd.n3125 gnd.n3124 0.152939
R18916 gnd.n3126 gnd.n3125 0.152939
R18917 gnd.n3126 gnd.n2627 0.152939
R18918 gnd.n3203 gnd.n2627 0.152939
R18919 gnd.n2879 gnd.n2878 0.152939
R18920 gnd.n2880 gnd.n2879 0.152939
R18921 gnd.n2881 gnd.n2880 0.152939
R18922 gnd.n2882 gnd.n2881 0.152939
R18923 gnd.n2883 gnd.n2882 0.152939
R18924 gnd.n2884 gnd.n2883 0.152939
R18925 gnd.n2885 gnd.n2884 0.152939
R18926 gnd.n2886 gnd.n2885 0.152939
R18927 gnd.n2887 gnd.n2886 0.152939
R18928 gnd.n2888 gnd.n2887 0.152939
R18929 gnd.n2889 gnd.n2888 0.152939
R18930 gnd.n2890 gnd.n2889 0.152939
R18931 gnd.n2891 gnd.n2890 0.152939
R18932 gnd.n2892 gnd.n2891 0.152939
R18933 gnd.n2893 gnd.n2892 0.152939
R18934 gnd.n2894 gnd.n2893 0.152939
R18935 gnd.n2895 gnd.n2894 0.152939
R18936 gnd.n2896 gnd.n2895 0.152939
R18937 gnd.n2897 gnd.n2896 0.152939
R18938 gnd.n2898 gnd.n2897 0.152939
R18939 gnd.n2899 gnd.n2898 0.152939
R18940 gnd.n2900 gnd.n2899 0.152939
R18941 gnd.n2904 gnd.n2900 0.152939
R18942 gnd.n2905 gnd.n2904 0.152939
R18943 gnd.n2905 gnd.n2862 0.152939
R18944 gnd.n2959 gnd.n2862 0.152939
R18945 gnd.n6718 gnd.n794 0.152939
R18946 gnd.n6726 gnd.n794 0.152939
R18947 gnd.n6727 gnd.n6726 0.152939
R18948 gnd.n6728 gnd.n6727 0.152939
R18949 gnd.n6728 gnd.n788 0.152939
R18950 gnd.n6736 gnd.n788 0.152939
R18951 gnd.n6737 gnd.n6736 0.152939
R18952 gnd.n6738 gnd.n6737 0.152939
R18953 gnd.n6738 gnd.n782 0.152939
R18954 gnd.n6746 gnd.n782 0.152939
R18955 gnd.n6747 gnd.n6746 0.152939
R18956 gnd.n6748 gnd.n6747 0.152939
R18957 gnd.n6748 gnd.n776 0.152939
R18958 gnd.n6756 gnd.n776 0.152939
R18959 gnd.n6757 gnd.n6756 0.152939
R18960 gnd.n6758 gnd.n6757 0.152939
R18961 gnd.n6758 gnd.n770 0.152939
R18962 gnd.n6766 gnd.n770 0.152939
R18963 gnd.n6767 gnd.n6766 0.152939
R18964 gnd.n6768 gnd.n6767 0.152939
R18965 gnd.n6768 gnd.n764 0.152939
R18966 gnd.n6776 gnd.n764 0.152939
R18967 gnd.n6777 gnd.n6776 0.152939
R18968 gnd.n6778 gnd.n6777 0.152939
R18969 gnd.n6778 gnd.n758 0.152939
R18970 gnd.n6786 gnd.n758 0.152939
R18971 gnd.n6787 gnd.n6786 0.152939
R18972 gnd.n6788 gnd.n6787 0.152939
R18973 gnd.n6788 gnd.n752 0.152939
R18974 gnd.n6796 gnd.n752 0.152939
R18975 gnd.n6797 gnd.n6796 0.152939
R18976 gnd.n6798 gnd.n6797 0.152939
R18977 gnd.n6798 gnd.n746 0.152939
R18978 gnd.n6806 gnd.n746 0.152939
R18979 gnd.n6807 gnd.n6806 0.152939
R18980 gnd.n6808 gnd.n6807 0.152939
R18981 gnd.n6808 gnd.n740 0.152939
R18982 gnd.n6816 gnd.n740 0.152939
R18983 gnd.n6817 gnd.n6816 0.152939
R18984 gnd.n6818 gnd.n6817 0.152939
R18985 gnd.n6818 gnd.n734 0.152939
R18986 gnd.n6826 gnd.n734 0.152939
R18987 gnd.n6827 gnd.n6826 0.152939
R18988 gnd.n6828 gnd.n6827 0.152939
R18989 gnd.n6828 gnd.n728 0.152939
R18990 gnd.n6836 gnd.n728 0.152939
R18991 gnd.n6837 gnd.n6836 0.152939
R18992 gnd.n6838 gnd.n6837 0.152939
R18993 gnd.n6838 gnd.n722 0.152939
R18994 gnd.n6846 gnd.n722 0.152939
R18995 gnd.n6847 gnd.n6846 0.152939
R18996 gnd.n6848 gnd.n6847 0.152939
R18997 gnd.n6848 gnd.n716 0.152939
R18998 gnd.n6856 gnd.n716 0.152939
R18999 gnd.n6857 gnd.n6856 0.152939
R19000 gnd.n6858 gnd.n6857 0.152939
R19001 gnd.n6858 gnd.n710 0.152939
R19002 gnd.n6866 gnd.n710 0.152939
R19003 gnd.n6867 gnd.n6866 0.152939
R19004 gnd.n6868 gnd.n6867 0.152939
R19005 gnd.n6868 gnd.n704 0.152939
R19006 gnd.n6876 gnd.n704 0.152939
R19007 gnd.n6877 gnd.n6876 0.152939
R19008 gnd.n6878 gnd.n6877 0.152939
R19009 gnd.n6878 gnd.n698 0.152939
R19010 gnd.n6886 gnd.n698 0.152939
R19011 gnd.n6887 gnd.n6886 0.152939
R19012 gnd.n6888 gnd.n6887 0.152939
R19013 gnd.n6888 gnd.n692 0.152939
R19014 gnd.n6896 gnd.n692 0.152939
R19015 gnd.n6897 gnd.n6896 0.152939
R19016 gnd.n6898 gnd.n6897 0.152939
R19017 gnd.n6898 gnd.n686 0.152939
R19018 gnd.n6906 gnd.n686 0.152939
R19019 gnd.n6907 gnd.n6906 0.152939
R19020 gnd.n6908 gnd.n6907 0.152939
R19021 gnd.n6908 gnd.n680 0.152939
R19022 gnd.n6916 gnd.n680 0.152939
R19023 gnd.n6917 gnd.n6916 0.152939
R19024 gnd.n6918 gnd.n6917 0.152939
R19025 gnd.n6918 gnd.n674 0.152939
R19026 gnd.n6926 gnd.n674 0.152939
R19027 gnd.n6927 gnd.n6926 0.152939
R19028 gnd.n6928 gnd.n6927 0.152939
R19029 gnd.n6928 gnd.n668 0.152939
R19030 gnd.n6936 gnd.n668 0.152939
R19031 gnd.n6937 gnd.n6936 0.152939
R19032 gnd.n6938 gnd.n6937 0.152939
R19033 gnd.n6938 gnd.n662 0.152939
R19034 gnd.n6946 gnd.n662 0.152939
R19035 gnd.n6947 gnd.n6946 0.152939
R19036 gnd.n6948 gnd.n6947 0.152939
R19037 gnd.n6948 gnd.n656 0.152939
R19038 gnd.n6956 gnd.n656 0.152939
R19039 gnd.n6957 gnd.n6956 0.152939
R19040 gnd.n6958 gnd.n6957 0.152939
R19041 gnd.n6958 gnd.n650 0.152939
R19042 gnd.n6966 gnd.n650 0.152939
R19043 gnd.n6967 gnd.n6966 0.152939
R19044 gnd.n6968 gnd.n6967 0.152939
R19045 gnd.n6968 gnd.n644 0.152939
R19046 gnd.n6976 gnd.n644 0.152939
R19047 gnd.n6977 gnd.n6976 0.152939
R19048 gnd.n6978 gnd.n6977 0.152939
R19049 gnd.n6978 gnd.n638 0.152939
R19050 gnd.n6986 gnd.n638 0.152939
R19051 gnd.n6987 gnd.n6986 0.152939
R19052 gnd.n6988 gnd.n6987 0.152939
R19053 gnd.n6988 gnd.n632 0.152939
R19054 gnd.n6996 gnd.n632 0.152939
R19055 gnd.n6997 gnd.n6996 0.152939
R19056 gnd.n6998 gnd.n6997 0.152939
R19057 gnd.n6998 gnd.n626 0.152939
R19058 gnd.n7006 gnd.n626 0.152939
R19059 gnd.n7007 gnd.n7006 0.152939
R19060 gnd.n7008 gnd.n7007 0.152939
R19061 gnd.n7008 gnd.n620 0.152939
R19062 gnd.n7016 gnd.n620 0.152939
R19063 gnd.n7017 gnd.n7016 0.152939
R19064 gnd.n7018 gnd.n7017 0.152939
R19065 gnd.n7018 gnd.n614 0.152939
R19066 gnd.n7026 gnd.n614 0.152939
R19067 gnd.n7027 gnd.n7026 0.152939
R19068 gnd.n7028 gnd.n7027 0.152939
R19069 gnd.n7028 gnd.n608 0.152939
R19070 gnd.n7036 gnd.n608 0.152939
R19071 gnd.n7037 gnd.n7036 0.152939
R19072 gnd.n7038 gnd.n7037 0.152939
R19073 gnd.n7038 gnd.n602 0.152939
R19074 gnd.n7046 gnd.n602 0.152939
R19075 gnd.n7047 gnd.n7046 0.152939
R19076 gnd.n7048 gnd.n7047 0.152939
R19077 gnd.n7048 gnd.n596 0.152939
R19078 gnd.n7056 gnd.n596 0.152939
R19079 gnd.n7057 gnd.n7056 0.152939
R19080 gnd.n7058 gnd.n7057 0.152939
R19081 gnd.n7058 gnd.n590 0.152939
R19082 gnd.n7066 gnd.n590 0.152939
R19083 gnd.n7067 gnd.n7066 0.152939
R19084 gnd.n7068 gnd.n7067 0.152939
R19085 gnd.n7068 gnd.n584 0.152939
R19086 gnd.n7076 gnd.n584 0.152939
R19087 gnd.n7077 gnd.n7076 0.152939
R19088 gnd.n7078 gnd.n7077 0.152939
R19089 gnd.n7078 gnd.n578 0.152939
R19090 gnd.n7086 gnd.n578 0.152939
R19091 gnd.n7087 gnd.n7086 0.152939
R19092 gnd.n7088 gnd.n7087 0.152939
R19093 gnd.n7088 gnd.n572 0.152939
R19094 gnd.n7096 gnd.n572 0.152939
R19095 gnd.n7097 gnd.n7096 0.152939
R19096 gnd.n7098 gnd.n7097 0.152939
R19097 gnd.n7098 gnd.n566 0.152939
R19098 gnd.n7106 gnd.n566 0.152939
R19099 gnd.n7107 gnd.n7106 0.152939
R19100 gnd.n7108 gnd.n7107 0.152939
R19101 gnd.n7108 gnd.n560 0.152939
R19102 gnd.n7116 gnd.n560 0.152939
R19103 gnd.n7117 gnd.n7116 0.152939
R19104 gnd.n7118 gnd.n7117 0.152939
R19105 gnd.n7118 gnd.n554 0.152939
R19106 gnd.n7126 gnd.n554 0.152939
R19107 gnd.n7127 gnd.n7126 0.152939
R19108 gnd.n7129 gnd.n7127 0.152939
R19109 gnd.n7129 gnd.n7128 0.152939
R19110 gnd.n7128 gnd.n548 0.152939
R19111 gnd.n7138 gnd.n548 0.152939
R19112 gnd.n7139 gnd.n543 0.152939
R19113 gnd.n7147 gnd.n543 0.152939
R19114 gnd.n7148 gnd.n7147 0.152939
R19115 gnd.n7149 gnd.n7148 0.152939
R19116 gnd.n7149 gnd.n537 0.152939
R19117 gnd.n7157 gnd.n537 0.152939
R19118 gnd.n7158 gnd.n7157 0.152939
R19119 gnd.n7159 gnd.n7158 0.152939
R19120 gnd.n7159 gnd.n531 0.152939
R19121 gnd.n7167 gnd.n531 0.152939
R19122 gnd.n7168 gnd.n7167 0.152939
R19123 gnd.n7169 gnd.n7168 0.152939
R19124 gnd.n7169 gnd.n525 0.152939
R19125 gnd.n7177 gnd.n525 0.152939
R19126 gnd.n7178 gnd.n7177 0.152939
R19127 gnd.n7179 gnd.n7178 0.152939
R19128 gnd.n7179 gnd.n519 0.152939
R19129 gnd.n7187 gnd.n519 0.152939
R19130 gnd.n7188 gnd.n7187 0.152939
R19131 gnd.n7189 gnd.n7188 0.152939
R19132 gnd.n7189 gnd.n513 0.152939
R19133 gnd.n7197 gnd.n513 0.152939
R19134 gnd.n7198 gnd.n7197 0.152939
R19135 gnd.n7199 gnd.n7198 0.152939
R19136 gnd.n7199 gnd.n507 0.152939
R19137 gnd.n7207 gnd.n507 0.152939
R19138 gnd.n7208 gnd.n7207 0.152939
R19139 gnd.n7209 gnd.n7208 0.152939
R19140 gnd.n7209 gnd.n501 0.152939
R19141 gnd.n7217 gnd.n501 0.152939
R19142 gnd.n7218 gnd.n7217 0.152939
R19143 gnd.n7219 gnd.n7218 0.152939
R19144 gnd.n7219 gnd.n495 0.152939
R19145 gnd.n7227 gnd.n495 0.152939
R19146 gnd.n7228 gnd.n7227 0.152939
R19147 gnd.n7229 gnd.n7228 0.152939
R19148 gnd.n7229 gnd.n489 0.152939
R19149 gnd.n7237 gnd.n489 0.152939
R19150 gnd.n7238 gnd.n7237 0.152939
R19151 gnd.n7239 gnd.n7238 0.152939
R19152 gnd.n7239 gnd.n483 0.152939
R19153 gnd.n7247 gnd.n483 0.152939
R19154 gnd.n7248 gnd.n7247 0.152939
R19155 gnd.n7249 gnd.n7248 0.152939
R19156 gnd.n7249 gnd.n477 0.152939
R19157 gnd.n7257 gnd.n477 0.152939
R19158 gnd.n7258 gnd.n7257 0.152939
R19159 gnd.n7259 gnd.n7258 0.152939
R19160 gnd.n7259 gnd.n471 0.152939
R19161 gnd.n7267 gnd.n471 0.152939
R19162 gnd.n7268 gnd.n7267 0.152939
R19163 gnd.n7269 gnd.n7268 0.152939
R19164 gnd.n7269 gnd.n465 0.152939
R19165 gnd.n7277 gnd.n465 0.152939
R19166 gnd.n7278 gnd.n7277 0.152939
R19167 gnd.n7279 gnd.n7278 0.152939
R19168 gnd.n7279 gnd.n459 0.152939
R19169 gnd.n7287 gnd.n459 0.152939
R19170 gnd.n7288 gnd.n7287 0.152939
R19171 gnd.n7289 gnd.n7288 0.152939
R19172 gnd.n7289 gnd.n453 0.152939
R19173 gnd.n7297 gnd.n453 0.152939
R19174 gnd.n7298 gnd.n7297 0.152939
R19175 gnd.n7299 gnd.n7298 0.152939
R19176 gnd.n7299 gnd.n447 0.152939
R19177 gnd.n7307 gnd.n447 0.152939
R19178 gnd.n7308 gnd.n7307 0.152939
R19179 gnd.n7309 gnd.n7308 0.152939
R19180 gnd.n7309 gnd.n441 0.152939
R19181 gnd.n7317 gnd.n441 0.152939
R19182 gnd.n7318 gnd.n7317 0.152939
R19183 gnd.n7319 gnd.n7318 0.152939
R19184 gnd.n7319 gnd.n435 0.152939
R19185 gnd.n7327 gnd.n435 0.152939
R19186 gnd.n7328 gnd.n7327 0.152939
R19187 gnd.n7329 gnd.n7328 0.152939
R19188 gnd.n7329 gnd.n429 0.152939
R19189 gnd.n7337 gnd.n429 0.152939
R19190 gnd.n7338 gnd.n7337 0.152939
R19191 gnd.n7339 gnd.n7338 0.152939
R19192 gnd.n7339 gnd.n423 0.152939
R19193 gnd.n7348 gnd.n423 0.152939
R19194 gnd.n7349 gnd.n7348 0.152939
R19195 gnd.n7350 gnd.n7349 0.152939
R19196 gnd.n7557 gnd.n7556 0.152939
R19197 gnd.n7557 gnd.n287 0.152939
R19198 gnd.n7571 gnd.n287 0.152939
R19199 gnd.n7572 gnd.n7571 0.152939
R19200 gnd.n7573 gnd.n7572 0.152939
R19201 gnd.n7573 gnd.n273 0.152939
R19202 gnd.n7587 gnd.n273 0.152939
R19203 gnd.n7588 gnd.n7587 0.152939
R19204 gnd.n7589 gnd.n7588 0.152939
R19205 gnd.n7589 gnd.n257 0.152939
R19206 gnd.n7603 gnd.n257 0.152939
R19207 gnd.n7604 gnd.n7603 0.152939
R19208 gnd.n7605 gnd.n7604 0.152939
R19209 gnd.n7605 gnd.n242 0.152939
R19210 gnd.n7619 gnd.n242 0.152939
R19211 gnd.n7620 gnd.n7619 0.152939
R19212 gnd.n7621 gnd.n7620 0.152939
R19213 gnd.n7621 gnd.n226 0.152939
R19214 gnd.n7635 gnd.n226 0.152939
R19215 gnd.n7636 gnd.n7635 0.152939
R19216 gnd.n7637 gnd.n7636 0.152939
R19217 gnd.n7637 gnd.n210 0.152939
R19218 gnd.n7719 gnd.n210 0.152939
R19219 gnd.n7720 gnd.n7719 0.152939
R19220 gnd.n7721 gnd.n7720 0.152939
R19221 gnd.n7721 gnd.n133 0.152939
R19222 gnd.n7801 gnd.n133 0.152939
R19223 gnd.n7800 gnd.n134 0.152939
R19224 gnd.n136 gnd.n134 0.152939
R19225 gnd.n140 gnd.n136 0.152939
R19226 gnd.n141 gnd.n140 0.152939
R19227 gnd.n142 gnd.n141 0.152939
R19228 gnd.n143 gnd.n142 0.152939
R19229 gnd.n147 gnd.n143 0.152939
R19230 gnd.n148 gnd.n147 0.152939
R19231 gnd.n149 gnd.n148 0.152939
R19232 gnd.n150 gnd.n149 0.152939
R19233 gnd.n154 gnd.n150 0.152939
R19234 gnd.n155 gnd.n154 0.152939
R19235 gnd.n156 gnd.n155 0.152939
R19236 gnd.n157 gnd.n156 0.152939
R19237 gnd.n161 gnd.n157 0.152939
R19238 gnd.n162 gnd.n161 0.152939
R19239 gnd.n163 gnd.n162 0.152939
R19240 gnd.n164 gnd.n163 0.152939
R19241 gnd.n168 gnd.n164 0.152939
R19242 gnd.n169 gnd.n168 0.152939
R19243 gnd.n170 gnd.n169 0.152939
R19244 gnd.n171 gnd.n170 0.152939
R19245 gnd.n175 gnd.n171 0.152939
R19246 gnd.n176 gnd.n175 0.152939
R19247 gnd.n177 gnd.n176 0.152939
R19248 gnd.n178 gnd.n177 0.152939
R19249 gnd.n182 gnd.n178 0.152939
R19250 gnd.n183 gnd.n182 0.152939
R19251 gnd.n184 gnd.n183 0.152939
R19252 gnd.n185 gnd.n184 0.152939
R19253 gnd.n189 gnd.n185 0.152939
R19254 gnd.n190 gnd.n189 0.152939
R19255 gnd.n191 gnd.n190 0.152939
R19256 gnd.n192 gnd.n191 0.152939
R19257 gnd.n196 gnd.n192 0.152939
R19258 gnd.n197 gnd.n196 0.152939
R19259 gnd.n7731 gnd.n197 0.152939
R19260 gnd.n7731 gnd.n7730 0.152939
R19261 gnd.n1456 gnd.n1333 0.152939
R19262 gnd.n1457 gnd.n1456 0.152939
R19263 gnd.n1458 gnd.n1457 0.152939
R19264 gnd.n1459 gnd.n1458 0.152939
R19265 gnd.n1460 gnd.n1459 0.152939
R19266 gnd.n1461 gnd.n1460 0.152939
R19267 gnd.n1462 gnd.n1461 0.152939
R19268 gnd.n1463 gnd.n1462 0.152939
R19269 gnd.n1464 gnd.n1463 0.152939
R19270 gnd.n1464 gnd.n1390 0.152939
R19271 gnd.n6124 gnd.n1390 0.152939
R19272 gnd.n6125 gnd.n6124 0.152939
R19273 gnd.n6126 gnd.n6125 0.152939
R19274 gnd.n6126 gnd.n1388 0.152939
R19275 gnd.n6131 gnd.n1388 0.152939
R19276 gnd.n6132 gnd.n6131 0.152939
R19277 gnd.n6133 gnd.n6132 0.152939
R19278 gnd.n6134 gnd.n6133 0.152939
R19279 gnd.n6134 gnd.n387 0.152939
R19280 gnd.n7387 gnd.n387 0.152939
R19281 gnd.n7388 gnd.n7387 0.152939
R19282 gnd.n7389 gnd.n7388 0.152939
R19283 gnd.n7390 gnd.n7389 0.152939
R19284 gnd.n7391 gnd.n7390 0.152939
R19285 gnd.n7391 gnd.n353 0.152939
R19286 gnd.n7432 gnd.n353 0.152939
R19287 gnd.n7433 gnd.n7432 0.152939
R19288 gnd.n7434 gnd.n7433 0.152939
R19289 gnd.n7435 gnd.n7434 0.152939
R19290 gnd.n7436 gnd.n7435 0.152939
R19291 gnd.n7437 gnd.n7436 0.152939
R19292 gnd.n7437 gnd.n337 0.152939
R19293 gnd.n7462 gnd.n337 0.152939
R19294 gnd.n7463 gnd.n7462 0.152939
R19295 gnd.n7464 gnd.n7463 0.152939
R19296 gnd.n7465 gnd.n7464 0.152939
R19297 gnd.n7466 gnd.n7465 0.152939
R19298 gnd.n7467 gnd.n7466 0.152939
R19299 gnd.n7468 gnd.n7467 0.152939
R19300 gnd.n7469 gnd.n7468 0.152939
R19301 gnd.n7470 gnd.n7469 0.152939
R19302 gnd.n7471 gnd.n7470 0.152939
R19303 gnd.n7472 gnd.n7471 0.152939
R19304 gnd.n7473 gnd.n7472 0.152939
R19305 gnd.n7474 gnd.n7473 0.152939
R19306 gnd.n7475 gnd.n7474 0.152939
R19307 gnd.n7476 gnd.n7475 0.152939
R19308 gnd.n7477 gnd.n7476 0.152939
R19309 gnd.n7478 gnd.n7477 0.152939
R19310 gnd.n7479 gnd.n7478 0.152939
R19311 gnd.n7480 gnd.n7479 0.152939
R19312 gnd.n7481 gnd.n7480 0.152939
R19313 gnd.n7482 gnd.n7481 0.152939
R19314 gnd.n7483 gnd.n7482 0.152939
R19315 gnd.n7484 gnd.n7483 0.152939
R19316 gnd.n7485 gnd.n7484 0.152939
R19317 gnd.n7486 gnd.n7485 0.152939
R19318 gnd.n7487 gnd.n7486 0.152939
R19319 gnd.n7488 gnd.n7487 0.152939
R19320 gnd.n7489 gnd.n7488 0.152939
R19321 gnd.n7491 gnd.n7489 0.152939
R19322 gnd.n7491 gnd.n7490 0.152939
R19323 gnd.n7490 gnd.n203 0.152939
R19324 gnd.n7729 gnd.n203 0.152939
R19325 gnd.n1290 gnd.n1289 0.152939
R19326 gnd.n1291 gnd.n1290 0.152939
R19327 gnd.n1292 gnd.n1291 0.152939
R19328 gnd.n1293 gnd.n1292 0.152939
R19329 gnd.n1294 gnd.n1293 0.152939
R19330 gnd.n1295 gnd.n1294 0.152939
R19331 gnd.n1296 gnd.n1295 0.152939
R19332 gnd.n1297 gnd.n1296 0.152939
R19333 gnd.n1298 gnd.n1297 0.152939
R19334 gnd.n1299 gnd.n1298 0.152939
R19335 gnd.n1300 gnd.n1299 0.152939
R19336 gnd.n1301 gnd.n1300 0.152939
R19337 gnd.n1302 gnd.n1301 0.152939
R19338 gnd.n1303 gnd.n1302 0.152939
R19339 gnd.n1304 gnd.n1303 0.152939
R19340 gnd.n1311 gnd.n1310 0.152939
R19341 gnd.n1312 gnd.n1311 0.152939
R19342 gnd.n1313 gnd.n1312 0.152939
R19343 gnd.n1314 gnd.n1313 0.152939
R19344 gnd.n1315 gnd.n1314 0.152939
R19345 gnd.n1316 gnd.n1315 0.152939
R19346 gnd.n1317 gnd.n1316 0.152939
R19347 gnd.n1318 gnd.n1317 0.152939
R19348 gnd.n1319 gnd.n1318 0.152939
R19349 gnd.n1320 gnd.n1319 0.152939
R19350 gnd.n1321 gnd.n1320 0.152939
R19351 gnd.n1322 gnd.n1321 0.152939
R19352 gnd.n1323 gnd.n1322 0.152939
R19353 gnd.n1324 gnd.n1323 0.152939
R19354 gnd.n1325 gnd.n1324 0.152939
R19355 gnd.n1326 gnd.n1325 0.152939
R19356 gnd.n1327 gnd.n1326 0.152939
R19357 gnd.n6224 gnd.n1327 0.152939
R19358 gnd.n6224 gnd.n6223 0.152939
R19359 gnd.n6223 gnd.n6222 0.152939
R19360 gnd.n6048 gnd.n6047 0.152939
R19361 gnd.n6049 gnd.n6048 0.152939
R19362 gnd.n6049 gnd.n1428 0.152939
R19363 gnd.n6077 gnd.n1428 0.152939
R19364 gnd.n6078 gnd.n6077 0.152939
R19365 gnd.n6079 gnd.n6078 0.152939
R19366 gnd.n6080 gnd.n6079 0.152939
R19367 gnd.n6080 gnd.n1401 0.152939
R19368 gnd.n6114 gnd.n1401 0.152939
R19369 gnd.n6115 gnd.n6114 0.152939
R19370 gnd.n6116 gnd.n6115 0.152939
R19371 gnd.n6117 gnd.n6116 0.152939
R19372 gnd.n6117 gnd.n1367 0.152939
R19373 gnd.n6184 gnd.n1367 0.152939
R19374 gnd.n6185 gnd.n6184 0.152939
R19375 gnd.n6186 gnd.n6185 0.152939
R19376 gnd.n6186 gnd.n396 0.152939
R19377 gnd.n7377 gnd.n396 0.152939
R19378 gnd.n7378 gnd.n7377 0.152939
R19379 gnd.n7379 gnd.n7378 0.152939
R19380 gnd.n7380 gnd.n7379 0.152939
R19381 gnd.n7380 gnd.n363 0.152939
R19382 gnd.n7423 gnd.n363 0.152939
R19383 gnd.n7424 gnd.n7423 0.152939
R19384 gnd.n7425 gnd.n7424 0.152939
R19385 gnd.n7425 gnd.n303 0.152939
R19386 gnd.n7556 gnd.n303 0.152939
R19387 gnd.n6545 gnd.n967 0.152939
R19388 gnd.n4371 gnd.n967 0.152939
R19389 gnd.n4372 gnd.n4371 0.152939
R19390 gnd.n4373 gnd.n4372 0.152939
R19391 gnd.n4373 gnd.n2164 0.152939
R19392 gnd.n4412 gnd.n2164 0.152939
R19393 gnd.n4413 gnd.n4412 0.152939
R19394 gnd.n4414 gnd.n4413 0.152939
R19395 gnd.n4414 gnd.n2160 0.152939
R19396 gnd.n4420 gnd.n2160 0.152939
R19397 gnd.n4421 gnd.n4420 0.152939
R19398 gnd.n4422 gnd.n4421 0.152939
R19399 gnd.n4422 gnd.n2143 0.152939
R19400 gnd.n4461 gnd.n2143 0.152939
R19401 gnd.n4462 gnd.n4461 0.152939
R19402 gnd.n4463 gnd.n4462 0.152939
R19403 gnd.n4463 gnd.n2139 0.152939
R19404 gnd.n4469 gnd.n2139 0.152939
R19405 gnd.n4470 gnd.n4469 0.152939
R19406 gnd.n4471 gnd.n4470 0.152939
R19407 gnd.n4472 gnd.n4471 0.152939
R19408 gnd.n4473 gnd.n4472 0.152939
R19409 gnd.n4476 gnd.n4473 0.152939
R19410 gnd.n4477 gnd.n4476 0.152939
R19411 gnd.n4478 gnd.n4477 0.152939
R19412 gnd.n4479 gnd.n4478 0.152939
R19413 gnd.n4482 gnd.n4479 0.152939
R19414 gnd.n4483 gnd.n4482 0.152939
R19415 gnd.n4484 gnd.n4483 0.152939
R19416 gnd.n4485 gnd.n4484 0.152939
R19417 gnd.n4487 gnd.n4485 0.152939
R19418 gnd.n4488 gnd.n4487 0.152939
R19419 gnd.n4488 gnd.n1964 0.152939
R19420 gnd.n5618 gnd.n1964 0.152939
R19421 gnd.n5619 gnd.n5618 0.152939
R19422 gnd.n5620 gnd.n5619 0.152939
R19423 gnd.n5620 gnd.n1950 0.152939
R19424 gnd.n5634 gnd.n1950 0.152939
R19425 gnd.n5635 gnd.n5634 0.152939
R19426 gnd.n5636 gnd.n5635 0.152939
R19427 gnd.n5636 gnd.n1938 0.152939
R19428 gnd.n5650 gnd.n1938 0.152939
R19429 gnd.n5651 gnd.n5650 0.152939
R19430 gnd.n5652 gnd.n5651 0.152939
R19431 gnd.n5652 gnd.n1925 0.152939
R19432 gnd.n5666 gnd.n1925 0.152939
R19433 gnd.n5667 gnd.n5666 0.152939
R19434 gnd.n5668 gnd.n5667 0.152939
R19435 gnd.n5668 gnd.n1910 0.152939
R19436 gnd.n5682 gnd.n1910 0.152939
R19437 gnd.n5683 gnd.n5682 0.152939
R19438 gnd.n5684 gnd.n5683 0.152939
R19439 gnd.n5684 gnd.n1896 0.152939
R19440 gnd.n5698 gnd.n1896 0.152939
R19441 gnd.n5699 gnd.n5698 0.152939
R19442 gnd.n5700 gnd.n5699 0.152939
R19443 gnd.n5700 gnd.n1882 0.152939
R19444 gnd.n5714 gnd.n1882 0.152939
R19445 gnd.n5715 gnd.n5714 0.152939
R19446 gnd.n5716 gnd.n5715 0.152939
R19447 gnd.n5716 gnd.n1867 0.152939
R19448 gnd.n5730 gnd.n1867 0.152939
R19449 gnd.n5731 gnd.n5730 0.152939
R19450 gnd.n5732 gnd.n5731 0.152939
R19451 gnd.n5732 gnd.n1854 0.152939
R19452 gnd.n5746 gnd.n1854 0.152939
R19453 gnd.n5747 gnd.n5746 0.152939
R19454 gnd.n5748 gnd.n5747 0.152939
R19455 gnd.n5748 gnd.n1839 0.152939
R19456 gnd.n5762 gnd.n1839 0.152939
R19457 gnd.n5763 gnd.n5762 0.152939
R19458 gnd.n5764 gnd.n5763 0.152939
R19459 gnd.n5764 gnd.n1824 0.152939
R19460 gnd.n5778 gnd.n1824 0.152939
R19461 gnd.n5779 gnd.n5778 0.152939
R19462 gnd.n5780 gnd.n5779 0.152939
R19463 gnd.n5780 gnd.n1809 0.152939
R19464 gnd.n5794 gnd.n1809 0.152939
R19465 gnd.n5795 gnd.n5794 0.152939
R19466 gnd.n5796 gnd.n5795 0.152939
R19467 gnd.n5796 gnd.n1794 0.152939
R19468 gnd.n5810 gnd.n1794 0.152939
R19469 gnd.n5811 gnd.n5810 0.152939
R19470 gnd.n5812 gnd.n5811 0.152939
R19471 gnd.n5812 gnd.n1780 0.152939
R19472 gnd.n5826 gnd.n1780 0.152939
R19473 gnd.n5827 gnd.n5826 0.152939
R19474 gnd.n5828 gnd.n5827 0.152939
R19475 gnd.n5828 gnd.n1765 0.152939
R19476 gnd.n5842 gnd.n1765 0.152939
R19477 gnd.n5843 gnd.n5842 0.152939
R19478 gnd.n5844 gnd.n5843 0.152939
R19479 gnd.n5844 gnd.n1750 0.152939
R19480 gnd.n5858 gnd.n1750 0.152939
R19481 gnd.n5859 gnd.n5858 0.152939
R19482 gnd.n5860 gnd.n5859 0.152939
R19483 gnd.n5860 gnd.n1736 0.152939
R19484 gnd.n5874 gnd.n1736 0.152939
R19485 gnd.n5875 gnd.n5874 0.152939
R19486 gnd.n5876 gnd.n5875 0.152939
R19487 gnd.n5876 gnd.n1721 0.152939
R19488 gnd.n5890 gnd.n1721 0.152939
R19489 gnd.n5891 gnd.n5890 0.152939
R19490 gnd.n5892 gnd.n5891 0.152939
R19491 gnd.n5892 gnd.n1707 0.152939
R19492 gnd.n5906 gnd.n1707 0.152939
R19493 gnd.n5907 gnd.n5906 0.152939
R19494 gnd.n5908 gnd.n5907 0.152939
R19495 gnd.n5908 gnd.n1691 0.152939
R19496 gnd.n5922 gnd.n1691 0.152939
R19497 gnd.n5923 gnd.n5922 0.152939
R19498 gnd.n5924 gnd.n5923 0.152939
R19499 gnd.n5924 gnd.n1677 0.152939
R19500 gnd.n5938 gnd.n1677 0.152939
R19501 gnd.n5939 gnd.n5938 0.152939
R19502 gnd.n5940 gnd.n5939 0.152939
R19503 gnd.n5940 gnd.n1665 0.152939
R19504 gnd.n5954 gnd.n1665 0.152939
R19505 gnd.n5955 gnd.n5954 0.152939
R19506 gnd.n5956 gnd.n5955 0.152939
R19507 gnd.n5956 gnd.n1650 0.152939
R19508 gnd.n5970 gnd.n1650 0.152939
R19509 gnd.n5971 gnd.n5970 0.152939
R19510 gnd.n5972 gnd.n5971 0.152939
R19511 gnd.n5972 gnd.n1636 0.152939
R19512 gnd.n5986 gnd.n1636 0.152939
R19513 gnd.n5987 gnd.n5986 0.152939
R19514 gnd.n5988 gnd.n5987 0.152939
R19515 gnd.n5988 gnd.n1623 0.152939
R19516 gnd.n6004 gnd.n1623 0.152939
R19517 gnd.n6005 gnd.n6004 0.152939
R19518 gnd.n6006 gnd.n6005 0.152939
R19519 gnd.n6008 gnd.n6006 0.152939
R19520 gnd.n6008 gnd.n6007 0.152939
R19521 gnd.n6007 gnd.n1251 0.152939
R19522 gnd.n1252 gnd.n1251 0.152939
R19523 gnd.n1253 gnd.n1252 0.152939
R19524 gnd.n1443 gnd.n1253 0.152939
R19525 gnd.n1446 gnd.n1443 0.152939
R19526 gnd.n1447 gnd.n1446 0.152939
R19527 gnd.n1448 gnd.n1447 0.152939
R19528 gnd.n1448 gnd.n1439 0.152939
R19529 gnd.n6066 gnd.n1439 0.152939
R19530 gnd.n6067 gnd.n6066 0.152939
R19531 gnd.n6068 gnd.n6067 0.152939
R19532 gnd.n6069 gnd.n6068 0.152939
R19533 gnd.n6069 gnd.n1411 0.152939
R19534 gnd.n6102 gnd.n1411 0.152939
R19535 gnd.n6103 gnd.n6102 0.152939
R19536 gnd.n6104 gnd.n6103 0.152939
R19537 gnd.n6105 gnd.n6104 0.152939
R19538 gnd.n6105 gnd.n1377 0.152939
R19539 gnd.n6163 gnd.n1377 0.152939
R19540 gnd.n6164 gnd.n6163 0.152939
R19541 gnd.n6165 gnd.n6164 0.152939
R19542 gnd.n6166 gnd.n6165 0.152939
R19543 gnd.n6167 gnd.n6166 0.152939
R19544 gnd.n6169 gnd.n6167 0.152939
R19545 gnd.n6171 gnd.n6169 0.152939
R19546 gnd.n6171 gnd.n6170 0.152939
R19547 gnd.n6170 gnd.n412 0.152939
R19548 gnd.n413 gnd.n412 0.152939
R19549 gnd.n414 gnd.n413 0.152939
R19550 gnd.n417 gnd.n414 0.152939
R19551 gnd.n418 gnd.n417 0.152939
R19552 gnd.n419 gnd.n418 0.152939
R19553 gnd.n420 gnd.n419 0.152939
R19554 gnd.n3879 gnd.n3878 0.152939
R19555 gnd.n3880 gnd.n3879 0.152939
R19556 gnd.n3881 gnd.n3880 0.152939
R19557 gnd.n3882 gnd.n3881 0.152939
R19558 gnd.n3883 gnd.n3882 0.152939
R19559 gnd.n3884 gnd.n3883 0.152939
R19560 gnd.n3885 gnd.n3884 0.152939
R19561 gnd.n3886 gnd.n3885 0.152939
R19562 gnd.n3887 gnd.n3886 0.152939
R19563 gnd.n3888 gnd.n3887 0.152939
R19564 gnd.n3889 gnd.n3888 0.152939
R19565 gnd.n3890 gnd.n3889 0.152939
R19566 gnd.n3891 gnd.n3890 0.152939
R19567 gnd.n3892 gnd.n3891 0.152939
R19568 gnd.n3893 gnd.n3892 0.152939
R19569 gnd.n3894 gnd.n3893 0.152939
R19570 gnd.n3895 gnd.n3894 0.152939
R19571 gnd.n3896 gnd.n3895 0.152939
R19572 gnd.n3897 gnd.n3896 0.152939
R19573 gnd.n3898 gnd.n3897 0.152939
R19574 gnd.n3899 gnd.n3898 0.152939
R19575 gnd.n3900 gnd.n3899 0.152939
R19576 gnd.n3901 gnd.n3900 0.152939
R19577 gnd.n3902 gnd.n3901 0.152939
R19578 gnd.n3903 gnd.n3902 0.152939
R19579 gnd.n3904 gnd.n3903 0.152939
R19580 gnd.n3905 gnd.n3904 0.152939
R19581 gnd.n3906 gnd.n3905 0.152939
R19582 gnd.n3907 gnd.n3906 0.152939
R19583 gnd.n3908 gnd.n3907 0.152939
R19584 gnd.n3909 gnd.n3908 0.152939
R19585 gnd.n3830 gnd.n2332 0.152939
R19586 gnd.n3838 gnd.n3830 0.152939
R19587 gnd.n3839 gnd.n3838 0.152939
R19588 gnd.n3840 gnd.n3839 0.152939
R19589 gnd.n3840 gnd.n3826 0.152939
R19590 gnd.n3848 gnd.n3826 0.152939
R19591 gnd.n3849 gnd.n3848 0.152939
R19592 gnd.n3850 gnd.n3849 0.152939
R19593 gnd.n3850 gnd.n3822 0.152939
R19594 gnd.n3858 gnd.n3822 0.152939
R19595 gnd.n3859 gnd.n3858 0.152939
R19596 gnd.n3860 gnd.n3859 0.152939
R19597 gnd.n3860 gnd.n3818 0.152939
R19598 gnd.n3868 gnd.n3818 0.152939
R19599 gnd.n3869 gnd.n3868 0.152939
R19600 gnd.n3870 gnd.n3869 0.152939
R19601 gnd.n3870 gnd.n3812 0.152939
R19602 gnd.n3877 gnd.n3812 0.152939
R19603 gnd.n4198 gnd.n4197 0.152939
R19604 gnd.n4199 gnd.n4198 0.152939
R19605 gnd.n4199 gnd.n2317 0.152939
R19606 gnd.n4213 gnd.n2317 0.152939
R19607 gnd.n4214 gnd.n4213 0.152939
R19608 gnd.n4215 gnd.n4214 0.152939
R19609 gnd.n4215 gnd.n2300 0.152939
R19610 gnd.n4229 gnd.n2300 0.152939
R19611 gnd.n4230 gnd.n4229 0.152939
R19612 gnd.n4231 gnd.n4230 0.152939
R19613 gnd.n4231 gnd.n2285 0.152939
R19614 gnd.n4245 gnd.n2285 0.152939
R19615 gnd.n4246 gnd.n4245 0.152939
R19616 gnd.n4247 gnd.n4246 0.152939
R19617 gnd.n4247 gnd.n2268 0.152939
R19618 gnd.n4261 gnd.n2268 0.152939
R19619 gnd.n4262 gnd.n4261 0.152939
R19620 gnd.n4263 gnd.n4262 0.152939
R19621 gnd.n4263 gnd.n2253 0.152939
R19622 gnd.n4277 gnd.n2253 0.152939
R19623 gnd.n4278 gnd.n4277 0.152939
R19624 gnd.n4279 gnd.n4278 0.152939
R19625 gnd.n4279 gnd.n2236 0.152939
R19626 gnd.n4294 gnd.n2236 0.152939
R19627 gnd.n4295 gnd.n4294 0.152939
R19628 gnd.n4296 gnd.n4295 0.152939
R19629 gnd.n4296 gnd.n2222 0.152939
R19630 gnd.n4310 gnd.n2222 0.152939
R19631 gnd.n4311 gnd.n4310 0.152939
R19632 gnd.n4312 gnd.n4311 0.152939
R19633 gnd.n4312 gnd.n2197 0.152939
R19634 gnd.n4328 gnd.n2197 0.152939
R19635 gnd.n4329 gnd.n4328 0.152939
R19636 gnd.n4330 gnd.n4329 0.152939
R19637 gnd.n4331 gnd.n4330 0.152939
R19638 gnd.n4332 gnd.n4331 0.152939
R19639 gnd.n4333 gnd.n4332 0.152939
R19640 gnd.n4335 gnd.n4333 0.152939
R19641 gnd.n4335 gnd.n4334 0.152939
R19642 gnd.n4334 gnd.n990 0.152939
R19643 gnd.n991 gnd.n990 0.152939
R19644 gnd.n992 gnd.n991 0.152939
R19645 gnd.n1009 gnd.n992 0.152939
R19646 gnd.n1010 gnd.n1009 0.152939
R19647 gnd.n1011 gnd.n1010 0.152939
R19648 gnd.n1012 gnd.n1011 0.152939
R19649 gnd.n1031 gnd.n1012 0.152939
R19650 gnd.n1032 gnd.n1031 0.152939
R19651 gnd.n1033 gnd.n1032 0.152939
R19652 gnd.n1034 gnd.n1033 0.152939
R19653 gnd.n1051 gnd.n1034 0.152939
R19654 gnd.n1052 gnd.n1051 0.152939
R19655 gnd.n1053 gnd.n1052 0.152939
R19656 gnd.n1054 gnd.n1053 0.152939
R19657 gnd.n1073 gnd.n1054 0.152939
R19658 gnd.n1074 gnd.n1073 0.152939
R19659 gnd.n1075 gnd.n1074 0.152939
R19660 gnd.n1076 gnd.n1075 0.152939
R19661 gnd.n1094 gnd.n1076 0.152939
R19662 gnd.n1095 gnd.n1094 0.152939
R19663 gnd.n1096 gnd.n1095 0.152939
R19664 gnd.n1097 gnd.n1096 0.152939
R19665 gnd.n1114 gnd.n1097 0.152939
R19666 gnd.n6460 gnd.n1114 0.152939
R19667 gnd.n978 gnd.n966 0.152939
R19668 gnd.n979 gnd.n978 0.152939
R19669 gnd.n980 gnd.n979 0.152939
R19670 gnd.n999 gnd.n980 0.152939
R19671 gnd.n1000 gnd.n999 0.152939
R19672 gnd.n1001 gnd.n1000 0.152939
R19673 gnd.n1002 gnd.n1001 0.152939
R19674 gnd.n1020 gnd.n1002 0.152939
R19675 gnd.n1021 gnd.n1020 0.152939
R19676 gnd.n1022 gnd.n1021 0.152939
R19677 gnd.n1023 gnd.n1022 0.152939
R19678 gnd.n1041 gnd.n1023 0.152939
R19679 gnd.n1042 gnd.n1041 0.152939
R19680 gnd.n1043 gnd.n1042 0.152939
R19681 gnd.n1044 gnd.n1043 0.152939
R19682 gnd.n1062 gnd.n1044 0.152939
R19683 gnd.n1063 gnd.n1062 0.152939
R19684 gnd.n1064 gnd.n1063 0.152939
R19685 gnd.n1065 gnd.n1064 0.152939
R19686 gnd.n1083 gnd.n1065 0.152939
R19687 gnd.n1084 gnd.n1083 0.152939
R19688 gnd.n1085 gnd.n1084 0.152939
R19689 gnd.n1086 gnd.n1085 0.152939
R19690 gnd.n1104 gnd.n1086 0.152939
R19691 gnd.n1105 gnd.n1104 0.152939
R19692 gnd.n1106 gnd.n1105 0.152939
R19693 gnd.n1107 gnd.n1106 0.152939
R19694 gnd.n2082 gnd.n2081 0.152939
R19695 gnd.n2083 gnd.n2082 0.152939
R19696 gnd.n2084 gnd.n2083 0.152939
R19697 gnd.n2085 gnd.n2084 0.152939
R19698 gnd.n2086 gnd.n2085 0.152939
R19699 gnd.n2087 gnd.n2086 0.152939
R19700 gnd.n2088 gnd.n2087 0.152939
R19701 gnd.n2089 gnd.n2088 0.152939
R19702 gnd.n2090 gnd.n2089 0.152939
R19703 gnd.n2091 gnd.n2090 0.152939
R19704 gnd.n2092 gnd.n2091 0.152939
R19705 gnd.n2093 gnd.n2092 0.152939
R19706 gnd.n2094 gnd.n2093 0.152939
R19707 gnd.n2095 gnd.n2094 0.152939
R19708 gnd.n2096 gnd.n2095 0.152939
R19709 gnd.n4615 gnd.n4614 0.152939
R19710 gnd.n4614 gnd.n2101 0.152939
R19711 gnd.n2102 gnd.n2101 0.152939
R19712 gnd.n2103 gnd.n2102 0.152939
R19713 gnd.n2104 gnd.n2103 0.152939
R19714 gnd.n2105 gnd.n2104 0.152939
R19715 gnd.n2106 gnd.n2105 0.152939
R19716 gnd.n2107 gnd.n2106 0.152939
R19717 gnd.n2108 gnd.n2107 0.152939
R19718 gnd.n2109 gnd.n2108 0.152939
R19719 gnd.n2110 gnd.n2109 0.152939
R19720 gnd.n2111 gnd.n2110 0.152939
R19721 gnd.n2112 gnd.n2111 0.152939
R19722 gnd.n2113 gnd.n2112 0.152939
R19723 gnd.n2114 gnd.n2113 0.152939
R19724 gnd.n2115 gnd.n2114 0.152939
R19725 gnd.n2116 gnd.n2115 0.152939
R19726 gnd.n2117 gnd.n2116 0.152939
R19727 gnd.n4574 gnd.n2117 0.152939
R19728 gnd.n4574 gnd.n4573 0.152939
R19729 gnd.n4111 gnd.n4035 0.152939
R19730 gnd.n4037 gnd.n4035 0.152939
R19731 gnd.n4038 gnd.n4037 0.152939
R19732 gnd.n4039 gnd.n4038 0.152939
R19733 gnd.n4040 gnd.n4039 0.152939
R19734 gnd.n4041 gnd.n4040 0.152939
R19735 gnd.n4042 gnd.n4041 0.152939
R19736 gnd.n4043 gnd.n4042 0.152939
R19737 gnd.n4044 gnd.n4043 0.152939
R19738 gnd.n4045 gnd.n4044 0.152939
R19739 gnd.n4046 gnd.n4045 0.152939
R19740 gnd.n4047 gnd.n4046 0.152939
R19741 gnd.n4048 gnd.n4047 0.152939
R19742 gnd.n4049 gnd.n4048 0.152939
R19743 gnd.n4050 gnd.n4049 0.152939
R19744 gnd.n4051 gnd.n4050 0.152939
R19745 gnd.n4052 gnd.n4051 0.152939
R19746 gnd.n4053 gnd.n4052 0.152939
R19747 gnd.n4054 gnd.n4053 0.152939
R19748 gnd.n4055 gnd.n4054 0.152939
R19749 gnd.n4056 gnd.n4055 0.152939
R19750 gnd.n4057 gnd.n4056 0.152939
R19751 gnd.n4058 gnd.n4057 0.152939
R19752 gnd.n4059 gnd.n4058 0.152939
R19753 gnd.n4060 gnd.n4059 0.152939
R19754 gnd.n4061 gnd.n4060 0.152939
R19755 gnd.n4062 gnd.n4061 0.152939
R19756 gnd.n4063 gnd.n4062 0.152939
R19757 gnd.n4064 gnd.n4063 0.152939
R19758 gnd.n4065 gnd.n4064 0.152939
R19759 gnd.n4065 gnd.n2199 0.152939
R19760 gnd.n4327 gnd.n2199 0.152939
R19761 gnd.n4327 gnd.n2200 0.152939
R19762 gnd.n2202 gnd.n2200 0.152939
R19763 gnd.n2203 gnd.n2202 0.152939
R19764 gnd.n2203 gnd.n2182 0.152939
R19765 gnd.n4354 gnd.n2182 0.152939
R19766 gnd.n4355 gnd.n4354 0.152939
R19767 gnd.n4356 gnd.n4355 0.152939
R19768 gnd.n4356 gnd.n2176 0.152939
R19769 gnd.n4380 gnd.n2176 0.152939
R19770 gnd.n4381 gnd.n4380 0.152939
R19771 gnd.n4382 gnd.n4381 0.152939
R19772 gnd.n4382 gnd.n2174 0.152939
R19773 gnd.n4388 gnd.n2174 0.152939
R19774 gnd.n4389 gnd.n4388 0.152939
R19775 gnd.n4390 gnd.n4389 0.152939
R19776 gnd.n4390 gnd.n2155 0.152939
R19777 gnd.n4429 gnd.n2155 0.152939
R19778 gnd.n4430 gnd.n4429 0.152939
R19779 gnd.n4431 gnd.n4430 0.152939
R19780 gnd.n4431 gnd.n2153 0.152939
R19781 gnd.n4437 gnd.n2153 0.152939
R19782 gnd.n4438 gnd.n4437 0.152939
R19783 gnd.n4439 gnd.n4438 0.152939
R19784 gnd.n4440 gnd.n4439 0.152939
R19785 gnd.n4441 gnd.n4440 0.152939
R19786 gnd.n4441 gnd.n2130 0.152939
R19787 gnd.n4522 gnd.n2130 0.152939
R19788 gnd.n4523 gnd.n4522 0.152939
R19789 gnd.n4525 gnd.n4523 0.152939
R19790 gnd.n4525 gnd.n4524 0.152939
R19791 gnd.n4524 gnd.n2122 0.152939
R19792 gnd.n4572 gnd.n2122 0.152939
R19793 gnd.n4190 gnd.n3974 0.152939
R19794 gnd.n3977 gnd.n3974 0.152939
R19795 gnd.n3978 gnd.n3977 0.152939
R19796 gnd.n3979 gnd.n3978 0.152939
R19797 gnd.n3982 gnd.n3979 0.152939
R19798 gnd.n3983 gnd.n3982 0.152939
R19799 gnd.n3984 gnd.n3983 0.152939
R19800 gnd.n3985 gnd.n3984 0.152939
R19801 gnd.n3988 gnd.n3985 0.152939
R19802 gnd.n3989 gnd.n3988 0.152939
R19803 gnd.n3990 gnd.n3989 0.152939
R19804 gnd.n3991 gnd.n3990 0.152939
R19805 gnd.n3994 gnd.n3991 0.152939
R19806 gnd.n3995 gnd.n3994 0.152939
R19807 gnd.n3996 gnd.n3995 0.152939
R19808 gnd.n3997 gnd.n3996 0.152939
R19809 gnd.n4003 gnd.n3997 0.152939
R19810 gnd.n4004 gnd.n4003 0.152939
R19811 gnd.n4005 gnd.n4004 0.152939
R19812 gnd.n4006 gnd.n4005 0.152939
R19813 gnd.n4009 gnd.n4006 0.152939
R19814 gnd.n4010 gnd.n4009 0.152939
R19815 gnd.n4011 gnd.n4010 0.152939
R19816 gnd.n4012 gnd.n4011 0.152939
R19817 gnd.n4015 gnd.n4012 0.152939
R19818 gnd.n4016 gnd.n4015 0.152939
R19819 gnd.n4017 gnd.n4016 0.152939
R19820 gnd.n4018 gnd.n4017 0.152939
R19821 gnd.n4021 gnd.n4018 0.152939
R19822 gnd.n4022 gnd.n4021 0.152939
R19823 gnd.n4023 gnd.n4022 0.152939
R19824 gnd.n4024 gnd.n4023 0.152939
R19825 gnd.n4027 gnd.n4024 0.152939
R19826 gnd.n4028 gnd.n4027 0.152939
R19827 gnd.n4029 gnd.n4028 0.152939
R19828 gnd.n4118 gnd.n4029 0.152939
R19829 gnd.n4118 gnd.n4117 0.152939
R19830 gnd.n4117 gnd.n4116 0.152939
R19831 gnd.n4191 gnd.n2325 0.152939
R19832 gnd.n4205 gnd.n2325 0.152939
R19833 gnd.n4206 gnd.n4205 0.152939
R19834 gnd.n4207 gnd.n4206 0.152939
R19835 gnd.n4207 gnd.n2309 0.152939
R19836 gnd.n4221 gnd.n2309 0.152939
R19837 gnd.n4222 gnd.n4221 0.152939
R19838 gnd.n4223 gnd.n4222 0.152939
R19839 gnd.n4223 gnd.n2293 0.152939
R19840 gnd.n4237 gnd.n2293 0.152939
R19841 gnd.n4238 gnd.n4237 0.152939
R19842 gnd.n4239 gnd.n4238 0.152939
R19843 gnd.n4239 gnd.n2277 0.152939
R19844 gnd.n4253 gnd.n2277 0.152939
R19845 gnd.n4254 gnd.n4253 0.152939
R19846 gnd.n4255 gnd.n4254 0.152939
R19847 gnd.n4255 gnd.n2261 0.152939
R19848 gnd.n4269 gnd.n2261 0.152939
R19849 gnd.n4270 gnd.n4269 0.152939
R19850 gnd.n4271 gnd.n4270 0.152939
R19851 gnd.n4271 gnd.n2245 0.152939
R19852 gnd.n4285 gnd.n2245 0.152939
R19853 gnd.n4286 gnd.n4285 0.152939
R19854 gnd.n4288 gnd.n4286 0.152939
R19855 gnd.n4288 gnd.n4287 0.152939
R19856 gnd.n4287 gnd.n2230 0.152939
R19857 gnd.n2230 gnd.n966 0.152939
R19858 gnd.n6717 gnd.n799 0.152939
R19859 gnd.n804 gnd.n799 0.152939
R19860 gnd.n805 gnd.n804 0.152939
R19861 gnd.n806 gnd.n805 0.152939
R19862 gnd.n807 gnd.n806 0.152939
R19863 gnd.n812 gnd.n807 0.152939
R19864 gnd.n813 gnd.n812 0.152939
R19865 gnd.n814 gnd.n813 0.152939
R19866 gnd.n815 gnd.n814 0.152939
R19867 gnd.n820 gnd.n815 0.152939
R19868 gnd.n821 gnd.n820 0.152939
R19869 gnd.n822 gnd.n821 0.152939
R19870 gnd.n823 gnd.n822 0.152939
R19871 gnd.n828 gnd.n823 0.152939
R19872 gnd.n829 gnd.n828 0.152939
R19873 gnd.n830 gnd.n829 0.152939
R19874 gnd.n831 gnd.n830 0.152939
R19875 gnd.n836 gnd.n831 0.152939
R19876 gnd.n837 gnd.n836 0.152939
R19877 gnd.n838 gnd.n837 0.152939
R19878 gnd.n839 gnd.n838 0.152939
R19879 gnd.n844 gnd.n839 0.152939
R19880 gnd.n845 gnd.n844 0.152939
R19881 gnd.n846 gnd.n845 0.152939
R19882 gnd.n847 gnd.n846 0.152939
R19883 gnd.n852 gnd.n847 0.152939
R19884 gnd.n853 gnd.n852 0.152939
R19885 gnd.n854 gnd.n853 0.152939
R19886 gnd.n855 gnd.n854 0.152939
R19887 gnd.n860 gnd.n855 0.152939
R19888 gnd.n861 gnd.n860 0.152939
R19889 gnd.n862 gnd.n861 0.152939
R19890 gnd.n863 gnd.n862 0.152939
R19891 gnd.n868 gnd.n863 0.152939
R19892 gnd.n869 gnd.n868 0.152939
R19893 gnd.n870 gnd.n869 0.152939
R19894 gnd.n871 gnd.n870 0.152939
R19895 gnd.n876 gnd.n871 0.152939
R19896 gnd.n877 gnd.n876 0.152939
R19897 gnd.n878 gnd.n877 0.152939
R19898 gnd.n879 gnd.n878 0.152939
R19899 gnd.n884 gnd.n879 0.152939
R19900 gnd.n885 gnd.n884 0.152939
R19901 gnd.n886 gnd.n885 0.152939
R19902 gnd.n887 gnd.n886 0.152939
R19903 gnd.n892 gnd.n887 0.152939
R19904 gnd.n893 gnd.n892 0.152939
R19905 gnd.n894 gnd.n893 0.152939
R19906 gnd.n895 gnd.n894 0.152939
R19907 gnd.n900 gnd.n895 0.152939
R19908 gnd.n901 gnd.n900 0.152939
R19909 gnd.n902 gnd.n901 0.152939
R19910 gnd.n903 gnd.n902 0.152939
R19911 gnd.n908 gnd.n903 0.152939
R19912 gnd.n909 gnd.n908 0.152939
R19913 gnd.n910 gnd.n909 0.152939
R19914 gnd.n911 gnd.n910 0.152939
R19915 gnd.n916 gnd.n911 0.152939
R19916 gnd.n917 gnd.n916 0.152939
R19917 gnd.n918 gnd.n917 0.152939
R19918 gnd.n919 gnd.n918 0.152939
R19919 gnd.n924 gnd.n919 0.152939
R19920 gnd.n925 gnd.n924 0.152939
R19921 gnd.n926 gnd.n925 0.152939
R19922 gnd.n927 gnd.n926 0.152939
R19923 gnd.n932 gnd.n927 0.152939
R19924 gnd.n933 gnd.n932 0.152939
R19925 gnd.n934 gnd.n933 0.152939
R19926 gnd.n935 gnd.n934 0.152939
R19927 gnd.n940 gnd.n935 0.152939
R19928 gnd.n941 gnd.n940 0.152939
R19929 gnd.n942 gnd.n941 0.152939
R19930 gnd.n943 gnd.n942 0.152939
R19931 gnd.n948 gnd.n943 0.152939
R19932 gnd.n949 gnd.n948 0.152939
R19933 gnd.n950 gnd.n949 0.152939
R19934 gnd.n951 gnd.n950 0.152939
R19935 gnd.n956 gnd.n951 0.152939
R19936 gnd.n957 gnd.n956 0.152939
R19937 gnd.n958 gnd.n957 0.152939
R19938 gnd.n959 gnd.n958 0.152939
R19939 gnd.n964 gnd.n959 0.152939
R19940 gnd.n965 gnd.n964 0.152939
R19941 gnd.n6547 gnd.n965 0.152939
R19942 gnd.n6040 gnd.n1479 0.152939
R19943 gnd.n6036 gnd.n1479 0.152939
R19944 gnd.n6036 gnd.n6035 0.152939
R19945 gnd.n6035 gnd.n6034 0.152939
R19946 gnd.n6034 gnd.n1607 0.152939
R19947 gnd.n6027 gnd.n1607 0.152939
R19948 gnd.n6027 gnd.n6026 0.152939
R19949 gnd.n6026 gnd.n6025 0.152939
R19950 gnd.n6025 gnd.n6018 0.152939
R19951 gnd.n5612 gnd.n5611 0.152939
R19952 gnd.n5612 gnd.n1957 0.152939
R19953 gnd.n5626 gnd.n1957 0.152939
R19954 gnd.n5627 gnd.n5626 0.152939
R19955 gnd.n5628 gnd.n5627 0.152939
R19956 gnd.n5628 gnd.n1944 0.152939
R19957 gnd.n5642 gnd.n1944 0.152939
R19958 gnd.n5643 gnd.n5642 0.152939
R19959 gnd.n5644 gnd.n5643 0.152939
R19960 gnd.n5644 gnd.n1931 0.152939
R19961 gnd.n5658 gnd.n1931 0.152939
R19962 gnd.n5659 gnd.n5658 0.152939
R19963 gnd.n5660 gnd.n5659 0.152939
R19964 gnd.n5660 gnd.n1917 0.152939
R19965 gnd.n5674 gnd.n1917 0.152939
R19966 gnd.n5675 gnd.n5674 0.152939
R19967 gnd.n5676 gnd.n5675 0.152939
R19968 gnd.n5676 gnd.n1902 0.152939
R19969 gnd.n5690 gnd.n1902 0.152939
R19970 gnd.n5691 gnd.n5690 0.152939
R19971 gnd.n5692 gnd.n5691 0.152939
R19972 gnd.n5692 gnd.n1888 0.152939
R19973 gnd.n5706 gnd.n1888 0.152939
R19974 gnd.n5707 gnd.n5706 0.152939
R19975 gnd.n5708 gnd.n5707 0.152939
R19976 gnd.n5708 gnd.n1874 0.152939
R19977 gnd.n5722 gnd.n1874 0.152939
R19978 gnd.n5723 gnd.n5722 0.152939
R19979 gnd.n5724 gnd.n5723 0.152939
R19980 gnd.n5724 gnd.n1860 0.152939
R19981 gnd.n5738 gnd.n1860 0.152939
R19982 gnd.n5739 gnd.n5738 0.152939
R19983 gnd.n5740 gnd.n5739 0.152939
R19984 gnd.n5740 gnd.n1846 0.152939
R19985 gnd.n5754 gnd.n1846 0.152939
R19986 gnd.n5755 gnd.n5754 0.152939
R19987 gnd.n5756 gnd.n5755 0.152939
R19988 gnd.n5756 gnd.n1832 0.152939
R19989 gnd.n5770 gnd.n1832 0.152939
R19990 gnd.n5771 gnd.n5770 0.152939
R19991 gnd.n5772 gnd.n5771 0.152939
R19992 gnd.n5772 gnd.n1816 0.152939
R19993 gnd.n5786 gnd.n1816 0.152939
R19994 gnd.n5787 gnd.n5786 0.152939
R19995 gnd.n5788 gnd.n5787 0.152939
R19996 gnd.n5788 gnd.n1801 0.152939
R19997 gnd.n5802 gnd.n1801 0.152939
R19998 gnd.n5803 gnd.n5802 0.152939
R19999 gnd.n5804 gnd.n5803 0.152939
R20000 gnd.n5804 gnd.n1786 0.152939
R20001 gnd.n5818 gnd.n1786 0.152939
R20002 gnd.n5819 gnd.n5818 0.152939
R20003 gnd.n5820 gnd.n5819 0.152939
R20004 gnd.n5820 gnd.n1772 0.152939
R20005 gnd.n5834 gnd.n1772 0.152939
R20006 gnd.n5835 gnd.n5834 0.152939
R20007 gnd.n5836 gnd.n5835 0.152939
R20008 gnd.n5836 gnd.n1757 0.152939
R20009 gnd.n5850 gnd.n1757 0.152939
R20010 gnd.n5851 gnd.n5850 0.152939
R20011 gnd.n5852 gnd.n5851 0.152939
R20012 gnd.n5852 gnd.n1742 0.152939
R20013 gnd.n5866 gnd.n1742 0.152939
R20014 gnd.n5867 gnd.n5866 0.152939
R20015 gnd.n5868 gnd.n5867 0.152939
R20016 gnd.n5868 gnd.n1728 0.152939
R20017 gnd.n5882 gnd.n1728 0.152939
R20018 gnd.n5883 gnd.n5882 0.152939
R20019 gnd.n5884 gnd.n5883 0.152939
R20020 gnd.n5884 gnd.n1714 0.152939
R20021 gnd.n5898 gnd.n1714 0.152939
R20022 gnd.n5899 gnd.n5898 0.152939
R20023 gnd.n5900 gnd.n5899 0.152939
R20024 gnd.n5900 gnd.n1698 0.152939
R20025 gnd.n5914 gnd.n1698 0.152939
R20026 gnd.n5915 gnd.n5914 0.152939
R20027 gnd.n5916 gnd.n5915 0.152939
R20028 gnd.n5916 gnd.n1683 0.152939
R20029 gnd.n5930 gnd.n1683 0.152939
R20030 gnd.n5931 gnd.n5930 0.152939
R20031 gnd.n5932 gnd.n5931 0.152939
R20032 gnd.n5932 gnd.n1670 0.152939
R20033 gnd.n5946 gnd.n1670 0.152939
R20034 gnd.n5947 gnd.n5946 0.152939
R20035 gnd.n5948 gnd.n5947 0.152939
R20036 gnd.n5948 gnd.n1657 0.152939
R20037 gnd.n5962 gnd.n1657 0.152939
R20038 gnd.n5963 gnd.n5962 0.152939
R20039 gnd.n5964 gnd.n5963 0.152939
R20040 gnd.n5964 gnd.n1643 0.152939
R20041 gnd.n5978 gnd.n1643 0.152939
R20042 gnd.n5979 gnd.n5978 0.152939
R20043 gnd.n5980 gnd.n5979 0.152939
R20044 gnd.n5980 gnd.n1630 0.152939
R20045 gnd.n5994 gnd.n1630 0.152939
R20046 gnd.n5995 gnd.n5994 0.152939
R20047 gnd.n5998 gnd.n5995 0.152939
R20048 gnd.n5998 gnd.n5997 0.152939
R20049 gnd.n5997 gnd.n5996 0.152939
R20050 gnd.n5996 gnd.n1615 0.152939
R20051 gnd.n6017 gnd.n1615 0.152939
R20052 gnd.n4558 gnd.n4533 0.152939
R20053 gnd.n4558 gnd.n4557 0.152939
R20054 gnd.n4557 gnd.n4556 0.152939
R20055 gnd.n4556 gnd.n4539 0.152939
R20056 gnd.n4552 gnd.n4539 0.152939
R20057 gnd.n4552 gnd.n4551 0.152939
R20058 gnd.n4551 gnd.n4546 0.152939
R20059 gnd.n4546 gnd.n1970 0.152939
R20060 gnd.n5610 gnd.n1970 0.152939
R20061 gnd.n3922 gnd.n3921 0.152939
R20062 gnd.n3921 gnd.n3912 0.152939
R20063 gnd.n3917 gnd.n3912 0.152939
R20064 gnd.n3917 gnd.n3916 0.152939
R20065 gnd.n3916 gnd.n2179 0.152939
R20066 gnd.n4362 gnd.n2179 0.152939
R20067 gnd.n4363 gnd.n4362 0.152939
R20068 gnd.n4364 gnd.n4363 0.152939
R20069 gnd.n4364 gnd.n2170 0.152939
R20070 gnd.n4405 gnd.n2170 0.152939
R20071 gnd.n4405 gnd.n4404 0.152939
R20072 gnd.n4404 gnd.n4403 0.152939
R20073 gnd.n4403 gnd.n2171 0.152939
R20074 gnd.n4399 gnd.n2171 0.152939
R20075 gnd.n4399 gnd.n4398 0.152939
R20076 gnd.n4398 gnd.n4397 0.152939
R20077 gnd.n4397 gnd.n2149 0.152939
R20078 gnd.n4454 gnd.n2149 0.152939
R20079 gnd.n4454 gnd.n4453 0.152939
R20080 gnd.n4453 gnd.n4452 0.152939
R20081 gnd.n4452 gnd.n2150 0.152939
R20082 gnd.n4448 gnd.n2150 0.152939
R20083 gnd.n4448 gnd.n2133 0.152939
R20084 gnd.n4514 gnd.n2133 0.152939
R20085 gnd.n4515 gnd.n4514 0.152939
R20086 gnd.n4516 gnd.n4515 0.152939
R20087 gnd.n4516 gnd.n2127 0.152939
R20088 gnd.n4531 gnd.n2127 0.152939
R20089 gnd.n4532 gnd.n4531 0.152939
R20090 gnd.n4565 gnd.n4532 0.152939
R20091 gnd.n4565 gnd.n4564 0.152939
R20092 gnd.n6457 gnd.n1117 0.152939
R20093 gnd.n6453 gnd.n1117 0.152939
R20094 gnd.n6453 gnd.n6452 0.152939
R20095 gnd.n6452 gnd.n6451 0.152939
R20096 gnd.n6451 gnd.n1122 0.152939
R20097 gnd.n6447 gnd.n1122 0.152939
R20098 gnd.n6447 gnd.n6446 0.152939
R20099 gnd.n6446 gnd.n6445 0.152939
R20100 gnd.n6445 gnd.n1127 0.152939
R20101 gnd.n6441 gnd.n1127 0.152939
R20102 gnd.n6441 gnd.n6440 0.152939
R20103 gnd.n6440 gnd.n6439 0.152939
R20104 gnd.n6439 gnd.n1132 0.152939
R20105 gnd.n6435 gnd.n1132 0.152939
R20106 gnd.n6435 gnd.n6434 0.152939
R20107 gnd.n6434 gnd.n6433 0.152939
R20108 gnd.n6433 gnd.n1137 0.152939
R20109 gnd.n6429 gnd.n1137 0.152939
R20110 gnd.n6429 gnd.n6428 0.152939
R20111 gnd.n6428 gnd.n6427 0.152939
R20112 gnd.n6427 gnd.n1142 0.152939
R20113 gnd.n6423 gnd.n1142 0.152939
R20114 gnd.n6423 gnd.n6422 0.152939
R20115 gnd.n6422 gnd.n6421 0.152939
R20116 gnd.n6421 gnd.n1147 0.152939
R20117 gnd.n6417 gnd.n1147 0.152939
R20118 gnd.n6417 gnd.n6416 0.152939
R20119 gnd.n6416 gnd.n6415 0.152939
R20120 gnd.n6415 gnd.n1152 0.152939
R20121 gnd.n6411 gnd.n1152 0.152939
R20122 gnd.n6411 gnd.n6410 0.152939
R20123 gnd.n6410 gnd.n6409 0.152939
R20124 gnd.n6409 gnd.n1157 0.152939
R20125 gnd.n6405 gnd.n1157 0.152939
R20126 gnd.n6405 gnd.n6404 0.152939
R20127 gnd.n6404 gnd.n6403 0.152939
R20128 gnd.n6403 gnd.n1162 0.152939
R20129 gnd.n6399 gnd.n1162 0.152939
R20130 gnd.n6399 gnd.n6398 0.152939
R20131 gnd.n6398 gnd.n6397 0.152939
R20132 gnd.n6397 gnd.n1167 0.152939
R20133 gnd.n6393 gnd.n1167 0.152939
R20134 gnd.n6393 gnd.n6392 0.152939
R20135 gnd.n6392 gnd.n6391 0.152939
R20136 gnd.n6391 gnd.n1172 0.152939
R20137 gnd.n6387 gnd.n1172 0.152939
R20138 gnd.n6387 gnd.n6386 0.152939
R20139 gnd.n6386 gnd.n6385 0.152939
R20140 gnd.n6385 gnd.n1177 0.152939
R20141 gnd.n6381 gnd.n1177 0.152939
R20142 gnd.n6381 gnd.n6380 0.152939
R20143 gnd.n6380 gnd.n6379 0.152939
R20144 gnd.n6379 gnd.n1182 0.152939
R20145 gnd.n6375 gnd.n1182 0.152939
R20146 gnd.n6375 gnd.n6374 0.152939
R20147 gnd.n6374 gnd.n6373 0.152939
R20148 gnd.n6373 gnd.n1187 0.152939
R20149 gnd.n6369 gnd.n1187 0.152939
R20150 gnd.n6369 gnd.n6368 0.152939
R20151 gnd.n6368 gnd.n6367 0.152939
R20152 gnd.n6367 gnd.n1192 0.152939
R20153 gnd.n6363 gnd.n1192 0.152939
R20154 gnd.n6363 gnd.n6362 0.152939
R20155 gnd.n6362 gnd.n6361 0.152939
R20156 gnd.n6361 gnd.n1197 0.152939
R20157 gnd.n6357 gnd.n1197 0.152939
R20158 gnd.n6357 gnd.n6356 0.152939
R20159 gnd.n6356 gnd.n6355 0.152939
R20160 gnd.n6355 gnd.n1202 0.152939
R20161 gnd.n6351 gnd.n1202 0.152939
R20162 gnd.n6351 gnd.n6350 0.152939
R20163 gnd.n6350 gnd.n6349 0.152939
R20164 gnd.n6349 gnd.n1207 0.152939
R20165 gnd.n6345 gnd.n1207 0.152939
R20166 gnd.n6345 gnd.n6344 0.152939
R20167 gnd.n6344 gnd.n6343 0.152939
R20168 gnd.n6343 gnd.n1212 0.152939
R20169 gnd.n6339 gnd.n1212 0.152939
R20170 gnd.n6339 gnd.n6338 0.152939
R20171 gnd.n6338 gnd.n6337 0.152939
R20172 gnd.n6337 gnd.n1217 0.152939
R20173 gnd.n6333 gnd.n1217 0.152939
R20174 gnd.n6333 gnd.n6332 0.152939
R20175 gnd.n6332 gnd.n6331 0.152939
R20176 gnd.n6331 gnd.n1222 0.152939
R20177 gnd.n6327 gnd.n1222 0.152939
R20178 gnd.n6327 gnd.n6326 0.152939
R20179 gnd.n6326 gnd.n6325 0.152939
R20180 gnd.n6325 gnd.n1227 0.152939
R20181 gnd.n6321 gnd.n1227 0.152939
R20182 gnd.n6321 gnd.n6320 0.152939
R20183 gnd.n6320 gnd.n6319 0.152939
R20184 gnd.n6319 gnd.n1232 0.152939
R20185 gnd.n6315 gnd.n1232 0.152939
R20186 gnd.n6315 gnd.n6314 0.152939
R20187 gnd.n6314 gnd.n6313 0.152939
R20188 gnd.n6313 gnd.n1237 0.152939
R20189 gnd.n6309 gnd.n1237 0.152939
R20190 gnd.n6309 gnd.n6308 0.152939
R20191 gnd.n6308 gnd.n6307 0.152939
R20192 gnd.n6307 gnd.n1242 0.152939
R20193 gnd.n6215 gnd.n6214 0.152939
R20194 gnd.n6214 gnd.n6213 0.152939
R20195 gnd.n6213 gnd.n1343 0.152939
R20196 gnd.n6209 gnd.n1343 0.152939
R20197 gnd.n6209 gnd.n6208 0.152939
R20198 gnd.n6208 gnd.n6207 0.152939
R20199 gnd.n6207 gnd.n1348 0.152939
R20200 gnd.n6203 gnd.n1348 0.152939
R20201 gnd.n6203 gnd.n6202 0.152939
R20202 gnd.n6202 gnd.n6201 0.152939
R20203 gnd.n6201 gnd.n1353 0.152939
R20204 gnd.n6197 gnd.n1353 0.152939
R20205 gnd.n6197 gnd.n6196 0.152939
R20206 gnd.n6196 gnd.n6195 0.152939
R20207 gnd.n6195 gnd.n1358 0.152939
R20208 gnd.n6191 gnd.n1358 0.152939
R20209 gnd.n6191 gnd.n407 0.152939
R20210 gnd.n7371 gnd.n407 0.152939
R20211 gnd.n7371 gnd.n7370 0.152939
R20212 gnd.n7370 gnd.n7369 0.152939
R20213 gnd.n7369 gnd.n408 0.152939
R20214 gnd.n408 gnd.n375 0.152939
R20215 gnd.n7417 gnd.n375 0.152939
R20216 gnd.n7417 gnd.n7416 0.152939
R20217 gnd.n7416 gnd.n7415 0.152939
R20218 gnd.n7415 gnd.n376 0.152939
R20219 gnd.n7411 gnd.n376 0.152939
R20220 gnd.n7411 gnd.n320 0.152939
R20221 gnd.n7548 gnd.n320 0.152939
R20222 gnd.n7548 gnd.n7547 0.152939
R20223 gnd.n7547 gnd.n7546 0.152939
R20224 gnd.n7546 gnd.n321 0.152939
R20225 gnd.n7542 gnd.n321 0.152939
R20226 gnd.n7542 gnd.n7541 0.152939
R20227 gnd.n7541 gnd.n7540 0.152939
R20228 gnd.n7540 gnd.n326 0.152939
R20229 gnd.n326 gnd.n296 0.152939
R20230 gnd.n7563 gnd.n296 0.152939
R20231 gnd.n7564 gnd.n7563 0.152939
R20232 gnd.n7565 gnd.n7564 0.152939
R20233 gnd.n7565 gnd.n280 0.152939
R20234 gnd.n7579 gnd.n280 0.152939
R20235 gnd.n7580 gnd.n7579 0.152939
R20236 gnd.n7581 gnd.n7580 0.152939
R20237 gnd.n7581 gnd.n266 0.152939
R20238 gnd.n7595 gnd.n266 0.152939
R20239 gnd.n7596 gnd.n7595 0.152939
R20240 gnd.n7597 gnd.n7596 0.152939
R20241 gnd.n7597 gnd.n250 0.152939
R20242 gnd.n7611 gnd.n250 0.152939
R20243 gnd.n7612 gnd.n7611 0.152939
R20244 gnd.n7613 gnd.n7612 0.152939
R20245 gnd.n7613 gnd.n235 0.152939
R20246 gnd.n7627 gnd.n235 0.152939
R20247 gnd.n7628 gnd.n7627 0.152939
R20248 gnd.n7629 gnd.n7628 0.152939
R20249 gnd.n7629 gnd.n220 0.152939
R20250 gnd.n7643 gnd.n220 0.152939
R20251 gnd.n7644 gnd.n7643 0.152939
R20252 gnd.n7713 gnd.n7644 0.152939
R20253 gnd.n7713 gnd.n7712 0.152939
R20254 gnd.n7712 gnd.n7711 0.152939
R20255 gnd.n7711 gnd.n7645 0.152939
R20256 gnd.n7707 gnd.n7645 0.152939
R20257 gnd.n7706 gnd.n7647 0.152939
R20258 gnd.n7702 gnd.n7647 0.152939
R20259 gnd.n7702 gnd.n7701 0.152939
R20260 gnd.n7701 gnd.n7700 0.152939
R20261 gnd.n7700 gnd.n7653 0.152939
R20262 gnd.n7696 gnd.n7653 0.152939
R20263 gnd.n7696 gnd.n7695 0.152939
R20264 gnd.n7695 gnd.n7694 0.152939
R20265 gnd.n7694 gnd.n7661 0.152939
R20266 gnd.n7690 gnd.n7661 0.152939
R20267 gnd.n7690 gnd.n7689 0.152939
R20268 gnd.n7689 gnd.n7688 0.152939
R20269 gnd.n7688 gnd.n7669 0.152939
R20270 gnd.n7684 gnd.n7669 0.152939
R20271 gnd.n7684 gnd.n7683 0.152939
R20272 gnd.n7683 gnd.n7682 0.152939
R20273 gnd.n7682 gnd.n121 0.152939
R20274 gnd.n7808 gnd.n121 0.152939
R20275 gnd.n6056 gnd.n6042 0.152939
R20276 gnd.n6057 gnd.n6056 0.152939
R20277 gnd.n6059 gnd.n6057 0.152939
R20278 gnd.n6059 gnd.n6058 0.152939
R20279 gnd.n6058 gnd.n1419 0.152939
R20280 gnd.n6087 gnd.n1419 0.152939
R20281 gnd.n6088 gnd.n6087 0.152939
R20282 gnd.n6095 gnd.n6088 0.152939
R20283 gnd.n6095 gnd.n6094 0.152939
R20284 gnd.n6094 gnd.n6093 0.152939
R20285 gnd.n6093 gnd.n6089 0.152939
R20286 gnd.n6089 gnd.n1384 0.152939
R20287 gnd.n6155 gnd.n1384 0.152939
R20288 gnd.n6155 gnd.n6154 0.152939
R20289 gnd.n6154 gnd.n6153 0.152939
R20290 gnd.n6153 gnd.n1385 0.152939
R20291 gnd.n6149 gnd.n1385 0.152939
R20292 gnd.n6149 gnd.n6148 0.152939
R20293 gnd.n6148 gnd.n6147 0.152939
R20294 gnd.n6147 gnd.n6142 0.152939
R20295 gnd.n6142 gnd.n6141 0.152939
R20296 gnd.n6141 gnd.n381 0.152939
R20297 gnd.n7402 gnd.n381 0.152939
R20298 gnd.n7403 gnd.n7402 0.152939
R20299 gnd.n7405 gnd.n7403 0.152939
R20300 gnd.n7405 gnd.n7404 0.152939
R20301 gnd.n7404 gnd.n347 0.152939
R20302 gnd.n7447 gnd.n347 0.152939
R20303 gnd.n7448 gnd.n7447 0.152939
R20304 gnd.n7449 gnd.n7448 0.152939
R20305 gnd.n7449 gnd.n79 0.152939
R20306 gnd.n7857 gnd.n79 0.152939
R20307 gnd.n7857 gnd.n7856 0.152939
R20308 gnd.n7856 gnd.n81 0.152939
R20309 gnd.n7852 gnd.n81 0.152939
R20310 gnd.n7852 gnd.n7851 0.152939
R20311 gnd.n7851 gnd.n7850 0.152939
R20312 gnd.n7850 gnd.n86 0.152939
R20313 gnd.n7846 gnd.n86 0.152939
R20314 gnd.n7846 gnd.n7845 0.152939
R20315 gnd.n7845 gnd.n7844 0.152939
R20316 gnd.n7844 gnd.n91 0.152939
R20317 gnd.n7840 gnd.n91 0.152939
R20318 gnd.n7840 gnd.n7839 0.152939
R20319 gnd.n7839 gnd.n7838 0.152939
R20320 gnd.n7838 gnd.n96 0.152939
R20321 gnd.n7834 gnd.n96 0.152939
R20322 gnd.n7834 gnd.n7833 0.152939
R20323 gnd.n7833 gnd.n7832 0.152939
R20324 gnd.n7832 gnd.n101 0.152939
R20325 gnd.n7828 gnd.n101 0.152939
R20326 gnd.n7828 gnd.n7827 0.152939
R20327 gnd.n7827 gnd.n7826 0.152939
R20328 gnd.n7826 gnd.n106 0.152939
R20329 gnd.n7822 gnd.n106 0.152939
R20330 gnd.n7822 gnd.n7821 0.152939
R20331 gnd.n7821 gnd.n7820 0.152939
R20332 gnd.n7820 gnd.n111 0.152939
R20333 gnd.n7816 gnd.n111 0.152939
R20334 gnd.n7816 gnd.n7815 0.152939
R20335 gnd.n7815 gnd.n7814 0.152939
R20336 gnd.n7814 gnd.n116 0.152939
R20337 gnd.n7810 gnd.n116 0.152939
R20338 gnd.n7810 gnd.n7809 0.152939
R20339 gnd.n6041 gnd.n6040 0.151415
R20340 gnd.n4563 gnd.n4533 0.151415
R20341 gnd.n3923 gnd.n3909 0.145814
R20342 gnd.n3923 gnd.n3922 0.145814
R20343 gnd.n3205 gnd.n3204 0.0767195
R20344 gnd.n3204 gnd.n3203 0.0767195
R20345 gnd.n6459 gnd.n6458 0.063
R20346 gnd.n1518 gnd.n1342 0.063
R20347 gnd.n3771 gnd.n2374 0.0477147
R20348 gnd.n2968 gnd.n2856 0.0442063
R20349 gnd.n2969 gnd.n2968 0.0442063
R20350 gnd.n2970 gnd.n2969 0.0442063
R20351 gnd.n2970 gnd.n2845 0.0442063
R20352 gnd.n2984 gnd.n2845 0.0442063
R20353 gnd.n2985 gnd.n2984 0.0442063
R20354 gnd.n2986 gnd.n2985 0.0442063
R20355 gnd.n2986 gnd.n2832 0.0442063
R20356 gnd.n3030 gnd.n2832 0.0442063
R20357 gnd.n3031 gnd.n3030 0.0442063
R20358 gnd.n3033 gnd.n2766 0.0344674
R20359 gnd.n1597 gnd.n1478 0.0343753
R20360 gnd.n4562 gnd.n2040 0.0343753
R20361 gnd.n3053 gnd.n3052 0.0269946
R20362 gnd.n3055 gnd.n3054 0.0269946
R20363 gnd.n2761 gnd.n2759 0.0269946
R20364 gnd.n3065 gnd.n3063 0.0269946
R20365 gnd.n3064 gnd.n2740 0.0269946
R20366 gnd.n3084 gnd.n3083 0.0269946
R20367 gnd.n3086 gnd.n3085 0.0269946
R20368 gnd.n2735 gnd.n2734 0.0269946
R20369 gnd.n3096 gnd.n2730 0.0269946
R20370 gnd.n3095 gnd.n2732 0.0269946
R20371 gnd.n2731 gnd.n2713 0.0269946
R20372 gnd.n3116 gnd.n2714 0.0269946
R20373 gnd.n3115 gnd.n2715 0.0269946
R20374 gnd.n3149 gnd.n2690 0.0269946
R20375 gnd.n3151 gnd.n3150 0.0269946
R20376 gnd.n3152 gnd.n2637 0.0269946
R20377 gnd.n2685 gnd.n2638 0.0269946
R20378 gnd.n2687 gnd.n2639 0.0269946
R20379 gnd.n3162 gnd.n3161 0.0269946
R20380 gnd.n3164 gnd.n3163 0.0269946
R20381 gnd.n3165 gnd.n2659 0.0269946
R20382 gnd.n3167 gnd.n2660 0.0269946
R20383 gnd.n3170 gnd.n2661 0.0269946
R20384 gnd.n3173 gnd.n3172 0.0269946
R20385 gnd.n3175 gnd.n3174 0.0269946
R20386 gnd.n3240 gnd.n2548 0.0269946
R20387 gnd.n3242 gnd.n3241 0.0269946
R20388 gnd.n3251 gnd.n2541 0.0269946
R20389 gnd.n3253 gnd.n3252 0.0269946
R20390 gnd.n3254 gnd.n2539 0.0269946
R20391 gnd.n3261 gnd.n3257 0.0269946
R20392 gnd.n3260 gnd.n3259 0.0269946
R20393 gnd.n3258 gnd.n2518 0.0269946
R20394 gnd.n3283 gnd.n2519 0.0269946
R20395 gnd.n3282 gnd.n2520 0.0269946
R20396 gnd.n3325 gnd.n2493 0.0269946
R20397 gnd.n3327 gnd.n3326 0.0269946
R20398 gnd.n3336 gnd.n2486 0.0269946
R20399 gnd.n3338 gnd.n3337 0.0269946
R20400 gnd.n3339 gnd.n2484 0.0269946
R20401 gnd.n3346 gnd.n3342 0.0269946
R20402 gnd.n3345 gnd.n3344 0.0269946
R20403 gnd.n3343 gnd.n2463 0.0269946
R20404 gnd.n3368 gnd.n2464 0.0269946
R20405 gnd.n3367 gnd.n2465 0.0269946
R20406 gnd.n3414 gnd.n2439 0.0269946
R20407 gnd.n3416 gnd.n3415 0.0269946
R20408 gnd.n3425 gnd.n2432 0.0269946
R20409 gnd.n3684 gnd.n2430 0.0269946
R20410 gnd.n3689 gnd.n3687 0.0269946
R20411 gnd.n3688 gnd.n2411 0.0269946
R20412 gnd.n3713 gnd.n3712 0.0269946
R20413 gnd.n1520 gnd.n1518 0.0245515
R20414 gnd.n6458 gnd.n1116 0.0245515
R20415 gnd.n3033 gnd.n3032 0.0202011
R20416 gnd.n1520 gnd.n1519 0.0174377
R20417 gnd.n1519 gnd.n1515 0.0174377
R20418 gnd.n1529 gnd.n1515 0.0174377
R20419 gnd.n1529 gnd.n1528 0.0174377
R20420 gnd.n1528 gnd.n1516 0.0174377
R20421 gnd.n1516 gnd.n1511 0.0174377
R20422 gnd.n1537 gnd.n1511 0.0174377
R20423 gnd.n1539 gnd.n1537 0.0174377
R20424 gnd.n1539 gnd.n1538 0.0174377
R20425 gnd.n1538 gnd.n1508 0.0174377
R20426 gnd.n1548 gnd.n1508 0.0174377
R20427 gnd.n1548 gnd.n1547 0.0174377
R20428 gnd.n1547 gnd.n1509 0.0174377
R20429 gnd.n1509 gnd.n1504 0.0174377
R20430 gnd.n1556 gnd.n1504 0.0174377
R20431 gnd.n1558 gnd.n1556 0.0174377
R20432 gnd.n1558 gnd.n1557 0.0174377
R20433 gnd.n1557 gnd.n1501 0.0174377
R20434 gnd.n1567 gnd.n1501 0.0174377
R20435 gnd.n1567 gnd.n1566 0.0174377
R20436 gnd.n1566 gnd.n1502 0.0174377
R20437 gnd.n1502 gnd.n1497 0.0174377
R20438 gnd.n1575 gnd.n1497 0.0174377
R20439 gnd.n1576 gnd.n1575 0.0174377
R20440 gnd.n1576 gnd.n1495 0.0174377
R20441 gnd.n1581 gnd.n1495 0.0174377
R20442 gnd.n1583 gnd.n1581 0.0174377
R20443 gnd.n1583 gnd.n1582 0.0174377
R20444 gnd.n1582 gnd.n1491 0.0174377
R20445 gnd.n1592 gnd.n1491 0.0174377
R20446 gnd.n1592 gnd.n1591 0.0174377
R20447 gnd.n1591 gnd.n1484 0.0174377
R20448 gnd.n1484 gnd.n1483 0.0174377
R20449 gnd.n1596 gnd.n1483 0.0174377
R20450 gnd.n1597 gnd.n1596 0.0174377
R20451 gnd.n1989 gnd.n1116 0.0174377
R20452 gnd.n1991 gnd.n1989 0.0174377
R20453 gnd.n5601 gnd.n1991 0.0174377
R20454 gnd.n5601 gnd.n5600 0.0174377
R20455 gnd.n5600 gnd.n1992 0.0174377
R20456 gnd.n5597 gnd.n1992 0.0174377
R20457 gnd.n5597 gnd.n5596 0.0174377
R20458 gnd.n5596 gnd.n1997 0.0174377
R20459 gnd.n5593 gnd.n1997 0.0174377
R20460 gnd.n5593 gnd.n5592 0.0174377
R20461 gnd.n5592 gnd.n2002 0.0174377
R20462 gnd.n5589 gnd.n2002 0.0174377
R20463 gnd.n5589 gnd.n5588 0.0174377
R20464 gnd.n5588 gnd.n2006 0.0174377
R20465 gnd.n5585 gnd.n2006 0.0174377
R20466 gnd.n5585 gnd.n5584 0.0174377
R20467 gnd.n5584 gnd.n2010 0.0174377
R20468 gnd.n5581 gnd.n2010 0.0174377
R20469 gnd.n5581 gnd.n5580 0.0174377
R20470 gnd.n5580 gnd.n2014 0.0174377
R20471 gnd.n5577 gnd.n2014 0.0174377
R20472 gnd.n5577 gnd.n5576 0.0174377
R20473 gnd.n5576 gnd.n2020 0.0174377
R20474 gnd.n5573 gnd.n2020 0.0174377
R20475 gnd.n5573 gnd.n5572 0.0174377
R20476 gnd.n5572 gnd.n2024 0.0174377
R20477 gnd.n5569 gnd.n2024 0.0174377
R20478 gnd.n5569 gnd.n5568 0.0174377
R20479 gnd.n5568 gnd.n2028 0.0174377
R20480 gnd.n5565 gnd.n2028 0.0174377
R20481 gnd.n5565 gnd.n5564 0.0174377
R20482 gnd.n5564 gnd.n2034 0.0174377
R20483 gnd.n5561 gnd.n2034 0.0174377
R20484 gnd.n5561 gnd.n5560 0.0174377
R20485 gnd.n5560 gnd.n2040 0.0174377
R20486 gnd.n3032 gnd.n3031 0.0148637
R20487 gnd.n3682 gnd.n3426 0.0144266
R20488 gnd.n3683 gnd.n3682 0.0130679
R20489 gnd.n3052 gnd.n2766 0.00797283
R20490 gnd.n3054 gnd.n3053 0.00797283
R20491 gnd.n3055 gnd.n2761 0.00797283
R20492 gnd.n3063 gnd.n2759 0.00797283
R20493 gnd.n3065 gnd.n3064 0.00797283
R20494 gnd.n3083 gnd.n2740 0.00797283
R20495 gnd.n3085 gnd.n3084 0.00797283
R20496 gnd.n3086 gnd.n2735 0.00797283
R20497 gnd.n2734 gnd.n2730 0.00797283
R20498 gnd.n3096 gnd.n3095 0.00797283
R20499 gnd.n2732 gnd.n2731 0.00797283
R20500 gnd.n2714 gnd.n2713 0.00797283
R20501 gnd.n3116 gnd.n3115 0.00797283
R20502 gnd.n2715 gnd.n2690 0.00797283
R20503 gnd.n3150 gnd.n3149 0.00797283
R20504 gnd.n3152 gnd.n3151 0.00797283
R20505 gnd.n2685 gnd.n2637 0.00797283
R20506 gnd.n2687 gnd.n2638 0.00797283
R20507 gnd.n3161 gnd.n2639 0.00797283
R20508 gnd.n3163 gnd.n3162 0.00797283
R20509 gnd.n3165 gnd.n3164 0.00797283
R20510 gnd.n3167 gnd.n2659 0.00797283
R20511 gnd.n3170 gnd.n2660 0.00797283
R20512 gnd.n3172 gnd.n2661 0.00797283
R20513 gnd.n3175 gnd.n3173 0.00797283
R20514 gnd.n3174 gnd.n2548 0.00797283
R20515 gnd.n3242 gnd.n3240 0.00797283
R20516 gnd.n3241 gnd.n2541 0.00797283
R20517 gnd.n3252 gnd.n3251 0.00797283
R20518 gnd.n3254 gnd.n3253 0.00797283
R20519 gnd.n3257 gnd.n2539 0.00797283
R20520 gnd.n3261 gnd.n3260 0.00797283
R20521 gnd.n3259 gnd.n3258 0.00797283
R20522 gnd.n2519 gnd.n2518 0.00797283
R20523 gnd.n3283 gnd.n3282 0.00797283
R20524 gnd.n2520 gnd.n2493 0.00797283
R20525 gnd.n3327 gnd.n3325 0.00797283
R20526 gnd.n3326 gnd.n2486 0.00797283
R20527 gnd.n3337 gnd.n3336 0.00797283
R20528 gnd.n3339 gnd.n3338 0.00797283
R20529 gnd.n3342 gnd.n2484 0.00797283
R20530 gnd.n3346 gnd.n3345 0.00797283
R20531 gnd.n3344 gnd.n3343 0.00797283
R20532 gnd.n2464 gnd.n2463 0.00797283
R20533 gnd.n3368 gnd.n3367 0.00797283
R20534 gnd.n2465 gnd.n2439 0.00797283
R20535 gnd.n3416 gnd.n3414 0.00797283
R20536 gnd.n3415 gnd.n2432 0.00797283
R20537 gnd.n3426 gnd.n3425 0.00797283
R20538 gnd.n3684 gnd.n3683 0.00797283
R20539 gnd.n3687 gnd.n2430 0.00797283
R20540 gnd.n3689 gnd.n3688 0.00797283
R20541 gnd.n3712 gnd.n2411 0.00797283
R20542 gnd.n3713 gnd.n2374 0.00797283
R20543 gnd.n337 gnd.n321 0.00433921
R20544 gnd.n4328 gnd.n4327 0.00433921
R20545 gnd.n6041 gnd.n1478 0.000838753
R20546 gnd.n4563 gnd.n4562 0.000838753
R20547 a_n1808_13878.n16 a_n1808_13878.n0 98.9633
R20548 a_n1808_13878.n3 a_n1808_13878.n1 98.7517
R20549 a_n1808_13878.n5 a_n1808_13878.n4 98.6055
R20550 a_n1808_13878.n3 a_n1808_13878.n2 98.6055
R20551 a_n1808_13878.n17 a_n1808_13878.n16 98.6054
R20552 a_n1808_13878.n15 a_n1808_13878.n14 98.6054
R20553 a_n1808_13878.n7 a_n1808_13878.t1 74.6477
R20554 a_n1808_13878.n12 a_n1808_13878.t2 74.2899
R20555 a_n1808_13878.n9 a_n1808_13878.t3 74.2899
R20556 a_n1808_13878.n8 a_n1808_13878.t0 74.2899
R20557 a_n1808_13878.n11 a_n1808_13878.n10 70.6783
R20558 a_n1808_13878.n7 a_n1808_13878.n6 70.6783
R20559 a_n1808_13878.n13 a_n1808_13878.n5 13.5694
R20560 a_n1808_13878.n15 a_n1808_13878.n13 11.5762
R20561 a_n1808_13878.n13 a_n1808_13878.n12 6.2408
R20562 a_n1808_13878.n14 a_n1808_13878.t15 3.61217
R20563 a_n1808_13878.n14 a_n1808_13878.t16 3.61217
R20564 a_n1808_13878.n0 a_n1808_13878.t13 3.61217
R20565 a_n1808_13878.n0 a_n1808_13878.t17 3.61217
R20566 a_n1808_13878.n10 a_n1808_13878.t6 3.61217
R20567 a_n1808_13878.n10 a_n1808_13878.t7 3.61217
R20568 a_n1808_13878.n6 a_n1808_13878.t4 3.61217
R20569 a_n1808_13878.n6 a_n1808_13878.t5 3.61217
R20570 a_n1808_13878.n4 a_n1808_13878.t12 3.61217
R20571 a_n1808_13878.n4 a_n1808_13878.t19 3.61217
R20572 a_n1808_13878.n2 a_n1808_13878.t14 3.61217
R20573 a_n1808_13878.n2 a_n1808_13878.t9 3.61217
R20574 a_n1808_13878.n1 a_n1808_13878.t8 3.61217
R20575 a_n1808_13878.n1 a_n1808_13878.t10 3.61217
R20576 a_n1808_13878.t18 a_n1808_13878.n17 3.61217
R20577 a_n1808_13878.n17 a_n1808_13878.t11 3.61217
R20578 a_n1808_13878.n8 a_n1808_13878.n7 0.358259
R20579 a_n1808_13878.n11 a_n1808_13878.n9 0.358259
R20580 a_n1808_13878.n12 a_n1808_13878.n11 0.358259
R20581 a_n1808_13878.n16 a_n1808_13878.n15 0.358259
R20582 a_n1808_13878.n5 a_n1808_13878.n3 0.146627
R20583 a_n1808_13878.n9 a_n1808_13878.n8 0.101793
R20584 outputibias.n27 outputibias.n1 289.615
R20585 outputibias.n58 outputibias.n32 289.615
R20586 outputibias.n90 outputibias.n64 289.615
R20587 outputibias.n122 outputibias.n96 289.615
R20588 outputibias.n28 outputibias.n27 185
R20589 outputibias.n26 outputibias.n25 185
R20590 outputibias.n5 outputibias.n4 185
R20591 outputibias.n20 outputibias.n19 185
R20592 outputibias.n18 outputibias.n17 185
R20593 outputibias.n9 outputibias.n8 185
R20594 outputibias.n12 outputibias.n11 185
R20595 outputibias.n59 outputibias.n58 185
R20596 outputibias.n57 outputibias.n56 185
R20597 outputibias.n36 outputibias.n35 185
R20598 outputibias.n51 outputibias.n50 185
R20599 outputibias.n49 outputibias.n48 185
R20600 outputibias.n40 outputibias.n39 185
R20601 outputibias.n43 outputibias.n42 185
R20602 outputibias.n91 outputibias.n90 185
R20603 outputibias.n89 outputibias.n88 185
R20604 outputibias.n68 outputibias.n67 185
R20605 outputibias.n83 outputibias.n82 185
R20606 outputibias.n81 outputibias.n80 185
R20607 outputibias.n72 outputibias.n71 185
R20608 outputibias.n75 outputibias.n74 185
R20609 outputibias.n123 outputibias.n122 185
R20610 outputibias.n121 outputibias.n120 185
R20611 outputibias.n100 outputibias.n99 185
R20612 outputibias.n115 outputibias.n114 185
R20613 outputibias.n113 outputibias.n112 185
R20614 outputibias.n104 outputibias.n103 185
R20615 outputibias.n107 outputibias.n106 185
R20616 outputibias.n0 outputibias.t8 178.945
R20617 outputibias.n133 outputibias.t9 177.018
R20618 outputibias.n132 outputibias.t11 177.018
R20619 outputibias.n0 outputibias.t10 177.018
R20620 outputibias.t5 outputibias.n10 147.661
R20621 outputibias.t3 outputibias.n41 147.661
R20622 outputibias.t1 outputibias.n73 147.661
R20623 outputibias.t7 outputibias.n105 147.661
R20624 outputibias.n128 outputibias.t4 132.363
R20625 outputibias.n128 outputibias.t2 130.436
R20626 outputibias.n129 outputibias.t0 130.436
R20627 outputibias.n130 outputibias.t6 130.436
R20628 outputibias.n27 outputibias.n26 104.615
R20629 outputibias.n26 outputibias.n4 104.615
R20630 outputibias.n19 outputibias.n4 104.615
R20631 outputibias.n19 outputibias.n18 104.615
R20632 outputibias.n18 outputibias.n8 104.615
R20633 outputibias.n11 outputibias.n8 104.615
R20634 outputibias.n58 outputibias.n57 104.615
R20635 outputibias.n57 outputibias.n35 104.615
R20636 outputibias.n50 outputibias.n35 104.615
R20637 outputibias.n50 outputibias.n49 104.615
R20638 outputibias.n49 outputibias.n39 104.615
R20639 outputibias.n42 outputibias.n39 104.615
R20640 outputibias.n90 outputibias.n89 104.615
R20641 outputibias.n89 outputibias.n67 104.615
R20642 outputibias.n82 outputibias.n67 104.615
R20643 outputibias.n82 outputibias.n81 104.615
R20644 outputibias.n81 outputibias.n71 104.615
R20645 outputibias.n74 outputibias.n71 104.615
R20646 outputibias.n122 outputibias.n121 104.615
R20647 outputibias.n121 outputibias.n99 104.615
R20648 outputibias.n114 outputibias.n99 104.615
R20649 outputibias.n114 outputibias.n113 104.615
R20650 outputibias.n113 outputibias.n103 104.615
R20651 outputibias.n106 outputibias.n103 104.615
R20652 outputibias.n63 outputibias.n31 95.6354
R20653 outputibias.n63 outputibias.n62 94.6732
R20654 outputibias.n95 outputibias.n94 94.6732
R20655 outputibias.n127 outputibias.n126 94.6732
R20656 outputibias.n11 outputibias.t5 52.3082
R20657 outputibias.n42 outputibias.t3 52.3082
R20658 outputibias.n74 outputibias.t1 52.3082
R20659 outputibias.n106 outputibias.t7 52.3082
R20660 outputibias.n12 outputibias.n10 15.6674
R20661 outputibias.n43 outputibias.n41 15.6674
R20662 outputibias.n75 outputibias.n73 15.6674
R20663 outputibias.n107 outputibias.n105 15.6674
R20664 outputibias.n13 outputibias.n9 12.8005
R20665 outputibias.n44 outputibias.n40 12.8005
R20666 outputibias.n76 outputibias.n72 12.8005
R20667 outputibias.n108 outputibias.n104 12.8005
R20668 outputibias.n17 outputibias.n16 12.0247
R20669 outputibias.n48 outputibias.n47 12.0247
R20670 outputibias.n80 outputibias.n79 12.0247
R20671 outputibias.n112 outputibias.n111 12.0247
R20672 outputibias.n20 outputibias.n7 11.249
R20673 outputibias.n51 outputibias.n38 11.249
R20674 outputibias.n83 outputibias.n70 11.249
R20675 outputibias.n115 outputibias.n102 11.249
R20676 outputibias.n21 outputibias.n5 10.4732
R20677 outputibias.n52 outputibias.n36 10.4732
R20678 outputibias.n84 outputibias.n68 10.4732
R20679 outputibias.n116 outputibias.n100 10.4732
R20680 outputibias.n25 outputibias.n24 9.69747
R20681 outputibias.n56 outputibias.n55 9.69747
R20682 outputibias.n88 outputibias.n87 9.69747
R20683 outputibias.n120 outputibias.n119 9.69747
R20684 outputibias.n31 outputibias.n30 9.45567
R20685 outputibias.n62 outputibias.n61 9.45567
R20686 outputibias.n94 outputibias.n93 9.45567
R20687 outputibias.n126 outputibias.n125 9.45567
R20688 outputibias.n30 outputibias.n29 9.3005
R20689 outputibias.n3 outputibias.n2 9.3005
R20690 outputibias.n24 outputibias.n23 9.3005
R20691 outputibias.n22 outputibias.n21 9.3005
R20692 outputibias.n7 outputibias.n6 9.3005
R20693 outputibias.n16 outputibias.n15 9.3005
R20694 outputibias.n14 outputibias.n13 9.3005
R20695 outputibias.n61 outputibias.n60 9.3005
R20696 outputibias.n34 outputibias.n33 9.3005
R20697 outputibias.n55 outputibias.n54 9.3005
R20698 outputibias.n53 outputibias.n52 9.3005
R20699 outputibias.n38 outputibias.n37 9.3005
R20700 outputibias.n47 outputibias.n46 9.3005
R20701 outputibias.n45 outputibias.n44 9.3005
R20702 outputibias.n93 outputibias.n92 9.3005
R20703 outputibias.n66 outputibias.n65 9.3005
R20704 outputibias.n87 outputibias.n86 9.3005
R20705 outputibias.n85 outputibias.n84 9.3005
R20706 outputibias.n70 outputibias.n69 9.3005
R20707 outputibias.n79 outputibias.n78 9.3005
R20708 outputibias.n77 outputibias.n76 9.3005
R20709 outputibias.n125 outputibias.n124 9.3005
R20710 outputibias.n98 outputibias.n97 9.3005
R20711 outputibias.n119 outputibias.n118 9.3005
R20712 outputibias.n117 outputibias.n116 9.3005
R20713 outputibias.n102 outputibias.n101 9.3005
R20714 outputibias.n111 outputibias.n110 9.3005
R20715 outputibias.n109 outputibias.n108 9.3005
R20716 outputibias.n28 outputibias.n3 8.92171
R20717 outputibias.n59 outputibias.n34 8.92171
R20718 outputibias.n91 outputibias.n66 8.92171
R20719 outputibias.n123 outputibias.n98 8.92171
R20720 outputibias.n29 outputibias.n1 8.14595
R20721 outputibias.n60 outputibias.n32 8.14595
R20722 outputibias.n92 outputibias.n64 8.14595
R20723 outputibias.n124 outputibias.n96 8.14595
R20724 outputibias.n31 outputibias.n1 5.81868
R20725 outputibias.n62 outputibias.n32 5.81868
R20726 outputibias.n94 outputibias.n64 5.81868
R20727 outputibias.n126 outputibias.n96 5.81868
R20728 outputibias.n131 outputibias.n130 5.20947
R20729 outputibias.n29 outputibias.n28 5.04292
R20730 outputibias.n60 outputibias.n59 5.04292
R20731 outputibias.n92 outputibias.n91 5.04292
R20732 outputibias.n124 outputibias.n123 5.04292
R20733 outputibias.n131 outputibias.n127 4.42209
R20734 outputibias.n14 outputibias.n10 4.38594
R20735 outputibias.n45 outputibias.n41 4.38594
R20736 outputibias.n77 outputibias.n73 4.38594
R20737 outputibias.n109 outputibias.n105 4.38594
R20738 outputibias.n132 outputibias.n131 4.28454
R20739 outputibias.n25 outputibias.n3 4.26717
R20740 outputibias.n56 outputibias.n34 4.26717
R20741 outputibias.n88 outputibias.n66 4.26717
R20742 outputibias.n120 outputibias.n98 4.26717
R20743 outputibias.n24 outputibias.n5 3.49141
R20744 outputibias.n55 outputibias.n36 3.49141
R20745 outputibias.n87 outputibias.n68 3.49141
R20746 outputibias.n119 outputibias.n100 3.49141
R20747 outputibias.n21 outputibias.n20 2.71565
R20748 outputibias.n52 outputibias.n51 2.71565
R20749 outputibias.n84 outputibias.n83 2.71565
R20750 outputibias.n116 outputibias.n115 2.71565
R20751 outputibias.n17 outputibias.n7 1.93989
R20752 outputibias.n48 outputibias.n38 1.93989
R20753 outputibias.n80 outputibias.n70 1.93989
R20754 outputibias.n112 outputibias.n102 1.93989
R20755 outputibias.n130 outputibias.n129 1.9266
R20756 outputibias.n129 outputibias.n128 1.9266
R20757 outputibias.n133 outputibias.n132 1.92658
R20758 outputibias.n134 outputibias.n133 1.29913
R20759 outputibias.n16 outputibias.n9 1.16414
R20760 outputibias.n47 outputibias.n40 1.16414
R20761 outputibias.n79 outputibias.n72 1.16414
R20762 outputibias.n111 outputibias.n104 1.16414
R20763 outputibias.n127 outputibias.n95 0.962709
R20764 outputibias.n95 outputibias.n63 0.962709
R20765 outputibias.n13 outputibias.n12 0.388379
R20766 outputibias.n44 outputibias.n43 0.388379
R20767 outputibias.n76 outputibias.n75 0.388379
R20768 outputibias.n108 outputibias.n107 0.388379
R20769 outputibias.n134 outputibias.n0 0.337251
R20770 outputibias outputibias.n134 0.302375
R20771 outputibias.n30 outputibias.n2 0.155672
R20772 outputibias.n23 outputibias.n2 0.155672
R20773 outputibias.n23 outputibias.n22 0.155672
R20774 outputibias.n22 outputibias.n6 0.155672
R20775 outputibias.n15 outputibias.n6 0.155672
R20776 outputibias.n15 outputibias.n14 0.155672
R20777 outputibias.n61 outputibias.n33 0.155672
R20778 outputibias.n54 outputibias.n33 0.155672
R20779 outputibias.n54 outputibias.n53 0.155672
R20780 outputibias.n53 outputibias.n37 0.155672
R20781 outputibias.n46 outputibias.n37 0.155672
R20782 outputibias.n46 outputibias.n45 0.155672
R20783 outputibias.n93 outputibias.n65 0.155672
R20784 outputibias.n86 outputibias.n65 0.155672
R20785 outputibias.n86 outputibias.n85 0.155672
R20786 outputibias.n85 outputibias.n69 0.155672
R20787 outputibias.n78 outputibias.n69 0.155672
R20788 outputibias.n78 outputibias.n77 0.155672
R20789 outputibias.n125 outputibias.n97 0.155672
R20790 outputibias.n118 outputibias.n97 0.155672
R20791 outputibias.n118 outputibias.n117 0.155672
R20792 outputibias.n117 outputibias.n101 0.155672
R20793 outputibias.n110 outputibias.n101 0.155672
R20794 outputibias.n110 outputibias.n109 0.155672
R20795 plus.n76 plus.t11 250.337
R20796 plus.n15 plus.t14 250.337
R20797 plus.n124 plus.t1 243.97
R20798 plus.n120 plus.t24 231.093
R20799 plus.n59 plus.t20 231.093
R20800 plus.n124 plus.n123 223.454
R20801 plus.n126 plus.n125 223.454
R20802 plus.n77 plus.t5 187.445
R20803 plus.n74 plus.t22 187.445
R20804 plus.n72 plus.t21 187.445
R20805 plus.n89 plus.t16 187.445
R20806 plus.n95 plus.t17 187.445
R20807 plus.n68 plus.t13 187.445
R20808 plus.n66 plus.t15 187.445
R20809 plus.n107 plus.t10 187.445
R20810 plus.n113 plus.t26 187.445
R20811 plus.n62 plus.t28 187.445
R20812 plus.n1 plus.t23 187.445
R20813 plus.n52 plus.t6 187.445
R20814 plus.n46 plus.t12 187.445
R20815 plus.n5 plus.t8 187.445
R20816 plus.n7 plus.t7 187.445
R20817 plus.n34 plus.t19 187.445
R20818 plus.n28 plus.t18 187.445
R20819 plus.n11 plus.t27 187.445
R20820 plus.n13 plus.t25 187.445
R20821 plus.n16 plus.t9 187.445
R20822 plus.n121 plus.n120 161.3
R20823 plus.n119 plus.n61 161.3
R20824 plus.n118 plus.n117 161.3
R20825 plus.n116 plus.n115 161.3
R20826 plus.n114 plus.n63 161.3
R20827 plus.n112 plus.n111 161.3
R20828 plus.n110 plus.n64 161.3
R20829 plus.n109 plus.n108 161.3
R20830 plus.n106 plus.n65 161.3
R20831 plus.n105 plus.n104 161.3
R20832 plus.n103 plus.n102 161.3
R20833 plus.n101 plus.n67 161.3
R20834 plus.n100 plus.n99 161.3
R20835 plus.n98 plus.n97 161.3
R20836 plus.n96 plus.n69 161.3
R20837 plus.n94 plus.n93 161.3
R20838 plus.n92 plus.n70 161.3
R20839 plus.n91 plus.n90 161.3
R20840 plus.n88 plus.n71 161.3
R20841 plus.n87 plus.n86 161.3
R20842 plus.n85 plus.n84 161.3
R20843 plus.n83 plus.n73 161.3
R20844 plus.n82 plus.n81 161.3
R20845 plus.n80 plus.n79 161.3
R20846 plus.n78 plus.n75 161.3
R20847 plus.n17 plus.n14 161.3
R20848 plus.n19 plus.n18 161.3
R20849 plus.n21 plus.n20 161.3
R20850 plus.n22 plus.n12 161.3
R20851 plus.n24 plus.n23 161.3
R20852 plus.n26 plus.n25 161.3
R20853 plus.n27 plus.n10 161.3
R20854 plus.n30 plus.n29 161.3
R20855 plus.n31 plus.n9 161.3
R20856 plus.n33 plus.n32 161.3
R20857 plus.n35 plus.n8 161.3
R20858 plus.n37 plus.n36 161.3
R20859 plus.n39 plus.n38 161.3
R20860 plus.n40 plus.n6 161.3
R20861 plus.n42 plus.n41 161.3
R20862 plus.n44 plus.n43 161.3
R20863 plus.n45 plus.n4 161.3
R20864 plus.n48 plus.n47 161.3
R20865 plus.n49 plus.n3 161.3
R20866 plus.n51 plus.n50 161.3
R20867 plus.n53 plus.n2 161.3
R20868 plus.n55 plus.n54 161.3
R20869 plus.n57 plus.n56 161.3
R20870 plus.n58 plus.n0 161.3
R20871 plus.n60 plus.n59 161.3
R20872 plus.n88 plus.n87 56.5617
R20873 plus.n97 plus.n96 56.5617
R20874 plus.n106 plus.n105 56.5617
R20875 plus.n45 plus.n44 56.5617
R20876 plus.n36 plus.n35 56.5617
R20877 plus.n27 plus.n26 56.5617
R20878 plus.n79 plus.n78 56.5617
R20879 plus.n115 plus.n114 56.5617
R20880 plus.n54 plus.n53 56.5617
R20881 plus.n18 plus.n17 56.5617
R20882 plus.n119 plus.n118 50.2647
R20883 plus.n58 plus.n57 50.2647
R20884 plus.n84 plus.n83 46.3896
R20885 plus.n108 plus.n64 46.3896
R20886 plus.n47 plus.n3 46.3896
R20887 plus.n23 plus.n22 46.3896
R20888 plus.n76 plus.n75 43.1929
R20889 plus.n15 plus.n14 43.1929
R20890 plus.n94 plus.n70 42.5146
R20891 plus.n101 plus.n100 42.5146
R20892 plus.n40 plus.n39 42.5146
R20893 plus.n33 plus.n9 42.5146
R20894 plus.n77 plus.n76 40.6041
R20895 plus.n16 plus.n15 40.6041
R20896 plus.n90 plus.n70 38.6395
R20897 plus.n102 plus.n101 38.6395
R20898 plus.n41 plus.n40 38.6395
R20899 plus.n29 plus.n9 38.6395
R20900 plus.n122 plus.n121 35.2031
R20901 plus.n83 plus.n82 34.7644
R20902 plus.n112 plus.n64 34.7644
R20903 plus.n51 plus.n3 34.7644
R20904 plus.n22 plus.n21 34.7644
R20905 plus.n79 plus.n74 21.8872
R20906 plus.n114 plus.n113 21.8872
R20907 plus.n53 plus.n52 21.8872
R20908 plus.n18 plus.n13 21.8872
R20909 plus.n89 plus.n88 19.9199
R20910 plus.n105 plus.n66 19.9199
R20911 plus.n44 plus.n5 19.9199
R20912 plus.n28 plus.n27 19.9199
R20913 plus.n123 plus.t2 19.8005
R20914 plus.n123 plus.t4 19.8005
R20915 plus.n125 plus.t3 19.8005
R20916 plus.n125 plus.t0 19.8005
R20917 plus.n96 plus.n95 17.9525
R20918 plus.n97 plus.n68 17.9525
R20919 plus.n36 plus.n7 17.9525
R20920 plus.n35 plus.n34 17.9525
R20921 plus.n87 plus.n72 15.9852
R20922 plus.n107 plus.n106 15.9852
R20923 plus.n46 plus.n45 15.9852
R20924 plus.n26 plus.n11 15.9852
R20925 plus plus.n127 15.3578
R20926 plus.n78 plus.n77 14.0178
R20927 plus.n115 plus.n62 14.0178
R20928 plus.n54 plus.n1 14.0178
R20929 plus.n17 plus.n16 14.0178
R20930 plus.n122 plus.n60 11.9342
R20931 plus.n118 plus.n62 10.575
R20932 plus.n57 plus.n1 10.575
R20933 plus.n120 plus.n119 9.49444
R20934 plus.n59 plus.n58 9.49444
R20935 plus.n84 plus.n72 8.60764
R20936 plus.n108 plus.n107 8.60764
R20937 plus.n47 plus.n46 8.60764
R20938 plus.n23 plus.n11 8.60764
R20939 plus.n95 plus.n94 6.6403
R20940 plus.n100 plus.n68 6.6403
R20941 plus.n39 plus.n7 6.6403
R20942 plus.n34 plus.n33 6.6403
R20943 plus.n127 plus.n126 5.40567
R20944 plus.n90 plus.n89 4.67295
R20945 plus.n102 plus.n66 4.67295
R20946 plus.n41 plus.n5 4.67295
R20947 plus.n29 plus.n28 4.67295
R20948 plus.n82 plus.n74 2.7056
R20949 plus.n113 plus.n112 2.7056
R20950 plus.n52 plus.n51 2.7056
R20951 plus.n21 plus.n13 2.7056
R20952 plus.n127 plus.n122 1.188
R20953 plus.n126 plus.n124 0.716017
R20954 plus.n80 plus.n75 0.189894
R20955 plus.n81 plus.n80 0.189894
R20956 plus.n81 plus.n73 0.189894
R20957 plus.n85 plus.n73 0.189894
R20958 plus.n86 plus.n85 0.189894
R20959 plus.n86 plus.n71 0.189894
R20960 plus.n91 plus.n71 0.189894
R20961 plus.n92 plus.n91 0.189894
R20962 plus.n93 plus.n92 0.189894
R20963 plus.n93 plus.n69 0.189894
R20964 plus.n98 plus.n69 0.189894
R20965 plus.n99 plus.n98 0.189894
R20966 plus.n99 plus.n67 0.189894
R20967 plus.n103 plus.n67 0.189894
R20968 plus.n104 plus.n103 0.189894
R20969 plus.n104 plus.n65 0.189894
R20970 plus.n109 plus.n65 0.189894
R20971 plus.n110 plus.n109 0.189894
R20972 plus.n111 plus.n110 0.189894
R20973 plus.n111 plus.n63 0.189894
R20974 plus.n116 plus.n63 0.189894
R20975 plus.n117 plus.n116 0.189894
R20976 plus.n117 plus.n61 0.189894
R20977 plus.n121 plus.n61 0.189894
R20978 plus.n60 plus.n0 0.189894
R20979 plus.n56 plus.n0 0.189894
R20980 plus.n56 plus.n55 0.189894
R20981 plus.n55 plus.n2 0.189894
R20982 plus.n50 plus.n2 0.189894
R20983 plus.n50 plus.n49 0.189894
R20984 plus.n49 plus.n48 0.189894
R20985 plus.n48 plus.n4 0.189894
R20986 plus.n43 plus.n4 0.189894
R20987 plus.n43 plus.n42 0.189894
R20988 plus.n42 plus.n6 0.189894
R20989 plus.n38 plus.n6 0.189894
R20990 plus.n38 plus.n37 0.189894
R20991 plus.n37 plus.n8 0.189894
R20992 plus.n32 plus.n8 0.189894
R20993 plus.n32 plus.n31 0.189894
R20994 plus.n31 plus.n30 0.189894
R20995 plus.n30 plus.n10 0.189894
R20996 plus.n25 plus.n10 0.189894
R20997 plus.n25 plus.n24 0.189894
R20998 plus.n24 plus.n12 0.189894
R20999 plus.n20 plus.n12 0.189894
R21000 plus.n20 plus.n19 0.189894
R21001 plus.n19 plus.n14 0.189894
R21002 a_n3827_n3924.n4 a_n3827_n3924.t23 214.938
R21003 a_n3827_n3924.n8 a_n3827_n3924.t9 214.409
R21004 a_n3827_n3924.n8 a_n3827_n3924.t55 214.321
R21005 a_n3827_n3924.n7 a_n3827_n3924.t3 214.321
R21006 a_n3827_n3924.n7 a_n3827_n3924.t18 214.321
R21007 a_n3827_n3924.n6 a_n3827_n3924.t5 214.321
R21008 a_n3827_n3924.n6 a_n3827_n3924.t56 214.321
R21009 a_n3827_n3924.n5 a_n3827_n3924.t16 214.321
R21010 a_n3827_n3924.n5 a_n3827_n3924.t13 214.321
R21011 a_n3827_n3924.n4 a_n3827_n3924.t28 214.321
R21012 a_n3827_n3924.n3 a_n3827_n3924.t46 55.8337
R21013 a_n3827_n3924.n3 a_n3827_n3924.t1 55.8337
R21014 a_n3827_n3924.n10 a_n3827_n3924.t10 55.8337
R21015 a_n3827_n3924.n2 a_n3827_n3924.t43 55.8335
R21016 a_n3827_n3924.n1 a_n3827_n3924.t25 55.8335
R21017 a_n3827_n3924.n0 a_n3827_n3924.t24 55.8335
R21018 a_n3827_n3924.n0 a_n3827_n3924.t47 55.8335
R21019 a_n3827_n3924.n12 a_n3827_n3924.t35 55.8335
R21020 a_n3827_n3924.n34 a_n3827_n3924.n1 53.0054
R21021 a_n3827_n3924.n2 a_n3827_n3924.n14 53.0052
R21022 a_n3827_n3924.n2 a_n3827_n3924.n15 53.0052
R21023 a_n3827_n3924.n2 a_n3827_n3924.n16 53.0052
R21024 a_n3827_n3924.n3 a_n3827_n3924.n17 53.0052
R21025 a_n3827_n3924.n3 a_n3827_n3924.n18 53.0052
R21026 a_n3827_n3924.n3 a_n3827_n3924.n19 53.0052
R21027 a_n3827_n3924.n3 a_n3827_n3924.n20 53.0052
R21028 a_n3827_n3924.n9 a_n3827_n3924.n21 53.0052
R21029 a_n3827_n3924.n9 a_n3827_n3924.n22 53.0052
R21030 a_n3827_n3924.n10 a_n3827_n3924.n23 53.0052
R21031 a_n3827_n3924.n1 a_n3827_n3924.n32 53.0051
R21032 a_n3827_n3924.n1 a_n3827_n3924.n33 53.0051
R21033 a_n3827_n3924.n0 a_n3827_n3924.n13 53.0051
R21034 a_n3827_n3924.n0 a_n3827_n3924.n24 53.0051
R21035 a_n3827_n3924.n0 a_n3827_n3924.n25 53.0051
R21036 a_n3827_n3924.n0 a_n3827_n3924.n26 53.0051
R21037 a_n3827_n3924.n11 a_n3827_n3924.n27 53.0051
R21038 a_n3827_n3924.n11 a_n3827_n3924.n28 53.0051
R21039 a_n3827_n3924.n12 a_n3827_n3924.n29 53.0051
R21040 a_n3827_n3924.n30 a_n3827_n3924.n10 12.2417
R21041 a_n3827_n3924.n31 a_n3827_n3924.n2 12.2417
R21042 a_n3827_n3924.n30 a_n3827_n3924.n12 5.16214
R21043 a_n3827_n3924.n1 a_n3827_n3924.n31 5.16214
R21044 a_n3827_n3924.n3 a_n3827_n3924.n2 3.18153
R21045 a_n3827_n3924.n1 a_n3827_n3924.n0 3.18153
R21046 a_n3827_n3924.n32 a_n3827_n3924.t17 2.82907
R21047 a_n3827_n3924.n32 a_n3827_n3924.t26 2.82907
R21048 a_n3827_n3924.n33 a_n3827_n3924.t21 2.82907
R21049 a_n3827_n3924.n33 a_n3827_n3924.t2 2.82907
R21050 a_n3827_n3924.n13 a_n3827_n3924.t8 2.82907
R21051 a_n3827_n3924.n13 a_n3827_n3924.t6 2.82907
R21052 a_n3827_n3924.n24 a_n3827_n3924.t4 2.82907
R21053 a_n3827_n3924.n24 a_n3827_n3924.t7 2.82907
R21054 a_n3827_n3924.n25 a_n3827_n3924.t32 2.82907
R21055 a_n3827_n3924.n25 a_n3827_n3924.t52 2.82907
R21056 a_n3827_n3924.n26 a_n3827_n3924.t33 2.82907
R21057 a_n3827_n3924.n26 a_n3827_n3924.t40 2.82907
R21058 a_n3827_n3924.n27 a_n3827_n3924.t54 2.82907
R21059 a_n3827_n3924.n27 a_n3827_n3924.t36 2.82907
R21060 a_n3827_n3924.n28 a_n3827_n3924.t45 2.82907
R21061 a_n3827_n3924.n28 a_n3827_n3924.t53 2.82907
R21062 a_n3827_n3924.n29 a_n3827_n3924.t44 2.82907
R21063 a_n3827_n3924.n29 a_n3827_n3924.t41 2.82907
R21064 a_n3827_n3924.n14 a_n3827_n3924.t31 2.82907
R21065 a_n3827_n3924.n14 a_n3827_n3924.t39 2.82907
R21066 a_n3827_n3924.n15 a_n3827_n3924.t50 2.82907
R21067 a_n3827_n3924.n15 a_n3827_n3924.t51 2.82907
R21068 a_n3827_n3924.n16 a_n3827_n3924.t34 2.82907
R21069 a_n3827_n3924.n16 a_n3827_n3924.t48 2.82907
R21070 a_n3827_n3924.n17 a_n3827_n3924.t38 2.82907
R21071 a_n3827_n3924.n17 a_n3827_n3924.t49 2.82907
R21072 a_n3827_n3924.n18 a_n3827_n3924.t42 2.82907
R21073 a_n3827_n3924.n18 a_n3827_n3924.t37 2.82907
R21074 a_n3827_n3924.n19 a_n3827_n3924.t19 2.82907
R21075 a_n3827_n3924.n19 a_n3827_n3924.t12 2.82907
R21076 a_n3827_n3924.n20 a_n3827_n3924.t29 2.82907
R21077 a_n3827_n3924.n20 a_n3827_n3924.t22 2.82907
R21078 a_n3827_n3924.n21 a_n3827_n3924.t57 2.82907
R21079 a_n3827_n3924.n21 a_n3827_n3924.t30 2.82907
R21080 a_n3827_n3924.n22 a_n3827_n3924.t20 2.82907
R21081 a_n3827_n3924.n22 a_n3827_n3924.t15 2.82907
R21082 a_n3827_n3924.n23 a_n3827_n3924.t11 2.82907
R21083 a_n3827_n3924.n23 a_n3827_n3924.t27 2.82907
R21084 a_n3827_n3924.n34 a_n3827_n3924.t14 2.82907
R21085 a_n3827_n3924.t0 a_n3827_n3924.n34 2.82907
R21086 a_n3827_n3924.n4 a_n3827_n3924.n30 1.95694
R21087 a_n3827_n3924.n31 a_n3827_n3924.n8 1.95694
R21088 a_n3827_n3924.n9 a_n3827_n3924.n3 1.82593
R21089 a_n3827_n3924.n11 a_n3827_n3924.n0 1.82593
R21090 a_n3827_n3924.n12 a_n3827_n3924.n11 1.59102
R21091 a_n3827_n3924.n10 a_n3827_n3924.n9 1.59102
R21092 a_n3827_n3924.n5 a_n3827_n3924.n4 1.39948
R21093 a_n3827_n3924.n7 a_n3827_n3924.n6 1.34352
R21094 a_n3827_n3924.n6 a_n3827_n3924.n5 1.34352
R21095 a_n3827_n3924.n8 a_n3827_n3924.n7 1.25704
R21096 a_n7636_8799.n233 a_n7636_8799.t65 485.149
R21097 a_n7636_8799.n295 a_n7636_8799.t77 485.149
R21098 a_n7636_8799.n358 a_n7636_8799.t114 485.149
R21099 a_n7636_8799.n43 a_n7636_8799.t137 485.149
R21100 a_n7636_8799.n105 a_n7636_8799.t151 485.149
R21101 a_n7636_8799.n168 a_n7636_8799.t113 485.149
R21102 a_n7636_8799.n276 a_n7636_8799.t87 464.166
R21103 a_n7636_8799.n275 a_n7636_8799.t86 464.166
R21104 a_n7636_8799.n217 a_n7636_8799.t59 464.166
R21105 a_n7636_8799.n269 a_n7636_8799.t135 464.166
R21106 a_n7636_8799.n268 a_n7636_8799.t90 464.166
R21107 a_n7636_8799.n220 a_n7636_8799.t66 464.166
R21108 a_n7636_8799.n262 a_n7636_8799.t141 464.166
R21109 a_n7636_8799.n261 a_n7636_8799.t107 464.166
R21110 a_n7636_8799.n223 a_n7636_8799.t105 464.166
R21111 a_n7636_8799.n255 a_n7636_8799.t40 464.166
R21112 a_n7636_8799.n254 a_n7636_8799.t111 464.166
R21113 a_n7636_8799.n226 a_n7636_8799.t110 464.166
R21114 a_n7636_8799.n248 a_n7636_8799.t42 464.166
R21115 a_n7636_8799.n247 a_n7636_8799.t41 464.166
R21116 a_n7636_8799.n229 a_n7636_8799.t127 464.166
R21117 a_n7636_8799.n241 a_n7636_8799.t61 464.166
R21118 a_n7636_8799.n240 a_n7636_8799.t44 464.166
R21119 a_n7636_8799.n232 a_n7636_8799.t131 464.166
R21120 a_n7636_8799.n234 a_n7636_8799.t89 464.166
R21121 a_n7636_8799.n338 a_n7636_8799.t97 464.166
R21122 a_n7636_8799.n337 a_n7636_8799.t96 464.166
R21123 a_n7636_8799.n279 a_n7636_8799.t74 464.166
R21124 a_n7636_8799.n331 a_n7636_8799.t150 464.166
R21125 a_n7636_8799.n330 a_n7636_8799.t104 464.166
R21126 a_n7636_8799.n282 a_n7636_8799.t76 464.166
R21127 a_n7636_8799.n324 a_n7636_8799.t36 464.166
R21128 a_n7636_8799.n323 a_n7636_8799.t120 464.166
R21129 a_n7636_8799.n285 a_n7636_8799.t119 464.166
R21130 a_n7636_8799.n317 a_n7636_8799.t50 464.166
R21131 a_n7636_8799.n316 a_n7636_8799.t123 464.166
R21132 a_n7636_8799.n288 a_n7636_8799.t122 464.166
R21133 a_n7636_8799.n310 a_n7636_8799.t54 464.166
R21134 a_n7636_8799.n309 a_n7636_8799.t53 464.166
R21135 a_n7636_8799.n291 a_n7636_8799.t144 464.166
R21136 a_n7636_8799.n303 a_n7636_8799.t75 464.166
R21137 a_n7636_8799.n302 a_n7636_8799.t57 464.166
R21138 a_n7636_8799.n294 a_n7636_8799.t145 464.166
R21139 a_n7636_8799.n296 a_n7636_8799.t103 464.166
R21140 a_n7636_8799.n401 a_n7636_8799.t154 464.166
R21141 a_n7636_8799.n400 a_n7636_8799.t52 464.166
R21142 a_n7636_8799.n342 a_n7636_8799.t102 464.166
R21143 a_n7636_8799.n394 a_n7636_8799.t39 464.166
R21144 a_n7636_8799.n393 a_n7636_8799.t126 464.166
R21145 a_n7636_8799.n345 a_n7636_8799.t63 464.166
R21146 a_n7636_8799.n387 a_n7636_8799.t109 464.166
R21147 a_n7636_8799.n386 a_n7636_8799.t45 464.166
R21148 a_n7636_8799.n348 a_n7636_8799.t69 464.166
R21149 a_n7636_8799.n380 a_n7636_8799.t149 464.166
R21150 a_n7636_8799.n379 a_n7636_8799.t118 464.166
R21151 a_n7636_8799.n351 a_n7636_8799.t143 464.166
R21152 a_n7636_8799.n373 a_n7636_8799.t100 464.166
R21153 a_n7636_8799.n372 a_n7636_8799.t121 464.166
R21154 a_n7636_8799.n354 a_n7636_8799.t56 464.166
R21155 a_n7636_8799.n366 a_n7636_8799.t140 464.166
R21156 a_n7636_8799.n365 a_n7636_8799.t81 464.166
R21157 a_n7636_8799.n357 a_n7636_8799.t132 464.166
R21158 a_n7636_8799.n359 a_n7636_8799.t68 464.166
R21159 a_n7636_8799.n44 a_n7636_8799.t138 464.166
R21160 a_n7636_8799.n46 a_n7636_8799.t88 464.166
R21161 a_n7636_8799.n50 a_n7636_8799.t117 464.166
R21162 a_n7636_8799.n51 a_n7636_8799.t134 464.166
R21163 a_n7636_8799.n39 a_n7636_8799.t84 464.166
R21164 a_n7636_8799.n57 a_n7636_8799.t85 464.166
R21165 a_n7636_8799.n58 a_n7636_8799.t115 464.166
R21166 a_n7636_8799.n62 a_n7636_8799.t72 464.166
R21167 a_n7636_8799.n64 a_n7636_8799.t73 464.166
R21168 a_n7636_8799.n35 a_n7636_8799.t112 464.166
R21169 a_n7636_8799.n69 a_n7636_8799.t37 464.166
R21170 a_n7636_8799.n33 a_n7636_8799.t70 464.166
R21171 a_n7636_8799.n74 a_n7636_8799.t93 464.166
R21172 a_n7636_8799.n76 a_n7636_8799.t136 464.166
R21173 a_n7636_8799.n80 a_n7636_8799.t49 464.166
R21174 a_n7636_8799.n81 a_n7636_8799.t67 464.166
R21175 a_n7636_8799.n29 a_n7636_8799.t133 464.166
R21176 a_n7636_8799.n87 a_n7636_8799.t46 464.166
R21177 a_n7636_8799.n88 a_n7636_8799.t47 464.166
R21178 a_n7636_8799.n106 a_n7636_8799.t155 464.166
R21179 a_n7636_8799.n108 a_n7636_8799.t98 464.166
R21180 a_n7636_8799.n112 a_n7636_8799.t130 464.166
R21181 a_n7636_8799.n113 a_n7636_8799.t148 464.166
R21182 a_n7636_8799.n101 a_n7636_8799.t94 464.166
R21183 a_n7636_8799.n119 a_n7636_8799.t95 464.166
R21184 a_n7636_8799.n120 a_n7636_8799.t128 464.166
R21185 a_n7636_8799.n124 a_n7636_8799.t82 464.166
R21186 a_n7636_8799.n126 a_n7636_8799.t83 464.166
R21187 a_n7636_8799.n97 a_n7636_8799.t124 464.166
R21188 a_n7636_8799.n131 a_n7636_8799.t48 464.166
R21189 a_n7636_8799.n95 a_n7636_8799.t79 464.166
R21190 a_n7636_8799.n136 a_n7636_8799.t106 464.166
R21191 a_n7636_8799.n138 a_n7636_8799.t152 464.166
R21192 a_n7636_8799.n142 a_n7636_8799.t64 464.166
R21193 a_n7636_8799.n143 a_n7636_8799.t78 464.166
R21194 a_n7636_8799.n91 a_n7636_8799.t146 464.166
R21195 a_n7636_8799.n149 a_n7636_8799.t58 464.166
R21196 a_n7636_8799.n150 a_n7636_8799.t60 464.166
R21197 a_n7636_8799.n169 a_n7636_8799.t91 464.166
R21198 a_n7636_8799.n171 a_n7636_8799.t129 464.166
R21199 a_n7636_8799.n175 a_n7636_8799.t80 464.166
R21200 a_n7636_8799.n176 a_n7636_8799.t139 464.166
R21201 a_n7636_8799.n164 a_n7636_8799.t55 464.166
R21202 a_n7636_8799.n182 a_n7636_8799.t38 464.166
R21203 a_n7636_8799.n183 a_n7636_8799.t99 464.166
R21204 a_n7636_8799.n187 a_n7636_8799.t142 464.166
R21205 a_n7636_8799.n189 a_n7636_8799.t116 464.166
R21206 a_n7636_8799.n160 a_n7636_8799.t147 464.166
R21207 a_n7636_8799.n194 a_n7636_8799.t92 464.166
R21208 a_n7636_8799.n158 a_n7636_8799.t43 464.166
R21209 a_n7636_8799.n199 a_n7636_8799.t108 464.166
R21210 a_n7636_8799.n201 a_n7636_8799.t62 464.166
R21211 a_n7636_8799.n205 a_n7636_8799.t125 464.166
R21212 a_n7636_8799.n206 a_n7636_8799.t71 464.166
R21213 a_n7636_8799.n154 a_n7636_8799.t101 464.166
R21214 a_n7636_8799.n212 a_n7636_8799.t51 464.166
R21215 a_n7636_8799.n213 a_n7636_8799.t153 464.166
R21216 a_n7636_8799.n236 a_n7636_8799.n235 161.3
R21217 a_n7636_8799.n237 a_n7636_8799.n232 161.3
R21218 a_n7636_8799.n239 a_n7636_8799.n238 161.3
R21219 a_n7636_8799.n240 a_n7636_8799.n231 161.3
R21220 a_n7636_8799.n241 a_n7636_8799.n230 161.3
R21221 a_n7636_8799.n243 a_n7636_8799.n242 161.3
R21222 a_n7636_8799.n244 a_n7636_8799.n229 161.3
R21223 a_n7636_8799.n246 a_n7636_8799.n245 161.3
R21224 a_n7636_8799.n247 a_n7636_8799.n228 161.3
R21225 a_n7636_8799.n248 a_n7636_8799.n227 161.3
R21226 a_n7636_8799.n250 a_n7636_8799.n249 161.3
R21227 a_n7636_8799.n251 a_n7636_8799.n226 161.3
R21228 a_n7636_8799.n253 a_n7636_8799.n252 161.3
R21229 a_n7636_8799.n254 a_n7636_8799.n225 161.3
R21230 a_n7636_8799.n255 a_n7636_8799.n224 161.3
R21231 a_n7636_8799.n257 a_n7636_8799.n256 161.3
R21232 a_n7636_8799.n258 a_n7636_8799.n223 161.3
R21233 a_n7636_8799.n260 a_n7636_8799.n259 161.3
R21234 a_n7636_8799.n261 a_n7636_8799.n222 161.3
R21235 a_n7636_8799.n262 a_n7636_8799.n221 161.3
R21236 a_n7636_8799.n264 a_n7636_8799.n263 161.3
R21237 a_n7636_8799.n265 a_n7636_8799.n220 161.3
R21238 a_n7636_8799.n267 a_n7636_8799.n266 161.3
R21239 a_n7636_8799.n268 a_n7636_8799.n219 161.3
R21240 a_n7636_8799.n269 a_n7636_8799.n218 161.3
R21241 a_n7636_8799.n271 a_n7636_8799.n270 161.3
R21242 a_n7636_8799.n272 a_n7636_8799.n217 161.3
R21243 a_n7636_8799.n274 a_n7636_8799.n273 161.3
R21244 a_n7636_8799.n275 a_n7636_8799.n216 161.3
R21245 a_n7636_8799.n277 a_n7636_8799.n276 161.3
R21246 a_n7636_8799.n298 a_n7636_8799.n297 161.3
R21247 a_n7636_8799.n299 a_n7636_8799.n294 161.3
R21248 a_n7636_8799.n301 a_n7636_8799.n300 161.3
R21249 a_n7636_8799.n302 a_n7636_8799.n293 161.3
R21250 a_n7636_8799.n303 a_n7636_8799.n292 161.3
R21251 a_n7636_8799.n305 a_n7636_8799.n304 161.3
R21252 a_n7636_8799.n306 a_n7636_8799.n291 161.3
R21253 a_n7636_8799.n308 a_n7636_8799.n307 161.3
R21254 a_n7636_8799.n309 a_n7636_8799.n290 161.3
R21255 a_n7636_8799.n310 a_n7636_8799.n289 161.3
R21256 a_n7636_8799.n312 a_n7636_8799.n311 161.3
R21257 a_n7636_8799.n313 a_n7636_8799.n288 161.3
R21258 a_n7636_8799.n315 a_n7636_8799.n314 161.3
R21259 a_n7636_8799.n316 a_n7636_8799.n287 161.3
R21260 a_n7636_8799.n317 a_n7636_8799.n286 161.3
R21261 a_n7636_8799.n319 a_n7636_8799.n318 161.3
R21262 a_n7636_8799.n320 a_n7636_8799.n285 161.3
R21263 a_n7636_8799.n322 a_n7636_8799.n321 161.3
R21264 a_n7636_8799.n323 a_n7636_8799.n284 161.3
R21265 a_n7636_8799.n324 a_n7636_8799.n283 161.3
R21266 a_n7636_8799.n326 a_n7636_8799.n325 161.3
R21267 a_n7636_8799.n327 a_n7636_8799.n282 161.3
R21268 a_n7636_8799.n329 a_n7636_8799.n328 161.3
R21269 a_n7636_8799.n330 a_n7636_8799.n281 161.3
R21270 a_n7636_8799.n331 a_n7636_8799.n280 161.3
R21271 a_n7636_8799.n333 a_n7636_8799.n332 161.3
R21272 a_n7636_8799.n334 a_n7636_8799.n279 161.3
R21273 a_n7636_8799.n336 a_n7636_8799.n335 161.3
R21274 a_n7636_8799.n337 a_n7636_8799.n278 161.3
R21275 a_n7636_8799.n339 a_n7636_8799.n338 161.3
R21276 a_n7636_8799.n361 a_n7636_8799.n360 161.3
R21277 a_n7636_8799.n362 a_n7636_8799.n357 161.3
R21278 a_n7636_8799.n364 a_n7636_8799.n363 161.3
R21279 a_n7636_8799.n365 a_n7636_8799.n356 161.3
R21280 a_n7636_8799.n366 a_n7636_8799.n355 161.3
R21281 a_n7636_8799.n368 a_n7636_8799.n367 161.3
R21282 a_n7636_8799.n369 a_n7636_8799.n354 161.3
R21283 a_n7636_8799.n371 a_n7636_8799.n370 161.3
R21284 a_n7636_8799.n372 a_n7636_8799.n353 161.3
R21285 a_n7636_8799.n373 a_n7636_8799.n352 161.3
R21286 a_n7636_8799.n375 a_n7636_8799.n374 161.3
R21287 a_n7636_8799.n376 a_n7636_8799.n351 161.3
R21288 a_n7636_8799.n378 a_n7636_8799.n377 161.3
R21289 a_n7636_8799.n379 a_n7636_8799.n350 161.3
R21290 a_n7636_8799.n380 a_n7636_8799.n349 161.3
R21291 a_n7636_8799.n382 a_n7636_8799.n381 161.3
R21292 a_n7636_8799.n383 a_n7636_8799.n348 161.3
R21293 a_n7636_8799.n385 a_n7636_8799.n384 161.3
R21294 a_n7636_8799.n386 a_n7636_8799.n347 161.3
R21295 a_n7636_8799.n387 a_n7636_8799.n346 161.3
R21296 a_n7636_8799.n389 a_n7636_8799.n388 161.3
R21297 a_n7636_8799.n390 a_n7636_8799.n345 161.3
R21298 a_n7636_8799.n392 a_n7636_8799.n391 161.3
R21299 a_n7636_8799.n393 a_n7636_8799.n344 161.3
R21300 a_n7636_8799.n394 a_n7636_8799.n343 161.3
R21301 a_n7636_8799.n396 a_n7636_8799.n395 161.3
R21302 a_n7636_8799.n397 a_n7636_8799.n342 161.3
R21303 a_n7636_8799.n399 a_n7636_8799.n398 161.3
R21304 a_n7636_8799.n400 a_n7636_8799.n341 161.3
R21305 a_n7636_8799.n402 a_n7636_8799.n401 161.3
R21306 a_n7636_8799.n89 a_n7636_8799.n88 161.3
R21307 a_n7636_8799.n87 a_n7636_8799.n28 161.3
R21308 a_n7636_8799.n86 a_n7636_8799.n85 161.3
R21309 a_n7636_8799.n84 a_n7636_8799.n29 161.3
R21310 a_n7636_8799.n83 a_n7636_8799.n82 161.3
R21311 a_n7636_8799.n81 a_n7636_8799.n30 161.3
R21312 a_n7636_8799.n80 a_n7636_8799.n79 161.3
R21313 a_n7636_8799.n78 a_n7636_8799.n31 161.3
R21314 a_n7636_8799.n77 a_n7636_8799.n76 161.3
R21315 a_n7636_8799.n75 a_n7636_8799.n32 161.3
R21316 a_n7636_8799.n74 a_n7636_8799.n73 161.3
R21317 a_n7636_8799.n72 a_n7636_8799.n33 161.3
R21318 a_n7636_8799.n71 a_n7636_8799.n70 161.3
R21319 a_n7636_8799.n69 a_n7636_8799.n34 161.3
R21320 a_n7636_8799.n68 a_n7636_8799.n67 161.3
R21321 a_n7636_8799.n66 a_n7636_8799.n35 161.3
R21322 a_n7636_8799.n65 a_n7636_8799.n64 161.3
R21323 a_n7636_8799.n63 a_n7636_8799.n36 161.3
R21324 a_n7636_8799.n62 a_n7636_8799.n61 161.3
R21325 a_n7636_8799.n60 a_n7636_8799.n37 161.3
R21326 a_n7636_8799.n59 a_n7636_8799.n58 161.3
R21327 a_n7636_8799.n57 a_n7636_8799.n38 161.3
R21328 a_n7636_8799.n56 a_n7636_8799.n55 161.3
R21329 a_n7636_8799.n54 a_n7636_8799.n39 161.3
R21330 a_n7636_8799.n53 a_n7636_8799.n52 161.3
R21331 a_n7636_8799.n51 a_n7636_8799.n40 161.3
R21332 a_n7636_8799.n50 a_n7636_8799.n49 161.3
R21333 a_n7636_8799.n48 a_n7636_8799.n41 161.3
R21334 a_n7636_8799.n47 a_n7636_8799.n46 161.3
R21335 a_n7636_8799.n45 a_n7636_8799.n42 161.3
R21336 a_n7636_8799.n151 a_n7636_8799.n150 161.3
R21337 a_n7636_8799.n149 a_n7636_8799.n90 161.3
R21338 a_n7636_8799.n148 a_n7636_8799.n147 161.3
R21339 a_n7636_8799.n146 a_n7636_8799.n91 161.3
R21340 a_n7636_8799.n145 a_n7636_8799.n144 161.3
R21341 a_n7636_8799.n143 a_n7636_8799.n92 161.3
R21342 a_n7636_8799.n142 a_n7636_8799.n141 161.3
R21343 a_n7636_8799.n140 a_n7636_8799.n93 161.3
R21344 a_n7636_8799.n139 a_n7636_8799.n138 161.3
R21345 a_n7636_8799.n137 a_n7636_8799.n94 161.3
R21346 a_n7636_8799.n136 a_n7636_8799.n135 161.3
R21347 a_n7636_8799.n134 a_n7636_8799.n95 161.3
R21348 a_n7636_8799.n133 a_n7636_8799.n132 161.3
R21349 a_n7636_8799.n131 a_n7636_8799.n96 161.3
R21350 a_n7636_8799.n130 a_n7636_8799.n129 161.3
R21351 a_n7636_8799.n128 a_n7636_8799.n97 161.3
R21352 a_n7636_8799.n127 a_n7636_8799.n126 161.3
R21353 a_n7636_8799.n125 a_n7636_8799.n98 161.3
R21354 a_n7636_8799.n124 a_n7636_8799.n123 161.3
R21355 a_n7636_8799.n122 a_n7636_8799.n99 161.3
R21356 a_n7636_8799.n121 a_n7636_8799.n120 161.3
R21357 a_n7636_8799.n119 a_n7636_8799.n100 161.3
R21358 a_n7636_8799.n118 a_n7636_8799.n117 161.3
R21359 a_n7636_8799.n116 a_n7636_8799.n101 161.3
R21360 a_n7636_8799.n115 a_n7636_8799.n114 161.3
R21361 a_n7636_8799.n113 a_n7636_8799.n102 161.3
R21362 a_n7636_8799.n112 a_n7636_8799.n111 161.3
R21363 a_n7636_8799.n110 a_n7636_8799.n103 161.3
R21364 a_n7636_8799.n109 a_n7636_8799.n108 161.3
R21365 a_n7636_8799.n107 a_n7636_8799.n104 161.3
R21366 a_n7636_8799.n214 a_n7636_8799.n213 161.3
R21367 a_n7636_8799.n212 a_n7636_8799.n153 161.3
R21368 a_n7636_8799.n211 a_n7636_8799.n210 161.3
R21369 a_n7636_8799.n209 a_n7636_8799.n154 161.3
R21370 a_n7636_8799.n208 a_n7636_8799.n207 161.3
R21371 a_n7636_8799.n206 a_n7636_8799.n155 161.3
R21372 a_n7636_8799.n205 a_n7636_8799.n204 161.3
R21373 a_n7636_8799.n203 a_n7636_8799.n156 161.3
R21374 a_n7636_8799.n202 a_n7636_8799.n201 161.3
R21375 a_n7636_8799.n200 a_n7636_8799.n157 161.3
R21376 a_n7636_8799.n199 a_n7636_8799.n198 161.3
R21377 a_n7636_8799.n197 a_n7636_8799.n158 161.3
R21378 a_n7636_8799.n196 a_n7636_8799.n195 161.3
R21379 a_n7636_8799.n194 a_n7636_8799.n159 161.3
R21380 a_n7636_8799.n193 a_n7636_8799.n192 161.3
R21381 a_n7636_8799.n191 a_n7636_8799.n160 161.3
R21382 a_n7636_8799.n190 a_n7636_8799.n189 161.3
R21383 a_n7636_8799.n188 a_n7636_8799.n161 161.3
R21384 a_n7636_8799.n187 a_n7636_8799.n186 161.3
R21385 a_n7636_8799.n185 a_n7636_8799.n162 161.3
R21386 a_n7636_8799.n184 a_n7636_8799.n183 161.3
R21387 a_n7636_8799.n182 a_n7636_8799.n163 161.3
R21388 a_n7636_8799.n181 a_n7636_8799.n180 161.3
R21389 a_n7636_8799.n179 a_n7636_8799.n164 161.3
R21390 a_n7636_8799.n178 a_n7636_8799.n177 161.3
R21391 a_n7636_8799.n176 a_n7636_8799.n165 161.3
R21392 a_n7636_8799.n175 a_n7636_8799.n174 161.3
R21393 a_n7636_8799.n173 a_n7636_8799.n166 161.3
R21394 a_n7636_8799.n172 a_n7636_8799.n171 161.3
R21395 a_n7636_8799.n170 a_n7636_8799.n167 161.3
R21396 a_n7636_8799.n2 a_n7636_8799.n0 98.9633
R21397 a_n7636_8799.n410 a_n7636_8799.n409 98.9631
R21398 a_n7636_8799.n408 a_n7636_8799.n407 98.6055
R21399 a_n7636_8799.n4 a_n7636_8799.n3 98.6055
R21400 a_n7636_8799.n2 a_n7636_8799.n1 98.6055
R21401 a_n7636_8799.n411 a_n7636_8799.n410 98.6054
R21402 a_n7636_8799.n7 a_n7636_8799.n5 81.4626
R21403 a_n7636_8799.n17 a_n7636_8799.n15 81.4626
R21404 a_n7636_8799.n12 a_n7636_8799.n10 81.4626
R21405 a_n7636_8799.n22 a_n7636_8799.n21 80.9324
R21406 a_n7636_8799.n24 a_n7636_8799.n23 80.9324
R21407 a_n7636_8799.n26 a_n7636_8799.n25 80.9324
R21408 a_n7636_8799.n9 a_n7636_8799.n8 80.9324
R21409 a_n7636_8799.n7 a_n7636_8799.n6 80.9324
R21410 a_n7636_8799.n17 a_n7636_8799.n16 80.9324
R21411 a_n7636_8799.n19 a_n7636_8799.n18 80.9324
R21412 a_n7636_8799.n14 a_n7636_8799.n13 80.9324
R21413 a_n7636_8799.n12 a_n7636_8799.n11 80.9324
R21414 a_n7636_8799.n236 a_n7636_8799.n233 70.4033
R21415 a_n7636_8799.n298 a_n7636_8799.n295 70.4033
R21416 a_n7636_8799.n361 a_n7636_8799.n358 70.4033
R21417 a_n7636_8799.n43 a_n7636_8799.n42 70.4033
R21418 a_n7636_8799.n105 a_n7636_8799.n104 70.4033
R21419 a_n7636_8799.n168 a_n7636_8799.n167 70.4033
R21420 a_n7636_8799.n276 a_n7636_8799.n275 48.2005
R21421 a_n7636_8799.n269 a_n7636_8799.n268 48.2005
R21422 a_n7636_8799.n262 a_n7636_8799.n261 48.2005
R21423 a_n7636_8799.n255 a_n7636_8799.n254 48.2005
R21424 a_n7636_8799.n248 a_n7636_8799.n247 48.2005
R21425 a_n7636_8799.n241 a_n7636_8799.n240 48.2005
R21426 a_n7636_8799.n338 a_n7636_8799.n337 48.2005
R21427 a_n7636_8799.n331 a_n7636_8799.n330 48.2005
R21428 a_n7636_8799.n324 a_n7636_8799.n323 48.2005
R21429 a_n7636_8799.n317 a_n7636_8799.n316 48.2005
R21430 a_n7636_8799.n310 a_n7636_8799.n309 48.2005
R21431 a_n7636_8799.n303 a_n7636_8799.n302 48.2005
R21432 a_n7636_8799.n401 a_n7636_8799.n400 48.2005
R21433 a_n7636_8799.n394 a_n7636_8799.n393 48.2005
R21434 a_n7636_8799.n387 a_n7636_8799.n386 48.2005
R21435 a_n7636_8799.n380 a_n7636_8799.n379 48.2005
R21436 a_n7636_8799.n373 a_n7636_8799.n372 48.2005
R21437 a_n7636_8799.n366 a_n7636_8799.n365 48.2005
R21438 a_n7636_8799.n51 a_n7636_8799.n50 48.2005
R21439 a_n7636_8799.n58 a_n7636_8799.n57 48.2005
R21440 a_n7636_8799.n64 a_n7636_8799.n35 48.2005
R21441 a_n7636_8799.n74 a_n7636_8799.n33 48.2005
R21442 a_n7636_8799.n81 a_n7636_8799.n80 48.2005
R21443 a_n7636_8799.n88 a_n7636_8799.n87 48.2005
R21444 a_n7636_8799.n113 a_n7636_8799.n112 48.2005
R21445 a_n7636_8799.n120 a_n7636_8799.n119 48.2005
R21446 a_n7636_8799.n126 a_n7636_8799.n97 48.2005
R21447 a_n7636_8799.n136 a_n7636_8799.n95 48.2005
R21448 a_n7636_8799.n143 a_n7636_8799.n142 48.2005
R21449 a_n7636_8799.n150 a_n7636_8799.n149 48.2005
R21450 a_n7636_8799.n176 a_n7636_8799.n175 48.2005
R21451 a_n7636_8799.n183 a_n7636_8799.n182 48.2005
R21452 a_n7636_8799.n189 a_n7636_8799.n160 48.2005
R21453 a_n7636_8799.n199 a_n7636_8799.n158 48.2005
R21454 a_n7636_8799.n206 a_n7636_8799.n205 48.2005
R21455 a_n7636_8799.n213 a_n7636_8799.n212 48.2005
R21456 a_n7636_8799.n274 a_n7636_8799.n217 40.1672
R21457 a_n7636_8799.n235 a_n7636_8799.n232 40.1672
R21458 a_n7636_8799.n336 a_n7636_8799.n279 40.1672
R21459 a_n7636_8799.n297 a_n7636_8799.n294 40.1672
R21460 a_n7636_8799.n399 a_n7636_8799.n342 40.1672
R21461 a_n7636_8799.n360 a_n7636_8799.n357 40.1672
R21462 a_n7636_8799.n46 a_n7636_8799.n45 40.1672
R21463 a_n7636_8799.n86 a_n7636_8799.n29 40.1672
R21464 a_n7636_8799.n108 a_n7636_8799.n107 40.1672
R21465 a_n7636_8799.n148 a_n7636_8799.n91 40.1672
R21466 a_n7636_8799.n171 a_n7636_8799.n170 40.1672
R21467 a_n7636_8799.n211 a_n7636_8799.n154 40.1672
R21468 a_n7636_8799.n267 a_n7636_8799.n220 38.7066
R21469 a_n7636_8799.n242 a_n7636_8799.n229 38.7066
R21470 a_n7636_8799.n329 a_n7636_8799.n282 38.7066
R21471 a_n7636_8799.n304 a_n7636_8799.n291 38.7066
R21472 a_n7636_8799.n392 a_n7636_8799.n345 38.7066
R21473 a_n7636_8799.n367 a_n7636_8799.n354 38.7066
R21474 a_n7636_8799.n52 a_n7636_8799.n39 38.7066
R21475 a_n7636_8799.n76 a_n7636_8799.n31 38.7066
R21476 a_n7636_8799.n114 a_n7636_8799.n101 38.7066
R21477 a_n7636_8799.n138 a_n7636_8799.n93 38.7066
R21478 a_n7636_8799.n177 a_n7636_8799.n164 38.7066
R21479 a_n7636_8799.n201 a_n7636_8799.n156 38.7066
R21480 a_n7636_8799.n260 a_n7636_8799.n223 37.246
R21481 a_n7636_8799.n249 a_n7636_8799.n226 37.246
R21482 a_n7636_8799.n322 a_n7636_8799.n285 37.246
R21483 a_n7636_8799.n311 a_n7636_8799.n288 37.246
R21484 a_n7636_8799.n385 a_n7636_8799.n348 37.246
R21485 a_n7636_8799.n374 a_n7636_8799.n351 37.246
R21486 a_n7636_8799.n62 a_n7636_8799.n37 37.246
R21487 a_n7636_8799.n70 a_n7636_8799.n69 37.246
R21488 a_n7636_8799.n124 a_n7636_8799.n99 37.246
R21489 a_n7636_8799.n132 a_n7636_8799.n131 37.246
R21490 a_n7636_8799.n187 a_n7636_8799.n162 37.246
R21491 a_n7636_8799.n195 a_n7636_8799.n194 37.246
R21492 a_n7636_8799.n256 a_n7636_8799.n223 35.7853
R21493 a_n7636_8799.n253 a_n7636_8799.n226 35.7853
R21494 a_n7636_8799.n318 a_n7636_8799.n285 35.7853
R21495 a_n7636_8799.n315 a_n7636_8799.n288 35.7853
R21496 a_n7636_8799.n381 a_n7636_8799.n348 35.7853
R21497 a_n7636_8799.n378 a_n7636_8799.n351 35.7853
R21498 a_n7636_8799.n63 a_n7636_8799.n62 35.7853
R21499 a_n7636_8799.n69 a_n7636_8799.n68 35.7853
R21500 a_n7636_8799.n125 a_n7636_8799.n124 35.7853
R21501 a_n7636_8799.n131 a_n7636_8799.n130 35.7853
R21502 a_n7636_8799.n188 a_n7636_8799.n187 35.7853
R21503 a_n7636_8799.n194 a_n7636_8799.n193 35.7853
R21504 a_n7636_8799.n263 a_n7636_8799.n220 34.3247
R21505 a_n7636_8799.n246 a_n7636_8799.n229 34.3247
R21506 a_n7636_8799.n325 a_n7636_8799.n282 34.3247
R21507 a_n7636_8799.n308 a_n7636_8799.n291 34.3247
R21508 a_n7636_8799.n388 a_n7636_8799.n345 34.3247
R21509 a_n7636_8799.n371 a_n7636_8799.n354 34.3247
R21510 a_n7636_8799.n56 a_n7636_8799.n39 34.3247
R21511 a_n7636_8799.n76 a_n7636_8799.n75 34.3247
R21512 a_n7636_8799.n118 a_n7636_8799.n101 34.3247
R21513 a_n7636_8799.n138 a_n7636_8799.n137 34.3247
R21514 a_n7636_8799.n181 a_n7636_8799.n164 34.3247
R21515 a_n7636_8799.n201 a_n7636_8799.n200 34.3247
R21516 a_n7636_8799.n22 a_n7636_8799.n20 34.3237
R21517 a_n7636_8799.n270 a_n7636_8799.n217 32.8641
R21518 a_n7636_8799.n239 a_n7636_8799.n232 32.8641
R21519 a_n7636_8799.n332 a_n7636_8799.n279 32.8641
R21520 a_n7636_8799.n301 a_n7636_8799.n294 32.8641
R21521 a_n7636_8799.n395 a_n7636_8799.n342 32.8641
R21522 a_n7636_8799.n364 a_n7636_8799.n357 32.8641
R21523 a_n7636_8799.n46 a_n7636_8799.n41 32.8641
R21524 a_n7636_8799.n82 a_n7636_8799.n29 32.8641
R21525 a_n7636_8799.n108 a_n7636_8799.n103 32.8641
R21526 a_n7636_8799.n144 a_n7636_8799.n91 32.8641
R21527 a_n7636_8799.n171 a_n7636_8799.n166 32.8641
R21528 a_n7636_8799.n207 a_n7636_8799.n154 32.8641
R21529 a_n7636_8799.n408 a_n7636_8799.n406 31.1941
R21530 a_n7636_8799.n234 a_n7636_8799.n233 20.9576
R21531 a_n7636_8799.n296 a_n7636_8799.n295 20.9576
R21532 a_n7636_8799.n359 a_n7636_8799.n358 20.9576
R21533 a_n7636_8799.n44 a_n7636_8799.n43 20.9576
R21534 a_n7636_8799.n106 a_n7636_8799.n105 20.9576
R21535 a_n7636_8799.n169 a_n7636_8799.n168 20.9576
R21536 a_n7636_8799.n406 a_n7636_8799.n4 17.2555
R21537 a_n7636_8799.n270 a_n7636_8799.n269 15.3369
R21538 a_n7636_8799.n240 a_n7636_8799.n239 15.3369
R21539 a_n7636_8799.n332 a_n7636_8799.n331 15.3369
R21540 a_n7636_8799.n302 a_n7636_8799.n301 15.3369
R21541 a_n7636_8799.n395 a_n7636_8799.n394 15.3369
R21542 a_n7636_8799.n365 a_n7636_8799.n364 15.3369
R21543 a_n7636_8799.n50 a_n7636_8799.n41 15.3369
R21544 a_n7636_8799.n82 a_n7636_8799.n81 15.3369
R21545 a_n7636_8799.n112 a_n7636_8799.n103 15.3369
R21546 a_n7636_8799.n144 a_n7636_8799.n143 15.3369
R21547 a_n7636_8799.n175 a_n7636_8799.n166 15.3369
R21548 a_n7636_8799.n207 a_n7636_8799.n206 15.3369
R21549 a_n7636_8799.n263 a_n7636_8799.n262 13.8763
R21550 a_n7636_8799.n247 a_n7636_8799.n246 13.8763
R21551 a_n7636_8799.n325 a_n7636_8799.n324 13.8763
R21552 a_n7636_8799.n309 a_n7636_8799.n308 13.8763
R21553 a_n7636_8799.n388 a_n7636_8799.n387 13.8763
R21554 a_n7636_8799.n372 a_n7636_8799.n371 13.8763
R21555 a_n7636_8799.n57 a_n7636_8799.n56 13.8763
R21556 a_n7636_8799.n75 a_n7636_8799.n74 13.8763
R21557 a_n7636_8799.n119 a_n7636_8799.n118 13.8763
R21558 a_n7636_8799.n137 a_n7636_8799.n136 13.8763
R21559 a_n7636_8799.n182 a_n7636_8799.n181 13.8763
R21560 a_n7636_8799.n200 a_n7636_8799.n199 13.8763
R21561 a_n7636_8799.n256 a_n7636_8799.n255 12.4157
R21562 a_n7636_8799.n254 a_n7636_8799.n253 12.4157
R21563 a_n7636_8799.n318 a_n7636_8799.n317 12.4157
R21564 a_n7636_8799.n316 a_n7636_8799.n315 12.4157
R21565 a_n7636_8799.n381 a_n7636_8799.n380 12.4157
R21566 a_n7636_8799.n379 a_n7636_8799.n378 12.4157
R21567 a_n7636_8799.n64 a_n7636_8799.n63 12.4157
R21568 a_n7636_8799.n68 a_n7636_8799.n35 12.4157
R21569 a_n7636_8799.n126 a_n7636_8799.n125 12.4157
R21570 a_n7636_8799.n130 a_n7636_8799.n97 12.4157
R21571 a_n7636_8799.n189 a_n7636_8799.n188 12.4157
R21572 a_n7636_8799.n193 a_n7636_8799.n160 12.4157
R21573 a_n7636_8799.n405 a_n7636_8799.n27 12.3339
R21574 a_n7636_8799.n406 a_n7636_8799.n405 11.4887
R21575 a_n7636_8799.n261 a_n7636_8799.n260 10.955
R21576 a_n7636_8799.n249 a_n7636_8799.n248 10.955
R21577 a_n7636_8799.n323 a_n7636_8799.n322 10.955
R21578 a_n7636_8799.n311 a_n7636_8799.n310 10.955
R21579 a_n7636_8799.n386 a_n7636_8799.n385 10.955
R21580 a_n7636_8799.n374 a_n7636_8799.n373 10.955
R21581 a_n7636_8799.n58 a_n7636_8799.n37 10.955
R21582 a_n7636_8799.n70 a_n7636_8799.n33 10.955
R21583 a_n7636_8799.n120 a_n7636_8799.n99 10.955
R21584 a_n7636_8799.n132 a_n7636_8799.n95 10.955
R21585 a_n7636_8799.n183 a_n7636_8799.n162 10.955
R21586 a_n7636_8799.n195 a_n7636_8799.n158 10.955
R21587 a_n7636_8799.n268 a_n7636_8799.n267 9.49444
R21588 a_n7636_8799.n242 a_n7636_8799.n241 9.49444
R21589 a_n7636_8799.n330 a_n7636_8799.n329 9.49444
R21590 a_n7636_8799.n304 a_n7636_8799.n303 9.49444
R21591 a_n7636_8799.n393 a_n7636_8799.n392 9.49444
R21592 a_n7636_8799.n367 a_n7636_8799.n366 9.49444
R21593 a_n7636_8799.n52 a_n7636_8799.n51 9.49444
R21594 a_n7636_8799.n80 a_n7636_8799.n31 9.49444
R21595 a_n7636_8799.n114 a_n7636_8799.n113 9.49444
R21596 a_n7636_8799.n142 a_n7636_8799.n93 9.49444
R21597 a_n7636_8799.n177 a_n7636_8799.n176 9.49444
R21598 a_n7636_8799.n205 a_n7636_8799.n156 9.49444
R21599 a_n7636_8799.n340 a_n7636_8799.n277 9.04406
R21600 a_n7636_8799.n152 a_n7636_8799.n89 9.04406
R21601 a_n7636_8799.n275 a_n7636_8799.n274 8.03383
R21602 a_n7636_8799.n235 a_n7636_8799.n234 8.03383
R21603 a_n7636_8799.n337 a_n7636_8799.n336 8.03383
R21604 a_n7636_8799.n297 a_n7636_8799.n296 8.03383
R21605 a_n7636_8799.n400 a_n7636_8799.n399 8.03383
R21606 a_n7636_8799.n360 a_n7636_8799.n359 8.03383
R21607 a_n7636_8799.n45 a_n7636_8799.n44 8.03383
R21608 a_n7636_8799.n87 a_n7636_8799.n86 8.03383
R21609 a_n7636_8799.n107 a_n7636_8799.n106 8.03383
R21610 a_n7636_8799.n149 a_n7636_8799.n148 8.03383
R21611 a_n7636_8799.n170 a_n7636_8799.n169 8.03383
R21612 a_n7636_8799.n212 a_n7636_8799.n211 8.03383
R21613 a_n7636_8799.n404 a_n7636_8799.n215 6.93972
R21614 a_n7636_8799.n404 a_n7636_8799.n403 6.44309
R21615 a_n7636_8799.n340 a_n7636_8799.n339 4.93611
R21616 a_n7636_8799.n403 a_n7636_8799.n402 4.93611
R21617 a_n7636_8799.n152 a_n7636_8799.n151 4.93611
R21618 a_n7636_8799.n215 a_n7636_8799.n214 4.93611
R21619 a_n7636_8799.n403 a_n7636_8799.n340 4.10845
R21620 a_n7636_8799.n215 a_n7636_8799.n152 4.10845
R21621 a_n7636_8799.n409 a_n7636_8799.t5 3.61217
R21622 a_n7636_8799.n409 a_n7636_8799.t10 3.61217
R21623 a_n7636_8799.n407 a_n7636_8799.t3 3.61217
R21624 a_n7636_8799.n407 a_n7636_8799.t2 3.61217
R21625 a_n7636_8799.n3 a_n7636_8799.t4 3.61217
R21626 a_n7636_8799.n3 a_n7636_8799.t1 3.61217
R21627 a_n7636_8799.n1 a_n7636_8799.t6 3.61217
R21628 a_n7636_8799.n1 a_n7636_8799.t9 3.61217
R21629 a_n7636_8799.n0 a_n7636_8799.t0 3.61217
R21630 a_n7636_8799.n0 a_n7636_8799.t7 3.61217
R21631 a_n7636_8799.t11 a_n7636_8799.n411 3.61217
R21632 a_n7636_8799.n411 a_n7636_8799.t8 3.61217
R21633 a_n7636_8799.n405 a_n7636_8799.n404 3.4105
R21634 a_n7636_8799.n21 a_n7636_8799.t12 2.82907
R21635 a_n7636_8799.n21 a_n7636_8799.t16 2.82907
R21636 a_n7636_8799.n23 a_n7636_8799.t30 2.82907
R21637 a_n7636_8799.n23 a_n7636_8799.t14 2.82907
R21638 a_n7636_8799.n25 a_n7636_8799.t27 2.82907
R21639 a_n7636_8799.n25 a_n7636_8799.t25 2.82907
R21640 a_n7636_8799.n8 a_n7636_8799.t24 2.82907
R21641 a_n7636_8799.n8 a_n7636_8799.t23 2.82907
R21642 a_n7636_8799.n6 a_n7636_8799.t18 2.82907
R21643 a_n7636_8799.n6 a_n7636_8799.t19 2.82907
R21644 a_n7636_8799.n5 a_n7636_8799.t29 2.82907
R21645 a_n7636_8799.n5 a_n7636_8799.t35 2.82907
R21646 a_n7636_8799.n15 a_n7636_8799.t31 2.82907
R21647 a_n7636_8799.n15 a_n7636_8799.t26 2.82907
R21648 a_n7636_8799.n16 a_n7636_8799.t13 2.82907
R21649 a_n7636_8799.n16 a_n7636_8799.t15 2.82907
R21650 a_n7636_8799.n18 a_n7636_8799.t21 2.82907
R21651 a_n7636_8799.n18 a_n7636_8799.t22 2.82907
R21652 a_n7636_8799.n13 a_n7636_8799.t32 2.82907
R21653 a_n7636_8799.n13 a_n7636_8799.t33 2.82907
R21654 a_n7636_8799.n11 a_n7636_8799.t34 2.82907
R21655 a_n7636_8799.n11 a_n7636_8799.t28 2.82907
R21656 a_n7636_8799.n10 a_n7636_8799.t20 2.82907
R21657 a_n7636_8799.n10 a_n7636_8799.t17 2.82907
R21658 a_n7636_8799.n14 a_n7636_8799.n12 0.530672
R21659 a_n7636_8799.n19 a_n7636_8799.n17 0.530672
R21660 a_n7636_8799.n9 a_n7636_8799.n7 0.530672
R21661 a_n7636_8799.n26 a_n7636_8799.n24 0.530672
R21662 a_n7636_8799.n24 a_n7636_8799.n22 0.530672
R21663 a_n7636_8799.n4 a_n7636_8799.n2 0.358259
R21664 a_n7636_8799.n410 a_n7636_8799.n408 0.358259
R21665 a_n7636_8799.n20 a_n7636_8799.n14 0.265586
R21666 a_n7636_8799.n20 a_n7636_8799.n19 0.265586
R21667 a_n7636_8799.n27 a_n7636_8799.n9 0.265586
R21668 a_n7636_8799.n27 a_n7636_8799.n26 0.265586
R21669 a_n7636_8799.n277 a_n7636_8799.n216 0.189894
R21670 a_n7636_8799.n273 a_n7636_8799.n216 0.189894
R21671 a_n7636_8799.n273 a_n7636_8799.n272 0.189894
R21672 a_n7636_8799.n272 a_n7636_8799.n271 0.189894
R21673 a_n7636_8799.n271 a_n7636_8799.n218 0.189894
R21674 a_n7636_8799.n219 a_n7636_8799.n218 0.189894
R21675 a_n7636_8799.n266 a_n7636_8799.n219 0.189894
R21676 a_n7636_8799.n266 a_n7636_8799.n265 0.189894
R21677 a_n7636_8799.n265 a_n7636_8799.n264 0.189894
R21678 a_n7636_8799.n264 a_n7636_8799.n221 0.189894
R21679 a_n7636_8799.n222 a_n7636_8799.n221 0.189894
R21680 a_n7636_8799.n259 a_n7636_8799.n222 0.189894
R21681 a_n7636_8799.n259 a_n7636_8799.n258 0.189894
R21682 a_n7636_8799.n258 a_n7636_8799.n257 0.189894
R21683 a_n7636_8799.n257 a_n7636_8799.n224 0.189894
R21684 a_n7636_8799.n225 a_n7636_8799.n224 0.189894
R21685 a_n7636_8799.n252 a_n7636_8799.n225 0.189894
R21686 a_n7636_8799.n252 a_n7636_8799.n251 0.189894
R21687 a_n7636_8799.n251 a_n7636_8799.n250 0.189894
R21688 a_n7636_8799.n250 a_n7636_8799.n227 0.189894
R21689 a_n7636_8799.n228 a_n7636_8799.n227 0.189894
R21690 a_n7636_8799.n245 a_n7636_8799.n228 0.189894
R21691 a_n7636_8799.n245 a_n7636_8799.n244 0.189894
R21692 a_n7636_8799.n244 a_n7636_8799.n243 0.189894
R21693 a_n7636_8799.n243 a_n7636_8799.n230 0.189894
R21694 a_n7636_8799.n231 a_n7636_8799.n230 0.189894
R21695 a_n7636_8799.n238 a_n7636_8799.n231 0.189894
R21696 a_n7636_8799.n238 a_n7636_8799.n237 0.189894
R21697 a_n7636_8799.n237 a_n7636_8799.n236 0.189894
R21698 a_n7636_8799.n339 a_n7636_8799.n278 0.189894
R21699 a_n7636_8799.n335 a_n7636_8799.n278 0.189894
R21700 a_n7636_8799.n335 a_n7636_8799.n334 0.189894
R21701 a_n7636_8799.n334 a_n7636_8799.n333 0.189894
R21702 a_n7636_8799.n333 a_n7636_8799.n280 0.189894
R21703 a_n7636_8799.n281 a_n7636_8799.n280 0.189894
R21704 a_n7636_8799.n328 a_n7636_8799.n281 0.189894
R21705 a_n7636_8799.n328 a_n7636_8799.n327 0.189894
R21706 a_n7636_8799.n327 a_n7636_8799.n326 0.189894
R21707 a_n7636_8799.n326 a_n7636_8799.n283 0.189894
R21708 a_n7636_8799.n284 a_n7636_8799.n283 0.189894
R21709 a_n7636_8799.n321 a_n7636_8799.n284 0.189894
R21710 a_n7636_8799.n321 a_n7636_8799.n320 0.189894
R21711 a_n7636_8799.n320 a_n7636_8799.n319 0.189894
R21712 a_n7636_8799.n319 a_n7636_8799.n286 0.189894
R21713 a_n7636_8799.n287 a_n7636_8799.n286 0.189894
R21714 a_n7636_8799.n314 a_n7636_8799.n287 0.189894
R21715 a_n7636_8799.n314 a_n7636_8799.n313 0.189894
R21716 a_n7636_8799.n313 a_n7636_8799.n312 0.189894
R21717 a_n7636_8799.n312 a_n7636_8799.n289 0.189894
R21718 a_n7636_8799.n290 a_n7636_8799.n289 0.189894
R21719 a_n7636_8799.n307 a_n7636_8799.n290 0.189894
R21720 a_n7636_8799.n307 a_n7636_8799.n306 0.189894
R21721 a_n7636_8799.n306 a_n7636_8799.n305 0.189894
R21722 a_n7636_8799.n305 a_n7636_8799.n292 0.189894
R21723 a_n7636_8799.n293 a_n7636_8799.n292 0.189894
R21724 a_n7636_8799.n300 a_n7636_8799.n293 0.189894
R21725 a_n7636_8799.n300 a_n7636_8799.n299 0.189894
R21726 a_n7636_8799.n299 a_n7636_8799.n298 0.189894
R21727 a_n7636_8799.n402 a_n7636_8799.n341 0.189894
R21728 a_n7636_8799.n398 a_n7636_8799.n341 0.189894
R21729 a_n7636_8799.n398 a_n7636_8799.n397 0.189894
R21730 a_n7636_8799.n397 a_n7636_8799.n396 0.189894
R21731 a_n7636_8799.n396 a_n7636_8799.n343 0.189894
R21732 a_n7636_8799.n344 a_n7636_8799.n343 0.189894
R21733 a_n7636_8799.n391 a_n7636_8799.n344 0.189894
R21734 a_n7636_8799.n391 a_n7636_8799.n390 0.189894
R21735 a_n7636_8799.n390 a_n7636_8799.n389 0.189894
R21736 a_n7636_8799.n389 a_n7636_8799.n346 0.189894
R21737 a_n7636_8799.n347 a_n7636_8799.n346 0.189894
R21738 a_n7636_8799.n384 a_n7636_8799.n347 0.189894
R21739 a_n7636_8799.n384 a_n7636_8799.n383 0.189894
R21740 a_n7636_8799.n383 a_n7636_8799.n382 0.189894
R21741 a_n7636_8799.n382 a_n7636_8799.n349 0.189894
R21742 a_n7636_8799.n350 a_n7636_8799.n349 0.189894
R21743 a_n7636_8799.n377 a_n7636_8799.n350 0.189894
R21744 a_n7636_8799.n377 a_n7636_8799.n376 0.189894
R21745 a_n7636_8799.n376 a_n7636_8799.n375 0.189894
R21746 a_n7636_8799.n375 a_n7636_8799.n352 0.189894
R21747 a_n7636_8799.n353 a_n7636_8799.n352 0.189894
R21748 a_n7636_8799.n370 a_n7636_8799.n353 0.189894
R21749 a_n7636_8799.n370 a_n7636_8799.n369 0.189894
R21750 a_n7636_8799.n369 a_n7636_8799.n368 0.189894
R21751 a_n7636_8799.n368 a_n7636_8799.n355 0.189894
R21752 a_n7636_8799.n356 a_n7636_8799.n355 0.189894
R21753 a_n7636_8799.n363 a_n7636_8799.n356 0.189894
R21754 a_n7636_8799.n363 a_n7636_8799.n362 0.189894
R21755 a_n7636_8799.n362 a_n7636_8799.n361 0.189894
R21756 a_n7636_8799.n47 a_n7636_8799.n42 0.189894
R21757 a_n7636_8799.n48 a_n7636_8799.n47 0.189894
R21758 a_n7636_8799.n49 a_n7636_8799.n48 0.189894
R21759 a_n7636_8799.n49 a_n7636_8799.n40 0.189894
R21760 a_n7636_8799.n53 a_n7636_8799.n40 0.189894
R21761 a_n7636_8799.n54 a_n7636_8799.n53 0.189894
R21762 a_n7636_8799.n55 a_n7636_8799.n54 0.189894
R21763 a_n7636_8799.n55 a_n7636_8799.n38 0.189894
R21764 a_n7636_8799.n59 a_n7636_8799.n38 0.189894
R21765 a_n7636_8799.n60 a_n7636_8799.n59 0.189894
R21766 a_n7636_8799.n61 a_n7636_8799.n60 0.189894
R21767 a_n7636_8799.n61 a_n7636_8799.n36 0.189894
R21768 a_n7636_8799.n65 a_n7636_8799.n36 0.189894
R21769 a_n7636_8799.n66 a_n7636_8799.n65 0.189894
R21770 a_n7636_8799.n67 a_n7636_8799.n66 0.189894
R21771 a_n7636_8799.n67 a_n7636_8799.n34 0.189894
R21772 a_n7636_8799.n71 a_n7636_8799.n34 0.189894
R21773 a_n7636_8799.n72 a_n7636_8799.n71 0.189894
R21774 a_n7636_8799.n73 a_n7636_8799.n72 0.189894
R21775 a_n7636_8799.n73 a_n7636_8799.n32 0.189894
R21776 a_n7636_8799.n77 a_n7636_8799.n32 0.189894
R21777 a_n7636_8799.n78 a_n7636_8799.n77 0.189894
R21778 a_n7636_8799.n79 a_n7636_8799.n78 0.189894
R21779 a_n7636_8799.n79 a_n7636_8799.n30 0.189894
R21780 a_n7636_8799.n83 a_n7636_8799.n30 0.189894
R21781 a_n7636_8799.n84 a_n7636_8799.n83 0.189894
R21782 a_n7636_8799.n85 a_n7636_8799.n84 0.189894
R21783 a_n7636_8799.n85 a_n7636_8799.n28 0.189894
R21784 a_n7636_8799.n89 a_n7636_8799.n28 0.189894
R21785 a_n7636_8799.n109 a_n7636_8799.n104 0.189894
R21786 a_n7636_8799.n110 a_n7636_8799.n109 0.189894
R21787 a_n7636_8799.n111 a_n7636_8799.n110 0.189894
R21788 a_n7636_8799.n111 a_n7636_8799.n102 0.189894
R21789 a_n7636_8799.n115 a_n7636_8799.n102 0.189894
R21790 a_n7636_8799.n116 a_n7636_8799.n115 0.189894
R21791 a_n7636_8799.n117 a_n7636_8799.n116 0.189894
R21792 a_n7636_8799.n117 a_n7636_8799.n100 0.189894
R21793 a_n7636_8799.n121 a_n7636_8799.n100 0.189894
R21794 a_n7636_8799.n122 a_n7636_8799.n121 0.189894
R21795 a_n7636_8799.n123 a_n7636_8799.n122 0.189894
R21796 a_n7636_8799.n123 a_n7636_8799.n98 0.189894
R21797 a_n7636_8799.n127 a_n7636_8799.n98 0.189894
R21798 a_n7636_8799.n128 a_n7636_8799.n127 0.189894
R21799 a_n7636_8799.n129 a_n7636_8799.n128 0.189894
R21800 a_n7636_8799.n129 a_n7636_8799.n96 0.189894
R21801 a_n7636_8799.n133 a_n7636_8799.n96 0.189894
R21802 a_n7636_8799.n134 a_n7636_8799.n133 0.189894
R21803 a_n7636_8799.n135 a_n7636_8799.n134 0.189894
R21804 a_n7636_8799.n135 a_n7636_8799.n94 0.189894
R21805 a_n7636_8799.n139 a_n7636_8799.n94 0.189894
R21806 a_n7636_8799.n140 a_n7636_8799.n139 0.189894
R21807 a_n7636_8799.n141 a_n7636_8799.n140 0.189894
R21808 a_n7636_8799.n141 a_n7636_8799.n92 0.189894
R21809 a_n7636_8799.n145 a_n7636_8799.n92 0.189894
R21810 a_n7636_8799.n146 a_n7636_8799.n145 0.189894
R21811 a_n7636_8799.n147 a_n7636_8799.n146 0.189894
R21812 a_n7636_8799.n147 a_n7636_8799.n90 0.189894
R21813 a_n7636_8799.n151 a_n7636_8799.n90 0.189894
R21814 a_n7636_8799.n172 a_n7636_8799.n167 0.189894
R21815 a_n7636_8799.n173 a_n7636_8799.n172 0.189894
R21816 a_n7636_8799.n174 a_n7636_8799.n173 0.189894
R21817 a_n7636_8799.n174 a_n7636_8799.n165 0.189894
R21818 a_n7636_8799.n178 a_n7636_8799.n165 0.189894
R21819 a_n7636_8799.n179 a_n7636_8799.n178 0.189894
R21820 a_n7636_8799.n180 a_n7636_8799.n179 0.189894
R21821 a_n7636_8799.n180 a_n7636_8799.n163 0.189894
R21822 a_n7636_8799.n184 a_n7636_8799.n163 0.189894
R21823 a_n7636_8799.n185 a_n7636_8799.n184 0.189894
R21824 a_n7636_8799.n186 a_n7636_8799.n185 0.189894
R21825 a_n7636_8799.n186 a_n7636_8799.n161 0.189894
R21826 a_n7636_8799.n190 a_n7636_8799.n161 0.189894
R21827 a_n7636_8799.n191 a_n7636_8799.n190 0.189894
R21828 a_n7636_8799.n192 a_n7636_8799.n191 0.189894
R21829 a_n7636_8799.n192 a_n7636_8799.n159 0.189894
R21830 a_n7636_8799.n196 a_n7636_8799.n159 0.189894
R21831 a_n7636_8799.n197 a_n7636_8799.n196 0.189894
R21832 a_n7636_8799.n198 a_n7636_8799.n197 0.189894
R21833 a_n7636_8799.n198 a_n7636_8799.n157 0.189894
R21834 a_n7636_8799.n202 a_n7636_8799.n157 0.189894
R21835 a_n7636_8799.n203 a_n7636_8799.n202 0.189894
R21836 a_n7636_8799.n204 a_n7636_8799.n203 0.189894
R21837 a_n7636_8799.n204 a_n7636_8799.n155 0.189894
R21838 a_n7636_8799.n208 a_n7636_8799.n155 0.189894
R21839 a_n7636_8799.n209 a_n7636_8799.n208 0.189894
R21840 a_n7636_8799.n210 a_n7636_8799.n209 0.189894
R21841 a_n7636_8799.n210 a_n7636_8799.n153 0.189894
R21842 a_n7636_8799.n214 a_n7636_8799.n153 0.189894
R21843 CSoutput.n19 CSoutput.t202 184.661
R21844 CSoutput.n78 CSoutput.n77 165.8
R21845 CSoutput.n76 CSoutput.n0 165.8
R21846 CSoutput.n75 CSoutput.n74 165.8
R21847 CSoutput.n73 CSoutput.n72 165.8
R21848 CSoutput.n71 CSoutput.n2 165.8
R21849 CSoutput.n69 CSoutput.n68 165.8
R21850 CSoutput.n67 CSoutput.n3 165.8
R21851 CSoutput.n66 CSoutput.n65 165.8
R21852 CSoutput.n63 CSoutput.n4 165.8
R21853 CSoutput.n61 CSoutput.n60 165.8
R21854 CSoutput.n59 CSoutput.n5 165.8
R21855 CSoutput.n58 CSoutput.n57 165.8
R21856 CSoutput.n55 CSoutput.n6 165.8
R21857 CSoutput.n54 CSoutput.n53 165.8
R21858 CSoutput.n52 CSoutput.n51 165.8
R21859 CSoutput.n50 CSoutput.n8 165.8
R21860 CSoutput.n48 CSoutput.n47 165.8
R21861 CSoutput.n46 CSoutput.n9 165.8
R21862 CSoutput.n45 CSoutput.n44 165.8
R21863 CSoutput.n42 CSoutput.n10 165.8
R21864 CSoutput.n41 CSoutput.n40 165.8
R21865 CSoutput.n39 CSoutput.n38 165.8
R21866 CSoutput.n37 CSoutput.n12 165.8
R21867 CSoutput.n35 CSoutput.n34 165.8
R21868 CSoutput.n33 CSoutput.n13 165.8
R21869 CSoutput.n32 CSoutput.n31 165.8
R21870 CSoutput.n29 CSoutput.n14 165.8
R21871 CSoutput.n28 CSoutput.n27 165.8
R21872 CSoutput.n26 CSoutput.n25 165.8
R21873 CSoutput.n24 CSoutput.n16 165.8
R21874 CSoutput.n22 CSoutput.n21 165.8
R21875 CSoutput.n20 CSoutput.n17 165.8
R21876 CSoutput.n77 CSoutput.t204 162.194
R21877 CSoutput.n18 CSoutput.t221 120.501
R21878 CSoutput.n23 CSoutput.t215 120.501
R21879 CSoutput.n15 CSoutput.t211 120.501
R21880 CSoutput.n30 CSoutput.t200 120.501
R21881 CSoutput.n36 CSoutput.t201 120.501
R21882 CSoutput.n11 CSoutput.t212 120.501
R21883 CSoutput.n43 CSoutput.t209 120.501
R21884 CSoutput.n49 CSoutput.t203 120.501
R21885 CSoutput.n7 CSoutput.t216 120.501
R21886 CSoutput.n56 CSoutput.t218 120.501
R21887 CSoutput.n62 CSoutput.t206 120.501
R21888 CSoutput.n64 CSoutput.t219 120.501
R21889 CSoutput.n70 CSoutput.t220 120.501
R21890 CSoutput.n1 CSoutput.t214 120.501
R21891 CSoutput.n330 CSoutput.n328 103.469
R21892 CSoutput.n310 CSoutput.n308 103.469
R21893 CSoutput.n291 CSoutput.n289 103.469
R21894 CSoutput.n120 CSoutput.n118 103.469
R21895 CSoutput.n100 CSoutput.n98 103.469
R21896 CSoutput.n81 CSoutput.n79 103.469
R21897 CSoutput.n344 CSoutput.n343 103.111
R21898 CSoutput.n342 CSoutput.n341 103.111
R21899 CSoutput.n340 CSoutput.n339 103.111
R21900 CSoutput.n338 CSoutput.n337 103.111
R21901 CSoutput.n336 CSoutput.n335 103.111
R21902 CSoutput.n334 CSoutput.n333 103.111
R21903 CSoutput.n332 CSoutput.n331 103.111
R21904 CSoutput.n330 CSoutput.n329 103.111
R21905 CSoutput.n326 CSoutput.n325 103.111
R21906 CSoutput.n324 CSoutput.n323 103.111
R21907 CSoutput.n322 CSoutput.n321 103.111
R21908 CSoutput.n320 CSoutput.n319 103.111
R21909 CSoutput.n318 CSoutput.n317 103.111
R21910 CSoutput.n316 CSoutput.n315 103.111
R21911 CSoutput.n314 CSoutput.n313 103.111
R21912 CSoutput.n312 CSoutput.n311 103.111
R21913 CSoutput.n310 CSoutput.n309 103.111
R21914 CSoutput.n307 CSoutput.n306 103.111
R21915 CSoutput.n305 CSoutput.n304 103.111
R21916 CSoutput.n303 CSoutput.n302 103.111
R21917 CSoutput.n301 CSoutput.n300 103.111
R21918 CSoutput.n299 CSoutput.n298 103.111
R21919 CSoutput.n297 CSoutput.n296 103.111
R21920 CSoutput.n295 CSoutput.n294 103.111
R21921 CSoutput.n293 CSoutput.n292 103.111
R21922 CSoutput.n291 CSoutput.n290 103.111
R21923 CSoutput.n120 CSoutput.n119 103.111
R21924 CSoutput.n122 CSoutput.n121 103.111
R21925 CSoutput.n124 CSoutput.n123 103.111
R21926 CSoutput.n126 CSoutput.n125 103.111
R21927 CSoutput.n128 CSoutput.n127 103.111
R21928 CSoutput.n130 CSoutput.n129 103.111
R21929 CSoutput.n132 CSoutput.n131 103.111
R21930 CSoutput.n134 CSoutput.n133 103.111
R21931 CSoutput.n136 CSoutput.n135 103.111
R21932 CSoutput.n100 CSoutput.n99 103.111
R21933 CSoutput.n102 CSoutput.n101 103.111
R21934 CSoutput.n104 CSoutput.n103 103.111
R21935 CSoutput.n106 CSoutput.n105 103.111
R21936 CSoutput.n108 CSoutput.n107 103.111
R21937 CSoutput.n110 CSoutput.n109 103.111
R21938 CSoutput.n112 CSoutput.n111 103.111
R21939 CSoutput.n114 CSoutput.n113 103.111
R21940 CSoutput.n116 CSoutput.n115 103.111
R21941 CSoutput.n81 CSoutput.n80 103.111
R21942 CSoutput.n83 CSoutput.n82 103.111
R21943 CSoutput.n85 CSoutput.n84 103.111
R21944 CSoutput.n87 CSoutput.n86 103.111
R21945 CSoutput.n89 CSoutput.n88 103.111
R21946 CSoutput.n91 CSoutput.n90 103.111
R21947 CSoutput.n93 CSoutput.n92 103.111
R21948 CSoutput.n95 CSoutput.n94 103.111
R21949 CSoutput.n97 CSoutput.n96 103.111
R21950 CSoutput.n346 CSoutput.n345 103.111
R21951 CSoutput.n370 CSoutput.n368 81.5057
R21952 CSoutput.n351 CSoutput.n349 81.5057
R21953 CSoutput.n410 CSoutput.n408 81.5057
R21954 CSoutput.n391 CSoutput.n389 81.5057
R21955 CSoutput.n386 CSoutput.n385 80.9324
R21956 CSoutput.n384 CSoutput.n383 80.9324
R21957 CSoutput.n382 CSoutput.n381 80.9324
R21958 CSoutput.n380 CSoutput.n379 80.9324
R21959 CSoutput.n378 CSoutput.n377 80.9324
R21960 CSoutput.n376 CSoutput.n375 80.9324
R21961 CSoutput.n374 CSoutput.n373 80.9324
R21962 CSoutput.n372 CSoutput.n371 80.9324
R21963 CSoutput.n370 CSoutput.n369 80.9324
R21964 CSoutput.n367 CSoutput.n366 80.9324
R21965 CSoutput.n365 CSoutput.n364 80.9324
R21966 CSoutput.n363 CSoutput.n362 80.9324
R21967 CSoutput.n361 CSoutput.n360 80.9324
R21968 CSoutput.n359 CSoutput.n358 80.9324
R21969 CSoutput.n357 CSoutput.n356 80.9324
R21970 CSoutput.n355 CSoutput.n354 80.9324
R21971 CSoutput.n353 CSoutput.n352 80.9324
R21972 CSoutput.n351 CSoutput.n350 80.9324
R21973 CSoutput.n410 CSoutput.n409 80.9324
R21974 CSoutput.n412 CSoutput.n411 80.9324
R21975 CSoutput.n414 CSoutput.n413 80.9324
R21976 CSoutput.n416 CSoutput.n415 80.9324
R21977 CSoutput.n418 CSoutput.n417 80.9324
R21978 CSoutput.n420 CSoutput.n419 80.9324
R21979 CSoutput.n422 CSoutput.n421 80.9324
R21980 CSoutput.n424 CSoutput.n423 80.9324
R21981 CSoutput.n426 CSoutput.n425 80.9324
R21982 CSoutput.n391 CSoutput.n390 80.9324
R21983 CSoutput.n393 CSoutput.n392 80.9324
R21984 CSoutput.n395 CSoutput.n394 80.9324
R21985 CSoutput.n397 CSoutput.n396 80.9324
R21986 CSoutput.n399 CSoutput.n398 80.9324
R21987 CSoutput.n401 CSoutput.n400 80.9324
R21988 CSoutput.n403 CSoutput.n402 80.9324
R21989 CSoutput.n405 CSoutput.n404 80.9324
R21990 CSoutput.n407 CSoutput.n406 80.9324
R21991 CSoutput.n25 CSoutput.n24 48.1486
R21992 CSoutput.n69 CSoutput.n3 48.1486
R21993 CSoutput.n38 CSoutput.n37 48.1486
R21994 CSoutput.n42 CSoutput.n41 48.1486
R21995 CSoutput.n51 CSoutput.n50 48.1486
R21996 CSoutput.n55 CSoutput.n54 48.1486
R21997 CSoutput.n22 CSoutput.n17 46.462
R21998 CSoutput.n72 CSoutput.n71 46.462
R21999 CSoutput.n20 CSoutput.n19 44.9055
R22000 CSoutput.n29 CSoutput.n28 43.7635
R22001 CSoutput.n65 CSoutput.n63 43.7635
R22002 CSoutput.n35 CSoutput.n13 41.7396
R22003 CSoutput.n57 CSoutput.n5 41.7396
R22004 CSoutput.n44 CSoutput.n9 37.0171
R22005 CSoutput.n48 CSoutput.n9 37.0171
R22006 CSoutput.n76 CSoutput.n75 34.9932
R22007 CSoutput.n31 CSoutput.n13 32.2947
R22008 CSoutput.n61 CSoutput.n5 32.2947
R22009 CSoutput.n30 CSoutput.n29 29.6014
R22010 CSoutput.n63 CSoutput.n62 29.6014
R22011 CSoutput.n19 CSoutput.n18 28.4085
R22012 CSoutput.n18 CSoutput.n17 25.1176
R22013 CSoutput.n72 CSoutput.n1 25.1176
R22014 CSoutput.n43 CSoutput.n42 22.0922
R22015 CSoutput.n50 CSoutput.n49 22.0922
R22016 CSoutput.n77 CSoutput.n76 21.8586
R22017 CSoutput.n37 CSoutput.n36 18.9681
R22018 CSoutput.n56 CSoutput.n55 18.9681
R22019 CSoutput.n25 CSoutput.n15 17.6292
R22020 CSoutput.n64 CSoutput.n3 17.6292
R22021 CSoutput.n24 CSoutput.n23 15.844
R22022 CSoutput.n70 CSoutput.n69 15.844
R22023 CSoutput.n38 CSoutput.n11 14.5051
R22024 CSoutput.n54 CSoutput.n7 14.5051
R22025 CSoutput.n429 CSoutput.n78 11.6139
R22026 CSoutput.n41 CSoutput.n11 11.3811
R22027 CSoutput.n51 CSoutput.n7 11.3811
R22028 CSoutput.n23 CSoutput.n22 10.0422
R22029 CSoutput.n71 CSoutput.n70 10.0422
R22030 CSoutput.n327 CSoutput.n307 9.25285
R22031 CSoutput.n117 CSoutput.n97 9.25285
R22032 CSoutput.n388 CSoutput.n348 9.09467
R22033 CSoutput.n387 CSoutput.n367 8.97993
R22034 CSoutput.n427 CSoutput.n407 8.97993
R22035 CSoutput.n28 CSoutput.n15 8.25698
R22036 CSoutput.n65 CSoutput.n64 8.25698
R22037 CSoutput.n388 CSoutput.n387 7.89345
R22038 CSoutput.n428 CSoutput.n427 7.89345
R22039 CSoutput.n348 CSoutput.n347 7.12641
R22040 CSoutput.n138 CSoutput.n137 7.12641
R22041 CSoutput.n36 CSoutput.n35 6.91809
R22042 CSoutput.n57 CSoutput.n56 6.91809
R22043 CSoutput.n429 CSoutput.n138 5.50223
R22044 CSoutput.n387 CSoutput.n386 5.25266
R22045 CSoutput.n427 CSoutput.n426 5.25266
R22046 CSoutput.n347 CSoutput.n346 5.1449
R22047 CSoutput.n327 CSoutput.n326 5.1449
R22048 CSoutput.n137 CSoutput.n136 5.1449
R22049 CSoutput.n117 CSoutput.n116 5.1449
R22050 CSoutput.n229 CSoutput.n182 4.5005
R22051 CSoutput.n198 CSoutput.n182 4.5005
R22052 CSoutput.n193 CSoutput.n177 4.5005
R22053 CSoutput.n193 CSoutput.n179 4.5005
R22054 CSoutput.n193 CSoutput.n176 4.5005
R22055 CSoutput.n193 CSoutput.n180 4.5005
R22056 CSoutput.n193 CSoutput.n175 4.5005
R22057 CSoutput.n193 CSoutput.t207 4.5005
R22058 CSoutput.n193 CSoutput.n174 4.5005
R22059 CSoutput.n193 CSoutput.n181 4.5005
R22060 CSoutput.n193 CSoutput.n182 4.5005
R22061 CSoutput.n191 CSoutput.n177 4.5005
R22062 CSoutput.n191 CSoutput.n179 4.5005
R22063 CSoutput.n191 CSoutput.n176 4.5005
R22064 CSoutput.n191 CSoutput.n180 4.5005
R22065 CSoutput.n191 CSoutput.n175 4.5005
R22066 CSoutput.n191 CSoutput.t207 4.5005
R22067 CSoutput.n191 CSoutput.n174 4.5005
R22068 CSoutput.n191 CSoutput.n181 4.5005
R22069 CSoutput.n191 CSoutput.n182 4.5005
R22070 CSoutput.n190 CSoutput.n177 4.5005
R22071 CSoutput.n190 CSoutput.n179 4.5005
R22072 CSoutput.n190 CSoutput.n176 4.5005
R22073 CSoutput.n190 CSoutput.n180 4.5005
R22074 CSoutput.n190 CSoutput.n175 4.5005
R22075 CSoutput.n190 CSoutput.t207 4.5005
R22076 CSoutput.n190 CSoutput.n174 4.5005
R22077 CSoutput.n190 CSoutput.n181 4.5005
R22078 CSoutput.n190 CSoutput.n182 4.5005
R22079 CSoutput.n275 CSoutput.n177 4.5005
R22080 CSoutput.n275 CSoutput.n179 4.5005
R22081 CSoutput.n275 CSoutput.n176 4.5005
R22082 CSoutput.n275 CSoutput.n180 4.5005
R22083 CSoutput.n275 CSoutput.n175 4.5005
R22084 CSoutput.n275 CSoutput.t207 4.5005
R22085 CSoutput.n275 CSoutput.n174 4.5005
R22086 CSoutput.n275 CSoutput.n181 4.5005
R22087 CSoutput.n275 CSoutput.n182 4.5005
R22088 CSoutput.n273 CSoutput.n177 4.5005
R22089 CSoutput.n273 CSoutput.n179 4.5005
R22090 CSoutput.n273 CSoutput.n176 4.5005
R22091 CSoutput.n273 CSoutput.n180 4.5005
R22092 CSoutput.n273 CSoutput.n175 4.5005
R22093 CSoutput.n273 CSoutput.t207 4.5005
R22094 CSoutput.n273 CSoutput.n174 4.5005
R22095 CSoutput.n273 CSoutput.n181 4.5005
R22096 CSoutput.n271 CSoutput.n177 4.5005
R22097 CSoutput.n271 CSoutput.n179 4.5005
R22098 CSoutput.n271 CSoutput.n176 4.5005
R22099 CSoutput.n271 CSoutput.n180 4.5005
R22100 CSoutput.n271 CSoutput.n175 4.5005
R22101 CSoutput.n271 CSoutput.t207 4.5005
R22102 CSoutput.n271 CSoutput.n174 4.5005
R22103 CSoutput.n271 CSoutput.n181 4.5005
R22104 CSoutput.n201 CSoutput.n177 4.5005
R22105 CSoutput.n201 CSoutput.n179 4.5005
R22106 CSoutput.n201 CSoutput.n176 4.5005
R22107 CSoutput.n201 CSoutput.n180 4.5005
R22108 CSoutput.n201 CSoutput.n175 4.5005
R22109 CSoutput.n201 CSoutput.t207 4.5005
R22110 CSoutput.n201 CSoutput.n174 4.5005
R22111 CSoutput.n201 CSoutput.n181 4.5005
R22112 CSoutput.n201 CSoutput.n182 4.5005
R22113 CSoutput.n200 CSoutput.n177 4.5005
R22114 CSoutput.n200 CSoutput.n179 4.5005
R22115 CSoutput.n200 CSoutput.n176 4.5005
R22116 CSoutput.n200 CSoutput.n180 4.5005
R22117 CSoutput.n200 CSoutput.n175 4.5005
R22118 CSoutput.n200 CSoutput.t207 4.5005
R22119 CSoutput.n200 CSoutput.n174 4.5005
R22120 CSoutput.n200 CSoutput.n181 4.5005
R22121 CSoutput.n200 CSoutput.n182 4.5005
R22122 CSoutput.n204 CSoutput.n177 4.5005
R22123 CSoutput.n204 CSoutput.n179 4.5005
R22124 CSoutput.n204 CSoutput.n176 4.5005
R22125 CSoutput.n204 CSoutput.n180 4.5005
R22126 CSoutput.n204 CSoutput.n175 4.5005
R22127 CSoutput.n204 CSoutput.t207 4.5005
R22128 CSoutput.n204 CSoutput.n174 4.5005
R22129 CSoutput.n204 CSoutput.n181 4.5005
R22130 CSoutput.n204 CSoutput.n182 4.5005
R22131 CSoutput.n203 CSoutput.n177 4.5005
R22132 CSoutput.n203 CSoutput.n179 4.5005
R22133 CSoutput.n203 CSoutput.n176 4.5005
R22134 CSoutput.n203 CSoutput.n180 4.5005
R22135 CSoutput.n203 CSoutput.n175 4.5005
R22136 CSoutput.n203 CSoutput.t207 4.5005
R22137 CSoutput.n203 CSoutput.n174 4.5005
R22138 CSoutput.n203 CSoutput.n181 4.5005
R22139 CSoutput.n203 CSoutput.n182 4.5005
R22140 CSoutput.n186 CSoutput.n177 4.5005
R22141 CSoutput.n186 CSoutput.n179 4.5005
R22142 CSoutput.n186 CSoutput.n176 4.5005
R22143 CSoutput.n186 CSoutput.n180 4.5005
R22144 CSoutput.n186 CSoutput.n175 4.5005
R22145 CSoutput.n186 CSoutput.t207 4.5005
R22146 CSoutput.n186 CSoutput.n174 4.5005
R22147 CSoutput.n186 CSoutput.n181 4.5005
R22148 CSoutput.n186 CSoutput.n182 4.5005
R22149 CSoutput.n278 CSoutput.n177 4.5005
R22150 CSoutput.n278 CSoutput.n179 4.5005
R22151 CSoutput.n278 CSoutput.n176 4.5005
R22152 CSoutput.n278 CSoutput.n180 4.5005
R22153 CSoutput.n278 CSoutput.n175 4.5005
R22154 CSoutput.n278 CSoutput.t207 4.5005
R22155 CSoutput.n278 CSoutput.n174 4.5005
R22156 CSoutput.n278 CSoutput.n181 4.5005
R22157 CSoutput.n278 CSoutput.n182 4.5005
R22158 CSoutput.n265 CSoutput.n236 4.5005
R22159 CSoutput.n265 CSoutput.n242 4.5005
R22160 CSoutput.n223 CSoutput.n212 4.5005
R22161 CSoutput.n223 CSoutput.n214 4.5005
R22162 CSoutput.n223 CSoutput.n211 4.5005
R22163 CSoutput.n223 CSoutput.n215 4.5005
R22164 CSoutput.n223 CSoutput.n210 4.5005
R22165 CSoutput.n223 CSoutput.t208 4.5005
R22166 CSoutput.n223 CSoutput.n209 4.5005
R22167 CSoutput.n223 CSoutput.n216 4.5005
R22168 CSoutput.n265 CSoutput.n223 4.5005
R22169 CSoutput.n244 CSoutput.n212 4.5005
R22170 CSoutput.n244 CSoutput.n214 4.5005
R22171 CSoutput.n244 CSoutput.n211 4.5005
R22172 CSoutput.n244 CSoutput.n215 4.5005
R22173 CSoutput.n244 CSoutput.n210 4.5005
R22174 CSoutput.n244 CSoutput.t208 4.5005
R22175 CSoutput.n244 CSoutput.n209 4.5005
R22176 CSoutput.n244 CSoutput.n216 4.5005
R22177 CSoutput.n265 CSoutput.n244 4.5005
R22178 CSoutput.n222 CSoutput.n212 4.5005
R22179 CSoutput.n222 CSoutput.n214 4.5005
R22180 CSoutput.n222 CSoutput.n211 4.5005
R22181 CSoutput.n222 CSoutput.n215 4.5005
R22182 CSoutput.n222 CSoutput.n210 4.5005
R22183 CSoutput.n222 CSoutput.t208 4.5005
R22184 CSoutput.n222 CSoutput.n209 4.5005
R22185 CSoutput.n222 CSoutput.n216 4.5005
R22186 CSoutput.n265 CSoutput.n222 4.5005
R22187 CSoutput.n246 CSoutput.n212 4.5005
R22188 CSoutput.n246 CSoutput.n214 4.5005
R22189 CSoutput.n246 CSoutput.n211 4.5005
R22190 CSoutput.n246 CSoutput.n215 4.5005
R22191 CSoutput.n246 CSoutput.n210 4.5005
R22192 CSoutput.n246 CSoutput.t208 4.5005
R22193 CSoutput.n246 CSoutput.n209 4.5005
R22194 CSoutput.n246 CSoutput.n216 4.5005
R22195 CSoutput.n265 CSoutput.n246 4.5005
R22196 CSoutput.n212 CSoutput.n207 4.5005
R22197 CSoutput.n214 CSoutput.n207 4.5005
R22198 CSoutput.n211 CSoutput.n207 4.5005
R22199 CSoutput.n215 CSoutput.n207 4.5005
R22200 CSoutput.n210 CSoutput.n207 4.5005
R22201 CSoutput.t208 CSoutput.n207 4.5005
R22202 CSoutput.n209 CSoutput.n207 4.5005
R22203 CSoutput.n216 CSoutput.n207 4.5005
R22204 CSoutput.n268 CSoutput.n212 4.5005
R22205 CSoutput.n268 CSoutput.n214 4.5005
R22206 CSoutput.n268 CSoutput.n211 4.5005
R22207 CSoutput.n268 CSoutput.n215 4.5005
R22208 CSoutput.n268 CSoutput.n210 4.5005
R22209 CSoutput.n268 CSoutput.t208 4.5005
R22210 CSoutput.n268 CSoutput.n209 4.5005
R22211 CSoutput.n268 CSoutput.n216 4.5005
R22212 CSoutput.n266 CSoutput.n212 4.5005
R22213 CSoutput.n266 CSoutput.n214 4.5005
R22214 CSoutput.n266 CSoutput.n211 4.5005
R22215 CSoutput.n266 CSoutput.n215 4.5005
R22216 CSoutput.n266 CSoutput.n210 4.5005
R22217 CSoutput.n266 CSoutput.t208 4.5005
R22218 CSoutput.n266 CSoutput.n209 4.5005
R22219 CSoutput.n266 CSoutput.n216 4.5005
R22220 CSoutput.n266 CSoutput.n265 4.5005
R22221 CSoutput.n248 CSoutput.n212 4.5005
R22222 CSoutput.n248 CSoutput.n214 4.5005
R22223 CSoutput.n248 CSoutput.n211 4.5005
R22224 CSoutput.n248 CSoutput.n215 4.5005
R22225 CSoutput.n248 CSoutput.n210 4.5005
R22226 CSoutput.n248 CSoutput.t208 4.5005
R22227 CSoutput.n248 CSoutput.n209 4.5005
R22228 CSoutput.n248 CSoutput.n216 4.5005
R22229 CSoutput.n265 CSoutput.n248 4.5005
R22230 CSoutput.n220 CSoutput.n212 4.5005
R22231 CSoutput.n220 CSoutput.n214 4.5005
R22232 CSoutput.n220 CSoutput.n211 4.5005
R22233 CSoutput.n220 CSoutput.n215 4.5005
R22234 CSoutput.n220 CSoutput.n210 4.5005
R22235 CSoutput.n220 CSoutput.t208 4.5005
R22236 CSoutput.n220 CSoutput.n209 4.5005
R22237 CSoutput.n220 CSoutput.n216 4.5005
R22238 CSoutput.n265 CSoutput.n220 4.5005
R22239 CSoutput.n250 CSoutput.n212 4.5005
R22240 CSoutput.n250 CSoutput.n214 4.5005
R22241 CSoutput.n250 CSoutput.n211 4.5005
R22242 CSoutput.n250 CSoutput.n215 4.5005
R22243 CSoutput.n250 CSoutput.n210 4.5005
R22244 CSoutput.n250 CSoutput.t208 4.5005
R22245 CSoutput.n250 CSoutput.n209 4.5005
R22246 CSoutput.n250 CSoutput.n216 4.5005
R22247 CSoutput.n265 CSoutput.n250 4.5005
R22248 CSoutput.n219 CSoutput.n212 4.5005
R22249 CSoutput.n219 CSoutput.n214 4.5005
R22250 CSoutput.n219 CSoutput.n211 4.5005
R22251 CSoutput.n219 CSoutput.n215 4.5005
R22252 CSoutput.n219 CSoutput.n210 4.5005
R22253 CSoutput.n219 CSoutput.t208 4.5005
R22254 CSoutput.n219 CSoutput.n209 4.5005
R22255 CSoutput.n219 CSoutput.n216 4.5005
R22256 CSoutput.n265 CSoutput.n219 4.5005
R22257 CSoutput.n264 CSoutput.n212 4.5005
R22258 CSoutput.n264 CSoutput.n214 4.5005
R22259 CSoutput.n264 CSoutput.n211 4.5005
R22260 CSoutput.n264 CSoutput.n215 4.5005
R22261 CSoutput.n264 CSoutput.n210 4.5005
R22262 CSoutput.n264 CSoutput.t208 4.5005
R22263 CSoutput.n264 CSoutput.n209 4.5005
R22264 CSoutput.n264 CSoutput.n216 4.5005
R22265 CSoutput.n265 CSoutput.n264 4.5005
R22266 CSoutput.n263 CSoutput.n148 4.5005
R22267 CSoutput.n164 CSoutput.n148 4.5005
R22268 CSoutput.n159 CSoutput.n143 4.5005
R22269 CSoutput.n159 CSoutput.n145 4.5005
R22270 CSoutput.n159 CSoutput.n142 4.5005
R22271 CSoutput.n159 CSoutput.n146 4.5005
R22272 CSoutput.n159 CSoutput.n141 4.5005
R22273 CSoutput.n159 CSoutput.t210 4.5005
R22274 CSoutput.n159 CSoutput.n140 4.5005
R22275 CSoutput.n159 CSoutput.n147 4.5005
R22276 CSoutput.n159 CSoutput.n148 4.5005
R22277 CSoutput.n157 CSoutput.n143 4.5005
R22278 CSoutput.n157 CSoutput.n145 4.5005
R22279 CSoutput.n157 CSoutput.n142 4.5005
R22280 CSoutput.n157 CSoutput.n146 4.5005
R22281 CSoutput.n157 CSoutput.n141 4.5005
R22282 CSoutput.n157 CSoutput.t210 4.5005
R22283 CSoutput.n157 CSoutput.n140 4.5005
R22284 CSoutput.n157 CSoutput.n147 4.5005
R22285 CSoutput.n157 CSoutput.n148 4.5005
R22286 CSoutput.n156 CSoutput.n143 4.5005
R22287 CSoutput.n156 CSoutput.n145 4.5005
R22288 CSoutput.n156 CSoutput.n142 4.5005
R22289 CSoutput.n156 CSoutput.n146 4.5005
R22290 CSoutput.n156 CSoutput.n141 4.5005
R22291 CSoutput.n156 CSoutput.t210 4.5005
R22292 CSoutput.n156 CSoutput.n140 4.5005
R22293 CSoutput.n156 CSoutput.n147 4.5005
R22294 CSoutput.n156 CSoutput.n148 4.5005
R22295 CSoutput.n285 CSoutput.n143 4.5005
R22296 CSoutput.n285 CSoutput.n145 4.5005
R22297 CSoutput.n285 CSoutput.n142 4.5005
R22298 CSoutput.n285 CSoutput.n146 4.5005
R22299 CSoutput.n285 CSoutput.n141 4.5005
R22300 CSoutput.n285 CSoutput.t210 4.5005
R22301 CSoutput.n285 CSoutput.n140 4.5005
R22302 CSoutput.n285 CSoutput.n147 4.5005
R22303 CSoutput.n285 CSoutput.n148 4.5005
R22304 CSoutput.n283 CSoutput.n143 4.5005
R22305 CSoutput.n283 CSoutput.n145 4.5005
R22306 CSoutput.n283 CSoutput.n142 4.5005
R22307 CSoutput.n283 CSoutput.n146 4.5005
R22308 CSoutput.n283 CSoutput.n141 4.5005
R22309 CSoutput.n283 CSoutput.t210 4.5005
R22310 CSoutput.n283 CSoutput.n140 4.5005
R22311 CSoutput.n283 CSoutput.n147 4.5005
R22312 CSoutput.n281 CSoutput.n143 4.5005
R22313 CSoutput.n281 CSoutput.n145 4.5005
R22314 CSoutput.n281 CSoutput.n142 4.5005
R22315 CSoutput.n281 CSoutput.n146 4.5005
R22316 CSoutput.n281 CSoutput.n141 4.5005
R22317 CSoutput.n281 CSoutput.t210 4.5005
R22318 CSoutput.n281 CSoutput.n140 4.5005
R22319 CSoutput.n281 CSoutput.n147 4.5005
R22320 CSoutput.n167 CSoutput.n143 4.5005
R22321 CSoutput.n167 CSoutput.n145 4.5005
R22322 CSoutput.n167 CSoutput.n142 4.5005
R22323 CSoutput.n167 CSoutput.n146 4.5005
R22324 CSoutput.n167 CSoutput.n141 4.5005
R22325 CSoutput.n167 CSoutput.t210 4.5005
R22326 CSoutput.n167 CSoutput.n140 4.5005
R22327 CSoutput.n167 CSoutput.n147 4.5005
R22328 CSoutput.n167 CSoutput.n148 4.5005
R22329 CSoutput.n166 CSoutput.n143 4.5005
R22330 CSoutput.n166 CSoutput.n145 4.5005
R22331 CSoutput.n166 CSoutput.n142 4.5005
R22332 CSoutput.n166 CSoutput.n146 4.5005
R22333 CSoutput.n166 CSoutput.n141 4.5005
R22334 CSoutput.n166 CSoutput.t210 4.5005
R22335 CSoutput.n166 CSoutput.n140 4.5005
R22336 CSoutput.n166 CSoutput.n147 4.5005
R22337 CSoutput.n166 CSoutput.n148 4.5005
R22338 CSoutput.n170 CSoutput.n143 4.5005
R22339 CSoutput.n170 CSoutput.n145 4.5005
R22340 CSoutput.n170 CSoutput.n142 4.5005
R22341 CSoutput.n170 CSoutput.n146 4.5005
R22342 CSoutput.n170 CSoutput.n141 4.5005
R22343 CSoutput.n170 CSoutput.t210 4.5005
R22344 CSoutput.n170 CSoutput.n140 4.5005
R22345 CSoutput.n170 CSoutput.n147 4.5005
R22346 CSoutput.n170 CSoutput.n148 4.5005
R22347 CSoutput.n169 CSoutput.n143 4.5005
R22348 CSoutput.n169 CSoutput.n145 4.5005
R22349 CSoutput.n169 CSoutput.n142 4.5005
R22350 CSoutput.n169 CSoutput.n146 4.5005
R22351 CSoutput.n169 CSoutput.n141 4.5005
R22352 CSoutput.n169 CSoutput.t210 4.5005
R22353 CSoutput.n169 CSoutput.n140 4.5005
R22354 CSoutput.n169 CSoutput.n147 4.5005
R22355 CSoutput.n169 CSoutput.n148 4.5005
R22356 CSoutput.n152 CSoutput.n143 4.5005
R22357 CSoutput.n152 CSoutput.n145 4.5005
R22358 CSoutput.n152 CSoutput.n142 4.5005
R22359 CSoutput.n152 CSoutput.n146 4.5005
R22360 CSoutput.n152 CSoutput.n141 4.5005
R22361 CSoutput.n152 CSoutput.t210 4.5005
R22362 CSoutput.n152 CSoutput.n140 4.5005
R22363 CSoutput.n152 CSoutput.n147 4.5005
R22364 CSoutput.n152 CSoutput.n148 4.5005
R22365 CSoutput.n288 CSoutput.n143 4.5005
R22366 CSoutput.n288 CSoutput.n145 4.5005
R22367 CSoutput.n288 CSoutput.n142 4.5005
R22368 CSoutput.n288 CSoutput.n146 4.5005
R22369 CSoutput.n288 CSoutput.n141 4.5005
R22370 CSoutput.n288 CSoutput.t210 4.5005
R22371 CSoutput.n288 CSoutput.n140 4.5005
R22372 CSoutput.n288 CSoutput.n147 4.5005
R22373 CSoutput.n288 CSoutput.n148 4.5005
R22374 CSoutput.n347 CSoutput.n327 4.10845
R22375 CSoutput.n137 CSoutput.n117 4.10845
R22376 CSoutput.n345 CSoutput.t72 4.06363
R22377 CSoutput.n345 CSoutput.t96 4.06363
R22378 CSoutput.n343 CSoutput.t117 4.06363
R22379 CSoutput.n343 CSoutput.t30 4.06363
R22380 CSoutput.n341 CSoutput.t34 4.06363
R22381 CSoutput.n341 CSoutput.t100 4.06363
R22382 CSoutput.n339 CSoutput.t119 4.06363
R22383 CSoutput.n339 CSoutput.t120 4.06363
R22384 CSoutput.n337 CSoutput.t50 4.06363
R22385 CSoutput.n337 CSoutput.t51 4.06363
R22386 CSoutput.n335 CSoutput.t56 4.06363
R22387 CSoutput.n335 CSoutput.t121 4.06363
R22388 CSoutput.n333 CSoutput.t20 4.06363
R22389 CSoutput.n333 CSoutput.t54 4.06363
R22390 CSoutput.n331 CSoutput.t71 4.06363
R22391 CSoutput.n331 CSoutput.t95 4.06363
R22392 CSoutput.n329 CSoutput.t102 4.06363
R22393 CSoutput.n329 CSoutput.t26 4.06363
R22394 CSoutput.n328 CSoutput.t74 4.06363
R22395 CSoutput.n328 CSoutput.t75 4.06363
R22396 CSoutput.n325 CSoutput.t58 4.06363
R22397 CSoutput.n325 CSoutput.t84 4.06363
R22398 CSoutput.n323 CSoutput.t104 4.06363
R22399 CSoutput.n323 CSoutput.t16 4.06363
R22400 CSoutput.n321 CSoutput.t17 4.06363
R22401 CSoutput.n321 CSoutput.t86 4.06363
R22402 CSoutput.n319 CSoutput.t107 4.06363
R22403 CSoutput.n319 CSoutput.t108 4.06363
R22404 CSoutput.n317 CSoutput.t38 4.06363
R22405 CSoutput.n317 CSoutput.t39 4.06363
R22406 CSoutput.n315 CSoutput.t42 4.06363
R22407 CSoutput.n315 CSoutput.t111 4.06363
R22408 CSoutput.n313 CSoutput.t125 4.06363
R22409 CSoutput.n313 CSoutput.t41 4.06363
R22410 CSoutput.n311 CSoutput.t57 4.06363
R22411 CSoutput.n311 CSoutput.t85 4.06363
R22412 CSoutput.n309 CSoutput.t87 4.06363
R22413 CSoutput.n309 CSoutput.t11 4.06363
R22414 CSoutput.n308 CSoutput.t64 4.06363
R22415 CSoutput.n308 CSoutput.t65 4.06363
R22416 CSoutput.n306 CSoutput.t93 4.06363
R22417 CSoutput.n306 CSoutput.t47 4.06363
R22418 CSoutput.n304 CSoutput.t80 4.06363
R22419 CSoutput.n304 CSoutput.t29 4.06363
R22420 CSoutput.n302 CSoutput.t105 4.06363
R22421 CSoutput.n302 CSoutput.t21 4.06363
R22422 CSoutput.n300 CSoutput.t61 4.06363
R22423 CSoutput.n300 CSoutput.t40 4.06363
R22424 CSoutput.n298 CSoutput.t43 4.06363
R22425 CSoutput.n298 CSoutput.t18 4.06363
R22426 CSoutput.n296 CSoutput.t92 4.06363
R22427 CSoutput.n296 CSoutput.t12 4.06363
R22428 CSoutput.n294 CSoutput.t52 4.06363
R22429 CSoutput.n294 CSoutput.t116 4.06363
R22430 CSoutput.n292 CSoutput.t35 4.06363
R22431 CSoutput.n292 CSoutput.t98 4.06363
R22432 CSoutput.n290 CSoutput.t59 4.06363
R22433 CSoutput.n290 CSoutput.t122 4.06363
R22434 CSoutput.n289 CSoutput.t7 4.06363
R22435 CSoutput.n289 CSoutput.t109 4.06363
R22436 CSoutput.n118 CSoutput.t115 4.06363
R22437 CSoutput.n118 CSoutput.t114 4.06363
R22438 CSoutput.n119 CSoutput.t94 4.06363
R22439 CSoutput.n119 CSoutput.t28 4.06363
R22440 CSoutput.n121 CSoutput.t25 4.06363
R22441 CSoutput.n121 CSoutput.t112 4.06363
R22442 CSoutput.n123 CSoutput.t91 4.06363
R22443 CSoutput.n123 CSoutput.t68 4.06363
R22444 CSoutput.n125 CSoutput.t49 4.06363
R22445 CSoutput.n125 CSoutput.t124 4.06363
R22446 CSoutput.n127 CSoutput.t89 4.06363
R22447 CSoutput.n127 CSoutput.t88 4.06363
R22448 CSoutput.n129 CSoutput.t76 4.06363
R22449 CSoutput.n129 CSoutput.t46 4.06363
R22450 CSoutput.n131 CSoutput.t27 4.06363
R22451 CSoutput.n131 CSoutput.t77 4.06363
R22452 CSoutput.n133 CSoutput.t73 4.06363
R22453 CSoutput.n133 CSoutput.t44 4.06363
R22454 CSoutput.n135 CSoutput.t24 4.06363
R22455 CSoutput.n135 CSoutput.t23 4.06363
R22456 CSoutput.n98 CSoutput.t103 4.06363
R22457 CSoutput.n98 CSoutput.t101 4.06363
R22458 CSoutput.n99 CSoutput.t83 4.06363
R22459 CSoutput.n99 CSoutput.t15 4.06363
R22460 CSoutput.n101 CSoutput.t9 4.06363
R22461 CSoutput.n101 CSoutput.t97 4.06363
R22462 CSoutput.n103 CSoutput.t82 4.06363
R22463 CSoutput.n103 CSoutput.t55 4.06363
R22464 CSoutput.n105 CSoutput.t37 4.06363
R22465 CSoutput.n105 CSoutput.t113 4.06363
R22466 CSoutput.n107 CSoutput.t79 4.06363
R22467 CSoutput.n107 CSoutput.t78 4.06363
R22468 CSoutput.n109 CSoutput.t66 4.06363
R22469 CSoutput.n109 CSoutput.t33 4.06363
R22470 CSoutput.n111 CSoutput.t13 4.06363
R22471 CSoutput.n111 CSoutput.t67 4.06363
R22472 CSoutput.n113 CSoutput.t63 4.06363
R22473 CSoutput.n113 CSoutput.t31 4.06363
R22474 CSoutput.n115 CSoutput.t10 4.06363
R22475 CSoutput.n115 CSoutput.t6 4.06363
R22476 CSoutput.n79 CSoutput.t110 4.06363
R22477 CSoutput.n79 CSoutput.t8 4.06363
R22478 CSoutput.n80 CSoutput.t90 4.06363
R22479 CSoutput.n80 CSoutput.t60 4.06363
R22480 CSoutput.n82 CSoutput.t99 4.06363
R22481 CSoutput.n82 CSoutput.t36 4.06363
R22482 CSoutput.n84 CSoutput.t118 4.06363
R22483 CSoutput.n84 CSoutput.t53 4.06363
R22484 CSoutput.n86 CSoutput.t14 4.06363
R22485 CSoutput.n86 CSoutput.t69 4.06363
R22486 CSoutput.n88 CSoutput.t19 4.06363
R22487 CSoutput.n88 CSoutput.t45 4.06363
R22488 CSoutput.n90 CSoutput.t123 4.06363
R22489 CSoutput.n90 CSoutput.t62 4.06363
R22490 CSoutput.n92 CSoutput.t22 4.06363
R22491 CSoutput.n92 CSoutput.t106 4.06363
R22492 CSoutput.n94 CSoutput.t32 4.06363
R22493 CSoutput.n94 CSoutput.t81 4.06363
R22494 CSoutput.n96 CSoutput.t48 4.06363
R22495 CSoutput.n96 CSoutput.t70 4.06363
R22496 CSoutput.n44 CSoutput.n43 3.79402
R22497 CSoutput.n49 CSoutput.n48 3.79402
R22498 CSoutput.n428 CSoutput.n388 3.71319
R22499 CSoutput.n429 CSoutput.n428 3.57343
R22500 CSoutput.n385 CSoutput.t151 2.82907
R22501 CSoutput.n385 CSoutput.t193 2.82907
R22502 CSoutput.n383 CSoutput.t134 2.82907
R22503 CSoutput.n383 CSoutput.t2 2.82907
R22504 CSoutput.n381 CSoutput.t165 2.82907
R22505 CSoutput.n381 CSoutput.t181 2.82907
R22506 CSoutput.n379 CSoutput.t192 2.82907
R22507 CSoutput.n379 CSoutput.t195 2.82907
R22508 CSoutput.n377 CSoutput.t172 2.82907
R22509 CSoutput.n377 CSoutput.t188 2.82907
R22510 CSoutput.n375 CSoutput.t186 2.82907
R22511 CSoutput.n375 CSoutput.t194 2.82907
R22512 CSoutput.n373 CSoutput.t150 2.82907
R22513 CSoutput.n373 CSoutput.t5 2.82907
R22514 CSoutput.n371 CSoutput.t138 2.82907
R22515 CSoutput.n371 CSoutput.t149 2.82907
R22516 CSoutput.n369 CSoutput.t0 2.82907
R22517 CSoutput.n369 CSoutput.t180 2.82907
R22518 CSoutput.n368 CSoutput.t159 2.82907
R22519 CSoutput.n368 CSoutput.t185 2.82907
R22520 CSoutput.n366 CSoutput.t161 2.82907
R22521 CSoutput.n366 CSoutput.t168 2.82907
R22522 CSoutput.n364 CSoutput.t157 2.82907
R22523 CSoutput.n364 CSoutput.t154 2.82907
R22524 CSoutput.n362 CSoutput.t133 2.82907
R22525 CSoutput.n362 CSoutput.t170 2.82907
R22526 CSoutput.n360 CSoutput.t184 2.82907
R22527 CSoutput.n360 CSoutput.t198 2.82907
R22528 CSoutput.n358 CSoutput.t166 2.82907
R22529 CSoutput.n358 CSoutput.t158 2.82907
R22530 CSoutput.n356 CSoutput.t1 2.82907
R22531 CSoutput.n356 CSoutput.t139 2.82907
R22532 CSoutput.n354 CSoutput.t160 2.82907
R22533 CSoutput.n354 CSoutput.t164 2.82907
R22534 CSoutput.n352 CSoutput.t130 2.82907
R22535 CSoutput.n352 CSoutput.t152 2.82907
R22536 CSoutput.n350 CSoutput.t127 2.82907
R22537 CSoutput.n350 CSoutput.t190 2.82907
R22538 CSoutput.n349 CSoutput.t171 2.82907
R22539 CSoutput.n349 CSoutput.t140 2.82907
R22540 CSoutput.n408 CSoutput.t155 2.82907
R22541 CSoutput.n408 CSoutput.t199 2.82907
R22542 CSoutput.n409 CSoutput.t137 2.82907
R22543 CSoutput.n409 CSoutput.t179 2.82907
R22544 CSoutput.n411 CSoutput.t144 2.82907
R22545 CSoutput.n411 CSoutput.t3 2.82907
R22546 CSoutput.n413 CSoutput.t163 2.82907
R22547 CSoutput.n413 CSoutput.t197 2.82907
R22548 CSoutput.n415 CSoutput.t141 2.82907
R22549 CSoutput.n415 CSoutput.t156 2.82907
R22550 CSoutput.n417 CSoutput.t148 2.82907
R22551 CSoutput.n417 CSoutput.t143 2.82907
R22552 CSoutput.n419 CSoutput.t146 2.82907
R22553 CSoutput.n419 CSoutput.t169 2.82907
R22554 CSoutput.n421 CSoutput.t162 2.82907
R22555 CSoutput.n421 CSoutput.t183 2.82907
R22556 CSoutput.n423 CSoutput.t128 2.82907
R22557 CSoutput.n423 CSoutput.t173 2.82907
R22558 CSoutput.n425 CSoutput.t189 2.82907
R22559 CSoutput.n425 CSoutput.t182 2.82907
R22560 CSoutput.n389 CSoutput.t142 2.82907
R22561 CSoutput.n389 CSoutput.t174 2.82907
R22562 CSoutput.n390 CSoutput.t129 2.82907
R22563 CSoutput.n390 CSoutput.t176 2.82907
R22564 CSoutput.n392 CSoutput.t196 2.82907
R22565 CSoutput.n392 CSoutput.t153 2.82907
R22566 CSoutput.n394 CSoutput.t136 2.82907
R22567 CSoutput.n394 CSoutput.t167 2.82907
R22568 CSoutput.n396 CSoutput.t177 2.82907
R22569 CSoutput.n396 CSoutput.t126 2.82907
R22570 CSoutput.n398 CSoutput.t145 2.82907
R22571 CSoutput.n398 CSoutput.t4 2.82907
R22572 CSoutput.n400 CSoutput.t178 2.82907
R22573 CSoutput.n400 CSoutput.t147 2.82907
R22574 CSoutput.n402 CSoutput.t132 2.82907
R22575 CSoutput.n402 CSoutput.t187 2.82907
R22576 CSoutput.n404 CSoutput.t131 2.82907
R22577 CSoutput.n404 CSoutput.t135 2.82907
R22578 CSoutput.n406 CSoutput.t175 2.82907
R22579 CSoutput.n406 CSoutput.t191 2.82907
R22580 CSoutput.n348 CSoutput.n138 2.57547
R22581 CSoutput.n75 CSoutput.n1 2.45513
R22582 CSoutput.n229 CSoutput.n227 2.251
R22583 CSoutput.n229 CSoutput.n226 2.251
R22584 CSoutput.n229 CSoutput.n225 2.251
R22585 CSoutput.n229 CSoutput.n224 2.251
R22586 CSoutput.n198 CSoutput.n197 2.251
R22587 CSoutput.n198 CSoutput.n196 2.251
R22588 CSoutput.n198 CSoutput.n195 2.251
R22589 CSoutput.n198 CSoutput.n194 2.251
R22590 CSoutput.n271 CSoutput.n270 2.251
R22591 CSoutput.n236 CSoutput.n234 2.251
R22592 CSoutput.n236 CSoutput.n233 2.251
R22593 CSoutput.n236 CSoutput.n232 2.251
R22594 CSoutput.n254 CSoutput.n236 2.251
R22595 CSoutput.n242 CSoutput.n241 2.251
R22596 CSoutput.n242 CSoutput.n240 2.251
R22597 CSoutput.n242 CSoutput.n239 2.251
R22598 CSoutput.n242 CSoutput.n238 2.251
R22599 CSoutput.n268 CSoutput.n208 2.251
R22600 CSoutput.n263 CSoutput.n261 2.251
R22601 CSoutput.n263 CSoutput.n260 2.251
R22602 CSoutput.n263 CSoutput.n259 2.251
R22603 CSoutput.n263 CSoutput.n258 2.251
R22604 CSoutput.n164 CSoutput.n163 2.251
R22605 CSoutput.n164 CSoutput.n162 2.251
R22606 CSoutput.n164 CSoutput.n161 2.251
R22607 CSoutput.n164 CSoutput.n160 2.251
R22608 CSoutput.n281 CSoutput.n280 2.251
R22609 CSoutput.n198 CSoutput.n178 2.2505
R22610 CSoutput.n193 CSoutput.n178 2.2505
R22611 CSoutput.n191 CSoutput.n178 2.2505
R22612 CSoutput.n190 CSoutput.n178 2.2505
R22613 CSoutput.n275 CSoutput.n178 2.2505
R22614 CSoutput.n273 CSoutput.n178 2.2505
R22615 CSoutput.n271 CSoutput.n178 2.2505
R22616 CSoutput.n201 CSoutput.n178 2.2505
R22617 CSoutput.n200 CSoutput.n178 2.2505
R22618 CSoutput.n204 CSoutput.n178 2.2505
R22619 CSoutput.n203 CSoutput.n178 2.2505
R22620 CSoutput.n186 CSoutput.n178 2.2505
R22621 CSoutput.n278 CSoutput.n178 2.2505
R22622 CSoutput.n278 CSoutput.n277 2.2505
R22623 CSoutput.n242 CSoutput.n213 2.2505
R22624 CSoutput.n223 CSoutput.n213 2.2505
R22625 CSoutput.n244 CSoutput.n213 2.2505
R22626 CSoutput.n222 CSoutput.n213 2.2505
R22627 CSoutput.n246 CSoutput.n213 2.2505
R22628 CSoutput.n213 CSoutput.n207 2.2505
R22629 CSoutput.n268 CSoutput.n213 2.2505
R22630 CSoutput.n266 CSoutput.n213 2.2505
R22631 CSoutput.n248 CSoutput.n213 2.2505
R22632 CSoutput.n220 CSoutput.n213 2.2505
R22633 CSoutput.n250 CSoutput.n213 2.2505
R22634 CSoutput.n219 CSoutput.n213 2.2505
R22635 CSoutput.n264 CSoutput.n213 2.2505
R22636 CSoutput.n264 CSoutput.n217 2.2505
R22637 CSoutput.n164 CSoutput.n144 2.2505
R22638 CSoutput.n159 CSoutput.n144 2.2505
R22639 CSoutput.n157 CSoutput.n144 2.2505
R22640 CSoutput.n156 CSoutput.n144 2.2505
R22641 CSoutput.n285 CSoutput.n144 2.2505
R22642 CSoutput.n283 CSoutput.n144 2.2505
R22643 CSoutput.n281 CSoutput.n144 2.2505
R22644 CSoutput.n167 CSoutput.n144 2.2505
R22645 CSoutput.n166 CSoutput.n144 2.2505
R22646 CSoutput.n170 CSoutput.n144 2.2505
R22647 CSoutput.n169 CSoutput.n144 2.2505
R22648 CSoutput.n152 CSoutput.n144 2.2505
R22649 CSoutput.n288 CSoutput.n144 2.2505
R22650 CSoutput.n288 CSoutput.n287 2.2505
R22651 CSoutput.n206 CSoutput.n199 2.25024
R22652 CSoutput.n206 CSoutput.n192 2.25024
R22653 CSoutput.n274 CSoutput.n206 2.25024
R22654 CSoutput.n206 CSoutput.n202 2.25024
R22655 CSoutput.n206 CSoutput.n205 2.25024
R22656 CSoutput.n206 CSoutput.n173 2.25024
R22657 CSoutput.n256 CSoutput.n253 2.25024
R22658 CSoutput.n256 CSoutput.n252 2.25024
R22659 CSoutput.n256 CSoutput.n251 2.25024
R22660 CSoutput.n256 CSoutput.n218 2.25024
R22661 CSoutput.n256 CSoutput.n255 2.25024
R22662 CSoutput.n257 CSoutput.n256 2.25024
R22663 CSoutput.n172 CSoutput.n165 2.25024
R22664 CSoutput.n172 CSoutput.n158 2.25024
R22665 CSoutput.n284 CSoutput.n172 2.25024
R22666 CSoutput.n172 CSoutput.n168 2.25024
R22667 CSoutput.n172 CSoutput.n171 2.25024
R22668 CSoutput.n172 CSoutput.n139 2.25024
R22669 CSoutput.n273 CSoutput.n183 1.50111
R22670 CSoutput.n221 CSoutput.n207 1.50111
R22671 CSoutput.n283 CSoutput.n149 1.50111
R22672 CSoutput.n229 CSoutput.n228 1.501
R22673 CSoutput.n236 CSoutput.n235 1.501
R22674 CSoutput.n263 CSoutput.n262 1.501
R22675 CSoutput.n277 CSoutput.n188 1.12536
R22676 CSoutput.n277 CSoutput.n189 1.12536
R22677 CSoutput.n277 CSoutput.n276 1.12536
R22678 CSoutput.n237 CSoutput.n217 1.12536
R22679 CSoutput.n243 CSoutput.n217 1.12536
R22680 CSoutput.n245 CSoutput.n217 1.12536
R22681 CSoutput.n287 CSoutput.n154 1.12536
R22682 CSoutput.n287 CSoutput.n155 1.12536
R22683 CSoutput.n287 CSoutput.n286 1.12536
R22684 CSoutput.n277 CSoutput.n184 1.12536
R22685 CSoutput.n277 CSoutput.n185 1.12536
R22686 CSoutput.n277 CSoutput.n187 1.12536
R22687 CSoutput.n267 CSoutput.n217 1.12536
R22688 CSoutput.n247 CSoutput.n217 1.12536
R22689 CSoutput.n249 CSoutput.n217 1.12536
R22690 CSoutput.n287 CSoutput.n150 1.12536
R22691 CSoutput.n287 CSoutput.n151 1.12536
R22692 CSoutput.n287 CSoutput.n153 1.12536
R22693 CSoutput.n31 CSoutput.n30 0.669944
R22694 CSoutput.n62 CSoutput.n61 0.669944
R22695 CSoutput.n372 CSoutput.n370 0.573776
R22696 CSoutput.n374 CSoutput.n372 0.573776
R22697 CSoutput.n376 CSoutput.n374 0.573776
R22698 CSoutput.n378 CSoutput.n376 0.573776
R22699 CSoutput.n380 CSoutput.n378 0.573776
R22700 CSoutput.n382 CSoutput.n380 0.573776
R22701 CSoutput.n384 CSoutput.n382 0.573776
R22702 CSoutput.n386 CSoutput.n384 0.573776
R22703 CSoutput.n353 CSoutput.n351 0.573776
R22704 CSoutput.n355 CSoutput.n353 0.573776
R22705 CSoutput.n357 CSoutput.n355 0.573776
R22706 CSoutput.n359 CSoutput.n357 0.573776
R22707 CSoutput.n361 CSoutput.n359 0.573776
R22708 CSoutput.n363 CSoutput.n361 0.573776
R22709 CSoutput.n365 CSoutput.n363 0.573776
R22710 CSoutput.n367 CSoutput.n365 0.573776
R22711 CSoutput.n426 CSoutput.n424 0.573776
R22712 CSoutput.n424 CSoutput.n422 0.573776
R22713 CSoutput.n422 CSoutput.n420 0.573776
R22714 CSoutput.n420 CSoutput.n418 0.573776
R22715 CSoutput.n418 CSoutput.n416 0.573776
R22716 CSoutput.n416 CSoutput.n414 0.573776
R22717 CSoutput.n414 CSoutput.n412 0.573776
R22718 CSoutput.n412 CSoutput.n410 0.573776
R22719 CSoutput.n407 CSoutput.n405 0.573776
R22720 CSoutput.n405 CSoutput.n403 0.573776
R22721 CSoutput.n403 CSoutput.n401 0.573776
R22722 CSoutput.n401 CSoutput.n399 0.573776
R22723 CSoutput.n399 CSoutput.n397 0.573776
R22724 CSoutput.n397 CSoutput.n395 0.573776
R22725 CSoutput.n395 CSoutput.n393 0.573776
R22726 CSoutput.n393 CSoutput.n391 0.573776
R22727 CSoutput.n429 CSoutput.n288 0.53442
R22728 CSoutput.n332 CSoutput.n330 0.358259
R22729 CSoutput.n334 CSoutput.n332 0.358259
R22730 CSoutput.n336 CSoutput.n334 0.358259
R22731 CSoutput.n338 CSoutput.n336 0.358259
R22732 CSoutput.n340 CSoutput.n338 0.358259
R22733 CSoutput.n342 CSoutput.n340 0.358259
R22734 CSoutput.n344 CSoutput.n342 0.358259
R22735 CSoutput.n346 CSoutput.n344 0.358259
R22736 CSoutput.n312 CSoutput.n310 0.358259
R22737 CSoutput.n314 CSoutput.n312 0.358259
R22738 CSoutput.n316 CSoutput.n314 0.358259
R22739 CSoutput.n318 CSoutput.n316 0.358259
R22740 CSoutput.n320 CSoutput.n318 0.358259
R22741 CSoutput.n322 CSoutput.n320 0.358259
R22742 CSoutput.n324 CSoutput.n322 0.358259
R22743 CSoutput.n326 CSoutput.n324 0.358259
R22744 CSoutput.n293 CSoutput.n291 0.358259
R22745 CSoutput.n295 CSoutput.n293 0.358259
R22746 CSoutput.n297 CSoutput.n295 0.358259
R22747 CSoutput.n299 CSoutput.n297 0.358259
R22748 CSoutput.n301 CSoutput.n299 0.358259
R22749 CSoutput.n303 CSoutput.n301 0.358259
R22750 CSoutput.n305 CSoutput.n303 0.358259
R22751 CSoutput.n307 CSoutput.n305 0.358259
R22752 CSoutput.n136 CSoutput.n134 0.358259
R22753 CSoutput.n134 CSoutput.n132 0.358259
R22754 CSoutput.n132 CSoutput.n130 0.358259
R22755 CSoutput.n130 CSoutput.n128 0.358259
R22756 CSoutput.n128 CSoutput.n126 0.358259
R22757 CSoutput.n126 CSoutput.n124 0.358259
R22758 CSoutput.n124 CSoutput.n122 0.358259
R22759 CSoutput.n122 CSoutput.n120 0.358259
R22760 CSoutput.n116 CSoutput.n114 0.358259
R22761 CSoutput.n114 CSoutput.n112 0.358259
R22762 CSoutput.n112 CSoutput.n110 0.358259
R22763 CSoutput.n110 CSoutput.n108 0.358259
R22764 CSoutput.n108 CSoutput.n106 0.358259
R22765 CSoutput.n106 CSoutput.n104 0.358259
R22766 CSoutput.n104 CSoutput.n102 0.358259
R22767 CSoutput.n102 CSoutput.n100 0.358259
R22768 CSoutput.n97 CSoutput.n95 0.358259
R22769 CSoutput.n95 CSoutput.n93 0.358259
R22770 CSoutput.n93 CSoutput.n91 0.358259
R22771 CSoutput.n91 CSoutput.n89 0.358259
R22772 CSoutput.n89 CSoutput.n87 0.358259
R22773 CSoutput.n87 CSoutput.n85 0.358259
R22774 CSoutput.n85 CSoutput.n83 0.358259
R22775 CSoutput.n83 CSoutput.n81 0.358259
R22776 CSoutput.n21 CSoutput.n20 0.169105
R22777 CSoutput.n21 CSoutput.n16 0.169105
R22778 CSoutput.n26 CSoutput.n16 0.169105
R22779 CSoutput.n27 CSoutput.n26 0.169105
R22780 CSoutput.n27 CSoutput.n14 0.169105
R22781 CSoutput.n32 CSoutput.n14 0.169105
R22782 CSoutput.n33 CSoutput.n32 0.169105
R22783 CSoutput.n34 CSoutput.n33 0.169105
R22784 CSoutput.n34 CSoutput.n12 0.169105
R22785 CSoutput.n39 CSoutput.n12 0.169105
R22786 CSoutput.n40 CSoutput.n39 0.169105
R22787 CSoutput.n40 CSoutput.n10 0.169105
R22788 CSoutput.n45 CSoutput.n10 0.169105
R22789 CSoutput.n46 CSoutput.n45 0.169105
R22790 CSoutput.n47 CSoutput.n46 0.169105
R22791 CSoutput.n47 CSoutput.n8 0.169105
R22792 CSoutput.n52 CSoutput.n8 0.169105
R22793 CSoutput.n53 CSoutput.n52 0.169105
R22794 CSoutput.n53 CSoutput.n6 0.169105
R22795 CSoutput.n58 CSoutput.n6 0.169105
R22796 CSoutput.n59 CSoutput.n58 0.169105
R22797 CSoutput.n60 CSoutput.n59 0.169105
R22798 CSoutput.n60 CSoutput.n4 0.169105
R22799 CSoutput.n66 CSoutput.n4 0.169105
R22800 CSoutput.n67 CSoutput.n66 0.169105
R22801 CSoutput.n68 CSoutput.n67 0.169105
R22802 CSoutput.n68 CSoutput.n2 0.169105
R22803 CSoutput.n73 CSoutput.n2 0.169105
R22804 CSoutput.n74 CSoutput.n73 0.169105
R22805 CSoutput.n74 CSoutput.n0 0.169105
R22806 CSoutput.n78 CSoutput.n0 0.169105
R22807 CSoutput.n231 CSoutput.n230 0.0910737
R22808 CSoutput.n282 CSoutput.n279 0.0723685
R22809 CSoutput.n236 CSoutput.n231 0.0522944
R22810 CSoutput.n279 CSoutput.n278 0.0499135
R22811 CSoutput.n230 CSoutput.n229 0.0499135
R22812 CSoutput.n264 CSoutput.n263 0.0464294
R22813 CSoutput.n272 CSoutput.n269 0.0391444
R22814 CSoutput.n231 CSoutput.t217 0.023435
R22815 CSoutput.n279 CSoutput.t205 0.02262
R22816 CSoutput.n230 CSoutput.t213 0.02262
R22817 CSoutput CSoutput.n429 0.0052
R22818 CSoutput.n201 CSoutput.n184 0.00365111
R22819 CSoutput.n204 CSoutput.n185 0.00365111
R22820 CSoutput.n187 CSoutput.n186 0.00365111
R22821 CSoutput.n229 CSoutput.n188 0.00365111
R22822 CSoutput.n193 CSoutput.n189 0.00365111
R22823 CSoutput.n276 CSoutput.n190 0.00365111
R22824 CSoutput.n267 CSoutput.n266 0.00365111
R22825 CSoutput.n247 CSoutput.n220 0.00365111
R22826 CSoutput.n249 CSoutput.n219 0.00365111
R22827 CSoutput.n237 CSoutput.n236 0.00365111
R22828 CSoutput.n243 CSoutput.n223 0.00365111
R22829 CSoutput.n245 CSoutput.n222 0.00365111
R22830 CSoutput.n167 CSoutput.n150 0.00365111
R22831 CSoutput.n170 CSoutput.n151 0.00365111
R22832 CSoutput.n153 CSoutput.n152 0.00365111
R22833 CSoutput.n263 CSoutput.n154 0.00365111
R22834 CSoutput.n159 CSoutput.n155 0.00365111
R22835 CSoutput.n286 CSoutput.n156 0.00365111
R22836 CSoutput.n198 CSoutput.n188 0.00340054
R22837 CSoutput.n191 CSoutput.n189 0.00340054
R22838 CSoutput.n276 CSoutput.n275 0.00340054
R22839 CSoutput.n271 CSoutput.n184 0.00340054
R22840 CSoutput.n200 CSoutput.n185 0.00340054
R22841 CSoutput.n203 CSoutput.n187 0.00340054
R22842 CSoutput.n242 CSoutput.n237 0.00340054
R22843 CSoutput.n244 CSoutput.n243 0.00340054
R22844 CSoutput.n246 CSoutput.n245 0.00340054
R22845 CSoutput.n268 CSoutput.n267 0.00340054
R22846 CSoutput.n248 CSoutput.n247 0.00340054
R22847 CSoutput.n250 CSoutput.n249 0.00340054
R22848 CSoutput.n164 CSoutput.n154 0.00340054
R22849 CSoutput.n157 CSoutput.n155 0.00340054
R22850 CSoutput.n286 CSoutput.n285 0.00340054
R22851 CSoutput.n281 CSoutput.n150 0.00340054
R22852 CSoutput.n166 CSoutput.n151 0.00340054
R22853 CSoutput.n169 CSoutput.n153 0.00340054
R22854 CSoutput.n199 CSoutput.n193 0.00252698
R22855 CSoutput.n192 CSoutput.n190 0.00252698
R22856 CSoutput.n274 CSoutput.n273 0.00252698
R22857 CSoutput.n202 CSoutput.n200 0.00252698
R22858 CSoutput.n205 CSoutput.n203 0.00252698
R22859 CSoutput.n278 CSoutput.n173 0.00252698
R22860 CSoutput.n199 CSoutput.n198 0.00252698
R22861 CSoutput.n192 CSoutput.n191 0.00252698
R22862 CSoutput.n275 CSoutput.n274 0.00252698
R22863 CSoutput.n202 CSoutput.n201 0.00252698
R22864 CSoutput.n205 CSoutput.n204 0.00252698
R22865 CSoutput.n186 CSoutput.n173 0.00252698
R22866 CSoutput.n253 CSoutput.n223 0.00252698
R22867 CSoutput.n252 CSoutput.n222 0.00252698
R22868 CSoutput.n251 CSoutput.n207 0.00252698
R22869 CSoutput.n248 CSoutput.n218 0.00252698
R22870 CSoutput.n255 CSoutput.n250 0.00252698
R22871 CSoutput.n264 CSoutput.n257 0.00252698
R22872 CSoutput.n253 CSoutput.n242 0.00252698
R22873 CSoutput.n252 CSoutput.n244 0.00252698
R22874 CSoutput.n251 CSoutput.n246 0.00252698
R22875 CSoutput.n266 CSoutput.n218 0.00252698
R22876 CSoutput.n255 CSoutput.n220 0.00252698
R22877 CSoutput.n257 CSoutput.n219 0.00252698
R22878 CSoutput.n165 CSoutput.n159 0.00252698
R22879 CSoutput.n158 CSoutput.n156 0.00252698
R22880 CSoutput.n284 CSoutput.n283 0.00252698
R22881 CSoutput.n168 CSoutput.n166 0.00252698
R22882 CSoutput.n171 CSoutput.n169 0.00252698
R22883 CSoutput.n288 CSoutput.n139 0.00252698
R22884 CSoutput.n165 CSoutput.n164 0.00252698
R22885 CSoutput.n158 CSoutput.n157 0.00252698
R22886 CSoutput.n285 CSoutput.n284 0.00252698
R22887 CSoutput.n168 CSoutput.n167 0.00252698
R22888 CSoutput.n171 CSoutput.n170 0.00252698
R22889 CSoutput.n152 CSoutput.n139 0.00252698
R22890 CSoutput.n273 CSoutput.n272 0.0020275
R22891 CSoutput.n272 CSoutput.n271 0.0020275
R22892 CSoutput.n269 CSoutput.n207 0.0020275
R22893 CSoutput.n269 CSoutput.n268 0.0020275
R22894 CSoutput.n283 CSoutput.n282 0.0020275
R22895 CSoutput.n282 CSoutput.n281 0.0020275
R22896 CSoutput.n183 CSoutput.n182 0.00166668
R22897 CSoutput.n265 CSoutput.n221 0.00166668
R22898 CSoutput.n149 CSoutput.n148 0.00166668
R22899 CSoutput.n287 CSoutput.n149 0.00133328
R22900 CSoutput.n221 CSoutput.n217 0.00133328
R22901 CSoutput.n277 CSoutput.n183 0.00133328
R22902 CSoutput.n280 CSoutput.n172 0.001
R22903 CSoutput.n258 CSoutput.n172 0.001
R22904 CSoutput.n160 CSoutput.n140 0.001
R22905 CSoutput.n259 CSoutput.n140 0.001
R22906 CSoutput.n161 CSoutput.n141 0.001
R22907 CSoutput.n260 CSoutput.n141 0.001
R22908 CSoutput.n162 CSoutput.n142 0.001
R22909 CSoutput.n261 CSoutput.n142 0.001
R22910 CSoutput.n163 CSoutput.n143 0.001
R22911 CSoutput.n262 CSoutput.n143 0.001
R22912 CSoutput.n256 CSoutput.n208 0.001
R22913 CSoutput.n256 CSoutput.n254 0.001
R22914 CSoutput.n238 CSoutput.n209 0.001
R22915 CSoutput.n232 CSoutput.n209 0.001
R22916 CSoutput.n239 CSoutput.n210 0.001
R22917 CSoutput.n233 CSoutput.n210 0.001
R22918 CSoutput.n240 CSoutput.n211 0.001
R22919 CSoutput.n234 CSoutput.n211 0.001
R22920 CSoutput.n241 CSoutput.n212 0.001
R22921 CSoutput.n235 CSoutput.n212 0.001
R22922 CSoutput.n270 CSoutput.n206 0.001
R22923 CSoutput.n224 CSoutput.n206 0.001
R22924 CSoutput.n194 CSoutput.n174 0.001
R22925 CSoutput.n225 CSoutput.n174 0.001
R22926 CSoutput.n195 CSoutput.n175 0.001
R22927 CSoutput.n226 CSoutput.n175 0.001
R22928 CSoutput.n196 CSoutput.n176 0.001
R22929 CSoutput.n227 CSoutput.n176 0.001
R22930 CSoutput.n197 CSoutput.n177 0.001
R22931 CSoutput.n228 CSoutput.n177 0.001
R22932 CSoutput.n228 CSoutput.n178 0.001
R22933 CSoutput.n227 CSoutput.n179 0.001
R22934 CSoutput.n226 CSoutput.n180 0.001
R22935 CSoutput.n225 CSoutput.t207 0.001
R22936 CSoutput.n224 CSoutput.n181 0.001
R22937 CSoutput.n197 CSoutput.n179 0.001
R22938 CSoutput.n196 CSoutput.n180 0.001
R22939 CSoutput.n195 CSoutput.t207 0.001
R22940 CSoutput.n194 CSoutput.n181 0.001
R22941 CSoutput.n270 CSoutput.n182 0.001
R22942 CSoutput.n235 CSoutput.n213 0.001
R22943 CSoutput.n234 CSoutput.n214 0.001
R22944 CSoutput.n233 CSoutput.n215 0.001
R22945 CSoutput.n232 CSoutput.t208 0.001
R22946 CSoutput.n254 CSoutput.n216 0.001
R22947 CSoutput.n241 CSoutput.n214 0.001
R22948 CSoutput.n240 CSoutput.n215 0.001
R22949 CSoutput.n239 CSoutput.t208 0.001
R22950 CSoutput.n238 CSoutput.n216 0.001
R22951 CSoutput.n265 CSoutput.n208 0.001
R22952 CSoutput.n262 CSoutput.n144 0.001
R22953 CSoutput.n261 CSoutput.n145 0.001
R22954 CSoutput.n260 CSoutput.n146 0.001
R22955 CSoutput.n259 CSoutput.t210 0.001
R22956 CSoutput.n258 CSoutput.n147 0.001
R22957 CSoutput.n163 CSoutput.n145 0.001
R22958 CSoutput.n162 CSoutput.n146 0.001
R22959 CSoutput.n161 CSoutput.t210 0.001
R22960 CSoutput.n160 CSoutput.n147 0.001
R22961 CSoutput.n280 CSoutput.n148 0.001
R22962 diffpairibias.n0 diffpairibias.t27 436.822
R22963 diffpairibias.n27 diffpairibias.t24 435.479
R22964 diffpairibias.n26 diffpairibias.t21 435.479
R22965 diffpairibias.n25 diffpairibias.t22 435.479
R22966 diffpairibias.n24 diffpairibias.t26 435.479
R22967 diffpairibias.n23 diffpairibias.t20 435.479
R22968 diffpairibias.n0 diffpairibias.t23 435.479
R22969 diffpairibias.n1 diffpairibias.t28 435.479
R22970 diffpairibias.n2 diffpairibias.t25 435.479
R22971 diffpairibias.n3 diffpairibias.t29 435.479
R22972 diffpairibias.n13 diffpairibias.t14 377.536
R22973 diffpairibias.n13 diffpairibias.t0 376.193
R22974 diffpairibias.n14 diffpairibias.t10 376.193
R22975 diffpairibias.n15 diffpairibias.t12 376.193
R22976 diffpairibias.n16 diffpairibias.t6 376.193
R22977 diffpairibias.n17 diffpairibias.t2 376.193
R22978 diffpairibias.n18 diffpairibias.t16 376.193
R22979 diffpairibias.n19 diffpairibias.t4 376.193
R22980 diffpairibias.n20 diffpairibias.t18 376.193
R22981 diffpairibias.n21 diffpairibias.t8 376.193
R22982 diffpairibias.n4 diffpairibias.t15 113.368
R22983 diffpairibias.n4 diffpairibias.t1 112.698
R22984 diffpairibias.n5 diffpairibias.t11 112.698
R22985 diffpairibias.n6 diffpairibias.t13 112.698
R22986 diffpairibias.n7 diffpairibias.t7 112.698
R22987 diffpairibias.n8 diffpairibias.t3 112.698
R22988 diffpairibias.n9 diffpairibias.t17 112.698
R22989 diffpairibias.n10 diffpairibias.t5 112.698
R22990 diffpairibias.n11 diffpairibias.t19 112.698
R22991 diffpairibias.n12 diffpairibias.t9 112.698
R22992 diffpairibias.n22 diffpairibias.n21 4.77242
R22993 diffpairibias.n22 diffpairibias.n12 4.30807
R22994 diffpairibias.n23 diffpairibias.n22 4.13945
R22995 diffpairibias.n21 diffpairibias.n20 1.34352
R22996 diffpairibias.n20 diffpairibias.n19 1.34352
R22997 diffpairibias.n19 diffpairibias.n18 1.34352
R22998 diffpairibias.n18 diffpairibias.n17 1.34352
R22999 diffpairibias.n17 diffpairibias.n16 1.34352
R23000 diffpairibias.n16 diffpairibias.n15 1.34352
R23001 diffpairibias.n15 diffpairibias.n14 1.34352
R23002 diffpairibias.n14 diffpairibias.n13 1.34352
R23003 diffpairibias.n3 diffpairibias.n2 1.34352
R23004 diffpairibias.n2 diffpairibias.n1 1.34352
R23005 diffpairibias.n1 diffpairibias.n0 1.34352
R23006 diffpairibias.n24 diffpairibias.n23 1.34352
R23007 diffpairibias.n25 diffpairibias.n24 1.34352
R23008 diffpairibias.n26 diffpairibias.n25 1.34352
R23009 diffpairibias.n27 diffpairibias.n26 1.34352
R23010 diffpairibias.n28 diffpairibias.n27 0.862419
R23011 diffpairibias diffpairibias.n28 0.684875
R23012 diffpairibias.n12 diffpairibias.n11 0.672012
R23013 diffpairibias.n11 diffpairibias.n10 0.672012
R23014 diffpairibias.n10 diffpairibias.n9 0.672012
R23015 diffpairibias.n9 diffpairibias.n8 0.672012
R23016 diffpairibias.n8 diffpairibias.n7 0.672012
R23017 diffpairibias.n7 diffpairibias.n6 0.672012
R23018 diffpairibias.n6 diffpairibias.n5 0.672012
R23019 diffpairibias.n5 diffpairibias.n4 0.672012
R23020 diffpairibias.n28 diffpairibias.n3 0.190907
R23021 commonsourceibias.n281 commonsourceibias.t101 222.032
R23022 commonsourceibias.n44 commonsourceibias.t78 222.032
R23023 commonsourceibias.n166 commonsourceibias.t117 222.032
R23024 commonsourceibias.n643 commonsourceibias.t106 222.032
R23025 commonsourceibias.n413 commonsourceibias.t28 222.032
R23026 commonsourceibias.n529 commonsourceibias.t123 222.032
R23027 commonsourceibias.n364 commonsourceibias.t100 207.983
R23028 commonsourceibias.n127 commonsourceibias.t74 207.983
R23029 commonsourceibias.n249 commonsourceibias.t115 207.983
R23030 commonsourceibias.n731 commonsourceibias.t122 207.983
R23031 commonsourceibias.n501 commonsourceibias.t14 207.983
R23032 commonsourceibias.n616 commonsourceibias.t140 207.983
R23033 commonsourceibias.n280 commonsourceibias.t87 168.701
R23034 commonsourceibias.n286 commonsourceibias.t129 168.701
R23035 commonsourceibias.n292 commonsourceibias.t110 168.701
R23036 commonsourceibias.n276 commonsourceibias.t93 168.701
R23037 commonsourceibias.n300 commonsourceibias.t95 168.701
R23038 commonsourceibias.n306 commonsourceibias.t121 168.701
R23039 commonsourceibias.n271 commonsourceibias.t102 168.701
R23040 commonsourceibias.n314 commonsourceibias.t108 168.701
R23041 commonsourceibias.n320 commonsourceibias.t159 168.701
R23042 commonsourceibias.n266 commonsourceibias.t138 168.701
R23043 commonsourceibias.n328 commonsourceibias.t118 168.701
R23044 commonsourceibias.n334 commonsourceibias.t83 168.701
R23045 commonsourceibias.n261 commonsourceibias.t86 168.701
R23046 commonsourceibias.n342 commonsourceibias.t128 168.701
R23047 commonsourceibias.n348 commonsourceibias.t109 168.701
R23048 commonsourceibias.n256 commonsourceibias.t92 168.701
R23049 commonsourceibias.n356 commonsourceibias.t137 168.701
R23050 commonsourceibias.n362 commonsourceibias.t119 168.701
R23051 commonsourceibias.n125 commonsourceibias.t20 168.701
R23052 commonsourceibias.n119 commonsourceibias.t50 168.701
R23053 commonsourceibias.n19 commonsourceibias.t8 168.701
R23054 commonsourceibias.n111 commonsourceibias.t36 168.701
R23055 commonsourceibias.n105 commonsourceibias.t76 168.701
R23056 commonsourceibias.n24 commonsourceibias.t24 168.701
R23057 commonsourceibias.n97 commonsourceibias.t34 168.701
R23058 commonsourceibias.n91 commonsourceibias.t10 168.701
R23059 commonsourceibias.n29 commonsourceibias.t40 168.701
R23060 commonsourceibias.n83 commonsourceibias.t56 168.701
R23061 commonsourceibias.n77 commonsourceibias.t26 168.701
R23062 commonsourceibias.n34 commonsourceibias.t38 168.701
R23063 commonsourceibias.n69 commonsourceibias.t70 168.701
R23064 commonsourceibias.n63 commonsourceibias.t18 168.701
R23065 commonsourceibias.n39 commonsourceibias.t22 168.701
R23066 commonsourceibias.n55 commonsourceibias.t54 168.701
R23067 commonsourceibias.n49 commonsourceibias.t4 168.701
R23068 commonsourceibias.n43 commonsourceibias.t46 168.701
R23069 commonsourceibias.n247 commonsourceibias.t136 168.701
R23070 commonsourceibias.n241 commonsourceibias.t151 168.701
R23071 commonsourceibias.n5 commonsourceibias.t105 168.701
R23072 commonsourceibias.n233 commonsourceibias.t126 168.701
R23073 commonsourceibias.n227 commonsourceibias.t144 168.701
R23074 commonsourceibias.n10 commonsourceibias.t98 168.701
R23075 commonsourceibias.n219 commonsourceibias.t94 168.701
R23076 commonsourceibias.n213 commonsourceibias.t135 168.701
R23077 commonsourceibias.n150 commonsourceibias.t153 168.701
R23078 commonsourceibias.n151 commonsourceibias.t88 168.701
R23079 commonsourceibias.n153 commonsourceibias.t125 168.701
R23080 commonsourceibias.n155 commonsourceibias.t120 168.701
R23081 commonsourceibias.n191 commonsourceibias.t139 168.701
R23082 commonsourceibias.n185 commonsourceibias.t112 168.701
R23083 commonsourceibias.n161 commonsourceibias.t107 168.701
R23084 commonsourceibias.n177 commonsourceibias.t127 168.701
R23085 commonsourceibias.n171 commonsourceibias.t146 168.701
R23086 commonsourceibias.n165 commonsourceibias.t99 168.701
R23087 commonsourceibias.n642 commonsourceibias.t90 168.701
R23088 commonsourceibias.n648 commonsourceibias.t134 168.701
R23089 commonsourceibias.n654 commonsourceibias.t116 168.701
R23090 commonsourceibias.n656 commonsourceibias.t96 168.701
R23091 commonsourceibias.n663 commonsourceibias.t91 168.701
R23092 commonsourceibias.n669 commonsourceibias.t145 168.701
R23093 commonsourceibias.n671 commonsourceibias.t124 168.701
R23094 commonsourceibias.n678 commonsourceibias.t131 168.701
R23095 commonsourceibias.n684 commonsourceibias.t152 168.701
R23096 commonsourceibias.n686 commonsourceibias.t157 168.701
R23097 commonsourceibias.n693 commonsourceibias.t141 168.701
R23098 commonsourceibias.n699 commonsourceibias.t97 168.701
R23099 commonsourceibias.n701 commonsourceibias.t81 168.701
R23100 commonsourceibias.n708 commonsourceibias.t149 168.701
R23101 commonsourceibias.n714 commonsourceibias.t132 168.701
R23102 commonsourceibias.n716 commonsourceibias.t111 168.701
R23103 commonsourceibias.n723 commonsourceibias.t156 168.701
R23104 commonsourceibias.n729 commonsourceibias.t142 168.701
R23105 commonsourceibias.n412 commonsourceibias.t2 168.701
R23106 commonsourceibias.n418 commonsourceibias.t48 168.701
R23107 commonsourceibias.n424 commonsourceibias.t12 168.701
R23108 commonsourceibias.n426 commonsourceibias.t68 168.701
R23109 commonsourceibias.n433 commonsourceibias.t66 168.701
R23110 commonsourceibias.n439 commonsourceibias.t6 168.701
R23111 commonsourceibias.n441 commonsourceibias.t62 168.701
R23112 commonsourceibias.n448 commonsourceibias.t52 168.701
R23113 commonsourceibias.n454 commonsourceibias.t72 168.701
R23114 commonsourceibias.n456 commonsourceibias.t64 168.701
R23115 commonsourceibias.n463 commonsourceibias.t32 168.701
R23116 commonsourceibias.n469 commonsourceibias.t58 168.701
R23117 commonsourceibias.n471 commonsourceibias.t44 168.701
R23118 commonsourceibias.n478 commonsourceibias.t16 168.701
R23119 commonsourceibias.n484 commonsourceibias.t60 168.701
R23120 commonsourceibias.n486 commonsourceibias.t30 168.701
R23121 commonsourceibias.n493 commonsourceibias.t0 168.701
R23122 commonsourceibias.n499 commonsourceibias.t42 168.701
R23123 commonsourceibias.n614 commonsourceibias.t155 168.701
R23124 commonsourceibias.n608 commonsourceibias.t84 168.701
R23125 commonsourceibias.n601 commonsourceibias.t130 168.701
R23126 commonsourceibias.n599 commonsourceibias.t148 168.701
R23127 commonsourceibias.n593 commonsourceibias.t80 168.701
R23128 commonsourceibias.n586 commonsourceibias.t89 168.701
R23129 commonsourceibias.n584 commonsourceibias.t113 168.701
R23130 commonsourceibias.n578 commonsourceibias.t154 168.701
R23131 commonsourceibias.n571 commonsourceibias.t85 168.701
R23132 commonsourceibias.n528 commonsourceibias.t103 168.701
R23133 commonsourceibias.n534 commonsourceibias.t150 168.701
R23134 commonsourceibias.n540 commonsourceibias.t133 168.701
R23135 commonsourceibias.n542 commonsourceibias.t114 168.701
R23136 commonsourceibias.n549 commonsourceibias.t104 168.701
R23137 commonsourceibias.n555 commonsourceibias.t158 168.701
R23138 commonsourceibias.n519 commonsourceibias.t143 168.701
R23139 commonsourceibias.n517 commonsourceibias.t147 168.701
R23140 commonsourceibias.n515 commonsourceibias.t82 168.701
R23141 commonsourceibias.n363 commonsourceibias.n251 161.3
R23142 commonsourceibias.n361 commonsourceibias.n360 161.3
R23143 commonsourceibias.n359 commonsourceibias.n252 161.3
R23144 commonsourceibias.n358 commonsourceibias.n357 161.3
R23145 commonsourceibias.n355 commonsourceibias.n253 161.3
R23146 commonsourceibias.n354 commonsourceibias.n353 161.3
R23147 commonsourceibias.n352 commonsourceibias.n254 161.3
R23148 commonsourceibias.n351 commonsourceibias.n350 161.3
R23149 commonsourceibias.n349 commonsourceibias.n255 161.3
R23150 commonsourceibias.n347 commonsourceibias.n346 161.3
R23151 commonsourceibias.n345 commonsourceibias.n257 161.3
R23152 commonsourceibias.n344 commonsourceibias.n343 161.3
R23153 commonsourceibias.n341 commonsourceibias.n258 161.3
R23154 commonsourceibias.n340 commonsourceibias.n339 161.3
R23155 commonsourceibias.n338 commonsourceibias.n259 161.3
R23156 commonsourceibias.n337 commonsourceibias.n336 161.3
R23157 commonsourceibias.n335 commonsourceibias.n260 161.3
R23158 commonsourceibias.n333 commonsourceibias.n332 161.3
R23159 commonsourceibias.n331 commonsourceibias.n262 161.3
R23160 commonsourceibias.n330 commonsourceibias.n329 161.3
R23161 commonsourceibias.n327 commonsourceibias.n263 161.3
R23162 commonsourceibias.n326 commonsourceibias.n325 161.3
R23163 commonsourceibias.n324 commonsourceibias.n264 161.3
R23164 commonsourceibias.n323 commonsourceibias.n322 161.3
R23165 commonsourceibias.n321 commonsourceibias.n265 161.3
R23166 commonsourceibias.n319 commonsourceibias.n318 161.3
R23167 commonsourceibias.n317 commonsourceibias.n267 161.3
R23168 commonsourceibias.n316 commonsourceibias.n315 161.3
R23169 commonsourceibias.n313 commonsourceibias.n268 161.3
R23170 commonsourceibias.n312 commonsourceibias.n311 161.3
R23171 commonsourceibias.n310 commonsourceibias.n269 161.3
R23172 commonsourceibias.n309 commonsourceibias.n308 161.3
R23173 commonsourceibias.n307 commonsourceibias.n270 161.3
R23174 commonsourceibias.n305 commonsourceibias.n304 161.3
R23175 commonsourceibias.n303 commonsourceibias.n272 161.3
R23176 commonsourceibias.n302 commonsourceibias.n301 161.3
R23177 commonsourceibias.n299 commonsourceibias.n273 161.3
R23178 commonsourceibias.n298 commonsourceibias.n297 161.3
R23179 commonsourceibias.n296 commonsourceibias.n274 161.3
R23180 commonsourceibias.n295 commonsourceibias.n294 161.3
R23181 commonsourceibias.n293 commonsourceibias.n275 161.3
R23182 commonsourceibias.n291 commonsourceibias.n290 161.3
R23183 commonsourceibias.n289 commonsourceibias.n277 161.3
R23184 commonsourceibias.n288 commonsourceibias.n287 161.3
R23185 commonsourceibias.n285 commonsourceibias.n278 161.3
R23186 commonsourceibias.n284 commonsourceibias.n283 161.3
R23187 commonsourceibias.n282 commonsourceibias.n279 161.3
R23188 commonsourceibias.n45 commonsourceibias.n42 161.3
R23189 commonsourceibias.n47 commonsourceibias.n46 161.3
R23190 commonsourceibias.n48 commonsourceibias.n41 161.3
R23191 commonsourceibias.n51 commonsourceibias.n50 161.3
R23192 commonsourceibias.n52 commonsourceibias.n40 161.3
R23193 commonsourceibias.n54 commonsourceibias.n53 161.3
R23194 commonsourceibias.n56 commonsourceibias.n38 161.3
R23195 commonsourceibias.n58 commonsourceibias.n57 161.3
R23196 commonsourceibias.n59 commonsourceibias.n37 161.3
R23197 commonsourceibias.n61 commonsourceibias.n60 161.3
R23198 commonsourceibias.n62 commonsourceibias.n36 161.3
R23199 commonsourceibias.n65 commonsourceibias.n64 161.3
R23200 commonsourceibias.n66 commonsourceibias.n35 161.3
R23201 commonsourceibias.n68 commonsourceibias.n67 161.3
R23202 commonsourceibias.n70 commonsourceibias.n33 161.3
R23203 commonsourceibias.n72 commonsourceibias.n71 161.3
R23204 commonsourceibias.n73 commonsourceibias.n32 161.3
R23205 commonsourceibias.n75 commonsourceibias.n74 161.3
R23206 commonsourceibias.n76 commonsourceibias.n31 161.3
R23207 commonsourceibias.n79 commonsourceibias.n78 161.3
R23208 commonsourceibias.n80 commonsourceibias.n30 161.3
R23209 commonsourceibias.n82 commonsourceibias.n81 161.3
R23210 commonsourceibias.n84 commonsourceibias.n28 161.3
R23211 commonsourceibias.n86 commonsourceibias.n85 161.3
R23212 commonsourceibias.n87 commonsourceibias.n27 161.3
R23213 commonsourceibias.n89 commonsourceibias.n88 161.3
R23214 commonsourceibias.n90 commonsourceibias.n26 161.3
R23215 commonsourceibias.n93 commonsourceibias.n92 161.3
R23216 commonsourceibias.n94 commonsourceibias.n25 161.3
R23217 commonsourceibias.n96 commonsourceibias.n95 161.3
R23218 commonsourceibias.n98 commonsourceibias.n23 161.3
R23219 commonsourceibias.n100 commonsourceibias.n99 161.3
R23220 commonsourceibias.n101 commonsourceibias.n22 161.3
R23221 commonsourceibias.n103 commonsourceibias.n102 161.3
R23222 commonsourceibias.n104 commonsourceibias.n21 161.3
R23223 commonsourceibias.n107 commonsourceibias.n106 161.3
R23224 commonsourceibias.n108 commonsourceibias.n20 161.3
R23225 commonsourceibias.n110 commonsourceibias.n109 161.3
R23226 commonsourceibias.n112 commonsourceibias.n18 161.3
R23227 commonsourceibias.n114 commonsourceibias.n113 161.3
R23228 commonsourceibias.n115 commonsourceibias.n17 161.3
R23229 commonsourceibias.n117 commonsourceibias.n116 161.3
R23230 commonsourceibias.n118 commonsourceibias.n16 161.3
R23231 commonsourceibias.n121 commonsourceibias.n120 161.3
R23232 commonsourceibias.n122 commonsourceibias.n15 161.3
R23233 commonsourceibias.n124 commonsourceibias.n123 161.3
R23234 commonsourceibias.n126 commonsourceibias.n14 161.3
R23235 commonsourceibias.n167 commonsourceibias.n164 161.3
R23236 commonsourceibias.n169 commonsourceibias.n168 161.3
R23237 commonsourceibias.n170 commonsourceibias.n163 161.3
R23238 commonsourceibias.n173 commonsourceibias.n172 161.3
R23239 commonsourceibias.n174 commonsourceibias.n162 161.3
R23240 commonsourceibias.n176 commonsourceibias.n175 161.3
R23241 commonsourceibias.n178 commonsourceibias.n160 161.3
R23242 commonsourceibias.n180 commonsourceibias.n179 161.3
R23243 commonsourceibias.n181 commonsourceibias.n159 161.3
R23244 commonsourceibias.n183 commonsourceibias.n182 161.3
R23245 commonsourceibias.n184 commonsourceibias.n158 161.3
R23246 commonsourceibias.n187 commonsourceibias.n186 161.3
R23247 commonsourceibias.n188 commonsourceibias.n157 161.3
R23248 commonsourceibias.n190 commonsourceibias.n189 161.3
R23249 commonsourceibias.n192 commonsourceibias.n156 161.3
R23250 commonsourceibias.n194 commonsourceibias.n193 161.3
R23251 commonsourceibias.n196 commonsourceibias.n195 161.3
R23252 commonsourceibias.n197 commonsourceibias.n154 161.3
R23253 commonsourceibias.n199 commonsourceibias.n198 161.3
R23254 commonsourceibias.n201 commonsourceibias.n200 161.3
R23255 commonsourceibias.n202 commonsourceibias.n152 161.3
R23256 commonsourceibias.n204 commonsourceibias.n203 161.3
R23257 commonsourceibias.n206 commonsourceibias.n205 161.3
R23258 commonsourceibias.n208 commonsourceibias.n207 161.3
R23259 commonsourceibias.n209 commonsourceibias.n13 161.3
R23260 commonsourceibias.n211 commonsourceibias.n210 161.3
R23261 commonsourceibias.n212 commonsourceibias.n12 161.3
R23262 commonsourceibias.n215 commonsourceibias.n214 161.3
R23263 commonsourceibias.n216 commonsourceibias.n11 161.3
R23264 commonsourceibias.n218 commonsourceibias.n217 161.3
R23265 commonsourceibias.n220 commonsourceibias.n9 161.3
R23266 commonsourceibias.n222 commonsourceibias.n221 161.3
R23267 commonsourceibias.n223 commonsourceibias.n8 161.3
R23268 commonsourceibias.n225 commonsourceibias.n224 161.3
R23269 commonsourceibias.n226 commonsourceibias.n7 161.3
R23270 commonsourceibias.n229 commonsourceibias.n228 161.3
R23271 commonsourceibias.n230 commonsourceibias.n6 161.3
R23272 commonsourceibias.n232 commonsourceibias.n231 161.3
R23273 commonsourceibias.n234 commonsourceibias.n4 161.3
R23274 commonsourceibias.n236 commonsourceibias.n235 161.3
R23275 commonsourceibias.n237 commonsourceibias.n3 161.3
R23276 commonsourceibias.n239 commonsourceibias.n238 161.3
R23277 commonsourceibias.n240 commonsourceibias.n2 161.3
R23278 commonsourceibias.n243 commonsourceibias.n242 161.3
R23279 commonsourceibias.n244 commonsourceibias.n1 161.3
R23280 commonsourceibias.n246 commonsourceibias.n245 161.3
R23281 commonsourceibias.n248 commonsourceibias.n0 161.3
R23282 commonsourceibias.n730 commonsourceibias.n618 161.3
R23283 commonsourceibias.n728 commonsourceibias.n727 161.3
R23284 commonsourceibias.n726 commonsourceibias.n619 161.3
R23285 commonsourceibias.n725 commonsourceibias.n724 161.3
R23286 commonsourceibias.n722 commonsourceibias.n620 161.3
R23287 commonsourceibias.n721 commonsourceibias.n720 161.3
R23288 commonsourceibias.n719 commonsourceibias.n621 161.3
R23289 commonsourceibias.n718 commonsourceibias.n717 161.3
R23290 commonsourceibias.n715 commonsourceibias.n622 161.3
R23291 commonsourceibias.n713 commonsourceibias.n712 161.3
R23292 commonsourceibias.n711 commonsourceibias.n623 161.3
R23293 commonsourceibias.n710 commonsourceibias.n709 161.3
R23294 commonsourceibias.n707 commonsourceibias.n624 161.3
R23295 commonsourceibias.n706 commonsourceibias.n705 161.3
R23296 commonsourceibias.n704 commonsourceibias.n625 161.3
R23297 commonsourceibias.n703 commonsourceibias.n702 161.3
R23298 commonsourceibias.n700 commonsourceibias.n626 161.3
R23299 commonsourceibias.n698 commonsourceibias.n697 161.3
R23300 commonsourceibias.n696 commonsourceibias.n627 161.3
R23301 commonsourceibias.n695 commonsourceibias.n694 161.3
R23302 commonsourceibias.n692 commonsourceibias.n628 161.3
R23303 commonsourceibias.n691 commonsourceibias.n690 161.3
R23304 commonsourceibias.n689 commonsourceibias.n629 161.3
R23305 commonsourceibias.n688 commonsourceibias.n687 161.3
R23306 commonsourceibias.n685 commonsourceibias.n630 161.3
R23307 commonsourceibias.n683 commonsourceibias.n682 161.3
R23308 commonsourceibias.n681 commonsourceibias.n631 161.3
R23309 commonsourceibias.n680 commonsourceibias.n679 161.3
R23310 commonsourceibias.n677 commonsourceibias.n632 161.3
R23311 commonsourceibias.n676 commonsourceibias.n675 161.3
R23312 commonsourceibias.n674 commonsourceibias.n633 161.3
R23313 commonsourceibias.n673 commonsourceibias.n672 161.3
R23314 commonsourceibias.n670 commonsourceibias.n634 161.3
R23315 commonsourceibias.n668 commonsourceibias.n667 161.3
R23316 commonsourceibias.n666 commonsourceibias.n635 161.3
R23317 commonsourceibias.n665 commonsourceibias.n664 161.3
R23318 commonsourceibias.n662 commonsourceibias.n636 161.3
R23319 commonsourceibias.n661 commonsourceibias.n660 161.3
R23320 commonsourceibias.n659 commonsourceibias.n637 161.3
R23321 commonsourceibias.n658 commonsourceibias.n657 161.3
R23322 commonsourceibias.n655 commonsourceibias.n638 161.3
R23323 commonsourceibias.n653 commonsourceibias.n652 161.3
R23324 commonsourceibias.n651 commonsourceibias.n639 161.3
R23325 commonsourceibias.n650 commonsourceibias.n649 161.3
R23326 commonsourceibias.n647 commonsourceibias.n640 161.3
R23327 commonsourceibias.n646 commonsourceibias.n645 161.3
R23328 commonsourceibias.n644 commonsourceibias.n641 161.3
R23329 commonsourceibias.n500 commonsourceibias.n388 161.3
R23330 commonsourceibias.n498 commonsourceibias.n497 161.3
R23331 commonsourceibias.n496 commonsourceibias.n389 161.3
R23332 commonsourceibias.n495 commonsourceibias.n494 161.3
R23333 commonsourceibias.n492 commonsourceibias.n390 161.3
R23334 commonsourceibias.n491 commonsourceibias.n490 161.3
R23335 commonsourceibias.n489 commonsourceibias.n391 161.3
R23336 commonsourceibias.n488 commonsourceibias.n487 161.3
R23337 commonsourceibias.n485 commonsourceibias.n392 161.3
R23338 commonsourceibias.n483 commonsourceibias.n482 161.3
R23339 commonsourceibias.n481 commonsourceibias.n393 161.3
R23340 commonsourceibias.n480 commonsourceibias.n479 161.3
R23341 commonsourceibias.n477 commonsourceibias.n394 161.3
R23342 commonsourceibias.n476 commonsourceibias.n475 161.3
R23343 commonsourceibias.n474 commonsourceibias.n395 161.3
R23344 commonsourceibias.n473 commonsourceibias.n472 161.3
R23345 commonsourceibias.n470 commonsourceibias.n396 161.3
R23346 commonsourceibias.n468 commonsourceibias.n467 161.3
R23347 commonsourceibias.n466 commonsourceibias.n397 161.3
R23348 commonsourceibias.n465 commonsourceibias.n464 161.3
R23349 commonsourceibias.n462 commonsourceibias.n398 161.3
R23350 commonsourceibias.n461 commonsourceibias.n460 161.3
R23351 commonsourceibias.n459 commonsourceibias.n399 161.3
R23352 commonsourceibias.n458 commonsourceibias.n457 161.3
R23353 commonsourceibias.n455 commonsourceibias.n400 161.3
R23354 commonsourceibias.n453 commonsourceibias.n452 161.3
R23355 commonsourceibias.n451 commonsourceibias.n401 161.3
R23356 commonsourceibias.n450 commonsourceibias.n449 161.3
R23357 commonsourceibias.n447 commonsourceibias.n402 161.3
R23358 commonsourceibias.n446 commonsourceibias.n445 161.3
R23359 commonsourceibias.n444 commonsourceibias.n403 161.3
R23360 commonsourceibias.n443 commonsourceibias.n442 161.3
R23361 commonsourceibias.n440 commonsourceibias.n404 161.3
R23362 commonsourceibias.n438 commonsourceibias.n437 161.3
R23363 commonsourceibias.n436 commonsourceibias.n405 161.3
R23364 commonsourceibias.n435 commonsourceibias.n434 161.3
R23365 commonsourceibias.n432 commonsourceibias.n406 161.3
R23366 commonsourceibias.n431 commonsourceibias.n430 161.3
R23367 commonsourceibias.n429 commonsourceibias.n407 161.3
R23368 commonsourceibias.n428 commonsourceibias.n427 161.3
R23369 commonsourceibias.n425 commonsourceibias.n408 161.3
R23370 commonsourceibias.n423 commonsourceibias.n422 161.3
R23371 commonsourceibias.n421 commonsourceibias.n409 161.3
R23372 commonsourceibias.n420 commonsourceibias.n419 161.3
R23373 commonsourceibias.n417 commonsourceibias.n410 161.3
R23374 commonsourceibias.n416 commonsourceibias.n415 161.3
R23375 commonsourceibias.n414 commonsourceibias.n411 161.3
R23376 commonsourceibias.n570 commonsourceibias.n569 161.3
R23377 commonsourceibias.n568 commonsourceibias.n567 161.3
R23378 commonsourceibias.n566 commonsourceibias.n516 161.3
R23379 commonsourceibias.n565 commonsourceibias.n564 161.3
R23380 commonsourceibias.n563 commonsourceibias.n562 161.3
R23381 commonsourceibias.n561 commonsourceibias.n518 161.3
R23382 commonsourceibias.n560 commonsourceibias.n559 161.3
R23383 commonsourceibias.n558 commonsourceibias.n557 161.3
R23384 commonsourceibias.n556 commonsourceibias.n520 161.3
R23385 commonsourceibias.n554 commonsourceibias.n553 161.3
R23386 commonsourceibias.n552 commonsourceibias.n521 161.3
R23387 commonsourceibias.n551 commonsourceibias.n550 161.3
R23388 commonsourceibias.n548 commonsourceibias.n522 161.3
R23389 commonsourceibias.n547 commonsourceibias.n546 161.3
R23390 commonsourceibias.n545 commonsourceibias.n523 161.3
R23391 commonsourceibias.n544 commonsourceibias.n543 161.3
R23392 commonsourceibias.n541 commonsourceibias.n524 161.3
R23393 commonsourceibias.n539 commonsourceibias.n538 161.3
R23394 commonsourceibias.n537 commonsourceibias.n525 161.3
R23395 commonsourceibias.n536 commonsourceibias.n535 161.3
R23396 commonsourceibias.n533 commonsourceibias.n526 161.3
R23397 commonsourceibias.n532 commonsourceibias.n531 161.3
R23398 commonsourceibias.n530 commonsourceibias.n527 161.3
R23399 commonsourceibias.n615 commonsourceibias.n367 161.3
R23400 commonsourceibias.n613 commonsourceibias.n612 161.3
R23401 commonsourceibias.n611 commonsourceibias.n368 161.3
R23402 commonsourceibias.n610 commonsourceibias.n609 161.3
R23403 commonsourceibias.n607 commonsourceibias.n369 161.3
R23404 commonsourceibias.n606 commonsourceibias.n605 161.3
R23405 commonsourceibias.n604 commonsourceibias.n370 161.3
R23406 commonsourceibias.n603 commonsourceibias.n602 161.3
R23407 commonsourceibias.n600 commonsourceibias.n371 161.3
R23408 commonsourceibias.n598 commonsourceibias.n597 161.3
R23409 commonsourceibias.n596 commonsourceibias.n372 161.3
R23410 commonsourceibias.n595 commonsourceibias.n594 161.3
R23411 commonsourceibias.n592 commonsourceibias.n373 161.3
R23412 commonsourceibias.n591 commonsourceibias.n590 161.3
R23413 commonsourceibias.n589 commonsourceibias.n374 161.3
R23414 commonsourceibias.n588 commonsourceibias.n587 161.3
R23415 commonsourceibias.n585 commonsourceibias.n375 161.3
R23416 commonsourceibias.n583 commonsourceibias.n582 161.3
R23417 commonsourceibias.n581 commonsourceibias.n376 161.3
R23418 commonsourceibias.n580 commonsourceibias.n579 161.3
R23419 commonsourceibias.n577 commonsourceibias.n377 161.3
R23420 commonsourceibias.n576 commonsourceibias.n575 161.3
R23421 commonsourceibias.n574 commonsourceibias.n378 161.3
R23422 commonsourceibias.n573 commonsourceibias.n572 161.3
R23423 commonsourceibias.n141 commonsourceibias.n139 81.5057
R23424 commonsourceibias.n381 commonsourceibias.n379 81.5057
R23425 commonsourceibias.n141 commonsourceibias.n140 80.9324
R23426 commonsourceibias.n143 commonsourceibias.n142 80.9324
R23427 commonsourceibias.n145 commonsourceibias.n144 80.9324
R23428 commonsourceibias.n147 commonsourceibias.n146 80.9324
R23429 commonsourceibias.n138 commonsourceibias.n137 80.9324
R23430 commonsourceibias.n136 commonsourceibias.n135 80.9324
R23431 commonsourceibias.n134 commonsourceibias.n133 80.9324
R23432 commonsourceibias.n132 commonsourceibias.n131 80.9324
R23433 commonsourceibias.n130 commonsourceibias.n129 80.9324
R23434 commonsourceibias.n504 commonsourceibias.n503 80.9324
R23435 commonsourceibias.n506 commonsourceibias.n505 80.9324
R23436 commonsourceibias.n508 commonsourceibias.n507 80.9324
R23437 commonsourceibias.n510 commonsourceibias.n509 80.9324
R23438 commonsourceibias.n512 commonsourceibias.n511 80.9324
R23439 commonsourceibias.n387 commonsourceibias.n386 80.9324
R23440 commonsourceibias.n385 commonsourceibias.n384 80.9324
R23441 commonsourceibias.n383 commonsourceibias.n382 80.9324
R23442 commonsourceibias.n381 commonsourceibias.n380 80.9324
R23443 commonsourceibias.n365 commonsourceibias.n364 80.6037
R23444 commonsourceibias.n128 commonsourceibias.n127 80.6037
R23445 commonsourceibias.n250 commonsourceibias.n249 80.6037
R23446 commonsourceibias.n732 commonsourceibias.n731 80.6037
R23447 commonsourceibias.n502 commonsourceibias.n501 80.6037
R23448 commonsourceibias.n617 commonsourceibias.n616 80.6037
R23449 commonsourceibias.n322 commonsourceibias.n321 56.5617
R23450 commonsourceibias.n336 commonsourceibias.n335 56.5617
R23451 commonsourceibias.n85 commonsourceibias.n84 56.5617
R23452 commonsourceibias.n71 commonsourceibias.n70 56.5617
R23453 commonsourceibias.n207 commonsourceibias.n206 56.5617
R23454 commonsourceibias.n193 commonsourceibias.n192 56.5617
R23455 commonsourceibias.n687 commonsourceibias.n685 56.5617
R23456 commonsourceibias.n702 commonsourceibias.n700 56.5617
R23457 commonsourceibias.n457 commonsourceibias.n455 56.5617
R23458 commonsourceibias.n472 commonsourceibias.n470 56.5617
R23459 commonsourceibias.n572 commonsourceibias.n570 56.5617
R23460 commonsourceibias.n294 commonsourceibias.n293 56.5617
R23461 commonsourceibias.n308 commonsourceibias.n307 56.5617
R23462 commonsourceibias.n350 commonsourceibias.n349 56.5617
R23463 commonsourceibias.n113 commonsourceibias.n112 56.5617
R23464 commonsourceibias.n99 commonsourceibias.n98 56.5617
R23465 commonsourceibias.n57 commonsourceibias.n56 56.5617
R23466 commonsourceibias.n235 commonsourceibias.n234 56.5617
R23467 commonsourceibias.n221 commonsourceibias.n220 56.5617
R23468 commonsourceibias.n179 commonsourceibias.n178 56.5617
R23469 commonsourceibias.n657 commonsourceibias.n655 56.5617
R23470 commonsourceibias.n672 commonsourceibias.n670 56.5617
R23471 commonsourceibias.n717 commonsourceibias.n715 56.5617
R23472 commonsourceibias.n427 commonsourceibias.n425 56.5617
R23473 commonsourceibias.n442 commonsourceibias.n440 56.5617
R23474 commonsourceibias.n487 commonsourceibias.n485 56.5617
R23475 commonsourceibias.n602 commonsourceibias.n600 56.5617
R23476 commonsourceibias.n587 commonsourceibias.n585 56.5617
R23477 commonsourceibias.n543 commonsourceibias.n541 56.5617
R23478 commonsourceibias.n557 commonsourceibias.n556 56.5617
R23479 commonsourceibias.n285 commonsourceibias.n284 51.2335
R23480 commonsourceibias.n357 commonsourceibias.n252 51.2335
R23481 commonsourceibias.n120 commonsourceibias.n15 51.2335
R23482 commonsourceibias.n48 commonsourceibias.n47 51.2335
R23483 commonsourceibias.n242 commonsourceibias.n1 51.2335
R23484 commonsourceibias.n170 commonsourceibias.n169 51.2335
R23485 commonsourceibias.n647 commonsourceibias.n646 51.2335
R23486 commonsourceibias.n724 commonsourceibias.n619 51.2335
R23487 commonsourceibias.n417 commonsourceibias.n416 51.2335
R23488 commonsourceibias.n494 commonsourceibias.n389 51.2335
R23489 commonsourceibias.n609 commonsourceibias.n368 51.2335
R23490 commonsourceibias.n533 commonsourceibias.n532 51.2335
R23491 commonsourceibias.n364 commonsourceibias.n363 50.9056
R23492 commonsourceibias.n127 commonsourceibias.n126 50.9056
R23493 commonsourceibias.n249 commonsourceibias.n248 50.9056
R23494 commonsourceibias.n731 commonsourceibias.n730 50.9056
R23495 commonsourceibias.n501 commonsourceibias.n500 50.9056
R23496 commonsourceibias.n616 commonsourceibias.n615 50.9056
R23497 commonsourceibias.n299 commonsourceibias.n298 50.2647
R23498 commonsourceibias.n343 commonsourceibias.n257 50.2647
R23499 commonsourceibias.n106 commonsourceibias.n20 50.2647
R23500 commonsourceibias.n62 commonsourceibias.n61 50.2647
R23501 commonsourceibias.n228 commonsourceibias.n6 50.2647
R23502 commonsourceibias.n184 commonsourceibias.n183 50.2647
R23503 commonsourceibias.n662 commonsourceibias.n661 50.2647
R23504 commonsourceibias.n709 commonsourceibias.n623 50.2647
R23505 commonsourceibias.n432 commonsourceibias.n431 50.2647
R23506 commonsourceibias.n479 commonsourceibias.n393 50.2647
R23507 commonsourceibias.n594 commonsourceibias.n372 50.2647
R23508 commonsourceibias.n548 commonsourceibias.n547 50.2647
R23509 commonsourceibias.n281 commonsourceibias.n280 49.9027
R23510 commonsourceibias.n44 commonsourceibias.n43 49.9027
R23511 commonsourceibias.n166 commonsourceibias.n165 49.9027
R23512 commonsourceibias.n643 commonsourceibias.n642 49.9027
R23513 commonsourceibias.n413 commonsourceibias.n412 49.9027
R23514 commonsourceibias.n529 commonsourceibias.n528 49.9027
R23515 commonsourceibias.n313 commonsourceibias.n312 49.296
R23516 commonsourceibias.n329 commonsourceibias.n262 49.296
R23517 commonsourceibias.n92 commonsourceibias.n25 49.296
R23518 commonsourceibias.n76 commonsourceibias.n75 49.296
R23519 commonsourceibias.n214 commonsourceibias.n11 49.296
R23520 commonsourceibias.n198 commonsourceibias.n197 49.296
R23521 commonsourceibias.n677 commonsourceibias.n676 49.296
R23522 commonsourceibias.n694 commonsourceibias.n627 49.296
R23523 commonsourceibias.n447 commonsourceibias.n446 49.296
R23524 commonsourceibias.n464 commonsourceibias.n397 49.296
R23525 commonsourceibias.n579 commonsourceibias.n376 49.296
R23526 commonsourceibias.n562 commonsourceibias.n561 49.296
R23527 commonsourceibias.n315 commonsourceibias.n267 48.3272
R23528 commonsourceibias.n327 commonsourceibias.n326 48.3272
R23529 commonsourceibias.n90 commonsourceibias.n89 48.3272
R23530 commonsourceibias.n78 commonsourceibias.n30 48.3272
R23531 commonsourceibias.n212 commonsourceibias.n211 48.3272
R23532 commonsourceibias.n202 commonsourceibias.n201 48.3272
R23533 commonsourceibias.n679 commonsourceibias.n631 48.3272
R23534 commonsourceibias.n692 commonsourceibias.n691 48.3272
R23535 commonsourceibias.n449 commonsourceibias.n401 48.3272
R23536 commonsourceibias.n462 commonsourceibias.n461 48.3272
R23537 commonsourceibias.n577 commonsourceibias.n576 48.3272
R23538 commonsourceibias.n566 commonsourceibias.n565 48.3272
R23539 commonsourceibias.n301 commonsourceibias.n272 47.3584
R23540 commonsourceibias.n341 commonsourceibias.n340 47.3584
R23541 commonsourceibias.n104 commonsourceibias.n103 47.3584
R23542 commonsourceibias.n64 commonsourceibias.n35 47.3584
R23543 commonsourceibias.n226 commonsourceibias.n225 47.3584
R23544 commonsourceibias.n186 commonsourceibias.n157 47.3584
R23545 commonsourceibias.n664 commonsourceibias.n635 47.3584
R23546 commonsourceibias.n707 commonsourceibias.n706 47.3584
R23547 commonsourceibias.n434 commonsourceibias.n405 47.3584
R23548 commonsourceibias.n477 commonsourceibias.n476 47.3584
R23549 commonsourceibias.n592 commonsourceibias.n591 47.3584
R23550 commonsourceibias.n550 commonsourceibias.n521 47.3584
R23551 commonsourceibias.n287 commonsourceibias.n277 46.3896
R23552 commonsourceibias.n355 commonsourceibias.n354 46.3896
R23553 commonsourceibias.n118 commonsourceibias.n117 46.3896
R23554 commonsourceibias.n50 commonsourceibias.n40 46.3896
R23555 commonsourceibias.n240 commonsourceibias.n239 46.3896
R23556 commonsourceibias.n172 commonsourceibias.n162 46.3896
R23557 commonsourceibias.n649 commonsourceibias.n639 46.3896
R23558 commonsourceibias.n722 commonsourceibias.n721 46.3896
R23559 commonsourceibias.n419 commonsourceibias.n409 46.3896
R23560 commonsourceibias.n492 commonsourceibias.n491 46.3896
R23561 commonsourceibias.n607 commonsourceibias.n606 46.3896
R23562 commonsourceibias.n535 commonsourceibias.n525 46.3896
R23563 commonsourceibias.n282 commonsourceibias.n281 44.7059
R23564 commonsourceibias.n644 commonsourceibias.n643 44.7059
R23565 commonsourceibias.n414 commonsourceibias.n413 44.7059
R23566 commonsourceibias.n530 commonsourceibias.n529 44.7059
R23567 commonsourceibias.n45 commonsourceibias.n44 44.7059
R23568 commonsourceibias.n167 commonsourceibias.n166 44.7059
R23569 commonsourceibias.n291 commonsourceibias.n277 34.7644
R23570 commonsourceibias.n354 commonsourceibias.n254 34.7644
R23571 commonsourceibias.n117 commonsourceibias.n17 34.7644
R23572 commonsourceibias.n54 commonsourceibias.n40 34.7644
R23573 commonsourceibias.n239 commonsourceibias.n3 34.7644
R23574 commonsourceibias.n176 commonsourceibias.n162 34.7644
R23575 commonsourceibias.n653 commonsourceibias.n639 34.7644
R23576 commonsourceibias.n721 commonsourceibias.n621 34.7644
R23577 commonsourceibias.n423 commonsourceibias.n409 34.7644
R23578 commonsourceibias.n491 commonsourceibias.n391 34.7644
R23579 commonsourceibias.n606 commonsourceibias.n370 34.7644
R23580 commonsourceibias.n539 commonsourceibias.n525 34.7644
R23581 commonsourceibias.n305 commonsourceibias.n272 33.7956
R23582 commonsourceibias.n340 commonsourceibias.n259 33.7956
R23583 commonsourceibias.n103 commonsourceibias.n22 33.7956
R23584 commonsourceibias.n68 commonsourceibias.n35 33.7956
R23585 commonsourceibias.n225 commonsourceibias.n8 33.7956
R23586 commonsourceibias.n190 commonsourceibias.n157 33.7956
R23587 commonsourceibias.n668 commonsourceibias.n635 33.7956
R23588 commonsourceibias.n706 commonsourceibias.n625 33.7956
R23589 commonsourceibias.n438 commonsourceibias.n405 33.7956
R23590 commonsourceibias.n476 commonsourceibias.n395 33.7956
R23591 commonsourceibias.n591 commonsourceibias.n374 33.7956
R23592 commonsourceibias.n554 commonsourceibias.n521 33.7956
R23593 commonsourceibias.n319 commonsourceibias.n267 32.8269
R23594 commonsourceibias.n326 commonsourceibias.n264 32.8269
R23595 commonsourceibias.n89 commonsourceibias.n27 32.8269
R23596 commonsourceibias.n82 commonsourceibias.n30 32.8269
R23597 commonsourceibias.n211 commonsourceibias.n13 32.8269
R23598 commonsourceibias.n203 commonsourceibias.n202 32.8269
R23599 commonsourceibias.n683 commonsourceibias.n631 32.8269
R23600 commonsourceibias.n691 commonsourceibias.n629 32.8269
R23601 commonsourceibias.n453 commonsourceibias.n401 32.8269
R23602 commonsourceibias.n461 commonsourceibias.n399 32.8269
R23603 commonsourceibias.n576 commonsourceibias.n378 32.8269
R23604 commonsourceibias.n567 commonsourceibias.n566 32.8269
R23605 commonsourceibias.n312 commonsourceibias.n269 31.8581
R23606 commonsourceibias.n333 commonsourceibias.n262 31.8581
R23607 commonsourceibias.n96 commonsourceibias.n25 31.8581
R23608 commonsourceibias.n75 commonsourceibias.n32 31.8581
R23609 commonsourceibias.n218 commonsourceibias.n11 31.8581
R23610 commonsourceibias.n197 commonsourceibias.n196 31.8581
R23611 commonsourceibias.n676 commonsourceibias.n633 31.8581
R23612 commonsourceibias.n698 commonsourceibias.n627 31.8581
R23613 commonsourceibias.n446 commonsourceibias.n403 31.8581
R23614 commonsourceibias.n468 commonsourceibias.n397 31.8581
R23615 commonsourceibias.n583 commonsourceibias.n376 31.8581
R23616 commonsourceibias.n561 commonsourceibias.n560 31.8581
R23617 commonsourceibias.n298 commonsourceibias.n274 30.8893
R23618 commonsourceibias.n347 commonsourceibias.n257 30.8893
R23619 commonsourceibias.n110 commonsourceibias.n20 30.8893
R23620 commonsourceibias.n61 commonsourceibias.n37 30.8893
R23621 commonsourceibias.n232 commonsourceibias.n6 30.8893
R23622 commonsourceibias.n183 commonsourceibias.n159 30.8893
R23623 commonsourceibias.n661 commonsourceibias.n637 30.8893
R23624 commonsourceibias.n713 commonsourceibias.n623 30.8893
R23625 commonsourceibias.n431 commonsourceibias.n407 30.8893
R23626 commonsourceibias.n483 commonsourceibias.n393 30.8893
R23627 commonsourceibias.n598 commonsourceibias.n372 30.8893
R23628 commonsourceibias.n547 commonsourceibias.n523 30.8893
R23629 commonsourceibias.n284 commonsourceibias.n279 29.9206
R23630 commonsourceibias.n361 commonsourceibias.n252 29.9206
R23631 commonsourceibias.n124 commonsourceibias.n15 29.9206
R23632 commonsourceibias.n47 commonsourceibias.n42 29.9206
R23633 commonsourceibias.n246 commonsourceibias.n1 29.9206
R23634 commonsourceibias.n169 commonsourceibias.n164 29.9206
R23635 commonsourceibias.n646 commonsourceibias.n641 29.9206
R23636 commonsourceibias.n728 commonsourceibias.n619 29.9206
R23637 commonsourceibias.n416 commonsourceibias.n411 29.9206
R23638 commonsourceibias.n498 commonsourceibias.n389 29.9206
R23639 commonsourceibias.n613 commonsourceibias.n368 29.9206
R23640 commonsourceibias.n532 commonsourceibias.n527 29.9206
R23641 commonsourceibias.n363 commonsourceibias.n362 21.8872
R23642 commonsourceibias.n126 commonsourceibias.n125 21.8872
R23643 commonsourceibias.n248 commonsourceibias.n247 21.8872
R23644 commonsourceibias.n730 commonsourceibias.n729 21.8872
R23645 commonsourceibias.n500 commonsourceibias.n499 21.8872
R23646 commonsourceibias.n615 commonsourceibias.n614 21.8872
R23647 commonsourceibias.n294 commonsourceibias.n276 21.3954
R23648 commonsourceibias.n349 commonsourceibias.n348 21.3954
R23649 commonsourceibias.n112 commonsourceibias.n111 21.3954
R23650 commonsourceibias.n57 commonsourceibias.n39 21.3954
R23651 commonsourceibias.n234 commonsourceibias.n233 21.3954
R23652 commonsourceibias.n179 commonsourceibias.n161 21.3954
R23653 commonsourceibias.n657 commonsourceibias.n656 21.3954
R23654 commonsourceibias.n715 commonsourceibias.n714 21.3954
R23655 commonsourceibias.n427 commonsourceibias.n426 21.3954
R23656 commonsourceibias.n485 commonsourceibias.n484 21.3954
R23657 commonsourceibias.n600 commonsourceibias.n599 21.3954
R23658 commonsourceibias.n543 commonsourceibias.n542 21.3954
R23659 commonsourceibias.n308 commonsourceibias.n271 20.9036
R23660 commonsourceibias.n335 commonsourceibias.n334 20.9036
R23661 commonsourceibias.n98 commonsourceibias.n97 20.9036
R23662 commonsourceibias.n71 commonsourceibias.n34 20.9036
R23663 commonsourceibias.n220 commonsourceibias.n219 20.9036
R23664 commonsourceibias.n193 commonsourceibias.n155 20.9036
R23665 commonsourceibias.n672 commonsourceibias.n671 20.9036
R23666 commonsourceibias.n700 commonsourceibias.n699 20.9036
R23667 commonsourceibias.n442 commonsourceibias.n441 20.9036
R23668 commonsourceibias.n470 commonsourceibias.n469 20.9036
R23669 commonsourceibias.n585 commonsourceibias.n584 20.9036
R23670 commonsourceibias.n557 commonsourceibias.n519 20.9036
R23671 commonsourceibias.n321 commonsourceibias.n320 20.4117
R23672 commonsourceibias.n322 commonsourceibias.n266 20.4117
R23673 commonsourceibias.n85 commonsourceibias.n29 20.4117
R23674 commonsourceibias.n84 commonsourceibias.n83 20.4117
R23675 commonsourceibias.n207 commonsourceibias.n150 20.4117
R23676 commonsourceibias.n206 commonsourceibias.n151 20.4117
R23677 commonsourceibias.n685 commonsourceibias.n684 20.4117
R23678 commonsourceibias.n687 commonsourceibias.n686 20.4117
R23679 commonsourceibias.n455 commonsourceibias.n454 20.4117
R23680 commonsourceibias.n457 commonsourceibias.n456 20.4117
R23681 commonsourceibias.n572 commonsourceibias.n571 20.4117
R23682 commonsourceibias.n570 commonsourceibias.n515 20.4117
R23683 commonsourceibias.n307 commonsourceibias.n306 19.9199
R23684 commonsourceibias.n336 commonsourceibias.n261 19.9199
R23685 commonsourceibias.n99 commonsourceibias.n24 19.9199
R23686 commonsourceibias.n70 commonsourceibias.n69 19.9199
R23687 commonsourceibias.n221 commonsourceibias.n10 19.9199
R23688 commonsourceibias.n192 commonsourceibias.n191 19.9199
R23689 commonsourceibias.n670 commonsourceibias.n669 19.9199
R23690 commonsourceibias.n702 commonsourceibias.n701 19.9199
R23691 commonsourceibias.n440 commonsourceibias.n439 19.9199
R23692 commonsourceibias.n472 commonsourceibias.n471 19.9199
R23693 commonsourceibias.n587 commonsourceibias.n586 19.9199
R23694 commonsourceibias.n556 commonsourceibias.n555 19.9199
R23695 commonsourceibias.n293 commonsourceibias.n292 19.4281
R23696 commonsourceibias.n350 commonsourceibias.n256 19.4281
R23697 commonsourceibias.n113 commonsourceibias.n19 19.4281
R23698 commonsourceibias.n56 commonsourceibias.n55 19.4281
R23699 commonsourceibias.n235 commonsourceibias.n5 19.4281
R23700 commonsourceibias.n178 commonsourceibias.n177 19.4281
R23701 commonsourceibias.n655 commonsourceibias.n654 19.4281
R23702 commonsourceibias.n717 commonsourceibias.n716 19.4281
R23703 commonsourceibias.n425 commonsourceibias.n424 19.4281
R23704 commonsourceibias.n487 commonsourceibias.n486 19.4281
R23705 commonsourceibias.n602 commonsourceibias.n601 19.4281
R23706 commonsourceibias.n541 commonsourceibias.n540 19.4281
R23707 commonsourceibias.n286 commonsourceibias.n285 13.526
R23708 commonsourceibias.n357 commonsourceibias.n356 13.526
R23709 commonsourceibias.n120 commonsourceibias.n119 13.526
R23710 commonsourceibias.n49 commonsourceibias.n48 13.526
R23711 commonsourceibias.n242 commonsourceibias.n241 13.526
R23712 commonsourceibias.n171 commonsourceibias.n170 13.526
R23713 commonsourceibias.n648 commonsourceibias.n647 13.526
R23714 commonsourceibias.n724 commonsourceibias.n723 13.526
R23715 commonsourceibias.n418 commonsourceibias.n417 13.526
R23716 commonsourceibias.n494 commonsourceibias.n493 13.526
R23717 commonsourceibias.n609 commonsourceibias.n608 13.526
R23718 commonsourceibias.n534 commonsourceibias.n533 13.526
R23719 commonsourceibias.n130 commonsourceibias.n128 13.2322
R23720 commonsourceibias.n504 commonsourceibias.n502 13.2322
R23721 commonsourceibias.n300 commonsourceibias.n299 13.0342
R23722 commonsourceibias.n343 commonsourceibias.n342 13.0342
R23723 commonsourceibias.n106 commonsourceibias.n105 13.0342
R23724 commonsourceibias.n63 commonsourceibias.n62 13.0342
R23725 commonsourceibias.n228 commonsourceibias.n227 13.0342
R23726 commonsourceibias.n185 commonsourceibias.n184 13.0342
R23727 commonsourceibias.n663 commonsourceibias.n662 13.0342
R23728 commonsourceibias.n709 commonsourceibias.n708 13.0342
R23729 commonsourceibias.n433 commonsourceibias.n432 13.0342
R23730 commonsourceibias.n479 commonsourceibias.n478 13.0342
R23731 commonsourceibias.n594 commonsourceibias.n593 13.0342
R23732 commonsourceibias.n549 commonsourceibias.n548 13.0342
R23733 commonsourceibias.n314 commonsourceibias.n313 12.5423
R23734 commonsourceibias.n329 commonsourceibias.n328 12.5423
R23735 commonsourceibias.n92 commonsourceibias.n91 12.5423
R23736 commonsourceibias.n77 commonsourceibias.n76 12.5423
R23737 commonsourceibias.n214 commonsourceibias.n213 12.5423
R23738 commonsourceibias.n198 commonsourceibias.n153 12.5423
R23739 commonsourceibias.n678 commonsourceibias.n677 12.5423
R23740 commonsourceibias.n694 commonsourceibias.n693 12.5423
R23741 commonsourceibias.n448 commonsourceibias.n447 12.5423
R23742 commonsourceibias.n464 commonsourceibias.n463 12.5423
R23743 commonsourceibias.n579 commonsourceibias.n578 12.5423
R23744 commonsourceibias.n562 commonsourceibias.n517 12.5423
R23745 commonsourceibias.n734 commonsourceibias.n366 12.2777
R23746 commonsourceibias.n315 commonsourceibias.n314 12.0505
R23747 commonsourceibias.n328 commonsourceibias.n327 12.0505
R23748 commonsourceibias.n91 commonsourceibias.n90 12.0505
R23749 commonsourceibias.n78 commonsourceibias.n77 12.0505
R23750 commonsourceibias.n213 commonsourceibias.n212 12.0505
R23751 commonsourceibias.n201 commonsourceibias.n153 12.0505
R23752 commonsourceibias.n679 commonsourceibias.n678 12.0505
R23753 commonsourceibias.n693 commonsourceibias.n692 12.0505
R23754 commonsourceibias.n449 commonsourceibias.n448 12.0505
R23755 commonsourceibias.n463 commonsourceibias.n462 12.0505
R23756 commonsourceibias.n578 commonsourceibias.n577 12.0505
R23757 commonsourceibias.n565 commonsourceibias.n517 12.0505
R23758 commonsourceibias.n301 commonsourceibias.n300 11.5587
R23759 commonsourceibias.n342 commonsourceibias.n341 11.5587
R23760 commonsourceibias.n105 commonsourceibias.n104 11.5587
R23761 commonsourceibias.n64 commonsourceibias.n63 11.5587
R23762 commonsourceibias.n227 commonsourceibias.n226 11.5587
R23763 commonsourceibias.n186 commonsourceibias.n185 11.5587
R23764 commonsourceibias.n664 commonsourceibias.n663 11.5587
R23765 commonsourceibias.n708 commonsourceibias.n707 11.5587
R23766 commonsourceibias.n434 commonsourceibias.n433 11.5587
R23767 commonsourceibias.n478 commonsourceibias.n477 11.5587
R23768 commonsourceibias.n593 commonsourceibias.n592 11.5587
R23769 commonsourceibias.n550 commonsourceibias.n549 11.5587
R23770 commonsourceibias.n287 commonsourceibias.n286 11.0668
R23771 commonsourceibias.n356 commonsourceibias.n355 11.0668
R23772 commonsourceibias.n119 commonsourceibias.n118 11.0668
R23773 commonsourceibias.n50 commonsourceibias.n49 11.0668
R23774 commonsourceibias.n241 commonsourceibias.n240 11.0668
R23775 commonsourceibias.n172 commonsourceibias.n171 11.0668
R23776 commonsourceibias.n649 commonsourceibias.n648 11.0668
R23777 commonsourceibias.n723 commonsourceibias.n722 11.0668
R23778 commonsourceibias.n419 commonsourceibias.n418 11.0668
R23779 commonsourceibias.n493 commonsourceibias.n492 11.0668
R23780 commonsourceibias.n608 commonsourceibias.n607 11.0668
R23781 commonsourceibias.n535 commonsourceibias.n534 11.0668
R23782 commonsourceibias.n734 commonsourceibias.n733 10.3347
R23783 commonsourceibias.n149 commonsourceibias.n148 9.50363
R23784 commonsourceibias.n514 commonsourceibias.n513 9.50363
R23785 commonsourceibias.n366 commonsourceibias.n250 8.75852
R23786 commonsourceibias.n733 commonsourceibias.n617 8.75852
R23787 commonsourceibias.n292 commonsourceibias.n291 5.16479
R23788 commonsourceibias.n256 commonsourceibias.n254 5.16479
R23789 commonsourceibias.n19 commonsourceibias.n17 5.16479
R23790 commonsourceibias.n55 commonsourceibias.n54 5.16479
R23791 commonsourceibias.n5 commonsourceibias.n3 5.16479
R23792 commonsourceibias.n177 commonsourceibias.n176 5.16479
R23793 commonsourceibias.n654 commonsourceibias.n653 5.16479
R23794 commonsourceibias.n716 commonsourceibias.n621 5.16479
R23795 commonsourceibias.n424 commonsourceibias.n423 5.16479
R23796 commonsourceibias.n486 commonsourceibias.n391 5.16479
R23797 commonsourceibias.n601 commonsourceibias.n370 5.16479
R23798 commonsourceibias.n540 commonsourceibias.n539 5.16479
R23799 commonsourceibias.n366 commonsourceibias.n365 5.03125
R23800 commonsourceibias.n733 commonsourceibias.n732 5.03125
R23801 commonsourceibias.n306 commonsourceibias.n305 4.67295
R23802 commonsourceibias.n261 commonsourceibias.n259 4.67295
R23803 commonsourceibias.n24 commonsourceibias.n22 4.67295
R23804 commonsourceibias.n69 commonsourceibias.n68 4.67295
R23805 commonsourceibias.n10 commonsourceibias.n8 4.67295
R23806 commonsourceibias.n191 commonsourceibias.n190 4.67295
R23807 commonsourceibias.n669 commonsourceibias.n668 4.67295
R23808 commonsourceibias.n701 commonsourceibias.n625 4.67295
R23809 commonsourceibias.n439 commonsourceibias.n438 4.67295
R23810 commonsourceibias.n471 commonsourceibias.n395 4.67295
R23811 commonsourceibias.n586 commonsourceibias.n374 4.67295
R23812 commonsourceibias.n555 commonsourceibias.n554 4.67295
R23813 commonsourceibias commonsourceibias.n734 4.20978
R23814 commonsourceibias.n320 commonsourceibias.n319 4.18111
R23815 commonsourceibias.n266 commonsourceibias.n264 4.18111
R23816 commonsourceibias.n29 commonsourceibias.n27 4.18111
R23817 commonsourceibias.n83 commonsourceibias.n82 4.18111
R23818 commonsourceibias.n150 commonsourceibias.n13 4.18111
R23819 commonsourceibias.n203 commonsourceibias.n151 4.18111
R23820 commonsourceibias.n684 commonsourceibias.n683 4.18111
R23821 commonsourceibias.n686 commonsourceibias.n629 4.18111
R23822 commonsourceibias.n454 commonsourceibias.n453 4.18111
R23823 commonsourceibias.n456 commonsourceibias.n399 4.18111
R23824 commonsourceibias.n571 commonsourceibias.n378 4.18111
R23825 commonsourceibias.n567 commonsourceibias.n515 4.18111
R23826 commonsourceibias.n271 commonsourceibias.n269 3.68928
R23827 commonsourceibias.n334 commonsourceibias.n333 3.68928
R23828 commonsourceibias.n97 commonsourceibias.n96 3.68928
R23829 commonsourceibias.n34 commonsourceibias.n32 3.68928
R23830 commonsourceibias.n219 commonsourceibias.n218 3.68928
R23831 commonsourceibias.n196 commonsourceibias.n155 3.68928
R23832 commonsourceibias.n671 commonsourceibias.n633 3.68928
R23833 commonsourceibias.n699 commonsourceibias.n698 3.68928
R23834 commonsourceibias.n441 commonsourceibias.n403 3.68928
R23835 commonsourceibias.n469 commonsourceibias.n468 3.68928
R23836 commonsourceibias.n584 commonsourceibias.n583 3.68928
R23837 commonsourceibias.n560 commonsourceibias.n519 3.68928
R23838 commonsourceibias.n276 commonsourceibias.n274 3.19744
R23839 commonsourceibias.n348 commonsourceibias.n347 3.19744
R23840 commonsourceibias.n111 commonsourceibias.n110 3.19744
R23841 commonsourceibias.n39 commonsourceibias.n37 3.19744
R23842 commonsourceibias.n233 commonsourceibias.n232 3.19744
R23843 commonsourceibias.n161 commonsourceibias.n159 3.19744
R23844 commonsourceibias.n656 commonsourceibias.n637 3.19744
R23845 commonsourceibias.n714 commonsourceibias.n713 3.19744
R23846 commonsourceibias.n426 commonsourceibias.n407 3.19744
R23847 commonsourceibias.n484 commonsourceibias.n483 3.19744
R23848 commonsourceibias.n599 commonsourceibias.n598 3.19744
R23849 commonsourceibias.n542 commonsourceibias.n523 3.19744
R23850 commonsourceibias.n139 commonsourceibias.t47 2.82907
R23851 commonsourceibias.n139 commonsourceibias.t79 2.82907
R23852 commonsourceibias.n140 commonsourceibias.t55 2.82907
R23853 commonsourceibias.n140 commonsourceibias.t5 2.82907
R23854 commonsourceibias.n142 commonsourceibias.t19 2.82907
R23855 commonsourceibias.n142 commonsourceibias.t23 2.82907
R23856 commonsourceibias.n144 commonsourceibias.t39 2.82907
R23857 commonsourceibias.n144 commonsourceibias.t71 2.82907
R23858 commonsourceibias.n146 commonsourceibias.t57 2.82907
R23859 commonsourceibias.n146 commonsourceibias.t27 2.82907
R23860 commonsourceibias.n137 commonsourceibias.t11 2.82907
R23861 commonsourceibias.n137 commonsourceibias.t41 2.82907
R23862 commonsourceibias.n135 commonsourceibias.t25 2.82907
R23863 commonsourceibias.n135 commonsourceibias.t35 2.82907
R23864 commonsourceibias.n133 commonsourceibias.t37 2.82907
R23865 commonsourceibias.n133 commonsourceibias.t77 2.82907
R23866 commonsourceibias.n131 commonsourceibias.t51 2.82907
R23867 commonsourceibias.n131 commonsourceibias.t9 2.82907
R23868 commonsourceibias.n129 commonsourceibias.t75 2.82907
R23869 commonsourceibias.n129 commonsourceibias.t21 2.82907
R23870 commonsourceibias.n503 commonsourceibias.t43 2.82907
R23871 commonsourceibias.n503 commonsourceibias.t15 2.82907
R23872 commonsourceibias.n505 commonsourceibias.t31 2.82907
R23873 commonsourceibias.n505 commonsourceibias.t1 2.82907
R23874 commonsourceibias.n507 commonsourceibias.t17 2.82907
R23875 commonsourceibias.n507 commonsourceibias.t61 2.82907
R23876 commonsourceibias.n509 commonsourceibias.t59 2.82907
R23877 commonsourceibias.n509 commonsourceibias.t45 2.82907
R23878 commonsourceibias.n511 commonsourceibias.t65 2.82907
R23879 commonsourceibias.n511 commonsourceibias.t33 2.82907
R23880 commonsourceibias.n386 commonsourceibias.t53 2.82907
R23881 commonsourceibias.n386 commonsourceibias.t73 2.82907
R23882 commonsourceibias.n384 commonsourceibias.t7 2.82907
R23883 commonsourceibias.n384 commonsourceibias.t63 2.82907
R23884 commonsourceibias.n382 commonsourceibias.t69 2.82907
R23885 commonsourceibias.n382 commonsourceibias.t67 2.82907
R23886 commonsourceibias.n380 commonsourceibias.t49 2.82907
R23887 commonsourceibias.n380 commonsourceibias.t13 2.82907
R23888 commonsourceibias.n379 commonsourceibias.t29 2.82907
R23889 commonsourceibias.n379 commonsourceibias.t3 2.82907
R23890 commonsourceibias.n280 commonsourceibias.n279 2.7056
R23891 commonsourceibias.n362 commonsourceibias.n361 2.7056
R23892 commonsourceibias.n125 commonsourceibias.n124 2.7056
R23893 commonsourceibias.n43 commonsourceibias.n42 2.7056
R23894 commonsourceibias.n247 commonsourceibias.n246 2.7056
R23895 commonsourceibias.n165 commonsourceibias.n164 2.7056
R23896 commonsourceibias.n642 commonsourceibias.n641 2.7056
R23897 commonsourceibias.n729 commonsourceibias.n728 2.7056
R23898 commonsourceibias.n412 commonsourceibias.n411 2.7056
R23899 commonsourceibias.n499 commonsourceibias.n498 2.7056
R23900 commonsourceibias.n614 commonsourceibias.n613 2.7056
R23901 commonsourceibias.n528 commonsourceibias.n527 2.7056
R23902 commonsourceibias.n132 commonsourceibias.n130 0.573776
R23903 commonsourceibias.n134 commonsourceibias.n132 0.573776
R23904 commonsourceibias.n136 commonsourceibias.n134 0.573776
R23905 commonsourceibias.n138 commonsourceibias.n136 0.573776
R23906 commonsourceibias.n147 commonsourceibias.n145 0.573776
R23907 commonsourceibias.n145 commonsourceibias.n143 0.573776
R23908 commonsourceibias.n143 commonsourceibias.n141 0.573776
R23909 commonsourceibias.n383 commonsourceibias.n381 0.573776
R23910 commonsourceibias.n385 commonsourceibias.n383 0.573776
R23911 commonsourceibias.n387 commonsourceibias.n385 0.573776
R23912 commonsourceibias.n512 commonsourceibias.n510 0.573776
R23913 commonsourceibias.n510 commonsourceibias.n508 0.573776
R23914 commonsourceibias.n508 commonsourceibias.n506 0.573776
R23915 commonsourceibias.n506 commonsourceibias.n504 0.573776
R23916 commonsourceibias.n148 commonsourceibias.n138 0.287138
R23917 commonsourceibias.n148 commonsourceibias.n147 0.287138
R23918 commonsourceibias.n513 commonsourceibias.n387 0.287138
R23919 commonsourceibias.n513 commonsourceibias.n512 0.287138
R23920 commonsourceibias.n365 commonsourceibias.n251 0.285035
R23921 commonsourceibias.n128 commonsourceibias.n14 0.285035
R23922 commonsourceibias.n250 commonsourceibias.n0 0.285035
R23923 commonsourceibias.n732 commonsourceibias.n618 0.285035
R23924 commonsourceibias.n502 commonsourceibias.n388 0.285035
R23925 commonsourceibias.n617 commonsourceibias.n367 0.285035
R23926 commonsourceibias.n360 commonsourceibias.n251 0.189894
R23927 commonsourceibias.n360 commonsourceibias.n359 0.189894
R23928 commonsourceibias.n359 commonsourceibias.n358 0.189894
R23929 commonsourceibias.n358 commonsourceibias.n253 0.189894
R23930 commonsourceibias.n353 commonsourceibias.n253 0.189894
R23931 commonsourceibias.n353 commonsourceibias.n352 0.189894
R23932 commonsourceibias.n352 commonsourceibias.n351 0.189894
R23933 commonsourceibias.n351 commonsourceibias.n255 0.189894
R23934 commonsourceibias.n346 commonsourceibias.n255 0.189894
R23935 commonsourceibias.n346 commonsourceibias.n345 0.189894
R23936 commonsourceibias.n345 commonsourceibias.n344 0.189894
R23937 commonsourceibias.n344 commonsourceibias.n258 0.189894
R23938 commonsourceibias.n339 commonsourceibias.n258 0.189894
R23939 commonsourceibias.n339 commonsourceibias.n338 0.189894
R23940 commonsourceibias.n338 commonsourceibias.n337 0.189894
R23941 commonsourceibias.n337 commonsourceibias.n260 0.189894
R23942 commonsourceibias.n332 commonsourceibias.n260 0.189894
R23943 commonsourceibias.n332 commonsourceibias.n331 0.189894
R23944 commonsourceibias.n331 commonsourceibias.n330 0.189894
R23945 commonsourceibias.n330 commonsourceibias.n263 0.189894
R23946 commonsourceibias.n325 commonsourceibias.n263 0.189894
R23947 commonsourceibias.n325 commonsourceibias.n324 0.189894
R23948 commonsourceibias.n324 commonsourceibias.n323 0.189894
R23949 commonsourceibias.n323 commonsourceibias.n265 0.189894
R23950 commonsourceibias.n318 commonsourceibias.n265 0.189894
R23951 commonsourceibias.n318 commonsourceibias.n317 0.189894
R23952 commonsourceibias.n317 commonsourceibias.n316 0.189894
R23953 commonsourceibias.n316 commonsourceibias.n268 0.189894
R23954 commonsourceibias.n311 commonsourceibias.n268 0.189894
R23955 commonsourceibias.n311 commonsourceibias.n310 0.189894
R23956 commonsourceibias.n310 commonsourceibias.n309 0.189894
R23957 commonsourceibias.n309 commonsourceibias.n270 0.189894
R23958 commonsourceibias.n304 commonsourceibias.n270 0.189894
R23959 commonsourceibias.n304 commonsourceibias.n303 0.189894
R23960 commonsourceibias.n303 commonsourceibias.n302 0.189894
R23961 commonsourceibias.n302 commonsourceibias.n273 0.189894
R23962 commonsourceibias.n297 commonsourceibias.n273 0.189894
R23963 commonsourceibias.n297 commonsourceibias.n296 0.189894
R23964 commonsourceibias.n296 commonsourceibias.n295 0.189894
R23965 commonsourceibias.n295 commonsourceibias.n275 0.189894
R23966 commonsourceibias.n290 commonsourceibias.n275 0.189894
R23967 commonsourceibias.n290 commonsourceibias.n289 0.189894
R23968 commonsourceibias.n289 commonsourceibias.n288 0.189894
R23969 commonsourceibias.n288 commonsourceibias.n278 0.189894
R23970 commonsourceibias.n283 commonsourceibias.n278 0.189894
R23971 commonsourceibias.n283 commonsourceibias.n282 0.189894
R23972 commonsourceibias.n123 commonsourceibias.n14 0.189894
R23973 commonsourceibias.n123 commonsourceibias.n122 0.189894
R23974 commonsourceibias.n122 commonsourceibias.n121 0.189894
R23975 commonsourceibias.n121 commonsourceibias.n16 0.189894
R23976 commonsourceibias.n116 commonsourceibias.n16 0.189894
R23977 commonsourceibias.n116 commonsourceibias.n115 0.189894
R23978 commonsourceibias.n115 commonsourceibias.n114 0.189894
R23979 commonsourceibias.n114 commonsourceibias.n18 0.189894
R23980 commonsourceibias.n109 commonsourceibias.n18 0.189894
R23981 commonsourceibias.n109 commonsourceibias.n108 0.189894
R23982 commonsourceibias.n108 commonsourceibias.n107 0.189894
R23983 commonsourceibias.n107 commonsourceibias.n21 0.189894
R23984 commonsourceibias.n102 commonsourceibias.n21 0.189894
R23985 commonsourceibias.n102 commonsourceibias.n101 0.189894
R23986 commonsourceibias.n101 commonsourceibias.n100 0.189894
R23987 commonsourceibias.n100 commonsourceibias.n23 0.189894
R23988 commonsourceibias.n95 commonsourceibias.n23 0.189894
R23989 commonsourceibias.n95 commonsourceibias.n94 0.189894
R23990 commonsourceibias.n94 commonsourceibias.n93 0.189894
R23991 commonsourceibias.n93 commonsourceibias.n26 0.189894
R23992 commonsourceibias.n88 commonsourceibias.n26 0.189894
R23993 commonsourceibias.n88 commonsourceibias.n87 0.189894
R23994 commonsourceibias.n87 commonsourceibias.n86 0.189894
R23995 commonsourceibias.n86 commonsourceibias.n28 0.189894
R23996 commonsourceibias.n81 commonsourceibias.n28 0.189894
R23997 commonsourceibias.n81 commonsourceibias.n80 0.189894
R23998 commonsourceibias.n80 commonsourceibias.n79 0.189894
R23999 commonsourceibias.n79 commonsourceibias.n31 0.189894
R24000 commonsourceibias.n74 commonsourceibias.n31 0.189894
R24001 commonsourceibias.n74 commonsourceibias.n73 0.189894
R24002 commonsourceibias.n73 commonsourceibias.n72 0.189894
R24003 commonsourceibias.n72 commonsourceibias.n33 0.189894
R24004 commonsourceibias.n67 commonsourceibias.n33 0.189894
R24005 commonsourceibias.n67 commonsourceibias.n66 0.189894
R24006 commonsourceibias.n66 commonsourceibias.n65 0.189894
R24007 commonsourceibias.n65 commonsourceibias.n36 0.189894
R24008 commonsourceibias.n60 commonsourceibias.n36 0.189894
R24009 commonsourceibias.n60 commonsourceibias.n59 0.189894
R24010 commonsourceibias.n59 commonsourceibias.n58 0.189894
R24011 commonsourceibias.n58 commonsourceibias.n38 0.189894
R24012 commonsourceibias.n53 commonsourceibias.n38 0.189894
R24013 commonsourceibias.n53 commonsourceibias.n52 0.189894
R24014 commonsourceibias.n52 commonsourceibias.n51 0.189894
R24015 commonsourceibias.n51 commonsourceibias.n41 0.189894
R24016 commonsourceibias.n46 commonsourceibias.n41 0.189894
R24017 commonsourceibias.n46 commonsourceibias.n45 0.189894
R24018 commonsourceibias.n205 commonsourceibias.n204 0.189894
R24019 commonsourceibias.n204 commonsourceibias.n152 0.189894
R24020 commonsourceibias.n200 commonsourceibias.n152 0.189894
R24021 commonsourceibias.n200 commonsourceibias.n199 0.189894
R24022 commonsourceibias.n199 commonsourceibias.n154 0.189894
R24023 commonsourceibias.n195 commonsourceibias.n154 0.189894
R24024 commonsourceibias.n195 commonsourceibias.n194 0.189894
R24025 commonsourceibias.n194 commonsourceibias.n156 0.189894
R24026 commonsourceibias.n189 commonsourceibias.n156 0.189894
R24027 commonsourceibias.n189 commonsourceibias.n188 0.189894
R24028 commonsourceibias.n188 commonsourceibias.n187 0.189894
R24029 commonsourceibias.n187 commonsourceibias.n158 0.189894
R24030 commonsourceibias.n182 commonsourceibias.n158 0.189894
R24031 commonsourceibias.n182 commonsourceibias.n181 0.189894
R24032 commonsourceibias.n181 commonsourceibias.n180 0.189894
R24033 commonsourceibias.n180 commonsourceibias.n160 0.189894
R24034 commonsourceibias.n175 commonsourceibias.n160 0.189894
R24035 commonsourceibias.n175 commonsourceibias.n174 0.189894
R24036 commonsourceibias.n174 commonsourceibias.n173 0.189894
R24037 commonsourceibias.n173 commonsourceibias.n163 0.189894
R24038 commonsourceibias.n168 commonsourceibias.n163 0.189894
R24039 commonsourceibias.n168 commonsourceibias.n167 0.189894
R24040 commonsourceibias.n245 commonsourceibias.n0 0.189894
R24041 commonsourceibias.n245 commonsourceibias.n244 0.189894
R24042 commonsourceibias.n244 commonsourceibias.n243 0.189894
R24043 commonsourceibias.n243 commonsourceibias.n2 0.189894
R24044 commonsourceibias.n238 commonsourceibias.n2 0.189894
R24045 commonsourceibias.n238 commonsourceibias.n237 0.189894
R24046 commonsourceibias.n237 commonsourceibias.n236 0.189894
R24047 commonsourceibias.n236 commonsourceibias.n4 0.189894
R24048 commonsourceibias.n231 commonsourceibias.n4 0.189894
R24049 commonsourceibias.n231 commonsourceibias.n230 0.189894
R24050 commonsourceibias.n230 commonsourceibias.n229 0.189894
R24051 commonsourceibias.n229 commonsourceibias.n7 0.189894
R24052 commonsourceibias.n224 commonsourceibias.n7 0.189894
R24053 commonsourceibias.n224 commonsourceibias.n223 0.189894
R24054 commonsourceibias.n223 commonsourceibias.n222 0.189894
R24055 commonsourceibias.n222 commonsourceibias.n9 0.189894
R24056 commonsourceibias.n217 commonsourceibias.n9 0.189894
R24057 commonsourceibias.n217 commonsourceibias.n216 0.189894
R24058 commonsourceibias.n216 commonsourceibias.n215 0.189894
R24059 commonsourceibias.n215 commonsourceibias.n12 0.189894
R24060 commonsourceibias.n210 commonsourceibias.n12 0.189894
R24061 commonsourceibias.n210 commonsourceibias.n209 0.189894
R24062 commonsourceibias.n209 commonsourceibias.n208 0.189894
R24063 commonsourceibias.n645 commonsourceibias.n644 0.189894
R24064 commonsourceibias.n645 commonsourceibias.n640 0.189894
R24065 commonsourceibias.n650 commonsourceibias.n640 0.189894
R24066 commonsourceibias.n651 commonsourceibias.n650 0.189894
R24067 commonsourceibias.n652 commonsourceibias.n651 0.189894
R24068 commonsourceibias.n652 commonsourceibias.n638 0.189894
R24069 commonsourceibias.n658 commonsourceibias.n638 0.189894
R24070 commonsourceibias.n659 commonsourceibias.n658 0.189894
R24071 commonsourceibias.n660 commonsourceibias.n659 0.189894
R24072 commonsourceibias.n660 commonsourceibias.n636 0.189894
R24073 commonsourceibias.n665 commonsourceibias.n636 0.189894
R24074 commonsourceibias.n666 commonsourceibias.n665 0.189894
R24075 commonsourceibias.n667 commonsourceibias.n666 0.189894
R24076 commonsourceibias.n667 commonsourceibias.n634 0.189894
R24077 commonsourceibias.n673 commonsourceibias.n634 0.189894
R24078 commonsourceibias.n674 commonsourceibias.n673 0.189894
R24079 commonsourceibias.n675 commonsourceibias.n674 0.189894
R24080 commonsourceibias.n675 commonsourceibias.n632 0.189894
R24081 commonsourceibias.n680 commonsourceibias.n632 0.189894
R24082 commonsourceibias.n681 commonsourceibias.n680 0.189894
R24083 commonsourceibias.n682 commonsourceibias.n681 0.189894
R24084 commonsourceibias.n682 commonsourceibias.n630 0.189894
R24085 commonsourceibias.n688 commonsourceibias.n630 0.189894
R24086 commonsourceibias.n689 commonsourceibias.n688 0.189894
R24087 commonsourceibias.n690 commonsourceibias.n689 0.189894
R24088 commonsourceibias.n690 commonsourceibias.n628 0.189894
R24089 commonsourceibias.n695 commonsourceibias.n628 0.189894
R24090 commonsourceibias.n696 commonsourceibias.n695 0.189894
R24091 commonsourceibias.n697 commonsourceibias.n696 0.189894
R24092 commonsourceibias.n697 commonsourceibias.n626 0.189894
R24093 commonsourceibias.n703 commonsourceibias.n626 0.189894
R24094 commonsourceibias.n704 commonsourceibias.n703 0.189894
R24095 commonsourceibias.n705 commonsourceibias.n704 0.189894
R24096 commonsourceibias.n705 commonsourceibias.n624 0.189894
R24097 commonsourceibias.n710 commonsourceibias.n624 0.189894
R24098 commonsourceibias.n711 commonsourceibias.n710 0.189894
R24099 commonsourceibias.n712 commonsourceibias.n711 0.189894
R24100 commonsourceibias.n712 commonsourceibias.n622 0.189894
R24101 commonsourceibias.n718 commonsourceibias.n622 0.189894
R24102 commonsourceibias.n719 commonsourceibias.n718 0.189894
R24103 commonsourceibias.n720 commonsourceibias.n719 0.189894
R24104 commonsourceibias.n720 commonsourceibias.n620 0.189894
R24105 commonsourceibias.n725 commonsourceibias.n620 0.189894
R24106 commonsourceibias.n726 commonsourceibias.n725 0.189894
R24107 commonsourceibias.n727 commonsourceibias.n726 0.189894
R24108 commonsourceibias.n727 commonsourceibias.n618 0.189894
R24109 commonsourceibias.n415 commonsourceibias.n414 0.189894
R24110 commonsourceibias.n415 commonsourceibias.n410 0.189894
R24111 commonsourceibias.n420 commonsourceibias.n410 0.189894
R24112 commonsourceibias.n421 commonsourceibias.n420 0.189894
R24113 commonsourceibias.n422 commonsourceibias.n421 0.189894
R24114 commonsourceibias.n422 commonsourceibias.n408 0.189894
R24115 commonsourceibias.n428 commonsourceibias.n408 0.189894
R24116 commonsourceibias.n429 commonsourceibias.n428 0.189894
R24117 commonsourceibias.n430 commonsourceibias.n429 0.189894
R24118 commonsourceibias.n430 commonsourceibias.n406 0.189894
R24119 commonsourceibias.n435 commonsourceibias.n406 0.189894
R24120 commonsourceibias.n436 commonsourceibias.n435 0.189894
R24121 commonsourceibias.n437 commonsourceibias.n436 0.189894
R24122 commonsourceibias.n437 commonsourceibias.n404 0.189894
R24123 commonsourceibias.n443 commonsourceibias.n404 0.189894
R24124 commonsourceibias.n444 commonsourceibias.n443 0.189894
R24125 commonsourceibias.n445 commonsourceibias.n444 0.189894
R24126 commonsourceibias.n445 commonsourceibias.n402 0.189894
R24127 commonsourceibias.n450 commonsourceibias.n402 0.189894
R24128 commonsourceibias.n451 commonsourceibias.n450 0.189894
R24129 commonsourceibias.n452 commonsourceibias.n451 0.189894
R24130 commonsourceibias.n452 commonsourceibias.n400 0.189894
R24131 commonsourceibias.n458 commonsourceibias.n400 0.189894
R24132 commonsourceibias.n459 commonsourceibias.n458 0.189894
R24133 commonsourceibias.n460 commonsourceibias.n459 0.189894
R24134 commonsourceibias.n460 commonsourceibias.n398 0.189894
R24135 commonsourceibias.n465 commonsourceibias.n398 0.189894
R24136 commonsourceibias.n466 commonsourceibias.n465 0.189894
R24137 commonsourceibias.n467 commonsourceibias.n466 0.189894
R24138 commonsourceibias.n467 commonsourceibias.n396 0.189894
R24139 commonsourceibias.n473 commonsourceibias.n396 0.189894
R24140 commonsourceibias.n474 commonsourceibias.n473 0.189894
R24141 commonsourceibias.n475 commonsourceibias.n474 0.189894
R24142 commonsourceibias.n475 commonsourceibias.n394 0.189894
R24143 commonsourceibias.n480 commonsourceibias.n394 0.189894
R24144 commonsourceibias.n481 commonsourceibias.n480 0.189894
R24145 commonsourceibias.n482 commonsourceibias.n481 0.189894
R24146 commonsourceibias.n482 commonsourceibias.n392 0.189894
R24147 commonsourceibias.n488 commonsourceibias.n392 0.189894
R24148 commonsourceibias.n489 commonsourceibias.n488 0.189894
R24149 commonsourceibias.n490 commonsourceibias.n489 0.189894
R24150 commonsourceibias.n490 commonsourceibias.n390 0.189894
R24151 commonsourceibias.n495 commonsourceibias.n390 0.189894
R24152 commonsourceibias.n496 commonsourceibias.n495 0.189894
R24153 commonsourceibias.n497 commonsourceibias.n496 0.189894
R24154 commonsourceibias.n497 commonsourceibias.n388 0.189894
R24155 commonsourceibias.n531 commonsourceibias.n530 0.189894
R24156 commonsourceibias.n531 commonsourceibias.n526 0.189894
R24157 commonsourceibias.n536 commonsourceibias.n526 0.189894
R24158 commonsourceibias.n537 commonsourceibias.n536 0.189894
R24159 commonsourceibias.n538 commonsourceibias.n537 0.189894
R24160 commonsourceibias.n538 commonsourceibias.n524 0.189894
R24161 commonsourceibias.n544 commonsourceibias.n524 0.189894
R24162 commonsourceibias.n545 commonsourceibias.n544 0.189894
R24163 commonsourceibias.n546 commonsourceibias.n545 0.189894
R24164 commonsourceibias.n546 commonsourceibias.n522 0.189894
R24165 commonsourceibias.n551 commonsourceibias.n522 0.189894
R24166 commonsourceibias.n552 commonsourceibias.n551 0.189894
R24167 commonsourceibias.n553 commonsourceibias.n552 0.189894
R24168 commonsourceibias.n553 commonsourceibias.n520 0.189894
R24169 commonsourceibias.n558 commonsourceibias.n520 0.189894
R24170 commonsourceibias.n559 commonsourceibias.n558 0.189894
R24171 commonsourceibias.n559 commonsourceibias.n518 0.189894
R24172 commonsourceibias.n563 commonsourceibias.n518 0.189894
R24173 commonsourceibias.n564 commonsourceibias.n563 0.189894
R24174 commonsourceibias.n564 commonsourceibias.n516 0.189894
R24175 commonsourceibias.n568 commonsourceibias.n516 0.189894
R24176 commonsourceibias.n569 commonsourceibias.n568 0.189894
R24177 commonsourceibias.n574 commonsourceibias.n573 0.189894
R24178 commonsourceibias.n575 commonsourceibias.n574 0.189894
R24179 commonsourceibias.n575 commonsourceibias.n377 0.189894
R24180 commonsourceibias.n580 commonsourceibias.n377 0.189894
R24181 commonsourceibias.n581 commonsourceibias.n580 0.189894
R24182 commonsourceibias.n582 commonsourceibias.n581 0.189894
R24183 commonsourceibias.n582 commonsourceibias.n375 0.189894
R24184 commonsourceibias.n588 commonsourceibias.n375 0.189894
R24185 commonsourceibias.n589 commonsourceibias.n588 0.189894
R24186 commonsourceibias.n590 commonsourceibias.n589 0.189894
R24187 commonsourceibias.n590 commonsourceibias.n373 0.189894
R24188 commonsourceibias.n595 commonsourceibias.n373 0.189894
R24189 commonsourceibias.n596 commonsourceibias.n595 0.189894
R24190 commonsourceibias.n597 commonsourceibias.n596 0.189894
R24191 commonsourceibias.n597 commonsourceibias.n371 0.189894
R24192 commonsourceibias.n603 commonsourceibias.n371 0.189894
R24193 commonsourceibias.n604 commonsourceibias.n603 0.189894
R24194 commonsourceibias.n605 commonsourceibias.n604 0.189894
R24195 commonsourceibias.n605 commonsourceibias.n369 0.189894
R24196 commonsourceibias.n610 commonsourceibias.n369 0.189894
R24197 commonsourceibias.n611 commonsourceibias.n610 0.189894
R24198 commonsourceibias.n612 commonsourceibias.n611 0.189894
R24199 commonsourceibias.n612 commonsourceibias.n367 0.189894
R24200 commonsourceibias.n205 commonsourceibias.n149 0.0762576
R24201 commonsourceibias.n208 commonsourceibias.n149 0.0762576
R24202 commonsourceibias.n569 commonsourceibias.n514 0.0762576
R24203 commonsourceibias.n573 commonsourceibias.n514 0.0762576
R24204 minus.n76 minus.t28 250.337
R24205 minus.n15 minus.t20 250.337
R24206 minus.n126 minus.t1 243.255
R24207 minus.n120 minus.t8 231.093
R24208 minus.n59 minus.t10 231.093
R24209 minus.n125 minus.n123 224.169
R24210 minus.n125 minus.n124 223.454
R24211 minus.n62 minus.t12 187.445
R24212 minus.n113 minus.t18 187.445
R24213 minus.n107 minus.t25 187.445
R24214 minus.n66 minus.t22 187.445
R24215 minus.n68 minus.t19 187.445
R24216 minus.n95 minus.t7 187.445
R24217 minus.n89 minus.t6 187.445
R24218 minus.n72 minus.t16 187.445
R24219 minus.n74 minus.t15 187.445
R24220 minus.n77 minus.t23 187.445
R24221 minus.n16 minus.t14 187.445
R24222 minus.n13 minus.t9 187.445
R24223 minus.n11 minus.t5 187.445
R24224 minus.n28 minus.t26 187.445
R24225 minus.n34 minus.t27 187.445
R24226 minus.n7 minus.t21 187.445
R24227 minus.n5 minus.t24 187.445
R24228 minus.n46 minus.t17 187.445
R24229 minus.n52 minus.t11 187.445
R24230 minus.n1 minus.t13 187.445
R24231 minus.n78 minus.n75 161.3
R24232 minus.n80 minus.n79 161.3
R24233 minus.n82 minus.n81 161.3
R24234 minus.n83 minus.n73 161.3
R24235 minus.n85 minus.n84 161.3
R24236 minus.n87 minus.n86 161.3
R24237 minus.n88 minus.n71 161.3
R24238 minus.n91 minus.n90 161.3
R24239 minus.n92 minus.n70 161.3
R24240 minus.n94 minus.n93 161.3
R24241 minus.n96 minus.n69 161.3
R24242 minus.n98 minus.n97 161.3
R24243 minus.n100 minus.n99 161.3
R24244 minus.n101 minus.n67 161.3
R24245 minus.n103 minus.n102 161.3
R24246 minus.n105 minus.n104 161.3
R24247 minus.n106 minus.n65 161.3
R24248 minus.n109 minus.n108 161.3
R24249 minus.n110 minus.n64 161.3
R24250 minus.n112 minus.n111 161.3
R24251 minus.n114 minus.n63 161.3
R24252 minus.n116 minus.n115 161.3
R24253 minus.n118 minus.n117 161.3
R24254 minus.n119 minus.n61 161.3
R24255 minus.n121 minus.n120 161.3
R24256 minus.n60 minus.n59 161.3
R24257 minus.n58 minus.n0 161.3
R24258 minus.n57 minus.n56 161.3
R24259 minus.n55 minus.n54 161.3
R24260 minus.n53 minus.n2 161.3
R24261 minus.n51 minus.n50 161.3
R24262 minus.n49 minus.n3 161.3
R24263 minus.n48 minus.n47 161.3
R24264 minus.n45 minus.n4 161.3
R24265 minus.n44 minus.n43 161.3
R24266 minus.n42 minus.n41 161.3
R24267 minus.n40 minus.n6 161.3
R24268 minus.n39 minus.n38 161.3
R24269 minus.n37 minus.n36 161.3
R24270 minus.n35 minus.n8 161.3
R24271 minus.n33 minus.n32 161.3
R24272 minus.n31 minus.n9 161.3
R24273 minus.n30 minus.n29 161.3
R24274 minus.n27 minus.n10 161.3
R24275 minus.n26 minus.n25 161.3
R24276 minus.n24 minus.n23 161.3
R24277 minus.n22 minus.n12 161.3
R24278 minus.n21 minus.n20 161.3
R24279 minus.n19 minus.n18 161.3
R24280 minus.n17 minus.n14 161.3
R24281 minus.n106 minus.n105 56.5617
R24282 minus.n97 minus.n96 56.5617
R24283 minus.n88 minus.n87 56.5617
R24284 minus.n27 minus.n26 56.5617
R24285 minus.n36 minus.n35 56.5617
R24286 minus.n45 minus.n44 56.5617
R24287 minus.n115 minus.n114 56.5617
R24288 minus.n79 minus.n78 56.5617
R24289 minus.n18 minus.n17 56.5617
R24290 minus.n54 minus.n53 56.5617
R24291 minus.n119 minus.n118 50.2647
R24292 minus.n58 minus.n57 50.2647
R24293 minus.n108 minus.n64 46.3896
R24294 minus.n84 minus.n83 46.3896
R24295 minus.n23 minus.n22 46.3896
R24296 minus.n47 minus.n3 46.3896
R24297 minus.n76 minus.n75 43.1929
R24298 minus.n15 minus.n14 43.1929
R24299 minus.n101 minus.n100 42.5146
R24300 minus.n94 minus.n70 42.5146
R24301 minus.n33 minus.n9 42.5146
R24302 minus.n40 minus.n39 42.5146
R24303 minus.n77 minus.n76 40.6041
R24304 minus.n16 minus.n15 40.6041
R24305 minus.n102 minus.n101 38.6395
R24306 minus.n90 minus.n70 38.6395
R24307 minus.n29 minus.n9 38.6395
R24308 minus.n41 minus.n40 38.6395
R24309 minus.n122 minus.n121 35.4191
R24310 minus.n112 minus.n64 34.7644
R24311 minus.n83 minus.n82 34.7644
R24312 minus.n22 minus.n21 34.7644
R24313 minus.n51 minus.n3 34.7644
R24314 minus.n114 minus.n113 21.8872
R24315 minus.n79 minus.n74 21.8872
R24316 minus.n18 minus.n13 21.8872
R24317 minus.n53 minus.n52 21.8872
R24318 minus.n105 minus.n66 19.9199
R24319 minus.n89 minus.n88 19.9199
R24320 minus.n28 minus.n27 19.9199
R24321 minus.n44 minus.n5 19.9199
R24322 minus.n124 minus.t0 19.8005
R24323 minus.n124 minus.t2 19.8005
R24324 minus.n123 minus.t4 19.8005
R24325 minus.n123 minus.t3 19.8005
R24326 minus.n97 minus.n68 17.9525
R24327 minus.n96 minus.n95 17.9525
R24328 minus.n35 minus.n34 17.9525
R24329 minus.n36 minus.n7 17.9525
R24330 minus.n107 minus.n106 15.9852
R24331 minus.n87 minus.n72 15.9852
R24332 minus.n26 minus.n11 15.9852
R24333 minus.n46 minus.n45 15.9852
R24334 minus.n115 minus.n62 14.0178
R24335 minus.n78 minus.n77 14.0178
R24336 minus.n17 minus.n16 14.0178
R24337 minus.n54 minus.n1 14.0178
R24338 minus.n122 minus.n60 12.1501
R24339 minus minus.n127 11.8706
R24340 minus.n118 minus.n62 10.575
R24341 minus.n57 minus.n1 10.575
R24342 minus.n120 minus.n119 9.49444
R24343 minus.n59 minus.n58 9.49444
R24344 minus.n108 minus.n107 8.60764
R24345 minus.n84 minus.n72 8.60764
R24346 minus.n23 minus.n11 8.60764
R24347 minus.n47 minus.n46 8.60764
R24348 minus.n100 minus.n68 6.6403
R24349 minus.n95 minus.n94 6.6403
R24350 minus.n34 minus.n33 6.6403
R24351 minus.n39 minus.n7 6.6403
R24352 minus.n127 minus.n126 4.80222
R24353 minus.n102 minus.n66 4.67295
R24354 minus.n90 minus.n89 4.67295
R24355 minus.n29 minus.n28 4.67295
R24356 minus.n41 minus.n5 4.67295
R24357 minus.n113 minus.n112 2.7056
R24358 minus.n82 minus.n74 2.7056
R24359 minus.n21 minus.n13 2.7056
R24360 minus.n52 minus.n51 2.7056
R24361 minus.n127 minus.n122 0.972091
R24362 minus.n126 minus.n125 0.716017
R24363 minus.n121 minus.n61 0.189894
R24364 minus.n117 minus.n61 0.189894
R24365 minus.n117 minus.n116 0.189894
R24366 minus.n116 minus.n63 0.189894
R24367 minus.n111 minus.n63 0.189894
R24368 minus.n111 minus.n110 0.189894
R24369 minus.n110 minus.n109 0.189894
R24370 minus.n109 minus.n65 0.189894
R24371 minus.n104 minus.n65 0.189894
R24372 minus.n104 minus.n103 0.189894
R24373 minus.n103 minus.n67 0.189894
R24374 minus.n99 minus.n67 0.189894
R24375 minus.n99 minus.n98 0.189894
R24376 minus.n98 minus.n69 0.189894
R24377 minus.n93 minus.n69 0.189894
R24378 minus.n93 minus.n92 0.189894
R24379 minus.n92 minus.n91 0.189894
R24380 minus.n91 minus.n71 0.189894
R24381 minus.n86 minus.n71 0.189894
R24382 minus.n86 minus.n85 0.189894
R24383 minus.n85 minus.n73 0.189894
R24384 minus.n81 minus.n73 0.189894
R24385 minus.n81 minus.n80 0.189894
R24386 minus.n80 minus.n75 0.189894
R24387 minus.n19 minus.n14 0.189894
R24388 minus.n20 minus.n19 0.189894
R24389 minus.n20 minus.n12 0.189894
R24390 minus.n24 minus.n12 0.189894
R24391 minus.n25 minus.n24 0.189894
R24392 minus.n25 minus.n10 0.189894
R24393 minus.n30 minus.n10 0.189894
R24394 minus.n31 minus.n30 0.189894
R24395 minus.n32 minus.n31 0.189894
R24396 minus.n32 minus.n8 0.189894
R24397 minus.n37 minus.n8 0.189894
R24398 minus.n38 minus.n37 0.189894
R24399 minus.n38 minus.n6 0.189894
R24400 minus.n42 minus.n6 0.189894
R24401 minus.n43 minus.n42 0.189894
R24402 minus.n43 minus.n4 0.189894
R24403 minus.n48 minus.n4 0.189894
R24404 minus.n49 minus.n48 0.189894
R24405 minus.n50 minus.n49 0.189894
R24406 minus.n50 minus.n2 0.189894
R24407 minus.n55 minus.n2 0.189894
R24408 minus.n56 minus.n55 0.189894
R24409 minus.n56 minus.n0 0.189894
R24410 minus.n60 minus.n0 0.189894
R24411 output.n41 output.n15 289.615
R24412 output.n72 output.n46 289.615
R24413 output.n104 output.n78 289.615
R24414 output.n136 output.n110 289.615
R24415 output.n77 output.n45 197.26
R24416 output.n77 output.n76 196.298
R24417 output.n109 output.n108 196.298
R24418 output.n141 output.n140 196.298
R24419 output.n42 output.n41 185
R24420 output.n40 output.n39 185
R24421 output.n19 output.n18 185
R24422 output.n34 output.n33 185
R24423 output.n32 output.n31 185
R24424 output.n23 output.n22 185
R24425 output.n26 output.n25 185
R24426 output.n73 output.n72 185
R24427 output.n71 output.n70 185
R24428 output.n50 output.n49 185
R24429 output.n65 output.n64 185
R24430 output.n63 output.n62 185
R24431 output.n54 output.n53 185
R24432 output.n57 output.n56 185
R24433 output.n105 output.n104 185
R24434 output.n103 output.n102 185
R24435 output.n82 output.n81 185
R24436 output.n97 output.n96 185
R24437 output.n95 output.n94 185
R24438 output.n86 output.n85 185
R24439 output.n89 output.n88 185
R24440 output.n137 output.n136 185
R24441 output.n135 output.n134 185
R24442 output.n114 output.n113 185
R24443 output.n129 output.n128 185
R24444 output.n127 output.n126 185
R24445 output.n118 output.n117 185
R24446 output.n121 output.n120 185
R24447 output.t19 output.n24 147.661
R24448 output.t17 output.n55 147.661
R24449 output.t18 output.n87 147.661
R24450 output.t16 output.n119 147.661
R24451 output.n41 output.n40 104.615
R24452 output.n40 output.n18 104.615
R24453 output.n33 output.n18 104.615
R24454 output.n33 output.n32 104.615
R24455 output.n32 output.n22 104.615
R24456 output.n25 output.n22 104.615
R24457 output.n72 output.n71 104.615
R24458 output.n71 output.n49 104.615
R24459 output.n64 output.n49 104.615
R24460 output.n64 output.n63 104.615
R24461 output.n63 output.n53 104.615
R24462 output.n56 output.n53 104.615
R24463 output.n104 output.n103 104.615
R24464 output.n103 output.n81 104.615
R24465 output.n96 output.n81 104.615
R24466 output.n96 output.n95 104.615
R24467 output.n95 output.n85 104.615
R24468 output.n88 output.n85 104.615
R24469 output.n136 output.n135 104.615
R24470 output.n135 output.n113 104.615
R24471 output.n128 output.n113 104.615
R24472 output.n128 output.n127 104.615
R24473 output.n127 output.n117 104.615
R24474 output.n120 output.n117 104.615
R24475 output.n1 output.t11 77.056
R24476 output.n14 output.t13 76.6694
R24477 output.n1 output.n0 72.7095
R24478 output.n3 output.n2 72.7095
R24479 output.n5 output.n4 72.7095
R24480 output.n7 output.n6 72.7095
R24481 output.n9 output.n8 72.7095
R24482 output.n11 output.n10 72.7095
R24483 output.n13 output.n12 72.7095
R24484 output.n25 output.t19 52.3082
R24485 output.n56 output.t17 52.3082
R24486 output.n88 output.t18 52.3082
R24487 output.n120 output.t16 52.3082
R24488 output.n26 output.n24 15.6674
R24489 output.n57 output.n55 15.6674
R24490 output.n89 output.n87 15.6674
R24491 output.n121 output.n119 15.6674
R24492 output.n27 output.n23 12.8005
R24493 output.n58 output.n54 12.8005
R24494 output.n90 output.n86 12.8005
R24495 output.n122 output.n118 12.8005
R24496 output.n31 output.n30 12.0247
R24497 output.n62 output.n61 12.0247
R24498 output.n94 output.n93 12.0247
R24499 output.n126 output.n125 12.0247
R24500 output.n34 output.n21 11.249
R24501 output.n65 output.n52 11.249
R24502 output.n97 output.n84 11.249
R24503 output.n129 output.n116 11.249
R24504 output.n35 output.n19 10.4732
R24505 output.n66 output.n50 10.4732
R24506 output.n98 output.n82 10.4732
R24507 output.n130 output.n114 10.4732
R24508 output.n39 output.n38 9.69747
R24509 output.n70 output.n69 9.69747
R24510 output.n102 output.n101 9.69747
R24511 output.n134 output.n133 9.69747
R24512 output.n45 output.n44 9.45567
R24513 output.n76 output.n75 9.45567
R24514 output.n108 output.n107 9.45567
R24515 output.n140 output.n139 9.45567
R24516 output.n44 output.n43 9.3005
R24517 output.n17 output.n16 9.3005
R24518 output.n38 output.n37 9.3005
R24519 output.n36 output.n35 9.3005
R24520 output.n21 output.n20 9.3005
R24521 output.n30 output.n29 9.3005
R24522 output.n28 output.n27 9.3005
R24523 output.n75 output.n74 9.3005
R24524 output.n48 output.n47 9.3005
R24525 output.n69 output.n68 9.3005
R24526 output.n67 output.n66 9.3005
R24527 output.n52 output.n51 9.3005
R24528 output.n61 output.n60 9.3005
R24529 output.n59 output.n58 9.3005
R24530 output.n107 output.n106 9.3005
R24531 output.n80 output.n79 9.3005
R24532 output.n101 output.n100 9.3005
R24533 output.n99 output.n98 9.3005
R24534 output.n84 output.n83 9.3005
R24535 output.n93 output.n92 9.3005
R24536 output.n91 output.n90 9.3005
R24537 output.n139 output.n138 9.3005
R24538 output.n112 output.n111 9.3005
R24539 output.n133 output.n132 9.3005
R24540 output.n131 output.n130 9.3005
R24541 output.n116 output.n115 9.3005
R24542 output.n125 output.n124 9.3005
R24543 output.n123 output.n122 9.3005
R24544 output.n42 output.n17 8.92171
R24545 output.n73 output.n48 8.92171
R24546 output.n105 output.n80 8.92171
R24547 output.n137 output.n112 8.92171
R24548 output output.n141 8.15037
R24549 output.n43 output.n15 8.14595
R24550 output.n74 output.n46 8.14595
R24551 output.n106 output.n78 8.14595
R24552 output.n138 output.n110 8.14595
R24553 output.n45 output.n15 5.81868
R24554 output.n76 output.n46 5.81868
R24555 output.n108 output.n78 5.81868
R24556 output.n140 output.n110 5.81868
R24557 output.n43 output.n42 5.04292
R24558 output.n74 output.n73 5.04292
R24559 output.n106 output.n105 5.04292
R24560 output.n138 output.n137 5.04292
R24561 output.n28 output.n24 4.38594
R24562 output.n59 output.n55 4.38594
R24563 output.n91 output.n87 4.38594
R24564 output.n123 output.n119 4.38594
R24565 output.n39 output.n17 4.26717
R24566 output.n70 output.n48 4.26717
R24567 output.n102 output.n80 4.26717
R24568 output.n134 output.n112 4.26717
R24569 output.n0 output.t1 3.9605
R24570 output.n0 output.t6 3.9605
R24571 output.n2 output.t10 3.9605
R24572 output.n2 output.t2 3.9605
R24573 output.n4 output.t4 3.9605
R24574 output.n4 output.t3 3.9605
R24575 output.n6 output.t9 3.9605
R24576 output.n6 output.t12 3.9605
R24577 output.n8 output.t14 3.9605
R24578 output.n8 output.t7 3.9605
R24579 output.n10 output.t8 3.9605
R24580 output.n10 output.t15 3.9605
R24581 output.n12 output.t0 3.9605
R24582 output.n12 output.t5 3.9605
R24583 output.n38 output.n19 3.49141
R24584 output.n69 output.n50 3.49141
R24585 output.n101 output.n82 3.49141
R24586 output.n133 output.n114 3.49141
R24587 output.n35 output.n34 2.71565
R24588 output.n66 output.n65 2.71565
R24589 output.n98 output.n97 2.71565
R24590 output.n130 output.n129 2.71565
R24591 output.n31 output.n21 1.93989
R24592 output.n62 output.n52 1.93989
R24593 output.n94 output.n84 1.93989
R24594 output.n126 output.n116 1.93989
R24595 output.n30 output.n23 1.16414
R24596 output.n61 output.n54 1.16414
R24597 output.n93 output.n86 1.16414
R24598 output.n125 output.n118 1.16414
R24599 output.n141 output.n109 0.962709
R24600 output.n109 output.n77 0.962709
R24601 output.n27 output.n26 0.388379
R24602 output.n58 output.n57 0.388379
R24603 output.n90 output.n89 0.388379
R24604 output.n122 output.n121 0.388379
R24605 output.n14 output.n13 0.387128
R24606 output.n13 output.n11 0.387128
R24607 output.n11 output.n9 0.387128
R24608 output.n9 output.n7 0.387128
R24609 output.n7 output.n5 0.387128
R24610 output.n5 output.n3 0.387128
R24611 output.n3 output.n1 0.387128
R24612 output.n44 output.n16 0.155672
R24613 output.n37 output.n16 0.155672
R24614 output.n37 output.n36 0.155672
R24615 output.n36 output.n20 0.155672
R24616 output.n29 output.n20 0.155672
R24617 output.n29 output.n28 0.155672
R24618 output.n75 output.n47 0.155672
R24619 output.n68 output.n47 0.155672
R24620 output.n68 output.n67 0.155672
R24621 output.n67 output.n51 0.155672
R24622 output.n60 output.n51 0.155672
R24623 output.n60 output.n59 0.155672
R24624 output.n107 output.n79 0.155672
R24625 output.n100 output.n79 0.155672
R24626 output.n100 output.n99 0.155672
R24627 output.n99 output.n83 0.155672
R24628 output.n92 output.n83 0.155672
R24629 output.n92 output.n91 0.155672
R24630 output.n139 output.n111 0.155672
R24631 output.n132 output.n111 0.155672
R24632 output.n132 output.n131 0.155672
R24633 output.n131 output.n115 0.155672
R24634 output.n124 output.n115 0.155672
R24635 output.n124 output.n123 0.155672
R24636 output output.n14 0.126227
C0 output outputibias 2.34152f
C1 vdd output 7.23429f
C2 CSoutput output 6.13571f
C3 CSoutput outputibias 0.032386f
C4 vdd CSoutput 0.140606p
C5 commonsourceibias output 0.006808f
C6 minus diffpairibias 5.39e-19
C7 CSoutput minus 3.03921f
C8 vdd plus 0.096191f
C9 plus diffpairibias 4.4e-19
C10 commonsourceibias outputibias 0.003832f
C11 vdd commonsourceibias 0.004218f
C12 CSoutput plus 0.931998f
C13 commonsourceibias diffpairibias 0.052527f
C14 CSoutput commonsourceibias 45.462303f
C15 minus plus 10.7649f
C16 minus commonsourceibias 0.343793f
C17 plus commonsourceibias 0.290384f
C18 diffpairibias gnd 59.991528f
C19 outputibias gnd 32.465668f
C20 output gnd 15.47879f
C21 commonsourceibias gnd 0.181983p
C22 plus gnd 40.3669f
C23 minus gnd 32.60239f
C24 CSoutput gnd 0.115655p
C25 vdd gnd 0.440142p
C26 output.t11 gnd 0.464308f
C27 output.t1 gnd 0.044422f
C28 output.t6 gnd 0.044422f
C29 output.n0 gnd 0.364624f
C30 output.n1 gnd 0.614102f
C31 output.t10 gnd 0.044422f
C32 output.t2 gnd 0.044422f
C33 output.n2 gnd 0.364624f
C34 output.n3 gnd 0.350265f
C35 output.t4 gnd 0.044422f
C36 output.t3 gnd 0.044422f
C37 output.n4 gnd 0.364624f
C38 output.n5 gnd 0.350265f
C39 output.t9 gnd 0.044422f
C40 output.t12 gnd 0.044422f
C41 output.n6 gnd 0.364624f
C42 output.n7 gnd 0.350265f
C43 output.t14 gnd 0.044422f
C44 output.t7 gnd 0.044422f
C45 output.n8 gnd 0.364624f
C46 output.n9 gnd 0.350265f
C47 output.t8 gnd 0.044422f
C48 output.t15 gnd 0.044422f
C49 output.n10 gnd 0.364624f
C50 output.n11 gnd 0.350265f
C51 output.t0 gnd 0.044422f
C52 output.t5 gnd 0.044422f
C53 output.n12 gnd 0.364624f
C54 output.n13 gnd 0.350265f
C55 output.t13 gnd 0.462979f
C56 output.n14 gnd 0.28994f
C57 output.n15 gnd 0.015803f
C58 output.n16 gnd 0.011243f
C59 output.n17 gnd 0.006041f
C60 output.n18 gnd 0.01428f
C61 output.n19 gnd 0.006397f
C62 output.n20 gnd 0.011243f
C63 output.n21 gnd 0.006041f
C64 output.n22 gnd 0.01428f
C65 output.n23 gnd 0.006397f
C66 output.n24 gnd 0.048111f
C67 output.t19 gnd 0.023274f
C68 output.n25 gnd 0.01071f
C69 output.n26 gnd 0.008435f
C70 output.n27 gnd 0.006041f
C71 output.n28 gnd 0.267512f
C72 output.n29 gnd 0.011243f
C73 output.n30 gnd 0.006041f
C74 output.n31 gnd 0.006397f
C75 output.n32 gnd 0.01428f
C76 output.n33 gnd 0.01428f
C77 output.n34 gnd 0.006397f
C78 output.n35 gnd 0.006041f
C79 output.n36 gnd 0.011243f
C80 output.n37 gnd 0.011243f
C81 output.n38 gnd 0.006041f
C82 output.n39 gnd 0.006397f
C83 output.n40 gnd 0.01428f
C84 output.n41 gnd 0.030913f
C85 output.n42 gnd 0.006397f
C86 output.n43 gnd 0.006041f
C87 output.n44 gnd 0.025987f
C88 output.n45 gnd 0.097665f
C89 output.n46 gnd 0.015803f
C90 output.n47 gnd 0.011243f
C91 output.n48 gnd 0.006041f
C92 output.n49 gnd 0.01428f
C93 output.n50 gnd 0.006397f
C94 output.n51 gnd 0.011243f
C95 output.n52 gnd 0.006041f
C96 output.n53 gnd 0.01428f
C97 output.n54 gnd 0.006397f
C98 output.n55 gnd 0.048111f
C99 output.t17 gnd 0.023274f
C100 output.n56 gnd 0.01071f
C101 output.n57 gnd 0.008435f
C102 output.n58 gnd 0.006041f
C103 output.n59 gnd 0.267512f
C104 output.n60 gnd 0.011243f
C105 output.n61 gnd 0.006041f
C106 output.n62 gnd 0.006397f
C107 output.n63 gnd 0.01428f
C108 output.n64 gnd 0.01428f
C109 output.n65 gnd 0.006397f
C110 output.n66 gnd 0.006041f
C111 output.n67 gnd 0.011243f
C112 output.n68 gnd 0.011243f
C113 output.n69 gnd 0.006041f
C114 output.n70 gnd 0.006397f
C115 output.n71 gnd 0.01428f
C116 output.n72 gnd 0.030913f
C117 output.n73 gnd 0.006397f
C118 output.n74 gnd 0.006041f
C119 output.n75 gnd 0.025987f
C120 output.n76 gnd 0.09306f
C121 output.n77 gnd 1.65264f
C122 output.n78 gnd 0.015803f
C123 output.n79 gnd 0.011243f
C124 output.n80 gnd 0.006041f
C125 output.n81 gnd 0.01428f
C126 output.n82 gnd 0.006397f
C127 output.n83 gnd 0.011243f
C128 output.n84 gnd 0.006041f
C129 output.n85 gnd 0.01428f
C130 output.n86 gnd 0.006397f
C131 output.n87 gnd 0.048111f
C132 output.t18 gnd 0.023274f
C133 output.n88 gnd 0.01071f
C134 output.n89 gnd 0.008435f
C135 output.n90 gnd 0.006041f
C136 output.n91 gnd 0.267512f
C137 output.n92 gnd 0.011243f
C138 output.n93 gnd 0.006041f
C139 output.n94 gnd 0.006397f
C140 output.n95 gnd 0.01428f
C141 output.n96 gnd 0.01428f
C142 output.n97 gnd 0.006397f
C143 output.n98 gnd 0.006041f
C144 output.n99 gnd 0.011243f
C145 output.n100 gnd 0.011243f
C146 output.n101 gnd 0.006041f
C147 output.n102 gnd 0.006397f
C148 output.n103 gnd 0.01428f
C149 output.n104 gnd 0.030913f
C150 output.n105 gnd 0.006397f
C151 output.n106 gnd 0.006041f
C152 output.n107 gnd 0.025987f
C153 output.n108 gnd 0.09306f
C154 output.n109 gnd 0.713089f
C155 output.n110 gnd 0.015803f
C156 output.n111 gnd 0.011243f
C157 output.n112 gnd 0.006041f
C158 output.n113 gnd 0.01428f
C159 output.n114 gnd 0.006397f
C160 output.n115 gnd 0.011243f
C161 output.n116 gnd 0.006041f
C162 output.n117 gnd 0.01428f
C163 output.n118 gnd 0.006397f
C164 output.n119 gnd 0.048111f
C165 output.t16 gnd 0.023274f
C166 output.n120 gnd 0.01071f
C167 output.n121 gnd 0.008435f
C168 output.n122 gnd 0.006041f
C169 output.n123 gnd 0.267512f
C170 output.n124 gnd 0.011243f
C171 output.n125 gnd 0.006041f
C172 output.n126 gnd 0.006397f
C173 output.n127 gnd 0.01428f
C174 output.n128 gnd 0.01428f
C175 output.n129 gnd 0.006397f
C176 output.n130 gnd 0.006041f
C177 output.n131 gnd 0.011243f
C178 output.n132 gnd 0.011243f
C179 output.n133 gnd 0.006041f
C180 output.n134 gnd 0.006397f
C181 output.n135 gnd 0.01428f
C182 output.n136 gnd 0.030913f
C183 output.n137 gnd 0.006397f
C184 output.n138 gnd 0.006041f
C185 output.n139 gnd 0.025987f
C186 output.n140 gnd 0.09306f
C187 output.n141 gnd 1.67353f
C188 minus.n0 gnd 0.030269f
C189 minus.t13 gnd 0.508973f
C190 minus.n1 gnd 0.205851f
C191 minus.n2 gnd 0.030269f
C192 minus.t11 gnd 0.508973f
C193 minus.n3 gnd 0.025866f
C194 minus.n4 gnd 0.030269f
C195 minus.t17 gnd 0.508973f
C196 minus.t24 gnd 0.508973f
C197 minus.n5 gnd 0.205851f
C198 minus.n6 gnd 0.030269f
C199 minus.t21 gnd 0.508973f
C200 minus.n7 gnd 0.205851f
C201 minus.n8 gnd 0.030269f
C202 minus.t27 gnd 0.508973f
C203 minus.n9 gnd 0.024602f
C204 minus.n10 gnd 0.030269f
C205 minus.t26 gnd 0.508973f
C206 minus.t5 gnd 0.508973f
C207 minus.n11 gnd 0.205851f
C208 minus.n12 gnd 0.030269f
C209 minus.t9 gnd 0.508973f
C210 minus.n13 gnd 0.205851f
C211 minus.n14 gnd 0.128459f
C212 minus.t14 gnd 0.508973f
C213 minus.t20 gnd 0.569378f
C214 minus.n15 gnd 0.240661f
C215 minus.n16 gnd 0.235738f
C216 minus.n17 gnd 0.038785f
C217 minus.n18 gnd 0.034253f
C218 minus.n19 gnd 0.030269f
C219 minus.n20 gnd 0.030269f
C220 minus.n21 gnd 0.036172f
C221 minus.n22 gnd 0.025866f
C222 minus.n23 gnd 0.039422f
C223 minus.n24 gnd 0.030269f
C224 minus.n25 gnd 0.030269f
C225 minus.n26 gnd 0.037652f
C226 minus.n27 gnd 0.035386f
C227 minus.n28 gnd 0.205851f
C228 minus.n29 gnd 0.037917f
C229 minus.n30 gnd 0.030269f
C230 minus.n31 gnd 0.030269f
C231 minus.n32 gnd 0.030269f
C232 minus.n33 gnd 0.03894f
C233 minus.n34 gnd 0.205851f
C234 minus.n35 gnd 0.036519f
C235 minus.n36 gnd 0.036519f
C236 minus.n37 gnd 0.030269f
C237 minus.n38 gnd 0.030269f
C238 minus.n39 gnd 0.03894f
C239 minus.n40 gnd 0.024602f
C240 minus.n41 gnd 0.037917f
C241 minus.n42 gnd 0.030269f
C242 minus.n43 gnd 0.030269f
C243 minus.n44 gnd 0.035386f
C244 minus.n45 gnd 0.037652f
C245 minus.n46 gnd 0.205851f
C246 minus.n47 gnd 0.039422f
C247 minus.n48 gnd 0.030269f
C248 minus.n49 gnd 0.030269f
C249 minus.n50 gnd 0.030269f
C250 minus.n51 gnd 0.036172f
C251 minus.n52 gnd 0.205851f
C252 minus.n53 gnd 0.034253f
C253 minus.n54 gnd 0.038785f
C254 minus.n55 gnd 0.030269f
C255 minus.n56 gnd 0.030269f
C256 minus.n57 gnd 0.039487f
C257 minus.n58 gnd 0.011001f
C258 minus.t10 gnd 0.550454f
C259 minus.n59 gnd 0.238341f
C260 minus.n60 gnd 0.354592f
C261 minus.n61 gnd 0.030269f
C262 minus.t8 gnd 0.550454f
C263 minus.t12 gnd 0.508973f
C264 minus.n62 gnd 0.205851f
C265 minus.n63 gnd 0.030269f
C266 minus.t18 gnd 0.508973f
C267 minus.n64 gnd 0.025866f
C268 minus.n65 gnd 0.030269f
C269 minus.t25 gnd 0.508973f
C270 minus.t22 gnd 0.508973f
C271 minus.n66 gnd 0.205851f
C272 minus.n67 gnd 0.030269f
C273 minus.t19 gnd 0.508973f
C274 minus.n68 gnd 0.205851f
C275 minus.n69 gnd 0.030269f
C276 minus.t7 gnd 0.508973f
C277 minus.n70 gnd 0.024602f
C278 minus.n71 gnd 0.030269f
C279 minus.t6 gnd 0.508973f
C280 minus.t16 gnd 0.508973f
C281 minus.n72 gnd 0.205851f
C282 minus.n73 gnd 0.030269f
C283 minus.t15 gnd 0.508973f
C284 minus.n74 gnd 0.205851f
C285 minus.n75 gnd 0.128459f
C286 minus.t23 gnd 0.508973f
C287 minus.t28 gnd 0.569378f
C288 minus.n76 gnd 0.240661f
C289 minus.n77 gnd 0.235738f
C290 minus.n78 gnd 0.038785f
C291 minus.n79 gnd 0.034253f
C292 minus.n80 gnd 0.030269f
C293 minus.n81 gnd 0.030269f
C294 minus.n82 gnd 0.036172f
C295 minus.n83 gnd 0.025866f
C296 minus.n84 gnd 0.039422f
C297 minus.n85 gnd 0.030269f
C298 minus.n86 gnd 0.030269f
C299 minus.n87 gnd 0.037652f
C300 minus.n88 gnd 0.035386f
C301 minus.n89 gnd 0.205851f
C302 minus.n90 gnd 0.037917f
C303 minus.n91 gnd 0.030269f
C304 minus.n92 gnd 0.030269f
C305 minus.n93 gnd 0.030269f
C306 minus.n94 gnd 0.03894f
C307 minus.n95 gnd 0.205851f
C308 minus.n96 gnd 0.036519f
C309 minus.n97 gnd 0.036519f
C310 minus.n98 gnd 0.030269f
C311 minus.n99 gnd 0.030269f
C312 minus.n100 gnd 0.03894f
C313 minus.n101 gnd 0.024602f
C314 minus.n102 gnd 0.037917f
C315 minus.n103 gnd 0.030269f
C316 minus.n104 gnd 0.030269f
C317 minus.n105 gnd 0.035386f
C318 minus.n106 gnd 0.037652f
C319 minus.n107 gnd 0.205851f
C320 minus.n108 gnd 0.039422f
C321 minus.n109 gnd 0.030269f
C322 minus.n110 gnd 0.030269f
C323 minus.n111 gnd 0.030269f
C324 minus.n112 gnd 0.036172f
C325 minus.n113 gnd 0.205851f
C326 minus.n114 gnd 0.034253f
C327 minus.n115 gnd 0.038785f
C328 minus.n116 gnd 0.030269f
C329 minus.n117 gnd 0.030269f
C330 minus.n118 gnd 0.039487f
C331 minus.n119 gnd 0.011001f
C332 minus.n120 gnd 0.238341f
C333 minus.n121 gnd 1.10421f
C334 minus.n122 gnd 1.622f
C335 minus.t4 gnd 0.009331f
C336 minus.t3 gnd 0.009331f
C337 minus.n123 gnd 0.030683f
C338 minus.t0 gnd 0.009331f
C339 minus.t2 gnd 0.009331f
C340 minus.n124 gnd 0.030263f
C341 minus.n125 gnd 0.258277f
C342 minus.t1 gnd 0.051936f
C343 minus.n126 gnd 0.140939f
C344 minus.n127 gnd 2.12621f
C345 commonsourceibias.n0 gnd 0.010724f
C346 commonsourceibias.t115 gnd 0.162395f
C347 commonsourceibias.t136 gnd 0.150157f
C348 commonsourceibias.n1 gnd 0.007823f
C349 commonsourceibias.n2 gnd 0.008037f
C350 commonsourceibias.t151 gnd 0.150157f
C351 commonsourceibias.n3 gnd 0.01034f
C352 commonsourceibias.n4 gnd 0.008037f
C353 commonsourceibias.t105 gnd 0.150157f
C354 commonsourceibias.n5 gnd 0.059912f
C355 commonsourceibias.t126 gnd 0.150157f
C356 commonsourceibias.n6 gnd 0.007578f
C357 commonsourceibias.n7 gnd 0.008037f
C358 commonsourceibias.t144 gnd 0.150157f
C359 commonsourceibias.n8 gnd 0.010186f
C360 commonsourceibias.n9 gnd 0.008037f
C361 commonsourceibias.t98 gnd 0.150157f
C362 commonsourceibias.n10 gnd 0.059912f
C363 commonsourceibias.t94 gnd 0.150157f
C364 commonsourceibias.n11 gnd 0.007361f
C365 commonsourceibias.n12 gnd 0.008037f
C366 commonsourceibias.t135 gnd 0.150157f
C367 commonsourceibias.n13 gnd 0.010015f
C368 commonsourceibias.n14 gnd 0.010724f
C369 commonsourceibias.t74 gnd 0.162395f
C370 commonsourceibias.t20 gnd 0.150157f
C371 commonsourceibias.n15 gnd 0.007823f
C372 commonsourceibias.n16 gnd 0.008037f
C373 commonsourceibias.t50 gnd 0.150157f
C374 commonsourceibias.n17 gnd 0.01034f
C375 commonsourceibias.n18 gnd 0.008037f
C376 commonsourceibias.t8 gnd 0.150157f
C377 commonsourceibias.n19 gnd 0.059912f
C378 commonsourceibias.t36 gnd 0.150157f
C379 commonsourceibias.n20 gnd 0.007578f
C380 commonsourceibias.n21 gnd 0.008037f
C381 commonsourceibias.t76 gnd 0.150157f
C382 commonsourceibias.n22 gnd 0.010186f
C383 commonsourceibias.n23 gnd 0.008037f
C384 commonsourceibias.t24 gnd 0.150157f
C385 commonsourceibias.n24 gnd 0.059912f
C386 commonsourceibias.t34 gnd 0.150157f
C387 commonsourceibias.n25 gnd 0.007361f
C388 commonsourceibias.n26 gnd 0.008037f
C389 commonsourceibias.t10 gnd 0.150157f
C390 commonsourceibias.n27 gnd 0.010015f
C391 commonsourceibias.n28 gnd 0.008037f
C392 commonsourceibias.t40 gnd 0.150157f
C393 commonsourceibias.n29 gnd 0.059912f
C394 commonsourceibias.t56 gnd 0.150157f
C395 commonsourceibias.n30 gnd 0.007172f
C396 commonsourceibias.n31 gnd 0.008037f
C397 commonsourceibias.t26 gnd 0.150157f
C398 commonsourceibias.n32 gnd 0.009825f
C399 commonsourceibias.n33 gnd 0.008037f
C400 commonsourceibias.t38 gnd 0.150157f
C401 commonsourceibias.n34 gnd 0.059912f
C402 commonsourceibias.t70 gnd 0.150157f
C403 commonsourceibias.n35 gnd 0.007008f
C404 commonsourceibias.n36 gnd 0.008037f
C405 commonsourceibias.t18 gnd 0.150157f
C406 commonsourceibias.n37 gnd 0.009613f
C407 commonsourceibias.n38 gnd 0.008037f
C408 commonsourceibias.t22 gnd 0.150157f
C409 commonsourceibias.n39 gnd 0.059912f
C410 commonsourceibias.t54 gnd 0.150157f
C411 commonsourceibias.n40 gnd 0.006868f
C412 commonsourceibias.n41 gnd 0.008037f
C413 commonsourceibias.t4 gnd 0.150157f
C414 commonsourceibias.n42 gnd 0.009378f
C415 commonsourceibias.t78 gnd 0.166947f
C416 commonsourceibias.t46 gnd 0.150157f
C417 commonsourceibias.n43 gnd 0.065449f
C418 commonsourceibias.n44 gnd 0.071822f
C419 commonsourceibias.n45 gnd 0.033327f
C420 commonsourceibias.n46 gnd 0.008037f
C421 commonsourceibias.n47 gnd 0.007823f
C422 commonsourceibias.n48 gnd 0.01121f
C423 commonsourceibias.n49 gnd 0.059912f
C424 commonsourceibias.n50 gnd 0.011203f
C425 commonsourceibias.n51 gnd 0.008037f
C426 commonsourceibias.n52 gnd 0.008037f
C427 commonsourceibias.n53 gnd 0.008037f
C428 commonsourceibias.n54 gnd 0.01034f
C429 commonsourceibias.n55 gnd 0.059912f
C430 commonsourceibias.n56 gnd 0.010583f
C431 commonsourceibias.n57 gnd 0.010282f
C432 commonsourceibias.n58 gnd 0.008037f
C433 commonsourceibias.n59 gnd 0.008037f
C434 commonsourceibias.n60 gnd 0.008037f
C435 commonsourceibias.n61 gnd 0.007578f
C436 commonsourceibias.n62 gnd 0.01122f
C437 commonsourceibias.n63 gnd 0.059912f
C438 commonsourceibias.n64 gnd 0.011217f
C439 commonsourceibias.n65 gnd 0.008037f
C440 commonsourceibias.n66 gnd 0.008037f
C441 commonsourceibias.n67 gnd 0.008037f
C442 commonsourceibias.n68 gnd 0.010186f
C443 commonsourceibias.n69 gnd 0.059912f
C444 commonsourceibias.n70 gnd 0.010507f
C445 commonsourceibias.n71 gnd 0.010357f
C446 commonsourceibias.n72 gnd 0.008037f
C447 commonsourceibias.n73 gnd 0.008037f
C448 commonsourceibias.n74 gnd 0.008037f
C449 commonsourceibias.n75 gnd 0.007361f
C450 commonsourceibias.n76 gnd 0.011225f
C451 commonsourceibias.n77 gnd 0.059912f
C452 commonsourceibias.n78 gnd 0.011224f
C453 commonsourceibias.n79 gnd 0.008037f
C454 commonsourceibias.n80 gnd 0.008037f
C455 commonsourceibias.n81 gnd 0.008037f
C456 commonsourceibias.n82 gnd 0.010015f
C457 commonsourceibias.n83 gnd 0.059912f
C458 commonsourceibias.n84 gnd 0.010432f
C459 commonsourceibias.n85 gnd 0.010432f
C460 commonsourceibias.n86 gnd 0.008037f
C461 commonsourceibias.n87 gnd 0.008037f
C462 commonsourceibias.n88 gnd 0.008037f
C463 commonsourceibias.n89 gnd 0.007172f
C464 commonsourceibias.n90 gnd 0.011224f
C465 commonsourceibias.n91 gnd 0.059912f
C466 commonsourceibias.n92 gnd 0.011225f
C467 commonsourceibias.n93 gnd 0.008037f
C468 commonsourceibias.n94 gnd 0.008037f
C469 commonsourceibias.n95 gnd 0.008037f
C470 commonsourceibias.n96 gnd 0.009825f
C471 commonsourceibias.n97 gnd 0.059912f
C472 commonsourceibias.n98 gnd 0.010357f
C473 commonsourceibias.n99 gnd 0.010507f
C474 commonsourceibias.n100 gnd 0.008037f
C475 commonsourceibias.n101 gnd 0.008037f
C476 commonsourceibias.n102 gnd 0.008037f
C477 commonsourceibias.n103 gnd 0.007008f
C478 commonsourceibias.n104 gnd 0.011217f
C479 commonsourceibias.n105 gnd 0.059912f
C480 commonsourceibias.n106 gnd 0.01122f
C481 commonsourceibias.n107 gnd 0.008037f
C482 commonsourceibias.n108 gnd 0.008037f
C483 commonsourceibias.n109 gnd 0.008037f
C484 commonsourceibias.n110 gnd 0.009613f
C485 commonsourceibias.n111 gnd 0.059912f
C486 commonsourceibias.n112 gnd 0.010282f
C487 commonsourceibias.n113 gnd 0.010583f
C488 commonsourceibias.n114 gnd 0.008037f
C489 commonsourceibias.n115 gnd 0.008037f
C490 commonsourceibias.n116 gnd 0.008037f
C491 commonsourceibias.n117 gnd 0.006868f
C492 commonsourceibias.n118 gnd 0.011203f
C493 commonsourceibias.n119 gnd 0.059912f
C494 commonsourceibias.n120 gnd 0.01121f
C495 commonsourceibias.n121 gnd 0.008037f
C496 commonsourceibias.n122 gnd 0.008037f
C497 commonsourceibias.n123 gnd 0.008037f
C498 commonsourceibias.n124 gnd 0.009378f
C499 commonsourceibias.n125 gnd 0.059912f
C500 commonsourceibias.n126 gnd 0.009861f
C501 commonsourceibias.n127 gnd 0.07189f
C502 commonsourceibias.n128 gnd 0.080075f
C503 commonsourceibias.t75 gnd 0.017343f
C504 commonsourceibias.t21 gnd 0.017343f
C505 commonsourceibias.n129 gnd 0.15325f
C506 commonsourceibias.n130 gnd 0.132562f
C507 commonsourceibias.t51 gnd 0.017343f
C508 commonsourceibias.t9 gnd 0.017343f
C509 commonsourceibias.n131 gnd 0.15325f
C510 commonsourceibias.n132 gnd 0.070394f
C511 commonsourceibias.t37 gnd 0.017343f
C512 commonsourceibias.t77 gnd 0.017343f
C513 commonsourceibias.n133 gnd 0.15325f
C514 commonsourceibias.n134 gnd 0.070394f
C515 commonsourceibias.t25 gnd 0.017343f
C516 commonsourceibias.t35 gnd 0.017343f
C517 commonsourceibias.n135 gnd 0.15325f
C518 commonsourceibias.n136 gnd 0.070394f
C519 commonsourceibias.t11 gnd 0.017343f
C520 commonsourceibias.t41 gnd 0.017343f
C521 commonsourceibias.n137 gnd 0.15325f
C522 commonsourceibias.n138 gnd 0.058811f
C523 commonsourceibias.t47 gnd 0.017343f
C524 commonsourceibias.t79 gnd 0.017343f
C525 commonsourceibias.n139 gnd 0.153763f
C526 commonsourceibias.t55 gnd 0.017343f
C527 commonsourceibias.t5 gnd 0.017343f
C528 commonsourceibias.n140 gnd 0.15325f
C529 commonsourceibias.n141 gnd 0.1428f
C530 commonsourceibias.t19 gnd 0.017343f
C531 commonsourceibias.t23 gnd 0.017343f
C532 commonsourceibias.n142 gnd 0.15325f
C533 commonsourceibias.n143 gnd 0.070394f
C534 commonsourceibias.t39 gnd 0.017343f
C535 commonsourceibias.t71 gnd 0.017343f
C536 commonsourceibias.n144 gnd 0.15325f
C537 commonsourceibias.n145 gnd 0.070394f
C538 commonsourceibias.t57 gnd 0.017343f
C539 commonsourceibias.t27 gnd 0.017343f
C540 commonsourceibias.n146 gnd 0.15325f
C541 commonsourceibias.n147 gnd 0.058811f
C542 commonsourceibias.n148 gnd 0.071213f
C543 commonsourceibias.n149 gnd 0.052016f
C544 commonsourceibias.t153 gnd 0.150157f
C545 commonsourceibias.n150 gnd 0.059912f
C546 commonsourceibias.t88 gnd 0.150157f
C547 commonsourceibias.n151 gnd 0.059912f
C548 commonsourceibias.n152 gnd 0.008037f
C549 commonsourceibias.t125 gnd 0.150157f
C550 commonsourceibias.n153 gnd 0.059912f
C551 commonsourceibias.n154 gnd 0.008037f
C552 commonsourceibias.t120 gnd 0.150157f
C553 commonsourceibias.n155 gnd 0.059912f
C554 commonsourceibias.n156 gnd 0.008037f
C555 commonsourceibias.t139 gnd 0.150157f
C556 commonsourceibias.n157 gnd 0.007008f
C557 commonsourceibias.n158 gnd 0.008037f
C558 commonsourceibias.t112 gnd 0.150157f
C559 commonsourceibias.n159 gnd 0.009613f
C560 commonsourceibias.n160 gnd 0.008037f
C561 commonsourceibias.t107 gnd 0.150157f
C562 commonsourceibias.n161 gnd 0.059912f
C563 commonsourceibias.t127 gnd 0.150157f
C564 commonsourceibias.n162 gnd 0.006868f
C565 commonsourceibias.n163 gnd 0.008037f
C566 commonsourceibias.t146 gnd 0.150157f
C567 commonsourceibias.n164 gnd 0.009378f
C568 commonsourceibias.t117 gnd 0.166947f
C569 commonsourceibias.t99 gnd 0.150157f
C570 commonsourceibias.n165 gnd 0.065449f
C571 commonsourceibias.n166 gnd 0.071822f
C572 commonsourceibias.n167 gnd 0.033327f
C573 commonsourceibias.n168 gnd 0.008037f
C574 commonsourceibias.n169 gnd 0.007823f
C575 commonsourceibias.n170 gnd 0.01121f
C576 commonsourceibias.n171 gnd 0.059912f
C577 commonsourceibias.n172 gnd 0.011203f
C578 commonsourceibias.n173 gnd 0.008037f
C579 commonsourceibias.n174 gnd 0.008037f
C580 commonsourceibias.n175 gnd 0.008037f
C581 commonsourceibias.n176 gnd 0.01034f
C582 commonsourceibias.n177 gnd 0.059912f
C583 commonsourceibias.n178 gnd 0.010583f
C584 commonsourceibias.n179 gnd 0.010282f
C585 commonsourceibias.n180 gnd 0.008037f
C586 commonsourceibias.n181 gnd 0.008037f
C587 commonsourceibias.n182 gnd 0.008037f
C588 commonsourceibias.n183 gnd 0.007578f
C589 commonsourceibias.n184 gnd 0.01122f
C590 commonsourceibias.n185 gnd 0.059912f
C591 commonsourceibias.n186 gnd 0.011217f
C592 commonsourceibias.n187 gnd 0.008037f
C593 commonsourceibias.n188 gnd 0.008037f
C594 commonsourceibias.n189 gnd 0.008037f
C595 commonsourceibias.n190 gnd 0.010186f
C596 commonsourceibias.n191 gnd 0.059912f
C597 commonsourceibias.n192 gnd 0.010507f
C598 commonsourceibias.n193 gnd 0.010357f
C599 commonsourceibias.n194 gnd 0.008037f
C600 commonsourceibias.n195 gnd 0.008037f
C601 commonsourceibias.n196 gnd 0.009825f
C602 commonsourceibias.n197 gnd 0.007361f
C603 commonsourceibias.n198 gnd 0.011225f
C604 commonsourceibias.n199 gnd 0.008037f
C605 commonsourceibias.n200 gnd 0.008037f
C606 commonsourceibias.n201 gnd 0.011224f
C607 commonsourceibias.n202 gnd 0.007172f
C608 commonsourceibias.n203 gnd 0.010015f
C609 commonsourceibias.n204 gnd 0.008037f
C610 commonsourceibias.n205 gnd 0.007021f
C611 commonsourceibias.n206 gnd 0.010432f
C612 commonsourceibias.n207 gnd 0.010432f
C613 commonsourceibias.n208 gnd 0.007021f
C614 commonsourceibias.n209 gnd 0.008037f
C615 commonsourceibias.n210 gnd 0.008037f
C616 commonsourceibias.n211 gnd 0.007172f
C617 commonsourceibias.n212 gnd 0.011224f
C618 commonsourceibias.n213 gnd 0.059912f
C619 commonsourceibias.n214 gnd 0.011225f
C620 commonsourceibias.n215 gnd 0.008037f
C621 commonsourceibias.n216 gnd 0.008037f
C622 commonsourceibias.n217 gnd 0.008037f
C623 commonsourceibias.n218 gnd 0.009825f
C624 commonsourceibias.n219 gnd 0.059912f
C625 commonsourceibias.n220 gnd 0.010357f
C626 commonsourceibias.n221 gnd 0.010507f
C627 commonsourceibias.n222 gnd 0.008037f
C628 commonsourceibias.n223 gnd 0.008037f
C629 commonsourceibias.n224 gnd 0.008037f
C630 commonsourceibias.n225 gnd 0.007008f
C631 commonsourceibias.n226 gnd 0.011217f
C632 commonsourceibias.n227 gnd 0.059912f
C633 commonsourceibias.n228 gnd 0.01122f
C634 commonsourceibias.n229 gnd 0.008037f
C635 commonsourceibias.n230 gnd 0.008037f
C636 commonsourceibias.n231 gnd 0.008037f
C637 commonsourceibias.n232 gnd 0.009613f
C638 commonsourceibias.n233 gnd 0.059912f
C639 commonsourceibias.n234 gnd 0.010282f
C640 commonsourceibias.n235 gnd 0.010583f
C641 commonsourceibias.n236 gnd 0.008037f
C642 commonsourceibias.n237 gnd 0.008037f
C643 commonsourceibias.n238 gnd 0.008037f
C644 commonsourceibias.n239 gnd 0.006868f
C645 commonsourceibias.n240 gnd 0.011203f
C646 commonsourceibias.n241 gnd 0.059912f
C647 commonsourceibias.n242 gnd 0.01121f
C648 commonsourceibias.n243 gnd 0.008037f
C649 commonsourceibias.n244 gnd 0.008037f
C650 commonsourceibias.n245 gnd 0.008037f
C651 commonsourceibias.n246 gnd 0.009378f
C652 commonsourceibias.n247 gnd 0.059912f
C653 commonsourceibias.n248 gnd 0.009861f
C654 commonsourceibias.n249 gnd 0.07189f
C655 commonsourceibias.n250 gnd 0.04697f
C656 commonsourceibias.n251 gnd 0.010724f
C657 commonsourceibias.t119 gnd 0.150157f
C658 commonsourceibias.n252 gnd 0.007823f
C659 commonsourceibias.n253 gnd 0.008037f
C660 commonsourceibias.t137 gnd 0.150157f
C661 commonsourceibias.n254 gnd 0.01034f
C662 commonsourceibias.n255 gnd 0.008037f
C663 commonsourceibias.t92 gnd 0.150157f
C664 commonsourceibias.n256 gnd 0.059912f
C665 commonsourceibias.t109 gnd 0.150157f
C666 commonsourceibias.n257 gnd 0.007578f
C667 commonsourceibias.n258 gnd 0.008037f
C668 commonsourceibias.t128 gnd 0.150157f
C669 commonsourceibias.n259 gnd 0.010186f
C670 commonsourceibias.n260 gnd 0.008037f
C671 commonsourceibias.t86 gnd 0.150157f
C672 commonsourceibias.n261 gnd 0.059912f
C673 commonsourceibias.t83 gnd 0.150157f
C674 commonsourceibias.n262 gnd 0.007361f
C675 commonsourceibias.n263 gnd 0.008037f
C676 commonsourceibias.t118 gnd 0.150157f
C677 commonsourceibias.n264 gnd 0.010015f
C678 commonsourceibias.n265 gnd 0.008037f
C679 commonsourceibias.t138 gnd 0.150157f
C680 commonsourceibias.n266 gnd 0.059912f
C681 commonsourceibias.t159 gnd 0.150157f
C682 commonsourceibias.n267 gnd 0.007172f
C683 commonsourceibias.n268 gnd 0.008037f
C684 commonsourceibias.t108 gnd 0.150157f
C685 commonsourceibias.n269 gnd 0.009825f
C686 commonsourceibias.n270 gnd 0.008037f
C687 commonsourceibias.t102 gnd 0.150157f
C688 commonsourceibias.n271 gnd 0.059912f
C689 commonsourceibias.t121 gnd 0.150157f
C690 commonsourceibias.n272 gnd 0.007008f
C691 commonsourceibias.n273 gnd 0.008037f
C692 commonsourceibias.t95 gnd 0.150157f
C693 commonsourceibias.n274 gnd 0.009613f
C694 commonsourceibias.n275 gnd 0.008037f
C695 commonsourceibias.t93 gnd 0.150157f
C696 commonsourceibias.n276 gnd 0.059912f
C697 commonsourceibias.t110 gnd 0.150157f
C698 commonsourceibias.n277 gnd 0.006868f
C699 commonsourceibias.n278 gnd 0.008037f
C700 commonsourceibias.t129 gnd 0.150157f
C701 commonsourceibias.n279 gnd 0.009378f
C702 commonsourceibias.t101 gnd 0.166947f
C703 commonsourceibias.t87 gnd 0.150157f
C704 commonsourceibias.n280 gnd 0.065449f
C705 commonsourceibias.n281 gnd 0.071822f
C706 commonsourceibias.n282 gnd 0.033327f
C707 commonsourceibias.n283 gnd 0.008037f
C708 commonsourceibias.n284 gnd 0.007823f
C709 commonsourceibias.n285 gnd 0.01121f
C710 commonsourceibias.n286 gnd 0.059912f
C711 commonsourceibias.n287 gnd 0.011203f
C712 commonsourceibias.n288 gnd 0.008037f
C713 commonsourceibias.n289 gnd 0.008037f
C714 commonsourceibias.n290 gnd 0.008037f
C715 commonsourceibias.n291 gnd 0.01034f
C716 commonsourceibias.n292 gnd 0.059912f
C717 commonsourceibias.n293 gnd 0.010583f
C718 commonsourceibias.n294 gnd 0.010282f
C719 commonsourceibias.n295 gnd 0.008037f
C720 commonsourceibias.n296 gnd 0.008037f
C721 commonsourceibias.n297 gnd 0.008037f
C722 commonsourceibias.n298 gnd 0.007578f
C723 commonsourceibias.n299 gnd 0.01122f
C724 commonsourceibias.n300 gnd 0.059912f
C725 commonsourceibias.n301 gnd 0.011217f
C726 commonsourceibias.n302 gnd 0.008037f
C727 commonsourceibias.n303 gnd 0.008037f
C728 commonsourceibias.n304 gnd 0.008037f
C729 commonsourceibias.n305 gnd 0.010186f
C730 commonsourceibias.n306 gnd 0.059912f
C731 commonsourceibias.n307 gnd 0.010507f
C732 commonsourceibias.n308 gnd 0.010357f
C733 commonsourceibias.n309 gnd 0.008037f
C734 commonsourceibias.n310 gnd 0.008037f
C735 commonsourceibias.n311 gnd 0.008037f
C736 commonsourceibias.n312 gnd 0.007361f
C737 commonsourceibias.n313 gnd 0.011225f
C738 commonsourceibias.n314 gnd 0.059912f
C739 commonsourceibias.n315 gnd 0.011224f
C740 commonsourceibias.n316 gnd 0.008037f
C741 commonsourceibias.n317 gnd 0.008037f
C742 commonsourceibias.n318 gnd 0.008037f
C743 commonsourceibias.n319 gnd 0.010015f
C744 commonsourceibias.n320 gnd 0.059912f
C745 commonsourceibias.n321 gnd 0.010432f
C746 commonsourceibias.n322 gnd 0.010432f
C747 commonsourceibias.n323 gnd 0.008037f
C748 commonsourceibias.n324 gnd 0.008037f
C749 commonsourceibias.n325 gnd 0.008037f
C750 commonsourceibias.n326 gnd 0.007172f
C751 commonsourceibias.n327 gnd 0.011224f
C752 commonsourceibias.n328 gnd 0.059912f
C753 commonsourceibias.n329 gnd 0.011225f
C754 commonsourceibias.n330 gnd 0.008037f
C755 commonsourceibias.n331 gnd 0.008037f
C756 commonsourceibias.n332 gnd 0.008037f
C757 commonsourceibias.n333 gnd 0.009825f
C758 commonsourceibias.n334 gnd 0.059912f
C759 commonsourceibias.n335 gnd 0.010357f
C760 commonsourceibias.n336 gnd 0.010507f
C761 commonsourceibias.n337 gnd 0.008037f
C762 commonsourceibias.n338 gnd 0.008037f
C763 commonsourceibias.n339 gnd 0.008037f
C764 commonsourceibias.n340 gnd 0.007008f
C765 commonsourceibias.n341 gnd 0.011217f
C766 commonsourceibias.n342 gnd 0.059912f
C767 commonsourceibias.n343 gnd 0.01122f
C768 commonsourceibias.n344 gnd 0.008037f
C769 commonsourceibias.n345 gnd 0.008037f
C770 commonsourceibias.n346 gnd 0.008037f
C771 commonsourceibias.n347 gnd 0.009613f
C772 commonsourceibias.n348 gnd 0.059912f
C773 commonsourceibias.n349 gnd 0.010282f
C774 commonsourceibias.n350 gnd 0.010583f
C775 commonsourceibias.n351 gnd 0.008037f
C776 commonsourceibias.n352 gnd 0.008037f
C777 commonsourceibias.n353 gnd 0.008037f
C778 commonsourceibias.n354 gnd 0.006868f
C779 commonsourceibias.n355 gnd 0.011203f
C780 commonsourceibias.n356 gnd 0.059912f
C781 commonsourceibias.n357 gnd 0.01121f
C782 commonsourceibias.n358 gnd 0.008037f
C783 commonsourceibias.n359 gnd 0.008037f
C784 commonsourceibias.n360 gnd 0.008037f
C785 commonsourceibias.n361 gnd 0.009378f
C786 commonsourceibias.n362 gnd 0.059912f
C787 commonsourceibias.n363 gnd 0.009861f
C788 commonsourceibias.t100 gnd 0.162395f
C789 commonsourceibias.n364 gnd 0.07189f
C790 commonsourceibias.n365 gnd 0.025003f
C791 commonsourceibias.n366 gnd 0.464917f
C792 commonsourceibias.n367 gnd 0.010724f
C793 commonsourceibias.t140 gnd 0.162395f
C794 commonsourceibias.t155 gnd 0.150157f
C795 commonsourceibias.n368 gnd 0.007823f
C796 commonsourceibias.n369 gnd 0.008037f
C797 commonsourceibias.t84 gnd 0.150157f
C798 commonsourceibias.n370 gnd 0.01034f
C799 commonsourceibias.n371 gnd 0.008037f
C800 commonsourceibias.t148 gnd 0.150157f
C801 commonsourceibias.n372 gnd 0.007578f
C802 commonsourceibias.n373 gnd 0.008037f
C803 commonsourceibias.t80 gnd 0.150157f
C804 commonsourceibias.n374 gnd 0.010186f
C805 commonsourceibias.n375 gnd 0.008037f
C806 commonsourceibias.t113 gnd 0.150157f
C807 commonsourceibias.n376 gnd 0.007361f
C808 commonsourceibias.n377 gnd 0.008037f
C809 commonsourceibias.t154 gnd 0.150157f
C810 commonsourceibias.n378 gnd 0.010015f
C811 commonsourceibias.t29 gnd 0.017343f
C812 commonsourceibias.t3 gnd 0.017343f
C813 commonsourceibias.n379 gnd 0.153763f
C814 commonsourceibias.t49 gnd 0.017343f
C815 commonsourceibias.t13 gnd 0.017343f
C816 commonsourceibias.n380 gnd 0.15325f
C817 commonsourceibias.n381 gnd 0.1428f
C818 commonsourceibias.t69 gnd 0.017343f
C819 commonsourceibias.t67 gnd 0.017343f
C820 commonsourceibias.n382 gnd 0.15325f
C821 commonsourceibias.n383 gnd 0.070394f
C822 commonsourceibias.t7 gnd 0.017343f
C823 commonsourceibias.t63 gnd 0.017343f
C824 commonsourceibias.n384 gnd 0.15325f
C825 commonsourceibias.n385 gnd 0.070394f
C826 commonsourceibias.t53 gnd 0.017343f
C827 commonsourceibias.t73 gnd 0.017343f
C828 commonsourceibias.n386 gnd 0.15325f
C829 commonsourceibias.n387 gnd 0.058811f
C830 commonsourceibias.n388 gnd 0.010724f
C831 commonsourceibias.t42 gnd 0.150157f
C832 commonsourceibias.n389 gnd 0.007823f
C833 commonsourceibias.n390 gnd 0.008037f
C834 commonsourceibias.t0 gnd 0.150157f
C835 commonsourceibias.n391 gnd 0.01034f
C836 commonsourceibias.n392 gnd 0.008037f
C837 commonsourceibias.t60 gnd 0.150157f
C838 commonsourceibias.n393 gnd 0.007578f
C839 commonsourceibias.n394 gnd 0.008037f
C840 commonsourceibias.t16 gnd 0.150157f
C841 commonsourceibias.n395 gnd 0.010186f
C842 commonsourceibias.n396 gnd 0.008037f
C843 commonsourceibias.t58 gnd 0.150157f
C844 commonsourceibias.n397 gnd 0.007361f
C845 commonsourceibias.n398 gnd 0.008037f
C846 commonsourceibias.t32 gnd 0.150157f
C847 commonsourceibias.n399 gnd 0.010015f
C848 commonsourceibias.n400 gnd 0.008037f
C849 commonsourceibias.t72 gnd 0.150157f
C850 commonsourceibias.n401 gnd 0.007172f
C851 commonsourceibias.n402 gnd 0.008037f
C852 commonsourceibias.t52 gnd 0.150157f
C853 commonsourceibias.n403 gnd 0.009825f
C854 commonsourceibias.n404 gnd 0.008037f
C855 commonsourceibias.t6 gnd 0.150157f
C856 commonsourceibias.n405 gnd 0.007008f
C857 commonsourceibias.n406 gnd 0.008037f
C858 commonsourceibias.t66 gnd 0.150157f
C859 commonsourceibias.n407 gnd 0.009613f
C860 commonsourceibias.n408 gnd 0.008037f
C861 commonsourceibias.t12 gnd 0.150157f
C862 commonsourceibias.n409 gnd 0.006868f
C863 commonsourceibias.n410 gnd 0.008037f
C864 commonsourceibias.t48 gnd 0.150157f
C865 commonsourceibias.n411 gnd 0.009378f
C866 commonsourceibias.t28 gnd 0.166947f
C867 commonsourceibias.t2 gnd 0.150157f
C868 commonsourceibias.n412 gnd 0.065449f
C869 commonsourceibias.n413 gnd 0.071822f
C870 commonsourceibias.n414 gnd 0.033327f
C871 commonsourceibias.n415 gnd 0.008037f
C872 commonsourceibias.n416 gnd 0.007823f
C873 commonsourceibias.n417 gnd 0.01121f
C874 commonsourceibias.n418 gnd 0.059912f
C875 commonsourceibias.n419 gnd 0.011203f
C876 commonsourceibias.n420 gnd 0.008037f
C877 commonsourceibias.n421 gnd 0.008037f
C878 commonsourceibias.n422 gnd 0.008037f
C879 commonsourceibias.n423 gnd 0.01034f
C880 commonsourceibias.n424 gnd 0.059912f
C881 commonsourceibias.n425 gnd 0.010583f
C882 commonsourceibias.t68 gnd 0.150157f
C883 commonsourceibias.n426 gnd 0.059912f
C884 commonsourceibias.n427 gnd 0.010282f
C885 commonsourceibias.n428 gnd 0.008037f
C886 commonsourceibias.n429 gnd 0.008037f
C887 commonsourceibias.n430 gnd 0.008037f
C888 commonsourceibias.n431 gnd 0.007578f
C889 commonsourceibias.n432 gnd 0.01122f
C890 commonsourceibias.n433 gnd 0.059912f
C891 commonsourceibias.n434 gnd 0.011217f
C892 commonsourceibias.n435 gnd 0.008037f
C893 commonsourceibias.n436 gnd 0.008037f
C894 commonsourceibias.n437 gnd 0.008037f
C895 commonsourceibias.n438 gnd 0.010186f
C896 commonsourceibias.n439 gnd 0.059912f
C897 commonsourceibias.n440 gnd 0.010507f
C898 commonsourceibias.t62 gnd 0.150157f
C899 commonsourceibias.n441 gnd 0.059912f
C900 commonsourceibias.n442 gnd 0.010357f
C901 commonsourceibias.n443 gnd 0.008037f
C902 commonsourceibias.n444 gnd 0.008037f
C903 commonsourceibias.n445 gnd 0.008037f
C904 commonsourceibias.n446 gnd 0.007361f
C905 commonsourceibias.n447 gnd 0.011225f
C906 commonsourceibias.n448 gnd 0.059912f
C907 commonsourceibias.n449 gnd 0.011224f
C908 commonsourceibias.n450 gnd 0.008037f
C909 commonsourceibias.n451 gnd 0.008037f
C910 commonsourceibias.n452 gnd 0.008037f
C911 commonsourceibias.n453 gnd 0.010015f
C912 commonsourceibias.n454 gnd 0.059912f
C913 commonsourceibias.n455 gnd 0.010432f
C914 commonsourceibias.t64 gnd 0.150157f
C915 commonsourceibias.n456 gnd 0.059912f
C916 commonsourceibias.n457 gnd 0.010432f
C917 commonsourceibias.n458 gnd 0.008037f
C918 commonsourceibias.n459 gnd 0.008037f
C919 commonsourceibias.n460 gnd 0.008037f
C920 commonsourceibias.n461 gnd 0.007172f
C921 commonsourceibias.n462 gnd 0.011224f
C922 commonsourceibias.n463 gnd 0.059912f
C923 commonsourceibias.n464 gnd 0.011225f
C924 commonsourceibias.n465 gnd 0.008037f
C925 commonsourceibias.n466 gnd 0.008037f
C926 commonsourceibias.n467 gnd 0.008037f
C927 commonsourceibias.n468 gnd 0.009825f
C928 commonsourceibias.n469 gnd 0.059912f
C929 commonsourceibias.n470 gnd 0.010357f
C930 commonsourceibias.t44 gnd 0.150157f
C931 commonsourceibias.n471 gnd 0.059912f
C932 commonsourceibias.n472 gnd 0.010507f
C933 commonsourceibias.n473 gnd 0.008037f
C934 commonsourceibias.n474 gnd 0.008037f
C935 commonsourceibias.n475 gnd 0.008037f
C936 commonsourceibias.n476 gnd 0.007008f
C937 commonsourceibias.n477 gnd 0.011217f
C938 commonsourceibias.n478 gnd 0.059912f
C939 commonsourceibias.n479 gnd 0.01122f
C940 commonsourceibias.n480 gnd 0.008037f
C941 commonsourceibias.n481 gnd 0.008037f
C942 commonsourceibias.n482 gnd 0.008037f
C943 commonsourceibias.n483 gnd 0.009613f
C944 commonsourceibias.n484 gnd 0.059912f
C945 commonsourceibias.n485 gnd 0.010282f
C946 commonsourceibias.t30 gnd 0.150157f
C947 commonsourceibias.n486 gnd 0.059912f
C948 commonsourceibias.n487 gnd 0.010583f
C949 commonsourceibias.n488 gnd 0.008037f
C950 commonsourceibias.n489 gnd 0.008037f
C951 commonsourceibias.n490 gnd 0.008037f
C952 commonsourceibias.n491 gnd 0.006868f
C953 commonsourceibias.n492 gnd 0.011203f
C954 commonsourceibias.n493 gnd 0.059912f
C955 commonsourceibias.n494 gnd 0.01121f
C956 commonsourceibias.n495 gnd 0.008037f
C957 commonsourceibias.n496 gnd 0.008037f
C958 commonsourceibias.n497 gnd 0.008037f
C959 commonsourceibias.n498 gnd 0.009378f
C960 commonsourceibias.n499 gnd 0.059912f
C961 commonsourceibias.n500 gnd 0.009861f
C962 commonsourceibias.t14 gnd 0.162395f
C963 commonsourceibias.n501 gnd 0.07189f
C964 commonsourceibias.n502 gnd 0.080075f
C965 commonsourceibias.t43 gnd 0.017343f
C966 commonsourceibias.t15 gnd 0.017343f
C967 commonsourceibias.n503 gnd 0.15325f
C968 commonsourceibias.n504 gnd 0.132562f
C969 commonsourceibias.t31 gnd 0.017343f
C970 commonsourceibias.t1 gnd 0.017343f
C971 commonsourceibias.n505 gnd 0.15325f
C972 commonsourceibias.n506 gnd 0.070394f
C973 commonsourceibias.t17 gnd 0.017343f
C974 commonsourceibias.t61 gnd 0.017343f
C975 commonsourceibias.n507 gnd 0.15325f
C976 commonsourceibias.n508 gnd 0.070394f
C977 commonsourceibias.t59 gnd 0.017343f
C978 commonsourceibias.t45 gnd 0.017343f
C979 commonsourceibias.n509 gnd 0.15325f
C980 commonsourceibias.n510 gnd 0.070394f
C981 commonsourceibias.t65 gnd 0.017343f
C982 commonsourceibias.t33 gnd 0.017343f
C983 commonsourceibias.n511 gnd 0.15325f
C984 commonsourceibias.n512 gnd 0.058811f
C985 commonsourceibias.n513 gnd 0.071213f
C986 commonsourceibias.n514 gnd 0.052016f
C987 commonsourceibias.t82 gnd 0.150157f
C988 commonsourceibias.n515 gnd 0.059912f
C989 commonsourceibias.n516 gnd 0.008037f
C990 commonsourceibias.t147 gnd 0.150157f
C991 commonsourceibias.n517 gnd 0.059912f
C992 commonsourceibias.n518 gnd 0.008037f
C993 commonsourceibias.t143 gnd 0.150157f
C994 commonsourceibias.n519 gnd 0.059912f
C995 commonsourceibias.n520 gnd 0.008037f
C996 commonsourceibias.t158 gnd 0.150157f
C997 commonsourceibias.n521 gnd 0.007008f
C998 commonsourceibias.n522 gnd 0.008037f
C999 commonsourceibias.t104 gnd 0.150157f
C1000 commonsourceibias.n523 gnd 0.009613f
C1001 commonsourceibias.n524 gnd 0.008037f
C1002 commonsourceibias.t133 gnd 0.150157f
C1003 commonsourceibias.n525 gnd 0.006868f
C1004 commonsourceibias.n526 gnd 0.008037f
C1005 commonsourceibias.t150 gnd 0.150157f
C1006 commonsourceibias.n527 gnd 0.009378f
C1007 commonsourceibias.t123 gnd 0.166947f
C1008 commonsourceibias.t103 gnd 0.150157f
C1009 commonsourceibias.n528 gnd 0.065449f
C1010 commonsourceibias.n529 gnd 0.071822f
C1011 commonsourceibias.n530 gnd 0.033327f
C1012 commonsourceibias.n531 gnd 0.008037f
C1013 commonsourceibias.n532 gnd 0.007823f
C1014 commonsourceibias.n533 gnd 0.01121f
C1015 commonsourceibias.n534 gnd 0.059912f
C1016 commonsourceibias.n535 gnd 0.011203f
C1017 commonsourceibias.n536 gnd 0.008037f
C1018 commonsourceibias.n537 gnd 0.008037f
C1019 commonsourceibias.n538 gnd 0.008037f
C1020 commonsourceibias.n539 gnd 0.01034f
C1021 commonsourceibias.n540 gnd 0.059912f
C1022 commonsourceibias.n541 gnd 0.010583f
C1023 commonsourceibias.t114 gnd 0.150157f
C1024 commonsourceibias.n542 gnd 0.059912f
C1025 commonsourceibias.n543 gnd 0.010282f
C1026 commonsourceibias.n544 gnd 0.008037f
C1027 commonsourceibias.n545 gnd 0.008037f
C1028 commonsourceibias.n546 gnd 0.008037f
C1029 commonsourceibias.n547 gnd 0.007578f
C1030 commonsourceibias.n548 gnd 0.01122f
C1031 commonsourceibias.n549 gnd 0.059912f
C1032 commonsourceibias.n550 gnd 0.011217f
C1033 commonsourceibias.n551 gnd 0.008037f
C1034 commonsourceibias.n552 gnd 0.008037f
C1035 commonsourceibias.n553 gnd 0.008037f
C1036 commonsourceibias.n554 gnd 0.010186f
C1037 commonsourceibias.n555 gnd 0.059912f
C1038 commonsourceibias.n556 gnd 0.010507f
C1039 commonsourceibias.n557 gnd 0.010357f
C1040 commonsourceibias.n558 gnd 0.008037f
C1041 commonsourceibias.n559 gnd 0.008037f
C1042 commonsourceibias.n560 gnd 0.009825f
C1043 commonsourceibias.n561 gnd 0.007361f
C1044 commonsourceibias.n562 gnd 0.011225f
C1045 commonsourceibias.n563 gnd 0.008037f
C1046 commonsourceibias.n564 gnd 0.008037f
C1047 commonsourceibias.n565 gnd 0.011224f
C1048 commonsourceibias.n566 gnd 0.007172f
C1049 commonsourceibias.n567 gnd 0.010015f
C1050 commonsourceibias.n568 gnd 0.008037f
C1051 commonsourceibias.n569 gnd 0.007021f
C1052 commonsourceibias.n570 gnd 0.010432f
C1053 commonsourceibias.t85 gnd 0.150157f
C1054 commonsourceibias.n571 gnd 0.059912f
C1055 commonsourceibias.n572 gnd 0.010432f
C1056 commonsourceibias.n573 gnd 0.007021f
C1057 commonsourceibias.n574 gnd 0.008037f
C1058 commonsourceibias.n575 gnd 0.008037f
C1059 commonsourceibias.n576 gnd 0.007172f
C1060 commonsourceibias.n577 gnd 0.011224f
C1061 commonsourceibias.n578 gnd 0.059912f
C1062 commonsourceibias.n579 gnd 0.011225f
C1063 commonsourceibias.n580 gnd 0.008037f
C1064 commonsourceibias.n581 gnd 0.008037f
C1065 commonsourceibias.n582 gnd 0.008037f
C1066 commonsourceibias.n583 gnd 0.009825f
C1067 commonsourceibias.n584 gnd 0.059912f
C1068 commonsourceibias.n585 gnd 0.010357f
C1069 commonsourceibias.t89 gnd 0.150157f
C1070 commonsourceibias.n586 gnd 0.059912f
C1071 commonsourceibias.n587 gnd 0.010507f
C1072 commonsourceibias.n588 gnd 0.008037f
C1073 commonsourceibias.n589 gnd 0.008037f
C1074 commonsourceibias.n590 gnd 0.008037f
C1075 commonsourceibias.n591 gnd 0.007008f
C1076 commonsourceibias.n592 gnd 0.011217f
C1077 commonsourceibias.n593 gnd 0.059912f
C1078 commonsourceibias.n594 gnd 0.01122f
C1079 commonsourceibias.n595 gnd 0.008037f
C1080 commonsourceibias.n596 gnd 0.008037f
C1081 commonsourceibias.n597 gnd 0.008037f
C1082 commonsourceibias.n598 gnd 0.009613f
C1083 commonsourceibias.n599 gnd 0.059912f
C1084 commonsourceibias.n600 gnd 0.010282f
C1085 commonsourceibias.t130 gnd 0.150157f
C1086 commonsourceibias.n601 gnd 0.059912f
C1087 commonsourceibias.n602 gnd 0.010583f
C1088 commonsourceibias.n603 gnd 0.008037f
C1089 commonsourceibias.n604 gnd 0.008037f
C1090 commonsourceibias.n605 gnd 0.008037f
C1091 commonsourceibias.n606 gnd 0.006868f
C1092 commonsourceibias.n607 gnd 0.011203f
C1093 commonsourceibias.n608 gnd 0.059912f
C1094 commonsourceibias.n609 gnd 0.01121f
C1095 commonsourceibias.n610 gnd 0.008037f
C1096 commonsourceibias.n611 gnd 0.008037f
C1097 commonsourceibias.n612 gnd 0.008037f
C1098 commonsourceibias.n613 gnd 0.009378f
C1099 commonsourceibias.n614 gnd 0.059912f
C1100 commonsourceibias.n615 gnd 0.009861f
C1101 commonsourceibias.n616 gnd 0.07189f
C1102 commonsourceibias.n617 gnd 0.04697f
C1103 commonsourceibias.n618 gnd 0.010724f
C1104 commonsourceibias.t142 gnd 0.150157f
C1105 commonsourceibias.n619 gnd 0.007823f
C1106 commonsourceibias.n620 gnd 0.008037f
C1107 commonsourceibias.t156 gnd 0.150157f
C1108 commonsourceibias.n621 gnd 0.01034f
C1109 commonsourceibias.n622 gnd 0.008037f
C1110 commonsourceibias.t132 gnd 0.150157f
C1111 commonsourceibias.n623 gnd 0.007578f
C1112 commonsourceibias.n624 gnd 0.008037f
C1113 commonsourceibias.t149 gnd 0.150157f
C1114 commonsourceibias.n625 gnd 0.010186f
C1115 commonsourceibias.n626 gnd 0.008037f
C1116 commonsourceibias.t97 gnd 0.150157f
C1117 commonsourceibias.n627 gnd 0.007361f
C1118 commonsourceibias.n628 gnd 0.008037f
C1119 commonsourceibias.t141 gnd 0.150157f
C1120 commonsourceibias.n629 gnd 0.010015f
C1121 commonsourceibias.n630 gnd 0.008037f
C1122 commonsourceibias.t152 gnd 0.150157f
C1123 commonsourceibias.n631 gnd 0.007172f
C1124 commonsourceibias.n632 gnd 0.008037f
C1125 commonsourceibias.t131 gnd 0.150157f
C1126 commonsourceibias.n633 gnd 0.009825f
C1127 commonsourceibias.n634 gnd 0.008037f
C1128 commonsourceibias.t145 gnd 0.150157f
C1129 commonsourceibias.n635 gnd 0.007008f
C1130 commonsourceibias.n636 gnd 0.008037f
C1131 commonsourceibias.t91 gnd 0.150157f
C1132 commonsourceibias.n637 gnd 0.009613f
C1133 commonsourceibias.n638 gnd 0.008037f
C1134 commonsourceibias.t116 gnd 0.150157f
C1135 commonsourceibias.n639 gnd 0.006868f
C1136 commonsourceibias.n640 gnd 0.008037f
C1137 commonsourceibias.t134 gnd 0.150157f
C1138 commonsourceibias.n641 gnd 0.009378f
C1139 commonsourceibias.t106 gnd 0.166947f
C1140 commonsourceibias.t90 gnd 0.150157f
C1141 commonsourceibias.n642 gnd 0.065449f
C1142 commonsourceibias.n643 gnd 0.071822f
C1143 commonsourceibias.n644 gnd 0.033327f
C1144 commonsourceibias.n645 gnd 0.008037f
C1145 commonsourceibias.n646 gnd 0.007823f
C1146 commonsourceibias.n647 gnd 0.01121f
C1147 commonsourceibias.n648 gnd 0.059912f
C1148 commonsourceibias.n649 gnd 0.011203f
C1149 commonsourceibias.n650 gnd 0.008037f
C1150 commonsourceibias.n651 gnd 0.008037f
C1151 commonsourceibias.n652 gnd 0.008037f
C1152 commonsourceibias.n653 gnd 0.01034f
C1153 commonsourceibias.n654 gnd 0.059912f
C1154 commonsourceibias.n655 gnd 0.010583f
C1155 commonsourceibias.t96 gnd 0.150157f
C1156 commonsourceibias.n656 gnd 0.059912f
C1157 commonsourceibias.n657 gnd 0.010282f
C1158 commonsourceibias.n658 gnd 0.008037f
C1159 commonsourceibias.n659 gnd 0.008037f
C1160 commonsourceibias.n660 gnd 0.008037f
C1161 commonsourceibias.n661 gnd 0.007578f
C1162 commonsourceibias.n662 gnd 0.01122f
C1163 commonsourceibias.n663 gnd 0.059912f
C1164 commonsourceibias.n664 gnd 0.011217f
C1165 commonsourceibias.n665 gnd 0.008037f
C1166 commonsourceibias.n666 gnd 0.008037f
C1167 commonsourceibias.n667 gnd 0.008037f
C1168 commonsourceibias.n668 gnd 0.010186f
C1169 commonsourceibias.n669 gnd 0.059912f
C1170 commonsourceibias.n670 gnd 0.010507f
C1171 commonsourceibias.t124 gnd 0.150157f
C1172 commonsourceibias.n671 gnd 0.059912f
C1173 commonsourceibias.n672 gnd 0.010357f
C1174 commonsourceibias.n673 gnd 0.008037f
C1175 commonsourceibias.n674 gnd 0.008037f
C1176 commonsourceibias.n675 gnd 0.008037f
C1177 commonsourceibias.n676 gnd 0.007361f
C1178 commonsourceibias.n677 gnd 0.011225f
C1179 commonsourceibias.n678 gnd 0.059912f
C1180 commonsourceibias.n679 gnd 0.011224f
C1181 commonsourceibias.n680 gnd 0.008037f
C1182 commonsourceibias.n681 gnd 0.008037f
C1183 commonsourceibias.n682 gnd 0.008037f
C1184 commonsourceibias.n683 gnd 0.010015f
C1185 commonsourceibias.n684 gnd 0.059912f
C1186 commonsourceibias.n685 gnd 0.010432f
C1187 commonsourceibias.t157 gnd 0.150157f
C1188 commonsourceibias.n686 gnd 0.059912f
C1189 commonsourceibias.n687 gnd 0.010432f
C1190 commonsourceibias.n688 gnd 0.008037f
C1191 commonsourceibias.n689 gnd 0.008037f
C1192 commonsourceibias.n690 gnd 0.008037f
C1193 commonsourceibias.n691 gnd 0.007172f
C1194 commonsourceibias.n692 gnd 0.011224f
C1195 commonsourceibias.n693 gnd 0.059912f
C1196 commonsourceibias.n694 gnd 0.011225f
C1197 commonsourceibias.n695 gnd 0.008037f
C1198 commonsourceibias.n696 gnd 0.008037f
C1199 commonsourceibias.n697 gnd 0.008037f
C1200 commonsourceibias.n698 gnd 0.009825f
C1201 commonsourceibias.n699 gnd 0.059912f
C1202 commonsourceibias.n700 gnd 0.010357f
C1203 commonsourceibias.t81 gnd 0.150157f
C1204 commonsourceibias.n701 gnd 0.059912f
C1205 commonsourceibias.n702 gnd 0.010507f
C1206 commonsourceibias.n703 gnd 0.008037f
C1207 commonsourceibias.n704 gnd 0.008037f
C1208 commonsourceibias.n705 gnd 0.008037f
C1209 commonsourceibias.n706 gnd 0.007008f
C1210 commonsourceibias.n707 gnd 0.011217f
C1211 commonsourceibias.n708 gnd 0.059912f
C1212 commonsourceibias.n709 gnd 0.01122f
C1213 commonsourceibias.n710 gnd 0.008037f
C1214 commonsourceibias.n711 gnd 0.008037f
C1215 commonsourceibias.n712 gnd 0.008037f
C1216 commonsourceibias.n713 gnd 0.009613f
C1217 commonsourceibias.n714 gnd 0.059912f
C1218 commonsourceibias.n715 gnd 0.010282f
C1219 commonsourceibias.t111 gnd 0.150157f
C1220 commonsourceibias.n716 gnd 0.059912f
C1221 commonsourceibias.n717 gnd 0.010583f
C1222 commonsourceibias.n718 gnd 0.008037f
C1223 commonsourceibias.n719 gnd 0.008037f
C1224 commonsourceibias.n720 gnd 0.008037f
C1225 commonsourceibias.n721 gnd 0.006868f
C1226 commonsourceibias.n722 gnd 0.011203f
C1227 commonsourceibias.n723 gnd 0.059912f
C1228 commonsourceibias.n724 gnd 0.01121f
C1229 commonsourceibias.n725 gnd 0.008037f
C1230 commonsourceibias.n726 gnd 0.008037f
C1231 commonsourceibias.n727 gnd 0.008037f
C1232 commonsourceibias.n728 gnd 0.009378f
C1233 commonsourceibias.n729 gnd 0.059912f
C1234 commonsourceibias.n730 gnd 0.009861f
C1235 commonsourceibias.t122 gnd 0.162395f
C1236 commonsourceibias.n731 gnd 0.07189f
C1237 commonsourceibias.n732 gnd 0.025003f
C1238 commonsourceibias.n733 gnd 0.221951f
C1239 commonsourceibias.n734 gnd 4.85761f
C1240 diffpairibias.t27 gnd 0.090128f
C1241 diffpairibias.t23 gnd 0.08996f
C1242 diffpairibias.n0 gnd 0.105991f
C1243 diffpairibias.t28 gnd 0.08996f
C1244 diffpairibias.n1 gnd 0.051736f
C1245 diffpairibias.t25 gnd 0.08996f
C1246 diffpairibias.n2 gnd 0.051736f
C1247 diffpairibias.t29 gnd 0.08996f
C1248 diffpairibias.n3 gnd 0.041084f
C1249 diffpairibias.t15 gnd 0.086371f
C1250 diffpairibias.t1 gnd 0.085993f
C1251 diffpairibias.n4 gnd 0.13579f
C1252 diffpairibias.t11 gnd 0.085993f
C1253 diffpairibias.n5 gnd 0.072463f
C1254 diffpairibias.t13 gnd 0.085993f
C1255 diffpairibias.n6 gnd 0.072463f
C1256 diffpairibias.t7 gnd 0.085993f
C1257 diffpairibias.n7 gnd 0.072463f
C1258 diffpairibias.t3 gnd 0.085993f
C1259 diffpairibias.n8 gnd 0.072463f
C1260 diffpairibias.t17 gnd 0.085993f
C1261 diffpairibias.n9 gnd 0.072463f
C1262 diffpairibias.t5 gnd 0.085993f
C1263 diffpairibias.n10 gnd 0.072463f
C1264 diffpairibias.t19 gnd 0.085993f
C1265 diffpairibias.n11 gnd 0.072463f
C1266 diffpairibias.t9 gnd 0.085993f
C1267 diffpairibias.n12 gnd 0.102883f
C1268 diffpairibias.t14 gnd 0.086899f
C1269 diffpairibias.t0 gnd 0.086748f
C1270 diffpairibias.n13 gnd 0.094648f
C1271 diffpairibias.t10 gnd 0.086748f
C1272 diffpairibias.n14 gnd 0.052262f
C1273 diffpairibias.t12 gnd 0.086748f
C1274 diffpairibias.n15 gnd 0.052262f
C1275 diffpairibias.t6 gnd 0.086748f
C1276 diffpairibias.n16 gnd 0.052262f
C1277 diffpairibias.t2 gnd 0.086748f
C1278 diffpairibias.n17 gnd 0.052262f
C1279 diffpairibias.t16 gnd 0.086748f
C1280 diffpairibias.n18 gnd 0.052262f
C1281 diffpairibias.t4 gnd 0.086748f
C1282 diffpairibias.n19 gnd 0.052262f
C1283 diffpairibias.t18 gnd 0.086748f
C1284 diffpairibias.n20 gnd 0.052262f
C1285 diffpairibias.t8 gnd 0.086748f
C1286 diffpairibias.n21 gnd 0.061849f
C1287 diffpairibias.n22 gnd 0.233513f
C1288 diffpairibias.t20 gnd 0.08996f
C1289 diffpairibias.n23 gnd 0.051747f
C1290 diffpairibias.t26 gnd 0.08996f
C1291 diffpairibias.n24 gnd 0.051736f
C1292 diffpairibias.t22 gnd 0.08996f
C1293 diffpairibias.n25 gnd 0.051736f
C1294 diffpairibias.t21 gnd 0.08996f
C1295 diffpairibias.n26 gnd 0.051736f
C1296 diffpairibias.t24 gnd 0.08996f
C1297 diffpairibias.n27 gnd 0.04729f
C1298 diffpairibias.n28 gnd 0.047711f
C1299 CSoutput.n0 gnd 0.048173f
C1300 CSoutput.t214 gnd 0.318657f
C1301 CSoutput.n1 gnd 0.143889f
C1302 CSoutput.n2 gnd 0.048173f
C1303 CSoutput.t220 gnd 0.318657f
C1304 CSoutput.n3 gnd 0.038181f
C1305 CSoutput.n4 gnd 0.048173f
C1306 CSoutput.t206 gnd 0.318657f
C1307 CSoutput.n5 gnd 0.032924f
C1308 CSoutput.n6 gnd 0.048173f
C1309 CSoutput.t218 gnd 0.318657f
C1310 CSoutput.t216 gnd 0.318657f
C1311 CSoutput.n7 gnd 0.142321f
C1312 CSoutput.n8 gnd 0.048173f
C1313 CSoutput.t203 gnd 0.318657f
C1314 CSoutput.n9 gnd 0.031391f
C1315 CSoutput.n10 gnd 0.048173f
C1316 CSoutput.t209 gnd 0.318657f
C1317 CSoutput.t212 gnd 0.318657f
C1318 CSoutput.n11 gnd 0.142321f
C1319 CSoutput.n12 gnd 0.048173f
C1320 CSoutput.t201 gnd 0.318657f
C1321 CSoutput.n13 gnd 0.032924f
C1322 CSoutput.n14 gnd 0.048173f
C1323 CSoutput.t200 gnd 0.318657f
C1324 CSoutput.t211 gnd 0.318657f
C1325 CSoutput.n15 gnd 0.142321f
C1326 CSoutput.n16 gnd 0.048173f
C1327 CSoutput.t215 gnd 0.318657f
C1328 CSoutput.n17 gnd 0.035165f
C1329 CSoutput.t202 gnd 0.380803f
C1330 CSoutput.t221 gnd 0.318657f
C1331 CSoutput.n18 gnd 0.181689f
C1332 CSoutput.n19 gnd 0.176301f
C1333 CSoutput.n20 gnd 0.20453f
C1334 CSoutput.n21 gnd 0.048173f
C1335 CSoutput.n22 gnd 0.040206f
C1336 CSoutput.n23 gnd 0.142321f
C1337 CSoutput.n24 gnd 0.038757f
C1338 CSoutput.n25 gnd 0.038181f
C1339 CSoutput.n26 gnd 0.048173f
C1340 CSoutput.n27 gnd 0.048173f
C1341 CSoutput.n28 gnd 0.039897f
C1342 CSoutput.n29 gnd 0.033874f
C1343 CSoutput.n30 gnd 0.145489f
C1344 CSoutput.n31 gnd 0.03434f
C1345 CSoutput.n32 gnd 0.048173f
C1346 CSoutput.n33 gnd 0.048173f
C1347 CSoutput.n34 gnd 0.048173f
C1348 CSoutput.n35 gnd 0.039472f
C1349 CSoutput.n36 gnd 0.142321f
C1350 CSoutput.n37 gnd 0.037749f
C1351 CSoutput.n38 gnd 0.039189f
C1352 CSoutput.n39 gnd 0.048173f
C1353 CSoutput.n40 gnd 0.048173f
C1354 CSoutput.n41 gnd 0.040198f
C1355 CSoutput.n42 gnd 0.036741f
C1356 CSoutput.n43 gnd 0.142321f
C1357 CSoutput.n44 gnd 0.037672f
C1358 CSoutput.n45 gnd 0.048173f
C1359 CSoutput.n46 gnd 0.048173f
C1360 CSoutput.n47 gnd 0.048173f
C1361 CSoutput.n48 gnd 0.037672f
C1362 CSoutput.n49 gnd 0.142321f
C1363 CSoutput.n50 gnd 0.036741f
C1364 CSoutput.n51 gnd 0.040198f
C1365 CSoutput.n52 gnd 0.048173f
C1366 CSoutput.n53 gnd 0.048173f
C1367 CSoutput.n54 gnd 0.039189f
C1368 CSoutput.n55 gnd 0.037749f
C1369 CSoutput.n56 gnd 0.142321f
C1370 CSoutput.n57 gnd 0.039472f
C1371 CSoutput.n58 gnd 0.048173f
C1372 CSoutput.n59 gnd 0.048173f
C1373 CSoutput.n60 gnd 0.048173f
C1374 CSoutput.n61 gnd 0.03434f
C1375 CSoutput.n62 gnd 0.145489f
C1376 CSoutput.n63 gnd 0.033874f
C1377 CSoutput.t219 gnd 0.318657f
C1378 CSoutput.n64 gnd 0.142321f
C1379 CSoutput.n65 gnd 0.039897f
C1380 CSoutput.n66 gnd 0.048173f
C1381 CSoutput.n67 gnd 0.048173f
C1382 CSoutput.n68 gnd 0.048173f
C1383 CSoutput.n69 gnd 0.038757f
C1384 CSoutput.n70 gnd 0.142321f
C1385 CSoutput.n71 gnd 0.040206f
C1386 CSoutput.n72 gnd 0.035165f
C1387 CSoutput.n73 gnd 0.048173f
C1388 CSoutput.n74 gnd 0.048173f
C1389 CSoutput.n75 gnd 0.036468f
C1390 CSoutput.n76 gnd 0.021659f
C1391 CSoutput.t204 gnd 0.358034f
C1392 CSoutput.n77 gnd 0.177857f
C1393 CSoutput.n78 gnd 0.761033f
C1394 CSoutput.t110 gnd 0.06009f
C1395 CSoutput.t8 gnd 0.06009f
C1396 CSoutput.n79 gnd 0.465233f
C1397 CSoutput.t90 gnd 0.06009f
C1398 CSoutput.t60 gnd 0.06009f
C1399 CSoutput.n80 gnd 0.464404f
C1400 CSoutput.n81 gnd 0.471369f
C1401 CSoutput.t99 gnd 0.06009f
C1402 CSoutput.t36 gnd 0.06009f
C1403 CSoutput.n82 gnd 0.464404f
C1404 CSoutput.n83 gnd 0.232271f
C1405 CSoutput.t118 gnd 0.06009f
C1406 CSoutput.t53 gnd 0.06009f
C1407 CSoutput.n84 gnd 0.464404f
C1408 CSoutput.n85 gnd 0.232271f
C1409 CSoutput.t14 gnd 0.06009f
C1410 CSoutput.t69 gnd 0.06009f
C1411 CSoutput.n86 gnd 0.464404f
C1412 CSoutput.n87 gnd 0.232271f
C1413 CSoutput.t19 gnd 0.06009f
C1414 CSoutput.t45 gnd 0.06009f
C1415 CSoutput.n88 gnd 0.464404f
C1416 CSoutput.n89 gnd 0.232271f
C1417 CSoutput.t123 gnd 0.06009f
C1418 CSoutput.t62 gnd 0.06009f
C1419 CSoutput.n90 gnd 0.464404f
C1420 CSoutput.n91 gnd 0.232271f
C1421 CSoutput.t22 gnd 0.06009f
C1422 CSoutput.t106 gnd 0.06009f
C1423 CSoutput.n92 gnd 0.464404f
C1424 CSoutput.n93 gnd 0.232271f
C1425 CSoutput.t32 gnd 0.06009f
C1426 CSoutput.t81 gnd 0.06009f
C1427 CSoutput.n94 gnd 0.464404f
C1428 CSoutput.n95 gnd 0.232271f
C1429 CSoutput.t48 gnd 0.06009f
C1430 CSoutput.t70 gnd 0.06009f
C1431 CSoutput.n96 gnd 0.464404f
C1432 CSoutput.n97 gnd 0.425931f
C1433 CSoutput.t103 gnd 0.06009f
C1434 CSoutput.t101 gnd 0.06009f
C1435 CSoutput.n98 gnd 0.465233f
C1436 CSoutput.t83 gnd 0.06009f
C1437 CSoutput.t15 gnd 0.06009f
C1438 CSoutput.n99 gnd 0.464404f
C1439 CSoutput.n100 gnd 0.471369f
C1440 CSoutput.t9 gnd 0.06009f
C1441 CSoutput.t97 gnd 0.06009f
C1442 CSoutput.n101 gnd 0.464404f
C1443 CSoutput.n102 gnd 0.232271f
C1444 CSoutput.t82 gnd 0.06009f
C1445 CSoutput.t55 gnd 0.06009f
C1446 CSoutput.n103 gnd 0.464404f
C1447 CSoutput.n104 gnd 0.232271f
C1448 CSoutput.t37 gnd 0.06009f
C1449 CSoutput.t113 gnd 0.06009f
C1450 CSoutput.n105 gnd 0.464404f
C1451 CSoutput.n106 gnd 0.232271f
C1452 CSoutput.t79 gnd 0.06009f
C1453 CSoutput.t78 gnd 0.06009f
C1454 CSoutput.n107 gnd 0.464404f
C1455 CSoutput.n108 gnd 0.232271f
C1456 CSoutput.t66 gnd 0.06009f
C1457 CSoutput.t33 gnd 0.06009f
C1458 CSoutput.n109 gnd 0.464404f
C1459 CSoutput.n110 gnd 0.232271f
C1460 CSoutput.t13 gnd 0.06009f
C1461 CSoutput.t67 gnd 0.06009f
C1462 CSoutput.n111 gnd 0.464404f
C1463 CSoutput.n112 gnd 0.232271f
C1464 CSoutput.t63 gnd 0.06009f
C1465 CSoutput.t31 gnd 0.06009f
C1466 CSoutput.n113 gnd 0.464404f
C1467 CSoutput.n114 gnd 0.232271f
C1468 CSoutput.t10 gnd 0.06009f
C1469 CSoutput.t6 gnd 0.06009f
C1470 CSoutput.n115 gnd 0.464404f
C1471 CSoutput.n116 gnd 0.346374f
C1472 CSoutput.n117 gnd 0.436776f
C1473 CSoutput.t115 gnd 0.06009f
C1474 CSoutput.t114 gnd 0.06009f
C1475 CSoutput.n118 gnd 0.465233f
C1476 CSoutput.t94 gnd 0.06009f
C1477 CSoutput.t28 gnd 0.06009f
C1478 CSoutput.n119 gnd 0.464404f
C1479 CSoutput.n120 gnd 0.471369f
C1480 CSoutput.t25 gnd 0.06009f
C1481 CSoutput.t112 gnd 0.06009f
C1482 CSoutput.n121 gnd 0.464404f
C1483 CSoutput.n122 gnd 0.232271f
C1484 CSoutput.t91 gnd 0.06009f
C1485 CSoutput.t68 gnd 0.06009f
C1486 CSoutput.n123 gnd 0.464404f
C1487 CSoutput.n124 gnd 0.232271f
C1488 CSoutput.t49 gnd 0.06009f
C1489 CSoutput.t124 gnd 0.06009f
C1490 CSoutput.n125 gnd 0.464404f
C1491 CSoutput.n126 gnd 0.232271f
C1492 CSoutput.t89 gnd 0.06009f
C1493 CSoutput.t88 gnd 0.06009f
C1494 CSoutput.n127 gnd 0.464404f
C1495 CSoutput.n128 gnd 0.232271f
C1496 CSoutput.t76 gnd 0.06009f
C1497 CSoutput.t46 gnd 0.06009f
C1498 CSoutput.n129 gnd 0.464404f
C1499 CSoutput.n130 gnd 0.232271f
C1500 CSoutput.t27 gnd 0.06009f
C1501 CSoutput.t77 gnd 0.06009f
C1502 CSoutput.n131 gnd 0.464404f
C1503 CSoutput.n132 gnd 0.232271f
C1504 CSoutput.t73 gnd 0.06009f
C1505 CSoutput.t44 gnd 0.06009f
C1506 CSoutput.n133 gnd 0.464404f
C1507 CSoutput.n134 gnd 0.232271f
C1508 CSoutput.t24 gnd 0.06009f
C1509 CSoutput.t23 gnd 0.06009f
C1510 CSoutput.n135 gnd 0.464404f
C1511 CSoutput.n136 gnd 0.346374f
C1512 CSoutput.n137 gnd 0.488203f
C1513 CSoutput.n138 gnd 10.1684f
C1514 CSoutput.n140 gnd 0.852179f
C1515 CSoutput.n141 gnd 0.639134f
C1516 CSoutput.n142 gnd 0.852179f
C1517 CSoutput.n143 gnd 0.852179f
C1518 CSoutput.n144 gnd 2.29433f
C1519 CSoutput.n145 gnd 0.852179f
C1520 CSoutput.n146 gnd 0.852179f
C1521 CSoutput.t210 gnd 1.06522f
C1522 CSoutput.n147 gnd 0.852179f
C1523 CSoutput.n148 gnd 0.852179f
C1524 CSoutput.n152 gnd 0.852179f
C1525 CSoutput.n156 gnd 0.852179f
C1526 CSoutput.n157 gnd 0.852179f
C1527 CSoutput.n159 gnd 0.852179f
C1528 CSoutput.n164 gnd 0.852179f
C1529 CSoutput.n166 gnd 0.852179f
C1530 CSoutput.n167 gnd 0.852179f
C1531 CSoutput.n169 gnd 0.852179f
C1532 CSoutput.n170 gnd 0.852179f
C1533 CSoutput.n172 gnd 0.852179f
C1534 CSoutput.t205 gnd 14.239799f
C1535 CSoutput.n174 gnd 0.852179f
C1536 CSoutput.n175 gnd 0.639134f
C1537 CSoutput.n176 gnd 0.852179f
C1538 CSoutput.n177 gnd 0.852179f
C1539 CSoutput.n178 gnd 2.29433f
C1540 CSoutput.n179 gnd 0.852179f
C1541 CSoutput.n180 gnd 0.852179f
C1542 CSoutput.t207 gnd 1.06522f
C1543 CSoutput.n181 gnd 0.852179f
C1544 CSoutput.n182 gnd 0.852179f
C1545 CSoutput.n186 gnd 0.852179f
C1546 CSoutput.n190 gnd 0.852179f
C1547 CSoutput.n191 gnd 0.852179f
C1548 CSoutput.n193 gnd 0.852179f
C1549 CSoutput.n198 gnd 0.852179f
C1550 CSoutput.n200 gnd 0.852179f
C1551 CSoutput.n201 gnd 0.852179f
C1552 CSoutput.n203 gnd 0.852179f
C1553 CSoutput.n204 gnd 0.852179f
C1554 CSoutput.n206 gnd 0.852179f
C1555 CSoutput.n207 gnd 0.639134f
C1556 CSoutput.n209 gnd 0.852179f
C1557 CSoutput.n210 gnd 0.639134f
C1558 CSoutput.n211 gnd 0.852179f
C1559 CSoutput.n212 gnd 0.852179f
C1560 CSoutput.n213 gnd 2.29433f
C1561 CSoutput.n214 gnd 0.852179f
C1562 CSoutput.n215 gnd 0.852179f
C1563 CSoutput.t208 gnd 1.06522f
C1564 CSoutput.n216 gnd 0.852179f
C1565 CSoutput.n217 gnd 2.29433f
C1566 CSoutput.n219 gnd 0.852179f
C1567 CSoutput.n220 gnd 0.852179f
C1568 CSoutput.n222 gnd 0.852179f
C1569 CSoutput.n223 gnd 0.852179f
C1570 CSoutput.t217 gnd 14.0078f
C1571 CSoutput.t213 gnd 14.239799f
C1572 CSoutput.n229 gnd 2.67341f
C1573 CSoutput.n230 gnd 10.8905f
C1574 CSoutput.n231 gnd 11.3462f
C1575 CSoutput.n236 gnd 2.89602f
C1576 CSoutput.n242 gnd 0.852179f
C1577 CSoutput.n244 gnd 0.852179f
C1578 CSoutput.n246 gnd 0.852179f
C1579 CSoutput.n248 gnd 0.852179f
C1580 CSoutput.n250 gnd 0.852179f
C1581 CSoutput.n256 gnd 0.852179f
C1582 CSoutput.n263 gnd 1.56342f
C1583 CSoutput.n264 gnd 1.56342f
C1584 CSoutput.n265 gnd 0.852179f
C1585 CSoutput.n266 gnd 0.852179f
C1586 CSoutput.n268 gnd 0.639134f
C1587 CSoutput.n269 gnd 0.547361f
C1588 CSoutput.n271 gnd 0.639134f
C1589 CSoutput.n272 gnd 0.547361f
C1590 CSoutput.n273 gnd 0.639134f
C1591 CSoutput.n275 gnd 0.852179f
C1592 CSoutput.n277 gnd 2.29433f
C1593 CSoutput.n278 gnd 2.67341f
C1594 CSoutput.n279 gnd 10.0165f
C1595 CSoutput.n281 gnd 0.639134f
C1596 CSoutput.n282 gnd 1.64453f
C1597 CSoutput.n283 gnd 0.639134f
C1598 CSoutput.n285 gnd 0.852179f
C1599 CSoutput.n287 gnd 2.29433f
C1600 CSoutput.n288 gnd 4.99742f
C1601 CSoutput.t7 gnd 0.06009f
C1602 CSoutput.t109 gnd 0.06009f
C1603 CSoutput.n289 gnd 0.465233f
C1604 CSoutput.t59 gnd 0.06009f
C1605 CSoutput.t122 gnd 0.06009f
C1606 CSoutput.n290 gnd 0.464404f
C1607 CSoutput.n291 gnd 0.471369f
C1608 CSoutput.t35 gnd 0.06009f
C1609 CSoutput.t98 gnd 0.06009f
C1610 CSoutput.n292 gnd 0.464404f
C1611 CSoutput.n293 gnd 0.232271f
C1612 CSoutput.t52 gnd 0.06009f
C1613 CSoutput.t116 gnd 0.06009f
C1614 CSoutput.n294 gnd 0.464404f
C1615 CSoutput.n295 gnd 0.232271f
C1616 CSoutput.t92 gnd 0.06009f
C1617 CSoutput.t12 gnd 0.06009f
C1618 CSoutput.n296 gnd 0.464404f
C1619 CSoutput.n297 gnd 0.232271f
C1620 CSoutput.t43 gnd 0.06009f
C1621 CSoutput.t18 gnd 0.06009f
C1622 CSoutput.n298 gnd 0.464404f
C1623 CSoutput.n299 gnd 0.232271f
C1624 CSoutput.t61 gnd 0.06009f
C1625 CSoutput.t40 gnd 0.06009f
C1626 CSoutput.n300 gnd 0.464404f
C1627 CSoutput.n301 gnd 0.232271f
C1628 CSoutput.t105 gnd 0.06009f
C1629 CSoutput.t21 gnd 0.06009f
C1630 CSoutput.n302 gnd 0.464404f
C1631 CSoutput.n303 gnd 0.232271f
C1632 CSoutput.t80 gnd 0.06009f
C1633 CSoutput.t29 gnd 0.06009f
C1634 CSoutput.n304 gnd 0.464404f
C1635 CSoutput.n305 gnd 0.232271f
C1636 CSoutput.t93 gnd 0.06009f
C1637 CSoutput.t47 gnd 0.06009f
C1638 CSoutput.n306 gnd 0.464404f
C1639 CSoutput.n307 gnd 0.425931f
C1640 CSoutput.t64 gnd 0.06009f
C1641 CSoutput.t65 gnd 0.06009f
C1642 CSoutput.n308 gnd 0.465233f
C1643 CSoutput.t87 gnd 0.06009f
C1644 CSoutput.t11 gnd 0.06009f
C1645 CSoutput.n309 gnd 0.464404f
C1646 CSoutput.n310 gnd 0.471369f
C1647 CSoutput.t57 gnd 0.06009f
C1648 CSoutput.t85 gnd 0.06009f
C1649 CSoutput.n311 gnd 0.464404f
C1650 CSoutput.n312 gnd 0.232271f
C1651 CSoutput.t125 gnd 0.06009f
C1652 CSoutput.t41 gnd 0.06009f
C1653 CSoutput.n313 gnd 0.464404f
C1654 CSoutput.n314 gnd 0.232271f
C1655 CSoutput.t42 gnd 0.06009f
C1656 CSoutput.t111 gnd 0.06009f
C1657 CSoutput.n315 gnd 0.464404f
C1658 CSoutput.n316 gnd 0.232271f
C1659 CSoutput.t38 gnd 0.06009f
C1660 CSoutput.t39 gnd 0.06009f
C1661 CSoutput.n317 gnd 0.464404f
C1662 CSoutput.n318 gnd 0.232271f
C1663 CSoutput.t107 gnd 0.06009f
C1664 CSoutput.t108 gnd 0.06009f
C1665 CSoutput.n319 gnd 0.464404f
C1666 CSoutput.n320 gnd 0.232271f
C1667 CSoutput.t17 gnd 0.06009f
C1668 CSoutput.t86 gnd 0.06009f
C1669 CSoutput.n321 gnd 0.464404f
C1670 CSoutput.n322 gnd 0.232271f
C1671 CSoutput.t104 gnd 0.06009f
C1672 CSoutput.t16 gnd 0.06009f
C1673 CSoutput.n323 gnd 0.464404f
C1674 CSoutput.n324 gnd 0.232271f
C1675 CSoutput.t58 gnd 0.06009f
C1676 CSoutput.t84 gnd 0.06009f
C1677 CSoutput.n325 gnd 0.464404f
C1678 CSoutput.n326 gnd 0.346374f
C1679 CSoutput.n327 gnd 0.436776f
C1680 CSoutput.t74 gnd 0.06009f
C1681 CSoutput.t75 gnd 0.06009f
C1682 CSoutput.n328 gnd 0.465233f
C1683 CSoutput.t102 gnd 0.06009f
C1684 CSoutput.t26 gnd 0.06009f
C1685 CSoutput.n329 gnd 0.464404f
C1686 CSoutput.n330 gnd 0.471369f
C1687 CSoutput.t71 gnd 0.06009f
C1688 CSoutput.t95 gnd 0.06009f
C1689 CSoutput.n331 gnd 0.464404f
C1690 CSoutput.n332 gnd 0.232271f
C1691 CSoutput.t20 gnd 0.06009f
C1692 CSoutput.t54 gnd 0.06009f
C1693 CSoutput.n333 gnd 0.464404f
C1694 CSoutput.n334 gnd 0.232271f
C1695 CSoutput.t56 gnd 0.06009f
C1696 CSoutput.t121 gnd 0.06009f
C1697 CSoutput.n335 gnd 0.464404f
C1698 CSoutput.n336 gnd 0.232271f
C1699 CSoutput.t50 gnd 0.06009f
C1700 CSoutput.t51 gnd 0.06009f
C1701 CSoutput.n337 gnd 0.464404f
C1702 CSoutput.n338 gnd 0.232271f
C1703 CSoutput.t119 gnd 0.06009f
C1704 CSoutput.t120 gnd 0.06009f
C1705 CSoutput.n339 gnd 0.464404f
C1706 CSoutput.n340 gnd 0.232271f
C1707 CSoutput.t34 gnd 0.06009f
C1708 CSoutput.t100 gnd 0.06009f
C1709 CSoutput.n341 gnd 0.464404f
C1710 CSoutput.n342 gnd 0.232271f
C1711 CSoutput.t117 gnd 0.06009f
C1712 CSoutput.t30 gnd 0.06009f
C1713 CSoutput.n343 gnd 0.464404f
C1714 CSoutput.n344 gnd 0.232271f
C1715 CSoutput.t72 gnd 0.06009f
C1716 CSoutput.t96 gnd 0.06009f
C1717 CSoutput.n345 gnd 0.464402f
C1718 CSoutput.n346 gnd 0.346376f
C1719 CSoutput.n347 gnd 0.488203f
C1720 CSoutput.n348 gnd 13.9948f
C1721 CSoutput.t171 gnd 0.052578f
C1722 CSoutput.t140 gnd 0.052578f
C1723 CSoutput.n349 gnd 0.466156f
C1724 CSoutput.t127 gnd 0.052578f
C1725 CSoutput.t190 gnd 0.052578f
C1726 CSoutput.n350 gnd 0.464601f
C1727 CSoutput.n351 gnd 0.432921f
C1728 CSoutput.t130 gnd 0.052578f
C1729 CSoutput.t152 gnd 0.052578f
C1730 CSoutput.n352 gnd 0.464601f
C1731 CSoutput.n353 gnd 0.21341f
C1732 CSoutput.t160 gnd 0.052578f
C1733 CSoutput.t164 gnd 0.052578f
C1734 CSoutput.n354 gnd 0.464601f
C1735 CSoutput.n355 gnd 0.21341f
C1736 CSoutput.t1 gnd 0.052578f
C1737 CSoutput.t139 gnd 0.052578f
C1738 CSoutput.n356 gnd 0.464601f
C1739 CSoutput.n357 gnd 0.21341f
C1740 CSoutput.t166 gnd 0.052578f
C1741 CSoutput.t158 gnd 0.052578f
C1742 CSoutput.n358 gnd 0.464601f
C1743 CSoutput.n359 gnd 0.21341f
C1744 CSoutput.t184 gnd 0.052578f
C1745 CSoutput.t198 gnd 0.052578f
C1746 CSoutput.n360 gnd 0.464601f
C1747 CSoutput.n361 gnd 0.21341f
C1748 CSoutput.t133 gnd 0.052578f
C1749 CSoutput.t170 gnd 0.052578f
C1750 CSoutput.n362 gnd 0.464601f
C1751 CSoutput.n363 gnd 0.21341f
C1752 CSoutput.t157 gnd 0.052578f
C1753 CSoutput.t154 gnd 0.052578f
C1754 CSoutput.n364 gnd 0.464601f
C1755 CSoutput.n365 gnd 0.21341f
C1756 CSoutput.t161 gnd 0.052578f
C1757 CSoutput.t168 gnd 0.052578f
C1758 CSoutput.n366 gnd 0.464601f
C1759 CSoutput.n367 gnd 0.393571f
C1760 CSoutput.t159 gnd 0.052578f
C1761 CSoutput.t185 gnd 0.052578f
C1762 CSoutput.n368 gnd 0.466156f
C1763 CSoutput.t0 gnd 0.052578f
C1764 CSoutput.t180 gnd 0.052578f
C1765 CSoutput.n369 gnd 0.464601f
C1766 CSoutput.n370 gnd 0.432921f
C1767 CSoutput.t138 gnd 0.052578f
C1768 CSoutput.t149 gnd 0.052578f
C1769 CSoutput.n371 gnd 0.464601f
C1770 CSoutput.n372 gnd 0.21341f
C1771 CSoutput.t150 gnd 0.052578f
C1772 CSoutput.t5 gnd 0.052578f
C1773 CSoutput.n373 gnd 0.464601f
C1774 CSoutput.n374 gnd 0.21341f
C1775 CSoutput.t186 gnd 0.052578f
C1776 CSoutput.t194 gnd 0.052578f
C1777 CSoutput.n375 gnd 0.464601f
C1778 CSoutput.n376 gnd 0.21341f
C1779 CSoutput.t172 gnd 0.052578f
C1780 CSoutput.t188 gnd 0.052578f
C1781 CSoutput.n377 gnd 0.464601f
C1782 CSoutput.n378 gnd 0.21341f
C1783 CSoutput.t192 gnd 0.052578f
C1784 CSoutput.t195 gnd 0.052578f
C1785 CSoutput.n379 gnd 0.464601f
C1786 CSoutput.n380 gnd 0.21341f
C1787 CSoutput.t165 gnd 0.052578f
C1788 CSoutput.t181 gnd 0.052578f
C1789 CSoutput.n381 gnd 0.464601f
C1790 CSoutput.n382 gnd 0.21341f
C1791 CSoutput.t134 gnd 0.052578f
C1792 CSoutput.t2 gnd 0.052578f
C1793 CSoutput.n383 gnd 0.464601f
C1794 CSoutput.n384 gnd 0.21341f
C1795 CSoutput.t151 gnd 0.052578f
C1796 CSoutput.t193 gnd 0.052578f
C1797 CSoutput.n385 gnd 0.464601f
C1798 CSoutput.n386 gnd 0.324002f
C1799 CSoutput.n387 gnd 0.60202f
C1800 CSoutput.n388 gnd 14.9575f
C1801 CSoutput.t142 gnd 0.052578f
C1802 CSoutput.t174 gnd 0.052578f
C1803 CSoutput.n389 gnd 0.466156f
C1804 CSoutput.t129 gnd 0.052578f
C1805 CSoutput.t176 gnd 0.052578f
C1806 CSoutput.n390 gnd 0.464601f
C1807 CSoutput.n391 gnd 0.432921f
C1808 CSoutput.t196 gnd 0.052578f
C1809 CSoutput.t153 gnd 0.052578f
C1810 CSoutput.n392 gnd 0.464601f
C1811 CSoutput.n393 gnd 0.21341f
C1812 CSoutput.t136 gnd 0.052578f
C1813 CSoutput.t167 gnd 0.052578f
C1814 CSoutput.n394 gnd 0.464601f
C1815 CSoutput.n395 gnd 0.21341f
C1816 CSoutput.t177 gnd 0.052578f
C1817 CSoutput.t126 gnd 0.052578f
C1818 CSoutput.n396 gnd 0.464601f
C1819 CSoutput.n397 gnd 0.21341f
C1820 CSoutput.t145 gnd 0.052578f
C1821 CSoutput.t4 gnd 0.052578f
C1822 CSoutput.n398 gnd 0.464601f
C1823 CSoutput.n399 gnd 0.21341f
C1824 CSoutput.t178 gnd 0.052578f
C1825 CSoutput.t147 gnd 0.052578f
C1826 CSoutput.n400 gnd 0.464601f
C1827 CSoutput.n401 gnd 0.21341f
C1828 CSoutput.t132 gnd 0.052578f
C1829 CSoutput.t187 gnd 0.052578f
C1830 CSoutput.n402 gnd 0.464601f
C1831 CSoutput.n403 gnd 0.21341f
C1832 CSoutput.t131 gnd 0.052578f
C1833 CSoutput.t135 gnd 0.052578f
C1834 CSoutput.n404 gnd 0.464601f
C1835 CSoutput.n405 gnd 0.21341f
C1836 CSoutput.t175 gnd 0.052578f
C1837 CSoutput.t191 gnd 0.052578f
C1838 CSoutput.n406 gnd 0.464601f
C1839 CSoutput.n407 gnd 0.393571f
C1840 CSoutput.t155 gnd 0.052578f
C1841 CSoutput.t199 gnd 0.052578f
C1842 CSoutput.n408 gnd 0.466156f
C1843 CSoutput.t137 gnd 0.052578f
C1844 CSoutput.t179 gnd 0.052578f
C1845 CSoutput.n409 gnd 0.464601f
C1846 CSoutput.n410 gnd 0.432921f
C1847 CSoutput.t144 gnd 0.052578f
C1848 CSoutput.t3 gnd 0.052578f
C1849 CSoutput.n411 gnd 0.464601f
C1850 CSoutput.n412 gnd 0.21341f
C1851 CSoutput.t163 gnd 0.052578f
C1852 CSoutput.t197 gnd 0.052578f
C1853 CSoutput.n413 gnd 0.464601f
C1854 CSoutput.n414 gnd 0.21341f
C1855 CSoutput.t141 gnd 0.052578f
C1856 CSoutput.t156 gnd 0.052578f
C1857 CSoutput.n415 gnd 0.464601f
C1858 CSoutput.n416 gnd 0.21341f
C1859 CSoutput.t148 gnd 0.052578f
C1860 CSoutput.t143 gnd 0.052578f
C1861 CSoutput.n417 gnd 0.464601f
C1862 CSoutput.n418 gnd 0.21341f
C1863 CSoutput.t146 gnd 0.052578f
C1864 CSoutput.t169 gnd 0.052578f
C1865 CSoutput.n419 gnd 0.464601f
C1866 CSoutput.n420 gnd 0.21341f
C1867 CSoutput.t162 gnd 0.052578f
C1868 CSoutput.t183 gnd 0.052578f
C1869 CSoutput.n421 gnd 0.464601f
C1870 CSoutput.n422 gnd 0.21341f
C1871 CSoutput.t128 gnd 0.052578f
C1872 CSoutput.t173 gnd 0.052578f
C1873 CSoutput.n423 gnd 0.464601f
C1874 CSoutput.n424 gnd 0.21341f
C1875 CSoutput.t189 gnd 0.052578f
C1876 CSoutput.t182 gnd 0.052578f
C1877 CSoutput.n425 gnd 0.464601f
C1878 CSoutput.n426 gnd 0.324002f
C1879 CSoutput.n427 gnd 0.60202f
C1880 CSoutput.n428 gnd 9.09676f
C1881 CSoutput.n429 gnd 15.7036f
C1882 a_n7636_8799.t8 gnd 0.144247f
C1883 a_n7636_8799.t0 gnd 0.144247f
C1884 a_n7636_8799.t7 gnd 0.144247f
C1885 a_n7636_8799.n0 gnd 1.1377f
C1886 a_n7636_8799.t6 gnd 0.144247f
C1887 a_n7636_8799.t9 gnd 0.144247f
C1888 a_n7636_8799.n1 gnd 1.13582f
C1889 a_n7636_8799.n2 gnd 1.02096f
C1890 a_n7636_8799.t4 gnd 0.144247f
C1891 a_n7636_8799.t1 gnd 0.144247f
C1892 a_n7636_8799.n3 gnd 1.13582f
C1893 a_n7636_8799.n4 gnd 1.77238f
C1894 a_n7636_8799.t29 gnd 0.112192f
C1895 a_n7636_8799.t35 gnd 0.112192f
C1896 a_n7636_8799.n5 gnd 0.994289f
C1897 a_n7636_8799.t18 gnd 0.112192f
C1898 a_n7636_8799.t19 gnd 0.112192f
C1899 a_n7636_8799.n6 gnd 0.991366f
C1900 a_n7636_8799.n7 gnd 0.879091f
C1901 a_n7636_8799.t24 gnd 0.112192f
C1902 a_n7636_8799.t23 gnd 0.112192f
C1903 a_n7636_8799.n8 gnd 0.991366f
C1904 a_n7636_8799.n9 gnd 0.363542f
C1905 a_n7636_8799.t20 gnd 0.112192f
C1906 a_n7636_8799.t17 gnd 0.112192f
C1907 a_n7636_8799.n10 gnd 0.994288f
C1908 a_n7636_8799.t34 gnd 0.112192f
C1909 a_n7636_8799.t28 gnd 0.112192f
C1910 a_n7636_8799.n11 gnd 0.991365f
C1911 a_n7636_8799.n12 gnd 0.879094f
C1912 a_n7636_8799.t32 gnd 0.112192f
C1913 a_n7636_8799.t33 gnd 0.112192f
C1914 a_n7636_8799.n13 gnd 0.991365f
C1915 a_n7636_8799.n14 gnd 0.363543f
C1916 a_n7636_8799.t31 gnd 0.112192f
C1917 a_n7636_8799.t26 gnd 0.112192f
C1918 a_n7636_8799.n15 gnd 0.994288f
C1919 a_n7636_8799.t13 gnd 0.112192f
C1920 a_n7636_8799.t15 gnd 0.112192f
C1921 a_n7636_8799.n16 gnd 0.991365f
C1922 a_n7636_8799.n17 gnd 0.879094f
C1923 a_n7636_8799.t21 gnd 0.112192f
C1924 a_n7636_8799.t22 gnd 0.112192f
C1925 a_n7636_8799.n18 gnd 0.991365f
C1926 a_n7636_8799.n19 gnd 0.363543f
C1927 a_n7636_8799.n20 gnd 2.68328f
C1928 a_n7636_8799.t12 gnd 0.112192f
C1929 a_n7636_8799.t16 gnd 0.112192f
C1930 a_n7636_8799.n21 gnd 0.991366f
C1931 a_n7636_8799.n22 gnd 3.09255f
C1932 a_n7636_8799.t30 gnd 0.112192f
C1933 a_n7636_8799.t14 gnd 0.112192f
C1934 a_n7636_8799.n23 gnd 0.991366f
C1935 a_n7636_8799.n24 gnd 0.432838f
C1936 a_n7636_8799.t27 gnd 0.112192f
C1937 a_n7636_8799.t25 gnd 0.112192f
C1938 a_n7636_8799.n25 gnd 0.991366f
C1939 a_n7636_8799.n26 gnd 0.363542f
C1940 a_n7636_8799.n27 gnd 0.493296f
C1941 a_n7636_8799.n28 gnd 0.051991f
C1942 a_n7636_8799.t133 gnd 0.598113f
C1943 a_n7636_8799.n29 gnd 0.267129f
C1944 a_n7636_8799.n30 gnd 0.051991f
C1945 a_n7636_8799.n31 gnd 0.011798f
C1946 a_n7636_8799.t49 gnd 0.598113f
C1947 a_n7636_8799.n32 gnd 0.051991f
C1948 a_n7636_8799.t70 gnd 0.598113f
C1949 a_n7636_8799.n33 gnd 0.264084f
C1950 a_n7636_8799.t93 gnd 0.598113f
C1951 a_n7636_8799.n34 gnd 0.051991f
C1952 a_n7636_8799.t112 gnd 0.598113f
C1953 a_n7636_8799.n35 gnd 0.264404f
C1954 a_n7636_8799.n36 gnd 0.051991f
C1955 a_n7636_8799.n37 gnd 0.011798f
C1956 a_n7636_8799.t72 gnd 0.598113f
C1957 a_n7636_8799.n38 gnd 0.051991f
C1958 a_n7636_8799.t84 gnd 0.598113f
C1959 a_n7636_8799.n39 gnd 0.267129f
C1960 a_n7636_8799.n40 gnd 0.051991f
C1961 a_n7636_8799.n41 gnd 0.011798f
C1962 a_n7636_8799.t117 gnd 0.598113f
C1963 a_n7636_8799.n42 gnd 0.164254f
C1964 a_n7636_8799.t138 gnd 0.598113f
C1965 a_n7636_8799.t137 gnd 0.609434f
C1966 a_n7636_8799.n43 gnd 0.250733f
C1967 a_n7636_8799.n44 gnd 0.263443f
C1968 a_n7636_8799.n45 gnd 0.011798f
C1969 a_n7636_8799.t88 gnd 0.598113f
C1970 a_n7636_8799.n46 gnd 0.267129f
C1971 a_n7636_8799.n47 gnd 0.051991f
C1972 a_n7636_8799.n48 gnd 0.051991f
C1973 a_n7636_8799.n49 gnd 0.051991f
C1974 a_n7636_8799.n50 gnd 0.265045f
C1975 a_n7636_8799.t134 gnd 0.598113f
C1976 a_n7636_8799.n51 gnd 0.263763f
C1977 a_n7636_8799.n52 gnd 0.011798f
C1978 a_n7636_8799.n53 gnd 0.051991f
C1979 a_n7636_8799.n54 gnd 0.051991f
C1980 a_n7636_8799.n55 gnd 0.051991f
C1981 a_n7636_8799.n56 gnd 0.011798f
C1982 a_n7636_8799.t85 gnd 0.598113f
C1983 a_n7636_8799.n57 gnd 0.264725f
C1984 a_n7636_8799.t115 gnd 0.598113f
C1985 a_n7636_8799.n58 gnd 0.264084f
C1986 a_n7636_8799.n59 gnd 0.051991f
C1987 a_n7636_8799.n60 gnd 0.051991f
C1988 a_n7636_8799.n61 gnd 0.051991f
C1989 a_n7636_8799.n62 gnd 0.267129f
C1990 a_n7636_8799.n63 gnd 0.011798f
C1991 a_n7636_8799.t73 gnd 0.598113f
C1992 a_n7636_8799.n64 gnd 0.264404f
C1993 a_n7636_8799.n65 gnd 0.051991f
C1994 a_n7636_8799.n66 gnd 0.051991f
C1995 a_n7636_8799.n67 gnd 0.051991f
C1996 a_n7636_8799.n68 gnd 0.011798f
C1997 a_n7636_8799.t37 gnd 0.598113f
C1998 a_n7636_8799.n69 gnd 0.267129f
C1999 a_n7636_8799.n70 gnd 0.011798f
C2000 a_n7636_8799.n71 gnd 0.051991f
C2001 a_n7636_8799.n72 gnd 0.051991f
C2002 a_n7636_8799.n73 gnd 0.051991f
C2003 a_n7636_8799.n74 gnd 0.264725f
C2004 a_n7636_8799.n75 gnd 0.011798f
C2005 a_n7636_8799.t136 gnd 0.598113f
C2006 a_n7636_8799.n76 gnd 0.267129f
C2007 a_n7636_8799.n77 gnd 0.051991f
C2008 a_n7636_8799.n78 gnd 0.051991f
C2009 a_n7636_8799.n79 gnd 0.051991f
C2010 a_n7636_8799.n80 gnd 0.263763f
C2011 a_n7636_8799.t67 gnd 0.598113f
C2012 a_n7636_8799.n81 gnd 0.265045f
C2013 a_n7636_8799.n82 gnd 0.011798f
C2014 a_n7636_8799.n83 gnd 0.051991f
C2015 a_n7636_8799.n84 gnd 0.051991f
C2016 a_n7636_8799.n85 gnd 0.051991f
C2017 a_n7636_8799.n86 gnd 0.011798f
C2018 a_n7636_8799.t46 gnd 0.598113f
C2019 a_n7636_8799.n87 gnd 0.263443f
C2020 a_n7636_8799.t47 gnd 0.598113f
C2021 a_n7636_8799.n88 gnd 0.26168f
C2022 a_n7636_8799.n89 gnd 0.294776f
C2023 a_n7636_8799.n90 gnd 0.051991f
C2024 a_n7636_8799.t146 gnd 0.598113f
C2025 a_n7636_8799.n91 gnd 0.267129f
C2026 a_n7636_8799.n92 gnd 0.051991f
C2027 a_n7636_8799.n93 gnd 0.011798f
C2028 a_n7636_8799.t64 gnd 0.598113f
C2029 a_n7636_8799.n94 gnd 0.051991f
C2030 a_n7636_8799.t79 gnd 0.598113f
C2031 a_n7636_8799.n95 gnd 0.264084f
C2032 a_n7636_8799.t106 gnd 0.598113f
C2033 a_n7636_8799.n96 gnd 0.051991f
C2034 a_n7636_8799.t124 gnd 0.598113f
C2035 a_n7636_8799.n97 gnd 0.264404f
C2036 a_n7636_8799.n98 gnd 0.051991f
C2037 a_n7636_8799.n99 gnd 0.011798f
C2038 a_n7636_8799.t82 gnd 0.598113f
C2039 a_n7636_8799.n100 gnd 0.051991f
C2040 a_n7636_8799.t94 gnd 0.598113f
C2041 a_n7636_8799.n101 gnd 0.267129f
C2042 a_n7636_8799.n102 gnd 0.051991f
C2043 a_n7636_8799.n103 gnd 0.011798f
C2044 a_n7636_8799.t130 gnd 0.598113f
C2045 a_n7636_8799.n104 gnd 0.164254f
C2046 a_n7636_8799.t155 gnd 0.598113f
C2047 a_n7636_8799.t151 gnd 0.609434f
C2048 a_n7636_8799.n105 gnd 0.250733f
C2049 a_n7636_8799.n106 gnd 0.263443f
C2050 a_n7636_8799.n107 gnd 0.011798f
C2051 a_n7636_8799.t98 gnd 0.598113f
C2052 a_n7636_8799.n108 gnd 0.267129f
C2053 a_n7636_8799.n109 gnd 0.051991f
C2054 a_n7636_8799.n110 gnd 0.051991f
C2055 a_n7636_8799.n111 gnd 0.051991f
C2056 a_n7636_8799.n112 gnd 0.265045f
C2057 a_n7636_8799.t148 gnd 0.598113f
C2058 a_n7636_8799.n113 gnd 0.263763f
C2059 a_n7636_8799.n114 gnd 0.011798f
C2060 a_n7636_8799.n115 gnd 0.051991f
C2061 a_n7636_8799.n116 gnd 0.051991f
C2062 a_n7636_8799.n117 gnd 0.051991f
C2063 a_n7636_8799.n118 gnd 0.011798f
C2064 a_n7636_8799.t95 gnd 0.598113f
C2065 a_n7636_8799.n119 gnd 0.264725f
C2066 a_n7636_8799.t128 gnd 0.598113f
C2067 a_n7636_8799.n120 gnd 0.264084f
C2068 a_n7636_8799.n121 gnd 0.051991f
C2069 a_n7636_8799.n122 gnd 0.051991f
C2070 a_n7636_8799.n123 gnd 0.051991f
C2071 a_n7636_8799.n124 gnd 0.267129f
C2072 a_n7636_8799.n125 gnd 0.011798f
C2073 a_n7636_8799.t83 gnd 0.598113f
C2074 a_n7636_8799.n126 gnd 0.264404f
C2075 a_n7636_8799.n127 gnd 0.051991f
C2076 a_n7636_8799.n128 gnd 0.051991f
C2077 a_n7636_8799.n129 gnd 0.051991f
C2078 a_n7636_8799.n130 gnd 0.011798f
C2079 a_n7636_8799.t48 gnd 0.598113f
C2080 a_n7636_8799.n131 gnd 0.267129f
C2081 a_n7636_8799.n132 gnd 0.011798f
C2082 a_n7636_8799.n133 gnd 0.051991f
C2083 a_n7636_8799.n134 gnd 0.051991f
C2084 a_n7636_8799.n135 gnd 0.051991f
C2085 a_n7636_8799.n136 gnd 0.264725f
C2086 a_n7636_8799.n137 gnd 0.011798f
C2087 a_n7636_8799.t152 gnd 0.598113f
C2088 a_n7636_8799.n138 gnd 0.267129f
C2089 a_n7636_8799.n139 gnd 0.051991f
C2090 a_n7636_8799.n140 gnd 0.051991f
C2091 a_n7636_8799.n141 gnd 0.051991f
C2092 a_n7636_8799.n142 gnd 0.263763f
C2093 a_n7636_8799.t78 gnd 0.598113f
C2094 a_n7636_8799.n143 gnd 0.265045f
C2095 a_n7636_8799.n144 gnd 0.011798f
C2096 a_n7636_8799.n145 gnd 0.051991f
C2097 a_n7636_8799.n146 gnd 0.051991f
C2098 a_n7636_8799.n147 gnd 0.051991f
C2099 a_n7636_8799.n148 gnd 0.011798f
C2100 a_n7636_8799.t58 gnd 0.598113f
C2101 a_n7636_8799.n149 gnd 0.263443f
C2102 a_n7636_8799.t60 gnd 0.598113f
C2103 a_n7636_8799.n150 gnd 0.26168f
C2104 a_n7636_8799.n151 gnd 0.129589f
C2105 a_n7636_8799.n152 gnd 0.89918f
C2106 a_n7636_8799.n153 gnd 0.051991f
C2107 a_n7636_8799.t101 gnd 0.598113f
C2108 a_n7636_8799.n154 gnd 0.267129f
C2109 a_n7636_8799.n155 gnd 0.051991f
C2110 a_n7636_8799.n156 gnd 0.011798f
C2111 a_n7636_8799.t125 gnd 0.598113f
C2112 a_n7636_8799.n157 gnd 0.051991f
C2113 a_n7636_8799.t43 gnd 0.598113f
C2114 a_n7636_8799.n158 gnd 0.264084f
C2115 a_n7636_8799.t108 gnd 0.598113f
C2116 a_n7636_8799.n159 gnd 0.051991f
C2117 a_n7636_8799.t147 gnd 0.598113f
C2118 a_n7636_8799.n160 gnd 0.264404f
C2119 a_n7636_8799.n161 gnd 0.051991f
C2120 a_n7636_8799.n162 gnd 0.011798f
C2121 a_n7636_8799.t142 gnd 0.598113f
C2122 a_n7636_8799.n163 gnd 0.051991f
C2123 a_n7636_8799.t55 gnd 0.598113f
C2124 a_n7636_8799.n164 gnd 0.267129f
C2125 a_n7636_8799.n165 gnd 0.051991f
C2126 a_n7636_8799.n166 gnd 0.011798f
C2127 a_n7636_8799.t80 gnd 0.598113f
C2128 a_n7636_8799.n167 gnd 0.164254f
C2129 a_n7636_8799.t91 gnd 0.598113f
C2130 a_n7636_8799.t113 gnd 0.609434f
C2131 a_n7636_8799.n168 gnd 0.250733f
C2132 a_n7636_8799.n169 gnd 0.263443f
C2133 a_n7636_8799.n170 gnd 0.011798f
C2134 a_n7636_8799.t129 gnd 0.598113f
C2135 a_n7636_8799.n171 gnd 0.267129f
C2136 a_n7636_8799.n172 gnd 0.051991f
C2137 a_n7636_8799.n173 gnd 0.051991f
C2138 a_n7636_8799.n174 gnd 0.051991f
C2139 a_n7636_8799.n175 gnd 0.265045f
C2140 a_n7636_8799.t139 gnd 0.598113f
C2141 a_n7636_8799.n176 gnd 0.263763f
C2142 a_n7636_8799.n177 gnd 0.011798f
C2143 a_n7636_8799.n178 gnd 0.051991f
C2144 a_n7636_8799.n179 gnd 0.051991f
C2145 a_n7636_8799.n180 gnd 0.051991f
C2146 a_n7636_8799.n181 gnd 0.011798f
C2147 a_n7636_8799.t38 gnd 0.598113f
C2148 a_n7636_8799.n182 gnd 0.264725f
C2149 a_n7636_8799.t99 gnd 0.598113f
C2150 a_n7636_8799.n183 gnd 0.264084f
C2151 a_n7636_8799.n184 gnd 0.051991f
C2152 a_n7636_8799.n185 gnd 0.051991f
C2153 a_n7636_8799.n186 gnd 0.051991f
C2154 a_n7636_8799.n187 gnd 0.267129f
C2155 a_n7636_8799.n188 gnd 0.011798f
C2156 a_n7636_8799.t116 gnd 0.598113f
C2157 a_n7636_8799.n189 gnd 0.264404f
C2158 a_n7636_8799.n190 gnd 0.051991f
C2159 a_n7636_8799.n191 gnd 0.051991f
C2160 a_n7636_8799.n192 gnd 0.051991f
C2161 a_n7636_8799.n193 gnd 0.011798f
C2162 a_n7636_8799.t92 gnd 0.598113f
C2163 a_n7636_8799.n194 gnd 0.267129f
C2164 a_n7636_8799.n195 gnd 0.011798f
C2165 a_n7636_8799.n196 gnd 0.051991f
C2166 a_n7636_8799.n197 gnd 0.051991f
C2167 a_n7636_8799.n198 gnd 0.051991f
C2168 a_n7636_8799.n199 gnd 0.264725f
C2169 a_n7636_8799.n200 gnd 0.011798f
C2170 a_n7636_8799.t62 gnd 0.598113f
C2171 a_n7636_8799.n201 gnd 0.267129f
C2172 a_n7636_8799.n202 gnd 0.051991f
C2173 a_n7636_8799.n203 gnd 0.051991f
C2174 a_n7636_8799.n204 gnd 0.051991f
C2175 a_n7636_8799.n205 gnd 0.263763f
C2176 a_n7636_8799.t71 gnd 0.598113f
C2177 a_n7636_8799.n206 gnd 0.265045f
C2178 a_n7636_8799.n207 gnd 0.011798f
C2179 a_n7636_8799.n208 gnd 0.051991f
C2180 a_n7636_8799.n209 gnd 0.051991f
C2181 a_n7636_8799.n210 gnd 0.051991f
C2182 a_n7636_8799.n211 gnd 0.011798f
C2183 a_n7636_8799.t51 gnd 0.598113f
C2184 a_n7636_8799.n212 gnd 0.263443f
C2185 a_n7636_8799.t153 gnd 0.598113f
C2186 a_n7636_8799.n213 gnd 0.26168f
C2187 a_n7636_8799.n214 gnd 0.129589f
C2188 a_n7636_8799.n215 gnd 1.54004f
C2189 a_n7636_8799.n216 gnd 0.051991f
C2190 a_n7636_8799.t87 gnd 0.598113f
C2191 a_n7636_8799.t86 gnd 0.598113f
C2192 a_n7636_8799.t59 gnd 0.598113f
C2193 a_n7636_8799.n217 gnd 0.267129f
C2194 a_n7636_8799.n218 gnd 0.051991f
C2195 a_n7636_8799.t135 gnd 0.598113f
C2196 a_n7636_8799.t90 gnd 0.598113f
C2197 a_n7636_8799.n219 gnd 0.051991f
C2198 a_n7636_8799.t66 gnd 0.598113f
C2199 a_n7636_8799.n220 gnd 0.267129f
C2200 a_n7636_8799.n221 gnd 0.051991f
C2201 a_n7636_8799.t141 gnd 0.598113f
C2202 a_n7636_8799.t107 gnd 0.598113f
C2203 a_n7636_8799.n222 gnd 0.051991f
C2204 a_n7636_8799.t105 gnd 0.598113f
C2205 a_n7636_8799.n223 gnd 0.267129f
C2206 a_n7636_8799.n224 gnd 0.051991f
C2207 a_n7636_8799.t40 gnd 0.598113f
C2208 a_n7636_8799.t111 gnd 0.598113f
C2209 a_n7636_8799.n225 gnd 0.051991f
C2210 a_n7636_8799.t110 gnd 0.598113f
C2211 a_n7636_8799.n226 gnd 0.267129f
C2212 a_n7636_8799.n227 gnd 0.051991f
C2213 a_n7636_8799.t42 gnd 0.598113f
C2214 a_n7636_8799.t41 gnd 0.598113f
C2215 a_n7636_8799.n228 gnd 0.051991f
C2216 a_n7636_8799.t127 gnd 0.598113f
C2217 a_n7636_8799.n229 gnd 0.267129f
C2218 a_n7636_8799.n230 gnd 0.051991f
C2219 a_n7636_8799.t61 gnd 0.598113f
C2220 a_n7636_8799.t44 gnd 0.598113f
C2221 a_n7636_8799.n231 gnd 0.051991f
C2222 a_n7636_8799.t131 gnd 0.598113f
C2223 a_n7636_8799.n232 gnd 0.267129f
C2224 a_n7636_8799.t65 gnd 0.609434f
C2225 a_n7636_8799.n233 gnd 0.250733f
C2226 a_n7636_8799.t89 gnd 0.598113f
C2227 a_n7636_8799.n234 gnd 0.263443f
C2228 a_n7636_8799.n235 gnd 0.011798f
C2229 a_n7636_8799.n236 gnd 0.164254f
C2230 a_n7636_8799.n237 gnd 0.051991f
C2231 a_n7636_8799.n238 gnd 0.051991f
C2232 a_n7636_8799.n239 gnd 0.011798f
C2233 a_n7636_8799.n240 gnd 0.265045f
C2234 a_n7636_8799.n241 gnd 0.263763f
C2235 a_n7636_8799.n242 gnd 0.011798f
C2236 a_n7636_8799.n243 gnd 0.051991f
C2237 a_n7636_8799.n244 gnd 0.051991f
C2238 a_n7636_8799.n245 gnd 0.051991f
C2239 a_n7636_8799.n246 gnd 0.011798f
C2240 a_n7636_8799.n247 gnd 0.264725f
C2241 a_n7636_8799.n248 gnd 0.264084f
C2242 a_n7636_8799.n249 gnd 0.011798f
C2243 a_n7636_8799.n250 gnd 0.051991f
C2244 a_n7636_8799.n251 gnd 0.051991f
C2245 a_n7636_8799.n252 gnd 0.051991f
C2246 a_n7636_8799.n253 gnd 0.011798f
C2247 a_n7636_8799.n254 gnd 0.264404f
C2248 a_n7636_8799.n255 gnd 0.264404f
C2249 a_n7636_8799.n256 gnd 0.011798f
C2250 a_n7636_8799.n257 gnd 0.051991f
C2251 a_n7636_8799.n258 gnd 0.051991f
C2252 a_n7636_8799.n259 gnd 0.051991f
C2253 a_n7636_8799.n260 gnd 0.011798f
C2254 a_n7636_8799.n261 gnd 0.264084f
C2255 a_n7636_8799.n262 gnd 0.264725f
C2256 a_n7636_8799.n263 gnd 0.011798f
C2257 a_n7636_8799.n264 gnd 0.051991f
C2258 a_n7636_8799.n265 gnd 0.051991f
C2259 a_n7636_8799.n266 gnd 0.051991f
C2260 a_n7636_8799.n267 gnd 0.011798f
C2261 a_n7636_8799.n268 gnd 0.263763f
C2262 a_n7636_8799.n269 gnd 0.265045f
C2263 a_n7636_8799.n270 gnd 0.011798f
C2264 a_n7636_8799.n271 gnd 0.051991f
C2265 a_n7636_8799.n272 gnd 0.051991f
C2266 a_n7636_8799.n273 gnd 0.051991f
C2267 a_n7636_8799.n274 gnd 0.011798f
C2268 a_n7636_8799.n275 gnd 0.263443f
C2269 a_n7636_8799.n276 gnd 0.26168f
C2270 a_n7636_8799.n277 gnd 0.294776f
C2271 a_n7636_8799.n278 gnd 0.051991f
C2272 a_n7636_8799.t97 gnd 0.598113f
C2273 a_n7636_8799.t96 gnd 0.598113f
C2274 a_n7636_8799.t74 gnd 0.598113f
C2275 a_n7636_8799.n279 gnd 0.267129f
C2276 a_n7636_8799.n280 gnd 0.051991f
C2277 a_n7636_8799.t150 gnd 0.598113f
C2278 a_n7636_8799.t104 gnd 0.598113f
C2279 a_n7636_8799.n281 gnd 0.051991f
C2280 a_n7636_8799.t76 gnd 0.598113f
C2281 a_n7636_8799.n282 gnd 0.267129f
C2282 a_n7636_8799.n283 gnd 0.051991f
C2283 a_n7636_8799.t36 gnd 0.598113f
C2284 a_n7636_8799.t120 gnd 0.598113f
C2285 a_n7636_8799.n284 gnd 0.051991f
C2286 a_n7636_8799.t119 gnd 0.598113f
C2287 a_n7636_8799.n285 gnd 0.267129f
C2288 a_n7636_8799.n286 gnd 0.051991f
C2289 a_n7636_8799.t50 gnd 0.598113f
C2290 a_n7636_8799.t123 gnd 0.598113f
C2291 a_n7636_8799.n287 gnd 0.051991f
C2292 a_n7636_8799.t122 gnd 0.598113f
C2293 a_n7636_8799.n288 gnd 0.267129f
C2294 a_n7636_8799.n289 gnd 0.051991f
C2295 a_n7636_8799.t54 gnd 0.598113f
C2296 a_n7636_8799.t53 gnd 0.598113f
C2297 a_n7636_8799.n290 gnd 0.051991f
C2298 a_n7636_8799.t144 gnd 0.598113f
C2299 a_n7636_8799.n291 gnd 0.267129f
C2300 a_n7636_8799.n292 gnd 0.051991f
C2301 a_n7636_8799.t75 gnd 0.598113f
C2302 a_n7636_8799.t57 gnd 0.598113f
C2303 a_n7636_8799.n293 gnd 0.051991f
C2304 a_n7636_8799.t145 gnd 0.598113f
C2305 a_n7636_8799.n294 gnd 0.267129f
C2306 a_n7636_8799.t77 gnd 0.609434f
C2307 a_n7636_8799.n295 gnd 0.250733f
C2308 a_n7636_8799.t103 gnd 0.598113f
C2309 a_n7636_8799.n296 gnd 0.263443f
C2310 a_n7636_8799.n297 gnd 0.011798f
C2311 a_n7636_8799.n298 gnd 0.164254f
C2312 a_n7636_8799.n299 gnd 0.051991f
C2313 a_n7636_8799.n300 gnd 0.051991f
C2314 a_n7636_8799.n301 gnd 0.011798f
C2315 a_n7636_8799.n302 gnd 0.265045f
C2316 a_n7636_8799.n303 gnd 0.263763f
C2317 a_n7636_8799.n304 gnd 0.011798f
C2318 a_n7636_8799.n305 gnd 0.051991f
C2319 a_n7636_8799.n306 gnd 0.051991f
C2320 a_n7636_8799.n307 gnd 0.051991f
C2321 a_n7636_8799.n308 gnd 0.011798f
C2322 a_n7636_8799.n309 gnd 0.264725f
C2323 a_n7636_8799.n310 gnd 0.264084f
C2324 a_n7636_8799.n311 gnd 0.011798f
C2325 a_n7636_8799.n312 gnd 0.051991f
C2326 a_n7636_8799.n313 gnd 0.051991f
C2327 a_n7636_8799.n314 gnd 0.051991f
C2328 a_n7636_8799.n315 gnd 0.011798f
C2329 a_n7636_8799.n316 gnd 0.264404f
C2330 a_n7636_8799.n317 gnd 0.264404f
C2331 a_n7636_8799.n318 gnd 0.011798f
C2332 a_n7636_8799.n319 gnd 0.051991f
C2333 a_n7636_8799.n320 gnd 0.051991f
C2334 a_n7636_8799.n321 gnd 0.051991f
C2335 a_n7636_8799.n322 gnd 0.011798f
C2336 a_n7636_8799.n323 gnd 0.264084f
C2337 a_n7636_8799.n324 gnd 0.264725f
C2338 a_n7636_8799.n325 gnd 0.011798f
C2339 a_n7636_8799.n326 gnd 0.051991f
C2340 a_n7636_8799.n327 gnd 0.051991f
C2341 a_n7636_8799.n328 gnd 0.051991f
C2342 a_n7636_8799.n329 gnd 0.011798f
C2343 a_n7636_8799.n330 gnd 0.263763f
C2344 a_n7636_8799.n331 gnd 0.265045f
C2345 a_n7636_8799.n332 gnd 0.011798f
C2346 a_n7636_8799.n333 gnd 0.051991f
C2347 a_n7636_8799.n334 gnd 0.051991f
C2348 a_n7636_8799.n335 gnd 0.051991f
C2349 a_n7636_8799.n336 gnd 0.011798f
C2350 a_n7636_8799.n337 gnd 0.263443f
C2351 a_n7636_8799.n338 gnd 0.26168f
C2352 a_n7636_8799.n339 gnd 0.129589f
C2353 a_n7636_8799.n340 gnd 0.89918f
C2354 a_n7636_8799.n341 gnd 0.051991f
C2355 a_n7636_8799.t154 gnd 0.598113f
C2356 a_n7636_8799.t52 gnd 0.598113f
C2357 a_n7636_8799.t102 gnd 0.598113f
C2358 a_n7636_8799.n342 gnd 0.267129f
C2359 a_n7636_8799.n343 gnd 0.051991f
C2360 a_n7636_8799.t39 gnd 0.598113f
C2361 a_n7636_8799.t126 gnd 0.598113f
C2362 a_n7636_8799.n344 gnd 0.051991f
C2363 a_n7636_8799.t63 gnd 0.598113f
C2364 a_n7636_8799.n345 gnd 0.267129f
C2365 a_n7636_8799.n346 gnd 0.051991f
C2366 a_n7636_8799.t109 gnd 0.598113f
C2367 a_n7636_8799.t45 gnd 0.598113f
C2368 a_n7636_8799.n347 gnd 0.051991f
C2369 a_n7636_8799.t69 gnd 0.598113f
C2370 a_n7636_8799.n348 gnd 0.267129f
C2371 a_n7636_8799.n349 gnd 0.051991f
C2372 a_n7636_8799.t149 gnd 0.598113f
C2373 a_n7636_8799.t118 gnd 0.598113f
C2374 a_n7636_8799.n350 gnd 0.051991f
C2375 a_n7636_8799.t143 gnd 0.598113f
C2376 a_n7636_8799.n351 gnd 0.267129f
C2377 a_n7636_8799.n352 gnd 0.051991f
C2378 a_n7636_8799.t100 gnd 0.598113f
C2379 a_n7636_8799.t121 gnd 0.598113f
C2380 a_n7636_8799.n353 gnd 0.051991f
C2381 a_n7636_8799.t56 gnd 0.598113f
C2382 a_n7636_8799.n354 gnd 0.267129f
C2383 a_n7636_8799.n355 gnd 0.051991f
C2384 a_n7636_8799.t140 gnd 0.598113f
C2385 a_n7636_8799.t81 gnd 0.598113f
C2386 a_n7636_8799.n356 gnd 0.051991f
C2387 a_n7636_8799.t132 gnd 0.598113f
C2388 a_n7636_8799.n357 gnd 0.267129f
C2389 a_n7636_8799.t114 gnd 0.609434f
C2390 a_n7636_8799.n358 gnd 0.250733f
C2391 a_n7636_8799.t68 gnd 0.598113f
C2392 a_n7636_8799.n359 gnd 0.263443f
C2393 a_n7636_8799.n360 gnd 0.011798f
C2394 a_n7636_8799.n361 gnd 0.164254f
C2395 a_n7636_8799.n362 gnd 0.051991f
C2396 a_n7636_8799.n363 gnd 0.051991f
C2397 a_n7636_8799.n364 gnd 0.011798f
C2398 a_n7636_8799.n365 gnd 0.265045f
C2399 a_n7636_8799.n366 gnd 0.263763f
C2400 a_n7636_8799.n367 gnd 0.011798f
C2401 a_n7636_8799.n368 gnd 0.051991f
C2402 a_n7636_8799.n369 gnd 0.051991f
C2403 a_n7636_8799.n370 gnd 0.051991f
C2404 a_n7636_8799.n371 gnd 0.011798f
C2405 a_n7636_8799.n372 gnd 0.264725f
C2406 a_n7636_8799.n373 gnd 0.264084f
C2407 a_n7636_8799.n374 gnd 0.011798f
C2408 a_n7636_8799.n375 gnd 0.051991f
C2409 a_n7636_8799.n376 gnd 0.051991f
C2410 a_n7636_8799.n377 gnd 0.051991f
C2411 a_n7636_8799.n378 gnd 0.011798f
C2412 a_n7636_8799.n379 gnd 0.264404f
C2413 a_n7636_8799.n380 gnd 0.264404f
C2414 a_n7636_8799.n381 gnd 0.011798f
C2415 a_n7636_8799.n382 gnd 0.051991f
C2416 a_n7636_8799.n383 gnd 0.051991f
C2417 a_n7636_8799.n384 gnd 0.051991f
C2418 a_n7636_8799.n385 gnd 0.011798f
C2419 a_n7636_8799.n386 gnd 0.264084f
C2420 a_n7636_8799.n387 gnd 0.264725f
C2421 a_n7636_8799.n388 gnd 0.011798f
C2422 a_n7636_8799.n389 gnd 0.051991f
C2423 a_n7636_8799.n390 gnd 0.051991f
C2424 a_n7636_8799.n391 gnd 0.051991f
C2425 a_n7636_8799.n392 gnd 0.011798f
C2426 a_n7636_8799.n393 gnd 0.263763f
C2427 a_n7636_8799.n394 gnd 0.265045f
C2428 a_n7636_8799.n395 gnd 0.011798f
C2429 a_n7636_8799.n396 gnd 0.051991f
C2430 a_n7636_8799.n397 gnd 0.051991f
C2431 a_n7636_8799.n398 gnd 0.051991f
C2432 a_n7636_8799.n399 gnd 0.011798f
C2433 a_n7636_8799.n400 gnd 0.263443f
C2434 a_n7636_8799.n401 gnd 0.26168f
C2435 a_n7636_8799.n402 gnd 0.129589f
C2436 a_n7636_8799.n403 gnd 1.08666f
C2437 a_n7636_8799.n404 gnd 12.216201f
C2438 a_n7636_8799.n405 gnd 4.37732f
C2439 a_n7636_8799.n406 gnd 5.67932f
C2440 a_n7636_8799.t3 gnd 0.144247f
C2441 a_n7636_8799.t2 gnd 0.144247f
C2442 a_n7636_8799.n407 gnd 1.13582f
C2443 a_n7636_8799.n408 gnd 3.01156f
C2444 a_n7636_8799.t5 gnd 0.144247f
C2445 a_n7636_8799.t10 gnd 0.144247f
C2446 a_n7636_8799.n409 gnd 1.13769f
C2447 a_n7636_8799.n410 gnd 1.02096f
C2448 a_n7636_8799.n411 gnd 1.13582f
C2449 a_n7636_8799.t11 gnd 0.144247f
C2450 a_n3827_n3924.n0 gnd 2.31453f
C2451 a_n3827_n3924.n1 gnd 1.78938f
C2452 a_n3827_n3924.n2 gnd 2.10086f
C2453 a_n3827_n3924.n3 gnd 2.31452f
C2454 a_n3827_n3924.n4 gnd 1.56597f
C2455 a_n3827_n3924.n5 gnd 1.73104f
C2456 a_n3827_n3924.n6 gnd 1.73104f
C2457 a_n3827_n3924.n7 gnd 1.73104f
C2458 a_n3827_n3924.n8 gnd 2.08302f
C2459 a_n3827_n3924.n9 gnd 0.78335f
C2460 a_n3827_n3924.n10 gnd 1.31751f
C2461 a_n3827_n3924.n11 gnd 0.783353f
C2462 a_n3827_n3924.n12 gnd 1.00603f
C2463 a_n3827_n3924.t14 gnd 0.095164f
C2464 a_n3827_n3924.t8 gnd 0.095164f
C2465 a_n3827_n3924.t6 gnd 0.095164f
C2466 a_n3827_n3924.n13 gnd 0.777219f
C2467 a_n3827_n3924.t43 gnd 0.989053f
C2468 a_n3827_n3924.t31 gnd 0.095164f
C2469 a_n3827_n3924.t39 gnd 0.095164f
C2470 a_n3827_n3924.n14 gnd 0.777221f
C2471 a_n3827_n3924.t50 gnd 0.095164f
C2472 a_n3827_n3924.t51 gnd 0.095164f
C2473 a_n3827_n3924.n15 gnd 0.777221f
C2474 a_n3827_n3924.t34 gnd 0.095164f
C2475 a_n3827_n3924.t48 gnd 0.095164f
C2476 a_n3827_n3924.n16 gnd 0.777221f
C2477 a_n3827_n3924.t38 gnd 0.095164f
C2478 a_n3827_n3924.t49 gnd 0.095164f
C2479 a_n3827_n3924.n17 gnd 0.777221f
C2480 a_n3827_n3924.t42 gnd 0.095164f
C2481 a_n3827_n3924.t37 gnd 0.095164f
C2482 a_n3827_n3924.n18 gnd 0.777221f
C2483 a_n3827_n3924.t46 gnd 0.989057f
C2484 a_n3827_n3924.t1 gnd 0.989057f
C2485 a_n3827_n3924.t19 gnd 0.095164f
C2486 a_n3827_n3924.t12 gnd 0.095164f
C2487 a_n3827_n3924.n19 gnd 0.777221f
C2488 a_n3827_n3924.t29 gnd 0.095164f
C2489 a_n3827_n3924.t22 gnd 0.095164f
C2490 a_n3827_n3924.n20 gnd 0.777221f
C2491 a_n3827_n3924.t57 gnd 0.095164f
C2492 a_n3827_n3924.t30 gnd 0.095164f
C2493 a_n3827_n3924.n21 gnd 0.777221f
C2494 a_n3827_n3924.t20 gnd 0.095164f
C2495 a_n3827_n3924.t15 gnd 0.095164f
C2496 a_n3827_n3924.n22 gnd 0.777221f
C2497 a_n3827_n3924.t11 gnd 0.095164f
C2498 a_n3827_n3924.t27 gnd 0.095164f
C2499 a_n3827_n3924.n23 gnd 0.777221f
C2500 a_n3827_n3924.t10 gnd 0.989057f
C2501 a_n3827_n3924.t4 gnd 0.095164f
C2502 a_n3827_n3924.t7 gnd 0.095164f
C2503 a_n3827_n3924.n24 gnd 0.777219f
C2504 a_n3827_n3924.t24 gnd 0.989053f
C2505 a_n3827_n3924.t47 gnd 0.989053f
C2506 a_n3827_n3924.t32 gnd 0.095164f
C2507 a_n3827_n3924.t52 gnd 0.095164f
C2508 a_n3827_n3924.n25 gnd 0.777219f
C2509 a_n3827_n3924.t33 gnd 0.095164f
C2510 a_n3827_n3924.t40 gnd 0.095164f
C2511 a_n3827_n3924.n26 gnd 0.777219f
C2512 a_n3827_n3924.t54 gnd 0.095164f
C2513 a_n3827_n3924.t36 gnd 0.095164f
C2514 a_n3827_n3924.n27 gnd 0.777219f
C2515 a_n3827_n3924.t45 gnd 0.095164f
C2516 a_n3827_n3924.t53 gnd 0.095164f
C2517 a_n3827_n3924.n28 gnd 0.777219f
C2518 a_n3827_n3924.t44 gnd 0.095164f
C2519 a_n3827_n3924.t41 gnd 0.095164f
C2520 a_n3827_n3924.n29 gnd 0.777219f
C2521 a_n3827_n3924.t35 gnd 0.989053f
C2522 a_n3827_n3924.n30 gnd 0.897154f
C2523 a_n3827_n3924.t23 gnd 1.23041f
C2524 a_n3827_n3924.t28 gnd 1.22888f
C2525 a_n3827_n3924.t13 gnd 1.22888f
C2526 a_n3827_n3924.t16 gnd 1.22888f
C2527 a_n3827_n3924.t56 gnd 1.22888f
C2528 a_n3827_n3924.t5 gnd 1.22888f
C2529 a_n3827_n3924.t18 gnd 1.22888f
C2530 a_n3827_n3924.t3 gnd 1.22888f
C2531 a_n3827_n3924.t55 gnd 1.22888f
C2532 a_n3827_n3924.t9 gnd 1.2292f
C2533 a_n3827_n3924.n31 gnd 0.897154f
C2534 a_n3827_n3924.t25 gnd 0.989053f
C2535 a_n3827_n3924.t17 gnd 0.095164f
C2536 a_n3827_n3924.t26 gnd 0.095164f
C2537 a_n3827_n3924.n32 gnd 0.777219f
C2538 a_n3827_n3924.t21 gnd 0.095164f
C2539 a_n3827_n3924.t2 gnd 0.095164f
C2540 a_n3827_n3924.n33 gnd 0.777219f
C2541 a_n3827_n3924.n34 gnd 0.777216f
C2542 a_n3827_n3924.t0 gnd 0.095164f
C2543 plus.n0 gnd 0.022575f
C2544 plus.t20 gnd 0.410529f
C2545 plus.t23 gnd 0.379592f
C2546 plus.n1 gnd 0.153524f
C2547 plus.n2 gnd 0.022575f
C2548 plus.t6 gnd 0.379592f
C2549 plus.n3 gnd 0.019291f
C2550 plus.n4 gnd 0.022575f
C2551 plus.t12 gnd 0.379592f
C2552 plus.t8 gnd 0.379592f
C2553 plus.n5 gnd 0.153524f
C2554 plus.n6 gnd 0.022575f
C2555 plus.t7 gnd 0.379592f
C2556 plus.n7 gnd 0.153524f
C2557 plus.n8 gnd 0.022575f
C2558 plus.t19 gnd 0.379592f
C2559 plus.n9 gnd 0.018348f
C2560 plus.n10 gnd 0.022575f
C2561 plus.t18 gnd 0.379592f
C2562 plus.t27 gnd 0.379592f
C2563 plus.n11 gnd 0.153524f
C2564 plus.n12 gnd 0.022575f
C2565 plus.t25 gnd 0.379592f
C2566 plus.n13 gnd 0.153524f
C2567 plus.n14 gnd 0.095805f
C2568 plus.t9 gnd 0.379592f
C2569 plus.t14 gnd 0.424642f
C2570 plus.n15 gnd 0.179485f
C2571 plus.n16 gnd 0.175814f
C2572 plus.n17 gnd 0.028926f
C2573 plus.n18 gnd 0.025546f
C2574 plus.n19 gnd 0.022575f
C2575 plus.n20 gnd 0.022575f
C2576 plus.n21 gnd 0.026977f
C2577 plus.n22 gnd 0.019291f
C2578 plus.n23 gnd 0.029401f
C2579 plus.n24 gnd 0.022575f
C2580 plus.n25 gnd 0.022575f
C2581 plus.n26 gnd 0.028081f
C2582 plus.n27 gnd 0.026391f
C2583 plus.n28 gnd 0.153524f
C2584 plus.n29 gnd 0.028279f
C2585 plus.n30 gnd 0.022575f
C2586 plus.n31 gnd 0.022575f
C2587 plus.n32 gnd 0.022575f
C2588 plus.n33 gnd 0.029042f
C2589 plus.n34 gnd 0.153524f
C2590 plus.n35 gnd 0.027236f
C2591 plus.n36 gnd 0.027236f
C2592 plus.n37 gnd 0.022575f
C2593 plus.n38 gnd 0.022575f
C2594 plus.n39 gnd 0.029042f
C2595 plus.n40 gnd 0.018348f
C2596 plus.n41 gnd 0.028279f
C2597 plus.n42 gnd 0.022575f
C2598 plus.n43 gnd 0.022575f
C2599 plus.n44 gnd 0.026391f
C2600 plus.n45 gnd 0.028081f
C2601 plus.n46 gnd 0.153524f
C2602 plus.n47 gnd 0.029401f
C2603 plus.n48 gnd 0.022575f
C2604 plus.n49 gnd 0.022575f
C2605 plus.n50 gnd 0.022575f
C2606 plus.n51 gnd 0.026977f
C2607 plus.n52 gnd 0.153524f
C2608 plus.n53 gnd 0.025546f
C2609 plus.n54 gnd 0.028926f
C2610 plus.n55 gnd 0.022575f
C2611 plus.n56 gnd 0.022575f
C2612 plus.n57 gnd 0.02945f
C2613 plus.n58 gnd 0.008204f
C2614 plus.n59 gnd 0.177755f
C2615 plus.n60 gnd 0.258648f
C2616 plus.n61 gnd 0.022575f
C2617 plus.t28 gnd 0.379592f
C2618 plus.n62 gnd 0.153524f
C2619 plus.n63 gnd 0.022575f
C2620 plus.t26 gnd 0.379592f
C2621 plus.n64 gnd 0.019291f
C2622 plus.n65 gnd 0.022575f
C2623 plus.t10 gnd 0.379592f
C2624 plus.t15 gnd 0.379592f
C2625 plus.n66 gnd 0.153524f
C2626 plus.n67 gnd 0.022575f
C2627 plus.t13 gnd 0.379592f
C2628 plus.n68 gnd 0.153524f
C2629 plus.n69 gnd 0.022575f
C2630 plus.t17 gnd 0.379592f
C2631 plus.n70 gnd 0.018348f
C2632 plus.n71 gnd 0.022575f
C2633 plus.t16 gnd 0.379592f
C2634 plus.t21 gnd 0.379592f
C2635 plus.n72 gnd 0.153524f
C2636 plus.n73 gnd 0.022575f
C2637 plus.t22 gnd 0.379592f
C2638 plus.n74 gnd 0.153524f
C2639 plus.n75 gnd 0.095805f
C2640 plus.t5 gnd 0.379592f
C2641 plus.t11 gnd 0.424642f
C2642 plus.n76 gnd 0.179485f
C2643 plus.n77 gnd 0.175814f
C2644 plus.n78 gnd 0.028926f
C2645 plus.n79 gnd 0.025546f
C2646 plus.n80 gnd 0.022575f
C2647 plus.n81 gnd 0.022575f
C2648 plus.n82 gnd 0.026977f
C2649 plus.n83 gnd 0.019291f
C2650 plus.n84 gnd 0.029401f
C2651 plus.n85 gnd 0.022575f
C2652 plus.n86 gnd 0.022575f
C2653 plus.n87 gnd 0.028081f
C2654 plus.n88 gnd 0.026391f
C2655 plus.n89 gnd 0.153524f
C2656 plus.n90 gnd 0.028279f
C2657 plus.n91 gnd 0.022575f
C2658 plus.n92 gnd 0.022575f
C2659 plus.n93 gnd 0.022575f
C2660 plus.n94 gnd 0.029042f
C2661 plus.n95 gnd 0.153524f
C2662 plus.n96 gnd 0.027236f
C2663 plus.n97 gnd 0.027236f
C2664 plus.n98 gnd 0.022575f
C2665 plus.n99 gnd 0.022575f
C2666 plus.n100 gnd 0.029042f
C2667 plus.n101 gnd 0.018348f
C2668 plus.n102 gnd 0.028279f
C2669 plus.n103 gnd 0.022575f
C2670 plus.n104 gnd 0.022575f
C2671 plus.n105 gnd 0.026391f
C2672 plus.n106 gnd 0.028081f
C2673 plus.n107 gnd 0.153524f
C2674 plus.n108 gnd 0.029401f
C2675 plus.n109 gnd 0.022575f
C2676 plus.n110 gnd 0.022575f
C2677 plus.n111 gnd 0.022575f
C2678 plus.n112 gnd 0.026977f
C2679 plus.n113 gnd 0.153524f
C2680 plus.n114 gnd 0.025546f
C2681 plus.n115 gnd 0.028926f
C2682 plus.n116 gnd 0.022575f
C2683 plus.n117 gnd 0.022575f
C2684 plus.n118 gnd 0.02945f
C2685 plus.n119 gnd 0.008204f
C2686 plus.t24 gnd 0.410529f
C2687 plus.n120 gnd 0.177755f
C2688 plus.n121 gnd 0.814491f
C2689 plus.n122 gnd 1.20072f
C2690 plus.t1 gnd 0.038971f
C2691 plus.t2 gnd 0.006959f
C2692 plus.t4 gnd 0.006959f
C2693 plus.n123 gnd 0.02257f
C2694 plus.n124 gnd 0.175211f
C2695 plus.t3 gnd 0.006959f
C2696 plus.t0 gnd 0.006959f
C2697 plus.n125 gnd 0.02257f
C2698 plus.n126 gnd 0.131517f
C2699 plus.n127 gnd 3.2133f
C2700 outputibias.t10 gnd 0.11477f
C2701 outputibias.t8 gnd 0.115567f
C2702 outputibias.n0 gnd 0.130108f
C2703 outputibias.n1 gnd 0.001372f
C2704 outputibias.n2 gnd 9.76e-19
C2705 outputibias.n3 gnd 5.24e-19
C2706 outputibias.n4 gnd 0.001239f
C2707 outputibias.n5 gnd 5.55e-19
C2708 outputibias.n6 gnd 9.76e-19
C2709 outputibias.n7 gnd 5.24e-19
C2710 outputibias.n8 gnd 0.001239f
C2711 outputibias.n9 gnd 5.55e-19
C2712 outputibias.n10 gnd 0.004176f
C2713 outputibias.t5 gnd 0.00202f
C2714 outputibias.n11 gnd 9.3e-19
C2715 outputibias.n12 gnd 7.32e-19
C2716 outputibias.n13 gnd 5.24e-19
C2717 outputibias.n14 gnd 0.02322f
C2718 outputibias.n15 gnd 9.76e-19
C2719 outputibias.n16 gnd 5.24e-19
C2720 outputibias.n17 gnd 5.55e-19
C2721 outputibias.n18 gnd 0.001239f
C2722 outputibias.n19 gnd 0.001239f
C2723 outputibias.n20 gnd 5.55e-19
C2724 outputibias.n21 gnd 5.24e-19
C2725 outputibias.n22 gnd 9.76e-19
C2726 outputibias.n23 gnd 9.76e-19
C2727 outputibias.n24 gnd 5.24e-19
C2728 outputibias.n25 gnd 5.55e-19
C2729 outputibias.n26 gnd 0.001239f
C2730 outputibias.n27 gnd 0.002683f
C2731 outputibias.n28 gnd 5.55e-19
C2732 outputibias.n29 gnd 5.24e-19
C2733 outputibias.n30 gnd 0.002256f
C2734 outputibias.n31 gnd 0.005781f
C2735 outputibias.n32 gnd 0.001372f
C2736 outputibias.n33 gnd 9.76e-19
C2737 outputibias.n34 gnd 5.24e-19
C2738 outputibias.n35 gnd 0.001239f
C2739 outputibias.n36 gnd 5.55e-19
C2740 outputibias.n37 gnd 9.76e-19
C2741 outputibias.n38 gnd 5.24e-19
C2742 outputibias.n39 gnd 0.001239f
C2743 outputibias.n40 gnd 5.55e-19
C2744 outputibias.n41 gnd 0.004176f
C2745 outputibias.t3 gnd 0.00202f
C2746 outputibias.n42 gnd 9.3e-19
C2747 outputibias.n43 gnd 7.32e-19
C2748 outputibias.n44 gnd 5.24e-19
C2749 outputibias.n45 gnd 0.02322f
C2750 outputibias.n46 gnd 9.76e-19
C2751 outputibias.n47 gnd 5.24e-19
C2752 outputibias.n48 gnd 5.55e-19
C2753 outputibias.n49 gnd 0.001239f
C2754 outputibias.n50 gnd 0.001239f
C2755 outputibias.n51 gnd 5.55e-19
C2756 outputibias.n52 gnd 5.24e-19
C2757 outputibias.n53 gnd 9.76e-19
C2758 outputibias.n54 gnd 9.76e-19
C2759 outputibias.n55 gnd 5.24e-19
C2760 outputibias.n56 gnd 5.55e-19
C2761 outputibias.n57 gnd 0.001239f
C2762 outputibias.n58 gnd 0.002683f
C2763 outputibias.n59 gnd 5.55e-19
C2764 outputibias.n60 gnd 5.24e-19
C2765 outputibias.n61 gnd 0.002256f
C2766 outputibias.n62 gnd 0.005197f
C2767 outputibias.n63 gnd 0.121892f
C2768 outputibias.n64 gnd 0.001372f
C2769 outputibias.n65 gnd 9.76e-19
C2770 outputibias.n66 gnd 5.24e-19
C2771 outputibias.n67 gnd 0.001239f
C2772 outputibias.n68 gnd 5.55e-19
C2773 outputibias.n69 gnd 9.76e-19
C2774 outputibias.n70 gnd 5.24e-19
C2775 outputibias.n71 gnd 0.001239f
C2776 outputibias.n72 gnd 5.55e-19
C2777 outputibias.n73 gnd 0.004176f
C2778 outputibias.t1 gnd 0.00202f
C2779 outputibias.n74 gnd 9.3e-19
C2780 outputibias.n75 gnd 7.32e-19
C2781 outputibias.n76 gnd 5.24e-19
C2782 outputibias.n77 gnd 0.02322f
C2783 outputibias.n78 gnd 9.76e-19
C2784 outputibias.n79 gnd 5.24e-19
C2785 outputibias.n80 gnd 5.55e-19
C2786 outputibias.n81 gnd 0.001239f
C2787 outputibias.n82 gnd 0.001239f
C2788 outputibias.n83 gnd 5.55e-19
C2789 outputibias.n84 gnd 5.24e-19
C2790 outputibias.n85 gnd 9.76e-19
C2791 outputibias.n86 gnd 9.76e-19
C2792 outputibias.n87 gnd 5.24e-19
C2793 outputibias.n88 gnd 5.55e-19
C2794 outputibias.n89 gnd 0.001239f
C2795 outputibias.n90 gnd 0.002683f
C2796 outputibias.n91 gnd 5.55e-19
C2797 outputibias.n92 gnd 5.24e-19
C2798 outputibias.n93 gnd 0.002256f
C2799 outputibias.n94 gnd 0.005197f
C2800 outputibias.n95 gnd 0.064513f
C2801 outputibias.n96 gnd 0.001372f
C2802 outputibias.n97 gnd 9.76e-19
C2803 outputibias.n98 gnd 5.24e-19
C2804 outputibias.n99 gnd 0.001239f
C2805 outputibias.n100 gnd 5.55e-19
C2806 outputibias.n101 gnd 9.76e-19
C2807 outputibias.n102 gnd 5.24e-19
C2808 outputibias.n103 gnd 0.001239f
C2809 outputibias.n104 gnd 5.55e-19
C2810 outputibias.n105 gnd 0.004176f
C2811 outputibias.t7 gnd 0.00202f
C2812 outputibias.n106 gnd 9.3e-19
C2813 outputibias.n107 gnd 7.32e-19
C2814 outputibias.n108 gnd 5.24e-19
C2815 outputibias.n109 gnd 0.02322f
C2816 outputibias.n110 gnd 9.76e-19
C2817 outputibias.n111 gnd 5.24e-19
C2818 outputibias.n112 gnd 5.55e-19
C2819 outputibias.n113 gnd 0.001239f
C2820 outputibias.n114 gnd 0.001239f
C2821 outputibias.n115 gnd 5.55e-19
C2822 outputibias.n116 gnd 5.24e-19
C2823 outputibias.n117 gnd 9.76e-19
C2824 outputibias.n118 gnd 9.76e-19
C2825 outputibias.n119 gnd 5.24e-19
C2826 outputibias.n120 gnd 5.55e-19
C2827 outputibias.n121 gnd 0.001239f
C2828 outputibias.n122 gnd 0.002683f
C2829 outputibias.n123 gnd 5.55e-19
C2830 outputibias.n124 gnd 5.24e-19
C2831 outputibias.n125 gnd 0.002256f
C2832 outputibias.n126 gnd 0.005197f
C2833 outputibias.n127 gnd 0.084814f
C2834 outputibias.t6 gnd 0.108319f
C2835 outputibias.t0 gnd 0.108319f
C2836 outputibias.t2 gnd 0.108319f
C2837 outputibias.t4 gnd 0.109238f
C2838 outputibias.n128 gnd 0.134674f
C2839 outputibias.n129 gnd 0.07244f
C2840 outputibias.n130 gnd 0.079818f
C2841 outputibias.n131 gnd 0.164901f
C2842 outputibias.t11 gnd 0.11477f
C2843 outputibias.n132 gnd 0.067481f
C2844 outputibias.t9 gnd 0.11477f
C2845 outputibias.n133 gnd 0.065115f
C2846 outputibias.n134 gnd 0.029159f
C2847 a_n1808_13878.t11 gnd 0.185195f
C2848 a_n1808_13878.t13 gnd 0.185195f
C2849 a_n1808_13878.t17 gnd 0.185195f
C2850 a_n1808_13878.n0 gnd 1.46067f
C2851 a_n1808_13878.t8 gnd 0.185195f
C2852 a_n1808_13878.t10 gnd 0.185195f
C2853 a_n1808_13878.n1 gnd 1.4598f
C2854 a_n1808_13878.t14 gnd 0.185195f
C2855 a_n1808_13878.t9 gnd 0.185195f
C2856 a_n1808_13878.n2 gnd 1.45825f
C2857 a_n1808_13878.n3 gnd 2.03762f
C2858 a_n1808_13878.t12 gnd 0.185195f
C2859 a_n1808_13878.t19 gnd 0.185195f
C2860 a_n1808_13878.n4 gnd 1.45825f
C2861 a_n1808_13878.n5 gnd 3.69301f
C2862 a_n1808_13878.t1 gnd 1.73408f
C2863 a_n1808_13878.t4 gnd 0.185195f
C2864 a_n1808_13878.t5 gnd 0.185195f
C2865 a_n1808_13878.n6 gnd 1.30452f
C2866 a_n1808_13878.n7 gnd 1.4576f
C2867 a_n1808_13878.t0 gnd 1.73062f
C2868 a_n1808_13878.n8 gnd 0.733487f
C2869 a_n1808_13878.t3 gnd 1.73062f
C2870 a_n1808_13878.n9 gnd 0.733487f
C2871 a_n1808_13878.t6 gnd 0.185195f
C2872 a_n1808_13878.t7 gnd 0.185195f
C2873 a_n1808_13878.n10 gnd 1.30452f
C2874 a_n1808_13878.n11 gnd 0.74059f
C2875 a_n1808_13878.t2 gnd 1.73062f
C2876 a_n1808_13878.n12 gnd 1.7272f
C2877 a_n1808_13878.n13 gnd 2.51438f
C2878 a_n1808_13878.t15 gnd 0.185195f
C2879 a_n1808_13878.t16 gnd 0.185195f
C2880 a_n1808_13878.n14 gnd 1.45825f
C2881 a_n1808_13878.n15 gnd 1.80025f
C2882 a_n1808_13878.n16 gnd 1.31079f
C2883 a_n1808_13878.n17 gnd 1.45826f
C2884 a_n1808_13878.t18 gnd 0.185195f
C2885 a_n1986_8322.t0 gnd 0.126101p
C2886 a_n1986_8322.t18 gnd 0.09348f
C2887 a_n1986_8322.t7 gnd 0.875295f
C2888 a_n1986_8322.t11 gnd 0.09348f
C2889 a_n1986_8322.t10 gnd 0.09348f
C2890 a_n1986_8322.n0 gnd 0.658471f
C2891 a_n1986_8322.n1 gnd 0.735747f
C2892 a_n1986_8322.t3 gnd 0.09348f
C2893 a_n1986_8322.t8 gnd 0.09348f
C2894 a_n1986_8322.n2 gnd 0.658471f
C2895 a_n1986_8322.n3 gnd 0.373822f
C2896 a_n1986_8322.t4 gnd 0.873554f
C2897 a_n1986_8322.n4 gnd 0.766087f
C2898 a_n1986_8322.n5 gnd 4.03761f
C2899 a_n1986_8322.t6 gnd 0.875297f
C2900 a_n1986_8322.t12 gnd 0.09348f
C2901 a_n1986_8322.t9 gnd 0.09348f
C2902 a_n1986_8322.n6 gnd 0.658471f
C2903 a_n1986_8322.n7 gnd 0.735745f
C2904 a_n1986_8322.t2 gnd 0.09348f
C2905 a_n1986_8322.t1 gnd 0.09348f
C2906 a_n1986_8322.n8 gnd 0.658471f
C2907 a_n1986_8322.n9 gnd 0.373822f
C2908 a_n1986_8322.t5 gnd 0.873554f
C2909 a_n1986_8322.n10 gnd 1.39817f
C2910 a_n1986_8322.n11 gnd 1.58981f
C2911 a_n1986_8322.t17 gnd 0.873554f
C2912 a_n1986_8322.n12 gnd 0.871824f
C2913 a_n1986_8322.t14 gnd 0.09348f
C2914 a_n1986_8322.t20 gnd 0.09348f
C2915 a_n1986_8322.n13 gnd 0.658471f
C2916 a_n1986_8322.n14 gnd 0.373822f
C2917 a_n1986_8322.t16 gnd 0.873554f
C2918 a_n1986_8322.n15 gnd 0.370237f
C2919 a_n1986_8322.t13 gnd 0.873554f
C2920 a_n1986_8322.n16 gnd 0.370237f
C2921 a_n1986_8322.t15 gnd 0.875297f
C2922 a_n1986_8322.n17 gnd 0.735743f
C2923 a_n1986_8322.n18 gnd 0.658473f
C2924 a_n1986_8322.t19 gnd 0.09348f
C2925 vdd.t263 gnd 0.040588f
C2926 vdd.t249 gnd 0.040588f
C2927 vdd.n0 gnd 0.320123f
C2928 vdd.t275 gnd 0.040588f
C2929 vdd.t259 gnd 0.040588f
C2930 vdd.n1 gnd 0.319595f
C2931 vdd.n2 gnd 0.294727f
C2932 vdd.t246 gnd 0.040588f
C2933 vdd.t269 gnd 0.040588f
C2934 vdd.n3 gnd 0.319595f
C2935 vdd.n4 gnd 0.149055f
C2936 vdd.t267 gnd 0.040588f
C2937 vdd.t254 gnd 0.040588f
C2938 vdd.n5 gnd 0.319595f
C2939 vdd.n6 gnd 0.13986f
C2940 vdd.t273 gnd 0.040588f
C2941 vdd.t244 gnd 0.040588f
C2942 vdd.n7 gnd 0.320123f
C2943 vdd.t252 gnd 0.040588f
C2944 vdd.t265 gnd 0.040588f
C2945 vdd.n8 gnd 0.319595f
C2946 vdd.n9 gnd 0.294727f
C2947 vdd.t236 gnd 0.040588f
C2948 vdd.t234 gnd 0.040588f
C2949 vdd.n10 gnd 0.319595f
C2950 vdd.n11 gnd 0.149055f
C2951 vdd.t241 gnd 0.040588f
C2952 vdd.t257 gnd 0.040588f
C2953 vdd.n12 gnd 0.319595f
C2954 vdd.n13 gnd 0.13986f
C2955 vdd.n14 gnd 0.098879f
C2956 vdd.t2 gnd 0.022549f
C2957 vdd.t142 gnd 0.022549f
C2958 vdd.n15 gnd 0.207552f
C2959 vdd.t136 gnd 0.022549f
C2960 vdd.t137 gnd 0.022549f
C2961 vdd.n16 gnd 0.206945f
C2962 vdd.n17 gnd 0.360149f
C2963 vdd.t49 gnd 0.022549f
C2964 vdd.t143 gnd 0.022549f
C2965 vdd.n18 gnd 0.206945f
C2966 vdd.n19 gnd 0.148998f
C2967 vdd.t11 gnd 0.022549f
C2968 vdd.t138 gnd 0.022549f
C2969 vdd.n20 gnd 0.207552f
C2970 vdd.t47 gnd 0.022549f
C2971 vdd.t0 gnd 0.022549f
C2972 vdd.n21 gnd 0.206945f
C2973 vdd.n22 gnd 0.360149f
C2974 vdd.t9 gnd 0.022549f
C2975 vdd.t10 gnd 0.022549f
C2976 vdd.n23 gnd 0.206945f
C2977 vdd.n24 gnd 0.148998f
C2978 vdd.t1 gnd 0.022549f
C2979 vdd.t139 gnd 0.022549f
C2980 vdd.n25 gnd 0.206945f
C2981 vdd.t141 gnd 0.022549f
C2982 vdd.t48 gnd 0.022549f
C2983 vdd.n26 gnd 0.206945f
C2984 vdd.n27 gnd 24.3046f
C2985 vdd.n28 gnd 9.22561f
C2986 vdd.n29 gnd 0.00615f
C2987 vdd.n30 gnd 0.005707f
C2988 vdd.n31 gnd 0.003157f
C2989 vdd.n32 gnd 0.007248f
C2990 vdd.n33 gnd 0.003067f
C2991 vdd.n34 gnd 0.003247f
C2992 vdd.n35 gnd 0.005707f
C2993 vdd.n36 gnd 0.003067f
C2994 vdd.n37 gnd 0.007248f
C2995 vdd.n38 gnd 0.003247f
C2996 vdd.n39 gnd 0.005707f
C2997 vdd.n40 gnd 0.003067f
C2998 vdd.n41 gnd 0.005436f
C2999 vdd.n42 gnd 0.005453f
C3000 vdd.t35 gnd 0.015573f
C3001 vdd.n43 gnd 0.034649f
C3002 vdd.n44 gnd 0.180321f
C3003 vdd.n45 gnd 0.003067f
C3004 vdd.n46 gnd 0.003247f
C3005 vdd.n47 gnd 0.007248f
C3006 vdd.n48 gnd 0.007248f
C3007 vdd.n49 gnd 0.003247f
C3008 vdd.n50 gnd 0.003067f
C3009 vdd.n51 gnd 0.005707f
C3010 vdd.n52 gnd 0.005707f
C3011 vdd.n53 gnd 0.003067f
C3012 vdd.n54 gnd 0.003247f
C3013 vdd.n55 gnd 0.007248f
C3014 vdd.n56 gnd 0.007248f
C3015 vdd.n57 gnd 0.003247f
C3016 vdd.n58 gnd 0.003067f
C3017 vdd.n59 gnd 0.005707f
C3018 vdd.n60 gnd 0.005707f
C3019 vdd.n61 gnd 0.003067f
C3020 vdd.n62 gnd 0.003247f
C3021 vdd.n63 gnd 0.007248f
C3022 vdd.n64 gnd 0.007248f
C3023 vdd.n65 gnd 0.017137f
C3024 vdd.n66 gnd 0.003157f
C3025 vdd.n67 gnd 0.003067f
C3026 vdd.n68 gnd 0.014751f
C3027 vdd.n69 gnd 0.010298f
C3028 vdd.t284 gnd 0.036078f
C3029 vdd.t73 gnd 0.036078f
C3030 vdd.n70 gnd 0.247954f
C3031 vdd.n71 gnd 0.194978f
C3032 vdd.t81 gnd 0.036078f
C3033 vdd.t19 gnd 0.036078f
C3034 vdd.n72 gnd 0.247954f
C3035 vdd.n73 gnd 0.157346f
C3036 vdd.t223 gnd 0.036078f
C3037 vdd.t119 gnd 0.036078f
C3038 vdd.n74 gnd 0.247954f
C3039 vdd.n75 gnd 0.157346f
C3040 vdd.t293 gnd 0.036078f
C3041 vdd.t98 gnd 0.036078f
C3042 vdd.n76 gnd 0.247954f
C3043 vdd.n77 gnd 0.157346f
C3044 vdd.t15 gnd 0.036078f
C3045 vdd.t12 gnd 0.036078f
C3046 vdd.n78 gnd 0.247954f
C3047 vdd.n79 gnd 0.157346f
C3048 vdd.t65 gnd 0.036078f
C3049 vdd.t280 gnd 0.036078f
C3050 vdd.n80 gnd 0.247954f
C3051 vdd.n81 gnd 0.157346f
C3052 vdd.t25 gnd 0.036078f
C3053 vdd.t286 gnd 0.036078f
C3054 vdd.n82 gnd 0.247954f
C3055 vdd.n83 gnd 0.157346f
C3056 vdd.t105 gnd 0.036078f
C3057 vdd.t126 gnd 0.036078f
C3058 vdd.n84 gnd 0.247954f
C3059 vdd.n85 gnd 0.157346f
C3060 vdd.t31 gnd 0.036078f
C3061 vdd.t97 gnd 0.036078f
C3062 vdd.n86 gnd 0.247954f
C3063 vdd.n87 gnd 0.157346f
C3064 vdd.n88 gnd 0.00615f
C3065 vdd.n89 gnd 0.005707f
C3066 vdd.n90 gnd 0.003157f
C3067 vdd.n91 gnd 0.007248f
C3068 vdd.n92 gnd 0.003067f
C3069 vdd.n93 gnd 0.003247f
C3070 vdd.n94 gnd 0.005707f
C3071 vdd.n95 gnd 0.003067f
C3072 vdd.n96 gnd 0.007248f
C3073 vdd.n97 gnd 0.003247f
C3074 vdd.n98 gnd 0.005707f
C3075 vdd.n99 gnd 0.003067f
C3076 vdd.n100 gnd 0.005436f
C3077 vdd.n101 gnd 0.005453f
C3078 vdd.t118 gnd 0.015573f
C3079 vdd.n102 gnd 0.034649f
C3080 vdd.n103 gnd 0.180321f
C3081 vdd.n104 gnd 0.003067f
C3082 vdd.n105 gnd 0.003247f
C3083 vdd.n106 gnd 0.007248f
C3084 vdd.n107 gnd 0.007248f
C3085 vdd.n108 gnd 0.003247f
C3086 vdd.n109 gnd 0.003067f
C3087 vdd.n110 gnd 0.005707f
C3088 vdd.n111 gnd 0.005707f
C3089 vdd.n112 gnd 0.003067f
C3090 vdd.n113 gnd 0.003247f
C3091 vdd.n114 gnd 0.007248f
C3092 vdd.n115 gnd 0.007248f
C3093 vdd.n116 gnd 0.003247f
C3094 vdd.n117 gnd 0.003067f
C3095 vdd.n118 gnd 0.005707f
C3096 vdd.n119 gnd 0.005707f
C3097 vdd.n120 gnd 0.003067f
C3098 vdd.n121 gnd 0.003247f
C3099 vdd.n122 gnd 0.007248f
C3100 vdd.n123 gnd 0.007248f
C3101 vdd.n124 gnd 0.017137f
C3102 vdd.n125 gnd 0.003157f
C3103 vdd.n126 gnd 0.003067f
C3104 vdd.n127 gnd 0.014751f
C3105 vdd.n128 gnd 0.009975f
C3106 vdd.n129 gnd 0.117066f
C3107 vdd.n130 gnd 0.00615f
C3108 vdd.n131 gnd 0.005707f
C3109 vdd.n132 gnd 0.003157f
C3110 vdd.n133 gnd 0.007248f
C3111 vdd.n134 gnd 0.003067f
C3112 vdd.n135 gnd 0.003247f
C3113 vdd.n136 gnd 0.005707f
C3114 vdd.n137 gnd 0.003067f
C3115 vdd.n138 gnd 0.007248f
C3116 vdd.n139 gnd 0.003247f
C3117 vdd.n140 gnd 0.005707f
C3118 vdd.n141 gnd 0.003067f
C3119 vdd.n142 gnd 0.005436f
C3120 vdd.n143 gnd 0.005453f
C3121 vdd.t46 gnd 0.015573f
C3122 vdd.n144 gnd 0.034649f
C3123 vdd.n145 gnd 0.180321f
C3124 vdd.n146 gnd 0.003067f
C3125 vdd.n147 gnd 0.003247f
C3126 vdd.n148 gnd 0.007248f
C3127 vdd.n149 gnd 0.007248f
C3128 vdd.n150 gnd 0.003247f
C3129 vdd.n151 gnd 0.003067f
C3130 vdd.n152 gnd 0.005707f
C3131 vdd.n153 gnd 0.005707f
C3132 vdd.n154 gnd 0.003067f
C3133 vdd.n155 gnd 0.003247f
C3134 vdd.n156 gnd 0.007248f
C3135 vdd.n157 gnd 0.007248f
C3136 vdd.n158 gnd 0.003247f
C3137 vdd.n159 gnd 0.003067f
C3138 vdd.n160 gnd 0.005707f
C3139 vdd.n161 gnd 0.005707f
C3140 vdd.n162 gnd 0.003067f
C3141 vdd.n163 gnd 0.003247f
C3142 vdd.n164 gnd 0.007248f
C3143 vdd.n165 gnd 0.007248f
C3144 vdd.n166 gnd 0.017137f
C3145 vdd.n167 gnd 0.003157f
C3146 vdd.n168 gnd 0.003067f
C3147 vdd.n169 gnd 0.014751f
C3148 vdd.n170 gnd 0.010298f
C3149 vdd.t45 gnd 0.036078f
C3150 vdd.t94 gnd 0.036078f
C3151 vdd.n171 gnd 0.247954f
C3152 vdd.n172 gnd 0.194978f
C3153 vdd.t134 gnd 0.036078f
C3154 vdd.t34 gnd 0.036078f
C3155 vdd.n173 gnd 0.247954f
C3156 vdd.n174 gnd 0.157346f
C3157 vdd.t106 gnd 0.036078f
C3158 vdd.t83 gnd 0.036078f
C3159 vdd.n175 gnd 0.247954f
C3160 vdd.n176 gnd 0.157346f
C3161 vdd.t4 gnd 0.036078f
C3162 vdd.t17 gnd 0.036078f
C3163 vdd.n177 gnd 0.247954f
C3164 vdd.n178 gnd 0.157346f
C3165 vdd.t230 gnd 0.036078f
C3166 vdd.t8 gnd 0.036078f
C3167 vdd.n179 gnd 0.247954f
C3168 vdd.n180 gnd 0.157346f
C3169 vdd.t277 gnd 0.036078f
C3170 vdd.t225 gnd 0.036078f
C3171 vdd.n181 gnd 0.247954f
C3172 vdd.n182 gnd 0.157346f
C3173 vdd.t285 gnd 0.036078f
C3174 vdd.t38 gnd 0.036078f
C3175 vdd.n183 gnd 0.247954f
C3176 vdd.n184 gnd 0.157346f
C3177 vdd.t96 gnd 0.036078f
C3178 vdd.t287 gnd 0.036078f
C3179 vdd.n185 gnd 0.247954f
C3180 vdd.n186 gnd 0.157346f
C3181 vdd.t36 gnd 0.036078f
C3182 vdd.t75 gnd 0.036078f
C3183 vdd.n187 gnd 0.247954f
C3184 vdd.n188 gnd 0.157346f
C3185 vdd.n189 gnd 0.00615f
C3186 vdd.n190 gnd 0.005707f
C3187 vdd.n191 gnd 0.003157f
C3188 vdd.n192 gnd 0.007248f
C3189 vdd.n193 gnd 0.003067f
C3190 vdd.n194 gnd 0.003247f
C3191 vdd.n195 gnd 0.005707f
C3192 vdd.n196 gnd 0.003067f
C3193 vdd.n197 gnd 0.007248f
C3194 vdd.n198 gnd 0.003247f
C3195 vdd.n199 gnd 0.005707f
C3196 vdd.n200 gnd 0.003067f
C3197 vdd.n201 gnd 0.005436f
C3198 vdd.n202 gnd 0.005453f
C3199 vdd.t107 gnd 0.015573f
C3200 vdd.n203 gnd 0.034649f
C3201 vdd.n204 gnd 0.180321f
C3202 vdd.n205 gnd 0.003067f
C3203 vdd.n206 gnd 0.003247f
C3204 vdd.n207 gnd 0.007248f
C3205 vdd.n208 gnd 0.007248f
C3206 vdd.n209 gnd 0.003247f
C3207 vdd.n210 gnd 0.003067f
C3208 vdd.n211 gnd 0.005707f
C3209 vdd.n212 gnd 0.005707f
C3210 vdd.n213 gnd 0.003067f
C3211 vdd.n214 gnd 0.003247f
C3212 vdd.n215 gnd 0.007248f
C3213 vdd.n216 gnd 0.007248f
C3214 vdd.n217 gnd 0.003247f
C3215 vdd.n218 gnd 0.003067f
C3216 vdd.n219 gnd 0.005707f
C3217 vdd.n220 gnd 0.005707f
C3218 vdd.n221 gnd 0.003067f
C3219 vdd.n222 gnd 0.003247f
C3220 vdd.n223 gnd 0.007248f
C3221 vdd.n224 gnd 0.007248f
C3222 vdd.n225 gnd 0.017137f
C3223 vdd.n226 gnd 0.003157f
C3224 vdd.n227 gnd 0.003067f
C3225 vdd.n228 gnd 0.014751f
C3226 vdd.n229 gnd 0.009975f
C3227 vdd.n230 gnd 0.069642f
C3228 vdd.n231 gnd 0.25094f
C3229 vdd.n232 gnd 0.00615f
C3230 vdd.n233 gnd 0.005707f
C3231 vdd.n234 gnd 0.003157f
C3232 vdd.n235 gnd 0.007248f
C3233 vdd.n236 gnd 0.003067f
C3234 vdd.n237 gnd 0.003247f
C3235 vdd.n238 gnd 0.005707f
C3236 vdd.n239 gnd 0.003067f
C3237 vdd.n240 gnd 0.007248f
C3238 vdd.n241 gnd 0.003247f
C3239 vdd.n242 gnd 0.005707f
C3240 vdd.n243 gnd 0.003067f
C3241 vdd.n244 gnd 0.005436f
C3242 vdd.n245 gnd 0.005453f
C3243 vdd.t23 gnd 0.015573f
C3244 vdd.n246 gnd 0.034649f
C3245 vdd.n247 gnd 0.180321f
C3246 vdd.n248 gnd 0.003067f
C3247 vdd.n249 gnd 0.003247f
C3248 vdd.n250 gnd 0.007248f
C3249 vdd.n251 gnd 0.007248f
C3250 vdd.n252 gnd 0.003247f
C3251 vdd.n253 gnd 0.003067f
C3252 vdd.n254 gnd 0.005707f
C3253 vdd.n255 gnd 0.005707f
C3254 vdd.n256 gnd 0.003067f
C3255 vdd.n257 gnd 0.003247f
C3256 vdd.n258 gnd 0.007248f
C3257 vdd.n259 gnd 0.007248f
C3258 vdd.n260 gnd 0.003247f
C3259 vdd.n261 gnd 0.003067f
C3260 vdd.n262 gnd 0.005707f
C3261 vdd.n263 gnd 0.005707f
C3262 vdd.n264 gnd 0.003067f
C3263 vdd.n265 gnd 0.003247f
C3264 vdd.n266 gnd 0.007248f
C3265 vdd.n267 gnd 0.007248f
C3266 vdd.n268 gnd 0.017137f
C3267 vdd.n269 gnd 0.003157f
C3268 vdd.n270 gnd 0.003067f
C3269 vdd.n271 gnd 0.014751f
C3270 vdd.n272 gnd 0.010298f
C3271 vdd.t21 gnd 0.036078f
C3272 vdd.t229 gnd 0.036078f
C3273 vdd.n273 gnd 0.247954f
C3274 vdd.n274 gnd 0.194978f
C3275 vdd.t108 gnd 0.036078f
C3276 vdd.t122 gnd 0.036078f
C3277 vdd.n275 gnd 0.247954f
C3278 vdd.n276 gnd 0.157346f
C3279 vdd.t100 gnd 0.036078f
C3280 vdd.t117 gnd 0.036078f
C3281 vdd.n277 gnd 0.247954f
C3282 vdd.n278 gnd 0.157346f
C3283 vdd.t135 gnd 0.036078f
C3284 vdd.t91 gnd 0.036078f
C3285 vdd.n279 gnd 0.247954f
C3286 vdd.n280 gnd 0.157346f
C3287 vdd.t89 gnd 0.036078f
C3288 vdd.t13 gnd 0.036078f
C3289 vdd.n281 gnd 0.247954f
C3290 vdd.n282 gnd 0.157346f
C3291 vdd.t278 gnd 0.036078f
C3292 vdd.t294 gnd 0.036078f
C3293 vdd.n283 gnd 0.247954f
C3294 vdd.n284 gnd 0.157346f
C3295 vdd.t90 gnd 0.036078f
C3296 vdd.t140 gnd 0.036078f
C3297 vdd.n285 gnd 0.247954f
C3298 vdd.n286 gnd 0.157346f
C3299 vdd.t283 gnd 0.036078f
C3300 vdd.t292 gnd 0.036078f
C3301 vdd.n287 gnd 0.247954f
C3302 vdd.n288 gnd 0.157346f
C3303 vdd.t129 gnd 0.036078f
C3304 vdd.t131 gnd 0.036078f
C3305 vdd.n289 gnd 0.247954f
C3306 vdd.n290 gnd 0.157346f
C3307 vdd.n291 gnd 0.00615f
C3308 vdd.n292 gnd 0.005707f
C3309 vdd.n293 gnd 0.003157f
C3310 vdd.n294 gnd 0.007248f
C3311 vdd.n295 gnd 0.003067f
C3312 vdd.n296 gnd 0.003247f
C3313 vdd.n297 gnd 0.005707f
C3314 vdd.n298 gnd 0.003067f
C3315 vdd.n299 gnd 0.007248f
C3316 vdd.n300 gnd 0.003247f
C3317 vdd.n301 gnd 0.005707f
C3318 vdd.n302 gnd 0.003067f
C3319 vdd.n303 gnd 0.005436f
C3320 vdd.n304 gnd 0.005453f
C3321 vdd.t104 gnd 0.015573f
C3322 vdd.n305 gnd 0.034649f
C3323 vdd.n306 gnd 0.180321f
C3324 vdd.n307 gnd 0.003067f
C3325 vdd.n308 gnd 0.003247f
C3326 vdd.n309 gnd 0.007248f
C3327 vdd.n310 gnd 0.007248f
C3328 vdd.n311 gnd 0.003247f
C3329 vdd.n312 gnd 0.003067f
C3330 vdd.n313 gnd 0.005707f
C3331 vdd.n314 gnd 0.005707f
C3332 vdd.n315 gnd 0.003067f
C3333 vdd.n316 gnd 0.003247f
C3334 vdd.n317 gnd 0.007248f
C3335 vdd.n318 gnd 0.007248f
C3336 vdd.n319 gnd 0.003247f
C3337 vdd.n320 gnd 0.003067f
C3338 vdd.n321 gnd 0.005707f
C3339 vdd.n322 gnd 0.005707f
C3340 vdd.n323 gnd 0.003067f
C3341 vdd.n324 gnd 0.003247f
C3342 vdd.n325 gnd 0.007248f
C3343 vdd.n326 gnd 0.007248f
C3344 vdd.n327 gnd 0.017137f
C3345 vdd.n328 gnd 0.003157f
C3346 vdd.n329 gnd 0.003067f
C3347 vdd.n330 gnd 0.014751f
C3348 vdd.n331 gnd 0.009975f
C3349 vdd.n332 gnd 0.069642f
C3350 vdd.n333 gnd 0.287272f
C3351 vdd.n334 gnd 0.008613f
C3352 vdd.n335 gnd 0.011206f
C3353 vdd.n336 gnd 0.00902f
C3354 vdd.n337 gnd 0.00902f
C3355 vdd.n338 gnd 0.011206f
C3356 vdd.n339 gnd 0.011206f
C3357 vdd.n340 gnd 0.818823f
C3358 vdd.n341 gnd 0.011206f
C3359 vdd.n342 gnd 0.011206f
C3360 vdd.n343 gnd 0.011206f
C3361 vdd.n344 gnd 0.887535f
C3362 vdd.n345 gnd 0.011206f
C3363 vdd.n346 gnd 0.011206f
C3364 vdd.n347 gnd 0.011206f
C3365 vdd.n348 gnd 0.011206f
C3366 vdd.n349 gnd 0.00902f
C3367 vdd.n350 gnd 0.011206f
C3368 vdd.t224 gnd 0.572603f
C3369 vdd.n351 gnd 0.011206f
C3370 vdd.n352 gnd 0.011206f
C3371 vdd.n353 gnd 0.011206f
C3372 vdd.t37 gnd 0.572603f
C3373 vdd.n354 gnd 0.011206f
C3374 vdd.n355 gnd 0.011206f
C3375 vdd.n356 gnd 0.011206f
C3376 vdd.n357 gnd 0.011206f
C3377 vdd.n358 gnd 0.011206f
C3378 vdd.n359 gnd 0.00902f
C3379 vdd.n360 gnd 0.011206f
C3380 vdd.n361 gnd 0.647042f
C3381 vdd.n362 gnd 0.011206f
C3382 vdd.n363 gnd 0.011206f
C3383 vdd.n364 gnd 0.011206f
C3384 vdd.t125 gnd 0.572603f
C3385 vdd.n365 gnd 0.011206f
C3386 vdd.n366 gnd 0.011206f
C3387 vdd.n367 gnd 0.011206f
C3388 vdd.n368 gnd 0.011206f
C3389 vdd.n369 gnd 0.011206f
C3390 vdd.n370 gnd 0.00902f
C3391 vdd.n371 gnd 0.011206f
C3392 vdd.t30 gnd 0.572603f
C3393 vdd.n372 gnd 0.011206f
C3394 vdd.n373 gnd 0.011206f
C3395 vdd.n374 gnd 0.011206f
C3396 vdd.n375 gnd 0.669946f
C3397 vdd.n376 gnd 0.011206f
C3398 vdd.n377 gnd 0.011206f
C3399 vdd.n378 gnd 0.011206f
C3400 vdd.n379 gnd 0.011206f
C3401 vdd.n380 gnd 0.011206f
C3402 vdd.n381 gnd 0.00902f
C3403 vdd.n382 gnd 0.011206f
C3404 vdd.t103 gnd 0.572603f
C3405 vdd.n383 gnd 0.011206f
C3406 vdd.n384 gnd 0.011206f
C3407 vdd.n385 gnd 0.011206f
C3408 vdd.n386 gnd 0.578329f
C3409 vdd.n387 gnd 0.011206f
C3410 vdd.n388 gnd 0.011206f
C3411 vdd.n389 gnd 0.011206f
C3412 vdd.n390 gnd 0.011206f
C3413 vdd.n391 gnd 0.027108f
C3414 vdd.n392 gnd 0.027689f
C3415 vdd.t167 gnd 0.572603f
C3416 vdd.n393 gnd 0.027108f
C3417 vdd.n425 gnd 0.011206f
C3418 vdd.t169 gnd 0.137864f
C3419 vdd.t168 gnd 0.147339f
C3420 vdd.t166 gnd 0.180049f
C3421 vdd.n426 gnd 0.230797f
C3422 vdd.n427 gnd 0.194813f
C3423 vdd.n428 gnd 0.014792f
C3424 vdd.n429 gnd 0.011206f
C3425 vdd.n430 gnd 0.00902f
C3426 vdd.n431 gnd 0.011206f
C3427 vdd.n432 gnd 0.00902f
C3428 vdd.n433 gnd 0.011206f
C3429 vdd.n434 gnd 0.00902f
C3430 vdd.n435 gnd 0.011206f
C3431 vdd.n436 gnd 0.00902f
C3432 vdd.n437 gnd 0.011206f
C3433 vdd.n438 gnd 0.00902f
C3434 vdd.n439 gnd 0.011206f
C3435 vdd.t210 gnd 0.137864f
C3436 vdd.t209 gnd 0.147339f
C3437 vdd.t208 gnd 0.180049f
C3438 vdd.n440 gnd 0.230797f
C3439 vdd.n441 gnd 0.194813f
C3440 vdd.n442 gnd 0.00902f
C3441 vdd.n443 gnd 0.011206f
C3442 vdd.n444 gnd 0.00902f
C3443 vdd.n445 gnd 0.011206f
C3444 vdd.n446 gnd 0.00902f
C3445 vdd.n447 gnd 0.011206f
C3446 vdd.n448 gnd 0.00902f
C3447 vdd.n449 gnd 0.011206f
C3448 vdd.n450 gnd 0.00902f
C3449 vdd.n451 gnd 0.011206f
C3450 vdd.t216 gnd 0.137864f
C3451 vdd.t215 gnd 0.147339f
C3452 vdd.t214 gnd 0.180049f
C3453 vdd.n452 gnd 0.230797f
C3454 vdd.n453 gnd 0.194813f
C3455 vdd.n454 gnd 0.019302f
C3456 vdd.n455 gnd 0.011206f
C3457 vdd.n456 gnd 0.00902f
C3458 vdd.n457 gnd 0.011206f
C3459 vdd.n458 gnd 0.00902f
C3460 vdd.n459 gnd 0.011206f
C3461 vdd.n460 gnd 0.00902f
C3462 vdd.n461 gnd 0.011206f
C3463 vdd.n462 gnd 0.00902f
C3464 vdd.n463 gnd 0.011206f
C3465 vdd.n464 gnd 0.027689f
C3466 vdd.n465 gnd 0.007486f
C3467 vdd.n466 gnd 0.00902f
C3468 vdd.n467 gnd 0.011206f
C3469 vdd.n468 gnd 0.011206f
C3470 vdd.n469 gnd 0.00902f
C3471 vdd.n470 gnd 0.011206f
C3472 vdd.n471 gnd 0.011206f
C3473 vdd.n472 gnd 0.011206f
C3474 vdd.n473 gnd 0.011206f
C3475 vdd.n474 gnd 0.011206f
C3476 vdd.n475 gnd 0.00902f
C3477 vdd.n476 gnd 0.00902f
C3478 vdd.n477 gnd 0.011206f
C3479 vdd.n478 gnd 0.011206f
C3480 vdd.n479 gnd 0.00902f
C3481 vdd.n480 gnd 0.011206f
C3482 vdd.n481 gnd 0.011206f
C3483 vdd.n482 gnd 0.011206f
C3484 vdd.n483 gnd 0.011206f
C3485 vdd.n484 gnd 0.011206f
C3486 vdd.n485 gnd 0.00902f
C3487 vdd.n486 gnd 0.00902f
C3488 vdd.n487 gnd 0.011206f
C3489 vdd.n488 gnd 0.011206f
C3490 vdd.n489 gnd 0.00902f
C3491 vdd.n490 gnd 0.011206f
C3492 vdd.n491 gnd 0.011206f
C3493 vdd.n492 gnd 0.011206f
C3494 vdd.n493 gnd 0.011206f
C3495 vdd.n494 gnd 0.011206f
C3496 vdd.n495 gnd 0.00902f
C3497 vdd.n496 gnd 0.00902f
C3498 vdd.n497 gnd 0.011206f
C3499 vdd.n498 gnd 0.011206f
C3500 vdd.n499 gnd 0.00902f
C3501 vdd.n500 gnd 0.011206f
C3502 vdd.n501 gnd 0.011206f
C3503 vdd.n502 gnd 0.011206f
C3504 vdd.n503 gnd 0.011206f
C3505 vdd.n504 gnd 0.011206f
C3506 vdd.n505 gnd 0.00902f
C3507 vdd.n506 gnd 0.00902f
C3508 vdd.n507 gnd 0.011206f
C3509 vdd.n508 gnd 0.011206f
C3510 vdd.n509 gnd 0.007531f
C3511 vdd.n510 gnd 0.011206f
C3512 vdd.n511 gnd 0.011206f
C3513 vdd.n512 gnd 0.011206f
C3514 vdd.n513 gnd 0.011206f
C3515 vdd.n514 gnd 0.011206f
C3516 vdd.n515 gnd 0.007531f
C3517 vdd.n516 gnd 0.00902f
C3518 vdd.n517 gnd 0.011206f
C3519 vdd.n518 gnd 0.011206f
C3520 vdd.n519 gnd 0.00902f
C3521 vdd.n520 gnd 0.011206f
C3522 vdd.n521 gnd 0.011206f
C3523 vdd.n522 gnd 0.011206f
C3524 vdd.n523 gnd 0.011206f
C3525 vdd.n524 gnd 0.011206f
C3526 vdd.n525 gnd 0.00902f
C3527 vdd.n526 gnd 0.00902f
C3528 vdd.n527 gnd 0.011206f
C3529 vdd.n528 gnd 0.011206f
C3530 vdd.n529 gnd 0.00902f
C3531 vdd.n530 gnd 0.011206f
C3532 vdd.n531 gnd 0.011206f
C3533 vdd.n532 gnd 0.011206f
C3534 vdd.n533 gnd 0.011206f
C3535 vdd.n534 gnd 0.011206f
C3536 vdd.n535 gnd 0.00902f
C3537 vdd.n536 gnd 0.00902f
C3538 vdd.n537 gnd 0.011206f
C3539 vdd.n538 gnd 0.011206f
C3540 vdd.n539 gnd 0.00902f
C3541 vdd.n540 gnd 0.011206f
C3542 vdd.n541 gnd 0.011206f
C3543 vdd.n542 gnd 0.011206f
C3544 vdd.n543 gnd 0.011206f
C3545 vdd.n544 gnd 0.011206f
C3546 vdd.n545 gnd 0.00902f
C3547 vdd.n546 gnd 0.00902f
C3548 vdd.n547 gnd 0.011206f
C3549 vdd.n548 gnd 0.011206f
C3550 vdd.n549 gnd 0.00902f
C3551 vdd.n550 gnd 0.011206f
C3552 vdd.n551 gnd 0.011206f
C3553 vdd.n552 gnd 0.011206f
C3554 vdd.n553 gnd 0.011206f
C3555 vdd.n554 gnd 0.011206f
C3556 vdd.n555 gnd 0.00902f
C3557 vdd.n556 gnd 0.00902f
C3558 vdd.n557 gnd 0.011206f
C3559 vdd.n558 gnd 0.011206f
C3560 vdd.n559 gnd 0.00902f
C3561 vdd.n560 gnd 0.011206f
C3562 vdd.n561 gnd 0.011206f
C3563 vdd.n562 gnd 0.011206f
C3564 vdd.n563 gnd 0.011206f
C3565 vdd.n564 gnd 0.011206f
C3566 vdd.n565 gnd 0.006133f
C3567 vdd.n566 gnd 0.019302f
C3568 vdd.n567 gnd 0.011206f
C3569 vdd.n568 gnd 0.011206f
C3570 vdd.n569 gnd 0.008929f
C3571 vdd.n570 gnd 0.011206f
C3572 vdd.n571 gnd 0.011206f
C3573 vdd.n572 gnd 0.011206f
C3574 vdd.n573 gnd 0.011206f
C3575 vdd.n574 gnd 0.011206f
C3576 vdd.n575 gnd 0.00902f
C3577 vdd.n576 gnd 0.00902f
C3578 vdd.n577 gnd 0.011206f
C3579 vdd.n578 gnd 0.011206f
C3580 vdd.n579 gnd 0.00902f
C3581 vdd.n580 gnd 0.011206f
C3582 vdd.n581 gnd 0.011206f
C3583 vdd.n582 gnd 0.011206f
C3584 vdd.n583 gnd 0.011206f
C3585 vdd.n584 gnd 0.011206f
C3586 vdd.n585 gnd 0.00902f
C3587 vdd.n586 gnd 0.00902f
C3588 vdd.n587 gnd 0.011206f
C3589 vdd.n588 gnd 0.011206f
C3590 vdd.n589 gnd 0.00902f
C3591 vdd.n590 gnd 0.011206f
C3592 vdd.n591 gnd 0.011206f
C3593 vdd.n592 gnd 0.011206f
C3594 vdd.n593 gnd 0.011206f
C3595 vdd.n594 gnd 0.011206f
C3596 vdd.n595 gnd 0.00902f
C3597 vdd.n596 gnd 0.00902f
C3598 vdd.n597 gnd 0.011206f
C3599 vdd.n598 gnd 0.011206f
C3600 vdd.n599 gnd 0.00902f
C3601 vdd.n600 gnd 0.011206f
C3602 vdd.n601 gnd 0.011206f
C3603 vdd.n602 gnd 0.011206f
C3604 vdd.n603 gnd 0.011206f
C3605 vdd.n604 gnd 0.011206f
C3606 vdd.n605 gnd 0.00902f
C3607 vdd.n606 gnd 0.00902f
C3608 vdd.n607 gnd 0.011206f
C3609 vdd.n608 gnd 0.011206f
C3610 vdd.n609 gnd 0.00902f
C3611 vdd.n610 gnd 0.011206f
C3612 vdd.n611 gnd 0.011206f
C3613 vdd.n612 gnd 0.011206f
C3614 vdd.n613 gnd 0.011206f
C3615 vdd.n614 gnd 0.011206f
C3616 vdd.n615 gnd 0.00902f
C3617 vdd.n616 gnd 0.011206f
C3618 vdd.n617 gnd 0.00902f
C3619 vdd.n618 gnd 0.004735f
C3620 vdd.n619 gnd 0.011206f
C3621 vdd.n620 gnd 0.011206f
C3622 vdd.n621 gnd 0.00902f
C3623 vdd.n622 gnd 0.011206f
C3624 vdd.n623 gnd 0.00902f
C3625 vdd.n624 gnd 0.011206f
C3626 vdd.n625 gnd 0.00902f
C3627 vdd.n626 gnd 0.011206f
C3628 vdd.n627 gnd 0.00902f
C3629 vdd.n628 gnd 0.011206f
C3630 vdd.n629 gnd 0.00902f
C3631 vdd.n630 gnd 0.011206f
C3632 vdd.n631 gnd 0.00902f
C3633 vdd.n632 gnd 0.011206f
C3634 vdd.n633 gnd 0.624138f
C3635 vdd.t14 gnd 0.572603f
C3636 vdd.n634 gnd 0.011206f
C3637 vdd.n635 gnd 0.00902f
C3638 vdd.n636 gnd 0.011206f
C3639 vdd.n637 gnd 0.00902f
C3640 vdd.n638 gnd 0.011206f
C3641 vdd.t3 gnd 0.572603f
C3642 vdd.n639 gnd 0.011206f
C3643 vdd.n640 gnd 0.00902f
C3644 vdd.n641 gnd 0.011206f
C3645 vdd.n642 gnd 0.00902f
C3646 vdd.n643 gnd 0.011206f
C3647 vdd.t82 gnd 0.572603f
C3648 vdd.n644 gnd 0.715754f
C3649 vdd.n645 gnd 0.011206f
C3650 vdd.n646 gnd 0.00902f
C3651 vdd.n647 gnd 0.011206f
C3652 vdd.n648 gnd 0.00902f
C3653 vdd.n649 gnd 0.011206f
C3654 vdd.t99 gnd 0.572603f
C3655 vdd.n650 gnd 0.011206f
C3656 vdd.n651 gnd 0.00902f
C3657 vdd.n652 gnd 0.011206f
C3658 vdd.n653 gnd 0.00902f
C3659 vdd.n654 gnd 0.011206f
C3660 vdd.n655 gnd 0.795919f
C3661 vdd.n656 gnd 0.950521f
C3662 vdd.t18 gnd 0.572603f
C3663 vdd.n657 gnd 0.011206f
C3664 vdd.n658 gnd 0.00902f
C3665 vdd.n659 gnd 0.011206f
C3666 vdd.n660 gnd 0.00902f
C3667 vdd.n661 gnd 0.011206f
C3668 vdd.n662 gnd 0.601233f
C3669 vdd.n663 gnd 0.011206f
C3670 vdd.n664 gnd 0.00902f
C3671 vdd.n665 gnd 0.011206f
C3672 vdd.n666 gnd 0.00902f
C3673 vdd.n667 gnd 0.011206f
C3674 vdd.t20 gnd 0.572603f
C3675 vdd.t72 gnd 0.572603f
C3676 vdd.n668 gnd 0.011206f
C3677 vdd.n669 gnd 0.00902f
C3678 vdd.n670 gnd 0.011206f
C3679 vdd.n671 gnd 0.00902f
C3680 vdd.n672 gnd 0.011206f
C3681 vdd.t22 gnd 0.572603f
C3682 vdd.n673 gnd 0.011206f
C3683 vdd.n674 gnd 0.00902f
C3684 vdd.n675 gnd 0.011206f
C3685 vdd.n676 gnd 0.00902f
C3686 vdd.n677 gnd 0.011206f
C3687 vdd.n678 gnd 1.14521f
C3688 vdd.n679 gnd 0.933343f
C3689 vdd.n680 gnd 0.011206f
C3690 vdd.n681 gnd 0.00902f
C3691 vdd.n682 gnd 0.027108f
C3692 vdd.n683 gnd 0.007486f
C3693 vdd.n684 gnd 0.027108f
C3694 vdd.t145 gnd 0.572603f
C3695 vdd.n685 gnd 0.027108f
C3696 vdd.n686 gnd 0.007486f
C3697 vdd.n687 gnd 0.009637f
C3698 vdd.t212 gnd 0.137864f
C3699 vdd.t213 gnd 0.147339f
C3700 vdd.t211 gnd 0.180049f
C3701 vdd.n688 gnd 0.230797f
C3702 vdd.n689 gnd 0.193911f
C3703 vdd.n690 gnd 0.01389f
C3704 vdd.n691 gnd 0.011206f
C3705 vdd.n692 gnd 7.89047f
C3706 vdd.n723 gnd 1.57466f
C3707 vdd.n724 gnd 0.011206f
C3708 vdd.n725 gnd 0.011206f
C3709 vdd.n726 gnd 0.027689f
C3710 vdd.n727 gnd 0.009637f
C3711 vdd.n728 gnd 0.011206f
C3712 vdd.n729 gnd 0.00902f
C3713 vdd.n730 gnd 0.007172f
C3714 vdd.n731 gnd 0.018311f
C3715 vdd.n732 gnd 0.00902f
C3716 vdd.n733 gnd 0.011206f
C3717 vdd.n734 gnd 0.011206f
C3718 vdd.n735 gnd 0.011206f
C3719 vdd.n736 gnd 0.011206f
C3720 vdd.n737 gnd 0.011206f
C3721 vdd.n738 gnd 0.011206f
C3722 vdd.n739 gnd 0.011206f
C3723 vdd.n740 gnd 0.011206f
C3724 vdd.n741 gnd 0.011206f
C3725 vdd.n742 gnd 0.011206f
C3726 vdd.n743 gnd 0.011206f
C3727 vdd.n744 gnd 0.011206f
C3728 vdd.n745 gnd 0.011206f
C3729 vdd.n746 gnd 0.011206f
C3730 vdd.n747 gnd 0.007531f
C3731 vdd.n748 gnd 0.011206f
C3732 vdd.n749 gnd 0.011206f
C3733 vdd.n750 gnd 0.011206f
C3734 vdd.n751 gnd 0.011206f
C3735 vdd.n752 gnd 0.011206f
C3736 vdd.n753 gnd 0.011206f
C3737 vdd.n754 gnd 0.011206f
C3738 vdd.n755 gnd 0.011206f
C3739 vdd.n756 gnd 0.011206f
C3740 vdd.n757 gnd 0.011206f
C3741 vdd.n758 gnd 0.011206f
C3742 vdd.n759 gnd 0.011206f
C3743 vdd.n760 gnd 0.011206f
C3744 vdd.n761 gnd 0.011206f
C3745 vdd.n762 gnd 0.011206f
C3746 vdd.n763 gnd 0.011206f
C3747 vdd.n764 gnd 0.011206f
C3748 vdd.n765 gnd 0.011206f
C3749 vdd.n766 gnd 0.011206f
C3750 vdd.n767 gnd 0.008929f
C3751 vdd.t146 gnd 0.137864f
C3752 vdd.t147 gnd 0.147339f
C3753 vdd.t144 gnd 0.180049f
C3754 vdd.n768 gnd 0.230797f
C3755 vdd.n769 gnd 0.193911f
C3756 vdd.n770 gnd 0.011206f
C3757 vdd.n771 gnd 0.011206f
C3758 vdd.n772 gnd 0.011206f
C3759 vdd.n773 gnd 0.011206f
C3760 vdd.n774 gnd 0.011206f
C3761 vdd.n775 gnd 0.011206f
C3762 vdd.n776 gnd 0.011206f
C3763 vdd.n777 gnd 0.011206f
C3764 vdd.n778 gnd 0.011206f
C3765 vdd.n779 gnd 0.011206f
C3766 vdd.n780 gnd 0.011206f
C3767 vdd.n781 gnd 0.011206f
C3768 vdd.n782 gnd 0.011206f
C3769 vdd.n783 gnd 0.007172f
C3770 vdd.n785 gnd 0.00762f
C3771 vdd.n786 gnd 0.00762f
C3772 vdd.n787 gnd 0.00762f
C3773 vdd.n788 gnd 0.00762f
C3774 vdd.n789 gnd 0.00762f
C3775 vdd.n790 gnd 0.00762f
C3776 vdd.n792 gnd 0.00762f
C3777 vdd.n793 gnd 0.00762f
C3778 vdd.n795 gnd 0.00762f
C3779 vdd.n796 gnd 0.005547f
C3780 vdd.n798 gnd 0.00762f
C3781 vdd.t193 gnd 0.307928f
C3782 vdd.t192 gnd 0.315203f
C3783 vdd.t191 gnd 0.201027f
C3784 vdd.n799 gnd 0.108644f
C3785 vdd.n800 gnd 0.061626f
C3786 vdd.n801 gnd 0.01089f
C3787 vdd.n802 gnd 0.01781f
C3788 vdd.n804 gnd 0.00762f
C3789 vdd.n805 gnd 0.77874f
C3790 vdd.n806 gnd 0.016882f
C3791 vdd.n807 gnd 0.016882f
C3792 vdd.n808 gnd 0.00762f
C3793 vdd.n809 gnd 0.018081f
C3794 vdd.n810 gnd 0.00762f
C3795 vdd.n811 gnd 0.00762f
C3796 vdd.n812 gnd 0.00762f
C3797 vdd.n813 gnd 0.00762f
C3798 vdd.n814 gnd 0.00762f
C3799 vdd.n816 gnd 0.00762f
C3800 vdd.n817 gnd 0.00762f
C3801 vdd.n819 gnd 0.00762f
C3802 vdd.n820 gnd 0.00762f
C3803 vdd.n822 gnd 0.00762f
C3804 vdd.n823 gnd 0.00762f
C3805 vdd.n825 gnd 0.00762f
C3806 vdd.n826 gnd 0.00762f
C3807 vdd.n828 gnd 0.00762f
C3808 vdd.n829 gnd 0.00762f
C3809 vdd.n831 gnd 0.00762f
C3810 vdd.t186 gnd 0.307928f
C3811 vdd.t185 gnd 0.315203f
C3812 vdd.t183 gnd 0.201027f
C3813 vdd.n832 gnd 0.108644f
C3814 vdd.n833 gnd 0.061626f
C3815 vdd.n834 gnd 0.00762f
C3816 vdd.n836 gnd 0.00762f
C3817 vdd.n837 gnd 0.00762f
C3818 vdd.t184 gnd 0.38937f
C3819 vdd.n838 gnd 0.00762f
C3820 vdd.n839 gnd 0.00762f
C3821 vdd.n840 gnd 0.00762f
C3822 vdd.n841 gnd 0.00762f
C3823 vdd.n842 gnd 0.00762f
C3824 vdd.n843 gnd 0.77874f
C3825 vdd.n844 gnd 0.00762f
C3826 vdd.n845 gnd 0.00762f
C3827 vdd.n846 gnd 0.681398f
C3828 vdd.n847 gnd 0.00762f
C3829 vdd.n848 gnd 0.00762f
C3830 vdd.n849 gnd 0.006724f
C3831 vdd.n850 gnd 0.00762f
C3832 vdd.n851 gnd 0.687124f
C3833 vdd.n852 gnd 0.00762f
C3834 vdd.n853 gnd 0.00762f
C3835 vdd.n854 gnd 0.00762f
C3836 vdd.n855 gnd 0.00762f
C3837 vdd.n856 gnd 0.00762f
C3838 vdd.n857 gnd 0.77874f
C3839 vdd.n858 gnd 0.00762f
C3840 vdd.n859 gnd 0.00762f
C3841 vdd.t156 gnd 0.349288f
C3842 vdd.t237 gnd 0.091616f
C3843 vdd.n860 gnd 0.00762f
C3844 vdd.n861 gnd 0.00762f
C3845 vdd.n862 gnd 0.00762f
C3846 vdd.t247 gnd 0.38937f
C3847 vdd.n863 gnd 0.00762f
C3848 vdd.n864 gnd 0.00762f
C3849 vdd.n865 gnd 0.00762f
C3850 vdd.n866 gnd 0.00762f
C3851 vdd.n867 gnd 0.00762f
C3852 vdd.t260 gnd 0.38937f
C3853 vdd.n868 gnd 0.00762f
C3854 vdd.n869 gnd 0.00762f
C3855 vdd.n870 gnd 0.647042f
C3856 vdd.n871 gnd 0.00762f
C3857 vdd.n872 gnd 0.00762f
C3858 vdd.n873 gnd 0.00762f
C3859 vdd.n874 gnd 0.475261f
C3860 vdd.n875 gnd 0.00762f
C3861 vdd.n876 gnd 0.00762f
C3862 vdd.t243 gnd 0.38937f
C3863 vdd.n877 gnd 0.00762f
C3864 vdd.n878 gnd 0.00762f
C3865 vdd.n879 gnd 0.00762f
C3866 vdd.n880 gnd 0.647042f
C3867 vdd.n881 gnd 0.00762f
C3868 vdd.n882 gnd 0.00762f
C3869 vdd.t255 gnd 0.33211f
C3870 vdd.t272 gnd 0.30348f
C3871 vdd.n883 gnd 0.00762f
C3872 vdd.n884 gnd 0.00762f
C3873 vdd.n885 gnd 0.00762f
C3874 vdd.t264 gnd 0.38937f
C3875 vdd.n886 gnd 0.00762f
C3876 vdd.n887 gnd 0.00762f
C3877 vdd.t261 gnd 0.38937f
C3878 vdd.n888 gnd 0.00762f
C3879 vdd.n889 gnd 0.00762f
C3880 vdd.n890 gnd 0.00762f
C3881 vdd.t232 gnd 0.286302f
C3882 vdd.n891 gnd 0.00762f
C3883 vdd.n892 gnd 0.00762f
C3884 vdd.n893 gnd 0.66422f
C3885 vdd.n894 gnd 0.00762f
C3886 vdd.n895 gnd 0.00762f
C3887 vdd.n896 gnd 0.00762f
C3888 vdd.n897 gnd 0.77874f
C3889 vdd.n898 gnd 0.00762f
C3890 vdd.n899 gnd 0.00762f
C3891 vdd.t251 gnd 0.349288f
C3892 vdd.n900 gnd 0.492439f
C3893 vdd.n901 gnd 0.00762f
C3894 vdd.n902 gnd 0.00762f
C3895 vdd.n903 gnd 0.00762f
C3896 vdd.t233 gnd 0.38937f
C3897 vdd.n904 gnd 0.00762f
C3898 vdd.n905 gnd 0.00762f
C3899 vdd.n906 gnd 0.00762f
C3900 vdd.n907 gnd 0.00762f
C3901 vdd.n908 gnd 0.00762f
C3902 vdd.t235 gnd 0.77874f
C3903 vdd.n909 gnd 0.00762f
C3904 vdd.n910 gnd 0.00762f
C3905 vdd.t188 gnd 0.38937f
C3906 vdd.n911 gnd 0.00762f
C3907 vdd.n912 gnd 0.018081f
C3908 vdd.n913 gnd 0.018081f
C3909 vdd.t256 gnd 0.732932f
C3910 vdd.n914 gnd 0.016882f
C3911 vdd.n915 gnd 0.016882f
C3912 vdd.n916 gnd 0.018081f
C3913 vdd.n917 gnd 0.00762f
C3914 vdd.n918 gnd 0.00762f
C3915 vdd.t266 gnd 0.732932f
C3916 vdd.n936 gnd 0.018081f
C3917 vdd.n954 gnd 0.016882f
C3918 vdd.n955 gnd 0.00762f
C3919 vdd.n956 gnd 0.016882f
C3920 vdd.t207 gnd 0.307928f
C3921 vdd.t206 gnd 0.315203f
C3922 vdd.t205 gnd 0.201027f
C3923 vdd.n957 gnd 0.108644f
C3924 vdd.n958 gnd 0.061626f
C3925 vdd.n959 gnd 0.01781f
C3926 vdd.n960 gnd 0.00762f
C3927 vdd.t268 gnd 0.77874f
C3928 vdd.n961 gnd 0.016882f
C3929 vdd.n962 gnd 0.00762f
C3930 vdd.n963 gnd 0.018081f
C3931 vdd.n964 gnd 0.00762f
C3932 vdd.t182 gnd 0.307928f
C3933 vdd.t181 gnd 0.315203f
C3934 vdd.t179 gnd 0.201027f
C3935 vdd.n965 gnd 0.108644f
C3936 vdd.n966 gnd 0.061626f
C3937 vdd.n967 gnd 0.01089f
C3938 vdd.n968 gnd 0.00762f
C3939 vdd.n969 gnd 0.00762f
C3940 vdd.t180 gnd 0.38937f
C3941 vdd.n970 gnd 0.00762f
C3942 vdd.n971 gnd 0.00762f
C3943 vdd.n972 gnd 0.00762f
C3944 vdd.n973 gnd 0.00762f
C3945 vdd.n974 gnd 0.00762f
C3946 vdd.n975 gnd 0.00762f
C3947 vdd.n976 gnd 0.77874f
C3948 vdd.n977 gnd 0.00762f
C3949 vdd.n978 gnd 0.00762f
C3950 vdd.t245 gnd 0.38937f
C3951 vdd.n979 gnd 0.00762f
C3952 vdd.n980 gnd 0.00762f
C3953 vdd.n981 gnd 0.00762f
C3954 vdd.n982 gnd 0.00762f
C3955 vdd.n983 gnd 0.492439f
C3956 vdd.n984 gnd 0.00762f
C3957 vdd.n985 gnd 0.00762f
C3958 vdd.n986 gnd 0.00762f
C3959 vdd.n987 gnd 0.00762f
C3960 vdd.n988 gnd 0.00762f
C3961 vdd.n989 gnd 0.66422f
C3962 vdd.n990 gnd 0.00762f
C3963 vdd.n991 gnd 0.00762f
C3964 vdd.t258 gnd 0.349288f
C3965 vdd.t271 gnd 0.286302f
C3966 vdd.n992 gnd 0.00762f
C3967 vdd.n993 gnd 0.00762f
C3968 vdd.n994 gnd 0.00762f
C3969 vdd.t250 gnd 0.38937f
C3970 vdd.n995 gnd 0.00762f
C3971 vdd.n996 gnd 0.00762f
C3972 vdd.t274 gnd 0.38937f
C3973 vdd.n997 gnd 0.00762f
C3974 vdd.n998 gnd 0.00762f
C3975 vdd.n999 gnd 0.00762f
C3976 vdd.t248 gnd 0.30348f
C3977 vdd.n1000 gnd 0.00762f
C3978 vdd.n1001 gnd 0.00762f
C3979 vdd.n1002 gnd 0.647042f
C3980 vdd.n1003 gnd 0.00762f
C3981 vdd.n1004 gnd 0.00762f
C3982 vdd.n1005 gnd 0.00762f
C3983 vdd.t262 gnd 0.38937f
C3984 vdd.n1006 gnd 0.00762f
C3985 vdd.n1007 gnd 0.00762f
C3986 vdd.t239 gnd 0.33211f
C3987 vdd.n1008 gnd 0.475261f
C3988 vdd.n1009 gnd 0.00762f
C3989 vdd.n1010 gnd 0.00762f
C3990 vdd.n1011 gnd 0.00762f
C3991 vdd.n1012 gnd 0.647042f
C3992 vdd.n1013 gnd 0.00762f
C3993 vdd.n1014 gnd 0.00762f
C3994 vdd.t270 gnd 0.38937f
C3995 vdd.n1015 gnd 0.00762f
C3996 vdd.n1016 gnd 0.00762f
C3997 vdd.n1017 gnd 0.00762f
C3998 vdd.n1018 gnd 0.77874f
C3999 vdd.n1019 gnd 0.00762f
C4000 vdd.n1020 gnd 0.00762f
C4001 vdd.t242 gnd 0.38937f
C4002 vdd.n1021 gnd 0.00762f
C4003 vdd.n1022 gnd 0.00762f
C4004 vdd.n1023 gnd 0.00762f
C4005 vdd.t238 gnd 0.091616f
C4006 vdd.n1024 gnd 0.00762f
C4007 vdd.n1025 gnd 0.00762f
C4008 vdd.n1026 gnd 0.00762f
C4009 vdd.t200 gnd 0.315203f
C4010 vdd.t198 gnd 0.201027f
C4011 vdd.t201 gnd 0.315203f
C4012 vdd.n1027 gnd 0.177157f
C4013 vdd.n1028 gnd 0.00762f
C4014 vdd.n1029 gnd 0.00762f
C4015 vdd.n1030 gnd 0.77874f
C4016 vdd.n1031 gnd 0.00762f
C4017 vdd.n1032 gnd 0.00762f
C4018 vdd.t199 gnd 0.349288f
C4019 vdd.n1033 gnd 0.687124f
C4020 vdd.n1034 gnd 0.00762f
C4021 vdd.n1035 gnd 0.00762f
C4022 vdd.n1036 gnd 0.00762f
C4023 vdd.n1037 gnd 0.681398f
C4024 vdd.n1038 gnd 0.00762f
C4025 vdd.n1039 gnd 0.00762f
C4026 vdd.n1040 gnd 0.00762f
C4027 vdd.n1041 gnd 0.00762f
C4028 vdd.n1042 gnd 0.00762f
C4029 vdd.n1043 gnd 0.77874f
C4030 vdd.n1044 gnd 0.00762f
C4031 vdd.n1045 gnd 0.00762f
C4032 vdd.t195 gnd 0.38937f
C4033 vdd.n1046 gnd 0.00762f
C4034 vdd.n1047 gnd 0.018081f
C4035 vdd.n1048 gnd 0.018081f
C4036 vdd.n1049 gnd 7.89047f
C4037 vdd.n1050 gnd 0.016882f
C4038 vdd.n1051 gnd 0.016882f
C4039 vdd.n1052 gnd 0.018081f
C4040 vdd.n1053 gnd 0.00762f
C4041 vdd.n1054 gnd 0.00762f
C4042 vdd.n1055 gnd 0.00762f
C4043 vdd.n1056 gnd 0.00762f
C4044 vdd.n1057 gnd 0.00762f
C4045 vdd.n1058 gnd 0.00762f
C4046 vdd.n1059 gnd 0.00762f
C4047 vdd.n1060 gnd 0.00762f
C4048 vdd.n1062 gnd 0.00762f
C4049 vdd.n1063 gnd 0.00762f
C4050 vdd.n1064 gnd 0.007172f
C4051 vdd.n1067 gnd 0.027689f
C4052 vdd.n1068 gnd 0.00902f
C4053 vdd.n1069 gnd 0.011206f
C4054 vdd.n1071 gnd 0.011206f
C4055 vdd.n1072 gnd 0.007486f
C4056 vdd.t152 gnd 0.572603f
C4057 vdd.n1073 gnd 8.27984f
C4058 vdd.n1074 gnd 0.011206f
C4059 vdd.n1075 gnd 0.027689f
C4060 vdd.n1076 gnd 0.00902f
C4061 vdd.n1077 gnd 0.011206f
C4062 vdd.n1078 gnd 0.00902f
C4063 vdd.n1079 gnd 0.011206f
C4064 vdd.n1080 gnd 1.14521f
C4065 vdd.n1081 gnd 0.011206f
C4066 vdd.n1082 gnd 0.00902f
C4067 vdd.n1083 gnd 0.00902f
C4068 vdd.n1084 gnd 0.011206f
C4069 vdd.n1085 gnd 0.00902f
C4070 vdd.n1086 gnd 0.011206f
C4071 vdd.t61 gnd 0.572603f
C4072 vdd.n1087 gnd 0.011206f
C4073 vdd.n1088 gnd 0.00902f
C4074 vdd.n1089 gnd 0.011206f
C4075 vdd.n1090 gnd 0.00902f
C4076 vdd.n1091 gnd 0.011206f
C4077 vdd.t227 gnd 0.572603f
C4078 vdd.n1092 gnd 0.011206f
C4079 vdd.n1093 gnd 0.00902f
C4080 vdd.n1094 gnd 0.011206f
C4081 vdd.n1095 gnd 0.00902f
C4082 vdd.n1096 gnd 0.011206f
C4083 vdd.n1097 gnd 0.921891f
C4084 vdd.n1098 gnd 0.950521f
C4085 vdd.t5 gnd 0.572603f
C4086 vdd.n1099 gnd 0.011206f
C4087 vdd.n1100 gnd 0.00902f
C4088 vdd.n1101 gnd 0.011206f
C4089 vdd.n1102 gnd 0.00902f
C4090 vdd.n1103 gnd 0.011206f
C4091 vdd.n1104 gnd 0.727206f
C4092 vdd.n1105 gnd 0.011206f
C4093 vdd.n1106 gnd 0.00902f
C4094 vdd.n1107 gnd 0.011206f
C4095 vdd.n1108 gnd 0.00902f
C4096 vdd.n1109 gnd 0.011206f
C4097 vdd.t67 gnd 0.572603f
C4098 vdd.t50 gnd 0.572603f
C4099 vdd.n1110 gnd 0.011206f
C4100 vdd.n1111 gnd 0.00902f
C4101 vdd.n1112 gnd 0.011206f
C4102 vdd.n1113 gnd 0.00902f
C4103 vdd.n1114 gnd 0.011206f
C4104 vdd.t70 gnd 0.572603f
C4105 vdd.n1115 gnd 0.011206f
C4106 vdd.n1116 gnd 0.00902f
C4107 vdd.n1117 gnd 0.011206f
C4108 vdd.n1118 gnd 0.00902f
C4109 vdd.n1119 gnd 0.011206f
C4110 vdd.t59 gnd 0.572603f
C4111 vdd.n1120 gnd 0.807371f
C4112 vdd.n1121 gnd 0.011206f
C4113 vdd.n1122 gnd 0.00902f
C4114 vdd.n1123 gnd 0.011206f
C4115 vdd.n1124 gnd 0.00902f
C4116 vdd.n1125 gnd 0.011206f
C4117 vdd.n1126 gnd 0.898987f
C4118 vdd.n1127 gnd 0.011206f
C4119 vdd.n1128 gnd 0.00902f
C4120 vdd.n1129 gnd 0.011206f
C4121 vdd.n1130 gnd 0.00902f
C4122 vdd.n1131 gnd 0.011206f
C4123 vdd.n1132 gnd 0.704302f
C4124 vdd.t85 gnd 0.572603f
C4125 vdd.n1133 gnd 0.011206f
C4126 vdd.n1134 gnd 0.00902f
C4127 vdd.n1135 gnd 0.011206f
C4128 vdd.n1136 gnd 0.00902f
C4129 vdd.n1137 gnd 0.011206f
C4130 vdd.t115 gnd 0.572603f
C4131 vdd.n1138 gnd 0.011206f
C4132 vdd.n1139 gnd 0.00902f
C4133 vdd.n1140 gnd 0.011206f
C4134 vdd.n1141 gnd 0.00902f
C4135 vdd.n1142 gnd 0.011206f
C4136 vdd.t32 gnd 0.572603f
C4137 vdd.n1143 gnd 0.63559f
C4138 vdd.n1144 gnd 0.011206f
C4139 vdd.n1145 gnd 0.00902f
C4140 vdd.n1146 gnd 0.011206f
C4141 vdd.n1147 gnd 0.00902f
C4142 vdd.n1148 gnd 0.011206f
C4143 vdd.t28 gnd 0.572603f
C4144 vdd.n1149 gnd 0.011206f
C4145 vdd.n1150 gnd 0.00902f
C4146 vdd.n1151 gnd 0.011206f
C4147 vdd.n1152 gnd 0.00902f
C4148 vdd.n1153 gnd 0.011206f
C4149 vdd.n1154 gnd 0.876083f
C4150 vdd.n1155 gnd 0.950521f
C4151 vdd.t26 gnd 0.572603f
C4152 vdd.n1156 gnd 0.011206f
C4153 vdd.n1157 gnd 0.00902f
C4154 vdd.n1158 gnd 0.011206f
C4155 vdd.n1159 gnd 0.00902f
C4156 vdd.n1160 gnd 0.011206f
C4157 vdd.n1161 gnd 0.681398f
C4158 vdd.n1162 gnd 0.011206f
C4159 vdd.n1163 gnd 0.00902f
C4160 vdd.n1164 gnd 0.011206f
C4161 vdd.n1165 gnd 0.00902f
C4162 vdd.n1166 gnd 0.011206f
C4163 vdd.t54 gnd 0.572603f
C4164 vdd.t41 gnd 0.572603f
C4165 vdd.n1167 gnd 0.011206f
C4166 vdd.n1168 gnd 0.00902f
C4167 vdd.n1169 gnd 0.011206f
C4168 vdd.n1170 gnd 0.00902f
C4169 vdd.n1171 gnd 0.011206f
C4170 vdd.t39 gnd 0.572603f
C4171 vdd.n1172 gnd 0.011206f
C4172 vdd.n1173 gnd 0.00902f
C4173 vdd.n1174 gnd 0.011206f
C4174 vdd.n1175 gnd 0.00902f
C4175 vdd.n1176 gnd 0.011206f
C4176 vdd.t52 gnd 0.572603f
C4177 vdd.n1177 gnd 0.853179f
C4178 vdd.n1178 gnd 0.011206f
C4179 vdd.n1179 gnd 0.00902f
C4180 vdd.n1180 gnd 0.011206f
C4181 vdd.n1181 gnd 0.00902f
C4182 vdd.n1182 gnd 0.011206f
C4183 vdd.n1183 gnd 1.14521f
C4184 vdd.n1184 gnd 0.011206f
C4185 vdd.n1185 gnd 0.00902f
C4186 vdd.n1186 gnd 0.027108f
C4187 vdd.n1187 gnd 0.007486f
C4188 vdd.n1188 gnd 0.027108f
C4189 vdd.t160 gnd 0.572603f
C4190 vdd.n1189 gnd 0.027108f
C4191 vdd.n1190 gnd 0.007486f
C4192 vdd.n1191 gnd 0.011206f
C4193 vdd.n1192 gnd 0.00902f
C4194 vdd.n1193 gnd 0.011206f
C4195 vdd.n1224 gnd 0.027689f
C4196 vdd.n1225 gnd 1.68918f
C4197 vdd.n1226 gnd 0.011206f
C4198 vdd.n1227 gnd 0.00902f
C4199 vdd.n1228 gnd 0.011206f
C4200 vdd.n1229 gnd 0.011206f
C4201 vdd.n1230 gnd 0.011206f
C4202 vdd.n1231 gnd 0.011206f
C4203 vdd.n1232 gnd 0.011206f
C4204 vdd.n1233 gnd 0.00902f
C4205 vdd.n1234 gnd 0.011206f
C4206 vdd.n1235 gnd 0.011206f
C4207 vdd.n1236 gnd 0.011206f
C4208 vdd.n1237 gnd 0.011206f
C4209 vdd.n1238 gnd 0.011206f
C4210 vdd.n1239 gnd 0.00902f
C4211 vdd.n1240 gnd 0.011206f
C4212 vdd.n1241 gnd 0.011206f
C4213 vdd.n1242 gnd 0.011206f
C4214 vdd.n1243 gnd 0.011206f
C4215 vdd.n1244 gnd 0.011206f
C4216 vdd.n1245 gnd 0.00902f
C4217 vdd.n1246 gnd 0.011206f
C4218 vdd.n1247 gnd 0.011206f
C4219 vdd.n1248 gnd 0.011206f
C4220 vdd.n1249 gnd 0.011206f
C4221 vdd.n1250 gnd 0.011206f
C4222 vdd.t174 gnd 0.137864f
C4223 vdd.t175 gnd 0.147339f
C4224 vdd.t173 gnd 0.180049f
C4225 vdd.n1251 gnd 0.230797f
C4226 vdd.n1252 gnd 0.194813f
C4227 vdd.n1253 gnd 0.019302f
C4228 vdd.n1254 gnd 0.011206f
C4229 vdd.n1255 gnd 0.011206f
C4230 vdd.n1256 gnd 0.011206f
C4231 vdd.n1257 gnd 0.011206f
C4232 vdd.n1258 gnd 0.011206f
C4233 vdd.n1259 gnd 0.00902f
C4234 vdd.n1260 gnd 0.011206f
C4235 vdd.n1261 gnd 0.011206f
C4236 vdd.n1262 gnd 0.011206f
C4237 vdd.n1263 gnd 0.011206f
C4238 vdd.n1264 gnd 0.011206f
C4239 vdd.n1265 gnd 0.00902f
C4240 vdd.n1266 gnd 0.011206f
C4241 vdd.n1267 gnd 0.011206f
C4242 vdd.n1268 gnd 0.011206f
C4243 vdd.n1269 gnd 0.011206f
C4244 vdd.n1270 gnd 0.011206f
C4245 vdd.n1271 gnd 0.00902f
C4246 vdd.n1272 gnd 0.011206f
C4247 vdd.n1273 gnd 0.011206f
C4248 vdd.n1274 gnd 0.011206f
C4249 vdd.n1275 gnd 0.011206f
C4250 vdd.n1276 gnd 0.011206f
C4251 vdd.n1277 gnd 0.00902f
C4252 vdd.n1278 gnd 0.011206f
C4253 vdd.n1279 gnd 0.011206f
C4254 vdd.n1280 gnd 0.011206f
C4255 vdd.n1281 gnd 0.011206f
C4256 vdd.n1282 gnd 0.011206f
C4257 vdd.n1283 gnd 0.00902f
C4258 vdd.n1284 gnd 0.011206f
C4259 vdd.n1285 gnd 0.011206f
C4260 vdd.n1286 gnd 0.011206f
C4261 vdd.n1287 gnd 0.011206f
C4262 vdd.n1288 gnd 0.00902f
C4263 vdd.n1289 gnd 0.011206f
C4264 vdd.n1290 gnd 0.011206f
C4265 vdd.n1291 gnd 0.011206f
C4266 vdd.n1292 gnd 0.011206f
C4267 vdd.n1293 gnd 0.011206f
C4268 vdd.n1294 gnd 0.00902f
C4269 vdd.n1295 gnd 0.011206f
C4270 vdd.n1296 gnd 0.011206f
C4271 vdd.n1297 gnd 0.011206f
C4272 vdd.n1298 gnd 0.011206f
C4273 vdd.n1299 gnd 0.011206f
C4274 vdd.n1300 gnd 0.00902f
C4275 vdd.n1301 gnd 0.011206f
C4276 vdd.n1302 gnd 0.011206f
C4277 vdd.n1303 gnd 0.011206f
C4278 vdd.n1304 gnd 0.011206f
C4279 vdd.n1305 gnd 0.011206f
C4280 vdd.n1306 gnd 0.00902f
C4281 vdd.n1307 gnd 0.011206f
C4282 vdd.n1308 gnd 0.011206f
C4283 vdd.n1309 gnd 0.011206f
C4284 vdd.n1310 gnd 0.011206f
C4285 vdd.n1311 gnd 0.011206f
C4286 vdd.n1312 gnd 0.00902f
C4287 vdd.n1313 gnd 0.011206f
C4288 vdd.n1314 gnd 0.011206f
C4289 vdd.n1315 gnd 0.011206f
C4290 vdd.n1316 gnd 0.011206f
C4291 vdd.t171 gnd 0.137864f
C4292 vdd.t172 gnd 0.147339f
C4293 vdd.t170 gnd 0.180049f
C4294 vdd.n1317 gnd 0.230797f
C4295 vdd.n1318 gnd 0.194813f
C4296 vdd.n1319 gnd 0.014792f
C4297 vdd.n1320 gnd 0.004284f
C4298 vdd.n1321 gnd 0.027689f
C4299 vdd.n1322 gnd 0.011206f
C4300 vdd.n1323 gnd 0.004735f
C4301 vdd.n1324 gnd 0.00902f
C4302 vdd.n1325 gnd 0.00902f
C4303 vdd.n1326 gnd 0.011206f
C4304 vdd.n1327 gnd 0.011206f
C4305 vdd.n1328 gnd 0.011206f
C4306 vdd.n1329 gnd 0.00902f
C4307 vdd.n1330 gnd 0.00902f
C4308 vdd.n1331 gnd 0.00902f
C4309 vdd.n1332 gnd 0.011206f
C4310 vdd.n1333 gnd 0.011206f
C4311 vdd.n1334 gnd 0.011206f
C4312 vdd.n1335 gnd 0.00902f
C4313 vdd.n1336 gnd 0.00902f
C4314 vdd.n1337 gnd 0.00902f
C4315 vdd.n1338 gnd 0.011206f
C4316 vdd.n1339 gnd 0.011206f
C4317 vdd.n1340 gnd 0.011206f
C4318 vdd.n1341 gnd 0.00902f
C4319 vdd.n1342 gnd 0.00902f
C4320 vdd.n1343 gnd 0.00902f
C4321 vdd.n1344 gnd 0.011206f
C4322 vdd.n1345 gnd 0.011206f
C4323 vdd.n1346 gnd 0.011206f
C4324 vdd.n1347 gnd 0.00902f
C4325 vdd.n1348 gnd 0.00902f
C4326 vdd.n1349 gnd 0.00902f
C4327 vdd.n1350 gnd 0.011206f
C4328 vdd.n1351 gnd 0.011206f
C4329 vdd.n1352 gnd 0.011206f
C4330 vdd.n1353 gnd 0.008929f
C4331 vdd.n1354 gnd 0.011206f
C4332 vdd.t161 gnd 0.137864f
C4333 vdd.t162 gnd 0.147339f
C4334 vdd.t159 gnd 0.180049f
C4335 vdd.n1355 gnd 0.230797f
C4336 vdd.n1356 gnd 0.194813f
C4337 vdd.n1357 gnd 0.019302f
C4338 vdd.n1358 gnd 0.006133f
C4339 vdd.n1359 gnd 0.011206f
C4340 vdd.n1360 gnd 0.011206f
C4341 vdd.n1361 gnd 0.011206f
C4342 vdd.n1362 gnd 0.00902f
C4343 vdd.n1363 gnd 0.00902f
C4344 vdd.n1364 gnd 0.00902f
C4345 vdd.n1365 gnd 0.011206f
C4346 vdd.n1366 gnd 0.011206f
C4347 vdd.n1367 gnd 0.011206f
C4348 vdd.n1368 gnd 0.00902f
C4349 vdd.n1369 gnd 0.00902f
C4350 vdd.n1370 gnd 0.00902f
C4351 vdd.n1371 gnd 0.011206f
C4352 vdd.n1372 gnd 0.011206f
C4353 vdd.n1373 gnd 0.011206f
C4354 vdd.n1374 gnd 0.00902f
C4355 vdd.n1375 gnd 0.00902f
C4356 vdd.n1376 gnd 0.00902f
C4357 vdd.n1377 gnd 0.011206f
C4358 vdd.n1378 gnd 0.011206f
C4359 vdd.n1379 gnd 0.011206f
C4360 vdd.n1380 gnd 0.00902f
C4361 vdd.n1381 gnd 0.00902f
C4362 vdd.n1382 gnd 0.00902f
C4363 vdd.n1383 gnd 0.011206f
C4364 vdd.n1384 gnd 0.011206f
C4365 vdd.n1385 gnd 0.011206f
C4366 vdd.n1386 gnd 0.00902f
C4367 vdd.n1387 gnd 0.00902f
C4368 vdd.n1388 gnd 0.007531f
C4369 vdd.n1389 gnd 0.011206f
C4370 vdd.n1390 gnd 0.011206f
C4371 vdd.n1391 gnd 0.011206f
C4372 vdd.n1392 gnd 0.007531f
C4373 vdd.n1393 gnd 0.00902f
C4374 vdd.n1394 gnd 0.00902f
C4375 vdd.n1395 gnd 0.011206f
C4376 vdd.n1396 gnd 0.011206f
C4377 vdd.n1397 gnd 0.011206f
C4378 vdd.n1398 gnd 0.00902f
C4379 vdd.n1399 gnd 0.00902f
C4380 vdd.n1400 gnd 0.00902f
C4381 vdd.n1401 gnd 0.011206f
C4382 vdd.n1402 gnd 0.011206f
C4383 vdd.n1403 gnd 0.011206f
C4384 vdd.n1404 gnd 0.00902f
C4385 vdd.n1405 gnd 0.00902f
C4386 vdd.n1406 gnd 0.00902f
C4387 vdd.n1407 gnd 0.011206f
C4388 vdd.n1408 gnd 0.011206f
C4389 vdd.n1409 gnd 0.011206f
C4390 vdd.n1410 gnd 0.00902f
C4391 vdd.n1411 gnd 0.00902f
C4392 vdd.n1412 gnd 0.00902f
C4393 vdd.n1413 gnd 0.011206f
C4394 vdd.n1414 gnd 0.011206f
C4395 vdd.n1415 gnd 0.011206f
C4396 vdd.n1416 gnd 0.00902f
C4397 vdd.n1417 gnd 0.011206f
C4398 vdd.n1418 gnd 2.71414f
C4399 vdd.n1420 gnd 0.027689f
C4400 vdd.n1421 gnd 0.007486f
C4401 vdd.n1422 gnd 0.027689f
C4402 vdd.n1423 gnd 0.027108f
C4403 vdd.n1424 gnd 0.011206f
C4404 vdd.n1425 gnd 0.00902f
C4405 vdd.n1426 gnd 0.011206f
C4406 vdd.n1427 gnd 0.578329f
C4407 vdd.n1428 gnd 0.011206f
C4408 vdd.n1429 gnd 0.00902f
C4409 vdd.n1430 gnd 0.011206f
C4410 vdd.n1431 gnd 0.011206f
C4411 vdd.n1432 gnd 0.011206f
C4412 vdd.n1433 gnd 0.00902f
C4413 vdd.n1434 gnd 0.011206f
C4414 vdd.n1435 gnd 1.04786f
C4415 vdd.n1436 gnd 1.14521f
C4416 vdd.n1437 gnd 0.011206f
C4417 vdd.n1438 gnd 0.00902f
C4418 vdd.n1439 gnd 0.011206f
C4419 vdd.n1440 gnd 0.011206f
C4420 vdd.n1441 gnd 0.011206f
C4421 vdd.n1442 gnd 0.00902f
C4422 vdd.n1443 gnd 0.011206f
C4423 vdd.n1444 gnd 0.669946f
C4424 vdd.n1445 gnd 0.011206f
C4425 vdd.n1446 gnd 0.00902f
C4426 vdd.n1447 gnd 0.011206f
C4427 vdd.n1448 gnd 0.011206f
C4428 vdd.n1449 gnd 0.011206f
C4429 vdd.n1450 gnd 0.00902f
C4430 vdd.n1451 gnd 0.011206f
C4431 vdd.n1452 gnd 0.658494f
C4432 vdd.n1453 gnd 0.864631f
C4433 vdd.n1454 gnd 0.011206f
C4434 vdd.n1455 gnd 0.00902f
C4435 vdd.n1456 gnd 0.011206f
C4436 vdd.n1457 gnd 0.011206f
C4437 vdd.n1458 gnd 0.011206f
C4438 vdd.n1459 gnd 0.00902f
C4439 vdd.n1460 gnd 0.011206f
C4440 vdd.n1461 gnd 0.950521f
C4441 vdd.n1462 gnd 0.011206f
C4442 vdd.n1463 gnd 0.00902f
C4443 vdd.n1464 gnd 0.011206f
C4444 vdd.n1465 gnd 0.011206f
C4445 vdd.n1466 gnd 0.011206f
C4446 vdd.n1467 gnd 0.00902f
C4447 vdd.n1468 gnd 0.011206f
C4448 vdd.t87 gnd 0.572603f
C4449 vdd.n1469 gnd 0.841727f
C4450 vdd.n1470 gnd 0.011206f
C4451 vdd.n1471 gnd 0.00902f
C4452 vdd.n1472 gnd 0.011206f
C4453 vdd.n1473 gnd 0.011206f
C4454 vdd.n1474 gnd 0.011206f
C4455 vdd.n1475 gnd 0.00902f
C4456 vdd.n1476 gnd 0.011206f
C4457 vdd.n1477 gnd 0.647042f
C4458 vdd.n1478 gnd 0.011206f
C4459 vdd.n1479 gnd 0.00902f
C4460 vdd.n1480 gnd 0.011206f
C4461 vdd.n1481 gnd 0.011206f
C4462 vdd.n1482 gnd 0.011206f
C4463 vdd.n1483 gnd 0.00902f
C4464 vdd.n1484 gnd 0.011206f
C4465 vdd.n1485 gnd 0.830275f
C4466 vdd.n1486 gnd 0.69285f
C4467 vdd.n1487 gnd 0.011206f
C4468 vdd.n1488 gnd 0.00902f
C4469 vdd.n1489 gnd 0.011206f
C4470 vdd.n1490 gnd 0.011206f
C4471 vdd.n1491 gnd 0.011206f
C4472 vdd.n1492 gnd 0.00902f
C4473 vdd.n1493 gnd 0.011206f
C4474 vdd.n1494 gnd 0.887535f
C4475 vdd.n1495 gnd 0.011206f
C4476 vdd.n1496 gnd 0.00902f
C4477 vdd.n1497 gnd 0.011206f
C4478 vdd.n1498 gnd 0.011206f
C4479 vdd.n1499 gnd 0.011206f
C4480 vdd.n1500 gnd 0.00902f
C4481 vdd.n1501 gnd 0.011206f
C4482 vdd.t43 gnd 0.572603f
C4483 vdd.n1502 gnd 0.950521f
C4484 vdd.n1503 gnd 0.011206f
C4485 vdd.n1504 gnd 0.00902f
C4486 vdd.n1505 gnd 0.011206f
C4487 vdd.n1506 gnd 0.008613f
C4488 vdd.n1507 gnd 0.00615f
C4489 vdd.n1508 gnd 0.005707f
C4490 vdd.n1509 gnd 0.003157f
C4491 vdd.n1510 gnd 0.007248f
C4492 vdd.n1511 gnd 0.003067f
C4493 vdd.n1512 gnd 0.003247f
C4494 vdd.n1513 gnd 0.005707f
C4495 vdd.n1514 gnd 0.003067f
C4496 vdd.n1515 gnd 0.007248f
C4497 vdd.n1516 gnd 0.003247f
C4498 vdd.n1517 gnd 0.005707f
C4499 vdd.n1518 gnd 0.003067f
C4500 vdd.n1519 gnd 0.005436f
C4501 vdd.n1520 gnd 0.005453f
C4502 vdd.t62 gnd 0.015573f
C4503 vdd.n1521 gnd 0.034649f
C4504 vdd.n1522 gnd 0.180321f
C4505 vdd.n1523 gnd 0.003067f
C4506 vdd.n1524 gnd 0.003247f
C4507 vdd.n1525 gnd 0.007248f
C4508 vdd.n1526 gnd 0.007248f
C4509 vdd.n1527 gnd 0.003247f
C4510 vdd.n1528 gnd 0.003067f
C4511 vdd.n1529 gnd 0.005707f
C4512 vdd.n1530 gnd 0.005707f
C4513 vdd.n1531 gnd 0.003067f
C4514 vdd.n1532 gnd 0.003247f
C4515 vdd.n1533 gnd 0.007248f
C4516 vdd.n1534 gnd 0.007248f
C4517 vdd.n1535 gnd 0.003247f
C4518 vdd.n1536 gnd 0.003067f
C4519 vdd.n1537 gnd 0.005707f
C4520 vdd.n1538 gnd 0.005707f
C4521 vdd.n1539 gnd 0.003067f
C4522 vdd.n1540 gnd 0.003247f
C4523 vdd.n1541 gnd 0.007248f
C4524 vdd.n1542 gnd 0.007248f
C4525 vdd.n1543 gnd 0.017137f
C4526 vdd.n1544 gnd 0.003157f
C4527 vdd.n1545 gnd 0.003067f
C4528 vdd.n1546 gnd 0.014751f
C4529 vdd.n1547 gnd 0.010298f
C4530 vdd.t281 gnd 0.036078f
C4531 vdd.t231 gnd 0.036078f
C4532 vdd.n1548 gnd 0.247954f
C4533 vdd.n1549 gnd 0.194978f
C4534 vdd.t51 gnd 0.036078f
C4535 vdd.t221 gnd 0.036078f
C4536 vdd.n1550 gnd 0.247954f
C4537 vdd.n1551 gnd 0.157346f
C4538 vdd.t71 gnd 0.036078f
C4539 vdd.t222 gnd 0.036078f
C4540 vdd.n1552 gnd 0.247954f
C4541 vdd.n1553 gnd 0.157346f
C4542 vdd.t77 gnd 0.036078f
C4543 vdd.t295 gnd 0.036078f
C4544 vdd.n1554 gnd 0.247954f
C4545 vdd.n1555 gnd 0.157346f
C4546 vdd.t44 gnd 0.036078f
C4547 vdd.t86 gnd 0.036078f
C4548 vdd.n1556 gnd 0.247954f
C4549 vdd.n1557 gnd 0.157346f
C4550 vdd.t56 gnd 0.036078f
C4551 vdd.t116 gnd 0.036078f
C4552 vdd.n1558 gnd 0.247954f
C4553 vdd.n1559 gnd 0.157346f
C4554 vdd.t226 gnd 0.036078f
C4555 vdd.t79 gnd 0.036078f
C4556 vdd.n1560 gnd 0.247954f
C4557 vdd.n1561 gnd 0.157346f
C4558 vdd.t124 gnd 0.036078f
C4559 vdd.t93 gnd 0.036078f
C4560 vdd.n1562 gnd 0.247954f
C4561 vdd.n1563 gnd 0.157346f
C4562 vdd.t123 gnd 0.036078f
C4563 vdd.t112 gnd 0.036078f
C4564 vdd.n1564 gnd 0.247954f
C4565 vdd.n1565 gnd 0.157346f
C4566 vdd.n1566 gnd 0.00615f
C4567 vdd.n1567 gnd 0.005707f
C4568 vdd.n1568 gnd 0.003157f
C4569 vdd.n1569 gnd 0.007248f
C4570 vdd.n1570 gnd 0.003067f
C4571 vdd.n1571 gnd 0.003247f
C4572 vdd.n1572 gnd 0.005707f
C4573 vdd.n1573 gnd 0.003067f
C4574 vdd.n1574 gnd 0.007248f
C4575 vdd.n1575 gnd 0.003247f
C4576 vdd.n1576 gnd 0.005707f
C4577 vdd.n1577 gnd 0.003067f
C4578 vdd.n1578 gnd 0.005436f
C4579 vdd.n1579 gnd 0.005453f
C4580 vdd.t53 gnd 0.015573f
C4581 vdd.n1580 gnd 0.034649f
C4582 vdd.n1581 gnd 0.180321f
C4583 vdd.n1582 gnd 0.003067f
C4584 vdd.n1583 gnd 0.003247f
C4585 vdd.n1584 gnd 0.007248f
C4586 vdd.n1585 gnd 0.007248f
C4587 vdd.n1586 gnd 0.003247f
C4588 vdd.n1587 gnd 0.003067f
C4589 vdd.n1588 gnd 0.005707f
C4590 vdd.n1589 gnd 0.005707f
C4591 vdd.n1590 gnd 0.003067f
C4592 vdd.n1591 gnd 0.003247f
C4593 vdd.n1592 gnd 0.007248f
C4594 vdd.n1593 gnd 0.007248f
C4595 vdd.n1594 gnd 0.003247f
C4596 vdd.n1595 gnd 0.003067f
C4597 vdd.n1596 gnd 0.005707f
C4598 vdd.n1597 gnd 0.005707f
C4599 vdd.n1598 gnd 0.003067f
C4600 vdd.n1599 gnd 0.003247f
C4601 vdd.n1600 gnd 0.007248f
C4602 vdd.n1601 gnd 0.007248f
C4603 vdd.n1602 gnd 0.017137f
C4604 vdd.n1603 gnd 0.003157f
C4605 vdd.n1604 gnd 0.003067f
C4606 vdd.n1605 gnd 0.014751f
C4607 vdd.n1606 gnd 0.009975f
C4608 vdd.n1607 gnd 0.117066f
C4609 vdd.n1608 gnd 0.00615f
C4610 vdd.n1609 gnd 0.005707f
C4611 vdd.n1610 gnd 0.003157f
C4612 vdd.n1611 gnd 0.007248f
C4613 vdd.n1612 gnd 0.003067f
C4614 vdd.n1613 gnd 0.003247f
C4615 vdd.n1614 gnd 0.005707f
C4616 vdd.n1615 gnd 0.003067f
C4617 vdd.n1616 gnd 0.007248f
C4618 vdd.n1617 gnd 0.003247f
C4619 vdd.n1618 gnd 0.005707f
C4620 vdd.n1619 gnd 0.003067f
C4621 vdd.n1620 gnd 0.005436f
C4622 vdd.n1621 gnd 0.005453f
C4623 vdd.t282 gnd 0.015573f
C4624 vdd.n1622 gnd 0.034649f
C4625 vdd.n1623 gnd 0.180321f
C4626 vdd.n1624 gnd 0.003067f
C4627 vdd.n1625 gnd 0.003247f
C4628 vdd.n1626 gnd 0.007248f
C4629 vdd.n1627 gnd 0.007248f
C4630 vdd.n1628 gnd 0.003247f
C4631 vdd.n1629 gnd 0.003067f
C4632 vdd.n1630 gnd 0.005707f
C4633 vdd.n1631 gnd 0.005707f
C4634 vdd.n1632 gnd 0.003067f
C4635 vdd.n1633 gnd 0.003247f
C4636 vdd.n1634 gnd 0.007248f
C4637 vdd.n1635 gnd 0.007248f
C4638 vdd.n1636 gnd 0.003247f
C4639 vdd.n1637 gnd 0.003067f
C4640 vdd.n1638 gnd 0.005707f
C4641 vdd.n1639 gnd 0.005707f
C4642 vdd.n1640 gnd 0.003067f
C4643 vdd.n1641 gnd 0.003247f
C4644 vdd.n1642 gnd 0.007248f
C4645 vdd.n1643 gnd 0.007248f
C4646 vdd.n1644 gnd 0.017137f
C4647 vdd.n1645 gnd 0.003157f
C4648 vdd.n1646 gnd 0.003067f
C4649 vdd.n1647 gnd 0.014751f
C4650 vdd.n1648 gnd 0.010298f
C4651 vdd.t6 gnd 0.036078f
C4652 vdd.t228 gnd 0.036078f
C4653 vdd.n1649 gnd 0.247954f
C4654 vdd.n1650 gnd 0.194978f
C4655 vdd.t102 gnd 0.036078f
C4656 vdd.t58 gnd 0.036078f
C4657 vdd.n1651 gnd 0.247954f
C4658 vdd.n1652 gnd 0.157346f
C4659 vdd.t92 gnd 0.036078f
C4660 vdd.t114 gnd 0.036078f
C4661 vdd.n1653 gnd 0.247954f
C4662 vdd.n1654 gnd 0.157346f
C4663 vdd.t288 gnd 0.036078f
C4664 vdd.t60 gnd 0.036078f
C4665 vdd.n1655 gnd 0.247954f
C4666 vdd.n1656 gnd 0.157346f
C4667 vdd.t133 gnd 0.036078f
C4668 vdd.t109 gnd 0.036078f
C4669 vdd.n1657 gnd 0.247954f
C4670 vdd.n1658 gnd 0.157346f
C4671 vdd.t33 gnd 0.036078f
C4672 vdd.t132 gnd 0.036078f
C4673 vdd.n1659 gnd 0.247954f
C4674 vdd.n1660 gnd 0.157346f
C4675 vdd.t120 gnd 0.036078f
C4676 vdd.t121 gnd 0.036078f
C4677 vdd.n1661 gnd 0.247954f
C4678 vdd.n1662 gnd 0.157346f
C4679 vdd.t111 gnd 0.036078f
C4680 vdd.t88 gnd 0.036078f
C4681 vdd.n1663 gnd 0.247954f
C4682 vdd.n1664 gnd 0.157346f
C4683 vdd.t113 gnd 0.036078f
C4684 vdd.t55 gnd 0.036078f
C4685 vdd.n1665 gnd 0.247954f
C4686 vdd.n1666 gnd 0.157346f
C4687 vdd.n1667 gnd 0.00615f
C4688 vdd.n1668 gnd 0.005707f
C4689 vdd.n1669 gnd 0.003157f
C4690 vdd.n1670 gnd 0.007248f
C4691 vdd.n1671 gnd 0.003067f
C4692 vdd.n1672 gnd 0.003247f
C4693 vdd.n1673 gnd 0.005707f
C4694 vdd.n1674 gnd 0.003067f
C4695 vdd.n1675 gnd 0.007248f
C4696 vdd.n1676 gnd 0.003247f
C4697 vdd.n1677 gnd 0.005707f
C4698 vdd.n1678 gnd 0.003067f
C4699 vdd.n1679 gnd 0.005436f
C4700 vdd.n1680 gnd 0.005453f
C4701 vdd.t63 gnd 0.015573f
C4702 vdd.n1681 gnd 0.034649f
C4703 vdd.n1682 gnd 0.180321f
C4704 vdd.n1683 gnd 0.003067f
C4705 vdd.n1684 gnd 0.003247f
C4706 vdd.n1685 gnd 0.007248f
C4707 vdd.n1686 gnd 0.007248f
C4708 vdd.n1687 gnd 0.003247f
C4709 vdd.n1688 gnd 0.003067f
C4710 vdd.n1689 gnd 0.005707f
C4711 vdd.n1690 gnd 0.005707f
C4712 vdd.n1691 gnd 0.003067f
C4713 vdd.n1692 gnd 0.003247f
C4714 vdd.n1693 gnd 0.007248f
C4715 vdd.n1694 gnd 0.007248f
C4716 vdd.n1695 gnd 0.003247f
C4717 vdd.n1696 gnd 0.003067f
C4718 vdd.n1697 gnd 0.005707f
C4719 vdd.n1698 gnd 0.005707f
C4720 vdd.n1699 gnd 0.003067f
C4721 vdd.n1700 gnd 0.003247f
C4722 vdd.n1701 gnd 0.007248f
C4723 vdd.n1702 gnd 0.007248f
C4724 vdd.n1703 gnd 0.017137f
C4725 vdd.n1704 gnd 0.003157f
C4726 vdd.n1705 gnd 0.003067f
C4727 vdd.n1706 gnd 0.014751f
C4728 vdd.n1707 gnd 0.009975f
C4729 vdd.n1708 gnd 0.069642f
C4730 vdd.n1709 gnd 0.25094f
C4731 vdd.n1710 gnd 0.00615f
C4732 vdd.n1711 gnd 0.005707f
C4733 vdd.n1712 gnd 0.003157f
C4734 vdd.n1713 gnd 0.007248f
C4735 vdd.n1714 gnd 0.003067f
C4736 vdd.n1715 gnd 0.003247f
C4737 vdd.n1716 gnd 0.005707f
C4738 vdd.n1717 gnd 0.003067f
C4739 vdd.n1718 gnd 0.007248f
C4740 vdd.n1719 gnd 0.003247f
C4741 vdd.n1720 gnd 0.005707f
C4742 vdd.n1721 gnd 0.003067f
C4743 vdd.n1722 gnd 0.005436f
C4744 vdd.n1723 gnd 0.005453f
C4745 vdd.t291 gnd 0.015573f
C4746 vdd.n1724 gnd 0.034649f
C4747 vdd.n1725 gnd 0.180321f
C4748 vdd.n1726 gnd 0.003067f
C4749 vdd.n1727 gnd 0.003247f
C4750 vdd.n1728 gnd 0.007248f
C4751 vdd.n1729 gnd 0.007248f
C4752 vdd.n1730 gnd 0.003247f
C4753 vdd.n1731 gnd 0.003067f
C4754 vdd.n1732 gnd 0.005707f
C4755 vdd.n1733 gnd 0.005707f
C4756 vdd.n1734 gnd 0.003067f
C4757 vdd.n1735 gnd 0.003247f
C4758 vdd.n1736 gnd 0.007248f
C4759 vdd.n1737 gnd 0.007248f
C4760 vdd.n1738 gnd 0.003247f
C4761 vdd.n1739 gnd 0.003067f
C4762 vdd.n1740 gnd 0.005707f
C4763 vdd.n1741 gnd 0.005707f
C4764 vdd.n1742 gnd 0.003067f
C4765 vdd.n1743 gnd 0.003247f
C4766 vdd.n1744 gnd 0.007248f
C4767 vdd.n1745 gnd 0.007248f
C4768 vdd.n1746 gnd 0.017137f
C4769 vdd.n1747 gnd 0.003157f
C4770 vdd.n1748 gnd 0.003067f
C4771 vdd.n1749 gnd 0.014751f
C4772 vdd.n1750 gnd 0.010298f
C4773 vdd.t276 gnd 0.036078f
C4774 vdd.t290 gnd 0.036078f
C4775 vdd.n1751 gnd 0.247954f
C4776 vdd.n1752 gnd 0.194978f
C4777 vdd.t289 gnd 0.036078f
C4778 vdd.t101 gnd 0.036078f
C4779 vdd.n1753 gnd 0.247954f
C4780 vdd.n1754 gnd 0.157346f
C4781 vdd.t78 gnd 0.036078f
C4782 vdd.t68 gnd 0.036078f
C4783 vdd.n1755 gnd 0.247954f
C4784 vdd.n1756 gnd 0.157346f
C4785 vdd.t84 gnd 0.036078f
C4786 vdd.t220 gnd 0.036078f
C4787 vdd.n1757 gnd 0.247954f
C4788 vdd.n1758 gnd 0.157346f
C4789 vdd.t128 gnd 0.036078f
C4790 vdd.t110 gnd 0.036078f
C4791 vdd.n1759 gnd 0.247954f
C4792 vdd.n1760 gnd 0.157346f
C4793 vdd.t69 gnd 0.036078f
C4794 vdd.t127 gnd 0.036078f
C4795 vdd.n1761 gnd 0.247954f
C4796 vdd.n1762 gnd 0.157346f
C4797 vdd.t27 gnd 0.036078f
C4798 vdd.t29 gnd 0.036078f
C4799 vdd.n1763 gnd 0.247954f
C4800 vdd.n1764 gnd 0.157346f
C4801 vdd.t42 gnd 0.036078f
C4802 vdd.t279 gnd 0.036078f
C4803 vdd.n1765 gnd 0.247954f
C4804 vdd.n1766 gnd 0.157346f
C4805 vdd.t40 gnd 0.036078f
C4806 vdd.t130 gnd 0.036078f
C4807 vdd.n1767 gnd 0.247954f
C4808 vdd.n1768 gnd 0.157346f
C4809 vdd.n1769 gnd 0.00615f
C4810 vdd.n1770 gnd 0.005707f
C4811 vdd.n1771 gnd 0.003157f
C4812 vdd.n1772 gnd 0.007248f
C4813 vdd.n1773 gnd 0.003067f
C4814 vdd.n1774 gnd 0.003247f
C4815 vdd.n1775 gnd 0.005707f
C4816 vdd.n1776 gnd 0.003067f
C4817 vdd.n1777 gnd 0.007248f
C4818 vdd.n1778 gnd 0.003247f
C4819 vdd.n1779 gnd 0.005707f
C4820 vdd.n1780 gnd 0.003067f
C4821 vdd.n1781 gnd 0.005436f
C4822 vdd.n1782 gnd 0.005453f
C4823 vdd.t66 gnd 0.015573f
C4824 vdd.n1783 gnd 0.034649f
C4825 vdd.n1784 gnd 0.180321f
C4826 vdd.n1785 gnd 0.003067f
C4827 vdd.n1786 gnd 0.003247f
C4828 vdd.n1787 gnd 0.007248f
C4829 vdd.n1788 gnd 0.007248f
C4830 vdd.n1789 gnd 0.003247f
C4831 vdd.n1790 gnd 0.003067f
C4832 vdd.n1791 gnd 0.005707f
C4833 vdd.n1792 gnd 0.005707f
C4834 vdd.n1793 gnd 0.003067f
C4835 vdd.n1794 gnd 0.003247f
C4836 vdd.n1795 gnd 0.007248f
C4837 vdd.n1796 gnd 0.007248f
C4838 vdd.n1797 gnd 0.003247f
C4839 vdd.n1798 gnd 0.003067f
C4840 vdd.n1799 gnd 0.005707f
C4841 vdd.n1800 gnd 0.005707f
C4842 vdd.n1801 gnd 0.003067f
C4843 vdd.n1802 gnd 0.003247f
C4844 vdd.n1803 gnd 0.007248f
C4845 vdd.n1804 gnd 0.007248f
C4846 vdd.n1805 gnd 0.017137f
C4847 vdd.n1806 gnd 0.003157f
C4848 vdd.n1807 gnd 0.003067f
C4849 vdd.n1808 gnd 0.014751f
C4850 vdd.n1809 gnd 0.009975f
C4851 vdd.n1810 gnd 0.069642f
C4852 vdd.n1811 gnd 0.287272f
C4853 vdd.n1812 gnd 2.87816f
C4854 vdd.n1813 gnd 0.660976f
C4855 vdd.n1814 gnd 0.008613f
C4856 vdd.n1815 gnd 0.00902f
C4857 vdd.n1816 gnd 0.011206f
C4858 vdd.n1817 gnd 0.818823f
C4859 vdd.n1818 gnd 0.011206f
C4860 vdd.n1819 gnd 0.00902f
C4861 vdd.n1820 gnd 0.011206f
C4862 vdd.n1821 gnd 0.011206f
C4863 vdd.n1822 gnd 0.011206f
C4864 vdd.n1823 gnd 0.00902f
C4865 vdd.n1824 gnd 0.011206f
C4866 vdd.n1825 gnd 0.950521f
C4867 vdd.t76 gnd 0.572603f
C4868 vdd.n1826 gnd 0.624138f
C4869 vdd.n1827 gnd 0.011206f
C4870 vdd.n1828 gnd 0.00902f
C4871 vdd.n1829 gnd 0.011206f
C4872 vdd.n1830 gnd 0.011206f
C4873 vdd.n1831 gnd 0.011206f
C4874 vdd.n1832 gnd 0.00902f
C4875 vdd.n1833 gnd 0.011206f
C4876 vdd.n1834 gnd 0.715754f
C4877 vdd.n1835 gnd 0.011206f
C4878 vdd.n1836 gnd 0.00902f
C4879 vdd.n1837 gnd 0.011206f
C4880 vdd.n1838 gnd 0.011206f
C4881 vdd.n1839 gnd 0.011206f
C4882 vdd.n1840 gnd 0.00902f
C4883 vdd.n1841 gnd 0.011206f
C4884 vdd.n1842 gnd 0.612685f
C4885 vdd.n1843 gnd 0.910439f
C4886 vdd.n1844 gnd 0.011206f
C4887 vdd.n1845 gnd 0.00902f
C4888 vdd.n1846 gnd 0.011206f
C4889 vdd.n1847 gnd 0.011206f
C4890 vdd.n1848 gnd 0.011206f
C4891 vdd.n1849 gnd 0.00902f
C4892 vdd.n1850 gnd 0.011206f
C4893 vdd.n1851 gnd 0.950521f
C4894 vdd.n1852 gnd 0.011206f
C4895 vdd.n1853 gnd 0.00902f
C4896 vdd.n1854 gnd 0.011206f
C4897 vdd.n1855 gnd 0.011206f
C4898 vdd.n1856 gnd 0.011206f
C4899 vdd.n1857 gnd 0.00902f
C4900 vdd.n1858 gnd 0.011206f
C4901 vdd.t57 gnd 0.572603f
C4902 vdd.n1859 gnd 0.795919f
C4903 vdd.n1860 gnd 0.011206f
C4904 vdd.n1861 gnd 0.00902f
C4905 vdd.n1862 gnd 0.011206f
C4906 vdd.n1863 gnd 0.011206f
C4907 vdd.n1864 gnd 0.011206f
C4908 vdd.n1865 gnd 0.00902f
C4909 vdd.n1866 gnd 0.011206f
C4910 vdd.n1867 gnd 0.601233f
C4911 vdd.n1868 gnd 0.011206f
C4912 vdd.n1869 gnd 0.00902f
C4913 vdd.n1870 gnd 0.011206f
C4914 vdd.n1871 gnd 0.011206f
C4915 vdd.n1872 gnd 0.011206f
C4916 vdd.n1873 gnd 0.00902f
C4917 vdd.n1874 gnd 0.011206f
C4918 vdd.n1875 gnd 0.784466f
C4919 vdd.n1876 gnd 0.738658f
C4920 vdd.n1877 gnd 0.011206f
C4921 vdd.n1878 gnd 0.00902f
C4922 vdd.n1879 gnd 0.011206f
C4923 vdd.n1880 gnd 0.011206f
C4924 vdd.n1881 gnd 0.011206f
C4925 vdd.n1882 gnd 0.00902f
C4926 vdd.n1883 gnd 0.011206f
C4927 vdd.n1884 gnd 0.933343f
C4928 vdd.n1885 gnd 0.011206f
C4929 vdd.n1886 gnd 0.00902f
C4930 vdd.n1887 gnd 0.011206f
C4931 vdd.n1888 gnd 0.011206f
C4932 vdd.n1889 gnd 0.027108f
C4933 vdd.n1890 gnd 0.011206f
C4934 vdd.n1891 gnd 0.011206f
C4935 vdd.n1892 gnd 0.00902f
C4936 vdd.n1893 gnd 0.011206f
C4937 vdd.n1894 gnd 0.69285f
C4938 vdd.n1895 gnd 1.14521f
C4939 vdd.n1896 gnd 0.011206f
C4940 vdd.n1897 gnd 0.00902f
C4941 vdd.n1898 gnd 0.011206f
C4942 vdd.n1899 gnd 0.011206f
C4943 vdd.n1900 gnd 0.009637f
C4944 vdd.n1901 gnd 0.00902f
C4945 vdd.n1903 gnd 0.011206f
C4946 vdd.n1905 gnd 0.00902f
C4947 vdd.n1906 gnd 0.011206f
C4948 vdd.n1907 gnd 0.00902f
C4949 vdd.n1909 gnd 0.011206f
C4950 vdd.n1910 gnd 0.00902f
C4951 vdd.n1911 gnd 0.011206f
C4952 vdd.n1912 gnd 0.011206f
C4953 vdd.n1913 gnd 0.011206f
C4954 vdd.n1914 gnd 0.011206f
C4955 vdd.n1915 gnd 0.011206f
C4956 vdd.n1916 gnd 0.00902f
C4957 vdd.n1918 gnd 0.011206f
C4958 vdd.n1919 gnd 0.011206f
C4959 vdd.n1920 gnd 0.011206f
C4960 vdd.n1921 gnd 0.011206f
C4961 vdd.n1922 gnd 0.011206f
C4962 vdd.n1923 gnd 0.00902f
C4963 vdd.n1925 gnd 0.011206f
C4964 vdd.n1926 gnd 0.011206f
C4965 vdd.n1927 gnd 0.011206f
C4966 vdd.n1928 gnd 0.011206f
C4967 vdd.n1929 gnd 0.007531f
C4968 vdd.t178 gnd 0.137864f
C4969 vdd.t177 gnd 0.147339f
C4970 vdd.t176 gnd 0.180049f
C4971 vdd.n1930 gnd 0.230797f
C4972 vdd.n1931 gnd 0.193911f
C4973 vdd.n1933 gnd 0.011206f
C4974 vdd.n1934 gnd 0.011206f
C4975 vdd.n1935 gnd 0.00902f
C4976 vdd.n1936 gnd 0.011206f
C4977 vdd.n1938 gnd 0.011206f
C4978 vdd.n1939 gnd 0.011206f
C4979 vdd.n1940 gnd 0.011206f
C4980 vdd.n1941 gnd 0.011206f
C4981 vdd.n1942 gnd 0.00902f
C4982 vdd.n1944 gnd 0.011206f
C4983 vdd.n1945 gnd 0.011206f
C4984 vdd.n1946 gnd 0.011206f
C4985 vdd.n1947 gnd 0.011206f
C4986 vdd.n1948 gnd 0.011206f
C4987 vdd.n1949 gnd 0.00902f
C4988 vdd.n1951 gnd 0.011206f
C4989 vdd.n1952 gnd 0.011206f
C4990 vdd.n1953 gnd 0.011206f
C4991 vdd.n1954 gnd 0.011206f
C4992 vdd.n1955 gnd 0.011206f
C4993 vdd.n1956 gnd 0.00902f
C4994 vdd.n1958 gnd 0.011206f
C4995 vdd.n1959 gnd 0.011206f
C4996 vdd.n1960 gnd 0.011206f
C4997 vdd.n1961 gnd 0.011206f
C4998 vdd.n1962 gnd 0.011206f
C4999 vdd.n1963 gnd 0.00902f
C5000 vdd.n1965 gnd 0.011206f
C5001 vdd.n1966 gnd 0.011206f
C5002 vdd.n1967 gnd 0.011206f
C5003 vdd.n1968 gnd 0.011206f
C5004 vdd.n1969 gnd 0.008929f
C5005 vdd.t165 gnd 0.137864f
C5006 vdd.t164 gnd 0.147339f
C5007 vdd.t163 gnd 0.180049f
C5008 vdd.n1970 gnd 0.230797f
C5009 vdd.n1971 gnd 0.193911f
C5010 vdd.n1973 gnd 0.011206f
C5011 vdd.n1974 gnd 0.011206f
C5012 vdd.n1975 gnd 0.00902f
C5013 vdd.n1976 gnd 0.011206f
C5014 vdd.n1978 gnd 0.011206f
C5015 vdd.n1979 gnd 0.011206f
C5016 vdd.n1980 gnd 0.011206f
C5017 vdd.n1981 gnd 0.011206f
C5018 vdd.n1982 gnd 0.00902f
C5019 vdd.n1984 gnd 0.011206f
C5020 vdd.n1985 gnd 0.011206f
C5021 vdd.n1986 gnd 0.011206f
C5022 vdd.n1987 gnd 0.011206f
C5023 vdd.n1988 gnd 0.011206f
C5024 vdd.n1989 gnd 0.00902f
C5025 vdd.n1991 gnd 0.011206f
C5026 vdd.n1992 gnd 0.011206f
C5027 vdd.n1993 gnd 0.011206f
C5028 vdd.n1994 gnd 0.011206f
C5029 vdd.n1995 gnd 0.011206f
C5030 vdd.n1996 gnd 0.011206f
C5031 vdd.n1997 gnd 0.00902f
C5032 vdd.n1999 gnd 0.011206f
C5033 vdd.n2001 gnd 0.011206f
C5034 vdd.n2002 gnd 0.00902f
C5035 vdd.n2003 gnd 0.00902f
C5036 vdd.n2004 gnd 0.011206f
C5037 vdd.n2006 gnd 0.011206f
C5038 vdd.n2007 gnd 0.00902f
C5039 vdd.n2008 gnd 0.00902f
C5040 vdd.n2009 gnd 0.011206f
C5041 vdd.n2011 gnd 0.011206f
C5042 vdd.n2012 gnd 0.011206f
C5043 vdd.n2013 gnd 0.00902f
C5044 vdd.n2014 gnd 0.00902f
C5045 vdd.n2015 gnd 0.00902f
C5046 vdd.n2016 gnd 0.011206f
C5047 vdd.n2018 gnd 0.011206f
C5048 vdd.n2019 gnd 0.011206f
C5049 vdd.n2020 gnd 0.00902f
C5050 vdd.n2021 gnd 0.00902f
C5051 vdd.n2022 gnd 0.00902f
C5052 vdd.n2023 gnd 0.011206f
C5053 vdd.n2025 gnd 0.011206f
C5054 vdd.n2026 gnd 0.011206f
C5055 vdd.n2027 gnd 0.00902f
C5056 vdd.n2028 gnd 0.00902f
C5057 vdd.n2029 gnd 0.00902f
C5058 vdd.n2030 gnd 0.011206f
C5059 vdd.n2032 gnd 0.011206f
C5060 vdd.n2033 gnd 0.011206f
C5061 vdd.n2034 gnd 0.00902f
C5062 vdd.n2035 gnd 0.011206f
C5063 vdd.n2036 gnd 0.011206f
C5064 vdd.n2037 gnd 0.011206f
C5065 vdd.n2038 gnd 0.0184f
C5066 vdd.n2039 gnd 0.006133f
C5067 vdd.n2040 gnd 0.00902f
C5068 vdd.n2041 gnd 0.011206f
C5069 vdd.n2043 gnd 0.011206f
C5070 vdd.n2044 gnd 0.011206f
C5071 vdd.n2045 gnd 0.00902f
C5072 vdd.n2046 gnd 0.00902f
C5073 vdd.n2047 gnd 0.00902f
C5074 vdd.n2048 gnd 0.011206f
C5075 vdd.n2050 gnd 0.011206f
C5076 vdd.n2051 gnd 0.011206f
C5077 vdd.n2052 gnd 0.00902f
C5078 vdd.n2053 gnd 0.00902f
C5079 vdd.n2054 gnd 0.00902f
C5080 vdd.n2055 gnd 0.011206f
C5081 vdd.n2057 gnd 0.011206f
C5082 vdd.n2058 gnd 0.011206f
C5083 vdd.n2059 gnd 0.00902f
C5084 vdd.n2060 gnd 0.00902f
C5085 vdd.n2061 gnd 0.00902f
C5086 vdd.n2062 gnd 0.011206f
C5087 vdd.n2064 gnd 0.011206f
C5088 vdd.n2065 gnd 0.011206f
C5089 vdd.n2066 gnd 0.00902f
C5090 vdd.n2067 gnd 0.00902f
C5091 vdd.n2068 gnd 0.00902f
C5092 vdd.n2069 gnd 0.011206f
C5093 vdd.n2071 gnd 0.011206f
C5094 vdd.n2072 gnd 0.011206f
C5095 vdd.n2073 gnd 0.00902f
C5096 vdd.n2074 gnd 0.011206f
C5097 vdd.n2075 gnd 0.011206f
C5098 vdd.n2076 gnd 0.011206f
C5099 vdd.n2077 gnd 0.0184f
C5100 vdd.n2078 gnd 0.007531f
C5101 vdd.n2079 gnd 0.00902f
C5102 vdd.n2080 gnd 0.011206f
C5103 vdd.n2082 gnd 0.011206f
C5104 vdd.n2083 gnd 0.011206f
C5105 vdd.n2084 gnd 0.00902f
C5106 vdd.n2085 gnd 0.00902f
C5107 vdd.n2086 gnd 0.00902f
C5108 vdd.n2087 gnd 0.011206f
C5109 vdd.n2089 gnd 0.011206f
C5110 vdd.n2090 gnd 0.011206f
C5111 vdd.n2091 gnd 0.00902f
C5112 vdd.n2092 gnd 0.00902f
C5113 vdd.n2093 gnd 0.00902f
C5114 vdd.n2094 gnd 0.011206f
C5115 vdd.n2096 gnd 0.011206f
C5116 vdd.n2097 gnd 0.011206f
C5117 vdd.n2099 gnd 0.011206f
C5118 vdd.n2100 gnd 0.00902f
C5119 vdd.n2101 gnd 0.007172f
C5120 vdd.n2102 gnd 0.00762f
C5121 vdd.n2103 gnd 0.00762f
C5122 vdd.n2104 gnd 0.00762f
C5123 vdd.n2105 gnd 0.00762f
C5124 vdd.n2106 gnd 0.00762f
C5125 vdd.n2107 gnd 0.00762f
C5126 vdd.n2108 gnd 0.00762f
C5127 vdd.n2109 gnd 0.00762f
C5128 vdd.n2111 gnd 0.00762f
C5129 vdd.n2112 gnd 0.00762f
C5130 vdd.n2113 gnd 0.00762f
C5131 vdd.n2114 gnd 0.00762f
C5132 vdd.n2115 gnd 0.00762f
C5133 vdd.n2117 gnd 0.00762f
C5134 vdd.n2119 gnd 0.00762f
C5135 vdd.n2120 gnd 0.00762f
C5136 vdd.n2121 gnd 0.00762f
C5137 vdd.n2122 gnd 0.00762f
C5138 vdd.n2123 gnd 0.00762f
C5139 vdd.n2125 gnd 0.00762f
C5140 vdd.n2127 gnd 0.00762f
C5141 vdd.n2128 gnd 0.00762f
C5142 vdd.n2129 gnd 0.00762f
C5143 vdd.n2130 gnd 0.00762f
C5144 vdd.n2131 gnd 0.00762f
C5145 vdd.n2133 gnd 0.00762f
C5146 vdd.n2135 gnd 0.00762f
C5147 vdd.n2136 gnd 0.00762f
C5148 vdd.n2137 gnd 0.00762f
C5149 vdd.n2138 gnd 0.00762f
C5150 vdd.n2139 gnd 0.00762f
C5151 vdd.n2141 gnd 0.00762f
C5152 vdd.n2142 gnd 0.00762f
C5153 vdd.n2143 gnd 0.00762f
C5154 vdd.n2144 gnd 0.00762f
C5155 vdd.n2145 gnd 0.00762f
C5156 vdd.n2146 gnd 0.00762f
C5157 vdd.n2147 gnd 0.00762f
C5158 vdd.n2148 gnd 0.00762f
C5159 vdd.n2149 gnd 0.005547f
C5160 vdd.n2150 gnd 0.00762f
C5161 vdd.t218 gnd 0.307928f
C5162 vdd.t219 gnd 0.315203f
C5163 vdd.t217 gnd 0.201027f
C5164 vdd.n2151 gnd 0.108644f
C5165 vdd.n2152 gnd 0.061626f
C5166 vdd.n2153 gnd 0.01089f
C5167 vdd.n2154 gnd 0.00762f
C5168 vdd.n2155 gnd 0.00762f
C5169 vdd.n2156 gnd 0.463809f
C5170 vdd.n2157 gnd 0.00762f
C5171 vdd.n2158 gnd 0.00762f
C5172 vdd.n2159 gnd 0.00762f
C5173 vdd.n2160 gnd 0.00762f
C5174 vdd.n2161 gnd 0.00762f
C5175 vdd.n2162 gnd 0.00762f
C5176 vdd.n2163 gnd 0.00762f
C5177 vdd.n2164 gnd 0.00762f
C5178 vdd.n2165 gnd 0.00762f
C5179 vdd.n2166 gnd 0.00762f
C5180 vdd.n2167 gnd 0.00762f
C5181 vdd.n2168 gnd 0.00762f
C5182 vdd.n2169 gnd 0.00762f
C5183 vdd.n2170 gnd 0.00762f
C5184 vdd.n2171 gnd 0.00762f
C5185 vdd.n2172 gnd 0.00762f
C5186 vdd.n2173 gnd 0.00762f
C5187 vdd.n2174 gnd 0.00762f
C5188 vdd.n2175 gnd 0.00762f
C5189 vdd.n2176 gnd 0.00762f
C5190 vdd.t196 gnd 0.307928f
C5191 vdd.t197 gnd 0.315203f
C5192 vdd.t194 gnd 0.201027f
C5193 vdd.n2177 gnd 0.108644f
C5194 vdd.n2178 gnd 0.061626f
C5195 vdd.n2179 gnd 0.00762f
C5196 vdd.n2180 gnd 0.00762f
C5197 vdd.n2181 gnd 0.00762f
C5198 vdd.n2182 gnd 0.00762f
C5199 vdd.n2183 gnd 0.00762f
C5200 vdd.n2184 gnd 0.00762f
C5201 vdd.n2186 gnd 0.00762f
C5202 vdd.n2187 gnd 0.00762f
C5203 vdd.n2188 gnd 0.00762f
C5204 vdd.n2189 gnd 0.00762f
C5205 vdd.n2191 gnd 0.00762f
C5206 vdd.n2193 gnd 0.00762f
C5207 vdd.n2194 gnd 0.00762f
C5208 vdd.n2195 gnd 0.00762f
C5209 vdd.n2196 gnd 0.00762f
C5210 vdd.n2197 gnd 0.00762f
C5211 vdd.n2199 gnd 0.00762f
C5212 vdd.n2201 gnd 0.00762f
C5213 vdd.n2202 gnd 0.00762f
C5214 vdd.n2203 gnd 0.00762f
C5215 vdd.n2204 gnd 0.00762f
C5216 vdd.n2205 gnd 0.00762f
C5217 vdd.n2207 gnd 0.00762f
C5218 vdd.n2209 gnd 0.00762f
C5219 vdd.n2210 gnd 0.00762f
C5220 vdd.n2211 gnd 0.005547f
C5221 vdd.n2212 gnd 0.01089f
C5222 vdd.n2213 gnd 0.005883f
C5223 vdd.n2214 gnd 0.00762f
C5224 vdd.n2216 gnd 0.00762f
C5225 vdd.n2217 gnd 0.018081f
C5226 vdd.n2218 gnd 0.018081f
C5227 vdd.n2219 gnd 0.016882f
C5228 vdd.n2220 gnd 0.00762f
C5229 vdd.n2221 gnd 0.00762f
C5230 vdd.n2222 gnd 0.00762f
C5231 vdd.n2223 gnd 0.00762f
C5232 vdd.n2224 gnd 0.00762f
C5233 vdd.n2225 gnd 0.00762f
C5234 vdd.n2226 gnd 0.00762f
C5235 vdd.n2227 gnd 0.00762f
C5236 vdd.n2228 gnd 0.00762f
C5237 vdd.n2229 gnd 0.00762f
C5238 vdd.n2230 gnd 0.00762f
C5239 vdd.n2231 gnd 0.00762f
C5240 vdd.n2232 gnd 0.00762f
C5241 vdd.n2233 gnd 0.00762f
C5242 vdd.n2234 gnd 0.00762f
C5243 vdd.n2235 gnd 0.00762f
C5244 vdd.n2236 gnd 0.00762f
C5245 vdd.n2237 gnd 0.00762f
C5246 vdd.n2238 gnd 0.00762f
C5247 vdd.n2239 gnd 0.00762f
C5248 vdd.n2240 gnd 0.00762f
C5249 vdd.n2241 gnd 0.00762f
C5250 vdd.n2242 gnd 0.00762f
C5251 vdd.n2243 gnd 0.00762f
C5252 vdd.n2244 gnd 0.00762f
C5253 vdd.n2245 gnd 0.00762f
C5254 vdd.n2246 gnd 0.00762f
C5255 vdd.n2247 gnd 0.00762f
C5256 vdd.n2248 gnd 0.00762f
C5257 vdd.n2249 gnd 0.00762f
C5258 vdd.n2250 gnd 0.00762f
C5259 vdd.n2251 gnd 0.00762f
C5260 vdd.n2252 gnd 0.00762f
C5261 vdd.n2253 gnd 0.00762f
C5262 vdd.n2254 gnd 0.00762f
C5263 vdd.n2255 gnd 0.00762f
C5264 vdd.n2256 gnd 0.00762f
C5265 vdd.n2257 gnd 0.246219f
C5266 vdd.n2258 gnd 0.00762f
C5267 vdd.n2259 gnd 0.00762f
C5268 vdd.n2260 gnd 0.00762f
C5269 vdd.n2261 gnd 0.00762f
C5270 vdd.n2262 gnd 0.00762f
C5271 vdd.n2263 gnd 0.00762f
C5272 vdd.n2264 gnd 0.00762f
C5273 vdd.n2265 gnd 0.00762f
C5274 vdd.n2266 gnd 0.00762f
C5275 vdd.n2267 gnd 0.00762f
C5276 vdd.n2268 gnd 0.00762f
C5277 vdd.n2269 gnd 0.00762f
C5278 vdd.n2270 gnd 0.00762f
C5279 vdd.n2271 gnd 0.00762f
C5280 vdd.n2272 gnd 0.00762f
C5281 vdd.n2273 gnd 0.00762f
C5282 vdd.n2274 gnd 0.00762f
C5283 vdd.n2275 gnd 0.00762f
C5284 vdd.n2276 gnd 0.00762f
C5285 vdd.n2277 gnd 0.00762f
C5286 vdd.n2278 gnd 0.016882f
C5287 vdd.n2280 gnd 0.018081f
C5288 vdd.n2281 gnd 0.018081f
C5289 vdd.n2282 gnd 0.00762f
C5290 vdd.n2283 gnd 0.005883f
C5291 vdd.n2284 gnd 0.00762f
C5292 vdd.n2286 gnd 0.00762f
C5293 vdd.n2288 gnd 0.00762f
C5294 vdd.n2289 gnd 0.00762f
C5295 vdd.n2290 gnd 0.00762f
C5296 vdd.n2291 gnd 0.00762f
C5297 vdd.n2292 gnd 0.00762f
C5298 vdd.n2294 gnd 0.00762f
C5299 vdd.n2296 gnd 0.00762f
C5300 vdd.n2297 gnd 0.00762f
C5301 vdd.n2298 gnd 0.00762f
C5302 vdd.n2299 gnd 0.00762f
C5303 vdd.n2300 gnd 0.00762f
C5304 vdd.n2302 gnd 0.00762f
C5305 vdd.n2304 gnd 0.00762f
C5306 vdd.n2305 gnd 0.00762f
C5307 vdd.n2306 gnd 0.00762f
C5308 vdd.n2307 gnd 0.00762f
C5309 vdd.n2308 gnd 0.00762f
C5310 vdd.n2310 gnd 0.00762f
C5311 vdd.n2312 gnd 0.00762f
C5312 vdd.n2313 gnd 0.00762f
C5313 vdd.n2314 gnd 0.022729f
C5314 vdd.n2315 gnd 0.673791f
C5315 vdd.n2317 gnd 0.00902f
C5316 vdd.n2318 gnd 0.00902f
C5317 vdd.n2319 gnd 0.011206f
C5318 vdd.n2321 gnd 0.011206f
C5319 vdd.n2322 gnd 0.011206f
C5320 vdd.n2323 gnd 0.00902f
C5321 vdd.n2324 gnd 0.007486f
C5322 vdd.n2325 gnd 0.027689f
C5323 vdd.n2326 gnd 0.027108f
C5324 vdd.n2327 gnd 0.007486f
C5325 vdd.n2328 gnd 0.027108f
C5326 vdd.n2329 gnd 1.57466f
C5327 vdd.n2330 gnd 0.027108f
C5328 vdd.n2331 gnd 0.027689f
C5329 vdd.n2332 gnd 0.004284f
C5330 vdd.t154 gnd 0.137864f
C5331 vdd.t153 gnd 0.147339f
C5332 vdd.t151 gnd 0.180049f
C5333 vdd.n2333 gnd 0.230797f
C5334 vdd.n2334 gnd 0.193911f
C5335 vdd.n2335 gnd 0.01389f
C5336 vdd.n2336 gnd 0.004735f
C5337 vdd.n2337 gnd 0.009637f
C5338 vdd.n2338 gnd 0.673791f
C5339 vdd.n2339 gnd 0.022729f
C5340 vdd.n2340 gnd 0.00762f
C5341 vdd.n2341 gnd 0.00762f
C5342 vdd.n2342 gnd 0.00762f
C5343 vdd.n2344 gnd 0.00762f
C5344 vdd.n2346 gnd 0.00762f
C5345 vdd.n2347 gnd 0.00762f
C5346 vdd.n2348 gnd 0.00762f
C5347 vdd.n2349 gnd 0.00762f
C5348 vdd.n2350 gnd 0.00762f
C5349 vdd.n2352 gnd 0.00762f
C5350 vdd.n2354 gnd 0.00762f
C5351 vdd.n2355 gnd 0.00762f
C5352 vdd.n2356 gnd 0.00762f
C5353 vdd.n2357 gnd 0.00762f
C5354 vdd.n2358 gnd 0.00762f
C5355 vdd.n2360 gnd 0.00762f
C5356 vdd.n2362 gnd 0.00762f
C5357 vdd.n2363 gnd 0.00762f
C5358 vdd.n2364 gnd 0.00762f
C5359 vdd.n2365 gnd 0.00762f
C5360 vdd.n2366 gnd 0.00762f
C5361 vdd.n2368 gnd 0.00762f
C5362 vdd.n2370 gnd 0.00762f
C5363 vdd.n2371 gnd 0.00762f
C5364 vdd.n2372 gnd 0.018081f
C5365 vdd.n2373 gnd 0.016882f
C5366 vdd.n2374 gnd 0.016882f
C5367 vdd.n2375 gnd 1.1223f
C5368 vdd.n2376 gnd 0.016882f
C5369 vdd.n2377 gnd 0.016882f
C5370 vdd.n2378 gnd 0.00762f
C5371 vdd.n2379 gnd 0.00762f
C5372 vdd.n2380 gnd 0.00762f
C5373 vdd.n2381 gnd 0.486713f
C5374 vdd.n2382 gnd 0.00762f
C5375 vdd.n2383 gnd 0.00762f
C5376 vdd.n2384 gnd 0.00762f
C5377 vdd.n2385 gnd 0.00762f
C5378 vdd.n2386 gnd 0.00762f
C5379 vdd.n2387 gnd 0.77874f
C5380 vdd.n2388 gnd 0.00762f
C5381 vdd.n2389 gnd 0.00762f
C5382 vdd.n2390 gnd 0.00762f
C5383 vdd.n2391 gnd 0.00762f
C5384 vdd.n2392 gnd 0.00762f
C5385 vdd.n2393 gnd 0.77874f
C5386 vdd.n2394 gnd 0.00762f
C5387 vdd.n2395 gnd 0.00762f
C5388 vdd.n2396 gnd 0.006724f
C5389 vdd.n2397 gnd 0.022075f
C5390 vdd.n2398 gnd 0.004707f
C5391 vdd.n2399 gnd 0.00762f
C5392 vdd.n2400 gnd 0.429452f
C5393 vdd.n2401 gnd 0.00762f
C5394 vdd.n2402 gnd 0.00762f
C5395 vdd.n2403 gnd 0.00762f
C5396 vdd.n2404 gnd 0.00762f
C5397 vdd.n2405 gnd 0.00762f
C5398 vdd.n2406 gnd 0.521069f
C5399 vdd.n2407 gnd 0.00762f
C5400 vdd.n2408 gnd 0.00762f
C5401 vdd.n2409 gnd 0.00762f
C5402 vdd.n2410 gnd 0.00762f
C5403 vdd.n2411 gnd 0.00762f
C5404 vdd.n2412 gnd 0.69285f
C5405 vdd.n2413 gnd 0.00762f
C5406 vdd.n2414 gnd 0.00762f
C5407 vdd.n2415 gnd 0.00762f
C5408 vdd.n2416 gnd 0.00762f
C5409 vdd.n2417 gnd 0.00762f
C5410 vdd.n2418 gnd 0.618412f
C5411 vdd.n2419 gnd 0.00762f
C5412 vdd.n2420 gnd 0.00762f
C5413 vdd.n2421 gnd 0.00762f
C5414 vdd.n2422 gnd 0.00762f
C5415 vdd.n2423 gnd 0.00762f
C5416 vdd.n2424 gnd 0.446631f
C5417 vdd.n2425 gnd 0.00762f
C5418 vdd.n2426 gnd 0.00762f
C5419 vdd.n2427 gnd 0.00762f
C5420 vdd.n2428 gnd 0.00762f
C5421 vdd.n2429 gnd 0.00762f
C5422 vdd.n2430 gnd 0.246219f
C5423 vdd.n2431 gnd 0.00762f
C5424 vdd.n2432 gnd 0.00762f
C5425 vdd.n2433 gnd 0.00762f
C5426 vdd.n2434 gnd 0.00762f
C5427 vdd.n2435 gnd 0.00762f
C5428 vdd.n2436 gnd 0.429452f
C5429 vdd.n2437 gnd 0.00762f
C5430 vdd.n2438 gnd 0.00762f
C5431 vdd.n2439 gnd 0.00762f
C5432 vdd.n2440 gnd 0.00762f
C5433 vdd.n2441 gnd 0.00762f
C5434 vdd.n2442 gnd 0.77874f
C5435 vdd.n2443 gnd 0.00762f
C5436 vdd.n2444 gnd 0.00762f
C5437 vdd.n2445 gnd 0.00762f
C5438 vdd.n2446 gnd 0.00762f
C5439 vdd.n2447 gnd 0.00762f
C5440 vdd.n2448 gnd 0.00762f
C5441 vdd.n2449 gnd 0.00762f
C5442 vdd.n2450 gnd 0.606959f
C5443 vdd.n2451 gnd 0.00762f
C5444 vdd.n2452 gnd 0.00762f
C5445 vdd.n2453 gnd 0.00762f
C5446 vdd.n2454 gnd 0.00762f
C5447 vdd.n2455 gnd 0.00762f
C5448 vdd.n2456 gnd 0.00762f
C5449 vdd.n2457 gnd 0.486713f
C5450 vdd.n2458 gnd 0.00762f
C5451 vdd.n2459 gnd 0.00762f
C5452 vdd.n2460 gnd 0.00762f
C5453 vdd.n2461 gnd 0.01781f
C5454 vdd.n2462 gnd 0.017153f
C5455 vdd.n2463 gnd 0.00762f
C5456 vdd.n2464 gnd 0.00762f
C5457 vdd.n2465 gnd 0.005883f
C5458 vdd.n2466 gnd 0.00762f
C5459 vdd.n2467 gnd 0.00762f
C5460 vdd.n2468 gnd 0.005547f
C5461 vdd.n2469 gnd 0.00762f
C5462 vdd.n2470 gnd 0.00762f
C5463 vdd.n2471 gnd 0.00762f
C5464 vdd.n2472 gnd 0.00762f
C5465 vdd.n2473 gnd 0.00762f
C5466 vdd.n2474 gnd 0.00762f
C5467 vdd.n2475 gnd 0.00762f
C5468 vdd.n2476 gnd 0.00762f
C5469 vdd.n2477 gnd 0.00762f
C5470 vdd.n2478 gnd 0.00762f
C5471 vdd.n2479 gnd 0.00762f
C5472 vdd.n2480 gnd 0.00762f
C5473 vdd.n2481 gnd 0.00762f
C5474 vdd.n2482 gnd 0.00762f
C5475 vdd.n2483 gnd 0.00762f
C5476 vdd.n2484 gnd 0.00762f
C5477 vdd.n2485 gnd 0.00762f
C5478 vdd.n2486 gnd 0.00762f
C5479 vdd.n2487 gnd 0.00762f
C5480 vdd.n2488 gnd 0.00762f
C5481 vdd.n2489 gnd 0.00762f
C5482 vdd.n2490 gnd 0.00762f
C5483 vdd.n2491 gnd 0.00762f
C5484 vdd.n2492 gnd 0.00762f
C5485 vdd.n2493 gnd 0.00762f
C5486 vdd.n2494 gnd 0.00762f
C5487 vdd.n2495 gnd 0.00762f
C5488 vdd.n2496 gnd 0.00762f
C5489 vdd.n2497 gnd 0.00762f
C5490 vdd.n2498 gnd 0.00762f
C5491 vdd.n2499 gnd 0.00762f
C5492 vdd.n2500 gnd 0.00762f
C5493 vdd.n2501 gnd 0.00762f
C5494 vdd.n2502 gnd 0.00762f
C5495 vdd.n2503 gnd 0.00762f
C5496 vdd.n2504 gnd 0.00762f
C5497 vdd.n2505 gnd 0.00762f
C5498 vdd.n2506 gnd 0.00762f
C5499 vdd.n2507 gnd 0.00762f
C5500 vdd.n2508 gnd 0.00762f
C5501 vdd.n2509 gnd 0.00762f
C5502 vdd.n2510 gnd 0.00762f
C5503 vdd.n2511 gnd 0.00762f
C5504 vdd.n2512 gnd 0.00762f
C5505 vdd.n2513 gnd 0.00762f
C5506 vdd.n2514 gnd 0.00762f
C5507 vdd.n2515 gnd 0.00762f
C5508 vdd.n2516 gnd 0.00762f
C5509 vdd.n2517 gnd 0.00762f
C5510 vdd.n2518 gnd 0.00762f
C5511 vdd.n2519 gnd 0.00762f
C5512 vdd.n2520 gnd 0.00762f
C5513 vdd.n2521 gnd 0.00762f
C5514 vdd.n2522 gnd 0.00762f
C5515 vdd.n2523 gnd 0.00762f
C5516 vdd.n2524 gnd 0.00762f
C5517 vdd.n2525 gnd 0.00762f
C5518 vdd.n2526 gnd 0.00762f
C5519 vdd.n2527 gnd 0.00762f
C5520 vdd.n2528 gnd 0.00762f
C5521 vdd.n2529 gnd 0.018081f
C5522 vdd.n2530 gnd 0.016882f
C5523 vdd.n2531 gnd 0.016882f
C5524 vdd.n2532 gnd 0.950521f
C5525 vdd.n2533 gnd 0.016882f
C5526 vdd.n2534 gnd 0.018081f
C5527 vdd.n2535 gnd 0.017153f
C5528 vdd.n2536 gnd 0.00762f
C5529 vdd.n2537 gnd 0.00762f
C5530 vdd.n2538 gnd 0.00762f
C5531 vdd.n2539 gnd 0.005883f
C5532 vdd.n2540 gnd 0.01089f
C5533 vdd.n2541 gnd 0.005547f
C5534 vdd.n2542 gnd 0.00762f
C5535 vdd.n2543 gnd 0.00762f
C5536 vdd.n2544 gnd 0.00762f
C5537 vdd.n2545 gnd 0.00762f
C5538 vdd.n2546 gnd 0.00762f
C5539 vdd.n2547 gnd 0.00762f
C5540 vdd.n2548 gnd 0.00762f
C5541 vdd.n2549 gnd 0.00762f
C5542 vdd.n2550 gnd 0.00762f
C5543 vdd.n2551 gnd 0.00762f
C5544 vdd.n2552 gnd 0.00762f
C5545 vdd.n2553 gnd 0.00762f
C5546 vdd.n2554 gnd 0.00762f
C5547 vdd.n2555 gnd 0.00762f
C5548 vdd.n2556 gnd 0.00762f
C5549 vdd.n2557 gnd 0.00762f
C5550 vdd.n2558 gnd 0.00762f
C5551 vdd.n2559 gnd 0.00762f
C5552 vdd.n2560 gnd 0.00762f
C5553 vdd.n2561 gnd 0.00762f
C5554 vdd.n2562 gnd 0.00762f
C5555 vdd.n2563 gnd 0.00762f
C5556 vdd.n2564 gnd 0.00762f
C5557 vdd.n2565 gnd 0.00762f
C5558 vdd.n2566 gnd 0.00762f
C5559 vdd.n2567 gnd 0.00762f
C5560 vdd.n2568 gnd 0.00762f
C5561 vdd.n2569 gnd 0.00762f
C5562 vdd.n2570 gnd 0.00762f
C5563 vdd.n2571 gnd 0.00762f
C5564 vdd.n2572 gnd 0.00762f
C5565 vdd.n2573 gnd 0.00762f
C5566 vdd.n2574 gnd 0.00762f
C5567 vdd.n2575 gnd 0.00762f
C5568 vdd.n2576 gnd 0.00762f
C5569 vdd.n2577 gnd 0.00762f
C5570 vdd.n2578 gnd 0.00762f
C5571 vdd.n2579 gnd 0.00762f
C5572 vdd.n2580 gnd 0.00762f
C5573 vdd.n2581 gnd 0.00762f
C5574 vdd.n2582 gnd 0.00762f
C5575 vdd.n2583 gnd 0.00762f
C5576 vdd.n2584 gnd 0.00762f
C5577 vdd.n2585 gnd 0.00762f
C5578 vdd.n2586 gnd 0.00762f
C5579 vdd.n2587 gnd 0.00762f
C5580 vdd.n2588 gnd 0.00762f
C5581 vdd.n2589 gnd 0.00762f
C5582 vdd.n2590 gnd 0.00762f
C5583 vdd.n2591 gnd 0.00762f
C5584 vdd.n2592 gnd 0.00762f
C5585 vdd.n2593 gnd 0.00762f
C5586 vdd.n2594 gnd 0.00762f
C5587 vdd.n2595 gnd 0.00762f
C5588 vdd.n2596 gnd 0.00762f
C5589 vdd.n2597 gnd 0.00762f
C5590 vdd.n2598 gnd 0.00762f
C5591 vdd.n2599 gnd 0.00762f
C5592 vdd.n2600 gnd 0.00762f
C5593 vdd.n2601 gnd 0.00762f
C5594 vdd.n2602 gnd 0.018081f
C5595 vdd.n2603 gnd 0.018081f
C5596 vdd.n2604 gnd 0.950521f
C5597 vdd.t253 gnd 3.37836f
C5598 vdd.t240 gnd 3.37836f
C5599 vdd.n2637 gnd 0.018081f
C5600 vdd.n2638 gnd 0.00762f
C5601 vdd.t189 gnd 0.307928f
C5602 vdd.t190 gnd 0.315203f
C5603 vdd.t187 gnd 0.201027f
C5604 vdd.n2639 gnd 0.108644f
C5605 vdd.n2640 gnd 0.061626f
C5606 vdd.n2641 gnd 0.00762f
C5607 vdd.t203 gnd 0.307928f
C5608 vdd.t204 gnd 0.315203f
C5609 vdd.t202 gnd 0.201027f
C5610 vdd.n2642 gnd 0.108644f
C5611 vdd.n2643 gnd 0.061626f
C5612 vdd.n2644 gnd 0.01089f
C5613 vdd.n2645 gnd 0.00762f
C5614 vdd.n2646 gnd 0.00762f
C5615 vdd.n2647 gnd 0.00762f
C5616 vdd.n2648 gnd 0.00762f
C5617 vdd.n2649 gnd 0.00762f
C5618 vdd.n2650 gnd 0.00762f
C5619 vdd.n2651 gnd 0.00762f
C5620 vdd.n2652 gnd 0.00762f
C5621 vdd.n2653 gnd 0.00762f
C5622 vdd.n2654 gnd 0.00762f
C5623 vdd.n2655 gnd 0.00762f
C5624 vdd.n2656 gnd 0.00762f
C5625 vdd.n2657 gnd 0.00762f
C5626 vdd.n2658 gnd 0.00762f
C5627 vdd.n2659 gnd 0.00762f
C5628 vdd.n2660 gnd 0.00762f
C5629 vdd.n2661 gnd 0.00762f
C5630 vdd.n2662 gnd 0.00762f
C5631 vdd.n2663 gnd 0.00762f
C5632 vdd.n2664 gnd 0.00762f
C5633 vdd.n2665 gnd 0.00762f
C5634 vdd.n2666 gnd 0.00762f
C5635 vdd.n2667 gnd 0.00762f
C5636 vdd.n2668 gnd 0.00762f
C5637 vdd.n2669 gnd 0.00762f
C5638 vdd.n2670 gnd 0.00762f
C5639 vdd.n2671 gnd 0.00762f
C5640 vdd.n2672 gnd 0.00762f
C5641 vdd.n2673 gnd 0.00762f
C5642 vdd.n2674 gnd 0.00762f
C5643 vdd.n2675 gnd 0.00762f
C5644 vdd.n2676 gnd 0.00762f
C5645 vdd.n2677 gnd 0.00762f
C5646 vdd.n2678 gnd 0.00762f
C5647 vdd.n2679 gnd 0.00762f
C5648 vdd.n2680 gnd 0.00762f
C5649 vdd.n2681 gnd 0.00762f
C5650 vdd.n2682 gnd 0.00762f
C5651 vdd.n2683 gnd 0.00762f
C5652 vdd.n2684 gnd 0.00762f
C5653 vdd.n2685 gnd 0.00762f
C5654 vdd.n2686 gnd 0.00762f
C5655 vdd.n2687 gnd 0.00762f
C5656 vdd.n2688 gnd 0.00762f
C5657 vdd.n2689 gnd 0.00762f
C5658 vdd.n2690 gnd 0.00762f
C5659 vdd.n2691 gnd 0.00762f
C5660 vdd.n2692 gnd 0.00762f
C5661 vdd.n2693 gnd 0.00762f
C5662 vdd.n2694 gnd 0.00762f
C5663 vdd.n2695 gnd 0.00762f
C5664 vdd.n2696 gnd 0.00762f
C5665 vdd.n2697 gnd 0.00762f
C5666 vdd.n2698 gnd 0.00762f
C5667 vdd.n2699 gnd 0.00762f
C5668 vdd.n2700 gnd 0.00762f
C5669 vdd.n2701 gnd 0.005547f
C5670 vdd.n2702 gnd 0.00762f
C5671 vdd.n2703 gnd 0.00762f
C5672 vdd.n2704 gnd 0.005883f
C5673 vdd.n2705 gnd 0.00762f
C5674 vdd.n2706 gnd 0.00762f
C5675 vdd.n2707 gnd 0.018081f
C5676 vdd.n2708 gnd 0.016882f
C5677 vdd.n2709 gnd 0.00762f
C5678 vdd.n2710 gnd 0.00762f
C5679 vdd.n2711 gnd 0.00762f
C5680 vdd.n2712 gnd 0.00762f
C5681 vdd.n2713 gnd 0.00762f
C5682 vdd.n2714 gnd 0.00762f
C5683 vdd.n2715 gnd 0.00762f
C5684 vdd.n2716 gnd 0.00762f
C5685 vdd.n2717 gnd 0.00762f
C5686 vdd.n2718 gnd 0.00762f
C5687 vdd.n2719 gnd 0.00762f
C5688 vdd.n2720 gnd 0.00762f
C5689 vdd.n2721 gnd 0.00762f
C5690 vdd.n2722 gnd 0.00762f
C5691 vdd.n2723 gnd 0.00762f
C5692 vdd.n2724 gnd 0.00762f
C5693 vdd.n2725 gnd 0.00762f
C5694 vdd.n2726 gnd 0.00762f
C5695 vdd.n2727 gnd 0.00762f
C5696 vdd.n2728 gnd 0.00762f
C5697 vdd.n2729 gnd 0.00762f
C5698 vdd.n2730 gnd 0.00762f
C5699 vdd.n2731 gnd 0.00762f
C5700 vdd.n2732 gnd 0.00762f
C5701 vdd.n2733 gnd 0.00762f
C5702 vdd.n2734 gnd 0.00762f
C5703 vdd.n2735 gnd 0.00762f
C5704 vdd.n2736 gnd 0.00762f
C5705 vdd.n2737 gnd 0.00762f
C5706 vdd.n2738 gnd 0.00762f
C5707 vdd.n2739 gnd 0.00762f
C5708 vdd.n2740 gnd 0.00762f
C5709 vdd.n2741 gnd 0.00762f
C5710 vdd.n2742 gnd 0.00762f
C5711 vdd.n2743 gnd 0.00762f
C5712 vdd.n2744 gnd 0.00762f
C5713 vdd.n2745 gnd 0.00762f
C5714 vdd.n2746 gnd 0.00762f
C5715 vdd.n2747 gnd 0.00762f
C5716 vdd.n2748 gnd 0.00762f
C5717 vdd.n2749 gnd 0.00762f
C5718 vdd.n2750 gnd 0.00762f
C5719 vdd.n2751 gnd 0.00762f
C5720 vdd.n2752 gnd 0.00762f
C5721 vdd.n2753 gnd 0.00762f
C5722 vdd.n2754 gnd 0.00762f
C5723 vdd.n2755 gnd 0.00762f
C5724 vdd.n2756 gnd 0.00762f
C5725 vdd.n2757 gnd 0.00762f
C5726 vdd.n2758 gnd 0.00762f
C5727 vdd.n2759 gnd 0.00762f
C5728 vdd.n2760 gnd 0.246219f
C5729 vdd.n2761 gnd 0.00762f
C5730 vdd.n2762 gnd 0.00762f
C5731 vdd.n2763 gnd 0.00762f
C5732 vdd.n2764 gnd 0.00762f
C5733 vdd.n2765 gnd 0.00762f
C5734 vdd.n2766 gnd 0.00762f
C5735 vdd.n2767 gnd 0.00762f
C5736 vdd.n2768 gnd 0.00762f
C5737 vdd.n2769 gnd 0.00762f
C5738 vdd.n2770 gnd 0.00762f
C5739 vdd.n2771 gnd 0.00762f
C5740 vdd.n2772 gnd 0.00762f
C5741 vdd.n2773 gnd 0.00762f
C5742 vdd.n2774 gnd 0.00762f
C5743 vdd.n2775 gnd 0.00762f
C5744 vdd.n2776 gnd 0.00762f
C5745 vdd.n2777 gnd 0.00762f
C5746 vdd.n2778 gnd 0.00762f
C5747 vdd.n2779 gnd 0.00762f
C5748 vdd.n2780 gnd 0.00762f
C5749 vdd.n2781 gnd 0.463809f
C5750 vdd.n2782 gnd 0.00762f
C5751 vdd.n2783 gnd 0.00762f
C5752 vdd.n2784 gnd 0.00762f
C5753 vdd.n2785 gnd 0.00762f
C5754 vdd.n2786 gnd 0.00762f
C5755 vdd.n2787 gnd 0.016882f
C5756 vdd.n2788 gnd 0.018081f
C5757 vdd.n2789 gnd 0.018081f
C5758 vdd.n2790 gnd 0.00762f
C5759 vdd.n2791 gnd 0.00762f
C5760 vdd.n2792 gnd 0.00762f
C5761 vdd.n2793 gnd 0.005883f
C5762 vdd.n2794 gnd 0.01089f
C5763 vdd.n2795 gnd 0.005547f
C5764 vdd.n2796 gnd 0.00762f
C5765 vdd.n2797 gnd 0.00762f
C5766 vdd.n2798 gnd 0.00762f
C5767 vdd.n2799 gnd 0.00762f
C5768 vdd.n2800 gnd 0.00762f
C5769 vdd.n2801 gnd 0.00762f
C5770 vdd.n2802 gnd 0.00762f
C5771 vdd.n2803 gnd 0.00762f
C5772 vdd.n2804 gnd 0.00762f
C5773 vdd.n2805 gnd 0.00762f
C5774 vdd.n2806 gnd 0.00762f
C5775 vdd.n2807 gnd 0.00762f
C5776 vdd.n2808 gnd 0.00762f
C5777 vdd.n2809 gnd 0.00762f
C5778 vdd.n2810 gnd 0.00762f
C5779 vdd.n2811 gnd 0.00762f
C5780 vdd.n2812 gnd 0.00762f
C5781 vdd.n2813 gnd 0.00762f
C5782 vdd.n2814 gnd 0.00762f
C5783 vdd.n2815 gnd 0.00762f
C5784 vdd.n2816 gnd 0.00762f
C5785 vdd.n2817 gnd 0.00762f
C5786 vdd.n2818 gnd 0.00762f
C5787 vdd.n2819 gnd 0.00762f
C5788 vdd.n2820 gnd 0.00762f
C5789 vdd.n2821 gnd 0.00762f
C5790 vdd.n2822 gnd 0.00762f
C5791 vdd.n2823 gnd 0.00762f
C5792 vdd.n2824 gnd 0.00762f
C5793 vdd.n2825 gnd 0.00762f
C5794 vdd.n2826 gnd 0.00762f
C5795 vdd.n2827 gnd 0.00762f
C5796 vdd.n2828 gnd 0.00762f
C5797 vdd.n2829 gnd 0.00762f
C5798 vdd.n2830 gnd 0.00762f
C5799 vdd.n2831 gnd 0.00762f
C5800 vdd.n2832 gnd 0.00762f
C5801 vdd.n2833 gnd 0.00762f
C5802 vdd.n2834 gnd 0.00762f
C5803 vdd.n2835 gnd 0.00762f
C5804 vdd.n2836 gnd 0.00762f
C5805 vdd.n2837 gnd 0.00762f
C5806 vdd.n2838 gnd 0.00762f
C5807 vdd.n2839 gnd 0.00762f
C5808 vdd.n2840 gnd 0.00762f
C5809 vdd.n2841 gnd 0.00762f
C5810 vdd.n2842 gnd 0.00762f
C5811 vdd.n2843 gnd 0.00762f
C5812 vdd.n2844 gnd 0.00762f
C5813 vdd.n2845 gnd 0.00762f
C5814 vdd.n2846 gnd 0.00762f
C5815 vdd.n2847 gnd 0.00762f
C5816 vdd.n2848 gnd 0.00762f
C5817 vdd.n2849 gnd 0.00762f
C5818 vdd.n2850 gnd 0.00762f
C5819 vdd.n2851 gnd 0.00762f
C5820 vdd.n2852 gnd 0.00762f
C5821 vdd.n2853 gnd 0.00762f
C5822 vdd.n2854 gnd 0.00762f
C5823 vdd.n2855 gnd 0.00762f
C5824 vdd.n2857 gnd 0.950521f
C5825 vdd.n2859 gnd 0.00762f
C5826 vdd.n2860 gnd 0.00762f
C5827 vdd.n2861 gnd 0.018081f
C5828 vdd.n2862 gnd 0.016882f
C5829 vdd.n2863 gnd 0.016882f
C5830 vdd.n2864 gnd 0.950521f
C5831 vdd.n2865 gnd 0.016882f
C5832 vdd.n2866 gnd 0.016882f
C5833 vdd.n2867 gnd 0.00762f
C5834 vdd.n2868 gnd 0.00762f
C5835 vdd.n2869 gnd 0.00762f
C5836 vdd.n2870 gnd 0.486713f
C5837 vdd.n2871 gnd 0.00762f
C5838 vdd.n2872 gnd 0.00762f
C5839 vdd.n2873 gnd 0.00762f
C5840 vdd.n2874 gnd 0.00762f
C5841 vdd.n2875 gnd 0.00762f
C5842 vdd.n2876 gnd 0.606959f
C5843 vdd.n2877 gnd 0.00762f
C5844 vdd.n2878 gnd 0.00762f
C5845 vdd.n2879 gnd 0.00762f
C5846 vdd.n2880 gnd 0.00762f
C5847 vdd.n2881 gnd 0.00762f
C5848 vdd.n2882 gnd 0.77874f
C5849 vdd.n2883 gnd 0.00762f
C5850 vdd.n2884 gnd 0.00762f
C5851 vdd.n2885 gnd 0.00762f
C5852 vdd.n2886 gnd 0.00762f
C5853 vdd.n2887 gnd 0.00762f
C5854 vdd.n2888 gnd 0.429452f
C5855 vdd.n2889 gnd 0.00762f
C5856 vdd.n2890 gnd 0.00762f
C5857 vdd.n2891 gnd 0.00762f
C5858 vdd.n2892 gnd 0.00762f
C5859 vdd.n2893 gnd 0.00762f
C5860 vdd.n2894 gnd 0.246219f
C5861 vdd.n2895 gnd 0.00762f
C5862 vdd.n2896 gnd 0.00762f
C5863 vdd.n2897 gnd 0.00762f
C5864 vdd.n2898 gnd 0.00762f
C5865 vdd.n2899 gnd 0.00762f
C5866 vdd.n2900 gnd 0.446631f
C5867 vdd.n2901 gnd 0.00762f
C5868 vdd.n2902 gnd 0.00762f
C5869 vdd.n2903 gnd 0.00762f
C5870 vdd.n2904 gnd 0.00762f
C5871 vdd.n2905 gnd 0.00762f
C5872 vdd.n2906 gnd 0.618412f
C5873 vdd.n2907 gnd 0.00762f
C5874 vdd.n2908 gnd 0.00762f
C5875 vdd.n2909 gnd 0.00762f
C5876 vdd.n2910 gnd 0.00762f
C5877 vdd.n2911 gnd 0.00762f
C5878 vdd.n2912 gnd 0.69285f
C5879 vdd.n2913 gnd 0.00762f
C5880 vdd.n2914 gnd 0.00762f
C5881 vdd.n2915 gnd 0.00762f
C5882 vdd.n2916 gnd 0.00762f
C5883 vdd.n2917 gnd 0.00762f
C5884 vdd.n2918 gnd 0.521069f
C5885 vdd.n2919 gnd 0.00762f
C5886 vdd.n2920 gnd 0.00762f
C5887 vdd.n2921 gnd 0.00762f
C5888 vdd.t157 gnd 0.315203f
C5889 vdd.t155 gnd 0.201027f
C5890 vdd.t158 gnd 0.315203f
C5891 vdd.n2922 gnd 0.177157f
C5892 vdd.n2923 gnd 0.022075f
C5893 vdd.n2924 gnd 0.004707f
C5894 vdd.n2925 gnd 0.00762f
C5895 vdd.n2926 gnd 0.429452f
C5896 vdd.n2927 gnd 0.00762f
C5897 vdd.n2928 gnd 0.00762f
C5898 vdd.n2929 gnd 0.00762f
C5899 vdd.n2930 gnd 0.00762f
C5900 vdd.n2931 gnd 0.00762f
C5901 vdd.n2932 gnd 0.77874f
C5902 vdd.n2933 gnd 0.00762f
C5903 vdd.n2934 gnd 0.00762f
C5904 vdd.n2935 gnd 0.00762f
C5905 vdd.n2936 gnd 0.00762f
C5906 vdd.n2937 gnd 0.00762f
C5907 vdd.n2938 gnd 0.00762f
C5908 vdd.n2940 gnd 0.00762f
C5909 vdd.n2941 gnd 0.00762f
C5910 vdd.n2943 gnd 0.00762f
C5911 vdd.n2944 gnd 0.00762f
C5912 vdd.n2947 gnd 0.00762f
C5913 vdd.n2948 gnd 0.00762f
C5914 vdd.n2949 gnd 0.00762f
C5915 vdd.n2950 gnd 0.00762f
C5916 vdd.n2952 gnd 0.00762f
C5917 vdd.n2953 gnd 0.00762f
C5918 vdd.n2954 gnd 0.00762f
C5919 vdd.n2955 gnd 0.00762f
C5920 vdd.n2956 gnd 0.00762f
C5921 vdd.n2957 gnd 0.00762f
C5922 vdd.n2959 gnd 0.00762f
C5923 vdd.n2960 gnd 0.00762f
C5924 vdd.n2961 gnd 0.00762f
C5925 vdd.n2962 gnd 0.00762f
C5926 vdd.n2963 gnd 0.00762f
C5927 vdd.n2964 gnd 0.00762f
C5928 vdd.n2966 gnd 0.00762f
C5929 vdd.n2967 gnd 0.00762f
C5930 vdd.n2968 gnd 0.00762f
C5931 vdd.n2969 gnd 0.00762f
C5932 vdd.n2970 gnd 0.00762f
C5933 vdd.n2971 gnd 0.00762f
C5934 vdd.n2973 gnd 0.00762f
C5935 vdd.n2974 gnd 0.018081f
C5936 vdd.n2975 gnd 0.018081f
C5937 vdd.n2976 gnd 0.016882f
C5938 vdd.n2977 gnd 0.00762f
C5939 vdd.n2978 gnd 0.00762f
C5940 vdd.n2979 gnd 0.00762f
C5941 vdd.n2980 gnd 0.00762f
C5942 vdd.n2981 gnd 0.00762f
C5943 vdd.n2982 gnd 0.00762f
C5944 vdd.n2983 gnd 0.77874f
C5945 vdd.n2984 gnd 0.00762f
C5946 vdd.n2985 gnd 0.00762f
C5947 vdd.n2986 gnd 0.00762f
C5948 vdd.n2987 gnd 0.00762f
C5949 vdd.n2988 gnd 0.00762f
C5950 vdd.n2989 gnd 0.486713f
C5951 vdd.n2990 gnd 0.00762f
C5952 vdd.n2991 gnd 0.00762f
C5953 vdd.n2992 gnd 0.00762f
C5954 vdd.n2993 gnd 0.01781f
C5955 vdd.n2994 gnd 0.017153f
C5956 vdd.n2995 gnd 0.018081f
C5957 vdd.n2997 gnd 0.00762f
C5958 vdd.n2998 gnd 0.00762f
C5959 vdd.n2999 gnd 0.005883f
C5960 vdd.n3000 gnd 0.01089f
C5961 vdd.n3001 gnd 0.005547f
C5962 vdd.n3002 gnd 0.00762f
C5963 vdd.n3003 gnd 0.00762f
C5964 vdd.n3005 gnd 0.00762f
C5965 vdd.n3006 gnd 0.00762f
C5966 vdd.n3007 gnd 0.00762f
C5967 vdd.n3008 gnd 0.00762f
C5968 vdd.n3009 gnd 0.00762f
C5969 vdd.n3010 gnd 0.00762f
C5970 vdd.n3012 gnd 0.00762f
C5971 vdd.n3013 gnd 0.00762f
C5972 vdd.n3014 gnd 0.00762f
C5973 vdd.n3015 gnd 0.00762f
C5974 vdd.n3016 gnd 0.00762f
C5975 vdd.n3017 gnd 0.00762f
C5976 vdd.n3019 gnd 0.00762f
C5977 vdd.n3020 gnd 0.00762f
C5978 vdd.n3021 gnd 0.00762f
C5979 vdd.n3022 gnd 0.00762f
C5980 vdd.n3023 gnd 0.00762f
C5981 vdd.n3024 gnd 0.00762f
C5982 vdd.n3026 gnd 0.00762f
C5983 vdd.n3027 gnd 0.00762f
C5984 vdd.n3028 gnd 0.00762f
C5985 vdd.n3030 gnd 0.00762f
C5986 vdd.n3031 gnd 0.00762f
C5987 vdd.n3032 gnd 0.00762f
C5988 vdd.n3033 gnd 0.00762f
C5989 vdd.n3034 gnd 0.00762f
C5990 vdd.n3035 gnd 0.00762f
C5991 vdd.n3037 gnd 0.00762f
C5992 vdd.n3038 gnd 0.00762f
C5993 vdd.n3039 gnd 0.00762f
C5994 vdd.n3040 gnd 0.00762f
C5995 vdd.n3041 gnd 0.00762f
C5996 vdd.n3042 gnd 0.00762f
C5997 vdd.n3044 gnd 0.00762f
C5998 vdd.n3045 gnd 0.00762f
C5999 vdd.n3046 gnd 0.00762f
C6000 vdd.n3047 gnd 0.00762f
C6001 vdd.n3048 gnd 0.00762f
C6002 vdd.n3049 gnd 0.00762f
C6003 vdd.n3051 gnd 0.00762f
C6004 vdd.n3052 gnd 0.00762f
C6005 vdd.n3054 gnd 0.00762f
C6006 vdd.n3055 gnd 0.00762f
C6007 vdd.n3056 gnd 0.018081f
C6008 vdd.n3057 gnd 0.016882f
C6009 vdd.n3058 gnd 0.016882f
C6010 vdd.n3059 gnd 1.1223f
C6011 vdd.n3060 gnd 0.016882f
C6012 vdd.n3061 gnd 0.018081f
C6013 vdd.n3062 gnd 0.017153f
C6014 vdd.n3063 gnd 0.00762f
C6015 vdd.n3064 gnd 0.005883f
C6016 vdd.n3065 gnd 0.00762f
C6017 vdd.n3067 gnd 0.00762f
C6018 vdd.n3068 gnd 0.00762f
C6019 vdd.n3069 gnd 0.00762f
C6020 vdd.n3070 gnd 0.00762f
C6021 vdd.n3071 gnd 0.00762f
C6022 vdd.n3072 gnd 0.00762f
C6023 vdd.n3074 gnd 0.00762f
C6024 vdd.n3075 gnd 0.00762f
C6025 vdd.n3076 gnd 0.00762f
C6026 vdd.n3077 gnd 0.00762f
C6027 vdd.n3078 gnd 0.00762f
C6028 vdd.n3079 gnd 0.00762f
C6029 vdd.n3081 gnd 0.00762f
C6030 vdd.n3082 gnd 0.00762f
C6031 vdd.n3083 gnd 0.00762f
C6032 vdd.n3084 gnd 0.00762f
C6033 vdd.n3085 gnd 0.00762f
C6034 vdd.n3086 gnd 0.00762f
C6035 vdd.n3088 gnd 0.00762f
C6036 vdd.n3089 gnd 0.00762f
C6037 vdd.n3091 gnd 0.00762f
C6038 vdd.n3092 gnd 0.018311f
C6039 vdd.n3093 gnd 0.678209f
C6040 vdd.n3095 gnd 0.004735f
C6041 vdd.n3096 gnd 0.00902f
C6042 vdd.n3097 gnd 0.011206f
C6043 vdd.n3098 gnd 0.011206f
C6044 vdd.n3099 gnd 0.00902f
C6045 vdd.n3100 gnd 0.00902f
C6046 vdd.n3101 gnd 0.011206f
C6047 vdd.n3102 gnd 0.011206f
C6048 vdd.n3103 gnd 0.00902f
C6049 vdd.n3104 gnd 0.00902f
C6050 vdd.n3105 gnd 0.011206f
C6051 vdd.n3106 gnd 0.011206f
C6052 vdd.n3107 gnd 0.00902f
C6053 vdd.n3108 gnd 0.00902f
C6054 vdd.n3109 gnd 0.011206f
C6055 vdd.n3110 gnd 0.011206f
C6056 vdd.n3111 gnd 0.00902f
C6057 vdd.n3112 gnd 0.00902f
C6058 vdd.n3113 gnd 0.011206f
C6059 vdd.n3114 gnd 0.011206f
C6060 vdd.n3115 gnd 0.00902f
C6061 vdd.n3116 gnd 0.00902f
C6062 vdd.n3117 gnd 0.011206f
C6063 vdd.n3118 gnd 0.011206f
C6064 vdd.n3119 gnd 0.00902f
C6065 vdd.n3120 gnd 0.00902f
C6066 vdd.n3121 gnd 0.011206f
C6067 vdd.n3122 gnd 0.011206f
C6068 vdd.n3123 gnd 0.00902f
C6069 vdd.n3124 gnd 0.00902f
C6070 vdd.n3125 gnd 0.011206f
C6071 vdd.n3126 gnd 0.011206f
C6072 vdd.n3127 gnd 0.00902f
C6073 vdd.n3128 gnd 0.00902f
C6074 vdd.n3129 gnd 0.011206f
C6075 vdd.n3130 gnd 0.011206f
C6076 vdd.n3131 gnd 0.00902f
C6077 vdd.n3132 gnd 0.011206f
C6078 vdd.n3133 gnd 0.011206f
C6079 vdd.n3134 gnd 0.00902f
C6080 vdd.n3135 gnd 0.011206f
C6081 vdd.n3136 gnd 0.011206f
C6082 vdd.n3137 gnd 0.011206f
C6083 vdd.n3138 gnd 0.0184f
C6084 vdd.n3139 gnd 0.011206f
C6085 vdd.n3140 gnd 0.011206f
C6086 vdd.n3141 gnd 0.006133f
C6087 vdd.n3142 gnd 0.00902f
C6088 vdd.n3143 gnd 0.011206f
C6089 vdd.n3144 gnd 0.011206f
C6090 vdd.n3145 gnd 0.00902f
C6091 vdd.n3146 gnd 0.00902f
C6092 vdd.n3147 gnd 0.011206f
C6093 vdd.n3148 gnd 0.011206f
C6094 vdd.n3149 gnd 0.00902f
C6095 vdd.n3150 gnd 0.00902f
C6096 vdd.n3151 gnd 0.011206f
C6097 vdd.n3152 gnd 0.011206f
C6098 vdd.n3153 gnd 0.00902f
C6099 vdd.n3154 gnd 0.00902f
C6100 vdd.n3155 gnd 0.011206f
C6101 vdd.n3156 gnd 0.011206f
C6102 vdd.n3157 gnd 0.00902f
C6103 vdd.n3158 gnd 0.00902f
C6104 vdd.n3159 gnd 0.011206f
C6105 vdd.n3160 gnd 0.011206f
C6106 vdd.n3161 gnd 0.00902f
C6107 vdd.n3162 gnd 0.00902f
C6108 vdd.n3163 gnd 0.011206f
C6109 vdd.n3164 gnd 0.011206f
C6110 vdd.n3165 gnd 0.00902f
C6111 vdd.n3166 gnd 0.00902f
C6112 vdd.n3167 gnd 0.011206f
C6113 vdd.n3168 gnd 0.011206f
C6114 vdd.n3169 gnd 0.00902f
C6115 vdd.n3170 gnd 0.00902f
C6116 vdd.n3171 gnd 0.011206f
C6117 vdd.n3172 gnd 0.011206f
C6118 vdd.n3173 gnd 0.00902f
C6119 vdd.n3174 gnd 0.00902f
C6120 vdd.n3175 gnd 0.011206f
C6121 vdd.n3176 gnd 0.011206f
C6122 vdd.n3177 gnd 0.00902f
C6123 vdd.n3178 gnd 0.011206f
C6124 vdd.n3179 gnd 0.011206f
C6125 vdd.n3180 gnd 0.00902f
C6126 vdd.n3181 gnd 0.011206f
C6127 vdd.n3182 gnd 0.011206f
C6128 vdd.n3183 gnd 0.011206f
C6129 vdd.t149 gnd 0.137864f
C6130 vdd.t150 gnd 0.147339f
C6131 vdd.t148 gnd 0.180049f
C6132 vdd.n3184 gnd 0.230797f
C6133 vdd.n3185 gnd 0.193911f
C6134 vdd.n3186 gnd 0.0184f
C6135 vdd.n3187 gnd 0.011206f
C6136 vdd.n3188 gnd 0.011206f
C6137 vdd.n3189 gnd 0.007531f
C6138 vdd.n3190 gnd 0.00902f
C6139 vdd.n3191 gnd 0.011206f
C6140 vdd.n3192 gnd 0.011206f
C6141 vdd.n3193 gnd 0.00902f
C6142 vdd.n3194 gnd 0.00902f
C6143 vdd.n3195 gnd 0.011206f
C6144 vdd.n3196 gnd 0.011206f
C6145 vdd.n3197 gnd 0.00902f
C6146 vdd.n3198 gnd 0.00902f
C6147 vdd.n3199 gnd 0.011206f
C6148 vdd.n3200 gnd 0.011206f
C6149 vdd.n3201 gnd 0.00902f
C6150 vdd.n3202 gnd 0.00902f
C6151 vdd.n3203 gnd 0.011206f
C6152 vdd.n3204 gnd 0.011206f
C6153 vdd.n3205 gnd 0.00902f
C6154 vdd.n3206 gnd 0.00902f
C6155 vdd.n3207 gnd 0.011206f
C6156 vdd.n3208 gnd 0.011206f
C6157 vdd.n3209 gnd 0.00902f
C6158 vdd.n3210 gnd 0.00902f
C6159 vdd.n3211 gnd 0.011206f
C6160 vdd.n3212 gnd 0.011206f
C6161 vdd.n3213 gnd 0.00902f
C6162 vdd.n3214 gnd 0.00902f
C6163 vdd.n3216 gnd 0.678209f
C6164 vdd.n3218 gnd 0.00902f
C6165 vdd.n3219 gnd 0.00902f
C6166 vdd.n3220 gnd 0.007486f
C6167 vdd.n3221 gnd 0.027689f
C6168 vdd.n3223 gnd 8.27984f
C6169 vdd.n3224 gnd 0.027689f
C6170 vdd.n3225 gnd 0.004284f
C6171 vdd.n3226 gnd 0.027689f
C6172 vdd.n3227 gnd 0.027108f
C6173 vdd.n3228 gnd 0.011206f
C6174 vdd.n3229 gnd 0.00902f
C6175 vdd.n3230 gnd 0.011206f
C6176 vdd.n3231 gnd 0.69285f
C6177 vdd.n3232 gnd 0.011206f
C6178 vdd.n3233 gnd 0.00902f
C6179 vdd.n3234 gnd 0.011206f
C6180 vdd.n3235 gnd 0.011206f
C6181 vdd.n3236 gnd 0.011206f
C6182 vdd.n3237 gnd 0.00902f
C6183 vdd.n3238 gnd 0.011206f
C6184 vdd.n3239 gnd 1.14521f
C6185 vdd.n3240 gnd 0.011206f
C6186 vdd.n3241 gnd 0.00902f
C6187 vdd.n3242 gnd 0.011206f
C6188 vdd.n3243 gnd 0.011206f
C6189 vdd.n3244 gnd 0.011206f
C6190 vdd.n3245 gnd 0.00902f
C6191 vdd.n3246 gnd 0.011206f
C6192 vdd.n3247 gnd 0.738658f
C6193 vdd.n3248 gnd 0.784466f
C6194 vdd.n3249 gnd 0.011206f
C6195 vdd.n3250 gnd 0.00902f
C6196 vdd.n3251 gnd 0.011206f
C6197 vdd.n3252 gnd 0.011206f
C6198 vdd.n3253 gnd 0.011206f
C6199 vdd.n3254 gnd 0.00902f
C6200 vdd.n3255 gnd 0.011206f
C6201 vdd.n3256 gnd 0.950521f
C6202 vdd.n3257 gnd 0.011206f
C6203 vdd.n3258 gnd 0.00902f
C6204 vdd.n3259 gnd 0.011206f
C6205 vdd.n3260 gnd 0.011206f
C6206 vdd.n3261 gnd 0.011206f
C6207 vdd.n3262 gnd 0.00902f
C6208 vdd.n3263 gnd 0.011206f
C6209 vdd.t80 gnd 0.572603f
C6210 vdd.n3264 gnd 0.921891f
C6211 vdd.n3265 gnd 0.011206f
C6212 vdd.n3266 gnd 0.00902f
C6213 vdd.n3267 gnd 0.011206f
C6214 vdd.n3268 gnd 0.011206f
C6215 vdd.n3269 gnd 0.011206f
C6216 vdd.n3270 gnd 0.00902f
C6217 vdd.n3271 gnd 0.011206f
C6218 vdd.n3272 gnd 0.727206f
C6219 vdd.n3273 gnd 0.011206f
C6220 vdd.n3274 gnd 0.00902f
C6221 vdd.n3275 gnd 0.011206f
C6222 vdd.n3276 gnd 0.011206f
C6223 vdd.n3277 gnd 0.011206f
C6224 vdd.n3278 gnd 0.00902f
C6225 vdd.n3279 gnd 0.011206f
C6226 vdd.n3280 gnd 0.910439f
C6227 vdd.n3281 gnd 0.612685f
C6228 vdd.n3282 gnd 0.011206f
C6229 vdd.n3283 gnd 0.00902f
C6230 vdd.n3284 gnd 0.011206f
C6231 vdd.n3285 gnd 0.011206f
C6232 vdd.n3286 gnd 0.011206f
C6233 vdd.n3287 gnd 0.00902f
C6234 vdd.n3288 gnd 0.011206f
C6235 vdd.n3289 gnd 0.807371f
C6236 vdd.n3290 gnd 0.011206f
C6237 vdd.n3291 gnd 0.00902f
C6238 vdd.n3292 gnd 0.011206f
C6239 vdd.n3293 gnd 0.011206f
C6240 vdd.n3294 gnd 0.011206f
C6241 vdd.n3295 gnd 0.011206f
C6242 vdd.n3296 gnd 0.011206f
C6243 vdd.n3297 gnd 0.00902f
C6244 vdd.n3298 gnd 0.00902f
C6245 vdd.n3299 gnd 0.011206f
C6246 vdd.t16 gnd 0.572603f
C6247 vdd.n3300 gnd 0.950521f
C6248 vdd.n3301 gnd 0.011206f
C6249 vdd.n3302 gnd 0.00902f
C6250 vdd.n3303 gnd 0.011206f
C6251 vdd.n3304 gnd 0.011206f
C6252 vdd.n3305 gnd 0.011206f
C6253 vdd.n3306 gnd 0.00902f
C6254 vdd.n3307 gnd 0.011206f
C6255 vdd.n3308 gnd 0.898987f
C6256 vdd.n3309 gnd 0.011206f
C6257 vdd.n3310 gnd 0.011206f
C6258 vdd.n3311 gnd 0.00902f
C6259 vdd.n3312 gnd 0.00902f
C6260 vdd.n3313 gnd 0.011206f
C6261 vdd.n3314 gnd 0.011206f
C6262 vdd.n3315 gnd 0.011206f
C6263 vdd.n3316 gnd 0.00902f
C6264 vdd.n3317 gnd 0.011206f
C6265 vdd.n3318 gnd 0.00902f
C6266 vdd.n3319 gnd 0.00902f
C6267 vdd.n3320 gnd 0.011206f
C6268 vdd.n3321 gnd 0.011206f
C6269 vdd.n3322 gnd 0.011206f
C6270 vdd.n3323 gnd 0.00902f
C6271 vdd.n3324 gnd 0.011206f
C6272 vdd.n3325 gnd 0.00902f
C6273 vdd.n3326 gnd 0.00902f
C6274 vdd.n3327 gnd 0.011206f
C6275 vdd.n3328 gnd 0.011206f
C6276 vdd.n3329 gnd 0.011206f
C6277 vdd.n3330 gnd 0.00902f
C6278 vdd.n3331 gnd 0.950521f
C6279 vdd.n3332 gnd 0.011206f
C6280 vdd.n3333 gnd 0.00902f
C6281 vdd.n3334 gnd 0.00902f
C6282 vdd.n3335 gnd 0.011206f
C6283 vdd.n3336 gnd 0.011206f
C6284 vdd.n3337 gnd 0.011206f
C6285 vdd.n3338 gnd 0.00902f
C6286 vdd.n3339 gnd 0.011206f
C6287 vdd.n3340 gnd 0.00902f
C6288 vdd.n3341 gnd 0.00902f
C6289 vdd.n3342 gnd 0.011206f
C6290 vdd.n3343 gnd 0.011206f
C6291 vdd.n3344 gnd 0.011206f
C6292 vdd.n3345 gnd 0.00902f
C6293 vdd.n3346 gnd 0.011206f
C6294 vdd.n3347 gnd 0.00902f
C6295 vdd.n3348 gnd 0.007486f
C6296 vdd.n3349 gnd 0.027108f
C6297 vdd.n3350 gnd 0.027689f
C6298 vdd.n3351 gnd 0.004284f
C6299 vdd.n3352 gnd 0.027689f
C6300 vdd.n3354 gnd 2.71414f
C6301 vdd.n3355 gnd 1.68918f
C6302 vdd.n3356 gnd 0.027108f
C6303 vdd.n3357 gnd 0.007486f
C6304 vdd.n3358 gnd 0.00902f
C6305 vdd.n3359 gnd 0.00902f
C6306 vdd.n3360 gnd 0.011206f
C6307 vdd.n3361 gnd 1.14521f
C6308 vdd.n3362 gnd 1.14521f
C6309 vdd.n3363 gnd 1.04786f
C6310 vdd.n3364 gnd 0.011206f
C6311 vdd.n3365 gnd 0.00902f
C6312 vdd.n3366 gnd 0.00902f
C6313 vdd.n3367 gnd 0.00902f
C6314 vdd.n3368 gnd 0.011206f
C6315 vdd.n3369 gnd 0.853179f
C6316 vdd.t74 gnd 0.572603f
C6317 vdd.n3370 gnd 0.864631f
C6318 vdd.n3371 gnd 0.658494f
C6319 vdd.n3372 gnd 0.011206f
C6320 vdd.n3373 gnd 0.00902f
C6321 vdd.n3374 gnd 0.00902f
C6322 vdd.n3375 gnd 0.00902f
C6323 vdd.n3376 gnd 0.011206f
C6324 vdd.n3377 gnd 0.681398f
C6325 vdd.n3378 gnd 0.841727f
C6326 vdd.t95 gnd 0.572603f
C6327 vdd.n3379 gnd 0.876083f
C6328 vdd.n3380 gnd 0.011206f
C6329 vdd.n3381 gnd 0.00902f
C6330 vdd.n3382 gnd 0.00902f
C6331 vdd.n3383 gnd 0.00902f
C6332 vdd.n3384 gnd 0.011206f
C6333 vdd.n3385 gnd 0.950521f
C6334 vdd.t24 gnd 0.572603f
C6335 vdd.n3386 gnd 0.69285f
C6336 vdd.n3387 gnd 0.830275f
C6337 vdd.n3388 gnd 0.011206f
C6338 vdd.n3389 gnd 0.00902f
C6339 vdd.n3390 gnd 0.00902f
C6340 vdd.n3391 gnd 0.00902f
C6341 vdd.n3392 gnd 0.011206f
C6342 vdd.n3393 gnd 0.63559f
C6343 vdd.t64 gnd 0.572603f
C6344 vdd.n3394 gnd 0.950521f
C6345 vdd.t7 gnd 0.572603f
C6346 vdd.n3395 gnd 0.704302f
C6347 vdd.n3396 gnd 0.011206f
C6348 vdd.n3397 gnd 0.00902f
C6349 vdd.n3398 gnd 0.008613f
C6350 vdd.n3399 gnd 0.660976f
C6351 vdd.n3400 gnd 2.86555f
C6352 a_n2848_n452.n0 gnd 3.415f
C6353 a_n2848_n452.n1 gnd 0.285666f
C6354 a_n2848_n452.n2 gnd 0.492471f
C6355 a_n2848_n452.n3 gnd 0.664435f
C6356 a_n2848_n452.n4 gnd 0.215942f
C6357 a_n2848_n452.n5 gnd 0.282512f
C6358 a_n2848_n452.n6 gnd 0.546457f
C6359 a_n2848_n452.n7 gnd 0.526038f
C6360 a_n2848_n452.n8 gnd 0.204894f
C6361 a_n2848_n452.n9 gnd 0.150908f
C6362 a_n2848_n452.n10 gnd 0.23718f
C6363 a_n2848_n452.n11 gnd 0.183194f
C6364 a_n2848_n452.n12 gnd 0.204894f
C6365 a_n2848_n452.n13 gnd 1.0063f
C6366 a_n2848_n452.n14 gnd 0.150908f
C6367 a_n2848_n452.n15 gnd 0.580023f
C6368 a_n2848_n452.n16 gnd 0.432289f
C6369 a_n2848_n452.n17 gnd 0.215942f
C6370 a_n2848_n452.n18 gnd 0.492471f
C6371 a_n2848_n452.n19 gnd 0.282512f
C6372 a_n2848_n452.n20 gnd 0.438486f
C6373 a_n2848_n452.n21 gnd 0.215942f
C6374 a_n2848_n452.n22 gnd 0.731535f
C6375 a_n2848_n452.n23 gnd 0.282512f
C6376 a_n2848_n452.n24 gnd 1.17886f
C6377 a_n2848_n452.n25 gnd 1.91568f
C6378 a_n2848_n452.n26 gnd 1.14458f
C6379 a_n2848_n452.n27 gnd 1.77783f
C6380 a_n2848_n452.n28 gnd 0.377489f
C6381 a_n2848_n452.n29 gnd 3.11576f
C6382 a_n2848_n452.n30 gnd 0.377488f
C6383 a_n2848_n452.n31 gnd 3.20158f
C6384 a_n2848_n452.n32 gnd 0.008361f
C6385 a_n2848_n452.n34 gnd 0.285666f
C6386 a_n2848_n452.n35 gnd 0.008361f
C6387 a_n2848_n452.n37 gnd 0.285666f
C6388 a_n2848_n452.n38 gnd 0.008361f
C6389 a_n2848_n452.n39 gnd 0.28526f
C6390 a_n2848_n452.n40 gnd 0.008361f
C6391 a_n2848_n452.n41 gnd 0.28526f
C6392 a_n2848_n452.n42 gnd 0.008361f
C6393 a_n2848_n452.n43 gnd 0.28526f
C6394 a_n2848_n452.n44 gnd 0.008361f
C6395 a_n2848_n452.n45 gnd 0.28526f
C6396 a_n2848_n452.n47 gnd 0.285666f
C6397 a_n2848_n452.n48 gnd 0.008361f
C6398 a_n2848_n452.n50 gnd 0.285666f
C6399 a_n2848_n452.t28 gnd 0.14978f
C6400 a_n2848_n452.t39 gnd 0.708223f
C6401 a_n2848_n452.t27 gnd 0.696704f
C6402 a_n2848_n452.t21 gnd 0.696704f
C6403 a_n2848_n452.t17 gnd 0.116496f
C6404 a_n2848_n452.t3 gnd 0.116496f
C6405 a_n2848_n452.n52 gnd 1.03243f
C6406 a_n2848_n452.t5 gnd 0.116496f
C6407 a_n2848_n452.t6 gnd 0.116496f
C6408 a_n2848_n452.n53 gnd 1.0294f
C6409 a_n2848_n452.n54 gnd 0.912817f
C6410 a_n2848_n452.t4 gnd 0.116496f
C6411 a_n2848_n452.t10 gnd 0.116496f
C6412 a_n2848_n452.n55 gnd 1.0294f
C6413 a_n2848_n452.t19 gnd 0.116496f
C6414 a_n2848_n452.t18 gnd 0.116496f
C6415 a_n2848_n452.n56 gnd 1.03243f
C6416 a_n2848_n452.t2 gnd 0.116496f
C6417 a_n2848_n452.t12 gnd 0.116496f
C6418 a_n2848_n452.n57 gnd 1.0294f
C6419 a_n2848_n452.n58 gnd 0.912817f
C6420 a_n2848_n452.t0 gnd 0.116496f
C6421 a_n2848_n452.t15 gnd 0.116496f
C6422 a_n2848_n452.n59 gnd 1.0294f
C6423 a_n2848_n452.t7 gnd 0.116496f
C6424 a_n2848_n452.t8 gnd 0.116496f
C6425 a_n2848_n452.n60 gnd 1.0294f
C6426 a_n2848_n452.n61 gnd 3.15028f
C6427 a_n2848_n452.t20 gnd 0.116496f
C6428 a_n2848_n452.t14 gnd 0.116496f
C6429 a_n2848_n452.n62 gnd 1.0294f
C6430 a_n2848_n452.n63 gnd 0.449443f
C6431 a_n2848_n452.t11 gnd 0.116496f
C6432 a_n2848_n452.t47 gnd 0.116496f
C6433 a_n2848_n452.n64 gnd 1.0294f
C6434 a_n2848_n452.t9 gnd 0.116496f
C6435 a_n2848_n452.t1 gnd 0.116496f
C6436 a_n2848_n452.n65 gnd 1.03243f
C6437 a_n2848_n452.t16 gnd 0.116496f
C6438 a_n2848_n452.t13 gnd 0.116496f
C6439 a_n2848_n452.n66 gnd 1.0294f
C6440 a_n2848_n452.n67 gnd 0.912814f
C6441 a_n2848_n452.t46 gnd 0.116496f
C6442 a_n2848_n452.t45 gnd 0.116496f
C6443 a_n2848_n452.n68 gnd 1.0294f
C6444 a_n2848_n452.t41 gnd 0.696704f
C6445 a_n2848_n452.n69 gnd 0.302425f
C6446 a_n2848_n452.t35 gnd 0.696704f
C6447 a_n2848_n452.t37 gnd 0.708223f
C6448 a_n2848_n452.t75 gnd 0.711378f
C6449 a_n2848_n452.t58 gnd 0.696704f
C6450 a_n2848_n452.t62 gnd 0.696704f
C6451 a_n2848_n452.t52 gnd 0.696704f
C6452 a_n2848_n452.n70 gnd 0.306315f
C6453 a_n2848_n452.t67 gnd 0.696704f
C6454 a_n2848_n452.t73 gnd 0.708223f
C6455 a_n2848_n452.t24 gnd 1.40246f
C6456 a_n2848_n452.t26 gnd 0.14978f
C6457 a_n2848_n452.t34 gnd 0.14978f
C6458 a_n2848_n452.n71 gnd 1.05505f
C6459 a_n2848_n452.t30 gnd 0.14978f
C6460 a_n2848_n452.t32 gnd 0.14978f
C6461 a_n2848_n452.n72 gnd 1.05505f
C6462 a_n2848_n452.t44 gnd 1.39967f
C6463 a_n2848_n452.t29 gnd 0.696704f
C6464 a_n2848_n452.n73 gnd 0.306315f
C6465 a_n2848_n452.t31 gnd 0.696704f
C6466 a_n2848_n452.t25 gnd 0.696704f
C6467 a_n2848_n452.t56 gnd 0.696704f
C6468 a_n2848_n452.n74 gnd 0.306315f
C6469 a_n2848_n452.t65 gnd 0.696704f
C6470 a_n2848_n452.t71 gnd 0.696704f
C6471 a_n2848_n452.t70 gnd 0.711378f
C6472 a_n2848_n452.n75 gnd 0.308932f
C6473 a_n2848_n452.t50 gnd 0.696704f
C6474 a_n2848_n452.n76 gnd 0.302425f
C6475 a_n2848_n452.n77 gnd 0.308933f
C6476 a_n2848_n452.t51 gnd 0.708223f
C6477 a_n2848_n452.t23 gnd 0.711378f
C6478 a_n2848_n452.n78 gnd 0.308932f
C6479 a_n2848_n452.t33 gnd 0.696704f
C6480 a_n2848_n452.n79 gnd 0.302425f
C6481 a_n2848_n452.n80 gnd 0.308933f
C6482 a_n2848_n452.t43 gnd 0.708223f
C6483 a_n2848_n452.n81 gnd 1.13204f
C6484 a_n2848_n452.t55 gnd 0.696704f
C6485 a_n2848_n452.n82 gnd 0.302425f
C6486 a_n2848_n452.t61 gnd 0.696704f
C6487 a_n2848_n452.n83 gnd 0.302425f
C6488 a_n2848_n452.t53 gnd 0.696704f
C6489 a_n2848_n452.n84 gnd 0.302425f
C6490 a_n2848_n452.t66 gnd 0.696704f
C6491 a_n2848_n452.n85 gnd 0.302425f
C6492 a_n2848_n452.t57 gnd 0.696704f
C6493 a_n2848_n452.n86 gnd 0.296933f
C6494 a_n2848_n452.t48 gnd 0.696704f
C6495 a_n2848_n452.n87 gnd 0.306315f
C6496 a_n2848_n452.t59 gnd 0.708378f
C6497 a_n2848_n452.t68 gnd 0.696704f
C6498 a_n2848_n452.n88 gnd 0.296933f
C6499 a_n2848_n452.t54 gnd 0.696704f
C6500 a_n2848_n452.n89 gnd 0.306315f
C6501 a_n2848_n452.t63 gnd 0.708378f
C6502 a_n2848_n452.t72 gnd 0.696704f
C6503 a_n2848_n452.n90 gnd 0.296933f
C6504 a_n2848_n452.t60 gnd 0.696704f
C6505 a_n2848_n452.n91 gnd 0.306315f
C6506 a_n2848_n452.t74 gnd 0.708378f
C6507 a_n2848_n452.t64 gnd 0.696704f
C6508 a_n2848_n452.n92 gnd 0.296933f
C6509 a_n2848_n452.t49 gnd 0.696704f
C6510 a_n2848_n452.n93 gnd 0.306315f
C6511 a_n2848_n452.t69 gnd 0.708378f
C6512 a_n2848_n452.n94 gnd 1.33845f
C6513 a_n2848_n452.n95 gnd 0.308933f
C6514 a_n2848_n452.n96 gnd 0.302425f
C6515 a_n2848_n452.n97 gnd 0.308932f
C6516 a_n2848_n452.n98 gnd 0.308933f
C6517 a_n2848_n452.n99 gnd 0.01225f
C6518 a_n2848_n452.n100 gnd 0.302425f
C6519 a_n2848_n452.n101 gnd 0.308933f
C6520 a_n2848_n452.n102 gnd 0.786935f
C6521 a_n2848_n452.t40 gnd 1.39967f
C6522 a_n2848_n452.t38 gnd 1.40246f
C6523 a_n2848_n452.t42 gnd 0.14978f
C6524 a_n2848_n452.t36 gnd 0.14978f
C6525 a_n2848_n452.n103 gnd 1.05505f
C6526 a_n2848_n452.n104 gnd 1.05505f
C6527 a_n2848_n452.t22 gnd 0.14978f
.ends

